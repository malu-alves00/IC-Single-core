`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PZHlLaxuFbwAc9iHdlkB4j00wTXVFJTi8zR0TwqkhocY8YRD6TGkLEqKJRILrgdz
f+qJFNi1w1L21fAm4/42CX/Jd/03d/Oi7FJto3osrVlLhCMxFX6bCI+q6A43pbZ2
wXyEmTydhP3snn4MaMBxZOOt5FRNdMcdUeMAVIhMlXgLHVUTr20QhNllmE4+CSHh
CxtksaAcTdXFQkmXJi2JSm81/ZMcCOICVh4GyaMC9wZxnO9pu9Z94q+nFX2dv2z6
+lL5pxeeNqli8yMkae3xOi7qoeBZbv/UtLzhThLdKhA8jhn7rYRnx+4CYKLKycbf
aLou7T9X2tzw0Ip1sMBNeG33E+Yz1l9gXTZXKG4URyS1Rkn1Dl/fxFuB2R7mdMKc
s3RmdhCjSeo7xlxwMsf6w0OGZQIKusauMDrDaFMV+xLnzEmJo8u+TPv+xVfSyee7
uU/pD5dTA4IvLn/ksbp+acZJMdRTM7pZLSfuXKAJF8yqCNvkurjUnlxLrFu3k+O0
XgG4RV6PfOvEtQDM52sKZOaQZ4c4KmfOy4PfUdD2DU5fJrila27GQTa/HRUi6pSb
eyS9G3YDGNPY8T3q0KJeSVb4IHN+4QPmT2dylPBIX6cScSrThBJybIGmSp+vcnAV
aZfSxJJuKskcJ2gr5Foy+vYS5thOo8lhIpDgbDBYC6TDmn7rsiE1xUU977ZmQRr8
ZEaOekHz/C8Pb8EVZx/EOxFRevzL3zfz35rJ4wj1uI3xN5iO8ZtVAA2YAnIlsHmr
0nVZxSNSzrFhitFFv9WQAsKW6gWO0hnIi+c2OquBfYODHjj0F0DVSthlxwf93ST/
updeDM4pf4EzERA3LArcTBm5JfZIjeGJHTJdGi8zqc/yEKTc3/3mBf8cZIQZPCfL
MNwz76jjGGLAXEfLqo3C/3pJDSlKd2xWm5H9Pc2GBkvJgfZk4z7eFGFwTWm3yHVA
ig6iTqf7pdb4Gg9U5pZL7tUNaLFEZXVOuPD3GXmiLgojfbaO8wJPZZzoPPH+Nr7S
dRIzr+6LczkwtIP9eQUmrIrv0lCbLD1pPPIeyrXTTMg=
`protect END_PROTECTED
