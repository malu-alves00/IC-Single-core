`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BsAFuieY15A8ZZ92KcVJ4bqKWm7IqviiQkX+KFZL0NdwQL0YkBhlaDplEhxGXAUu
ZEG6tRs8IzdTfQTjVrfz+/7YINysKL4Y8iEHcvjzHp5AH/M1wCRY/vgyHp3Dv8Sw
Ld8NmI3e3urrjxUSPuiy99ronKtHTVkIvUSHIrVRSH20SD7dAXPfE68/9dic6L5w
`protect END_PROTECTED
