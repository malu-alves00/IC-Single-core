`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OeBNhmMlz+fAg8/48oEYBPBiXwIsYiaEg1KlxXvX3kOqNKSKtMS2C2UpbXUcwwfG
iRDyYQS/Q4e8B/MW47BLoLc8JcOcESE8OXEMSSuwuRoz+kqAvnoUESL+F6JGsUyj
Pnuehx7bFYnHwihsTBnNEt83HjuQ1Hc7uNklYJ45DXgtoWg/YW0cyriaf+GNVbDp
1D45sEjQ9EcjIZ4XwQSMc0vTiY7AZR9/1wZIveKGwu4/tHtePTWhUzGbiPpjA8gq
KNltPBoqADQPZNeTdfBMNXnQ1khOtw+bpeJ2WG/W+87aGXpMViOULuUBfIxkWNVE
IzQAdFB3B8XfWoOrvh/+R/Cwv1yhbbnyV5RlShw/hef+F05Y/+FAH0z/Vuv6ySsn
qUcTvlRGIWNuAj68sXYRW2ILHTEYFq+aUb7QcsTJ1RpJOGEURQzIJCY2lbaUn1sj
2bZtGKOGM4uan0Vp5UMx6XDICKqmEED2kG94JlPdMCvYnvORNEpJYfuOl+SxZAAx
5cuV2URZ/Sc9HHs1Ip6mEasAZQ02Om6T/h5cp2DDbLnXr0r3Zaw7fFGM+rp5tS6B
Veocbynd2DW1Q9T4iQrstEKYCq7hgEgrOTlTYTvknXROlZJhbyFRc0OgM7fKI+8Z
J2XGX4U+hyP7XFj8Uqg/8PMsHtLhRncw2OhmxVDEju0VfhIMnbMb5B+YYVwAeYWI
jURwv02opf+Jma8ftyIye8gjAgNY8YuxWglOR+Tq6RFucrgQ3fSlYeLk7Lton+Nd
RwhmyWLtWr3GFx0iiXRiTWi5WhVGezjNaznzOXtiCf6rVBmAUrw9+N7W42U73CBN
466gTPWF7SsTOsHMMyKq8SJ1dfYDdslPi8yGPr7eowx+CKqRLGw/JXtUWcrY08ke
MqanY+IDaxc6/L968Cumaj5cr2j67O1XULfs4gGfLqi0cEw3UEFDLEPxhIpfx7M9
PC7+OVbETWgcCCpMssFy3Ebowc2s4eDe5ovrgIsVXKrxf6O84tIRlvf4TNWNICgq
RWH1HDM9IQdDC92jbxfZp16SckCuA4iFhvLsIVkjGvuPIfKLFEJ074bTB5GZUVDk
jXFfpEW7cG8RKkgbydvkBn0ArWIruXXZVmW5uLLX3TXxuX77S455TvfUBrXo3wPv
jRCsYNd9btyRiJ0HvkPWRpLG30vSW7ytNtGAPL1UVDlRREh9gnngiBgof1BvrOzc
YaatUDedMsKP2ESmEv3wQGZbP39+S56lZxr1MdUVw/t3T6vB+P1ND1r/YJC1xpvu
9CicqfGJ5PekK69fOtSw8IIolFwgQ7P45LDTth2onT/c3pavQKQsX60HjQk8I1mG
pvaauWN8kwnBbGN6F0cNVUGCpV6S5wfFB97qb9g+ovi2CfojTYbSxy8XbT6n56aq
IvztuShzOHv0fJTC3TQA9A6G/mrMlCcqIDG5mb41E/oD0svbO+UaaWbtCjhjQCEB
duCt863mJMUxlPAfe5jblL9RabB1I6Mx9EbAzy6hs+9COf2iO/8COg65oOKcXFkM
1E/W3MhpXbdK+vOjf/HI4LUNHcw25zr4by5HF8qQHYSyb+ZENyhLvDry39myai0y
wfr+zl16N3yA9w/6uhBNND0ZZgfMoDeY9+XYpXl36TaB6lFE8ve7ZIGb/UAVQOxA
B5OsckG+6biUYAdqhXsTUQU13W4mxYt9PD2foR7FEOPE4/lMyfPnptxhL0NailRf
gQ2BR36x4qeXchCvju4/RwcORkev0z15lc6HHIAXHRzqFMv6Z1J0WCOVo0taPNeV
uqJX8MK/pTl8lsVx5B1BLuMklID3Cu8tEqqAZTykS0QXrXxGqnG1yB/E9Ccdjkjp
OW9/blM/JM0Vm+dCgsGulnogH2Nfd5LPHgTEvaEUds8el0E0G4Eo4CXn8lRoTynH
UU2UGy8UoUlyygZ36m3cs5aIfuMsjQXRRrH8Wle1S89DwlPRTKzJ93mKWy1/sOur
Kt8Kgap0HcpmbkdI5dwBYXAGDHiYQO42uV2CTLN2CmEwJO9NYBtR7CuTsfcIXqtf
kled00EtmnUpX3QXiURO/bysngLLX2ZxMYGPTeqnjE6eYuohgdP1sjTCGTrzrMC7
iISjqB98QwjzPibmbXj7YQZZ/sEk3eikcsBriWQvU0M/eW30qopfd4O0+36VbeCu
9EjOtFG1mjErRvYJBwTnFqedJ/PAq281tVxxl9WtmrzN6Jt5z+cCeq1JzddaSIvh
peLprGKIVXHuPrimRcud8oUZIPOckspqC/eDJ8SBJMFB/20qA7/uTEW3JDCOmCjj
/+bXFLD3rYMyhFdHKesfdq/4UK5aVFEXMYJlMtrTm5+Se3Y6XLx6x0Mk0QrmJIJa
lDg+sLhJQXpPif3GNkkxyabDE3vk6WERKqMLJ77k3YPnHh8NeYq1+ZdyhZozv49b
AC0HTmNmfZ/pY3+WjY9Oy37wBf23YBfDsiapDLgk1voEoLTCpQ9zrsdyZGMuzuak
zUqaftibRRlPRkBrgDhlKB0ncHHSpd4QjVXx24YV8ZWvxIzX1AXox7coIQHoP1ZI
6aSUegE6w9bcxx6KlGeS/jdVMIecaeWfMaGAaNvDddUhzABZ7jVm15DmoZhY2x+X
F5lBNJ6/8LXvhgevH/TH0I+p3s8pHeuyvX8kfvs6SSnEhmx/hpt3enlbcI5U8s5T
JnRlUz3NWHOyAY5b/hndR8oQHBhNRQTutQJygQ7GiOW4vsLSIple2/uGQ5pQgo+D
OLVfo8t+w3MdGZU+rZCQb4wr1tVYQcayGjaYkrNeRpHyJsF/KlC4+kRTVSJCOK2z
x6su258jbEzTMcJYQT2Ts94iHY2IRJVvpBYhzNVKAhLkrhnc/UWMeAHkLR4kFmaY
u+e0Q0boAZTUjXOP7cKPODHXV+CAoql/X92l1+JvDFYBYIwWlyvBikijYEhv1tPc
0n850NYAxfw5t8tQYD3QxKXvmkXy5kEn8GE2JfmQ4Dm1uESoclLIRsk4Jq4g3mkA
TMqCBkiqNv9Qog/8sCXsp+T/gFkDkEQmULC85nzRHb51mdXm1iBXqUsG5QS92eWi
YYJHf+mCp5jSMMvHubB3F9EasPRQ9By1/MQmkpS3Zxv6r5ggiyGSIUeJxrnC0As8
LKlk2YMG7znSpGg233jtZ+KEgTUBIU1LFD3WebWRNrUJyCjyO76qdWbnIyvARfbQ
+Aiuo4OZIG2eeXihcmvGEhq6V+ho8xAONhZPKrJHQe0GS1tfokqdXwae02S6Rh0o
Q2oJqq9shA8UTQAlq5iwnqo0BqTpWAT6x3Hgu0alFBpNFVI061sD8o/hyk66Nh9J
Ho94YAsLCJ2s/2zlcZEWDYpizy1qZ2t8KeZ41GxN5j+gY8YV1QZbrV/drAPSM4PW
0kx/7pkJiEB9m//9p8XSC5NZ4TFNTlNAGjB2QyN3xq8KSmH5JCZfPEDWLFL5QKmK
88Pq40tIk0tmEfHT+toNuPIl7VBc+qlq2ymn94LDuMLGLFMdeqf6kwBIAXFtSml4
R7dEdf6mF9/MRmZ78fWuoYH7bnM7oiSxUyRLiu8YXvoyOUkEgVoK+1IGzQ526d/j
XAHhMF8dfL25MZjOnAMlLeYTwmJN20OI+8eyam3txj5O+fuws48TBqK6/SSPXMpm
rnhz7/YxcX+DX+KzErNNQHv2KM5YUu84XMT5nLb7vJXSIEqGl9EvoOIhwBq8g2/Q
wGT2DjXgBlEWzrQkfgd6s1/T+6j+GS/SoSElfyHBBj/cplLmD8O8M4xuDDitjOtc
AQZZrScfcsb+PgKPBc7Mjhasoad/4gxrmqbT1DiirNh1j8Y3pPyjGwKkhBa81K/N
w+0K+ep2Ii/effQsFsehudP/jD1nsuYazOEsy1RdMXeFecihR4AjOUEaRxrQzCw2
p3D2IFa1At+JXgDanJN8dfXX+N9HirjpNEHp3MazIhjZukN1P0jevfEFdpg1XyMK
9CngAcvn8nlaf5+BEVY3t9tll9kjsKlGjuNrEf5Z05kpSdV6OoGbjJHJNucUFp3a
15R5gtnHpafPYAve7uvdqKfjJtxaRFjrQuLaJBWzxsYciN5z8ln3xyR4AmDW6CZr
SBkbOj06slM48hUUHXyM8vQ1+1OxkdNYIRldNVnP1hQTJ3tLc4bHgldUpXjwTJsf
ArfW/5pEy8GSmsg2R+/skTx5DEjToR+7sFmx2197/X+GgGlG3ZDJhlTGLhNM8Old
Nw1/vDlxOZPGDAqmi+uDQ7gDElD1dvHZVgGcMAjZyN6X6CeYVfXoKw6pc8XL2uXk
1bYDHLWobX+1pUsuUfxrYIYIr3GCekrY3+9ugNpr1+KvU7Wkh/ByYT3mj01yoiYL
6p2S09fF3bnkutBLEGnL3zVAIZUWSRAXE4krJhY5y2HzJ4yzahPaAQcd22eJJSxS
nEt7vhdGCHFfB5d0/k7rDC89bEEViAUPksjuxppt3/jXo/L06D/W/cdj3lCMXdMu
Suu/hfiOgi3zGAUKmMRxdSZz470q8HZ4/hTFyo5Gl1q6yFunKInglDySK66xj/St
gOeTtF/phn0+SO3oy5I53t5OdRPbcVB0ikNctJIbSxXSrPZZOdemGBkpyK4UCRmH
H1i/OYYRqM3kzyEBuSud1aPdtc4YsbGePoh5pxs4P+fm1v1dYEVecvF/k0/jt6Jt
RiTJmXaugK6IJngf/vsDBYCYQWuW/aPO32v6sw5GEy+9S1OFlmHXSsFsLdy60n9V
tsluFTVQkAlfb5X5SyIle7zkYW0kKHmRNMitH4JMgYH0jUgOOSxfPx6Ucj6jr9kK
zTAjFtXYB4mpgnM5t1xQo6yHMkscp9CoAV28N8rZYzEQ/PyK5fmAhJUtcvddTxs0
dguomPLTqdHNHBGGFtQ9n8WEptaJ3QvpDW4YK30pS78MhXOumRl1ewbjWg2eiq15
WLyqudFVgjtr89GKHt8chLYkKzgi//SadLvibrIAoOEHdzz19zqqCH9VuNAO6Ti4
bitQVt0d8TpzuYeLsT6yhOQFLK6qYVqSjbvrgc4UP7wcTWNxio/N9wra4ocgrVRF
nxvfhzzPEmXMmoj0JSRMiLxJgTTnBAXyE4YGx5OqERr/7TjIi0h1U2vJye2y1sqd
5MtRfPz4U5rLYEoTNFp8vTOWH0YuJJPKgVnBurkFYCgx6kFJQnlT9Muwz/IaEAx3
gKQSuv1UvtEkxid44z/WljmdU2RJRJzsttTaLzQjdDHmfh3QSQ9YNR+wByNAEIi3
jnMbjN07LVUuFQcDpkHz465wYOgWDE4qmn3BfwzP1bN/3sAvUpsVIdIP/ykXUrs2
0M9LxtfUxeuZ0xiEg9KPnz5c087iCPo6diILE06nQbfp+7wGUng0b6Jfx8m/rJYt
wAK53umqbEfNdyhS9o2OoOJ05yTwO0by7qaqNapwzp702d2ppgCJiUG5+9lt0v2q
lJP5wF6ntV4X66O6Zz1Z5g9jXK1yzrL7LtrBXYSNrVOnLDcIF4ign/uRLXccptVF
CX0oN0RbgG5aMordZxA3kU5zqXrEcQ8iniAbOfkPEXm3K+5QxxFZxHxdPUd3/de8
uvXpRiGm2RtNitdqaiBDWoVQu7vZaSpfw+sAmm1Rr4bXLRivbZEYnSU7hGnytsQo
idGNKWiQKc2viZdwQKhyX/JWzGmSzuqjVtYXLYn4ZU6/29KewXeRUup4VoAuwVQg
xjN81zJoxHauEqdQYg/7kcv9bpuzlw6miYQQGKe1cutiKFjbpCwm47/RnRzU5N/h
DBGB48/iVQ8Ityh5MdyIOOOlWP4tIlhlAFJ4kGlGwKRfEN30PSDIu8sPZu/vX7Bf
mujNLxFO+/tSymRZ1kEWPcviVv5o8w2MhvnyxvKwVCOx310iIEuUpHaZ6Uje41GN
DNujdvPF4PffUQCGQdEGbMcFyJzySfckQuBCuKnd0ryHQV/n7Yajfozi1H8u6eeV
`protect END_PROTECTED
