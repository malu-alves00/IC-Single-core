`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3bfnZlSonEHrYGgF/oaHanhVEWNfy0A56zNBcFVda/onUVZv3csIJhyvqTkmvslM
OcQHcW9w5NjY0iLo1eV/hop6J2wfMxSBVIiLizpQse+pjhb25fb0Kb9CyH7xdd7e
8TjwWpCQdBLSbPUKKycETQCBtRk69kPOY9ksCqXFgt/6/BxEnoYIE6JfvgMK3snY
FimrUOcqRpVJ6YeASxc/geVmoEB8BpEEE0HKqawCBoOUieVI3NH4p1jmz7EfRhGQ
CQ9BR7gS7k4EiUjTITQ3LEpyRG7LtBGs9cVclGCmt6MvCxTgsBVeN0zJNneejZZB
3KjIF52ta1LwsgVeWvwnD7FCY0/YgN5J8qAfDvpBb6T/IYmsp8fuFtWcBKjbstbR
ToCyXsoOy/dqtcWrY0zz9CjyZ0/dhWWQ/7w7dvIhOaDhm6TUM3nmmWzzOXYEMa2k
k5xgUWzLTcX7ZVvtBiL16/3OrGQLUYqkNQgDQ2qAaMozCWZKuhNto8/Hur5K+Po1
DO3sJ4HbLr8d7Jk2E8QNixY2pTWzFnn+E3bcbCrCIJ8jwUabOKoXnhcNDCC2nrX6
Bx0lq3107StjWMPj/F6BUCJ0Nr1AHYitA39NNs/WFVBLNSg3At3vuJjLwv8uwSLd
Al8LWjQ3K/0yfj81i9xonsrE7YyYmuJ/9QLg9L6x24YuM4vf0+uxB1X9iKrosNMR
HQSIA5sltuvFPccU5qcGPqUDC8Ov4VpCKvedSSGXhxbDWHiXoouJNycIVy5mij4P
ZpxK8xmMbGD9W3RsRRLQxYHckYQLoZ3v0IBE8u8a2/ifZU7h1M9iMqHH3KhcFtor
yFB4LGIM0is/TuviVWswX+KWQvxyR3LsALEQzwjheBLYRZjKrIRvAfNLqef/CR6N
6Vz6aTyNcZQsioAZwiAE56sJ8CwIIvg7uWRtFLVojqDSRr+hLRophKvOKyavks7v
3sF9q98RaKFel7bq8dMm1LgvHSiHiv+CUeG5lyXk587G5aXPvqW0kJi1ah+uE7nI
2PlD8Jg7IncBzFHjGcFcSjJ2JElYqtzLiqm+dX8Ahb2RhTCMVqNvXtercn2GIxc1
+7TqsJE9FjronWqyClYfH+/6EnBlVkpsJXvLp5wj5rXu15FIW6GaYEy79BL4LoAg
qZU1V5qVZ+SqxrdeX6dMBWClaRuNzJdoBOwURLR2QvEyMdtiiPY4x7/h89hGLHKL
W9McfZYWTipmxTrhZRumwyeQUW8tjCEGwpkL0GN3iZe5CTtER1+P2D4xOqU+QFzb
sR8Y0do2RCDL0FFdSChKJzrsrfYhee4b69B1eG52xJxoAbQB5BIfYkYSLu3CMpU4
jQ+WpEcKXrzCMyZfqbDGMFiMA7u6uqbg3KG8Xx8Hv9U2hOd8IUP5N7uOjKcdXz3t
W8mbnNtmEeg+DEmXEMlc57SByWC2cLGxBm761ERYdTveZfufx+EXIEfVsBKzCdou
rp+w8ZfU2YnDoc/LW5Aixxiwx5+UkHAjFc9iuJC8ktcY6mf0PSbRcNtWTnrMYb1m
Alq12ZzbB9RoJrM+f809mGXlKIPd7xVSMZq5PE6V6qy+/6bk3fxa0rDAJ6+QPkw6
SiMT8oma8txd6XAPOkT6nrEiGEeTMtK+6mREqamnLEIi/FASARE0WpXujJS0vP2V
ttPTEbQqYrH6TUSTEhkHTJIOyOczNhMkp4t1/gcuZ8SKcp8WbzhkXo+yNFtkkvJr
UsNsJz9qaJipgYDsFj3HQrru9/bqQZvICkH+25v8Ah53Wudg9a3dE0NtyZIPgT1y
ale27TeRtzrUJkfe3RKDWOHrl4iUa7+FsBDyMxjcRIVVd6isqcQ6p2pqxFMtrDbl
hGr7U+ODeBZvFR4aLQ57o5wLkpwqn3Hs0bU06Wp7sr4DXbtfmHDKHMiV1lVGS7Bc
5cJW6fiiS0GpTLd7HfI4lRXCQSo/2ngYTRfxZv6LYhn6O/9AZALvHgUfNpehSr5f
bSaW+5uXvQJxFgFdLJy6/0EaHJxpA2uLx1j7C1JnEQxu8BIM2wTWDWj40R9JrcKQ
StCnnZwDbvn2veMeXNWIoJ3xKL33rJtK43U2txE9gFwGTLTB7BTU7RGWDfPGStMg
xfftAfEhrSZEP5LxQRd/eGW2gtsF5EYrHWJ2SXZHNrZ3mKqWOncOtaUrYmqbC1Qc
U5uN9u73zBYdxjZ6NavoG8WAVP4B7j3vimJWH+g6ygpwo2xlS6YiXl5I5rI/dWCb
1DDaktfIO6zmvW+DFlsz55EaNnnmCj1GObX+RyIKof5cWOoTtpqWUyswIW2Ybbi3
rrnoVrPWgUPpyiyWk3mn+ETe+WGu8Sszp77PgWsIjsqFGgTkd9MQOv6FrGT+RXbJ
cMFDvoO20X51Yeeu3DRue8OrjnzEw3UFFoECogcochChIt2Hp82Q6jW97DieJUPP
RVcPUCH0SsVIHZVQnIsKkW5I5hkmmXLGjj9vN3ICIOY1/hqNyFHVzE2PQg8kifUm
uIS7LrizbMq9C7JMEwvWLsH6C215j+zyU0AxKCN1ohNvNQDTf75M7dJxYSzXgwr0
YaeBe9K4w7lZvSdw5ZSN/3J40v5Cm0qxJylcU+VTEjX5W5+J/UIvRGy+wD6hlMEc
/Nyw35RRDZ2g9tyjSNlQQZCvL3QG0alKNKar7o+P8uS4kP63j92nsrenT+i2JcBD
gNGAIktMtfZYfRfSwmHsm9kHVJY7vVwavKy7w757IP9v0tm3umOCqziYFK/CZICy
NTaTGpv7/9v/zpVmuc9F5BwVNNEcf0XvO02TWo2omes7tXes52YDF0cwznvv5C+h
4jgO8CbdWaNHTVoe66ohOtPkFriz0ofIF0BXxpHqISHeQYVd7ja4K/kc5wf2okLB
KKqY9TupQjyyC8KRqoIcpNzlD3e2VnEj/3ccN8QDgj9xyOsc43TccONgja4/d2th
aoyFrthB+G4YBFrvd62EKFcKl3bleceZeu614d8y66wb8ZiinwB02ctf4PCoCTF1
btqMsSSkD0aujPPSZNyw0+ynNbXynSM/Uyyn2iImwAVrIUTGbD3yjREW9Ru8vh20
XEF4eKtdxsi2bQWVYzPI6xVNBOa3jEHJbevZHzMB8dC4eAmJTRp093cFopSCadNc
zPzKCp1BiQVEoudrmuAt6fZtQtPFZVTumHN4dsgsKltv36z5c4ZBpSAOmI1GW7K8
qL2V51tXccXEcuDaSUlAn1iTTLAywJDHMldgZ/0vcBrc8bfewuaWxQWBOdlg7ksT
kqPXesJOUajgU50u3jjFm9cycz2uUydlr8HoIbfkGu0YtFF3wJOAa6T8/ppOr5ka
34SIACIZKbBUCEz0iOFHHjcZP7TjNEKjUs40BYRQogxJ6L2qcDKiYiO5+Nct1PCX
Y43sfCAla92dKX0AcwcAbOZRLxivtMYAM2vNCAawmsqPSJHR6oHvXCebOUy14yvC
qq8Bxu3DXBxvki7nKRdLJnEdbq0GlX5Q9qIh5OGYhzHlL35Xq8vH/NvxBoEe1VO8
kMeA+BXVN2IIOJPg0tTGg77kn/v7Fz3sEbcywi0up1l9WOakMrMGcjqoxpXcJL4x
1mxtX9BGaBCAzOV3RZ/SQX6xIjUa5OU1iKP2SqQdPvOdnlG6APRaPj14+dLh1kYu
Ri0QjAXpPDDpuEpa76N/K+rOBzsm5qHoKq0YvkCI4Z3KjJP4BzOmMfsNS30cKj98
omKBYvmQXwZszEl3Ua0bb8tJfjZZSepS+O82HzDj78DE0BGPokQ84RCDDBRd2q0B
F7m9teygvm2KfqKkfV+R//8l4md4SiCU1KEwQ7g5qVul05oQWjVptbsJ1i7Q2sX9
hZ4WL1gmzuXYfqqet6WiGRYLJBqS5ehJJfvsRu8c2Nc8bs0VrbCbsubRIMG/ZuOV
w7YpCGniHvuE6tDd0XzuQKJuk143Se5H3RRKHOAM3bbsxd8YZ56MD4+9CHL6ziy0
GUGvZJVzwwzumkG9wQp4h/Orf+7YGTyCV4Vn+TFJdRXjDQ0Z7emi6q/fBVtLewbn
boSnFTp4LZRy2ALUDqQbTZziwGeXawfZG3iOOTL3QjtkJ4cShBG+rDVA6bpFCJ8m
mCEARBmI+C/uzbInPHSmfMVMNptXgptO7ZPTD2+sIWwtks6ruWSX4IaSDRZJPipy
Tvij2Zth0adAGbn4Br1QylYar85eKnq+1ynqM/msWS0NgzHusLkCHHFaykubMdje
ErgcLVFixEEx72xOL4oBsDsdwTzi8CMt/dF9HzBRguxtfUwBNtJv1qrUnvOPz6X4
YfmgbUN6qPvw5QB0irnk8tbsLONHkQWc2a5J6ZVOwo0CPwK6ii16/FeNvWdG2qlG
gFxgDIyOkWE/QP3TznOOlwY4LpmatutSZHdaxcxTFK4el5gdvNpDBOXLscp+XS1Y
Den3S/cV4/l1ZM4fJCztAEMvYHEx4WAHqGuTqfspQ/nrQOqt4SiCUAnORjSJNRFa
avgvyBgmdJkqGEJQi8r13jB5Cp7fqPBnaK5xThLHF3z7ri5WN5qkOZ1VIs1sfuc+
IQ6ndxUVseMhup4/5dor9oURBC3PpHG+ppF8XzZSvOaaLR8nFfyNlulYxA+Yr9bj
l0v4xDLb247Osu0wXdM4A1xhshtmbwBAPXB4yjhGBnyYFlDn+8OdkaDeK960fkn6
BW3P0xCO1e+YZVuXknXhteuKC/BQdBHbSVCjsrNHQXehDHztBsggEY5eMUWuVRkL
+j0fnAy5Dh2VzPyPs0PW+TfrPsUy+rakwioFcaYyGPPqomOqbyu21itXFAcCd3gZ
MV+7nv/l2V/e/aetEiU0HgH3Epno2Lsq8dza61b0VtdCZIBRPMVJeFqJukS/z9AT
UNZIeb4wSLpp44vQSR1Z2MeNLdjRAz7jqloFA01yw7mKhqGRTbI25uuHwna9cXr/
vO2M0RwxoBBQFyf59GkafbkmEKld8o0iHPFdkEYYyddPl+phf4eqZ03k/Rrine6z
kh3/ND6AdZ1GqU/RJG+45cbMjZUGWurt0rwYfIqV+tlLHVzvkH8550+I3d2g7Bq4
j1UN/ZLYt5bbEeNFNsMsCw8G5pHNJAH4ZoAfmjtIjUXPXkotfz4/B3dgcj80Pkq4
SrE2BoSMnh2WW9yBmTLt/2pq/vTuhycvmSeKO1/xPT/l/m18AWKdvXa7oZ1qOBEV
Xp7nJtE7yg3jmhn62A3epvc4BnIsZkBNGjct6XXluYI0CqeoY5xovYem1Q9wGOhW
sVg8LulJsJV2ECoX0ZRtLVobE53kgwUhh/UC/1yyksMLkGaGvdRMnVh4BF8KSmpT
xjCkgVO0+ULtJqu6HPKVr1iK0Q4hZoVJWZMso/ekN6XM0LQx2s6L2gbNn4e/QcNZ
96RhUM7Bisf2hhC2UV+tBOimXW6pYO1sQwM6pSAG/3HrkJ5qsP0FFbluUX8oy8oV
AivN4oxtGxyHWNsxibMn5tC6KEIW4JoJ+om/DrozhwM9jTWtIN2lTJ2PGnPN9CD+
S1ZWOZcG6e30OlCUsfUST8hg8Ji+rz69v+NCruKcop72XsEo+uN6PZVkW1y8sJTq
Nf7dT6aUPQnCztyqLiDp5TVqM0SGW5AwZxGXFQwo1UbwT57mNbpMhmHvkOb8OD5n
mfpdGtZcL9zJ5x0Zim737D0UOjecyAo1RyG/vQerMSzG33entjANEzIVsKyhwcqI
BGA3YZFx3oLrZ+ES8d6sVfO+uH3usI0J5/sm1ld/BufmwJWGMsupw3cQnhPM1Svf
a32EQlYZRHAphO/2FEssZAqFK+yiq162ujzV/JEuCU6rDYekYrWmiLUO8R6RWger
iIFMOEHJ1KmJ4nVEl79Q9AxRcYLix09qwIt3iZ/MZM49oaJhNYFdD4Rd5tyUmPVj
wRqabdlUtQqKS9Veiodf48ZTI6lMZLm/vEGLBEIScr4Y1BM1plU3NMQGReYk29HT
vmT+g8UwtCtZ5aYkjZkvQI3FIV5QMG/FI9hc2iciVzU=
`protect END_PROTECTED
