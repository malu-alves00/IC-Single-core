`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ow9xCvQDwURg0Ng6YMnyNJmTr+BZ8UcmS41ITtGzoUGzcOnLyygnDovPZQW6T/hG
fEZ1U31fqeIpmZUvOG3lLYNuLs8iQGsLA4yzQJgCTPLzs10Gr7WNMv0dUst1V64x
FHN04tkZYNAO+o+3yiTwZhZAwhkLvxX+qXgl4Hst5uWFWa3xJC+SbYRqr5E26j80
6EJCCpMy2aJ89jr4GWGuuJyFuWlACoBHOlFqhjCEK/bzcoNpVqLkX7qqRI/Pbsq+
rZ7FxrG20CDun53PombtWNQIsHH7z4UsTfAt+tSpiAf9p3apb0N9JOx8uARSptUT
PTdRAFFBXd//SD5txdWy/bhO2ROFdLu2oF24xyWP5EuymnVtTbS2ChOi2a48yKmM
3ox16qNZYjXW5jReSXfjVsEXOseAJZGKMm95X5nmXWar4pKbRB2N0DbiMlmKOctz
ct3R9jllXZ45xhh+AHLJgcL7RA+uop20st4vKaVNlh9poEjlWMa0V6zkVWwIz2eR
UbKzV9Nv9prPNBqZbkmgrevqYupfRKTcnUsDvqJC1MXRh79/t4BuZnl6Ksl6kihw
GIADYlxcvRbtOctN6BRDJjKsNl/+9G7EOBn0yleGUTcr523eVSqF5slXdtJLsezp
D94F8CAdw2VJ/yiMzaodsKO6cHTDV2pB78gpyEYSWK21+Tc/FQHD0NppYjsz5Z8o
AotOGp8aB67Dg4FUbPG+tdTbWchTBWHPKycEpBIijeoOM/9HgY0ZfRxYdsKrqBgS
lOKH3afy9C0teeVg/1o+gBry55LNxAfBCQBcemgBWbSfMPN8jReRZmotQGgTP1Sa
0AOasxGrtKMjUqJjMMiC3EqKxDTUSsrMK7GtLQxtHNu8tzJLd8kGglqZ2kN68uZK
yU7MmKiF8korRjVb1UrvdGMltNIXYHFAEKXu2NBrVkGQ7kDnNSwxiFEvKHKtL46U
AHgjExHdPQycnxB5O90E0SixKs7HxqKmZIDxzkGdc/6AsMpguK+jwOIMxdf8zgWe
cATAn5PwzlXKmbjXS3RYvObGsNzRkrTwb7MsfRMicxmkX9bWV3DcVVut5WPcmleQ
D8AbZwUpvUBdd/c9As/FZ0ti0vnahlXC9k4lxP6yyzA8W1Krt0XvuEa4HFba4GfV
D8gZObPOVmJr7qMHyjvk0dCeYo32Qbrj8MFNb1JoNTtHHHY/Uoso2r6vr73Chq5G
LehqcxNsY8VPg9jWjM3VjXqqWdMS0aJDf1qix9r0OckcDzTsgv4jYGjnNKdmckK4
gCSC84Hq/cJMuJmDNwfOE/H1hrb8RmDOMMyRVzklCAh/lL+1rGlC4wj/TJWuySK9
Zzc/ulJXkVepAUz4WWLxM+nftbY09JMtFsGjmTzFnrrkE9hvFXKdOqRHoHLKUafk
8n3KIzZ/ru07WkYaziRwVDe0N8XF5e9s81Cu9Uz+LpC6o61sNraI6ebyA+kEUED4
JWVfpX0PPwz6OmuNkbMVtp/C+n/KBD0oIY+/KVEjaTEj9sGAi2RNbXJrv76vGrmo
k0PlbP9O78NbWzBQY+hT24jP3ZgaXVLFs5IdDZv7X72MDdEwqIOGB5EE0/xwjb6U
Ls6MNGlqDZSLOMY8mUtKSQpU8QZcafJvsUUgjsQEWJaQOVkQgpoTp3ZKdx7pWpfo
7/Gbo/qTUfN8eFNfEeuqLVbIWF8P8OP1QiZZH9FAyCs1fltdt7ok6/8HDcKJbOMl
bOAkZFiYdy9lR3qyud7kwLnyr15ZbUPsZf7W75pg0Rund/uzfs9d80+XMsdcpazZ
Y0ei44Ov07N2aNJq76uMRQpmWdOhr0XndC8vlkwJR5mKqor3XJkz5Ax+WkdUrceX
+osFVBKsFcc2IeR0s9TbBRHFtLaCKk2xG9BZHOKw9I+Lt66DRGMlQyUQ8jYvHWbZ
HjkNEGtmq0tgmY2hY26W2wMpLCnId44r6h8OUvL+JZHpCBcfFREaXGfL28BPgBrI
Y5LO474WcByQePNMap+bY4yI2a1rhaVpGIpJTN9/UDSxjHbhAtm8P6qlR/PEfSxe
xsbJruuoydxFEUbAhPOvMz0ZtpzyIyU++h1sJrOAKweQbw8GFw2qgC8acGSVGG4p
e1Bb5rmCHZ1Tmc5BL9jwWO2KBu8ME1z/QGfoWa/XJ77lWd4Rk13wyFFPTZopPJK8
7hFJUtRXxU7pOdgbd+ZFCdfZGOaPHpVHNo7mMU5Zc1vxAaSQKZadQTg+nBtwxVwI
7kWSV3zzcTg8W7beooyrDeFhRD33uUKZxEzx1VSQhxV9ocS9qeJ2n7rINzScQESz
7ttEMQ3yTn0ycx7EW0zUASsjGVp1/AiKLpgSE5tt74Y2mM1nTqSySRDwWJGVHcdo
8gUVpWtGt7mDc3L1SQxdboeN1+lEMxi+YaqQb5bfM0VBKmwBnehdz3FklOETJjp9
Fxh7LFBK/lr71wFxBt+h38GL3S+TyNcwcIDYRMOMOeo0f/TeOydbDBGlhSIZQ4lv
rwArLI1CDmY+GEJmsF4mGcQxQrQNM+ljekhsL9PEPExxb79JWismIksJrJJBfn5N
Uv4uUAcs4uEHVL3pnXcrTJhCoIU58GA8x3vqK7FvTJTbs9GpermICdgV6obG4TYA
3GQNkc7MMHok4Imnh1jqT6qRgQvz5zmw9fhhDsNOVGAgyFV0fz7eRemO+1ypoY0v
KrJHW+lLhxmaDmBE3HwADYF+Ic5rzBCbauUyyaRyyFkCtJDzms81RjcgCzivbz4z
s3hb+gUGm7yqv///1ganL1A4HNK2MGdpBxDTAkaDQmtGTHOv1Lj5GwExaqxw5Z7Y
wFmRgICiwLNhZevw6lpcRqb8lktcqKGRYSodedpEbxADIwt5ht8VvOvCptVeBahK
YgfF9A4eEmC5JjM7/d1hc033Cun90BEUvgh7eS+j4ZQ3AKFgg8pxLhoST6r1HiTF
G14I6kKrIRhFFdi8DR9w0xFThxEe7oN2UP4Sw35CPgv/n6qr0Mg0oIQZkDP2f468
RXRi8U+HDrF4hEr5b+jrH1HS8eh58CnjauYecXvm0ZxRgzQj4s7JcoWO6rIrnT4T
6/LyFd/XXNzGI4++FOfgBf/eaCgm/fZOiark+xjDB/LYjxsd60bqpWEOpu4hM5ho
lUiF9Gp3TVHUsweMFLfbWVhdNKBzzZ1srByRI2X5DIF5PSSJgLxnc9BbgNAoHwot
sVwudxjCZTja8RpFYtJUiB36AzLTKZ3A8uVsHSs5yvNX7i3IZr5xk+7jPDepXWIT
9Ni/w4pRZkTtt7aFBKItcGnGomZpFWnZ03gMMGCyAU2ViISxK1/SJh1HmuViUv93
dX+6KbHZmfSx7LQ3ws7aUqZubvAhn3y+LHq1b7ITZYyHivaMM+7U6/vpqE8O3Ktw
+j/P0hvQYyQtwZmFEHqwaB4BdcZjCHilykKuqxWEAPPtDPXuWMYslE3dXFgg2WE6
oithl8EFxcVfGI+sfbFnOVyxIXLxtX5iS8bPs5WLYlMVGMaNB9lJ71uQhLWr4B4R
1l6EwC/tp5rf1K6+51Pw1mOQvW1+NaddRN7m6n36lQ9ujE+hjpEXoxMdVXwE+MKA
HK8gKc1XM9r855pleg6YqKbH+V244l9WfuI5nWbi5ujNhux5xYE40Ug8m2wssrx1
lo/jjvBjIS5HwPbrDNhrbmrdx3/y+0U41kcEtkPWEv3q8vpnjlvP3T4p4A3sMQvH
P4enujSxlfaJAXbJJ620nR7UzJhao7nhVFN8Jq0HVsX+7qC1idgkr3eZnOqM2Mhm
XTj+5khvbPE/11pz+6vk3aFar7GXcrvJl6UbFa7FEj6hKIb0JasGf9NwgwADomyi
uEHUszuuGAqZImkqnWiJYOpm+bwa24pxgQQ6jd+v0RizFkQi6WLCeL4LH/SG41aa
DxuPgupOwx8EnaDDAE2UP1iJZPvbJXRCF5gAFgEWV1gQ2SEeKGdeMydi3NF/caXd
JqTjxAt0iY8J05egbZvL8gCTWrSOGLNwx0MNKvR7c7auyx0+s+8aKhz8gkdr2mMo
yTkKVAtcd8Y5aCXQJM+ljiIL0jIl3Ghj1gh/YxMBbg06JSytMx4QsN+gEqk6YmqJ
pltjMhfwUBGtDJg3hXrQYqz+541t6xWprKlulEsWAbwkPeOBFLDRG/rY0V7OIQGs
Wankn4uotYhoGUlwO/UTaJB/JY7QqO89c2Gua6U16FFuzUSZbBKGm1HY4dldaMQT
QsZSuRY0POxr64I+upXsiX1zMmOs8qylw1hdTUSN4GnwT+yerHdiDq5EPdB30Faq
ksX1FoKSoIMXrkIzZ9htmGiWitoBhW68KdhL+eBQh3ornBHaT5yEAGEesB/DG1L/
qVzD+UFtDkOUkP7RYD/pzXBs+czLpsmq8ylJgBq/9Ym+7x7zq6QsTzSxAktal7pA
r4RSZSob/uJrcKESkRhKEi/wcu4CBMUDvHyUBzO4ibkQ0I22NlP0SdTdm5s829RQ
Sffk3uHkun7ADUagOtTJXLl5595qASXFw6QD7fq0GWXpisH+JtvdAcgun3OVORyS
H5ViTL9T6EG2LKImJ5VXjwp5iTupGMiaRDqIlt1vxAx3Z3M+l5KFkP/gV1HeuCOB
6DNx+gdDx51nDlitv3NFvW3QQT/AIIYYR7n3Li8uIYdAq1aJn1N+mI7IAnC6KnDA
3ci8Ld65/AoV61iTLijTknm8uV6zAN0mUxKqFBReNLCXQCkMtiFpUuldJxfYzl45
hS0rfHiXV5HsHvqgbYSQGwTBpgrIrxns5buVEoGUDqigBHjb6y9vLOg05HfRPQ6I
xgxduAeAAhIzzC/7vdXEAUc5oVHw1lerQ+MqieDciyXl+A9XQbOKG4Drk7sJrzsj
X3gJKYW0BTdOXND+gN5xhotXnDdfl7MVVcvc2yKpLuh6bOLCrHEhJQkiU9XB4niG
5gP8ge3j2HfV2H5yVhzx16s1iZgv8VaLYfhm5pPsjWhPrZ8so8i8vSD4b6YLnwvJ
Ett4A6npzV+caBEEvywPhNnB9u+X19aPbL+TbNkEAvcD3rprwOojUOTZiSYxHVHT
WZzpftAvszIa2n4aH5v3wZKnvzqE4ndRzlaeR/r4+59+8MAllZ1FmyX9cIKUvSjh
zXapG1t6liu01xuXJSRlQ/8Umx3VvIDGAtoKa1+I4qZKXb3xhBVABpkrFTTSskLg
L3vwJGdLBpkwBcSzYj/aVuILjfFdKqjANchg4PbwHwipxWoEAxvAk/5G//COX4R6
w2Y2VrMAJv/lPkLc6w3BKEAL5S58KVrkWwabx3Lwevx+MADBI63LJmgiRD1USBYI
0uVFD/F6RakYuwR4yPztzrGTW+7VZacqkLwt/BO8+quVlElz3lVCSdrAqxmVS5i8
aavGhcrfC39TnC5VuWTWsYA/T8J2ilZom1tL1ZUxHGAK3r5r3bwqbUCTETKUK0Jj
XaK/82Q0dRUZBKpj3yHdYS2V2zl29xx/Mi1/PmJKfQSvqthjs+zCo4op0vFebu6t
e2SqMP8vouAI/YrNiYK6BkynkrIBq9UEzgHVSymQWyOuGpdYi87nRDfi4rcpLvet
8JqqczJPBD3EqeZ1P5e+v4HPMTmKQH33nwPDlCiZ0NwGyXl5zD/BmnLZ/FIOVbJs
TyPGimzO8cNlUjTP31izJos//qJLghYTQ1S0eTJKCUKZaiYYvzPZLZk/qVNc9zln
4O6RuVCOY/paZjmMw7VYzKaIUJFl2uyfbvZAqomY7fZHuob/ou+6R06OBOiK3+6p
ZmNM/wuX+AHG14AHBZCx369a9IB/1AA5Xd4gSBPZoUot3NSxj/H7bbwRvsSkAILI
zRNrX/j6yN9jkv5HmZK2J3MVZmiclgy+WbD3WXEHEnJE0Ex3wlVuemjcIE2/3Lnn
wWByQteghvmaVJoRTmZeYbIA6aaLJnkbseRnW/LQpFJIe+6a0CXbCbRzRxPxPIk+
9i/7uB5MLalRra/+gIckBSBowv5hPEc5jCs8/r6mkKFKWx+Bp27TSk2YLM7nDkqg
owUXsRILfg2hS/STH3P3mnFdYPrmL8v9sqEMvrd729lI5i2uYuZk7wZTwqznhVIe
`protect END_PROTECTED
