`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/REZs+sV89YiUSUGwAJHevqpeSiV31t3SHQjaSNNrtfg2MnXyXCYfabnPAOs9ZKN
I5XnxCNc24/9zpnPmhc4pag7lYrcbuppEGr5bSMPqg9YmJ77/0e/XGwtdyJ7TQMY
aANQUfv+acCehfIRAN5xMnhyIG0BIPsOonpAO+j4YrtlfQzfXPKEMwTkD/2e6jFI
+27nTXyJi5hnrBoQbtEIMEKOhIVNmRnteeVaGlAjULEArMD0rRp4kOVPes2rk7aO
YxIojLcobO9R7MAI9o88WW3Qsvo/Q+k9MQZEdwVO218byvKnm8ctg+S0rKc4o8jO
6lS18nCmBQCjhRNcq2spjq3RMl7rVLumwHo1ByIZXts7ZNXotyhaYsOzaEcdyVa4
ouao18rJK/9AMErjTR6SDSkQFevEP1FVF/PhwSe+cwjeCbjkbf5lWTySara4xur+
XgagPXVVQtYJHn0auQJEwMPcSGeCnCKAZDf9bFF1u46JpdNMTRw/m6qHEqTXb6jW
Ugr0tYjB1Y+wTkhtssO7ga/xW7skTkP280PyKsCbWd66bWeJNOS8fsPs/kLyvNjS
JaUazBsOmP0szcvv8vrXmjse9lB5iRmieQhKL3nPnYaA50CcwP4RWl0OToTl/yFH
EUp2BUE8qSPdH0SpGSc5YeEbruyvhBroM2yzxIKrvavHRay18872j9S46lfQW5Qj
7n3AFOUTAiNTkRzISt7K/X3MYS8XtZmoh+oYvufxmeaMAbBcZ/ZVH5xINzexpy9J
oGjCHFXyYE0YcOKRVfQXBfGha4jJeU2M/DiZYHlqxuBoVMHkjI9HqZijJ88j44j4
xUNHRmFmjPJ2LuMoXMbBSkvaNGMAe32YEGeJH7S3eQ+rE2OIE3MHcPxiXa3kEvDZ
VVr1+AOfYlR1B3FvCYDoa0Y9dO38akowSXfghG/4qwEXSacqUA07M1yGju+yw/p5
gsPrZI465pQvDOQkanc3qKlLPq3qjaON6sVwV4r+I3H6bac2YIWuAMffZfU0tdVh
Wy9wT/UdnCAfhUfxVmY6cWZ7xRHo+SdXoFsK3YhbglPoklezhZzdgiUEArOQomtv
U1ThByxJfHNsXuhbzGX0vmoQuHBAHyoN3oG9g3aL/uiGZcUEf1ABuIzsWpRJdMFy
FXglcVk3exW8nv56jtyI+TJum8eRpQ+9uorDYab+557iRw2JS9Loyr6cFYHgBF8B
Kyg9POD+pcOnPRhQg4VrotfeF+pd23O33pWQcYbfBEocKHy8fjKsBAgaj+P5DvmH
ChfiHLchbOjBzK8hVMbirNfNRxyAfZg3uxZFuDqIm58GRi13pjLPVbzcFxjnl7XE
ajHcXeANXBIi1y2e6niRPDx93cpvbKdOCju0FOEXGX3XZMeR70bVjXgaKQ7ekqFg
8N6PWmGsrpgmVTweucMXF6k2RhFSLG6+PccGzpKEeH3wofyCA8GYmM0hY/AKKrqa
UDSioIbPWJXm2Q14Am4JFOjAEwEsBKZRvgoeWcm1t1NVDAAr58+jiI5SqXiWJQ9Y
yeJnxZVhBUb0D4LeslHT2NF4mu59n2DHkzYJVx5yJX8iGoFvvTp37DukUeMRiHx9
B4dHOW2kaE5/ugvOes67wQqUCpaJ8UzWwo7gpJiMhRMlp27vg5mmquwJ+6TX2WJ0
E7ybeCMc7Yv7AHpK0OGW8ZIRF4cvAvRV/qIob/2jW8ZZO2E509TzeHGPaDTskqWt
ecPEYRvbcIwVd9OUD16gnwD/3Y4NvuK7oHAbxEn2eems16qz6EUdje0psw+PRdty
gv7+VMl7KNjQwdi8F6SZr+SPG2MMKSkdyHmre5EnY9yyJgBzXsWJY8k4nirEzm5w
spf0Kmi30vsyj8l9xCiL8ETIPUTe9UNoO0cP6liw2KHFjBEueBoEzxQ4Ayo8J5U8
C3vdjNLxDlfSSgwf8/qRr56JcU7sFbNyFevfwmU9uq1Kxs4OoXrDXmEnvLrjStvo
Aj5umUtQXsOCaknY+/5mIVUiq/9g1TyVL2V5Y4XjJsKUvQ6oWQlHKquKkDjN14xZ
Kd4mu08Qvh2Vz3r1LSDk3D5QRju7TxcV9G+tpNbLo+hjRYJ/IvYwNSr4mnIzoRqa
zb3u13+Ia6428BqdR1PO+fdMRFsiqc74KPmwZ8HLzwSySCsCP3AMvXWjpa+215u/
ZZnLW6g3hyvOeUVYG6Ov+xJ/tQDOt8P20FDIL/iR2DBe/m91hBtCQIl59WvNMdzD
AUMxyRIgFy2y9knK+SFMqPZnIt9nA/11aFl3w4rKSYyNUjt27QLInNC9JoHtECKE
PL4vvRIzPt/oQ+lGvGpUbKE95MbS84yi/fda55JiJqhfkttZ+lpFgVlrWKkJA5AF
j/ODKLlXgoVWI6vgUFXI4VbkC2zsHXcc1mg3B0rFbGaWJLj/M/pUh1gYVpE6Av0F
T5nTYZX3bLPEQz6TofB+ORETvPoebrjEDtxEs3ObnbYtkVWaLFtRBUxDB9WiYwg9
7lj8NzcCw8bv7j4v+nNNv13FmlUMSMpWAIbfOwEgWP6i35sN2PbojVa2mAnEpB3x
WhcbKsqcv0qd+biUUtbVzXJU3IPDmyionpVHXQo/RDasi06ndqMdb6Xi6Ys/SxBS
0ThdwuhOt+tUkdtQF7RdzOA/8Hpz22akwh4dU8+z3P7umSMuq0lytIiBkWb1rtqG
ZqnLqon3dD0PFagRV7sSW3ss20+rAfw+LXcP3yLNCegJTr1MzEmd4MZ2FQZVQMXU
rDv9yU96g0I9l6pGdZmrVhfRhmZ0iEM8/QSKAiNmspYdKBE9XXH9R/5F6n9W9Wcd
M+3uwinaD0N9XR2Lcj7diJP29pJ/pjR/taXOQ9hy3dxSr1isJofFJf02d8/nE1GW
PPUr/wFqLRxSicU/3zGT4l9zIegmgDfVDZJsidOMISJJ0GytB0ap/I8DpdQOy67C
j54UNt3P30o6MTLr1ZQ9h8/lPPvzG5j4r73yj7N1g3ibwyPyuqFEBURMwvJJoexb
HJk3aaZEbF0/iln67ezroGaPikfaY0wgoXlRd3NfqmIQ+OmE7LmuSZ5X5nTN/7RW
tgYGyOZ3MmkIuGTjNlmeX6zoRLeuiV/PEumMAgdCmbayYDZGlbAPtTK8yRMxExNL
c6sTnuAOzl0F6LbJVCYV/MrflcTSf6LgP8K4qWqsvYGYnbH3+rMBMGpnK6tzKM2L
cKzU4GQOBQ70ortXbmO4lA==
`protect END_PROTECTED
