`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FHx2KzjdB2kUn8j2PzxUR7TJxbpHn8Kb8YR8hmc1aHHA/+S/xyMxrHsHgJkwr9qx
vj+m5BI/azbFk4lHAtGYfx/4DysxdxvmK64nVG2xO+4RY5tacAY7AI9JPVo4XNVr
3jievaWXqKXMqe53WZnhyzT5SmhMII9nul10x40BvFDYg1BK1gmpSKUNPQBcxmYF
oVDkJJvHrC13WHuBbuSAj0zZlns9NhjrsFOauG7lw97WDgQIZS4b3lKl2DjouxWG
cw2BVs+fH7LdVyY2rY0+sA==
`protect END_PROTECTED
