`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hREgdbTERbAIx85E/MpEykpDA3Y7/12UYudrBg8wV1kXxbneJHMUmo51ioecofRw
ehtxM1gBbp7iZSFRgtJlDqtR+FsLgQ3rU1ArzVNA4uSTxbvjM3VPsCHkme/Dwg84
hkwWwDUZu0wWe/9catUZRnwBCXX3opVpZ8pEVEvU+aO7M1FcCY1RQzwus69hIbIR
8XQuF4QTmanJyAbIjXvcOZyvFowJcuWPZfzMcRALZ4SvcXutTUQJbYdQbA+CIxpO
ooJ7jMtt285pX8JaL9w13O2zdOA72OeztbohOrJY3aGE5JZO95wWGiehPVrJWtns
EBxS4DZALDXQkyEUBK+7ecvVNLSfawIDmoeCim4/J6/RpJYSsh6yvLSqa4u6oS9b
kEcLUgminTIFZTtdygvjhcuLzn/k3cBl6cLKbIpoA7B4gZEyZzq0aQpGkOcdChJ2
DrYq4IVLtPBPcLN3Ku0rM3A2+icc5xp0fPkCjmOWhSNyQTjt5peq5A/zTrK0jWu1
1gf7LFPF0OWoUq8fT8MqwyPG3oJua7xPgmKJYHX3Km2oGHIL4pIxGDf7jbWqSX6Y
ZdgFW9BCLA6NI102ROlEdNwH5yfUxEMtB6nH76GxDIegeDoAr6JVkeenXrolaWMd
NYOcjrr3ZkMUDM9kOa7jybIkJzVZEXa8PlctuDyapUkEzGI3Y/EUdKXnbc83USYx
r7479DdtT1ddjzePf++XvloqymbUBXLp7G2yoiw/Y+5ov5eLMZwx8D0HAB2Jdeqz
kN7E5Ap+eTH2vYbpuHZlH4OIj8bhLQVAK+K5F40fngnAcsZCuyAojvSeIdgNyTkS
psNSiInRONYomcfGbXYhD2Syh9t9629m3j+deNRSeJcwvmzGqZtQ9hRADPwU+DKl
6qosDkI0qoEXeFVceA48Rd6LDf5KiWoHAlkmigeQAQXz/QG2mqgF4GO8WXWP5gIW
LUvsifA/QXVCa8Jm9RmG/58DT9DVTWh1O7zkczFBazAg04Buo3xLte4AHC+tzu4n
So9plvT65HFaif7rMe2G5g==
`protect END_PROTECTED
