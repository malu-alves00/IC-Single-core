`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+HmyPHIbAe34R07Qo3dMk8GTtnZqyBnJYSXwkmMkRzPF2J9CjdZuvu//8NdjcfDq
OvXpV2ZeHX52zKj/UesyXlhuxQP71IwWM+kwgSGMRVXqZBDr2gGMCu9AVKFZR3Nx
Mw/2Mn/SX9gPLr7+vIp0eLwj2rfd2Qc8RjlglZ8IQOaxA7xSL78n07lss8Qo3ElC
CszpL0mt7bWM7miknj9Q9fVRjh8tsPzLoQk+ER98vO4KABD6oSjLqcBfECTicsic
FkmcYZ1PHcFqlqudJPoDKIOs19coeTfueQNc/woRsrVSoGbXpVF1GYvfrFsmlhUS
DCn0F+CM9qqVSd554KtzqH67vwFLjhPmhZNIxDdzhiZLmcWofJWVV7V2qLfKuYK5
kmq35uyc+k8ILytdPb5q/5VJfJZ5JLIzzOmx8ga8500paL6n57f4pUlZCVLqrs6k
g8iqUq7jzhtHmytqLCK/GvII1OWCsCkchYgsZcbV6EIwC41YMDXM8l2hWq0NtfUS
0dnCNPQdieV9rIoPWzgfCDJjFktjzuwUk6Tswkb9A1Iz6wupMV36ykXCOGWPlLHd
1IlQFiIRM6KFHOvngAFfnlOR8eMIs7suorMcoTnhjzCkv/NbzsxBZ1u4TXGhp1rY
e6mFxeF3R95v3VoTxkgGJmBb/102IuymrhrSb1SHMGfGzV3PssKTY9QCpSM81a2o
6VFilRunoMZ4zqsbiSnYxxMqXu3aZqhV4rYDtbwDbRzFWMnWBFPYXCVSBewQuiJk
ordjOddfVU/ao2E+1QiMlNALsYQREI/kjCFJaTjgShxOG28o5Nd6TgL4LDJIDcJv
rAbwrgyjt08qCR2eT37tVau25v6RwAtYeNR4D8KA774C7XZtox5w+odvbgFcRTio
WvPiaYSVD73rsK0ZNaFustSHFBNbk9wvwLdSlnxsskkPV/fXamC8ondLVa5YhTqH
j3429pVKW/qRjRMUEFi68qrbU2r1PGGlWzDjDL1D9g5NZ0MpNk3WhMaLhQNYbYl2
XXJKFmWz6m9F/4UrieMF7x6qynOoqQWDjDoeCGA9kMDLu720Fu82ki8P1ZzUsGwB
w+hHbocdI3ZmApkPO1u0BSnY2D1pi8SGpPKHEpA5nB9OkqqyPI4/5yIyls9eewfj
8qdVPEQcfefOiTpK6ZUxKzkD5Xzfu2Fno9fn9OHNisVRCZZCJ7rEQZgGmkJaJ8xq
P8VC1O5V7fZwD5EtvoPi5yc3ArPdfTpeIEBoFyZUjoLxAn6Sym+Q6aJsllom2WFB
M68TVcrzBw+aTtsXDAPjq6tYrTNtJxzulktxpgmSCc6rED1rsIN1nK2TeVIIdjTP
tNeLS4NhqHIE4KtvljBuJRazAId3VJ6tMHp8uXrzHA2PwRf7stp6RIGLL2gh1GBa
asQ+B3xTyQxAue+F/63aLg==
`protect END_PROTECTED
