`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
x1Bx6QcR2vqnaFU1rO+l8+qEumFU8fQueDfZNNSs+8snt4zFacyyLNiGFo1i5qT0
ve9nDvuDN0CfZS8tmTkyFlDyIxchoVtgUlYDnV77kVkkDulBVsTYsos+YOcOUdAv
hqWz/F0Ub8x2bHqSJfIIYXusxZxwwVV203750vt/Kwnmydpcmo3geODz+QuRFAuk
ThgiGvzVOA//t3JkCIfqoZt0lgToYbADaNNGbSVpk9gVfFiBXTlTCHoFa0f3yLOr
Hu0UvPia2r7uV1BibjjHX3cQzHdPfCScFY3im0YNXB+j1ARP0key7c9QYL/qt4FI
W5TB7okMqZyFe/VZwte/uH2yjZuGZJct2YNDicT4esQXWpTDEXsNGE94MRqCwfAU
lWwFMaEjiGy0XxRZwmx1J1rB7CyGSRkbd2WkvjVsQeIyA53eYh5X8fJFwvno41t8
SegiNXa5fc27Hp6PnpHJzKQnArVWqdMtyAOSh7W+orfzdZ7kjpXiuUwJyzdE5Mjc
Eo0Q5l0SOgr4WPUOQA7WiMXP6EwBLnhkhCfD0ErwDpD292lJNSXEBgVcrm0N3SvM
wjBq4bKySey9ghel2ZMbMn4gSDc1xGMJwfXCKc0qT8m4YE/miq080J+4QhsZzyq6
XlsEIYaG597wm2h5aVsfeQ==
`protect END_PROTECTED
