`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
R8h/wi9BQKcRC/k0q0T8K0UYIPWVSAyrx7rEMLR9jHwoHv1sZBaohO1wesqD5lUo
XBG7Bk2YhFAyinoatCDDOezq+nvIukNOV4LAgUP5Tk4/dlzEFDGFZ0ZdXpw3Wjrx
kk8OjINfco8Lk9VGrjPhPiBuvqyTrjSWc+QbfKN1YWx92AOZCqOMUCAEO87uHVN7
SpEPErAQCJ6CW6vvUoVY99ns66J4czcBWkEZCpvBNXvWJStDbCGObZbcNxniJy+y
FNaDiqtB33liCudEVZ6aKrYTxcfl8GQhmxdIbWQmq5w9R/1ZzhgdhfWzbQaHNTG8
lX09Cb1zTNGAH+hKAHvo1jE6eZOsR60/6Tu0hv+3cHM1VpWf5KRG6EL90GXdHhuH
EivqsRoxtSasCIR49bivGdNnzzxmpL5AcAdLFeFArix2es/tJRi+jPbQkTefsErS
t+Q4e6jF0jhAhjHKGAoY/+w6WG7hamO6xfNw5nMVKyY1i0NmqTIYHrALC9VHAhUX
Cs0ljlSGjnEI66rcuIGcJcZHVJt+RRComcqbjFwTzp+jn3FQtWk3XUCZCnIXHKms
iBaQwh4y0KZ0aiGEndpntKW+2GCY086f4a1jSRCkUVkdrbUi0KECKibC8CQzvcXd
/aaIHIswKvVRavhdFfEqRjPQJZuYvLL0rUBjCIlZxFOHPK+ipHuzgXNeh6u2f8w8
Zqm9jPtv5tx2gj2qgOHqRzRraAxzvkOb+ZyC1ogTJ8bNXQBRVC3AYX9NQjx632ns
l+Wl2c3tMwOC2ZsluE3dDbxa1TDXjnU8BWVluJ0k2qIbUl6xl2YDJoDTfHpaK+pV
UGXXRw4YGWbwisL8bgT263a2LBSuK8vaVV8mEexZMaC6jb9wVcztMpS8tCVqjL8a
cTXWqQUmABks3rvUcNSlXK3fzZlyPAe/9wJ05C0K/QVTJ8HLLWQFYspbYjnCdXLO
+b3NBFGicvObrDIy3Ytl3RWf1MjPQGZpb7gH9kxRPz3+g7tBCVY8t2UqAix4j00V
Jajms0wYrzvpG14g7GgsSPqaSLu7U1nFy0HQFr/RubMRIdIehad1nlEIQ6zh8LCW
YxjAIZphFlrSTNzC9/QcXHbNo48m1fzjSf3sXy5+mlJ8y6ttXPoM+bCLEl1GmRIg
5ymUMD0OrhkHqLQebqep+Jf9ZtuOh1oBlJ0lArb/UT5Ds6uIpMi1s4Is1h41eFm0
DAbJd4OZ3gkJWiiZ+Cm026k/Q6Sa2OeTZDRB2L3dwwsuc3sZrG1FvV6tZu7H66H6
y0kHwwwFlLoo8NIZVq9A1KO8Z9VLQYauzJS1/SVWEIwrjE4+tedz/tyNxeOcpcWH
b6VSYgVwk6Oz00YxTuok3S0aN8GJX8LIht6DcmMXrqOzJJ3S242Y28vV0rzEkIlf
Q2xzbwgyWcqhO7Z4UQyWnI4iZysjmQ+tic8r+xQlt1XGtIVUt3/PMuctijCZBnxe
dHGdxx1/dqaNSDM7NyERjcAP55qkzFpmJIlGWtOFzPqlQV69ZrZqsam5TMFQv64i
Q8MY09zhL3Sd3xKJUk8UTc70R0Jb1eAOfketP3/FEvE1B8ZCnbZ7MImuonNiTGTK
GXqnqSGQ6IQrwSwMR7JZicgzJn/SX6337R59UQa6/1uDd3eIaC1CIjFlawO1zmOx
wlbaEIgsx+IlgNRsH54bS86XBcT6n6mteysu8Qq5+rYA+cEfkCagR0qpx437Agvq
/RxZ+QCVSR9TY99URKLIF4kQ5laKqhoyYSqElMYtOJ9gE3JavlEmBdnygmw+254H
B5CuV/gI9BsEtIxDTXv2RsemmbymeyxtdShmOMfsr9ZsmfZ/0F8VLu3N23EI9sIg
gCIpHmZxUgY76xQzhgITu2sjLn90xfOv8dvI7cjdCWHUSKS+JEZgfSbb/bTDLTyf
OW6GPPSaiuOtSlkxEzkPqcQyEiNN4bCpd6JNXog/Il8urFco+ebInwEcDtQ3oNug
H2mZovdWMMaO7/dnVP11WMgvMnHnT8UL6QThPZB0VNC/mOKIEP/rSQrVw8UYJ9R0
o331eEezZYsiQuLrUZyBAfNYsm/nEnYXq+wVbdG0MFh+q4gt6KMGcDYZQXO6yw73
OIHmyxsQ9L9PB+u88wZCBu2Ws8ZpV/+mhohzW3s5pgoVemT5dWSDwYhTIVHcsP+V
JEEOHq1q2rjOnszOEhF7guLl6TP7GT4lPfqdf6UBW6XuEhfLfIsn80rvRW9ThugG
+05vDlEGwTLtNRBxx3L1ndjQSJnaFpSV4t/CY4cNVE8VchBMSDJbpbEqaWJN2VBQ
Wo0UkkIn/vmD/RGyprfbp8VLvxG6uRh7Db1w/7HRHkHnufAZgFuJLzTX14majGK0
xygpd+Uw+n4XUbTS/YRpnNa2JIlsOUQ1hVvlkJbLQ6wZDDYosSviXdRQ3upWc2Jm
F3cF6NxLdXVZ0JoxDU9+8XSsubZmzsqpl1EulD+EHnIib3zT+CM2TN4r62WVOFHk
1HvXsLbH1CzZOTJUQEZNOo+IuZsIXgGX9d5N4ewPOqo=
`protect END_PROTECTED
