`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9GtFtqelclZLzBHb+RDc81Q+Ki22eQBcyD/4zdCXPJMeODV+2CX1p8nqglSthyOl
aLrs69VQhXNO6R4CugccWyGRTPz2jHYPfJoc6RvhyKXIjM1Ny+lkeAtxlq7/gHg6
oUdAY5ZB82huj2yhE1piMmSkPwjajrvj7AvuW9JGNQXp7kAnq+CQAa/2VWRePnZ/
dkMXVCKmZhFYe9JUqFt8KbrVVKtXkHPmlEkjFrjIAYGSykamX51rj8DiGsFV2VxN
erl9csNCfJgVHuMzDhz8CGnnrugP4U9IkgTWOVubTQ/DfXH5ktZVhFL3oc3fcCjI
AcdJ4SLAJ9ZhT1OAV1MnQ6Wq5n8hR4pd8VcNqXH+bc1KmouM4uhFsvz0R9yHjYbJ
feaJjtRZ591HTYpTKGjLS5EcnMgZWyyE1xCwkQiCNmgl9OSYnJ6BANngrwCwiUOm
Ho0hIGEWMFZrLuShdw0uUnattJfGVdO/a5g5Mng1tuOV+WT05ix3Pp92fJ9SZWTj
dULNqBTM0xZMfkTOULDewiVgIl7eDba+PaLDMYV/EYxpkTjWIBbNnY04L1UozMo0
kKKUvYBAKwfAcl+CjG3M0wkGdd9jcT6fs1jkx0ehB7azdGV9yuNNSfchQ5HRkGbT
vBtPpzK7bFMPRPqDDuJbp0GhR0s3NehYAi/fCS4niPnkFD4Bi6rNJIRiHQDI0Atl
6F0hF70SvNxhGFjii3sNZ9ijb14oOIkEPMbyjwJ0n/ngKSHrKDU76M2AYSHpWQfJ
W5Orrfye8krR5N0ZOng8eqN/eQlogu+uNQNm8gVkuxbEPMZ0bp3X3HFVViDdJHhq
GJtnOCUxPBfZKev5QMpgQ4sbJ6jfR++PwnI3RORT2QlUsDNe+b/QNYdrmd5j3MOe
fFzGNqQ2EKkZZUYcoAaEUkuwecRS307wXMeFRi7L+Q+0rj4Zrsb/ojXf1zN1pKV2
ycayvWuZq5GFM/zF4MAgaPrEoqyoyzobZkQhyQOVu0kct4O9Up3DY3pQSJaONGYH
UC0HqVbCT4sCOVsNwDjQsWBSVsCPDdZ6wG9f+2q2pOYW59geCOEKvKA+B33OYNdh
pTUTIB/PGprQb+DpEfMiTqEYDArY2N1LabvhPeDJS4MnIYFXBUCvmswSTm4mY/t7
rbGbsxdZksXWEzHuuw2wqMSkZL399a+gjrug+V2X3RBnEtwvp6SAHTH4OeB6FRnQ
zPUv6VlJjR7lEOmm7e7QC/rjvLIaFipOOFh9gmczAqN0tRFOZMZ5pRW6vGRp3vRP
mfr0XsFftUk+P513g7LYmCQiejlLWYaHfKqxw10Wp/+1ASryCpi+5F6DosqYH7p+
BJed7ekKWDtR/hywPmZ5MABaTEQNojqffPGiYpogKGyX5fFY1oQROEiY7qbD1UZf
znxNffv+l1TBXrr3Hd510o8Jo6CNtoWgtiS5a2mOkoyUo2VqMT1s/E46DAMTlKde
wZQgFDlWN/uO/jabSInAkUh7mXjcwYBUJ+kmQUlDlpsl2474B0fik2uibOxgMmEK
Qn+J05Yy3vv4z1qtcPYchM0IvuIFUZSLREtmRo8fjKd2F4qSGn09MDmWnWVDeQbi
pSJsoRNjrr1HXHeF3HBQRSA2bWoAc2sY7J8nM8HHT9Jhv0bNRJbVXgtlFTj6Pucq
OTI9MHIeXrKzPk/a4/n+cP6wL9CREPgt1hUwHFOOlUWsH6nkvv8Cb8pNy2CFuHLt
CYEkELPbyABZD1oZCs7ApDaSkNcSxKc+ycc2VxrTbvn8mwVD5FjyNH2ftXIBsk7d
w/2iaSU1+rGHJcJGI8AMNaGQ6nu7VKSpjhGO5miz7vpP/eHyJVeaR+aLQ6ZLf0N7
2ldzAZ4Tr+5fany6LcdBLww0xRRTPhnb2vpZSovgjxPTskDwX82C6RXFbBYq/Ogn
hAmvBwLbPgXH1oj1yYgCTXC7HvelpxveHkGrr7WLNh9plUtKo8x5eyjd+uKS90p+
FlmKh/HrIONctNKlCnO76hlBF7c11bU0rMSZBlHGeq8LeaLstFK744PLkkkudcTJ
7eyx20jsjeINKE/+1PNmGRdl/YHb+RWJfFeUnr5QrBGzs9ylnecgwDR4JVCxhjxN
JI9y6EKwd+BptN6v+fputLEQ6fHiDVpHDH4Ckx0G9IE5vdzgA6p5semPFW+/7OM/
rW+rHPtavXP7ihV4gh2V4wu8AHLpmph5ADGC4bkX53nc6uwadO1Q8by5r4wFux/P
8x2LtQ3WRhljhwbx4xnL6R7VEobi/axtKy+7qKNnnETekTTdM9SwlJt2VoMzTAI2
2wGm6ThPAz8IlIbMWiC67fEt66hY+tfRMd4MpJj2dWT6bCKtZ5UQQ5wZs3vXevb1
zlXTPLGZfj0tCwL4HTX3eLFj1QHFoXX+JuhuRckb5QASnmlJDPr5WEi/TolqGR9t
BA92edz2PemfaOHlhjblxe9V5RrUYaR88cX6GLgCCSQgXof1MBgXhSbpBL/VdGja
zi+GJf9DKqMcKhX/RKlovZsV1t+z51aAvLu2sWmpEWSF8D+tsdVN5OH+JTE7R1oD
RLh4PxSsMZ7YuRusRp7YH5KWz5CCsrQcq49dnGYRKgfJgGiyn4TWK8YSvADhsxZN
zT2opA4yo6omaUPhTjZ5hAycUkfXjZdhOzw0VLvQZuwtit8T0AG3c4HdVQWvlEuJ
430X0PUpezFWp9W/1y2z1A==
`protect END_PROTECTED
