`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AYdVlzH0gQ+wQCATrJ8vVK7Kq0MXerUk53Q+hrxW5y38x2N2+0riI3tZI2kDmlVL
C62f+krLHKD446o+BfYCWlC1RIDh3Mz7hQhDHdedeOo+f/pLQd1R2XD+fAQTEzTp
aVh0IrfcdT/Dbji22zQjV/zNntscl+iY0wS2AhDCwPWEu0kX3ryjrbgaFghtowxd
8aHkY++5tUXvkNBP57cdFTZf95isJDtg6o7R4BZjbGD2Vs86BjQh8scejUbkU9XO
vUAZ58hZz1GpqQjQpaj4SYVo2zpGWfqcJiuKp5qK2qUQyxNjGv1ENePoD4vJYuZ5
4aWngXr2Y94S8M/gxYpUhNMHOcpYEUkpKj8cISH7HcxD+Ux4hUvJ94nLrpUAO0zm
vH9UeDf3iGN4rBA7WUmZglw7YHbyplLCB8uy+XhGwVeZrPynW5ZXh67hRbUbXl4c
`protect END_PROTECTED
