`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WNSoPMHuOBAyaHtCTYTZc54D2gVt2ecUntaxI8C20tCpLGmFCoKJVM7WzTYiUzwi
/ZAxwhvRjnSz9QEhdO1dTbntjVpKUePfeBXcKfgyt2l0LGA5Ryfj6NgY1Hd8i4qB
bX92LmkRWvJTBA7s+ZnODFG3oJg47kLU0VNFQLwYfXLUvyd7Xj1UAx5LJ1ry/Mwz
CTA/DJddAyO5/MWUVvnYgn1ysWhQ4en+OgMTCYVtPGcg48To5KiPErWgbHMrWmol
S1BNGVQ6kU0XmkHB7KAW/A2B9a/A/FVwQLFlnmGtXCk5151BS98sZLkX3qlC30KV
okVzVwmPvdckLgXxPlr6tEggGZ177PePmgXnntUa75xkTzOFMrI5wI2Kb2TVCP3b
oNdT4DO9Cx/HsdjAStzZ4ZM/ntqVwqIRMTbLS+29dSHnAD97vIzP6vFs4oBW7+XB
ZCyl4p1HMv1pkEZbWj+eUnAHk8KGllQtYOYYKMbCYfZ1H4Y96gWZFRQOWyvua4q0
VOrT60H+dDs/jDCebMKzWJIJ6ELAkrnrpEGrhBBHQWvzkAzkXfcjW7kpVGAsV1PD
I3EBHeQW4uo/A6cEWvhrarMFxtvn+LOB9XbMaKkrleG3PENE7DySNZypReFCDqGu
sPWrWEpKh3fY+Gr8rhqlEWsXq9mGh0x4IM9g2+2grIS7+7PL8V6Su3N0TAVz1JgM
315aTEe/k0lEGkBy+NhJLUba8eP035FCzd83jNTygME=
`protect END_PROTECTED
