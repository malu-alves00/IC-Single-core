`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OEb2EyiHRKNzHKTw/pc+ymc0R+slmPV3QghdpGGtJomctmy22r0GzpVTZOrAOHbv
KE4/RG7+IqGJG9b/qRdEWJjhu89gY+XmOujjBgU2GGb3XDbbFIzhMXL6RIsau8F0
NfkmwGa100mC1C+/zVgXo1WC4bbn+bGfH8paYGDlxtkW+3R30lsvxOB7GlojZCMX
KIzvXGe5bdePpBMBzF1+EMsJKSS/oV820FtjXipvqAoFautq0navDsuRWJ4WCLZu
nSuehIOM2i7No7WOVpJpBhPXyuHgvehrsFN9U/X2zg5Ue0SmO2tYxfCmRP6XESLr
Qli8+pKhlOlFEK7Q66FHGAhbIkd5ekN6/8skhti7m3+5zJMUhWD5ESMskArcu2On
oT+iMDJDZQZqIplpjdrw1VFY7ADJKU/QtaJDnAvb9QcKYnBCNuuBHPQX5KA/RXVk
uXXYrRgTuFP7ts5XGF2DLAsP5X3I1JlC2wYUIysdP5XSbe/V1K7p6mUjxgMnkPtM
Rz5DxDbPCeF6uYqMR60VpnaWG1fI+b8kyEDdoM2yuDn9hHRfWG7pLwqkzekqwuSz
8LvQ5JQ1LNk4Gaxiy+StoMkMtk6bXOyFVsGHNvpVdNTAuvO1nnJhoHhobOWZ4BQj
rtQTZvj4oZ+Je/n2dWW/gadIt35fLbbySWaTIWC2m28mlGL1oxM9E9NV747+vE07
zbmEuyijjfSkavK6xMEYd/mQg7/KDfFRNshYo3GFsoQM+MOumEdVE5VGvFtfI9dU
x+0OUm7ubXebdqRp4gUwWrTdFpTLK97nX4gd39cpJgsLaASVwIhgWbOkvrPmADrj
rrjggvVOLIWwubkhdDuLnP/Won1uhgeK0yzbv6m03cyx4oVlNRiLJIldYSCONo5t
qSE12Q4elXVBorx4jA0cdg0Lhe4ngCogMsZ1z3r/Dpjt0vLMUqd25SMv0i0kcLta
s4M6xbjQN49861iSXB/fCMdfbvBWWU0P96Tt7D6IdYYfd+dc8chTVUd81lNdGtrT
3wxwmaNfsLefl++dWn19PIscwVjjs+EkDis19p4r+J0w+7PS/6vs7+7EMnLVbqfE
Cghprtuv4e2/adisHAGy2NpM4Ht+ESLy7yqHUxCo1VcHifObtt6mDOGXwmtqWxEY
zJrpXij5jvSrI3UtrTmQhFuEcZDRb74Net0mWZ/jo+/P988Z+UxVCoV5yXKNbDMc
aVtA9doNiz21dceDRv15dAKRZ+5Zq57ZWw217SR2qqq9aPHmZ+D5IFwGeiYSjQmZ
6XNha6Z84EmtYbJ3utq9zwQ3GrwYKL7rTurDwRosBsjJbQaTmP8/WSimqtDWMFei
U9y5kP6Ih335P1Y9c8HpI+ymLX0e0mjnzAIgkrEeCLAJ2+BZFzUQaAQxPEMzPCOB
zlZzgYDQDDyyWn8xB061zlLLzItKZ0s0UrP3nJ2nQ/gIVGzmkODSNamvFwJOK8iP
gwpPUObPIp0sCAOC4LK68Zp3cipS0e4TMKHk86Zgsjsg9L5Yy4l6fRihiEeTk1mF
McKQg7ZfXCeuQQ70TJFmaYsSzGZYlQ9TPWdnI5pJRGE9Ywkjjda72lORyLk4aoMy
m9KFDNb2/YgC3uDYgCYHidDi+KV60p5Pra8+/Xkb+a1ux8KomZfoS8DXoafJx1AD
XfIrpswgbH4Zo7LclJybV8fa/P1vg8uWfqg/JoW0Zfmuk7UxTG0u3p1PpwvALrBo
zf0+zb16j/QiX584ow8N67W3Xib/O9hK2EG922bOxU9GY6O1WSoRKAd/QIP5q1u6
R8pW1p8h2T/f5YCOipxmww==
`protect END_PROTECTED
