`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wxYt6BMiPPip0RJrLoJRatJG3CDWqQNCdcrTtZ4zB/ScoscINHlSiF/tHzpLKkz2
Nt+JOcnStUpGTTyswDJwm2a4lMbQgcJdnUV3fA9plEeuRzj5SqenKlviKrjBIxBU
OcP/8HQa2CYddOCgIZSrkvmzwCBDVl8b/JLBpnCgzYGlXP+pa16wPC91b6/qcf3O
YrtD9ix8LRrhoFOsuxAXIDiI8W0+i1flk+F0oK+Us9r7XOlY+GUW67qAV/axwyPL
Zpdb2VN0DYGEMphUssxPCt3i3REuMb7rz91e9SSpPQo+B6EUylYYhvbdoYUm41Bz
8CZSSOeB0UnVeFQSg4E1nI10o1HsiuGOgQCw06PA4tCr9Jxtb+HoqTbBnqPYZ4+o
RQejlr6RGjy4PEkhPA86MyvkzOmrpjGx0FN53HJmEeTlc3eyWF4+OrtV0qzgyMYk
t3nz8GhOOG+1Slk9IrIZ76Zz7KPdQ4ebeWdGyqf3455puBzPPHG4xisjiKjiDxZs
fekdKKvVyrHwnbAiWkxt3LegIgIp0CMvUnzFpFUXSfVrzKQphnUQHIB+OuKGoU2I
JOThyjk1M40rZZjySQt7rN63VdPrbDDvLcYGNGfp1b2RsL0P6qE1CUPcmA1Viv6q
uUwapWY34BnEX1iqWo5MV6UNQQG0fWPHnX7oXmVdc7phLApLxeqKFGe1EKeUhKh6
f14JhtH3sLQ7wrilps4GytlnGbkVL39BZCcA5yRyV65+kGyRTg/KHUIlCXGXwpIh
UpHL2Xk4LKy1D6H4dF9aOxp2QfUxkkIF3okK9gJejfs=
`protect END_PROTECTED
