`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
S+ACRQGjCynFGhlSc3BzSgI5e/KxvOtbfDScBzBNyOBRC1NwcDvcUIwkeeqocNR1
M8IEcsH4vuF2ygZ4N2RsAsqaFNyIipT8rd6/JDbrJle2QWhC+KacBiHv9jpIQ7CP
YEMgYJisAPwYHty3S6/Yy/qC4+Dpu+ZZ/edNmb+HNlKACnqfetUlHBl89vKEfiYv
gm9iXdrUecp4CFVUmzbK9SVWKA0OG4jWPFNNpxmt4TPEU9gzK0JkhnFtc5tHTnGl
L+cV/1SpcJmtST98jjYYQk5CqygUlRkFXXbUXS4M/Nd9X/b8sBEaLeblBG6OgDbZ
myrTJ3ce1RwMYNDZ1XBa4Th5UdPHOHinfSU8ETsPhWv6Rns/8SBw34VY7qP/qX9/
Ivvx+lbDg2SU/tJBs60OF/Hsx7rHbXiodTAZ1fWSE6jpUrecGwpuX8rdfgC0sE9d
P5oW8cIdluGLuro3zq+1QmbwTPmvoYKcu9q+4YGDopIbwr0Bm3vZtRngBpvdAGdc
9g1oxPs/XyJUsU7DG3Nera+sYFG6WA1EXTe4gGsM0SQI3zy5VpZxZdWtvoME1EXA
ugT3uKuowcsQEGpZC2gzDIShigSw8Dj+xh5JaI0G7RA7jTFIL1Gy1Kagn9vxgE9q
EwM7ioZ5LfCn4RNSbJNoZGxwYo1UMekDrXFchpBmPGDEKYMnrEpFPdgt+pT1g3K8
g671UYxh2bZZ51z7JHQrtmPV7HV7kd0yyiXvErT6s4kLAIjBh8Qo4n3bi1faWFmj
YZIQr3v9fwskOKkznkJF/9ytqrQYSRpp633Truolwq3OzRxJ3sf5lpk1HpFUg79j
N/UI815U5HG2D/niQjUZYLUCD6N5oJtzEdYazRi6u/8ztJMorG0OCKxVHAF2++Hj
8aqMWzY70T2so+Vl2qNm4ckZKBNda9BrIBHXK6+wrj2x/H1V3im5QMomXySrWlAR
ukWuk/2q+ygWW8/beCPlcThy6Qpbxl2FQqnJLrUYNzQREoEN9/klOBPVWXfESv7q
HaqKKbcPw221LU6y+zQd8ynsPVkObHfd8Silu/FcWloP9qvxii5xoqzycqH/PIG5
fKiRC4IRFsQddbXVariblndS6V4QrwAOmKXpu5oU9NncFsEn9Nn7KPWfdINmGDA2
GEE50maGOZkpHOV69FjPawW0ozsKCe8AsKFoUZkemXIVTHxToz6v0OU6TOqvubw2
7c5rOPQ+nYEceeZnI4trzzCIaGFrOB9lxvliz0cdJU4uwzZUYKe7XZqZrJfzdgPi
PK7PX/jJe3kMuBoGqMtgWEhfUmFabK/X8FuL3BMF2UPR9Bz5Ew5fdnWgLIAIEGDQ
DR8vV+nMYHe+fD9GAS4ao0qIoSWTWYjpIXgLU4DOg2M9+n/53RdE4JRIKMYd/vDs
cFAAEQGi3dNgDBevuLax6W2eil+2d0LC0QEbsfY3Q9hnDmsWBlSBh7znw57WkmTY
cebheUhel7BY1PrCsJa/83obfj+GgP+3E5cbkguCKOh5PjkPUmZF/eYY/KXQ6IZR
zCIKTp+XRaGvHPvMPjaHPOgYZbRgm5J50rWZ7YWJT8lgAhNpayJoYE7ceKIKDB41
jMbRoBENFdawWoTUZeY9XWzcVksePl0ekA+qlBXIvFwJWCMb2ZpVRV0MqnztVzD2
MX6ZeWX+M1xCmu3Y41yDQqPeHNEE6ObuylWYWhMMt9ObBUFrwVIOv444WqyAAA7I
eE7G6No7mIeWHKDe8BN8K59o97TiUFWlLZuYKQF/jEo9QzAjFcdlWRO4CAjUIeFG
DYjLmO/SrtLct0wPX88k7+WTDgv/X/Ki9+Nit29vtCbQxvBjp8j7l5CZDFodu6vS
0aiJ2dNl+BYn62UVXdQPVBG0unSCpSBear8kL8voDd9aLK08nQmK9CYLfEqHX9nM
+ZOp1NSInvBsLGE8nGJSw4jexZ7yd3iBLQ6etQ0yNKeRE4IRHIP4mV/PRWN4pyzX
uQY7DyNJalV9RZhVm3xZfJyHwJsmGsWSEhGSbaZ4wShbylA2XWBDnsvan2P63XCF
Ri9/aAWyYuJdowByPE3yP7mj1y6DP9kAPv77F9NYIAzJ5GJk2XaqqbLQvKdowqUe
YPX7peDydyHUxudf214NzNTKvkizFh2szypHKkXSU1PEztbA9iBkquMvLCBx4Esm
Z/UD1eHjWdrRhF8x3UcNsVdkJ3X81ZV4WT2Ig3Ifd9PphlsGB8uASaa/w+KEWvnE
UsNR7P4GKmCR2KRw5bCQeIXAbvmPbSnQDj5UgeeteaYf157qFzo2SFVXWQbPxcT4
VxcycwL3k6nGspaLWUX8N8Sbn5LxMflXGfnn2OyE+qfLLALaiv/CcVSJn5d0SYAI
oEirS/Xr2VFH78092wZVFtEPh/TqqBMvnq+wF5DwgbPHXeJxC01t+UUwsZ3Jf2Ib
tYEaBnSWdZAzb5vkgUGzKLz+WyO8YmcALtONidu3Z/NxxN6TDJlplXM/kbcYYiyM
8OX2Enhgl9LeVSvXlABNabG/a2KMkN+AkOP8Gvzmtd4n8U70fqWOw2OqSmwY3LtW
0RpLiQYbtqFvXQZWNAyKwtOxBJrPCDwqYVxLXIGL8qEBDhXy+RYNRlXlscJi367a
VIBIAbGMe66yyDno3bPh3qu0HDCM2UnLuGc7dSTRinzUnYOLHs9kzMj07wA8IgaH
sbtoRhxLxwez9LEUlG3S2EOurKBB/NpwCRWHImY216DtDJxWPP3Z2tpzA7cD6QYO
jDCukz4f5Ta0xcDObnfPNAdRFyUwQcpAwJOepdb8Hwdh1pUJxSYq0Jdw5hyUfKj4
ns9o7nGrGBbBr7M/NBFvysAEmVg/SFtbujIH/PBLXM9jZ598e+IP0TYHK3WoFemg
KtJxVeMZccjHBLY/jS2gTP29smT1h9C3Gi+2yZnlGUAdmDtag87Nz7lGzR4bL7b1
d4pi1d0yzy80ZECbSS9DV09cvCM4fjvBNSyQlsoabbs0mKNiKrwCGOPLlXH2QIO2
EMZsJWm/sw+sZm9HKptAHhGf00IxHggRaE2JDblNYwojZl15jQdJgAx6mCVjzjUZ
MRZLpyQOOIDL+1zqE75/CsviAjbWz5WumQc0ZG2ZKKeYwIVIkh+U1hbjaK1lMe/V
JZU5MXFDyZbFvnwhvhtIy+oQqboOs8NQ36cIiopbla1yW57AuR7PbPMwlHdnZSTQ
alCRd7r/nWzhYv707yiYtDAMeXAUcVlSrMqs9UsaDTnpmvOMD0FsssGr3wul8HDe
/Cx9Mf2xmQpF8PeNqnEhVmc5i6Vj1VQup6UgOm3jyew2RdmusHloaB5d+8gmm+f3
0otQjuN6oBVNyw7M6ZGzmwlBp69oln+EQ53WUm8MNbWDZ/WjlKNxlrKGHuL+40f3
PqDXMaNmLkWdy1Bb8NsvRZsZpqOSRGzrPzvpa84J3N1FXAC/ZpbnDryug5mmxyD+
ymjLY1XzIUKAyxYz/5+bhhkGH6z2XR0YxoWp8/huvmoA6xJfQmMsJQfk5pMx/LDk
lkGImXf6rwhdo/M3iZHGH8lvqMuCbFEd4xJx1pTv7vcNApJAIwuXZo+axHC7bDfa
uHFWuY2FP5hSYulHKLyoSp4hqTe4HR5RGbb4LHC9meMdKoWBErZ9n9XoHCEMn+BI
5nv0P0lDKwWBA3ysGELUb8FcxsW7q51KJ4KWxa2e2x+FurAZ4LupoLoxVfNABJjU
kwr4ZgL9C98EHSflK/C6E8VwHtEvWo6+SABQ79r5RbKvxqLzXN0u6qNrYEA3tX+G
03Ih+QyXOaSqB182A7AHiw==
`protect END_PROTECTED
