`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7c8YqktjHKnMWXbmuzk2BWmVTCpTHrYqzR8hcSwGCCVs3fcyWIRF9JVJPvjtvNF9
4oRmAAf+1u6QUi8SyQXBeYVkajuf3aB5vYEHsRW32jaoJCIXvhYIq9nqz8et7eTA
ZPSg+gpI7E0MR6LBqzZyOWEkykZIobvjuQtC93eIX2urt1Okqh5dKZZ9P+0yI4g9
GHk0Xnfxgw/yz9rJ4QxpDbR/Zhl7dI94l4JdJUB09yl/oMfLXqo7JGges29HgzsT
s4nsqBL8BVh6aPQ+M8OoO9tswkDgmrF+OP5JvfOdPNdFZdLuo+BFj9uzVGZs8Uhw
y/fNUf3qGEq8DoI5+/nDpjhjDnwKbzxWLVIXi4IbWoxZJLBqcbEmy5vPl32+oEpU
vGEzOr6HelOxOunS4PDvw78kBuHubhn20q5XgbadOIOhBUcntfyjadeeJRj+Vs0X
7fM0Us8Jzph5r/AvCd+NqxbGOGE6EJ2X4ORcowLesjbTOohOXKMD8F9Hh6sVMmj8
VsXkIwKRkEsUpX9F6tJThEhThhqyCN7oIdwVfZQ3j+vpmrouLnMVPy0FqZl6loM1
wsGEeL9qOTuuha2nTtFY+12rXmfTAiy56kmj/65bUPILf0Nq31DCYYG/092PP4Nn
oqnOwfdzhsgRRs04NOO9NPKErmrTYMWTLP5oLPDgpRxzcQP+gHKrYqvRSFEK4yJg
QNuHrixhacjgoXTaq0Xm3a/rRy3FlH7SL1Oy5/i+mWgW0fe1nt6koFE3hpthEHW2
0n5LMikVb9hJfk+4nUVEDR1os86TvSisU07omLF9SiuWQL72A2aV8J28bMx4OM7T
DtEVEMKg/vB0GGaqLdYQONxTAoE8ssDZLnRj8mDflkDBhgyK5SM6yPBl+PGeBybe
J3xED0BJKQkLNpOVzHtWCHZCF3HQguUnjqhCgq8pPOJsmVEczQiCKKyREPMucLrN
cvAY+VfcH7ypDOacdtGx+aoFr0YoupP2+M1cGEGLh/H77x5CX0aP4YhSFAsRETsE
VWJZnuS4EdsPBkt4fohYm7gmdod6zV9/VKMtBDaQ2zLcZ+PuTiiMZOsMBJVK729z
ZE1UkcJSa4aa5jpAMSX+EGt2iQvw65L2gidbcqg1FPexe7TCxayaxQohCSU6v6ue
pPUL3rqSmVs7YQoiOkCcDaQtTJjBUxovTmB8CmIRNFxuV/H6SWCyI+Xx8swoBIbd
jVwSpg/aqog0EumeI+ggtBEapih7DY/JinD7ru8ClXCXDuWCQGRL0QxH1hi1t+LS
CpO+KYNE6WJbG41HrNbqGbTNiayXryjWB57n/vF63WuiZn1Mxukm62zyHbw0uhtc
Mk6HcXQfK/f7W0x7W+Vi5r9N80sCHA/XnEm8Czpv8g37Ih8hGDgEDnMBO8E6tUN/
LltCM5u/xXyy5ALHgocSH1vnIwc7t7ECX2eWURi/yVkzcNfkNISWGt6f8hlSddg4
dbtLbWSi/I3MNDXIUXguJDd59JbnKbYBOsnk9XUGukDYzaUvih/NXDOotd67gJ0Q
NNJV5BhQJ5dbG6DWn75Z5B81dauCNzXy/yA0v/bP23XcfSSmQwjeVAsnwXkFOW4p
5ujjbPUtgEgcL0lhDWbL9ebDchadxJnmgtgNV/iwQXJJ9NJ8LDZaSFnkhl1nOZh7
SuVQ6e9fu8L6xHLnjHrMcWggI3SKdTOB04g2lfVuLcmj61Z1Sz4qZ/sUYgViesov
VuJMHVYiSdylDmMLoNNEWglN1beXl6Xlyh32FAVlhGMVb/7JDZb36Lucj4nTVcGp
fQ/h/sZdI56cQ0Caz0Nhadbuk5AmhdMKUrByDt6G9hOMGu6BtYX0ayDU76q9uSE4
4569+vndAWa/RnwsL3RXOUi1h+EbycpGyFup9xZD7WYJzrFmPoDy+Z+8YTN2uOaG
cER4ozqNFU1QXLBIEsXx5zuhMKNYUvrwN9+PO+dLRq6NmOo43A2UkQ9Zi/7FBsIW
FC3AEdGmrZM+zhADXR55baitF0LMYe3R66lglkLu1qs3+1gBuylPaTsQzJ4i0zbT
in3MvsNTVP/h2C8WIPEY3COt4P+ASGyNXuuniO2mors0w9U/2vjcfNvWEnM1qH3f
MRgN9UtBoEDRgrmdjj+rFrEYnnrRsXXDbXvpHsp4rjYPwLQAy5iOuGSsyDnwjroP
V7Bzxm094AsVlmrU6f3IujKEdk+B3q1zmgUyvZ6odL6SZjxvNQ0g9GgSZDfFuqxT
okDooFEMBSUu957GXLAojePnMSNaxqifp6qj9UfyFO/i0fHPk9RJO09nAcloy3Zw
osrBfU9UBKkDX42tI6frWqpF3akohFgv9XrdnhEzr+WKMBj/KX/0QsFUtlQrSjO4
MFZFPtw2awOpNghNGIOB/41vcoCfrAOIKrxnri4/36QuSrfE4+wMKdiD83cmNZXS
6m3XUut+xVaovILsJuEKCYNhul9bSzT/P0Hudn/3QH8grIwmoOh68cln+5esD+6g
shJRwrH+OA5NM46VCfWprA==
`protect END_PROTECTED
