`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
R5WhxFGBzpTQzOEo7rlBcZUCb3okZfIohC3/+fv66e+88j6Lo/+0JzPIdJ/RDIXo
eR3rjMAm82GhVkXpjIz60FzSGPcQ0GYPFt63qjIHKBZX+pHqy7Eycn3k39+SCSmi
ulyGWNDaATVKW3dzbwA1Mm9/bOKZO34thGbEzmoiZZhJJW3oe8i0QM1a1Y3KFCBn
4QyWKDekTkg68R8KtOO9FBv2OiL2Pe57ruD4yb20uVlSWEAOt16OZAswBwXVH9Ue
KMFjM/s7E+OBMABGQKR4BI9WA2j5lXO3r1AqZfGB3Jl7xu4rHOJwXKtNuwcVb9r2
RhaGhlbzOTk5SqfYXIbJd6cetR4Lq/CXawHCZrv49i9PvxaifGOjNZKUqlnXkbFi
FfxhUnywFUI3/VwZ2ePh6zSqImY7YIAnOdLFvsZWENy+hnJ7e7aR6Sn3FMVL2TR3
a6jw46193vOnPr5QcilFjg==
`protect END_PROTECTED
