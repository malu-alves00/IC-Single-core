`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hpmp0OqshaXSNqXFNS805DOgujvRrXvshf0at4KzCAeoyEFpNTBTW1S2VSfZ+e+I
9ULuopEHNAduIjibq7ZbalNEVvjyQCyuAHqpsQfPkFfMQzeDB4SJnJAMALKSnJxh
Yhu3xg4UQM56nUOCGjJbrHmKVFC1iw61xo4oVUbL9OegCfzj+zrYiuKqmPID/Hyp
ig4LQBYd8Xp15kNGLQK9GM1ivLzEZA1Bt6SeiGYbiPPBDqPhRkwg6fvmoxfEA1C7
QVEskS9XDcAMTXw5QQCjUAWYeJXC1wc3KeOUtl/HDUyJGaS/6W3GCqzREd0Xcixc
o/i2dx5YllQPurWt2nOalcM5s//t1fSFN0IGoDZ8IDeCj/Jx5dIEA1nHNsJqX7qQ
mxZNXvXfuYluFoZdWF0ahU3Zhf39Oma880a+ixhFqcEMmtveBN9BIZpP9Ey8jqQQ
kjOHenEl81dD4xmhRYNZ0VpN/iG5RTfopF1UiZ+GP0GdnYuki4AplQIIpQaRHB+m
4TJAtKZjYok306vbCf89/dIjy8Ouq/l3nWPY+0Xymu2Dsd276BlqiS3lQBKZNDa5
6sm6vo6j3DERDGoKq138x/JdcxA1nmbAeJbww5ONl8Ms5Dcp4PYnJ1DLUwwdVfv4
tTYNTf+jkG4dnb5MZdFB0hfhK8RIpvrPmxzA7m4JzX6ROvCHGMDDCuNRJO06p+TA
VYNg6+kKVODz8d1vbY2nVAmeLKJ6YER5ldWTgGioT1lq0Hvrft00/ux4ueH6rak7
T2q5lBIaU5oPCFUowYSkIWYeMlCySWuhFpjOhsi8CpOGsOC8TXR+9DVzBcLeyefs
dyc/QG+9BhqbNkPMDW3l6g+4AK05Vtp3Bg6M2b4h4L+TIhzu9xerj5GEXVmv+rtV
z7YEoE7trsjKjtO1ofeT7fIgsZmU204M++H/EPmR4DQDPoqi5TFNVn7Uxlrd7lEV
JkQ340BYUvzv41Jd32Zv+lb4Q2h3BhXw2HhIGOB+PI1SVrAvvucoH17qu410xFe3
f67UhRec1bqlWdQdoiIhJMgsvq4oj9AdN9LkfVJpBsg1/LSOQlN9BYIZjHOnljm9
9fFxgLx/Tzm0FWJKEdIv3avT1ktnrRkCwsRtoTTY/glcPRkdMn/TNLc5cLuccyYo
we4THC97HDL09cbAhMAa4d7LE+WkjTxMbM56XDi6AdFpuFuYEF7jyUMucfoWnVPq
r0yeLmeKgDF4KMrf2tP1edbZLGHxLO3EyGSWTQeMCRquMZoDbI2AEUCsHrM0tVzF
TafFIwxcJVEusfYTF88wrsYNGme5g8byMNIaqhAbiKoDrjCLNWJWCCLlZJFt4V13
pIk+guE8ORG4cGgZyGuolV2ggBx0RKfifwghfWNYl8fVjZGWvXElKOpMi8v1pFKb
P4dRk48iOy6S318IfA+Nzn7o9GoTWZZ+00Kh7BQDRCu8JTm994UPxJDrSZS81No3
w1T4W1y2KJN8hxAXszKMmUmtmFQ3BQBon+VUAw+RwdkbfvyB66XtUVIZS1GbvjVp
JfGO2PZgSbS0gpzG6NYW6CTPHfCykU7AEMzKNNeFRwv0rrUna7CvlD7Rzfe14XVD
F0vezYfNNVsfpqi+rNyiV5A9Mys5gWrgogeTMgG72yFGlegnwLZo+X++h4ceSmht
fRZCykOFARuqQNxp/g4IPflcWk95ZTsh1m65+B4F0Sg+Bw1DcZpegITfcpWXq3oT
FYX8ek3rJpnay0wVv4/aTvkeq9tDPIYRRb6KAGS2BGQ7n5ZZFNvRMUAlZa7F6joB
auje5fQm7na7thfjSvDuNyOvEMYsnzo/704h7Gcyo4uoQJJS3gPNmB4KBhhvug1l
oPN43Cm4S1bvT7MV/DnxrifG/YZEfcF/8aAkR+fuHNC2KopZ/eyW9cugIq8YYLMz
yo7XC4m0Kjls70R2QtPT56WYvxA4CBc5JnDRrnDZn5NsygiclRGt9Vf5n+uvtEQp
uXOT3g+kUCZd9CoiotsFCwEskD7nXSNwZ5q1EESioe6DpHPLB3zRbBwgBn2XJ506
b44ZGMlrwNjsMWnXpgHuYiu7cQK4DbkPoLaFmzwWCs0p/AGvwrIoKHYELseOhfVs
RYl58EeZQQzvU+zWsUcSnGj+GxLz1Pz0DntOGNEhN72Bn53AfHL/DkCl1UWyjeJ0
t6ZOzoF9BRZPd3QJebYvKlrW+Edl5yswGSUQnhhv/Iol2aNwSCdf2wQyqfPBqaRb
RXZNbmJayAB3e/zcaBRLN8CRqLeNHpyGGgF5MM+wVDF1Tj9O5+nicjhn6zIv0/vp
rvJK5d2JY0C5P0xzuMNXvlS64tZLRZ0whLJU5w1Xkl72mRSmqjgcL8AUkgrcXnyx
333kv1O4jUKH24lFF75sx/YT+6q+6ymsk1Vz6eIvKE+fUyZkCsFN7Q8HSAntT2Mk
4hgstWexdre8vlBGY7UusJWOsBmk+J4esJMJx6szB1UQAnO1NNJl+r+euT+kqWa1
zEYJ82g0zwOi9HE1Khzs3itfbuUfo5AbR2IZIOanimP3GRT1Sw+LhtS8cmwGo1sC
083Lyk6Jb9BCIjDGWAShtYdWFU390BNXU7+09qsRNKfCKzW68mSgZplmm2L0EPLN
0G3U/MmaznHFaVktAZouzJjIaXvZc7GOnQkS7UySGrbjEJXZr2ZS0Qu28SSx1Szk
hO0bzKL+HgnVePDnSWDYRTZEz4pmHRkkjApP3X+oCYY3EyTwNKcDgpf5RtBFqgld
IRpuXEqOdEJxyHHCnEhqzpQqFmH4K7/0dZ2AVYYu9f52X/3jEUQS+yLlDlKBfsx2
uU0sODEpHHUlJbezI9G0VVXZsU8qmmvwOXp+S1715I+GlFX+xuO8U2g//woPYKGE
x5JAhkvCzGRpCf9rvaxf1s7NR5Qt2x2SV8oYKZklmIfFUe7uaaJOTb7ySDZD812V
4TfjJT4hjUChZ1BS+7Q0n1J8yIiLryGO3IjsptGhMNDi9qtvlff3HVj2+6G5Jhvg
sIN45j36N5jvriZbeJ7maZSnFQnKORnH3O/7W55JlIYMrGMrBdERrLpblNPR/gFp
nBODFjPzlryBkHKg+dJHnlQPKDDVZUDn3RqmeIpL8y4qHMiNyL5/IurI+fUfVUis
axG+qCB4jM7HrK8coBkEg5r1gnnlbkVWPaQyYI4PmYgZh8PmGCWRGyhlD1HWYsPo
2FOEspa4HY8PtMMqi+3E5jSEq7Zb4LMiZ3VIN1mHdiAv5z+lXopY56HXNmZ8olPM
YE5aIPzVYOZwrBTu1QHQljLrwlu4u2ufo3guwvQz6GT6kHED8PfFyT8DRFVVpr/T
/qOM54BkC+R8/hbnoz4QPRLvPrP+F8xm+7vZLsMts5mgVSWvCSoVnTj18iXJNV2I
I/iBVXAnE4us4MTEMpywDuGCTZr4G0VjHzrIw3Nv0p4g/lkdNCEszR0GpE57JG/w
A/b9k5MQB5sBfGsmYKPM0ClP1RmA9cc2ShihnnhA/rDsBRZtjLeulrtQe3eUXrCD
JfaJB20aCvlfecgnwaqFsoFem2ovQjsjM3bbacQ0NRVg1f5dI+ZuMXspljt8TMWB
7Xy5NavD4nZL3WOUBayWFl1gyZqCgVWsOMTru3SPN8x4GFhVrwif8yxhArC2Oxf7
jWtiGqYMFVoqaF9uOu9SUuhrRZgqcvFIU6Nqs7rgmhJU4Xlaa4qc33T5fy8wj5ka
sUax8T8kduKzV8dJh86GDS+SjVCLc+hBqyKnOIKPsPq9KumoT4+gGRHFGLfFsN0I
yFlWl6C4/ZOYvd4+izUCjzAGJFk4ZFG82POZI1AysKB2+XUx+6k4I6sj9YmkAi0X
BS1sRgb+8ki54rz9VQsdnTQ+mOthFLOz1cMS5PXdYsXoRqwAsLfvxtTipMTaRK7T
D0FlsapUavi9ZU9NP/eHxXn4aiZvCPneMg9UkPkZj0ApCCsHgaLr2KoF9KSIXUJW
OaJ5qxywIUZlOnG/aiHycT7kK2z3Lx1zM642jubOgnOZkzv1Yl6PppAZ4+5j3Ny/
eEpz0hwbupsxOFarjfqYkDlzluvCulm7m0XtPPpdE+bOpJTCbilhZ7h2HdssN2AK
QN4aAyXlDAJolVkVPRJ2fgaT2ZdxW4wvLcTWq8TKuGKVlxJY+6V2zHYDGazn8CtR
oyetefDxh8pn/WrzYMwBvSFyr5Ki4CDQRqhKs13ikZ3KtuozhRvAV0RQhg5VCmdy
2zQwEIF6vv7/ub53CFZGKQmnwWrSW+KUAfgh+p0+JCcpr+oIGhhu4o5E6Kwh/Fhw
KoBYpMvIPAjYkBnFcCm581zEQ+90edDmXBq0ea6qf/y0mHD42DZtDFGG2vO3AKzm
LXl6pEMjzE4pVYr2AulJhc0GCyQbuZz3lSpTmCyocHtcKkFo/ZOg8OUra8GAlYSi
0gJmx/4h7Qj4V0nmOBUObLQLihLBW/j9ksLXjE9XdM4mmIumBL7S+6hKUZEFwwFP
r7dR7u9t+UpydvidR707mNe8wiX7pHBwmMhPSk8d9WJ3kqr/9W3WPiH5//HVmQY5
HXrGZuU7ZH11XeI8vnjj4j67BiwkMYbpBypo07r2SIlerMEG6OsXqtbKq7q4Gz64
cZJR/nhbN/2whIdUPMD1PIh1wc98hTgDdqEr3WFmg7Y7iuATQ6OJOEq5V/G06wqR
Dy8iExb0vB9/kLbOg/P1yMJezaJiuZ6p/s01aaqVMwVn4brt0Nh7onrlC7lQERdh
V80hbue63YGQZ7DAMJxt2xB9pHu9V7kKdQfZqa7tnbS7vaFHhTkiRR5wVl7LbixM
0jZPCR3+b7wz4XyFI9/gbR8hnSd2kjSNUW1nPfIJtakfAtLlQfX9lLwDGPSfRv4j
AvbyWopFLHppLYsHzKTM0avgLdEEFMIWLYfUTsdFaD7iVu7MbHOi6pa8zlxUS0yY
ClnOs+H77t7LTfptVkQwxZXZS0X7U1VRLENRRqiYkk0HQB1DNhBFevK60fjLB6x6
evYo4cVmzUR8M2fE8tZZEtnYAUuCVlVbN4/W6Uf8aaArf8LXf0EqaYUhjb19HERo
O58iMGhB48eMAvotm4fngcYMN7OkvOMtTPtqdA07Dz4kGe/Q5j5EY8vRrHRcNH0T
/vvuS97iIOfNeKRfYmZf5So0WEAYUCxkk3/1Zz9B2MuNgsBTcc+K5RsUaisdIynR
C9fAa7ngOHeZ0GiOyuMijqBaM/dQbDa2M+O/Ei7rwVbnHE0DjmL+TJ04fsY447nc
X0Z5wp4sIMTHR5Tkk4s+f8qwJgYYsNWUMBcwidmHy/IKy5neW9SfqSv150thn0Jk
GTyGU+O8UlHRySgRxvrzfu435zYUzAiPviWLQyRgJ2hjboPNYc2LWZz9kN8vJfc+
pE6QfGoyqCdCReL8RQe8y3yogNgh22RMmawkCqOsnJZkuIQC0LYvHlJFsa3/X+BZ
UHeIzbwa8crP7ISZUQjGNdB6nRa3KfP36Z+SoNMIm4dTBNO+sMGu7cQ7k0tJlENw
nSXM1ztH3W6FUdgqM590Rf+Y3v1KThHVF1zI2A32877P0SkpGZonlPLfstPhDjNn
84WgI5XGBKfh8zBH9mhFThPUD6y3t8vXtWur/a/7JGdsoih++soo+B12WPEJ9bHP
jJPljG3EghtXVTIFfWh/8f8ql+v57g6SfwG1AXriOrmWktOgLCecCK3MgwbasME5
QZ7eTEPfebb/CK61YwVoqaxsc+3V26bpl5UoMbPkVOWUNzohdUCcFGVe0Ul+YZaF
iP4RIpLKLE86NZdPaS3ojYX3lWEchtEE95vr93pGg0AwTI7wmaM9TbXknkduY0Zh
HQ7G4Wkxo/wSF27Pp2IiR6BSQ8RMBciSbIFVN7RAzFA4ntYA7NuKLeJ/wFZuAxj8
mBk7VJlpwzbpOpQJgj+3J/NH6AbnWmgZQaE/8eC2svw5pxheMmN9twNScaygs6Pa
8auil6UbEExAYzm/jBebI1o/Zlq8ud/pEKzSBpV+wEjzh/3U98gCpcm6MrssHhxI
k2fcqVDY+CXcM1h2+h2iRAWUFS4wRmk2c8DKvSp3hemGK1h4NAw+ZpPkedn5mIXZ
CbQIXj2SYB0YVcGb3pxAKTTLX8gORWS10X0XOWXX5Y2BjPIkLshJAWvQofAEJqJQ
VP7en8mkI/pqEpEcn4F4Hqxqg/WBvpU6iBxNSx8LtxOLcGlnvpTUMm0KCWb+RNy7
aJRXWjjxWOe8cukY+y/Suk4Ht6CiWvAiE1qS0WLGASVOe3wtOJmsXHx/Viq3XhP8
iJzImJFRCKXdcLPkeYOJvBkFF66dhgad2pXSKlAZt81uZR4tc4nEnLB64jANsRh1
M4kgctvXO/6k8dHGJaBZ4O+1pc68xibsAeMeQCGgiklKz2AokscW6kRyOTCyzweC
nNt+e5XNnKhsV2PfuSzRR4WzFvYe8sM8zAPDh2elHiqRd+BL+PZg3DZWCKHKxec2
1HX00NcW5clEb+cZ1+RtwwxhRiLFM8NNT/u+ZH07UDjJAswyS8kUN5Q0XxrEim4n
a46n3h9fm4648UgvRoD9FXsXiA3lwd4vsIIM6QpwXblIK4PgeXcEskpba2ZMMwEC
NZeN/qWE0ZiMYzD+KsXF/wrpyxqQV9STK1Udc9O/yCc3zkQDWdDrU22WlF/9uDJq
XLM8ILwqcch6Ee1qcokjjPT29OOUHdj13Gm3NDawi4zqjSh7pE5D/WtxwxWFKonr
t9A09YFMuV6VBFdxavCd3YQ9IuHur7hyURzKdj4CxMLyRYzsg27gLxqmDRopUJgJ
2Iw9YiWAbyzBDRP1uL89xqmiLkMBM4g1UbhZAkMGLxRkccmCkWOBthcuiqIhXMsm
1oHCf9/CgUt5NiyAbJP0X+2dHtYwJGyQVe9TFIcJrYrRl8UYr/MhH2LlTmpUkpAq
ydhNtXwZMsKsMExYa3Had5X+M6FPf1IHJ/Pxo8TMBf637OwSdV9aXJ1CtYUgz4RX
rTryHBgsE61y+snvpVVY+wnmtF+sFinazFP0BeYMkwIv241v7VOlwGt83yrypHqz
XzpdhABAiiPk0ppV4OmN8bNBHqCg/Osyly0vn4WBhjHyPvKF9/lAVUo8aF+APVQ9
9fRRZLUNZbYiWHUU4UFN0zpC4n8s/O/mU4KPXb9kV7yvLG2aU7I05JPXoeP+XIdQ
h4Z3RbCJ4lDSdfIbmzQ+3ORjhNXfPEgiWYQ0DP+w/UyxhulNVcOjLC6XxI3X/nae
PmNkKmzlbeEbnoYAwrnrOr9yvp7sqi/9C6V6X/XCmfktSC3f2lWI9pN+6f13JZo6
CNTAGRLbBZqiE0JOyRqFKtQ0+5ExtEsMZnB1JU8KL+eklpd487XNlRoM4OyazGxG
oNjZu46Hrz1B2cAg/VAoOC4scKgARc9JDmZdrwPmJxs33FCs9eZjU94CETZ1Pytz
cYjfK1ly6dxVI3tvrO3nKfDWzlCwhCyaVB970eqqPqwHOYJIuGlTPFbh+XGG1YPN
t8zO/+d7uYWwE2q5z7OluHrOC5QuI3qdQkVuDO7t2iFImw+TR8qAetNwq80HkIh3
Nmv32eF6m1Y82LSkcbrkrJz4i8tUCNZJxjutOBuQIKPLrS5aGCYTeYLqiswzwv2I
8Mg9d+y9Ll/zq0PztbAwbxP+sq9yWGYEVd2D1nZcCeK1SG65Nkl6lQOUVJL7nXqC
GfSvZ5QQkmxs/rfIH3owv+6h+VPZ2VAVNR1SfQNSlG6h4wbaPj79qK0pVQgIodSI
WGRFXd3uMwV+l4UYUwvQ8oh/bOwI5IObWKoOHZi3U/C0EXAm2eHNjb9Mhmsci5Pg
ewoNnS9T5i1sV06AVXP5dWvnPizQAgvtAEn911aMJz0+nJqQ9YE1RQdqL2Sm5UHO
3kjTRteldC0B80ks3HOUz2ax4C8JhldYakCNtil+0k0BK1BMTO6CcKzvtyfn6Sv+
86L/1HkrpjGmAVzYeSIUAXbmV1GFPjWIJGo++vSR4+yE8bUB+nWk9qL7F+06/4ro
jB/KwbWVDKRDsGkvYG7+lR2s8BaroU4XD/BrOV75P+9OYZ7D+4IJs3TL9udZn6c1
uoW6WYTl0Xb3GXTUPqgmdsi1HAwRYZzjUIDdDZOaELegsUDpCHuDg9zkvdd+FlXk
kDBNgT+RB1Mqk0VO9/oCG5Y0SsH5uPBXkNO8Pyqwj8XtSCdcjnTqhAyzi5RCoPKL
ZwxnERUjV53vn1fB1NJQdlZKwa8dJXpgroR22hDQsOHZWeWCb+IzONNcZMEMCAuZ
lpgx3FShX0+fcj8P+haxYaV1hm42Rg+XyTGd75+eFDEmzzbZjlUU+bn8sZyUQo9y
bNN1+A6lLfO34hZ9F03bsI6vExpHuPC+i6NKgQ4HJ4H3JNVDHcJdBTQGWBVEFi5a
e2w7nivnwNRwHvdPozTHj/ULXX2BPFQTDHgmU8pJF5az9fpIeu3ha+K+R15qYDb+
VNuUlPYfbmuBIgGige62Vnoo3Xj6RtHUIOJVtAarJd2chuum6mNGLHZWDrwr4fm/
IQnyET0oSAcDNrJtRwNKTJnUZ5BxHpENIhpig1LyRwcjfyjWF+N4/5x3M/u8Fygj
YFYvZ8g+Zfy+/EiWky8bNtpE+qBLARksR35r1aU+vTdndmQObO+Bz6IzuBSoDfDv
YbKOIbYaC1R1rihw2ThQh216+C+zRJWH16wpwvW45IeEAGCSlfmH/KiFw0HhHoXV
7/OZJPZ6JK4zisUNYHLLstN0T5dqk0gEaX/pq/w9z3KCfSMRFl1RJYfk3teRUd9P
MQ2UeoF728FfXp41nqXLylE0P1AIneegRwcZTBPjAW+5y+BSnPnwbQmbxYGGzza3
QNiWJUNX69uIvQod46ChXKJ8kJWQq98zg+poK+AocI4=
`protect END_PROTECTED
