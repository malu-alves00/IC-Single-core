`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
glCTNXsA6w+6/vPE7ip/S8b4nPNxYGWWJvbGlGzPoU7R47hXcq07W8Ixma/vEach
qDb1dwnYblt5nT/7mniWWeUiNQXV36j+fn0vsXmPZlbLALUUMZ4FrbBW5PiFZaQ1
EbupcBNNhGrRqKGmqJfvJdO+Y/9BQW/Qm6k4jjaoXxlzseDgkbjHkExtc4nthsqa
2thL2QHjSKhjOxSay/w8sYMhTBTmhs5vCBNEGNJjILFl7ZRc+qr35i8YNEDTBSqj
V+DeA2WVhxjbUt0OB0d5z2u3TgTXPBOv/U9xLFIcilXG0AUAM0ASnw53cn+veNOa
31aDw3zbQ7wnFm/J5SxJM0tP5EASoaREU1rSACy7xVniQmm+Bxx4kDYKJFvk6BSP
C53pW+9ahe7MzqxwPE8UVSz6Vlw+oo3OEArVRUo+i/hEFDTSFydwYcU0ziS4MYc4
ybzlKMYnxCNHeM8Ug4Vm+6Gp8tHUb42ikam6Vq99SKA=
`protect END_PROTECTED
