`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
P2q71evRcamBlbnk0AOgpYc4C1q6cytyDiv5M4U9bOQEuI+nKSVvt5Z9SmkfBPQz
mKSatUrgBYFCJBkjPi3/mp5Q3C+bDrEzNc4oi9Njmr57YcnhCTeN9HJ/fXRUO6QP
ln21wAr/VOy/RLV5opYGt1HpqznQrhBJ/6c7qfO5YDl5UU3UGJI09NqweqP22Uhg
Q1hifGn/W59l2a7m/3snTIWah9zTkwuaBQJJrVj6C8e0WqTPhugzJO78zui9EBSM
Oe3YRCNWkmLVX0ExKCPGWHFswAjeLOWX9jtLY6iIFb5dTwl47UAFLkplxpOKTVWt
Zd0uKxSYYUaEWUdL5+sgizld2Z0HlPeOnBWJWUiAppUhrIRiJSKu84yeqLOhKfj/
BN7Km3pdHPJvGmIo218BazfZZo7VAxv/Klp1bLPy/xceiUZnIOjOfDl+qjkJgkik
p823FzMQ4psAFrUt9TKUYBWbnmbsJfSvfz3F3CNq8dUFZ6OlwTkkfX8DEKNgfOOz
mps4ZlMdSkn6F/7oX64joGqjSvOY/k/d92uDRbz6C7HRr3Lb0k/4ffYH0jT5t8nH
ThMWk08cwX7LhAg5CB6GGMArUWtT2WMhnXtpwqFuCtfoLUb+t9NNCH02gLZjWNzA
ejW1g+ibD3WoR/Vws+Feze68aP8UiYWL1z9zo36Q07rLHNUMJJ2AXmPmi2ufBbm5
NnCIgaT7gLxNQPMVg4+qoyJZtloHu9q8SkajMYnp50luJUgM2UajUN+L/xsGW+Ax
TdfPAVxkQznl72FL451OIwjNAdcD/IhNl2TnaCtLgjpSOFj81gd7IoCyIpkKL5OV
J6KvoEmnSEhtvz02brZORFt24rcGsTB+5hmhDO/hGoxBLO965bAMs9/51tfqP7Oc
MJGiurdszMISB5v90+77HYKWPkd6/TXqJeVVtuvHvzAwmXl7Xc5cvzokqlk1GaKf
tkoHGysmZC7F634d5L9a3eqNWAO9CKnFz5bji3yTjLfwHIArg//+XzWugAm2ES46
n4nQyMlmG3Eej5pc1OAeU1m3TpSDFDpbB0KkfkeZ1WNRDRyGXO+T8EfhzoJN42C9
Ak5QPSjYfkgjgoWLEW3T8SoSuApO1qm1alsvHcFRFX/hxoIPvBlAY4iE3eVAElno
ylVaT8mw8vn503vcZ4UViiMiSvp8L1YqDChF9Zmhekn85j+ZiQunPerFClpe8tbw
VrXrLax9iOPlP9jQTzjbVuTKHd0USGTgl6l6P5+bSYagUJgbVwhydDUwfv9E5ZRJ
xhmYpyVVVjySlG0ZAcEpllf0yRj1NDx0Itfk4ykn936y4NUoOnHpG7knqXgL2Z/q
kKPUgm/Jl/wF7lTkVOeWYZIvXWGeUFWdxlGpG6cQhwiejwxQpKUU04J43KP4X+f1
Hnpk4N33Fu8aE258JX12edbr4feA+GzBmt+Xp8TQbhzJoW4N4ZBUOxhvEjnQ4wsi
wLXNrRwvMpKCIRw5U7+slYEahwEjXElTXe+0Bd/23fyOOxj1ZqM6Qet3vey1Yn1l
vTCdxqKtH6D4qtSnLYnrsw==
`protect END_PROTECTED
