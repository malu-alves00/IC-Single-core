`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
krngDw+1RN1ZCy3VBjATX7MlQkPvjaL3ie5rjxn7SdENVrMisapJBr6zXcCH28Sk
nqLf75h3+nBtPsC1karujB1iW4P8D9+oUSbFYUPUGpZhHTnLT1ie5wCLOC1lL8zK
80PSh698QSoqKV9Us7iItH3EFD99ganXBJ0pJJjAn2YPrZ17AFD3a/WziP80Uv0H
cDsSyzj7HlanNJQYrU91BugHAbXKFQaDn3TOI2UXrBuMice5jSQtL7Ipj/73V4wu
G836kCby8Exzsa6lIreeIpPjnL2UQJTR5W7fCx0Lu/rp+e72Pj9GVXiqXWECMyqP
RiGSeRxvgsY6E8iL683DMR8QtgFW/TEaXdGhw+RF32feoOPozFoJh9VKcMZ+JTHD
ysrSVDZjHN2317zGo3VuEmT3x+Y4JpxQF/GAhUBah2gfPOUTSkrc1iFil74LXxGh
nSFvaDw7QzwBV7KvveBB1TwsKtKhbDcpBkHHoPWGCTyubTOMI1NYCrR0rb2PhG8Q
lpzp9GVH/dBL6VlByr/F0wxEGfx5Bwyr/1CXrAgIBD3LU9og1HP9aAou8zYlNf3W
TOgLez9gHlprvzQxgx9a3Nm8M8ax+hAlniG/Z0ZSZbSO6J2XXap+KbtnjcTDD3vO
TvmASdjAP/wRdYQmCewmuMHU3+a/Gb8tHqdvuBy8Q7PRe29ZVJXVUMgaodnIxCyg
KH59+Di7wTV38Pvf47KlrWGsNl7ipFfbeOp6LMpcKxTe87u+/zbPvlLsk6asFjn1
qo+a2/xA+IrnEOTMRGwZgTQVaONAWcIcGF5yQJ5wCDXgJptAMr3wl30fYUDt7wLP
oIKlrAOcBMkx1zuduImJH5mvyhKq9J7HZe2sIovvSeBDMzTQGdVh+Q8b6YswG+3D
Yz91dXR8bv8LEea9753078QBN2QxKNM1Qx2uVih/HQGR9EJywW/0yHBZuEjOcH+E
G3Y/Y9HN23SnaS4uIq2dylaBkIN8I2ORaRwqg52Dvkeb3JaKflHQ+3cxEl/6/Rqd
ECXtwRiEmk3EMgVh2qaZIE13q72lHUzl2YdhVPiqafejp1M2gqwp9nwfuyrtU3FG
o5DNXWIXtJeCdfw5rKZbLOJqMKr4I4lMS7tCt84W+aM=
`protect END_PROTECTED
