`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Qh9ifuqQZB0LQ+U0QtMyZ4HYSedfAuGhXwSM3UEcJpqYkcAwVnSmws/8QysW4b4S
mQAN6hIJb/8DVgDrd+RpfiA/GC+ktqfko+UGrzdKQpU5s1LCi275e1fuTlV+BDe6
Ngp2IB9CrmTm4vbLOtjAPzHokFN38DZG2zAkOB48O4bcC4vDjWwOJS/gibOZO8Qp
xfC+M7BtelvI6drJ2qt2oJzT4W/717QPFX8Iq7PxLJmtvZYCcIfuFBQUf1wMrzwK
nfHT75xje84gxvDA9Z8TgmCktnkjOgcSlKnx9gPbYnRbsZVtTqRqHO78DSZNJUVO
m5dDwreMn1T/vA2KvMOFXmCO6QXRZoSmLEvKS8v3JIJaq0iGZlVaJjGNnQrfsG8o
vizjbNnym3PlNkcg4NBy5xL8pHtd0D5Cc1C6jHGNu/N1mxaZ1mH4RYr8QEZsr7o0
AGXz/h6m4OofctoIoYmOg8y6c4bv9S/4NTfpAg4gG0E=
`protect END_PROTECTED
