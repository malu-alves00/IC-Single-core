`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Km4I92hnOawLYr+NqSwmFEnAV2cla6LxyKxKuwy1CJknw5m49p8oqopI8YhpfA36
C+M5AGd530BRfF+ZyS/ls/7VqxFCpTp/mWmUOfXHyvwhH109cu+MG4jtgowTuKds
ivZE5m9T9y5dth1f/GiQv4ERpLZRNRlYF3jgK8ajWGcbJghHz7kr+jWbcoeD2Rci
CTxz4sOhuLmjPGusDMuxnIwZfLBSf1/iMBAHZSpXpSPRt9XyoBqAgwQe/22Cx1VY
vHrMXgPVrkFphtbJGJ8DLc8V227byOat/gFNMKacDVT+uk7TC/eO35+AQbiPs74E
X5vJGlniKlBcbE+VHP+df6w4c1qSnTEYxVgvsNFni8lqJ2X6M5ypC0itHIE+HB2P
gMY5Ss3XroLxg03DD32KAxjV/v4KmADfsT6c1otmR5YPxOZ7eaCgD1QyXi7MEYtO
ovXqy/+iWl5Q1hAZwUJU1eQJwWhKwrcL0IzYxpuerlKFI/Y7hpdfmGimgdLNdEJr
Cvo3E1Axmslbv1wsOKxYgnzjVdUvucT1FF/E/arFyuEie4y+HoS2v0NTDNwVsjyH
QM2KGvpSDbz+EG5Rrv6ZMVB9XqjcIe0bFhBgn8IiuujP3IkYVTQIUSe0kdtw36ol
N+e7CPOn67BMB6lL+HTQViXz1JHM5gcfJxvWwidpHXfL+96Ghrs5iejiDcDZ3BAx
fIpQribVLLuk8NRT4a95TytWDQOOvYYIM3QUgDIGG96CirUsVjUMIQw7w6oIUC+8
3J/xBXXnYMN1xNdVpC+vO+LdOlFY8cNYTYAo5QQo9dsMXeEPX/KJBHc2CrDWOsKD
oAm82E6ZS7aw8b8rowMTwiGKS9VeE9tZhjUVFXNoNz4K55h0KiusBH3xA43aQ5c4
WmDLyUsyZv86h3zXtzTbbOTUXaqjAX3OOmMKToSpbpuAFMM7ZAgxJhh984HPltBT
NPFIxFHOjCtuTBqHMvHyjLrrcXcY2tRZ6d5CP5YehzM5YZaXphJ0Oge6OZEavJdv
95py5MiSZV9wneBt+DHgRSZGkHDjPx+/z00qXKR3tXdYJ3/85UHZssoMubfnWTUO
zF4j0E1C17jRc5zDq5UJsf0hQK1P2/RLSNG3aOZ/q0GQkOAzrin7kSfF+acNK6HM
cJOEkkkJXI8WlZG3ttsXjy/GEMjqM6nQ6c043z83vF4re3d/bR5bZxioUdUbc1AF
c3Re4++r1n1foJGoDCguzMgqkrq5v3+o56cgjA43Blm2ZVwkNMzseUDUgfNSMdEv
OC0uwItFW1WVaf6dJOUdxYBgAZnl/OGX+A2TcXozQ2zEcaifYgKw+g37lxEhPM1y
SpI7W1C6nlp97CVXucAX2lDGG3P8DMBUNGClB/XwqNNC8C4KDDQ20PBYwFu6x5SS
PGeGmJ2WQbGPUJ5xuGHONdDZphCgf7tk2CF8lSjlTW8x2+fSkZJicMzwSEaxF7K5
84/BYYHxhZq3WOhKH2Zr1Biw5SjzHHkbxBe2HtAk36Akl3KMjUwqAxsGG+iqLHa1
88wETm5lsRP4IlfoE9f13VZ/VxIhmMS4G81QuoHlb8JOZ0xKmoECpC6fOqT1lrQg
hPGAYnPUlNZQhAq7zZG1W2gZe3xDZnfqjeuOR95bHynlM+f86SvfBHCyLNDKiZL7
g07/0gtUt4X1DcXsuT8aYqYNarXoF5BLnBxlPBIxcG3uahXf6cfm8sL2PAnn9uUP
YZDjwsEd3cwhQYhV0lOqMu0ts4fqALl1wYpTx6fwH7mm55gMq5yG4ngmWzRmRmU+
lX3BLvQ27jVJvf8bAIzWUyVrGZVTuR2L1f72o08+k2Y4FbqXlzYF8IobAMTVhW4l
nEPUm+E9b/enPjK+FNebQi1sjmM9BZecfHgf07F0dxdeZK5ulsrp/u2tgweELQqz
Hi0GOa7KumVq3dq2IWgQE+osbnhGBZCoFfiCegXrROtaRPYL6YpZfiHefjd2rNJh
xCbq/VZ3jnfisitIm/ALsJcCNeGaBXkITVyWdXLuygs8rSm8hjrCc/8OxWcmgF9s
hfoqSdsvSICVY84C2pS6iKNaDIX1bm4OAf8v6O7mHo9/iQzWAdIxKGLiDASUPZ+F
5J5Fnx59cIfnF2G5LvACgP7s1NUworVxwWbO4j8rUr5ndWXcOE5omJ8SonV2lu8/
VG0aUQVpQaXmqR2rBcOTCqN44TxBd8GSGipg8EACCSe/tmjVuh0Lwbuv+HxHssUb
OryMSel/eIlwWLFA+ABjvNvBAcNiGIvQPibdFxWeZdYzbbnPgNB1Ka2dC2jYFCQI
Qf7RPLmCWu8nz/xdKL8zKtSXOdgMpTMwWE0WEER6bf8JEuWz78lVFlnhIFEMtjD7
3BBkJ1ze+0U+H+kQZib1ncNhUhtYYAQmDNnwAoNpG8DYmTNzY148U9ayFj09oTWd
PXoPVwAeJdUI6tE/vcaetK8Go+v7eOh7V1EG6iAIWBGc/bQaG2rTZaPFycsMi7/u
fZ4jyhjgPbBEFedIHY6/BlOm6QXgXNpVpj2fRC5DtU6LhosCXf6iuXCAIEGfg+dO
4zj2Shb0ADHwaY6O+zFEAReRH3GmNN2HXplSiK3SuSCw1fdAkwvinOh5ntGcroZ9
RMHel66jEn5YSpNAGczFpWgQJEmieROAeHLuUxvan5ye29VklD9HSxTWS8m21sbk
PYPTZl4gbjM04SyOILiOkKCZsAxNWs8gbe/Bbx7xXYhSZXykVWPN5Wqakrtqsknr
Di1hmGrpuyoVOAIQzhFq4fNfx4wL2aSdcuQRblYDK7eYeoflpUGcVSBifkoFJxgo
yeOc/6L6OzYCZzvCjWJfoX4msquscvxy4bksrCP1W/UcU95CuujHxDjX+/7GUCAC
zyy7OiNFnIU6mRII8qwROXCCS2OjXBbyRsllmINjNuoc7AQoBh59CH5yu/VNfAIa
9KPnMTOEkO7UqUwmWvCh2F4PZrDuKtumHkKVEF8/IMvOkZBVDr/V2S+1MiScd4bR
L4nxFtrXFFwpEfxcbOMyf9MD4Ec1SbRevIqjNg5+weNi7BCBnUgquv5k5WWiP9NR
wvDkG+CxfFAmyCoodhjRpXbIrDNKRndK+9zEVe/SrydBC8G/43kPTMQabqU+SmAr
QvKSTmXk2TaqPn8SChlql78LrqCVOacGZHmxRpv41xQDlvfLXS4ga2aPyNJupw+i
IpImDBlgHhZE1f1ukwzO1JRW3Fx1LZIzce1gFCvwhjCOiV+SU3QJYWvcRpJF7trP
HQn++DK92YlO4ewRtWFonoI2h+uO07lC2FXPsbEPQrZ4R6FuVn9OFW6FzQFBApqL
mdsDqRlGPf5UaU9pcq0O6Iw5YsWCxwlLJa7vCmARgGDwoI69TR8cyeB+feCRZKNp
roQgh355mwRZlxhmwGzAdKrrGQgw/iKolROyUe44eOnKXCZ/fhFGBccftSb1SlnB
bzSZ0RAfBJeNf7O/xye0uXyqISY0cOTO+7ay6EGsSjHI6IMiLfGtQhCLd29s5nZf
v+Vat8YROWB62AY7TdfTI1fL44Uyv9tIUzXSPXdzds1CJ+rctTXOa9TBfUNUXQEL
5e9FL6CoGuGD72h/0Y8BN/bue8LqzTgbOTLkf+hMdRqtkVlC780AMgjYbGKi83W3
d/46WjIpchDkLklmLoLUA6x/kIjDR6AFiijKdRiU0+VXjf2n/ss4CeItnBvdmJaZ
WMQGxPQRlQNbe/RfW0XW6sxgYXuylO7LZ30M8Hm4gUifckYFC6xkFM91CJvpvgE4
jaYfrVHqxVbH/mKdMPP8ycJnOiN9Sa4/u41BipgrraRjVjGhbZjA1lghL+DWMAOo
M58swev2jOZmXw9shpEv8U2UWUeUoxKTgiPnu/SH6pVmI4FB0vkcpVQebrqOMJr4
3yEGJ65VCxAMRHbrP+KWgWWAYBMu6umMpw2a0ilfD+n9Y23TCN89i6JTZBVvrQ1t
RxfMfWiclVhg/Iqnj0JOt1riQZk+QG7ID0p+NBWQAxFvDDX9MXtgpxrou7oFwcaI
KXQI68AULjSPJfKhNjZ4J4Db4YPJNq/Qkn6LKMHK8HaoyxnSgPXz0/t5lPC/eqr+
DETORM+dHUmxPSjCfMFKLmHa774dn8NXNKH1/I4+Idg6aSOjhZTP39+ciI1XkvJB
KIX1BIdynVuJuH9x9cX14vihkbLQdjymZcjwuEh4ES+eLxBcPO2jlbmz+cXZ1f/x
JAStjCFXgDHAihVyin3//VHUqr5dSBIFvFWoMv4q4mLMtM30PZ76Sf/KYE6I5vbj
gjZbFX1hC+gXteOr0gaFtcvv1T+sTgpSHs0m8OxU7kgQfZMwH6dZkVGyYeWv8efu
diS5S0NOOPaERYO16jKJBS/dc4LN/cdqzGADFurp2YlNhwk8ZPzEPLJdp22Hzklc
7nmlRVCSBw433ljJjcuVU/gVoBHjAHIvxmzY39wZbqyH7T8Db0ms5c/xTJME9qk+
q28N7h0NvIdML2c0VFxew9ToxZ392Ih52AdYR2MMngneSQD8YVnmECMq3/z9mUfX
F7TezN7IpywtT2xOxRLnVJy1kg/wirafB4uT4P+24uLrU8FIQeEHjPizp2chijES
60qxOPjzcWtP9kIOFReojBA97nl9RfPO8ZxciH1H0i3cI3+VhZTmGuSCrVaTa76t
70iIaIWOlnFq/+a+tKyfv2htAC/LDkb4vRqviFBFLlgK+k3RZQ4IDFnUBZFWOhDN
A8CYP5ZKPRMQR8hMav0l/pBHTYJh7mkVGd89M+tq8pB8lg0vWT1bAOBuitYFq+DT
O+TKjpKCPxRg/xHOpywg+qj0xSgc5MEuuMMrVfW2pOO5MfKikcFipi9+LSElXbtQ
yGYwCl8l1o+TQGu0BJtJLqbf+YSeO+Xkb+NgyWfIPk+xM/coeH+XOhc6XI5+CPua
mxIHwlJTWHqeBu4FREYmS41EPOWGgy88VjZarrUAjVDkrt+Y8bc4qzt6ggLyPgtX
0ix0m05bDiufCKX69mkcwQLhT4V9A9BZPK7lvDbGTO2dMpt5wGU1/XNhJQFwjYy8
4xveUH0GAEeUwKy5rRIGjPT1WQsFPdhfzxKAD72WAiSttmFpZps79TjXiwi4DAzh
Oz8ulBX7hRDXk6SqvZ7zwVUwK0Hy/uW4IMgVfDjqAOwkSPmUXsdaPXNicaPGflrt
BMRHHjwWAJAgJ+dGFEo40kOqXCwe6ijC3dgldaA0iQ6RFiDDZYIOiaywTyBJvTkW
LUwtJjAzY6783oP9YOyg3riBAn+EMJQK5EOcOcQGmQWKEj/tdlqBrsEKBcq+A0jr
Dux6Yd5nmpPepvRRJfpp+UMpL3um1yIir1hJdYj8TbmpaNkqJsqz3xDfw7L8NPlt
nlSKcCf19X/HWjNNcjEWzUKPNatEmmTpMFHaSh9i3WzSUPUu3TD5L++qFV/p0hB/
+MSPLOXhNuh4V1UAX6T/Ox4HST10WPMsYpDecFkmVm91qZ96SGhCOAsBqZKbQugm
AZWuV6D7S/8vHEkhAyH4TsaBgpVELIrs3bp3ERKF7MLpg35IWyxAB+A5YUYgO0zf
bVKeajncOjB+544Hd+W2u2ITH4ZbBXxgCzvZTyd4cvODUtsQIOglu2riuf6wnd8j
1hzdB/0RlJBpsKhBEX9ecv6jns22srr+m0jH/UT2vEkMIjPg6uGgp/GsAm8zEPMQ
wRrs6ph7Q58r4I/3OzMv9W7pPlpp3fwJ2ONvSC24Th1dx/EDWA4C2SDql5vrii3e
hACL/2co+V+ifqDHlEKGkZfwUmdww2fsTKuwLM7FMcgi6CdfQin2GTtAlToaUc3s
rfMToAd0JAzhmkyPHuGMTYF4RR1ITBZEBEswlTcBCTA=
`protect END_PROTECTED
