`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
J8D8zCf1G73kivOgPq8dLzVCPQkDTl4sFP7tiZjsj3L0P1z4URJZXml5Fxd1FMYl
NM45aHKuhT6aLacFejWNq5Ni7xL4wgMkix4PRYeY5DJF/oEPONgir5awcE0n/XBN
cRtJHjBbtTKYmfBm9Pn+T6u+PjqqsNHJx+yq2E9EvCvknZygBeshnWg+bqudExrI
omtJ7SS8/wqETnkY6g2F+UucFEkCxURwI0hkaP31l43j7DlNPHSRboSae5QszsT/
hI2jG7j53qxOGmI9aRf+rV9yfvlpR52ZzcaoBta2eIQrY4h0innIKtQcYK/ULLEJ
bahhLODizF2un2y+fgks4BWfF3oxj+TnYbOQ3c9vp53SC0X7XWZXYgxdyXEti72w
QqTwDoRqSliodeD6drjL2LO1BbB9/0qPA3RQdu/yq9PxnfTNME2yAHVH9Uuq6JQM
pa2kbGpXJHbNMaL+16/LkVYcOdsFWTsB9LCxypc0+lzH+XR41J8zrQYcnYe6NV+e
2o06l6iELso7Sg2FGH4VqNqDQShxvVYp+GsCiRrqtLull/gt6q5DYD9dzsgysJAT
0kIw2QZ0A8K3ySg4w3gUfhdfHFaAvrZ/aemEcMEnA79eGTd18mlHueV+SpogX+uy
qfdd1ZFXbRL6M7btXJC5hoqRZGwxKw/zeZbIJDbQdekKaHe2s+5W7J0bxDxjQKGc
qVfCyetPb68QhHWLcFz0DJZAUwhKAzOHE1dXnzQTt/bxqq6MN23h7xikhr8C1k4N
4eEr53ZuC35DKRuQ9oaR/aKOn1CdpNICVLBUph1wVqXr+roqIE+i4Xkru3KJMawc
pjuhu3WBXP2f6yEn0Ca0GiBcFRpkpck0APBKCb4s4F3CNtdn+LAZEq2nGoT4yj16
IX5ba3Zk9WxyYwZcnIL5ZMFgckOkFRkYeUVR/5eAzf/TA9atBkCh3n48pzCMaZQs
SxPUp/Eqx2kuMjSfYGxpZhe7aHT5wila87eq3Vli4lDoVyLpBajv0i3+1HwmTFHV
6585etnCRZ20WZYO3xqTw/6FBmeIsESb6Gzoqob82lDWcaNWJa18UgqikfE3yAng
6r977oFr6tc1YotuUwgwhH9WX2B4t9dDHzpvSh2IU/ciq3gRToSnuLrDqc/7ATfZ
yi73VBmmfxX2Vkvti081jON4hAv5gTSMjPBdbDRUGBn3SRi51YR9LhiQynNo0Wz0
6OEonYz8kUri5+01j95fABBsZpxTCTjbfZl7keJ5nvwM6wO7N3WaHXI++4qLlRTC
vl34xhgVkFhAZuMTwAu5W9wyuEfglvGAqOQBlECNPPOTHL7ltQ4tIUw9P6PMTmFP
D0fKGI0EiP1ONbHrMBmupwRQdtszv0K3bBvaBhSqa1STvXZl+H8s0lPVFvC7Pcds
8wANqBfrsB0Gar87BlGH4ikgiPTWO2SoH0n5IuzrnM7X4ZsvsIX1jRf/MqEyNJm3
m7315HiY9SFlhhgL+wcFkbGHW1ypuh7DWPq1jJ75kSPpGpiYTkEHYwN7VapmK48n
DZGyE92oQ+PU5+JGTO+IFp5LY5guuG092wQEUwrcAlL5GFbpw54jboIMIqD71jRI
5wP5JEdQ+TVHdry7GpqFMKrdqEFyYq2NrKbkteOEtYJn9dDj/ZrvWeUOEa5kuba+
ML7QMmJ0cCsgpHRTQ9SwDggX0ePfxkzGhpU74mLFmT+U2DBw8cdlKzq7tplROdAw
DJCWroA9jVFJ44D3YYaJdmNtO2yeNRDrHaPksoLqwPWNZzXfg19zCdnEmYh22WyO
vpoGuhrqTdYa2bSW5bllzTVTDIseV0zXAGX50lhyaJ3OZE6b5F0IYCBbOqSTH3Vh
xQ3BYPme0rnOjma3gNKmDXKmWPbP4TyW4qTmzvWCCFRHY3LY95mPpDdot6tp70fg
U8FVXBa5IsO3+A09nRYyNzQ6Csr5RhUJmAnaqu7NaJmX23jRRrWxT/uTzjJiPIic
hLHbsT9lpBB5Y5H3VMQ4SxdsJDSOReRDuP1ba0T0QbXa3+6cakN+0CnJPVKXhyBb
VipHdQG27I9Rn7BP3YuveUvsbQLE6DdaWR58duvs9ptskR7Oydgf8mD9OwspmQi7
YsVnHcoMMMiHcjOhm3aLw0nBGq1+QngAevft+uoTtCamu/d/1L3GRddimH3l6rLx
cZ1Qaucp3XgCvk5dFwYwuWc/283qdOOD1omAa7t2eEGYBUT5zGuitf1cbGYbnqhY
U6lxGKdlllltO/sxphz8rnPLZQVCTzC9KkBGeoW5AR2iFPLUyzNfufDukShLdWMi
LOL0vj/AtEtIptX5nHD03Q==
`protect END_PROTECTED
