`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/tPntxONnSfI6d7J0RmURh7gjPYQqacN0YuPTMCPTCUMbd6yVpKT1HiOq0ZyCYN2
9p2DBFKeliF4XBdh6vJ9GHjJV1sPaBT9hBhW79CWVq5kCu3NUnbO8ao5Ee82fEj8
0Df/l7fexfHZmayqVm0KDjw7YqFGT8W1jAwSsR65Faax5At6YUg+2vmfLZVYwdva
nMz7G0We0rfL6GV9jSfwroO/aaFz/quiAYbkExJHdLQsJKcfyzGMmX9yhuitOWM3
sZUaZGWksjfWzGOFICeU+YewTZqQYZRrpPUVtEOBW811bUoHEMLy37iOFNOuQQFX
3xcqkekTEzhdv74toa8spmYkL/mkNf0VhEHIuRc5jBGzS5nLtphEcprvAAMChj4+
HyjtmuCBqyOlRn2KMrXzHKAUiZQYgzf9uihvErUEimHUOdTXb1Q8wC2gFITWaOFj
YiHu2b5j/sVK4phfs3El7NU0UXd7XyE2ce2vNXA29cA23pVKCWvc9FN9ITplNgg6
NzrsGjwntyPd8zJU+r7IRn/PvFj6JQJ9kgLW8WVFCWvu0KY34y9RxGpvrKRzRiyR
tUdiMPIo4CER5RW3T3OhkFTWFMWJG+vqNjkpjhwFQUntLzmaFVvsbDgYp+KWnHDd
GPDQr4r2DPrnlx5ZoXWNuxtnHAIo3kf+LRhQfhbLliTIS0hbh+I5omhtUkmNyiHI
oQb3U69G/BG37oHum3KRLOef8hAfZGI5XheajcxllZgDuiyf2VOMTUzhXVXuAVZR
JZoScSgSgVWcb6TbrSkDRcDbndNsSbZT6y1ZjgTLw8ZedDrZXtqadNrUDtGf5BgP
m3QKD8D+ied3ObubBsP7c/YqfBPFsqWVHrlza4bsxhoCxjjRdctwRG3vFEpR41GW
CY+vhNKaiEmfngxE4aD8GJdIEpyqGPz5tleXRtgJQTZmOAb//HjpUlvJsOBLmOT+
/So+ZG1sR7aEruWtoOURRRbrNCm1Sdj32WcBtWJqSnUzZXmVkryAh/xbmOGq3QFV
R0ntSabhEjn7BmlE9CGOYJcYZe+CyoKvu4sSowRu1a6Cu6+BXH6m2cTl+Kw2wdwe
u6Us4UrThl1BCU9UFYEzYTnps/Q9Qhf9+p5u8pAaj45XRdxcslfs5uOOfiva818M
MmlTttXYjIZs3XST6hXCg0irwuRnLFCjBAerXBByul0HgjNU0MzPMjIkqpvCWkpM
lyZUau1cHyrc8QSnVKA0Y/HvIvT2taG3gd4H8AYDmkXItYLOISSDU+KMjQRbaYGn
n4n7VQYN6Sk3pwX7W/dstdrYjmm24ZDvmSB1vjdlEQRn6qME8Hr4urD528DKhHCG
qyUKRHtScEH5xC1QqN7TkqMZ+zxG4snGha8les1xGv6ytGURh+HcO0vpg7Stg4OF
S4AIA62yf01/zRqAhJ7MkOy277MuosunpM5tg5iosjC1Wi/+FYlV/fv+LppTG3a5
DseLVD+WdiMuXu6ygAQmzdETGKIZSqSEOzvNt/b5r7FdaFanatqs6iD9JcqjKXmu
iAOZ6/HMFiOg7mOpfWU1p1jYMm9ZYBJQppbSPEFdXwSn/wEv/OeIFTcH4awdB58j
G6rnQ0L6Le/kSlHnZIntw2GkaOGY6E/acF2qZfDRsEKEmoGmURz5laEbnwvIcKGG
u4EZoV3XyqB9H7Wy9HW6gFIIPBMODxaM3Y5fnT3OijoZrMHvLkFxedN7+IvTOyiH
7oBL9wfDMGtFFsKfwZMcEO7a0v7T6RiiMMvQrsFt9UlDinY4okxOmJ8Vn1LHzEgB
3AIuswbPYT9IfU3tQ6Qkb30cyCZyTVsQ8CGgZUogIpYT3goJjGzVAuo+KcR5KkD+
NwCCVcn12hLN8ASnReH+BRZAUCY3Nd5ydXNp0quQRCv6yJiKaEyZupWezDRQryDL
6PPZPefenCQBKQjk/2gwPypaZMHQzTJz8pJXsIP3NHdYpb/A7SfyBKvSA8bpC4wg
Ip+P1wE0l6IeWxKvfrsZJ/0/4wa6pex2hq7NnRjv9eZpvZjUiuIMaIid6a5+f/4I
IioHp6dcIx0aRVQDU4gVe7pyUUAQiDRf7GAwBa0hHfcCLG0KRANqM0JbrtfLwanw
tcUhXdie8mVwWIBN86Dw7Yin807wm42hSMjhxEJIqq8r8y76IqOsig2cokiZpgxV
ZyZLxO05DqZu95kYswEXtFW15Qsm/hWoh4QBj6CsCfImf6mqD34CSB6HC0H80P1p
b+aCiFlkArOqY7/tE0mfHGFgPGp9xendfX6E1fgzaCuNHKgI+4lbM2Czhio9fQV8
nN2dGVG48JYFO1bGofY4Q6USZfLN3hdRvgpqToY/fADMLKO25mkdRmdYkICdwpEF
xWB25wfEWjPPGyB5fMjk75xLiSD2Hg1nfOYhjZmVLQjh6HARlASgC33QlkBsstPY
KQePeRs4AarzRT6SXaE1bQiGffKp9JVbUJsaWTnYVFjWQrVbkNq+whaUowH10WKs
63BZvnj8geb1B0owNqw3Q2RANK0DqzrwVkBxjMppc/vBO2rhu2Wvbc5i5TDScGc/
hT3zVm6NXz4XdP+Anuplf642FwSuaqQA7b22DmslyBYfRAMTffFzI0avC/5dBB4F
q2I6ArXpvoQYTURY8gdH441OiHGsp+fVAsIbuuSNRYOJIHmZwQSZXF4ifNj0rv8u
1vZQsvqLo2r6ajIYK+AJJYxNo3J/b7KgR07FbLvRN0IQDYd9PoYS4NXiPhpJEpc0
bEbwZBIUih0N1NHBxdtaI+fTW+8WxUfNS1N87KedKhKRcNqhemLN7BSQJyHoXiRz
z+OMowDOoRwVRxBbhc+eP8Wdn0nM3OcRC9CX8xBIAOJ56z2KDW1+9hgvmd3pBstr
ciIwyFqBJuNGKwXFajlMtXDz0xagCRvHtLHFsM52mf4gMmd87EoGYpkIEP06sA6s
nll8EG63u3XgnNo8BGjjV8275/8Z82tOhem8o1Ik6KP/ZcMQ9rf51ipk339sw3NR
`protect END_PROTECTED
