`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ak3jhGcjArRg2rAu8+RRvNY7qWl2Egq2BFF7afdO+lHYIZlvXy1kwunLrCy0BCgM
+ceeQh1EYrMc4g7Uw1lCOKMtfHGVi4emQuupDY9cxF6BA7yzEYBhkehNWns8Y+mo
0kSZatYO92D9uQdFemI17dMb4yEiDDJhA54LduNRgwKslE2y6AO+JzcFcIl3p0ab
TApu76GGDo+ZJDP1jUTdHNOLM/iX+o1VtpGdl65BaVpomdenCtKMTocxA/t8dwb+
9mG5KRPqezD0NJHf6cdbLv698S1lV/rt8/Yb/lZP8DSPpeQYAWc2WCIxC6Y/MuRC
dE0MXA4gwWSTGJFdQddD9UOsOFVrkXtHRYCnqIPg8sFPFVgqX7QPl4j05jaiKdDL
iNRR6CZfbvDhH+O4RYA2IiFuv8y55iJpI3ivzo4XFN+trONbI5msel0rosbOllL3
L3/IApx1czSyNPBcPiHLDeI5ZRdCfHtVGib4y0xIPcKV88Ana7LIO7b4mLulg5c+
L18o18VvNT+g5fFwVT1WqFLuAF5VlfewfZs71/8Gf1phpIh5StoFd6jasjfq2XhQ
hci0wTiX9O5XeTPvGna7nIc9xA4/dm/wf674SXZwtKvN6sayIbNqhQzcqiq+4tJk
sAZ+HrE/GjAGLeXNocS7sbtpopPSzJt7xvJDIAvphw9gDeFO7S33g6I6mtfF3wT7
BpwcAVZMbAhbdTPUDW+oWADPLfQkmqo551BWhPA+P8+lmymjIfITwggZiN31z4xK
WiWIP1MFjay9C2RtBXN49HPw5YQOmqbzVx553/UbVwfMfJmNdx1akKNrUbsJtEsh
1zqD7D2tba+QawVPpmEwpFIaQGhQjJg0kF4JeooYAAh+VTCaKQW3aFyHObNttjtN
8dN1A9owYMb6rGXLDFbnpdOG+3drZPMrdWccxf4fu8Oc0iJp/cj2UJ+zm49SPACA
H05zwv0Zt45GTGxbK8KksaE5lGXSs3pFMVsbTgdtdLTsLNDoGh6C8VM0agPmIUvi
WgF28Dy6QsowGtmEFdear0gFruWyAgKufk9mNxOWEelTonIsiLr3D+Lm+nKua1kp
2w8KgJ133E+/Gr/UvG63fPBHno5I1jS1ZCLCadSrwqms6QYzDVM/gQQ4zlDKLIWC
H2Pl1AuvfKPfQLKgIwf3BIj13eQAGM6yMY9Pxcru33F6dglXvyL9ocZEpDGnkUhP
kh6VjMofJlRCruAMF+/fkcE8uIdFfyvhKbHdn1WH3tmZTcwvotGvpQQwG8JAQNkT
XlYvu7cQQBYWdI+keHnkQxwKZy7i52pIz0+yA7nMocj/uEZBE4GXg/1u879iIiZi
66KnGTT/rTBedp5AjnIpTg/M3JW2i7YdvKd+6M8SLjzdzO5PKTo0VLuWmJUynmbv
RVKTc+cxO0e61LhlRAPJBHCTJns4KJY9U5oaPQHK0OfY8hC0OOxINFc6+6tZjDHT
7h4lgPjMpJA6Muq7aSxqRa+7jQE2YhutxMNLeYulK+4XwQXdhiPwIcjC3XsxxCd/
PA1+0QLbKv5dPVwaTiOWynHP2R6rlKuJtWq1gVPZZT9IgdGSxtNsuq5slfgEBBkZ
L6aiHACpR3CZ71N1t4bUl3dzPrZB2XUwunDs49mPZLUETlT9EWe4bVqYIb1ze9+x
4Qbdwi4gjD0GNmepMvIPNXdKbZ0o4wSM6oEPFTFZnUpaymZWgfsBvI/lCuVDTfVX
YeIikvNu01xV2Q8JsCehz+f3ucX59aP2qwMFVWnnxYNtvX7/nMS632AH248WS4LV
jdsoI4EhRXt7PPfiPc1wYvKf8GsB73eO43uGIY3DKdpFRQLtQjtsw0jJB9O3xXhq
ciJMDFbbNBpOcA+9gc83bjalJHoB0CwVKaxKBMvCdsFbA9w2fQ/3uE0eqxkSQV2i
IId6hsDVlD7HhVPFrwiuRCI5kR/LkXNhp6mYKyrNsoE4fre2M3ezTgC4M2+NjAS5
Af+QfsF2b5DGRC/blqP2vdqrqG7Su6m+JLotXUZwkNjssKVV7noy/hXV1xXFYv/X
snxSifQ4/V2st7nEooLcsraFEICndqyv81ZCfhWOzA/kauvKvOkQbvMWd8FyFyjv
+pbvcgF2VxxpXKrfar60/X19cS91HLYShYH3PVWxBs69fIluWAOmPcoj/c5CBE56
WLooKgwOxxYgx0BYMgOHIwFxfC6uiOCWiYMghpxpDujUf4a51PP36U4yAwuMvJhy
N30WuP/hCF+Hec7hd7ssCoCtBDn3u7gf6k+g0EYAoi8LCQdKlekZiK9Zwe1NM2pv
UHgpBa2aMf8K+crx2tyeRu8CxnGmGrdvUnPz+NYfWwfC5it+B/I+lyJfM1q7vGb4
a4F655ocm+dv4T5KelJV5e//aYG7Xj6etimXXiw8zQg4m61lXzpR9FG1oR+C88Mw
sh5Var640U2wMHZ/e8g0rB/OAObi691aPey0UJdSRtWSULVtW2ybMmWg58FjDSUD
PYYzDML6T0ipJGXxHHQDMU15c+HpjI8/ky+brsRW7byG3SRqQGZtiVi1HNMY3jIR
DtCZDrz7KVIkmaHwFfwlQSzBYb/9iyeCzdpkgXHg5gb6CVTyCwSi4v9ydZFEQ8qR
pTnGr2w8RpHnnJIyiGXyZ2Nh3jjcreV1nVud81jSbv1cdaUK3FKEU1E0+turqUxp
UpxWWXhVy5XAFkoIggRnN2CvTwouInhyVEa05pFrccaIwjHbzT2DDE93JEvr3lty
KKhOGna/OValOwF+gVBkHp8OK8gaC1/FqtDev7etYtOGMV5fdxfxlxq8MCc8OpRJ
zCSVTvRAxLGWmG16YfUeinVbaIcdNsHZYHW/0vSoBszxbK+6YZQ1h32D9T/eiB6r
RLBGQ3QXOHkq097/V9Lzz1xUbC+3q66nFJ+wIQOGlc0CFYzmoi7oFJz70s6P7vr9
5MVnSOXK/QWN56HY+6Hk0ozMS4MQYltt47Na6mi2hWA90r1eOl3BbtUDOUpfLMgo
/SuT+uokgLVY85Y3UMIY2tSSGpQo6Kpgy1HsLPxv5X0Yd4tpyLZnCfIZJZy3K9fQ
41DWHVJzVTzCgkUyX1LpHPBVndMTiZtqRGyx2PHh3kaajGqtWh5wqe2RJpo4e2S4
2VCNa3CORf0yPIoV99eBQm5iyV88H5yZNmParg5RrepiofAwumP1bR+nzXncsJ2A
D+kyi6MHHzkY32npPptCejhwqoAu8d2VNGENDR4B1HFbS8Yd/gWl6zC7lbbPyqCe
NSmCqDPI3pFXGAa9Gdy1jkV8K3is3jWHXmg2T2sgC19oWUuobtcszAG8vZWhe+mR
Akonfj+1Zvv/2WgQQw+XoFdaKhIAA+js0Ky+L+F4BH88hbClFDfTkvJUdEo+XwZN
wPnY6URog82HBoKn+XKj8xq5PGVxl9qjVax54tjjjJisOhygRlgUf464Yd6LVafg
oofK6chuYogaR9xCY0bobqdXBesYmAETTuujZiYI0sM7VQn7nu6U9d5lgHHO/E29
m/qHkzoBcWXPi8dAA8fSEeU/5FvJsxaZKBUji4nlhfM+agKznFbZ7wqQku69Q8Qm
UeyvouYtx6a6ALjO8jdqAgG0kJ5MQgRZhAnzF8W22dGZokwpkwJ/O/fhmjTxc5Dm
IrGR14hH4WVeDHq7UB7ru4g3sAZwkoEfaOf4zZphR9C24gOOJ/FwW5XjVtvAojXt
ryLQKD/skarr475ek/ha4UXAiT7zwT9yMbUHTV+Fr8ZT63JMtCx1sdod+Y7VydV1
MJyMXf/0fs460ROoiBzUAQ==
`protect END_PROTECTED
