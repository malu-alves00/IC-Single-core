`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LIisKbbvEfAjaRMvlhdKzT+mdKK7VlITRfxJugZbJGtSBgJOLctAXy6iecQGuWAV
dwNY8AcaZMN1i4cmWlmcTJDZ+65gr2K4QPWkKkcwhly6FnNB+4ppcdkXPrvIzBsY
4ZoG4hYA7gVGOCdwgZUepEJhkwFXe4l7Locosu9ArtVwT7ZEjBrSE22gSM0irxlS
3L2E2ukJMrxqZpgLBwVpBoiC5WoatbShakHBaYlZv0A2rrl2CjAmSH55RsSgLebh
0dtHGjAHHId6+96jHhkNSCVb/6aEqcoqOGKqXW8PnwriUZRNTFd2Tk7CqTlk/zGc
709NmDqhSoCNTQgFhOMYqkint1lM50Yw5kiLwwAR/Yb0i895m7XC3IcKWdiMU5YF
UwafCdgA3HQFk7qT25LRimBu4EKqH1sLfIUo0Hot3bZb/IF3ybj682FBR1GCjRCS
p0eteCnsWAr3PbXmahF4VCr17dIz4cWD5XFd/OacUhw6UTa9CcRyuJO3iJkoc12F
upDL0NmzDZFeZK0mULBptbt9N0+bpmB4D+I4VBk/hY0c8rhN63J2N7zNnNw3wuiR
aPlw0GS/tImZcJJAaEOq28IRi+sGZ3K+MX5IwUczV1zzKHrGmFmM2cpUbDNzDseQ
raIiTJv0To5sprq/MNlbNNWwvDQNq2jJLly01x/gfnAw7SWpskFgmByXkFDntgQJ
hpLhX9XG0E33iiuCPFdmSMZwRJpeyyh7YRTQ3aYANDh/88JoW8nVfsYaXeUs9v2b
rJswxdmTCe9I6PwBKTEGTYhXIMjrBD5/6Fd9vBAshNNZaWcxH+PbAhg+14zTuzBq
auEsiZDutgOxbYiPSZjVbZAwQ9eVy1JoE+nibzon1bw8QVHlFsp8/J2448lL+Pj6
uoAF8zKTYvIkLAAOtAz6C8al2O9Jq1zWLTL5QQKsvBqCo9MnDQSWMW3w9kpNEJiL
pPrpNdYVJs+/vYrG1Zk/7Cii2iZCeG06y+10eT2ol5cLCHXu7RPU1gipuEzZ29qG
4Xcp85sdjtQYwjYISnmjwiagxfLTCQvXiQ1w+pBTA/oPri7iQRg0Sq3697khyH+T
t9iZ7je2XbgBRp6TK2k1SfN1rCxt3BIrbB1N+8bGlvieCpsVFuUuyW6bR8EoTwQq
mdWky4326zyPICp5+83qr9WjqndmDVrHmvbexWa7F505uY7ukJ+XTEjAUZTgzmQd
D4QP0CwIDcqxAfXpHdPRIJ/Z9IpVa4KhaFhnHirquJgt9Rc1KCPtSsxn2tslvZSD
oA+aBm4cfs+lFYn6+/+7EoMDTvlP5Tpmlmr8YEA+jczb1fItPPl4yjzQYtomgu5B
R0IhQQr0LxmjbJB+gwAEfQ==
`protect END_PROTECTED
