`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ev2Yn0PwTkvun/388iBzdMsMy86w9oOkUKq+lHkmK9G5N4zSfjnTYvkdM/y0Aigj
ph3jmo2KmsDpnFw5Bgr9ARwIfSR4UEJTs3Uf/tcTp1wH3wZtBTmpP3Dz6qsRzMcN
FtSLwnex1lpVO5kn70uzt3nmccxIERLHM5OjsblF7kZ9pjoQfvQvbCz5V9Zy8ctf
b0eImNybS9EIeEGPx+4bodHVO1sOEkORfx1lx5JZlKmYi2Aa6X3y6cQnFmHnTIG8
5ycshXgRCCQ+SstzndekyrwHZ/TV7hm5zSGi0ZJYepYHOliWPDeOt8f/Hz+/2j7Y
QIbThpeI7aeU31nmwzGVSKi2m8aZSBb4cTy2FkWdiRjERRddFkF7eSQVI4lSIWog
fYDNbEjt2i5BDk/OZQO7pczGiYyh8VsbyxO7dIZALUv4RHL4mvvHuctyScyura91
TJ33JHbSVtowzPnYwEmLFDJpD3GdTJU6AxjNz8EQlkWD/vwVzsAbUaxf3PcGxemZ
4pClAcAIVkj+UCSs61iNArFff0r7R2ElRT0UBN7N0bC4JqbwDnPnIS846ULPl1hb
vMHI0uYi4oCv2pjHJ6J9D8EjHRgbhhaKXDfeg6e8Pa6OpSMdLjswLqq2i9zgQfss
Rfz/nyA2O7bdsDxLRnHenUVywVDfJ6doz/9RYJSyK1v2OcIm7DY2eY8fG1zKvW3u
/DNiITGst2LqB7v9f3zFkjk1IOofyo0Hm6svyT1YbQs=
`protect END_PROTECTED
