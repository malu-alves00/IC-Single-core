`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SQ2EHg5/1fc6jXyjfUDaWrLJeCDRdIrLDNriZxkZytP1peFIY08AcNXM7Mp5Dzl7
CuJyjt2h/K5yM7yJdm/k3eNE8S6MtPy41tB3Zay1ydU4Xj8z0fpoypuv89BNpZgq
tXSfuxGkVaz5ixRhY7DQdognewzq3vHWw+AGcxY9W8zpUJ66qp8z0v8aJj9Wxkkp
quEYmHrRi5IWPpe/Y3s07R1ztTAvr4fNiNx7VIntF8i/WREL/9VfccBVSE4y1SFq
sSqgmhgJVDqCXQzvqj2aABDj8Mi1lSRpF/QPAyvaZ2VxktfB1upbF2CfkHjefE4G
B6KvTC/TcZA5ZACuT+YroY6yY0NW/HbURWE3sUNEkoas/F1xag7DU5mozyTHxb4L
UI81ZaEgAUwMOCtealQoyS2ORwvxpYgVXYG+wzdYBqai7iIUIrzRxo9e9rotFW/F
Bi+ip7wy33ejoiVzSr0W1iTyDrSDZ211znOo7F1FOtb0GKcScomQFRu9RSt2IP+7
gZRDwIzFZPjXVxOCSG7L40p7N1LMZxna9MJ5/VktPyLEiJhwLX1sL0DaMGwAJwO2
alhWUFHADnKDcfpyS+DZ6YUZCccYgWGw3qiOVn9gD+i2KyX+W7koHRl1FMal2XXc
yqS0LkfoBZYrcWp88x99RqTOhGYlCWdkRyBYak+K48NjsnFa5ussevFyi9eM6tXi
n/GxZhXiQQK89ejZrBcMEaT4aTWLjwW8nyzzssGOFGzeBRcMoremfjKnU8It/6ic
ZBBoT1R2sN20gpZkwKfVvKKkXc78hx4OluZzmdGeEif96J0oZdJvO9hz2dbIXOPi
HktrDb9TQhx40Xo23y70dzwaJXglgGl9WzcjMtkFfksaHIdqR/6zxXfXNbmp6TC/
QknBE0i1kST74whKIWLJEpVgVNe/R9FhV2NbPmrjemmktFmVGkBwzQE4W+VfaolF
MAqDz7GsNgAKYBaBmmQI0tnLNyku3ZIxp8OgFRNnBNB4PGXNdz3Roh6VBTa/ackv
p7k4J/qtOeDIG7KNkJyC+viheFNeLYxJafcaeL/LXqmmCH8DwPZvxYABuTm0Ar95
v9JGDfeAi08W6MOmeq6F+X+SFdM1rgEK+XzK2go9J6aXo33tqK9zFqaihmFxY2Hh
wt9zEWYlg22HlUB2YswnxXzeJlH5dDklv67t09eNxsZpAC9Tl1QyzUODP6hONM3B
5bRU8rW+4XV6EO7xTxVnKNlQ6qwlG3i1YWcTUvLaC41OqMpt4tX+huNgZyQSW4f1
ky02sN5OO/1ryzyMqMa8xMRss0MaQGOCLCrHO+he9uoFTvtgi1LbLNpZRUKFMw+6
9u3WwNaXk1nrGHrYtsevOkCgveFfsNkQ2VQPaS7D05mz8JQ9vvI/QtaQeLSb6QKz
c8G3J2SogAbM/+7pzWjMguO83T5AKsrFiDNZqcgBJZ2uEMmGmARsuqOa0LYrjN2f
CYBDA7kYC3XqRA9Gow3x3gbKNUzGr7dp0IEtipqLVtliqfNd0B08jQ57Z+9wzAxE
7Fd/MlTsWkHgSrW9+puHPfjD3KB0hYgSdfnaXPbkLsTBzoB9YRQUjk9yogJHN/G/
L6XgK0n7krG+qcHMa0r7uNyLJ4t54QtnNqGNx6pDtJT5UuzgtoDjWLJ4iMW5VIyX
AU9FoLASUB95qi6tuIug/i6DZgO48XGUTJiXp3I1pzSIP6Zzpi6A9EmtsO967rhx
rl7kSiD+Xes0BlBag/1HQFedMJY4HKjI7pYHsMXesHG+7NLn2EhEzmWWxeSTVdNT
PBdBetR9BZKFdJdyIbs2q7yOP/6vYwYYMUBGVUE4NjHsarvfEFm0i2qsWQe8I9/C
lUwSXY2+ZJu3hy0skycMDI0Kef+BMuI28uuilZ7vZwUasFIbQJMb6ZzjHexBARhJ
FSkBLdAfWPOjSAtatinfjRJ6eon61aPVY2zu208m5I7KC4rw5YcDjA+yAU+2ngFj
UCXNkq0pFu5AhoUzruiCkMaSXJSJIrnKixeZ2dPs+wmjeCBknV/+2beu4Z9Bv2Ah
AHjUGZi0pNo1Kh1P8gU9c9LrqwWO0EXcYUESuxu0xLyn6vXnovyjz+tHHwSZqHjS
VleRy89yVZtWRWYdhNTSqwS6uKpxlTCDmGG3vRmMXDj8XuX+pcu+CycDYUZgocUW
2gSC823nqnGeqs+gbPOUSF78Mupab+IGrXzma/GU/JRx4YLq1W1M1R8HY3psG8dV
wlOAlbpz1gZQE7N9C9tMSIYjX2M+9DfoIdKCuMZGPBFiduppVp9OGFMRkxTlzkxz
cwLKVH8BvyunuJh0vuseKgz5bgcUSQLtIU9S+T/hzKANUikD8N50id3S+Q23YavT
ZEmlcLiPtsm0KDPejK2wP/3RXFV+fNPzWe01aev8HmCe5Vx8K4JvoSKTn6WaDRsr
En44jiN09Q0/f85C6sAzhwmNVTnVr8DNvTvaQAV8rZgeX6OXcdeKG0867jHs++VX
3bjFUhc5uH0IDW+QSlvQG5AVMJDlDzCldLx06P9C8fV3J8N98ETHEFjsI2ZBBIy6
hF+ewTfGmcY5SD5r5va+Z/JAJnLmlApj3fajUsxU1fQAuQ7LLK1fTUmS/X2Nx+M0
qa5BgAW6nQiek0vO97J5VfQ2ymluT/4TEd8c7GBpocZsZqkK+I9nPwanHk2k5qYv
hY8+jnnxMdCWhoIvavY9dPGKuSpK5ULa8uoFEiFVMmG65PRkUo5u+LOii5COSPQs
ovp9naUzJraK8p1zBF6n3YPUGxkSkN7hT0RtUT/DhJ3IvNPrfKyLLrKeoPoLZyJF
oIjr5B3cmH7MLkgdpgCar6oqWLYsJkDRVHFAqOPWasqjUsQfsSZajknl8jloQBpf
KJ9ZpdDgsJQn7+dxdf6fk54Je7CgEQ1NMW5Vv3jBe/3XJ+brA/OJlPVeE4rPmjuc
gNrbfr+73F1CMegDHDNlpXurHqinxh/35fxKEQ/1H+0yI9yjG/q8di1uwIkbjOux
j1QCJDyDkro/guXqvGNNug+81Mgux5Uw0d/BNDABt01hZ46ncwblyG7vWYxah6OH
t6SqBsPeq+J3g1uLvS2UP4qs9E3p9W8cwQNfqWRGur3w/Emu2p1SG5/RnlpPn8No
3BjYB/N9fr2VI2ob1L/g8d5guhzsEa4BA33rU1fHh+Xbon5unNIKzFnsEyHAwuuq
gX98fYilLB2CmsnTk86IEAVs3E0sUnw5OzJea/NBn/QYeGcGUQVDtt3WOYvc+OvE
1eZ0QkMtBFmrdbLCSoQJvdGZqhD/GIrqN2biMbxdlyzR2F4goXIP5YVecol4A17V
RuAYf4I++Sg+oaIUXhKxFXjb2ZUvpbX2cvu9bIhCshgaQK2GYFkJek0xFA/Cwq51
VLrC7vTXMICGHh5x0mL4QO07C+sr0tMu9h8yoF81zSxTiO6x5s3LdZ1J2FeCsMjH
xNQDiocpwFlCkVRiHyVvg17KiV/8EQ7gskse9FSqbW19YBEXbFD7LEDl+JGCwQHT
hQDOe0gvKvMt+0LWVj/Wzyn1RKe53uQYWnwDdCZUFwvTWG+S67Y1I65G8skmwFNS
BooQs+narOB1GzLSL5Ol2/o2J4R5RuxSSwLbp06D8g0=
`protect END_PROTECTED
