`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7ZcrsqVQlX6xrGY6CQ9kFsPHU9h2AvVGB1ODEHrhs67dVjGwJzMRwpHBp+4ECHR6
UqiPvLROKn8IlPAh0ACBsIMVtfBiIPX700ZEKziH+EdWhajn1GktmcNmPTbACDXJ
r+Yr4FRp95xZhYIVckZfPMRjOMaF/QJDvxupa4ZAxxcLxDQGLmhmzZ9BfqCH4brq
DEaumWyM73de10QutnxRQMTMp5Xg3JOxpGdK5rLfOAJVgIetMCKlxM3Pq3nXeIoO
YnxdS4NhfwX7ouEsIB4nyt3/awy9Q/mlYQan1dnADpH06xcChV3mUgTCoy1YRbpY
SkuOpnpxXdrR0vxZxXfctzL2PotPLYtHZNIGKUR6iDKR6R0spylbfm9VSgzL7Ohc
TfD2RIqigAcmxZY+1Mqu98tEwJCUSa1cR4c4KOjr7fI019GVeDZ+C5F0WU9iMoVj
ojhL3A4/zt8dPMSnrIuFdfFkppYR7G8n+fH8N6+LM/mnNZPhMCNy6SYKNEIDNAri
jq7hHPdrxs/1fkp7+DJ+Sg+wG8qHPLHAMMhwKqPcsqn10eJpbTzmsmKDO1RVn/xx
O9ShiyjCrg1v2bznO98+Ncqdj6xgmAPH17c80sNie7V3/7ZGAxDieej89yOXkLNl
7RKEkMnwA+B+QGlZhE7C9Q+hngXlMRBPbav0m8S55A3mtmYUXAvy/T0XQD2ofkY0
Zi3rXoJq163JJVQsGMkS3PBHIh0GGAeL+peGpAc3HRz1RG6LCDn/p/TWhfMzVloV
d3B4ui5bYnsAJiO4RIJD14Hhx+2YwLhTLVqssHUoT2II3G2Wb060n+lCTj6T986a
O7JZ98mCAANruYtb2hlLNGqXuqXLy6rQEcwgyO/Kdqpx99fcuyDAL5zDAoNoiOC4
dEwYhPFpilDG8FFVpv6hGvLU3I8rZYHCMdCyKo6ntqjcLCwjNGdtN332HEcpbyPq
AnNsqq4JZZENYVBDIiF9SF7Da8pGxEnFVQPOX7Fyuwty6X+VmUq8UC/43fk40dm9
RWnEDUCUZxnoVAHQT7JAfEXc5CcXbuCnrWHMV4k1pPRLgv60/nuk1MAWgJFjLuYy
Afsfsb7q0WyfXGlqBxzieaARV7VwequgRwXkmKoIBb++q+hxEwAg5FkxLrkGuS8K
QcjrxMkmTEmjibWy/WHn/7iLL32Y6CrQedvB6MGhZFbMgJxEVgUycgyMLbigeu4j
PKoSsjQs4Rr/UNyZYIRXWRcnJ0O69CLDSxZPfnIm0Gb6FPYDJnh7ih6q2L4S5Iy7
R65lsLWjDEHip65t+VS+6mbClxwfO+fmc6o4u3btGl3f3amYPROoiSnoKVpXARcd
4mlZXcvN7+A2IdTCHAMlpQsXPj0aUPWXYQXYUW2qu3f9MoS8NbUuDYtLhIxPURpz
O2p2aqEpBKzV21A0TwQejPzyQlb/r5evbulTKbSPLJM5AddhIStkH/3QpC3kIZzc
`protect END_PROTECTED
