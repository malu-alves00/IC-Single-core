`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
utib0v5dvR/SWJa8CmS/RrU/uDx4r08T/8mioo0qXwjc+WdiSGzpDSieprqGhkI6
MCSjr5b1xqvvf896KAPZv2bqRwjs46GbuhdNS7da/iN5NXWeq0kZuEupovqp2U2D
MzUMkgA21LbpgzlfgJEnpbZQdjyCnePrNk6LpNqf4nPFNTL6hfPQSPKpEp/XGQNC
3Q/ptuVjgACXnUlmseO7n+6PT+1CKTgoDOIlLLkRHmIRSxV0TQBWZoTKJ8NXIvJf
YpxvUcwdAv2u6AdGc1rqWM31hbRSbKOpYolxgA+S3LyQ6iPx51cmYqM3gT2Vk+jY
byfDks+fd1m7lbSRqFelqJSc8GhrQbEBT5zrbsSUy/kY6E3V4WG9rVB6mluHcOwr
Rcf6m6Q2I2WIM8W/P5ZdrjgognCPO0llpok4UiFac4u4qMUCcNVgrAvnEMgwhRYQ
6Gtra2v28fp5j9qDu2ovrZZZ3kxrDxKC2RBVRMny3x/n7Zershus4cM+uLB0TmF8
lWKDLrQGkIFX7lABKlYodpGFHEeLwvUiev+/TvltQAiDSNzUXZO0nqX/4OEY6Nbj
++IUoE0UWHLKngDWqexedRwlJPnWcjFaIUjYPSbOQwubT5VSeGSTWKOTc2YUezuH
kxxXmotJBEOg94ZzuOP/U57Oey/js98WTUskOlpFVdOB7JhFwpFUd9acPZy2Lf8Y
RW8BRv29zJOL5rQ+xTd7Q4hacUoLLBcvoeJgK5x6ymO5jTPIjET+H1jupvwWt2vL
I1CeV3O7LkSDDgzikoBSNsB/fKIZgvnLcnKeI6rTWIOS/IEhUUEwyBEfYuBjL8UD
Rmte0lWde80vv2YkJZILvPGWcTTRfhLtKt6Fk/uc3r66IYqeHXhNEoEjyTeRDcoN
PuSKYRB8CcjaaJQMGSxI1HMOlZuFMYe+l5KYsr20NrZufyyKZTC4qA2bLN8ZBIZB
JkjjkTOmZ7FeANnasySfzsey42iPiIYvK8Nu3dMWc74xI4ENDeq1NvyOB8mF1LI+
tkPJieqhze37Wl8oBDrraZ1zflbZxxCMNjAeOGdjxc5/TO82yOxCkj6Neu/tyP54
LoTxUrNgNBeMp4vSKN64ExE87Affy3TO+x0rkvzPIgzH9dvkFdo9wjJFYEMAUkJl
SXNzv6sheE8diQG48Yp9g+VRVX/K7K7LOjmoFqqBH3ZGi1ePh1tVa9EV73spV6Fw
IEjIg/oxj3G9PoP0rP+kUa7eXDSAO2laKwFFEQKxz1Ia90tBym6ZrfLh4qhZubqx
OEYoyzYHpqbZ6dTtixAOXfLxNsRB4kH9efzir2qpM4lRNlV0C28Q9aG71Jc5NKS1
+Z55PIyaZ8eF9w8Vo9yjhUmUSxCp8JXwsS4TxalFYPATdRODojRV9DcWCtkfp2PR
wZ40BRqtZeL+PPsO6uLinc7dnYo4vDsc4sKkJWTM0bu0lyfCWsJjeNLbbNsb+KtP
RD4mRIAj0OFbVHF2Hcudqr1nTFLiSL68tPU4F31e1ZJFU3PwWcUoqhVGO4IQGCzX
9bEt9PevKjPj8f3+FOYpdmivR6F3JFpeEgg6kQ3gMHksG0GHZwE6rv5tKHLt1JR6
nHHRRYZizbfdN6jzplX28bfjtpeOOyleXJqmYpnYnUOpLEsQ5gyCZ/CDP4Y9ffnp
JbHpNhXkdnbJmPLkphAa+d3cP8OgI+SUMNMR+JEiPCItAoZBa0WUtOSsgEKR5kXn
6gwvPBXu/YnSAMLppXYGjQw85nOmrAsBWhLXaBZ34KPSgXdkc29EA+hwtGvIRJey
Hi6EL7TWjINhGL7ARHPjP+1JF1EtZc+OMc5Bjg6G+0LXi4QUhs/biwHtZl1HY61C
152PRRc3Uj/XJhqD82Fn+eBQhQvgln6LHEvu/+FMoGnD2sAoUWddmvIwZss8nh+8
4yO4zPHK0KDTxj2+l7pJdKBaOzIR+VPA9JG7eB00FVjPKeNx6Q6ZzF6E1izZcuub
Wsvp0NLw/DgbovtvpPSaSeUZhIU64ZKePSA/ISCX6uGwskdJlLiWSIryQ9Uxzr1D
BZMG7yl5KETOdnhJ3LGuMK2BWRG+hpUnIknOVwozvQKmMFM0CrCPITxKt53AwbLT
0vpyp7fzLJpIZq2fbk6O/hsb+KTP9aWopb/avgOmf2lr6FNzs054aUg/2T8Fi3BM
6dEyWKvl3C14Xze9V0afUK7CkhtdZFixagKcYXPfXvPnL7tQPx1McvFGvJQPF90b
6BkAPeUa+1jvCs0hhgy3wnD6qZVklacAcC1hSdQd84xoDv60X24H6VEWiRsCAR5+
oaCUmrSHguFVkver5CnOzhuoxAmox907oMW59DY5DaXgp11hBnizIhKfM9kB8AY6
qKxyczBGL8/NroPzJKIH7MTClo5IWDOCE+Gqty2Hoya1ba4BI5t+6NbfWb1YgQN3
/ISxnmPBw9woQqKG/TtwIsiZYhGq1cdyRD9W1GFG1B29HLDNCrsyWM8U6Jy7x2o/
Civz/xurk7PFrTYp8YrnGGddsYhl/wAcECoQfvTqRUvV4RCFFkAsmI1tI3Y/iYEG
4VVGxBpdPMx/yzw5IatdbtKjTWqP0UG0vafyxze5jquT6C1hw+S6lKTdeOjy9XX4
5j7eSzqxey9jMtsqi5iD9BdNHweqV5F9KA5f23kSeBjcr3B4szTQ9I/s6cF4Di0X
LYm7zQk4pDrkTHIQfyob2eeiaZMH0ICtR7uW0V33lSAghwx2evHnOET+qy+s7sE4
/Wfb75sGzkEm0VOYaXh5yQrxC6wtiTEupnk5Jj5GACsKkSGpmF18U/gnAXYeUfPA
K3s3fUQGh3OOybmZRvRtFhu4K6e8YLonHG8Uoa7WAlHbySELC+Ft/2ZhtUtZJpF8
OHX5OeB7vXRsfV6YTY3WbBl160/8pkLkPbMnzva7j/s=
`protect END_PROTECTED
