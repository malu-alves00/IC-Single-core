`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VSStCKUi5S3DRYnMEWo2SV6DqCled8XfK7f5sasXwOK/Nl8SIK1HeYTeFFdt4gSO
Llwdp38Z/LtBNeD3cYC1VvPaCC78FhJqEHOZQ6qK+3/cJ9u8yQsdKO6ZT5MY30Vg
m4Wfs/968prrm5AL6GdwSRnWvr6MPDRPpYckWCHkFdOCwhgqux/xS6DPJFPW1DWZ
QRVoMOSWaWPNQGgL5MHLaGKfowpvKRnOxlQTDxcwGgWkrdNfDS6Mw1Hrd9BLF2Qt
suSCeJ3Myh8j+C9Dj/aMoonXndoDZyCoBPWF934umYDqlTLGfBPxYgN6nkaxyTeA
b1N2oziEpwx3VXRR7XoyR/F3ggkmBYJqFu0D1Wt4FIgRC/wX2cTUXM+OJUTl7eBe
RokfjMC4fi1uxVbfX8Wt2MPAt5CbUzNnMrnJCIBmZcvSYHROwaSu8mDODd0GXoDf
Bbiegl+coX1TnTCQCAPcHvQyrQudByjQyOqSf0yZD4duDJOpRTMq6vKXIhJq7R1M
L/0XPKoUEWHecHJDs1prLEw6tpTp0zOdV9h5NuXaLRd52UxzG2/UPPo4kLp6wkXw
Op1br0gRxbvccuKsKROjoQpNw2SuTCLLnv4PG6HGBkFztKSMcJr83/K3i8X+mjBi
J4FY3UpBu/AmhtqsIZnWGIH0oqUh+SPHr9RWsG7JyIC5OfFfoem2tj5AZeMWJ0Mt
g8OIIJjwRYf6BpD7c8VrMWQr1sqvKnzmlJhI/Ag/EX1hdQdA93jlG8LkHPp2srSI
vXhFnGBORQWE04bewVyAsylfbIC2LWREauOO2pmfrCDcxICt9lYQ6JvZCul2JPzV
oboThompfaq1xh0vB1ronoOTJF9eLb/C4ETOHET14S/bOCu4FBsLOKQ7PUnbsOLZ
h3UIJiD54aAwcw1+zD78CsT/f8j91pTzjCJYdPvQH0yUJ4J6pXsW31xdTeLZ9b0S
gUdbxckG0pryzyELMqGpheqizeHRXnZoNp9LsQDwxeTdPhtl0Y6CJJW0RnqsEYg7
Nutwp+YlS/Hs7cUPNqwBJ2lWXZeJwScYlNEF/P9ng6gF3UtA5rN9OEOTzvZbEODq
UY4nbG0+szuIfzM7zTiKK6mx2UiJv9JGKvuYvVy0uqo9agVpLbL9ZoLcEGW7D6dH
0DG9YIxg/L8gDVqcd/Oaf8D6Td1QE8utfSgtz2RYFZ5jqCgD8K/G9a6F868yZV1u
6kC0jXQ9yfZg2D6dY+EDT6miw7TB4DOu4XO5+a1dUJOyacZPXbOxbUtd5JIbOiWH
GK1od4/JPVNAb1pWlUGttAIPSBG+2JII1mofGw+65CYMLIwWv+g4Id8kh5HQ0Au+
A3b8KyJEt/RuNIfR7ihTxvwIKidgkA/wNOWNKoMWTf/LvVe5brEf3vneZQlC7RZz
9cDNQN2X58Uq7xFAe4meeIRuZcHIlC9yx/KI3T2UUHGIpOlkwE45Y8x+91I+265y
o1jTDVYFJNgqCSOYZLN3LxOV2b5BZSb3DbuDdxitZy/M6NrhB8toLwL3p6R/W+Zb
3gzjaLGCR0KvyRsST2yH7sy4TDrDGig8MBLpnCacQ+DO5cJycPX0hN+0CbXns8rS
bwhyiqtD+8QnxH2/CeEocRajzHt8MpHEfXYzIYsp0yBQTdaEY7siNmvCDdD57mbZ
VqZa4NQDh2X3d5nVAJRK5CMdJwlmNx0mhO49b0XGniubkzrCZT1rDuJZRFZRzTMx
cEmbIgEYjaRut3NVQ9NZ9lraQxYFqMbA+GC1AziunUpqXWyumOniDlk5iXmOqfTk
/OBHKhNfZ+GWpPHSmIHru65OBj13NsjKn7z65Q2l78jTgaeBVpYTTgD0x7Ln1+AR
BBdzqLoHYgpQ6ozMZX6CNArd74gh93A91BBgq0ll63AwlRf2NPby5DzW+Na5NYtr
j2aV+4HHrswWMXvMK3rMxGGh5+9XSdoonlaJ7UPVSZl+2ISP1TXBAjCIz8Vy5AAp
nDPFNdZBo3Ba9iUDeXHr/Lq0Enbwp/fx+JhA/kptJLRonFqmj9hFIUK8C+a8qlXV
Uez8tXggO7oiLObvGzRaiitNS5bs3oeWBXajluARmGilSNe0XMCjeCH5f4+UTDwk
cKYvUwiEXs7Uxy3BsrxE+MCx4XvoVwGJRQ+I6EvSae/VxDvbt7t3CY4jl7/gsvGF
o8C4kbpa9ELK0EVrnL7/8ZiE+uuaz4jnE3vDca+GAivzBzFfSB4wepjGFUvpX48O
QUkaQ0YKYjqlnqHIwXAJ77v7OagJeJJN13RMa3meWVKfJYmIVm/E5fnD/bacN17l
RbOoFLy3DLX5vrFfi67uVobrPZY4uNhCeIOHTxmE6Y5Ya7LUzhe0Aa0/3GLwedbl
8+m61Re38ypK0/uVOYgTQNVSOfllCp9/Tg6UV+tiPi0RRo1rMFF8UpkV3O+xpAu9
JkoDnC9/fDyHr9eWwqLItbHdVCGHntpvM14j1aezUvRcYkVaFG5tx4+42OrlTXgN
h3Ph+KVa4fUMWBAMgG6evzCG6n3pE+os6Mb4f9oxMbM0sCugzm9gGX97ohv2oUSG
P2SeK4Fx98v3HG12Q7Qiox7SGPb3wpEHwe02xpT6zQjtiRNB7gw4cYuB/Pesclui
KT8PuOgfjpvbRrMQR1zV5cj+ovYMYfY2m/Gk4H9AyLDzr82BCxK2+HqB6jdKbE76
HT5gLv3G3R/tdLbMoB/vBJPnMcHA6yHmyAGulC9Haamr36QDbc/NzV6o503ohLL8
CRcr2OXHelmizIAUo7C9y6AeBw59+8z3COs5Rf5vd23tgx9zffCrbVDJsAYZ+aXj
9iWiXiN+wbzYa2+xIV1hbjVPnwzfRiTVGCHiaFQCf7g+U/NQSTiNFwJel3mTBuCq
iad7URNeQsn01sfPVinbz396iRPtyF58Y9a++4gdyssZU2vLe1AW5BKVqQvor2dg
e+R5/IcAkPYffCNuo/3/WL2FWhJelM2e8hoUbunPDSBtjTCyrnin1yDwivXZ6c/q
ND9LUCz/Pas28QQbUluDkb10p10G60Lcvrp30EULVan+mgBFVsS/JU26ka7v9ZgT
h7Lph/107g+qpHkOdqiOsw==
`protect END_PROTECTED
