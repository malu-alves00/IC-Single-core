`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8cp8Ywjq8Y+GPwJ6N2tpLahilngt93pCuRPsgJRBRfnaharJ5Qe8B/PFrwNWKAvJ
w8rHxAZxdwMJEZSVRyypL1qYno08+5lVSxi2RYymVFeTFxYqoAOFbWA/+w/8Ajnj
yUnr4dLSC7fpVbEGXHqE/8Befy4TqoR0dOH8DoX+hxMqtUsyzBSGlG+9rCvqNHVP
yOXJtmNKWreBrcVpR8iM3Wp0UhCfHJklT+isWxEIDv4Z3V5zEtRjomiNRM/ww6yf
TCNXxAwjt5oqrQ5DvPHB0GDUDOl5Vzf3FZIyZ/UivDPi1miZhQxTzJ5HRdY6Zjzi
5B4YHYMs/VKMKTJ8BrUdd6NeybSVPS1IzJAaQW0YeJkvzx7fi8hr1vw4Eel2lp68
vNkZHVizETLZsgq7DJ5w7hTfslna248CH/LHjeQT2uw86o+usH2jUtZQJJPGzKnE
c83hwo6xsoqQicLjVrdMdm3j0sDWZhtGST46l9qaRd8+b360Ba2gKQKPAd1ruMlv
eC6QlccF50r83vBjfWnlfuKJz+WF402B3wjKcMNYQjeOG1bjbfX1LdO0l0AhPgcH
ZgpNuw0UL3SZWiK56EGvU/zbP49GrBMUQjyTzEUTanygLFIRmiTJGmR4jigdgks4
r/xbpElJ89Z1OfcYUIjeI0vVNrGPv5GJYWoDCFAZa5EpB9wIatj0V0fXo7uM+qv+
07G167RMJrA6P2f8PRjXRWaBXpfYBhWByYJxLpL3XuT6o9+uRbkbvjzxQ/TD8kMD
k1LZ3ICFnqp8cPE0U0/Urbqo3tlPdm6Mt3Uux4Rpm2bV2/LFISF239PBXWbgblkR
Gs+gf56qAQMrXElEZoyPaoWk5sSkwrfo952rkHQRXFaw6BzZ5eMuG8v+FLMDabSO
Aqg9kJOGSTU5BYF+EGcyz9Z02WS0Fx9f1a5vt4TbOVz7JNKao14QbrVwLRNds7+T
m3AjN81U6fWPgX0MOg+zYp6Mb9rQKTgQvWO6Hmsx6w+K0bS1hZDhlPlMSCD/ZaAY
GXX+lNzuBSGJjCvMCE+zywjXkwj/+VdRAYc5zhXYrNQFHEKEYNpuKJL/W1+t+UKh
2CRycwDDAolqciscfHHM2ammT7OeWQmtYPr4C8mojsEUAVIxVndUfRnzDVNiqp5F
vnXlr0yD3MhAaEtFhD8Z4m5kTG3SKueAylvGasDreWky0lh32JEqPVYS/DfxvTJ4
G+haBV/aAGy6ksHteOzFgRmAjRcxuzj2OFZr7l6juoqTpNHVNxrVFU6MjonOutzZ
TzQQANuCVIrkXD/DO+23XBsgeMTZc0o6yzyeEz/akBqHfu+/Phe9wj5nrIcYDKxz
tyBzVpMyrrgTsM/KQQaQJzxDzaQtfIE4PVA7yWbYj9K9FItg4SpLhMi0eZfvv/Uq
5PDQPiWt9J1J6++FeYdua+qjlWsBjQj+8tEse42gIUOLeV6xUk7uAGxmXL3gYOrc
IXeh4jfW29Wv5D96jtyqomRrPCi6XUP3gdyfRGOBlQTi/LWsBzM4ifloizeitFli
9jqn7PU4dPmjktVmeNFebtyPDUozU53ZHdCdTPcPzLxLowUjH1CZYJI9tqZEaQUB
QtIcpnFUBB18DNeXA+sOdk0+Qf+HL22EpHrxXZjU3bKtGhuwkSj3YewPNu5APBS+
72JA/uzbIjxVvuUT2Xzllztrg6dHKhIHdLn/hVKZV/agJWBSGULom5NAzK2CGCHa
Srgpz8ovuJRKR6HglXUCZEuyawi9RwEtbbB5RONYvl7Uhn88cD2GE9vXL/1JUlBc
HLM/g3wvLusVIK8BD3dx43usb+Fc2gTLr87o2GLMuRFFtMDnAjCrHC8OinsizJjP
qk5aMzHRcUnyp6rpoFlEpnNofRT7BEzpbk6RrBJPtlqoN+4wOhXP3qR2PY9PysWq
sK94fJLcYSZvweEOJGqlhzVCJHOe5kwHS0H4m72myU39JrBmujZ/TGEKYIM82FIk
6+D5Dbf0wApg38utW0XoRzlb2pM43Rs2K+gf+ihfNW7taAugjE1rmtC/CFxUP8Zn
F744rmnam2tU+cxPwr1jpo+nikVt9gxfaUu+DdMk580PjmAhGc55wNh5h4dQRaTM
6Um7nzHuXGOKOTbbQZWshbulCco++BCQluf259WgDNPTsATIguT2TyqUJOwXGg48
p74uV1lmC7s4bT2DnNh3rG+ytlEG6MVTOVOEf/LBxDuhfvcuaeB9SSvsRtr3JEAi
K4hXLZCCSjii91dncDblB4J1HWHxSsboQ8jzvb9ze3paa8Or2Ry985DmIECaKGEe
Ri3dM9LZQO42SQ2yd4SjSHtsMh/jyL6c5G8v25LL8RGpteYKkO5AxmIaEE7bJmld
WuMw9Gv/JqidLFohdessrnyHy6UDHAZ1ZbdXT8m/k1/LMsWv+rrDHJZibuocpthD
5eMsIbB/wyHok2ZMt+Rb/JAswSDtuBiSTH2lD8yOeWUNVDomNwXfSp4vKbckMlXk
hpZzuTJqquix1byFiue3J19R8IoohUeP2aLA46fhvpy128c9eO1YWY/BdVJ6fEqn
BYE7FCzSHgwPFylCA0gnQQGethWIsG4ytKKrsI9wCtrhe1OdzdIZn7D6ZmMd5C7S
dB0tL1YvVEKUJWeJ6XmmT9YMISF9MbZufaWRxp7rVdaQIwJsXWUAtlXG5ujQAyWH
qI6aBsLfYjk3R3WYkRYnqn4h/JgGievopg79QFE0/YnhdBo49YO2jgmQFihewgps
7Mw7o6Lb2Y/5vHO8CFu49D0fpNTeUjKPrx7vK3ECo0ZHCs0HG/Hds3d92+x/MifW
LVQthnTk38g+YwUl1uWaqNMMMSWD3iBs0foLU6wvlmxkeNS+iP45N2iKRrdfTs4W
PQnEVOMu52/7/teJLkKUkJIFztlR7/6u9J1W6PUnh9UaMrI9FfE0KJg0Mwl1g71F
/Ttry8eMfyB7nuJ+o7chpKtZKyAS5J8v1kR+GZRuAQ6M64lOtq9c1IiHWZEKUZYp
7ZRK7+tZ+GxeyXXC46zneJpn2eQB8PoHa7achYDtypmDkgaK78ewQHqeZ/5XOsF8
9uV8Go1mohzSDWmqz0luuibybIvoAQeJCaIUbrHA0+QeKRiis34H8ViUe1teBXnC
yXrl5gJV+TPYR3G81ZIOk6OH2MCfHJrRG0/MEtqyZ8RsRR+tp5idjeMdNNQLXAYG
rZd1NhKsmH6E3Uxep+YIS4DV63YtlfX6zOygzyyfjRhsqVP1uPoZ6D6iRxAT/aU9
I8eKsvA4YZCHjemGjYGPtZjNMC6fsdVV65QJERbPSSWTINsClq+nvWFg9C5ebhOd
eag8zuLVifpzEfRHL/Ts6HNOUqXcnj70LWZPg136bM4=
`protect END_PROTECTED
