`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
R29kRfOqdDw/V6yM916ClaAIY9L7FQOzV5JrXoui1F9W3X2GKhC4LZAkXIg1TZG7
25x0wn1HL6/UndZOmgx6uKlziGOZ4FtFBfJFa7i2asRdcME4LJ0TntY0wt4OJCxy
My4MXvf0ch55fqo2qwrKygGpiA3PMJSGdaIHGl+to7qpiqyOz1Vjb+dRHuNdDuZX
GKqUBqeu+WY1yV9UXHy9GpMau+i6Cb96kJpje1jUZ7M5TzcKGPQ0iUxz95mrxeX7
SzJOflmyq249YhyXZvqLJh1ZC2egUX5hNrbfHfoTQwaGbHLFZH4EHWKKvJxFvcKK
+OZ+Iwa3CWa+22x2Xs+Tg6pHQwxhybD5aMDYf6oVKvdVwgBrOiOy7soZygmJayIc
OxMsgqI/O7CRhFHST3F+eKLoeySssRQMf8ZnuyU31ndlvvhlpi0rf/CXBJTX5xUt
wvfkoUblWBbtXRAJrwIMDBbQft/uyutqdAyXkxw/qT+lyo87+Yc54phJ/VcYg//O
kq0pByf5JO7fXwWyvDOgaHvOlGYbYsqC+k7GP/TqLenNXKxv2U2dvWPdK6chijCc
Tga2YAjxvUpZbiXLksAJC67PPALU7kqAYBZBlHFhKnOlNivUi2vEKbIsxA4Joe3g
8psAohdH2ZxRn9VW0cG/SgZW1cxJwz3gppflkI36rpTiO4isKRmx7BUwfgjOI4n1
Om6+KRMnBJtiy+CzSjMaIkmEVDxHF5N5FO0W1LcQWyNvDmZ/CmpwWaQ8ikN8n3Wv
qpm+YJtZl4x1/gF+EOs/cGcW2LGXdjgw9jVmD345SDhiHkWuJaapfJIRZe5pE3ug
kvVHhJAZhf9XAupNFNI9cVN4RdfaawDfljuoN0GG89ngnaYrMnRk8HKRW0de7M4P
gIQIf7aUCpd6RPDoEnm/UNrwkgRDmeG8KNVhBWq1RgP+J0rzQbRem9LCLdlAcElO
LJeND9PZ6LCfGz5vaM5RQ3gWfb7dHZOqLN49Z06xqkV3mqxNDPqb9pcF/89bETEH
owtUI7L1fkD1YJxjWiEJJlSaJTjgbu9cnG4JYbXth2nvzC/eqP0tA5CMKlvIrGxK
g9490ZMlPOFK+aqiuoU6K/LYwfbQ19TdElCqypsQ2SiuetbDrQprTOGAnBSg4/cw
Uyr2JKeZKfJYmVIrEMaF/hJL42XdSY+KfOmM59C2T+M5Zk9Ud8Z8ebjKcVEnowqD
2ndwJF41c1sHafnooZootxQU/ifxfKArIZ5PwETnJDU=
`protect END_PROTECTED
