`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yBFBNi5+Gz9rRqzIbT8ee4WrNzg90PWb9ZnbgpOkoBEX1KKWed3MMWGDgOrgkHRQ
ZyiPnuMln3TcE+T6xZ4Sh6Mh3XlgFDGF+5dnuKPRE2omB46N9zrRVhUKLlQGEmbe
H4hChTff3iK9hokAIooordv0dFzvyl2mQg0vdBpo5d4j7kExtlF+ju4a2v9rFlqw
nIlrwc3+GIVXghSy4FGrxrLU2BeQ9wGLkSdFDl65g6VVgZgLsETt5WMHW8tQUlLy
LFQ/+tCUUGDjvNxfZ4NoWpsTnaJgYxiNPoYUmg9i8odXpHnbRkaSduC3xyS5boGJ
DIim9Ox0p9SZj6AmZKh6ae1AL4UCD14RKs3w0CMzIImrW01pOvA9MfhRt/Z9lKaX
PoUIx7Ymw81/CQjIQWWn1MyZ2el9RBZ/SQSsCpwh0/ayrfUTkcCvq7ln5y47JC4B
eeMsnV0uXo7wYGMsUTq+i8Ze3/wUaKwlXoR0QqVSMYrpyDywPb6Q83c++IJKzGyi
cXgcckwZm7FxUC2wDLiv4oQrS32bMO6APWaI9BDlRxymjJeLBbe5B9QkHSt9WVG0
YBqR8vLdZiNFI+Ry/OE7E2I962M24t9GnvZbjEtYlu9+pzOqwrTG80gGXwCCSdGd
OLre9YXPnsqVDvsa6Dfg3tNfbZF2k+rvoITcffhJrBu4qVynUO1eTfsrh7XPHmZG
h/a3hgBiru9Kl8vWMbJaTuctuKcxVzoHaEZOr+Hw9AamhZRGqB4qtEqb7ZXcvqOU
etQlvXrU7sY0ru5HZAap3Yoy8o3GxTSHwONAWUiw/fBuU17fu5rQKYjsL8lgpbVS
SnphjxiImBclh6UXqZH3PUvpPv/OQzWtHBAs02IhGj+xqin5+bPHweGsP9PmSFDd
`protect END_PROTECTED
