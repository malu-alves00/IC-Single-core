`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GSYA4hpQBrJiDAfjzPIqGnp2c7w1umd8B/Kur/8YCCXZ6m4162R8QqrIU/UgPch6
CDkNvrR3h504KRiTLCU26FjdoM+g2L6+FygEksRL8o1bPdzFegMLEKJLC+xTd1U2
kZ1EqoYFazsqDWJlheSKwgbPlMSAlRidIJYBIYaacLnrUj407ILUiaC2uK59t5ns
VGGzPB9IB/Vprf2LXjJJ5VrKqiwkhbZ1Nxw+KSSgMc+cnUy4Dhp2XjCX/C5FzXWB
Hc7l2LxQeBuPtrBLqEzNsNn1jE9KUSUPM5ed6LJP9yp09IzJC4U4UW2eVqAnvwve
C1zd+Es/GK34KaORSJPg6IxRvVMrXRI0xqBo1appRRTjvGTOVvb+z85TKDWmnhR+
DYRmuIRsZ09GEpLvMg6CNU2Rl+t/b4JfIF6nS1j7N0TeYJ6vtOJpcYd/sdO0QUq5
N7m+p+IAgcg9440u106rEcH+SxK33faHCnLA3fbywNP6aU1SBlrpswTfVFUexNVv
KrB3T5OrSYGqk9SA5kT8IA==
`protect END_PROTECTED
