`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
T7DWCzFxe2L/19pPGGC4aKfupZb3xlIiaFZeoV07omclwZKqC7ZbxZEx2uteaGaW
gLByYfNMdL7GzNe5/L5tsSOGzEYWuekBgYjl194d8hKGcTF6uOxstbcYZFHmsCo0
f6IxLABP6ArkQkLq7VQ2oCmLLGe1yLppbjByR3FywRrT4MhcVPl+ta7V2deL7BQR
F92IshEmLCVeMVOhOVmElCu9Qd6PqDaMAxhf9TGMqjAU4rSpruv9/znVhQbLXbQn
E+82SmOWx2zTESn2QjtF3e3tJMmcyzEDN8arUSRopptmTRtkhiEbLqIG19Z4isrY
sRTtCpmMr0R1NlaeYBcBMr3rdeE0nhrwOCV4mqZVT3Tp42zbAkh2nbx12pHLmhf5
60bwxanK9Q7t8kYj/l9/EtKp9JEVbmYPlLkbNZ537kgqS0D0dkQVbP9WTwqcQWuO
vCpifVWKfl6rXpURHorEa4hQfvWN3X0oztK6ZrRRRX+SoTtUeeF7E8m7t+cocvf7
g6HAbRv55Msn2yCF8ck0Y7dDOjWEYh/qG1ACG2JdrFUhBABQlOWxpWdkz+MtWocl
C6+bRxaHgaRShXsKnJf+MI5BrKXqVIL+Qcyk4H1RAXsc4F0qqN0JQhsddua5a5qP
ETXfcSB7PcUc60SIlFSZxqE+cYhixDxhrVFVGCPhIAh+ubQE9+/tpqCbNXzk2Oub
lnaEWvw0IacR3NnMAYpLhR9zxtzfyjj+g89cNYDdRZQLybaZEmtzntFDbpo9yiW0
RxaXMguGzY7sKBZ4GPN1Va8ZJmONSYp+FhhZE+kl3pY+Ty0Qgw70PxH3K0lRaZFY
M9Lrhzhx6gJVMxqgUksHsfLeWua2LLMm2oO89PWPqItQg6wDcfzM02jeb4sih7r9
ckboKElV9Yi95LBqQjR5UVKkabS+vsXlOl/OU33pUYhqAS2vL2FZ4Fv9SgEiAj9m
tov8sY2w9Atusvx5EU4SQVXNPIiysnyGAcHCJj+1+YNVNG9sRYiKOLqgm01PQlL5
ev9YLAbHe2pXHs9cFcEMyIO+rQGPyyWffu2u/uMiTS6BaKLkj/oqkOXh6jQG4TTj
FLVZkfoh88ydnPv6YmXl1KEYhA/+SjXjrt+WL4di+5+eWY6cM/akxLNch3Smnu1X
wymxLC1UJRfTd/SKsONCcR8YE+XINCZn+5e2tga855X69Hb9IcmPE0pX0Lh38GZW
jybKSZg7e/av9JeqE2B3jzcMwStblATynKbFpNB4BIjTiLXRzrU9TP1So4WaO1z+
DB7peklbEkSPVNFM9ohjIwwNlktD9Z+5I4tExC0c2Zuc7a+qBFtF5jRXxo2Dq9cU
nOVjeQen7zSz/q579aseXgxw9u8FI2GDvxkb+DhZmTHojkEW++UWfbedda64BpRL
oVY8j7PJfv0ACIjwh679YGZPEu8+nAnCncJMtQGfUmeL+vrTCXP/Zws8HcIpIMJc
JlsQzXmsseoRGJAqiXXfDjMInjrzD0W1KC3BH69zQSmbOtL7NLYi9FjwoQg6R5OI
gyTCAoLbgu0iGtiLR/NMX/4ixIn5Dw4f5VlT3CibPj8UnSZeauOP1L7p4Eej3GDs
pTaMSAPEgc9Ny1sx+4qhZyLHKyv7j1pBlwPOuyGy7M1PjfpIukx8RrWDSQEo6xMC
HXO+bQNlpYpn1kIBBcmb/eoq/HBQAF3Mf3sOSDWaY5ZMRfdkr+0ZWszM6u5uMu5Z
id1JaBlX9xgfsRWN7aYFvIeRtz8JnjkASIq73QR9QgDi/2hI1gviR9bbD1hzua18
KQXYSKJVJ/X12FeykCzBt4S9++j3mbBgD8UUOZMkMGkUOo71ioC0+uqaNQTudL/9
QlPTi7J+jLw+jVm/gaKD3hVo1gh9nK2OSrFbI3oTEtN2zC4ykMWPXZJwXj7h4JWN
SbuiZ77Y0QaajoW+fY67x6clQ9lGWQHlDTCXqPGAR7jJDVw0RQkWqVkzrvzHVVO5
3okB6iI15kY68+vzjXLejpp2/rqHofDwkikJ93RJo1p76+mLU7oKsMlzxKpKb1b4
E8KZOo8GTIFVlEmebtGAzliCJ16BvdvwiQIpqKMN3s4pPkTlJ3ObJfJU5wu8sBZ1
X7SZZH7kiq84zWGOYKPO4vGi1NDuseWsSN9Hmis4w7twLN1zN3B3oKgyGFocVAYJ
7tqpcaFqD+fmxZgpmo2h5Dnk4FxIeyDdBqpyVZ40hCS2hsPc7A3jK6MkSc/nSO6X
grl7Y5rTk9IfKcsoPzseJzxdoK9Bxt7K8/hpeEJGwXUv1WJD0s48y+dSqC6a7Yx0
MUl8Bm5YP3NPgGGgPFHF+Rp+v6r08LGS9pNwNUiNcmnSF4fOtHhWcx0HNHzoTv1l
krOZjetfXcf0Yo3bpSpJyvzRuQkcf93niPzJHrrTPAfT42vNAqlR0zgeMzmRuahh
`protect END_PROTECTED
