`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XcgygvM8mxyeONgzfzzelj/7QFCemnDSVuHTIF8W44S/fjVFz6/n87BppQEngpWy
02f3E+z5g7huWdy6zlkPwiHRnBgUwLnpTbuTQk9P20EzySjAG1wvqKqWkuFKD8u1
RjqEUKhbmxxOoKo1AZE4lWRxkuweuJY4Sd3Gq60YKCHU5LZ5sbvgxqtIZwmj2zRO
IHnvKZketcwznOOgdAUBuWDAu6Xt/fFiTJeSHNjXAP8egbA/59l4AK1kUDhCk/R9
tXIyznmX5ri2SDZNX/AvFD6Cv6cRDy/JzxbyunhwvDojSbfuCeymiab7D4T4zHi6
U7bV75Dy6tdsu/N/dwAa9VI4HfnpcP9seMUaV1mbZRYSiyk+vHi5qf43aAgukH3T
QBIDmaRqTwwGbO2S4kcQA6+YkO6rPA4PFUNXKaBX6QAc0RrAjs2FveozrHF1x9Gc
Sj6c2sP+NRwNO9p5EUesAw9w+coSnbJy7qpP3BtY0tnvhkW3sPCcCTNTiDma1Isc
IhKdcg3wNaV5mI5j+6pqpaOrANqFQcDlFz06v82SQUfQCyBhvuaUxmEq66kAQWme
XGO7VWKVCe47GMXX6zDxtlvKT9P4+ceqJsVWDZ5DwURY63x7i9h3IjaCMKTBc4Of
LI4hvxaTgxiGd7Nfgf9UbKL+I5SKrE+9SFloPoyDsSsJcJ7lvbZx1I+VyMtS4AaL
0aZ404t6vA8ATiJAQxGQmRPfdJnVtR/vc853G8JccJwDQAUois2phF/S6PO/1Ki5
w54mmjU0O7Ukn3yOdE/fzinyi6EJA+4s7xl7wMagq3hinmeZeGmBM1q6lK2H8gr3
DxP1e7mYBl8BEi60drFoyUsajdCeDQ2dRvY04qa389Qh+5vVO/47Yx/vZOb7XXpf
+aSUYal26AjR+nYfzRsOZ+3oxaRc9YSbcTu5VQ9wIW7RjLAHh8v7Oq96BGh4+Y0w
TzqbaoMHoUQF/TeekCRavfzKSlUWdYfa4ZArGM1SQmJV5zIwOZVsUWMo/3YgPbq6
1QJfGL+RsWwHygA/w1+Kbw5UMVWpFhmCyBcUhW93Tr0l6/WsRucgaLWnuYrcT2NV
7/sHA9Y4a52fFbZ56bEWjN4QaVOX0kGRO0TtLVxc6w4bbdP3WVCd1GewKm1mjaPv
IOVgURcxpLi8ZpAWtj+2J2JOvCVD8nvTNQnJMkmvHM4A0Fbm7G9hCd60BKLXy4Ve
8o8JW0zKLd7rCIQ982PiWDIN0Wumxl4G8PujIrfffRBufbjz/dmip/ksDA2HmgUV
Z3xwEKPkM4OFULuRrdwZ4tEnDJdbqqoaNwGwSe5NzTnIHv5sAz5V191fhe8R29ck
EqTaNwxfEqCXbXfyR+oh8ZPDCuSd56bpLPdqCAq462ifvOudo9aT4hiR1NYs6Nvl
u/ekOs0SIqrIQ1duasr2AglAB6M1Z9dE1zy8IDbvF/jpEhCZ0s0fUxcLfLjoQzVv
gKpQ4tdYqMYTWiMCGg/rLgskVYO+2WhvFNUapPJs7J3uDJpXa6OOusE/9YkaQ8NL
bnGFHtxT//TyicFyM5LvblDteJL9IGLMqbs3yXOWJqBoL+mI2dFAqdhNP0A2Axts
HYVdLDB2oE3qx4M67wTQ2QysQisfievesfqgPKPf8dthbo/6Q9iRohy+u83ysjNk
t9hxAVC0xvJc+V22l1Wn37e0uHKWHVy15croNM83MSOjCdEF3oTCNypkGACXSpWi
xdBn5MjYY0y1DT27Ntsa+PnNgP7wDz/5FlPX8e5JVXdXAR9Rfobqjmx7nHTFmvHp
KEel0REo2bv2CUTcNE1DLjn8Ngbz0LNUW/XelvG6mlSyIdj4raPta8AdWcDLBbms
4u5Qytn3GPBompJpp3Jpe2tFKdXIVIBcKZ028eguZrGML0UGhu0WGVo0KpzdwcFe
TDBtLKJI5BYyK8/OB4Ipcc6plVMaFuYKyAg3PCfb7WoPDLTSIccZwqIisThwE10Q
1MmOnUmo4B93GyTHtom12L/JBxxDxRo9exwLOTqVpf9JgYkVx/sWMCSPDcg4t3Cw
bOBUpMzYAkfU6elw+OPOoC5ercrMty4FFwISLYx4qccdVTQEXUZ5R+7WUznXV+MA
NVEzBEiyVKxrL+1++54NiOKs8TiPF8ukqKgcOGXqnfM0sqIRU/A+frSnfQD/NDs8
AgmUFDeK74Gm6kumLE7nt1fXdAHPJ+FkG04lL0hz3FSN0VNpo8YrSt/2ZwlcdLsN
5sAjymFg64peDjGeYZNhXzED6MAFY5KHGKqv3TaaLDqAr+Sc9SeK8AHG+A5lI/VQ
lQGQEg6EG03ZgS5ne4qReTbtfnG0BncaA16sklDagoaoHD6fz/Sg/sMFaJ1XcaCk
eWdds3QgE3hDeoY9N8epfSfW3GWLDWhEfzrSJ6S4NvChE/ZCiLmAlcAG1JMh0vaa
36Xaa2/iNSPz4ePaep6VJ0vb3m4j43rS4SerRuzSRc7LVFoHU1C+PMlHUO9Mhau6
ecDY1/BqlNZpTVbREOUIfWwkFFFbe8iulaZir6g2g+o9Tn0u5zVNPqGtKQftfsjo
y7RTCa2Y5o32Lrrx+ik/k58kCUgqUgRihVk4MFOk/yO9tOLFbT3sfQ5txdoZByYR
xxoiEXbXYWPbQRhuAsR25RX67TQMxatKzlvSXa2x5T1vGSxeMWCN8tYtutg2wKv3
POowM+SGyN/KCMHSWrAjGdEknwDn/6xU1qjlt5k1B06o+k3n+Y1kqUoL2yAzlQai
7JmDYC6ORyPY/Xg1BX/vCAaLb+YS0vv7f94zAa9KN4SJUv8AB22oPrlZcPxeA7o5
WhIrBzuiSQYZ5YCJ1axyrZTgr15Q8rSTtqafC3x4iIu50wprThvvsLFcXZ8I64Ch
yPFFU47ZxPuCCf0SennHOmMgdNcVrGecKmNrRseeVfQcfbjqM+TxId8rWDavmDQP
MOCGleObl/GoY2nLA+Ynd8Km6NsKpJ2qEI6JPNFTu7qs1SfZE6jbw725Pb5MYzRD
VJcsMHJRt0ZR19tSaNVwqPNFmlQg89tCPMBF9oYJbaWneyKrtlPipj4RS3YHWm1T
WBjsP7Jmk47cHD/fINzHeZtJbKMJzugNs+jC8wk+x5l9r4kAEXasSUsfRnVBvkPb
7bISle7Nd2xHk9sDb1YtDM0IStAFyFH49C+8Jrg4pn+YIh2ESD6FFc9XSdWWxQDr
AVrfM1Z7mjfIbKgb57L6d9Elf8FE4gzlR8lwOM23oZRRbeBmKhVVU2EGwhoAn9g+
9dnjKQECpKWJHh2E9fXebIS5fzc8RYo/qTbXLZAYl6zJu938eMIlUihEH+y9pMG+
gUvLxF48P1YEmc/sPWl9XKlQPAaVUAYRyb0cbqgQE3kayDWYjsF5x3XIDRUzrCjW
6dFAMfbtF4JI8uHy6LVHXgtqiAx5duWrBje9G/vqt9h7GrbAex5j56SEQIfyt/KU
LPaRw2Fj1286198Kkh7Kk4gULr9nO03S+1nEWrMobsyjKrSMWU+RQ1zP4VU2Vi1I
3mVFG8CnsT98Tgo/fBpq6mXfdRZxl2zctpnYqqW1gHgaoQStEKUdZ49BWGtCow7v
FK7RlQf39NdV6y/O4fDiLfSs64o5bAcNpwN9iUNebyH+qa4mx640pgV1x1KM9khj
xZ4/fGDlJ4eywSE4ipxIb/MQNItCKKipkNHKTcUzzXTL2ne7I6OU28H5TrfKLFS8
y0AlE6IdRZZCjHJBo6XXX0XYPnax0N3KHZmniaQ8M5EXYBNO0fqaUinqUrSjJEFr
XIqn2PN0JyY9he/KcLizLZET0IkVqK5Kei1yWFzDuuwyPr8XAL64Sf897nOemVS7
STUi/yEgI/SwtuDlQO/nBdrrtN4y+BE0z+qEe8H6oY243UcnWA4Lsu8QAgTBOaDo
s7f39GNvH51tGWjNb7yGSJGPliqqRTaveZeemLFZbYwDXvzQp3mBLRGGTPxkIyFu
kFy0pOLBhJQZy2VMvSGlZd+rX0s+JfO67fx+AlkbQVKtckNqk+lcnf9bEPbK/LJD
fMNhs2DjZowl3MkIZT7KZ47enIL0H6brVTHt0gQt8MTZfPP5Yeo+7BlRhHjXOJjL
uF/HfXkAHvDSlqMbclFpYBA8LAdN4ihKxB8x4w/VGLBHv4Laxw8muN1L1/o5sVlZ
HMA5cZOaRSXofjmoBiP6ZFtYR6bD49VIMZfeWJH0kXhRGSbBjatwHU//DsTiiyC7
epea8+tr7QZJ6Oy2fubYQ/CqLaDD/NqP43MT4HjjpvisBFeci18vIgBpsQAZaRVi
OfYVggiSgoLvSOCxBKuxHwNhQ6dVQWDdRcl7xXWZRwFqXFY1vFLJkdR+tEdAxLHC
ILfZA19KIfsFodflTdnl6lcer9a+1NRC7u9nOp9JJoYkQGf6AYIAkxgslyz0lczH
xke54A16Ct+OZBdl1C9YHAJsCOz29ChOhu/9aDaLIahSPJ2BD8+/SLWDKhBVKBAn
r/xrKCT1WYz64Ep6N2vm2olKnRHUtdDKKS0aWP957m4digXwiWsxrCvlyXMzDNno
zA3VeCn3/5PGmoOE1MSrpkjUZWu43MmIjAOzT0JmFp/sXsEe48s4y6GI/D/+9aKk
7LF5bzUqvbjqABPWS62fWxTfb3njJpci357KgRuHQIJQEklu3UdTzqwi4ubaqckN
spzGepwD9r7cE10jivI4bgQ9ddnzzIEm0l3D5NCT0MZgDjXG/kXgBObjggGAR/W7
ClxAC5kO9fG1uM6tz5TftHFUSJOrKgXsZu5U3EGNzDRrjFex4Bj4YOzfDFuzuaSd
bjVnWO3c61/qiUQmA75WCoPw1SkVKYNlGBpwHCMMkXTCn6OQREAb+7IMN5WFrxIT
sAXLGHWwlGQRGsiEp6DVCLqrbVAMlWKxRdu4fyN6TGr402WHrnxK9i6BmnrBV9RE
vc7CeUeT6n25fn+61TaN61hAKDmCOGfcbKVtC9azjHk1oF5PCH40aL3rChjv9LJ0
KkQIoRPzBG+qKIL8SY0iL3n6pkhW/33xT6ftdXM0KEGFKMtaZSUA6drxx/7uE77D
SB/i4CEJNb54txU87cwKU34fpYoO11UXJMRXB+s43QQkSNkmTpIzxHcMBRbNC17q
BSJ6K9eupodONSzzWm8WX6Z/jvTVhTLG2NKsjzMR8WcG43/07qtL0S/u1iiw8gmi
4lZCQJopKpJyMgiWkUYDn4EGMqZq0jrnO5NQhdMnqW/CfzXsIQjFP+88tX5QxfGw
6StWobfs9yqwmw/qQFz68okvQ4eEpkdMGkMyNqEh8f2oO2g6VfJQAa3iNgGaCAaC
IiHR87tZYWoFe9klKoHsKT9h2YNAnlcgpPM7IJsW2WSLOqN+WEf/lGsJkrGYJlc8
ECpimouu99egtkYi0ZCi8r6Md3RJzftuEBel/QjHwYii2uNiVb9BWH5Y7cUpOWCB
9j/ZbWAq1fMODf/E63oQrImgwahvq4CnnCrf4oaIEI0dNz6jkF3TItEFk+lkR+cY
lfz2GhoMsi8KT/4q0jyi6rmX9XuGb4F++8USf5ApzUPlmAaLw0889HMrgeEuYpGI
lXx/XJcVJLEgmzsWq/BUZSbyoz4Gf01TJFk2ihuQXnH3LvAOXGBlzbKCcPQQ6JDa
H7PwxILzhNsUaXmcYwxwi1TiRJziYZuLQA5obQBvP1XL77l4O6XGXVSS62TtLCcd
JuYIkCRWwlvEFWXMC/KzWRUKPZz0OLXEF5lBf/qo7MjWlrwhHQZOWUL3GpcAbBQI
87PKBeL6tPLlSyvbd+UcKun7PDF/iNnb6uCPDSLpptOLVHnbUQON1g6KymsK67SV
nFm9zpYZPW1O38vZyz0oIDPRaY9eO9awvyFUGSGen1YvMSsoTot/PQY2WeAbhrBN
xGVZlD3hXjh19S6C+dTZr8p7bW1u5qPB7Wp/RO/xFwcX8Q61Oh0fRc66Nu+rBmKf
ILq8RNawbiVFV8Hjz3DKBK1Ef/a/E0MS854m4LvCT57GRgyWY6Nyv547fRyCD9Ty
IrxEszOARmxkFQP6DN6+cHGgZMLEIoK7HpnFRVfcGHUzERjE8vF1xrguSw/cnHh4
+qURWSOAhzKzgc/n30PReH8tZD4+FkRKOvCSQ3N3BS+HIQ1Aio16wJ4Bs/0B3voQ
jNW5aGA2rM1OD4P0CkAigb+Pk+b8BvZZMowYq2Pymtutmkdx2Wp6tLpWubIMdgHo
SJrFml8umXnEsF+MvDM169LNZdDBbzJg4rTY69CiCgs8S4HRgXR1qjSOzMqqo4a0
pXLMMEw0NX0STXUcj+1isUqfVtUCqWqytLi52y+iF255avpkhHjB+lNAvaJRS/NI
aHpgXgdIWmrKmvbbyxfsTv2XTeQtWNlNkyIzqxR5V9SYcUWmLo/3iV3Fb82GbT7F
iVZn3IHEhF/0BiRxNwhyJPFK6D26Uw/Ak1nv5wMh6A/4pAWDOrfxNZKumdx/2Yem
DO/GOPQvMAsT6SE65Kv0dflImJN9U0HU0G6UMszIs/8BTnQ/dpttAUvh3B4vVd4v
tjj1BBWpJ4M8ytdMYNCWG9KUzfPqUwQK5kDjeUjVlLo0C5x85eClv9L6xXrnyHBY
Y/GWNU9v+S2czwNXwaMTvuf6wCQVS8xDvjMiSgO2WClH8rXZuFJNafJaDKfqd3+0
tpUhLag9D6sbAVsU/wcmdhNKKHzkmAtPnTYG5c9f8zFmggX9LqCC5A4cD0/KxI7A
/5Y9+v91tf+5mk2/LXJfNuSnVbeoSG1kZrO2KgpAEkbqsndTMm0ks1QsvvfHNLlE
JAxU0rb44Gr8dK2DyEAaXqGO9i1ngTl+T0B4aX/ObkPRXrZZZsq7UQLhpYsiYRKY
QgcucUzluq9jP6msMpadPC2LR567GyvzkhX8h6HYYVl9cEmQh/CCirDUz/9LptG4
GCpRIfg+Cbxkiq+LLJmrKkPEcuspuZrCcfX2gJl971KWYtGsQON3zaf2KV4N2+Pe
4FazBJiNQkNimBYhkTjIt9p48gpiPKFbKcO+0bpUAHSxtX6PoYXXjNnQHVY+c6q1
RagP0jhtdEoNVb6pCW4ef24o8KW75aDCJilcjhWhdrlxG7FoPwG/e56tcyyNSOIr
8Tp0VR7o5+0Fc39nuioRsrqBTrR/GvAclCeDcWY/NreYjwEbaWhuygmI+KYYSav3
YXlBMqGZ+3XAhbgtABK+A2GYYTlCmx0QmZ7gS8z0Wdf9PWh+W7kuokahZp6TMmzd
D8UIO5f2+KysgU0EYOn5rCSkcy7sjcJwWDKBiRHZCn/K82wSYCdXhu1UXXal8JvV
dLm04EjJ+sU+CD8ra8dW+19kbpRyfRIk4HbacnQ1qcv8SUMHe6sU6B8HFHhdRWQf
q2JC79Rlp5W0in9/cWtnXtsINjJ2UsAw0wxE7DEEoRKyZUGt1N8x/n/rPrsRgEW5
Ge/W0di2caFETJbl1KbWYLUKS5toBq143lzG7cBRsD3DL5lExY/YfGsPpO3Q/adZ
BjhY9g1DTsLWj1/0FJqBHy1qwYte4oOSEXwSnb1nEejKZ5jXkm8I3MFvx6PofJzN
a3SnZJSzMVTXbnuabRU+YUZwupZ9h42owOcbyo3+2Fkt9roh/Iwthq3ujuVbiPh0
EcJAjFy3e7igB21EoAJYjH6eZzulaZ2i2PbACQ8H7ltbcRa1Bqn04e5AdP0tpJf9
xRgyS7z5sHn8LCxtl3x0mq6XNcD8/ACvARKAAO/wSashCK7XOi4DAd89gHvHHV/y
e04QMVIVD1iiS/uSVFK0D5KBRYJDiqt0q1QMwSR9bt3UifhR6Jau3Q9sG34sFQBU
Tb2rhKMr2semjr+xnUb6wxOlSBOtoe7isP6zpSn+N22rgXd7pR6jyjrB0ZBk3MHU
lR/sGiFEfjUA1IHZtr4KaPLDmhNqr1NLDbmEDnUcbWNljjdrIaq8YuRp/rBhFtOA
RW1xqZzgLWds54uIeqYfQC8g9P3UAh/pj4BNpSAbf9hILFsgL7mpxNyJbgX+LtIQ
Lcqdie1sDBk7ERgGPzHXbBF+KCPK0GiYRFDLqYknl/TxE7ky3eUy5EO8GjI/LgpM
fwt5ABERFbKkXr/IndO68gmgKJRS9gjQ6ZisHGnBg5jBt9BdrIdarjzUh2Wcxc4a
kPkSqyO2QsQYoX6ac5W621o4dyjY29LT33jRrYLt5dg2W+8qL2BGFmdNK0+D8GU8
IJRboTnrH6WzuM7D3WYfZ74/Z5LS5QWBC8rsilu9wh4aCTrgi4K+msVKZvS/aQ15
soW97JIKgXrwJQ14mYL3NFHeW/Y3m3g+nyDAJOP73iEnHwVPWsbEx5TWbzWPoIY3
8lnTyi6V8VB2s9eombRyg1i6wAaWGyyzRiszSIPoYowDa96CMSFPiGBTUXtH17rh
C/XEbhKv7AMQhKjj7+xLrzoPqV+MKHMO1yBg2r5wFAUGqUSYfNxhk2Rp+0sH9xHx
JlrL29MCRCi4yB6jzwAFJ3WcCQtPytM1UORfjXCNveCPjUwkMAIDhohBGHFAaDkz
pfOX7lmYgpmJbecmoosqG7EVzGvVcNGM++/nX9vbvHP6oyeoE6COECcGK0B53623
E3ow9cSZgWzdbEB5veqe0TENJzn8lNdKLU2fZe0/WqYl8v5RSehwhQTXkSWjuVMg
te6xzNjJfm2cAkgyPsOEOgNHnB6TmQPD6PGFd1J4wnMzmLLZW9UWQUSwJlandjgm
WK5v5FGChP9hYNE+AI6Av2KG2vis8CIYF0BbfugTO+vymjepxV6zb0auazNFgzE9
UDtEo0UbEfcB+qZvGadMELzQa464ltNB3DqhmoG3WhI9YZU1p+XYozqqDfu4bo6w
mhkFOCXPfN23yDLew6XIc1lGzcfkulPcM6DpGy7uXzXqL7xTTNoQIeNGCHLbCcZH
C5IBa46UEEyW+yDQL3Fxr/R91lWLtdzePXYgrPr4nex26j+oHOg82T6BbW38C/O2
fnmT2Wg8XT8L4AT1NZjGXk03YlPP7+0m1xpXdABP/+xHkRIGZSJLD4mn+g5eBL/a
s4tWbC6SecoJKfNlLhBK2bKYEgRH2Iyt0P0Ga1qPdinj7qd8Q7gxhxCb0ROxdwkc
eeKqLV0d6YtBEWYaVMMSpGHsAIL3Cfn//mkwhmfQX/C8WgDfyAj0FZVi3G5kJm32
LCskmYwVIay5g0Rdx2lX2YTNv0Ts9t7/m1xig8qsaVOpc8XoaN9hQ+WdrZQ20Tpg
N5Dd3jrc4jGSqmH+C7kOSlwCiK29qaOfXe9GfJtVNilwAjReaeVe5zsWpyC5Evmv
sgx2nQkfjHjYArr/yFm0X0nHK/oV3Oyx5lL94/k/Rl2/vLQxkwhzf4hJetfq8l4l
vMzO1ko65b7PlbdZLnK3pMFtJDsjybpxHOUwb1caEZVEh54VusUh8zHHo8v0w3Z9
YZVjvQLqURWXOMvss6Dw5WFbUZliappbxIvREAnVmYIYqEsutZwynwXZEWES9OBC
Yo3VQQvYX9YuWSbND0wZmpM4NrLgnHQyt33dwt3fLRLI2HthJYDDzzwrubs3Vq4L
e2A+xyIHH37ZwW8u7Utkw69/Lf4ZdCkteztY5q8Mbs7OjPAbKn71AWyLptJtY8V4
NMRBT8rHunrHJUStqTzqJ6yPP78bVWNC1tG6PrjM+Eqzi4w781hqcKANGBAw5g8d
czO0Gx53rc3SITaUItEV9YuOd+RpMj4ibFo3QUG+jYKSZ1gmg863i9HhUGuM3cG8
5XLqG+RtJXVMpaXQ5zC2whiLajgbZIFTwpjG1i7QO48NHmromxC6pi4dS3lBnSxj
ySchXlgMRlrCBUN8HRqZ9FNdx43TUMS2DEzhQZqm+huFOH+dG7V6F5WUR8q4T+JQ
/Wg4HZNrbIGl7nF6dr3k12JrXPRUjeckNjYVxFW6tbLEgCLwF+p2/OsnFLTV0LHi
HbQ24UCUMLSfzGn27bvn0aGBav0n9nxnnySreofx1dGzNJFH/dA9I4EjtX0EPFzf
Z01BDP/aRej8Ixm+Z1EiPVMyZ4tkKX2OK17a5IeQYNVahzmGVUElnSOFz96bzY29
nAd9Rn6rQF29n5ESjGFYCCMAGq5eYkzrelzFZ46C5zFFmgTLhRVJLSCh5y5XJ/Om
E2hlrTlojtvxr9L6Nnh2Rk9aW5V/d37RXjAYGR/KrEVZwZwOCxX/5sCjFwwBdMVL
tdRjObdVZ7dTr/5MWeCv72ZbHBiEsekbM557aFLnr4J2HH2YtKQRon1kKK/q9RvL
TIm90x9TcDy65CAAMI4It2NQSkQD7Y5hm+qabOfYhVBVnBP7xImVY3Tvp59SMxjS
MgrMy40ztiy5rdZRqd7/rcKyn7PykUL90oaaqdMglR0T5rmxr+mJIobGDpfCSANs
wN/UPX4zq/s3Y9il1xmA+ml+alOPz1GkvsHdeqF/LQ2/Rb/NG50/ZigZMdm/jOJT
B9DCQZgLjA2Za0VYm2VoMQjEvs2r3ugqFuAB4VfAH5310O+3MUefQ1dIVkWeifTW
jPdUYLi3LL3moupdt1YepOJVVV34aiNdDWKtsow23+ekwC6hhnx0s08ti0v2GPBC
aiTjPEf/vM0nI8s3RBiXmXvzRiz3jQaXld/PIUxWfoWAgNdaaMcMxv7d1BPIprWx
5xtiNEKJCwo0Uv7l86vyABC7Tb/HkhzGUJ7XZCvJMaZ1gjrOiNHjMO75kQ6Fzh4U
Nz3YL6NdIUKBeIraEsl4VOrvWmtQs8DGnydqvts8NNP+8IXqRfJA9lCGrPU/Xqft
cwpwG6qNoe8c9W8xkwpIiul1v4DRMwD7gl/iutiews3zQ94S9wM9QStJDxnn9UMy
p0v+P0R9uzvbztFlrCqxsHw+C1lm18W0RNBRKPIPJJHf4nNO8anVTaXb0Xg9NksF
A9+YszyewGX42oJ8y6XRlLEPFFV6D5WlGMbWZGVV/e1agsDpmvpnle96YItbHO2I
5URz326g3rZIrkwndtU0/2X0B9bzni7O+Aw8W91bxxUUNwBAxN4Xrl+VSv6iAq7n
78KOM5KbjAAalYGLm02KUUBa1mq6n/kn27ZicZHflsJJUfiBPC+EtdVIWM66QEeW
/OGp4hxh6QnQ9ld3nI+GcpbMk7NjAr32iiSygD1/GH0pYYdgHQrXNGNl2VThVGPy
aJBTbBNL1MLTuA6Uok5n9EsqEF5JzPKqrIMTnmLSfBhmH/0ZQg/eZfoEpZ06YzqO
3pBM3uM7Ihe0SZ9IWxDbW3IwFaEJkgJng6KqSvKHIAT61QKOkGiHvuX7l3Syeb0G
A62uVcQOyGVKYjAeVUblKfCGFycF9GRR79xMbDG4Tixnt47f/Jiai2Nsez/iwARf
agsHTWxmDC8dxkOzAXKYbbXomYLOPTuArxwjTyNK3FIt1sSTx/r/E4UtB3eA9Wx2
UD7dT66rKQhE3DzqYrIEMRQLq5lN2BryB++H7qEpZcGadPWGm2EBgyA54F5RZsgS
8P1d0sVsCbxqoj7kV22fx6z3RQ5W2hl6O3ZGV0I0AY3A9tTaHpajzmIy1CK3Akcn
Mtm0JZlKANh5WcIawOp5FJHu9uZF9CikzbYveqaSUcIBntJIZRQpxs24W+GHEltH
AAqTHXj7YcLucxm4XWlLJNSQ2ghT8HjoTbuNIY32AbO2i1koHx8MS4IxpZi7MYbg
BuPEs7hwZFhttvLgvVsIMYCoDLB7XsxadJoDWtzrdY85ySrKsTpn6hM5HllC0b2+
E9ivsJh/nYaECuGoUGP804Wha7q8NgV2CxT6D4cs01zSmdVdZyLJD9hrJgdfNt/r
WcQEbHdvILStZ8HsushW+DwdMQXrBO+R+OX0EeecEVn3/nlmenx+tzj/YmiEll+u
A/DjC4527zUQy2nzULnINPXq8QiiR/jk0ro+xzuOg82m1N7nxvBODzu6GxmX10Qf
UO5Wk2iYN7gntxojgHCebkaYuhAOXCVLkncJW8APdzS3xi5WAVofeJPe6TTxCbPJ
PBaGwSSOnjJH6q7NGF+SnAKlbDY2hPcYx65qi9d/AS5mvhkilAL83x3UjBJrut/z
hdxczel9hJIaO1GaQqXeIYLoTS1ku/FpJPXDaDlLvgsJyxHjhxQ8g6J5t9d9gPyj
RW/Vz5s//MY4j/C0Wwki992hLUGVoQzurL9UDabg9R2Y1RPu6Tlk+HLyp/7HPGau
skXDHkXMTT4npNSbOmcfhRyUYk6VIN1dDk3FsLXu1VMhl7lh/36MTUYTjXPI51t2
WRJFXIU3bwWWBaeaJ87yP7bUqyQBIbFlzRJXUatx8YfSo203sPYMfSeHU6jYCDLL
4jQO/x3n3UFhTXvdW5ZXI7oiElhYHX/svEykJ2JLJasmcIzMvqoBblMYe+aJmWCJ
vn564hRveolFN++lcz2CukblXH7Gcjp747vR9dOHtGLnkyZAwA45AbNFrjl6ztV5
yRxfsXr8gul+LtoR9GA21BTIDo79xDOjUAUuGSUdC/u9/cI6FbhIsmLNQyHeKiU8
LwyWq6awlyRkBtZ50WEH+H679+Jt2bjJVwu/ZHzgVpirFU4m9y2PWGq9UyKvGjh4
yX9Q6deEIszVTUBiaSmyOrKmIz0iMtqRl+neseucj0uPB1WhMrrm19a4OqhoaNEi
2TRDmsAaWbiMbsPfahDj2E8vnONW5vOOLGLWSDAg71WXvWCooVLpotkENxjVfJUu
Fvamdp5n4kbmsrqd6x/CL+th4mei3XV+2llxDOLvgksH/LQLh3VgNsCMWYpJ2so2
fyJQCPC5/sAIw+botR7JNZhUvLjJGEWD/Zo5AjKWu8MByXAppV4nk24wDeGrpLhQ
CmCu7i5QAdfSJ+RgBfLEjgCkOtOQDUlkAmY0SN284J7wpcuyaxj8uJk9kQQkUxqt
UwCpClxvOAwaL8/qaGbWo7P05XCxs1wng11oR4yCCwv+aTJfISgiFBU0f5RO4Uz9
n0FNmNU2Ka2Ymmm7QA/31Emm/jfo2iZ2YpMzJyd6nLpNGf64Oey5tBlWzE15YRqj
HUNNS2koinX4rhTIf/ZLuVIcalpNXNuV/YU3TKj3Ew31EwwS9nnx+8qKIIbYekZI
I4RFXTGSH+Zbmn5AKtFVE99yo6jLaCBYb0Sve/74WPNyAz+FmCMnTFxt6i05QrX0
noldtngv/xyRNuxypSPtPlj0FAJ58ZE/aGE0/Ra0e00MfHjxWywMxcj8vToqDZ5I
VssqJyDi7Xq/HEErfHfKFzi0GmmzBwBfhIEICD7gKtOieoxoJHRwGEwAaLtJELuN
J/Bag7rR4NjZuR214nMb+ZC5tnJNdevHRLdqtR9vLFZc19blu9mQg56um+TbtG+6
wVPv3RckP16s7WEpS+AC3Hs6FSFVk72Tr8Rb47yJQQI0iQsyhXhivXXYx0UC2BqV
kq4+Wh3pKsaVbSiaC/yp86awd7lFvFJ8JcXLSWvmdcA1fpBMU846CpVV2AFi3YpA
o12WIUUSUAbFDNdNqRkEoy8gn9kSg8InzW7dXVxR337uV0fk5kM34mtZtR31kddC
Tca6+Z3hzYfWS/Ac+vHI0C/dH7yOrJ1gKd6s3Osf99TqX9u0F68+6EKZgck3CA40
4cZK7kzfBkt9pRccY5dM7WQS9Nmit1NhfYY8xYy8ScgO3yQMienJOzsIN9f9K3qB
e6zKGkAbbbZWaGBQnXd9k3ZBwUIEC1JHYxnvT7XA7isWI/3lUbPKiSnBGu1sle0F
Y8zec0pjhVUa6uEyI0R0Gs/8UzpVXGEutrAalnRb6U5ynF86J6FSJi/xol16/bpl
qDBRPE1QYifVfYfP7l08w87SpkG/QWQfQO2CMFPGHBoVxIwzCrqy52Il49BYioKt
UzVFaaWaTE6c00Vl4Y+JLEtELT/qf2mOq2GS7CEFt1DaDddmo4EyavM6iURBpZ9H
FPhMDS3ulpHTjYck1jOpYAttsa7jc922GHtbNCspP47JiCWEEIEp3RXyucOeYdOI
rUU7xi8Is38Ak458zjYsrbIugb02P5JDXp6tytAwz/bxeQKupqyQLDqfbgsGrQZQ
KSF/mNuMLLPrGKbXDj13E4+yC7LlUzBH8n4WFrwsuUj6FPHigOfjB4tgvQH1gPVr
ao9OVesTLUA+aG3fyl0hwPxOxr2DhggPK49n7iyvDrexiukAz3xoF+Qwif4e5FcV
iqxorC10LNkQ3/EGYW3t6IdpHeRv1xiv7SrZgt9St76libO3Ap0AmzTZORokiuPS
cYbmbj6zS8qU52bYrUoUv3Tus8ew/r+VEExmEut+EwCPGPvB508lrLE8ewnxMYE3
qfGdyyayFXGu5FD0YT45Hjy7j1L3G+Ek4Kfjwxg8P7gOMCuRU2oPhcad1/o7yBRl
SLV4MtPCrdVOWjW3ystrYu2O8VJ7EaVBNFvqkk2e7BG7+4VDPoskJf66Pm52/0X9
8cGxcD8ee0kcQHDEZyJFJY96hCcbGtj9mAaJJi+obCWK7g2dVIOR2Exq8YiRuaFy
6tZ0Jg8UJnOlZQRq/gwD/uYbU4JyFXcT3asC4+ZUtke4RGsGJrtb7bpK2y8OQ8gW
if4kErUVv7tN3ZvhDhJPL96YS3SrEjOUsrxfgwxB/x86AgfiFr8xNJvk8Ujescw4
JXFm36NzeEa1CJMVEPQeliJ4lrIdoSmMY5qost86dgbYb60GNZ5vBt/bRv42Cirs
ZefYVGoDkJzav4aiUzzsP7dEFY/PA5xPi63IdU5AmajMJohbYopXEhdKSRyGM7gm
ZuknDEiuiv7iovIg0xjlPlD6tFn6vHDPj/a5QtSCvYTqE9g2KySN1OnXGDOU/wrh
D0cBvchpxp6LW8dMW+L4IzpXcoKlIKQJU3NvfsnQzGWjHWb8CafXjJJMwcyWp47v
Sn0rFcq/sYQpKuTV7gMfCSFjDBlR79aW/QmBT3nXJe9nRIOYbrQ5daH+YBayoYzX
SSfIzHoVooOom2UPqsoslAuR8EOg6El0E9ODeUMy9NwUoAJG2T4G7baD39FuS6wy
r2eneFdJ5ImSh0aHt2i+yL6YEyZ3rBok1GJ9yzSdkwqFlLWOEVLsS0CN+XVVyBKk
Ra1nQzFFrj+/z5B0W6zSCrQzJA2EnytovqZsHVBBla5C6FjmDbRzePHJwp5mU1Eq
NpaM7p6YPXfZI1IZxav7CR9swi9uKWZXdddIlEM1GOYkpcbXZVlMn3lua0L7eY+r
/bvuuOiCdyvjrskVEUAK+N1PpqnykRixwFe6lDN3IY8iEhogclEfJWd6jSloDwpA
p+hwbtwIOlEOUFH1FZG18QVWfDv+jWY7GMNY5yleSTE4jc+Y7rfVvQ3BfMkqKp4m
sw0n96Wp5aXfIZmRsCgFZ3h+4r2/hYio9jRoWzoEDHzY3C6SSIOWuSPz1QT8pEhh
UiBSql7tM2KD5ycIspPiK2pxXj3ZOrcu8X5LFSnWApWRnAfuvKdpP3qKSVquRzcO
IjMXO46jNkKzs7VZxswvuqh/6JWvNJx8086KPXRaq5RvrNgKTJ9r8mni/K0gFwy+
8Cp7lnXrXg7cFJUrVvIJOgCC5uf3qjmjJESYHKjcKv4+aL+PDjURQJoT3GCsOS6C
NdCSQ+QrDIHqzYjyhEzmmc7zWUIRezo1MlFMbz3xXZ/dicGg7njd4EgKbmZiY4ce
Ffb/E2M6ChS2MLkjQ80Bu2QPCqDmyC22NL2EJM90kC6ZdQqg6Mtt9gl+LiFTnflq
T/Sq2FEMmagQhlw9s/ZOirBScGlD6XCsFewOwnhzKfWqjq9f1T+2vT7uxomPkfAD
vwRM+AlCHMft97CRO3hzRY472dvOsZG5PTeXiiErtT8ObkrBbfECvWnxHj91deQx
+m46LwM+rF+jed3W4FKcMSfzMDC+moXxztDU+Ynv7Lj9lbzNyThWA70d6hu5K41A
5wEjYIYDuypn/onYDhJrKyR/LDvbeeoO+HsWYIoqMBLa1J695BtwZ9Pcgp6AP7sY
0+vfBLGGRRsig7HqWrdBTB0I9u9traAmr8yK5H1dCc4I4u24ncYsl0Nh/jFd3jCS
PRPdK80a1sS8Xd0OkI+Izq0YVF1fKd0LE5l2R13eW30BbBDLU8j98vb/lmD4AJNy
sHOM4DWAasOmNbSrAcN1q7KMhgnKiFEqAm7cwq070MaLs5ITuXWo7hTBGYPtpFpA
diQL6Suym7OeW8XIPBI5CK9Ya3Bxec+LkaPCNZBItVJnw63HMdZBcHBXFO5gsVlP
XURyooQLT6RQXmm1WktYiQm4LAZmu3SJtuzXNFbuUupeNUOU66OwI4ZHF1Jft3nr
h4W9C1pT0XDviZKU5b00OEXRAIe8kM2f7eBWl4XF8LjsdHVX/+g34H3HuC21KUWL
x7MsZIo9RFsTlpLGDXl1EIwdEyTf1zjIAPqIQZqBX1ZlF5t1K1A52hn9FGk9zKf4
RzLz2WflEJ1dDQTdgYaA09svzo0Z4H8m0aesFAJlirGr6qGG7+LE/cNsK1/6l68Q
Ys1vR1ldBaIxkYD3F9tG4p5lkGZyAO8IjvAD59AiYUHGksC5DW8iOfl1AHDihGxI
OOntaAuqIBs8IvzJXfsvm0guFMiglwWDTvM6jm4P49MG59zoHb69RHZodHlhCOq9
/E0JN7+w5+ZmSYoGl0ozdLryeDuGWEXWiyyrPR6VLpUcJANZ3rX288Vod9VGKykM
1dZbYtpYI/+mU/uJSL1Gse9PmK/6in+yl8Oo7FZJ8RORQYo9gltHUA/H8ySNLWoA
4exQp/LL4V15Fs9VCJyy3xjhgw5ngj8TsDLJ7diKk/QNZA/9kl4F/bFbvgw3A0Rk
TbEiWdw+XZyXzOCpB7YC0cQPGPEHdZaXcbFT153CNLVQPmFh3T3NJF+aqMGlO6Wi
qUgPrQ7pm9GEMzgK4cO0NKhEZHjo6HCKmfe57ZrWYQvWBsR+i+bcY5ZXnoJsicz4
EveXWxJmMg/+PGgItyPtEfNnLOXAEArsWL4JsIBy0oHhnwR4YOCsf+VVocG6szQS
Yo1gHGAxC97o6Tentv298q9AUO8Khney8qc/bGwTBhcEEYRqMnR/zwXmLzkp+7zZ
1WEvcpWHsQeaXxII1hb+ieczn5iazfU/30WZvfDUCC8cLJ0ir/KRGBr4H2YW4DXL
7d/xl5HJE6sfg8MaI6W8n/EWYladLo/s0z5g70snii9+cZMhLwRGT8harC+1tnAE
S7vGU3oYNTnjONQ3tAM4FBz2hJnZy2pNL4W7cECZJ9Jd0/U3jJ+53YarZQGoyWQv
qT88uFnVHTOm289l+oxZD2sxUN7wRC91qzHjdNP2+YJ10YGeU6GuNU1DtlZgASDp
RATNIwELgcCEXrwRJj73HmQHyQHB2H+VeLnhgugHGanQeWaa6VpG3zA5zB9HreYw
nOyTlR46Fnj/zHu6O9Xqhb0WzG1WsdKY/on3etdVjksdrgLd51c7tjQrIe/w3uPF
cAjc00MyVSUS/tFv3J2J7ODz11IGSz7l5yiw0fiK7pgcRdOv1QBJ015gD0auMZzZ
sTKiltxVABv2ILb+34sR9Q5Dk133TXqUZFAfU14Xx6+aQuo9IJ1ctNCvhXDAOjFY
fLGqaNR5vHMDd0hrEWaRZWrdj3Djs+rIJFIjkQ40kFf3eOZh0vzWXxehz+sBZLJ2
y2fKqQLxlKT9d5HoLtalPOOOs4Q/ry56EN+roDnDJtZAZfmkpmezGBX95RQ0HYTz
SQX6lHkV8Xs+KNUL2Dq/cFuXzNY+9HunLJQX4BaZPSrZWMH99D+do8psYbjrfk0Z
Z23Yc5A/yITo+wTIHmbORPLmdYjh5PpLckKa8PWpzAOtBgmCRpv1ssgFlj3/s2Vr
W/wYYA+NxaLmHVKQksm+0pzccnR3m/K8Cl3b+dFhAN9oaI3q/6YRbbI0H1rBp4HG
WySkLUsZSyf0ClAFyRSgktHMES2Hm4Mo3Dxx9PezORTR4xBhvFchOmzQ3gf4Ftsj
fpsLwFcyA3yP2+/4VP+/Ly+mAC9TYDgCWb03kLgylchyw0Wpwtyj1Yd3Aqi04p+R
OobehQ5tjm1pkgLK49PAtySc5gQIJJk/azVyD2Ws5sDC8ZN1BoplDJ/CR2SOb/gc
QBaGhpU1ZqPCdNh8qNznXxBwcVKhb9XJNyi19xTuWZsH9UNDFAaE7rrPUm21nMEw
9qfXckFnL7J47RrAEi1uO48gkNa64JIKo78a+ukMTuPNw7qtUYAbR60ZntoduIrB
x+cp5s3M8y7q1L03PZ3Tw6NEbnqBy6sPvScJtdppw0mJO1QvKVGomHkyAiSjsXjh
bOrMXlJ/dRqvKrbqoReLImbjckrCKspZ54g+sqrqgm6CKuMTjaT5JDugKl4geqa4
agAQcazEr4GLwOEZPKJNV3gBU2vsCZTHNNHrZ0r1EZ43Fk1/prLLMY27IqLy3yF9
zqPRKWRXY8OwvszUKe8a5Rd770FGG6dutruA1u0CnF5/hY5W9XBq7L6crkcARzWE
Hw0pboKvWDRgFvrCmhwXak275zuesNAauT/+BbPu/oIKvzdbMUABU7Pj5G0WuSth
QK0AjitoKpahxbkHYX92Rt5egfNz+WsZx2QgpLYYPJWToE616FZamVNU4yB/19s2
nj8x7svH3I1tN911EWew6rrqltbzda1W8UGeIphqTsPGHW3VRgCO17tGtNGVOiup
qrepUvaVoHR4qBnSagOSN3qFHvbNPSPwto19thRtXWT1G51M/ZaW8hzFxcrYCeC9
5GZYnT/YsEYq8t8i1hv4onj6uSP7m0F3N4XKN4jTCsxCfwZ7ISiS9tmSl2hH/tCH
18lYCDD/cZhqn6uQmFZJGA1NgtgwqI16W/BbqsCp4l2oG3CSUcuO3mudWH9FLhhg
oIqxWjN3f9Ib9V7B+rNDkZBFA9JxaAlmPWJ9AfQx1+gszObqgqHuNkFHOXn0k1bM
dx09LRsS1fZ5MAtD907ebFnWdW+slyDIAF+bNxWRCPcWj4S0mcYK/PQ13uJrBFkf
stv/WyDPqsJwTTaqVYnoZQhSapd3bIVyx9TshZry+wuc57ncty0bTCfDiL1luEAk
ZHUTF2pXiAGWwrk1i3bAFxzOPXZJyOU0BUfSp6xuzCKXq8tSC8yh2WJMvHNoyx1K
BboA8fael6nnN/gWfgPTGei99k2YXTmME5fwFAWeAJyuYPOe/w1X+wZ/XQp42KvS
CLj08aEgxypjb2CxkLwvSOz5sreYeEr4+6c5RjcykImu49ggVqq63uuYL9zDff1u
Mzjp44kKkNNgl/njEjwCef50l20lGLSvBHZc1gS45K04CZzyc7BPKZ+lMRcXnwZ3
nZ/UDfRkvKARPYQFMtKMkPTqr96qpi2mn3qYdOEp0R82JsOrywwM+OI647e0XsAp
ZyxFXF3M1sW901qduLu5qHIWZGrQOXSkIVqiEBtCZx9FkVvvT3p7q4SEuF6AKEfm
Q9PGgbYz7jCFiLTqxJ4ZrZEkQPDOmi75TiKisuXWwd9PKf1jHN65Uzc0ziNsgE2Y
FVvnuahFO9Oa0MtKoYl8cON7UlV1jlRJnUZRu5ncW5f4ZhhzAZuL0JcI/Tudn4xZ
lVVZdMsd87t0rauOmqw0D/drBn3nNl6QrfZxifhoiOMXrnsEqgEft5fvRo8eZz0A
T19Jb5JZPEAHsQ2NhkjikY7OoC9htVvWiOsa3oS+pcQ2S2rTPIuBlEkspqgKjyLA
yCK87/EIyw8OG/AZZcA5n6+c5b/3D+oN7DFnQ8L0C1ylb+HD2ZRl23elym5ISTOy
L2wQO+Tum4IYBEkd5p0V+CUHg83h7hd+gBhPwOJAbP/ha0gI/Ypx5Lw/JmzBxqCa
Pn3fUWN7NItXrFlhFE0hw1MPEKv8s0ypAnVB2CtBja8IukoOsH+OcluSqeAdODyE
ETXvSIIGozrpbFZNumOui5fWgwvAtC16xmwjRO80PUWf2lh1rFG/58RrkCbdnQMc
F3/pep3pI4Qa7GFCgLg/VvoFZ2+sha6zwG5TlnmSBL70ph5dIKh8QxJebsXss0FQ
6YZGAHQHhrOrGR46NnBryCD4pxJPXHqIVtaZkGWfffgGy/6OKiGF1nzhfvmZA1Ge
BFf/75H1u6V3zxwUPn1A3ZcYTQZf3cjgooxom9EQrHGvxrCCkYzNjyUJ2/3KwslZ
VwYcJ5RWrkV7deTN9wsjKCK/8WyxMfP3tDpwx6cSZYV1X/h3k9745JFluqn3AZsW
7UNsuRxc7MniisdT2c2peCldS1V8Gyo8Kdk1gjsyM2P2ouV1NTd2u3+kRvxRep4Y
w2Fwk3r0MruQY5fD2rdGjvedaEkJuYenQXFCl3Sh55SR3SvBp3XIeJ29sU3vYnS6
wyb9mj41urtcTWxOtierFjL+QSfXyd7010YtjedrhXLQjxvORQsdypSmOfZ2a3B0
Q9/3aECb7tWS0XAXuLVRJGY9kEXKSpeV0E1xrJpDIyHuQeIXDyEfZa1CdTOmjggk
qCc55E5dbbhkRwVmDc+JQqTICG1shHYI1xCIyrsB24b8zyPf90SOvzZ35eR/aXcW
toCKb1RcgFC6aESQlFqN4Ef8zm+YFwLyLBoCShHojuwxaetiJ3uEQx0X7IrEbB24
GrL8VjIbJrYO7BuO0Qs2dc7HDtZGAmpjO5THvuRlygWejUyGybvL8qZmLTzBaOUR
Ps0kejsnpDM8zS7xtAHM4cV0GjkbnYCqez+fmzEkQzpsG+g8eDm6R4OS013/lLmV
KJUmtb2YnCVpj5WS+Avv1vEC9P51GbUd39NgyqSy7mav0BvkO3B0JNr/haBM0y1x
VvqQvakMHDSxyyO9+6TPXbK6JJKZTAgS/b+lM3GmSUZLYAV0FuAX7JzFTyTC6iOD
EDP24gMUT57rP7+2U6yo4MHguhusMxpcQ9+gP+o5H3UgL18bpJOGk2bvcc1qMJMW
o48WdFWYYd5WM1XwIfZLH7TNti7v55+g+7LcZ1KQTrmDbCZFmF2mlqtDJEBtWoZU
gFiEEkdR9aUEplOKOIZJ98lpBKx/NB6UjgDszL680ows1hnlXiKywMrAwq83Oym8
IfPqvUGpR8H1CMMoR9Q89cUZ5HtrRCoCl3A1LfimEOjzZrCBOXrU4GrbehDSkFwX
m43msan7kAj4PylG9qbjF+RYn48lWh2q03AnlzSWhhtXGh7mu6xwlts2zAb9NBJG
nLNczmUG3ieeGRbDoR1JWjdH9Nxm1+mQKHqoeQp/uU+XFDY+4JxJhAGnoxj49EH6
1dT5V41Awm79GreG44jYlb4XrWq5xE6oJSBmUzSO2U/whjm7pGBIJQM4R75YjXRl
RLCi8Mp3TZ7Q84wro/s5zwRNZ2WNDovhx3XzljdEw3xADs1r7k6qydiPQ6Xm8Lg/
EWQfDxr4lXLPeM48EjwXPjst//8TdDcZrJTNpY/LxMjyNrjaYSFuM22KYpd7c02n
0XT/hbHV1DVmfdIkZybxq5rxUR4QKNr6aHh2R2Nb0GTDm0dvZjAQ0mqQdanVtu9Q
3UykGAkOQty8p1fS4LOSVCJbaHepZWuO09G6yzH2xJAcxvlgcZSoz1pCoBZUPj0h
UpyivspPTsiLL4bdXkV9hug6sRJv5Z97acSSxk+PUAN59rJrL4OgQtJriRSVWW4c
nqfLPbQCCuONibxaZry39y286No9EpZBGLLqPVDFlnaZcQ1RjG7JJcyCkgVLW9Fi
PlFBVP+raRigRz496odwq15Q3HMuh6uXdkVyBpgeON/FtZ3SKR89oN8lt2r98Nm3
USf1w8zfKdb9Wk4Q5SOLMCSEdCy4lY6yexSru1QXKN0Hd6+NU3eoOrqrt4tTMc/1
vPTagaAjq3snKV4+5vD8GoEHUbbMQ8DRMXNoG+5ivXlIpmepRHZwGLp9pa+KgRzZ
ZLJw6Wm6sBxJq5mMaRZ/EcBKQMiRAezIELSy32s/jPnRckC9+R+Pd65XDylCpz8/
5+n8WUlJRUpW5c6Qu4hUtzkR+XBJW4H2EMP9vHjfdp8VPQci/w4eiBMP2vNWH6LW
V9XQRs5b9d6zt1PVcjOs9jWFcpQUcJVierHj+lkYitV8fpNAzGowR08tnXrgs+A1
6WJT6YDz09qm62QgPzaYMGegy9d2KpS2UO8qhX/80q8ZVyb6QSXhty+jdSNJ0HOo
h8nmkHpKa0GQlPkDNo6WotwYnSTcJWT5sARxvmszjrshcwhJ0GtF5FxZBHuoclgs
Rxrf39hhzC4Bqcqvkx8BinFSyhGV9VrOgfoS1wv+LqezlwaJhRfINw9fLKzoRswh
MqYIdn2O1hI+IGE0PpQ67jQd/W2kdGxpmT0d8b5FRMD1D51GSm4MAPgk0JlknvvN
7VLqVjImW7Qw+iBD2mzF3Hzmd6+hXnwBODSvqk4C+CKyoIDhP8sS11leEfHT8Rq+
x0V1e2Qa/Yp7LUg5+e95Uy3gGmgACimBkdwOu42Rx8uMYJemgWidd7hxB7sCZuJe
N2Dzlwo2U2u/jNFJQGRrWqSrq4a3bBLMmuATO0P1kz4Eif4izd9GIA/sCVF1Iyx0
byy8VFS2Y6wO76cFs4DSvCO+7mqWWAf0Q8v7vOmm6SZXdvQcBVTxEqKGIM6XPYTX
RiiOXdYmmRXl38zs1cRugTVy5neqVTLK8V8gC87c4LxZ3PRuuUtE5qtnwe/q84ID
XQEvXRR5OhRgqLdZCnwuR05vhTUNuHo+SrdMHNvSqK8qwy7F5c5p+U46JN0NbLVV
LCsMtMZIEY6TqzVs0br57Pg8SM3Cc5gxBUBX9ijKxV9RjQXPD0zuDpr36+fHSzeJ
1NEh7QGizOiEg50eiiTTJd9XtHyffMVNVI4EhLLFIkkPL9w7EIv7GfGD63pugDB8
OPgvESZrVA4I5U5EXm1tRFBZZVc4HKKBci/CeYPNATIm9EL1/MVxABXpXfJYLEMV
w9Dh2Ch5U0jvXR9ZoYO1h0BBfPIAeEXjHJf4ftll7jUSVE2RzkEA0Rt19dwU0xKM
lr3lOinNLLhsmr8O5NqPfFGJr8sQ4pAiJau0Xb+Ncog3PT8oDcslSmvkFsHFSe7y
M8qNwD1lSjF2WNRygNWC3qEK0wmd9PWxT35MD0d/DoCPpf3VzYi+NGni+5apB1KC
iCPgjrWm9wXqXHbeyA1FEgq3EXgs+N74pHE20y+0OkBzRq7l4bub3sq+1/99qkIc
LeM0bpFaTAag6oaI8keTGLZvc5aRDmmu2uX7WkDwb0QDGkQCTdNk3EyGS6W0as07
T2EKji1U4gs6I2SfKiw3PApEQy8lHa4lGaDp0fTOZJmXzfeI8Z4U1EyS8gU+2crn
BrecZBlHH5DOVvQe8Jx6svKTZVd3QtQJ0yYYZ/GrpBHl0kuJbmzwVDo8OoYIZusw
WU4e0kbKrN367Vr5pdAXMC8fYV/wLRxtGP5jBU91EponEuQz2UVseZCAmu0XA/6U
dcqB6+OlQw2pyuINL5USUJMhZhoXq9Upssoj60kBfo919a6YCjUyUkAFFuz8nFND
NnCk0+u/fMEuLWRHAVls/EQ9mzIy8i04UkwPpGAzXssn/SqYLLVkI75t7uNBeKgr
rtaShL0BTktxWZVK80YPT/dL8qiMZzMsv9nzwF1YXeqxxUE5WdjZu5d5egu9v6ZX
rAyAn+X1VXwKh7zVJhHLyFz3PIkynN4aM7VMIP+hrZVhlekBWU+F0lbpuRaN4iXY
nEyuy/WTRgl11BRr0ynd6denNxghdFsy+PI5BufnjgrHZP/kYRe5k6IcIihVw/d0
zanUbB7sgQb2r2r0zxJ3CZq8wUGc+59cCf1ZmxX0h5as4dEbGEzoWbP8gYBg87zI
u2B1IHISN7cOxqEyDwwavNEdniBWVLr/s+XBF8j4KbUGVmWd61KihtB+4FHx9bBd
VhVfyvont6/waHKlLTJjczdVDbbrTAvz8npFC/dwZaHmGcfQVOiPnYsSPTpmzv0i
fJkIMmnC1sKQ4Y0xDUfj/HuX6AWFSbmQLCVjniearn6wUdIoql80WDA87OK41l4c
v65UfCYMgvcS9v8UGLUcxgHCBRxrH5XS8fQabP3rNhB93Pp7v1jOqAP+7S6nHkqt
MdWIItuk4xvFya1oMdmLhcDoIwYRFKyejdF45ody6efdjpfiaprrSIQOFdycxknv
2O9shjWvd0gN0LZupacsp6cjhLeGocXlE94MDgt0KoaKnqcw5h+R5Qd2VxOM6grN
5FSeRB/+4zZtT0GqrL+/8b6LdUB1gLEPFoTcVW/1mo6d78Rop6CCSwReA/o2GcWA
BJ9kO3cmzNX+KuDtPgR//0TYahKYUCN1/4NFPZkHZmSVwaQDRfPNN7c8tn4Yod7+
eJ2cW/25BtJW3p/mHipTrfGnWauq6CpXzNFMnfOp/IxD1Jy6GiHdfAm70PhtJU4Q
64xJKgyWHvoo50Zhh0ZUudzEKmIL3DZukKrCvbWkzDmo/F53ilZYJMXcUHViJ6qu
D7kBS7yq9tXqtfSuqvtbMtCfsYsrMRWpVsJ2CvSXOL9+Mji9301o7dCEFWr5dS9I
IU5IJkS944/0sjSewHzqnGCVldBg2RFtkYl+QPHHIxAFI4YbDMYi+q7qOY2xJs5D
RXpkOph+3GNiSrUY3x8bYqbms6GSEg8JAmLKWuTLRBXaVNha9UjZlf8GaAxNikJK
ji+zl1rQJCEOwQE8bs2CXHXoTZUxLIJy0Kg87QDdGvs8DTPYd2wXJ7Vrk9knlZmB
3xrUEYSiWq7493gXrwRd5fRUBFncsHsw2q3m5ahiXw2gN278ayvFkQ4YmREJMAqo
c4H+qeJvzt4GnaGK02F8F16nQ4XpGQyF4NS+TsKIJLP3+KmRW4j7BoO9EbCOFcqg
vUGOXElXo5qXPm5h/N2ekuzjtprb7XzjSVPxTiFw7sBiLmW2ThxNaSFRzZWKBXlo
rjDAcaLKO6ZdwoRs+VJUZkSk1iY8hnXR+GoEz1yCrDK/St6aFv3BZde7jxVMArNm
10QxuSRDSnWKwwogoSufZQ0ZPFAz4uiLlQyeDWFXoMu+o3+tW10NFClkGAUkIlFf
aaE+2mIKcE0Zzo6BS5ZmaQqJiqV4fvXtP/dWzudM11Fhc4IXblt//IMQ2IE1p7ve
/vb50Rn51upeW1tTbrBdYhNBvBhYCp+mBaZ9RemwyLFQ/Ybb1XUrHREyPONTdIZj
GBCPjFkqqpuGBQ57F6GS9NGzRYcMzbMEguGjHfBpLFumjgAdlgAupabsnpEY8j3z
44Jh/er770JIP366Tm0HbAyD9PA9wdmwO9L5USkwcdmNc2HcZiIscvAaOxVNx9v8
kuQ0b5Ph+yfzFVGEkC87y85kFcbhrxku/rf293pi5JlKhjmFr/GVHWR9jFpBznhD
Bqe8RMPnYbOtVA4eLHtA4CeMC7vb2YQCQoIM1ThJP4NrWqK9USl+MX1AvR8++1mK
v+N4mgoGBjyKJppyYr4jpzvung9Iq8mX9Bx9AcmiJJLyjuv+BMXnmqQPvWgTEhkU
Rx+5F/l/7xZTnB6RZx+EEEu+ZglAwDPycOFSRsWx6iv0EiIKmU3B2NChP+uo0iAY
fWzDmbDG5NiCtsklYr3Zwqy2NIZhiYKVX5yvAog1vo6kD2JFvecDbPbwPe8n0IMR
/x2nSUzGmfB3atbxiwXt63BgNoIivtWmQV4A0HxTcLJGZuLJoCiDk4XrVhz3+ukQ
q4YH3qOc8E7nJUMnF20YJQWARdJO8RzUMPGGPZihLobCYWoWz2CTi1cV3KYYhw6U
01U2Qn732KfuoxpEUiEy2QZVkXhPc+7f3OtQOg1FyxRNk7Rw7Mah0E8GNgasdIeL
M6j+dGZcK3FTwt765nzPF1zaqvKBtd0bxHpRTnUgqKZgtsU11Ju/GX4Ya9Sc4tWU
7+k0Ix2HN/BpGPLFQTaqyX6QToYEPUEvS1OeDChoiKMvl3l2y1DHBjimY/hBN3Io
gYNgsl6pYcmn2aGy9qwpkDeDhGIUYLsVXAH/bIAeWao1Z0+oQGjGfDGauuzyMRMQ
NL5uwMp0TLvbj74KpGpnC7pokdIOL8Kvj4UKRwqmpL9Mdfs/PaWTOrKCeUS9I4Ns
AxtfJcQdXP4UFY3ny4FLk1iFpQ2MF0Jw2fEQHXnsn3qrgCepo6J4wDyUjuwGUtER
HwNjHPuHqdRZGEYMAuCKh/ibrooEvuSVPTlXQqoRvW+oRJhy9iMqKdxxxxYtxzUZ
K3cARBJGKnU6wHm+7x4li4XigkuQOzay48zQM7xZ6ZU/xHzvVq4dgaOkoQjEbHbP
6j8K/PBojKr750HxTN4mRHvbu0DujlsJjLwdyjkap10V9pMVC+F8dpYeq5n+moSJ
VgGLYVmHaqGx+JmsAWqJcpcgyEx24XYP04JFlK6sJE+2d6Wc7JhOV7br5KbU1Le3
HhWTDts2oDB9AwQ2ulCPJ3ykpu4tt8wkmaaGzJFg3ideCMVIrynLXAt0yGX4CR16
LgiNGiF8EScYW5yPkyMcqtxGGwBr5G92UHz8kSSFCn5L1X6L6puf3gIabzOkfKpw
myvyyS7b0DBsZ3zfO4fK7rYrvb/KyRNhroF/+H4ZKnk5+MRrU81DKVGn9XBhYlE1
5xcynLAxDCF9jc237WNVlZt9THQ88WLIXxUAYF2AiKVSiANxlegViTRqYqL5qR+e
ycVc2htKC8t53SXA6yl/jkVruxkWFHesWrRc6duFpGidvXGrt1M5Ly3DHqNrPhhe
1F3upJesi3wIFuNv0i7NMEC/miLZZIegRsLFOxL5t7/XU+Mx86V1Ir5VRNgF12DQ
G55AwgFVXLhVEIx9l9bYQ9733t+T5CckiyPImLhhwibBhNShhoK2M/0OP1caSSYo
A3rrpOlZrDT2J+uWKa8+NCscS+rC0F/KPHrKuciSJJQgLiWqMgheGBxnjpb1nIL3
deJ/yVMrl8Fy51Wh4bWIU0/tFMlPzaIfwwS+RXmD69WpG9sNLrMBYqiUYEYnN0Ye
SV5Fff6YSfqbNg432nX7IwNxirretEw7CbLqJiJVRxw7bG9puv8e/Qj+0U+brlOy
JZSTHmOr0ztklvRHvFa9bQt+RN/sIFz2mKPfxBVGUlESeq1W1WNZLk4OrAVI0iiv
WYDQTEWpN3seuJS1Rwoji4Eyn8QObyxRSoSRmzcoJubUQMnR4cOZWF0OGXF2oQ8q
RJKRYQogEN8alB1Bq77Mim/QWkyhnc5hqlJr3n8RHN0IQ7cBLZr0kqdniA2Tx/BN
X9Irxd187Ybg4lkDC8ZyIMrCmZA0tZv8mKYNgI9BfEHUTwBT1qHqyx9rfwXg8skK
qEEqzSXkNWBpIeTilbJs1efOL/l2KSCW86ON95QR8+OYGE+nNRdvaSH5K4DrR3ac
pR/zqZ31ID1FGb78ESbOltdK/vJPoCs+Bz1KUc4NokVwzebRnDEA7TBqIOKAGTGI
9pjrhGRMgx9rhMip+Xg3fd5EOFMryD/vmekjwEFtXDBOUeBpmWWRle9Y1udfaEUb
KyjSVgn9x0vOtWEKh+pcfNI2rNXm8t6musIXpAiN11uStBKF9RWZ2QXIhzLTB58N
xY6XjePcVCZNJfIOPeN8SutUbWfoYIMRVBG7jHQKI9cXDXikurulRldFbze5o5Lk
gyIqZ5aEqTd+ZA0CTzrfSCuJ2+mcR5Nl7Wtr0she1n2eZBt4tkJY2i3O43lrsXY+
BS+JtkjC2ImEk1xroqA+3Zm/srIaNnMaxiABSJHEcWjA+iIpEspPEpESKBHsu5gx
oG5tnwyXsJ0EA+oWqJlqicjkik/4nICEsSRlfYnFyaR8MrfzCd4IN5amTBNIzM3J
MnOYmwUSFcUvoEMVfBiNYEA0DKXXflUmNz+BBxAN0czt4lq2aLP2T2ssxcTCuRTO
mCoMedud8ZQoyTzArdBytWbYbA6PQWpUSk/2BA2rxzT93yhQYX/7nfS+uTf7q7KU
znpCsu7hdR3boK6dkO5d7HYya5EkzRWMFwincWhcS9a05+uqI90Babt9AJDm2aZH
3Vawhems3phiCN/vH7ygVO6ucYnnJImHbyFE4ZWNDtwovjvxohSHjGhW86DkpmHw
WHJoS9vXhKcSYtStNAVtJP4aZIZa8VZJ6NTmSFgsuSyMs/kSejmjPy5lUe66Gpx4
+MHLNxx+8wc4tquBSoo022viFsUj6HSNiRQttDtFyPd6k9KuCntC2avq4Dkc7uGV
E5xlgsRhtuwZlmhbCGOLIKeun09F8rTJs+Y8LPLo90DCwgPVuEWZSq9iLdwTOi6N
eUu4hgeQks18PzECP57IujAgDWEifFvodNM/WVZ/tKWUx8ef1tiyDPbJsIvZK7bi
Y/K2NWTEWsTKrc5LRMX1FPjNC6iJ9brBWlji/fUDq7bk2paVUO0ULyvgXzmljFn3
lFpHOkc6OWjy3OAX0XhY0BtY7Jqhk+H5Lqm0qG0WiUKMRLcu3VDs2lSc43NdZKxP
wa5PgQUbB0gQ0GRihb1xddFT85Qy5CusXMckc5z/r8QWYkxOVfTUxq8csOlU02+g
w0uef/OrguhhHUxufrKZBjvkMGAGZokg3niQ6XyUm6m0cPkxOGXnYRW2gURBPM9D
6XORIM5QBZ5O2z4RUrhiUyCUNSHISski5AdGISr1b9++7tqbu2yLj1dAEkPhYxhz
RX1jRTp1Fge5j8dxvcAXWW5IMLyfxbAVQFE4xSGyQbjNhYlSUlMG7Ogvlpab2nKD
0GNRAoG+TSzjykXPcxK3NFpaamtJvQrt7R/ULxWOL9pK0GHYmfTe29eQHDcFlZDw
pMOlRw6fj6ZgKBkWrlA3C3s5XXs/VfIOt1abxWKjxYXVXDtZjmaqo80WScqRjos4
u5KyP67u0kkoEq8cPjstX7EWwlF3/ZDwCrriF6g0Mk5yyLfY4AdIdI1cKTtaeRBy
pwLzDmd8wM1SLDqi649FYu5EvbdPgYMfrXAO3g/o490lpaAppyUX/CS2UZB+oQnq
ezvXsQDl4j8edsshXqCRC4f68InlELXoYClpxnml8PuDcBixR+MV2ttFRdPt8/ym
YFTMRAPaV3ZcO9LLUQGuhP4xagc7c8Az9a1gZ26z5+cOkiOlMyG0qIlXK5/PNlhJ
G7VqoNS8ZFZ/vEi0pEbvgW4z6KU+yaGMxyJboOCwmPunUWypSBBrKys+5lM5En14
9G/7crGSH3h0PDu6iG7fjsPLBE+rZxkC1U6YJy0+20DXNmFahzKcWmu54YN08Q13
uIbq9tm7qIZ2BFa2bKwzAKQ77Ehr22Mik3agMMRWRUZOFmM/Wq2m42oZL48XwG/o
W5MUAUTq2ATtmEAIjJXP/k3bfxRKuFqtSCiUGu/o8h6kJzQke9H9UYqpOJYYI6NY
7yjXZKOizt38fRmIcJrTbuMllFUsxKmDNa5fqcV8gltzpNmiSfkxB4xYSWiRJ738
CsEuID6iWWXZ5pOE8pGsLJDjJgsU57cr275hzk2Nn/FEHkBP4Zy4hqBJ6NfHubWI
X8193XNGVAWHPInySwZD6yTJ56QFu6LT3gTC1Q1MwJFjSev6lmV1aC5C454e1VT2
1xuyTppPiXxC/PpIn2Q3dRO4rEStLD2Fm73x9W9PyagxYIUzEjD9WHRlXjRUej4z
nnxq5Y+r6w3+Xy4tlvt8pX981HHqhmHiqnK3CdgVBfbXHEtOetOcRKUKkBjFHn6w
3S+zGkfZIRTMTAzKuptYRUDp3ynlQ6d49CeKCTcJw1k9N0yer6h+NJMFai8BxSOQ
EzlHcY9qYifjfHyZdMlwQ42iAk0Q6Vc3whuJjIC1nwMZVCdlDxdN1bkjHphJahoq
HiIj1SD8l2rt8hRDlp5w3j1jiq/pAgv81sz62dLrFLDQmQzuy5XEGjHuT+WHM0ZH
YwFZ+SyHKNkI1xUAu9Julu3tAPixKeQQv5HKfhyIsAV0Zsl394i0Knqm8WfVZCHV
5D5YUUOs3rP3VhYYv7C9Jadu8uQFVsXJB1YWy1qR2e/HhczK7o5XVdIiRByGCjA5
WMrViycf4lbRZhv74vpaVtIkgTZSM11eXUxOhWynAYwb/0PLG1u5rj3eQVb2lbjr
23fDoRdevyddN8F5p5dkMLPdgaDiA2rLblUf67AuppR9h7J/I3OTZhncHj+UOidp
ECYEDjp156E29dEVVugHp54ho5ICO+bMWudSMBYhv6B7odfppNtIalmwYp4/zAFE
pEvf0U9sMB0G9vUgIaLXLCu80BKCvW+SoV/HklJtk8ys7FqiQknT/1VG766D/NbB
T92MvP8RuoXVdohl/MD8c2zSFTWoCmBxFYJpgp1Ea3jYozvMUmf7J1YeO2XKSzuM
GWV2atKh56mN7YSbtLEW+g+ZSTVhRWhSwR64Nw5w6mLlZLbcfHBXZZvKgaGZmEth
CzMxGAXK6zm0AOxRQoS5GqSGqUYNZLjKEWznHGb2Zdf5akyhFn1Nz8MpmAxqzjRp
BZX8etU+IWEnTh2J/bNVcKdPB+pDnGYsnsppt2NoF14URr0axlNVDuVn2aeitBhn
0IEwcZaNhtzpZ+K42XhLxusvBiDerk7Fq7+0+5ZMGzPXticVcGqSEM8uSvZ4A4Bt
rdPFcFFXpIrkNLvUlkkDDZL9r/YQwDc1YflF64m8QzYNOjGUDulVvlLvBUj1dG59
T7emUlQzaH5GiiL5jKjqeEPDxin/N2r/mimawN0Ct/yjVbEDCPta6ERf5+WiK7jL
bfmDuacgZ82A3mzh6dbAQLFcQ8r9j/+PKSt4Zm0UyPUehvgh/bj4XxhTiy1WxOVm
cwlG2EVAwl2jZMXyzsi/BUuAhngsAnSNdeNpnj61WfOLPTuiSS2vfFpPidSbplk6
wpiokwtJnTHlxPToOoQHRInbars4VnIgsyS71m9SPladQUEOdN+AF9+fXmydnA+M
yNSh224GmYWWj4aXRscZEd79d7q51XICDRr39aAFMXaKN3pNng7yWwz2v4AAXgc8
5tbc5yx5HOjbbp82GJfYlq1LrH6C0BpP+El8Dw3kmNFvILKY8NN9+PGInFvrNAUg
tmRZWl0SLYfQtrQSJsEu0YcrsIGS0N3zRgEymlYcoZIcAMwp+doAIzgnA4frr8yx
8MnsFUTkJ5Tzf2cSQYRqjj1hnywa+qBUhjfA27R2ZHeikujyqXIskNg5CmFq7zH8
yhrv2Szuyd/Is7khWpjoTmpJcq8lSi5kD6HmRZ/BZf9AsJY9CR36p1jiVujkP+8o
jLCxbsGwo1T9G5n6kp3IvwllQXTTdeNDHBnQi1r3HzptINRowGohiaQVjaWCKSpM
BNC3wW/v8QAKCz2aUSe2C555qQ8HCEKzunxcH4+MxTLIU8X5xYztrQg82JExcX4/
2EO5Hd+w9H9gerdiVMCYQAOgnVrBPMpd3j3wUdmhFVPALcQXlhZ6UJoshU5NXlug
199ECaltNiJJVOELzEF1OHNcsg5+JFIb5fLhpGGv8nvZTbXBsyjlhXfVdl57A022
Fq7t8Ei/CtmP4FhZSsuUMKinU91nDl5Zi8alWrZVShsGjxa42DsK49+L7qT5UxaC
QNDUnfW0uLh4qitAjGysfSbbLZ0KPL673rKnCuF9eMScg2K8nQFLd7wEnx+WnB6u
K4gE5Ga3zoWejANSsRTOfwZOrJRDrT6W/hPFA21XUwaemW9hCVczgvEgHlS14Ooe
IMvbDbY/1XBRY7IlLhes1qcKdtx09EYnH0arW+aqX6JmSi5mhDL+ipwGqQQvDAU8
aBHtRHx02E2SF9ZlDWVlHCqJRU1UrveGkGfgu/FrueX0gZX1krJMsfQvUaI9NGap
G1Y4Qm1gLfqtZDESGkavzvX4C6peekiLlOUAZ37FboXlBtoSKXmolfpdq9uIL7jv
JTGzi7KY4e5FisFMa2JG+HT0qvk1uGHUgV1GHF1aqgUoHJLsePopcBK5Tr1s32Gr
d+l972/TmioHZMur6Zn7rbuwXB7Zl5EjzJ54Qd8lFXkjyfU7ok/4bEjj0m8xk823
Acvd+bUOko+wTYOKaXFzaayDP3J5cgcCbKJ9dxAUVgrAuqc2jTKQLDT9HejQ1eyd
0Qjl3p1XwHbKLvlIV6rlmuxq98YKhV5G2Zhq5dlzkG1wqq8NbdsAtfu4iYv2NiZ+
53Lzy3qXOFiEqIu+RhNdx46gx3qGlynsPHlmuZHEJvz9/7+FhV0CSyrl+3Zq/310
2KnFVEAgtLQGijvV/USQHifGNOuFBblWV7s5wrEF2zAkG6EpnrliopsW5uL5yXGz
+p9o1KObxr/SF5PuQlv52jnpMgA5HQd2AObvbG0tD3RXxfAa+jBuZbZBLORTwvs5
CndGYBBeBSNU7oEGShW7mjG1T3r50Tae6SxiEiAgh9IvSYP4BMsp15f3PhL9jP6D
xCZJlrSN4FzkV4JWW1GXd+NPWNS+sIxbyR2dCL5Q6zw9K+osWoLomTbyVt//WQW3
CbG2uTNkiJMpSf4Z/YcGO+1FANn6kXEg643iFIWrDYskFvcFSH+Ja7QGERHRy14b
ZOC1TfB/OSoe9JgPNHCt4fm7przhncsLu4bjyWgn+S47SG5tp+e7nL5wtQBrXEHf
fFa0cI0Gmv3sBZCWgJULrNnCAnMWTNccdA6DQfw/JyKXQQQQZHT9EsulXhdklmos
udz5G/bXFjuZhb++Fc0V6XQoqr8pGAZBOoIwhTWl6pyk/bs94hKssSEk2Vgy2cbn
sBSfTuEBYvDEQRzfNfca+lnG0wOiqwgbw3OC9jWjdWWmQ1Ak49/ZB0MwDZ7wDm3R
e832mbYUXjfm5ll0OPpx4Vif535OOVuVRHV2KTOhpKvDmr5zErl3TzFPKRo70hRt
lo/QlZXzIFb3kZD8QqSb6Dq/VMlosJBL5R851ufC6IXhTA0lFlbFLs8WkHdfJ4UZ
T/uixSoOh7QSwu0A/4LwxpWu6Gj2Lv9ZnfzjB5hdO1X3+feahyi7/nDph1+cHK27
26eFRYRlcEd3VSDvbWhZbcH7m4D2Rm/XdaufGMP4MTu761jharPL9pIf3dGC4M6n
sXKUMNwVVjxUUTBJpR7n20QplwiNJWkQzHG3jG8pDY4LW2nQBQbdAhSC6UdMhDYX
kHtLUA/qlt+zkMIrM2dYoiPhUbPKCXEZax/KBbe6Hc4eSyllrf22Wy0gk+/ysiy9
avPMlKokCs0+DcqnHpELJeF0pyPxzyc0Fgl/VmUVUxFVz7CqYdoIn5uBLw+7ls9O
YdNNhy2PifcVbuhUeIi+tDn7B1NVG4mbeRzkQSMIuFpZkGvo+zUGQGobmHwllFG4
wItX3fcfdU6/x1ZHkfTkkzVXH5h+USa/LAjzkBoMh3rHxiJmXrJhH8BwXI1Yppvh
zm6YAd5FD49phCTNIwqHIl39673P2REn4Sdhhs7SJjhNergwRZm17s4jlYZv2Bba
WEDXtnO0VtxGBys0q88b/mShZ5c0ivjdqGRlkh07TMhyVByyozSHIPB45qIkggpu
IxWeYNGmCvMhmMd9GmgkVD2vO2CW71oeJFldJsPBc24T6sJhp3srplks+go0YShX
Bh7bMLk1G7KSVcRgR2z5X4YLbItWWd1IsWqzyx1uU55GpvFagyeAnsYnDuKsgEnu
pAtpYcLNIKHxPEev+cvUchyVu8oRQx7JNocG+lK+GpCRroZquw+gixQrQ6/yTAOt
cyyHjFgrzfpHK7GTyEuYYHnNZg8lSVXJzjlaTojnzuVSOC8CJOk9J5uDJo5R2mkR
MIsNJpXg/NSvpcdcJGNg+FNve0NyEaljhXJAxUnZ7madfMiACHel8qS2onwzI8KC
t+Oj+trwstARcxYFXlaDkXJ6eQSBIsUPTXzeH5E2kLbY18/63UZDXgMiJDua3s61
e4HYdY2WrOuQdFvA1VinAyqWSHmQh2tX2VQv8CbljZTy8AHtdncAAJ54Y2G8+aPL
SkpB9aMbupB1Tjc7fsdZWtVJJKNv4aeaiQUcUt8WZTwB3XPpej0Q7u9JdVXayAIw
BlhML7YqNkPyASPsY/8aMJKMYvF458rdMjzDXmBQn5ldjhLOIyIBYpfLOSS3+v6M
d2VRfZnDffUveZkEd7NstBW809YUNDgwgQ/P/EYpJrptub5KH87TYJedxOgFCnYp
rvrcE82AsG6ZJvmuZMzULAF1WjOVPY6NXiAEEatu4ilLTX9TP3K/WUf0z7MDBbMi
lZFaw6ca0YQVf1On25MaeD6icq7E0VQ8S3onR+l1kNRKuN3AoVp5gs2FQq0UHosM
0IgDazM6sAJPUP38olXbSLutE8dDP8GmEZZhDrjbdsdSdGMtvi1w3A8rwFBleGi2
qRte0ciDq1Y2z74Jh4nTqYFHzkDa37dFK5KfpLOH55VDSD5QAgmxhsoYKDACQIMv
6zTDnYYYumW1i10BLBB4jvFmLSfZv9MeSrW9SuWcJ7D6proNkPQlCXjci3Cn3OZA
abzLm5nJWJUtZnBi0O3S3LVzuqDrqE21nSqI76bRXakDzP8SAmQGwWPwb39g3i6T
QfzHUYoBodI3d2CC+P6t38FdCXx+l86B5vg4ecBs9hZ0133tVUuwUer1eJbCe+9o
Ni0+b9fZpQviN+5DaZ+HAKFRmAaWxEQNsoRA9YtyJOYQK42cLuaBJQJ0ZPT0z05X
6upOYVph0T5fnAHKF9TnfD47gRl3PpGtztjw8pmZ8l1RoqI7nV/IskWPIa9ZPcru
1uOomyGEJ60wMMX8IXWvSuqYLIFQb4bHHGRPoD1XeiCiXGR98hRsbullk1zrjree
ScrrEmTjXxrJUb1+7V8excLX4ulxfDCvwheQN4EYqh8SVZa9qwAgHgq8gV2x70XY
rV5cmSdwXengNBrrd5PiSpVKLQkNHNaFysyKBwjqf0+6yyrywG+RxNy0hCoZRVei
YxFdPPxXuxBTq/b5cNv6Nnd7YjN9rk6chQT/mUoiaUTLX8yZfU78bkNimMcykCHx
iZOd3S8oJLsGZaz96ALGTsMrwTmTr/zsxnlz7zgGftgPv6aBjI1u7FKr0eRPFNaG
FC1c+7ALgzJwZwwyMf13CgNt5sOAWRSkfT7IUkZnmDq8NN2XxqP9QJEkkifHgBiR
1qnzHvwI/R9fMmOgEJFUW0ZfG6tMl8coTa7PUHb3tSJ+eQd7maCyE99KTULUsX7m
DuXBQ7Pe7DoLK6YqATbDIo1ZiLtGpoRmsOFDCTxq659OBlAOPFGEO2lrFM+5MPkg
zVQ1IzQdIP+3GdIa2qT3zRd4RZifjZmooCyyzXxzSjKaEklTo9HnW5CxkbRvcnHk
UVdH9DfBnxCyIdDwObtFPqApm3SiTz+aw433DosWHg6EhCXq25DAn1tbyABb/lEs
T6UQ49NuYT5+YLkwnw5hT/AnQNrm2lOUdz2dnTKRRvXZYiD6+h18OJH5p27gXURT
Iwq69YuAKN+Sro3xUL2twOXqp3TwqxKykUOI4dh0b0HlPe+QthwVioVI2l8pBPd+
AfDDH6DhzJFszKH6YvMpAqhRUQBdOGTw7xjvnluqrOtp4/H+6o7cIwM3Y9Nu3mxw
puyD9PYpTGL1P81jFANQzGlqsvZLHXZltAEe5sito5AMuaP2eGpnjIMf4xgAqIZ6
eOVAYTBAm+9yZ5ee1rJYwVR9c7m7od812QmWSgBuEZgOexPHQrkU+BP/o+KcdaV/
clIGDR/dVgBmG+/XnsseRilEKOnpyutvla1qpVGDC/gi6T6GrBQ0FoqhQt8J9tyh
y7wLt6Zhv61YcIWGyyUVE5GX6VCrgXauzs7MggBH8I9Evz3A2lM0aMapuIwjWejd
v/0FTMcU+Xhx8/EUQmsY8uBhqEYopps809gx0Y2l9KRUZ+Guz90/ifEA78dVMtI/
6mrD3NOWgy5xT7zNhj3oXkWIPDJt1NQ3NnBhVBlBzOCncYKfayFo/aZNxPguUm9k
ql1t0dwdsUT4Pa+q1HHu3m9sHB/SmFWPbKLlcb43d6rkCsVLiz99D3Lxi3s+Hz43
pstIQFbAJBgTnmb7RRZ3Jh3vokY+/ScGuHM/bqPV/rzoys+Zcwjj7loFZmOdy7zS
th2cs/9MDFGZhpWPNxz1/5FTlZBq+CfZiJmk6hMw9FJRATNn/OtTGAcA3+lY95nD
4EhWUbHkxoBy+nFT4bn+wbk+OwqF9G7B0YmvCT5XtcG2aw7IjXjG/JY9HpXBnOmu
+NScomVQtms2h18WHAC00TBu8YMKd5BD2/yS94lugF3WhIrk0+HJRDMPLEnpCyh1
/iWcLGlSuJB14lGh4P91/P8zp327etU3eWeNZ+YfBiiJyY+4HRkeL4McC8gTKUmD
L17ZXgQSQXHpFVVDhTK3TJ/iamBBsAKhltgY2GyGr7qLdMISWOhqr8eXHN0a+Pk1
5S2aHdJOp6H+psvJ8LggkfjPdE38+s9FXRCY3x3DcLUNa0qKVeIQcEmSjwSl/W+u
XWxKQS+qLhxWayaxMU/7D+BwPOA3bTpuOLTFgS19nijUP0xtHYDB7zadfCRzUxSD
QbwCBfTcaacNGqM+bLYmHFs2NiUiM4fYJnqWzNj0dPT7JBHnq+No1wUVJETYuiQ7
LtnV583qPnvYo7TqpDHZaGFARSNTxWQorsBMiencjgKC8gWWBRXTaxTfBO/ANfES
SX2ajf5uJysZZRcCESC6YUuoIs77IKQTlgNjrPAb4GT2KXwdLStdg5bX4I+PLOf2
eBHY+0s5qJO4WDTNPFRtxAC4sCOlQk9a609n7mIvAxrg5FChNO6hWD+/L8WeUl7O
oU62t3S2L/jvR8WKrjCBeG0K9WEH7JToP9hXD8XMucFURrgU5hli03ui7U0KV/Op
IeU1XJdI1XjIt+rZXyBLVAzO7lwNf9fYfg4OHzkxEIaxtWhpeXyFXvDlmF3FnKY2
asYbrUqVx5Uy5O4l5unFve0vNOOXxer0RyKEs1dc4jFkZix14yJliyKum9NaNi/A
+KoUTUeBUJkskDd1YXNaNXQafdSZN9qpwNHaX9C039/BrBP+hfbdWgREo/WuQD6G
7iSAXGJ8UOF1mXh4T9mhBsNMFn1ARrMJUA3u7oXadYZANEnjRqrUi1aHWS3qosZo
yssoFxxgE+KFgoKLaTyWc9a+sBPMuiSZZ+/p/YfLO3VHgoR1TcWKQ+5eaKqcUYNE
bM1eg41dtIsaHs+zZRgxsnTtViRUVU/F3TdqUHUhfMEWfn6877hSBzf4G0gmAGtF
qaudbfJ9JADOCV6XaF8RYR2h7tuUMY1fnJt/yqEiAIvzEIJRbzy7tvXn9QIxcqop
gb+N+45XypM2lBmslwgFvTPM6xjv/NJlfupFmlAwzfGFG9hTzesdu87fKhWJhbXv
JFNr0npd8XMmN92/s3/0zUrsoUVUcAIDiBEwyV92KBAw/Ez3f6bio6p6jQ5EstGs
6uFGwjuadTN9fZNS2CpWeaZYZLqdOM3KxXDPAynxUIqW2O9CiWQ1VLEH6J80YslR
BIAiT+aee3+B/7xg3cNU6BOxeQkaz876SIGV5gnIaVFJby2Yzn5kJEYJz5slucf0
XPQ0TpXRzw6u7UC0DLKrecQQLjB75CzaTpg0sh7Oov2KaDduikuzDXjIzVuusqHn
EUDugGMT05jtLMmBllWGRXiyCVUqX9jj6CUQnd0lKt9b85OSyuC8PrE6UX4NLITs
pIqMA3YNXnstL3GKye7XLOfJZVSFLLA06OSiauMZP8rbHVnka2PWv0JuKkS3LBq0
vSZcV51vXqr79hGHpWBTm8T768wuuMhnTBoqsSqsNfOiAcM8XhyDiXPXBE9IDzq5
DRj+YLX/va+bGB8Lixf7JR6NHmdGTJbb82ewRsNJcYHsqybtgWwgoXDrPdFyImP9
R2IioeGNqrKyhL0Oe8OfW1ISW20QwDq5kXcu45ljJTQd1yXvBLwN6n7OLYujcRbK
j58muzs0dThfIj8KyOlBJyLkpvs+nT4ksdsgT7krsFweQ8+f+D+Snf8RqCoJhtfM
z50oRFFVL42cIgQTtn9BCfVMmxsowi6zWbj12OCBm3wqUnAtbtFILXLKQva7H9id
9XWkMO7vVc9oi5q/JqatIjQGcXbBuGzDvbVD1bn03+aL3T24tasINlgb1eQGu1h1
M8n8/rDthdaGhORKVKKfXmXyVnsIQ4HSlCDajrvywzMu4kYQ+N6+YU20gKdKek9d
IODe8w80tL7uD/jlqHpmv7sn+ogTT6Ks6KEK/gGkzkVS4WWcxyOIGQec+3UOX/tl
s+jvpnNTIW6IVyfxVrH6o7uNUsgAFhJ1zvxZAJP+BXu1zd66FnZNi3YPL7F8OWlZ
xcwe3L0VtkbVojKyrFJZF/kNxgrGKSK42rLvvUM1WwJ27cAJkMsiupTPUn39cf1N
WNAV6qQ/qwrfO4aRe6TEWhRjFXWkvilo7S2k7Yxe5ueN4gdwKxlfGNc0xTAkKpYN
8DyibzjS6AF82afnKLa0yWf1O4i4l8A5jDrG1AEretFOAcSB8UjLC0MyNUnigniL
Qpg0DY4N8CxyS2nvx3q+b+0T4r/A+gtrWx+f4aSxn6RQzrxGjPrTLF1y7Gvixcbt
QINwihY8u9Bsj5bTIPVKuOyoE6V7eYnLtGbnIGeGKFPmPLq5aJF1HWIv6jtFrYCm
U1zCLU+Ex4VM+Lzb4hREBkx6K2l7V7RcaX2A5tH0fd0THoYF+OCKOYwzJipLrSvZ
AywneUve6W7IY149ILPh8ssnvz0BybX9WTBROBKvIP7kr6x8+Mxf5NnWMsoFQacT
rel/OedkbloJO+bt+g3Y994yYwBJ8EzPqK9EavkQnz87SlVHKcLHpdhKBn9GlWHn
KYEXgSbfZ/QKlNwkt+k9xqa26t9vB607IAv8yGBdJz0EiPPWwNwd7FRG2K3CsA1R
JI15sCO+mk70slaicsAXpb4cQKsONCZXyly2ldoQGtvHbN5GzptzdNzJZaG3q7I3
fxjtPEP4Ct3qS1kbYAV124z7J5ZO39d0FIZdk43Cy7zMxR7LCPEZOFYEEOZ6Nhfz
OVrIUw9dHCQYgQbIDzOwsclp2IY52tkhoIEYMwWp2sjW6KYQtNkbmHDEhSfh/5ki
PuV1Emz5otke+yV0twonKd1RHd/7H2HJ9QLsp1gqdIP9ZFmBshgOaraLa9nM+DcC
h0iniJYew8HYY2oALs0jiTMmqxIYwczSgmwyBMze/4Nc7JRgb+GkuiurQzx/1HtC
+hMGSRwt8tRJ4n6Og2FzNxJoWmo4qygw7DXZG2NaEFblcY+JxZRoviapf6mnA9dk
FNQVCvolSx7enZKfubuGT601FhP3zSCVxTZDg/XJw2r0xoq7WA2QxnIvZDRlL8Qa
gz/TX6SoOHB0NxEqUEkWKGMYt9gW2tRenF8ENEcBhoIMjJAmbxX+nX3wnWhiSnc+
E+CliBeYiZfdfh5eGg7mZ7K8z3bndmh3OuxwsVGTe1EejjzrpLvStS29imyT9ZJQ
02v7MUTidQ52iexVxBu6+zf2HtdDSxDcRH/hryMlUstQrxCzlMk8Sl5oSgeOvNYV
hil71GORkdqTg6Kua9QMVxspOHOD5A93JgbiSj3awz//DX/b82M/l8b8CNbFKjRJ
7vgUWKIigTCE7I/T4n/ss7x9V3hsdBBEUhhf7ZJkay+wcQpw0VrAcouFDhTHqUp/
3A3AA2fPxx2WHn+zH1sphbQNTdloBiZvWS83oEPxLhPdGLQqNNed02rZRJKnCanQ
MB7WBm/P+g1xd5co6fqxg+UTKmkUaIo/pgEe2yYpcyEhcYOWRoqffR7LuAzrLEM2
T1jkoqYEQWuy/HRWHJfmM7ahxyi/IUD+T3/i8CaVeXKMOp02i42MneTC0dx/eJb1
IcmiCXVq2dRrIP0lBVRgaFQ7zYvAzts7TJgPwULeL6nOVxMLAoASpi+KoMZwSEkh
O+Crejpfeah871pk0Rp7d9un6IdCaQNiXArZBipQGIb7hRlxOfKZkYeDPpg5nTZ6
3WYqEpTD1uT4W+qlPtKtsY0ks31n4IE4PNKiR/PglXXMnhiuegUoLI+4e21+4azf
A+C9L7XMEg4yJtrHdkjgzBSGx5fokvhrNvv4HnNCNTX8D6KNSOMtHcSL8K4N0e2Z
k68PWbPMyBFRKYGSyh05AELUMKjC9kr1FNbhGPRaa1RYvHIaQY4xhcDMTYI2RN7w
XC0RPr8eO1r3ihzQ1N759LXOP80+bhJOxGV9dAahAp8=
`protect END_PROTECTED
