`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
t8AXwRbl6GAgjb5alPErg2xCEkMqd02+oAlDKih3m97srG8Y21JwRNXh3nRPKDOs
DO20PQtshBxgnNu4VXm35CSHkTRCjXKHx24om5AK7h1zdAoxVLIqycUyfJRuanh+
oRoJ68XD+2igVrKok/QFmFq9MKbqakDcCeBxGhXZtudVs4aVo6rV6LwRroWG1s4A
ab8Tq2eqAmczjCoXsOGgmfJjZdhrItYI8wdPVnh/+RfTT8/9RSZi3cVFKPcmDGii
3CXY6byKSyk+LmXz7igQuZj2ObgKWImCfAvzc5SmCk3GNdlYjAMzghO285WY66mS
xSHW0KDTnYn1Bu5iYHQ/0SqAAqJYc+7KJz/3MKFuxHr6wQ3cfKQWybOS9TfdCqkM
2rG5SGLLWSDkyWs/qA+mfxgPrG8atJaN7vbBNQ+qT6A3kOx0ntZRsGWA+7wB/p1i
bp+Qi8b9ZzYpEW+SQXobfQhTRvNXMu8qt/TFdBed3S32QR+XTQ+XDhAZgVlOqPSC
rrsY8OsB0FXfrflJ9idZpldH17Kmi7/N51Par6jDRbT7jKl/nw0pT3LuRCE1Upn8
xu21OIWzi0txKs300OZvtAbmg9VSA+PvddNeCnuv35MMZTJBXXLrT9SDUsC3CMYT
QzYXSZ4QyCnrWKNdHlTUh+MTamrIgpEN0mWh3gKr8jEbBoCRURwdLfnWjkn+0tKw
Hg0KSCBSzt5wx4WLleDR10ADXu2VrH8yZ+/NpghG2TKLZEvzRn5v4mPnXkiUTIqr
Tjnd8PTkpyTg+jFPZxRAdZIPXILozfgLe5nnuYPamvf4zUapRNqAPKlY5brG4Rsw
DRqoBzE3pXtzVhpZncuRKpGLu77WC9TQtIzPDMT+MS7+w5McInpXrHKp5Xm18jrB
Exwvy+4Gw/+XeULkoWx9qhTnJLWVK1IPI0MSLh6E9u3/CpWC4VG34hUfTBKuDfOC
mBA6UhFKhslS/YcXCH4UwNFTtak/rNFBPBf8KJ1MlzD8eYMDbhbFB51RW6brVVji
nVuxqtZ+wmiQIQigKrqbJ5GY4rLKw5WCl1gxjn76DKLu1aO1qmP/nbK7bXYavtuK
Rho6153/vlkKafJ/tzpKk7A/vSAyIiqOSzYRlEs7OxFFnoREeJDZ9o0wX/HnDNhX
n4njx/kgaeENZNUgmxPDeSBqna1Ly1q7gqMvBhZLlqj9SQPEqIoyXuAFWLouuq17
P78/waK5M79eulRO8zotnx/65re4YScs+sngZKzS9llM9dRQV9sDUyHc49M4l09c
gksku93vrLw8UeFsJabY0FdI40NNH5gQNWU/g1BQi/9dOxGWBS5hxfhlw1guN4gf
i/DI+iePP29oWo9aOUguMw==
`protect END_PROTECTED
