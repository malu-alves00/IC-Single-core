`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
z2cUpwBcIyz2EWRsMuj0QSnUleAGF3Fp2OVo0gGf6UkcHW5tdl4g7hXBkO6H949R
TXi0GAABSA8OIHfrhNb5WjFCl9GT0e0tSrYH3rKy+XrUBHpEHcrXCQTHwvWTKcuy
IcnyHWs7/p9FHC66RGTdgft7Ynj5Cnml6A6nz18OUdt7XgqjAM0Xku9N4UomiyyE
ygmQTSqjS49P+P4gw58dqf/iiYddy5hPstJlfL/fMrdQJf6KIljNLhggS75nn8JI
xPLwZWTh8itl2n8XffnlRIc5LyjGg6mku7l9W3rRTu26tLau4dL1cpe2tzlc/RjS
aK9orsSkmLwT8L6RjrIB2CuRb/Xy16cGSIXjMB95IXHQK3eo8bRpFIRK7S+C35tg
m2l7WDDqjtPk8esZJAhu2JPq/FceGF6mHk6lWk2t+p5xclaNNE6+nYY5PjaYYkqQ
/CjN7eBohrfC46A5tRZukKQFmRlBUpVi3cPxjkxFkzEnjBcASdHiWKLFALWAP1C9
Vu1uknzyxUPb9QiMmyzWvnfjw2pZqhyNIiQSt9+ig5r6KbDPDDfFNTEEWyRXwiak
kJ7OIsp7ZUOuroYe2LjtOo9ADbag9eYejv16xUOi8vT2e69xeDp+/5LjsF5nD6Hl
/JYDC7ZptacxBqY8t2cfuuFIEspvET+od+YmS1/ZKn0qB17UpEmBA539o71m8yLL
Es4kR4d1Ro/PtdFYlAO1AszgVKAKILLELtDJ+uTBD20OtIHx1DsyUlYi5CvXjHtV
0sUruV7s90+lEfhEt4tBtVwGbuoqf/W2Ep3pp1e084No3ivc2TdX38fd05FkSTbE
vCM+BLDUgeaz1NirIt8Ps9Njh5dl28eOLLVm8CHp2H7SLFuKP/c8pGKEczmEenr6
Q4RRxYOpHvKl3igN8wFp6sDL3lV9QGmEmtZc7H7mumhpQJG/5E3y+X9jE3JNY/E/
23sI6rUcfqBP1t5cVpuRdeomqrE9DIwkEcjlmmO0BPHFrT/wKcxoH8EBVcOuutay
8dd4FsJi6VUO105o3pJVXZyK8CElJKKOuoPMa64wDNlzafYr3XTak4zPLCKz5iUw
sjl8h/E4PxwX1wsU1ZnktbL5qBteDjgO9pjMgt2CzJ3vpHziV885zEixHJtn+lyh
YDInP5MykrvdcsI/ncczexdl0knmzhTvoFpGITv6+kBnNKsoC+SbT74dK/usFBE9
ZYNGX7Y2BLsJ9YJQIGS3fY0ZSYrTjzqBBpiwAzkCjB4VfnUkjRvCfi3t+9Tr80ap
Y/+b3kr/zqm0k4E8zKRpK0YejKioSI1PONa/mHFyZFQcqNA8vb13uCXRpL7bjVgk
Pp7g4o9mu8uhsReWkEgyH7HQ/Ezt1pgUXrvnQWI1bYopcVY0T//oEcMpKhjvc6ui
5VtOpPAlO9UN8zC0Sh5mvw==
`protect END_PROTECTED
