`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OsC6ZDi2OQA/0hUowkV3btdxiQVpeD6HOBgQKVswbL8eQ6Gzbs5zKok6FNNqGNr4
DBnp6t3bhf++ME4ujX98hbaVqGG3M9mpQ3qfkZNCMWHCCyopy6TBLRMg/oIkc6Re
rYh5WgRI4sG8j7D3qAOTdUYB00hdfLTbw9U5gSYNLmPL4GRTFO1b8x733Vr9D0Vk
zlDU0HIhdOOJUllIIXB8wY0YbrwW9Z/qJBzVI52Pcv6KaroD5k3JNMrgILrovL0H
M1for35NKxgY+uxDcBuomKShmaF5TX0bgMllZzP8kMj1CPx5RB7pJnTPn3qQWFhk
lJ630riww5dUEyw/y6hDLHIu2+GTYNfNI2kd9JLDnjPo4w+E4z5V0l5qyP1vdOIa
mwHvshxTuspJvkg3hL/bjFcqD4jLHf9JI0wQg7ZP3cMxb2D3GNC35uPydUI/aqS4
Kud6aAe/CTGOFrhugU2i0WiC5cuR7+3Op8NVtM+RFTFSOXHUlCmUpHaSJ4dbWLkA
7gnZWM6W4Qjc1YSvNv4seZE/tP3FiNBNw0V6X/c5FkREybo16mEXtXx61zcpyP1D
R3kbF1bMkPFW/ZD6Kl9KkPuwA65IFz09Y11QWPmvZ4DntbI85SQfgNiRdSLGyuQu
AjeYRDe14HMkfUtKOX89L+pTCh16otn7c3F006tlV6Zs0UR9HNtTEOdTUNpY6kp9
fOuJblczZq1c0gUU54zlIWJrXllnzNWX1anzC11TTVTJKemER5INPaB3sSxCeo9p
nPow7gt/KXpEKUNYLt8D2vQ7YfmDw+LCC5mh7Dkl7rPPW5cbECKFYy07LbbB25Iv
tl1+4GBEChOB9p1iO7VkcRLXxE7/QKxgu0u2HwlZBPDF0bKTRlXFv5OuU0605SSt
`protect END_PROTECTED
