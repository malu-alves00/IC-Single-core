`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dgXogml7eOf0QkM7XxEC5BfBo7k0IBGoEXQhQmrY5i9DgwpcaMrCax7GfFaokPhd
uGNLCF/2BxwEULFs8poIXY3VDCBh7DolVJ6mVLCNVpIYF5V3SbuTEQEPdhHnEgpk
FIn8sI8tgxXdiOv9/jVEva6lBGKUGbwlN4gtZR8dqLD388eCev8CLCYetRnG/0Tt
qDRj1HEwCvPo1qjhpVtJ6XsyKGbwaFnlqSIpXvACatOoiRBNYp8QGRK1GFGXtMOA
nFwWvbisVJoSpoaUNPbJRQHIVgUNBLGlA4nERbhfcltCpxyJEYCaFTKIlOotKf9E
izZgOzTH5JePbfxjtOmdyxqnnbRlSTwoG+/cRFDTJJd0uTVrQX+XW7i7Lpt7g7mr
liVLeUsl4sZKSZZJcAnv6TchnjyG4Zwbt4Wgi2edeLfzFAI59wG3vh+9tsjxFeIK
Dz6FX2Bw8vX6/dUXzUhFC/AzJRkN7ncrPa2NIYJelt3I62YOy2CxaWdv8NcSUDOL
rsREVNQXC5PSYb0eyMJ4/95MrTdb2WF7crmLgpOYoutPdU9e/Mvi0KtsJb/S92ug
VKLb/qFlcaVOJARhSqcIgVZSCPC+PVvz3qyAAWHjolbe3MAN+tfx3iEJr+2TlEWE
uSs82yg9M5HnF1q8WhyfZZMTZK/HUBmuGYLqDebhCjMqdcVEhlQQGaHV6FQKQr++
8ZdUlKurgOd1bjY9LTnfjV5UjW//J576pPZ+rc1hCIPgDC7ReHeBeve3PY2MWTs7
Kz6JO40AwJicKErnKYxFTBgUFSa2pqbIuhVtkdn0HPIXokOhZdlt9GS8CdTdsJIk
47Dl922KZ7Smg+hbj5+f0G6eqDwWYs59t0tvDN+RIjW5MBSQJlu0NALMPgQRBxeJ
jGsjUs2lG+0HHEWqcxk5B8Adm88GfAzsHy4RZZfFa0yJVNK1hf2uW5/wRUzqxke/
HoTvJYwyTo8h+KJybRm/phgTOlsBbYpN/fOTWeGVykbi9+QopnzcZNUoLO3IHSne
lDSSpuawbABpgauZH5r35w==
`protect END_PROTECTED
