`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
M6G5H7Tgdt/BdrdQlg0080qN+XOpmU+0Hat4ZjRZwTbz8SbYEXEJo/f4Mxztzdrr
KFMK60ndiB4UDm/nkFn2vX/Rr0LrWtdaSzHAP672oqCwrG02u9QL4vFJexBzWxwV
bGvjTdC/vLqDAJXt6W4ZFbb8MT+TjIzYPsj+1NWqeN29SVbmAX7k3E5JdAvyPdha
kE+0uEsregEXSRSDHWdrQM/w1m/YL1i5lFFnEpfMSWHv23V05XOLdhzKzv84yku4
iCYKNyonlpvAX9Qey9MpRMiIxHaU5jD9FoEWzKRQD2OeubzOe3HAVTcM6I+a3Zni
f339o20crpLkD0OHlNv4P8YL8FKNDvDPacuMbRyOStYY4VSaLhzgppQi3eNXG2YJ
1d7XLJDy+fGzBt4cIxKBaYC4HcYOWaJbrnDTY9KwUKaBdjLeXNT0gaiD7LCoI4Xo
fFzx7nTRra1+RQtOMsbxDnhIvJFl50gsJc9QoHULG8kcvQ/8AlvIOJi7+hAWue1d
TVQThvJ0zl/qrKEUQY8ISCmTSZjwmp4SEB1SmUXx7vstl9zul6A01fAso3P0J4lk
+YQaJPEkH7Fbi1yDCQcHvA==
`protect END_PROTECTED
