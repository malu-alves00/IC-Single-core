`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
T50zREZ9uUBr7K/rfL3JyrXpSj1Bur2cS3vqIHLzvY09GB3Noe7dHvAE1+w9Tjq4
ZRm4Q3KIq29VMHaVvnaQ6jgesIsfOJWPvgzfjs6fAOG52Oe8RmzfnuncgK0QOVFd
thxdCtSm2GmEgJNKnbjIPYrIuRs2IEBY5atDx6mpQmzr5+QFNSOTv9fQCmCl7W6b
anmPAcBaoNKNCgOb2w7Jf1RzSL4nQ5wqJ8kf/XLuwypBcHWW+rhm1BaoEZ+7HQWt
Ph0hpYJ6NL0kMErGRc2u/gPJfyDf2BOxERGO0DpEl+A99bdFtf10RE50ikDtLaAf
c34yY/kQAn6647oPN4QDlpZhKrqqht5MQjj+8i2+VTeuQJaaFJFRlHdqhhI4SJJs
ZFftpqpvxuRuUPkMdqgLbwr+dwe8AnSJGRilXQJDkBG1DhLizgOL/ejuBRCLOfmb
9WEBqd67dmucWgoogmSSsHzgx+c/ValJBbUaRGVfrSb9tiV7CqX2EebALP9konzK
oo4RekwE1X/l2nvcvdJCguSlC/vM1K1C2BwcpENzZI1num9SlMEnyc0NBE/gEBlE
m0/iL7dYyKEefJVcQNxySrmMCzoAtr73ugEQTsdTFpKd2us3xDlA5ltSOHA5u7Vd
0iq6hoPkYmvbhcpK9X2bvW62Qoe9eHQp8b9d6yRYJSQq+VmnkOwA7dIkZH4qLpEI
Gip6f2Pk7s2EEFEFdoca3+dzANZ/2pw1FgAiuUbnTTtUrr6KNiJPT7jajurQI10C
5WxNSIzhpXuSkpw16KU89699zCrJYwT4oFUk4fNV/cEdkRSgbXLyfhc553kqT8GY
iJzQ8mCQR6WtYW8O7TYi57ntZ9iooeTexQPcnQIL2hfG8OpvhwnD8IAT+gJcOHxZ
yZBxFyNeDFEbscLGuyjONwJHp/lkQ12lDplDYLPFHYtHxrq/hCQElNYL+6jESjlr
kMrg17Uj4iPrYFUvH5DtYWtpLFmgsvphLDRIlteWExOpWXp5NJLIS41j1PtQOy7k
SxwZ5itB78dSqDDfirrUOMZP0E5kpZTj6ntynB5iPfn+Dzqt5zMz2ayXzbTu0/Ub
bsH5VNQKJeKG6qzGr/MTdAjRR2WNmfLpgkvD6KIUSQYdGQ+goundukgQzu1VGaHc
e7Sfd/XP85sueDgpXb+WwJ6+boFYXn9GPcPIWHbJ33fpBxmgrWvKt7inyJCH67aS
ElXMe5S8k9/5JSddXLDk6mq1T1fuCwMu40TBquPpgqUB26SdA0rr94S2sVZTd84j
+WbXolrWSOo5TCQTSc0suWfF5oeP5bt25lpW92lqiQIyhiP3fNV/W8KLzY3tzeMK
HtyPpoS8GTx/MusavWpY5w==
`protect END_PROTECTED
