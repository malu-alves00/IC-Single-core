`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aryaXkfJojZ2p5PtTXYYwkCVqvvN6OHFA9tnqk+8iYhEZR1lnuhd9aymlCxT1dfP
EobC/FgZXBPMiip2eY/oRwilZOToTPPZzCEcabNfwzKrFE00GcoTtpmGOK3MWUQa
JNEZSdZfsos1Iltg72HUKtnmMG//OCPEvuhfdCE9tBY+MunORf7AiZ74PJ9wvefJ
XsMQUDhiNwFbn9pCFYAnqEgVKuYBfAc4Pag8rWPb9ycwfT44b4inqMpI5sPB0a5b
3w4SkjBwDPzGUUwF9EMtluUHrb9/eX4WpCICyGRM1gk4o746jB+QGMDkPMB4Y60I
P+qjc6jiKKas+7ZGTgUdLzm3J3dRTODQVSAVdIBKC2r2mPZFBWuTtalbZFGveQKf
jNrUw5l4m3ParQyG/Cwmvq7hEqN+vzurDTyLj1+reLkRpUukMEcua5YDD5sS/cj6
P7aWuK3NEvyU1CMw9FeqgwA3X/nK2+bq8scsVn+OxIj/FHEn2bjRzEUWxn73FY6o
w0Wxw2M7xellrMWQDZEGf+/Lg//JEwrj29h9yFxgTwFfocDjSt3Xii55ClMqbDd2
enbbmKhs6dZkwaPPD0K0OJpGsubRwxr6zTNciqYgiqH+Mn0ophNYxDiUttyR/V8a
nKLXkvO0raOJciVPY4QlvD02Kt4PsUAHbJLBVq8cvz0Lc7AgEJ2Zu8LWpAOdk8CV
4MNalcclbpFMP3CAI7zsAXiVeI520xf1AoAUarHS2v/8Xe37K40rfD6PlaGs5T6H
nXXVBNKYK7doLOGky1WLXYrtSLbrveTyLMq0xE6/Dvq1a7oeahezedFfFlVZG9FM
`protect END_PROTECTED
