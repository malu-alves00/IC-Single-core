`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
apYqtO99xlMILlfL1+XCJuwFDOMlg9AXsfcL0fHkIu0rAWIp15V9gm40gtmNhFt1
xtV5soon2wiuJpvhJLf1xAYEw1TetwPixb6zLCXBv6eMfAkOtmEafTZO6vV3o32P
ZiGmouUYlxLQh9+RNYKOUZMmTttlzq0ZINGLSI7to0f12i52MF/ctMgSvl4Io10J
vJrd22X071sFDpmwcsm+I7igQjrH2tcho3Bc66AX10taWimcB6wtLhl5kzb9hhvs
pcWchdDw1dgoV/HTlCxJLHtqkaDftsSOHsJY/fdyobmM7KS1B6exiLkpbB5BYG6T
/E93vwBP2vrq1OfMtezMmSuNKIjuQGeVg1UAxgxbtwiyN7gKYIFtOnE/+4yLuuoX
K/ELB/Zi2T3kYKYkUOTYPwuQGqwS3GyWYQJFccqz7XliijEkKL5h876QW/Ufdq3c
O4D92VGClEQA2PPr3fuBB9Fe5gRgQQ3vl9KEh9445jtuA08sIaMLfGkApmMZ5Dmm
h5ykvED2WtBd/Yqm58ZBdW/DqPE0F6v7K7LoeiiFi/LDpbcv5qWpX3M5Ld4ldBXd
GfEleCTpW6gnfpz+5m/pvM1LcBHpkNCpLrnBFmtGqhszOk93OAXk0OljhxhNoetR
d4rs54rgKA7iFMi6ChcmDVxWoa6oiESEdNB+nAlvuA1zWF3XO7R4iLINVkF+imQT
PTJQOwjNWaiPfukwWj6PAHF7EuIkxNewJfLmYn9hum/sf98YlJmxDVa/edOZyYU6
X26s5vOhy4gRpNYSSnjMkfnqO7x/HOx4kiK8yhRQKxlnjYnhePj4nQE2LMO/puEc
O2EZsvNr8eCVMHAiscqMcrHWF31UVcKrT2zUo517xuu0LLCArNLirUxE/DenMhvZ
a7pGFx4t3dlAFgVZnz/YDyUsjS3M7g0N74w5vxBE50vIsJ3sQmpSL2eqGSrlVVhy
15ABj1GuekbCzo/IcIhjmab2mFogGzWKgy0Vpg8SWuPmi8jrD8GWPZ9Tye7k8DLe
pBJCps44GeHvztNqcmk5WG5A3w9xYHip9XH7BIBSeQniaNI6TjHTG75v+sWyBiEP
xJ3D7VETwqJFUQ8c2anwSFjPyl50IEolQZpkYVo7csXd7CvI+7BbNDvKw4kEvzSM
5w2Q/uE/gTVI2gINd5s/Xx9TaDiX5WBiRQNzSoOZRBrTV/cD6RJz22mnl7EjsVFj
LNNBpto81ffa2q8oe2uAMcRdNRAxhBYUas3mKzTabnzI4Cld1uOu3fd3GCQoikgu
TVjsYfCAu8W0b5VBDX0J9pZ1FU5jYmjVIHPiiKjH2UuA01i4afc9a7SlRwyA6Ugf
ucGlHz03v3qm9MTJPj+qQ3Em9u+Ug/uhoKG6ZuerqDs9Pbz6cF4bIl89JJdPRvbJ
Jskxb158+veqlZfRtY+HD13T1gHxjidEyJlsdl+QjoxWGa5M1+PLeVMUEV1amGEX
4jRigcm76GMTt+xW8N6SLLkEJ0CXMWwQBejM+Mkfd8RJYZWuF2iDj8DzhBEJsehg
2RyACsy9g+2Uhg2KocqhTnJnKAyuuBunkW5GRVbk5P2nucX/ljXGBjmsa0qb1SLA
0LUkMfMUihlTycuSwBWOommWoQT4uEpPFF1YovtJTtSzgqWsGi2DghhfeD2+Ad7m
Q6z2KKa/ZyNPRHqRDwKtwVRSZwp/fkj4GvMh3LpZ7ERDmcAEjuG/zymmmAx5T+q0
+3QusC4FOzae/64xV6NMddoKnuFUvR1lRXuqOEv/feAubxvZW6H3cgNBLEkY/uVS
NAH9oq0/DGMJ04RSIBVBzC2qDfHFaqsZa8oFBs1NHj0C1A+vpUK0WLhVLVmgvWsB
irrYNPbOs48lQCjUVUrW8Q==
`protect END_PROTECTED
