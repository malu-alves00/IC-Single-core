`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
x5m7K3MGLREYmt9BHDZjhsjEE1IcgED7dMxglKKJLy0lvzGxz8CWUFE1ypU9aabE
Wq+iR6wMpQVR0+JUatbFfhkLcHIuZLXXZs+n0fNPanvPVMyyUstYis5s0us8DZaA
jeKk4GgqxQ6gsZiYFtoW4h4CSdnGfqHC/dLkVJXPMGbOKEVMsPUY+FWYDKDTISow
5ggGSrSuXXQ3BpPmLsBwn4Q6NTd1YQ+5aNtJiAfgkfPiF2elBPkEWfuomTmyqUMF
dAGejyrB9g5saY+UfVBjPHPsus284Gc2SMvfyShyFhCMH00YC5iNb1938cnq/3i6
jM1lOPB93N8Dqovw6lQOXPmHwdU9RkC4ig9oCRJHXngRXuuOq+VuUJZo6sRBAVyA
1fbRJXSlLIaCTpbDO+n6YkTUIEwjU5BrcVVbxRCd10/D64kcTuUsv38PDw4aQYnu
OMIrD/597G3bYEBK2/h/9toVQeMG/IP5aGJBn3k02VGTq6wOgMirXidE524neGRS
3hewPgXY9oGeYIe2fZp0l8IbxZfOY/dkUuXDwa6oNDyqvlymxW3w8fTKIRLOyTNr
fhleJhyZaytWIKMwWqjZxdvM6304BsNzs7ebFVHo5zDLzqDrGwej3/QFLz3ea1q7
LOQd64h6XZg49gYFJliwmWLRveWFgaiyqU+oXN8OD9PTs5yPKgkn0oOSt9etLAGW
KNmSF7g01Xxr7UKTUp9R1/U9VPtNkVt5cCSMcpiXR9a17CTOxoFz3FtT5I1xz0x/
jzT+psonW+bsI11q9K4UtnuDrXzMPRgtJOvbha+6kaooXkMvCiPCJt4DrqaaEa0C
qjp6DSTH5m6YSN/qBVWcfE8BKrysoYePaFeHmZfa1rFZeTViHF8S6O1WCxQgzCs9
6Skn/XWFfb3sV2W8U0gPaDBnD6pjuBgWgUInkEwFh8F1WnnwT5OiHPL3z2fie2DI
FqSuENmJ2vt9rd7QEtJA1lpSAdCDG4WY+qwOn3/nqiNEGckuOJfhHqSpo/tAxh4W
u9Z/nP1xZ0m4oQwBl+XAetDcSEnmwpfsT2IMvHnT475z8vZGdFURbkcsZOWQLz00
`protect END_PROTECTED
