`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
V+5JBy0GQMOXqAxRShJcMgrkhHaK2TXYv6VY6DjttlaowhR3wePkVeLbBjp6FpD1
WaxJE+VBffgqhYHb/HIzQtMidCfxv/eMydT9ntHuKmOzkFIecpd3f+buK7gIaL6b
V1Jx4KnGfZAsjDlLoqOZWwR5d+mNnG7E+1ezIq+a6+TxhmdBoWikoGpIu9AgjaR4
QYiwi95m6zVKLbeLycuOxdZ9E1gVq6/luuLBpQg0TPzuKtH1eaVHwqXW3VoNfU8n
LiV9kWfdNFJCAdI8ibPwdKoQbzJNoE8HSWm+lwT5I6515JEIfyuqldRZUpKVdpBE
Mc9zS5rA9aJegC+CD8643w6mh96b3L2Y977wv9ox/wn7SO5F6dXbZtEfE6hQb7uM
rniKEWvp3hbZVEZfEiOdbyPVaouw2JKP3TjwNME1UjO95YiFI7FmbV425WMzhYhR
EqaPFCszoCC/QLEe591BnNmCpoqJssQfrrDXw2LR2Y8algc+Z64qN051JHpre7Dy
V4YRTw1AJEKsXtRnj/ewL3emHNwrzwxDvZrHGYMQ3L5uBVtGXXmo5I7+6ya6PZCs
OwVJ8zyZsAq15SG2oj44UZ3lkjkMZw9BV9OiQeiZ0qat8HAFO0ldvC2UsM7kQNXZ
xyNuaWGR1oORixtPs+2ukQOs3s8D+EihztdrGI07190AbYEDT40G4r94zRzddpg0
rx8agm0VEuaNgWRa/Yu6TdQJmGyiZuIRTUCg5jDK6aRtuYIe+OYxUNFDjCwO5VmQ
Ap12sGDLSOeNk/UlbsdQDhNjTzBs7oZZ6Yq7hNzRwHm05O4YvclHbLLTxCrD78DS
df541hYAmWzyCMqYq2k0PfxNCV9UpTpQ9Wpd2fF0lePX8n8RePwE3CQnezbBrdfC
QTqnX+PAqdxl67a6eIUZpAHmsLGNJaxQvk/v1ZwyjaFJ7+RHQZ0wIxTzzR1zVT/H
64UhiMr7syqPTVkHoBUJ6FsPJ4zW3+ndbfo9bTp3IwqtxQPapRJxca4Xz3mxcrjc
JQef/NIGw9LX9wsQu+O4KzFnDD4HrSsGs4QVDkK9YLpAH6a19sCyTvpWbicRJKtp
gujuITa81LHEt0lB0h0GGQvl9832QOI+l0ktZAD06bzq5zQcLUNEfOo9yg75ZbiD
na3zHv/Zd0+VGCnQOKHvGGMcIThXyFP36WufNy0u+ZtfsITrVT2yvQHHDTl51Epo
Z7q0da2DiIyVMkdbuw1UQrmsZ8ExXXCd0oCfjiVFtYW5va7jShn9rbeq9ZSF4BgH
BMyTdKIv9Pn5YtlT+ikIJqqdVp+STjC7rxd07RkbaP2bDMjp2LINSshjC1mWQpnT
+oDQmckvffw1yXasn8ugG9T7X1RT3gZClJG4XebK1xOj2/x+T1BlnAoPswpA8Hn5
hKDDcMk7Bg/qM1zGib/jz289X/YOGsjcP2ScX7N+Qel3S2RaKpevPIiTpfJxIzmv
zmFb2zb+l66tFZ4R1M/jbQgG/JIbrLHN0qlIEaXvml6XsMqdu4m1ZWv613EahwNH
7dp6kXwVGF/O10fs+wGuGdChRsbb6cKnFzfOBUi3LOeA6O0WaVP+13SrwG+4J3wl
KC4Y2D0oAYmy2Lzda1QACRSdS0mBDqXuBnXGbTTg4Q5itDP6EdWK56GyHVA5LJb8
4LqeNyi4e37fm0UhoLsg42MzH9WFqzLmDlDDE8cL7+CXgxEFwTptpLm0Rev+A+Be
hT2L7jeEt8HFhGm4uwN8JRDdIV8YnDN99v0LL9gPFsNegpNuLHd7CcNCB1jKSaEm
ADcJhZY96JbjnFBiOWh9r9RuQxt6Ch/wn3B6TZQWLEEvc1ttrHvk9Xt70s6lhoOK
eUxnEk2KILkPxmmkBYby8i2WUyYOUS546m1YApURWP8Zdercwi2Up1sjSTxOaP0p
skdDeEFsp+vuwFtv9UMBgUKXe7R7lqm9/9Xx7fdyE/lcUPRdcLTkVnv+vvsNHxPK
hXxlJr0rBtM4IbyuFJjWNcWGAngbTMt/NUzJRom6VDGSAYM7txGo7XxtjNE1CWJw
bSpHmi++U5SmTAJiW2whkxLlX6Pzbu5+hcLcJAm/PdhUw9L3wc5/Lw0N5KkNkXLP
BT0pr7xx1p48KjcV9+4I7g9anmOMj0M/HFRW5ZVasz17hMkZr/D5i6DPolhVzpdM
ifdJ9NxYtIbVubtM/8jKSeslxU4UepUjlzwKHpZnzGMs2lMn/9WDMLLs2Nmy1XEr
GFxUk4OJQx2sYaDeuMUGFqOXn8SILm2yhvxjfrzeHpAsD5U57+olmk37HFfyrN/Q
/9drSEyF8AKSHWsUCXfBuuLbauiLiJ78rP9JVUQm1lm86pks8tXSQtbQ4Uo4slyj
aFM24BITY8lgyMWVRvgc3K1wLtaH7YXWI0NOQnYFEH4PvivMG4vH557p9squYr0Z
GcHXW1ptVdYzI1XyZxfrJHBKTeVaSJc+fcjRb29VcdH5zzUIowVAnZba7fihzYhv
C+4blc2t5d6Oi0hY2NviUzwgLF5Ll2Yxd3rkbkeH74OeFEOKCn49mmavW4DoAw9w
UzHTCU2Op42p4lLi1mG6CqrEzkzkpW8FmHeIqW0SyOoIJa5iRSRpxtPeXynsTWZj
/Hx9N3pzqBOaWZKQuVPxqlQKcgdZ/Pru7NasEoFBmWTBzDBjCuaX1mnE1eF/5rGC
UXXK5DuQr4UUg3bIIaYWBjfj6ckpUS48fzCCnVrToeQMf60+cp36VKNh8OlqdoEZ
QhjdcTtKCXeKdH1bkiVe3FFub+6pGz71YErUyEAVVMc4NRsL6wbxCqccOytqEROb
iQXz8VFmx3PA97w3E4KuFLwKrjK97ZotMsyqcbxLfxID3Px0DazKjnyriSkdufBN
k6ssM3hnzE9+2kkCcnEa5ICdP7yCDA7gV9dDHolfJ1GWrBqJZRwZhp1ulweGuyEN
IG9QvuWqU6p3ZMmLwW8zmfcfp+EkfU9g5XHPaWS0bEAle3n8u11t05NA/Gfo7ioi
50kYhP52MNf4+aP9oDCaU4NHKJRjrykSt7V+bqQWlpAk71c+lW2Ct2np6LuBX0YT
nuIWw6vGAIpSF09MumZmsA==
`protect END_PROTECTED
