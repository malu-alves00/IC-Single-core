`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
t3pQvM7m5Ex26fNgiezTvku+Yhvm0rMA3vlCcJ0eTTOW1FA4ofRonG9VoNdQcQJE
QxSmaRlOjXLNA5W20iAWzrE3+w4UKEmFK651g1NKn32TChYXyW0uaQWojmvWGIV5
lqrMQoE03/vrmfPaCKvLUzblYpY5id0aAtxvAZqmy8r1v8K3p1qBaP8iQtPUrlYg
IkSye49gAMBRWjLVL25UeZgEgOmJ/sfv3+MhCW5ovdBocQT5exfN+1Dvrbpvm4l3
jG833/gFirgoLnF8xVaeXXKY+vvuABwA7dLXVlPR1hfYWhOlis1F29hKg2phCWXi
hsRQSfOg9F7yLW0QljNrzBrQ2O266Cp5R0vquy932aGKoj6HKc7Ia1R9vzlLNp4b
`protect END_PROTECTED
