`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
H2s0NAv057Bb5mu4o9K5RzdyZL+YVL36brZ/rW3A2gi1FrGrO0alCyuIkwoCttLP
OXp9+Ao+U1Zc30TQrzDAEyc7EEfrPZl+ILiW85Ubz3uWaYHpPsfaTcP0CUZwrG6j
yQDf/QW+pSLCHSbLYeuTpvMbP+/9Do2jzGbZORO1XgCM5NzwVXfPItsfBcxy6xA2
QUO0uCGu882RzOXzTrz7GiVX4jDOHaVaJD8XaMUqlHpTGL32NGOWJIW4j3jQTWqu
XgRA6IXeObaUthIlJfBiPLhWsjyILH9lL/DlTyOnf+Hqz1p/QStAEf5eR71P1lcP
EmJXMmrLbuJCQEg48sL9kO3xF+02RCkAyjWCJyxPTKg5MQqDA84qsf8mWMKtAP8p
oJkh8ozQ4DAZxKv15OyIiQauGy58QggSFBit+2KP7IHFNq359lDoO470nwMCtwEv
XpMde3fRiLmQIOq+Zqj2+4pW0smqpt7bscS8yVqGnOEhC3TqYc17mmdjUbf4qMnR
fxfexXoo38Yr4JABCadoFkbZjOiTm6YPLUR4OuprovKJtlxHry/d54XxmPsoU1/C
JCfIj9A7cKyPp0gFfdDprN7BxFZJDNmz90DF6sP/jiadusW7CQNSP60k2wyf8hxO
Gv/uJnLctEnfnzRxIfVa8im/DNhn9UGq3mqOSaF38OzcLu8wUwccAoH9RlsqBuzc
7Zkr3km+jE14rOuqTfpECEG2FJ51ETlj1nNEI577/JsKFDwpYiqEoXjLN4VRoehU
gyebNwR06WQSZUAat1uwo6Qa9ov/4X5wbDPJ+S0REB7Lj7waf5Dl4JpngYM62VMe
i3URstPqrjBe6goQMZchPr0lIT7r5Mi+dg6QTU3F3SsPjWL5gw4D1dJvuIxxrcPE
Zu22A5KywQvVqdrUPkxgG0X/eQ/nrtcmXW36XKygIuocZxRna4DrfGWxqY/YO9bT
5YYhBT0Px3vTRtFQXxtHwIkX7iHTyCnf2hSGVyWEAZSP6odJ5vCNlmVAJgJppD46
2FRfqZy22A3wEGe7wJIz6DsMu1rKDfFvwmn9LwLfSpR8BILegiqlbBb55n5iuFaP
zBHWyx7MjcpD0P+H4xhQP2dX2nzGpCR0il5CSppyPiIYI/nIIvGu/CSWeYGizxED
2a1TTttp7/Gp+TpWRr3vkISPSWIYI3f1T3VE0D2r8izE/0Cl5ErChr9oCLPPLOkG
viT4ZLpU6kQZ2dbFpR2+DG3BuwrGmjC7S7I5s1yG9jFJVQOqDM//iF69xIFmRK0E
m2zvpUZiA3FXq4IgQosEAFRKFF2uQ/xNYcgN7QdDBAkPt3xz57I3SWgNOlwgH33H
nCmTmTj9TZHumcmZ88CXHDvsiltQxN6ucNGvnvm8HzcPAqfew4WY85Eo1kSFr80j
tkgWErV7vIW2xDH9ZyV6b+7TvUEhKs9yt1KcTSZKDeI3XctruOoA2KDY2vG3B+gl
Cf+liXBJK8KARAIY948Dta7AmJk9+1voCFijM9yL6tOoLPdHqbh4UfYvs7Tvh9fw
jA5kD0V6V1L12/+X26gUuo6QNl2o2sou7n3K22Xpc12XmORkb/nWtA3/AHx51P65
dfvY4mybVpCSJhDTAP7PjFYgIrjhNsaHj8YRk1BpEIgfPyyzPOGDGWPEQL5Dt2fY
77ix9uvW433LKjNwqh32c+r1yBD4b671JM5MQbqRmL7iDLHyIPRo43W2L7izLsGd
LM4jalhvCa0e1NMYO70Y7zRAtX9VO9ZLt2mFYTVAftezudiUylnHjcggI51W0g3S
dKVw8SdDJkux7qbpDAMfkqnCajtUDIxEPoBzU36dU7QLvde0Yon/gCnsobCgX/9X
bignqGpDT61is2c6iKjw6A/LzpN8vBnU+Epwii7B7aSHJ94i+7Dm/qhM1RsgAH/N
`protect END_PROTECTED
