`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
D4Qu6b35p/AMFKuEl6Ir7eEQ8f+ARuOH9+x5W4kILCLjpOdn4GAoHMHUOR9ElQi2
kAp/kCw1JjHz9kiqLhNM5GKFYpjRbwe6IXugL5XBL9fwpJ1ufbHJ5AFhzdLtArAu
kgzCciFkPrUf7VCRzBejB9RRWjqUQRlPXT7vu80lsY45davwAdGLUvJGxIt5CKZH
6MhDIf85mgXmKpOOV8OS9pRu30MY16TojdeVRUfixBKox2SQaOtd7chBqhPYruxL
mfAfdxlFyJ+X6VYaJY4AewwSBiQ3VRqVUJTQnIQ906kutCaIR3P4T0+m96LEMSvg
w8TrOFfyDL+6Uw+QswanSDACcD0gHzCtoHbs9YPOWVPbWYPQo4WmlpEKrRncp4OQ
b+bEbWhUVa2wFORfY0Qido+tPrU6s+gzhkqhArBnAlfVF1jV8mIYHicZ9wO4r/9G
jw3cFbrV6Ezpd3KJJ5JgHfIHzlhJuMzonJdaNMPjcjTq42vRvRVjSQa9/DjbpXQM
qHeV5dIQ9EIOap9VoHB0IPqP9B0YkY8z3fkDnNqmMqC5EpG90ldpSLoITUb4BLaV
bCC3XUWtG2YJYO4GYq8VDjCrbo63bxbPqjusOnhVL5FQgOGOUPoKObka15uH2Pt6
aRYHsqVXsl+x/bK71sLo794Bp3tVmAQzSuW3K7Zpau4QTJ0RJTR8D/dmE98a4GtU
+CVrQU7NbWRNAqiXtSpoh/jmQsmFMlo22YpbTisQHaZQ+Cds8XuEEDITcvt33LYN
abv5Ua9bIM5gaXy9O2YDTwtWz5L4+USzGIxzNJXToQGw9Vrq4bn9IorGB94RaE2N
CxjQTnhkUBk3wVNhVEIzoWXtXAL+tUAx0wowZ+BdM4xwhtlkVMl068w5I89gNq0z
95S8lb9OctS46ZIhEWZkkK7V5csGXrDpCi6fOrn9QvwxNZo8msMUc8M74YhsIcTq
Tzz4DQSYhV2FbK1WvduutZBa2300giagOwjqnO7A5VA9hsFMAmVMQQ50LV9WN2D4
NuO3TP1T4av+Q1dUh3adAjYmBBHMhlRSbK1Xjpa2tqHAa4IG83+IgLfbzPlbZAs6
97pB3uadTFcrd+Rm9vrMGgboJefbnAMccfzsSeBDbXMQzAG3bUC4JNuST65wzkP/
NUXiOQKY+qejlodR6ZFK0B590d7UoORlOx9x3P0k6A/Tx5TI1VXJMlOy0waC0Az7
yRCmW3VO0SGpVdkDgVCl7E3rd6z/3HIjjUcKFzj7uqU1BA+h6ADO8U0lFhJznVWI
MTygGdUTFeZJinynKFIrqk0NZgJ4Vp0G7Sviao1bx6zFLK3Etg47bBU1Ge53P2O/
j+Ug1DTgSL4B3sGqd0kKbf9ugbmArh/Ji5oV0fvHmpaYai9mbaKdVfHOqYqRF6xC
QQgwJPf+D89ka3jrUoZPNtLdTH+ac7w3s+OuM8O1WQMc38vH5OYTV5XpbyBub/ij
MfEr/IBRdZyXJ71ehRqbUA==
`protect END_PROTECTED
