`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hZ3wtgSkmkv2cy+Le/CohuRaYf2vNoDms5Cp7o/suB7GErOkedfAB3YoDaXE6Bul
vLEM1TW6Env7JOb0EZkmgPJM7qTKDmqpQcd366NpvtbpjJao5bw0QCuMy/PjsZ2a
8fqcadxqjXWuSsPFxkcJf+oDP8MOiJ1R/7N7Z4fVbywbq2cvJJPq61oXMTshQ31v
OcRsGX46Vuny7iiNEbKUfkZGRRwUdLjffGuyMB//3wpJis+JakCG0Bd9yHvsxBhd
wo1AqsWvU4wnPlVknhEdPYHIMzfoV1TyXrhDPLnWlRZCr1mECXP+JMNdIhC8jO9h
ZTQqO6J3I4aHiJjTRZzhIa1YFROjCCdA3Oy30TZ4TH8bDgRB0+g/d73Y0mADNTdC
C0Mw7KnXZ/uOicU/UUAWJ8EG0YkpkLaC78VuYi7FRO2/ElETtsGLh7ggQ66S0Noh
vq1d9S9j3030pXtG7CadzgTa1c3hmz7gwaah4Fs6IrAVuuzzInnY7YIFYtNPGmCX
sUfQHdg7Rb0fjSodRpmgoSTwLZnSxMMnOElFJojLJhSnzdc6oRtuxpeHmKZT1xiI
u8FDhwJQnigZ5JDZAdaGDTtK6uuv8krFEjBgt7Xzxy/X7XF/VYbA0Pchign6GMoG
S1+WryulVmbxvkJRu2+OkBiNOzwSLFsFj6k5ONycYnl6GEbygllz0OOJhAHuVSKy
l7vHQ9RtSUTf0nTTWRPJRSnleOpZ/Hs0vCSOYp9z95XC1MlcMSWF7Rg48a0ae+sN
BbcweZ9AdMie2Y8DpNtgm463fURKeQiWCQjJQpi1T/q9mQKGO9M94yScvTllBwJ6
LzBY9kgtA5KazQnDo6N7NxUzB5I3XqQUvXy9k6xqxFr7k9PCwpMIn/IQ4zPvJn5t
qFKoI4IWYWoXGcMtPEqtew==
`protect END_PROTECTED
