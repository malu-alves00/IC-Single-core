`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GkBrJETXcwjWTJRBFlO0mLMYqw0AFom7h1CErenaykx2gERbHCtWSepOM8icgYOM
emCwd8Q20UjYtXK9U3KmNNLKv5QMvYOoiWIek2XMvSyLUZfUelahtSMzSshgKC7K
VRSueCScz6w7ms5N1uktLPk64BSXpop74MIXRZWgZGXy+2WPEQpeyjdzpDzvhzwG
flwUnSozzWt1/DnYcbfqTyXZ3/L/SnZ4gx5Q3VsRHjN0s82DUjVuDU2+RWigcc9U
tbXWGYOK+BYpYOp6jY5sk/ZLq+q2UDwhTpjteWxA0eKcc7O4zuGYWFUgQR/p8dFU
gB5E/nch9/7qlqnxJkELhHEw/eXWAeKxNOq6absX3dnb9gRveAj5SDfDeodbRdLR
Yax1wCI8k6pCc3fTNWAhm8xs8knfQB543EBibTq4rcArzvsWn7YQ8q0kN073vzgR
6hj7jzit6PWNS8KNV25pltW/QbwzkAGD31hMB3bsfO7aGSOVEYDx9Z+QzR3FpT2S
DppBZeHqZIOuOD0WXVdNtYL7Jm5jl6iSuD9blX3qpaE+2uJHw9ZTkjpQiwwYPgxX
1v1l5fF+Yn2vUDUwbPa2Mtu4rqnB3WyQbJq+PSuDk/MwhtSF28He2gI7kndtaoY1
SCcsBXIre0mNrvL42i1w/jOaurkpIGU/qhjrEzBc3i8aKLDSCiNgdbaGNY8jUBME
4EBnBkyLkarEMC1GUz9S+A+wsKIYCbVv4YLHKjj7HoZoOIbcF8bUJPJLAxGDPxPt
aB8Mtz2eywS+tTRyyEG7SdLUoAhCq02XMgq3yz7zsw1IyoMYFVSAwEiYsg6iPE6+
w0p6QudgzQ0m0iard8aYOEcLwc1hQGX0xB0HDRJUdc0XfDyDRhD8FRJZ9rDP4IuW
HYSk0cwg1ZefBPJ9znTM0KWru/HWA+dRZVi39b733u/um1XMZTjNJemchdtdTW9c
GLQWw0CqFcO0gEhr2nK30AHv10c5c+8XDtkg24FmmFbZgvRH89RBv2usJgi0xxTK
mBLz4QXIbF09WVEQkf351539aO8ay9fCNIobkxVSbSJuvY4X4k7m5KFwcugvHFcv
kJAYCd8ahKec/koEzZJBk/6ltIKPGMSAyDcZ79061xb2ddwAVjQCn0ak2farav5E
ZqbVaQSfbsUgzcCnQ1D7bMOv/I1pE3gitp4LDetf5Qf6D22V2G6TmbJkTQDim73q
LLCYn1T4JtVnErLKX1s4Nzy138ZaY3IO6Mt0p72HPl8H/Ekbw4e9p+GuinJ6bGVe
9t9LgCxVBGdPZ9xQjg3uHBYoowexAWH7AK8sRLcqyOfx+DPCUpijwLbcHQgF0Sgp
w6PJ06oeMj4EEE6sO6ZCw5lmeIZYTGMrSRsrhEmTkUxjc5QlghohMTwRSCWOb91e
JoIBqRQ791aXQYc0bPifh0kyAlEKiCZKg7bhkdFCy//VGM4wKoK8WogBPG3Z+tNu
ZUKddUFd75RcG2qkfB71+rs7LH4lH9zIJ3jlbAVtDo82Qj4ochZdHA1h8RcOxbPJ
K5TEkiYtxzjPuZ3qs91Zgg==
`protect END_PROTECTED
