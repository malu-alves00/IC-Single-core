`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FfXCMmyKkYWvWL54IyOtbyqwgUHwYo6R1TVHxNei91PrSzCnm1bzawOLabu9Dvay
ajroeEN24O321mmnmN3K+hrLWcvCh0st2bd1H0tUzBUsQ8iHvnAv4aSpen/yJANR
eM5jfb8LVrVxKzSTJzkX1gHaH4CDkuclHqmcwnWcVQ50VCpAI7iAMAgOTA9aOTA8
1OeuO6m+9aEOq0l3cs1LVBIHOerNeesyhsoAMXQJO8XTtWxCV8JV6f612b6nkFX7
BYC2ej7k3FCkYPhNHH06XYrrvE1zoogKbJYmYPThbf9CL+qxHsNj/10D7Zw6PbnZ
NFruuRs5RnSVOxvNWyYZG4cV/0JciEL85r5ro08Aky3cY2pggWgRAe2DWd3m4dFJ
yJ8ruhh2MarK35x2K3pJt56cFFjHSY1TilO2nPI121OULWuEWQO0lXnRf1I+Fk/G
XItFULR4a2x4a+fo0+OpIHUDcYbFYoUXSiTn9WlJTeEwjkvBjUpLyk3kH3tI+CKv
1AETim4fpKftSvU/06G2MwoI2TfLALikD+YLuo3OYA+dDsY0iYB4rKmMHOzrIvX6
wD6X02TnzumzK/rxeKAP4Rlp3ECszDQHFqxCrfpyGn/jvFERLmg2cPjbGhR9W0AR
RxAzVKeZmUmi8zDABho/TQewKG7rxWQvYMuceu6qN34EUl80vDyJ1q1JuYJEn9dQ
pFl09hUlq2rardml4dUz9cy6ZoZxbyxlr4dhcaQUQJK8PO4YmDAKMpFoGpRUDyzr
eksl+cIgpT9beiA1WWpT8RN2V6e/gzvR9ZuVRzsSM1nFnoDjgx7owRiBpyrszd8+
T6ukRSbyWF/UH/+jl6lbNtJ3obVNRY9o6j3plmvFayCN52rZpMqy6SIJlopcbdO1
TawkBuCAgyxkYpQjoenrIl8NroESE7ljOVTBZFqY1tHrGa2iP2NMxzZqTiIErL0f
MHeOLwApfRAeME0P86TDqdSKoS65gvAu0gqt+6YYnTfGzI4m9ygaHqNjJYTFXsUm
VgCeR//GzjmfaXgIV5WiNksy7vFN9mTu2oMGtoSCU3PUAUMvAoickSf0WYthzf8B
uNkIqLCfAh1M6SCmPj0Bcw==
`protect END_PROTECTED
