`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZIjQf8/KXiTVFmFFIbfSdlBpxRjz4/kUAeHb+ip9ZVartook/Q7hl5PtGH5+xr5O
IRhvXo8/ALtc9i5IOalSIrywLi1u6W/qbk7Xpc1Qmv724gsA57e5FbXrZ47rBMxu
myBhUi7l/wUtecJzYUxVKgJn9tOdCWHo0ULR7QRTyuNuU+kL4oEkjI9nuO1gO39L
2e+O/mQFTVovlza+gPZbg2F3tOIPaX/XEYSi7wdgSLCRN24S8b+si7WVHPpLrMjj
2kY+WgWuIE7jWISpbaCAVPt8OaBvXtkPQo09virK04F3pZDl5x5TiiVGGQUaKze/
jhdO+QopC+WAMvwL4Nq3V8BsenCwuICQmDt3XYO4gGsUg2Xqces9Df56ctnODvVN
FL778TCFL9RWz+VDOK0wbjOJqE+d0pC2zIsXRL4fVw3wN39oz9HCgwSEtJoF9GuV
MPkQ5O0K0N33O+E26db4IVVmKb3RXDVQgpnUDSCrrvlQHmSMCuwKU02UWDf1ud84
c7e4RdJ+mqrfFu+0HzUkcZsvBzmAruD/ie505QVlEkf/8UZqJcsqEBJiuTeQ7Cdu
Ria8ob4LAfkr6y55av4jPX5Lt1CVw15ir2AZaae2YfX/av0Ig93BEmLDXmRJnvdn
8lBGy9tJAPutMGezYJGlhHy1OQxXRh6y7lKdCEibyRnhXaYwtQuWINJdQ1Xt4WBq
ecLgX4gM8uiL97n1PUx/dVzbmIJzPY/OPfKZ+7MBV/d3beUFy6L0DUdIJlCD6HgU
Fxpp3shHsBTsnVGQJD+WR/Dz7FZzZp4WBQsnvyLnrU28z8PfO5rZy8APwOy8gmbO
xx9tesrJFfznrXJBJ7KgvlNwTIyyztJ4msSkP0H4ec+TR+Zasw+yFeoDJ0TM73ys
OTpXvHz/z2uXS61GGd7XiyN5lyvfL6He929k4JqCJsp0b0QuYIAaEOpMQf/cRdOO
kQL2zNmJfqsNwtg//2IN+vSDP3H46KNrQzAXwhckyFcfTCWJqggkmKsK/aFdQpSs
dQNVNZOytglgEZy5+DULz6BNZijU5Q19LDuCVorsG9T/WLA85+6SThr0C5wPz6ka
x2L6JF7PoEswr6tN6AkaZrsB5voCWuqiOe+rB/TKEl3Y3Uib6sYJKbPyLAa4ke5d
xroXNdcF194MKe9dYQdVQ/v+rNCVYT8uqA4auH1URkuGw2WYO86ORQBz5B8dc5/3
+ErC8yKx2oJGNLZ0KbCkinZqHz9WSL+dBzWiEegf9d3KH2QJCy0ufgK7KJtt1O2B
A4c2KEmccffvhpuetXr/ETKhe9GIyEhh4K9jVOz8sO24axM0gWGktMpjurzARTJb
G605qWjT5ge9hqWc7bDfCRvlOMnuwqKtaQp6ozvt7FXnbEhnjIYECF+dOawabreN
QHecuIf3oAb0V/iyzH3KQl0s03sbrRrWYJ5Z2eClcX6s0NpwxUS72nAYqy23ipr+
ticXX/embA7ZH/yPmXgAsmBmT5YqiVCEzU5LFRXGjv47tBr+lDrhDVQWlWdf74x9
rKDqdwX7zBylNT/lFT+Sfvv1hODLcua9r7tpXU8C93ZEdK8PjCMY492Xf+a6FeRg
CCznUmbGEPGch/pQvY8PWMa/2IOKa5xwG3OaIpKdkHzHkNb0XscHC+Y4kl6W7qw/
sKF8b4bDuqnMHHq4Feui+vL+7aqJdoIcpG/cV9px7maRmD7RapJmAiQSC2/MKWGf
8/s5TdpzthEbtwpfFfnUiXUFXlZZfbud/DI3SH1s4M0sxfSn7AQQYf6knIP2M9EB
bOefJNwcU5ZHaB9xx39YTROCn21DB/iJ2ep3C23/2bY1jIpwJZ6Rln0TMjgX8P4x
EUfaVgFmy3U6H3ZxAGsk4ECsCKjEzW0wlcXBqfgNr2qzaHQTVPAROivI5rJplAvw
1zx/B5df8e1jZTreDszVH5JnkxhbBzB0x1qp/BYXN0FAdxOQqb34Wfjts9r7CrS/
lIygjS2wKfF0WlE3rDgjprrftJO7A6Nxon+IXav+4FdoVwslCcM/d6R5pKbf5H5l
zCwIG1ZqQy+MQVdN35bjKZcWY1Wmoub1OdPR/YsVoWH/FQ8YIX/3KJU4hfRUHDBm
56ozcpV9r9a43diGmHBDFmRK3KL+r5/Rix657kdCCBNRweRGQBsrH0efxstKJ+Yb
V92o05mJZsvt2LREFH9e9nYf28PDdfJhbUP/5CEPRS1rS7FFlsOOUa0Hw7iQ3CyB
La89oMCEZlRy6fx63l45xLbfbLDPsvUvRygQ5jNwdWgdQ1T0mHZAO06DXG259AkJ
kULdGeju6YcmpI/FufapFyHPiErziK/Bhccdp+6oxVyUaUVrSnXhH9PKmRT9tR4Y
5mTzNB3REi+1NC7JRKaLh/T40MhyVYw/QJv0ijctG/ajFNMRKXeiZkmdOWIfZoVW
3srt2lkO3c85DG5teCsJjXqD2AfTo8A8BRRzIwBNPL2Yn0YDqhMKe8A1Xfkc/W4z
7XqQ44J9bgLzyweIOiYLEyMtZQTy2MshRZ/gme8tRSbD5cOyxzgDaOsYkfOUfubf
CpN0WZ9asI1tHL9AUjl1Fvw6SygZUCO7RWZPBosZPAGNNr18qgwNpVBTdxSiBQxA
n9fsIGsNHM0YFdgpJTFIdCsjSn+J7DDTepmMLn1Yi98fIidkOMvMQBYrQ9Bl26jD
NZz6iB6dbC+YL8wOSWKOiIVLmDBpuI7Hw5RPr6ORxF18UupFxBR07t7yc/Lim20s
NobEziH+IlOpowiwqzklc0Wj/bIptdek7KWrvyMKb0pXxVt3450OSj9yAOGgIcZY
BSWuS8opvT2YwSuFb/4I5gy2J0HTdy1M3V2p674kcUOiWaIeKhEeR48I/99edlmY
xr0VgWxMKtVP8oPC5gU2VRUTtl8al4cvD6G4uXacBbFoMS8YKf3tWsjv1GRvm7Th
3dzKlR/WkOWChIxFBJiXB6M773ugXQZp6FmkAL8VZ0Pdn0fbXvbPp1qmqTaVxAYC
RRaUbOoBXbuAeRAi+1IqVQkWYlpAp6pC6CeACxtn1GQ2NOiO+fTGpBHp2Of1ay4M
qdqeJwmIrnBrjCOHKwtR7N/1VtWZhcxbSITK49yg7fpkpCc3XetxyNn1syfgb2Nd
CxrQBxMuprMoKfY4TWjGIYDOY0gGqlzIS+vOeBe4PCDKATVTbXZceCpUTbi0KFpT
RF6hObuu6izfE5cUdyJpfGHrsN3CBF+lyvoMgnQDV6fqzsabZNCRafvQExmvMV+Z
twvmCW5xUVE72Y3Tfifx1EUNSAjJeeHTjDO63i0RCa2wQxeSu1ikQKRkUZRkVXr1
BcXAj0yfg7TiGnWwGcGkwIPVOoaN+KUhq7VdJYWedMa7lDDkhKIqKQ+U8a0xsJU2
3J6bHE5sq0ho+bXC96A7Ob4b5vITKQPnEEHH3yU3DaHsq7cwAYV6sSCQXrk5lrUN
IBbSukvrArqlMuJVUeNqODgWIdbopRgVksQk48/SHPuuDF4uEEyy5BmAXPqQrad8
dMUy+ftT56vKCl/ZmogM4UTV/LOGqa3orMwVNB0aJX9BDHklKCjiQi+VI5dX+74V
PV1KGusL7BEWZO1qwka2bY4vOT1k99PZKP7o+fZVzN2Ax+cb9YLhoxRBnx3rhYtR
ZDxeh/m32T73S1Ijk65B5oH6DbU5s47NMtqnZHz+ZKGwr6UjKpDp3cFk9PKqivjD
dgaZfCdAEGvl50VHhWqtarffipX6oqA92l7CCf6pwdaWZICGxXZwDHpfnVTVIclC
0fg1DdlbIZ2xYzkBU2WPl6pUkWRbOr3NpGZNkuh97fTNXyrCYAA+yoEw9IoafS2q
PFtN20YVsI13ooTZg2Ep+I3wOZvmzWEyTz66GFifVEhv8TKcruQhu2XYbycG2e+e
6A0yRFxzeen4oLOPYCPT1aMuBrvyvGx0AFegqg9j5zbltWaJ3JBdaOEt+xcIEOAH
KwBfe4laiaqzEvPSp1TQ9xn/Bmo+quzimz+dnVsksWd6b8E7x+PpNlL41l0L45dm
0l4gru10PWFabC9d7OrhRHPHQ7F1c7RGeaR8cD13DgIzn/ASA/P/teh9KhmIZquO
4qff2j1XLKQ0Ceh9hx1HTcIuLUgiHaUhSrSoROdT8aSpEIdpEw8XgYKmco0FqFhK
fdTUVr1DzmepzKKBkWWYQxKOoA+qzRmtVzEh8Hb1NEaLemOx0Cr9eSTZpm9Rucvc
yKm57xZiifgzQMmrtaHr8uFngJyQOAGgstdgGFnPGUaCNqekIexGVtUi5AX/xB8y
LXXl3UkrWmgH6VfKdhMVEoqzaX1Rr8XbJv9Q2pJ5RPMB8kdjtuKuFEwoobeOk5eA
GQ0i2OHdPk8Htxh/4+Kqmfem1/C+wR57IXWcZCBgw7ux4m5yjmaPpX+h0NO0etl4
5JxidapetoEdpv8E+chYS4OUX4XkAdg8lmFw8s1CRyjW/HshTkh+1cemBYn2ORA6
4EPh3g4xMimkx4klssWMS9wQlqOfb2WtXPb9WFIYbapUlKxLPIK5DBJEDUcnwdlj
KsR/19MeOgTiW9j7bZ5yMyy7/rch/s5bXah9AmIM+dQD6kQsiasw6E73tneNZ9Oe
/jjKUS63atBa77yCwA5dCh0/fRPYw1nawQdgQrkkHIz3lPOuYH36hzwj7Da/u0QH
Y8YNqyBhjnl9f9zY5qUaOInCrwYXjgfc+SS/Md615LSKw07DyKclnsdbl4EwS0vZ
VhhlEBunLgRyaLsQaiPKsw3cA0XCZPjhwsKMfFtEzbDwtVVrm3Kol1GkeWdjl6Ot
YevyI09yeqh2/iWNwWIc+uu2YfPdGtxk02Gf4Fi0UREPRTTKv+8zKJ2wC1/rP0MS
LM1P/m2ypk8msW6qziyWJd0pLGI+Rgyau/zYPMEwaakqBamQSoq+/Red9ykSenfz
l8JRiVRpU3TtWOX4ijSXhGaDC9nagqdNctJk0xOGixDzmJlVy2+xmvVJLjsE3yqI
ngyDixK81PIpLIBn7Rfg0urSQurjL6M1LqEQ5s3b9sb+oEctCUIurcTVzoF6Cpbb
tOgYdQpCwG/hD8dg9/9ysMs47d57hhfyR0kz2SP3tMz6k7hDzxnXelI+YP8e1LCu
VeAi2tHoZHUL44sHQcHkt4Ry5bW1tv3f6DrxWaY1/H+5QXQ3Yx2FS9KErF2rguyL
ajDBOoM2yIEIJRncFZBEpANZo2/19xQYUpSqmDSL+D8A13k/z7pmGjVjFwJcJjnM
eG3zUf4xtKvb3qlwfTsWT88bE8U9rc87WWaA3rUTURIGT3Rn1N4uu3rkxevrtoHE
qeqEKoHcQ0KqIngQra12iymJHHAP3WGMe7+6ncdA9BuETiBk+ZZdtF27O7JcsQ4c
clfddc/nRkW3vyrcZTxrAcCX+Bp/Qf6vZzUx5d1di8OK+4cEU7bch08OLESJkSBj
bu57FlowgOCzjuR50YmSBBGjb3NyfT7XTsd8WAw7kOLiS7cjaninaD/cKKNn8h49
4nvXavIlAA3nD/TDnS31zNSUmLCn/dOnp3jxMG8zilsf53ErAuvVy03tTI/pVku+
qQoJw65OjsDjgr5vA6pbE5wxpOx2owRys7rMvfw2BPkoO9neIn/D5cRtwl5wV/6Q
ptwAZOnyInKaQjXAcRIE1WYzF41bDSfRMHCnEndENL0+FFcQecFuetH7MdrvH9FW
xZI8wHwaPmeuX9fA99dSMHI7kSooO7FH+7Q5gCUZDIM/EfZxs/q0XNgIRLmLXaUD
ncMNMyevCwcAnvWTQBDCJf6FYaLd79qoO5BMIxBH8RXEb4SJIfvPJXG4SX7NXnzj
WeH93KEMJVJRSp6t2jcZhg+IsHk7NMDhB2srrKC1nb7zHP4T53h3AkCowgB/Km1t
csHCm/5O/Z11do+l5teQOycByKt1H60IHmyGDe29Z5Ibb/hMItw75xxeIIuxK2lr
UjOAcnJpdcBBDgmdZaYZ0/Hx+hL2S9JfX3nBRW7rD9S9M7c4ZVu0C6lo4t8NJvGZ
1Q1hcvbAvSYvTmJPm8bJm9FoHy4KiBK4JEJKFGccnL+iHOh/8/2i3fMF3GeiBTxH
GIyyf2wRYiotVy+/T7QdFht6+MhcZn4pgt4hRLsA200a2erP9vjzzHapgZVCDMhS
Jt4ZJUOzCL0Vic105SLhaWtEl0iXaBq+8etikA4+69UtceeaHicLw4klVqSIsr2t
CxBZQBdUOBSvp63+SWh8abONzyU8eqqbFvkSu+aAPfUVsM6LBMK1DnHHVSx0HNd0
ACyAGD3kiHVZn4zQdYqgMh0o7ok2NM/FwMJxDjPjsMN5Cu8j/aim2N3HV2H6lBWc
KodtKGqhESgQfZUw8e1zJ5Q/+yAbi1FO1Aqs6MjNYZJ2BC2WvJ1oGpMbiqtOxygc
48Oc7T7wGxx5p5utMVWqHJxfdmohvoVG4aaviYrNWfyuXkgFLFkHX0LAts1FYUha
kQclIDwR5+DRJAISxqYmzRKo1Qw/vbkAqOG8kFB729I2FYHVBTxKgbjlElIEUCsM
lE6GBCAZJ0okW9JZydOlo+O6/i6wMs3pPRm1U2dzBE4oI3VZ0Hh/3YoES4eeG84z
8Zw7SDdPwZPBf74c2UZ3bnqJYAYNaSsV1lolNbPPC/LgSAbqMVdkxym+9EMCD1HJ
2eUPAsLikfBDWBuKhLzA5ZXIdnPkRCKtRLYVUFcurzB1J95tWamF+InEwz7suO1f
/vEOfYFqMp3yJcWWGOzx4pAWz1bKS7eC4uZikGGQcskwqR6Q0WRbe7/tFvGNfY7i
5yNN4TTpyw6PD0yerRguQH0R+wXx8DcV2ab1DjcNAQ/SiE7KXR/WXFTgORqeegOB
o1fXpiuhn02bdLnwun9DSUSW1fvjO4/FvP6iN82ljccm6R9aDEsmf/AOJwsrLrCV
RW8duGJYvm8fRAlQkaV7wZYv5mMBo4HR7pIy1SDMKOkcwAxSNLsYVRrz+Ui6pZN2
dJcYj/+nGrmLYvvBnwbEt6vXrsicHJHvV9vqgWecYubpodaXl1pfmDwlmJT1kWkA
BOpp2GEU8QsPZ2u9K7z6utPQYGIuZSoC0M4RTvZf1seOys7Hf6H3yAOVhhzLYkla
CHHauoBSOIvgi1yqimPcyEBpkUJBM1JAGMtbxRyJN3AJV6QHvnRh3tnv1HvwxPdj
kCNi2JFSTD70IUzu4fIorlUe1MOBjLMfNA06v/wNKV0XkO9A6z9rRWt40oGR9kNe
YBZNbRrvbjFXdHlchSS+iJSjA9Rj4VSzjoDma5uZcGw0YD9Sy5R3fJU8hO1GnoG6
o2EcLc75ffEU5MFsf07u7kS/AducwuH4SNSEW3ZIT22kOnDQ6iHzKRoDSFfTsxse
r2Oojk2JZFBzLXWKhB+4fLDMMJtuT4e5yTXLYeSQ6wo0TIctQ86vBAcgjvINuVs8
7l8Gk7xAnEd5UYCLONZbFVD0owheJC+4UGcqfd+dYS0SAGjDzyy3h3xAQDJbx0Oq
k1M6sOMoVdEGf/HQlPc+ZHRRM0T0VIMh/G2ESIkxF1zVXXKX+3+CwXUhryjzL0hM
2XiqlbaoN42is2Oel/d+g9vtWAnjreO7aB6vVFeyNgg98dc7vR6K0ZfWPd10CfmU
Dl9s6MKHcKjstQ5PpBSe4WfGzjThCLu830wA88LaeXn+awoOF2+Mcq2k1In9ECDz
c89IPFufC7HipIbTvvgMDy033H3AX3EK3aT2+ZxHwLhosvjBGYjlGSYBAAudFpTi
wz9hvr/KHqnYtcqt1GKb5N8/gKYH58/lS8rnl0drUJ/LYYu+rLAlEcdzWz4lzJ8A
zdgSV9Uf0PYjrRU+NHKOjseRPZh9RxZe2X6I/GYuIdEUoNHQn8xWitL27uSx79za
dTLg7JvGMqVr0l5GyOSpScKtbu2LzeZKAHe1f/MOQqewi1bMHGEQpenkFyUo2h6F
rr/w88f40MKUKWgT+zydgKzpcKyynS910cyuw7DVYUIUN0OmNQH4rcfn9+9KphZo
P/d6y1cxAKKRP7rpWfP7QfZ1RtZS9f0COpbi5aHrCt7gaIW0d8/2WeGEjn8h4g6I
C/ZW/szwkXaqyYumJxmpivHuqkiC9YtG1Rd+My0M/z9VPP0JBOJqFIQ6MQcNLCTp
Sn86fjxZjF9CVdEskah42Q8RFYYgIbtXKiuWBf+f2g75sdui8x2yJc7P/3CiyUvp
653GsBN2+V3Vr1oXRwr0rwLa11HBrASjXnYHxeqvHpDrUBo6sc70DEAzysK6Y7XR
yrmuhzOx2LYc/NT6yQsw7YUkTOY2+vXvMRMzKrAo+Gn3/Od3XQDtoBMcAvq1aiQM
RgMO+2dU/OBz65gVxbRSioqGE4ugOM4J8IVZoO53bb1ZQB70pWdpFZTiDlIV/bFi
zwLenO6MjSEPFI+xxU6mKlBpJiF8o/DL8j5DohHokgnSwXcxfeJdjUaejyUeDBH8
iW4GNq6Q1ZdfgvWU685oeMZKCP7iYWyTs9+ULta+KD0NOvOk0V9+2h1icGY1/06b
wZvO6n6huxDKf263C6OvO0psWrMarPY5e0FxsUv0eufTu3mDU44zOws3XCZPtlyV
iOyX6vj3XOwTDC46KbRjfK0TauYlmoxLFVhChYvngBN87bjMez/TTrS8A33u2k8w
PWJSPQNlgq6LybYfvUTGm3rMiUQnWTYmFXkKmD3fdFMTLZS1uPFWkhE6NG1YQAbY
V5Y9eFDHktsvHbMtkuVbC7pTeTMqFK4LoPh2wO27vFtyeejEGRaLU+PYQugrMBeM
2YTEQhP2a1jqK0dztYReFQN/84bTFQ3FwUVCUdE+r6+V1cRaWcGTD1fJhxJMvZzb
oqjo4jAAFyl2YjvnlfbCYrrx0/V33Ie8Z9cPNggu9juDTenjT29T/9JhLE2y6qdb
oI60SFl9MXCdwGk9CdOmVk3loafbxtom1eZ/Ovo5h2NlUypdGZXj0yTyL1X6UTfE
gu/BhCKxHaxQO9Vn6iMnGJChaBtSWzkBXh0+G4vPUhuf/TENjjdBAy/gYuYSCNBX
pUC0fYPLV1MM2RvmuCOBpbXu+E9NigvaN+RPWEFYbgLh0/CF3lgLiJ+IPc8PjWVE
vQt+jegl2olmqvYZOEszCfBkLV/IppXIDh93K3XtlhUofUabbgEaLuQYxDZEAAtm
egZkFJv4k7ZcaCGq1GCIYxcnk1rG/JTqfch+R8m7RvJbzWNjZm2IkroTUHk4R7v4
AsknnV5B/o6Qz7MLD1wQ8/AtwTsxZJntt4feW5rKgxLkXh/8q3NZ7bhfzA/IlaaS
Yy8fm04PCmvo1/0MpSxYPFnpeGuAti79DgWelH2jwxy8oZLLzkD/cL16mq9fG5nA
ibrtfdJiAm7hlw0/AyaJZnC+EHeJtJXaK2cKJ8RYf0MP2cEz4FLAoJbcOx6g2NgK
U/xac+I/bNpcKLe2PD/rGFvIKQ8wi4cDW+V3UPf37f6ho2jqig19E/hWPOPw3Zuu
kR2DK9Zz4SAcVnOziYqraZBKBr2oBROI2xClvQVfVM/sCwMcGX801bVhFgwbUrJS
2LKGn7e6NkC7po1nggA+UtZlq3rEFFJHh08p05zzkWdp0CGxJbH2bWqF9Ru8SBgb
BvUj3C1ENltuKykPaVJ0ayJd62h/zNbIVx1VQF7g1LZVbQ6ctDPin0JYOfoTH6Tg
V+8xcq4AnWxKNpwppfsfCcKrhQRr7bWCD+LWUxg+HdtBCOjuyEspbpI15NdKbjkd
FqUp3IRQFqxxPsHWMDysyVPwglsJuMFcpzYmyqzB+Th2MxeuBJ1W7MhLacByAJ10
+CQUkWYMDLA0VDiISw1mBdS17h+UVMCXmZ60XlgPRU+7x+Yq9f8/ejKURWbWvKNF
VqQAr7sq0bI0vrnCaOc2dg/Pu2dk9IYnjNKVnutypEPDppLFcTPumMEniPB7AAH4
OOv4iYtSm2jj93zmtlogFeImgUgD5GIA5u/ssCvQlJglUdJo0cyl8XNJRxK5nirj
lriWfz6HUaywkXu5o6gd9+14at9gRVys6ofIpiVR0x/xOg40FBzWggNEtEYugDGX
5AhSM0Us4DNS2UUMZhQtY0XAi3vcnSJQ4tcRxW0y3OjhH39Off4ZVvJoiv/ouQGU
fALbVFNvDqq6znCxYUccfsgslwqtanHYR23WPICV3i8hxeuiV+maxCFJoJ1S3WIF
MmIDK1b0c+fQqjbe62uKHKDRsgTHykoh2mCZnCAeLsVfcWxEX9d/O3Q2SQ/M2+tk
QsxUnDSYRVsQJ2UqNcnDqlgArtfBlyEUblFTpfu4IWz9RAEFeufW8CcxRLr91fqr
hg30uTAzNb1cx+YU3Wyci23BWq6unCRnkHFoQBKpQ5pDwQlvOgSbtCHtx4s1xS/T
ftXCiXkHBpZeZD9NWmTxCiBeVDPqUBzjo+eadFm538vOEmTwdBWqZuBLwsWCUDwF
QwqwnpwuQ8jO+W2jpugK0lEfDvG5Iva1Ak7T07Aca1XX0QQ6JTIepz5R/ALxZYS1
2vX8FIyUjjdJq1nIvtzSWiP9mNJJtTsxVH+bWzeGRZ0k+CNhf9uywx56BKKRs8Xz
moKs2BuVLe3hhOwfazf/KQ0GZkv7OqXE7VECUlXgwQYsTq6nLepTv1qhVcHYsPxX
46HyxFP8ysRJgh9SItG+S+5z8RFNgD7neChGEJMvW2TjfUF/BNVk1HxLapKdjZyr
im8Xce3NhKK1l8LVxKi/TT1S4UUMfwj5wjtwykOqjBOvlJxZUSRlwN6ydmc5haYD
NJ/66SvoU2+j3OYLSZXJoesCdnEz9oT1tOT7sCFFOw6CclgxLXyTFF46r7WQYHZn
cBVp8V5b4Wd5cQskdv7w7bn0gT4OXOhbewPLee09JmzOGJI6ao8+5aj+mbWOkOVZ
6o2NW/7aAq3NQaxtrdRRigMRZmBImb7Fun5oVfxSpep9uj/XmsvT54eveID6W8qt
MmivL3sD2UdEBDgd971dg69+gQM71Vt2JIumkZ8BEfUpnN3wIE/0+pZ9dqzgyjIj
VDPO3eTsb3o5CCZReDtFWxNekuAmvxRRapLk0xtLRnPhB1G8KqnmRepF9cX+SOzi
TmTBKcK4fqsYWryRSMXvSajHNJUy991EuZB2NpexghfyvF6J2/CuI+Ptaz6RVYxo
wXntTw9OEgKovWClqrfoTJfEZtSfGEphQb1DRBSh5SCevGnEzDvrxXr+QAWb7vRt
hJ9U3qlWyQa3BWe/NUxQk23Zt8px0GkP3Q0oAl7sWqjyX3GAuc9eJGCOlxlC/jtS
BuHZ9nDWgA/RLwTIUtHlMUh6ltqCls5LWCpc6SizWqirwK6ByI/w5VKe/NFRU71J
qYbj2bifZIeM3dvqPfd6GCu3ayn5RlA2kxGqVZ+N+LOPKKs+wwE/hmTB+nn+vjjW
1tqsENfzCY18ZoMKt0YMOPz3FOUr8yosy65ObTahGvJUFXomC/asl0Bi7n99Pqwf
Lyrug8iBTuDFMluNy5iy4VCr5sPSN/Rrq0QkjrtxwgdR/kGi1PNI+PFZ5A6s+m3a
rAwlCgE6tZit8i0heVsaBnpVFlDhMfNgVYfASAzhULu8DsVYz67yBf/ifXYQcsDF
bT0VbM7fUtrUwbKsOm94ZDu5urqXHx//V5Bbt8SdqXsqZI3hfcBLc3j5N99Er4hQ
saWgb9w8gShVbijGw/RNTP8g5uGXfizjIFAv74gjj/D0rhNo7Ru2iuA+M1g0ZWpd
bcCXsB8JtgixkLk3IEclaV3zfySU1fgXwpWn5ZzVgjbsCg7waYT0SteBhujiUF27
5fJEuAN/gYM2teqbOLos93jpyRLjr5cHANA0mGZcDECrLdHVGMECq476Tm9Nc80S
8BCp7gTBOewe/+7jAIefFTBOYIi17cHn0dC4n62FibXt4rXzYUdeHRstFaLd9Zve
2lJxKpN5cBOVT+wUXv+8EAJUIzeBPLx3MiRMu25dEKMTTQmHeoC2P9fhzj+SqNka
dEhH/nCUvcV9T9NxLlcpfRQ/IEyimCd7yr4p8DtrwJvDxwpygXtvBU+ak3N7zxfA
/+rDE3quoKvBY5Yipv25BLYtYCBoQspDZ8VZW/A/3hP2giq46fGx66DY7oTZ0M2M
slZX+zx3mvkGW8w9CHVPO24NUjnFdHOCXEQRdXypKU46E+ycfnfGOHzvbBG1TgsU
QWZZHQ2ypBrbn3onbuz1fpLJY9Fht1HcUqAD19r5x+QDc9KfNHCDEBlI7BDeK1tL
o21u5gT86MKpJVtgrGCCKUjvnjANRhBPw863UfHD/TCb6dgpLr0oXtf5DMpoRXlh
QjRiRcHZuQCXgdv1zXAhD2uxPh8nD4LbEyWOD1H3pK8IenYcwiCHf7dbDriGDSoF
PikwtuRbe5Pm/BEly9cKK0IRKX/7GuQyHKHyoaN39bkElQTjWrMUwiAQ6+IWoORU
Rina3Cwfhx0V2R4T2ijzVeEAvk2FXvOypHh2iYPewP9s/zWxq+xiSHs45SecJ81O
8mRg2duew8N+3Fh6KSEjST2oMf/aKGryvMrr655plY8KZfsN+IHFtU5Orz+k3W3B
s412aOp+NlNzT7KSyZqa+yi7r2LeegfXBTazxPAVGnG5wr5QyFzKdDlc2Jx8OmDV
XHTA4OA39jG9IHZLtOvwCbXIF2rcXerWSDTi41A5wcUsvf50yE7HsokW5sijQKI4
GACdFfhz8aPJAdppcMpq9g==
`protect END_PROTECTED
