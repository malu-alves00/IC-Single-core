`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WXK62h+w1Eos6zfGIwwa51XbjXBenCtLXnL/5QK7u+ZY4conOG2oAc1APUr8UcsT
QVPhSJyWGD/O3l4cr9Ht/1qXm53uvoneLjVyl75W1yx8RHamFXUBMLC1C90Rarpo
iQ/enMCnuC5d3qMkaabHHGRRqKJmzqEDmbEvAZZZyGk9aqt+6AZr+R1EZqPt1eH7
uRQ3+ZggltAnC/M/WGkKpqzdqrEDkhlTe0lEVhaZnAJdsieklSUvwV4Tt5oP0uu/
ums4flftptLky4kju/Fvwi8yu2xkokHx0O5gAnuVcus56fborlUhnfZ4lMfQJct3
o1cUThIBshW8LuzOmfwFaAEM4BmW8KNXBded94c9rjN7gNgowl4BQK0KCA+NTHAs
3TbAP27Acf0cXpwhZoMWog==
`protect END_PROTECTED
