`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tDdYwj3HXtfh2fr1Ey0WaCeBP7bpDtrredugxPeXgU2akYeMQPDAElLHZaR/9Zcq
qb2v64lhcGGXS8vRWo1jzQ50iacLpMrgkNLCYKlBRbmIwKZLS0NBGJkFEV9TPNru
/5enx0LzvwRrrz42qNTCC+6zRtvh0GPDVxMMGgqhQ+NIySrauO1c0933WDtUdMki
iLvXD9YEsO3DKNchZNGLHDtIc9KHtYWBd7NzVVOCtolmMg94sNs2KMSMR8be1+H2
7tK5Xf3dQ3cknCkjiHQAo4sb9+mNPpXv7NxzWBXOmUUMrMd1FwSNg+KOVFG/oUKN
e34DzFMxRe0knRFw1k/x+4COksEQnxr27Wt+WKJhPn7TfgRQtiLN9gpW/kjmpLsE
lfNYuIIQ4DMpJoIx+WUTK5LwxK9RqERa4+1RNlMapg9N0aLJaOegQrAiaILBxipx
7k6lyb1pPEWdB2qAacTyA3aNzkZyMjUD9VAMZAwGffRFT/pYd7O4JRJSUwyGzbY3
avYQVqXeXuqDH4O9Qx/c4NY3nyrrhmYEGEA1RrWs4ikvM2HjFmTx7Nj7Us8C9tKJ
NIjRN8yGD+QyPw0ySziR8RxwFMqfsTGPGx/1rkhNLqOoC+fiAClYjwJYX3hOYjKH
OFrL2dVcS0p8d6T6nFonPK+NKHGA9GypqJqL793ddy5uyBYM0ihZS8HuBG8TUfU1
96Djx0gd69XjUCzFMkzsarp0b/awKXjvoGxSyOnMrZJ4D75FsUXfKyRV0pnUzPrJ
W35F51uLDXSn1HirDVj/aUYF/zEVWhAbdj+r8yweX9Ag2GOF3K2aaax6rrZ17jBf
jWvuJR36GoCDkdZiiv1HXnmme7xez/kDMphvRDyaEccG/ykgpmyMCPRBCBoZIWe4
f9fWMAc8xLYr8LNLmkPNpHQS1UDsidEK4DSotR+DrJ2Z+fUJXIA6EOysqDiwxFcu
qXiAOn150c13omQoVvirBhZLJ5HFTkrZhumsGglTyGk33HRVQI/aPn+tnqrPp/n6
PfFnVYDWCy6ijT1CIvUqEq5jbVt4v/7SqEUVxgSRJlxfx5TBUn3pnaz4wRz3UAzy
Upk4DZNCgKvMff+syOBXX0zJDFTYyXq48VmR3s902lZ+oqqkw9/NDwo/b1iP+FWe
4pqxXE47T6dFJ1ADqBosmfJvHRJAu3cWuCQbXJKmGkY86Bb3pCZjHZ3TGOdbnO4W
fuinOqvvwqU+5Zq4CtiHOMvQI/2WViSDzSbwaQ93Hguex6x8e6Qqo4iD3JgbiGb9
Ci8TMsR+Z08IN1Xn77e597QOcGLB3Mz73XeirnxfDrDMk7vQH6pO0Dark9B8fzMY
N1TJn/I/0s9dlrDQBIZg9ZnyGEwmB9dIV68IEnyNr6Fqp+I+ct6BPEJQpp+dwBh4
ywI883aY43MXvBhoRD8jQNLw8sENSPOZkOCCkS32rYp7ShhkTIfKd3pO17WDp7+k
MSWw1VpRYaONazbT9MgkrUoI4yKiEQzJISjdah1P3L3MpavTNaRHJMTUvZ1EDO1M
M0rxoVvK8JBlAyr5Sos8cuVV+artwGjCJgpxdFK50pzONeH0lGYPqwiw+2df7/gS
BnYmxg9KBIw240M7YZAY0+Kc/XTTPu9e27mv+51j4rD6OgXnh4nird2fO+PBbQ+x
t+3sgUy8Ct6N/13eZJozDnsRMWR6dgC/yblMN2Cn/rjawDi5mgq/2u1wAeH3kZNs
d/VTVapIK8wCz8UoB6LyG7on2TDWUyHk4r/OlKJcPsJpS4btrFjDIASD0Niy0cqP
qevNwyBiu0C/Y0L8dyaSGuBB9zmL7zIicpgfcwxPhXElJzAats0qZGo0BWN96eUD
9Qi91XNMjVbipM2YWpvhdrH3urGKY9U1S5vD9JogAz72p8xfSDD9ovFd6ACacOvs
JcgHU5um5gCYwYnUFGrt2LJpsGPWIaCXhmlsjVYIcSrzULhaecyn0MXDhsGzSm9r
3W9Ixz+D4eslSg8RH6iOJ7eTQGaYTAr1iMSF+MZ76IZSU4Xy7YnFIHCE8R77xv4j
Lc2ViaPIfWt3ZR38476E44nWJMWevfy1HtKhMygv+CjUlPgWxNttu2pHQIPHdivg
yXdjIVli9BeCBnlBSSZ77mORZEWEgSTqmRuKFiT5tI0GGwdmwHTh6tOQ/8bjXoZU
77OuTqhS8/cp5E7cbDXG1NOUrLa+MecRlQW3zLoJ14aR5L7kYF+AKfimesPnWx8Q
zlhbx/2KS4cycVINgSGynDKIRZfFJdKogNXJJmZFrDH4s4oIwxRQBAdgA3UZ3vQ7
J4Jy2QoP0N9mbJMkuoaYDuu0usNMqJ44B85ZdPCw56Yhz5wYLyRV+XYtfDJM08JO
gqhh87b0nJn25Z6jxXYpwHuJuuWT2xmcSh3sDTOkOsp3fCfy+KO3cJqtyAXagJi8
zp3bXtOfbHXwZVg9lRS6hkGr2+DuZIQ8jhHdazcz9v30SwlSRwtFwjY4VvIajGMU
nhQJOeD0lIvJC6qsbe6Vtr8BkYnR58ns6m5oYVYIFlmCIocg5ic2cAusjggF1upg
/eEtAMXja0ltbKfcSWK8fh+c9502pwniEuTOots7I5WDrM2E2N7dVwJ6PF8Gx2FC
k6beGRVHLwi71fmKyTZeWx1sBIYoT4p+zsoj5n2Q/aOgzyK7sSuucYe8ZjPC+Pmq
27EhqPv2HAcPNHUPhKU9P7lAae85Gq2KjmQ17nwhJJD4LDGzNWVn4INFLyUPUKZL
fnCPauQUBzukBl3uOMhnGO3Sq6onVkoHfV7LtB6ZCufpVfY/LVatVHQp1/lkg7v3
1reNWFG3iUSBK9JKmqHA3RhkK17HVULIQ1OJ6MzeNWby8sV2TViS+G+go0ShjgvB
sYWbcAv+LYbu48s+Hme4wzGqDoP7D9T3ju79pukAh75/bZFCRKn9NBC6whZX+U65
G27mdm1nJex0Acntk9Clf5egl8SLXrVGsTAFeADJEN3PC92lo97IwLJewF4r3Rg3
Cvu+1nh7vlUV99Agkiv1afHK0wOE8P40WRrwgc6XMrozZ94OoPUbr1vPrOF3FSWv
ysklwMtdVntUZKXnoVXYPG6laogAVImjuZJFnUxLkX1GI6NPESW/9wtD4mO6iDci
Q3y75TckXYp0Cw00gEqUakSon8K2g41iTxWp1jvnhKvSdDmiK9RiWFe/EWIb9paj
78iFPEEaU9h16+viGkILNfz5jB+bavBqWXVHW7MJNQOYyQnczRr0Wb+yRhPM1yWQ
A/OY01RV6K89nyn3Lkaxic5hOHROmZu+jKdrt/a0aaH/g1pVtMzh6+Zmkxl9cPKv
Leg1m83GL8U8df/5hiI6UCzrAg1xgD7yJbDekmj54cnKfLRPB5TitOxxtDhNZvpY
r0221f1/tlFbUpFm5flPXF+4V28LUIKo9P5ydz4l+pVMh9bhHyXmpjqVt68jgXX9
WYBwIaK4Rg2CL8CsnDghixTjnZyufWn/IknfaTC4omLzhR6KKEa/o5WUgRkUnDmH
MWx/3Ln2CjpuNW/RdNrqOyHUlwCkiOFmad3QMLRW/uZuj4VE1a1Qf+lDCcsWfUVn
pSxCv7lJLrjpdNb33vaq2LmTgzBVarxjlDL61mKcfhAwn46FYHMSicSepKd/2uzY
0ybqfhkeHv0/SxhmylccLcwbkfkjpBHG3OHdO1/f1aNpFe2sOhuy34fKqcdQSlvd
MHB5skpJMY0lmc13MQoQ5pCfMBhPgqy/MQmln4E3i2qxhuq/e9OwuA6ka6uSD/FN
9CbaZyfciJLfKiQEw+Mum03wqb+Jr0NjlYR6yXLwMnLIh0VwWRwLcpO2Pbie8u4A
n9he1sERHuZRfX3GmfwPsPW5T66VamWio1EO6fxzZyfPrNlr8jCien5L51ykqSgc
byghk97jmPSYk/wSEV2k72umlpHhxmi7s7wGN3JnhEXAndncajaXHFaHmt4GGSju
0w4roC9PecmTqtzrqQ+xpJsOviwyUaH6T0wLYyKcqNvd9tkJufJjrkZT+LR0sk8y
B6pVan/Npu89JKFrdY8CBSJ49VYnsTrL4uDgWD48kwtDAcqCvkUgBu8t/Uuy/QH2
oKWyCqSYQsmikHLej27E9kCfau9FY7qDmeefvyvpV3ewz/6j2F75NCioLfqqpSP9
NwDmZB1triqjZrbE2zcep2IDM7RSSzKTBn4kiy5PZjj7vbEXiF1Ggp7Mq0JM5tYf
d1yxFOw76U59RgCTOCBLLYhYloPz/Z317K/yonSh0nUo6p5V3sHzG9725hc6zcwp
p31bFVDIKX//62toAxFJYSnxYNpuCWYkHY7p28DDWl3sZcnXONIxkJplBXcxPwon
Oe81ZFutUXgQQoBzT0TUsOnChWSnX7X/pckC1HvvXl5OQE6p014YTVEyqFx2jWx5
P7r+gdUTdoPjgYWDdIjUU8jdJ5oVGkjC6U96jQQB905DyBpR1eIejMHsnAH7lFjP
U104SFGf/Vz71TRYAqHoUBvVoFPeQOkprLdt+2nsVsH15+vWM37RgRXjvWeP2fu/
0EB/BBQLwKctIzHWs079l0CVtyVX6HZRXVeKihgrRiqh77LHxUpfmT8wbTOkrxIR
YlqyOauHXe1amTZowzz2fZyoyuooqjWuLI345R/4kmH97ZwF9tXNlsc/dDa2QWTX
lnF6scT0D6kwVA0CBjqMNugd9Kii5D5sINMPciai2N7kzHI8doGMXC24cGpYAMC/
2nkhPK3fNM1SkKgKroqZixk1ixzPRLXb7nD/p7oGhG+jqd1jHziMbNZhiOX2IeAQ
ubiN+wGckHP6RMg+RpUAMAW/dvySWcCo77t5jDOP1jco8ALMcPUtbq0aiIdgcnaK
3m2Z5RiQzPjHJ5SGQFKnyCfyRkuDCJwln3E0aG2hVU8ytfuzlIJphzaWeaMb8lG1
30bk62bfT+I8gx78caZugu8TTtRbxTOWqKDX3w9ean3AMyvD0Q5Pv7ht2OtnxZ4Q
9dZfXSBWHKK0MgtnE6hHWsDJWRQUBmtvXXvtgBn3KQtsUvFYPjPeXcUsCBexF0Ob
1KRUkABffA6zOytL2e3zlcZiw89lj30RE+abs/xiAavumQVgmAtWpFglTvbOPwOz
i3pjAessAGRQQyjl7uXYICH4xz+Uuv5LHtBf/3rTBe/gZngP8CAt7FAZMcG1AD6l
UNy1OCRclVju1pJJ23XQplXXBjsBaSd9AiqDJh3zcir+8jkp3Bzg1Ee/7fQryyHX
pc07YacUtXKCyMrO00lvidlfbfbvUhNSHasnvoqheiKGpi/gfcEOi9eBLT5UZNUX
YhcrNLtE5rssni6FyNcY0ZTtlA/79b+1ku0PsyEb4ep1F4F317JbObxZeIPuZK86
wdnoal/al8wiadUu/UlDbofP1wq7rVcYHHQSbzV8rnmyRCy1yAq3aKy0U1UHDM7Y
vdBvshudiEoBsDY/FJvskstrHhaTJMKIVEWbweS5i62JjVhmgoFBojXTpKGsoZBs
c9XPtwfOQRxhznmsODw5Xh4ui3JAtsfbc3/7Dcj+g9/ysR/bXpHCwbuI67wPlNmw
zdv2urmvU7qEJ/GCHcFFkDoADL3ly3EnZFIAeZiP18+ImAUEOzkhGllO0f4m8m1g
TNsfgz3HeLRFrKhvAK4I49C0ZztRQcvCMTpMHjxQr5Yxbjr0O1MCCJ5ylza/BiMG
Xk0A3QaVblA5d1pnag0tjppeTomQy7I8Ms7EA45ijVV6hF7OQh0Enc2vPkKlkqzw
takj92c7Tjz1mD+2yBtlv9UmkaQn46KPjrlE7+yFqvuqVdbF8/htQ/RuEWhJ97nq
NxJzbdqOnH12zSGhUilMb3Q1AHackNCdSCKnzMhISsxFBWzINli/x75JSOMiNTg5
1RXTx/aorUjJA+ylBI7N/shPqa2QC0rtX1GyCbOz5lbV5bf+6HAPJpprYOi5bpgw
+RAiFu8LLmFb/RA8Gi8OPLoq/fVCaLW0uKJlkSlg0MLnjXwtMlXAKLQQ8a/Vj1pB
+DMi2Jc2g90sPQstdBXjgoA9kNy/9TSVfr5Lt2QzUJyMadBhGCmdmfXRWcw8N79/
EMj9RBCsgFaOoSR8jhrcB5adqShhsMOomWRvWT+ZWK7na3poX+j0dPLBob+92FJX
LnE3ve440YuB48FrOPhLrBFfQC7nT2qtRYH6r58V1RtC32jkb4DxTJ9MHWEoV8h5
ly721pa5xhHWJxfSjOw4masmuT/sJq04x3SluNN8Kzw7lJS9Fm68/x+Ex0jg1e4O
CuLJOIsJMCfxTvcVIYA9z8TdC42bQ4epD5Ju9LmPK+IgEZUm4MQGJeoreZOUnIw4
gmnOgpZxiOClDeGVKFuE1qJMLgELdydIqqDT2EsFhSsBxD5k3MyhkdZy/Gsp/PCq
aTF9lnRoEAgtUyPbjv/yqN/hlnnxONRe8y+spaNRM1n12mR+nLQFiCCqpStlvMd8
PlQzaKJVjlqbgy11rGw1zY1ujS96uumf5DMCBP3hnAbFYoBmQoN5ia/TsAwTiI/v
kLH18Mc2Mscx4Lo8fgy44oGCspSi+dHPVgKTtmat85CIbddH30t7C0lwIhHeJFpV
qRjzi4Q1cF0EPcwbfLRkVH8JL6HvaLT/h1LoRW9b7HyN/VrV5ugLB9BRLuvkylIl
vcIKMvJwmeJTvuWChIXCAMVV/QlbA/S1pRVOAF3r2TW39FjkiFCv5hczij2sYJtc
2frP6PA9pjyf/eMbr02kMhE/FWBloMJEEtUNKM8T7QK2TR5RU7OL1RWzcOmNrYZA
3QW8SGhRYET8VQflwmHq7O1fZLyOkPP5nSFUA6Rnfj84y9UVH1aOLHQ24Bl6Zrjr
V9hPYesyxTbCAO6rcaoaNY++P9YjesMFau4PT9XqKI9ugRxWHhhFFkyEuNSwXAZg
qoJRmVu/4UNrJVKytiHJPpEy/1uL/yzG1SUZvpXkU5ddH6/JRc9zWF2Aaxrx/9iT
KmqJJxnA5PKTpgohKDSedWaIcLv92Q8h/jQKzR5QanehJQK/sk34jS59vWgEaj89
db4zMVzeTuwEe5EwQrfT+sI8OFrOJj4YUyOPLN8IvymisMdjTxYkeXIz21zoX0TG
s1cfXZSbHHvb6DzQoCyrUs0+MPOwMZ8ihINk7Rk1TcBEJQZbuV2EArpz6ezAEcUC
/nYyNt5kY5lqMVhoDhDmhpPE3WExo66KKX/tsdZGr86kYCEM9DxVbfCRJ5i1ZYRe
YQuW2YzBYY7GxzOGSpGU+bGDVdkQOct6+b0BugDHOqX5B6tCIzkZMMOtcZNmYme/
C9qbkYpRNv3/RYx0WGeDkmKif78Psw7ggIbmynXk14NialmA3Tr0tZSYbCVOyXaZ
UBC31KVxrBDX5Bpt7+kTYQmDSknI+1XhNES0Hjdj+gwCjeZzcK+sWsOiFlX7html
g8+IMoa6Y0lKv+wNdU4WaRkz7XxLZgwAj5ykqOS48DBPGdlKtaf3q74HEKeZV4pb
oC+eMhc4NhKJmciI3ElCoLx4uyBsZYrbM2XJgL/MDafgFu/uW9jiqX4Z/ANkPh2y
EfZDsVcYq6kAc32QDm4yQHjmqmb10F3CmK6GV/Mp4qZWrSfNvtBQ0I+117bZVUCp
bmuMAp6HHQJk+gaT4v2QN3U/sQMHmuntdee843+R4N1VKAw2Xts183IBtXrCltSO
0F9fKoFYPQhuDwQnL/97lIA30Isy6MnmbCoBlXXrXqmEPwumTXiMJ5NZmxJ9Y4pz
n0B6YpckRE9GreV4bxWMGlNJe2OY72AaHHt/JC/sAMTuyRNqSBUD8KvwGRKD7MKz
MIZz3ZTN2E0Erzq9t+BlchsURUL73jUqxL1IpZOpLTUteJnc1g7u0pSyzGSlnj4x
0tvm6OkMeG7usZ2alQ0hhr7AOXNN0w22RSfSrT2WDw4QR1HscCgdW1OmWHwMJMSb
AdXHuUwydtDk0/bQ7s6v/1qRPEzoq4r3FM8Pt0ptNVHvRZ1KGQK3bQQHxlE5HtF0
4fzxxWCUntE7ESaHSvBgKBltvyqETv2NQddGpLRjj/k6hejTiTUBb8gGIJIe3Cjb
y/IXOR2Ou3IERx2Narne8APqJaNPwx1mayZGaqoRwlL+iAKEvoiMyIn526W3Dseh
QJSU2ZRLo9ekSVX2n3nz80V4BVhk+dhGz+ESMv770T8hSvDkfASFMhgE94zhobsV
9/IwXM917jFXv4rvARDIqX0ExfyponmtLjHD7yHVsRrgtDS9jhZMeyb/WXVwr1vS
nM5CRr7gHUC0rt7/Js7icEiiAvXnkLasoLwOSKEG1T9G8o50t/h0xntNT2VrVM9w
NvzUY+z7JSvOCnlQOFO7jPlO+vT8DU5nc0oim8a/301eS9NBv6OSQ0uVOIzAEjOl
G8WMN9mGuvjB20LASH1QUBJJdDA/N3tqftJeucEi28Fjj1oRlcRgbDeXRIBap0vs
aK4khqjqLvhMPQxIdmT/tdPkecY+JFBKJrWvi1tG/4MMO3wmIbbrxtBBAzqELjmc
0UIIgV6YaAvytM5JggsQrs+zx/9n4Fqt41EkZcHNTZ6nB2MnxY5RWIiVXGjGqbOl
07LlVmT8rFCBKpVDUubmOkK1buhZ/klgbYS/OTzG+yQK5gt6TwhDdpn+cBMARsDJ
tRZ1JQ9wlbfGFl9CfOzyqAb+gnXgvEaswEfwpKuXB6im4cH5AW0qPXXREZNyBJX6
r6k+mBUf0xRw9jWiLyIicumETcIyHb3wBRmFH1R6VnkF6kGpU7Ujb6n3e3ZD8i5g
glbvDFy+qNIAoSDD04ExpdS5ngnZ5OA1DfdF51ECqGtN4LCLEm70o7mXvNMz7lpd
lytbxhub07TT7VDoFEQRe74Tu/wLZCdsiare/In/JM/mCQK2smyUNcl8jCbvgDZX
ZamsFKzejsPZiP0Wlsd86ofJgPiMrflrOQzSDRyFQOUtas/GN/sl4GzCVzliGMFY
IWuLsIlcNTprNOqu0xH0Bc8XetLUpbcKGqCOLqlqlPtcNf4G9ufp/lonQI71U/o4
EIZ90ai8k/LoKfeYNVWZNfpvSlrIP36VzkRkKpRAkTmiOGylgRsNwFBvzNaOUHR5
adGUuraqgJH5vkKzqqTgV1pUjDA/ntQ4bXPy98YwJ7H1ILTtOsZ+8aJ8ihd5Yb8u
TwntyWMvTki/VCqnzq6wtJfol0KczKW4L/2dF9ncJQ3fRjnt7IFgnKDES0Y10OnL
ajGDgYQscGsEf1IHt8e+hFEwuAERlp+EbhBw77KfC+ybG+zmxWHenJm8Y6h+Wwpu
cbQswdva0tzc+uskNI1rVDx4TQUJQoLmOg8TkB4NeBfk8L/+RTxwzgPpSsB1mZN+
WtKd2x7ZSmSc4U6karYOOWzTCqfr4KCYKov5W3JYD7mwmPPy+NwJpy5yy5vzEXqe
eQ/NvdHXBMlyo+bY+GiPZHBL0a5VUTXeMchCg3l/mC/4ZGtrBWhQTlxJMBgHvx+h
H2GeHiJ44nU8OTcXt58Qobl/fIyv7kT8iG8RbNx0BiCZNSf8/K+8ZvunZPp8zXPq
QxhKhpq2oQ9rovF35z0QLNsnnJGMCJQERsaWq90aGb7LF8f8vtgKDA1tRnspnBaP
2ObVb74Ck5Ry7PV0QeisnqRnew5r+ZiURpNCdxDfHBdNKGnVJmnFRE35JmDHac8x
VaGu92rnizfbLJDgzv+xQb+aD7DPYOrKo67f37ziKsyZUx5X67rFvsUKN5uAOgUt
QnGaNhTk+UgCN+Y0dCCsZBCGFt1NyKiL8NGNvDA0sN+uQ1V46Lgqkbha05NbfZS2
HrkehJK+sEXaQqfBGg80qL3rBKQAbQ3ZOFmIFRI9KPO2EU0ENNSko84SfFCfu119
kK86TxUTfnQH4gFhHUF0lwdH/diPi45O4b/GvmabOmd6gHN3tBlEDtJ8mPo0rKja
uzp7T2N5dczOfLEGpuQHxQW+rFbSbCk3LJPiVRNTvf8rnPvB+pfNsn+b/HVLPtzw
njCrsdyIxh/r8QpRT1b4Sxd8aUvOG8giX52hlDyqvVm9UYHd5qQZR8+WjvXgDByt
pKCgm2+oc0PpXJN47vbcjdcrCgYDWzaHq8+MVu1ZVCOIoJE93Umv7VS/aWF5IND+
+l63GfzxvpaxRAMWm/4m0SxT8K9AP1wMqFW+ZUXBNK8oUnbQP2s/C7tL3kj6Ifkd
0XnSe7kUrZe2yYzDtH9SaFygEUzNjzN4DbvU5BCF4mRIRbcV4pjH3Y0G2SX51wP/
WSLERypCRDrNW/RkGV5iDBpkfrNmvnQuf0QJQD1PpSZgmGsGWOUGZNjo87UfU3ZO
tPlFKf3ycvlba+MYsvkgvXsPhLEKSRMumNU9ge226FM7ARing3GQt3NeifKSxoyj
QwNGGvoIG5+OwWBw96XaoyvP2iJTSD/QF5Dz05WK4bRRez2263R6kRbCZgMM8qha
Pf5Ir0WCqwe8qt6D7hZHZZL/XuxP9oBTuVYdiWBXcc2VtYCjWlPQArK+WboIyANI
oGnt6lEnhMHiOpi+r7DOZ9pZmecHNpxzsZPwR94rg7MzcruFWhU7KZ0akgrgck3g
s/fvTXivG4hNDNdZ8FoFzGy/10aICKn+kWLSVaWVBNouFIfUVdAfBlxksPg++0lw
4QQZRJHTiagdc7dQEtS8YHyWpW9V8a6hK9atyBTbYxd7YWez3zFj2eWZsV5xBgQT
sFf4x4h5deVEIJDY9W57Ow==
`protect END_PROTECTED
