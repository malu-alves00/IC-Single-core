`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3r1Aro7Itg6ZHxHSv5L50lyEX/P5uQAfYzV7BTLnD6SSDe2ZMccfMktSJopvtSu+
FFna2A4ayaRKK8RSqp1Lu5qOtc87Z6eE/VTJjVlVpB0ZONNlbe1uh6dK6bu8NICC
/13ojjKPYLv54C3X1GA3waTIMZxr0+nRdmUfPfFRAhhUZttcaxR3D8P7rHw0+cyw
8m5W3Kagt1SinC330/mD9IVpTCFQ/ynW0QKoHZr2shiVJ+/Hcjpe/kwzgaxPHao4
x5FKDAl5MLb0GR+qkS8D5ue+S2UKj6tISrZ4SVPi0lnFlHc+nX1HKg1Uh2mIhX1W
LppBDa5WRb//sQ1ftEq0HOWkErGTQLlDOv+0O9/veok=
`protect END_PROTECTED
