`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qNXEnO8TKykKs1n8ue8+2Kpo9vZc5dPmcRmbTyn/qA+rEZm+cHtuHawl2aoeYz08
Dr4gsXzUcoo3YrJDhTyFWfCb7rr18xWyTa7suDHe4yqyLFn8LrgtoPM1N+7yo3p3
wktfgzGs+uJdP+fqpS8wzLO6iwrWIVeuRGC9c/xA7LfaR9rxIgJjX4b19F6Bldss
fa2QeQp0w7H9O3jD9qBbplP5OIXLQc4X/t0pHVcS+Pjh3Ev6pXYcJlGq4Cl6vlng
QMjTEGgoh+ooaPghEXX7Kv3EC7KNzi0v/pIAwnH2ThaZDzdIDCiSOwbvni7gtXcd
OJKQL0KuoYNRr/q2uxgRjpIG2ivBZ+8u+CQL8BwfknmIG5G4XmYOVZtusFLF9ztg
n5ScJ8f0TzDd/22qNQhkq1imnIN77PgA5Mieuzj/pB9g+7Ffe9f8p61GdpQCJndS
I0XXPNYzw+rs89VjimLcVwORURjsGIGvjgx1RMLM9tp8gMmyvjEW8oN+f7CBexZM
FkM3w9EYQ4YpMcro8h+bHwL2VB7QhEVY1D+L/Aqs6bKXJAsBIlWXnZicGa0ea6eZ
gdv/Y1u25bw7SYYBGRMrbEe8RcU+rpL5jDfXIjXUFNJsMN3faLLT/hyNTKirMaF9
JaNTxgpi5CSMzE+3gWuFP3rcFFqL1iYUmM6L5mUa1lSIPgp0O82uuZfDmm822eCZ
yGG+mtwoJJz+thPG0F7rXhPDF588hbUwqlVH1fw/huMVUpTNamhWivWcp9W20yJ0
CRNSWUL8Eg8PdEZqCo3XCQzPo0M+djlmDK9LWYoQEtyvOadcZFF4Y/sD13Pf58ww
K/RkQO58oZw6o7VPvj7OQOljK9YVmMRLVMMK0xFK/Zf19I8AQ4lSUKYfPelgf7GY
9cmeJm9NJIfREySWF/p1WX5KkXAaQFsQhKNtm28MPNjsNKuj+fVdqHgX86IxM1zb
YHdMkaXBnLkrwBVJyaSEnVuSK0FD05WzLjuCzajpkPZjLWnIAYxUVycpdI9P8PPv
7vxlIi+ZwqbBNcsSPbO52Y4DRByovbt+k4Zk090MmUYnUsdYO3nMLc1FcDhrLB/6
RFaI6AZWLpx4jLAXeUekwXgRvFBvEL8/Tw2yJRiLiO5Dbia78tIiqMIXu3eFER86
4xUAjZGIh/+PEif1zEhSJwKlaJwmJpXUga73Gz7bypt5OG00blI6V98zbAxlb0RK
h4WIRMGtJYZmZfBXoRKJ6tc7zAdQItK+akUsR03vQFy1IdxaUXc8UxT4tdjAnLgO
0fh3EXaGM2wSLxku1bx5ZudjK8MAjoQCzKWouBekdWd3vkZ1divoQGT+jU5kHHQU
AEnPqcibG38V2Fgiu/6+uxpOGqbFrmuBCa1c6vRRWUqQmhRCTSuaGUj/+Ql0Oxfw
1TdQ1O9qbRZ0UIZkNV1XMbhLMZNJ+9vuexjaowNetEUY5/0AL0VW/s5PygIkbsEv
LsBl5klWO26RhW7+bcg4mkbFQsLMKC45gwmWQ87pAS1HfavKOk+Jxp+3+RSvkbLd
O21UFKZ3nSF5MnvIbmdV9lVtPQLnfW15zx+o7cqrtvCFbUxwJ5vUTF6zJuLTRlMe
fjDXe8NkSD60OGxUHC2TjyOHVs517rLIZz2Zg5GQUGxkxlXBMFCbn6XTwtEcxeFO
QonKcRhR2pZPnbI6vM/a/oaA49oz9di6jF6+0k0iby5TgybCHlbZH6rInVFz8SYO
XrcOAGtQSYzS3l286a+pWQw3QiUfB26GqnrsZn3hNL0SsZqCIZ4YN7ZD8zBaDvp9
9Uzj+U2l8pp7KunlTklDXJTk6UNSzKSs0yfPGQVDPfbQu9Iv9FE9dJgLXiknnq0g
3ZS0ETZ6EE7gB70brYwIL5j/YldMjvislCLIzePp5qbBgtjEUcA5++u4F/bHy5Vn
j/rbi6OthnsxSoFQHDJ5B+V43QHDwuifij3AOMwkJJBRcpVcqQpm7QgWKuHLuR48
zfZ74qWZCXfdc3ZVs4LGTyviG7T5fRHjr3zm8zpcIgT52h8bS8J3ShPwioC/5Ppe
0NbxeFgUMKjr1lvT5g55rNvQnL/nYKawXyhCHTzygFVa0RN/TSshjCx1WH01TmNE
`protect END_PROTECTED
