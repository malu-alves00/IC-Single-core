`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gB4zCbB11gm0uiasPZyLf2kegrf7lteeELs2xkE1hmrAHo1BuFM9BrFgO4LC97vC
Ks8rfN0/b2d/SXUw/kaujuewTLzx9zKmV4LEEj0aFizCYIefV5XjIGQnHUU1iaBB
a3oaK92UnXol00o2Fyp6jnsGy4A+h8q9ekzKR0YRGydC9eq51nQpgaHpV05OiP+z
6wywVtD5fhLLFbCl/+JsqS+POjjbOp3vggPmfXW2NR0/6JIxD+FctPUgX5rnEiFO
Dw9+lvi0to9CkBH1s73UMrZ8A8bESGORvOtMZtNmXsGYwZ4Z9oPtgpcHGNqhQMpq
m61IDlyiGRmoCROcUvv1qVN4EZZsCOlVAi8dW125bGo11rxlGcx0AgQyBVzNkIxU
o5Vt0fmFFyXVUXvI8vl0aTYVukS36q/6EM/a0tSHn8U8XuMpCjJ3qVXmy/9GzwVK
MWjj98IdobZyeu7AYhesRIScGkT64NrY0ee4x1S19NKeJ2b72uREb1ycZpjGhxib
HckQo/wUF0Wy9orBu04zbkqw4CTZuP9y5079Rd5hNrsOhJgyp75H4dev1nCeoSti
1yGp8VutgpQe6Dkei9o9H/Or4aHTqoBLhE7NeN2redHP8Nq49msG6eHobqsxI+tt
LiQPRzWVRJRb3qCR2V1wrFRHMMlB0mLyqWR0q4AHfw1pe0/zZSwT26rvcKW64kYe
O/hcUSntAii87oyiPJ73KAGD4ooj0xJivrj9NPv+KL4RvQKQY3GrrZd5nb5Znd6h
FtQw2h/5/8bwKOPUTih0IYSV870HjxVauKXQmeUQ+vU4PVLQjUjJZuygY8XEEd5B
L98v4Qr8fnhfdmd9XDtwqGts6SudLVU4tA71KWheY47Hbv5wXcSWWkwfZoNnfDUd
`protect END_PROTECTED
