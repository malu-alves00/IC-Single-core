`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
l/hnSDT/t3pAiqgvPGxGkBohfjETlAwTZ0Z0nWN2O4uh0cR7ChRAVEWtD/7wgcsD
QXXUz9pPjddF/10FbzRgdg1iyD3V4M64dnBfdycUitkltq5XFQ2I1Ir4BlnnsOqg
MUjpKhlA6jyPyhPXEKd7ilEoRRJcIgrvDH51asGh2xZyQNIcA9xHQAlPKIoVp0Ni
CfZcD/jJZoa1FyIbckmvqVNTyZQGsokDryxZybVbSOxQZOcXDcWCKiHcVa5NTuYL
xZpegUgH/TKzCcl2eAFXLhR19jplcZWHNgCmkPWQdPHhzAP/XUCyC5+KL89RMQYe
yLoIkMPZUoWRcNCZ1qJrncK4eZa9Qd6NA+2ezS9X94QvAvTBMR0i4vCjAhilI1oR
ykXJjw7qwgpF6UKoX0oX7/hIu3GsTcYv4skyPOuVakM2dbWy3LOMm7X4935F0ENz
dNPQ34r32v9hSYFpcQvmIkw0XNU3Mg1qhXnkspP30Y5xgSql4sDU/kZ2qxdPR9i4
BxlfIIgb4/lJdWVeNHsPlWcsk2qK22p1jFcTjbc22+3lgS8i3Tspi+2p832vebMu
n7hQpPBGmiJVdcyLkR3BsnqOpk62M////URAuehFSF2r8BUbhxZim8gbIpDnuS5P
YVxqMT8Xwzlph1q8UqzD0UG84O0POd35wVq91A2U0gqw1rPE1HPHA/95M1q7rlOJ
kjvaJstR8JMO2Epx1NySw6h885+oL57nGUCIBqYbwlE0bV7QRypa/WdJUZruwNrj
7LABwAGIrUndTvMvQSOzb4spz/XylmS4gfLPIeEt4RFCQKS0gQCMAEtra7PfINJR
oj+zdTd4OYvYM3Ukx8FZH414gVxRXKdosmwZQ1E16e4=
`protect END_PROTECTED
