`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
82lVooHZ3or0MUIEgGHURGvZDr+K+UIOYvhT7MoSp+o77wP4Co+CLRusZppTe1cA
bWYiBXN8j5Gbj9+39dBZTHLtzNO4BExfHee4DR5FDcw+yZoKwJ2EjDrKtDwk5SaR
esAq420foOmdBvBtYFSt4HU9s1hZpEWBkPPreZ4BUcJ9xVAqMno6O8JtEnYb2F2q
3RQnaaxX2CY0SS3T+NQ/jrt8SgeKRzA9MeHD4+NiRfU5Fny8R2nE5UbQWdL8eRtl
zliG3+k2YW/h9dDKvb0xeK3IeHIefaG/33EK0wefneVmtrGxnpyXQSyFD5DHpreV
ezmQDuNMTjyeXSowgV3pyt74fQCaHhXU2xrXFfrKn5r4L/ceBjsWx+NkK0c6ybYp
29m9J5q1TgHUZbLyM1I5aqzZiYLRCJvEKZTyPZO/eZgbRidsB7gZnoXg5LjUy4uL
4Dv64B/h8yWb2wYh89ApyDNST+yHHFf2HSG/1yU85mFJYx4TL9mi4RBYi0E0TNY8
VdeawMss/IiW3Cp8n/mEx9U2wBJV+sattHjQ4iXpMQBrzO3Y4KhZLW2RxVTe7o8E
Ep7plM2Ai3dSA+/JmFjJQTedPS7xg/yonWby5KoIJPRG888fh6a2heE65dJPrL7m
8eIjgo4B991SZ4QoklDVEFSeWHX0xKE79rBuYZsuzzgAqtghDRF1rqyQIv4pvUDk
gXGc5cHFGpTqBJ7y4nM4q0z0TucGAl6zNr2PS2zoeRQRdHZ+839qD4id+ooDRP7u
O7tB9OcfG7Y63DLdCCmVnLlCbuVUEasL6shPuVcsxKcDGl6O7RFxIAupKQ7w9hfq
`protect END_PROTECTED
