`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SUcW24JnvJb92ENor+KDa55Ott+5aE2AtJ9M+B5dB5Yrbl5vOJgTMN2NXGkJ2fCf
waNKojIGbH2GSmIR0pLP+1zxpxmL70djzLZaYZmO5meDyh1xx+eOVYvvtYcG7I6n
tf5KqdL/c9TkA75vsnUmOEobNMyo8qTeBrIFmHP94Wygb4DorGzjd/oVRuvduTSb
PnZfUFS2hJtfgdZnls17na7ClBtMQmH0F8bM3S0SQjyxQhXrz6/a2QEn2/YHfQj4
FESUl9CIHBVudeDE19Kpw2RKfkT27hzEc023XkLYraEFYVUIoZ4xVSLt6loO4h2V
+Qymo3OFQsF1fvSCoeVmEgv1yXD/lKbJm7Kap4B3XTBElXIsY5caGnzM185uqtPu
EJS4wR5YHoSjDYDQQkXhb2V59df13JGohKnr8aEqi85VQSNBfLGoS2vvqNmTjc9V
nam8fdXfOLz0zuD9+0G9TlMeSyZepZDgEnePUp9KMDURWThE6T19YyeOHGayP5um
1BO6NFCDTHaszuj45slPSsKPN9YqIgjISa8lwHJ/iAPvOmD1NuzQoJxM5KoeGbse
ptEPBG/qSdSv7+ghYj2cmyUTJk/66mLKl0JKdNW/ixBtjCQs/F1ybo2yV3tk7qfm
rs5cyAwSZ7ObJ3cvSo/DvTleuwkyVBrYwgKnjYuDhmWL/8YAuRUoc43lj729nknZ
Qs7XFcjpPXJeJ/6zQHg6lOCm/g4jvagzDaJmyDxqI6O3dcAMyx+Ah+QXDKmpTbH8
ARp59khwWn8amrn0Oif9Nw==
`protect END_PROTECTED
