`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iYp+ZOHtlS5RlL57mogec0+qe7kGpwLBjsLZGWCuGu3FW+9DLA+Cs+UqwxtJRRPx
AqSQFfUSf4BAf3qZTzoWHuo6tt8iyi0nDLh6ax124UGDRqU0OXNT8BwFR68dndgQ
ljG2mEfAKMOnq5GR+uU73QPx0u5485xYkK+DcffMCEbGmuzWUVUyNkMux+3WwM7I
st6U7LiZIHBNBOYWKsNqg/tToPys9cVMrtoz2+14cQpZ70bPQBnPGwZb4viAgU0Q
nNtr2snAAuFA5B5t3ZngNp7wYeALLHtRAfzphDw2QhmPM5tTD0fHqNT627DeJZVN
eCoRbdI7aDf8bzdg028QZCHet3M2uUlWYyV1uZAwkSBvYm6fFxY7CKXx1rrANVXD
1tegNuiQDk+JWDcVqsMgDQU+BSY6S4V/eDlE1Tz6vW+wjsY3ZciJ8hpI922teUWI
RUVXjw8yBlrcJNbhTgzaJlcMeZ4LmmXLdptVg92rSrdjy32eyH5z3B+1RStOGR4n
6zN21z7Y6rlFR9E/3gcVLmxS8btmMc8Uf23Gd2YlDR4c/LBwWMMqcj6RUCuxzO+o
Q+geQunzmSFcTs4J0IoiNxKFsYR213VVYn5GQTS+bw3XCNGx7teBAxBmcibmf6Fk
khDw2ghpW5wHhEMgV1d37PkKrtMafMkq9En0Lfs5SQVw7f3x4JxIe36ETK0uh9H/
sdb4c5X16VCYV4jT3C61qym0wsNhgisdCo3z+08tPNTKphMFrC3W40NcScuBchPa
EtQJ/Jg9HN1STRq3NOFCiuz6Zm9f7Jiiexz3AY1IJW4SNSIbyxNu4VlfaEzLr2Dk
fPYpsJmCQ7dCWOGRmECWobtjctGs0HDkhSTOZYquhwF/qRv6oDd40cXVDRVZ7sKm
84g8BK1jBKO15ZHQUsRXSdzVKAycVQQewpd+Jp2fIi4O9n3LEqeUJLOo/MVwuum6
Ai5kvUMbiLEoJ5Cw+Sxm9ES+mZJYj2ZFS1Dadv4mrOBuQjQhQOrqRCq1zLFF6Dao
iHfhBJ6BXXm/2OhCy7x8nTUO6vSH4WgMFIFVXxP61gGiUzjw58gLI244uFQLwMIh
bCEiNiW5ZooLaFUaDRe9/YBBGjyIAkYQ2WueXz1PFnOUQ3Nv8D0yQ6nrgdh0dxVj
7RVGnENwYMa4U0wq0RSCzQy+gylXGo0nZmY31mXO1519HYTiuf5onH8GKZIA41Bk
xUtP/ZjfBOv5fhc2WgmAD9VmNmq5Q84lOdYRvZG1YSs1HyKdK/MJYB+GFIpI+Ah6
csI424usz1V5Vy0/t3I7UHUsXoxbUt3zM3+tcrNflQjAHeSOgxNw75kiAwmR9JQS
qoUzLgGccVfHXRzUL06jVQ885JSFPEPdAa4DP7l28ioUe/KfWlcnB3Mlzg95SZBt
RgVIcSMLeZJScxyhctV9guCRM8ei6yOlV+mjqOME2eI=
`protect END_PROTECTED
