`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/LIkDqKihxOppwUjbottuxiNUvOngffH4V04aeBx7zlmw458xHkLx7jBNd5XAPt7
VMXnKg8uRmUfZJSHptyunlGPNL58FcnGnr5XGu11rylfFjZSgYjggWM5a/sfoZ+O
9S0573XMTtM+1fLtEuRDZrPy9f7xPVhGkyjZOcgrf09A1nVVnC5PQaIzv0zd9BbH
SkQgXMhJaFuVmK/EfNooJpnkrx6qeNvBr7KTjlEgdiDlbfnLIcDV7sbkg6IoaN4f
Tm7UKvydfjVuf67mHDUuMBkHPAqDW/PLkDCiTYtm2ingws8IlVdReYkRQd7ZHMAY
NsPGctxCS18StXpwIPjg0s2AZjIEmrWirMgmvf1DrVBJltIX8PLeZ/DxZPyZo/ou
I4H5gY/PNUERHR1saVnwntb3gwXEG8sPrHKQl49LItCxCqq2zmwMp0oPfbtdmn8r
t3B5GhvLi0ZnDogvfNeJYCd6+ImMmVsAK5O6zISf6Kp7KrjLdD4RrbKu/lRJ81Fr
3ygfRwcf4LCa99K4gUOOZcQByTfxyx/1ohEjJZbrojWJ6iqHi9iW9eZWH7yDJLV6
jnfNdXpGm0ztONOeQGmkGMEwm4WaAh0rLWUlG5pRmHkcI1XYpEXaw7UUO8+QjcQI
avqf+TibF6t+2SKhWWrv3xBxPsgyLnn1Rm11EmojCnKPSwrjXWKVN3HaBzosb/vv
sb4GwIrAncN9AVxEsr32S0+Xy1sUEHGHBappQRpC94Qjf1DI1LGhcEliI5mjCJu4
rR4B+5LskITPPzNRQ/1sUB2jIKV9PHl+jT9NuDZIpUcNaW7a7K60NokF8HTlKHHP
s07W6Dru743kIBPLS+r3dU18ZFPWWEu92MmlylQ7D152Ba4pf+C4B46ra3KVBNmk
cskF0qX3FEACHBpEt6TH1I58+oQJToomvp6E3iVVTyZM+htUHlLt8DziOCAndCN8
lwTMpWyMKIMXQApM15ApoTGD3b1c8BYdd5gBek0RGbuCm24kRrOsEUg7gvIU9AMD
JorfA7yIxBj4xVyM3ZFJWT2HnBO9gQiB2LxoApV0ewtHkYCj+L1tro1JnoB3SPR9
sXzhH4x7cxhg3ddyVykRzd13HSYJ9lKAxdpbKLka7my/WKoYmYZBAe1upPTVP8ek
vU/ttUMg7MYFYJaIhpXv4cqe/dend3uE+oQr7F/aaXaRMeARK1nO90dDIAf4BxrK
Za5kTH55w2iBlAAHvXxOYk46hME3c504wvRbGBxFlm7Qh0BpE3Bma2943dCKPin7
Z2mmFS8UjxKqBPoJa897522GbDTGVcgxr6b1iHOpilAWTbkvDoa3U0bpmWxJb6rR
rMkcUYvgCG8PH3T4cVadrh05G22jv/TTIbFDzjn9b4BpdP0T8/BsU2FDOGjCvZq6
LHXCi8bogs4nUHtBKFYPX6+slzEHxGsB5IIOAJ5yuB6PaamNlYY/JqWeyiFE60qf
3Rflp7d+rI/I0gNnWzVGo8SKtLuhSWYi7lTJCzRFiWvzGmu9aDb6qhAC9v+OlfuB
kC7MPHiq8hatPsxZWgG/bWnLLF/6BWu3n5n+9iVoElcmL5iw+8sYKL+UB1IGFYlv
rRVWkbErbIsicoX+Tb7qgDgOwwKEB5FobUdCYApNyZBY8/WDlonruk7Olv2c40aI
nSaO6NGt1XVWn1TWgRP4RScWzF7oCAA9LracHjOlmG5r07I/20tGl2BEC5P85eVi
TEvKbvib+qY5X9basUVNGL038iL73JQSIbZfORVRcLVHn01fLyjVYMFWtrden/CC
EVfJe4+AkqKdwC6Jc5Um98gWhjvX9B6ft6BNCYHaDIefUmPVZpGLJQFSvgzzYyCH
A9t96vT7gUREq1zaoFcdph0QAPlAVv5x0ZymDDTJ0WYL272WtHcA9DoVaD+lLiln
o0dQ3J+A/Tvda7cv+zX0xtpN/zOopv9/W4JNSRDjhnzjv781DNr39Apm5C4SNKDr
Ox+Q+p0+VoGSNyG+ZhT8A5/eZjAkBmuoUZgElPUMrB4ETHVCEzudeBjF6MoEPAon
MPyvWliwYcfirxNMNpyoCG3bjBLZawo8fYDf/2RYNCbNe6cCW5Oqmizgj71gJ+wi
2tNb4Ko0LcJvk544BQ0EV73ueQ/07s4E/0EEieF/spE5lecdH3Xy5Xl2GydsXUUU
o12L8T3XNekE6uN9wPAUqoyyrrvniL6xOQdU7bJZwNoYJSpHQWfEzERAClRtupre
cUQLeXE0rW2hbVJbq9+zURcJuyuTmgZBcclJBc1O/6yozN8yCuWAGSaDpekNQ/St
Ihn6165BxL9ye2mEeBbf3+BcUCMo40CI5l+24bqjyUXNJF2io8fYt/bp7DruaDab
cM1zpXNrkaUzobdJr5VyTXO9EzpcJcVnWXyqeIN9bv294BKeAYo9jc+tuYAc6bWA
a6PGE4VgohIlKAUaVr5Dp6A0HuEG0LYHNS1T2+hifsE5/Fz1AoRSvFvD0FNZYHdm
Ak948euRu3Bm29WDOEDuZLu9wgxcgr/V4qS1Eq1Td0kWl5P8oweR7lRpyQvmW7xB
YI71btueRixHuUx7g8k23i7uT0SXktHbLvEd576cPtdEeWCmXXmkV1HioW5+QSX4
ZBfI2L/LKf0aqdh9On5yIN9UarPKDRjpaj/WN/pPmQEHumzsk8vN6PNJyMRZGTOc
M5NOz5pTY2FEwlNwPuwGwqs+enqYt1NuBwhgGYXqfczWiKjYv15/SswdEwZ73/1J
adqjBBO2I9QI0D/xPGN5zqs9hdWqBmS4qqIdl69CF4n5d6XrCpmjK3veK/QOyaPW
ZQIsXQKXIZiPhC587bGKXPbgjfLMbzhucJsgZr72L2QgOgE0sSJF4PGdjRegNn6O
jhAARFbDlyHwELHCCta3zA==
`protect END_PROTECTED
