`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CZVXJnGCDgyP6TMCdZZajwzsGVLvXYk3rpcGfHx0/2dRvttCc/XuuUG3vKv8F/rF
13HC6mJFcu41K9Ihv8SuQzltOUexv44cm2V25TwcaTQRMuw3n89Cx5O7ZVixGn80
X0jE8DkqRHtj1esgJlpuoRUntsQ3v9OvUfADNxFjlHPVVCxRgGZh2GazLgeYL9eL
6Vfv3O1+iZ6/B74pLWPNUuV7+1vf6+a6FmYkltyUzIF4uvDFTg9X/THIPwov5CI/
DosEn332CqvpVBSzH4BJ72VhHbG5QLIhDzuxdWx1D7ITL6+m3t6+N8WFQqt2bl/o
p2REdWeKthkuI4v3QcgMYKzeWFkS5GHFZSK8/QUhuoVezJyXvoxH+08RSSroe2xe
Pxom3WMSQTNQGuEan13lGOc+aoERBvBmhppYRez/afUP4vljyfIGgD+P+acglcs+
1iCNlGfJDPITiL/7GX4VKoQ5XiSq0GTJ6ezZ+5sCXEHTl+CBKmN3y2v9Zy3gScED
OdgdQ0lMgpORng+hFl7AfpUhQFlFHRQp6zsHLh6iRehgbYF6cdczCCiZx+DBzjrT
AtAuuuAMD1OexP9UlXMsR3OsQzLKVs3LWVLzopwIQfVxI0NJaM2lhqicI44ROTOd
kwEyYV8UN9WZP2I7Epqxz9PYdhqi780tzkfU+76EItLc5LuelCTNBKTLMnNRp8+0
C1nMNnCYuC/cO2clpehvFvdQnlba1uoK1CVMYblJBIfOe18iVJ+HgN4i8pwc6uiR
xE4vGOxyfON0VFtzVv+HaB9LelmkjTCHowsPbwEm6WYj9ks5Vcpn9d/StDwxT6qM
dKKn7OynRG2/uw/iwRZVdvWR3BO8J1/EgMNKtBLZWZ1nykqjvEpOig7SBuBENNAE
NhkVi+fJw2T5WCK4ut9dvZEAVLypdWA1EGCm9xCvRT2l+r57Y8mhJ5fA+c1YnoHh
2xJhRv14pjWCEuuzqHEwI2DOrHIwepohqSc9TtcROHHEJqc3ViJvqhDB/z19MWCg
81gj/Y/tEqNMIbkjSlrnaoBK58kj/1bu2PJNQJiVScBRjAigucdbblz3O7eClvqR
HFTdls9soovIuqNmdhxl5WRujmq29RtgHosMDe2W7f4PRM4U/3ZxDz/5+/SV+wYl
6n83XpXm+TTEuyK8po+H3/qptb31G1Z9QDdcmF+zJE5Gxb3pdg5gBr63IJdicVFf
cg4J7zQ1e521dSYbbC5WvM+/sawJfOX9D1sB0ZGYCaYI7fZ/caAMg1dtC56za8rS
fnKxGFlJYzW7iLY6PgmhvC31l5yjb6+xtvO14Hv8XrhAaX5ZNsgupN6gL3Wt5m+P
Q23WToXP59gj0bS546Cztntf7Cm164vG4UMlyYxwr5s=
`protect END_PROTECTED
