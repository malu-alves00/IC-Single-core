`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Xh9RMGydmzP5HXyyRYpenHM/vEpCw4YbHhHnlCzYiKsiMFbPqTmPjixcw+3D352U
9rszB19zCNmpKFMrHi31J5IrsgVGjlQQH+CgMqS4IRCnhCihusy1ngu9ZHQV1QHT
xKrfVDzqJRjUNL17LWmP8Y5U0iZqohFtC7tNWbbhu1CYTkYXEAofvINDQmHT702F
yI1uf81tW1TQ1P+ytJXHXCgLXuK2DvEvv1tShHixPFLzpXfPwn6zZB0v7rCxEnF5
4GmmOfKEEkB61dp+OHL9xolgBpSaXVyf0XKpUnUbRBldzsA2nVwMZk3oSz3Ttk8F
kO3fwM4WiXJpzHkSJY6jHxw6HRH0JB/ABq6WJ4sPeOiYOsivtvYyuok+1Toa/fqJ
KMFGBaV1TEgdYt3TOmkgE4sVVwWGMKmpz6IJyp5gqzoQyph591JUp7Xo0pJdPlx6
vlUhX1JpHAx5E0BKThW2PJirQxgHQvwXdibIS3vcPdKpDtnsYorb+hSRLZYT0+TK
GT9tZxDjBoLx4Pdnb9FN/IuZbjAXUo3ahWdO6wnPhPwCRWJ7DXji3euh0KEq2DX1
tkIVd2M4nDPqY93zPBknwVqs6H+hiyGRPcYHtc+9rkvelS4seCgcsVihQVEJLLTt
+zmrNI3nzCUakI2TaTMREYhMjnT+L8dzVCkG22sUwdP8gDzqUaIAK+rtNerez2E+
L57/x7PTr8+zBxv0925k2PEJj4n2MHNR2GoQbQgSHfr1DlNHhXuyIJtrrISACh0K
8TCxbi05PUU1/TSX13CnaIxHUsR4RyED0K/qAjVbVN1lgblX9aGDasRWUmYx6JmD
Y9tGVgW3u1V3vXUe19rr71qUBa8Fv8OKTBJKwH7C7JIR3Qqh8hyASOJBmtX0Q+3g
J7++/AgI6lkjgJPKqxVRVDzA+DxE61tW/y6B6BQM/g0wxMhyvK8NauAL6F0ifC79
qCi7NQRVPBmzQjsv+a1KcqdfUQ0anXmxiJdz+YOUQ7fVQNO1H5//Ruc88ZS8Y1vN
vKJeG8QGB9YYCdvYx0bVPHvHxQpVmDqx9daHPvVngK/GuZHqZ8Q+h4CqP3pX0jU7
af4eCf58oAcXhkPHjA1uNgLYcwm4qPZBOsPdoOn5abYkFwonjbVQHSGfshyCLCPX
tArWOxBQYXwGMjJRRofRSPCHThm3P4t0ndpyYiZ5R1D2oRxw+6LRLpVrUNajPxZw
V3UdASZcxFwUEBNFuTsujpFEd90hBKp1noCZ0GSftAOkQz1AEDEBdHGCHoiepGC4
SERi4n4TlZFwCe2Ph//b2qh531ebO+J9AiGS3P8pf2xp2rIaEs+IoFnXmcG1p7PA
5RYvZTy4sTFXP+pMX/Xiz5EnBsFNYpICRzGewRxiu3ssLHjgx3bfY45AyHSUB+rp
lkrDlF2ZVIHPbYv3ujnrQdW24XuUwiHbSgH7U+8OqbTQj46LTZgc+885wLjxEKK2
CnWjnc1ITcY+zXqqnBKH/ybDeupdhPCJq9k6Pesqw3o6IyGIkPFXHpFp3XZGZvsV
tTcriB0HEjzJ58ZRandBxfVdoY5jf0VWBciwXhYSAzHuI4VS4joGKB6lOtYJ3O7t
ESkBYCjFNvdepWL87y1buTBgANjkSY0JtLIgfHFU+/iXs8V5w+EmJUrVcTDP5UgU
F4UVHla/QFwFiZ49rHbTSKq6wU4Su9xAio0fGqJVo2MNoUBa/WTBeAXWvtz4xJyI
O9iYl79nZHAQhPa/AvXQf361aFlI1gJKM1KbtJrHw+Ai2P0o0M2c5cH3GC7Oh7tB
HwL2IDXd92qj7kXmIIA3SGl7nSC2O1JJIZR8oPdgHLLe+3uqsG0WsjY/JE4q3CRI
yaLr1YUzugtgkWro7Y0wJnfN0G8aoPBgaoZBZFjBBDgIWjbL//6qBfEJpRfnT0nC
nFzdaV7rDhGIC1iJCkvAhMC+ddf2aIqPur5wMu1FgxjET4GVZ59tlBApfCGLM3d2
3kQJiX8Y+EJg58QFbfTzA0Q9ZL72sikc7n6R2LSrJC0joTT4yyULBfjkYS5f/XnO
KfkHVvNXVcKII9SBt6mnc8TWkhOtwFSuPvnYGedccHNdCPUPIhE5Kx+ulROJXHbr
KTdITrMmqWqGyHTm9h2x+0o8+uRlgBsk5aegJqOY2+5dVFV7HRAKfT15gTEquVTI
xg72BAQD/HUhshie6Ud63eY8FhARWFHpI7pYO/FxacaX47T1F03E3+aGP3MD6vmX
T/hYDLL3SJ9fFJ6cVUxZ0x1fhEWqa5DX/C9ldhkZd9XRBwU16vgGaFB4tzlSXLiS
hvNMU9yFv4fdp8Ut847GqOnJ5sI77a4GVL73gI1iClhlpENnxe1DmPy+WkeCuBsL
aXVA1PtgSEMHCY0lRt5nIoupPItMO8EoQ9xvq6qYzZZ7X8UNeFWaDGyhcV48BjVO
rC/DsF3gHOja3XgUlaUPg+oKy7NHJyKlfVHNzCbT9Bqmj3O465zYrQ1QIqcrQiNt
IkTBHsSOGesXEE7WLIQOT2fQzVg11hi+x8ROpWa/QK5EezuBswABz83JmdxgzzGb
DqDO8eu6j/kVSwiGXlMpIzX0bGD6AN2hfpRlo2WWNd5aOypiinqQCG5CLBwjuMuX
Hz/IxlsSuVLFU93qrYKDrYJHLk7w+HxuSi3n62booeDTySQMjziq8VpGRDVvcSzm
HD9hSHdxwBdIQ6GJLHRhGcQ/MhWbl0D8EOK6teEJnuNxz4UA1SyNgccf8uUY6SGe
qr/1sK9lf2KzKp6G6/m53cP8j0YR5kt2KUS1MuH1Aqrt0GvlfiGYLFkJpxH/rqAH
wPYCXnDo6WilDWW8EabfMum4GkEKAyWMgGcsxX/9iPLgolmypatqbY6BMa3ve/CW
z0DUBtCajaumQIFn2Iht9EcIh6++bSIJjoebnrysiROEEUKq/NRI2zujc4zlZjOJ
9mGTSjJ2fz+s5+m6Fo2bPK1H3tDu1eRVp2DfK27zeetsoOXlpB+OLx17zkGk9NCC
njGupv4YED2YHdfuwDh+0PnKon7LKrQCYJJVAbNK71V6kVdmD4i1vr6p4++y6/lu
15mYBr92ewPLYV/46MfKzLZ4WctbTV8iXrQvNHcnD38dhCeVgup+OSG35tjvfV5I
CZAMUgACP6GHSBU2Ty7jjXp/2L9dwN4EaMNVfgCrmAn+U2nYnCULlqySxY3KJutY
gzq/A2os8JU5MUm5MCC/dWn6CV7NNbS3GBjWP1FoXDA5ehAcS1ISMgfr1xGZ2/j6
PO+EaIqJXEfEBd/B7TN05p9HY52meepQ7e2T/+RWteFsMynNs/BV4EM0TIIF4MXv
J0ZDHHOJS+zKZsmNj/JMxBE5CwO/H+w01Tein/dw/Jfz46rbkDBWfFqh0YGRRde1
Nypnm85La9KoNwNryZTXhN3wtqNSvguVljvIV3FPV5eFwOZFK9fRgy5LwPDxTOb+
2SsZWKp6o3fvwy34n/QhSbKohwz/OF/8jREfQdIhHzbZ4U5bvO/wO+CES/S/iFQB
1pMNhfL+zrbrbVoAJIpOKPDgA92POXmGzfBAoyxl0yeskVSW2wIvsTaUp5zuMuhG
+VFK3nL7jhN+tmUv3wN5CRUZnN6ux4SENCz2IzEQC6wXfGQves/bl+ocVf4UdWFA
/97+e0esJhYetoR5TKAANczGr/gU9aaKipfgMluuLAQLs8UaOU+Rxv/2wozCygIH
WLHZk1LFGC40EhVN17/xEd2jbMb919zeRgO5+gOnxkSXFOcnZ2Iyw2fCEUWKlaDc
QParPu46C4wznxajZObuMffFSeq0P+N+H8zHQJDr/gr0CsYwjT6K2nIH0geUEhr9
m14A2hVZE+mR3vEHudMh83w8w/iag7avbj9GUbkmPY861xnL7w/xHCu7ZB9A+W96
OsZZgW2+sUj/+69tOP2NjGnUmhXuchZqLAqGKOkSQdplBPWvaXQ0bkBIReZ8534E
u3nSw8EMJ29bF8HLJTec6A1Pxy89LDWSeMRt8JyaX6HgFVIWcvfK5OUW1fuwd0/s
zmQqjaD8oPsvypB8ufJCY3x7Hf+Tdq1eAXCMIhZ4l8bn1vgeotQqVrRiMA/eh/Ba
huI/rEgCV170iFr+zVq6Bvo4VfIwYlIpDsr68Ee0B3IjLClsKtMARkjqKvuGbeec
40RbYU4K4yXyrGF/KBODEMF7TmZydhJNlRvssNqPHapc8QbfW07YMIf+TBR2FrUl
DMHSHx+8K6iG+bavgnkzTmVO91OeVdXNhyIk25Sc4ngR7AcEHIht2WTfa9RXAi3K
1vR9UA4vdlllhviM92OagE+w6d2AdXgo/RDCUMXqekYQEh+gbcw1VCevGEDLk6PC
dL5Pis+xjC8b7nWfTz69OcpddYwO9/r1xU0mLLjA4NgZpjuyvl7jmeKu6BzGG7s9
jzlltGaImX2Ih15O8JVAk4FY2+oLq28BfYVVpzsXSWs/p2x4Xc9xeyeTyGIO2l5P
gPMOLqsJX15kU2/4/yEBTg7HQ+8o0DhDxCi+plD63pmO4BOfYpOlIlyFE7SqLFRy
KaxFxqGuZK7agyD7MNzrgbTNA0ScRuEc+hnuAfIywpYfJ/LroPeItXVGuAi33zmx
jIMItQg6Tp+5v2AkyeXXfLU04oKMnYoXwLmHgfKvimRow/wirlhsxqn9HydVDGmu
bqnekTWtJHBT0XoS5lNqALBG565Hl02uUpmongSYIZNlM15SjGNLbQHn9Ry6tVnR
Y0PP6hwaTD61Db+nKQWfzWznunmcnmUJ+BITAqyQnLc3IaJpfldGm98R2LoGwrkU
uBtK3TWMVTxXW1HAEAcWfGKKwqZOp5xX3myAv2tDM8jxCG+XsO+S2l99jt/H+8VD
e80hfOwW/xbVWoE39qev+TAYcTJ0ataZfKp8aA+yKayXLchPrs6WFhtD21tqASyh
5OuX7JAl4bxAM6Y6+O1sZpT5GlkoCtT4hmpuC5nwWmVwWWWL3rx4ePufbiAUwGfh
dJefacuAZYgV4okQ9xHfZOy7GWiGQoAJq2UtpbTsHS24cPMgYchGJqSBz+9ynMen
zYyYDE/+2MMfGNTqMjHAflVYAlXYrnvMAsPx7tPb8Lm6rciz46HR1G6FLwHfXE1R
5kD/wYHNJpa3hVFDlGOXHLrnKgTaYhBMO7d/sdQVcpX9gneWAg5H01MNgcG/NkiM
b0IrGzmU8J6ER1X3CM6fHXuJFPtc4+Z8qTO3qb2qUa6/o7nsAEPT2EFPDXRwQ7oh
DRFKYHVzuMNyLPUJrL1YWy0yqb7sR6FCRAdiXgGQmrpiv09la1sYzkza25jfbmdB
d4iSvpiSOpuifa1KRFBbMVrCrptqmu1U/v9Dwi/MhKpHt1h1vCqrQxR2/QQDpzFP
j+taXJcTrY1hz/VtrVyiiAF5pGzQuxgEuIZ3ArP5A+2o1gmyY20WTiFxn4JsvGZ3
OaqYXnj29YZlbo1AW1vljU4GF+mLXLyKMF1hcoPa7kYwI1tFaSgrt+Hbq1NBDWJN
M5Ng5HVfu47iXCbiGzV0lJcCAhZy4v5sff5pxuHsjdG6cVDmtDhCwvBH0cQsnTtP
FAfOE2pCbq++ALVSyz8T8yeLvfVSRjq98vKrto574bfIteha3pIVKkl8cyB7WINc
SzU8WkUBRUl/9WV2+SC0fhpxr1cb1Gq/KYgRZQhN8XCQCK6tk9E9QuIzQSQFp8HQ
bzAqrMK+HveRnoHwLtYMuHndnWrX6ByY2eWasJu7CuWUfb6lhLC/FMExu16IjFog
vjs6GavGRT1yztPWbe52sinne7P+oyMnbVMWvTcQnQvnyRMkVHdFlYfVv5N//Aen
miWAzuD/0VLV1kMZrO1azzNeIhiJqy/G+P7zFaat6BqLpHIOA3PoTpbtkYtYzqaZ
yJgSyNNETH5oij74iERmcOiJONWZnsgQBxjTC+C8LxFD3BxbiYkIU8KJqrYzkCLk
yUVfeSy75u6TaX6Q10w6URn62jNGsoWc8dxmZ++EmXYm2/ZNhaJ9hm8MlJ6pN3se
u3IZB2lZP1dnNPjqw7+zdJTvBdFo3GYM/eMBbEwtPhTMeAPpHywn8/qh6cB91NKb
UHODB4QEsl33QWAJ8JtLIyNxrg2KDidb2t6FnCzMEfoapEFh9Hoc0iHNfWsBdYzL
llNXME+c3JfIZkHi1pWrJTbd2Pp1/MGmwLCEsLNUgNe5NCGSmvLsoLJGwSXDW2YJ
hUQd9qYNeL803IA/Al8I8/qLQeiHMimECZVDLag5oihCr5dsqbLW8qg1anr7WY8p
WmB30cBBWV5FAwwRcsvgciY+ZpUvRZdYon/hr3WDqkMN/n9UjKSZzKZPevjNh8wy
4hFBu5M60tHw9CsMfC6XX8RVAnz/0NafeBka4fVabSAEj+bvAS4yiEThfceuYhl5
vAVQuT+BSQFZFR8lKqEzdJuvet0TWa54lyCMQFWI5sHQ0F8RRqCCWjAwnK9iv4YN
uyd1275PxB6jpYMLG8J06qSAwZzFMnEG03LagPbnjp4ltdSyD/t7RQ7IP0k2tA/6
nN1PzXJettf83UbwnvcB0Hod+VVsR+36/oyrzrWtNnncoDZn2ZWrURs96v7DrQ+3
11t4OiFrLMQfi1FhWbI4Df2MNr/a0eBeqOc9LANgdHkQfrsdvJVuY1nikpWowvtu
IrokLsn3liJvbO/Zl//8/d5wtmxZ79fDtwtSvzaaZcXRbQYoAIc4rOCswuz1niaX
jSln/YkI+R0AOYDKeMdg0lu6o1Gh9Lx8c6F4u9edQY4Y/uS+48RLSkso+UGYuHs6
y8x9PMPZzY9F5Tl9GC++LuPsX4dDjPajnyCym5yhqVNf8gYzrclUy6lnlXjYAzDU
NLbMLAwcxnVOk4jXhtaSjR1Qsak2ySt9pUvxSYSr+eOamVI202oPlRjRnFolpqaR
FcR1rwwlEjlHFJV2QLG4EIqiA7emFeyoVP1Ad0wC3n5f0Rjp4RNR0zQ9L10L2PvS
JR0hZ2rXj88cuvI6HA2bb2pv02EuZpFyGyJSbsY8heiep5cKnfIvbkAeTyq03TIg
4CjOm2T1w/qTJKfraQOT/kINecxET3z1ROHzDsvsN9dy374R9PXRfuk+18OCfA1H
eATXZJEPK5Hww0jPryFdIXdeMP6ZWNuIWEniNp9HkJQENXRtlBdXqunEzAxLNgvh
N1MTZSDrJWn23ICdmm9soJlA3uAk6UPkULBX31S2PZ/a/8qnfQz8YqZO/2LQFQsm
ipA9SV/sx7xggUvrM/WlMSmSS8Htr01z+ES8MpPV8xUTF86C016qceS5PW6Dow0z
T02IBr2Zlf6vkG0S0XhJu4BosiKs5kLqqZcx69X3ijnr/+CicSx22pZan+T2eu1N
Fye3y6c2BVnYUyYOAXT6z6pVjg2bXtDmrBrUqQk9ro5iOTUqUmhXAVT39FZFjKNt
DPr4qOgmUrEVGZXApX7MCb41OXiR0aBgdyjDRTRV9s3Zjpwhiwv/MNXFvv5Xt9SD
Yu0CJdMGibi+ObOm1PPbL8fgbuuBQAG7sWfRhyXpK2uPQcrAIRVU38Dg7S3yYKtH
jmbsO8Fg8KX+k1zgb2Cd3mB6UPAa2Sp0KaiX/YbuilpY/gOrdGaZPfYtcaD3cWnK
yn5JjKE9JBm0pdicINPPK7lrJ+kVDttIm1QW2hP8QdxACIDqmiXSeBm0zpd1BoKL
tX7qBpaYvstWWPLYYuKb5wRRd5HKUbWjPqByGl3BcMcdxR6IGxf0Y4/zZekQcWUY
Xy+6mXXkLFECYOvzQ64Ww4zNvXzYBF3FfcWvs2gz5FBzN/XonNcZZpZ6jPPtCoTU
tN9dH5GaQZ39EOY30NtgeYctK2UckgVuStxE6p2krbsDjdSPtdRL8s552aE9Va0e
rh2XBYV1nhQkw+3Ku15nSoRkGwpch4EAtT13hmPUMRCcQi6xnjP+tk6CaFLf6ZHO
2/4pADIla2mQdp3gUx02Ty4HPuPJzcDa/ESLgsdGgb+TIqLn2hR4i3UI09JtI//q
/3r+2f2oSkrOVgxDbL6kkaUY4APIVY6Cg4pValgTVbvyfnK8TeYvMbqENXSMpMOs
rvdSL3r8DdgZJVj8kjekX8vZcBEFzyW3AQwMdk0rDGTRONKvu1mRdO/QkON9dCWq
6ivMOjFNDSKPxZhW2FJtZ2BM/Yea555AauPUId6USCErQPrDQjGUP2lasRXkcA5P
VhRHARJhOwauFkv/DRlyiQ1Mj2mA+X6WYJSqIWV9Bwz2t2+br+VqlIxTgJL24Z0D
MECfeACgGFTfPzVLwrbnyIEIHbH3zUDjVPsVU3bUXpmrxb3g3E0G8Z9iI3kLStlD
+eYLOoglPvQxvZgPa+8oDWEvmdsWoP1uhydqTDcjVQCEan9Q4Dl2u6P7Y06VizjX
DP4G/r+FkH2cjXO4aELdSwx3QodLOj9uHHP/9D/Wrz8vzm95JmGaYdNXbyRIUBvt
I34J3Mw/EJfHEH/oAribgl7ASCX7K8wBAU7w+xaee0H5WcfpSvV803I195FPOJuO
sc2+SCQvVY+L0q0iBGCwUBIEoQ5/FZX3oWmCRjQPjv61kt94fugcW+tpKmPErBdK
MLN2hsxZbSLXSzxhqhfQtT94EI8ofcmc+xPawytvaNi1dCvjppLylEg2YdAAV1z0
1IXOGR+IUQ0WMFgY44su3NeL/jwAJEoMaesjY5eaknZo49JXCxvmqgsCfoV8URSP
jBJzSWrB7Q0m2OxQv3bULZrtOtANC3BrdOX4e1fIGgZ1xKJQivIqJakoat5NEdNV
9UAVnVpJxq7d/RK3nPleNGeMmEcefdMLR0vEZCA51HxEfy9G3exF4+MyV4ClW87h
iqCUUIIJh2fvUB7FXw/r1sVO+iFy/osROkb6/1HUrFUl1w3ao4+WpFQY7FBxU3/I
h2VIFFN9uUEpvUvziNjY59oKG/SJAmYZe/ikQE4iA/AWkcjpf6m8E0cUYJoMB6AG
LMA018dsYghutGeq6P1ZxcSOeddSRU4NRwxyba0bXHtJQc7TvYHIo0zF2gmdCWvC
4h9HObSXRhnE3grV/2XI2bjNQY+aaRV/7N4cxDv5/aygsUdzsyymaTxtdgOjg+/5
BJIqHT7qPXgLVe3egxgEblcq56k4tK5bCtEKgy3QTghHBguswlHL4q94ZcvkdusU
btg1Z4CY/YseiZ0s7WvASkfFpMyfzszCIsvhOrfy1qac6XTSZYIlHt6RnVaFhyj8
lFbyF/ERBdWMuawnIiFhtYCJR61xrn8uogmsoWe7uop0dXuKWAu6rhzNdpCpv0UO
7qWgdu4BuT53kfIo8P+qWYKVtVPISBNQFLQfBtIu19x0Dg5klSlH4cdxyWpDBhBf
dlOginK0pIUIWlaFZDLZblCmaIpfdDify8E5dJOdQ0Y2dQ18DpRe7yvorOvuh3OM
GkLTdUxm0iOhb3Hc7EHYELHrufyDJHc/fgOdnWZkl3Gc3F6T4u7ur0Z8Oelasvam
WRfJ01H7nnbPzGuGELw7ba+oU+27A2v+1EEWqgI/Mp2Qi2mGv/ka22Ew7QYeeOQv
sV3636vbZcIavYEyrWskyFFvwVpusUIvVORapmNSSurF/iDBpZ7u6JimHFahGRug
ICmqePQNBxxzOFGMo8YGGdqg1zkpo0ZDqlAMo2UhO0TFwQp09B9Rq/gg8nr8DYvb
FUSPtAPYcunqk085BuyzThZYcDnxOMatXEIBRa3QIY8INGUbQkshGdZjCkSCmtmP
0F+ZP2v6AKGiV2lbxTR1mImBfhQ0wer14tusfQEYuRDpwSZZ7iP9HYjMR2klTPMB
GCRoOgLItbXJMPIdAPBvP0P3I/Hz3g6R7JdlnuQR2Wo0SQgA7LTUEtqotnGE1zrh
lWxqHVE6UQLN7r2wXzAcnKABr9DCx4CKCmaPwkViyKoYgduXprFpHznVpU7yEB5T
M4a2PBWt9xs/ZbXHBXo0DTRn+udW7R5zU4DOBqbVF0PhY9G2IFVtyrc+Q7RE2oi4
SlHWeGuAJ4OTvsRwMPSxsVgFt5Y5e7V/wkSo4vWX5HrPzpQuNYBHqYF+bgNAQsyF
qmtORSUhnrp0NKdWoAvJM/h4+JRIdcT96g5Jv6B1/EzcScrdV537rqNsyg/X2X4o
rTykspBOqKqj/cYRud1+JX+j38yFVuo8w5t/ZVSpG5csDY0MQxasADum5umQxMYZ
qZ/D24Yoa/jDJIvFtB6sTIShkmTINrf/5wGIkV5SdVccAIb9V+IQoVdPuB/PHbH3
rFxB7s1A8kyWiSXxNVhrUNZBKzNh/l7WF6F/XhGHo8YNcb9OvC6KFq9OR+Aus/Si
HYPBK1qrnWFhE5p/aIqmDskc0yNbWiHrgy9iA0xKtazSC/hssg+RGa/ARtzRve9j
OS7Dm9Z+khbjrUWOOcKkDL4hZ0acrkHXBWXGmcBNDKA5vR5Bi9VB0+NAd28x6ope
1+JKTKXEMOXXJaufzkzCLiFHUUjZr2z1iki1Vj1lJwRipU5UyoXFr9m8ut9Edo/p
DdDs8TZM6kv2qTOUE7sibapohNMmjQcUOYn64MEwlPYQiimguBhOnAou7KyHFoMo
Qy1XYxdBGBcL9aJm3ZiYAZMFM8CaCK0e9s/2xKm8FeP7T+Pacv0e8p0XfvwFLluf
Yco1U2xRnUNRX2NH3HYkMcXIR4nk/dj0cQ6Z9pYp7a8816zHT6vYlSZQwFWbZgNO
nN0Vp4gcj+kKSmVpn2KAsctRlaWHGnSJ8X6S2Bw876mgAekhfDyBLmFr6Tt0rvbu
gJNGn944N0PnmEgUMwK17e1mdfJq8/Nk01hx8f3xGFi6jnQfX2QxduH8L6vFS/sS
prheyRjFe9Ha+96/xBGm3NqI0E0TOa85io2Q+Lh0c7QrhbmQHXgUODPAZ/lU6+HB
93TU7Zl6u6c0dbsnJ/+gL5rMHyrDxmP3OrMcs3oygXnLgCzvM6a3b0k3DU1f6Clj
XuXMCAFeeKjBFZoeWfjBsKaHDic0dpFJMFaP2HplEWJBoTqBe7pW6KweFkQ9Juie
Ymoy7BKrH030dAsJwR0iiKfjKmXkm3SN0/wqiFxoCxxTAg7UJerZ5VWJSl+vl3sY
wlzxYZZR0kp7jUTgBHpVyNOtu6k9P7JYlz0FouLcNlfI5EvOnnhmeW2dJB7L9Oi7
+LEsT4dseRWU5O+BEfJ9PUyq+YkWxfJlfN5GXXoMx4gDqwLAKEZa2orcdKu8lBM6
W8SVLTlEBgUYvqJoAVzWrancU5DpVDEoBhoMs0FQjn8zAx+jtQJYOfiQUgDBog6L
XviSO+aGfSV9mg2O69jMpNpuSw6K3AErteBGJmixp7H21Xm2++dscGrGZIiUWy86
7jQXc2b9PPRGYF4r/HAJ2A6S0KM4tkM6sW2DQyQaNwLqZl3kU1h1Q3ao+eHcA5Kn
GH5R31e1VReybFHoQJ6wEO/LVbwualX7C6w6kFKQtEBx2Dfj1B0OEwu6l9mpMLRU
L32zafXJRV9MEOf37W5e4SYv4tllYX2D1VT/94jWaNw1RkfaIiE6aEfScbkNLsZ0
6cDbGe/pe+U/nP3Z6IQ+G6Bb8bR/FR9Xx5aCmdW3miZ0M/GvqmCJ6V81HTnMhRuL
Wen0hr4gM/QbFAkbJS8JMjrSdJ4zHK5OmfskM/ktk8ugqsMbU391f5ztzCtgDv4U
CyyqvYAXB+QQjBNbXI714TrH30FY32DAQAXxYaH7vUeyuhRAIW3V7y1PByINgzyP
ivKkV6ImqiBA4Q3y2gELhP2WYgzgN+ovP6xMn+YdzkKqia35ErSOxL3VGhTWLzHS
sdu2aORaJ4olQapdrGCzreunbr+LlbsxOLFy8/0toCg5/EwxsEx1geX++r85W4lq
GKbYlPHA2qCrgVnJ3F5RYdObTTevmXeSvbQkHAkEMLRB6Kaf5EVajqdmdXD0jPKf
oQwW1CjXGzI97ncrf3mBDiDbkNLJhmecOkxC6b58ypmdEH72b0ihRBKuGl46sJOt
F5heQb0UkRg8pVg+WfsuO0nRNuSh8qK55UG6szeqOtjvGLil3htfXMj3wg+K8gJR
F/6oBnVy+t1WP5vbVM1GgzlxWx8vaFwcWfnMm0qyZOSTPHkv6nEymm7mCIx19iwV
EWymoSEL2fwT7Pk5YstGdB22MA5hmbRwseDLQIr2UeZNtE96GeA0D7NAl4E9S/E3
2MRs0Bm8yB+DHqxVv7x7lF0HkcZXzu62nbZN5Le2qS/EzjEXdy65SZvf4IUHEwWE
8luERxzSUaXEuvJub3ZjPYt8mvmGgRaAmGgXH4SQlf+IeLaGv1gb6CP6rLiO8uGy
rBLnjG3ZWcath9uK+jwDUVfveRxucgWtcG/739yxD868efL+mQlTqeb2XF86o1FH
cJ5A8j14TYvvGo+RZxnfrjeiac8BbRacp5xBitdtx6NGvqdNn/RRl+EM7KWbt9KM
W37ueylF1jeFucKUNyGmnFwm32LrURrM5dLFR6CvrZOkgtlLLu/Aenk6po2gn+hv
JoP9ig9Bwvissz0nbkD66w5JzZrUIeXOt8oWhQiFS0IHK9o1Pkf2IEawLG8sXINz
iDW5ARlB7YrkMcMGZMLKNtYMSYiUHWjApYNjsUcgV4CYTBrniksinDR8MaVjrM8o
Lb355/09zI2i9Ve7ENSp+xWWPvLetGLtiXzDwBRq5zgk/oNjU0LUQbKDuHiSVsTR
7jNh58B7yAkSlGt9fTfqqWFSR4hznlXARen8X0RoIKyI7YDIZXsz136WyODMRIoJ
beyrxW0RBCFEzhiowl9dJosFvS2dkcIN7tUDnGPeDLgx2MZfRQLZraIdcqrO8N9l
+i+J5Vfm/stzA+KyALKU1YN9lsGwyWOKvQ+usszGMXQCfsyfRDIyWwbi1b1UsxUS
+lluJ6SO3oSllyq7GkXa66Wo8x9BEWGM/e4E2AV1Iu0LavFgwPzJGEXkdmX9enFX
T731pWpeKiCFTnWPGdepvRIbkSyEvDTn1RJyh5qGZknNRomJo5j8At/EBr28PT4P
lbJuSZjDcMb9EX1KWghTBMjsRwPko3eU/g6S/oD0o3IqmdrEAlej3bxfmUCVzAzb
4Imbp/5305ECjFQcWhGDmNjG1k6YzU3bUPNLWJpI1JUPxr7cEbD8T6yHuzCz0CxH
lxwWz+aHSg1EK/nBnvsw3AgKjBiA/FTyg54TmsIqQALeQEyQQhLZUGgJQWd5DHTK
9fGxBFeTkvL4wWX+4tUguW8EpArfSQ9UK9KRMtZKTk7wfh0Y90eK9HH8GQI0kKl2
IPJGQ15ge5MCkh+Na93m6q9VCUUiboquGHfDZUWUdep5nAg/e2q21uvQyygUrJCR
9SxKBf2yWfr324CgeL/q2HNZpd0QLV4Ozu0teV2F10hjVZSU4jtfMIitBoAUm8+0
8LcrXxHf7jome1r/N5vCnYnPDF2s6oD0+GVm0ZB6uI70Ry8ZHbSvevysKqDRYLIo
dAMLAsdXs+QNxKOWWkTqgR1h5S9dHRxrOjY+tXXWlvlSMhRP8pNZ82tJurGAdgQy
GH0UDezCU9aNu2nxciXlYDp1P/c73/5X6zCFBKOXZadrQ5eB7fcwliQYWMYOxfg/
CowiOG8O1ly6pP+uKrqC+cPbbCWFW+7mQbF+W3n3mWd83/BLqqGxXDXsJhI/wecG
sOFPj7PBNxYvjWFY/DYIewLnpfJW+08QXVDWd3hLLR4/3vMRCK+MwrxoyCNqy3OZ
HhNBb9Zqbr01f6izC2BKi5igbmtRCcTORbxKA4zwhrtqSzJsippb8DvKaPhYBxiR
yIWNwo8wXaBRptCVGjJm1W8pgQc4DpBdO5HtV9TVJyJJQUmtUQWt5WehcVQjGRNj
otUAlcJywuOdh0IC0VoTYXhOHscFj45jUYiOMHJlecWrwI4ATl/AMBuV7a3sCnMv
VtrkoSCRt229RXgCccVNW1EgJ4SBGQtWnzZIzcvLllU8cG+lszffve6nEhDCt7s5
pKkdxCdd1xy38wpUuEKPNzcbqhaEkAvTFQukpvmdahP3TMdIN+RtqlOBhHcAvaK4
MZc58oXUFg/X8nChFYEqPlyAp4lZdXvF8TW9WuXqpbtJkksoD50Jf1DkPeYFqzcR
WVh+P+/MpVc8gGqRT0XwTsxKI1iNQH51F7gt37d/8p2xcGvIY9AKxbIBnjIQDFa7
YRBqYu2kMgdAQe8JJb7jV006m3PgivApSA2/2mXsghFbAwko/zg914+It24ozjvb
gwk9qLrFs6GclJWCy99rYAVRmy6CvMczxAD4cx/+AyCA1qEsSAC6CXKKgbM3iDud
fG/LGdVpGf5wn881aY0fQ6Ua4uGkMwD8kpZXU4u83d44k0+dJETbnweL1S8gByjl
Z7jd1QoAQjv8lIDJlP+soksNoozpTDby0rm/xxQZ63uwrlwSJUOXdLAnbAntTJbq
nUTsr7dA3+Mz8VDrprj61ORObUDd2a2yfh5Ex1JSrlFpO+iY+Y4/hN4HQIfucOU5
s9pz1SxjpvY0JrsdXSUxPNA7a2GAS52XBcHDbineCkooxVCX8IjIupc+6ZnYIcl9
o0fymwvcQzSgcwNR4h5gzcJubu2fazDvGWdR6xffJZdzOLJsJ1+IcFjjvjHbrrB3
GgK4AyVR5g57eBqPiR1wg8MNVpNZxYdq4adbJ+5PU2mZkJiQpdgg7/HmxpG5fB7C
ww5UE7ik7PAyqa3Kl14Y/fTjmAgt9AgEymE4u2VT+dTn9RdBXfmgUxFSfJgwhmg8
FDDMh2XkKmrgnRq1AGccsAeE9yAobU7q37TUGPl8qUkQpu6a5IaQgl0OunjW1XEt
ny0PMgk3L8FzGrVAFXSlnMzvsQ/lEvPfw917AI2gqR/DhAzFkqYtfyJw1BhzFZx+
49xgYcxrZZxa44N8TUuRQrgtsNkjEOKpInpaWCaOLJy1YcL1VldniweuJBjr0+Rn
ZCeIayBWkJJLmq5ehhvCHOw3sX8C8yNioSSJkKVRbJXdiVAoIfmNrYvqnw4hUMZS
xH/sBcG+3YOrIJsPOi6FK9r2ujyut0zafHNMtORPcXrLywDMTDAMnHB+/4OefR2+
Zg9X9Ho5ijtP08pxFZS+OMacAET7xyfN6CV0ITv+pkjTyPd5dv+I0U0cJIB/xVde
CLntxbKhtFnA8F5r5oGe3JKWlJ2VoVUr7+SiUc89NmPe4+S5djEfjOtRv9wKIYJC
zLVnIgMRh1x4ebdHTB8C8j44pPts3hTmvYdZefAc/scZoHM8fAdYUVaAnafrACOD
se9wzREtLr9osObfUEoTRl1KG7KtgOR5XRRi+rj8er/dj5BQ65A/skvGmJdY4Zmm
zKLkgYdA239pUiC+F/ztcXDyZ1uS8h7dYMaXmRu1OTkffdV+6U9HU6NiaWwE3ZZt
xXsr1UpJApjD+3UM/lGrpOF3mNjb9oIEbrp+hWBed7jiqu0I7kon4ng2QfoxcwF3
Dcog7W52NmASF+72gbSoq0Hi9wwVN7CXZ3/hEXCz0fXnH202u5cV/PMbdYzrNYZY
rJM2Kd3wdJrZJTBmL4wWDF3wgp/e4/+f7S/WncktPhsv1eBhqF1XKTMLP8nWZede
fwp9BBgqcTH1tCn2CJeKCPoEBs9gPWwOCVV6z1aioRJ6EQQKkNZfqCEcXjD+whbF
256T/Ix9b3rKrVDLXcMUqN5vTboqQtG3cgaLoTNpQ2QQG5TP68iV2GuUXmbhGexK
dwdSPVwGkyNbGj0auS2QQRwF4hMp5uGK4gitxlxJDvwhHxNN9OoHr4v69yhXggAe
WEFiQiOO6SrJ+Ts0VKekkiI4TtsW8EIzQGJXsefs4rwWy8+m8v74/GIZnrbzkrKO
nwWcj9+UUyNPkzumYLYusMX6447kVDiGzcLK1ob5CTQBoP8HQQ0nHFM1mLVg9KmA
tna+MkXKpS2BA7vDlONRh3WnnYpZMBHbPduw5O+4hogjv3Wn3CsCnHUmuE1ogWwg
B6FvnuxGpOP2kp7oYAIdoYGYP2YiQKv9MW0jn0j3Tst7bwFTxRpurfPydHDQyTdZ
UHZuNCW2m8woHvqhR4MJJnWRD9JLhD5XcJjDkyROoT+EmnvkQG4XJzX1bi+7obYn
dKzWTBHGS6jUpK7HqmQyTvhc9PsGIhcDgmgT5+1dptWwZ1+6fy02jGFujU3Al+8s
CBfdgzj/aQd8KqscIjWKOZOI0szPl1v830xxLPDcdDxkixCBwvW5P2tQoAL34vgz
kJTbNKYR5IeBxwgBQNbTYyeju39tmjlXGFxqrd7yYxagrAPFZsGgOMVSzlBJmTbY
nhQVF6RWhm0G7J/XwLSMGGn7SUPH57Cn+EwrRa1d8CA3RaqPl/rpVimlW7Nud8p7
pIyfiaPcFFsW2+vtmle8lPP6a7DpmE/AAnhvk5lluyvBqhHFvQ4QHQyruhiPkISt
fczWEy2YFzomTJtcYUhSKRnoTh0utW2E72KZjlmyVT5svAybDZp5uA07jZXpqk7g
yoA2cjLhMkvPO1jykuCmxnUBfO9+S77nGUoPpSIIAsg9hA03jMvE5c46dkR4hHsp
EaYxFkJ2tISbfZ7zcdjqlSkZzaaEuFOinSgylaEtt67VpmzHHB5SbKK0E1w/htWY
dntTd2y1+bsE+TvqUkRJclArXjCM/YtQNl4hKVAkl4beBOXYxKbaAGK4N3CX1iR0
NnMACA2wueAG/Vxoo9kqqLPkXoEiEzC+LUywnYdPsLzDXuOcRLnRBHGzPHxoU6Uy
RxJ2kuy9MC1MaUFlqDMPxBqj6uQtb9/IiSc7rFKhVTiDq0EiR2wFzZRyp3yvbQEG
hCqopauCux664nTJbnpSGK6MdP0X4RSv0rKo6NgeByQDzhr+zUBMzObeEstsuSd6
TCweo4H1A6Dz8laHdvyUTHERKa8sG+N0TgguiF2LPvuKTJjZc1sb/eBgQ07Ckm5+
9ywtaPdkjjOjGQrmTikiVrD9jescmFkCZcSkrTFp1RjjOVX1FaWnfV7efHNRiUx7
RNMdnjt1+YRPg9C9oPimzxunb/ct7066uf7zOgL6mpv9hsm4MU0+4GLYFpAy6UbA
OLPWUaDG9ieSAkNz8Bew0gFNWy0hk7caRF71ZNMXIiAhY98r660/ihs+1SFmQoH5
TBnY3VXnlhOeJUFHEw0Ce88RaCFmyO0qqXmPpp9lqw3pO1aNJBuDz2HIKcoy6EvN
JQpzzrtziCI0HXbJ82p3dCudRGSnkUbR0tzBr81i5Vr4TM9tnwYZ2BLXGo7OZxyC
lW1hIbclWgP4cvDCkvhLwao4dg12anWzgpQrQ8WSEmC6rDSZuUEIjAnLqLtHnDbc
nkGw+/Y/YO19X2dW/nPBqdaurqSjXSCs5w3d6zNl2I/IxV2EzEBkk+6lrA2NuQp+
+ov6OkmnB3sXIJ1J0GAfzIs/eJUFDWQPIKUPtC+dS8Kjqw4Tsa2LqjsfweLAxR71
9Q4NkkkpIOgEEXG5bqjGASUHrcHU9JXM5DVoCpbsa1t6nkvUOVmOeFiq/twIqvPU
LqMpdLMUmEVHtLXEorPjcWraRxnqY3hpUXF3XJcijm1SWA5YSFo9fb/TQaM/r7AX
HRRKm+iagVpFcXz4wJeLXYLnVetZw8M6YLGdRGX1dgd7pJSKcE1D6JpWTUcLbkUf
nTFq5c//nVkEJlv+TY1xXw/niNLUHrPfOKIT0I23HJ62C7fjgjivUhkDTw5D5y5e
szz7dbsKC2MEbvslTlCl1rCyZhUKGHcA9UxCdUeeTnOdBxDXg+Ok+ApLM8gGNJM6
PsSkTHDOFYSYzAFENqfFr0Elu25YMpHYd9jfd31sx5PAwjJLxsti2q4ZBVM1BZj4
CVpi7rjxb0AmcpTcuYGhhBkeNSMxcOMTd2q9L1ZRsYhY4HuAYcnmjfauxcoUd/HU
LsHSk/UxIuco7BWXmV+RqZ94zUywHqN3iq42JlTtIAtXQ7QJcF6/niEwwp/79Ovc
bKkPKydwdpwfOhMIX46JF4a3FjMAFjmpSLYf7TFO91hyHixincHQGtU+jVu7nBUG
G/cLYuYOAyzxiqnZ+c4bIkxOukEAlrOiFUwXdZ2DSyjg2371aXR38dZfABhUIwEM
Ih8brvhZatQQZEObGO1YCqmjdAI1CgUYwY1MdWn584D9T/FccnL9rdE7ShawN1L0
tctPucSCcgxb9V0y8XHR01nSne1HIUXIPRrdGXgvE2kYJd922CIlGniUUL3rqlk1
04YuTZP6LTqKPvemIdqLhtvxOxUhrRL7DkFTPrnXYwS399Cq9C/str6F7KK/BdXJ
A3j8M2nZgArJD9OQUAl11jPlCaQZbs5oKIxcWkxbHTR915NqbJ69NV7mNzLJ8MxZ
QygDLSa7URBlX6Pg8/5gAdUo+naPkL6HgPF91uGRDGfFbf7Ifm7KoNk/4fqfwE1b
GLcUIRnmLj7fGsP9WZlxlag/k8FlPc1JM1MKbTRKJNaasAQ+YhlSikhpgUA/Fbmo
Bg0th+g12qNK4YbkjcXVV9vxa11mZazbTY3foW44FUICymnvU7sV1dIvgKAUwNHy
5lNgCGajuLn7ye59bYIleW/dglObE8aEcB8FkUCh6IHJUYphVVpFlF59UxHkNx2P
JqPgvmUwKXYnBlRSdvn147u7p8DYV9yPyFfn4KIoum6Cn1z/3w/ukOCml5DjlLZY
p60PTR+Zst3j0Ni9bx033iqUDxILfVrkkiVQixw5Ke/FJWFz8c23a2wKZ0wDFk40
2vhp6iLJYD+lMYo5bfNR3u/2yyuIZrob0f0/Vmh/B5vDdFp+IGOPmH77ezwhzGMd
/Ic2k+E/YIykaBTtSphzkPlhbQ73fi8O1Y9tO7RlYD4yvouCZjGYCTMk7ULd8PHO
zFYiP/i6aKWvBPY1pIYq+MY7O5QryT/4kFrqk+9MM3eQBzourjCMa5cKHM07e0Hm
kLJgTAMqBJsnLaHsvh9v86cysAlCHJo4vD5KkXSGrXHR33hTyY/awTLSHBTx+D7g
tPHXiUj3glDCfJBdvQA7z7WQWHp9Ek3xaR2JjQ0lMAKbEvfj0iUsqYmZ9fZ6msft
wiurF3oO4JZkAUh5s+L7uUR9kDEcY2qKojRGw+71LAP1y14Yzl02UxIHfSD8p3zA
AGCR2dpynFtoz4OoNwbYyHt+VcfckbkHGRlENLbxwm6qprZTa5TNR508ZCzW6aLp
i802ebkeRWg8rBAWBD3zVPGd3ehZXcXptq5dE6qB8Ok7u+guUP/bCsFMgLaciWTS
lP2yMRMh4sSs80CaKdaZ0KdLcT3jQWMOWmcrdv4/akiC23k+MfZw7IN5HAqKLrcm
Ag8XyGlOhPPVOcxkp81gTDnA6O5QjWmHJzxsba671wqHMTZ/UEWXRDAN86p0NmUv
NJRgMU/J+7v/vV2lKU80XilAypsSz6e4AiyVATiF1MN/UKwR+kI4jC3KsqKx6L7i
GxFbhRGP76lP7/lErORSSqEE1Q4niFehFYDuc6LatNRv+nAiTmnYeY4jFy33DSAU
/b3xES93lEEJYF+AlUIGaNOZka5tSUGqQ7Vtg1pT5SZoQsOMEe8OI84rlYGMLfLn
o4jA84orrGHz+981zFlewkwqLnh5Ffw8EOvgCF4FzD1fTAazRg7RAS/ThDFqW9Qo
NywHtkZIMFHHyVRtL1Cya6iN04ubjStV84Crnzf/cLil7c6ITsIV2kAtu8DRvp+n
Cl31kewuWlOb6ptxy1xUE3GLjSlLm84YNRwDBD6rtmPHDXz5rJdXBeVDcBO4faKF
7/GNV5QTKC5uLIxgB/q5RBkuyx7su9L32iFeBiK1XFZnrm9LxZJZO1argPEWWjEY
cN4PdKyNVwA3iJy+dtRcEaxO/yL5VVEXWFxNq3fhnKtSyYJoX5vbuE+V/4UQ6/4w
zs7y5JEYmB2wsORpY7+MU/zqewqMep5DDuPtbKh3thDk8PpgLEy8ozDJ4ctBhBdj
U7s3he8PRLDlg5h/yzaRZJTqGOUvsceL7ksSad572wVT8GSPuE+p+6j+joU/+/zx
SfXiHoQcFqfOjTPNBhuTkNSkYsZNzbB0BX9KNYtZTfTySsWl4vYe/RXj0KRimdZX
VAklXjfPAF1OzRm7/BsXu0KluFJdtIfSJoc4X9CKOk49lkXdQMzb3j0Ha2Vn5C3u
NH7bRo88mLVahumrNWDD6W8fMRMn+Jgi9ia80XSV5fPFCSqfHbZRa9x2PndoONZl
06IS0iGJaTz29HPtOI5NJzW6rJNUqXhsa7N9HzHuPp8tQv2pDZoo+fTENUZHgjEz
IX2k4t+klvoS0m7RjMgKXAMxBruk3a7JvDlSfU/YcfpUy8/FGF9a+UhVTXxneW+8
hPGC2GgdgOLwL3vZGBEoA8SXfH3vKFnuLCajLSua1ocMCDIsieHi2Zh1hhblwpfJ
mrQrTo9ipOb8tCeh6uUkUGjmsKI0Wgn2HL9UBXjRg772pV4d7iZR0Sxm5QyAMZJc
5+RtPvkrb7vbQFVIE+pdcYA4+MvQkYZzXFvCR6syCzn8IMitFHwQQYA0FboyjQCS
eMyrHBZJkxgSEV+T7SV+Wf5R/6wsV6YSRT4qx0jqlBLVCDx2UX8+8R74Iv9Z6E7R
zzb8XC8K3udFKDNs0TkJPxvnINGxZf4TvHDTefp+kKx+RKx7lsOhQ/Iu2atIATwz
S+h2fFHtEZ4RX4EwLT7XO2YvScqnBUjDMRlbhffU8cKNPoboWPLR9/9Y1cdnCP3y
Vhn80Vuqiq/QaJy7JRUc2qvAJoAeFYcESPozKU7Z2jMpCEoccMNy0ZqzXr+j0eip
P3vA0GAmjd/dBT8X7HVZlMbFN+n4R06zikewPvbvOJOc2fK13YT6c3wXrvvMfnrv
OqES2HMQNObALaqWZ8stitU+rBOYoPZ6OzmUVvgfxsYwLxQv+2VgWW8MQHsFvEBq
p/RuwcFuFLR9cTHx59+SWsp6z3cFC2QaWMH2Qx1cHOHwD/c7emohtPY58va5uu8K
5S2DrNUsNtx1TT3ycgpxJMVK7Tu1bHtpSVqiMa0gqQq4oG/62IGh6hh73R+79PhM
KE9c7V5Ugy9Uz4O0SQbvcZNb2XM5DbalejLUJRsir2nl0dbDnCcdglCJCG0q1KfG
rz52KSzomHtz/0JrDjIIFrItZnwzWTO9WRka8bp2aLp7GRmVNt5jbnizGUEF8xlG
WBnITT3++WBiZdnp2f1+S2j9LOpMLQh4Mqcuj8fm7eE=
`protect END_PROTECTED
