`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UzS53N3JCGuN+RLLIsWKgCZSbCLBV89JzAB1Xxn7NKVNT/2pn2zXnF+sN0cR8wBA
VHOG75m6Qffa513gAS4koqJKcW6IaQ77ipI/qK9zt2TwomvCJ5IgywSHF/OuSfmJ
2x4lsQizpfLSvBNmqSq31jLY4NTOdYSpsIE7HJRKl1DUBZlTWJlkyb+QdUjKgnQV
wetYrpjk4c9/CF2lTSpcc//VzkjZPR9i8127nt2biBhu6wllbUWWq6N/WoBAszfQ
k9oI4ND+Y3zxaZYtufSOKdYCJjXYyEFH5fdJyzfTuCnsZmANE7Ib06lzherkJfmu
YOPVjOQJtgsZBDIc+ine+cCIpRWWGX0Di/KTZTZair+I+dPa149ZVSe/TOh6ewYz
xpPohL0+pQmrWl+ZY4hpceyRwYK3cHZyOhriwkQWW8RCdTRksw9srUpRf6Q4ke2w
Vc+HE6VaaQlAJfTc1Y6widSa89iVm+7GDP+drQnoPyTPL6Pf+u7zp5kQY7LkFcVP
V5z/Cr3Qg8+9nOpAg9gmY7A8gPKx/V+9ncK8is/95meb3Oy+RG1i6D+EpFKQTa5v
hqSIOB1VLtMszK8yvq32X0aLPqlM6JIMbD5ToT5c67X8jbvcdYNvvIJWIsb4BiDg
9snZmNZpzoXr9jr1aiiu1cMrp4Vhaeey1bmyWmZSPLIRceiFjtHr4bJpjTjgnD3R
a+3j7nqI+69udQfEpszYLSV9JW1NaqOzQMn43OVyPv10f7QPedeLOUbinZIFlwlH
PMEQUxEzLanHKUWbSTlBLLh1RF9mJ2DDWKKtuSV9iAxB42nFiakE6Aa9Qb2E1JWo
vXOpgeOvSEF+FAAkSwAI28vj44uEPkVwdd048ZSZxBqo3kW8xtoLND0oid8Hjsv0
FVQxpgtKrPIbXQgBPkJqCx9xLnQC17kDmkH3EiKGcaXVkFNZwFwH96xbJOrUA/ZC
sZMQ6Usd1Zoq3Q6N94Iik/jf28zXeR/F7XhAtXLA16ulb/LlQQBzgv8O6/hO6feB
fxs6owWES8AHnurm5i6LWPPuFAmkg4lVEZD2XtB6ji253hqie5mfHrvVoxUsp1zl
odvc59qrpBHCDVxtA/aa8ddNARJU8JM8bWpjp8BXOq9BRONtOxe0J7xjtEkaCMKw
cc/2r+qR6Ew1WVM2VovNaTq8nUkAHSSZOP/ciRQMB75dsYz9dI/fJ9Y0ujId67nW
O8EsX2xtbvK+cIaY6fRI0TvH45roBEY4uBz526opwnI57TLJGuTyUg2eL2+w5kBM
ZXHy4SlJIsXFy9i01/Sj7WLQ2lViOuwZC9Qk4dZwlINM3C1JGQxPnrzqBfuAoBPP
1zf/LrJVbc4NlY2BlXpzdDYFLcdXyQ11SYv/Wmf2xRqay7FOMj3jXO1fPizRH/Nk
Wf58xBQGvouSm4JUaBnBOAN6SilyyPlGe0tt3zIfrJjTEJieEwKDgE5QefgpeZ0Z
TULXlBUF6OIJKvOgdsk3NpSse/JSpWeRd7nnvLMQ+2Lacol3JfsqJ7OEBkQOsRnN
kiHgkbTMztF6c0MCu/F5L16qnTBkArAQrLfMFcOIjSjU9DT1rqVKYTsE2kechoDU
NV4+/UL44uEYA4iPYc5GB4Ig7xkdix5OdW1XhdROFa7wZxsZEBOSSGZnVf/+VKBj
f+RKZEr5p5TzxBmkBxV5/owNmK/KkDOrlsKXUjl5BKmKz3Z6Cb4MDhQb8r+7ySbe
86sS9vf5ATuLziYFfiMoq+aShIXh1dQDchqHTByIty7RjEAf1B8T34EnOZexv0au
WJxSektE/FxwG+NGyRaXezqv4xDAmd+JgbREGrpDz3SWxmJDJl1RkWd5Ix/cNGaw
CCkzRsz5yoRQ2HCn5pwJSzAVr9FOHOY5ptRiqovrkSA6eSv+mOK33TwdsE77oqCW
cSL9z3UnksBKcGvhpTjtyGu/sAafamJCOk/MYTwNFT5KQkxZa2giEQAtmG92wpSt
xmjRcMQeqL3huzrAEpob/a123Fv+r4y4xBp9wtcxc29u8mb7SKsm16SLeDCU8y1H
z0NT3NwuUnuZjOgYCwxvvnzNMXKLsyuJhkmf8Nmze//3PMOQBfjUlYDKqvuJ+AtS
YaFQmRhj6hkjXTbagleYVxF3hw2BgI/SXlkDfKHJLkoIyMyy0d0DPUmPxnTP6f9c
ofKPxABoxxOKfnmlaWh69SzSbBm/cShM/Sk/nwgz5wSJ08Va7KsL2aQsRHjho/tp
gVOHqoSkM7wcUKIkovMO9xFN6eJwb1TOxN62sqfzUxmzrnlj4Mr1w2tAkxA34qEl
PgH9IFYVqBsjm/u39cBNLoNfOYYXFho+dr0EeUCQDRfiljGr/Dds3v6boOA/DN+m
rdwp6lOZI2fjA71XnyTpG41bWVCJq6ZIjooVmvsFI1gsZ5/VJ08DIYfexQIBOM4c
V9raEUs5HAP49jg+puwJVMdElan3y4X8ngrnYqU1041x7PflI0JCsgzAxiaYcfPP
qiCQr/ZjYN71wGP8Gwg+XLjR9uQHnxZNyqOkw73j/1bHUV4UplZzFBMEFJXMgAlo
69H9g3/Dm/MVDDrQUpLDUbr1crHhmuq88PRUSmDbxLt2lnih498/Tr5krZntpN+Z
OLvMhPVTGnLWy32pYpTi+SX19Dv8136ZqECEfjp27CGWINdGiXgDAiReahFoqaPq
gLyY3ONn9YJqdp3svPNXCanw9bl9cvJQHBK2y9EXOiIfXWtJCBR6CmhiIW0GGA0Z
yUx1otGGO4/aVbaXBUB08EW16qJmkDazHhv/nS4xpY3potvtiECiS0k0EO2FhC06
6jJw+KMprlQjtngwWA5rA2LQM/sz/wHJjK7TaVlvlfjDIT6b40KpiKG02u2KTazk
JzohS1n3WIuXBe94cOJT3dxGL1MDzBmhaxyD30F8tZc07N84OQEg8NJCad5AtTVQ
IL4MBs//Gvbiq4yqt884OsPBzgkmkJNxdBZ1FrjhRQ3buxO19Dx43Us61AIExv65
qwfskBmMfd+BGbaxv5M2QaizVAI+lBC+z7sOgvenfrNcV5kCGxMQhNOYwQK+p4ON
GnhMUQOsy0nLy/ia6s/EJTa76fR/TEgW/acug8BIMs6eyjM/DbnrxyoDwBEmJQ+k
+WfM6hzFYR+QZt4Ovogx7hlJCi1uNzL5XMoFjguZLQrotr4r9LltfvRi3yxGKqg0
qGthupG/KsJbP8SeuwE/zNHOrTScon7+M6BE70jY0uZnceSn8aC0l+3nHafH2Jze
RnJYqVTVyMQKVXoJUczzhkv6JdPOorzDQOno9CCZlICW+fTQXQkLKH2w10cfEcyU
OsXrjWWcQPmdqIDrk6GOkd+nv879RneJs+ZkZvp3fdiOtGEtXUhLVByOvluTt8HN
iU38LcG3417fvlBXiVnBClhtQBq0eSmQrZaL0TzuUeM75OYggy2ssPsN5ok+6H6j
44OUuN+mDKCRoG5wdCAXjjNJUNdz4xUbFoMWUwjsIiY5eqJG4ffPcKIwF5aVbDXV
Nvywd7biZIt+fj0kYtUeHTyphvTHS9ar1lFZ6Jx4YmC5xSsgl4x74EUOGZOczMW7
2x6fJhy+M9sHIl2zcG5SsRDWJbAruvn5EzPandqUhH8QFs7Eyhla1eoMsquIGYmL
5G7WCn+ooCMFj321304yDT/hJmET6njz9qxjVwximUI=
`protect END_PROTECTED
