`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iuI9H+nh5F57LwXIqDPoxnQla2fnAtSr2I+Q0pfxHJSIPyoMZ8b+oeAxXD8n07zl
2/yXVwDW086JnjME6FM8fgHvxMyGFoSK48FTHGol3kpVQoCRC2/BIRzGzC2txFQP
3Re7I6sTMYZ2DRZjfIp6D3Mdo9SPLvjJuwVK5kPbOZiORCa/MltrNMhPDQ6ZdRJ7
BcncmeG+zI1t93/KGitXNqu7N3YAeEq+q28agdOWs7pFdaj8LPfBOnxqTtAawjG7
OxWjZ+7mRJ+XhbvOIH8NjepaUJEfCgY/dmMEl3OhLpkxEmhppCuXkhncfm/QF3m1
OKLjSkwXVFG+mxsTkWc8TtSJaj4PiFti0MUZcuhylrXYqM2vGJKZMFBceggn3jx5
SeLe9fONzjk4O1c/CUd6z9B36oUFvEPS51ypf64unkhQCr/27k0LpxDZJl0x7pMg
zfX3CjRNJ5sMlEsxoZneysS7qWUBvnnAuFEL+9PA8tVwbDYdrsGyEzVcp9yKA86F
IvoJKqVtVQMaBV4kiH+q1lR+u+AgDaobrq4a7BABVy/oeYgCcvEQ242JQf9eSgQI
6bRTNYIci9BNj0FkNrIgxvJeifzg1YJeYcBYCqjSiMaNrh+68ZjnZvwMgmWduSHt
t7iUBj1bZ/UKeTrmBnHJUGfgCCs2EKxBnequf3/6SqztrXX729U021Ma16dBcVD1
gksoWNOE2FEbKtGqCKCQS14RW6dlp/E4d7RqPFro/65iq6p4ZH0D98HdEUIsJekh
VzYEWbTUTONxrvLB2+k80zXgPoW7IBMiUbkXEYa9TN0ykjShYBRyWIZvF1pZGmLd
G9c4y6a9Jf21/h6lpYYPgpeOqaywsSh6d+/hVmRmO3MoP33gmDOHvanlnCOqWW3u
osnkcS1oKMqvuBqUM1QXn9vhoync8dN9QtuZIb5IQv6rH9CV6FqdsoBpmBWbehq9
xAkzjygKJpwDT3tsBRe0cRUyAyj9S6GeqtRkwCBB2q3WqktiRykufwjBTAJRh7lF
1DnrKBS3gWzZUpZ7EKwFWdiINTIphnjL/oWgKo4sOwkfF4mfVGkM8U5ORNfjOhwr
kq1UPXa8WhQPetOT9sK27Mt8FTipcN6tBTs+qbUgytAcWybjUAaCozePwDA8U7PZ
h/6/dxBVN2kX9SVL7PpXkvBFzeSILBHzlEJo6AoGFfL6y8ea0nxWnRJO2DVz+diw
FTu7qLjvNSbbg05+jHU7pJyjGaUwEImaedBZiT5WqaS11va8kDaVbC3jWj9Ofheb
ipiNWahlyhUxn3UAnakgLnX4SI97DZw16ZYSBHcD8zqkq0Lpl8078v8nVt5Tj+mU
23WHxxVdIiorzjCzpUe1MBJI64a3R3q2jxe3WG5sCorJAWr5eZTh20iGzd4WBU6J
6hBtNWQOpQoCVpPatEmoiYiGUDosJAT5/U9QKGHnRRc5nIajmcmIa2x+aXG2ZGn6
+UQ8veDD2eVWV4qPcc8R92u4ctGKIODWcEi+wOxsCM80o7aINRujTmDALpz6q/vi
bXNdH2DRbxKU5lnlhP/uyEmCJ1QZXpgy4EQYY4YxPg11R14DscqbU0YNn41sl9gH
a7tMPk5sXjmjWqC0iYEGnVOFA2aph+Samd1Z5iBEwdm8CJauwN8x225pqUhCcgvr
3s00zpY3QZRsI6EwVX8xW+Ha8+b49qhf4iQZb1iYHtxLDQGpbe91GTE9m7OY+cog
TwV0X+wgLKv1NqKiTDw3Et9h2aTQ73tXnBsXGQXvEXsUK53MD/0eiXjYDsryKrF9
97YAu2hwTCKkEUCEDlvK/kVRG20R48WEESfmuJJCGRRqu9UbQG5/oXJ/xXwugOs7
W+o8qpJA7LAgbrYEsmv/4A9UgnXORfxnXDmOj57qzFvXBzF9LHxMZmIY1kw4fbzG
dus/xY5X7qsb3NP153DqOCqCNtLDktCQmsBk8Bj9+yu3VRABWFULlHaAa6jFcphL
G+QUup2jlBmazjr75zklIONUptL9MV7G2kf7muwhAZdeFKsLa5+qmy3l5/9uGhuR
s980PHG5tKrHFm0xSYLb6dut8qx1DVeki8MhcEpXzbiSbqwKwbKdv9yoDw35tD5u
6svyU6sJLkv/djmWYG+6fFx85b6s/KCjWKXCXsklYykDfvxkAY/kUKqctxb9Wh6Q
idET2HFzGOeJ3WeR1jb3KYclczVZjd/reMqloNTNFS8L3X0l9U+/9Jw388qDi3Wr
Rr6NLpXH96TujVMBtInBdAReSbjhH1ohU8XU3miXyGwl001qdvHWBCzPVyWUmi3Q
hGfa1keAawHlULSvtEidAOS/LnE6bgEIi9EWMIkVZIQWbkOvv1bNNhkyBbnKWctv
UF75iiDKKk69Q1bsPTUIbmXENtgosIZAUrFt+envyOKpaLB5NMgXqSaIJUD+RJAJ
ta/oKsYXFx3oS0jpzsua6z0imfRAEdeZi5Q9kyEO1zK2k6sLeHonMy6n+0oDhthv
mZewz/7EkshZSanVC4U0K+lqf/KOpE3VxNkpw3YMggln4PIgZBL46nFeldLg2QbB
KgTVLIidf8PkNeXMcy1kdVBh3dQpCt5HlfzM115MPlMevPV6AePoYpp4vDp/XEhj
42b0Yk/37g0tra1Zk+IxBzZtASJKSXRKhOibIo+O63PB9K1Z6jgmP36zcQXaUufQ
0pI7sLwiX7optMj7QabrY75PTTTFM+FnVYvFT1qyE1ZjM+QHo6x8kYg3/YaaH+tR
7U5EodSKEiVz12wRxGvhmklC4KZ4ti8P3YJePKgVaDx0mYYdZtDC1l2ATsM9o2du
wU4lstesCzj2d5agWNraax4qBYMdEC08sAyshMjFSnLju2ASAYCGz/2HU+Dd3fJj
3g0Jtk1h8ajjDx6063jNQrGU/Rg8yjXyc2GYoGv5Q4pw3hLdI18UWT5h9Nhpwgm0
FmYqsLZT2KYueMFQxO2xBjOVZ/qron4OGqlMuh0QKRadqOk0XgiUOOSyBgfT7jf9
umE9dO7b+so6WuIl5DQseJ9fsfoJu/uWBcRyv4LSve+lo8byWGi0WPQTBJXSmr+J
jfXjquyTPMu6ciGIhfMhzMkkMHWTRVaRH4ZnrbKMaeI2sKtMl8jWTM5f1KVpNo8q
9MGe+K+We1ucntFnBREBqdNvN/jTNYN9zFhE1Kdxtk011sj9NkeDc1bA4jf1z1XF
5QdV51n/9BamH4W/1RgoAa5mel6QgwCtiOUTZPWEbF2jEGFnK/rDyr0Vak8c9Swp
4+M3usjvAh7psxUVQUol6cyr+s7FmM4QfCIPcV3hcsTTVTKV/MTk5TpMcOCiS5fk
fx29z1BxTaLREdqHmAh6JwcM1A9Ke28VA+nfN3KLSoRsixDue2fK5TS74nT33q/r
qsZXD8KGWEfF8aj6reB+QI7X5VsE+CPJNMQ3Rohdy38G5nqp+00Y4BAu4QKyBfaO
j1oSHJMJBbtv6Q7/VjiOtn85yzNQ7DeKBuCwo2WoCN7g1oV/x/MtAVg2N9Ut07d/
xC/B2U1BFBS3Lqb1VkBKyoMqEeIBRanMMI+8e8hrmONXJvLsZMroSJCUzCUDKoWx
HrIyEw22tjBZHF7k92pX9dhH4NQBTodDWFwCtGcAkBGIvhIQ6A8Fff1ewp0bMyrQ
jI2oNQqCITpnyBHZYpafPivCbx2idycd9X/x9VusQjLQ87Ql5KNAbNF1UEYR6D1T
qsmNsB1aYqNIr/0RANBgdCTbB9d+A+UCX3ayMCuvvr2uhaKDJ3QvFZg9ObpA9/Rk
CnZWrAYMgxkbdFHcJIf6UXtncb2l9lqjOUOV7VjonolF1jvyG/dqGrU+Ozsdsari
LrI+ZCr4aG65CtfY7xO1+qZtxlLslGLtEeCYlNNwpLTi/U5P0XF+DKMeSGX9h0J1
wK+WHDGxTyfKw8b9JtfZeO7Cl1z7lJXyenNe8jC5qYfvBJmTw+Jumb5NKnQSXHzi
VIhgxp/BeT5RMX96LXuIE6VGlzsj2NQY7zmvGoLiYeKHxMZU+PhwFa+vAqeUF+ge
OntVbeHe3HfsfCLY3SBLckheJOMK6buZmJgdyrACKthA6i0rDWzn2sHbc8Dmt8st
kWb1jyWssRpmE7eBJ/1F1EM30qTQWOegK2ufTN/xTOUkE2p2IGfP/DKKMlnup0Pb
VVfaycbF37yULXrqM64HwlZVjIDuBw2xiquDOZopnvc88Hwh7C64TJddp1IC3zXj
7IsuE5x0fkevhXh7wA6yXbNJDxBv0A607xhDI1KEPOQC2vEa0qe2N250wBvlWvsX
iVSDCnfRGfTL0z1uBb6HZVty3Sa6+2MJyvHmdmXJDjefeFO345yu9iA+8ZwAJaIc
zGONzD7GHXchO4u8+yUmOMJGP8HahczXlQmRsylaoR85/YHzKQ8zZmT8eHwBnZ18
Bmly4BVN81mOCAHT0DY9gPgU58QVbzO1Wy5PvIWPpiKu5rxo9YE/90snC1YpfnKr
4amrlTouH+neI4iQOZ+UjyR+KRjmGlliYfEGf9ruG0mJkvyLXBtwvVe+FrqofKLf
bVKLP8QyBLEs9ekze7GeO87VuuRrF5nnmpzSzO0t2BnCr88WpIzHZWudRgEuW5s1
eMLCbFq+cwx75tOHlVEgnvW6k/QJ//sibxtbvDkB1lPq/lmxVWa/Qz9stwdDMr6R
E4b1KMVr160duDzpWz7BXIJpQ/JzbXgd0/ED/7XB+M5EIbS6T0nWrFxRbJlaCd+t
24QNDdmW4m1dSXFTe3MPFBRS6y1ucfyi6lAJ49HD4VJKmoNExf46YY+pK6PAw26h
tLd5ljRIpZkmwk9f9jQGh5sd8XXvgV147+DutkQH3eAUmcS/CBA5QCcgG5SUqcWg
Zdh/Q3TyvW1zxkDoxon0E8CbgKyDMUSYhN7uyM1uot0pL1EpfE2EkJE2lFwCtMHY
Rcj2rX+UaYwXPON6DuB1KjTwTXVCGTvkxN15Pc/snkScV0LhgxPp5CK/yksDEuqD
UyQ190mbsYDjle9HzE/FdZebSxLSaOhtvCZtIO4TeQMTPdfsCXqrmKIx28IjJtcV
9+5epDCUT9ceno01qNn9/06KxkEQzk/jYRUow3ymS/OF0vS9d85AIcxyyUJngSTy
fgMntgLl+JKjLbgCm8wj5/oNtWPCVrqDoWg2uZYIEyIhBF+JRuNufCcfUEcG8pHj
Ygbvx5uvQroOyWJ0ZrCvmGA2LBKZgFOCDwRqabd0YdrS2J577IK4Hg51tZ6ttT/j
72RfsM87eu+j+190Pmt1s0ZDAHCCaUIRitjiAadIYSwZyozjZOMO0jnMEfV2EO6x
ytmmlazKtqFSJq3sP8q8lV5exnMTzzM9YFOgNWl9qeO5YFsU4op99Sh2mehvXEy+
Im529vzjIVNyRn6mRsRbKqIVlZxrmqLOm8GjlJr1EiuExUkSd1Pcn7x/juJcgH7h
Yehj5HnPIY5OLeWWvzRHGnZ9drftEMATr/QYArgjaMNyyx+pmwWH6XkBU1NEO60R
HcvUyrYUKrb+6MvoOG3nHMqNSWJH/vhOuiQWAUdkuKIXQKU9GNnpDBugUD+FtAVe
Y4P3HRzAGp48Hef/8Z1VeXva6tWlESa5TqzlvMHEWFdmMcj8uWkXhUAekp7mksIV
g0e4boxRcih6Z8h+VttQEZz02PGCuQBk96Zf478P2oxiQ/DaOH2dlJuWOsRWVfid
by4y6Wd74JETsVpg5wFKls4UhVbNfS3lwL3zneRvcsixRAbx2qtaaVcX7amGTK6b
5B2X6LeLpxGTxfzUi3knCWr71I6CBgPUafLFJ7y4T/tIpLI0fqP2nuuIBahNbEbb
Lym+oV34lwhFWnO9eo5FZtyMoE57U8Rb78td/DKm7i4MPkvun2CDL7m+Q2ubEcLg
H8s+uzFWvNhaFYghRmOho8szNnz79Y9JdIqLtl593ECJ52f1ICg4j/+RaKuiEUQj
INZQ3UGoXAQoq2dfMdicvmQLWRRIeSAJYiUqdqAJ0YSegCMIbDco6nI+Td6WO6Oj
vXmFo9f67fo10Y6c0hA07/+iSIGvncXGsHfcWMCX3S98rQWYMLszpZRBcISDo/sB
3Kgj+TdWjFJyxohc52MAQaTABuEP+u0zyRoZJRJFhN2j9b+Uuaa9ODvOfk//sS3h
3/vsjae1A5ww6WIfXgChhU1RWz6Yx/ZPKP48NRW9eZ/kjHKp0WppD6/fYzRULslA
ToktmMakzzp/8g9sGartEgDm80VuaI2Z4GY3DPIGryqAiwcdlaORY5Z9XxKabimC
YmZqeW6LtjFKj0/8I2o9ncphPbZ/m2yR1/aMnicUBf6ze+21PoBUNi7BpXVildJm
+Hc9Oxx49RpSIlYMC+xXHloI2NM1GCQmXQPNnPo/N/VYc1yXYe/H+peoqQYnelO2
zVbB/yJM3dBirT2lyij4VuOgoD2kTcueXVVy4qWN0VwsUEIen05wODPvrShfLjpN
zrRklMgpRv/dDa9CIOk6i2O5Yd7ycTuJwKcAxpbhY0mQY0ZzxTkY+NwA/abujoQE
tff/bZbjpKtkfq3CZZEu2ct+uzDD8C9RYPuQYVQmkxROly34x39+m+U8JJJTd1Qi
AISVMpW5IJ/EcKbGa3mj9yrrad+d5EfkZNAgO8fg5xQVbRXESm0mVFY7OrjG5i0l
lVO/pmfShozlpcquX6YF7zrUK/VYVXvrHDDOu9z1qwBh6HwNN6Je5fp9fHNMXwDn
wZwdJTINXs8iYBNd3X8INz/pAElY6gfo6cG8dqThCvr1jFmoLrIUKW8DsbbR6Cjb
7SESx1OJxdajOLSvyj6oKHvs3ebP4+NchqhjnDIAkG7sCfjrTK798qIy58YNKJ3V
JXuaAkNoKLau909fZW3kbcful670VONIpGikxg5m1UpeJKiXIgG+ALAttsuUp+gN
KXG5VfJQNZJ2mCUUedmxVPiPu7HuuS1W5vACWrt+nNpfwCptxXwQAB7bxfPbfSqt
W7yqboKtg1nEq2WrreuTX+1ImHo5jFyTisiqpJwGkJ5M1mg5RAIiJGNMig303paq
uhp6DO2k9/zy1gmVQNaZhmZ/KIMiy/oGPsDolGENEyjRJXhG4cVm0iWV/y6189Sc
Lo7rUmSf8Y6pQZ/Ui/FvR8j8WVkJstSgp7pXyJ9+2S6w+n0NNTMFFgXzB+xnyhFY
tBUy2feMKMrYt+51DVp0kQesMVIpaKDCPOqJfpgYtp1ffnCwKBCtyGjolJrOzbGD
rkpSI5RUaeiiIIPdkFBRYMGBisSQMYATazLn/FZGhrBmC5Zs4MKYEoJ/hPj5XAxk
6Ic53k9yBT7nryW192nTA50gbnwPC9D6ArxiuEVV259DD9VT7+gFQe7gWsrfdEMN
0qbBV3EUL00VAE9PIXGTicKaDwL3cPUWhFhizjsafNybgPeNzILquf7XTm5MR4L/
9QkaWTVxgLmY6ngXbfqTbLVMufW6xn1u1piWlA8PVNHVrV1Uzb3NZB+sS61hUUN4
lJsHNBwaRsALcuKkl4ZuIqTwFwNMwTQ3JGKy5kKjlu0nT3Pz7I5zla6G4jRnaeic
7G8kUmmQHITPgZn5O27uM0qyjC3uS3NYdXc2fBl/8pxDzNd6YiSkIepatePal5UV
Z3WkXweb9Svhb7XsmwLOQYhX3o18csdQ35zi+cQJNHrzjsnSa1YtPhxDm1XpaDVb
ryPEejhboDJ1I/cL9cSWhxkBUhscV5WKt+LLfGBQs/ukbEPxF/h8fVLLLZ4Dptgd
VROae92Nd3NA6+RWYbRJCm3FobKCKZMl3dQEGPwJ1OV8zDTBc4NB/OcnEqiT3kCR
2TDiKcKXNnfSgRxVTaB+kUUiYikAxerSJD63KGRR2cGH8o+PEzHTHUu0RHJ1g3jR
Ie3i5fQ0gPNtzzlniJdDgOlB2X9AM+Pzq8KeKZbaAWr0vqglDBF9Yd9INIgs7SeE
3YUvg4m5A5ZmeVk6m079LuMl1mWZroLfvNJaRhbetMFalGRukgzDJhIHlyXqMajZ
GAqqh1eR//fD/Rvo8xvVzWHxfb2mfUPwfM5tm+NbyR9LOHV5+9vx2YQv3Y7AO545
BLcY5Qg3TvrjWxmyhga+98+FG79Gav8Nx79wPF37l+DhxoiDe5lJYr6gjwNsg6Hy
jO3i9Dv/0weDhvUnkW75yBZ+xuQt0wNhH7d0TJ3SCE5fR4esTKPi6IvL2Viec93z
sSi+T0c2jtJDFiz+CSDyZHcT/KY1Et/u9exdHIZlVagoD0YUGA0uzrkIUDEDiIRc
e+9r3p9pVDB8n8dnNIbDq3KlaMC8EKDc0+3/ND72Ok9b3EnZbyr5wjjQMUyu8lCZ
GofpJbfwg/LYNJawk0XDDC3rNMGv5wrxWpipSHJrgeCK8fXe77bYVz2aUNNk24mL
b8sapeTA+0yqjZVJcbqyLh1sl/KLzGlnx9YUvY/8tla2krNCxgRLyEvywFqkLb2r
vtbGniJ6hFBcyYXqwD43q5GEEt9shwLseJflpwZQxMivSc1zVR4Dsm+2C1Z7tvvM
ek5s3I1r03XwUCjM3j/bWV0U/jp9Yvor1EbGEnuwR/LunXfVxWlx0f40ZHFd6zbv
9yDDY4guoKuYI0cjhSI9E8uKV1Aw0iWHV6iCX0R81HRt08804W7Bw6cOesjLR9aU
++e2XG5rZAkGXyQhlkjAhLT8KjksLZNQUzQHYO3nKpPYhzghbEj9wHg9enTZAOBa
0up7sJzbBYG6k5Bg1HBmD76zzTy4v/bsXLzmGWKGduHdmQXtTJ4Mrq9VdcQDeaDu
v7/xm6wLrV+gGVoUq/xV0wB0qUDrCh3Dy/juuCFtnUsZzgCUu9sDAxyVsDD4a2tS
W3bRsALp020Wsuw4i9yC2aRBZcgQWXyjGEGjMWtBsREqQmYp6tjHtCvs4C5nvkAO
TiJ++5mNQkPFUTW+oexCDUHmkA5aB1TntJoJS41MbpeOmnBvFV3+DtP9/lECbzYR
MQLCDs3O9bYne+eSralcFqRbRcQVc0tvQa5rbw7GHAsnJRY5InDdxHauMGXDRH03
q8917RHy+dqz9/JsaV5bgBTl8TaVcFI2juFZsKELOS/EU0wRwrrjKulDkuLMmFA2
RHTBwSnxgOdVfW4HBBdXFaQNk5hEiSoRWmaJEtepBAqYTfXvZlrq5fulVzKcT+w7
6h62zv+57RViAmv8NRCZjSCN86LyydeCKeNiT2rC9u3mnwu5FsUN+NaXgAxfTjd7
szW+/xpp6tSz0hOBw2bN+12y+MWiR9R9XPdil7CQF4xJfY4wxjCELFrkAGIh7HQC
1v+W0bsdd/BNTzs7cbZ9RP5tQTrsM5QlouMTa+oGwXM97aB67T7rJAey9w1wYSS2
znnN8i/P1om1Hc8QxMgzHkaKg7W0wJr3Fkub0mSCakDQrxS3S3PX9uI3Ht1BDDIf
sdBETdmsVpO+Rscga/hylLjGLyuxUfoZPJ/HrYBY5rXh5rQ8fuA6mAeCcRMBezQq
lpQqLOoC9APW1z7/zx94W2VPjG4LqgmmWSkyCiscOnnAEQuv9/HAba5BMIz7qofJ
Qqv0JDk5c3RGNpO484rcFvNii9crox1Vd6i6oKCMsPzKaQq704PzcdoqKlzC/z7K
VjnbmyLGTOXi4GN9pF7rwbJ1+4oav+vgLpp4yzIMeIUUecE0tCMFpV+FUskMnvFO
/9BYLVTazEVgL7E/MKL42TMK6X6vTCkdOI7r2OLWZq70I7lsRYScEQdutdMQJb4P
66X+PJh+5O5fVMqKcLkSW+3+JNlennInd7kcHOPDbElruJXjAt7HJ94Vp15aG4Oj
89bASrrQmaNMmTQUvhLhW78l1jkGYs3m080JrND3NKG6/QX4no+org8UVbplm750
nThcLwzgneaYKGB+c6jD/Na2dYNoi+VyfAmcnkDQ91+JkfBjAd6ZF2zc3N/KKDg2
D/XvgWqewnjJKUMCeyJT5qBZmc6DBZBCSJx0ve+6yt2nW/DjppBHs+5FmEofItOD
hFhiTyeY5Q+E+trIAMTgGnXF0759eUMt7FenViojLtlxqh2OrgPQkqUy+RNmowXF
HzFwNnOqzH5vcFIf+COsUo6OAISSVbacTSxN8RM1HoISlUC3GOenBl6OIHVD75Yi
RQyAddJNgy5kY/wwCS2VSqNjar/b7VFaiZNTLOXU69WyGzG/Wp7cmF8gbJQG6FOD
En/WVGUPkg8fvgY4jI/9LjVnnf27llpL/mixP+BxOfhrzRbNgGy3O8XGYFar/rKs
hmWKQ2OzdmXL09EkwfkBGBGio9HcBaHGQyEon8vRobp1qLOPNogZf2UkhupNYzRB
TW/oIk0y3zUCLUIw3JouVOkJ9hdh80kdzxp9jNTyz+ryVSESc+Utr9zvQMvQj+gJ
7yNWgEBnGFE7CY2mUzpCixPfKUjHp6EkVDcBjmfof4hlfpLHy7v4vjKJuV5nqfrP
tvoxkFSRMYZD4BALIeV45qSVAHwNk/kHBx9CNasP3zAXnwcLqsl1cI/JDyXmx8k3
0i/EYATkxNGLZYsOEb1iEjt64G7Ke7XxZt9XxnUmTmmk9yyMBQSETP07ND8VsCaH
M1vlVvMeGx5T3zKfc3dtvosIOpxq9GyN0Yv3lFFavvwG1vmbkxacS5Oitx8CIIDB
e2Xh4t0pAmQ8/Iok83e2IA4778HXFoM5Mr7ctkYSXad84nKtlwQKgNJyWK0ECYF+
YJ8xDZgFGVqgqE58sGgQgallPz0o/cVEYrBq0W76VnamDNg1p9RDRbh0bNE+KhC/
i+q+E6jWt+t6EXPqkNJY/6qHJKrj4s0LKizWBkg7q0amfkT409z/Phnx9RHoFDcI
/SgKOMS+B5z28VwENOb4aAkuEolTK/2KojxyT1kk9NJYRpJXZr4E4/2SQkA2nqcY
PK9pfEOY080eIov0PbD+XII2CVeu8hrfTiOum93Oek82+xrTpmyv3EMVXY67kYqK
8oNIx1DHE0yLCcQjKzL6HZwd0ZbpPT+cH8MWqTxmhWjcGy5qqumBvW1DxFvncNzb
EkdoRnRRLqT6zdUi9S3pjZJEm7F+y5eH8cZo+JbSW1aYUeXWE8j5tmTOs6qjAW8u
Ocji9GHSMOzXKKA5nj5C5ix6J+IfGjBdvcWbMZFOIWQmGZkwar3nJiEJG1w6tdiZ
wRmZJX2B9ZJQ7a/yZr/7oMs+fq0YWX4NGELTA8VxzLCPgWjRybCiok1Ig9Se09Hn
kkKyNslvjNgoDcT+cNaod0eo9jJNs67Eu7wL0eAjofW9trLxpmHOeFIV9DEskNcn
G1xQXQcF8NxHEn6omrX33NW7XlbFKct4rC6OoUdEz52vgD55gQ8ReYv2HxHKEVUA
+wRWKAz8xNhQ48AqDCte9lzy4hgE8kNceYT7G1OgD1a1wvftovaDJOW6seEZeZsm
auWd+Um9nXHkCf0nnwegSQqzuVFU5gtEl0d1pZCh79NxDcYOTWPJVzEMRztHxMGV
pTvgcE87MMJ0/h4KmRHL5yN27uu1u2G1RxcFk8YRK+SU1dhzXVjfIXzq6O0kRhpj
QW3Yrrhh4+TwCcHcJmNX9IG5RCAan48weQxnNL0WgcNvN+bVJqI95QbqPf5MX+iK
WNPQcF2VFkg/DMYgqanadfU93lHIDH0GPysMEhSAxz00+2kdkni5mqYAkcSNw8vY
gIYh0XI6Z0UCnsOKI2w2Ms2a+jC59GiqhMK50nDnzHpyz+1lSRjE0/Oqb5O26YcN
4w6m/U8ZtLKAcNCvQQzZBGzwaje4AhiEIDEoLVrzApeocfI9JBrqHvTkBC9S0Fk+
1yIwi1v3HfO6wcbs0SeGS9DgwtoP3/Okm+e2d885RiF4J89jMyZuYpXB5L5zZNu2
N2n3JDYqAUm+A5J/S3jwTSUqh2gNP38Wwb7CkEXp3B+TWgbuPGo2tjLmZshk/VYR
XuZG39sHvuLPbzL4rg4LnurmI7Z9jtOdOb/b+C/tGxWez9SpreO4RVbprcg1ujyo
9cxoDP7pPdoOi2uQQxOVnoWIYkjO4Nu34TITrEQpPd4CZv8PYHSHFmr99FLriZO1
Mo1VPAW/sWpex8cNSlOVazqWiTyDbgGUU83j2qBChQ9sRXMbgxOWveR2Nc91jR0A
dXjMpQ2IyIWh177bhYH2mgyosK0xnwOydMcKoM42YBJN4v3ewjNUhd4w78tAeRLe
ciPWdrOk7FnfGsaIU+nKbmTzWuIMOAwMMp0L9lKUbJ1ajDGb6UjPe/4axEmFkh4o
XOILX5SGjcd77WQgSJe1souSpIyxFbkUc8HNtepKroYK5fOV0Ttum/FCOxeZbFi/
QUGl5Bvqlzto/oLvrzk/b1RuKtQc/Rwrc15qcusDUCcN/5R6O6TIVlq/jVaAM30K
BPvfywmL8SBJpT7Oh66ZTqoYkLeH9C1DNR5FLv+IfvY/gYiwdGRUcF6HaWLKKFqZ
9afRFlq6DnaYW91NBiZMsSJ/x0nkZQ9yxauMpILUCYhT383RjMzUgQZT3RvlxKVx
OXvTQj48aSs2aqVgY/ybVKJW5LgXEbyQIr2JSzDDbeoTgNCl+NjwXFwqE10yhOUh
vv1LW4dedWX7FubBYGDJV2ZyOmfgw5gH9uZ7ovuEiHby42CqmuQCALUhZeq39hIw
2mpvKw4zqohw4tUTO1Z+lE190FzJfFhY7TZL/FH4XoVwW1SRzqWycc9o6aqYJGg4
nglOjtiTRfOtj/TE7x5juEWt/oMHfPUngR0rswDnCEePxUnMC8H6252C1B41bT30
AXg9RqnvgamN9d8/t5c3yFfiXXcrMkvmNwXq1JV51oQucTrChNVp+XGZVTj1NOFz
J6h/jWdWFRCw9KO1IYDR+d/v3aBNrGfVjmrd3i+zwKioY+4eKpj0OToiFEN7JkFj
GNVAY3spuPshMb1VfNx9mauyQUW34oJeilgnqbB7HRVEw6TCt+NuamnZfnYIHb6A
+v/jfkqSv/EJusRg4UlN7klQTc8NA/FRUA+ZvQsxejxWtGj2y47tjzgvNQkCJCx5
mOT4KCTw7P5GSfY8zJsViMGaPXb7UGBLAP3txWUTZTzw6Iu7t4uFmB3otSkSwR7T
v/dA15rh/Mn6E2lQkVb1mTvmEdQEhTbhAHWfS70/7Y1DYAv91SGm4cNJsNrazNdc
QHxtjq6B28IAMm5ed5waWfz1re7z933JcFAXUEDiYmvAwkJP04EO2G7evinsQdYM
uMcotmlQjt2lDOh8C5T5OvE3gbBoYmtmlXwaZ97jfYddHT4DCZeFhImeyACnYLjL
6xSdLVaH2t+FLjE6Vv+lV9lICeLhGYnCKqHrJjuoULa7xusHley2BWZYo032L6hx
L5WTOyXl0NCaeWn1+gdf0BaxXGlitQJC5uFsMK1Vh+AUdb/JOpxRD7rlOSaJlviq
sKE6j0RudkNxXfEwj3ReOQyi3x2y43YxUXqhzpoZrU4D6XGjrZY3ZBZ748+OqvMP
z+VLBON691hbVRYpOG04/rcjgrmITgVm+dBl84x1n1h31jfEH1jFmVtAcZu0Q88w
2rcArbSzI+4vn4L1zHdvT7IixSiNY5IxwUpkqPPf4AIWySjEuLmXbqNqJFDhLpGC
8XmAbF076V07SVSUdstIiyl6QUPlR5JNkwsiFwEkx2DSjOmkrkz+x2bmMvWhyScN
I9p4HbG7eB009Wzywt7pxJxGP3K+Uy8pxsfYaTqj+j0+k2CSf+ipdWxaW6zk7N/c
UmL0fCxAFkLIJj6L4ZzkmLUI5rftj6cri82jQMvtOr7hGn0lOP839PcpufQ9VIZO
DHTrfjBnzZwrcP0iStCnDUAvy1hqaMmAP8rIoRlFMo1WcxdLoaJO6BipgNmqxSVT
ROhadMQ/gP5JRlTWR8F4UzhPK9UUQV+u7pkXzxbKse9nw72qiX+I6ExoXWzBivY7
44CggY9++lwts3+xIhxKDOs4QiKx4E0jE0z+BlkCEtv7hArH6xYYO/hENDwRPule
HA/G7QtXib9T8hDZD/rdZ0Su0MPE+denxZz3QiOvp8FHah2ySJZxHnCpi2ms8Jj4
BKuEqtBitsxmZsurHqVHDW0kSWizqP+2DcJ1ZISPs9QTO5BSBhABeSYd5xzAgn42
LV3U1b5kzbwKmVKRulFbE3p7wEFcOnSrejBV74IRIyu43b74XE9Yus5tY7Uuncpk
JlAsV94UmbS7vdMTidewv56sIV27D+UvOA4XKPuEs7sAoIqFgXg27QcLDtjLk1lN
uFD/YZ0+tLZMDJpbcqAgNqVsiolqnY04GNeJCccpLBMRtOOF5ys7Khq7apryDlx5
4/sCVcd1m6tRtVJXtl3s4MVBk8W71F6C0i7yBckNmrBpVjUXVIzPJdDD9twcR4B0
hNBa52ZUqGmH3qBJotCxn3zvhRcwXTspntbBb2URvzW1LMQF2SEcZyv+hO3mpjyF
Fk4iIHrEpfgq0RsbQePFNDWBrrn3gV54SF+Uk51YIsoGSdv1oRdtn3J8rOiqyluD
Ps0BS87GiG9AelvQKw2+1wLWzEVZe126LBztGbNFnFSgC69uLcwbfCnS6xRr1sxD
fo8ELEcC/rnFFi+3rXGpZet6KGQw26VnTS0IIKVkfkvr8sMFo/q74k6P8AmHCI/P
QEek8wmAkyN1L2Abr53cVjM6Huu6AOncbGudrLk0tQ4S/88pLTV1nv6K9i1Sseky
phdI6qyoIPuaqJXD2ZMiIiy0PZjsRBssOvfhlavuePdczb66NKeG9oVeeXRmzXhx
HXmYRm41zF1o9XongiiJfv/4DhMQb1UzS64OsgLexIUpekp5Ajs8iS5fxeqqG/VF
tdxmUI6EW5k4BMaWMvrGbjEe9bplD699WdLYwh/Tik4rfnWSwqrLQjJobcBFt+2d
b2EtERpbnWdjV/nwqEsd6LS/SkOyqDXdC8hjHSzFY5ysLivedoj791LtvlKYdUES
NdjBYJLaX9UjNbxddmIzmCNkMtvOI40GAY+Kf9EaZtjBQ1VR04hXEaynV5gVMJPZ
tLTuDlAarcZnkn5jHkbl2iy9Ss+w5/6BFAcmgvAa0nWj6RyuqU0+hMlw/juqjpAS
fs42Dyo1pv/b6GIwSXxnLjNFhOQi61ondN1pBZmnFCcSU6yoBO5g61FVJDbb/MFi
W6GH43YPwTCcWq0+6Eh+PpWkgAMZvjqyTBkFtMHHMDZCGzY6lL+S4pdrUNBfKyAO
ygLAcOnOoVfmURTkXo5ldbns3vm1ph85EMgTbQYCQgFvrw3vvPw05KyTSzRhta9k
HqKweKZeaw0szuZI5YuCtSFnym2jYOCKsn2Tef6se8eJ06CxrLNLlIykEQC+r920
qnkm4ZPCiyF2wpnXN7W4idtqWu54SwQ5MErqXb6he+g7Kv4vNhDKrDzsOHa5DDop
MGcikeyKRz9ncw/dLuGDVA/NDSSUKdd2oXFy4n/9oR9ztKNhyzhBCuJqX86sFgq4
30/quPb64rv+lQCh3jsFEYuTEEc0dorvt0dpnLGKtvpsRO/PbU+i1sBFbrWVCBjD
+1pMN3uoS+n9NiLyV1XZHh8te11xarYq9DE8zLwkZ98g2/cm7ysuMnpoc0LzmW6z
jZHPCMzfjVwg+d/ugjwf1WKrGYLsWfS0p7c/Z3MedjTkqhwx8f6woUNSd8uzdmga
AUARCq/xSBI4WMPlsJw+kIzY0ZKKMcXA7sW8lVqod1daM7/fZhSAIxKgljdM6izT
iPdC1ye5hlSitWUI/tQseyHM6x6WEpFJBk9GAEc4gC2DTWIipY3btLSBLSyMb0Ns
b5sMY0UXlCoVT60UUN1TP1Kmp/thr3fsYMpbW6FpTg+i9ycQZHAW6cExOrUZeuUu
Yxj+a3ZySy5N7osQD3RIJ3sU+DEOHw0hyZpANgfzbcJQUazUal6NOXE0C9qeCoI/
lHpVplhOeqEJcM5uR013BIzciAPMuXFF29xtFge0KQwBAQ0WZa6XTwco75CmJZyn
YSFQd93sL8CsYSxhYlJ+4EEPJnqg4GfY4R0ZLOym7ZjY8gKSR486jMX80L0c8WM0
PdClOuJfUkDSwmyj3VETLDmwX/E86JuQgP/nspqfBfXpj4RD4tjmdLJltt3XCwAx
AtOWquqL9Kv+hbzhzja03olixT4YPLZQMBn1AmzJAedbzTeWE29bBduWdCssJyKl
g95MnXfN1c9iu22a9txCwai/BEzDl8IbDLW3grN+mtOA+rTZepsfhbzficWwiD73
l78D7KJyK9+zIx6+51qzFnBSvVBNA7HCcTpyi6PvMXTKn2rEUFidlP+6qVldsElX
APOJP48MjhEI/wKdQVEmia8ufKMmfI56yTWWwqnSdoWknPUxkyE+VgPsTX51CpA2
ZPmcQO2RIKhCcFalmnDkZ4IvkV8d4Ga3LjTA/OQ2Bws3diEYDl89A9kt+HlU3E4v
6l9zpRBYl7kXEmcLMEc3s2KI23a/axzmevFB030G5aABxIYYBu+3Mbfj5vkg8HUg
OMraJJpBhtLhD+mBSrQPa1UA4NyuSh4et5nnF8hd3MoP0KvtyqtRyjBATti6bNrg
lLFZjiUU5J5seVmnaUmKdma6INN09MJcYzniqOC5FEWJbJAq8VHAKwkdr1c9gCPc
V7f4bDny6ni/jB8WOtcY61z9FbHQws4XO1tygbRtUifqX4Z0cydPH2kED0/W6aT6
XxHbpIuZRO8DjZ8eWJESGL8GXe9RGwK97NYob/Mk2f4abJEYdC4+pkTIshVJlPXr
Vqx1zjfNIWjYjZmFYq1H7L6pzVaiGBuKk8lO51/IuJELy7Vo7NuumEW+Z0VpG2oi
5r0JQG9Xtipr65ytWoJUSdILsXOKzoonpUR72crOfBE6hG6rrPgtxV0Qx0gGU1kf
ax4Sdo9JDnsLJvryAmlDYCl6oeiVLa0fX9uxE1DVGE6zIrVvTFs8dCFqgrayCU+v
pXP19TqcijjZSuXz60cKCM4FL8GKPt0DdCCLIVtn35m+zPU/RNmoJaCuzzZa0gDe
j7xaJl942kCBBAHmhkRAysxEYQpycHbzUHIiG9az7aar+knltRt10mT9chAH/Cfx
eTtqdi6tVXOCCnTVqF4dOkP3XRNRr9upl1lCp/yYmSE1qpni3F0eBwxt78BDndIK
OiPozLa1gtdn3ADtkpqO9K7ifb64HfJ8//mdVgNW+V5KuBwunbv4ilDAt7NiWG7C
QmEY8PXE7VTGgyihFNU6WNNJCuZBLQbQtgHIC9voC/n04XT1eaKdY5+AuIKCWFpq
2vGZHcDxM6iUxIiBZ0Ef55RRRNfuv1sOLZQ1zBCkc8332E6dnvDdepF88LPzwATV
RZtFBtgXF9lGOSKKqUbFo1kJP6T7nS8ycgLvE0yQ3aToYlMWFytDg0ULKG5iCtE+
qbmINyOonh/2dSbltQPEPUXTTjo8+KwejNHcCzo9W0ZCEGFt5T1Ji7+ahYKRqGe9
LRnRgxTZ6nqGimShA0borTQzUimK9pY9UTd9xt2wrvUOBNweSu/J8CYadUZ66XY+
QjAzUrMfVe665I2JStUHS49jqTYBp8+Gyq89vKtFpc7vUBEPUoKyMQAs+SuJI528
qCE/b91tcGMAntYfU+4ARxRvCBojsXS31E1RPfLq14Ba2ubOyO4OBRHKhy6A0sJe
pRY+Kg6BKuihNM5P6SZ5KboTAJ5X0LCtyDzWeUkVwvB/dwcnzx5aVKdqEZd8EazD
SBqi39gieFan67H7qWyhnxuhgcItkccLRaoFB1LgrK/QMfvsy5e8K68ms10Y0Jb0
EGpfJDZ9a68DZVuwDJivqxIQvb714rcY7LW5WlyxlkdYg38qDI+7MpBWKKxNvGh6
ffmmcsvzeQ2yILmDB5csU0Rw51nKoMihoMHOAgly9OuruLva1Mw3Yi19tjT0vuTN
2ICwIVt25+hNLMUi52ySKpITNJ5YH8d9S5wMVVh6fo0sF2sbOQ2xrWZxua5lcsd/
jXxvOf41VUWleYD8AV2vaB6GHlt2G69I9K6t/F0UfhHyp/DCC8KOcET9yBrsfoab
9yfpfy+ODWb1FoXE/LScR8pHwDYgMRQ5lMDMVjKkyTNCs5EGidqM2VE0Z/TSXZQW
TA0H4XyDey2PflWaJMu2yFnGYwlwJ6rZQFgY0Q4zRFOF0RaObiwu0tjFYfQ9Rswk
dSL6Bjn71e5qAlpyqu3SwkHVJMFyssB7eTJ9hjrALAeKNhFbtcEB511r/YKbrAcD
IBWSf959edf42ggcPnnQvTPRv3QfxeXwbJdCA9L8tBJ59f8Pnah3w+HUi2cKtCCO
7M9eOD0k5opmIHfLTWYDUIYLEzIDnORbUHetnFysPPycbqEW6bBPjgBNtWQSweeH
telFpxD9JS4FQqCIkaD0+HLo8VcMZd1hM7wOZyMhCMniHWWQfWLkkM0E2kNV6Wvh
qk6BYh55MaNWhGycl52Dw37ry2wBXO2SMOCyBG2ivV1Q8fTVEl+xBqZJY0PuX2Hw
1z6XlsaUtSTS45aUf8Nz1dqsC/c7RrJEBnI+flsVdftHqNE2xsQFABql6R2xEUBE
CqH3A5XA4e0R/BUeXlGcmp1H36iR4bo5Jv8kVZ1dmretjP6yfaCP1NUkFVEWLlNb
iZYqN3do55yNrdcyYySqk97AS4DsWN+OmpTgd6Bt06vI7ZfG4aCUMvlcdZlvLDq7
G24rrklZZKqMTWPNVeCx/KExNHwXKfBEE+1iIyb8ZsAxIx/P4oluDyhYrd8/ymLv
gCtahgPr72tLgaZePk2VDdI4q2sv2ro2zvxFkcsrnfQWHDoIjR97uxYQfusD/1HC
MZpcPMuxq4WCNkgTr9oJ4noG2ysBZhNtyqGn1APxeWkFoEpLNn7/ECQzex+wsnK1
qGoRjGDJFOZooD9WoegYJHU325Z1/rgV7u2P6puG7v3EJJIiFVXW4KgD4o/dnwVA
se5oMz7wqmCprdahih0xCN+Fx69c4sXTzG5l7daOb5k/jHOKHburw1Rp0BvGPyQR
QSQGU9FLnRNjXYKKoMK8WtLc74UKZKeBINL24jgxNLbxkHCKpe3QkGylbkX40NJj
gMeHbTaYRYOGjSpLQSCjDUshuXEwHefYqWpyVAOpxIabdWbXhAMoZ7WMUETEDjd6
YsynmfhJqxdGMpWx+5DYX68Qs+c1rniLjC3qdhx10gVs8cBdN/77//4uIrOCun9d
o97lJwE6WYj75lN7zlaTAY019NIJpfPVSWOc8MYELu5XMnoea6DqKZVeOZ96xe2z
a78EF7M/XAA1lQQHKTz7Rvu1nOuXIlFcWh7vAHjR6VtJYkuNJDQ74uV4g1UowAWX
lNlHlKdkq9PZXbAN7E49H273XBXXnEVC7mQvtsucNSJJWbZTj14TX7IOrUjHKVHK
souoqJmFTuwd9YJ5OiUzB9cuyUcPZ1Cc3g1JesDkqTbFv+oFnlowK+SfTCre8YB/
3ZsCXXBwpBJgI9WfnQAxurAdtT/pwwfvTXIh40DUka8IzgYWoNNOhKaRFQuK0Ik4
fPcdtu5i8cC8kQk6OpNTXpOEyOae7Zj+B+i4dJxdI+Cj1czdqnfAHsrbCOz70Fzo
F6yb0imr5j8mEStO0hWZc1KNbF2HddwljfW9WCb7a01Q1MtG1EAfTD98NUj67ThQ
0SyemrDIRrTON0u1a6crVdRt8pEgNYtNrUVuQDMCsAKwPWUveWwxmQxV4MgFfmcA
IT+pWzKE0AxUTIOYs7/wouuiHtr6ujE22FHHNxQwYcye3n2rNcYYGYmCy5gbnLOa
ns9QIGx770RwBGvPh1f5R9Y2OrXjjgLAdJ2HBxXqaAKW4QaIbMmqanYkAcPc1Rhr
EV0BkC4tXCrWAOw0VXSHYxsfDoIonZI68pVB9TIkjBzbJagvM3445e6Os/6mo47f
ziIIM3DbTjYOl5qGNpExazGpXZPOaa5QULt20XQ2Jkob8MmNpZo6v0UuZprBSpmE
3uAATFlLBAHhE9UL/EwJZhGNk5vlbPvVTd3G3vo7sDpynm4SQ7hMQBcilLYMCk+/
++pdvP7OokJGMxSfsDttWS6iyP2ZNOzyA9K56Y+SBBiM1tApoIC4GMXm0QUPLORd
4KEiJEcoVQgxBKEjw1zmV55+FfScVqS/kjl61bDaRwg/ngBSwnUyx8Fc7OpZVYMJ
An2ir4g8X+QfjN0t5dPtBsbpKTMMSEzrpVmLYEofe2g1PaydVjnt9d8Roohh4QsS
8Hb7BfUgFoPWZP1Z1TPRwgasNsCsbVD2LCHgLMG1nt3U/i2RNXD5xbMXwSf0XFOU
LXTIh3gruL/yXpA8Wk5DBodUsN1CA8rQdZsp09X9xUb0WxJ6alqD26fv3dRJT6Qh
+Z+NYPqsfHJdP4JRGQt2JZQEGBWU4PZ+6K/m7XmRmYp3Erwk8w928E0aT7xmg1NS
B+HQDzus7tjjL8qbX08iBSVSBE1nb/5450xQkM8z7636Q4h2xYEyxi/4i7j+yP5F
lLGyudNyAAIJ/14H1+A9Dl0C7nZnQhpQoRa47N0TBCO3iC5BWJ3IU25ZqmrL2Enx
gzvQcxSBqR8FoX+vyQa0psJp+2U1LifYHgNJWPZEmRIwLmnItGayo0czFMKpStvi
YbqbdT5wX+n+6TUxEVOVglR04yStCIrmY1O7JVtIVjMCsfgdU4b0fuUDRg2ieX8s
5qETaIWbDjYBLoHlA81bL8041BJq7CZEQsgLpe3KzWUddjIhdpWuM1M9MJCxmxx0
IahljFh+/R7ZRirycphpbTEV/Yp2XokplZPRWsWiXjbd6icb4blzqfXiLT+8U0z9
VrCTq+sbCpOjhGPtX4n6+xIdnUIZXLRKErvsXRnIvh0VeTF5HN5Uzop3LTpxfaVb
jcYqwp31b9dQiOCG1j5zWFkTaZo16dXxTwgSnTq8TuVWRRw3xQhySId//BZVt6hE
Ln/DulUiEESPytWbgUIF2uFekDGvigiDTHm+xYVA92bzymOSzZKTOAJ1wh/6uaq0
LwS9c95NU2+Gn9Stg3WtGOuEfPHP5gcCaJ/8Ztc/C0Tc1w7HGTjUjv7WrbEEMRoi
zYXHrdpUeJe58V04ePxYXklpwvjjgx+FJX/Ylrb1QvLNdpq74BgQ9m6NIIBPWaDq
/rplCRs1MdzouIJkezDzYxagkRCBeocWAPZjTnDTxOm8ZYhirjkE6KR6koSHFKJz
8NfF6TTWmQSvboD4T6xPdhiP8x44BnX0K4FwMXIluOwAJ851SwzeS+LiFXeC1c6T
4ErdSJJkkZGI3lOxxWqoTSzzj9z912qJe1utuCujyIMo9r0WN+y6vZTMy0KtMrLj
hUPCtrvMU7Ij04NhxrdrYB2msZP1REf1ZRb2O1fvJRB9cCOJxD2J3VpFz7JJfw5c
/u1avzlQrb5/DJ5oXt6259IESua887/tX2foAKdQ792/lVgTXmdSSG2dPdbOEGN+
jfQbVtpp8ipC4pP87bVBmtO9hsdK+ssvA0atdcX58rlhWdRaYWqBfMBayx65IK8Y
WD21S3LSNB0LCRvHsTYgCni9MqRyLQE8Nyo/4U0Wgn8QnS4ff/BMEeI6lcIEwEql
++KBD9kXQS74GbPDE/R+QQH3ofw2usNj1oTva46fydDyx8/wT86hopdG9t4fdi0p
U6jXXtAAFruVXVLbzrsUdmzLum4wKcVas2/akJ/q1l2i5U41iYWgddmD5AQZ4EkU
bdwsh9vc4D/Y3OXqy5Ic+kiQHBLHMqazJnAL4NVpCYZ/VrDV5vMtI6gav6/XcnRH
XPgNr9Sgi+zdMwVLcEjLsq6GuIfP0t8UK+vZe+3BZlwgyOyRYi+wTM+wGTPoGrXx
rn7jmgBRTAt3RSshb3Tl7rEks8WOvb/NlcUmomnz0CCoGxkwAZx454fF8T4x4mO5
o2hMkEyjNPp0GHfEVYdCCnR1xrgmz46RUDipWUzYsBzNVGaIMpQq7E84uySJqy/V
5Xs8GSa8MoMZs4qcv8EzW2uSoFNLjlSj+bCJAvvAXGELJ+/a02WgeojxBeS2koK5
o5dqtdr9OlMnNZHeurSYeWswLJ/l8ysaU+c0ZqPF0tRiLn43tk/Hws2BlbB0l70E
O/2MIZ+wT82MLCC9ZrkX0LYpMyxWE6OZz+0glUBBg136AlecvuRtyT6nWwyqnnRS
dgbaPSz147oqpu33UNhEC3kVJiO1WJMRi5DDhEpfZiJTZtI45nNDRyjAuU6jIN5B
HwxASh3LDlpEMF6hsDdvkJaHgUZ/ZGvHm63ow2iGUVdnh0Awokwkxmrto7i1InJ0
vcj/ICCJiQylodweS0Ww1PkVgCuyqHCSK37xNilBQal5SIlrMMlneoGeTywTMW2C
aDiTrGSpeuCwFOR/M+JIki9Sj5Uf9Uv3Bpw0BgPMheCgzte1Bx7Ut8HngG6x+nbC
8W2vGgOsMxp1Z7Q94B4iFszovQjOZLnH9fiT6FQoThv09sw0LZo1UIn7yROnRu0X
7uEXvV8YXFDkDN+PZKM6KIlWyPSyyZEKzpLmo/ATvX73DXLXHRF7we8/XIlo+Gu8
R170rZMZzaNgYlFejSdLdPCEOMeukuFNCSRGhRw0+Yi1asC5BDUqRzuuVqIGnn+I
b+g0RGYG0bTI+f4n2fIm8k6v/O5AG5yoqOrfRInNDlYGMOnIOYAVhEx6/SB8A6+T
lTLIa8QSWzGHw3fW01BIBMGYC0Gue7EXOxLsYkUeYVMneKVt6pHNRIZHx/wAovzb
O5JhwIYUXbF9XWU++WcsKmfV4Z807wAViadvU+M4vMTNRCChQYLESonHdq8iqXaW
tQDxDazrFbRSaK6Mm7S8SqBjnP1wlcoY/DTzRwHp1n/r/JYO70LaEsShXy901PXt
9kPah40acTast9Z0wEiz01UHxQ1mjMHn28CkrojSJxzQCvfu+c3g1gWiv7+CMpkE
01LOQUmvsu/Kr+Lm7JJ0jsPCqEtljrVelKERvSfC2OB1V9rQpUcErUQ/WPTL4Xej
F/wHq/eI8VV4ZXaAndKSOQvQNB/mTDwqwo5weAke3cZ5LN+rhm2/kjKBUsJvBpap
SVz9xIjFJZq21NZ7lb9czwW39yC5PA5B6V8rIBe+/nNne2dLqcnK7KkZb5XylP9I
U3Dv5yh8x97iTtH04m1ESeK/5q7ka0Z6tgAdqDRoShrzUbYqTdQduMzkEciiD4u4
XP1tUTwGMJcZlFckdB2R46GgHr2WHrbJ9+DNtNboxLzDTMk8thWBbv1Cvb0tL2db
X95ze3ErcYuuZDLQIDvP7OM95MDhkGwu49Eq7NNy/Cp3nExUOcc6VdAdIkJO1JoV
X3FDfmXI9eU+6ylAfAUi/8Vh4u7T1xnOgnJuteNSfWA7gHJiAi9Y8PRVI5rVyQ+Z
51u07eclBvk/lRXBp3noARgCw4p5Nz2v3bfvgz8LjAGf+EUpfSG8i4cfWT9Y3ZIQ
zMNPxF2vONIZqJJ7fpD7RK+gLkoaScg9KmD/9QaOnsPTX3a5kshPRvt9Gtue7Rd4
49WukG4AXX9VShHvKMaLMVuEr/ysiJURFa2iAgCTdtqJiOc4OoTm7JNmhOedP12B
Om88wqrSpwzgsSKPW+RINSVi8eT5TGKHkUHXWX3w7t24UPeQsAt9+r5A82zgwuDB
RahbPHbKUfxJMAUJ2hQu1hGAddtWF0iOUnifu+KzghmLgLNy4QiQy3YsbYwjbj8I
nPodlg3XxXhBDPf2Dvyk5zo8uREBquLtckka3VMe8R+bhZANitGHk1gZZZrGuTS1
NFRSdM7UgX0wRPFvemP0JTBcbkWuPya05MB/Btu7GvEhp7j+MILUp4aRTDkCYMxQ
QA3ynH9jN/FaGqPCgJqMFa4tTBgLL7NimvwNFXylv4ByMbeDGszu9TULJHXggWWM
WKOxRvmGWmM+di7wTIdUvUaij7MSJnKOSV4gGnyJA7fZrLLbcfcxnxTX1of8SXXg
CCRTRsGYbkQCsAIbhAc+oBq7qUl/Dligww1ynSzzqWSOzgGyrpRNzUehghTgAlGe
rFAkn6QnFGNmgLfkiWVAVKQY65pRRTvl/+2BecIrk001c2WDYkfhw98mZZoU/zBt
3vP23jE6ZTV3kZK7KdKorw3XzFRkmAAa/hfQDRKuxUtBuLVgF+cc1yPqkPtBMKj7
41uW/icQas6RPh0jYx59W5Dn/MDwVrwQC5bXSWEbHjl6TpXt3Mn/Z/DZJBnth3li
CbtYmmt5UjSFBzCGLHc196wvqc8CRQKvf9MRR70T1VLLQHvvRQb9jMG2uaN/5awe
j2WGPGpOEkmKjEWyTHzkiJXiJ72ruaInKPGvEO/8qnksC3jYyCLF5xCUT7v9N/v6
NSNs4lyUasj3YQALBzXM1cNCtBzuLB+sFLhAtjG2EJJZLzbhyzUODDt+/arlRgBa
00RU9xwHx3gsKsZhel4Sj7Ds4PyVvcwWvR2/6OAMSx8sITIqb4YZQgSRWYRHWtUH
o+wjPFQfCSaHIaM0fjPEsJzMPG/c90HtJIzyyzV6TJhdaU4EM3w/VHMFAHFhMThf
H9pjfOm0et40J54iMwMwEXAsnsi+4fa3zG7OPy9+T2ZLhuLPcekZPS5Z3E/AWjAM
opI0IQLKND43XrB6UBio0s8/JyqR1NEmx+Kti9hF+kVQrMa61rsa8tF/YhNkZufa
mOAHwcAoDLpnrUAyQHjTm2NW5Ej3tJQvIKgRzN3YIkWUJtwXPht2o2ApQWtIhVpU
ofozkkmdawF805rYDBIQ7JGEvmpxi5TaCto1AgDfvVY6iVySM2mPxQ2vL/MK1WfN
qwV7BWUTG3bDZdoRTh1KzqTwTHV3vXL1elgg8yxpLC/s+heNjkseKVe0Ld9zD0WJ
FI6b021gMsLU6dsFwH8bDBkND4QU7O5OOZ7yTjmd0d8LzV8QzSw1t1GUpibih7xw
U5SumzYY+hjBVOrjZ+qUe756z0M8otJStn0+TqzM2YV47emIjwHgAfsltFZf3WYH
ipAmWSjrp9wRcKJnpsnTvHWaUXnX4lMsSX8pd9uMV2t3byvBDclu1WJfonrczAK4
ZTlB+kSfErxzFnCpL68DEQV6bfLWtmxmfsJOVaruIfZn5ndY/nueocOHj9KgLraS
rdHpIw/eMix42Lu9grAxYBAlpzhzuKHGrbhy4DpR6DNsMb4ocpxleAgmKxLILxx7
6+ob0DQ48plwbalReEEh+nO8MRwJMLnUERmtxEN+kwdWyNNGqZgieDUOX3UiUjQn
M4rBV36wluXn5Sj/iqcqGLo+znM1mex2yGKUerm9S1o+OORjmLCQGtiP2ZoN1yn+
XGBhlkyAuSd8K0x754ADY2k6tD2jaa04HEieAeOF1QIwAgkgfT9pOacxrDtMmFnp
rcWyxr1d3Ho81RGII+vMzX4XN36tlTNVvzeJqM8srsy2+VZoeXrn9IMNdgEw1TbA
v4jwfSUpB7/YHAfyrc07HDyB4bOc6CgISyBqhUKp2I7pGjZkxl5KH0+RJcbddj3u
wxoROcvpixPd2eHhlJRkVKEMluwn3gyjap2npb3rlQ9bWE5jT3/nRXa4jLRWtILq
Bdm1BMPYm2Z8bc/LfoHDaEJ7Rp+zHgxRUshdLWCEhSlRHADO43Cm99V3RkGXz5FG
EBvspaz8vB2qSWBmSt5UPJ7gzBLrISh8DrkEMiWDkghZMs/gOy1uRkIIm8oTUw4r
M3JMJEdQ7qG7nzubfqwnp10IfzYYLYSF6FnbzGvJFUON3bLouKLV7lWXfQP5Ihnl
5uO662c5TfrTtVn+DX/RKZlikWcgjENN9EyZQEHHPwUI31DwU+7z+n8L4lNYM7dw
Kc1G2EqLZ+B+LCpTO1olzEgphJmlB3kUCErtV3QKzqpoNquEy8zxyFYp6rVE7qMk
Z0BHLR+uxFbTVOINCg/muAlKT33ggYzjqYDQUR9R/lwTUE/5ZMtXUV/jUDkUweB3
z/bROBg+MIB1LsMuEYAnhN8Ua3KFqI6pl7Dx6lfh8j1bdgIXSOeSLYBi7t2Wg8C7
vxcZYDXLM3ZhL6o9y2tDCbmEA1IJCtc7InDSfRFifnb3l/UjJd64wFiGgJzI6vRD
iIUgw9zeRWQ/fgYILx/A3XXNNWTFHeT8IIn6a1+2fwxl0BIElH90ma9mH8/GLSAF
v7AjQjoulvUZvMfZeNeI4nYgeCYAZm6diwNBROghOGtqjNB9xvWmYPyxxPhZ7MBx
4ZluSV+eQJS9SLv29mI22vsf9FDc24pG50hs5DjLtBQ8EUL5fhdBXTVwqgpZ/C8H
vvO3FAhiOXnEOzRotOTpEvMq6rPVUpMQmbqVD+V7pswzmzLIvgrqPxNGBILAbWaa
+tygBh+EBSz+gp7WZr6Rpt6dSnguA0OEySvHXtTNluVOV4yNecGdhVKAw0y2j0LT
8CwMW0qOnkUh04bo1MNBsIx0ZKYvjt++CdXNom3egPn/A6TmUyPbQp4kuMgDo2KG
460UMGOWaWDiqI2Jg/QK9sgw3Mx4parsWxt8eAeAqQ9xZG8zO+e4F9StoJJkXL+H
zuBBc9UpO2TNMaJba6pefBdZGJKw9VxDU82u0wNPC2J7PWAOEc8YS2l+nTcioDaZ
Wx6WNhvegiDbAvR/DR04ixEAMOQIvasiZ8NYWtrm7hlgPl6EKQJK6AHOb+rLQnfA
CmqW8jOUxtSWB6/DhdYHQrw0eS2o/ue+ZmpMSnnhsPDO9/qNnStTKY0hs8lGFA0r
q+BNxkdRhgbfuBISLlcJywSRtDa5hSbpvIbq8gjDGW88VuyRoY09mGMZbtjTctUn
r1+r9FFpufz8XHW38zqF2Bvk0h8ongCynF0XDpG+aPvNS27YKS2NRfVL8Enr8Ywq
rNKQ98RtyOH4Z5r2aOF4iDrmVKJorMJZqUuFgZjacbszf+HF0BxysoZPahT9/li6
F7AvHYb/qsCiAYEM4b6Otyyl70Ebxyrg3RNJliD3XxJ2ahPGVGgGkwu0ziQkgA0i
657OZ9VLeZxnvcEmPTZYhpQ2xlDK3FmhtmE5dcNQOnKRCgYCrMKYWIQY+ilwerkv
3TyLTKopbZ7DqEREtI1OhMIMQtabuWtR6RBvdy8w5C9nA2c4e83Exu9FCrtDRt3q
ACuJZxuLo7zMUNRsSCKr71YrlqWFVrISuDk7bCT7alDW6I1jQRhMwgnUkiEg4XQq
3s+8a25VtXFhBmwTPNzNkzktK7Cb/EMN0sIWImAuabGuYOCLxd6udHI8BqJK3crJ
Uc4GutQ+4ZEZGpr9EnsMyc78bRJJ7Pf1dMgHFdF/Qrh/sfvkC7M/3e6wMzWMFZil
/dE6a91D091DEBB2aTP/kfR1+UzBfKwKdro5+EhQcRTQTrFfukN7wYoUxsZ6tQFE
S4bv7LpOg8W2wCxJ/IyvSPcvzcUvuz0BKRsS2SDqAxh3tUpKpKhcjoyhUyx4V57S
fMAn4hProRagBpSp+mg36SDUimInDpeVoT9UHrh/40ykpRW8KNBgG4tJh8QuMJVG
RHIweYuXsme1NuVMOtl7z+y2wia73tp3uR1KTCPs8bJHfzM6TkG7KrOUDx1TG39U
PbpyCPG6GAsWwoJPOA71Zfq6CI1jhmjf7qrwFrLe5mRkGL2qMPNfbuMFfddBKtFO
xwvReo+6j//muDlU3hx/VA/KVSjV6nrFkW7TMtpoSo7f7r2fmI7tq2xou2kYQWmW
5LXQY+a899EVRCdyrVM79iFQ/VaepgbFttOUZynNy4Yo+zInfHZO0euxGb6CVRAF
/1veQUzS29klXcgrivUXtKG20L4I889Qlwb0AdPpJolsZgxqP5y23h2fC2MDY1l9
3W/OxnKZHgK6VLTIWEEQ8YZxYlgZypyTERe0ew9h5n0j/tQJKKfj1GIoCKGn/3c6
8B/Xtpo7E/pdnnpShHZQLROtZCVTUV7jLjSxZP5qYjpgvlt81+5WhEW+UlyrTBLf
cwXPQDaqncGS78Bih3smKAE1fgwy0Ai2ar/5h9G3zVp96w/80fEv2XQHSdhhPwCH
TWARlkfvG1o2w6TVU+o2QdJ4TWcR+UziM3TO4C26+LXZgeW0SITrviUvwmVlf7yb
o/KfGg6chA/CKK0NV59DOaIkA1G3AtQ3NN8qCTDbGhBX0Nixxs+BsZoYVNIXk/9s
60RuH5Sd7Tmb3Pa4Dc+8AUufsztsdVXiux6WKR9q4Nyl4b+yqIlrp61GXpJO/pLN
95qRe+iBNzMUrva2UPotsKnr2AKwfZ3JrecplCcETv2us2LhmVo27VEbJgWSh53e
GnYxf1KwB1cuQM1UB9nxRbgt5FhfJsLJHfu4W/cpSd4pM7fZnkPerxE8wfV285z7
kMyzUlhNYLW+AqOqmbt7gtMbMsDGPqJNyPbbgYoyzjvzD2XO/8QezTPn9rqSZESE
VZNGBqY9OpleYlsDTYil9Pn8EJBXRpFbrorryB9b5k2DpqhEfnPsUH04dMDZr5oT
tRwNP3PA+SG+EzJBjttf9tGGbbEOhFkBR/Yan2yT/Syk9X3ADfVMFaSAog7EEMxk
3eE27LAP5m3Bl1Q/+mrFPRXe9lu9UxGLZmgooq7Y+vZsge1Bpl5fqgNZaYcHBXsm
6fUVRS3B/Ae5gKnrNSwd05tsgO2C3+nPtCy5aK8sZJFlz88xCHrPaVqs6H1fjpgk
6LAKyeggDl5CnuSv+vxnNx1m2X9SHEycoVaNkmL5zKa2I7lJmHiinzpgJ9PQZEo7
XWDs+t9facCew4019W22MQWq0rbZhjryHQ26bfkF6RM/VSrKW0jK87hArFuR/H20
qYYIT8uGM2rIpUc+tYphYz09DW6ZPEFbORmuBRqAuG367WEPPID3F6bfNehc295h
Lw0X4XqYBM9pgVnVfuUeW1yLNF5uCj/CnEAcGXSYyP6UhGkaEHtn5bEP0UhidXHF
dGfpis8ACfPL80UeQ8EprvgRmKoFqmsbnPB96Q2PXtCKOR+a1WURi7o+02ypOaC5
X37oddOSFtxPLFxWNdtlt47MCPeYs6X3dMhrg+fZ2Bi5TgL4f8Kgyqqvnw+1wlYN
HOAbhUr4PlgcbxYNj4kzXR6KyWJyBpufH7tRXHhT8pG3yt2r061sAv1OUt7E8oje
W35dBjcNJXRtEjViO2rNMvfE3ij+Ib3qw8oy26eEC9ehUjDUV4paPyhVI3+m+JTC
DeRIqan/2Dz6TSwzVcN6l3cLgWNmyTw7xD0ve83xMPa8osjitl3ihm6pOhSGGUap
8Oj9vTm9DNAqwUivNQbnfbHzkZwmqqMDrdyxLiy+dwElCyVQVxAZ5gYIvB3oyNQC
0JcYOATYclayJmwmcTLJDcEiVGr0AD/YcvHO5Yu+Yt8vdfMK9Ns+uLA3PQRMa/DP
O6ErUgD7JyTj+9eyXJZmYYFEvZg8IsForRC2IfW0msyMMF/iAbAWPi6qHKmV4IJ/
H9J5Xb5/LcmzPHSs/dqRzT4O5UDMo9lKPlx0VJ0tTDxKaMgZJKLUlsgfvkCFnknw
rYLj8QK3sGpgWTjySwQ+GsNT1hvzXWPueEemDylfq+2Iff3JWI+hqSG/ZIXV59vc
kG08MabRmXvRnVsQtdyutkx5DAWwAgCUkf5SOEv6rZyefh6B+rv1f/6pCFfKn93l
GDTRfF2BGw4qMKDGxUmOTP/DLCVIU3TSnudFjJ03T0y3J0R74foz6Zg7WTrylP1F
cKPIySlxjkBAAeULLJoqVkABOwqzLLSgeWraVTLgpNFNbWBczJzD7kL+6DtMEiB/
Y9wzW47cQKiF8GD57RAfWeOY2DQAo3bOnLIjb8MYLoCApj9teF+Mjzm37CnkY5eh
Hh7iPmeOdgDlGpM7tbb20C+nSAp5wD99fx4gDcrSZxSnf56EzUfIkj6IWZ9ofomz
wkMuB680zXesKJJHOJvdKIqIlM9Zxgvm/lg/QHvzTt+KoUU7phT20BNYGXwrG3O7
xPdzK+DmcvS8G557/VDTUko3SSaKSi18/uwmF9/hyUpaI+6K53Kctdfv7Lh8lSir
rRX1gWoVgQ38rHROSizVeasuteMeAEelvBH4qNQfvfxkUOvoqrql1iOotS/DqTE2
4POYxrqP7XcHVbUdKP1K9TL3lNiEBE2h6k+F9CrBG0lBXQ4doWGoh/1K+L+33Tj3
zm+/764QsBwtDrr5YPZfRVK8JLhnEQbuV16qMCZDbrQ8MBRL+DhEiAfiO7R+MnFD
NRByut9ynfDqXXMR5Dpn1UzjW7m3Df74N1d0E7PaVYM8igCSRnHBxpb5rNsUyYwz
kKHwuH3HtIvOYaFGK0+vZH8AQr2UR6O5hUcEtrXOSi6JT+FoIKawePuwvpKL5rVi
S07p5rN/hlRZnIHadWejauC9GwtK3Qwd/ikrnQXxL1izAtMP7cGwIrI/5W0H0EGW
WLkHUFGC65w6tcYZDFH4OCT/3yfn5xGIWgE2fCamhBFZQ6EV17eVDkeg6Oyx/dHt
oFSx/t/wJyXr/NvQM5cT4qRsv8f2t5Mm7MBJnoiwjii3oHIKMPplI2PRkNQcXMzU
4DnTjTBWkvBm8H/5X9b1FhM7tw3oWNZZ0N+I6S5LKUfqP2EheFd8Q5tdG2MufBEb
9ih0tKli74WY/OJb4BhOLro13XzWGqLk5fNq0TK6cAcMwlwTsB3X/T77ki/Nv8FC
yluIcKdcp4MVVvHnnVH8sySaCdlRORUYWGg6fL84dKhYBngZ5bn5ARAqWOhiLI44
uJHIaQBqRzJtbfblPmXXaqNQgWxka/QTNVp7g6zRKYwHhMBxEhKUjKbscQEmKtc4
6aXctI8Dnt66VFBhTtGa+aqDZ+Y5jpHI/fKg1h+cQkXoS9Eas99l6hhWLyBvKBsV
iPzjf1tODuoA2MuYJgR3RoXeEDBimoYDLmseTZ/qnSVLF8kp6YTCKXdcafHHb16m
f0HrG+yd0So9E2pvmdEReK9SlP3vmIzrp/f1AXoS+ypHQmBqAoq+0H9XHhf5mr9N
71LgZX5QP3bGWKudzIjo5sN845M6DV9hLgGIwdoA8llXO0uNX4F9HbHH7SYPTSRA
R28+4TnNSWXU5ExfREBdBK6ron0LpqLG0IQrS+2kroUkYc3oQaN+qbDjMuDDsAkK
pq8UiEyeZahavZcCxoB5YvaK6KDcbOOFLdmxfH54C1eIoHBoVXhYkzj4Zqjufarp
lEXxY0fbzNEf6kRf+QCQZFNgk9PJJJTw+5IbY6BMYfIErgfsOtRPUuL5nLxlHka/
epLeNiQunyrx525oKMETGs7w9i6XFANdzZqSTogvM8M85uPDcZPLnTynNvtwUDQj
1FrAY6CD3ldSrE5NCfs9wXy1pmPBoo+6/ismVoK/gQnBwfr4vU1cLBYiqeO8l9u5
oWU2Xm9Y9/EvEzCtMMGE4Qr0VsW8Up9p7T3Zqc/46Hx2PeoenjjqPKZ3wvAau4h/
XxMlSg56N+fIPwKiyAaHW2mXug5U5d3hhFny7qvK6NGA7CvsHmImJ2G4Tj5kNtUD
qnaQ5KPwcTyXY2IQ11rnlQrPUvEmqL2JPCfkj+3WOsg1QWfCXEwHfZ7kQ934L3tK
rhwY7lKwTQPr+RFuQBmA0eTKNhYQgyaZy+H5hukKa0+0itSFgdiq6u9VAJvIT3NX
yZKSaA7w+oU0aIuJblOZP8yIXk9N6yWp541JKLqqIlR/GYlK/sKKA/NnxjktIrCN
Hj7Mc6lyqymGIrZYssekbRfFla6ChbkY6cqDivrDuqaCISWzz/N6MEYenY5WFdaZ
9X5+gCyIqDxSnfxihHIkBBlB0aiarEI40RYVfSOyl/ZVHTcM30s6GpcVRjRo4CqK
JqLP9JvkcFZw48KYxwCUxkQtOXzz13N/tPrFeHYjE0Pzl2ABUrSMr9/tzCjLmr97
ojOcSqHx1rQmet4fOA67Lm7ZJI/6vXculckmpDJkagFVVcGDgpnFu6HqX6MEEpLA
uqyk8SHLQWeUApNRnLkyqFGQQWysOI6RIvL5WxYG9wWQ0A8W0sUCrQknQiKUuC7i
K8mweNci0GNoHxdpn7ZBL5ziv1tVuRWkiI7p1N6OIGJSCA02y//iHywZ0DHnA8le
7mee5E+iup7Iz37lT853J8kv2SzrNkYM4QagMB0A+H8v+expxdMw9QEHMhmhVG0D
5f8WxdzSQFawvEGQmn++mNSj/JZcfC8pFCgBybYfZVBT4zekT9aFy7KrVqsbrFd2
TlkR4xh25CicDK6sYmDpDJCPI2tOds0PeCGmcSu3zzDUnDVLfoYG97TU329bUVAK
ChN+3V4RL6wU3u713GM2b7Tic+hrr2j9q1WkyDfo8XUQt15v7tY0vnCRoOlOEqAL
sA8AVMsNbibbwLsDtuZ9RLzT4VWhHjLCW2DU01cxtNcdfFhEOoL3WUob6tgcng47
6k0+Xv4fM39wa3non4ujOHC2RFauWkdUEGIBoCM7uL/KpUsxaoIqaLkHtw72QVpa
Z2rtG44YezeLjOCDCG035LdUDOaSGH7yDA0I2dhH+JnwJlMODyy3DkLSiGX5DowT
KRLxq0eVFylFI/EopUO4auaW0gY3jYAvjun8qUSxGuBipkLLEz8+qTzyO33eH6VN
NktrKxbsrCcWNogizcxzGm6LM753uS0kX0np9E7j7kPf+wlH4k34ny9niwxt9Qmt
ViWnE28Q9Ow2KfQ7rpv/XxIadopP7/YDAkv8xbypJF3Pmp3dCE7oLFYPfaToi13e
LcGm/VdcSJPkx1TmeQSS85pO/d6DZyhA84SlYBoFY87CZGWzH5TK7toZxp71vqEa
XKy0YEstAOcx7hAOylcSxvJUt2mJ5fK1tfZwhVYfBikyO4Civs+lSxo9pIIAoVQj
EZrwj1elMtyA1JZxCD3RlmiVFQ50i5Xx50cIOykaBVxPQHOi5qz9mqzJjvFw2J2X
GqJBgU+av+wuXoiZUwJpQDfMsQvBdIjbkN9RYLw8mGERgn8pK3/0Wk0r+dOfLFr5
38FNrXtalhwYHQVBJS6D/oPLRvgXbvh4FJL24muGoUjbm61sXsO89TZwzzdC2HJI
ylFPIuGTJX5QhblPJ/e0Xatn8h/GljTlbZllOwAQrEBcjR2gv1VzzMCkqt3tzm+9
Fp9oscaq6/2OoPSLEA6arlGTzDcBia85zbmhtGoAJ8bntrnBivb1ioX0mTmDiQVj
Aer2NgpTTIQelXfoYbvKyTfZ48PneS6zfZUx+HZaNIICWngZ5QWycxZHWAC8o/38
QSy/RCEFKGHpv8J2JbAJlBjnPqpNRIwKsyQ7iax1gstZdu2YEjzntJ1SM3uRzEsh
oxumS4zdbZr6VpKouQwl7y3MFzrehnOL2asMA3ttECeFEVBsIKfbS6TT7TsHsDz5
OER1mJFWUKdN14EmMvwqalj4osE8zY7ye4zcu2eVdkzx+OI+uSryARmFI37Fl8XD
frA+5IuW7ahloYFEW6KogvILPa+i0HIo8O5qHlwFCBeiEBFIAe3fZpdwKkIFsxJj
/9wIKePgezsWA/vyCN6EVGxSegVmHzJ3L0YQy9YFAaJzSKH1vo44Lw3GVijNxjy0
MDpJRFqQg/OQIZzj6ty/m3F34B+rRoqC7P9Ek0Mcd5bceaSZr5hu2RblpQCTZCQz
cgFBYqtNQBTzgzoTQJynkEiVEjNK6LclDkBiXK0mVDA1DRri+5SokOQc8epKAsvd
4ebGli0Pa8X/N0MynytjmjSV7lb1TgHxwOVTSXIdYZNNmGv+Ksbg6tW5l4Z54+LB
7u9JBX7t1PoQZ33K2jVhdcPtmlDx6upjHvGWmEiQ7sN6qEmQJCrrpWqQaNSlAD/F
657ftjvOnYjHO8T8cMfri0u9vZATMkdT+qYS84Qy/ddf2T7eGJOVa9lPQTn6ErFY
Wrzncf0mTAGT6BleAeE0EUgAbQnraYkVJiCqSbXytJVgUMsl3PrPw4YuDKKKPCQI
HJZdOVzm/Hv0YQK3VBBm7L5BjpnAi89+ZdSg8gRJHaAaxNmCXiJ1QG0PQ86yxL57
BBdNjdn5KBCzqpbX8YLguQwzjXCMFJiw+URzkm5jxf9UHLFaSCkhYcKuie6ELg3z
WlmHf3dYtmKyfHCx3Mp9cTkED4lufXcNGwnbS10lvSeHopTCa3ikGoeh46bJTnSi
N6aMHkIvDv7ZQeayLRZq01tsU9K4n/yWnGg+bTOKojtlJMM8k9OwKDjZZLylEucq
noDHYGtgSkwh4+PxfBjU49GSxg/y6rI1h1BeMmTF2B2E1rmUIjW7IjAsnJBHiw6Q
Z5bCOl3goNEt9MhN6wLlDIEdYkh6p30FkCC86icm49y1p4y8N8rn81zclLbP083R
25JKHvx3bqfjlvgbYvYFuJ8mlX6Zzut53w0+da9BDlT8uxbzp7uI39PHZix6zVO4
H2r9/FUy/+9o8K1bOAbsaE3Cz9cWjpUSx1X513TYFUr/Ju1U4csnAqfF9ZSUQG+J
912PExNHUZRzBCLhQW5va7RDL+ppklQxxsE+KTYRs3l7AgMpgnKOgSmOrUApO6H5
M8005JlxlH9hAKl4/1xx6V1+/Mspiu2A+7QF3IJxYOdJO6sejdXTIgBH6FXFAHu2
IYiL+3HoyecW9zWu+Xqv+8B6mMp4/thwYgu3L7HnXlUo2uoku1U5JSrkEBc5JuAV
5hHLo4x9hB+tRBi/aRTzODUCmHIx3VMyeoXGFQT/Zb2p3B3U+zAt5nFoTtf7id5D
YYM0LYDoV1ODrj7H/IS8cGY82ub0ngCWQsQ5cu9U0DVqMlaN//AYCfrf4idbKB7H
ajS48Pl0RyyHv+Qxh8svhViNRAbjNCbqWMtdDAPTlJWqiqtua5Wz2A2ZtC6Rwwyk
NWqGKkzq42BJtvFA9XGh4aXfuvwNcamyTp0FbW9QY8SR+70iI+t2PgLaUbyxpGui
JW/PKUa71BLJlxdF2lEmmO1SMoTbl7AuxuQq0UAYYd00ugjDRiOmdRZAuTgArtYz
Y8ilJ1QobDdR+ZkFEB4YjEzyTassSvxc/m5ZPCic4v7micvAeyDr/LAvwGR5Cqlb
iU50pdT8cyo/pF3y+bXi4W+i4uzII7OdesEAYT2pxOpS/GBPGy6T1cwX+BgRBlvR
HookOJyNsGzROKvgmYKJ2DMWmM2fHcZ8y5flQ35kPJVguL07vFVWFyBSQ+smzw1L
YaL8clM5UroyyDV+Mm30vcuRkpICKTP7IUYCd5EMSdf5L3tAOlLsdjesmhKf+mJf
9LOL62BPNXJFQvJVmmKmekmPH9EL75Eo1Z20irIYQOytKKy5+L1Q9RO/dLeb7SqH
4ahXl7qNZbXeyV6myLpMrBJRatFT7kgjoG7VHpKpdt39BCsrcdG19CIZER5/6wZ0
rJpxfSfQLVNJVV6CycXpW4DZqNsuJmjV6VpAqMtt7GgNDEtjhYcR7tDpyMVXcaJy
UlzLZJtC84Dp6QoTgUoSRvI2zjLU2GNGgDtRmYybvea8I1VakgeoTUvd25b8hPa+
FyoHWbcRcDD1sWpdobub8CnCucezcB0JJUtwaDNAVqds+ySa2ouRfwwAFQESky2g
RLTXr+JQmkF7hjX10TABLkUGdiua8VtInz5A7zEdR88mqAhQvdVnA1QqSi2tTWar
pNnU4kGlrKM+0dFi0IvXD/c5GSirTyQvhO5JHcVc5MFNPoP6C9J8C6ax6N+T+oBv
E4+OSEqQ3RveyOzW4dsgFFXFj29EKaGXdCw2wzHf40/rqbUxpj5K2o4vwlCQYox6
dRwThKx4qRgj3YC95mNH08+RjiJbqTYUC/COzMa3QNv8r+1XrW9QG7bwlniRvaoD
V2oZbWUS3WnxZS2awuVZig6CpU2Zv6tDQu32XPHRa4NUyhxhnyoqBJXZwP8asEIM
4IUBhEMWy2eyy4hCpajQV5Tuy81xpo8tbdqGe8wJEq3MlaputgIBqfWg6cuktVe2
O0w6NKh1044fqOO3ALQwbLy+ZIo34yemgYWgLPf7cxkEFmf9aXT6TlxcbQwKb5dD
CTZeD5TbwPYh71J326Xd5ZXSVt16IGcPec7lPn+bPt1vV2HioTAIClTppI1PxrxF
OdNN39oj1lTEdC2uABvqD3r6av2tkOOuHdGnf7MUSmQfv300e6KiDUcLG7SIMYSs
3tml06ITNgeTBMhhgQfRPfe42hf2DlomSmA/93AI6PaoIZMuHvsh3j0fltQGDDbL
7t/3ZqpMo88v/HmtCDSrIhBGLigu561Nud6ALOndcjh+VW/Paui/OOG4kLnoZVkN
bOcTfqe95GPjAPEbH+ELUAksrTmwE1wW4yNKFH3B9fh5utaZxk+QdnZvrJtFbtaV
3nhBZqpOgTPA5CLpup4cfVzjz0O5n73gm67DdPT5v7LlqUClNFkA/+R4NQvLZMu3
f6GW4vKZhdQZozwvf1h37q7vkV6TKP/Ny4wBbSbbZMdiOFxP2hiHD8IR9h2SuA/D
fK6/0z6hdIUCG7v9Xo2m174gvDxbNzkbkt/GsMyXJTs75PMpXw75lErMIm4CUCKk
/WzVanPutclOChLdRJZoKKG4nIMqUFTyzUATEeSd+K4e7VZo59w1bmrM4nVL65cB
zMyIGHblVAkJ2MrO8hxUOywu9zqvm7KAaBlhXSYthmGpAtJS3J4YvGVJzuQV1+yJ
JmXVN1FK5XJTEFvDrLmolXhoX+kn/uUXs1c6XJYNvmGS8+McC36ZWkDgXpDG3Pbl
qBAS5kiqn5+U16zk/T/E67RtTakL+i6KjhZv4JHpMHRYHaqGHOxeS87Tas5WUmQf
bDoPs+03rwXwnE7xB4E0Yli0FWLrWn7GlfPvJyhx34B+Uf6f+3Kq2J0EuLargeP6
76Gq0CfK0VRidlYqQovT+MwiJSmijgqetvacOfk+Xzlkiz9mfQytiUtK/T3yy4EY
tSEVSLq2gBiYO/1/AnnEHj4Bz4y0TahHP/6Jq/SGBHKz94c/0bLVRU361n6cDquc
wrNP8enMSeb4naV+d2a80EI5vGSOrV5Vg7/Hj8VjU++5OUmDJ3y+ubbnlEuTUhsq
X6k7OSFgwfN2UNigSgcn/P64sYwlnipsmwoQzKIsMC7GnokWWCYi4CNRsC1Tsme8
xokKG5Ri43OkWTsoEoeyn9Jkk1tV3Gam84t6raBVyK6EU+PMj4iKqUKmC6xr7aSq
2ruGzUNAjc4E3naQjZY2fVT9FCVqUPoiQDlRdW7HoZF+W0zSt2U4GnZFKeVhOuFx
l6xc3ejkPMkAe1PGdCv3sTCQ2d2HPFEM4/0axUX16MksPK5bJWpzmyGnDlcj3jwM
/WP4qxw3ie+6O0Dpd4Qlv31M45sYk5Bj/e5npUKcyvE3u4ZWg6I/FbZgj7vm0nPT
T2gg7UrrH/dyEOl42oUxzcP4b1jMlHvXmabABwwcIIPC7+GONdvcZDTgOv5F8Q3L
WXbYbkpDLsK4laDur3Tk7PLCzqrB9Gkqo0QNNy4+HewBLa8l2zKdlTiIru4oohKQ
r4FmeAWkkS04joQkO9lrt5pH+2130HL20a1jzXV77dsE4nWF2ATrIIiMxx1szWWQ
iym0lZEfb8hW82u9iZN+tzVxexVOmLxr0GNVh2pVUp7YnSLHnIELxhjc/2MUytsO
wE8gIykqRmX7z7PWsKrBxi03cbFecRWfsWT9S7Qc81OcPnElChAny3DOWvE95JOl
F0DAL+lSY6S3SRfwMOs3K9TL5+6rcmvKby+GzCqPhDS078opyuoV3VsQ+WNew1eB
OFsQ0hfImKzRV5RHUovNdOMrFY0EuX1fJiUMI1SzESCwLlmKQ5odvOG1dTIvES83
kWFR2MNIHIPNFa9meRJ7fegXua4BfsZaZMuxeWJrvFP5NSEQlfDxgcxj/4lNWNkj
4MF3iISCvKp/uMXNNX3zh+bLz0EsVs5mKbBIrhuJxPLSqnVwN5mGBDQNuhmF6lky
EwymqoMz0o94oNQkpj9c1HAWsiS9CZgVqR3CtmdNc2m4QdRwg7K7syhHmNATNxMR
CBLjtsGMBIsQ/tsTyX2I0uYLyhrJpAcZUeGgztvb3Cf3W6i37gTTpYm2kxfWPp1k
n/Ur2xEIP7P9bKndjBwpHFLRK5vDlBCgL2Isi9YdJF6NiSCkV7yVnpalUD91w9yj
Je2FTkphjHZ3H08dLS1bFsq2riwz9zLEOwUy+G5Z29ClLz3mDH3YvFbd7NWYm0wh
xb3LPx6owXVx6J80czjuN6vjfD4F03Nvw6oH6EFLSTAYlkdA0XHomb+ABNcQdEOa
vaG7mMW6uQ0lP3RnqILcRLycXCVdmcEgM2XMlO1ibi7+6YY8Mquag72MG2hVcn0a
cCWYn9TSA4yLaVVPaM9+LXBCidplfpZpDmhyIAlONyE2sXNoNhk1BLUrmOZ7xJAU
CnsB2eqEd/dflEhR73hhoJJ4OQssGtYIim9x9FZYagvWOBsY44lr3zd2u8HdcxH3
vfZWDg8zQpZhV3SLG162hqmnjQXAqzO5jKUL0fT00skrmJD7l1LwTXPW58qGhvK5
xaXtvjI5WJ6//wAG/ZTGlzKlMmKOw8ILQT787rSibVmLALybNG0hHTbP7qzSL/vP
Rzlhl+hbAZJUDJYsdvlDBH2bgBUtlJUVQYcCw0Dlqg5PBC6CVIrEX3X3+aqP0gBH
UGR5J6864QrHL55UVQiFdTxYya4JSQ98wUjP2fON7TxlCQDw94m6uOUqrG3pblMR
xWXvTsiXgAdhsJXSZK40ZHSfmJ+kGpjtanLU6SskRNBamRN4+FR2RaSiF1cxlrHf
gscZk4/KYBaVZ8G1DEVSeJYhuRa3OsnXRR5VCma1wkVI22/QUFHeLpivD9OsnIQK
LD1F3N2HpAWJhTes9xfTCEMufDE6DpLM2yrLVHMij53sx6q0dKcqWAEmpwUATlAr
zREbs+/va/e70sfRq5RcvSk5bJa4vFuSdm8oTySF7tb6Upry72PW2sBEOsOGAF1r
C/O9oh58WRrS8AfdAauh7wnfhc6eM7Bv6P8/jAbX/M5ffPX400fgAhCacIxtldXh
0AJYlb+jnSfrylZjQPTKz3Q3DGkRhjuaJ1AT2cKapk2cUyv8k2tgAEudaNODIUNC
N0uOp+hCOSx91NFL2yTv7G5J0Y4aMLUd5BhhDt41SU1/A7eJ9wJaLb9LyM3ipoAu
zMkJAgQNJbEyqLyHzA/thr3fw5Kd4qKjdtporkoNMZVz16/4tAGbpEUPXktiSCt7
qXMTLD1kUlwAqCN8aO/aPDBmkzp6yd4onBmqJzKjRSI3IMsQxRUlb+c6WjiDp+G2
2N2Sng32ZW9sAaGhI5+40QSwHFbJNJcFPNZIV0ZKG+32qh4AJZgpepUNgJ6krTPy
njiK+nFxIzN/BNIysmvgmGvXq/U42CG0baBKv6OpcNFqatKF4RNP1IzoUV5CpluD
2o1WB232lE+9ygvquNvtgPE/C+ZjCX/Zfb1oXi1tFBe1A6RoMhjwMHGDBLvmQGMJ
2rIQGtW7o4f5fPnaAeNPtRgMNzPhBhrCQzpNCss5WV4INcFCfnjXKlHovFTNszD7
2TUu/jfYNBlooRK9Z80uohzr3zRphkCKSZVRTyjo2t2qb19/hN/rUjj/OWkXKRQo
d3HSz2oV2sD7IPLhmsjSoujSAuRNjB6Mg0o3klUORkQKgAvVGpU8kxBMzMOl0zux
POEkr+iC7y0/KcNYhY9jf40OTWrLYeGIAO3qTvVjAjqGVb5VTtBDp6PKxB0/f1qR
xmxX2hYvHt60e8coDPliZwoQUjZvncSElWVkC9xbHInohCAx2e0fnvwYw5ikRA3f
6G1IxiJvKKamgyOx2i0ge5+6TKSMQ9q35/j2Vy9fVWIIkUCDVCfX571P2cI12vJO
a0n9VhuSRhJ8TlZ4uZcIv0raidnRv5jL8HZgjc+4gfk4R3Tnfh0uQXaHPIGzGn12
JBvOrY4YTah75drXKBhcukmQdueDvJWDqxuLRUuMdpXG7naYnTwlib5mD0XrH3z2
z4QYsrZUPSa+mjN81oZrBJKI8HSlqVo57zHjux2h6ELjd58jdNKAVg+ilMAi5mMN
mVBUdlzuWVIVhuUfCVf/wXA87JdoXP29Dxn1UBoKV1f9xk0SxaLfoBOpm6KCQJD9
iZqrLQDXs8yiZfUTnkJfnMeIGhHtxtklpO20L2F63s49tVWhar6S4F5ThhqdhFwh
KJyzs+D9ccYWdrAsz4X2bcw8x9SKZQISv2sO5gNNTen1p+ReeYJEGSm4lCEoJK7Z
DtFwv8Na8cPo3Z2WiiIrbDi45u2V5GHGI5Co2XhXt08ZT37yKUrgmSeZTLqz7auj
FJ3Swf+DsvDn7yOjFHYTKWS/r0XAbUSY9O4Kh+BNn2AO9eN6LEYPQnFyvHUYLeCD
/2mAvq+uI3LGcL2FgZCzNB6qiq0/1RHpxkUKhkxx7ABRu3i/DuXW27M+aoICcERq
zhTvj8U9Sn/alQtw6gJLavvE6c0lr/xrrNjfs8G3NwI2B2Mw9VpcM7dze3/TlCDO
BsGkjLAiQM4f5qa1wBNWY7v0c9F6sqka7kVNYIZXUjUx5+iIMOvELJEoSPgx3uZe
/wroyshgaZPhJUVo0NiGvFcoEajU0F2HPl60G3ZSHleeGq8JxOcgPs+9Am4ka2aI
yufm7GYOKtQZYPNtz8NtjEybksClQEB/4GKPja9P2/ULdyR02Yxe3JP28TUqOs/a
k/WxJpv+veG5DfeueC8gn9T43tCSoJGk07vZQqXpdbKsyyAuAXahDFhKfLDpVlbI
VC6ywaCvYs5FhAbTik938BVDqSteaJAVJgOHAsg+UeT21niNwjlK3xqSEmo4HBbi
wo9cJ4B3XRFLjenr6cYpqswM/A71aba2Ir8nvS8OnUUSHc38insBG0zNQe4okPcK
qx4EdLGrtTufYysti0rbJ4TZHS9F5PMZf3JwW4KouyQ4CcvJ/DoU6k6Rlei1oVEk
fIZ7j6b7lghFZpkSH1q+0mNSTcjwnVFHhrHTNlQwcM0Eblu3CR3TIQEpK0bdOV2K
VSlxu1H/diJZBCUftFj3oNf/zV03vbhBZzQU1+4fK2RTURRFPLfG01jdI5PocFYU
gab7HmbCfbmKmGwbDmbxjXj0ZSVQZCGkkDD46+g99uBUcDTNIdAED4umC6uW4GSW
lOQEcDtCrADKTfJZAblG8KIUZPgS3252/uMdr10UwCV1sQHLaRawUvvI5avB2PHG
m+u/810WGJMKuaaHULj4nur9j6szcExKJIWKnxoyEG3PLbNWyjO25LAEVDEMdWrF
XGeblvjyrLd3OkMrZJKiYNbNN0B9w5L6cXlVihnX2TvJxnMBKfdqporkZo0x/CRn
6ldkpWwRnX7WSOtJCrrUllsxNlDVBpLO2r3Vow/uWXkJxJ+o7CwlwryaSWbd6frQ
HBmts/e4jdP+uwfF5x2+CXz1B+s9wedcXSpLhrus0JJadCX4is3Z7l9lP7yNSgi/
++NUXYCBVxQToxhQZGEUh/JWB/v8+nuObF8o0aIKCCRcxcF2EiNFqRiLsQt3pjRl
XYAnhWoYTykX1Xf81iNDeuj8cKCu7AWXlfdDzY9r1WRnAsdqpxg0foqzeGYhfgrg
5h0PD01QEDAQtqBTdquoRzacsy7hTWMAv8dkhnzAi95tdXtfUpeE1Gh+KkTwRqwh
d3ROmxHLef1POhGKpug1kwjFD14XAAvo5ryQbmHgZ/z2tRqSD2dGnPkbo4Jebjh/
psywqxBVaeDDGikscndJ+5l1YGBmUygEUWTKvPm+3mqQfSkT0PDnVhQs0Z1wt9B5
KoQQWZhSP8hPI1OeEVEDOApcw2F7rH4CsbDzlODqZSrbV2v7Cwzr483bz3Wli3fG
DRI7axv4h6jddr+1ukbOSlolsttpjP0QXfRSJMm9hyjt3mHVxPxlCZ7asAe1Ldcg
6ToYe0Qt+4uHk1X417ISWrtBbOtpt2H6U8FoiWOF6MlPYbDb0xVX6bBL0HldzL6S
MCE0OBEhw8ldhl1VwZLcb+aTELta/QWdLA4X8DsS7p2VgB9PMe/P2kHDAIWzpw3+
M0Mwh7tmQN60Iud1xdPYAaVgnMYTag+JX+tI8gF2VggLKY+Kx/1Cwm3biwat58Nm
bNaLxAMrxGsCGHvMmndnQSAeKekNXBjIEbvCk0XDjfxPRnxTqVA3sjmhIZ/VC9gc
aXhatcbH26TEB1BcQkaYgUKjrrMZXpcnhz8xNcl39Bd3jXqgl3FzRK7qrTz1z1Y2
lxeJq6UxmsX210FXFsn/gY7/ce5ChV9LRseRY7OiMZe5jGu0qw1bdHb91R0ThChx
lLdUE3DFjPlvlXUmWTvUSfyf5RVVf91b6y8RxGv8ZBzvmssqj7Nw7xHCnNZpT1bS
VVcagk1DKYoAZ6Mo7+Pe4y0NfbDNXmhGNBp/0SZDuXvANHcZe/vW0gBHX09bHHQo
5MPLf7hEXx83HBymquly4uaZQ9nRGNkjyVhj74BP77R7i+fSAHwB+b/zZ30oBpFJ
SzKNVG7cHimG/3y3pHpU9c5XPfJQgUBYwq0f4GOFhMwXUli9aN83KZrvRrznszAN
I8OEQYxs8Znp/fKx5hMjbQIA61G7urXVhtvV/uXHDKRN6pycrA4sZ1awml0KS69h
FqKtTgLLsiOj7cuGkis5AQBVYwRhvtFZAlHWitR9XhV4ziKlb78QuP62rYYL77ri
0D/6eNYhtCef9LZz7srr0CklxrzX5FDHrXo92Defj6FimAXle8YFInDam5btUZMx
V+Bs6eoPfe+OCQ1cvsgyygkxuSBD1AQuRbUpAIAgMuxShvaxF6SX2h2xTzL6xVKE
sMDiK8o+g42lauNFaQGLNpkq9NQcaUaskiVfeJ6d0nBu1SA0T4umqufpdoGPDj4a
NGlL6Ixpz1c7+o8v2mErxdCvDnSXaRdagqeiQutfPBmzmrWVe23spzj58UPzEHDX
Tm5pkDmn7xY6+KQ3/XvfJYBxtITj8IgMWnwNMedtASUFgwpjQtE71j+mAl+0BBOq
sJj2wIErou68qmX06EAbZat5lYDVHjBqOhAhtSeu7Ii4ygkcu8FKHKjXvwBwe/Ay
mzOlK7HO0CIdA735D92v/jr1OncnyATPUJzxEZe7rvNBHq+62vZ+MKgIjQvSlLpc
k+FkqNualc3sH8ICX66VnTuGI+NjHO249qrwUzLsx0TUPocS1JYYaGb6Nwg2zQwo
OZ045YxFlz9Evfx081+qmmPPWbbNs9KEJr/9DLEw1cSnib4NIJSeQIJCK0331Q9i
+x1hqMhzABuItkYVmJRY1n/Er3G4xMbNB0JrmYZO/pNsNvdvv0b+OltjpnnZNc10
ICCU1N09su5VJcR6b9gU3s8yBWiDgsUrkForsLFjVKQsDUPTqffJPNpNsVA5khyC
izvjz+/dGKIphzwJYji6HV29x96U8IdWZrH0lmLox9dDJzlfvm7suMWqgJfLHDvh
b4vbUWzg0TtBM3hdi0DaW68bWa/CdZy2ZwwD2n3nlnaWeq8Q57zCMc8mJptl99VZ
RtP1L+oEqkANjBRh2fxcwMhPXq1P5irZasB75m61uGAi75P0Jr+ORDQiLSYQKckE
1pircRjs1WRatZoMHGEDLwCd5b7F0vIXMV7ucGfJ8oSy5Oac5PYAABZaNDE5un+g
msLqO7y9lev4Czmm3GUv1MOrQStuJBv/iyaf21s7rxfaGUFPiS9YlisH88ocxtWd
qwc9vcjFEZRg3cHPOwwon2FDoUWRvtKxwDdkT5l/JfR59IW3uCDeEMpcw4w/1INH
fNPg0C/lQeydfMJLIgr8EoNRatX1IX/w+NVd+6WWaoRLwWse+ZPXE8dKNUVBWU+U
JT4+t3jUlvwfQPbMICnTOjwYyjYrE4SRoBUrwIRbOtQB4NkCTu18PjpweNAfG3II
wMN7s/WZDSX6vnK3Ffl0IbaV/8RsVUNQ6W2awfVWAIjY+IyegEmFxx6LEvvOHFQA
ooVLSHaNur7U2kC431FL8fa22Mr2dphMTu+tErXuKvNjcNj6cUe0VwMRNKktTGui
mw/1e17bewF7cM61imwNTeLjKFZf76P7vVtKuIhm0qviuByOZrIRv5zX5c2RQr6Q
BgnHsKTgrsKwrHuHswm2zP10axORCrgG0Av9crt6/QjdlFWeLwA8vzXp/olw40pQ
akMDbaRxWA8W7vLgYDRis90wwmaZbO9oWE8ut2c8FSpCDDFCkjMmEIWUnNrxOf8j
opI5fF3KAUiZ9oP7TXbL9HddpsbFIUqiR7R0Loag038g6YXnwuq2dsv+/RUveNhu
Viwi0uBWA7VGV3pS804QFJnMxFu8OSO3WDNNIj0iVLtV5v6ORLrHstY3+qxsRKEQ
bqj+/5/w6FDdF5H4sNN7NADgRTKGbivRe1XrxRp8Hlg/W2ENxBZICZ9AdCATWJSJ
93qVZMeE6RsExDRBFIoBA+x1KKj/AhCC2P8oTOo3JBakr4Tp4YcpoyKyBvlfPJpJ
41bORbb6xZB5iKkADU2n+Ut55mpnImhoOAgEkwNmC5Vzow2XLIuvs4wsm0HuYg62
H+YT+n+ad24xIjqKKToxwYtZbXKpbz4vpq7qpoQVd8fH2J+FQ928YqN+aXWrwe9W
3IAa8LQGh0ekeEc054sF8ARJ3BVN6AVtgx5x2hFDVeoRcxdI6voE7n+s259DkYXG
xEdGTGIgVhSGGjqrsuz2utllxKXiV6x1E5W9dThWfcQ4PNZUlXXz5TCmDx3lGevc
kh4H8f8KXTkyzDMCXCnnuiURMALVr+PlICPtB96dmhGmiNowjYmG2n6erb75pQc3
ylKnybwQEZF2FNp8LiJAqK4s4ntRnRBo2PCxskDQgTWvF1dLieguByeGUrlOXhlT
oYwSBaHjNS9qwrZESdKKQqhbKa/D/Jvi6G6o/WWr5OI8lGrkfXlenB0kqNkC35hg
4WQNShS2uomlWORWtfRseCopaejAipZxzAKqB8sDjKCdIsHAarOlwZM1kq32FNaf
8q7MGdRoOUTjqSiLDztyi69aFWA03+HKBL8HkLFvj4Yleui9MCQMkDejluw89z2W
/cK5VJ9Q+GbUFpQKdDSedIwHsEpgFSI4EX+7iGyirdQ+gzI1QmouiGsn8IKuUF+c
rbAoHbsHH0gU0Tb46afgjHAUfGHSN6+4iIHY4dKl90etsL8ohY3ZESvZ9pM790hW
qbSHvGAZjbGgNZAGaMuyaEc08N0R0IdjkQ8tYW6208nVWfXLVvUUphwzkt0C/5Ry
QfllLZw7zQcKS66kb1t72qQUBIC9Wkl42zEOIGRs92/KfspOf3a9vfpk2XGUHwf5
2Ojnk3ivm1awP01p9AesvVoq/kNYJztJKrtL4kUygN0rq2GR6WRClHb98Fy+F9o6
fHb3TCCmGRTn++A+MwyKOrIORuBEa1vUiZ2fR21NpxSNQJX1ZvDzV7jzVko0kUb4
sblZU56kBcVmGEdqdbSbhYbPQHPuiaRSoWQSCzjUGO+YNzpZpBFLnbO42SzYU0Fg
XWb9WboKvb+L/KhsuT2Ryi9TvijLGgx2Vjegf+XLzlxQu4H0gQ3kZOSqr019FjdU
gI8B6iCLMGHwAf28kJ7gl6xIeyCFYxXohgdB/Zq7BbcBgRhhDa9+3UGco03vBAV7
R5hv0/eI8wzLCBmJniqkcuW8Z4yw8Edwzfng09hsx7ys6Vr7k95h8bz85Qgow0f6
nPMEmmi64yJb6TI/zI6eBHLFiT5jujOcQI11mrpPhbqh/t9YDhgIC5Cq0zWxumzm
LtH7DB1OrAFQ2fydOCeRq2Teyxr02Rq9p5q4qzW+0dfvtxR2FjZQ1VPiMFdOqeIM
5DnHJADyn9n8WfkqpTWyHmtjuL/6y5dJO/LsZBwlKZAX+7thFWHSe05cvpwhUFGm
YQhRcs/iFlxEJOw1776tiXdUkVjjBY1kFIJBdvtJ2d6sIYjWlWD8KvnCoBAVCDKQ
+2P7uUIbeaDQiXPsId4EA8CpLyTNQQmh8TCimINjZWgxIvME1arX2SxNFTRWuS0l
coAKvKN+kuOwO9UoUQF6CVrFO+c/Fm4Srkuz+AYu/L0tcuOoQLhkToI6EXxIXqrG
xJznfyztx7WVBJI75Rye1RI5TJDkqjLEJubB4m0hUppnLKNzZ61enhItMqlDv3Vi
r2yGg1HnBysZbA/N81yCTjYg7PRjKk7g0VdVv0izJKagnL/QBaaZHtSoWR9UK+Ui
H3/cEdeavyAJu89tdxxbStQpufRhhgDEtiv+qIilnwTgmpeMInkDFwMZBBt65PEG
J1OWrOAjQoJf7s1DNk5zCBJILpa9UgICoJQSFbn8/zIGzXEFODTrwOodu4QiwP2+
MuiKlpfJSxQoNdZXmudR2s1HVuVu+hlOzki3t1GjA3o1pK3kXn2TqtUntoKREOGd
YWR0UnahpHYalDI/6pdUL2mF7rabJXGi8/Hv+6S03J52ikvOPeJZ1RGMm7H0trPR
MMzdn9QtFNTXxS3FFKt0fWN0rzA2/rP0j5Vl8AuQAoFPpHAyatY+OxNdX/Tn0NwM
5+QXOEoki3asN2GjplwcplUKsaHNW48Afg5zhaDQlZVteOWKFksWIZvvO/IWtrKa
XsrMsd4RrwLX9ZUsjSymduk0yIps10sD+DnMkygNINhu7Lg8Oyv5VHi2K8W7EmhO
eHH/yV7+rwSrsSJlJIS1aiNFHq0ZouhHDQrzX6aniwO/eC8uq8gCff5/2tD6nIRy
NBSNTemO1tFH1ZkeekfNZq5mcEzDR85egyaV+clTl5yyeyOpzJPx71hYU7Ndv03i
HF66irgcZZRReDhy720SDJDLA7kGIMSsOTAPubBaCv93fpf+fQT/5xs56vNqhrd0
t0ujJeI8TA62w869FL1UU+uekcyy1XyXbGQSFhaNxrMvT5RzQ+C0M86wGgS7z/5q
I0TaD2WkJF5II2zLTY1j+aqQpRYWz+0Prsn9TKXQv73ubchw1FCJ+i/5Mqy1MIV/
+UyxLjoLmAsglrf2W7pu49KGlewCjSrxW0Lywum4cpAKU25k/uRrYuHhmW+Tmh4q
lN2s6Ty5m+xWaJyqjt4BrCKg+c06KpGVe+QO5HoUFnTaW74oU6zWAWzKAFJ1uXJ9
1AdIAx3Q8b3TJTr9Fb1mZ/yD16MhpBHee9NO3L9jB9/QhszarQKXuzp64cZ/f0Y5
knXpirOeGL0kNUML5Va2l76DI6IO/Puo49o1DPjWeMGWaRUbPjEqszIQ0vurTxrB
E50ZAb0Yo0QditVsNEcb7U0tQHtJ9yjyTVPyJ/+7+D8c6q28J4gyXw57ioi5BsqQ
ZYCI3vfzSRixpxtxCzz+iMN6bG9HHfFVkghH4tIAcLe3dET2Z00tTJujmDKHqJPM
eHg5IiIdneXhphTAxeCfZ5Q3FXMjbIq38dJfswWGDZ6zSwlzOHa0fjGXVaLoVlRi
/9Oe9/UJZnnACBgoQpH/tccNFKtRwQFFy/2o+p7Hp0q9VEUzCVcpFaR65rYd07cX
kfEJw60c9Lj8u65SaWJb7rG3xDj+zrAOcKj4BP0Ovx7rYAmU8GXtH3HwE6fTDrEq
Io5yfDZWaOhnxpnvb1yQkOYJUA1Y5ACjVOmKRqrP3+Sz6NscX1jNoM3bCTbSq8vs
vmKxatrWETvVDfJC3BEW9gnECjo160gfadY0t0Qq142ti8eQTDWiYMYTDQ+mxZ3j
VHvnuxeU9p0nwxhp9EnUvp0P7smpwDMQwzaIK0B4ZS19RfmrZ2Z4F4XqpdFu7jLI
/h7iac/EdRzR0pRJqKFa8LX06n9TL2PIM7/ScZHkNwzffKScBBmCjDn8iVCP4IP4
nN9WzvxJabBmvjG+uY55sSsb4RPPiPkLzBJ4UI6NVkhSxSB8wljeKP6OIW6x7Js4
yaB8XrJaSU9yFLrV3fAuquJoFHSOyXvZrNpKdOjDP2u2JB33dev1ak8HWBgrAXzG
2yq9eXaZSD6T8jiPkoQjnapVVfbrHLz5a7gkrdvO62Ogy8Vssxc9d85z5iWM7X0T
xd4wfeabNQf6Cv4Ww9+IhuUAICjDI8ElxMw4xpOQrpfKz1I+JvyUkKG992BuZUNk
RdPuTZ/w4hYvT0FBGS3eVDN9/y2VJcZzV9A+9j1wwL5yDMcxwc41EItErr7MTQ6L
d3wamZiHROd8DM+U6Xw9OZqfI0XiRL3mdNJ61+quWDrTnXM23i0cb8gxqRxWpoGa
sva//xmc5hetV5SiMRRfSHyK1b4OVsycQ6aG0liN7gcJadRvZ2dfIP5LiklIrOo3
wKvAQwN3V+YzG0OxORURW0XRItYbvbxAuLn1qH6cpA6EWPSerpZZSt+Mk3K+bXff
CyEeiQmAu+XQ5r3pEkJzuKMwpc//lVucQqwuA7UK6JxS8MEA9OuuYhtWc9NGMloS
NGhJwtzA+uqBzvLlFTxW9HW7gzXKAXOEIKHztJ1yLFcTTkao6HnVELFr88boMwhb
KpEAtmO1NCFOdgOENroPJRU5HIuK5l1rcuwQIIOMak1Zpwy6Y4cwOhzULpG83/+t
FBSSZB/grlbnNdAEHLxJr7SPzV5t/v4wY0ESSgJMcmqWQCr/+6MP161H3o0hNGWX
3bZKt+b/UlLIAVg8d/R3AYO/KGa7jefeyIW1uaQiI+4Nwjd64mkBA5nTdcdhj48A
70KeyJO0HiYE6JtLOk74HikHnISiGWLUBCKE+gTl4r4n1SQvuf2SCbsT0DO4zevg
78AtNmPSE7zf1s6FLqpTGS+ZDo6rYAul65K7DOk6gCqBTb4+TC7OyKH1g4nesIPJ
ctUA0QhjQsMmw7+zBQkP/DvKMFfONLCgxUAC0C0uZPKAGEUYIrKHJNXLY4ofcmhM
81MNSd1vylWTgQ0/mXQpagYU19vBFYZEaSauy8Uw0iPElL/ovktDZO7n6mSKKM9S
qF+U0pGpBhZy+JrFj/RwMFeSPloeJLEN0C0ZC6s8Bq0EtWYYzxF7IutohShs9PKw
kS6ENH67qF0SP10mIIpNdYJVa45DjPG+cHvQ7GQ8xMlmuWkJZMq1mcfx8uV6r92Y
2XnGrgYcKJ5tKr2y0doJYGByCi2np1g2lCsHtdX+kL06R/eTfRwT5/jJLNkTMMFD
SwCbMvPT/l+kFOjGt2xGLxnBjtEa/clNf1JrYctBOGImVKQB1EWnGCSewf3hR3BA
w49R2gBxhlWc4cybc5bA7XgQ9swna5CMhfpSQCphCdJKh4edBcSuPZP6oEI0Vn+2
wPo/vjxVZooGscUvW6ex76xRSWDoXVjKVC6rFZJaKPD+SjLLjhMMrPehfhUbVe40
yppOLrjR1aVWtoxJh7otCjI250Owdnq6mT3YhDxArphU0j6AfFrZiaKpA2SL4THl
re1DJ26ScISnjSdlgrGxiqlCu4n6ZCuNWd5UX56MRX+A+yqjBrQRlSUsiTpiK1XH
6UvIjY96BQJlWIsDdGQHndeedZ4AC72ooG7MOYVtbM4SAwbwfnxddlHrUBbdTmKo
ThSe4j875HVfAFNHUg1p7+ENQeNsfcMtYV6sAU8CQ8ICXffFkkhdi/xoNtclvh1m
m6MDEPfL2tQ3Jaix6PLMQUcYsw88UOGLKWgcZET12xb1UXrzWisQ9I3n8RcBGmST
SmyycQ6yvGRGWch9e9tXJ8oEPzev6CZoPMIVlf07FcN87mgC0YEe6uTxYEk/lLcf
MYUI6NXWtp7WwWjmubCdLLrqdGUyJ4HXwXS51tKWTKMPB0gOgxAhR6Bj85YbPJxJ
0jLYt2xHXNsLbxIH4I2u631JHe1WlYZ6/40ODY10tXVFRL96eJG05gFf/PIkCdqr
5IVn2fQbl4VLVY3fOqwvJ4L7NyPB/4bbiA5xR9oP8uzCxoidGMYarmD+qJ/FcEaN
GYRB7gpRhm1LyGQgCTPlIWAcX8ZRNDOBej50F4dkJmq10pfRAwc1B6HFP5CkabW1
bRH6t25yeJNLsvBZ2KDWYBjnJNSfEX0/3Dv3pygyyo4rmqTwQIOdStvpOXvUxSIt
iVP9JPJ0mgNOKjllMLhrHF3ABsb+399zFvyezocu+RDbxeY+7xKrZGBzpZLRck2F
SGqFJEFwVhwRuWX0hPttaqoXUSB4K3vDHFsb9+5+qXAEbDdmKbuisgoSVHeLsrPY
P1Mc9/A4eEOQ8zGw4LhxpirSug6kAaG2U1QYTdpwhGPRgm5GiptpMnb+UiIndxFU
ZrE0fSWtVpOUInpn26EMhYu7sq81P190l2g8C/a0ybEHBPXxuXXrnpnA7jilKa/x
LbSPgmTxEGKiTf8mYOBFWZFT+VLLBpT3mMfEWgqSvkD1X53xB3rHq2++oZ8kPjbm
QZSiakTGMPtEtKhiNzwOb3QWsESsvYeg7yDgENzR0wr+dBlTMx/CgUK5SSLfaLPZ
1j0gbfRMXordbxOdjbV8+Wpgqg7aL0gau5PIeqHiWHbNc1vigXLZX/hiJ3Gmr98p
GEQPY6hrt0as5UNE/bTe6wHvx3qqEltLIZxYncp/cJeWykqXTFK4lVFmhzkzqyjq
iBS7yRvb6vuU8GXYLOf8KqIcfTKMHpuYxLcWCTkNM//DYfcgDgpLtuThfSFwNJWH
soqAmT5drlBxXFpv9tSiXbm1pkDNd8d+tcBBRLZd75KHk/RNrAy5kYCWEg6fe+qj
wqxuN8B6drxdHtCIQ5OzqCl/sra6ROXYUGCnbbmli5W9EQJgWyBOsF+097Tka8Qb
x6yPZM6lrloUqY0n3OY/NAEernptzG1JuLX/X9yeMHlYPr+6jJOjY1KcJEI7B5V0
Zg4Wb3VeoSPJHeIB9jhBu8QJKlTCaAZOFhn987pR4ZLJF22AO87fKljulUDxiArR
FiEnxEdr2Qs07NbbKoWXkI7JvAMElPgDJaWsEDiQqcVdaTFhev+TSq6uZtPsQRo2
0ihx0rAFnKlQ17kvwVGY2j2Yv4cLi9sdFTt0w+I4QlfMQX5eWyvAdxiI/nBR/edE
IEK5TnBEsjRQ4dGnyUKoGHOFbdcGNcIxq/Ex6rxhrTP2pZhPFcL0hMfCEok5FiZG
+Q4mNZkTFrfxfneeJo8qyd8U+DwxDMidoLflcmtgo+EPhFMk0MS85a4uKBxR2sv0
q+6Q6dmAU2qEHNbQ8kW5WGyGLeHofWA7Nt7zZuyvCQgvuKsM5w3bUJl9COHogld6
NkgziPoe/AhJ+WtUwH6YPUa2pWtatTqTplwIsvOrcygUO6swO+lO1AMNmhCbt8Gf
CMmjsgd5OMY/AXklBhRGmCwtseXpE084dEqOnCNd1vS1sdXBT4woWyaEMgWfpk+x
MzLYshd4z4jCJzVPjBgvWsSrsH7xkGR9d03hOA71cvhN9A5ymEBtSPd1Ime8Cn4v
pqs0+taBi9hiNI8HNxtWsYSzaLJV3AAcWuiwdsSZ0/Kv5aRnL5GtUQTsXvYmngyB
0zhcKcGJYvn53iOim/spqaTNWCeXSFdU1bAhCpwqgZMkuCwWGFBA658C3SodqKgk
HrW3TAnB+EIDh9aCXT1LD4vSCQwwwYsk45+m3n37tERP01dSCO1nhMim8r2YOQMQ
aHPFTbfBkzBE35UEFrXepf3NELU7trSiSLUMMs60vpx+v/+FAUF27GXqUqThhASr
GP6Y5E3LIVYlkBZ9uJycezRjFeK/HnM3MAD8vXtn/VV2cyZwrxeehzXKa7px2VnC
R8wWJZk5jfdVdEcIzKo04zI9dPf5zeijrTGCpIl/ORkPiWwCE7/PI/3YV7HY4M2U
ymbU4FR81LDxvT9HIPgpGqNmqIQ2tNA9qYqD/esM3wSZOGlKF9eRcxzzvXU9PEsy
X2TWD77N177s8lc2gwLncipue7KauPZA0iYlyQwgXeM3pjlu2xkgImsijDwNQNny
wNIiDTBt6H2p2dmckOHUOiV0A9noOCnSN2FDXcowcprdtvx66gP3L1rjiKsDIUmx
ojvBaldarqR6jb370M2DhpUDPXfCu0vScAdZZP/Op2ZxdhZpxgjdxTOt8oCCid9G
SZt6CqucBk41U5DVyrSRtibX9wtelKYchVeRp7SBMu6uoQHRIS/miz9WjnQmD5Ha
9pB1ZtNf6+kLi0nzAy7t/ZefPfBcGO5t9WOKysF/9k3mJFz0xRR3NRCecoSrRT/w
q33TTWVZYyt5gFkIZg12lrnj2VetarHtjDBHStwwbU5LSdYjwWylzNX17YQOJvgE
w8JSWpKwHpZO4BPyi+A01lCT8/sCUObIQU1562xVq6gR2EKNvZwSR8dHrwoeUwmP
TphOKWL9K1K9yzRgjIQhSaPEccCpIQiFPyM4/uX68q1dDxY2SBKU3Gvvum0fooEE
zLRYAL5NAJ/S15jegBowDJqRvnXno7vowrxKx8ZYFKNBrQsLJctRxVNCCmPw6gL/
ai1Qt1kFwwcPi1psTHjR7t/PLOmPWzqn1TCjvy5WiWHfgw9ee1LukSStJJE7GSyh
DO0qSqJQN4VLXrPnNTt8wsjceB5T2fKL+Ku/Mkg0w9Tq61ec81+Ad2pFOKL9QA05
JqJ0G5Q4/F0I/W5DJAgGL3tXCSidd+aoeFFjxo0vcijK52AVwcwBTEOd7rnx+CEE
zCwk123hPXnH6yN5iBc4tvIdhtZ3TXphfXe34JSZgFdQU4R+nNInJkAoSyaTtD5A
SuLMSco/n7B+615ijKuLopH0U7xuszO+rLiIuWNwzXImsiN6VICtUWJms2gAMdzB
cMGgRnU7+sxkxoet+HaryNIYpY9Qqn7dbq+7/vFRGjS+kV9Bdz+hWUmL10uAqa7m
S17d0warpjqFNoMmjzQ+UtpYik3iqCuckcJmsCWokbjc3ESjz2LThJvobHOCJerc
PWovo47D7MlLMkdA6tLBuPvRq0o9Bf6xxg5xSg8oEW9O9quWRWflLa1r86Nth3K3
Qli4bQ6ZsVSTYOV3Y9kJRAJPdvA3QzVsfiPOLOOLFnOoXAteaqFVhVlIQLe4hJxy
DWNKuRMvFeCULolaGcLozY7e2hLLRltTPu6y4myy0Kjd2hfvfHoLfhibU8+4GbZ8
c7CWFa1MN4AuFVzIMd9zOPCKW33uLpBZvGpemd3bKC7Yoo2E2/O39tTUd+cTXIIo
BFJ2ADIC+yaRAdrJczB8sHz5vW4KQgHZkUoS6ciim1m62k9WFS26+VlK9WmX4FMb
ZfrGxvEgCyskRu6imKht7NhGcAxlLvEQB883hIjymgfifjvOx3tEGaaJC3ozQ3qg
B1Kax1JmOy24y3agFOoj7hxE81Rpwzb3cPNMPOlvTSBCJne7fot++7OLI7GSDDtX
i5DYbmvUaqH9t+0fDf8VIInQPQbz3k/MHfQxmCjpzID74lf2ZBY0tZBlMRNkk4Yw
P1UbN7QXMEj6iwCX45F9zXg4Y9zTnQsfKAffWW31z6UPc1fwKSkr5RO/5s1sKltB
lqPQqHNKduJJ45ge/vNMHi2vEVa8haDc2SeAq6judwxcvTILPhQdWWjAW7u/7i40
PNkINu0AancbP0JJm1OsbHGN8VawZemCe/6aWKoXyivHps/n0wn4UMPsI5AGz8o9
bw72hu3y0zUZtSQ0FDna7UI6kbplQRkfy7XnlIf6iS3ZdfZFTEUYUxB/g5gc4cR4
E0RsGwxyBCAHSfriLPxC1DAZi7gXGQmBCPn1InhNWryugjLmgzHv8b9g4QgB790I
XOx5EmepigDiBUQgSb9znbtYWs+t/oZ/4fEbCDsU2s3/KSOqFRW8wsbHfAUm/brk
SViIAdbzQLAGPMtZF7h3nTHQcw5dbn3JzA4kNNDiaUlMKzffjyaa69gLTsWFndUD
snmoMnpHe76JQDERd++/zwAInhJ2XRvJwR0QU7/vqpz6aCMfQW7XClJHPOwOH1R9
tcYZG8AVYqt4/ABUW48czb+x4RiylSnZ2CVc9T9xmisZfozEAMKd1HNkggzfH2H2
qNT06xK/9qbah9nyaiKCtD1q53DjAF2lkJAbY+d8p9trrT7VxcIjHVOoxTK3fpHd
r1s4OVZbrthOM3X9eaWVl30NBVGhMu/at8RW8DTlz6F6q8Zu8oHZRWZLBOK0/OTc
2eCIgMmyQDrX5n1+w5nyIJBhirGuKusj1REffggEkAhuXGvJc/Zzby7jK0cbYGv0
LVHeAwf/lx/cHyn/ffqqNiA1DuoKATbCWb5QzjFR8W8+RaNJWUM/1VgaTaGPkB+6
oipmY07Z+CnxxVYffxaObPYcnWGszjaKT8rfjphtUYhgxJ6VCtlk5YC6eDOY+kkw
+yQ9dkwemRw1ltdLDYbzjBefluIjDZOp4mxKCiGn+AAZcu+BkP4RVTRkfnTScFZY
zz6F46N78/max02Z4VvQ+c/FpXv2ubx1S63WgPlXUdzdzDgZwlthcGt2O95ekHcM
4SGV1EB63/ILgGuXrcQoNEo7zT6xpGFtOuoU/A7/N8XpQMQFoMFrOaFQ4RpZK1ZT
UbCfrovkzccL67cFOVwNHvMImHxlgvhg8Q6eLvK7L9BaDov42SMcrXGirH9QuSMV
ESVFPCu1wA0E/qyLX/VSxLzsKbs1Lstpt2+5JMvfOXA0y1Hj8aQdM57xuowIxEX+
oM9EKzcZMsHOZuQ+1EKNzN9tfQvLocm15AVHGsRjKjIii6n6HRACsYOvBa8XChB8
by3pku6wZee6EcwP0BBiQUKq8Ok2+iRe30F5cowz45uP2vJbyXWOoCiAnLKWSWMW
DBVoVwBuM6/o9pz1XgnhJauM4/WOW/5zxx1g5nbmmbr2tkb9zayJipIce94zDwdT
N0Cq5yd3VLF58/TD4Qet2ZUppvV7TFiLwCu8PgY3yQavFPFfR3AhkmTTO8M3IWXe
Yu6XUXX7oyjsLk2dedffOWi9EZaW0v6uI7lFTPWU4irUhBvmNibfl0EKwrrb0pzB
dUptWAiX4po7uqQEJob3lRx37GEdaUGzCxnH19mBgcXaCGY/o/94EV2Z+LNpqq79
1JNPomCAp1NMRO+eZaY81iWGCKN3l+g8OuhaDbUwDzVSFBIxMGyXuA01k2DTDV39
Piad8TbggzdWcKzrYiJNFuacTv6ohKI7k+ciekHoIfgnoYYlPXlAqTBJDA+riMCu
F+kQDjWTisSNSQE4PxzE6Qc4G+Vn0FefuzqOWM8IpaRlgqssfVt8lv5hbht2X6P5
OLw3xit8S87+s3qSORTNuEx+UoZcZe7d++fpJnuWrb/dZZn99ZCYqOf+8Pit2Qd3
4PEzaiiPPPoiodC3AUY2RRdT5lg3HxFkp+rUpqZxdk1LsVoeV45FQzg1ZfF9ivKE
khM0yHHJ/GS8QOIEQr5fSKE7nKfLbha6iI30X0ioRthyaUO4V1AGi0aVhaP8UHBS
kbYcSL0zr2o0bLjgmKplRSf8TsRzFgaCQQxPFdihpeWUJ5sxVUVmlJ07PlUm+w5q
X6YB2ZKzzyF1V+sU08GGb3cRsqIua475g0zgbdSyt7SW0u1ULJ3slJJ897NHw/Vh
PwhDPNcjI+bSd1wlmId2RbbYQz/gqVlv3g+YAWFDC8X2AB4tyZus8r7hFs0/kL+Q
UYGgItoSE+HEdUJt0dDDTq6XIBgE24+1SnTyNqhKCHKMsVO5SuV/3vM5jNh2SVI5
DJxAgnB43XzdoxJKDdLn2oVZ+DTKpjHUDo7tZJYB092amSHNo6NMZFGCZxS7IQ2A
QQQ85hRxDcLFJg00qXa6YstoSbqzR2cwp51MaU1KNtTYUwLhqbh0PoygWGzilm/n
D+ZMLRXgOPSzjn6PNpfaSj4uhWbNjjWFAStZ2aMpy9WiHzTpC1OK43diW1Vv60Nb
cxBBMT2PjWiNi+knXff0HnpoZt7CQdddd3U/qrJ8xzhUIYcbbd48Fi3PWLYsB/sc
e5ZV0wfsOXq88HpNS54xGR3JTh0F3vyM5j5kkNh31UeIt9ezSc+FP7Q8s6hIzmuz
BUL/kAgS3XIYeoIHKO5BoeD4LXoQr4gsyWauUCpwQpbjbmTDwLW+0a3wcybmKysZ
NjX467e95N2LD7ItkQ1TaG1Z6BWR/MJYsmPPzJ1NGAQ9pvCfoRP10M3YLgon4tDn
NaD4ALSKGU3lWCtZGo5W3JoHMdZNb1hH0RkTFlZDUuSF/JIrqg1VLwrc/vPc+P4F
TCW7jaH9iQJepk4vXl8Dhu/kermM2D71eNl6LHVUqp5D+bu1n3RTp78HwANNsMMr
kDQtiRTSE7tcT1kFhNGzwxQbhXy/P5gxpZ5OgcCOKFhs6IBJ9eZTBHBE7bQ8qauF
luK3VjSCNlZ4oZM9dQedYqQOymaUMlfA1qV5QJJoYJ1yPj58zDNT7Lw54Rm0lun1
LJ4paIPge+6acNkdSeAmOLwZsP/pB/k5hkIy2oq454M+K+oV0Tv5AQS+HWfa1jlB
wuPb4t4Ttgk1HbnJjhG0gyYNc5lC7OTnwuCgML/sNECFGLQFrGUQRQZR4NcjPO+S
hHUHNB1IstdP/U8A2VL1a7I9o8lGeXLaQTVbUebgWxhQz5wDGsXH6R1mnVXOqH8M
Rbz1NMNzwK2LmB+kNmWmn6jCNTX1mA+q3wJBCElQAYp5Kw6fFAbKIv+1b7k6kugR
C3xx1RDvcIfKdIm7jB6ox7tTdaEAPLP3K+GlJDEplUJf7ZkE9wqyjDsclOdgbBKt
h5PK2RsAwXWphp03Ol+0frCml9x8bBHWQ1PC1RY7HLlNb/M9s74I0ZJNAAtW/nXw
0C4gPBmogLRHxMgmEin7YQS4G8ao865NqBQvimcMd2GA75qFMwxq1U3naG5CTc+z
wMieddvg33lRAbsm2IwyvppOBNMEf1c4A9nUaJBuHmI9wbEi/DAQM7dJrnO3FF0I
JkN4LLaXlzpthLpyL1i0yQ2ukJnypXUDteLRHpm2T8GRPh4oRMYb+/g8J/CCXUcK
+7aNQkxKPlWu5yEWO+L1bkr8Gle0tLTna0lSgjWzXuJej5/w0peXHnZGKI/HLm9Z
mB7PjAk1XA6PK1JAK7xpDA+c/3xQL/7JG/4upjo+8XsBFJDsXYhYSnviHUmZUkv9
VjelmQ67eMki354FWb7yxWgeCPIlpMmR9I8kcDjZks/Yyp9/NUTP59bJ+Rz210Fy
ptsSn4AJjwDTDu0PHa+NOYdR+ojEOx1FXEVF2XXdaDkvmZQh49Zm8efhVFPwJCVy
/L4DtHQ0pfoXKtxDiwSLde7bJKJ88y/ACdCELNYKnO/+0JgVa2uivCqC4Xi1Etsq
mVUiIrhqSbK2rmCVF0bcZ/HDk08ecuwbVA8Ne88BrhVHbCTntCxjQrRbvXJ6xU+T
LZS62pq1WawYIrl/or4g+vFnz8fHfngx4abCg9WRlKFrLfDCpeDUmG8OPf7qlhxL
CZdgjSM+shFsBugaLWpNEMW0kTgau6yM5ROm+fc3HIm3gTEeab0SZLkkRU7dcuSd
ye2hMuf+lljyVTuTKf7ldzBFRqB3vpD1uhAA4e1eoG+ORYkEgVjxUwkJFDA20IEQ
X20/qagga33IeKWvodPrfTZuEwAL4Tm05Yo/NzwCsKCsdbpkH2PiQYWQug2Bepb4
2biLH815kEcYd2v9TC+9DoQSCaivPbancxaC3PDuUlIHGoPWTDdzUH0IPxgphUeY
7RKSA9vkxMxLmrxs0NGBPQ0nywIvCu5QpC0ySFnd4IoXDtuanbxWT/33nF2H8/AG
4vs8agbmz3H7zuFVPstxx5LyMEPFjSNoVFSUVisqpN69ngWOwMN7NpHpYI3ys0ER
Gcctg4Sz4b81sc3F0QUkxamZoRhhjCdYFHdAFysWIuTArkpY5X0bRBmBl1y4WZZ7
xI6bWHa0nSbVKvVFqJXkngdjXaM26sR2e7wJ8N6vAXnUnZXHpGaZsLOETKTUnPzR
1R/qN0FXIfaDbV/Aqn4BNf6OWK6NYg1TxO9fteJZTEw/lOM82eoJ3gB3S+CR8V1X
Ie2bHoLaZKb9baGSqDASC+ScdXcMbpvAOiOtA+N/ZHZLQoHFwmDtH/yngXphfnQL
3rx/P9ht3/xP8sPB6xSiggz5m2igN/SoDp81wBfUW2jTfNzydZOydGeIXwLREb/H
+YgHsr2J676LrZ7aXwlsaqHCg7WocyySdhxZplhjxTZiwjpz37FSkfpBtw6Ihsjf
glUf1VgZSYbUl9spQkW8dL8bntQwzFXHIUrxc0VZe6K8CEC2HKUx6Qoj+CrigkfL
RZnJaZaXIYBBO8SXsRYrRYS0f3biGnOR+7IYlG57W6Z1gp2/K3UDAGKfiSjmZSrI
dkPxUqiBCCujuoDktOj+i3SxIsksPRsByw6gc/wFXrgbTU83HBg6o7h4GW7W1/dP
VT2Q7v3rs2F056sWqjKIXdubjET1EyJRStI4TAdNOlvw0FG9upKxCCgPY/+5Njaj
CMcsvAWu12N2qVZSWZplJFsluKo3pfVZ26n6sQ6sZqndf1a7EKRaDiHWM1/hoRkV
cqSYpVM8eo6x24kkbUEGbV2QGaUtPil3lCs2dEqYtXf/BrlEQ6Pd3yMherIV4q0B
hyLpkS26asv/DqG2mPhLUtqpndFeBNWRmSkQbc595p6J2nTpLZAdNHfLTtp6YuOh
aFpdi+/sMdB+5ak9zZoPYHAmdfwRURU5060coOritmDzkzT9iFGQPyuDhhoxMBqL
IIAiMxC35gMBhpq8grXf7vboeZplLowGWz8jmfLs5+1R7DU7va25aqrcfrzLIX3g
iZDgZQ9nzDdvq09fqYznEGEbIXzY6gg5gHAGI0Px3EOaDQaDiuu8CzRfnIhotc2v
VpCeLd4g9m8tDjJWBewuuCWEX7quzynxzieJIYgjkFeBrQvb916BE9TFBEL1fHup
nT0WMK+zKjIwPCrldA+KpwlJZLVbuNfaT3lVKPbkfbeyDSHhCOaU1zk+VGIhEKDS
hMI6snCGK66bobo7st8LPJwP7bsTac6G8mtkvMa+IrfVGp1i7lSYjDJLfY9FZgYj
LSNWr6DaYoNr3lqKaqbEIw8VE3kSwYyMtM6ZINl2JxFetKyzIfAnnOdugmYE2U2D
0PRkJCWa2exQR/9cdzohM93mJsFqdme5J6irEnKMCySddHMPVDuXXdhHmNJ1v1Kf
Z6XqNfw87bgHlQXQKFtHbHPn18wD+KH7DI0hMuVXvkccZ/YXJxzghlRAWvxNx8Wy
pu4qfPxIJWOvQ65qz8hA0PGRYOt1hVxfJEyzoWuz9EpN+y13l0jTICb+5SSsjqOd
IIlwnDRDVCFlyv0hgxE/qsJwt8O2DmoF70pUNRXn+Rk+sWuCvtXzvvYh+orvFE1q
noRaHzKxChQ9nd3ECvBbwynH7ddTFvO6aHjVfjqGwmHl9pi3hZorzqLyhJf57WNx
DIhdLrQYVfYD24/cEni21A8ggBlOsH6cngwajOIbxf8/+XuA18pq2/l2u/nESpcF
eBMxsiHc9VXPr4ab8M/uFx8ZUQDcW52knOMLb9HXj2zgB3+pyAf508rVFqYdLYyS
WLUGhqzpAvyzOTJk0IzofGRrLbBp1DLk4tsMMH99C+Qz6piCYY93qRb1xzjyNvMQ
3q0iUpVeCuof6hXZOxxvXP/cUSEfYUvr8ZiWjZ0ejQC9cEqxrxLBlUkV9I/5+Pve
6RNZCglgEHtywLAmqMJ8xZ4HXhX7hw820bS4K5ePm1S08qdBaDmpuRyy+Ff85sU1
izjMchIjzi5Jv9wjnT0hyJr+S9yTHs932jD60WcR/O1wfMg5T5K9P4m4TZLssIBM
B9YYVsvq08u1nV8Idd3xoJKaLUAezRJXiXmNEPfgIXAwf8Qn49l/VBo2z3MkVIwN
/7LRPqhg4qpM5kfRbGiVoi/XNMUW+nYuu8h2G7vAK0H2Hs2yEPZiMCR0/0j/81AH
nPF+/nMsNBpbqRx3dARyTDEJCeLYOmJ4p4lsSUvcHe+osG/OsrNHfvRdGStDux0C
IWFlHb8JSr2+kx2qJ96a9O8OoV9mm1S9JTblTykoRf16VHrz1UDl7QHk6Lh548+f
8eaJYGTY68kiL9wgT12baTvhWrDuzZQtVrXcMWJ/FlT4yOENskPFvUF1Pr2u6JmV
szdhupAQITM7ah69vLiifg7LeNV786US9ERQB38fOw+sj/Jr3Xf/iJ/65vwvlSCp
QVieOeBFxPnq0iXK4Rl5ZzV/voTjRNzKi84c3o/MIBVFpsRJ9YgU0fy5SHrS/rtz
oFBOyJ68J+mXsxFEeU4ec5HnM0iHHfe3U2hWvuUbp8/k0Nt540VSA9TQSkjxVKCV
zji5Lkw1ggTgbLDaRs+fIMICq4qBGOipX+JIrUDeM0IZyzmhKvtdWs+tk9GMyk9s
ukCAii2oKK2BNXV8/nfqaUrB2cObZ6LnqaF8Hum43ZV5tjhOpTvQPhh8broegpNx
b43I5pOT8elUbhv+ALVQYJcjCpqWM+nFDzZ03JjwFbyamtppPVmuAMABnxEWJXs6
sekpCLoTybQUS8g1ir6uuUBXnTWYuvIu6GyNKiI9q0Zjf6lsySmhXLvekqdtkwD8
lFgfeD8z8x1PhzWY3q42QbFoZuOCvMy47lGLT5v4H0L+RsTtJa+pYaCQxFYUfWCk
b4MLtVG2Cs+l41ZnFXtIFvJVJPZqfuyYsAZGSYMGy3cuPUSA40rvE5mqBvnXejWp
TNVUNgYHwhGnZUupg6K669Fvyznbq0xVabVNfjtosEs39xyy/VMcKKlj2dyjqHkp
ObVsa0sR5ymHDHQyZYnG4d7OKZHo1DxVZSfLPEoLrFkgkoT+slYP8b+OTCaroa8R
aKCxfE90jWz8sAw0Kih/KOqneJpZ1iX+tTLSB51k4w2L86ybQKDRz8pHxFv+XjBD
BNTY/+mtcxMteX+cndCWNmpnSBCBX31BOWfFLwxnINqsCMU3MELGrWzpp66Okjxo
WZOEGA9pUyjQ6T8ZbDX2cOYfpB6cjs/HXsI+VmGh5uUN0OFFL21qU0rp5IU48rgh
69q2xPd9spWgLcFmbV3N5e4+WR3HWIQuh2e4MVxrtrXf4Purb2ME1E8rKMu5zFmz
7jUY5XdLmXSL8nIjyNqLTZiSMxil6/kJ7TIsXEDpfTWfXisIgPUV1GJ84EAO3OCG
o8sUuTL9OjlFhQwKU8Ev1XmLItfenk9A70kF8esNC5L0nhMHi8X/eA2efz6ldYAK
QH8uA+eK41DvRmBRyf5fPZXsvTYKBjbaqyW9FfnMBJ5a/t4jZRl10EiQ/GcaLxZq
QRV1qyB/0oQ+D9aFXF/hgafdJT+XJz+BWKFF9rDtYBcVF4xnyUSTK537ITj8p23J
V6SX9GoK3g/Y/B++TF98HdvOgVL6GstxwoUhYPIvPHRmNkJ/fyKe/UyBLKsY/Kf1
wOPEaiPBPatjnyQPHt14gpoXyODvQg6rJ7bJ4z6GiMROSQ34we/AR6ayZnsi2pCH
/mTu0tkr+p3yRqRucdn/UafZ/Q7uTYKjuaTbz2fZ+v0nu3/RdvGXUTNLwsn5o5JV
oW4dCbGRDLxjlMxSOUvGn5wklA9ejZkMi44ZoTwdRXsArLOuolIgX8SQ958Fq7TP
ljbz2nJzBO/ApWrLPC1b7fhuZrpM4CWc07oD1M04mIUDEkGY3G9TozOcS4WFU82c
lk1clio9V7goNjLcvRoBm5MywFbj7s/2xGUZaLV3L7v26OL7NI6+7/1vww7HF1js
S+/VbyJK3JYA2Ea8grvug7E1GcHB6hTU3pNvCrhPYgXLlv4AyaNmPSlu78ZiFdgB
qgI68QUy1ePXQDckZoi2YnxREBWYKA7VEyjET3xPw5hffIR+e9iF1Gs2dMOWDBMm
cz+Rsu8q9QAWGLgqeJ+Kq6jCFUYbwoaxsKs033wAY+HgE2R1G+2xKkWQJaaqelqT
IW7MQRmEnNpbyyf+p+FpzqkqdBKDZFKf+Rr37CR2TIsQfu+RuQtHNRps4qW+Biw/
zd4PBe4AB09FWn5fT7eFAuAxKnYqHesQ8H6KtGk1vZHDfCEkxg+T8hUNLTxOdPz1
HGXn0yufvRJbFi8AOymdi39R189e4bSbI7xnd4V8roQI51mpH0GVdiryiNin71f+
cAO4Lb63Atk+SJv0/+TgENwLiNZy6GGtI+uaYVAoxpbQqzv1MUS7YAHaXe7psXR1
kSZQbBJBWQuXc8Vwu86Li/IDqbsqyiEX4XYwuQ6G3eto0xPXUN10eyYCdOso4Mm4
EarMu0aZ2RV37EJovFt0lkVLLQnCxdCjnQ4v04CVofgQc6yjUX2EguonUwT5ov7S
iuuM5BJLbgMoXAWCkNIy8EzYDklhnf0kPghQQTIRsn4wdLXQ9gbc+seh818//Vmj
vZWojNY0m4PUEq9ehn5AiLIHe18sydOdofp2PZiw8y3/q6Ms5DBs7coqVfGHm6j9
FB8HAI0eZpZH3zSDpvtMaEloAp4nEHyrnGBc1gk4TdXQcqVJcMD90s0xrozzVxKg
+LOmOAGYQArMtv+zm7fRlc74MIfAZQGcLM0YD24blbgutt4GAZA0dQa1eQtrUm8e
/BBv4ETznXdaOwDPECnGRZbrJ+/JS72Inwlksm9+upALe0erzKdTKVRLaTo4ySjL
xgqcebeczFJVQip2qmTCWdXCM4r8eHDfCqKY8jk2gBbIZpWf9p4SSqgIIKy1I4QB
f4ppQ+/RlFRLaIbCiuPqFsWD7ib2QN+V9cqF9MKtn9aGJI3p4Uf2+lguGkbGUDc3
Br/Ngt7El+AYAYd63x1RhN0lNvwlaIUNfa0lag3BuiGyaOvN2gAC+f4rM4HhDU34
u6ulyLHRIkM001D2eRg+XmkI+/8gfihtdyyBvPKQsyJLpITuxRlwm/zYkYCO+oMe
6Qv3BMsG3kGJJvp/BVwIrIDlEY5wB4wvhVJlRqXL/ZPl3/hkWUEqfACD9BNt8LGR
sLVLj+M/ShgkuzgEjWSmLewymr2fcvXM1HXwpIc/HqDStp4ayywF15C69m17qq3r
4uhWYqep4wxfwr2qGhFhdgi8YehLV5KYT1JqJtqpi/M8pFEyxRakEyAFhu08p1Rz
RVddVvzsxWt5/2HJDd9DJfOPAqCwXA5xi2nZuQYwbKTyl1DLwQCWgDk7ZfxEBVtl
wujGx2cuxJFFKA6YVp/y7QoaumauLNFmC6W2YFIAXyqfizzqSRlouPMpMm+cmgQx
HxlDvVbHXuqVF/bvU5ceS2fy2E0hDVSmr7huoW8ZWk+yl1sTsKcu5s/ZUKsLPBXz
czBaswTgKdUl3wSRfwLyuThUtaqogqjU/A9NSlW4tK/ezHdYBFNTfea07c2jBptH
kM/pghOsr6lkZBU9ndxKEtXcssdBkB34HA8YjwpT/sLn5Ej1XNHXxPEe2vn/OPUw
cdKMJmQka66MezCiXpP2bLLstoTx+lDaEOo2/pWUUPS7t+eM56ZuFxwf8W2mQ6hG
rg1dpDyh6U51nrnfASPrG8zS1TSngVdtASDBzOupvOHc9FfyXLliT+H6t2zPB+ZI
D1ZBfHsmMCkxP3/zy6jET54rDv3Jvp1afHXw25aQRUNNntX9+pfjeutM82D1tBAO
O++uxSBAKbn7niKcb0fAvHm6f4WQRmnJTKr0q9mNS5d7tyUmBk3e0zaK4mD8BJII
z1GAE1gjqkr5n4thOWPEtcLj4EBPHqHqbK78cLorW8HTLu+jkSKD2z7PWF6dKt9P
BmepF5T8nIzGhmuTgSZwgF7bHI/32NvpAkNAlWA05m6QLA9bifAFAy9FIVyNfKCE
X18mE3HlcB00oKRj98u9qrltCn+xr6hcu3gpNqk0smkazKDBudnpKE6Cg7qNnjW7
tQwBUtvz7SaRmbhQmCX4YvXJPKUmky4uwXl+zdbWkfAOMMAc0LH+jwrHyjHKsQKf
hKJbTydAzcvQOOZeqxIzVQsXjjsVESvGoVa428SQSDiJN1biINyXYDHuLFiqjkaY
QhwaYKswkr4p9D3g08Ntu0BO+IMj9G1G4kdMIp4al7P4e9phwv9fM9Vsdh+pfVxO
lMttQar/wCjxCkn6xO8p4CuDzpbqJk8+w4gOrYhWD3/2LRhGW4Nb0+hjVRY+pgWH
yQ4XB+naTLD96gwb2Yyn4hYAlv767ANM5r0G10dSKXHXr0yjN9RLKQcppfw4Fra1
OOVWdPxoGRfs9vW03lZbpXDcFqxCRDen2cOkmiVONZKuH0zfPq4C0FNdo99OwiId
RJhbR6+hL1ZPVyZkjmOfdBZS7hHBHYeWKRGJkuQZO1w5Wd+pdrvoEXjKbRZLiFCo
BzwLUyYCFI6zxGQpjysH07JtztuH0ggIpHqzBG5hOIwmmRQOsGrhRcsx440F/x/Q
/+bxs9vi3Zm4JmvZbBtTdV53yByBHSaM/H95Uzjky8Cb7qgfYV0zvnbgdX0ZpnrR
5QehrGQ7Zd5PhNi/gDPk2GWqzRhJ6gv+G7BNKZw0ekjqZUXtAjZxP+mP6JiMQGkF
d7Vd0FoV7o4mZg1ZueyurNkL1HrYXUcrf6a2nUgT8Uqio2SLbhB7rPp8ryYjYHCm
F2oUZs9LAa7Ca/byD8kDxPJGoOdOpVwrfI15ESV5L4q3pU9mTlfJeHkNewgTes7X
YkyccCbqaft/YGwdTJj9ydl7hmajX5y2eTfYh7mkw8aMv0OJH7JcLnknfgjOTUUD
WFdSEsoEPIqyjLioUbE93BRrBFdR5llQzFJrygB3rgxH+GCZFnp4tEbb6xx1IESX
ytBGDx5LUdO7jmXqgwMbFLAiNISy0aIysnywdfy87cIoPKSGrZXNRABNy/JeOk6z
M0+Z+Y7vGG4rbhh5MQyPYkvlqsG/OSIKZF6X8WorwNJ5fhNyoxghrQ2dMpQgObEw
PS3nWTvuwkaouYrWJ5R230x/U3RvZIa4IekMjqC0An3fQjWL3pgEXglwUG/wq9QL
1B5xjVS7at15O6apZlba0ywyNQeoqXQB84XzFgQMV/W1D/Yz4jwYT44dPUExmdyo
Pq+nb/1J0oTQyr8kmAnrduAFxsK9aR9QabjYOEt6iJIfqJQwflUqKNYqNi5iT3uC
MU3qWhtYGJwTyh7kiKj3ST0W9eTP5+K1QXGGf5EsqQK+HE+GiShPTqvOXJgpW40o
rYzg3KOJHr6rKgkTkOdB39xOQJxrwJL+W37rEjk21CCdyX5/LAIkQvr8SRGbnrbT
LKHdGI7WDZQCbOtUz6Z8HAaFuFkX6F/k0YKRzc9h12tBc3ZtEwIdcIXB92MSP9p+
AK8xAkbn4X+WIKyn1auUJmtwIQBAIWg8Fmu3i4cVKJMk+KOc+4VTJNnLPI4Ww7xn
HvEQkCphrrwys4JLp5BWh8UaoB8ZfJUB85/NLq5NvKuRiWpRLYiBzUXSSjL6/zhW
Ta+c5tcycuHv4X6AvLtpqgdbzKR4HMTTmmzzMUR+9AvDrzFjult6ivPa+MLovpE0
K+OQiKXso2Q2BtDxbxmaZnU2lE68stqaf0KB7w9HZVf0y5/7paHWJ1JR6Vga5mF8
GTz2GJXQeAXwh2euebTP1/o5Kv/NdIfcy7QgkcR6oute1RTYqO1lcCun3jp9wDdy
bcqbOEEQQaW1bfrVEh0k/nO9X7MwCvxe9OfhShXYjPC3CuOObxb+WMgyeHyaP5N1
DI93E/T/Dnr6TBeljXAe2905I7ko8Phq+V61MQv4go9kGDooBfw1C26xsZ8noXjX
BEuZwUQ4UVIo4Q9B9QdSvoDk7Gcb1rZz3SaVKWW+8nA+dYpUu9m4VWgWYCkBBhQ3
Im3nnMG9w4CBZA8K564ZygOLO3bE9D6sI4Zr7MZbySym0aIRcxkZsUa9pJ+vFFxZ
QcnoGb9w2FKPsH+qs2Q5NggnmIXDIfQu6gT/hbqzfgfEdIQp2+vCoItTPOyr0FkB
w8cjdFz4IvpfSs4pSoVIAG+tcF0ZQqibPYfG2Ykea4OIUNCKXtLuiLIABNOgIb7N
/14roNc7saZfmP5TVph14I2poS1mkRJ58OoM/Ju3rz2SGD9GiSPZzxhz/MQ1xOl6
XhoF2XlbxGs14VoN8TE1dkwLgcWzn5NwwnsSOGGwzs8w3SeEN7UuggwzzOZu0a+A
jsKuMAVjqWTveTNTXJuW9bM726/dxfkfT17pHHGULa9nw1L7Kk32i09DjnLhEd2n
sWsu9h2fl5lFE3onzvdL6K2zn35tPR8udBqpeOA6qB3vT7qNMB9SJTSSGmKMXZaf
F/BtdrCbR5ow8ET/xQavMas7hi1W2W3XX1nA3Wrvh/KE5D/cbrFmK5XYIcs4fWk6
tLtqyT/hAvrJn7T+ZkEz3Za98IUgm8QYtnWQ9TrROsGvd+rqDotKRXibq4uqV3dE
RQybQKzwVfaEvzR8d9G0PU0TQRFDnNumnVe7R86VYuKVSUAvovH7loAArhHVhFNr
SUn/hqmwdozY6jrF0/DmuPdJ3b14X6/3hQBmJoj2geDvrvikX+zuTlN2os+tLl5P
OeqwybHaMWb6VHMT0V0rSu3zfG8EN38KBXaIwIsIifoLIMb2no6kJbY70kMaWCmf
90EqBNHZ4wz5/T15nNeUS/nBwz+F8dXEIPORJ/s2AViZmy8fbQXIgUroFo3XpAT0
ADVMeDVeSTpcVUiUk9yDBgI+CeFu7qvkCI/EWiYPXV6LKD3xeaiND2nvfHTqLXft
/PJzwoqDCuKI841tk/XEMUMFhyOYkf3Gv6RYQVbYke/blWWwX8OMTrNnkna46PTW
JR4m8dU6bNbAvVpZWI1G1UTV+nXoG/wC++DX9EJHzYdtIdLTDw00umCYzFJwlWMU
JSFwNXw4iBowhlIfxroP+dz/JGu9yG43LZW1FypozrwO1wbouH6iud6D5Iazc9ho
QIpPrT/XRtXe1V48nDPgcJmtaalaJzqVQ3ycXQHPHkLe2M0lF2B97DF2Em60nl+v
69a9tgGnY/kg08uRai9QXbLcOczEGthi+uBex3+QsZ9XFmCi/0tqr864X4WS6CY9
fR0Oxt9dwOfj8tdLZEckbDevclNM8UTb13b+lwJ0eYLa2eOY3/kLt/ZvTfMOefec
AXk56sHVKZ756+Mdvxt5dOhh52mazORAb9RJEIrpEBJCeqB41FhVWfirgXjRhKxF
k3qu84B/L4P//VGgAOwh/j2HHcnUzl1ojepHsWL9b0+Jaspu5hRy+Pq45IZFvD82
HZKw1lSVUSZcj9z60vzyrrPAZaxBY0u+oIld0LHGPsKM7SGa1BoB0R43f33kEf5+
yoI/qgK8m8ptfCQ9Pl9+BNLYNT4mTCyH98Fs45TRIcVJaqsonvFvmHR5OW4utZQy
51s/pISf4eAlDr79FPYaW+YgqqxHy8/GUqeR6S9WQIKolXSIbZJoAngx95P39i/R
epIxHtgEli4NCQTiN8M5nM6uEO0fXiZ6C4dJnhLgduJhN5euuU0Q06fjEw3WNqYx
C4QPKhDXbvVOZbm94/fP+WlVuiOJe7MTWFcwNFYBzcHMHeg3LHgdmzzvv1LUAHJ1
CfZa16qk86h6m+CPll86844ab5tqoxEmZ7ljqsKrsp65++rX/cP1ba7PazsLfoZl
iKD39/7uMYFNXrj9c3ONwaUoPUyYBvdzAPiLjPil7Z0kv7uHs+qLpJaxZaZ404Lq
v/usG5JLXKaixX9bZtrr4ccKQkf45Gsltl7hvinSzFhLoEYXlkudevwGOPdAY+x+
h7tXdhNYtYVB6yLTIg7tv9f8lNRVYLbeNU0MOcjtyrtV5ulXbCdCG8RJSNbOmtdz
XiNpf/7OaekywShKylIUO5Obbj0F2D1Ne+8Cm5QnqjAIJe66kPNJz2mcgkTxsOvG
lPy1bYFuBZy1tjcsFyc370rQlPcgLOVLxaEa4i4gOSQs8aS4BrosMbNLD/PS08f9
uFQVpOSN7GDKvt78XNbfuR6ZpwVy8DcH3Us6Z6DtOnLKWSy8hYBVtrcSJ5B35Okg
G3ds56QkhnzkKyhXPUjOQ6kmIEf5uHSjB+77wBm5pim/t02x/uMhBwwSfK7BX0ip
2i1THXfoqQfSQkaFV1ivIIRsVcReI8MXu82a3T6bKTLl6P2jsOfDTDAABAlffpX/
cIitzMycvpFozUGYoOSIIsmUTCJPJpQs1dRpm7hBVcrL5welxhXexzrh6JxB39P0
crP+Rd7rWGbywsrha4qo2nCKwU0qFKXVc9zj8KVR/KS7mXaNFFc2RRre6X9N+dZS
a8l/2emdie9Up6myphy+pxIFV5IilEkQMPJYAKZftARC1fBPAC5J5uRHippE3m1o
R8SH5uFQitV5xtTT86v7gyoV6oV2T0/pOs/2aCfDT7UkSEHgDb725/X8ykumNjtj
dLoeW144VHaNH+vXfMqQHclyq8ldbMVfgxqYlzRubAnVJ/uiR4ZEHnbawWCAh8wH
9q1rx6MEHzW7gMACmuUCFxdmbFSv+RM4ySVqE/qvDevL0Fp75MaIspWM7Rz88L0O
SOGLshJrsc9rBC8KCoYo5Ofyn8pfUKNwjg2ENIkjlWdE4BIIlWNFqmPMJ06zUjZk
1rl9SSJRgvCL+dlDH0y0Tk4IfScSyTmmiR9B35s730nOz0fwPeCoAkUOgC0Jd2pJ
t19uw9uqiTyPAfHSEsC1RqIr2EGKLSLMiKeVlcpBpGThB3dBxyHVvqFw9v3JN2Ae
Pz8UsPmofnOGsu+tMr811Wdv2vn7cYDNx7ySv+TKxfm4L+UBvHcSdcJbAnjnE5rj
ijZME/9ETbty+Bwze7IAvmEGJhxnKoqPnuJcsNn3sFwkHu3p6mW4wv25bp319asu
FjvyQH2G9T/o/ZO523Cu9mmmURnbLBYm+cPPUd/jkYrNt6jkM9jlkx5XCArs8MYs
ETo22+JpKxpU2anwxSP4cXucJmWp75Ha6S1cLuTkTTUQ9AOs7CPcU4T2X3dXXZmv
aqJpYkJtECbXyKKvkGv7IruNF2UnA3oF4XoEkHKP4JMZ1DxVvdJ5nm3Lp/nGWbyo
P2qIFVHDTnNUE78yRdetlbFaNqSqj3NoXB59ht7P9GyILXPKmXVPfbIlOQTE5Uaq
7KI9RuiSHNIaykd9cTeEtq26KUc+1guM8CGAl5hKHdjjopKZwdj6K1N3txjulrte
M8TAJ3sKzSLnZO0rG78ndDXvQ/ARuVgTAdNBY0qBNm4GUEN7KFfyiS6D6w+eNbf+
TTtwGz/3jlrh7SFAaVPGkyusYwAmcn9glrzifaGhqYKCa2ZlhVXBOSMXuRFH9ZZN
rWVsnEF8bjS9F9JGwrsJnO6MEhezLbN2L4neQBXbJrZMsjepXGgyg8cAn8UPOsX8
1As6laPOEtjVugXUv5nWur+UXQfPIgJNeNCM9ICeWlPA2PYaashBD7AL+5RPi66X
gnBc8uIoidBNdSXRTAO5JCyyvWAIu1Yt3not9Bn/Ua4+dupEp8Z6V5SgtrSOvfep
7HMkVhwrt4fkwnboWGkgjC6IksUx3CLjcV8VGMNLwRleAI9tvf8CbcCUKC7XO+Ca
eerSyDZidCtl2EPTeodr78bHipcdUIH0byu8gr10sTT1no3v08u3IHwuPMk6wKHu
Xfde+7A/J7ZdVYhjwTqyR3jKIOleD9ZBq88+sMmzpm9raYrpEnqRebbC8vMuXRTx
KyiOOX1DmfOYYdTRka5hF9aEMNxXlb0vj06+yPx533MtzUH3vO9cQ3jbwZiveU9t
TLnKj0hRrn/56WweEcZQhJiIQdhkBJYLc3fxAgI9M4VztxQZNVVciUmj0ZsnYzfR
H3kcaxlNPK+0eTmA6q/hCG+ts7x/IZD5lQ5yzEyO2pZS08cO9hnd7cjPiH4rDlhC
yASehlriDjHsZelHIxna+TtQSxeQDbdqKcfO722y3FAk1e8X2CJl/Em9mS1mKcAy
hoAwq/a2Cyadiyipgsxi0NJHUi8eg2MDZEC1UNXwlL10iYshF8Lm2f5aXf7EIqVj
3kKJJNvIh8fnIEJiSSYY6NtspwH4flwZRBNCGVapwWg3Q2jI1L9m4ynqJCZJUJSS
p29WvbQDX06sUv8+uu4FZPW+hganjf/usAdaLpXF5ksJ1nIN/l66fTtAPvBQFij4
OrilpzEL63MD8BxYmdV9z0L8EvBPWbmmsG2bjysjdqWg+uhWWKg4+zKgpv/t2aKq
i/gJj7v/zXDOY+OcfHPl90v+aRHALbB35KojAxhOcURz+s6j/01oZS5kHO3dQzfd
LgTGgq8Zl78qwTMHvvy4ge1gFuR+apAIxe1YK5lO8ZRswRKP7naS1Tf3RLOLOV6e
1BDARef7YWMqVxyX9eqa8xsR8V1ZB3IwgC+9J8PR2tea10op8+EIC12zqcYkOLwa
0oR0J+gBgvjAUfZ/kxbLJb5xVxw/Rx52QTa9zuRpRKuBEgyXdXecU7rMukNE1YXR
t65ArGbCW9IY50w0EXTwcHPUqxBoPT8WQaEbMCth8J1BVgneATeNjctRCOu+qckR
3zC/c5vc1A3fdYGiyArvXf2+gH6h/tJwVtMTgR1JkbCFEwv8nSlBI1lsXdjBOQeY
HbV3wXmhFXzdQ0A6LryPvPsZhMpcqtUVfPKmTv5loK4/GZnW1ke9twr9lbJpV+Sc
xUDOjSbW+qgvf1HN+g/4XVGjlC9MTxB8ffg2uPuinxWPFskgvYpG1pTeHf4ipZtD
O97ojn/YWEX5YxgzsHTyBm7HIUuAY7jaKapY+Erk8/xLjAALC2XCEQrpm8M0A5dY
RXAUTAYAa+Fl++OpOGszPWUkHu/sLQR1mo+B8DPSPo/re5ZpxWP0J9X4Rnx2C9Ae
3hhrvH52V7uWh2ZSxP7mhzDf3yY9HmNx2YeH2L6DwkRuRv3uy9hU3RKEHCaEjdIa
UohrJ5GSAUCUkBZ2aW8sm5vDxXkEovTFh3O2gw9HRRF59XH1btHeHSJozNEM7ZHn
yVGvfgOANkcFHNdsV3MNu8oy6vQ9MQDh0Awa571/uKyE5Tq4czpmtkGn0f96PZ3R
ZzRLdo6dhU4Idou/hN8Z9dQ4MNIO0UE4GtQ5JVzFP0C37hVFjkdUNwxU6oXGRnYy
nKoMYXB5Q3gYhuXfdp7MfIWj58E/Arkz7eN2+UQBCbGWg1PdTEnzjRIXVvROP0QX
P9HwvD3ZgHObrtDOqmCg6bNHWC9y0+f3Ipwn0sSk3Pibse80VewInCgRf2QKZBoA
tIio74TBsmBZzq60TSYa+34TNEhwr64A7EzlmJotwN16PN3AQ8NP6oIQX5wUvcLg
3xqpBVItXkcPDHNUm3PRYpKfYo/Is8vLNAiojqtqkQ55xRer4a+QMCc3sOieDqam
/wgBtrOZd/11MKusP2ANZ9mMIdw8f679gt+d8WsnVVHrbzOPfg4X3WfI2/6N5coS
GKljIOnjWDW62/UuPcvqX3xuild1dlPpU7xIFgSYjMbOBsM/lc7h69dHJ5BkQIOk
NmSOdj7eJlUtFKmVmP2g3namdeeEM4+tbnv8mj/uGC0VyBYF1LaI1Wz20ULPHv6/
uG3RiCYu3kTtAWRKYM662MH1wZSI54sitg73jc9RdECgB1tVo9pzJO/LXkndJiaD
Bi0h6ThHRlsiwt43uou8dRJPhBiG+oOVLbUJT9YvwrgqarjrascQPfGERHT2gX+l
9UBmAKLRAD118WASIC5vWHYJn1v7BXa8SMJjXBdoja1Us92ktH2NYgf3+THhyuDk
uAPA0ZJO50WyPkP+DA6ZQExik7LNMn/8vblPZJbFCMpWVOybcW8JRh/9qWQ0dPAN
udiYJrC0ejg40brKJOMHWpY79djLhL76QlOlwwj7YhsuPLA8VjcEfz1T7td63ScG
Dd8y7iKLWWH+gY41/wpIOd+QwqAfTW7k+zG/LCKTOaKPmqgiwnLjvcyJA9D0Pg/V
rbRfkZGtLONqoG/yIVxHqPthkARjy+nvvPePW9GupyVpYi7VKyesOZJAlLXRSJpp
bg+wbN04szbPLdDpVtVt+oZjrq6VsJBcYxs5qZL0SOAxXkMS0s2kFGRUVRd6HME5
h0OxaXhjGC2XudJ9vHnf6omM3UOYY1nb+UyWfCa4hr0kQ9l0LYCEqsGcGmt0hleK
23YVNG6nSufgH+oWKDlQN2rIdfSTfllJNuDrFtkUJmM53wgBq31efyFGBwNF+dY1
6QY92ZGZzRShKesnHuL3iQT1nYtcps7h5JDnzd82E/rFuctnyQCIkESbmKFzTc7c
dxYS9z4Wr87n19lhjzpckdJYKM2CGB4CvFV2Vcj5NIb56jjNtFcm/fMgcCFQ3A5f
IaBjCPTizbfxPI5dlfBWYD1F25QEpxYGdOJcd8PDqt12lB48vqdWYM0aME4SSuDy
ejS6hmoEsH4D9vWu++S7pwx0tTlS7C9rOwDDInxIAq9x4R4UdhpamKs54Sn9d/vd
MxD69NOHYUoCYm32wHeGcpprMRYThOwZLpxvvv3kYuBpUgzSpOvTs9jzSifWkwO2
F7T1BjPgsDDNjMmnCUwHeS6PLPBSxGk4Ncs5KsM1wL0oQlqMF1+mLlIkoFYIQlTb
SDLRMnzd1TrFncYxPQdiUnYN+U4HRaJzzfhAG9Pc9pxBx685moFZOp09jS7TekUp
R4yaoi+8yxK/Oxy+ivnJYL2ScqO8xMPpVi+ghOYeog39PcP8312RBb3Xsc2O6uv6
CbHS7jJdUD7OScU3f4ddUb+To0pmw2DDksLhjU35hAbYV2SbDIIBc1BKWaYlw7IE
qL0Jk78k1xgxhKEDHV4hqa2rz/6jsknuNeDFvYLSCCM7awXnMzHDN7yO5G6bGmvB
mt91T7oMZreziSZEyBQtuLf1VNtYs+ZjS8logh29PnRcGnP7W0M8ol01ZQ+Y5BhE
snHy+icBH6cgv2gCvmVD5ngM1/6NqFIZILF8v4Zq+1nJOuN6e4YuHbam7+8xwjrJ
xS+6GNDjG5FQCIlSeJyXa5UtVsc6WcufWtHeCS0RZeZzOJTf25hXMvKsfZkb8WH6
NN9Jfubs9skV5cYOY6TswHcWxahbx68ISxJNQwx4FO8ok05NETZsUQ9sg0AA7/lI
nh4suhZgnpN8R4o4dKWz0L1eSadmIgCXtnjhEfQTwO5Z6xLZDya9YWtyVxh0yWrU
P/Q9yppUlUPxOEWvmYX21p6DQfs89EUHiHX7/OvIJpUroGITfdUUCcEyBaeLF9cf
z0EfJkix733Moolku5NWc2y+2xdpuyeEYtk+zbPFvTuxAxwPHuuRLhCD31eBv6zd
Kn4wqKqduaFTI92QF93FFPX6DNxDIFHZoGvOA7lLoa/nwXLBRfBCK8sSLaeU7hSn
dwvbXMHm2z42ezxHW8VsNjYw5Xp8xiRUGts9J34/Z5LSz5gPGi0VkXBteqCTqErk
+j1w5SDXNFXNs76dn++I8FC9rTfPD9r/ErXXrzQnByPUVKtBm0Qv498xOq0i2gXR
tzfj6ttVJcgnLXfZ4nDc+duDrCaYqKxbDcXabwEHyzoFZRKV/buSRoX4uBmmEqM0
FTd/oWGETw1oyI/oza7A2DPRFRfOi+78g46SUIxSSyAxcXitkOvYA0eQgWbqnH6Z
0MUHbQSvaw4FvwDLrXCoOa5QlcwvR2X7rKP1SJkncRmJINIBwdYuYNhspxi8QWKV
FhhpiqD4lhHJPf1ovUqBn6pOoVx9osCV/bM4ac6AgpuxjZrZhPg91bToqdpEp9NR
nwou6NMOf115yMON/yYBEogvdrzUVSOBaiH/qTQdcTE7i8aD6SPdboY3cAsowbsA
MIVEmkWYZyed1AysGv1yaLyTusW70DlJCbDa23jHvrO6CM+ObNwAWKHy0yaBDwtE
FpWyhxKm39St7pcZo2YLMZaDaJF9b76oCmdHBWDF3W3PCH+7tRZtfQOWlYZPovax
ezIpDxP9BEvqACoGE5oZyWrdvlMyJCF4ZtHXSixAbVyKjYPFWCQA/dBj7SpNVg/h
jPhAe7I9OoYp0bey0Ix+IXy6J9g8l+eKVH8GTNSDcE7UCbg+xQBOshm0KPPMl2dM
RzFKUaNjFtDyZfaKPT/leVIMYsW1mY+qoUT4yiw1B9ODNujyOZAmNdnLRzP5iR5Z
ixhmgEG9QacoPrx7eyDjLYwHBeGJCpdBHTzK9lBVIroo5WtSBgaGcPPC+klxp7+U
aPfzq5D960VBU6lDd6InPAt3yh+2FS+ObzO8FL+UI6+cBx0Lh1KQmSQx0g66gNUe
hmwV0zii+TLyuNAqzDQ6/1cb/cXlory/weHT6cZWa1L5CSgTjt49uHbJj3Q3KXk1
Aq8Hjd+lmuL8dHgIOkSB+bduFWAiBsldWhdPBizRZ9e5C15H0cbf55q859fnaThX
fd5e4V4yOvtbpF9G9qgTzNaIqM7fHEKqQHy5FWg21evfg3bg0E3gOeEhgEJuHKAV
a/2K4T+jE9FWj8rUGdlNRoDBlTcvcyhPj9r6zOpRzHYyNnARSqZC/dDC+xG/4K4l
FTq7rZ+tlaIzgg93fzCiVDF95aI+ZCxgJaFcGY+9QnXvBdO6tlB7QANCN+1ji1Hv
5A6h1oVJtYv1tk+xPu0LTAH7OqDuo+xgkPqaAI47339rKgZNWEE3yg5s5v6QTz2J
NJFoYG3Ur+FfnytPBfMcoIreJWAwspF5EzgWlHqf6JPZGP8nss8UaEBcTFrYhemN
uG7lW/dh5mxDkrNxBHymv0PE0L3/0Cz2YCKYAgC66ipc8KzweiDcV10n3/B6oa0g
EZqgAVJG6vuPuyepNvKqq75OuC882qIAzyjqajdwcj1eylPxOsjN8vK7CGKNHzCr
Doqi/YKjCQ0+G8/sgtmPoCKzpfZVvL3R85x3VbdcXi5mQDja3Q3C2SiCCzq/zqfI
UGTKJ9BAE/aRPoqArLc76WCMcpFRhVtmEHNj0pzfA2YvlXf0OOY4VkEsnYn5IT4Y
Ybvcqnw+8TBqAxQlQOWhPrBJgtBt8JSgbDpnOznLJxyBN8loiOHS+lX1wTjxb37B
hPnnIy76hqknPFjiumok2Y/H/Xkiy0bFHDNC0NgYpUrW25nffqzrtkPJEI0goitu
FJPZeC6RP2KBu0Ygw5J45aCOf2sIDu0BO8Gumoj5ZZNt61zmGUSWjs6r56RX6vIF
/CqmTcrZzTb+a5tuyTmhKG2elxIE36z5RddD0B3ips8oeiCX+ewkyRLDhdk5f9IN
WBHX6ms3iXgcTWWQ1bPZnCQDTaUI5PaIIcvQi+NjEsj7DYYdiuyhKXQe/RRAvfLI
G3H/1ELbMV633h9qnZLNmOQeJyPxWSxLRisZMQzwqNA1V0n/pOkQh3Q16ZGppKCF
vmgs18Qwk8TACQaa/9eU94SIwVzXkgLg1+UPTodjIUJX34CZJGPLFy4jXYSaUM9p
shiGYVGkHfUkWgHt3W44YM4TUoLspSlJT/jyWGQ+mbdTxW2zOr/XRlCjTfejtwIa
a8+0qrDeh/5/kkQc6I3maKuKzs2MleLkVxjHdu4xIF/1F5dKMRyAHL3BdsQ4vBfC
6SBLiOyEKXq5aC/erSRKxIq1dOvukcGS0l3kYIf+URd0fnaavIpT1GLUoYLNIcQ8
PquHLAQo9nV0iOs6OT/5O1nG0f8kcgPl5dH4cx4Cw2QH/7e19d6BMadUOQ3Pz8cG
3XroMqJYRgsK1C8L6yv5ZpgL7pFF2FPK/xTcvRMw6KxIQv79jZSQeDsr9m8y9NzZ
O2vBIAS8OQk1SmqW/KFJjmjhWgYAN8NLSOt/uyVqMXk0LeyIwAM8B/UU+vqOar0K
O0PnUHsYtYO3B0V7kXrw8uYy62YXWPfl23kWNJ6f88R//LyaVed0f2IrJi+C+WDE
dBr/ZvYJ0vbDBzNqJi5Qv+IyG5bUJtTkBn1c9GeBcUtV2YQpIgoVaqTfhF1s9X/J
4F4T48L8THtEvx5LEb6suCzncYFKtsmEGi6xvoz769s1vu8rS5iDRTlkMVUqNXUD
jDwPP/M+2eXbqIvYbqldF+gSKZi64cu1Tlqq/45/9k9e5NcpbQfjF4//e2/adTrI
VhU22GVkQXZeTcqadFfK5KQ2i31LObJtlf2jKPZQW30by16F0zBkHMkhbC5miu9G
VsP5bXilJN89wBinPWX/cmUJl7M27oUIkfHyA2wzKC7WuZFBouq7Cw2TGAmAB4fz
LpID6vzNiDailk0oBuwxINUiqTMIQQa2/YoNVoCTzjnye1pg9/a8V/m4h7KASmTB
VyuVUhTs5KdE/SmlfQnZqC2XtCSyk6kKj1Wk2JM6/rj0hm6QWl616w30dAvjTnVo
2jwBKvbOndKVmTNio4l/eZikO4dNTKP6wJjDBL8GpmIJ2jEKmQBuT6rsqIu8Bk1F
dnInFSP68UdPrADqMihcSlqJr8fqhxUfc9aAcebvtRiPF7E474lSotkoux0rTJ/V
iAibppBoiGf+mE8mTmT+WxZsbo1Q/SZh5IHJLrbiymA5YJ4C+xOO+GkJNOxX119w
183+RVa1DGXvZZcQN+JkSdYTjUXf44azn/h97OtzpKVd99WFdJDIblqOrz9/Dgkz
q8eY3EeTGmi88hSjkI1P5q1+rVdzuBx3FhDsGJDJMZpLoqBFQYYNxH9TS0OPLJKo
F4WByjObnUKKbuTMLDlGrxM1k2l8/VvHEgXG4/+bLkiGE0XV1PiRKAvrZQcTr3yk
3TPC6ANdcn43/AUSCYSlCSnbaS/q7oqi9Jc5Vu+5bIpglmTyAC3BiaE6uU/YOJ+A
qQbr2DI28cdB9hmnSjtm0wzxRwqzAADkfCiiB6nJ1T3jYfJXB98wC7pCHXrlJoYO
6JXdZAbKr4xW2l6IZCmP+tmoThAENxS8nPRzfKV4+L7RX62j1655beii+M5QVaFh
xV4LniXzNZoQoYULZik37RTDW6jMcZ01wO33jP3Q6bsVs28irOHBL8Mon9qZnZo0
ofyQdg3nVn4Xa0TTjH14HDzys6aJ9dPgMX0IRCoV21vGhVX7lsHDBM/o3YPx7J0I
hbfknU/XApnUfb1PvrH4x3+SKcbwI9vLGAt+lkbfkACKMKbVlekHFNPkSskfWqK4
SENSCNsmV0WZmN+khpyOWIRV1971h7cB5CsiC5bivSnT/zRqt0jSOKC4Q8Kgxeeh
uD0wLqdNUllcxhDT+etiIxqGkBCeizxbBCq2h0XlmEuatmJXpGFDkCkvYD8R59RP
z0WBuv9ZwAE7zgaz/BiiTv8QoAHbk8KYNu2KANBXy/eZI0zuaDIoybU9PM10c3uI
U0UdEuT3/G+LsUCI5hRKrKMraJt+O90XOjiNdyhYrCv1mk8bOrIQDRcxnoHcJpy/
8AfEIgyjJi/SeSmD0qTZT+m+sQLRuYtazy7lHoxLu1M3qw9i+EAshMV9RuNwMHFp
z7AIcBAQeyJgry1ijp2wMDTgaYxL+sI+39lFNR3Az5Zn46nobDdw3yK7BiBBIpSC
Cgd4ILJnSYfQJ0lz3Fwy77V0oe13Z2yVDd+5QZsGKuZGjmupxpBtxRMnghz1RAUb
7nEYHNh5xyu0PIoCTRTu+D+eXXO5simlOHkV0iksNSsInnZDJ5Ms357F4XS0MtRT
Q1dNRGVcBE/8hfQ8pWJWVpn4BqI5Fpv+qGkdLh6+3wbXQPv/Zt93o3k/VPOiRd0Z
XSUq7dEOSuuX6vDqhSarxGU6JiMK9XTVJdeu5n0IkT+eJ+FFT+QAkcROT3tVeFxA
eiVE8LFSDhjuSwC4xYL67ciAqTg0xgvzoLFv4Ta0wZZprcnM2utme5v6L9lX2y0E
/sCySteUsnG/s3exmPWSGMYXPIP+PIsD7wtnkWDU43z1zvAGYjVr+gyGLiqMfb4J
TWlL+565QbCmHzSZcm/TW53QNLSGKw927FanlluhWMG+irjOMyyoXPVVSzYV4aVT
n9wFIYvuPAtqb+0sWm4/I7L3n7Ibgzsjo30VNRKrNRVOYJk5aEFbZU2AI5qEpFzJ
z9goi7g880lTPZtKCP/qlJVp6nIaCkAuGs0w1EFUz3He0wD87UKJxO8VqOavOkO+
g4D59ozQCAN0Q1jGPx51zLz8htgGFM77kKPRuw31XaoApP+nPoMeJy4TO+18vURM
owcLZgeIYzpsQoEKED2m5q6bW/qF9CcoDmLBFwPWKjM16zar1S5KchQdimXpMFqj
KUOlsHIugolGulWZtBrPeCpXyuBKwgU50UlbhovzRh+6NSBLdtRMCIum5h0XWmZv
7KQdJpPmxtR1ffXKwr7I7ZKDyCXZcRmVphkiqkHWFY+Wll6iNb1VyPTuBh66bXrE
d/xMfw3C9oVQ4gM1GMFs7MU27hU80EiCB3sKVqvfhgrjiNpvtiJhJ/DkSYum2b2x
vefSQe2ZaTvMSdQWiCOkI3qB2QKy+mVQS5Sra466qnhXxNTdbPQTyzI6npYt7GNN
1fs9lzpv+nm17YPpHbNpxTVqtthMETLsiPgawgpc1BAgnYTWJSWgLMckaMruOMSv
T3pjtDKuJyLNstVTaA+Vg2Hw1J9mzl/ItPEbzkX7A/B4cwi3AxZb6yEbaHZWhZoV
JjcsTSNeEbbdd3XMDwRRTFknk1IY7zHmCPtVIcXcoAM++oSMBhJqAjvzXCHbQF/G
FIh81t3PIZhQM14D4jbAXDN/5eanCdL7OH+SOVw4KFLklITI4921a00hJ0iWelfw
cjosXt2gFelLbUOsLgMnf9svao2qCAp2z8k6RTWsrbIxTeWhoBpMeNFoMcuM+AIz
Wi6WbEN9E4Ln6D/HLzdM6lMOnuvjXiLOS41iOvZ1U6+HUtuxi5DEbaXkH5FzSzPO
hsfamgmFkGhe7A56HI5iMcdOEjvPK+spsmHAjy2V7PSXpHyX4bWRlMXDbihU+lPx
dVuIjsi2I0wV6T3d1nKh+IEWqI/u61g53S4YeWqhZYllc2vPlzrhlU+vZVLAgMgE
0yoGiLrt4D9iVKgB/O7cIKwsvqf1I/azviPHzOhK5uHQFhw0qoBmKdUoAQ2+fxM6
UJ8Qw5QEbybadjAe7Cm6BkV1aiKUNvBDblRiHVM4Zozwhv5+VwqWI7HuW+aqNK3w
VtWLCESnmgkX+3ri5a1ebeKp/95SGKLdMuQ32kccoBBeWtngs17bgBYOexrRc3bB
ksw6z157lwBVqHnGzshVjs0vHPVB+DyZo1+5iiywi5dTE7pZQXUESxBSDQ5Bf51C
ieXvDtD8AJBTd2v6d9L/1MiLUBKs3y4f6PTLH9EnWyxbLMfh5vnLtHsVnwSIdhZo
lkWavOYmQCPLgTQMyYjM2N8tLz3T9u0r8AZRgP3b4d5c5gmBdroe6bLZMfbF3Yc1
7AaVEzTvk24FzFFpUMOV998DjwgSfz9Tpps4Bsy9Z4riG9/7x5I2i6cESc7wR/6N
aRZlx/VUxm68Vqna2MTU3EJELinRe64+QpLCqtsKsVdYv/Wo1FlVNHihrSx8BWLY
X1m3zOec6VqlOIqass1jRquhBnwLO5C+4LRLzfe+W3flpA2amDD0saOcgVlEjpT3
wriAmBIrdMlH8ECcXwToFl/P6ycSsVKEnH1SMuI59LWq4oYKp3H/eZM0wsPmhLM1
vrSvqlqF/1/bnlIEskVEL5nqNG+ojieir/qHVvw8oUY+in7mLMr/X9IEM1rgDQY1
zauMH2z+1UJWWMTJBS8yi+sBFVMld2CmmiF7Vo+SIH/ClEj+gp6O6c76knzdgEBw
/0UDC99eOy8IYga9xx0sOupDYBpc1weF8EXlYJqe/66nCHts90cVYpijOJi+dJ9S
UunXu0ahYoaYR/WwuouUlMXApD8mfEm3AQcogk86lmz/P8mwF7DojJeROhxFAH1M
5XzcC+/KFA31+h7CMMODBk0OP3YA+x+ZE9dbGDo6sjgzIdizX9jWxtHVDZS/KE1w
cOrDFvn2zepHh0n3o0z4CTDnduG2NJduFpjbxKUuhUuzZwWm8RyXurH6ee3C2Q6b
XfmMMLlxS0ABGLF5TK/0zITzs+hO/nZ3nlrGypD/UdN1l9HRyogp8YKMUYKrn5/o
ROhP67wVguC6YKHrNGIm1kv1NOl/5/H879NUU0iVq8PCIWiKRniXlnh2uwcYvfv0
MM/qTiYfVfjkxFs/ObSSH/i3fLOFIFKf2Lu6qJNjuUdGlc5jTma3RhPBusgFDfl7
xQGUcGksztLeU1it1iQIHet4QYK9e9Nq+ypNHRAxWPjvf32J45gks3jSv6KWYToG
U4+/NONwwVOhS6VGBc3LitDu1IatJ3j29B5kwrOcPhdRsgKfJ+7Qp7jvA7o4knZv
JMbdNSoO5ABbNn2YbrjRSXP9CTM3bj6fi3x3FRc/Zj2NRgpzfLH1m1WI1+TNs5NT
pqdUbA13onHiHFOtSo91SX4jXOqM4yNHir7LbMcVThOzOGj8GE9PSrd6CBZSRa+x
bOTIH/KRSDPca/QfAgaWRbLk+02/6B3knZXzvre9oLIT167TqHqkIHy6KPn9xMJc
PsA0PftmB1qzp+UaCJ0fgeS0+7Dkf6iXsmHce3IoV133pqEdC298x+S8ME1SgBVe
CC9KUk/0VlqCi/QmItfMNu10q9WDBKOdcgGRkZ5Y3+71a+OcAEtLBscP9AOZ8mEK
Dme8Jh7QTcDtnrq4t2GkC+TcMbtPiArm2MOyHrTnoP8q3IC+E9O5PXKO1KOxkoZZ
25EsL3mLx97iOVJ5oEgFlVffH65oaXWPXdDvs5P80s7eh/Hap7VkNtBhBo0wikpX
z8MNeVJ14qNwhryfDeuBHYj94A2D+UximuVtSWnMUR/vLqCDBGo4JhNNwJhTUCDk
1SnlCLg0R248iWWxOTrfilfP+ByH+eqgsXDUaR5AChUIMIHL/QPyOeLzOF2zUUp1
AT3hs//JMobfv5UNoj+XELOQUH2HTDsHlI7g+uGl9+NbEkWEVVKT1Eo4bd2fSI7u
oTLZbCX00JnVaUIJAf2p0CXW+7pNq2xFUoE9auvhTNj/hozWCvTMPVJYuZg5L82h
lBaZxKDnC4QkbaORQZyAnW4aPK5rBZCHPRlf7QzIIt1NEkUaOHMCGH2uszNE57n/
MaxoIl0vAep1ROHuqo4SuxBrbUqK1ew44yE51qjX+l5zsXIixyZlG6AE97fbdIWJ
5ap0OrlOW5yvmVBjeJfYJNlJne05rAIGEbkuFkDt4BO1uOqa1hyweYFLk6s1LQbk
kNRkW4Az1zDRBO6wZWZxjv/6gwlkLE6iz+S5JBsmquKoSItIKbB0AFO+y0F+ibAG
4/lmYPqTQhtbjSj7q+umOrdnFA67aFuLkRKUt3UlCqNjhq9iUq8SwmGVZGcvtncW
LDh1Xd7uGfv1PDDHQtCX7t08h05LnZoqydbahJtflRbPQhm798fLl0noouZdj5nh
uvvuZAI4KTcTimtsrVqbC76jYpKXGnB1yGQV6zZIkfg6XnbCGc/qkWMsrkIgKdSe
1wpQRPp/vN98g/4KkrMSjZcGLDx5TOm//tmXBPQVULmrXDCNLpJAz1x2Lz91R+AZ
Sw5BHYVJfNdku6RxSl69zXygxUWJPbYmPHKW/6g4GdYLJIdxR4dOqyo5f06ig8wc
PKT7d1sIFB6Nb3NqbBbnApUzF2Vf+axcEk7o18mVHwIB8tOLTQjXeEmuVYlV+2qG
FaD8txJsRE/lhyRw0SHXh2Q4873+EgYHojrsPGJDU5Lx02EC6pO1vuGZHc4d7/U9
57uhXqsR+X4Bup6S9uAVYgMj0xsq2wCqOqP7KRlWD9DwcWhGDhFtpyEqvJ7AXEgi
eD9aozikcRUbc14cudFHQGdkBr1ZCKdfs1EqRb67KW2/zRfuke5Ah47+xfVOH9qo
t4FXNbnauesCUjoWBpPGS2dtlBGHTYnUPgh7cIzmcmcoxaBI2BTJIHmWEItTWt5H
u9fytRFu6D0aSeFp5NZ0p5ckRpusarvxA/P+xwcw7k19ZeY4a7E/pxUWL9c2vkxY
vwHBwIsuSLvh9xAUrjhF0mEzUuSoj/bivV692OfcfsBcq1v5AZoHPEtZHNIaTzkL
KyCZX/fHNt9M/ux/5kDrIAw6MgJDTYIP1Tq5zT8wRzp8aLVCAk/098bvETML2WZU
SF8T1n4M5tSdw1f0XnXmtng54PfmeDMrj7qKBhBtnjq+6X+Icw7CNZfuvAWzRxXe
ik8Kmqi2Q2znzQ5IEG4kgNfbqmi30+CSaYahZfpjlouZIPkYTbDxk9s4SapOeoq9
sKGgh9HwyMOuxt9JIY5v7JH0OrmG/4zGIFz1PyhKhFklnCLxU40ZiGEgl3Lq35Bf
9U+ObpFANk5DfgsmIXlLsaYK3+p8wqaNRhEPGL0mTT7vSAnIcaSSCYtfCmhvb73j
znWVOQ53X41LYs4yvuAjLYSAoPjB8fswJOHHZYrhNcfGn/hLZyfYiG3ngkTQJv0v
7IIzOOEox0ABTSI7oLiTU8HkrC6V2F9pR8QHJronDfSwwoRxsq0UXYXNoRfKvRff
RBhPUrvCBkp0BbEFJ0D2Dz3Bb9HyOmtFYisfKEHGT475XDBsAurCDWSu6/xMjl/J
5to2pHA7es067o9pXjM9XENCAo97vtzGOQM7PttOfWHm/Qex5i99Rd0qQ8UXB0AC
wPmSCSDFOdzrIepN1CENyql6CqOVUUDaKRt1QAf8Z8m/6UywAt71KsHSWcaBrdFh
zLxQ0Ec6Urz2DLfAnt+woIskQjY8zPr+MumJvxL61O0pUtCzJWqtUorlrLWTEGzx
xR1q5mllIQtRZl9iExOyh3BU+7TJDGwnNYpyLV63etfE+jbdTSHRoWLDLp+fm/14
/sUa02BsBim+eYImjXDKBDrU2JfzqS1EMULspLI3zjO4nF/OOL+C0ztlOBDQtzxO
fuGqYcfKK4y7uUaNWnFvy6syrjgCHjCCbauX/XWrE8F3yd/P/MBTxlpZEV34fJau
StdQGOqoGYJ54MkVqX+g0SOz9GZjfS6jK6lF+qy+so3Cy24mvUCZrPH3RXiesbHo
+ygz1Yx3bFmP5n963Q0/dO2ub2MyoeeP69F5n23Avs/+fQguaf/WJPqBe8/VSXGv
JVRsEibu/xsXCSIumTQOHaETaCj6SxPjdpvHXLHz6qCLYnft0qu7Q5IAFuDH4FEk
JdoqxcYOI//RirnLMFkOAie8IK+O/KwjXsryXVuEyGM6KluP4H/oysrXawLCzV+C
ShFPQrkiDyqYTM6V8IUIgF2mEQrSAYQYh+hgNyx+OFGCKCluAIKTtdd08HRdcBWq
mSe53KYFf8pX1GZokvkRzfGYnyWV7ab3NyAs9pKLR51CoywIwBTU2n644j9eWppz
7D9qJLCOCohMZYHLOdqWabjTXOwXq3IjvcmdCb5p/klGQhZ6/Co/SkKKdgqWqiAN
QcTpQDbJaQ5Nk9vvSOaQq1Wm16tuTNL4/j1DeYc2QvPDbVwsgdY4jcj4SaCA5oFR
uwR4/bMLNV7lG82GrjVEo2XiA7D0CcDo6vIBlN4OlNMFbWWIZYwdR1g3Qyd/zDk0
MHli5z/IRBQ13JtWUYDtpVbK5OG6pwAdcM9n36/gFRh2g1IHQlXYjaZ8UTx9Psl0
EN3tRhpPGBUd8imF92ABCqdpmQW9L5XmRdqlGx/ayca7rxOwXtH3eOczEs9KWbH7
ebYO0lIK/mbgw4ZlhmbQsglqCbpfNUEJU+lcS/cT1397XmBPV3mJh1bQxehahIMV
5Nlf0V9b4N7RT4/b+uFWmsi59+yOwvDqkmpBmcasd2F6j0HigpS5zuOhKVmXy6Cj
Tx3wUIzrssRawfGgdR0kVUlfPyfTsqedg6deaHSviXAs9bJa75hfqZrW4S0Im8Qd
IxXCnP9ksjSjOMWeiccA2jVTjtZIizB3GCotPhCcp+RY3XJuMBHd9xLjKJPRLdA2
qT4TdMnEediSu3Agz/tPmNYxMRIc6URACDV76bo4f1oMT2vS/h4uKtpfufUy8YdN
RT7aA0rww/LjzLu1LsWJ+mZnRXbXkPF//o+OKZadzoNwoYnoiYg5NyoWvyQ3ispX
8lg1ezarOKmV+EmSL+Fgw4MoJVmwRGtJXYt9KW3GpySuVhZI/aganbW5HqxJOjkY
ANrqkTVmV2r/oZiOwMSQVTDTndSUg5cP+/h5/MqjljV25nAygndaKnC+1Klp49+u
vEnDdpruqtQlk+Aidf/IwhfSDM+ydX17XB53qwaCd/whm1HDauZdnmmpuAD5GCIz
a0gLFOvDm4FwHdXTV/8F5PppV8bnn/7BKjf9UgKoVB7l1ghKg1mSvixRtp1olbt6
+ouvW46oDF9e4ABUEOt6eOYoyl6xnCt4BX9/caV1T25GvEXBNyFHFHout9ryujmd
WZ0M76niiBkU90Ihmv5oScSM21S+YMn+NbYB6RwwoR0yCGZvoapxSp8oXqv1/Ybo
u1d39HGAePipUJPCNCK9V5XP/MwaKxBJgtRCl3CcwhUgKY8WAvgHzNgOpwHtbP88
ZNi06J991+eE1L/Fm3EK7BjunrpyO+Hzi1STLzHdh53eo1I41KEvV07GpbeAO7re
xa6sn+jvsOuQs3RowClESF+l6rkbSnGBfmLnY2bq2fNtixNRLzVSWkwh/HXRt4IP
SEwo1YcqbsFcHueKiRsvJoDTgPILwjOr7Ni6JemEpSNaB3w3u/tptS6utV4TKbsB
Lp8ir7Q9hfNH93VL1PYbYrA7x5yYlWXdcXLUvu4FKENjQead6iMwiBEpfwlW8NW1
t2RxEjT1lC/Rvqwq/NJaWAGL2VOG29PekvZYhS10jsGqrJ8s6VGiY2/Vff6bIgI7
qFqYr51/jnINvDmDlGFQFJYzKl5ms2qGBndvUoIZLfAfktWa4Zc2QwrxOOeYLlXG
Q/z2Ty01voFi1M5R1Nqo6iWv4ktDiBVcctI5fvz+AjNix1lxmv5lRTT2dwNRXBr8
LBrukYKLPwXbUpbfJs+NrgtcGRqZs3Lo1jPaqpp0MDyohw7zu6FqOrF18Qw4/ArH
zKhsxr5ngIGVkxLTcKZ7AIy6Mxxv2VapQdyoa40R+577+b/V7A/mldvpwSF1d2Pd
g0bKSnWg9WLKhCslFrghXY3X8Cn2zQu6UGuGDngur4ZcILKGfgs6OJvTPMF7+Wu3
kjr81jar+f7JYPgNWxyyKinQ2BwuRI62yZADsj+KVoqHiUfwhgqxYqR8TzRZPqD1
hNVi3xqZjnVoHMAleq6wjWSMI8g0aQPnAjiQeK2LZUBkJr9v77JeawPTvFhDtMPy
7lMzOzqAOj5ROOaaZzh7IQVRztYluUKqeiHslaXoFdNj+kz09HkKNM93dFZLaU1k
KYwlYEliZXspZ09FBdvt8I5SkZX+A69XybDqLvSgBm5bTmVzRyBUdhi0gGRGQHcO
t4nXBHO/0YJ6wpgHsOpBBSNE06ZQad+Iy1xrwB444D2TGfWHifprdZPS8MxgJotT
QEFhvYn0YP/7CsVKNt2bZ7UTBehkh3YIAP7YcGPuwgublPwvm6TWBtCL55odp1Kf
lTclV7yY7TY1SlHsNquK4Se9pFT4nMRCrcFn1VJmVbs//7daVcD9zDK8F2VfhNq6
yQcJAhKWijfcD9OSXKJnPjurJurxeXDAmhNZgjy1Tdn3d/IumdLCfd5h+Gt26fsV
P4MHRZI99Xp8i2OHq5xci7wl+KwLG9AAqmwukwsmnDOUQEZXznqk7e1RybfSv1Dy
wG6yASEDXmiCd82DZLTL1myP7w7u2Ztk50UlQlGR8KDn2YazEG+waQPgFg8d3I+O
0aZ6yS5pbN/MUnSvKz/lXIEySsFixmjbhYjYrdgViRJt0GKN5roW1Uz/dH3nblrP
XAhKOpHYZYf3sanG/5PhdY2oi2t5lB7fl1pwvWqyyYE9Y8BM8qVSF8T0nQYQyhFi
AIcQGKsVG4xFZKXccv4L3PucOzcAQWjQSKcydRmbRBB3uPlLFGUEAU/VghwVc2QC
EP2ivVnv99iPUzxqSx9qI598WlLuS+E9gcVw97i97zhAsprlpqwJc9qU53Pu6ISu
qWpS/uujvNad37oeSwnQBqEEP2bfQNWD9SpECUQU1XQIyLhhyhqq8IqeZ5IrX2W6
bQkeZ3VDnJ+GGvoQDLfNJK0pz2uySnSpx0dBKkRsrzRvihMWgUPGlJtqseyPfsY6
D3GZO8BUp/4dcEJN0QSqCPo0eEypKnnmkWzQxPPFc858temDceOalQGqQKpi4tYb
AOOpXtyQ8l8ml/DllWWCSHgnlXqaxAKNTPmvGikbTTkCGDgLl5hMjkVxhTrYAaSB
+ksf/YCPSiofsw7C0vVW9v/T9mCEFfstneyVwqm/D91lGMlwx0g+1RwXZ29gck9R
IW/cV9EvTalWiQWXY+yhlFhaVHSaUz9PSq4AsfzDNJ/mCdvxrGP5hoPRIJBdGbrJ
3Q4myn3+ePvyVE8vxuJ7V0FLTI15sakYu4CLjAsQM3CKhUBU4QUtLwM8W0mnEGgE
ptD5MDSOQ+nlgRyU5z3ISQgDeiikfb755B7DeHk9OBq7vIgb0sSo5PDaAvqUqtdW
3am2NgLJkKMijgjx8E+9IPrcte/kADgAL5fwngJOLZ91xTOr3S8x1nmJj4Ejq3ix
aQbGE4Jtn3Euke7bnB7tkO860k6O17PhWYqh+qABUG3RmlAt8eRxEyW7Os3o3/M/
A9cSlsG4upfc5qCSS1diCFqS5hq2jNZR+kOjRaU8Fsi5+8G+M91tvuV22n7TRx9I
wstwKvS2w+Jr9HLCiLCcuommIBfQKyqWiWZK7rRU3Jqyws38YMxbIChYn7Nyaqvq
MMCDtRusAL/+lEvwTwPz/gT6mOLeYGjPA2zpDv0OpWCkC/y1taEcF4qnfBERENnm
gbVLR/oYbj5LqoWVUMogNlcUXVQTT4c4auxoVb8vyg3Pui8SXvAKbsoABexA4w2V
pe0zbT5lOYDUMMSQwwa+ADoC2PeEgYjkABltwx9DMU4MRrUsijq6jEL+nOk/8VGj
7wNekhJIJnplHucombEsiKRur6+w14MJsFgTdqkzKzQXYtl73+ljmuy7Rci0CODh
iFrYzTaRcgWznEE6J649/qRj7X+BSE4GWO9EipfmLS/luVCM6ILtY3QwkbZlHMPS
NxZe0nvoe1TJwKAYrz7qAOCEEer0I4hHJTzpjvsjiH+VAnMEJdoJlmkwSWD7UYbD
3zbyc8YLsGQRbDdvp8MqKxWHmAXECyjdwJLQJwy8Xjfc2HbWVNPM84ps+C3kOgh/
Rn0S8wv/CTJIMH5Id7SMPJ4lCGetXtyVan2vZLNh5oTYTVy3JcS5Y6i+Why2K1mi
g9mN1HlYdk1JMehfeSE7c49ROryij0Pu61CEDE+zIDGFm0YR3bJWZdITv/gb01Xn
wb3d9kx2Bfpgbmk1nQfIzb4XL6RyLOKH0GIL4BRwH1eG/lK7ccA0ocXWmXCz8KLm
Lh3fxpWiJQ65WYpFOIjnWqEcl9Oj1xxZWmhA4rfzDsDMwKzhLZ2k3ScVIF+Kj3iR
oW5QFhcWFsUhgpzN5ebN25tZyph7GuGpyDbL94PejPShI832lFCTSj+qC1bqRsSs
eABEXS014ktsn5aHxaJz+hX8SoMv3ISEhKKUBIbAaAI22bAlmnl6mitLFvCFQ8TP
ydVzwLcSY2vUiru9HgsYwYyHfp6oI9WOiiu5hi9GTJQ22jvKIE+DFnBrzhWjml4C
PV4IywiiCN03UhXgC38PJdTDZiEqC6urxvpdjDVbrdQJ8jvq05INCehyvzaObjfD
oqbM1ZEhkyi2plcty2H1+KW7yff7GYbLVtItPUI+xHNas2G3FBB2rB/NT2Y2tuy/
emXcYx9p4CDfS3DkhUtO075FMTGb/tbuNNlAagY9C54MS/fkIHohVLR3IudaINSj
GwnExm4Yaf7jUR7MCo45GCHPePx1moTt7i0SypLueMQ4ZC50/9f/RmUpR1rMRQrr
1WXDKogRKVumw2ecYLy4W2TF8vMciTNzxVl2mv28AhmEJSoMQKPgGEivAQdwdMZm
QKhc3PJmI+8pF7ACamZOCHOwi73Tj0nwlTiNaKZYeyglSyIXvPo/TVd8xjo3bo0f
fEfGv9kRCLO3AvUebRZZT4yLjGUVUnGeZ1TNIByDGlS0MY94JHFriH0yPQJTPeqT
HppJ156albmb0wjdVeeB+50O+KaHTSXtMFUKuTPw2eO7GeYrsRPKX27lf7mf+tXR
wc3aNsntAXmva1f/YSqMpPxjgqN3Dvm228u9psrCqM3MpaWnVSqvhKXfS2lwhSIh
IjR3vZ8Lf4RWgp+F13081+w8rlk05INajXTI3d2d2d/la8FuIFM8cP8RtmHZuYpm
aDSivvSqRtWx5tNCDNRRf1Udq4Dbxcvgp/y6rrysuQnhPF1nbcyYpYWtJxRMYPck
WGH7n03faB+rkQT0Y8KiYSNVvMstNKxxrZZmVEcR/Or2cSMzsB3MdVn1GzPe1MIw
BT1+CTlNaR67J7qLoXj79nIlcenPcI9SdJNee5ySt0MeyecIXpugoBrttau7ML/Z
o0S7NKJD7/xi74m/JE9EST38lyvh2M614ZbjDlCqf4vtQsRZ/O85KRehbDGRG6nd
ruL07NxaOR+WyeT5hb5LMfbrjzrDuacI3LhJHglunPherjcuDoY5LhHa65x+aj1t
CyEN41PNDuDy8ADrYZAgvjwEFNMEj2/TsQln8LqanbuhPWPKRJ8ACXKD1iqukv56
DlZluP5KLGiwGw0CztbrRuXYr+XEmmS4jLS7aQVWxc3NvHN0DEUFKTK5edJmnQ26
syHmaeEfVNFr3gZyqAZJFuFOkH1aDB5cnPxIrfqUvdRfn0Sv7+oN7yTbiZ/qsgKB
upnVLC0zoSR/QmfIDtHWwfLxWHi2FyEpszqkeQzCDNJfFWjBongcQxGbqUrtPfSr
okYf7Kt22IZswDVjNiuCQZScN8xUOQqBQZu0pFZLQZl1Tt0YuM29BOTNSQCbP1Da
IuwEmuNKiAHi3/w6Mmr09X1Ak9GwzTx5pYkxy3xYKfupjxNUSrTrLyn0rsQK2+X+
w1JFNMH/sNl7UBFZnlcLAygtaniXMGYhtz5QMTGH7dDiJOaV3ZpKrl1aDEziVmwD
utBsEzQLzl38dnRD8NdlYheqIP16brdtV5Cm4UiBguJOsO8D+UmTDcqreanijZYB
JdWXIJftcXEI8Ew/b+uPld4yX7tA8r+EtWoyvje0P733pK797bc3zDQbiu3uauRC
/4MRWLWwJ5KHdQPvbfd+fvSZMK3/5Jy8Y8ogLZ26gpC/cM8/jhst/FAcQ3cKTySs
gHkknXy3BEKSKx7rSWM6loKjUUQZDJ/O3yVeWNq6c2JUu4vTaGVNzT2kjpnPiMkp
b9Zm8H9Y1YQU+cVczdbS4e1QWRQg1Rb5K/9Kz9KW3JYtZBKorU/Y0/x36PD8/9CY
dKIQixovS3eInFh6fJm/PgI531eVDWsRbVXNh/wu8t9YATJmhqYs3swB5vFijsfx
RM4Bz1Tq8H1FckD3CKI3ZEYOGwKKg0AVkH//6rwIMb6U/IP3pAPpq/iGKDu+0IOv
9Sgr4Yw7mrNowxRfurl01A4ztEtRS7Z4ALORvzi9c586X9CJsBnB8MMDcPm62vP/
HzTcK8KkErSjacpObcRVTJSHaAwO+DrtR2ngjLjfKvtxpmDSwXMlHQ+eUPeBMpUX
tDvtiaLmw/DpH9YwUPS5yDwnec+O57ur1cXwTpKvGsNznVjnn7g3kfHky/ovhJTQ
sTUKakPDomrC4QoCA2/Z0UJsnuvJEC9a0/VfFqlRcG8z7E7g4J6rueuznjB8Ym6/
k40kkwxSaDS2Z5Jsz6s8WbHeXmDpFhRwRUksUOKKv7VAM3fBL1nLNnsRsnnTgRpz
jm14II/C8OgDHmtHqNyw1v1fMX/sScKLYb3XZPMljCGwQVk2F3t+JXNsw0etBkub
kaKVq30S+TvNjAA84zNtSftnyjPmOZax7gOJaz7KCQPaIpiOiYOXoDcyVMfDTzpl
yadyc4x42opjlnhY3V2WgbrIKyc5bqx8npNxoHkVgy8j27RnmsS8oQ0MEa1mxPK0
nf5B1wxhYIVGPwmuRdgvASwdQJI6TaruTfKYV0+vdcXi8NZoVPEy97KDOq/ue3Uv
TGKg7rlJjwumkU8ycRt6qhYWwonkbEBb63jRqE1/nXjcjQTx1WmZH4rPSmvEzTYg
ZrnJ5hCjKwTtJkaOkC7HBfE+YD/NqBMhSvQ1cADzoh6y/w8+zHzzTnEBZfMp57LY
WelHX2xY4iidwfD+yY3e2MNlBx+zpzh2r0tymV5BKiEu28D3sziMQw1knymhCsp3
vuaE83N+Bu2nBBazXZ50c0WHvFCIgnNyRIfimkUsYwubgJbp/YfVc7M/5MG+39yG
qAHYkeyLEE+L7LM1fHt0DkSnXxe413O+ue4BihrXEpvhn/xTVeo/em6sGadTd6JV
Xz0fo+0JpSxNhqkfxwEj8vrttGMHl1wXfeNUOY7WRujR3qo/Cnpyepn7Wn20uD0K
k+WlyzghCEyPAyJWe9MTLpNbs6yKMDVqDgUtdVh5d1Stlii79FCw+5EPBgrfM5QU
syO4PucB+P6w/cq36AP9YEbx5wZAeVO1DY2PsT7HBrFEM/lxAfeeH/B6QzWnc6p9
bqJsipvbZt9LRjEt9mRwJY4bCRtOkXR/Ogni3IBHtzTSdeQ0X0z3bGeE7X3UagXg
Mm8OyuMVYbPV4p0Zcl8BOMGLi4OSX8+iRPino7stNGvEztFIkyadtTBe9dMSEWqd
iOWkejCIONNsXSJIXZuVBLWTLZ7fT0S5Jp1v/qRaEVDXbYDRG3/VOlz07wrlpOkI
by4UuT2CgkDETDYDC7KEbzhvdCVddWbjMywqUydWpoLNpsMV/41mK4yO07MDEuLt
IKPOFW421maHVaBci+CH4B7f60DaLpQKyjy2/OjeGydMAPUSI8nea/hy/qWccjNB
WYR5tdMcaDrBsHaS3kACeyuuYjkc/CRVq5PwCM7jfOxBK2T6CR8U3dDJ7jGuJ2lS
bybzPE16rnkZEsmg2E1GXudLlsTvc5oXRp1K+ZgYqNdROgACzA1k0+c5VDFl4igN
nsbzF2NXmnr7GK745pxQ59L1sPP/l33XaKpgifXvHQEX+gMHsxR27kxdbos2aBIt
wusHPqGRNvwFcVX4nkawcaksn74c3YS7U012i8dXpgHjEiqVfVf6VkI86467NSTf
eH8EjrbQep5J0/OmRoZfzFCuY7ONVq2Mav4NI/dF34Q6/6mGjOPmDuU5K0isHwig
lAKY1pF1xkFCgQf6N5IFN/ihO+v06ue8DUv4FkD5zO4w12/rkecu7o9qQ34HuHNt
ap3qWlqMU+p2DKtBsFCGI83QG6nwkX9tmigp8Q7jfQ6fgjMq1ScLBhYHpXYAY5tw
Xd9RwNhbytLhRFdNTak9dpzTSM/1sphj5EnBSNNEjC0mExunDt2Lop8NqZivjDCh
SzY+annwsZnasXfHwyNbC3GpWAOZaUU5srC14om1gb0RpEUEbDHHfZXESDNHLdIW
HNJrvGVvPzZXb1Q2I0einNqBaVfQsl0u0QAqGabymkcxKeJEgRxyNnAobgnRD7ET
WenTK/Lwz8Zs7RyiECWz+ik7ZhGR9V3WMJOIgwZAzzFDySFNF9piJBZGHJKmUNt8
N50Uc3zlLYNl+2tx1XESG2Z4qPJgXJJB9Iii43N4MVJY3v4UXgK5OA3wQReg3XHW
+e19QL09u9lNfnOWj64ncVaWG5D1Usuk9WzWYf49NsiD2yXvmAb1U3Vod4MaaGah
iF9uXEKZ0NCWa9IFesk+kILjgHrICKPjb+Iponc8x3YyFZtFItP+jKH8h9oMv1TU
CTFWVuVW2fOzGXoJ67j+WGhzOamxYfJeEjZCZcfGu5LO7iLIPNeEwGsr/ZNB0Vw/
ipgHdE2vyBks9XxJJ3nBfni+fNaQmB04GW+8NKchVOvD9OcoC4/Uh/l7HlYVvQWb
O8qFZu/OWTlocYwQoPwudzafszL3C1Giv6snvmnH4w7dQQ5emJCqNxAkM+Lc+d/d
JiFnCrGZJbXrF6xa2I5qp5WcWzg6sMpjKxizV3HocIbOf+z3HDw++1W4ysxrtjNy
7XsvthlOg5VCzzL2UEKF2S3xLKgH1+Ocez6FIPuVGWpYLCU9dmZ3ia2imV3hFJEq
nFm5cOKYCeMjq2yuD8tAhlhTFmL0IipDMgs7qvsxpdvoqdUp4SiDgXuJi0YD4f99
ndcDu00u7PnrmSsB+u9G+uPu9hGvv2/+iAPe68ZoFI85OkoOfeMEqvitrYrRwbco
wk0rdL1/7ETaTXywb+Csp3HFg8Tum9XOZzLaq5s0DNid7JqZnhnTuV9B7TxVNfkw
DrbTy2nvzX9idaqUeB3O81D3R59D8u/dEAAN2r5ld00jILJ76COJbo9YJ5UZ7NG4
8qTYWt5jbJ6SYm1Ou9FtDUP4J9RkrluL2jMirzPIDHViIP1kCXccvz90O+Uop8hN
A/HllpvqsTBX6KE72HI8dLOl6tjiuPYfvDgfV2sBUy1F2N2P74BsmzAwG2mKnrNc
IQvzFu1xk+TGjoAdvZyEezrlsRkMuiYxyGsjWLqfqTwJxMkDZn8DT7mVUAaZB4lt
Fkgcc+E36avp+lmUCJad7DbrVtx67P9eBlgyaS5EYpdp0kuIjaBW8Bxs3hzOCtDa
JJr/cSnIa1HDDDC7BO0VGmvp3LSg0Djp+us92XdGQOb1lcWzkZhWqC+XD7HYfIM4
3DoSSUOCpMIgJSwsya8GjV/16CM6rEW0UAz5qmLXlJOUSC1arCIOrNr6EyEMh6Z0
m0zh9h4NFAG0djn6rF1VGFMt9TSKvjy+m49p6AkOCjDFJnMXB9S+XrgsX4Ez4ZXL
0tb6t+Xe1xvULvx4dywRttT8051Ap9mIFsWi12Rs/UZXwf04HCAQnlPdVMrbJma3
Vr/uxOZDzUw3SgUdpVPmOjvnRxgLfUk7inDji0AI6MDaN8St4HiY3tuVue+Y0GI1
NQMYJ3RqerL08kMOOO6EX73+mm1vr7YXtu8r5Q2sTha7EDJsgd9IySdpmiQfK5SE
MWTzbIpXtny9PTPA3JCGHaZsHew7JRpECceZWl55xB7+r+58HTKCYEhS1HdkS1f/
46GYrCodDwCeakX/EGJWm8EywdUm4Go96WEi4eNq/nbMXMGmz4kvP/bBkWfE46Hp
a2awVK4twH6j2z/uxSZa+x3G3yUl/gst6EmzpInRwE56DxTyR1/NltL/kiKVgvEg
d+XgYGkS42eIYyMCthS+IPV7kVLcOkedbjNW+ohXDLGcqrcbK6IJyuYepd84emCt
JZoLw9bAyNiNtmIF3IB6v5DGmCmRoKLc3VfPXQxSBMi3txpY0j9u2J0iaOEmLB7l
LAp/1SYsU+QhGi5cOjzg54ruhitgIQitSGJW+Lt3Chg4UNQ/jKqrAFYLg9wZvwOK
rUYFHARd4UBh9lI/jc1Ll6787NdA3dF+FUeh7+vaLv3vpHFuhjVVD8ffubcVK9XB
ucA2HgsJtkTVNbqLhSWrCCUECZzYXIYWz/XRPentXN6k2xJBNm/YPkAFu8bojh0C
3GJ4XjvRc8rnplKZAWHtNgeUFs/OWbvUgD7J8LP4RD/tpcUV+oQXsYOPJrqaUXqg
T5xOpLydoZ7Vdxcuk2k7Wav0HyByOBw2GyOAIcsy+eYxFeR4kA+UffjipgwMENHO
dVQOxBRNNY9oNzm0F5wzOkHcZlHMvXf4rZn0rSvnJVc+1O63WcJKuZjtoI+JDrp8
gWuLLhvumQ6DE9dtiG9FvmoPbdgVrMMFF1kRs3xABI6L5LLXJD2Bqc2OPRQFeksS
i0xcMb89fwrDyU5IGQdGnHoK8H65wE1w39v7FyomZjLm7l90lJUjlcaXAgikPize
t53HpTxHqOyvTnRaeu99QWrSS8Cy2hZe7qxHBLDpJ185dk/z7ruUNwfHN4dqR9pa
UMfo8ugzN3uGr0QjmYnD6U3smOVjaoVkFszNWw8nmSIHU3es97IgB0c1vOpWOiiW
D5ePpx1O2VNQgUMGhB4O3xpcdh0dW+gZYbJg3Y/VI7gMrU7rnFN7x0NcsKN8wuUb
trGf+yUQhhZrhLhQ3qHEf4yWJYBR44gkSJUnLLAJIp1zJerFCxxRY88XgIKhpvX6
aUwMqt03XKp+nDPq1WDz/mProhlPTilfZsj37H6CXlGhOTgpAQ6FJ2wBwwb0EC9+
nYBF05+UgIRiUGrZnL0TSxinvcdkTQV3A6SYQta6eH9q3plpjvYCy90EDe4ISakW
fqSiTpfUNOBjg/BRwXvwdb6x7aSDP71hFaudZelkvycDMtMmpRCFfwgi/1n5eL2W
za7YmUs65ZPUJka0oIpOvRU/38Hx5YJIp+6PWEgc4M+Pa1y4wLxmJrY654EQEf4O
vKFfHMsbspBo7R6xODPrA8r1LHzyofFALszWCnCjbKE+bFO5DXDJzEeJHhunn/7G
bbBtFChFyd4lAjw5RxjfBMCES1Cr00J+zq+s8SH+9sgA0eHAW5vFDwOOsirjYUG5
ReYR+Eo7otnmdkDuIL60/BMEwX4qE0LrtW5Ofh316BhQqwS/onBygWn1IEKGQhU7
GWIHEtx6T6u9FdVON10eFt9pf2PZEt/woXi2WwkZtHx3REWsJEKKFFnwdQhnKoP/
uok1WFGQ42402xbuGdkoomTYJIxeAOh45P1Nd+NnfFm+/gpVeNF9Wo/NsjrILPFB
jbNxjZ9fCo+KW1LW7GMFzIIsMwiAVFTKyGIJ59gC3P/xRg6czl16WfEoI+HQMf2K
2SpHeD/iXawmcUCBRo7gqpLdCA2lFWx2dGa3TEXI8HemI1WN+HDKSgy9BpTWVOrq
QuVcwMkrr7/5ZPXgq5Ko7LMPS3A2/MabPyY9sjrlcicGNepFoduB3Mxjs5tByS+t
t76Y/27wY/2/6sCxaxKjn9T2+LHtie1yB6uTlFZ+NxjQIeEQejVUm3y8HjvmsxGy
zcAHRk9l77ZYwkAz/xlyF84E6enUBik3lVaipeF8dy8qXeDw2YF9grUV9jBM/xzB
qmQu2cG1XNZf7yEHBvJEj39o591btPwxcA4ZC4uSR8f6PeVG7mw2DfOARaaYzCua
93LaBo6QLFDzbbChC2q7UiaP0+7TM4U2fDP3gwpJAQj7pszfYh2I+BEUpDChf6xg
N3jFeVn9yDcpCGO3axlx+IeIHEpSKjQiCSasbZmIblxJZk3NAsCITi8Oa4KGE3mA
vXXnLU1KT6uxL7+ot9hOhoSuwlXJTNREJhEiaNneAEJn/Li3IrDk174dUMpOmZh7
3hnEtUxLGRfmyjjKirRQwcxudHqFZ4bphhs/hRUdIK4/HW4xjuAhUrpVybvEENms
emG7c4A7+TmNIHKd3hWSV3uaAeLwYUgzU9arKL7q7n7akL+JfiANpDYZHPyZF7zo
hM9uGNcp3/RU9GpzyQxP7vag1tVbvnBFehMrdCSelhYCIdICYDfTHRmBIoEQsYWs
GOUqbO+62OyvKnWVX7wadNdG3EE1nEZchpeLqM6Y5Ws0ixoS/iKwBR/EDrpGN33N
/TtiPfpQiedYBPzxSek2SVdy26ZWayjUx7KrEsQscevBpPEeQUAq3Kczx3qoccHW
cdaY45MvMkOow6tQWfWR9tJ82k4oLkceJZcb7xe3iyp4zXQGYdnm5T41FM7E78SS
l57G/SgZvo9I3jBLBmqNT7BSjWu2+ZM7DorMTpMWr7HjDgDLplxSmtycOuaovW+U
RyfO66xsapMDhX/lL/5PF+VS/Q+Y+2JYUp9Fne4SVVdk5oZb4dWme63Vk1MFnp81
vnChVFtN9ZXubUi82SR6DGA7Kly9nwnabn7qfVxaW6JlZZg2VTIRGniZuH2LYSmw
icv2wxWf2rCJTDvcrr5WoBnCl+6C0v54iq0usqsn/Qw6GjHAZZLxEE7zF17BdrfH
to7+BDXCoitH7lG9kskNHEuwvigeKMHzuDyoVeWWOQBKvcCpCvmm7z3sT6/tkLmV
jCwl0CDITel4hJBBJshiQLqU0PAqVWQ5+VIbX0Elx/MPPcCtJ6WoG8OMV7PwKwdz
RggQhBj3w3LR0eb+1F1mb/KRn1RlKmwWwIHlSS4xhYJxowK5xwhy/ZRh8ZmLxxFK
59ld+DqObxjHzRzigKSqe1Tg8qwsBL9XK4C1bnapHa/rvzkBpgoWkbJZowFUKMT6
7hrn1G+qJg0MQwYPPTwoe4Z4SlTeM0NkmdYXWn5zrA1g1/IedSDNCAy8DtlpsmNR
MauamydVn0QLf10EmFEjpS3ArCtwas2U2go+WrRgCLcfjZRVImOUJra3alQiUfB7
F0ofIvbU7XwK0ReI8SfGAZEC9OzcNjoAJKmgRVyFcQkFmO3wJjU100V1o2a5a1Vq
7DIl35ldJ3yYW9XRbPqRXLBrDqKNULs5OKcSB4Z/vCGMs/t4s6UO7quZm4go6OJr
gM8TIpK+//W4QgWFhp4EUO33bvdS6Mpk9SYsufCvgp0HpIAYBAncVgUUbtqk5BZh
2+bvFdD+wY2MH3JW92MwEzpjFmRBBBJ3XwQ36sBVXME3JykMDjYsIt4cQOd0LCJi
TsHMx91GOldfqIsp5jbwvZwelKeN7yBFxnpVZgKpNx/bAtbBORW0QNrdmSDFFriY
1gbGo4cqukah9Rnd8+jjNk6I4yC8Drfd4H4O3SLS//zaZBr6iOL4ljMTT3Fdc9Xr
Wqj99RxMaHG8JiN+IfCos4nrKobW8WDKRkI2WTkV+8iiQCH1+M/VeDcYxFxxbsY3
wnPQjSPaXEycTUrijsIIWo571avqtDaqMhHJbe8kKoCRylN0d66sHMSMIcrpDtmn
fvxqulp2e5Whtb63nMKVi5WBXrmscead5HxJDZGyn47I5vFtkNYwREPFAILFA0Vn
HnE04gW3NvuZvEHSfTwIufVuGhyrJ4rDjaOANZjkXNth5LvgsmR8uqxfeWaDDg3w
9GHL8jbzDukP6bakewEz3XV2xGJ/BWlrUtF70rBgofuOggbxaRvHSHQFhh9xlMFS
7TcDwHNCzaaOZ8+eFry3VXlimX7FhulWHpsVLo1EHE8dEgmI7yxB6ERiB190aBdT
nCt7EXuOLLlGJyru6H/XWuMiBvt9uGJzW3+NVpYgi90qMR6nVVfGsjg7FxlzH73E
QBL2NmGO5JGDNt5GG9kkrLlhkqEIDY5HnoOrF+c0JIXRKpxnWC6WEK9rJPKlG+Ka
DjCjSzcrzMbPaHXLvzvzX/uC8EOl6yABdICbp8Sr57E4AzSzQhJ9lSkhVP5T2+V0
UnX1Ksbo3YsFf7TGiFTLaFDU2vo/OSFVoDoa/Jv/lU0oLoZWdZa8qy60ON93dYWa
5vO71wbwvOViCMb/JOtqgVKMDVo4JJ/AlvqVPG4kBqO5eAzWEZRc/XQVtX1If/7n
fHsB2ekGCQgZ2i7Ntm41t99g0yJBqRtLymi+7BqbxoiNg3WuFvzogvtcrNQmMUq7
PNXut5qhyhiXfFGVarlAIonbU12LaFvOl9jmU+4GoEKG9biPVhyuOe9Tvm4jkdHW
faZqfgaF2pPAsDBQ9Ddj2PJbfBV5gYtDvVnsoK5zc4cdqTgE3zNGvqXpHLO6j7gp
tTF1cvjHPCdVXfb+8ZiuKtbk+zPhl7V/JkD+Z+FOx7Sj+7X6mMdvYIWQgAHou3aO
7iNA4BVh6yPBYwEYueRWtz6x4doPqCF7+7alEgp74fjgNhNaPQoLgWPjVkhLhcV/
QXpJXUqjctvWqI6IdICMXfYD27AJTy4Hr8TyoT0GfZMb/NGYO1SmTxRZAkJEoPI6
2XoDp9Oj37UR1f8VVBhrFv+V+4xnrHK8H7O+IL8FnKrQXKXVH9N3u5zNdoWs/llw
h9CxCvQnk9WcsKbalQA6/3IXdD3RPyA1JGeOZ1EwxpDRSkkvRKP7gEhkViQYOmcT
LDyIwq76xm58fGIEkTChjwaStWL7YjJtNMpYu2dJl47/QRiTMFXkZ7QM9g+LiaOo
hGRaCJKC1synDnCp1IY6SLH3jPnfbp/QBGFBweBLWfPxNPg2EELEFWJ04ofo42EX
JmIhBMy22VbDopyBF+Y+tHwhnFaFDAAEcoIJqa4k5rZUOtZ8eGSwv5OcDUAg7wiH
DETQUgDdTv77GwH84GpAn/XBEkKNAYJGGdgN+XCA4MCeTQlt9yQC+Vy9lbhlGN3J
dZcBHYLxT2s1hrrp0s+y+9eKak5o0/xcu71GmPCDb25nUVuRhyIut6j/26wchjde
EkRLjyg/ek5pnqESJzb+W0XdZs381nc4jbfI9ekBe5OLJVCnXMBa0KhGLOjyIxLo
ZPfi9510wEo63a5yWlkG+b7VQLItUVQ8K6uAh8Sdo+IAPHH1ikKWuOu12E0Hs8lr
gKuSzoXJmQ2ALvj/FHOjioS+eTYFETBIKaNu1dt7fXkE/kmTrtQa1rcr/t6Y5Np0
y9MeVjOw/+1hCigUmOLiMUHTRyEulmxZPmI+qz0l/E60oKsjhuK1xjKgWbVTf+zr
W+C1/MOW2WuU+57mSVB8f0CmIYUXfrW9y2KWy267lP6Ara4WWmHquMz7WBTL6fJW
ijxFosj0ZdGMs1Pwl2+s80c+qu02u0liYP6fIvBzqoHPreuFuStBDx1wslmTW7Dl
2ly9M1ITPeP1dzgJy68th3ixCAdouEZARrxMZO2D0VE0gJ+enJY9GCfloH3D2eDO
ITLQw20xvkDMsKCmbXRecEBpmpuHFp/Nqx3py+MzljNsaYKNBPsDPSs+EIH8v/hR
FNisk/nB/9ZJd8/eRcfdmzq3OArMLHPDa/u56QPy7eimwb2KQpx6YPfXlOqTT45x
9v2TJy8lWUeCrfAE92IqRdDt7QZN4P++Y8nQ4jz0RGZawmiaBgos2v7SKFFJGKFL
gTk2ttt7/4RAn67aw21PSfmJSmsyxdhJW5pw8hviHug08MUZKUp1uZYq0ZMhO0Wr
wkZ4DgWW9jsje2jsy8ZSPgP5HbHLGkX3jocy/rEL6Yz52XlbAWbcxTipeCmusEtv
7f9HodOT30XunxDKqYW/GhQ7vcDU/A2mzGxk0UoDAlFBMxqq14+/k5vr3cZl2DWZ
lVHQQ9q8Doo85PbiliJ1md1/VDTYLjGKrriUsAxi3Dd9l8ujwAwgBPoXHHkCXNE/
5KrJleaPSgioNeC8kPdoQyT4tBT8S9YWAG0SB0bqaOpwWqYOA9ro8KKMqOxp72iQ
Ovvse/cHiHITcJ4BKt4w+riwD/Z27hMBbtU1RQz6M1MVWYJAQLllGuCYa6DnGSUj
4jx+6021DGw5CZ4AlJZrGL1qYT2seP1836tU9masp2wBPXyAQEIrhZG+BVt04SUv
ogFt+Y0sB6Si1L4QQu1M3HZRrQ5g1z1FjDtRtTkSuY4BnQuaKL/kJJkRMjWUT5IS
Tyy0W2/0Rx7w9PFcFnsGkx3bcvy2bfY0NciOs3jBQUhJav2YfBIQw0+i6SzUquJo
brd+YHymQPgkRissNLF50dStYgfMaPV8Fc0FV/FnPEwjN8lprmuvJsKM5r6KrPMT
qWd5lgm0Yttbdu6jj51d2e+YHHFfPZN1bTWX6ClspsSRh+lF9nU0p2ttezMaB+b/
UqniQdNrKyuVDTDNf08mGfAZHxC14w+v4MBZnwxqSRc6OY43K7MVovhy+4cdAw8O
Tl/CLZNcLEy4yF/47CFX+Td/41sD/6gow99WI3Yc9SunL2JGPCWY38JbVzbtGUSy
wCuKQdIr3uBiI/EpZW28jHNEPCFeA6KzfMDfgAJPq+PWfvc5KiNcIznsm3EIi/04
uhNSvsdQWN2p8X2JbkqaSxScJ58YKvAxfUqeDTcLYYuMisn2N2tLcQe1+j6Cy2hV
YB7xlCC8M3qPjGjwuuqHo1AvWLlyGxSn/yiUJSfx/Xyxlh4gHUTRJ6RxsmYhzaqG
PAbLiVrYm70ewDugbYBSdCJ7XMrePx8ofZ/TAaxKtwhbTMgHuofwxCNoJCtOG8lw
gnF4nHhpRtH4XE+jm9Vos6NjrCngayoItdLAmwwM82mR65hkpWVcyyzZhLvKfY3r
qujVAyvBWWMEZl8pFuEgd5ZBIUiYTxuiDX+LBpdPfG8KYKda0QUrQHfFQ251Y3i2
zKK/6cuDiF5Bwrgmsacu3sqV9QtHNgr/TKizlP5V0qrkdJAMZAZOcXle9ZeTS+LN
DUD+GRsz0EbuMSFjKnmY0hFPdkw2B4wHgyruA2XN5r4966U1Wa65U+JZodpVxFbt
YjjeWLwlgvPi2GXTuC8hTGiIDRSoP2sGP3zDeZFXw9tHvJeKm7+aBON1423w9sde
h17ZNyhEqjYDsPBw5Ytqb3kAjmelYvZktbABSxYaCWycS7NIMryYdp7mTLUElQ0o
PSnPGZKY22uJqLgv1aLW6S6Z6mJzN4L7gReoTSFqcBTsTBZY+rK+s4Yx0qZeZJA/
V+aOf97EE0gwT/UgsGyptmFiKDKdG0cm7AGwIiZck7hU2HfTCtYKCrrtys6tl9ry
3VN5MLedRS3+r1sQjCZrZ/fmF6LX7LOX3FN6IUHKuJRwnEXCDf4bKHpnuGNb38fZ
Fn4B0WQt2pLLzY1+1UJu5DtQycGCFsJ9o6u3ZqmsBykJlr++7u1iRj5mprjpM0G2
pdYSD9Y6cqMmb4tHdbcFlqMfyWjj56UTCEJ+A35ym9ZSQ9q+dpyj3J0xP8Om7wPe
91bUWbdjo4uTu4AzgyK4Iy3Jn+qG5imBmqnjoRObrXtJPNn3wHlJMQh3wl8RUOYu
hurvwMwVLG6m43VQA7dmVIGQJ9JDIsVnPQVjlZDUqoYjHAbdTj7vUHCdQq6GcEw/
nddDIcblDQizm7XZD/A6oReXlP6mhf6HqobBlXDP8asccwz/sAjjfJfw2I9aLbWY
drXMkkAP2ocK6lUvbgbH3RMV5gBg/lxGHee+U3/5qvDa58KVRqzBF9olcQ019TsG
uRMc0Xw2VUL/xt1Tug9qOFGXM2opPKh25pW1wjk7wpIsg3RYFdE8LaZHTFleNZpW
UrEsQbm3lKECHN+scU2gCX8brLMu/M5JNf3X7FEiPoAcKHY58Q+ZfQt5Rq4EInoA
tmoLOCE8chQfhgC/PcmZCTYvO2gaZUsWkqjdPhm2Ot+tnGULNV/hHmKHezK2rU+T
cne9gjBQ5fS2OJJ0aJM0pyWsZiRp25vyCJbTWE3z7gF1pqtuOqEW6zA5G2XBKIaH
2YLIMkBC0S4CBM4iMc1Nkz4u5RD3kmV9BDaErDXcdNeDIwMYAPDyL2Ybtl7tqQW4
PhhGydD7DjBzqrcczu4WNlI2Ic1reTkuQ+xCrWoDplz4719zppQvsF97kx5NYA/s
dMoZ/ad76jcLkmfhCdA7BeyeERCV9qLo3roUVJ4l52xTJfzGAZC/tUU8dEVhkpa8
MhfrbS1LpEQVZ952QVccYoKD6XzhUXdJKxC18LkOu+SB/f3SyLBA+zY6BRCK45N5
n7jAv1QcUcRRJsPn1xFcF2ckmH/xZGcSidO5bnK2Bs5uva93p+X13VOq8HWQhmWy
OQsIalk2Vy+uCnANHtVdgpQ6UqYwz2X6nqbKlijv44HRJzSuUTRuEbKW2U56eLvs
OAdw7ICWGkEeWbqGbhK/djm0ABJpqxA4fLwcEfS3ZA2w0stBci5ANnA47hehhKI3
N9eGn1u/ZtrjFjaQwfOsa2RmrvXvgk/v6OGlO5rdxasDSp6DL4MZk0zdWV3pxPC/
vrB92gWkiked0vn1JgJotahcRV3bu/NOx9fasyRd1d/i6+HQTwHPCgr5mcX0KROi
ylTPStFXJpjfk0FDW7zFu/wwHzvYPsdf7JA1mkyq/9DqOJ+g7RCN3iQPE4yg6dOO
LCiefB65ULor+7yrcdgri1RS6EAUEMZc/bTnvHVkKIJnQ1dFVb8+M5hCKh+HFzvo
W8cBuur9MdPlu2iTV90q61N3cCqJrIZBj8ZQ3MIO0BM9idN1HoGC/txtQuJP2L2p
OEFmCOyCcV/wbLFZuG7s0ttGaJGch0PqgQcG3FP5YeP4Z2TjGwWt1AitnRvC2bpo
Wggk2ZL199j4MyKlDeliZWoFUiCIoxChmzVrLS1dGxsmDmpZ1RpsRd2YRMyxLazv
Y91T9jEJOXt+CPgwAXMAcOLpl02i+uHMFM/v2Lqcu2pJ593G52IKRPyCQDaVFFeR
Lmz6mdHyRUVxN7jpkr/TM5IdbX20vSJMbw6DlMqpKIzvX2/4i8BCXiwGIdpCiHTM
+2TtvD7iG32qIexV/M+mmtDlxzxNfY0WRwwtWltbx4UZgXdF3EQo17n/mzRuNK3r
KQaTB+ylHYYgfQ9r8YtRPrxjZGyGKIg4M8M8TEwfGLfl0LF8QufowVdhbFRFb95a
kzu1xBu/VPd75QBsOYPvfgUOVOqjW+cbZvZU9MWGyA8XlxvhPCx/UPQbLZmn5tG4
ZNl7jlG42LS4GbjpHf+3O0YE8MksB7UlhzoyhLjg5QFjBE3DGDgY4nsKUH3bwUzZ
yCn6FYJwONl3CDiMHEgi0qUdwOYjWwmb0snPXBl0UYi/zvrS/neETSeMlr+OOc87
HFWlC7MIa5Ew9x9jD72FsHWHhpveeYt1OTBloaR9T2KRkiikU8lKHXSJ9llVFre1
iLFxJ5TWQ9ykd4sN06HI0H9SzRFHFqyYnUfRmOOSIK8GpvnfPlJ80PD9ajh1O35A
p284v+lySggYd8e36LeNaz9Iw33/+REHGerQK+F6msYCWjtCFjNMOM56Fi9HhDc5
EeEeLaIcvk8/MqcxEEMvSyyM2gyXmQnxzu7Pt8U+lReUgS/Z2UXynEgKPjmoIqmh
ZUrTwOv3q03hZHfr42wsBNZRA/dU0hZYMGi3t+dfmrd55oAbSxL9brWrwv3zHTbV
zA422MIehaMQPv9oAtgDorWRYSE41loN9kNxKeCer7Uw9QWerbQmZkcInyekPyMk
hHzIg1MZdCm5mgYMHljwyspHf/xQdH9hlDHWCDQUSv+oit3Xq2WyTHQYSy7jIE/P
mDDV6SQZd0GALLqM5TG3PmBWum6v4Tbx3xVLgFi2Qzy4IKEMln55CfXkHyrP1Tup
+sXEeo3hxnbwKTkY0UjR19kXsv3xE8zFpkCDPQehnoQeR57xWTVqVPl8zSrmgxrZ
VZHVgCEIkVtS3tG0EV9mmWR7fmfFNpxbtBD7w5R3MA/5h+wQZZxleJLWauXuGOqc
ZTw56QHQelSxAn6kO9IMOxuMDU+cDoXqgVsuKe2bGDzkxKHV6EpchWbs2dzI+ODU
cUD5IgSuTgJmJ9I/dFZaV1RHjIyUFRj/WL6ElpbODN4YzgfrIwLymADn6sKIsTd9
kHJJZZtq3t19LWjv0GW3ClGNh12GZNSUt/pYyduu9FJlHttVR46FfGNDmfyVYvdD
oTFrxrMuWPcY+krIXgOm8Lc/j9s3sOPiQjCQ57psidOjBCxzjvQuMd+e+Rtg+T/H
sLtnIpPf6+7Oa80j7UB2420k7y6M1lRiAz2Of3oSsR1gMEWYHsIC5s+ld1x8CLCL
FiapFvDJwNXpglNKCI12CMUWH4vWpVBkGHleaRBqZFHixkxMAZlIPmqufuPyPs/M
pwWxg8AixSp02/jioZl+XgOrhFyXRp4H6NkQQaSVfIXcSdldSCGvDmKqsoE7Jpme
tmylYlAt1+g2niO2RC2+cPVm8/fEga/P6/5d+7nWbt+RdKQd7ieXlvgQUa1FToZF
KaHjK6haXvFVtqsuaE9ygldb2L4nTn/aUWUsTeh5toWqjNqVe+WT6pUcLEFuHtxO
c1GVrzCB3YvfHiH3aSsBAd1M3dq2EwHpR+m1jQ/a+EoeBjNU5xG2E1kpWe7TJaS7
zlUaSXw2yIBMu7iI8srRlQM4jZr8P6AtWjpCli6dHqz5Zod8qrhCjRaQbo28g+Eq
9pVyf5GRgDLEZrSz2d05rxWVguBe7tBphxPk6dIxENbcvQQclkP58KNEzo8SXE4B
pGxZSPkgXI4wJV+uLJWpbJqksywQwb02Cz8E1jJD5rLlAPRcNVQnRaM5zsKAQApr
Mubag1mx7s59sMi5NIodmaGg1F5BVDR7oXAVJEG5K/fx1ZuA9kYg+7Jm9HMENVqL
BmLg6NSeMjB6GEugtHZlI3igIWhcR+sA81hmR0Y9lkSOSHHkQMG49aUhM4Moixcd
hNtPll575nCzDw7TvNd8c/ey4ndx+urxopSdXVE8u1dUdSPuVC4JsmQgHxAxJVK2
wWxAtSX6g/P6GY5x8NV6zVnrZ4K8HZeIdZ/Lx64kGI0uKqfk1CZILJ/uMUQX6XkK
x7WqR7glmkyhq/VYvTTRf5wQzoXOAml/bZxthBHETAuFtg8gUk9QQLAAn3al82p3
Noioc2XYvQjOO61dWY6vFaa1n8ojMde+Zha6eJuX8kR2CF3wPaOx6HyBr8hdhrow
9vJN9CMI4gQeJiNtddIqyFXz3PlnEgdGnF/Mj76o5UrZ58QBy7l3ZEpU5hQ1mnXY
7cqO27DQ8UDOyYZZ1HUH3W9WAJy3ySMYXeByw1euqLakukrd+JaYE4ll3MKCyy03
9ooxpYzob5xU27SjCMlZ8WmnqorGIJ8OOEax7zQG9sMix6MIKcfSQ2+X7iq/5cqm
yTn8APICMN35sMLYUC2nJy0A1LUAU99zlqX/G/fXya1sg9Xmde8llfB6aR3ai8aq
HRDqDbKIm4u9Ai2jkFZo+OdWfrRxjJGSnrgrjIPWA1YK6+Kg/qephhbO0/6GHm9w
LnblUKRLrtuNKguCfPkMqrAynzPn12U/iSCmlATTY3BSe2KLnVYoDbv3h0Nx6Jme
ywQEqE47oIcaiZ3Fr8M1N8uCjCWPtcYmvLseZmD17X22nuUcj5Dia4xMno1Rcc5p
yRInWHEZ/qe4DyU4O3CuiXXQ1n+PuXPEfxMROZ/ZW5CForx+6WWFso5tdM7DSlUt
KlJ046GJWtQ1V7uNibtJH95tu7fJadwpWeDpucdTB/3rVKl3EVIhvS7M7S4Fudef
RF1xsKVMihS0g3zSdzA5WSDH6mLxfYu7IrsuD3PtGr2Wt95dzfYvqaHnwFKdQ8Od
tOkNNis1stvNzx+QZobPl9bMPTUoFAjM+1mNkWwgj2/on7zabOM9zGoKiWJTMqBW
afl0bKl0nK3fcDI2Wfuf7xX4gjmG7L4gz+Yi+a4jbNwdSkr4t5SRDVgVyW9qh7BP
gMMtJ+LMvry7hTVKbLQzPCIFImvfh2l80HWSHV5Z85yUBEc37Os6HBKmoiH7qIbh
c/CSoeAVBcYZ/RqIfGrvMyx0iI7Q5xsBKQAoFxQLcXWROoH3krh16EO+A3kQMv7q
cY7AGsGqCSkeeU5y4SnkS6ZyJbWZYUaJNBxDS5o6vQ4hJ9FoGpIPw+RBRSCIaoUJ
wMhZapfXWpF6vPAAe2cLGEfVScYivSm+IjlhXRZNAIJGNhLySxFTDmCuI1dw4Uqj
HBXmdmTDDHlvWyWmCTiSVuWlA25FHqPUBaI+e5qKttL4W7vaOe8nX/atXjEBs4Ri
XJF9X1nDiK9jcNX+eER/W9RDocdPc5rdnYdjSg+6d1SxYmY4kmAzGRRa1YOe/DnQ
6gr11wuuvuSziJaoQ1yNxQp3VBTtP6tGupgJ6It72T/BmZt7HjohNGFp+zEXz3mg
aKw2cg96LfDeUwZCbSbiBOGBvSeZXEEozF8yw1kxvvV6KgVlPNGxP++p+Rq8AGQ9
UGc/cY2pSWeI9B+LIhPaRdYaTN7T2m+64tCwJexhoDyrqcDDt0aNBTLlqyeLJoH6
c/MN/tqytog7xGeLLdwk1UdtnodJrHnDyaEFbFzAF6Pk5hbLGyJxqrpLSLUGavca
jXWsFJAr5+TbkDiBIZtTgE4GNMVPRCK4AJ0KbVpZKUB/UHYILpxfTQtXVN5HB8YI
7YB5ZJNsmbuyvcsaqauFw2zoxou9UMlnybOkF1U4vSUP1llNcR5YdnTFoh2Wd6pJ
2tbelgoDPekz+CUi1CVXjJaPrmpnxjycnjEKMfnKtNxn+tdPMn9yM/dBofgXW1jo
PdSohUURmKYNoX50kvUQAn46mVP3W/s6I75bwiZm8zQslL+9RMGrxBUHXvWDoDoN
2ke3h8LmqezL71nhRusZgZbqbCaPOyhNKzZ0jsqao2tMylJFrw0xmgbKxjwOjIZq
EDssnTGj/kTdc5cr/XSUEgUjkCV1YvcnTK8T1xWcSy9NtXN5WO+C8+1T3nnOYpbD
c0re+pwpFPQ0TVwGskAmmkhTulq2TWZIf5B11MU7gioT/EQ7q+PX9xkaQKvq5fwm
P0xtY09J6qxJ5K2fEwyG/WeEPbuRfsmZt6+dtPuHgKfRBJNcHC9fUtHEVliIvvFb
CFLzlc4D1PDeaNXuBhnUiYFhJ1OORwUxvThDBflN23X7dax+js8DqjDwvPFnsUaA
lEW3lFbkaWaCexli5wOd81aLbexk8SDVMpoH1VnhdDEYzAyqPYA7Hd0CnOr1hHfm
OR5q/a/4i5mZ79PHCOldU6+W3s9jtJLZ7xVtMpGJM7iqBb4qTq/oMc/+7fWUAHJ0
ynx+R4uU5uaBmQZGg8AC0C2ym8dEkdAq4yjHMYzqYi3fuzQ6EDqrv30U4ozpNj6i
l4bHLsE21WwQg7jO8ojD3WXlWckcT7rfoupmJRr51BI6ZmLJiyFY0uQ9MarYVQsl
q+r8ue4ud/GIMHSZ8PWr2vuWL0+viVFruh6SeVaacrd4GtrLnxTvIUMfc+fYv+BE
lv80jlhT7vqSoC9f463kMEyQdOP9H5kXxMVHh2/nc0mX5Fd0DxUpqYmFWkFWse/c
p2WnLORQUqxksOYqTfcQfyFt5UnMwHe/3Wem5kSyvceZkdrErlIVhAnCaNq/JzEp
Tv5/tYaJ1OCytfJz+zVKiGOoZ5mWjo+i+Tc7QKGtYXptJY6n0i0c2i5wputLMYuJ
SxNG3AztDkl4RBZKQb3x7jzXBQXKexIkgwBr2MQfaQJUmJfvFh/ylnpzdHW03Bna
xq+mOJjBwU2V2jA2JJ8gZ66GvpYtQ34vxrH2RkvnFT8BvzPco2khL5TtGeVUMhRk
wyPPXjA0BxTFJTOgveywtHHnFq4Na5dakSv0y/gBGq1A4+L2cVrXCx0NH+I2gmI6
KoTNByvoSdxr/byRfM4YGNeZ/h8m+qGwbOOcR4r0udiuJvqhJ+l9KmfyB9kAdbkj
nzsQdiqjAhZYKbP+7ygxtbjkpUmvWk5AS7fhzXjAFDK+juP/mG3wPJT2bwR7Joet
r6+76+y575SxQ9FbuQ9hWDRpmpC+3greABjejvQjoJalGa+Jcj344tFDXRk0wNzo
rdkhW7GFBneI9EkYSXjDxq0gYsHapxDiIBl8GNrD0MgtRUwf5wWN9mNCKA4/LhiY
wKxUyhoJBUJZ8VHmudDGrLDtzHt5skHrS6kFRsrK6OQwvQ21MzPTQ3tVPBbmrJTv
y6VoMMGw78GGYdYv3uFeds3N1GFJunXNZTjiMzg6a9pVCE6GkBNg/EP+SAAoU1YI
NOrdUJOpXLdv2MhLo7lQpfzvS/DO/Rsuc943vOtvoG7Zb2eDrdb1BhZm2r6YUgKS
+vxjhIm6pAV2KuYfsdFYOclQeNRlVq759WDr4FSNi05JOa/7h3OYeJd20XqJ6cym
O+MWORWUVG3JHQRJmBExV3G5va/iu3hIsihxiwk5wweS5mUvynWt5dglAxHPGjhq
pjimjts9JSat4uEzRL03n/3qGigsIZXzToMTj1LryAEyo1BxCmKfz8C937YHbptt
o23Zv2WeTcb23yrq2+RR8BkZP/ixHgdiDbKi62zq+u1mLptwF1aTxpQK1fSMrN39
6WEuhM6RXk8FK2UGCglDMzTGdmtIoSyzeyWpMHJN7/SQBmC9E7BOIIK0GlKV6kfD
9hhl7zBOOHbVDpHF87pMTQEVhuAWtdJqR1MgzMR/CWkqkyZTNQSoWPa3w39oZcYk
f1qWSL6ZVq3qSmSreaOfYQs6ZR2yh36pxuWw1wOt5hDoHwUc6vOgGKSeptDh3GUT
UC29SkeU+xGlILQMm0gtUn/gE3OtJNbsp1Moc4jyM9wa9Yqn8KYy2smJm1IM/rIj
lv5QZn6hEsUIjrUl98AGBsVuE7Q0gkRgc23vFHV17nzG6xTHts8iq11O/CfQ+Qah
00NpndneFHjzeSnULKG3LQYEuDEfT5kfhSog7Zy0Ur336/bS5dyQPjX6eQrzUjdr
9WdtUrDkW6S+/2n4pz7Y9h1d8MXZbEYyLpGqfiZIKzZ/sHqwC35PDPpVf7Wyn3xS
AR5LTmFAGDEABaKMJBun4N5/NTDNrKC7zKtJIYZW8VLB+PR0MfRPcFxkqer8HXr2
ODtXzABWkTr8YFHaE06GTVQOiFgP4Cr8iO4OzOjZRxEH/PurSD3aC/JsyCpGFr7r
Ueap2yLn47ke8PLRjpM1HE07B0KJmSYzkyFSw3pXkYQUD7QdGTTxjm45VllAzGvz
3PrGiJvlfZGlJ8c4pdn8Ng7WV/ngf5kWloiYSor3hK+7o4UKeJmfD81KWs+6O5OB
zAsp0Egubt68v3V9MohBZNaMqZ6i16jgft/hdw+JbV35gllds/MY+/zbNO5BWVo4
v15EYW8apVpOIxIJqWBqNMoKb3nNTEeXXvXknnNfz6+P3MUIm5A4uYwnKMRfz1wx
rg8F6Qyo8/t6NR4wcVV/rlV+f9lnp2uMzBbLPqVfYl0GqO7yMhpnq2qarU8yNMEm
VURXE3GEC3exoAH8DOiXj3/5vnNVvT5vM1dz9Sm45YTalbBW/nX7oqdduPkvAkgT
l/N3mARBm4Bh+jYpcllE9PhvPhEe4DuOUSChORu3c7I+6HJk49e+PV/qi/xhoAKy
cfZSbdjSUEr1lpxRS/2YFvxHoiY1OzDbHB9jtRvRGvUiqw+GEKwgSDg+S5TFkxt+
IrEpfLQF6YDCnnI/kAY6ZSZ1klFiw8jQ/oWuYGFTUGQa/z4VqVj+//tpb88oSoQi
ruYe/kPoB/Fb+wf86VbZyu/6QG+7MdOkl4qM1n68bAAhnpYMn2Y++VBaH2BMk3N+
oTxbkAL+RkrX21JWt7u4qg79wr7zim4VUe0VR26NOnFUj/GFPBeJGTkwb4/od1mp
zCbJoThJJRj3PPhdJ81QgAtFiMOJQb6IWP/3/zrKSxNE9S6H6AfTLTAGdzoYdPBO
V4BWecpq5H//lddmMQ+pxRgV7+gdLNU3WbttdfPqyVybYZ5V/+uZwsvanoAsOupF
h6+l5vL4eGmoAeT2xG4d/Gc74gQ3GSJ3XwuSJPj5DbcJqkB6x4i9zQPaqwybvNmM
V/4PLe2T0w8apPd6suO7IQtAX5QcjIOrRl5MA1cKY3a1us4fw7Y20XlS3x/cgXQY
ulMGf/StsisXh7V/nM2rVL4FcQ3KjXf0V8GuHvEs0PCzDWZffY7ZMhSX4867vs5p
FJ8kRCZ0X8iacXw9qJu/Mkbg79MbmZYy5S+gpi3XKAU/xDfyalZ/wfByebrYYgbB
R4kCSIKhtBGNnniZlq1KyvnCCo6wX7GERZ7r8mN80OeL1hoFLYqoKrMGBNgR3VTi
5m1mllxxILBDSdy62YWvU2msaIZfZxnKq1H6mg+3I/f9iqie3m7nEeBDQo2AMPuM
qCnrdXU0bwyoAHip3Ma6N3FSSUh1x62QVkXeW0Q20T2nD+2e0FPfnUFTC2K55uyZ
Qn3yX+7k77mIUO8JGqCN7N00iUErxKJ89dxnZwzsBwzzlszA9t8nXm4yM9L9rlTG
24QDx3s5UwlYxB8179ZCHtN9Xcos1Cm1mHek7XnN12N2R/E8VJouACsX+qYjrd7i
aJsXJgqvxokmxrfT6V2DTX43proNGM9kfYhWDSLzeVMvW0R3EIrcZmk7tsWcvfeP
2BZLeJEfZO588zucWHJBi6LQnzvu8VqgLcbS2O4WFIHXIPA4a1rqtI07ZN4ZeIND
FP50gI1jJy98pqsm/DolbdAnKI1JnIPwG7rG4Q5QPgwc9+Fk781FdlRO7CWh3XIq
5/3ZVBfoYwkzR9IS2tsDqJZoO7dZfm6PuNgHlciDUQE=
`protect END_PROTECTED
