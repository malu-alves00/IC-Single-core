`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
goGzG1aDgLg27G0e8RdeWJjBbtfTaBXF/4C7Snicfh5ETE5MvCGa9RyOH9RrHry2
QLGQPEIJ4tn07ny24qaUhhwH26bAtPzv0TR+hmtyyMiVah4fuxVqwQIODIVCaoIF
uGd7QiJbkIhB/XmF5zW1+7Dq/ent0PwQEOblxtXtf0DCvUz47tpDun3u770RC7sg
kDo31T+DM+Gzfn3+tQHxU4p0tzhMf76Xwa0Fc9qo1c/92F7poIFd1/X+JFRMdLyV
3Huzlhu234LoeH8+pcTBCoymj37EppGDarfQdID+A4nZbf65iewWrGcO4K61zSYd
nrEmENbmE6bracpE7njFEyLfYvkpG9Aiz9x28KrhY+Be/i20ocblfTGfn91f3ZiN
I+JLS2zNQCQoLm0Q7xZxar8oy4nbNrB9mU8n5TDN02znMrxK2IO9d7I+T0WFW1qx
ufw+iS5P84QgaAIT1fuSIX5xUOpvngsrKShKO9+N4ZE4cg4TgG05p89h7CUHf/4i
uo/+buK5yi71teQ/8W+Yr+K8cn1GUuJVEpyCdGMNK6am8dT2bowmQzmdUqJvsqOl
BLSrpEi2RXHS+2WZIUmNqw==
`protect END_PROTECTED
