library verilog;
use verilog.vl_types.all;
entity arriav_hssi_pma_tx_buf is
    generic(
        enable_debug_info: string  := "false";
        channel_number  : integer := 0;
        avmm_group_channel_index: integer := 0;
        use_default_base_address: string  := "true";
        user_base_address: integer := 0;
        common_mode_driver_sel: string  := "volt_0p65v";
        driver_resolution_ctrl: string  := "disabled";
        fir_coeff_ctrl_sel: string  := "ram_ctl";
        local_ib_ctl    : string  := "ib_29ohm";
        lst             : string  := "atb_disabled";
        pre_emp_switching_ctrl_1st_post_tap: integer := 0;
        rx_det          : integer := 0;
        rx_det_pdb      : string  := "false";
        slew_rate_ctrl  : integer := 5;
        swing_boost     : string  := "not_boost";
        term_sel        : string  := "100 ohms";
        vcm_current_addl: string  := "vcm_current_1";
        vod_boost       : string  := "not_boost";
        vod_switching_ctrl_main_tap: integer := 10;
        local_ib_en     : string  := "no_local_ib";
        cml_en          : string  := "no_cml";
        tx_powerdown    : string  := "normal_tx_on"
    );
    port(
        avgvon          : in     vl_logic_vector(0 downto 0);
        avgvop          : in     vl_logic_vector(0 downto 0);
        datain          : in     vl_logic_vector(0 downto 0);
        icoeff          : in     vl_logic_vector(11 downto 0);
        rxdetclk        : in     vl_logic_vector(0 downto 0);
        txdetrx         : in     vl_logic_vector(0 downto 0);
        txelecidl       : in     vl_logic_vector(0 downto 0);
        vrlpbkn         : in     vl_logic_vector(0 downto 0);
        vrlpbkn1t       : in     vl_logic_vector(0 downto 0);
        vrlpbkp         : in     vl_logic_vector(0 downto 0);
        vrlpbkp1t       : in     vl_logic_vector(0 downto 0);
        compass         : out    vl_logic_vector(0 downto 0);
        dataout         : out    vl_logic_vector(0 downto 0);
        detecton        : out    vl_logic_vector(1 downto 0);
        fixedclkout     : out    vl_logic_vector(0 downto 0);
        nonuserfrompmaux: in     vl_logic_vector(0 downto 0);
        probepass       : out    vl_logic_vector(0 downto 0);
        rxdetectvalid   : out    vl_logic_vector(0 downto 0);
        rxfound         : out    vl_logic_vector(0 downto 0);
        avmmaddress     : in     vl_logic_vector(10 downto 0);
        avmmbyteen      : in     vl_logic_vector(1 downto 0);
        avmmclk         : in     vl_logic_vector(0 downto 0);
        avmmread        : in     vl_logic_vector(0 downto 0);
        avmmrstn        : in     vl_logic_vector(0 downto 0);
        avmmwrite       : in     vl_logic_vector(0 downto 0);
        avmmwritedata   : in     vl_logic_vector(15 downto 0);
        avmmreaddata    : out    vl_logic_vector(15 downto 0);
        blockselect     : out    vl_logic_vector(0 downto 0)
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of enable_debug_info : constant is 1;
    attribute mti_svvh_generic_type of channel_number : constant is 1;
    attribute mti_svvh_generic_type of avmm_group_channel_index : constant is 1;
    attribute mti_svvh_generic_type of use_default_base_address : constant is 1;
    attribute mti_svvh_generic_type of user_base_address : constant is 1;
    attribute mti_svvh_generic_type of common_mode_driver_sel : constant is 1;
    attribute mti_svvh_generic_type of driver_resolution_ctrl : constant is 1;
    attribute mti_svvh_generic_type of fir_coeff_ctrl_sel : constant is 1;
    attribute mti_svvh_generic_type of local_ib_ctl : constant is 1;
    attribute mti_svvh_generic_type of lst : constant is 1;
    attribute mti_svvh_generic_type of pre_emp_switching_ctrl_1st_post_tap : constant is 1;
    attribute mti_svvh_generic_type of rx_det : constant is 1;
    attribute mti_svvh_generic_type of rx_det_pdb : constant is 1;
    attribute mti_svvh_generic_type of slew_rate_ctrl : constant is 1;
    attribute mti_svvh_generic_type of swing_boost : constant is 1;
    attribute mti_svvh_generic_type of term_sel : constant is 1;
    attribute mti_svvh_generic_type of vcm_current_addl : constant is 1;
    attribute mti_svvh_generic_type of vod_boost : constant is 1;
    attribute mti_svvh_generic_type of vod_switching_ctrl_main_tap : constant is 1;
    attribute mti_svvh_generic_type of local_ib_en : constant is 1;
    attribute mti_svvh_generic_type of cml_en : constant is 1;
    attribute mti_svvh_generic_type of tx_powerdown : constant is 1;
end arriav_hssi_pma_tx_buf;
