`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EnqV/FXuNr3hoMOzY4HQdPcZgnlDH32mZPBgPZ8MGOpRVaFkKgkz+nExd8ifjicu
wv7UDZl7S0Yi/UMMP4AIn+y4kxnzxANN9DrMOgd0SrQSf6V8uD0+i8iQocFl5mN4
BuisvQozaYhsGcqehoRI157gdLO3WCtJeWe47QPprooL+RdUUC7D5tq/84H3ANUV
0XSe6T3WL6o8WBbAVbs7b23g7E2cokHAV4VsVrM2G1JUlaHbkRbr9eQrEtCNSPS/
BKLG5POys2+Z/BeKzPuQk+7s65EJ2TUrq0cBmSRGyhtZxnOD4nn2P5XoIx02m3VV
GpMFlGg0yH3/ND0XUZEzYKyXs4Ys6Rkhh5R+PmpA4toWwu3AoC1XQTNcB2dsAWVR
AmZoYJOlwo8HGjVLtK6rqmbGrt49mNn8+cTgigQrryoCcvzwGORLn0R+XaOElHpC
Bc6bAAtDyftaG59a/IlPIeclbhtKEm/ofvMpqsRq+z6ympNb6mGlz21RZx+iFD7p
nOVmfZ2ct20jQSjlZlq/p6ORyX6nuehr1YE1qXRPl9qTbFKfZZYxj9q1gU/HLCFN
GzHrB8HzvL1iTIl3rZm8xiRJ9u28KOgjtN8An3Z/1n+VAExJsPCLjYatFoiGSJCS
9DodznJrzTo0Z0XJy1tEBqk6Cfq5uprcP6K32o6SwjYvkDhDywRS4CuYHp1DJPoR
fvy6VAuzBa7ni5T2o8+pfOSiH7PPq20BZRy6HtfdxSpdvA5egOmfRsO2qIBe6Q3M
xoUEexfZONhdt6P8ZucxmpXpNfTxqtpuhAeo54g4MQLyX57NeW7HOk6Xt0cwenRx
0lF1nmMkVfcSZP4sWgcktqP3ay7a4MVxnctgT5h0oBEKg+8aMPRCOYyRkXDB2DmZ
oydB6jBlBx+2rmBDcc43Ygf6Dk/adSHmf0R+GTtO0hfoNMJq9x6+OvJvyRhcuY9b
bTk28eqQ8CEEVzIIAn3CSKbhjKmepYYQElpJ6uTe7JajlnUaoo+VRbidDv5T/xlF
DG1dtVyzANiU2m53/gThEhNzcNZfVfOVDNTF8GMeyyC/e6dJ+d9W2+80kQJ9bRtT
RniIc41SZv3UDZwukjhIfOmevYceEee35szYjbj7R2t0CBZWSdKn+SZEEORPX8xe
R+ESBL5LlwUkmf6veLeG7GxsuAwmNR9QiaE5vIWAu9f50rh+lid/euGwc3Z6JXCU
BJjBOiPNFUEIhzmBoF0bOYFanvXU2vl6IeSRALa5NbB+YWygtKuJ9Bq0PhZT01Sg
IAYTBTdMgxYsOTra4nv2QEsJPUJIkQZc/Gi0fdU+xLg/c2674JwPCL8TFnLTMM1c
1vhBoN01Z+tcFd5ROQgAclaX8d1KtmcUb8zHo0BiudV9lD1EmRytfm9WznefKbOO
MJ+qDvjN78v8bK0XniOczMS+b50sBjWtzULwDkndjRvGHaStm/xtLTVkC00gceEn
4UukJkIC081LqH18ycSA0HVpCoQz75E5QEGCdu6hB4IXksl4QXCeHjTWrrK2NBi7
IjEVIQ+ufwn5TlA7JLEWQIC8Rm4K2ZoAc4maIJxKILkePsNAspWW8L5LPOWoCzuQ
dXmpQY6wqIvn5MGAyFF9Md7U75PqPkMRVDZjQ976Sou+c6mZIaQf9u3aNpD5VOeb
`protect END_PROTECTED
