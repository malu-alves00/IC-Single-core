`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EpLJKftoUnBFmWgvagzokcSsaHVCdnv7U5dzuE8jm/UKA6jLFBXJF97CgggDqrfn
8d7TwM+1TUBbG4eSLGnLdNPbHv41kqpm2bCEUVn2+2IA5+ufEzyqLMn76QMefuKW
dxsDyF7uOb8nnpvApO0Sp8n1ULp3NehOs+86qW/dUi3WDic8SGCiKlDJ0mIs+ICs
6ku+HAEvG8Yk0tJHNBIEUjpk9Xu4HOm9LUIpsLqtQX4JgTRvmNjWHIyqNVcvIU4q
okkMHZ322v0z9GiUownl6wOGnkS8mpzmR9OwzPlW/WRxVIeQKuvib5mhuiExTiXy
ucdqJFaqXjC8s07CBiX0OiEjfIgyxmFo22wKEH9clwDvYR0vqZO6sJyv91cr+Ke5
dAElgWkO9wDU98kRuvJXsTnoLK5mogjWVCRnyf783bI49Uy0/JrP8aa15ToI7B9a
62ki9Q85wKU69e2qJe7oxpsNpuAeA2XT0wR/uhx1A438dDgDvYHZO781TCSGgJ1L
xibtp68qR3GtQ4AkcS2yvc8PXNPdzCYUrrOnSINcnIXlwevPD6g/R7ZdVotjJN8u
86sXdQabNIDxUc+OcL08T//eMIF5LmcYxgAp9TUrtvSWymnNdihRhz9K4dAB/BX0
4rN8sZr/PnqpV3soyrq4VNQG2DHHUReZx3JnwJvRHEWy9XBTqTrLPNDt03Kpo3ND
eNAvmjood1+cc1/rzMaqxP35Bko9hQaXc17/c67ie/va6quEPNuxzLoIZkYnhFq4
78971iL95/KVLUjGDqJgYjYTsCuKJZ+rOcXggct1vSRJGZS+wn4qyVDfv0OFaaIf
2UKVjJRBxSb8hdNKft0GwRSpAjAFq1m7PPbSUV64QgKB2KxJ6NDCqvWHp/wWVtlo
hkP85dp2gZGLRHDGCw9f75wEY+V4qVc7caS/x5qMTQHhxE7/xkHQnBPDkwtJLtXX
cwJWNNupkoCp6CmrWikmrbjfx3H8UgFORtK8vc9xy4z+kf4rcMAGed9V8V2fm75P
7etwEycD6xlPFBw4siF5CUf9e8cSTltM9f3syUfF+yHqRBHBH14VT6tLwCfSL+SD
iK7eSVnwTFkxWhUVuBySrRkwFbGAjBpGNjczZxWfHoXoTS1iVBYQ318s+fHPPWtJ
Ct9g9nWPte4T68hw+6vPDzTwoZNSdrYOI+iZ3ZWpRtM+LeJOiheLYK6eEP7hxrGI
XU1M/3d9GLIDWtJQasWzOZNRjSddopeiZ6pN/wDDgGPMtHvoWMan35RPbKagwqj8
gzyZzO1NKU1bzQzQYE6j+MB4PN/tklbZcD6JS+0h4aq6SFAC1Qo8BEj9tsbMDmeP
ekdY8/95NMMUHH31EHMfXWkrxM7FgIU9m9OidWBJeTQbWwEjraI2I/CJOeOyTpjX
R80+7UMJM/Hw5M/WRCp2g4BX5rXkrToaTFbzCDO88Y3qhdTPQf9dGZzwFlcTVcs2
V54hMvq0+nciK5wTIKoAdIHG1nXaS8h49dMWqeSOTAGHbYlPV2m/jOrsUnGBJRsg
TniANPbUM5R4uDgdjmqwSQKpQDjodBCRYjlpzvCo6Ue0Djkxs/leEAQwqm4Q0tHP
sO9V5eI4v+JgmkNjcDfzJABb4rJOhihxaMg4OUT4ZRsfuU9HO9a5IXIUGFvKeYPa
S+IzuNdDVkDRl66qyGJVwkeMbcHQHURK+3VxdhtLYsg5EuElWpGyr1G04zKAVbcW
u5JBAwPtUcJyIOgpXAc462NZKfu63pL9UmC8yVAZO4Y1xORuriXfEKGG0daz/X8C
s3M6qvWODq1Tq1m1MXz9HcYYNPGb1meX9dbJ4/nM77MT8NeBuGv0aJSlCzu3s3LW
gpK8SOmok/VBXosL8UDcZ8kAtobxdPa14ysHjmoY8Y8IlNupe1NHhL+9xCoo+tC4
pzIIMDiO7edS114w/fWRci+avEMqX91qW45j7uY1DDLQUXpoGnCu8FZVG6SEriAx
TcA4UGRAnAWazHc2o9aGExwBz70JpxJdPhhALaCAnC0biumNprd0mL9ebtSjEYKp
/wGCNSaqsSfjR8W4icmPrpEqoJiQBQRCcN9QUUcXmKDZLG1CuewRklpYauUMUPvJ
IAunyVNLyZSiMX23U/wGqSdO1sCt0Q7nrsCgrnd1BdjVcYilHGw+hBU7sEbGSre7
jBavQHMtAseADMzAtJ8y49CUWosGOFg6U5WutEjMs+FhQYwAe+V5zMdVQHYgc4Ay
yNU9Yu15zv8n94ZmqkX/hJLGnEZDY8Jl007p9K7x8ZqQeAY7BzLlBXXm6yH2C8uz
V41wCui9IcwX7Ubv04uedNT81LqLRH1qjtiAS2uebOMVfehA3txTr4L873cJmBhb
2m63JleAF40q8kgaJB+Q7d33WHG49C0+wF5XV+CA2ar8eg3Jzz+lTpHmThc8ooST
/r5883qARpAdKZxZe4XUkH/8k9WgXby/HxFhBQOXwKuX9kmiQvXx2YtuxEoaaAoR
oPSkcbxjrq7iWG/or1eaoI0zNXq+cz/lF9P6uVS90+PiPpE7dJqDSpwj4pEYEPys
3V7/EfBs3sqsTO2tjuGahSFjxrBQZgAbr3yO1KxrcxLm8K18EjnWJoke1rxQVnMt
3zbwgZkNcOCBZ5f0Rsp0xBhvImp4h0C4dig3ExXyA4n6B1oYBNmofUKWxwCPplon
+YN0OnbSMdzhNfCTZksjtRQblqf763kvbTkI4+NRK5rgQyQkSQBqeWeRysymzbIH
phWwNTuBm4HnjSQ1CBbyCFoQL6cG3JwsRsZyDOBWvjJF3xgg1E02QTofUvoc45e0
OnPi7bCUTGlzU/kK4+u0C04B/zPJbNiXrV/KeqpCn64j3kPOLRHgxp3mz+l7DSOu
8ndkJl6AaFWPHM2wrmRH20SWEpViPsWo8HZPa7kUZUYjeZ4O3StNitLmKMJrci/Q
g7P1xNQfIr7U4n/20WZO9ZP43fNRLxbwj1ZIRqJTP4r8RvZ+kRuzHd6M4XKOzdom
gms4hS70qlxh6M5XC/rJnntCYbTqpCGnolsoRrmCa3hM//zTx3HtElACeCebtJC1
XNQ9zmmeidW6R1dxnqYcvicdTaIIfMr7VICiQJbTUFB4CsqmUU9UYYjdOsWZ6YDO
XR8jBmbbhUUuSRK/QbaBQs2lE+KwGNrH1weS/ch7Yg/FuPdTaRI6gK2lySkiIw5r
35np2c1mzCMlyUKwdzRaiQ==
`protect END_PROTECTED
