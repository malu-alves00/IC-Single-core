`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vhDByMqxYtEbs1fua/OWsNV0lfFyk47m0O7UlMP4Uto0BI5vBL8rXjZAyIDwyXUj
gbbmM51NQbNfjhnbdgZMTqUs4f4zShfNhHcZ1dQIOdegngtG6Av1Hkj5YIXbxsAA
ZvHlGMsq9czUncms3CAArwJsHXeA4AlZ5d4F7PlmUn5NIcfJvEGovS5nmOwb7DIc
bdHWmBA1dv2n6hkyAy2/UkA144/FVsM1qfE3Pfm0kB5CrS0cNH3tmlWdYepF64ju
+Km61YegSHt5hFA/MKbHlySTRK2wtCpYN8VI/KNDjwMkmnnAghdcxpbvxp+tWj3s
z/QZxXxTfQfBAWHo67dvrY3GAb3B7IWlxmlW0l4rdVAFKWM99FmBd/pQzyVrwzE4
RUH+/fZO8GNMEaR5Ql0VDFHNd5wQ0sq1FYFpwaI++P8BIucFtjYV6aTqankUoeLM
oUve2V8/n6vxVHX9RnMJa3Y/NVM9JXl8yH5XtDLZlmRtkY0bB9sI2FpfA3hfPtvK
iRgMzD1MiYV35PH8IsEpRFpRxMUQcQ4sqhml1NSZDUMI5EEae/UaoVVzmwIa/cb0
F2kDdfTMvuBUq6eID7xnTuddnQlQdK/qMjhpG3z/DgZbgAqBwFPK6zr99mk7C4uN
no8/5TQs61ZWGDyTD6845gwpKeVxfjnm+SoWE+TDDKC13CfV5xjEFmLZupOn+Sif
pYx8ozoP3pFuARgoZl+wPCLQASbCK+17chbq77vMQxxtWOe2fBhYbNHn4JWjbWVE
kHzSkZgb6ZRafMHzQLN11NoXPX487OoH1mb8SpUQDzeRSVYmuK4S/kPp7axCoi7H
lQoPEx6a37xfoekbptFXXIWQP26b0PpMYWTQNKQSQhQZ1wRlQNtvXazIZvKoi9jZ
FSRSo9jCwdhdDtFiua/9NqCIWHPbw0DQRB9/zVGag1PQAeNbGDPktUgIXKDtI+3x
0v1a91XNyBSM99Je2lnLt5jq07B2wSq4hsmd8DtNJrgTZIYFCc1mqh22o8qNqlHf
S0ybv0gqXPIJrqDcCgPahS69paU0N8PK3ygGskQ/ScuqcUatFSRmnIabg4Z1v9WE
5YGegXky12hXYmSA/nrmc4vv1PLrhNonPTXxCGY6cN50H3azx8arVYyLiWtasA8Z
B9D0DH5T3zvIvbioHeaQ4w9W15jXyOQzSoOJnbr+1VG8C3tFq1dbiAr9f8y1V82g
`protect END_PROTECTED
