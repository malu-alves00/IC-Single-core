`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oZzwE0pjsKNjnNMb1wnjyqWvTCfqbQSdbDzZkiQ023t/rMlLyyjRP1aOoUYJ4oja
qy8XrS9IFJO7HCZ98yzVQ7japMeDWs16yF27QFqknOdS85FUvcBGo3+xm9SoK4cg
hq3GQjZzfbscFByhGww+yWbMsbjrUhmOT67oYvrgcH/4K/mwm1vxmQfAC/buSt3s
SHdjGIAlbdXnA/VGpTDS3ctiTvfAd3Ahw+vK1f1ntnIe1VbL5MrmS9sktM9vFxQI
0TMk5R/ciWLELjC0EbOlnPmdNT1fo/MzwlSGiZtxQFgvaIbnGHT+JEQc/XvHYIJn
BORaFNIsSnld7vvX/BzJaHZiLy0jjEWKXVgnsT5RbiOiykEl9kkQlXltX4FleYQv
2y/kNFOdcP2i+yd3WsPoLilYzeD5m+msZwzi6kuicKkL57YKDB2qU/fxty3r39+S
Og+KTp5TQyOGbegYUfXw+HmvCzxGTHXdi+95UAJWKsPNT9i93WsmYupt38GnCHwA
s1gnxHiWWYxkPGd5hyfGR10y6JBD4Ogu/buclYiA/U/eyr4C50Emsgc+UhCH48s8
36tQz2RqCRxnWeJxdpM+Y1rfekuyczffKnox1qYI3/mPoT3NbXZe+ZSybwhOSdsp
DAWYEwDoKiuTHXGr2g7/BjFEJ5rX/cnvgK81PEZWrINkMX7GwaOErpRnaDNLuOvZ
/Ue23uDUFtKvhUbRFt1WfMHC5cpS+XJRGFK/U7pwXxrljzUorrDd/LfGLvhU7HhV
SJS7/IKW3UMvuGC7k/LtIsFS/JdipDnK7TR2lkYbu5k0mxFL1w30s1gocMrGcJWq
FbGhTmEvbs/OBXXsnHM8aD1MOa6srxgyGkxxFfL5AYURPPgsIA/AVYLihFlYQ2sE
EnQn3VwXYZUnTveadSEB4Jh1XNg4M8TI8RCd7A8IowoLJC9bnkxuMChlDd5rKqtE
FkJ9Gwe49rStE61uFy9KyAKobkwhsCiXshS/J+U5zqzTQcGUwuHU2QmzjNtawAXd
1HMOYcdQKRjMv5yYzSsGdjaY/FvmumqGyY4cDPj5t13vUP4Cx9Tp16whL2fJ7AdS
vjeCvjr8XvE80OpNDtjG+tdsSkWEagdX7lacFS41zWyyJLZ6HRlcx5EMqj2zVedn
5Y3cm+w02rejDCNoE1A2TUf2dkQ2Ov+ieLyvBHU1CDS1qSovewTQw+OMP2R7p6wt
gW2qBpqvJ1Akwn+U22Q21x9InNQelpT9fST9Ad7BAi/1PMzpf6AZQ9GxVNKmYV81
NeR84AguxeOCsWRPmDSbB9+Vkug4wG2FE5TferNhrdzOplqHKgfFsC108kuTikl6
It+CpQM80VUAFMlgY8nqSFuG5i42qAYvaMseQRK9Ah3HleuIBPEKWfRKgDWFJ1Xb
qDJeSUtQ+J6jmoADK6TnkJUuPG2VHgJhbXwM4B4erSBjn9l9mM5MqNn6Dav9tYLz
V2pAOfguPg/4dwteuDR4BoG4sO59RZUph+tG8sb+/dcWtMsJ3IPGBNMj67D3Tjrv
ViJ9UxsaVucxZyKMQO0aoCO3Rzkf9hIUoAaVDPOniyoib5TXeCWLw0cI7Y5WgjSf
tf3fmEwP7lb8Wrc4/SAVIavsDv1XzAvX3jbgb0AIwK8XeTEEGlTrqxYaFvl0gOOR
ropdncBC+aIpEqSDaipvm4ufpUQTswcwj3Ar7hJWurYGkRbrjLh45IRcr5l/CSdA
w3qygrVQbP4n6UzAUEYO9tA/3iaB1KuDF9Wk94p9rXyvxNh5CfkaeZZ+4pUR0RAw
NOmrkdTdjk4QK0nomE9FPwsJiPIDgqLUXL5FoWxE8SvVO1NHeL/xD9+5WyEx2PPq
ytbYqXDdmsJtzyXuJz11pz1uOzJqyUN2/HGKZ9gMYvKaTZcevSTYWll1YDlzB8fP
GOrErBmQLkYJms7i3rxKtVhY5ZCZ/gNg80+R/5fEIgWwOHoHxUGjQlo10HtYpaYE
gBBlO45wu6y+d3aueQmXWSlcdJckfz3oRApXokE6GF2TXxzZfd8JmwKHf/ue1p3a
lD9lfEi7na4HLEsvC1UmyT4g8N0Slck4cIDF5mG9X4hIGk5KBDpcbPBdNbJzjhhJ
wzOSCYayatAJJCmkDoH3ye6sK1pV2SqQsmHSzpQXBHd29KFE06jAS1ydZVpPHfW+
K9WFoiovIIsJjPuCZborYKgo01pyV9MOwLGOE8k/dUrztsK2BNh3kgF3MJiqTrDN
k6a+lWtXo6E1Yd0kUabsRPKw+AKCu47aWwCuh3bw/hG2GoPElRFDs+PQK4w9pnjB
eTvHGuI4I3OPFxRJWphEjr/R93Ryom+yXFAD7jKlcaxEaCGzHMoLU8bahqNqSDKb
auMGvXNjKX4suBAXQRagySxfdyUK/J1LAp/LqV6wYU0H397YxQ8Xd5Uf1+RLfcNl
Q26olteo8V0V+Dd/YyovMThnWH5RxESV40V1ttcxC+wyDsGrO6ETGO554wBZhGJk
L39ct+8ed3dvDILm0rGgkUyn+DVQ3RBUHVepYfS03G6x/1W7MYlMs3f5AC4UvdAY
yvqlPfxhJ58QujZTXhmFfzHG8Ua7vbQ0lfKu3SI8zxzY4Lm+m4T4qi7ev3IwcHk9
1TLG5mPnF4/nN5s7QvLP9gFyjqRTxr0i/xrO7cXxZiyG4yjj3fKQfN+Nkwkfo1Xg
7a0UVVryeR2LbQR7T/d4TwhIoFqE8xdKCJ2Dyxqjtkr4/Wsa8Vg5P5nD7E0qclBm
CmchUcEd7apDdkvQGYNJXkfgBx7MHzhwP8nPnzgJS0TSMzWYHmcBocbF/FpyDM6r
HGDG5Y/c92UC3ojRY+5OfC3q0Cmd9hGefo0ywSN042uu4jnAtM1rqszrr3DV7NgZ
QlUfs8WXgdhGEJbPGRjJm/QTs6Jir6MUyh9KbuPFNWU5/nAUdQzxvMICtdVeRCx1
8frlYW8Kea3y+1DiqbzNaU2CLVJIIwUkk3puVEVmMRU3ldmi2m5OMcFz+U5IAcT2
z9icCM00pbUVXPF8fvwPZP4MM/UkhK/oMHwfIIQ3YU/35uhS2xNW2bpbnzX2p32h
7MgzPddBim1Bfm1wyRPURFi24EjNsHgNy77JUAmTozWryQReW8pcrd2ENgzKr4Y0
n1tlyDQIWuFIKRMxrmUwSuXXPvNjsp3mm6T7Std+cq9+CqmjW4dRd1D2d1l0gnFX
xcjNbo/5DnKcYWBE0e/sfyOQnew8Jn7RLWYbnIhN19kSPDJZUrlodsL3jwZGWI7h
ktpSyPTRIbHmo7SXT8MNIBdiuXyFLvOF6hwymK6kxw5fI67IvNzOUbcID1iHV24l
nn1/+rGaKzf8Rz7BNhN7rg5ZC4arJKKW9PreQMNJwL5fCYuPKyJyxzIIA9OIhk6h
9b7EsBbxk6ow7TM5CxS67nMf6OfDntg4nDxxz00VfyFC6UA2wcJEkUfpj+XcoRsi
7hsZ/Gc9gP+V3xhpS9nCFJkEWDv/vh3NmFayDgF9vby1/LGYsQL4ae0vW3a+Mxno
gV144Vkaml9wXZ4aaE6oj8bbLbS2H97ktbWRlWwKezDUeMwSaY3yjYBxiDloSUJ1
DBH12lhGjva6iuO2hulQHm6S2VonxcPlcric3EI2SUBoVtsnBC/uaFfUyn3fSOZp
u8FqeYabgba6Vynfr2IKWveQl+5ovW74ClgSZBjqQi1fnvFS0o8I0L758eelvqWy
1zr2eGloRUvj8c/FTixLobnnXJzNqm6sVh818MXdq8RtzpqzjvGCSopMMTlgn3vg
aNgxTGiKosHWfTXgj+xaEYJAVEbzP57KTVQ5YLnk2B74RPO2tu86tJ0gnZUAWNBg
lcDxw52O08VmgHh/59AwZizieAD9yqvTa3gdra7/NCBfjSqmLbyiL4xUAndkSgug
x9CZA2JI8tEZv7k+D84iCd2tu/0V8ZilepGstA7lc3o9MUBNO+C7VlEshN6+U7wb
yYikv3DDtfgTXz9TLb2+mxyi2ykk3Qdbx/G9eJk7yhTz+oXbE5wBCYwOVDSpISkj
5U/KCo4MXglTfoAPVWVN1UC5qce5QZNfsQfQzfqla6qxZDpSMGWJqJRaO72AwKQf
3zY5tjnndVu14Hy6YFRJ2oqngPZ8JC1ZrvMAJipc5LNYZSFiPEEyXZA67jtv+4sQ
Uyazmgxup7rtLrTg0bHKjNiSpc4JaRgDyfOPb3gnQH9IIXjhHPHVps7ejW0h042i
LoioJoCvYByGo3R0XacHK23Em2kMv7pPcg2OZZGpz5MTVP27pv316oWCk6P6Emrh
JEGOeCKXii1cm9/G3ZLnIieIEIT89hRSN2Is1leE6omKFVYJ/eL9W+Tt6SQVR1jW
6cOj/NIGGNWrXhKAa89nTBir6yV16jAIQ3EEDgygU3XMvpev9C5BGxRdemvEJWC9
INgWCyPqGl6aBcwdHQzvCxbjbF5l9SbapMn66awt6KzLXeEoOXjIRL8pKwSrIu8p
WLKw5RRmvDKaBjP6N/27GOwFzFShKdaWe3YH/Ac6DS7Q+WLUVDn8Qll0Qrg8AZoP
fEHtQWo4qv1IirU+cdZnTDfDGZJC0RuO7iKBjlkDsATfGaNNFBhjRNS+CO8EKzpn
T/oo65Y/Uk5zInwUoc7aOMo2nCDDXxwG/MM/efzHvnWoh4JlAM7Puc2cdODZcdyV
o0AiFvKZgZ32F5z9fOgu1mevBhrP3bGm2dvnBssHYXg8/xH9VH7yuTeElfyIWj9b
IsinTyse0sh0YX1k3KgFI0ffpcBRQ3pXC/MMwQaw+5yoAP3L9VvYa+cmeUOzSe+T
w8WZiPMjPlJnUYSzLuk/xnxvHXcm0Wthh0W/D86kfg3Iqay8nh8AW3pmnDyCnj0i
dXR9eE+5wm5m7FFOsZtkFPgMXxvQrB5fnYkYuTJG3CDK1YC0b0b+ykbzXWenYWKY
0+wUtCDFGHxoiH6ELkWesLHL95PuBbhN1t5GZLr1eS3c8s5PXAXku/dqqFxv7ha8
5V/Pw/36aMm4/GB4qZiY+ekq6Vw4xSgVUEysN1yCP8S9uel0GO3OWPWWBnV0fEtJ
aTq2xMsB7He2mBOT1knZZ4wraPWSCZCtabcZA3gsytiWk4fmen+UIZV8gEbAuwTT
lp6hhmAKeePwYoHBULjIWXhJVfq3xdhfvAI26WBeB2hZtBWxUx8xpww6drh2zWph
NDA+FMtGOoM2zvioI4k32iGxlB68JLR1RlKWccaU90NpnWecAiPoJkCpTurCzsoS
d3JH3pYK/it14E6efOfkrGpxjdQmEZO35TZhYXZE1HU16J9L319rB/jrCbf7LZ4Y
0ywyd74zozQQtoQEvkUadfhayZ/zyFtb8dSokmsXYZl+3ttALWtSqlgNtLFZfWMA
acLKFHLU6JawwurHoso2jXIKXubR4WConclInjTK/0Vw5L3lq7nmgojnLnJCe5Kh
caemPE07IazswZArhzGna2v2T27LHhQqQFq/BboD0aXD9u87q6lDXRN9lIR72tvI
cyn4NwIr49/YwewDqKd2Nj2P0s5oOrO5c9bSW5KZxid7Vp09QhsAf2XQ7RKxTClb
3lTQF7HtMTYA7Pn7YVn+BVYRb61rHFr/PSBjTnUo7br/OeLbKwCS/9s9tbeNUncZ
1I5FsDuIZqJzm3ZJKw1WhNxYO0oBbrW0tp+a+lXqJaObs/Be1ubqaVaVNJfpJqYp
dQRGo7Zgov2ampxNP3D1joR0CnLoTI9yv/l3vgZlTQikcJvya2jxXk/93X1Zj4W1
k0ljBekDTKb88FdvygeTUpPacV7aQ6oKCPrvV0HC5uu8oiuV2JOpFRVVTuLMCn7V
TxHGxO9CF1DhWyuWJph280G898mNeyGferoNhXa5F1hu9FWehMJs97eMdFN3XZjs
DhDka0bCGgvr8Agmy3XVKgNZLm78ZeqXFgZDwhQCxRnQGJX4zHsWD52LZHq3IW7O
mG8+9kGmsG4TMsiCV/YOSQlV6TpllSQXPC//I8zm8L2pkAwfaZ5bLnobhrso2SCv
+lsbH2/wvs0gSKxs2HYJLKnQDNnWPH/vM7uh2PLKff5X5RHsSBBYLXv6XhknSdv5
3tYYYdPGO3AI6tDGGyJAXaVrYEK0/jHCLPTKut2ZY/nw/5aup1qliJ3Wtpj+9Tho
MwIWwbzSvH0zMK1HQdTi0APJt2HwlhmFpAIBY87Al2FZuQ24j3H6F50PVAnVZO5i
kDmNP8tX86io5e9ZIYcMtkAVeYkE31gHniQbpN+9atX1bdR+G1nptHTtSOoqh52P
/mav6sDpOFcbDAQxpssOvD5+rN/cWUdR/OjUhswmy/Euq6MTaZJZJ/l0dEOHxWFC
eN0/LKRAFoBk8dryD+BFHo8wM4l/n4bebW6iIbuKt6aKdlckMHNL8PDN82u+redO
BZcGMoYQaKhLBsoYRDPk7iU9uEy3vXG4FBMi4dIiqfjPbcvAEf2rqbIZryxejQ1J
3COna4YCJE8oxCDTYxjC0tf5AeDR29R0EGuvgIMJ+dpO/3z3gL3neWW3Ojym5cgK
k5LmIWFcpP9XVZDjSx08+Ra2VDtc1NdDJBhX8zfo6EHUFWHAWAwKD+XnqjUAHYZf
2ULybenfYphyQcLDn+PftsPtb3NYbz2Fqdq5sL6uRM26yCHyheOWOq9mlCx/p5vd
oAqDIiE/ThtNe43hEQp+GTXg+BhHdMO2tWaBwOxRmPeKwXxQWMYy5mp3RZg839+R
UcHkUEE9cqrSol+Gzd3KeeCz5Oe1o2ovOyCw5EQkJRrhsy3AW2KmhVsPR+iPehdV
Xscc1QSoi6mm8zxavoIEK6gwUHX6ZY6ng2Y4bxMJmhKR6QS2BW43Kb66krcrfj7+
NhNDKd005lPA53qLtiTAd8u3pEMd7OogcrFO46EiLF4wDm6d6qKiJOtLRzCn3A4t
rhE9VpqyX0mFyRpgqUIqoFgAh4xEVBT1SrU9QecJvz8BJ09ACoILqGju9OKsCCwf
vOET3UonSwGBpBwS420mD0Zr+Me8HWTDffHymRfGd6KgYNu1wQ+ErCX2UJKgdWlb
nafpv7er7t5FE3/HfTEFq3lbKKC5aQtMAhwszKw/1d+fj9Imv/loWaSn2CzJBy0q
p0ZZvhf1WoF4DthgL6aCBge+SbpeyjXfRp4hyZO5ve2ZKram30waYpE7RgpHSSJe
4cB66HOvL092jBpuK6z4DfUb70CKgQrxHP+QpRSFRLlUQDnm58M1Lqll5DXzP7BY
VfGTaAZbpDXIJy57hmxw/gsFmuKwsTr6NxibdTGNnrpgQ1dhhwRoiVQBjKAD4HsM
+Hi1E+m4sAClN6Wi1RKe13QiBAR7xhuTu62LXpr4kBzauGAawuQkGAxxrqQatx4r
DxpyUeCtK1NxQ/4B745Om+8JtvulHIHYxD6N5xGR1oipSNIShKKzu8g7SpvFf32k
sWN79q0XfqX/ScrXhMHk1blWjCzNaELTLvx7zoQWHQsK2X4yGO3ek0LrnlTnNUZD
Pclm9/HJuTPMi6kV8DpHqc3znhCVRKJSkkFAtvzMEW735TEHpz4wu2bEsyX+cjOx
M20umT3J4blHbFQm9KcpwOV+EWkvMLPwwMyjmEEemndrUEolKXcoMhnnu5OoOObW
MyNH72+VwsFvy1dJKN127Ob7N/FPvr/sbp7xbUEZUve4adwO93CixG66NZfLL/+e
FM9z+B13tqz9nVTYKxLwdWIqFYZdUTAf1aKyGxaMDWur8Xdsjq7pPqLZaNhUUhi4
hQ3PdQMYsSXkoNf12Q/u7NgmwB5XYk1yP54CvSG+ndAYTvAoOWsKCZ0Ny4BO1k6a
VXGitx2tXe6ZuiDSTHqeLHDFAVyQrGwJNjPohv0W8qPLfBycu5ajH/NeabNkTT0U
M0xoT3skghORRpLKXL56eiVXF81SyJBxt/QK7xVUbLzqNU0wQLzYlKhvth4hlg8w
8HXv6TUDX58FI1Wa0F4cvRpZaUvN1RTZvUD49phDUWQRpbUE9kaNq3lCj9qYlHgJ
4fbYqwbayR3RlJfCPq1pyNMZK7uWSCD0BUFcoSG216M=
`protect END_PROTECTED
