`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ni5wKxrHdGn01ikd9MNjyb7mrzWm8H9JwzLWWu9TUuWYOKeP+0K+TYCnlqHUpKSr
FaSiZ5mRsa40JN8E3G0NwLMM0X2mxZYl5KFhSYmuTPG00mNJxm9fPkA6K7P+Q+wg
Ls52oH4kLyckrPeq//v5BiVNYJzkcGiaXmHNlVgBieL6qSWXuqBkN7f21Y4djQ45
xK4pTVPi8buPIsDaNEFaAxWOt9LDIK6QGo6rzifahwwyhbckzwu8SXlmgb0kGEY0
Gi/Ro1E1hMJsAIs/R3RUZYuok6DkR6FmoEZ+eDjy01dm0etSm6B11qb3fHznDrMj
mf/wCR6p/2ZpWethPHVGXsBLmdSx1B3RePl+AYdLRd328QXDQsWbi78tkVOhoYE5
6tyuAfc3VceMdJN8WrpQFsIptLkdocSUyGhYT4KqrTDCAXDU2gP7acldEVxnNF4L
FYSUqtP3Y/xb86wOC6Mz7ax9LEK+D4YZ5/x2vC4sbB2CvuN4Q+P/vfurBYlPkyb7
fs56lqhM/YL06C1gm85EZ8mtDWlXE05On6b/Sg3LArMIjZ6RzttWKURxcSkD/ZHo
NvS9QFI7Iiip429FT7TDGCMROeB25cxyt8y1EpJQVKC2EHjc2MYNok5/O0OYhKHK
mbhLZm6mkmetImZvqhsfFCsSIaaSUFb9iU+lbmBA3KmWV6EKGF21AVFYKMVZB/fQ
iXnu7cVOvemZSG2FovR6Gx/dO53Hr8cDyuIjuQwGD3MdmzWOS5wxRlEjN3d3ao2g
T778+gEBmelCtl44VEHqL/coqv2MVEnY/gxycOQabfhHou7/T6edw2KA5r4NncW7
uzPz0QzRjsXWHkuX+yazBQSY434tpTDDVY2wRKgKLfcRcq3zDtiAlSIDKoi/i980
MBZ3wCjhUxS8KIF21JkCqikiPJ5DL1LkKKoXdcytjbHhjHEv4tTXdtvETlKTN+L0
zLpTfj2CqbHQ/g34/xXYYYdxSH/VGTKyLEPw2jofg27WMg5SdXm9HtOUXnRt9Rpz
5pCz5fcN1KVEUcu3R5K6913Lx0zX4JMEjbWEPbDXWaEA0BF3CeYLNAPzsmHoFMu+
qLqew1T5Ol65HOMnDcHotaEoSVvhkbxhkuwmblRhVD3NfSchMv1xzAK4aXTxrDVk
XE0eqN7ajKTvX9YGFNvYgfgYx3JlzdFBerpvBIVZ/FIfrQ8fl7+fK4UgGNiceUZW
tqKLY5NEN/wuvQIGKOtUYsegZ6J+Wi55mCAPwfY1TdXJPfm+TrLB7mOYHqBiAAkv
Q6kLT0ubj/wD6Y/lw2FknFEc/U2WQzp3EbWROJ266Ts+UYG+d3sxjvhJNOxCdyAn
TZxqAYkARG+W+dRPvct9QF3oadZweptVKIycCu3pt8jHm3Xjl2eUZbokGCSTuVCw
RWZhoh1DRmUNsEx0kX9n23OCnYRkFKRD17RrH4km/iJupH/yYAatiycH8Drn3RL8
wysjmeUgiIB7t+VUKCRXjhJd/PcNkNw7te6yskAr4GE3NXbz+R9gyaDYtgw8DgOF
uy27m5PTG9ffQCNn/RdiBlUwSJi/dDX6ZLBB6JTt8BZcIYky7Hwai4C6XDWdAumH
x8UpgjuA1ik90YPeh1WNlQV+5yVc4Kg/iegRn5Wj7DC62xAItH9MWyEGHR1BjibJ
91DTiw8qTNRzXPJ7wgIfYEsMZzpvMjvZ7uRptlJM+2SrnYyImdOnmu4sJwiV8vZR
bMIvOq7cDdBjYp9d9fYwTy1yJtJqN/HrVby2SRKlkUBi1Ea79EXJMyqOeIzN3G4Y
zBf1nInpn/BZ6JflRuQRUN4rvTYr0Z8Ula0mbwxr+MLxVTHb98/1aOaMObaSUOyW
90GnVqUL+thEcJV7SKn7d/z8q6UHZCejcYHLeananVOSYowLlgFhdRdxBca0ZY5q
MaBVUBl7P8YX1q917pujBCA60tED1MzhHTHt1EbC+Rr5iGd8MYA9+U84Z/c/pKPg
4ektONni7Ub4h1toRkGnHy+2LPthnMYGJx/uoMakCBfhPWQtK6cn09F4ujV5T4dw
nke9XtAdJ81SFLHlMgU3s9GyrTsgkM37c7tcNinimTWVbswHv0BCwNkhw9DS9bSN
Jz5qufMIcO3nsDKHvhaTMG8EeUXmT0DPV1fZkS0qx7ml1NK98Q/sVCNShveYh4m/
6XPH6xxq9VggVuRQOUspg2Gnwo3CpPWkAWoHTXyU2h0UBX7fIhn0Gwnc7hg317D+
71MKBEHL4w4Z8fN+v04h7eIFfg3aqKevwR1WpF/a+nCUChzaZzofVAuzMWkSSSIb
Jqn29ZRNFDeWCirWK6eHurOAinkhU208mdrKsqHT7fToo4/co7oy2asMwjFUsCvC
Y0/ysuxn+0C46NZ/fHuUFF3+u5tqp27eLd/MlTlLqMI9/Ib31oJJdkskbbEPr5ov
Doku256jld3UijBMBW7xLTamlwhZYs3rBt3Uc8m4YLD6YxRpzSzZhL3rZy08Mufv
2YZZnzeQHgb4eVEGeemA4wvKXvSKIU7XHMfhzW56sl+h1ZkbCL5QrenbgEWrVgoL
phk3GSTfmIfV33U5vJob9WJZ2OFvBq5lgpBCbRprpbDd271PheWRTvO5JxEef4Dl
begJCTGqA1zyQt8D4qwW7oB9qkQ5Y0vcPN6L+OqxInQsXQG1QKanyuuSNY1DaQIX
4b7scEKHWDgKZ/eNlC73GUVDT7efBx3VZC7F0q+PZMRpv2uWzQl7kLMfa4fWZChn
vyBCSgOWFHDjCjrVxZ1Ampib9/nJGcnIEIlM50+XMbEOFaf9JVR5KvyfJNW/zucZ
32oJBfobrMWdEn6eVY2IeZ4N94bE6Kt0RHfhV78rl8zg2x5uadq8HMpb3SW13zNf
zQqFByZQHTLcChJoeh0Gv0HgKinr74QiVE0mO3cWiwNohMvXg5k4fY7ru06+aW0n
nRE6J5nCOH9rcqxhB6NkkiEe+jHaQvKr3dZMGfKgLtopj514N5/9OoS2t/LwawSb
V7w7ydymnW95Y6WS2kyPinOmShFAlJetz9MFzfY/4gzTAcIRAa2Dwr9GdnNofsVf
/PwGiJ3yJSr4CfsV1z6kTpPJkxWPYILifdsg5MmAafb+OGgDpoCazJqvjxnfOBeJ
QEi6up4ernAfw4ItaHKWk8Gzuh9tMZyaNC7wUAw7g+rog+LfsuIV7I5KE8XKRciV
KdruruSqAMR3wmrqtX4IXLRSiEHPJ/6zfyO78YNZeqQMWaJCeTm/AGWGqApcT9S6
cy7OywYxW0kywExTSRrMKxmtQMT8+wAhj1cdzR10YFKxDOsmNke6VxEDjmKweTYw
TlrqGTGoZUMjaeP0zN1FtLn3PiT0UTKcG2jbJuLG027d7cgCuchRVKMJCEckSIe3
pITt97ufqBh8Bmgw3hj/544XuCG5B2OSpNzUcDGeFde3s+acIaFcOq3wpaV5FBOb
HxYOiGJBwsZRftXx2Lqu6mmr0MaZg0lBuwcLC3hK+mgnRhdIJ6h+qhg5pv1nvPrD
E1gm+q+5m6JrucQ0jmTaJzZoEHDJarBu+H3LHSeqVlkw/YQsRpTJjAkvebMNe63i
OYoZKRBui0kgIJr1N9zMJQH+5w1AM2Dg8V2t+SgzpJw1oP91SnRvmh6OXC+i49we
tfQAISu9lxZ7hL7YOvesAWQFtIREDPRInLz8dUW3nGnl3ykv4//WVauNAHxp9WMZ
bXBpdR35LrXaTML9tzwKb9FwzmTjioQOHYIDnRsB611+0WrjyaEl01OMSr6jTRf7
tVNMQNahM8yl2OdEGyltDahEVhWCB8f57dltGkVh0fDF5fmQsoJRqaFCsVDNe2G+
swliJ3Z3SCi3w3csbSQXWSmL07fj227w0Z7WCNuxFjNefKmf4v97D1QnjTO6LsVO
bYsuu0Y91X41kKlW4i1MkTVx+fWkyHe3MRsGeae24A3PYyCRJHt5mAXoJeZQ7yXc
kqBBg3L7iJu1FkS2jMzJPrT7CLeli/hNu1qvtjcat+KRzKkYhc7zEmlgyX6pkdIs
mAe4QIsY7cGIHUNrABJbz+3d5Feu2PpFnfewq57i9+/TBk2XKNW47B7XiiqhsZU8
WCDh/3raWRCrhRLEiysai2DHJIAetwiSXqaqB1cWOEPVFFO3IqiF8kcJEO4Uvjgx
YoqwCLjiwt+joMyUJIPEDvmX0p6ND1apOBxzONnKNcUNXloSg/dKtJD6tjC3OZhl
V5iUEPZuzUo/kpWoaL5E+KvjmAkUifz8zYS3spJA0S+w+DrnFwpcQ/fwFmNsVzv/
FRMiNycleea2Af0sdACYWNystHyCCt4I7+JTMj/k3SYjKD8jqzuacMRyctDVcvbX
4gKvYSzdQAYclpiIQM3QJ1rb36LYxyQjytzBME2cEJPzKO5ilLUBpKQ0Ewrf39fz
l85nV7RJBqAY0/+7O0P+FOcufW8LmlQyIjfEtaN0MhCwHcQD3iUEJ1BAtRZ1POsI
2lgiQmexrFtZAJBqlepNKIeRKZQf/Lo2f/61MuJ0zva3YX0gGSx5NOhV/aAU9CAP
s1VGe7AuW5nY5dxcu4Da0JMCbgLkjKTC0I9K1COWgVburdjQyER6z9XbQLirHsVv
5GZY1qq3yqd/+oHliF1HXwJDt9KLLdr6oJPnGNZo+4iGpj/60GaNavCug7jB9S2m
kPC71fWi/mQ9NR6+wjZWQfKHq9Agbx/3CBx8mCRTHhuZWjG36HxfS/k5d5r5Lf2A
mdCuej8t6m5I0W//O40lKskUwu2DEznxhjDicmkN7F9X+5mn4CsaXlN1GgZ7Mwsx
3QNBK+5v7Iy4QnDi9z8JY8WRtv8t1wEfKng4gIb4b3oSod0k2TMogL03/3a97YG/
DLknsJNGRYbpzP0vQ8Gu2WSFBNvJcY5/uhcTt8FddveNSWdNFZYW1Ad6RuwmYyUM
u4A8APh3ulebwdy00T1VZ1J887oyKG0JeAeJwgRSSomJb7QTeucRADNTkoBFTM/q
jDip2mqFo4PAqS3rn5Lmzl8z05sgDfQLqDIDv0Z1m4xm+CpXJFHogDwx4E+QGB7y
PjaeQyD7J3dclavkslnyR0An9sJE6uNSOhshBpuaeZo8ykZuKxh36oRipu8aioUo
T2QzOnopFjuimgsIkQ4E2fpyaDMyJ5nRejyYMqvMwVeVTIULB4mOKInFA40d4z/4
l7NqJMwIEpyCTSihgWDi92ocPIcKwWzYaOOWRu8x7xPy2ob49h2FzKVd3d/WV249
V1J3MYoajEy8I4/G25N/6qIGZdS8oIZKXRBlxSh8AlzAffNnYtrachvZJmf7h57u
Q7ZQ+xUki2I6LhpNLG7qxfkETxgm5/DyVR6juv3OpCBKCM6/OyqfsJfX+pUKSaJI
og3oTis83wLQp1q9pUjJKC0Ctf6bkQ5d4fv5pSwUPJFUMztcZmpTJaxOp1WmDjXC
nNr2aOZHaGKDYgxls8wqECc++USJjvJDTL3+srx6nAChfBTIyLs6FufsBZB6IIbb
gSt63XaIDI2PR9ocHWar8rgagqxYsiec65ITn7P+dTgqbiHJXhUYxxUHzQ1NdN8t
RPA716WU3nY5FsuN2Cbfx+39HLMbKuF/gKoNilRv/X43WVD1s1fwwIJtVZcOLOLg
lkvTH2I8AynQUEUi68vx/BvW6G5/ja6MRLdGMTNsHAPQ/+yYJVqECiNVpmyqeYxN
o6kCJXS7K0uXVydXe94wNylCl3pNuk2GtGBn6TG1vmsk3to3y3ej2QiOm342rR6m
NAs7LxzV2DzsDOFrCjpTT71gJ/uDqdcIqp58ncI9W9nAn/4PUc7EtXILMp4LjSRP
fJJjwZbMfED3AEQWUB9NX5ckRd6EH2Slb1W6u5sB5qZwccbxv6DJFBu3yEwEUX6R
xEFBjX/5UylrlPZSE/AonFOJmcrjZdWFGdHHYRQQ4dCUFVr879mY2DAD76yJLiSl
nc/AMO9iEgSBwsJB0QBgMITsO1IevHsPVtWLX9aFKXNgCGbRXfjRwZsVeeL0wvJe
HbS3kVOLE1vVQIvxu8+shTuL97VV75GclK0F7nzxt3Qm3F2XujiHG7ojB3NV8tl+
WinlxoL88MmOq+JMQ+Hw37plka5sUR8hBK0m0MaYzDqyc42s5208y5rqsndwTQut
hpn9fu2loJnmdadoIYXxFI4LZuqTAqceJiIJhKRdqG+LdPwotpuyb5u5lh58G1Jw
L4kD8qFFORLyFhTULKHmqyUNQBls6oPF/hJw5XApbNeBCkH+OOjQNfxPwHM9g+5+
beLS70QxtbEfr3I2f/AQ/eSVOgN2KlZApJhBwRBIJTsYGcvg737M4N1NMZK5ribo
euulnvuA6rBOx2JPTfQHMDpHoJUYNFaLzdQ3S2qA64Ge3AcZ9tHJM6CUXm8uyVm/
SGegQ601TDRpP/FVJK40g09J41Vp2QnIiO3C49CTmTcSSuSfATV16bgwg1YO4uNv
cX/rdDooJZckTh85vlvc+A0DoTzHZqEbx1uuY6yRiBYls3zArI6tn9QbBHarr0Ek
SmhqaJvjXx9sjwnj95TkZl1+Y0NV3ZBYDxRYtt62dw757+XaA4pnDY9+/xSM6ZDl
9SvCsergGKRjF8puaIyCFSvyJBj2ZNVI2LeOF1k6OOrreMsAqlnvXv10D0h06Im3
62vxOC5oVJztrZp9BFAHe5lT2oWQl/Tc+UAQaqZtvKpUeB4VDg2cAttiQouruvlp
i0RNlGG9mWJnRIkh/IrnfBv/hGOBrKfEjI3wL326EV2EfngCj1wp8XRNtcbaBc5H
kIM1iCsb5A952VUFmrK3JeDvKHlVuzztTHP5atWtYnDcYRO+HGXulh/mV6RM3W4Y
1guD69pm/hFFIBJI0+MEgOOakelFi0n+P/YI9ykchfAAro2bQznNg57TkPLKPhah
I+Ek4k/ILpx3FgTR9kUzxm9Pl6OO8zof5GKC8SR+3i7Asm17MXX6Ly7fXkWtewdP
29k5YBopcoBW1kdy2mNHHqrpuzK3VkLeRFnWH9rdwu2RNHF+mgdJ0rzD2a310aA6
1CBOxvXCa6Upw2oWr9TvXv6Dv4V7Jly9RrCE7+D+r31LsIzf4d3QK7crsJwqJxn5
HrK49GK/yUBOe1bN9uwPsp3V8TWtGvH8EvQnPHN1GV6MRuO/wDjJHySnEy+ptdJe
BqtzxxnrStYpoea7qP4bGvJ7yzhO2AzKXvfoAen756BmvSfTSb8MvBZ6FXkw0yAr
J7fuuRBEuEer8Py7wpK3aeF+iUO6rEA+kJWejJrVzsaeG8mU/cNOP8JG0e3wd3LH
eifmVdGKIhf5NCPlzT1p69rljZGW/0SIxaw84oKEwOjTx2KqOVK1hJAVZFBwBgSR
cew9HEKBcPSMxw5OMNNfqT22P1vMtRWJWGx2+/AF0NSl4Dr67T6wQ017VgARrhkI
NRb6sHW272rjEjkqnxVYQQVZoqKaGZ3yT2o8UUJrI74ZARy+XQMQmeOxutXv9VfP
PoJb+WTgSV7R51oz797n4d4HMA13PsdGCZKwWwGmYtYZtiK3L/kjncPxLwvLMGEo
IZCYE8KZKpn0ISUg2iKBGX8DmOIL3cz1gpYiR5SZee8fNKhcKvoIqH7+Fc6/k2BU
3P7oBnrdiiwNWkl+q9xQrM7RY7XM8YHv1arIWxlfrWEYrV/LQMy82TPdGZNmvLor
t8I0B4osstsuSP/i9zegFK3awxQ2vtwJ1Mxi2p0XLY1IWt8Iv0Y/+PCTooP873Fl
lR12i+AfVRh9/bJclLymwQJ5b/djI8B7kR1ZwpO556m55X4ZliO/9SGDa4Cb74+i
ZKmnj+xBLuDhApj06g3zs3RZdlpRyWbVUGiSZxfmZveljniUHFj9d+8aFccby1Wb
5aids5N1a6eF4KSjFsITomBBl63JDkGF0H4xqdAQgkP7hxPzr8FN34GYiUBYlfUl
DC+oIOLs8T9Fk3U6UXGNig/m6ljCEQTL7UIT/ktNYuYodDThxW7XgQpWWjm8rRbd
9KqfiGN5k/DPgMbtVnas3pmO6gkOD9al9dMLDHIxHUkeaTA6Ee2Scq/BYCPuhYST
/DvwJzbkVGxqwjlpdI/YO0EWL+u1u9kSZmJDXSEezsVyp2q+hpjoDFRIXy7x3pYd
79U801KfR6laBk/+u4/+aCg/FPARegCaWc/yJ6NMIyoMFTST1X+Ex6HpN846WLT2
CdA7apTGiisYIjdamxJEhN9yXcU4Y+YrVbMrKnqI9gdpzWR6qZPNbWSIyldXJ4QS
4MfY2OrkTxuBuLC9DcIqrCHk7qaDypM70lGILgWx/MHUpK1izHM1PcLjeG9gU59Y
bjkFn20mjQCOEfUK4I/YTbzreAL7cliOA1TbIf5DiwTAEGE7uHAUunQ7AsvELvc4
4kCvaN3A7jUYsZQ5m6BTlKzz4oD0i62d0SO0aIkjYPKuFKS5FtzDmGfS9Sx9tlSo
hC2etGyScoBbs3auA4TvDwjM8kdh7mwi6dUFdL0PuWwQ9Z1MRuucT2NBCK2KFSmI
g3N1T3eA0RyssnQ8IrlU+ijk1I+3IzZFym7LL15Qc01rQHP9tDQhOoHpvw+JbX5/
MfGpqBt8Cd28NKTgaZvR98iLmaLC8ruItFReh5/q0VYLh5EmVP1uscOeyVp7aUUD
1pTLUxpu5WCxzTKixKFmYclKgEwXzsjbUqemNzTVOKwlctfzrhUTeS33RNsGxaCU
iz1D7/WYaoToi6aT/LCDJV+GHtln5LMuLncwM335mMvHo31npUtLW/G+k4hPTp1x
4qVFoF46ROw2+cvQa4xqK9oVk894KCiYTrP2+vKaaKrfGSffCAAZuzIX1qFV5Wfm
++sOenpdgURMgnqc2JJDaSZKEqPQDJpDYdlRyc1URluwSaJVFMogGkfLfHlJswmz
We/JZCyP10U/gDn81nOYFkB8xs+MlBBC7CN2uwOHtRvM3D7GiLRwflNxs1RWemn9
0hQDC1K24X2twj8KBz3wUSapIiMqvU/YFFlxZF6l1DWRPRWN4UtztDksvU01NqPr
f3LfpWb8acprKYLv4kF9kIWyB1fAr4Y7L5Lf7Fx722tTfcLtAuATvZQ9nmX33Jvi
V5qh+iwqcJRygKgbO741n0POQpatB8uDPipUHJIMYkOKHlW+5dkygvmjYqw6nWaj
2Tn1JUem727tjusu9lqULwB1rPIn+ZabYzsBjJNDXmHDYe4XTbE/ObltaUJCKSkF
GN6gTr3PuK97DrvGeyoMuUa5fYilgL3WpIlpKt98WZLGxPGuBvHpSI6pY7rur/4K
3TLD+AtcBT+rKhGSGx9yPeyHIgdg/vE4rLWRYRClhl/r+TgzWRw5gOr0jrgf4DVz
VngujSnYk1u72MBaforaKKMEjhhLYrNMpqWqfIjuOiy6Bcp4AixldoJYh2InwIbd
tLAG/7JQR70gt7040gk7R/XQWVGXrEk6sNA0I4c2P0aFGOrl2wFkqjUPMJ9M0ums
1G4qbnLuWvNIcdNKsx91EqW8iOvdEU5FIJCztqKrcV7mbVXej2rvH2c6+RU3xWqZ
riJwzqzgszRxeWMHF/7pG7uBRyybPYukZuWz9HbnOwrWbK4mZWmCRaCeP3rVC0wY
BegkOiV/C20/QJyen64AnE6oShPRtK+hu7gSS04LX0fLZbrU7aqBZH7bbQKfKf2Z
3VQJ4hDwLlaZ4o0vcYEPt+MsFhky+AZeBwGawfrRgyWfQtZvSaBO/mJMbV1X3GQV
MA0g5bdyTzhcmmovjBrU9xWabVC0Lyz4BzWAQNVpQZJe2PMg+frGqeUFqjStMjRW
DYEcbTwaLShk4ZeC0UBLxhzL5wYVQrLQvwpE84og8kmJzmjbTbSWgruJtmwkYLRj
hPttK2WOrgqgkpCzE+ROR8mzqlqVb0yGh2BJzBj2dh4x1R+TNREg4e9Kt/zcMbCV
Fj2sy9ZnMdPRJh/5zZVjK++ujDhmHpLd+jOT4tvsYj35PMlJ7eEKVo4Mp6evciTJ
KBPJLQs15bNh1xOA2LanE5poDQODUDRmj0+dXj1VbJ31WYh0Pkf+SDUfznpz19xg
BQeS+V7h8RKxTQAyGjdVVkgSGtV420FCcopCBFSN6BxX/PF27LyOrwFxqg7fcdCv
lzx6XYLaogqGRsHaJ/J9Eqt4OFJtH1M586yRjrG63BOQs0SdX6jyvnmh5S+tPECs
eKr2Qrr94eBXqGm8Uj1Lp146xbd7UQ9+7aP4TLYzIlTcfS+dpzYZDzrfuxS191+H
8RqpnelHs6LF/lKt0/E7LLsA3TqkY0KtD0pyBe38G3QU+iRtIYDhu87CjXIFN52X
Z2DR0R9Xyjx7JwJXHdmNaGuB/eHrM41ut8wAkXeE+fEvoyhYqvRvjQd8kOfzmP9M
5FOcml1EnSAQ8t8Vqm3ljbQBUg1Nz8YMMYZhQsv0PJ9uPxr3JZbNVK1wZ5k/X89w
NOkv5TzSKLcQRHEH4bb7jBUUB5Iv5ydbaJ+lO0w7SpSBgXo4cjztxe+i7ILRyhhB
g985A/k0Pun6S4KcXQr5Rr3ptfo1b/wa2wRkcICgbWYOpynGptgYn52lLOMRBelz
XUjz0XQTdwV6A9bKsvcaH1CXipsqRAu8tX06vkAu5MNO2od0Qj44AQJECsjzLUwx
hMAui0g1/G2ZPfIRVu/plukZuL9dYV212ZRSztfvd6cbDMAFVLKLa8+6GIjyYSBi
VUeMd8Nk9YEJTuArZGarBBL+FmsVgIK9hm+bnmpdtVri8LIphmCKjIy2i7uPAIsd
PrbkHkeNev5HpDZR9hJRHC80MvGgRWoWqhadeOKl3pyNOc9HU0SxTwGayjRCMkQB
Wy1QuVR5z335S0kQyNU/K1ghnxA7KpEbSQhJGfWOz1cs59a+gEygqECKzw1/GCJX
AghUO7bx2vi4uZe74JNEN1fJcyMgUM6+0FE5fqaw7a9LcRzdCn5Az7Z9MO5djJL2
4fzIu5frG2CIrTnTYR9qmxyS8x5hkOVN6hlB4dr/IwYkPQATdbaS6BoWa/FDIa24
8IRuySR/zs5k92+2Sp4l+wbdk+rU1BJ3nZ+2IvPJe9PnhXtA9wwgQvMCpaJ5U7qg
WsSCBigAp1j4PArpgafi9UyVXOa8ptcOynuIMorw4KFlfLKpo3AhxQCuU3rcDzor
hs+jgVKmIpi42TccPVV1xv3wjut8bmyj5y+zxutP82LxavufadfNTSkNw2ad21Iw
sGWpl+Hynh3XcrMyADD+ryWdaH6UdL8dKvrxXDTx6QYnjCb/PLCUe/KQXB7OuyTL
1EhWZzfhdoMcjfI4+crBnuVpVRkq6cMQuoU6gmhnpz4/k297Xm6mSyfBH8ROi2hT
32Cg7w9YYoVkK66cueK62gGKQ6W2w+/FLBZGU3gECCvNVN1wsJG9A3aDrP4TJuYx
bVk7gLLzhR3WjardxCd3/L4XFsqBw8yFNQUTKuYPK9DKWx4V1yI8SqNCusJspWae
HblMiTXJlUtpgnJ4KuZDw9A0H8DVW0TExFV+/iu8uWrChEnYFdCTJnEMPfBQdFlB
wv/r2wImC+bez5HfqUI4WeEbRAyWSPSM/RQ1Hh70q1mXEYb/kyZQGs+mDDUTNdcH
vVh9fZnubAtREGBBtGVRoxaK4yycOnNHNbx6+pwW3WOVVygyAdicKVWhsZa3OcMv
Z1/CVKCZ/ztuWOQ1kp5NVdiRuM8I0NO4NXzrnez+j0DHxwXF0d/EUVy528QqjA2Y
P5pgk9jNoHg1XkehbI+1eeW5tkBLEr2HiEn18WcKK4oLlsxJnRxtS3XciO4uMljn
5RVuRkvgPsRXteTSRFJc/FwZZyy7Lr48qMkK1vEzQnjiK3S1oD5Y1wvlr0zpaJ4g
Za4KwTo0AXRaoznqPnGLMtkON+iQZYtxR/ut6rIq87iBzEzxH3CjgpLwWKl4fk1b
qAHnZfK8GCyGNaeeU69ofsOr4vD+jqT7aQ5Acgbk8gLbVcTL3l+z/fTdncSTVSfQ
tlXUVd3vPEPD4siWV/kjHc942k3/hsD1UNJnmXH4x0gV4DLYEXtUAMcjcuWIWg7f
QQufcOgROdELQ19001pqML5y3NDJlpwBva51RjJo6DwMGTRmcLUvhXGtfhrasqKy
lDF4gZhQNlLaHVQuiXHVuE/bm/9HC9fB/z2FKit/w3CrhD9624jSac+dBv14uP31
IW//17bEE1mc+FK4T+VSnbP90QY239TM2llE9AZYPhKlaNr77bL83SB1x5Llk843
Gnks2H3x2zi8qG7b+Nv9qrOjyOBEWkhPbpC9BtxcTz7KTKQi9As8jMS1WB3M+TG+
pk01qLjWCF0ZWmiq9XbNKPfLBiUp0C/o472rtO1z2KVJ2s4bsIuCsBUT/fjmi8NV
nfQxC0s7cFHhyY2UWZRrBPBmNbKFj7IJbV4mB77rMGVF3TyPzLBUN79Yu0XB/A+n
Otsxu0OjBw/9kXyV+1eiVrABTj6BOqHC2CTLiG5X2Mz0+JquPvBTuyeh05rRI80e
q2SkZHH5WR4geA07PWCNrCuABA2SXlkKM1zrGmv55aKPb9ZsntkjJiVOe9apYvRQ
/Tq/60D2TmGXvtMsdnObgpVo+fZvB6hNab3J4tbf9TEMcpOAzwzg5Z0fB8myQy8j
9bAIBtakxQr2WTeqa1Bew6vhfNuGDAF58Bysj+2FxPtUaokNR/stYXdNxfMpnlsw
vdaWIwapMfxbZu9M+pl79r3tg6BdLm/T2wqK3uAUImfEQ2vlqjkd36g5tThRygT6
EGfPS6TR97I+fJsZJm5xaEnXy412BBg5dDy4FMJ6mDlNdwgRmfUfGmyVJ6XnCTdU
YI/7391N4WruPOaO7RSE6wy8kpi5tiCxxP21H9QW7M2uDlGzvhnitoTKMLZjHrSr
+ZjJtzUp9pzHaFaBwdLZr5wZiAvvvzQQvPW7pSGAUfdlo6FhJSl3vCCncyVoR0sA
i9GxYZ/OBCuZALsvnedRqn7ZHgmbAa2ae0JoBoa+g7To40uUw4gR+egr1PjrXCyt
V9dkcH+HXwJKWNMrTfOaMmU+7+X6QiMslbaww2Fw/5RL3OWMQm2lpYVo9+g7DvDB
dk7TGgz1cLyVaRc2bVgZhFvfhMECoqeNR5HxJC27vt24HW2ml2FTq3Mhv+x9B834
W+jSqTIa+zOU3dR1SHlPy7ee86FeP1WYecxwmodx6G4/FPMaFsUSgTnK8/FXEp6t
7nRrZa8DDEX8hP+pfG5YYjyHETtHdM1YXheBL5BdCWbhLjyOUsybRQQZmQ1K00a/
J3QfLYkSSqmt0xC94bAkwkdacQbBbBXbGxfpHIIV0yO5FXNIYfRzk6KfAnMJS7y7
ydQQ39IhOqYbTCZl0zIMuFt8xbSNIekBwEbX8iKivheVR8u2f8GgQPc04HuFcq35
35Out2MTTWtwLrYBA+U4XSI0lZRUl6KWzcUmv1YAgqp9iMHkQuCVd80Xqq6ZIFLS
//NcyLeYcsS0aJbIr8FkNVgAKROfM042dOSPbE9bLscU8Y64BfgqEVZldRR0v9ui
TVLeIwxuQ2C4PBTa/mZGhWOrMoH/ijD9NhNBzsGNnW7i4pRk86e4v7NDWRpNr9Gf
tEAAtI0TnGQuLsCiLyvzSEIRIH87fyLAL7T1u9hYXGZGIGKU7KujFhFWWn9AWNkX
1+TNYRs8Hi1aydHD4CS4V4sDQdhpSNwtbQl8FAtrbaFN79hIm85S2URBYLl7BWLW
O3oS5bfGH8iWw9V9VoY4y7r6lVIxVoGG2XwrKETH9UBVsWPOKkGUgsuR+oc3DAbu
E+bBY+sq97k4H74bA5ZnzKRpe+HNOkVQOXbP5cL0/43vntzKH1WXIuqY/+1QJ6Mm
KLBdkTvuYVszdn+lx+ECqp0g5z8xba7RmCFjojCZdS30Tu6Wfw74I0Lw1Ux1jCxE
5CJis4jyxK1doVAR0+4j0LaUbzPHhHKKTjKbwJjLPYgNgT7aJI48ZA98HrEgGYl7
Buosfsib26yWL0SpLskeuIECj3XIIHvXNKFyS7ig3xhZ+oBCaJGjxoCibyQ3y1U6
YKGzEDjykUO1KTZ0UOI8A3jziV4LNlwDKO53MgJfS2Q556nFsquAL0OCQCFNRZbw
n/9wlhUUCoRIJdJWm5tuN81VGfuROYlJE2/Dx+Wkj8FWaGe5+5wu1B3p+K7OQ335
8UOLq3VALPc3OeGAwXOeYw56x8y/ZA5fCSOUnkdkQVjAf0MGl7pyA2ZMoKM3ELaq
28Nk8GYOC+BBq8G8gF7Cxd6IGtMSJFxSYz0Z865GlPZFzVNY73+gaO7kxIDeztIr
6h1edSNhRN2jAOslCRp74upe1P8nX+dDweb/NEWV0QCkfGka6SGyvzv0piGW4Ogu
jrDU7qXY2YNPapz+EDhj9SzwFAZKO6tpjiSeRZjnWTCaNhXA8TcJxx8wMXwCupJP
vDfzZlYIb3VcWH1R4IYhAP3uHtLv0741bN2aeILY4uQ4figtd9Yx4+GqesJ2y/OK
qnOk9wjhXQPAD0F2b7Mc42vp5tIyZi6aBy/TOzRujDK82zsX00059Ix1e8waKc3V
7MsvHWTYBItYeniUsD6Cp4eXiRQIrKjnGxeqQlQvYO+kd12/V+HyHSAc7l1x1M33
lBBBMC2gBiYBhVJpYJ1z2i90ftVBGxbkllbmTy9gk7b6lXi1LbYLb9L8MQ7k5P/5
c5xQxZfOh70pE/TQDcMzIVhR45FvXdXYWJ+fbpLROCkmBViwv+5q3/05V/Kbw5VR
/YtWVfhOkpdcyqJqcLHG1NN+mo40Td62JVItGClke/l9NJe8oJoRgSGW/GYVnHeq
W/l55NZ/ok/SBJMoiIt/PTFxTjgouxM4fk+6M8OkgYaC2a0zRIoglXp7vt/UxWUu
VE80Xd2OcXwcBRWyi9kH/pA8npRXY6FQvY5UlG6eXmweYN3GTltKktYEBu27HyWB
0sypJLmmk+jK3rLbX3WC4eqfmt0LDDXYUE7G4+n/Vo4pna6BIqeKi07z1AP8Jeva
KEcK9v9qHgZ+W76CZcOdWdASvjWLh+wWtJe8r0D8ip/yM/c3JvlxvzQLXDvazhlk
7PArY/KqCcIUsM1i8oQkpMF+fimek8CjiNWF4hbbVypm3kkgyu3wrc5q5pMTMEtq
cpt/2O03LfofH7K/P1/EZTSGOC7aLolQ8v64pZRi36L/GfjGcQwey2RREJmC+7S0
O4sntMxOgQU1vgbQWWji6cIsREUSkwvxLul/5en13HSgeCQkhdXQBPaExeRGcZkx
nhEdog5/ucs9Vx1lg3VFBeCKq1v9GdV7vLQi+z/TCoqHN8/gw881vY3z8cy5l+rk
DQoziBJzFWBTGy6KMG0gMzBLCysNI7ygJXyI8rrh7y9R8suOx2rr7Op+Npi+9o9n
RvBOyX3UDBR28LSLgQLG65NtKe08Fa336xq/7FymZWpWEa3qeIgsuZdg++VU1mYY
0iM9ft8POr2OVgJ6ojxAHJRTXGn0IwijcqkUesPZyACrCYwcdtXRSFX3DjUpIT2X
DDM+SMiZSLC/+k6hl1Gs+yHrjrDzxAafYlBXkvkzubhGuyUGjjB9U4KM8A+0jTgO
Jx9iuC+YtaOXuWhzSb4iCojGwuYMKQy7F6b6dcdUBbg+ZRdK35FfEcFz/ajZ0zIs
J2YWGQG21Y4ErceyS6TxQPo/zXHLVRPeqwLd3lcBdKhSmx9/E/G+w7a9Vsz2tWa2
Ub6kVQwCvWkV9LzjH0PsKbeqo/m1k4dRk/QzYtewGg1NKaurTsTQS+0v3PNqGAQK
d0tisPz363YMzupBS9j7COQnwI+opCRDCCP8KjcReWV167jxCThe9jGYWKD3aW1H
6nDF3IqE8UJ/qcAr4Qj0dGkwnM5I9ht+aJumrWAJ7h2TLW3FQ9BLuDxMLtbUy8Jc
8f9U2oVGZkI5LBzE75zefLcNwzkCQciuZOArZSFTUQ//1K6Yu5wJIHNxi5kwEe0u
yLdAEpog+kpBcKYBvfjACtiswDk+6HTCvQU/h41bKJXSP69ogRAvP0Vh5scchGF3
AESlZw3ldFtA8AT2B4iPzUkQFVUQbv8HtoysD4CQPz3PlQIuLWBryfqzyaMR1S/8
t/biOWyzBNyIaVaPCcQzLacwQLhVEWW2ZSnCmGd2fdCLTyU0wDk2q3kpTJJPaJ9N
eWX+etGURQkVczzAExvsMPqyp1WxJ14Qy0MbMDNArTT2zCg4et2DB8+1ffYAAAxW
EkEaJjTlnTWfStjyNg3zLKtigPnBBIuJWg3f3OxYcQJJ/968ENdJJtRpeCYBx0kP
TySeYD+IZlst1+2hMvF8G7wIbBOE83skYUKuHsKT/ZTqCSuXyXx62BbkfRzbvAph
YDcaOM3N0lWZJ6IhNj7G/IzNWv0pT6VK9yQa4tR/+N/W7UpIcsMWoSd4kzjxKaM/
3HqBzC2Nn7BhtHLW8Iht7zgjiKC+pMRBlNZ5/k//eDWS2DFzLf3h4xfR7VXsefky
YzbqIYKr9PVCZ9tbDmgu31QIKu2QCRl9LG/RhvqYN231Dxmal5yP63ynrws0LA+H
XNPEcnDGJqC/vfrVTYC7AW838UFvPRrJmaTtUwg8l0L9YpTOtZGCEbv3+Gg4Ufhu
Ytr8Q++H/mRRa2F6ezWccRKV5PYc9AXeb+rc6PwDSsvGQ8a0+hlGqACROTzDThDQ
fHL2+bRnsoDKLeZI9zg/qch4bZWzFm/yQRAZZBZtpESA9VXNM4ohBc2Dyu2v6mtJ
PAFR9yxqiSFQjNH7xsF6cg7yg05E0M4z8geEDkwmQN9TBOpTjdviNSnek+V+AY1t
1isAFu+B/YjiF8ByjfxdWeBe3+GiC9mBOYY8MSGIMM8I5QxbijC3nDfpkVifSRoB
v1IhPjMlCJfcScyq4+mtmHqIskT9HauaWvZegMs8+86m1KCOELwq/PEB13ZLDzHd
kL+mi0u8kYtp1gCvMuF1qrJW9PgbSUa+5PRyYUI+87nUr0eu/Osb7bfhg/xB4YDb
jxyGsVIIeLpPhg1GUjm2C8WxezcTgCHwOT8W1eqd986ZUJwPPFtqzomPCWk+sIGC
YCZNbEeS6kFQeBDkrBAr44wB80N7JZVSyObrL7B99810xhoQkt1sSOUVyYEJWKju
gFknJhFwng1wfu/H2ElN5v5wO7g9vMsF1B8WAL/RxxwJ1wlYaaFqs7ieghvG2X+6
a3Af5u+pEaGAxmq09q7Tg5PGq07OG+cFcw+u7V96OVe66Hl5q230Dedrs/tdgSLw
7+a/FZYdcPbmDf+COyTLmo/kW/lZaz2iDPsQkSJb7OwXbmeccPHjSJn5ituloQJW
3PqzghJNOnveoBRtxC6N02txOoylXFOlamW2/ueywe174KA7MnWZusSS3GYco3mT
7t330gLYp/TQ7aq0eBqZAmQxw35Zz2qPnzck6gSEeTs397wySwZVihy61ooyLKWj
O82BzxbMEApV8oKqKNWWxR51TaHM32F9wpYus7OtmNk4Yju6B22YYLle4CiKlLdv
01A65ROMi5m7wHyZqqkvPRoNJHbLQ9c+MjxsoAae315jmIJNCFYeZNwPEt8kormF
F58SCx4OJFX7OO6UyWH+iir6nAirH0gEeJ8sFrhuMqlAoDV2jFaKiljwNdb3L6xX
WK/dbc3ZfDjAPrk5mvP26dc1ExcUXxHSvCvEfqYPvVfStpGOxMh0XNYveiULir9/
U9RY+kzcJAVbfe97k7uU4bOT24DT06g/pF80UiXddFrq2gNJr+rqFFsbDSx3vY7E
yfZNCVfKNWSQwdnPWFfDDhaE/M7YUUANkY4vHeSGAQedxzsIy3P8yX9U9NyVvRvz
ikNGguKUKZA6JXPpnCNN1zVS576+LSHH9W08CVlVpSCaKe3geF0ObRmiFFvMk5Hr
43zxwhYulmU5pT0e2Yf+gJvYpxyGEwkUBg+Ufu+++0DIsrTPw/B0bPVnSru9Nqqs
6qT6d7f9p0mstmgjv8Qe5QqvJm3Wfjd0gHwkclCDZo/Z7y2AnuOkt8Wlvuilly4J
bl9CKUkyYI/NdrlXPzgj6AMyygH8uXvn0xA4PPKl8Vx0xZ2wySDuktcLYJLh2p9Y
i5bW2WpJfsIP0noCJGNBwLacLervI9AZQAM17398K1HxGmTG8cIqXBMA9n7tidJ8
402mOc5x7luKfosC7xALaDOI179BwHPz+lHU4kJUTOkSF5+Hdvjh3SWTGN/pzdtK
flelpTXQGkj0570Y2Ef9YeoCcQuO6McuGm0ZcztgCHWMzzMCTCqobP4VRWR9zOpo
Fe6ghH/4R683cqno5ElGedNsDUWT+xu8rVAMLl6lArHXoL0WYsC4qALpy/LXncr3
2gUhKgTeLgC1nzYgvwY+qq+Md3fr8/YyBJ9vgqD9hKIuoMFkhwrfhNPssTd5g77S
ZfHKrhYEzWa17Y6rOjbG2hoGnyVtoNbuzOxEQzuK7SfgjtTvyto3eV+5tXyQ7UGu
p/ZfJpFpFgFx3vfrx1XX1Xa0I6BAbWs0pUiXawohOSW25G0SUJAy+UAdWlx5QI3W
70MMf3h71wOLVmkDCccOgabdhhCz1XnNtrJm3Y8jXUqgHOaYpuZPg6fUqkGGsdQD
IBH8osLNaxed2rB20jOR6BeJkeldmHuMU6BkU3hkyFP7Y3RogHDGvwa0HGivDA62
+hsd3tBjUvHimKokriVgvSlAtQi/oD4qUAv92xKPx0mC70Gjm838WPn8we11dMBx
5wW7QwO1YKfBdd/kmb0CM1KzsL+I+RhBL+fJNRHvldFY2wxjnac6KiTtiQFUJ8bD
1FQywK7/YVIr1A7KZ7n1Td7cMHjq0xe+R5cKxgTExW0gCl7sUCASVtlZeD/i0O6o
XCPK8K6oMKu/xeh0rKIgASx5DhXH74ElmTAW4h0kvvPbXQmFLoSz/eIDf+WGV1Gl
o8xMKKIXM2BWbH2GOeuf9EcxKpJJZ0Qm0VGiiBUJwoSK/9KUNUlpTb35InGjVuCR
61PnxE5ky7AuBMg6yHs4npeqqmXLFgZrhlOtm7Pd+oRnuqjfnAdzQ+R+3VUnctJE
HWKdlyteI2BrDMxxTWnPav8Z4amKkho81Mrt5ccjGmHy+7CeOoBS4wMvi5tmER2g
VpZ5+wFPassuwS7DojeeyMFy9viYTpPZhVrwXWFbC6Lp8Wi3YVgwUoPNV5Hxg9iG
HJceVX45jAVKzz4GNdVD4YIdE42KOHBtzo0Wk59v27Cs9TpMZhnHKdhuwQOuIh72
k5fnSBG3MubsbMI1gIm2hOkLnc+2dIOcLORSXzT1NwwlbNEaBsMcIRLQfl7uXCed
zQARDoj0qKDQx/MLthPIzsrj0SWP1ImjyD7WpiTWs+1uWbngMkNPbQjgjWHD3KVk
i5R6+f0ysRhS+AgQYl4sOpDegp1cNMdxhKPlDRxZvT9fB6bP83IlMlsrDn6i7qWS
/WCcDhge/LSiIhbb/XnWJtimWyzh6FDPERQksufXU3/Sa004g8MzykY/hjl0AMFL
UHqKSE/mw1l4JGEk9oG4Ue8IgOd9ugqwth6UFt4MZ82xPITUkfJsJ9eEj1u1DWjQ
nTVJwnoYSlBgdLlBu+YZ5R1VZGX5l60UNXGetUflLXldjob1ivUdKR0EU5CBk84c
URl6NFVGK4bcWgVj8109gdSDWgvOZpiLy1UQvYB0xtarrCD1UPwH50A7a5zTK0Jf
5PNxJm0LWY0w/Fc8+0OSqIA9YLqP4bTFJGSfOgoOXHvQ2YbIwptSjo42k/hUSvS9
AdETq90fc/Yy/RW18/ZloT8OiH9DdgM57UaMxrOK7zkPuhOsEmkzztmYHac0kc37
ipfGJBn/7+mJlzCMO7SlMVSSHD4hunoTz7V0kRyWt0KRGM/P0Bca/kemH9sV4d0K
4BHiq/M1HUfsasHU5amfF/8s2gaojRdTDBtsSwB28ZWdRAnYeM2ePBfOUxxheczw
ZuYGDFLIa8kSNNHH5pmA7qjKNSgJX1woe2u5VofWFuidmqpyRZZ83L1XNnrL7kJS
7OzC9jDHhtvpwOOkR3AMtMYu2nYL2hGUTzNO85iXr1oM7RPpOUxYQAVCtVrx2rql
dC/SbypbI3OZPfl2ZtMRG0EKMpB7J55d+w/siRIEWFvF+9sIsdUIPR1w5MmRKcAD
O5oO8oZxa8e0rmzxrnUTR5U+phS97n7c1Aez6ywHiT/yHGl7MCXtpf78Sh9iZqQ5
Q9RczpGz8MHRh4JgsgGtnGjPUt5/bBiQb8Pf9qiJvN8AZQybBlyTY6eKgzToAhHG
3RIk8YKjLuOF362O5Llytc5w83u+ZnKHKCJ/vnO0IzBSDZCzNtJ4OF6YWUOTurk1
+v8V5AJEqUgGWOA2zovgwMJkaUWq+kWLZsyOKOCszKeZDnlpib6MdzS7wyK/cqfG
COYy8j1/D3wuHXo6N1e+20WjXTWlQU5A8YsI4q/MsfjH47Re9oODqXCTnQUXYuB2
c3AoDBQR5j/xXA9MKztOCqWoXqtiqEZxvuo6n/nEEdiXhyJmIG5at6y3CxlwWkDh
9dzUxd5sTh8vvK69c/Ib6qIWapi3I+4bfFMmUakHP/pfHxKXyZO0EPsmiGb/oe/7
4ies2amg5pXJHUYvT+NmrRpqsqob8FL3ocZb5cwQDNdmMv0Xz2IZqU73r5l8UQlZ
5aXpnFyB8wqL0j0lxuGZmh+Fw0ttZ5HNMDS74XY5cmGVZa74a1LUFbEjBCvenJah
cHOJMRLrvddHMEtLR110x5iulHGLljh+AlAGQOJ6vpvZKArmOYhXdVH19DiyBF+1
0x1e3FzypgCbtA1SP0ShMkV7z+K5y3NgrMIHvY0S9v7mx9CuoBJrd4TUc7FYz6Lj
cHMqzrZO68+DoAblCYmXG5TzuQTgT/hTD7quVM2AiajoCcB8HxIeeubeM+yLXLVh
+SoB+3iiT4XMCTjRvfAfJ7kolFghzyP79/ztv7gSEezdCbPUFpYYVkcV2QyMdRXf
Rm0szFBCuElnx7Xqusi/9dOAnJwpIIAcTkOYSnbnOdqEEFttA5B9hct6uyz93z8e
6JCzP43jdnADJmJdX5eSqX+EmrvhxmqdKMGPW5vB0ER2MiBOELOowr0Cd6J0yJYk
hBHZCJk4fG96eN2EK2LtFZYN/FZjlNb0rqH679SG7coJ5SsqVBEK/COCHyDUCTIj
l2EdTcLNf4RqVTOTY65Amu2Hgcp18Q5odAopfMk7YDcreBM7JFrd37Btxpsr+YHe
NIAZ3sHRj9xjFIY0g70VS5B8PQovjtXuTjwh/xBTYrPle2rzyRft9w/7S9Vk/arz
4obWg9wzV0wh0Lt+YWC0ZZwD6JONFi2cdLqUPnGgcnxOjaHXYuzD+H5dlS80uank
Ld/KTJbBjxS4WkcmrNDqVr6pvV3M2rKCtwLGXWaoIaUtkUFgsyxYrxphl88YrbUK
frnXgmJMkaf36VTnsfLh6gO0/mTJVlt2M7DnaKVxbrgaNBx7R/MKGyzlfLbzTiCd
3kuYLUcZWeXOSpLQR2hT/9sHx66iqwZ7yg13NGGj4ji6pGpTaeo63YS5GC2YYbCt
Dtm+Ug295Sr4TtrXfEtICSUoO6hFfc5kz4riBTtm2Tbz7FF7urrxDLKQFYgoKOCw
QTMmxQWKAZRibJVPHksVHv4r6biWA6ULaY9x/uZnA3VEMPUAM4KSHqXKGAe1o1AI
V0CkDxeutYwXaQJjQaZWkeQoMPb2bSRT9Btmybb25S24ftr4XxaCxLRbVi6WiqDk
DHzpPDugcVT9i9L6hy5lUuO14ijcCdNji1kqaHdkoreeE24v6dfXXJxmjkChhiJg
PsyBOLsn0pz7GH0Y3LTJSuyeH/0XE3OyJuHKF5wkpu1JJiY6nfzz8vXRcSG3Y/Ej
q7ffhvxJqMmx+kKmny/o+SNVobk/J5vHSDkZIUrmZW2ip7uvqfuPFCrn4nTqb6nH
AKPVSIQAQSLtNU8H1qhVf6A+EzkqsEVu7AnNHtCsTbNvcuIfi0qIB3R6GwukMLOf
9AEBQIDcrYRb7BSmxWu5kCc3LLcu89rrBhoR1JUNlEfcwwivO4gIU/pvMKAmTTZl
DucJaXZd6/TvGmN4piFSaWBHvNCvuHqbO6JIsYhE06lOU7l159Ym2L60zfb8igz3
vKYNpY38Hv67KZpV2e/Q1YnzVcI02MihSH6yxb7E3ExT6NjhHLfbivtoBbcMtoiu
Pot/sYrp0nBUuVUR6MEjd+yJEMV3y/lvlEifh1CNAj2gP8duaSySMz3CXoc/zz42
hnAcochPT9TOwmabCPU62fIfKpYxAVOLcWjThhJ1fkhlEK6pJZMpPHBaU7B7ia0X
ipx/bthLPAsiWAzmUvZAE2AKbbaw0LxRcARSwYvlLumUeNlhcmSKPb+zLFnk5/ZW
MAMhqd8eOTuLockX/97z2WUyoULZ1hLrssvcfGFdX244T91qd/rzfTQoaxfhv8GY
lyGRYvBA6QxYJ/bAOPANDgSLVSYRqo6nYxWmG6e4eFDn6olY/OSGer8Imzk30/kx
ULWdMqkInF50tV0IqvtiqX8FE1V5QwbI9Br3/VOpjOCC1uFFCvq6TsxISgtuBmdq
mtcDxX+2uBTXulHBBWAVzRjekxIj2/fzZSXhjc4x6tKYDYBPKHSWB3g0Ecz3TqVl
sY2FXw5wnAuo+w+U4VVftKHVIjuTiiphbOlUHIHl1o24NRsrq0YnZkwAoDFkg9z6
6zqerO4qRlgwWz4xE/j7pw6jmzAk3HvF772xlKptDeuSUmpHygtpXGxWwgLglEBZ
JBnucs2a65/9KM/O3YEH8yA+TGQ1+f1+EaeMVxFhxwW67SDIF/o3IgjCC3pQF2K8
5u/6bWWLcfDC3b8ijZdUdHiA22El06qALAWlAPvUuiALcl1/kf2E43FSo6Yl8NTJ
PKzamRP463/mzJiB+aluFCyWDjAsCIYutTQOHLT5pQJ9qIT6a5V1jzqHSY/L0Q2/
cC6dZaWoj9pe6wMGg6E4ITZKmUQahIM0Pv/ABxeW57/ZQ6Z0LtJCweRBrkel90ve
Nr/EEktl6EAmjhOyp8tjb2LqxgJManxYukbkhUJJKIy670m5H/tDKATN74PgxIPa
0gO4zij+m3cHi80lv8u+OWd48Px2x9fKzsfi4XDcTAngFH0HtqvTi2yoWv/J/HrX
Hb7a7nDR2TwwpCYm7+nfxW3AUvwWCT3kQszV7rAg/wiPlY0dG93ZmzrQST5UMSLS
ccnmS3W0FB0PBDJhlaASwf9Nry5lRFQELL/GexolCogv4QWFMshbA/Vmw+g6gKEP
yZ4+wC5K6W8ukNJR9kkWpQpkXHN4xNGuLx3l/4kguJlX7d3UljNlPAc3AppKByuM
Og5q6vPGvcGvY+emlpL9QDAg5J+fTL8gLLyG9NmMLNT3rZF96rcvMbYH9FFkNMs/
5oNs78Iu8Jr6rTt2jx0o3XoShAEU3jhoJm1A6N7B7z3J1B8fsJBe/PnY6CvupEZV
l0U4fT53Ob2DmSryAojN63EMAEJphzXNfWGE9QKcAJ9hbCRnEAfj0VYMbBB4hkwb
qcIlWuEM0+kx7iU24y1zlVhGwLpiRXJN6HQGBko71KxvTkgLgKRpz9UWmff8MbgN
GWH6qmyrkXa87vryLuGpBNDFDFa8qaloTjwQIN7q5T0Zby8GrwnttkzKOftvgOfA
7a4Q95jzpxNHbeP9ik3300RSTPMwgWLSuRo3DChcXr332UFqy9dEct3r4CwQBR+X
4kYpH/faQgfU1NMTvWiAKnSHEO3mJ6UAsDI6yBMog75vo/5e1Y2TSHfdsCRgoTuS
tXsGnZ0GDxSOhrRqRV9O6tyjA/iOqF0Ye7KWmn/sWKi/tu1wUZ3M6Hy65s7A+7wo
oUasEV1SZi7o7jnFMv3OB5neujHsv1B8Huu8r0r3zlEna24UbrTxdCvfkon+oX0d
SRWh29+LvpxFxr1gNHiakL3TCqnm3k+WV9dWEvVRAf3AquaPFgrrNyRxdYgAoRrs
MfSD4++3MwS7hghAfUTa0pDLE4i49QQYe3S1t6+TT/26TdmT3NWGySAMXY6nuphV
gWMkeXzWM2cRs+1wVCG2P0HTxkQG72N/h7EkZd8YmWXMjtFn4a+fGyLcwdopXfWL
wLdIPEueCqtZPuDH2kjQRCO7/gKDCktutuk6ozmLOL2ZI3o88FuMmqaRyrTZJPBK
TTf9v713F4dUHfB8PYJEIGdhFy1fzNqTY+IljMxDHoQCgMuAn0WXqTe9ZR9kiIkT
nT+GczmKcxTrk3E9JwRdSn1gO8YnXWLPiUwVzlbv/kj91uod2oIREc3aBgAdQmfy
S6sp59Si6SwW8umxGFMUMJcNQwFeArng2kjfKJwa5SmJCQM7A6FpWSrz2aCtqn9c
Su9ItjNWiJsX92GkNeFa/gNORYnjcvadQ+iMHdydsT+rUoegA6MWyFs2WIXDnCEo
O1bpB1hSDo14Lj1bYkgCB9LZg3n3TJ8ohhlA2FR+pyg7v9HbjjjxH0bZFxH3tX0T
LVthyWdZNkz9KKo4Spf0pYLk7MKO2fciu3xC45m0ZFHid/20w2Ur1a/PVx2SNfAs
UuLMQINRK+8F7YPcV1rfYNQjR3qhN5WwS51PAmBhmlzgyF+x9ERGL3Mt9Yhodep8
udU75wx9NmhwLBeggsgzmDIXvrj5/FGyqlEwIVY3mt6OtjSwpl3c7ST22GXF5qYI
WcQRLWSMB+fB0zX0cPawtWzgXEpdq4lSCFb4dDnfJhB1IqRhV8/GkqOQ8b8ZtG5W
vlTAUDZh4GkhKH89+XbmZ6VoaqK3ydHiTJpuu8osvG7PRsp0vooFsdjaUTscYZF5
nXTChUQWL1FkZawczDCAhkrvJOsQpvbDuRPYINX/W8gpN6CjFO6h8Bko9fHAocGB
Wfgmg9s03V3jx9FGczYqQb+M0NlsK2LhbsDnW8oYILkM+alzSj9hix4/n2HflpG6
ILNV1pCvhmwiHItVgYaHGrYJ1XpDApzy42lr1+68Ceo5pEgKNdF5NJKo3NU+YPXD
qjPsy1BGTw2pUchXdSd+474Qbd7Q+u+La5NjHXK4DRXeN5KvVsVqL/9ZHMXHWF/b
vAXbnQlnlvfQ8ZnxU4bwUKX5R+qa2OdCdK1lf0muvwJ4rNBB0/G6hh6t6UEt5oWj
i7w7MZ9JXd44YOy6EOnkcrvVJBIx47e2cxbVeVHEjcUQ48eegGNY0Onl47XY5AlW
+RYT/g8KFFv4VhMCJhGED5UYKEVDx8k++Bjj27SR4ADKPyxQksTMpXOIJSzGDAwr
daEffCUJRC4cxPQ+j+wTVSyt3U97Xg9yUIoNQ4JiVPg7R9cfjei/Ry8jTxZaPqr/
7GMs/RKD6wHeqOg9gf8Yr3IicdL6Iy+YL41DwhRoeokNEUgGWkKZlso7Xz1BGKus
s4pcbkVpfjDCF3YqHN2iwsLrH49CJhV32XO4EmUNZWQq/SLg/AlMqfErXZ5HafX6
FQL71yyXffUCHyVn612VbQ9j0epUESvLfEe/CIRL/F+J5U5T8CqHY1Mj2GLu0wqi
0io02Kcsz0Rjq01QHys/38Nrk/XvZ8PEVhzUr7SYHEcUadXJkk3l7PHW+6OILaYq
tceL0FWe3vCnYGf7BdtdzrPpaA88mdGsu9cToup0+kdl/LW1pxWUsAoxWY/i06Yv
PwBvFsMh9/de3/6WtiMjN6fUgz/znBV/QOLvUic45a0TrIUU0EztL9cTMujgPtxn
IkVOcwbraDZ7gwuuYJYuVplxd+FLhdv9VsKaHeupGQEQEQBZv2JUWzwkwdcMND/S
zI0jaCpZ7LPVu4Df+Ww50p9r/khVvCyRtcnaGXlryERFMHSgenkNjC11Fd52MGYa
QWHRkEP+dAIIbVBm7Ic+mZykcjw/aQ8QGHt5DKvztSsXmMZ4MINh2FefAT0DivY8
+6XjZQmuqmKHa8U3zAswAsAe0fNKSMb0v9L4rIwqpcuRCvUBFali/PwOXCb+z4E9
yTnVZVtkYfQkg4NF0jnsM6psCV4r4g5pK5Kc8+HC4DiBmsrQUeCFQu5WoFBNktAk
mwYHkrtYMbQiyJ/uR/W4ynuuDKbHyU0ZIxWcOlWxr6kvszgnxiVhqVKx6SiAssnf
W1kH+PlmPDp/2Og/q85YrPufrC4375uA1LcI5UrYMNA4M1JyqSBcenn9JJOdZvtJ
X18x0MDlbQhc/Yj7CKAIM7YMw6Cg1Mg5hVMmra8907MKIMIYqMyml7GrN1Rd/4FV
E9tRx1JmETmGqM8iOhOdV7wwS6QgS1lGvv2At85bWASHdjsf+ymTXdYu1ebR6fNQ
EXMGsJ04ICVlgxasxrQKcLUWalgYEUz/x2Xm0Pc187onYsSSgrwE9TwX0ZRQrn4X
CxVc68Ja+T0rkhowW3vNkn2AonqpW3687G+jv7MlTQ/WWzIxFL9MopUpyud8tbMp
6WW1tVxQ9+K9yH4QhR/obC22g7/6lyv+FYczD0UgXQHzpdW0uLh+a8TZbRXxlHVi
AQ+s2gmUJUV5XYBOvjbJ/SqV6Q+D8vUcg41j9fSqG/a3ntAY7o7cTXSWlVe0BDtn
gcek431AvI13UsaBXSRt2yEWSLnQs7zQivRnkRwErUbGFgjZ/5rUomBzQixgy2Em
m5QbB4DUg4BYXGQs4r4eOroBo/5TGdUc5bVUXdzO2Lf/RFH2XqT4PtK3SkF4lbn1
mwXvM+sHtl3zSOqasgCrgtd3GkolS4Esd/zrP8qmCtG+Fn5hz3fpeNSfP/HsEeiR
c3rbvmuUjhdZ5CjsiwFn1bS2asexRYaxTBF+ZgDebuLjf41xIZ6hvQNKK+iJajH/
NWqbnHY1RbLUBJRO31nBjTLtHgPMOxk4wFFieX7opuZE2Bc7pPT8dS8HDJyc77iw
N4y+OajCj5pNUFhfr3u/dSVGWuvyF+IcHBrINHckzxKSzuKfFXPeX0WGtoSGhdu8
2mLxhAkUsT60moukoEMJCuFAYodwK4+TZw/Llz9muIlvZV37nRntt4KHd/XVkcI2
hq5JmhCGtmcg+e85f7iGBN+XAcnHQ2MZnAGXmFndHM1CVKw86vccbxaiqAviUN7T
IuddIOq6+rxR8xgWbfHWmM6G3byGZLW5c3fZdSH1d78ZIFHLij4OwuRuxN6abaZX
/14Gt0e+/+VJY8JZZBYIzzcmOIwxEBUWJf3MB+pfbuyR0vUzKux63QC5cwjnG3jr
alrGc+C5CX2t+PbbkI2U31A8SU3qVUH6/X7pjrvZuTwKcHQIape90GO3AXxQwgpe
RGQQ9+n+jfL2Vvyw48weCPqYEZY8P+PIS+SWWRD8jcDpgdrn9mhiCOEyEgM3anD0
oQVHEMMa8f6MELCXL3Z05YRT3UsB6Be0i57P7jYvc0RBZZFItrGk4GFXikyrPA1k
OsTxxXivG690EvE7PqejUJUncWK9GzFjN/ZU0U7UhcxNXDeClTjvWdfPGkq3NG+U
4vVyE/9jhH5/5zyMQxL4w7rKHkF+1YisUjcTnNlBRFu3sJSJS3kthdrSBMxzfwQ2
dJ2tGS/De05R3C973UX57XMIPzzwOpwUgEjuzZXdDEi57+eVNgZ8pdfOk49RhoOy
fiv5v6VSz6OBWHFXss23/7SVtIC9RVi1ruwWaLQeKsXbbbEql5a/4xNvrHzw2lck
6eq5rhIJ2L8L28W2CruDmzeaP7eZarZSNGZyKelTdg+8wL1jVEn3O8TF/oILCSLr
BMDtnM17dDDMBANj4MPCChc3whvWrCxkCc8G8QYvvDfS72S97aw8mIBA++RKg0xK
+2S7tmN8U9FN4Q5mlaOaoZG7MXNr4CYBRSGZj2DE5RdlLqM0gL3Ig22WXrsESjCs
e7NRMm8plWBK2XZ2EYiryKRf+GHPGphKNkQ7r926+mIOArtPCPNlLMMgjgJZvRGd
weY8q35oz4kJVEIw2EQlEetFIfy3n4m2pzOd1T1qDgau0VwnB3pue7yKngKDwpYx
n1dXAdlkRU1PBRhjz+AwoFJq6QQ7BbMLGzGIkGYrRWA0lEWFMFp3WfN6+McB+bE2
EkxgS40noR6burrkLmNEHCacC9kb/+FBQwrzQ0UP73G5A5O/f+o8rXlij690ptqx
WUeFFwG7IyZRUEw8mijH3CBrEBpqXBMLCvkWW+mXDorke9EWaaUABnP3YU8tUHr3
56k8ZxtTHETOnYTbvS2aDxm3MgTClVRpMmUniUaWechxQ8uAz7FTN7/WF1YxbjxS
MCelh8+w6NWGdE1Gno0RdWt1rASUH6P3CjYQKmbTd8yit1pi6vtuSPIUZPZ0mn8z
zz0bP5RQCg4dyu8A6J55Ynzh8hrx7JiJEtSkeqquOFA4naAPTcQV7FLYxCCkpxAc
Ycv6GoMn8GkNSjnmiHOl45ycJ/w5s4DgPd0yrh2HWXzAgCzDwvN/BJlF7rZkn2ny
O92kqOEIo+SqZfiQEKLcQpvb95FiPlDuOTbZ0oxgZ+vUhwHbcOD8JnDejYfzKSYd
kowtA0yPTeUkoip1cuJhQ3feHAbeRMsgKnSexczhbW57bLnX8bwQoKW1S1NAAHfs
1n8IGpdy7Z7ip0izUmv7+MFbNL/04N556+DFtftbdpMm7TPRnAuCxLqt44lUv0wg
1PElg2hmssRkTPbxwKUpKzmsZVlF8OmyzQBIZQwtRRt/BFO9AGV590tLeoJUlTPc
dICNH3vJy3wyFG2r71OoQ4oncbvft9FNd12GY+mki83Xos8nhlQzkj0lnNgioSIq
3+CQfFtyqu5eWK3wj26y97dNdhyekalEvZBJvZIdQj2Hkz49B4NEPlCYyYJZZKeP
4hpsfYi9dhVh6EqXvuUBv/ML64a4dQ1MJGOtiFESRg86lvDBzKaAq75Q6M0tublC
K8YNsqQ6yYA/hjLr+tYepEsq2V+WyaVfV6fK9x6fAaYEmmPqsfcgDRXx5g8zk4Ws
vQ4jZywFc+SpIeb4ZiGjqbsPsbM0y7Nm8I/EGlhPY07Sjho29iQMru1XMKe/FIjE
VYGRSibe4b3BI11tPObZgVcASW7MzVL0kRpEyOckSmCIUwS6jLD9DE+GHU+JIDKO
bdaDVVTs+yvtKYCAPXdWhGeaaxE94td18pYndyuD+EtVkgc+ECoWwEkQwoAGH/3t
bdFM05HjlMa8ZFbd07uWxi2hzvgYkJf91h160+MM7eK0IGiYwixyvEsdyi/RYsyp
798LTQmT4j3426Z3yJ5nqD6BcY+Z1ScmTecuM+pVVV1m3RAYbKJ9YtGsg46EIG+x
ygTdSmda5kS9zg1S+B8TldCT/IHzBx/nm1alrJNwImNZb29JwSUQbG2+ypulKhVr
OKpUIfoyPwq1xL8l/E0iszPRXoiCn4coC8G3+8315cME6fajUVt0olWryUXPpVgR
eiBq+buYdorywjuyybf1xPqTJlbYeMkB8BPCuy/foNd0kKEOL2aL63ICL0sKVoog
HSzkqIHcUTyFJpziy/8ooE3uWL5erYMdQ9jtBUZ0EsTgU02Y97lKMCdHX1FLyqfk
/o9FHr0GaXNR8ASFGuXqntXUUjG8tAV9d+lypHVww8SeKz2SflrCyYELw332dhSf
FcNdq0eLUUGyC9pOHPw0pafqsYPfxOhMPifcOAtjgQNTyFu1DIX1qaw20L+mZ7Tq
1ivmrOpA1fHFNRL3FlV9Rdonm5IwHHA5WOx/mZ8EhXAadc5HMVYuxPYduKb+Rgn1
IdCOK2ozFnK4/i9WVVxE5fJRmhrsNGn/fiDxZlTYsjpZl0KQMfdRJDOOX8LVYJl1
BJ05wM5RmYpNDTdiNWEqv5VwOgAi/VRPx/206jWtzuEeZTOmDb/TbR2PiOurFrbH
HhdmetQt9nok1g6q70iKq7CgivTKmVUvQbjsZOdVexuGkjA/Rh1c32tgh7JoTZW4
8RWV60y8Ti4lLR6u8z14lQ+uGPRlA8gu+DBgj+/1HHglRtXaLeG+xMOzHyAVTarA
Yz+dTsTZ63xLDxlokfx4/HYian5K1pzfBBhLme5ZpqCZsMaA3ysAbM/CWh7WkQI0
Fm8zFgN2hcsoSvMXpg+4AGOQMwYf1wUTIC9ZEcDulk7aFu+P85QN9fed+z4Ig1lT
HC+zNv+aYLW9QtaNWWVwEcEK78KlS/BBsOmxoIxDuBOi/ADVHV7jiYdEW7knu2m9
ZYbZeQCSeKrQYtd4JyKJ9sJ7U4CZP6txW26Mx3er+K43SOgj94NV8EIq586mKVGb
7oeq2h+r4TmFAEGszFPp51WxRcNkTK0zcgJJCzz34UlXRSYBnhg1IVDqJoPGfEQT
IurFp+57fyc89yIWs8iURkD54kp4fd9wkOmAWjLtQTtQjjTCdIq1je6o/FgKxt+A
h7Jc7NJjpDlwk7oFdXH6yUiK5u21CdoeaDbR1IRKbdAjyTH1ELixL/ksymHxjo9d
zc/Mgs+0Y6KOzZPmSfr0p8MXOVlyKSeby1oJ0QG95YZV/QqtZqyYjyR/JjzO5vRX
I/TfPNXlzvsTTW+Xi7mz8XT7c45aeHyLQPIB4236bu5XbUsiqmmtdBZu7X4BUY60
byPDvKJeurgd35RIWUujxdd6iJuCQZ+WIsuXicQPVQTR9YAJIWBOi9TooHPJxcd4
2RDa+vf7Boi65UdIqiFFas2J7gp3LakjHrCDA6a8DoJrhSPeapmZPM+B8NpCfq/w
iKFJX647lwN7x0h5zWi1u2TUBan0oKOAGUzSz3xQS41CAU5Ocdp2QaX8lWzrmsjM
Yv2iiVwVyQQeQfSk0mV7l4YX97+BLNJtgCDpFjZQQGAdWuiQwRRP4Y6sjolwmmyz
omHznqcYmCpnvWxL3o4O6ubHg1eA+VVBnZJgnnv/6csZ0Ik2dwvUgMGDfGXyOEm9
kIT5do5rmgtI3L3DNK0sipJgYgZyL8d/xGPPipzvRb8qh1sqhx6TsndhKmUyJjgn
305MMVaE8l4c2i5Oi2USr2FRWS7k2giM32KzSG471ZvGFKjE1X313/neScF8Echb
TRjbbIKQgPSaHlIxAeD/lZfmZq4d3b4mJJPwlK20RmBKkN5GM+LohgCZgP9/JOT6
t5jdaJNlW74+xs5M0kr89dlb6+LmPswnqDiD7kLFGc0iKfzwucMbQ3F5uBXL5TNB
8487BvvESfN5voxMA45VeAEtZsGNMRjY41wJM45K5u8iefWOtI+oghSyNIK0XwnJ
xRy4tj/F4gOsz3rcfaCdZ2HOKm3Y0gE9BbRAhWEQoXTdLUkDOhNZ6lmsmmZtxdzs
zKSjJFUandMpTnv32b9FV08xW0kT8Bf5cPmWfhRl//C4eKlv85bNDavTlEdJmUNs
BbB2I2Tw6ApnZV/wlakGM/Lgsm7AzbM/mBUbJxExz2LfhAd54YKYkagihGCfYNTi
v3LYCK3wu1hr4gtHlhVnAMT0VdUl208tMv0+G5/MrdBHF1LqtgcB/0WiwrQ8cyAo
Z+VdY6icZ4uA31ImZfdxdvochMQnZtO5HPlBDy3VfPngbnlOqG7eap6/O7cIJnIN
Au85NnXHbIsslIFfhttDSJ10UpX5LImoJu7EAByLF0fpBaSbfEZgONj9WqRC1d8f
m4UqTy0cGV9Jn2mo8UEW4Rev8NM3fEyDjatzhn5eWQpkojk9rVvudZkutSmQf3lf
a2LDtC9bm7qWhRXi05C0OWURNfouc6D5aPtE6TywpTcob3XBqy2halINN3zvsy5/
KzVOv2cYYaPIiedNR98u3HNeOaF18tbSy9FpJn5vBqCuftlfrPDc/vExM2YLEkAJ
5Ly6DSiiemRNrXu6NiN3qntm1O2i/KLQZgofK8+rrM3tcxCegP3xYnTuicOFjZpv
caKthG8/SF8piYmCS6MZSWp5VymJkV3zkuvh/iiDVv0fuAWEpLWQRmZ4tFgVSYeB
nmfTKNJwrDhzm7d7ovcVVVryhM28UksMrGWzej4Wv6qxENxmDnA0KC3aQ6TDweXy
m4keBmm6qBX9JQqXrjz42HA1kIpQt96F2mox3Qq+Pi0s6WnDj+C8VrpuicEBwzH2
8LFmC65aAlGPHC8x5pSmk/ZLMfwDoxstdJiENABm1U16Zid71FrYFdNlP3zpWA/g
YXKEY7XIZ3xI39Y1bbItpb0omUtND+TSibXrj+BJEokZEAXqh+KqbcgQ+qeDlFGa
MKLxAWo730gZqIqadVyjdYxy3k1u9+Z0ABVLG7H7EFNQWOJn8pKjRxyUS+N+oLLh
W4wXXirIiDfclaYADpsyCoO+DClDF+clIgUQLZY7d/B4NtQTn6Vdpqc+31e1jEwe
dUBJVjbPkqRnQ4qD/+EuDZBXghY13AZwHblLkeB28pWI5VVfN8zwM3v4dwBuiJsN
Ne945edwrxtbkw1Zf54WXON47MMBlwtFToXERTJgRgZ9tgMFejuGpcNcW3eplO50
iZ79PcmDUpM4Kz7BZAHNb2upxmeRcc/qPVZpP4G6sF+kpdZ088DDxuy76UouST9D
TtGPW/rnWpCxU3CiJLZPzShQs1HE1ig51K43V//sQC9Xs2Tf9HhVqZveBzrhEhlO
i76ruHtAK93si7WNqcSHfKkDV8L/yjURB5DIeY/G9gV2EovuIUb+dK6v3KQ9eJEn
kyHwA2uqt3KiN0zsqg+bWKhOpTy7FFHubjHxtWbQnND6WINL6Tk96pT3Yg8pYWGd
OCfFsu9HB4z/DMZWrNFsEhBB0t9C3nzL4wCv0AHwwmsHj1Epfp9u/AjXIudjfRUs
ikOPzO4Wh2e4Ip1Bmu7Y9azKVDW25A5gxWEhgh7LXZcJ0HNUJYhB4eMgQdOhKGtl
zNU27l5VFIzO2FWxWj4YSFZWAj+N6JCdBBkzjOVV8Ss+eeOWm6Fzvutfs/emD/79
YDM4Z3HXSzqgMluXKR2IIMu+P3aZkf/dF7W+/d+KxDGVCs94nvMHF+sO10o8dssd
l+Dl5thvhiCTHk7pOt8ZKsXORwyQs9NMY/0+XaFhkwpRGjkS5C3+0zJGf2a1Z5Oi
UOnGZ9E7UdPUzjLMGvRW27w5P56WyHuPwjLRwEj7yC2Zjy+b7PH5Re7TzFi/PFf0
Bv5R4eQw4N9fAyfYPeCe+4BT6k6ogpQ3KoYR4iM9Hg544cYPctXpEYOM9qQnr6Sw
uK+ca1wMeN3Kx4TSHDazAmx7f7oAVZlKEzgIc345vYHB8J/GGV3H9hh3iX+Opv9e
mlu2aNxaji7MaaU2aYzRwovWFtjSmGK8U5OnKxwHcn16vhcVH4ogY9Ns4fYy749d
EC+sW9Mgot0iAqzYFG1+E3cVxR1jfVsVn1+ggmYvHi2uX9RdoI5syV3JI497zPOo
gzn1RLAJfCRT9oQfd9Jz5bzv15d3bNumearslQ0adatnFuXMH19KXyc91qCcle/e
GbIYw1yPgIsh4A8OgfZsaC3Og9T73s7/8RsYHStyws3FMxQhukyURekTP5+9vvQO
HoL8s/2Hg4Mxe/XKPYgk9MufnMXL+8gPAm5GAhDdPeBMfL2e/lbgszKXNTh/N4hz
IXhMFmDNjuBm5EFrT22opUq+Dv2dvgiwMuC2x9KnFxpta5tPmFWLlpSQex3t0/TR
uKj/N5N98JhRlL1ZxSyG/mqhXJdUx0G9S58AVsZqLq5cpB2ctqKRB+uzKKcSTdBc
5wdeMVAGhQrUxqIJ6z16Dx0/buNMiDCL0yHKKTVTQEwiyrPSUb364BJFam3JhGxp
ZZGEEk6q1LwfegmbFtJwV/OGmvHoj6HXf0u2oyQBfSZZOsxYcdKMMU7l/nHQSM9B
dHhE71OrJsp8gn3mDCaB887/wUNdkXS42fyJ55e95Gbx0rZ6eBl85WoD9/kNk6KP
KoTCUOHo0+Mi/WDVH/8As3y7ensvr7WxmZSPKl07HKIESlPgQn6SwOxUFZAS7HhH
Bv/MmLierXJI96w+e/nbYU1FbB/oTd9eqJVtdTByv2F/BlbbRRxViNJqOnhHwwZM
Ofa8LXNxISj658WLNEM5RrS64HP1ZEygINjvizcMvRBIXwzXZG0kz49VO1rnynJb
I6tM1UzzXsCv6AeS9KC/t63LNLi1qkxD5+RlxlUFj+GgQ8iq7/ttaqtVrG28hDyq
AASdxOJAsK3lI04oKJ9GZ8sWsLUR2IPiwfyjuX9Ik3pK94t+xWx8AYDTYQ6cxUrv
a50CPeIXLinOFmw7fepCTfy7HooADq8U2DMpHaDtrqxpeOr5nkms7AgG6o3uoG+K
MDafGMhUASLvPUw6moI+Epx/vRQNDz/lO62wWsgWD5T0KLekV3Tz3+RC+f0XIgGP
dTNmmyKtStoFo+s5vXymgXBZBW1NAE4G+Zjw2nBUngm92h/Y7gzy/RlIghrqapBG
tXX5Cjb0T7+wWUJKw6Iep1DeNYV/XHeiUAzk7f2/VLuX/lRV/jTlzdbhSJL15BNE
fWlMgzKCGaS95ZccwU4+EHSR9lNtRU7tXAzsi59WpV8lEjBkMgaHJglE+3tsvjdZ
f8nyPymcfRRkqDgp3OunaXhc4FcK7Eu05z5W5qZMPRxkNprU1vLE+mrLi9/hIGSQ
gHzXy2eSEsGp2e2/ok9ZeRvGOux4NkOOnRVWYBZnREe/LJ1iXuPcINBp6v63mlA7
Zj6rvAjWPiskDy/qk7HorK0xu9GkYwy3xsMlPTY77Yx9wS7qKmHCuKNoujIYS/35
oyU+IuunlohUIBN6Sj7qbRHWXCwdPSlDJL8xTZNnT3OHJIvvXzgFMWHgJJ8rmQrV
KA43vEt1aorLbc1+fW45r/UbcobaKYBK0Sv1a3lF8Z01JYBwEeLM6b6K83Redg6G
dXvVfLxwbJWQCk2uT2H1I0hbnWkDRY/GLnmEQKcBSY3j8mvRV+wuvUnqPCSfSitB
958zBTjKg1zA8QUIo3FYcqxyvwnc+mQv9HIlx9x3PXTGRode1jwSjHhsr1fl4h/x
fvmnBG6QlH81WZS/9P254X7Z7fEAl8ZI1Po33gj2dR7HdW3f+8sxSNcUW3tIQpHH
J/aOLIBd2QvcCubV+Py5URhT05W3m1GPtUfjPAoDjt7cyZPuYYPHxHxC2UZTy3xl
julrvSxWBwSh0E/U+u24zuBL7UbhzY+Yt1mQq+X847GyuvGVfZV06oHPMkZADtHk
WkVHptnejH67C2ATYuHh0aC0lxe+um/WUq5DlPzZihHLiaMWrEPhHcwYPc6tiE8X
7PJkvnsUj+3o3n2UM3GT0lSeEZ1QQjSCmlyy3Hpzn0grpVuDLkygeU7ZpoVigPgd
qsj63fR1Enj0geBYd69tUfWh38xnj7unKhPVLknWvp9o0gPKprtbVbt8vDUP0wfQ
xBr2n0tgla4gF7wao5MvXBYC34GjMA0X+B9qzU9R1zdpNesX7cytDSP5dj3TAViv
BBOfiiqzl4+ziuVnTpQIeaJbSA8QiZzrLkUMk2a2M8U7yFNBxBoB2CIRd09EAIwU
oidaPSS0eUHyby/xXHmlNtEDxlvDsGXeRIhiIHU1yaG9xbEs2t4m3sM7hHAGYYia
gZp0XI+KuL+AELYwsfLRJTP9TDqHA6jli7VwGzsVIsFids3yxgH/zFuXuBk22Z/X
1TA5+yYv8uhZhsVHW4RWZxGuhi/xuI7ykynuqGbqkcexCzlE73T+DI+IWnmCXq9S
LsmrBy7PYEz1uPqTL8C5sA9JRVemBnWNAQapFcOsFQt5SwPE/OfZQMjpvA3lR/mX
BblzoReNdX9amb8gLYRoLADUQD3iC6KIbwqdGbrYWiXcX7QEYqUD0T+Ac48plEsw
oko6au5Lp9cB0WKjoFxq8EW2hVXyager2c2TH990TcqI83maoBlTQ788C+jAObGk
IEcnYhVj0sSUhAFo3OGIYjlu6v0h2jLenz5C+QLIobuKQkEh6/d6gXRz2r1sejHM
XGlkYYXEFCmPI+C8WTSvXgCoUi7Pr0REQMeTNW73PLnEZNRKjj/MirIuZsrLhlfV
BeqlZzP1wsswJyhvzHLGQcpDT0m9WwUtLZVI/25czktZkhVkJyugOY63AaOlnARH
JeKwTVWNvWaA1dSdZjHe45pUluDL664Dm9Z2xosPmu2KAvG9MO4dDHOkU8l7Oyn8
6GPXbgrqgfq4IBFjcG7XQUdpc1dGOxptVddDGWnSDHad7IhKHl23OqU2FxOG7wXe
QW5O1QW8J3PQwHmCo7rLVIQax91tyApdLW0tPK0Q1izVTGNmgl50t4iUDUXURxyS
v+tfyHUdAiK7rtb/uis+xm2nSqSdpYoniEk2mD6MctwUuQHVZgaIvI6x6zS9VPmS
w3+wE8Cq7IRimmWkx/1x25mN8tfinz+n4yxTxvc1W0K8dDTHEmiqXv1XJBWhV6sY
kIvK+5wTiaLMo2WYtl4LMVn3IMjaqfmDk35Gxah/QppxY/fsXZlbhepmeMZNLqA2
g8J+hdOkBOc0qW0Z8TL4DB84W2jYz+n986eb4pPtGOPbvlMoTUxdCmIoAQhJUerP
wHMU8tg3P/VL+63vbAKyaA1s9tdSWEpiX/hD2IxlBBT0q7viGGKiWnB/v7p1Ydnl
1OJCvcIuWOc0ZThQUOxNuMMwwkupHm4YLuJYHMeLAomGfRR8SQs2T22nXtEMRYkZ
n+J9Qio4cXUiKTgU4xT6CI8AoIg4eKA3fKYPfXolnOuUZ9V7+I6QUUeAShzq4FLZ
a0i4Ock/jug+FvmOPPjw3F7zxRbLtuRyp4q+jkC4LOQdIxEWc7nP+N3luNfC6ECP
PvMXOfn/AvwQKERoJUg3LMSgFhnPvF+bcO0EUG8Aa4ts/RlFLxBnZ5YiTnY718Pr
Mrm6hSdAnGKURh0RXDAmlFz0HyDvrdkywL0Er/j6avLQrkBV4Q9oqvONM9ahgdQr
JlFs2pQ5/IpJjDY8OpBXcL4cxgoZgsYK7pmgc9M8PV7AeJ2pvmWoqF6i4jZuKqaL
VYl834Y6T8K8au4kgGNN93dciOh85LYexr3E4YRkpAufbx5XyXIm08NWMfXR+Baf
/dxrFm1ullHtbSJVm32BF/ky7RaMNzO4XImrsVygYLfsPdt61RzOh4kr/fqw9wkK
wWHZwwHKPSA4C0JKTV+av4KYb7zeRbs6vFu/lkZgX2bSCpvzvtulY8t9xRPyCRU6
ERFuJp+gjBWqKN3Qb3hkSOiniDeChGypI2g6wjHezUGq/0sX5FaLCOu+WXhQZB+Y
MuqBS1FDmyDE1vygriYwRUcV9gPGvN/JdfRv0g0A9WXkiJNaig4TmFkxEaBu+yQj
XQphoen9QES93/HNvlfu4VE0KCNjqx4h36H9vguJ3/ZJzq4lUTYpmPuML8wIgYo7
pnWdy3yaAU/zffaVMrSqrvZ9F44YID/nlNPbbbYA7O6pv3rUZr06jDPaC6RyF+B7
XkPbt0exdzeMs8k9u0U+bgUD8z/SDGrz3kguuF3Z898pF2vA7A+HhSWAEqvTcKgJ
IMnzH0HTjhY0OVjbXVuJuZHtkmmX2UpVlglr6uJNdfh1hFFJHysOQZ0ofFNsRr0J
cOKD24xrmDUgxYooQiRRQROSVo8F9I7SQzvVMPEvNQP0mTJ95fpj+Na9K8ko4CgG
hFAvCSGL3cT895dGN0Q+3bIMDMlFcK7X9ZIAf6H4NiVrg8pOxnil4uTga5qi0m75
MflZ2AQ44/jk6lmHppNgVcXRgNcTOgQ492qFEV4rFbidL3+q2jcG27B9l1yEIKce
SOakUMYzYCMKjfYON+j8TXz+WbY63fa/6ez8oe5McIekFx9XWJNlpyGbbFeBMXUv
Bc1j+8ctD70Y8ahyTWpA2EJJcuZu2486XExCKbUf9HZjShKFcHyDb/TOjYoBjAif
rbTC0xxxB2xLx2iyKlmt+3OiQz8fYl4AfsToS2U4SLALC1S7NihhjZSuySCRHgs3
JCwN5HKuxTORR6sIkHy8O3uGXl2eDjA9hqYntrCwfn2U91W6pDCfZri5rbhFwoVh
VCecNRKXEnwwatO/maVb025uVHphPt9g5WSXwC+ysmvJWOISzbmkf2xzqKnLgpxP
Ab1eQC/Io3sEQkuzPvvoK94oY/jiOKy4EUgbbw6bab8nadYoEqcown9Y8gDaj3xN
3Gzn7b43x3XheMhGhnAEz7zsi4AzGj0J4ngyAoPwVqQBRbnXH66sUIICagVrFTs1
1M45+BrXzYbJ1Z4tpszn/9zkL1cdgj9sD4fQuQcoTy+2LQt2Zdmqj3YwilXZdlOc
Wu6vDXYdU6QiK+rHQEx5AGk7KCpCZl6c8tfRVrXW2rYRnvKjeQdthRo1k0emRuBe
VomQRVirWDIdwNI/dD8vLiDwPWAsAHRWEduvHWmcwTeF6aOme4B8llag8aSHTwX/
XmR9Q1oVCOtYKO6XsDQYw6K+J3BvZl3FitA3kq1G/L/EvzivELv7s/FjWPwIY2ry
Ir2A4lsuhXMREljfSI7t8zuKUhpik55KXT6LKVj+Mw7/B+pSSqISvufx3Vjf0ga1
Jd807NBWbxgvv8i5YCXpeNRJ6qpBvXipqAW6mtA7432H7B6CaMyU7VlxccYSMnfx
X41J91N9wJpPqBg6mMjq1ePPHjKgr3KaBvwC9T9TaQbAiTIhXO2E6toQ9AI5nezP
n3KoPQkEocxN/gOkbrNcZTnkKdzSpTQZjtYc99sFf43LE7TbqsGImeeG1c+Tc5FT
52yDXsJWS6wWo1vnL4rR1RGUx4rBPHBwlCwUZfDAJ0mcjkNqqacru6GE7LxI0ZUW
TWJhGhsesihxSYrLMCjme1TlufdiHWABsd4/4Gxo0HDLw4S6amoNkiYf8GLEB66O
okFcacBe7STYhPYBPbI3Rabr/pfuEmZ0Jhp2W4V1Afyp2XuIb3HAlA8lRpT5jo8c
dWUSVypY+v1qhiTYc3N9ce6D6uOwMYQDt0ZYxy4GG5KKSQguYa+fcreKSthTsqRQ
lWHK+BilD4pCo/wtg7TC7OgxIw73Z7+SN0+NRETQ4CL5J0P3fKTBSn7ei6d4D6iz
UJAqh6HnJmCv3JsalACKY/aujDfTNn3pyFtSl9H95e/XK8PHZTPb/YvZKUx7H5vl
U7kSihaGJUQxNMZHm1dsNKDygFY9ZRVGzzhltDsbq5Z/tmlqQQwVmHhbeIIsSSL+
Rhtet0axC/m1pFZiOi5pfjecC9lNfTaLQGruT4bFQJbLnk6Tsn9qmzQRo/Lpbn6I
HpkCG+SDYxI6GGafkrollvXrIQEGUY2M2N/uc15NaQYtg9t8ws2VSZ9ELcTpxFEg
DikOgTybftXOthpcJvVsjJkH0Or/k7JjRrOegdFiLqo5CP3xE0jJBjiioM6hPrIC
stAzo+Z7rNhsZYm09erJ+paqgYwH/T8Fkh2wHERFsHlG3IbGxCdUmA/jCnWgnNuy
vPceZfu2x4iweNfBzrDBD6qX/KQH2SCxMwEQDeWQaoXkgq0NGd/ZR4R9wZjx3W7s
CmOKmOT7e6b/hPil15+DpzK5s9W/UMslA5+NILgTIH+N4IrawLsaN208eKGzVLA2
QN3OG3UIKTQ9tNnj4yOBmZ852xzOJ52Sohe5C2fUzsizxyQOvE+Q8zwuqjXMQv9g
r8i2zSQKpfW90cL/CCj3RvX/pi0CI80TZJ1iclgZuTA9IfMOntI06U0m3h++NBLd
1mr8LN/bo+LFevFCecrJQimnGhzBFfO6UpLO1yfJuNRvrSXZmD7RfGL/fgRXWg+s
LC24ipv+5ts7RwYrU6xFICNKuo/3P7pIory+gJO0RydFvwbWK6UWJJJQCHnB0hoT
4Hhrq3J7uITwqYj4+ybbrXoD2g3peSjuTgx+jFU0mP7nFuovWa/m5T8TXJF8Hig2
6P2rTpiWQu9ZShKSbKhzY7cHvRKsQAAjsHNWRObgbjTKi+tcs/PAjGWWayJnS7zn
VqysuLXpOWWINOWLquD23R6a/x7Skil96wEGdRyl7JOfVEeHdZ8ucBCgKzDvzHxN
6M33lSKGI1yfXlpIAygFAOrOL2+gzNmpbeS3BQfjGFWFHu/lahC98+/kR1N4qvU8
Q1k20WmzxbgknPWMYUJCa9dGYbnkIeEtX2p5VD8+VwgAWIbVC3Ho0MyCVK+gExIr
m/L0HOWDL8n+LWrRqYrkyCf4+s6bBvmRT08iTxWMyHWr0IWsrZVF6x4/x/Kt5YiY
nM/Utwd3GtBNHK+VUO3PEbfd2vfQS29CnsiQvM/6LyGN2HKDngdVhtvzoT7xplI5
HbSs1dJKgQLOukB3szNolTg9hqYDueZI6VtWDv0TrKW5TAql7DJlKH/tgNN7BGJc
lCJe2NrPEyFzli6UdMES6OXpJsTAlJ4r+ne6b0OtVLe33nAz6IhSpDnSJyS+Xqqa
rjNg61nsiVqzN4Ezd4wwF485hAW0Rm2mkSwjC6RMoyCeEZgpbn/g0YIK98g3gU5O
vMoCvoshnP/b7BlhyHCaACrUeOGKGHgYYNpnXGO5Z06q08SJj+0HMZ7BwzEUnEIN
xd0ARbUDXO4gIFUfMjm/7gwsxwfmhZa0TzhHgGRNwRxFtyS00b9D+ji8YmAMsRXf
SsNNNXXc3YCj3UUMHRcyVXR4/rPqWPKZMz5cE9fCQVpT37mL3rnzETWJ9uUXW+jw
HvC2Ret4nXyYH+3e+g2Xn8Nb/xLOmVSp3zkuRFqoev9Xs8WOYOgInb1GtiTOJVmx
U12tcDIHr+VJFHhlIuuA5I/Pufovj3Mx+NAwYoCVQpWoNpyfGAornPZDX6uaFNJ/
cvb5LCbEMTOhzR+yaSTaczumKs+75896rF0um+9oKk3gQteICBWmb0N/Cl3IBecH
xDDuxHt3AJnO83Rjmmec843s/ZcVz44rOyC9JRQjHuSMunrHt9r7KTpERzMHE4YY
ZFSVoR61xJBTiXSMnsgDgxcmqHPfZCUA2sWgOEXXieQh4vi8nZFYvj+FF78/NxsW
cCapiPTJjMn+ZnoebRh6gnoNppAk3bj0GaKo43P/bT/RITYMDSUoeRHYobfwODEj
WcKl20FzSdu40x4aUZbkYMmw//jzxXwAE22FghqGhcU7RLYZKTl9xnjCVTV5ZRvu
XRrGHgmjjOQNjMHSnJIXPPj159YelxfmgeFAhYYiHicF2INiKYzZ1/fBqxZ2hWgn
+sGCta/UuhrOemox9bolSxOPKPwfCT/qLLw+8XlkIodkx77yzIRm+So9Epxk6vGB
Ox3JKNoUaYMHtI1Dh46OlI2zLL3xhkuO8BQWhcoCZT6TtyhG7GHBoSHu3DcoRdMA
lbdl2lLPkXTtI7jROht7L6V2TtaYdZnc7MWxu9g8qFvrbTj8DEgXCM9zIL56BRqu
fr9o2n6dGBbOJJxSXlAhe9hq5fIRGHoahNlRsx6igHpiofZ/m9JpBRBbtf8Aed/D
SMHSRtmPp8GQgD3CraAe8SOwkHMKfpxTywqb7QaeE0DDOfT2jkc5tx43HIz703K1
sm+tEp8fydXxlIcKaUKzh9+RjEWvlSv54fIIHCe85PWp05V72EJMksnhF9UGHPRq
Z216YjI/B4dwHWNIuNKtqXKlS6ieqiT1tl07Md1oNX62RZg+QhFIeUGYpotEbfyx
fYK9XoWmbHxsfottByPFzjMFqR/cqtSaynk3BU0U4PGFzk2faUhAmjDJeEmXesCD
kKbFjMh/5ItfVT4Fu1NLsgzjixV2FQMoKO7pQzKfV7Vppbz1gKPiYD7fE6jYkYba
XcdRDWzJJdPvzwdxVT18bubYLct6WL3Sju+HLkpivJNvWeX3l2DyrFhZMouTFHRQ
Ka0g3xrFsMVWB+dBKwp/MFTNL5xP37oar/nPDYqP0X5upsT16JDxweP0pN2o3d7i
aTZLUgBtyafMsaRRRmyDa1l3O2ryZjOOV5UHKONqdH4vBNwTFPs+tg8Yg6dtMnkT
i31OQyrb2hHb0BzTh1/lVvNznfMMG/Tb31rYnd8rW+2difbfTAkVXhQ2cQzk9LS0
TE5Y+r1b99K9jFTd9gbivOKWMROIJpbUNfC/1Vb1XTl2d+NIsLEV0m9J59+LJ7sU
8+J3gCcyxvcWRCDTDMOaT8tOLVn99mRD4TdobfX0yREo7SBxGnFdhb7s2sPTCFgy
7dTZgbhHjZ9/Rk2cBYvHK2GKBnn2zhflheYyu2qJjuoFyCjIoSYPK0aGEDxHcB2s
2r8vBTHaKr6Y/VNv34Q+am1EC0OiocXmIz6Lnggu+9Npane8irUxp4eyTlmpSau5
NtU0pjn+IQhgSxWllXk8Emrfi+YPuKS0p4c0G/D/RXP1iyjS/wcbP08ig85pkIOU
9UPhyJU8iWcR1OaEwmVtQAag4ekron5FwOTuSCL79LMF/Wb8236CWaldrGkX5WQV
73uL41tz2nZcbwTLhdnjInSZZ9tRNWJW7B4CDE03/5lmKgsFhti5xtW9pXHa10IG
xIWDqrzaq6mLeP0QGDodsJZaJcXDh4xzH4x3kLa3khp90v0DHxoIVuyiyWCXzivh
IsPjzASLb/Gf3GeYiEu9V6yGp0D5spezyqr5VwvnDFKW9G8+41psY6Kvj7y7BNMO
uul9PDaEgqUARb+7UAACbhdoH7VqwiwYx+l2aM2+MLfuOdG7u19CffLzLuXeQ7Ea
ZtSjIAkbL+1+yQAipVgGftDSfg/+qbXenaIqbxGf6UHYon/9uid+4+OtrB6Lk+/9
6J4+AZqnye+i6i00JL1tJh76BS/8mfLuoDFPMFRZ/1Cxb8nFICNf34wtxj9a/FKK
14C+zO2+qwGaEgN195qxk2BHhEEmdeIvjEgjytedSIag/eEBtTDy0DyQ02TrNASa
tq/erP/N0vZdYp1gvN+61dvZiXnYhI2qXcyryhJ8xGw6BfF8tJ0TjGwwOi5Xs9lg
HZiS5Y7WvWGdCb7mAJ8Z8Dvz3Kkw4N8DrmGUQQTNNqS3vbkbO41AKY0fi/kK1EUp
Z/tDlFhFZJOjfPDJg8ptoAIqltaGauMRp8txKCJR+quSRji7C9Z6qDYhXvqslTQU
Aw+vKmPYXyDo/NKw8bYrzC2dwZt2Z4RoNoZARafy58hrBRa4RkDFYLdtH8crOoyd
saEXdJuyeEq7MLP4gEPNcMwo5Nomz6muIq7QexqpuvhMy3MW639elCrD0FFmJ64b
HtA8GrDfEQTdruHwzFJbkTKVYtNlRPp5MAN29gFWQwsHHwlzRTIBYEoaHtBgwCQQ
bt9Ha2rxY2gK9zviD9tg9iTKbS0k+x0SQvCsKre0v6X3g0RC+VfCoJoZF9g4tKqd
MGKZI1FCP255vPQZJaTQLWXfjgAnS/TFO35/5OWNZRKIk+oTXQLv9ik44ZZztgfs
QyfPUp/bsLbVAT6k4QCKE4UvWFEh0gQOn0iTgyegto1xK2w9OWItrH+IGK2uf+Oz
EkiM4q2FuqlFMfHwv91nO+bEf79kPhiO63JYPioNYPy+UkWYPQgnINx+l5KcUOtU
5pGtuq84w+NUS4BekmJMcH2RYs+kctEfmBnIwhh4gAiqc57pU5dpv3TgB9Hx6SPb
Giw7VZLhqpaUoitxKBsreh8Ne/YkAt1NSjphAY74V2RTZ2C6s8Ie3oDlT3YRdIzU
4W2stVRnSWzMtF5SeOwdNn1jIWHTdtwbT3LQcPnbtrgrv99VwjbEbwek7Rs9kq16
vQEwv08io5QQK2oLMfhdCRROlxTviz5zrTEPAWh3PcTVH9YCtlmvC11WfEU5Xfoz
PoMwRRofS8Sm8/a6f6hdqZw3wWJBcxeWRNdUJjbZOgClcFCdrtiRztJc40JpDyDs
/a3P/E0LzsU89U47lriHozgpHKsGAh9GAAokfouEEm2lLNCbD0K9Eh/+TqFen48P
7pyRX6DPM4NGlQn6A8h06ud2hIA4RjUtE7M/GO9onssOrWU2eKUuz2GeYQxUewNZ
jf7QW5OvSLJ/kMOrWF+2CH/qOOFsH35ILSoeIV+OvKGcTBCD7CqpP+Ug+xbkDwlz
imqxXLK7Q8xhsh2YbV8REbnXdAGlkUeOsyL0oyr8cZsw8a8KXhvmLsiQYrLZ8Vwm
3VwMKElkXTUQBW74/xBNtqIPDdRuCTCYAHHYHyWLRyYb/mSnhhk+cJvpgjGDkLZC
Eq8PMdi+gilcPK+i/9K7xY30Oo6gRk43mNFMZpAyuvV03OgaRp1xXfCcUok6Tp8e
qB9BBuJgTZg9HYJMlbYwH9WBb2vSDzD99wxBQejuur1Pk3ymGsDwvXMUhgC5RWQZ
SMwQIJyKileTXx1EsVu1We1YvjBv0PkRogIaLLyfXDVB6fAeWtKKiWf5no9qItMZ
wudTGiZMMFwNxPVYbo35t3on5C//UMZsJnz2035NKsQAFf1e2H7IGklamf/Bl0jO
y88xlocFmiPUhkdWkuRZaMxLHSockUc3tAL036lv08gVerkhQwM0lbyd4TfZHTUG
JU0Vf442QEU6b7rroN7KAe9aKV69HC2tIaat9Nsty88/zMZlwSEwlQDMDldz1zWf
8iPKFZc7ExlzQU4FIe+ZbXcF07xyz+TBkjdSOXgm/8RggitBxXEtjUGelKYymefR
6ij7Yo45bZfhd6S4lYl9dLfJ5b+bjHO0m7kiMUIKuD+i149AAxF+EGjYYUvNJnyU
30Sz8sbkBBJ9V8VjcQ2RkR2gyVNL6i5MTYYrfExKgMCZAjo/I6TRqvg9PuDvLHnz
GADwKkJvcTiZ+C0ECzq8d2Q6zGrDzfgGhnh4czJY33UT5wPxrPtGpJQgZEI2/luY
Yi8hJAEBXiLb3DRLRq0OgnLmC0Wdt9I1KeNR1o8PgsYgn+MhjMZFNQvO3DhB6is2
TcjcSp461l2XOmctpFMANJR97Z+dvAbW5ls4tMHU2nBkK75jbyGPcNJ6beHnqk64
mA5RJ5wOAh1riaU1j68IknL1Lhv4yd1JXo6HoewV5r0zsZCD6XFWRtSsBbSa0D4+
3ng71kctbrylg/dQq6a55UeUW1KQ/Xml2yxsN/TTp1+ZycUAekiPNz6zR9GxJXfh
wE5fC5KfQc7s2FG/NF7QMajSI6Qt+bpissvD0AMNWrGlEW0my9rWGCuDMjXLNAgk
IO5QEkrVd29Z91uABI9qbzIrvxiXVAcZpEjyh7zI9mkfGkmSxn1eAiFxpU5jZP1M
ftB0EI2Ey1Z/sO1IKnLpZt8gPJUXWqdhoF3Gb6tc09bLVOjq7lonyDO8HuVGmmL5
ejYRxQ8U6WhW1AILyAM1S29rYigVng3SC4q1FbH60cLIEwZsMYydO4M4R/143Fn+
d3JR5HXUNkw4I2tEkIOGucOLtO7k2PC1RNd2zVX8hxFJXQh/zYpZqsAK6R+M0Gbs
4Vs1cZEymmhZEynxE1g316yE885v1vVFxdS8aq303Y/b5uxe0D8d7P1NGXd6wR6q
4L39S4sQvkiZ164ev4ojesA6FuP0kweDGy5PwsAQTsU71v+xotpT0TDLvwJ2ssaz
wTs9Tgbmw5KWNjzm/dP3X60WAf/X7fSgI6nZGTyZY3azm+IVFxeOry4kvJNl9Ttm
qJfQB32BD9F2qOj3KIp+adgx3HJnQaieElwKZ+n80VPFMjInEseNPUCrOCjDeMMl
KvFPoF0q4RTUVEh2d/oz5z41wPZ/vj8MG54b12P+9BmjVI4s6fCi3cF6c4CqYS3y
EMFOyGEeFy8/LncoW4hsXD/KIvOrSgcOS0BK3MpUWAFb41CCMf3fsOUjR/u0o1RS
wO1/TYXQMl2iu5MvkqYcMrQ1O/b3/04EfOAVeRD4quFia4311ScrJ0vYdiGy88I7
BAXSiA4rwOj+RBpa4r26+K1tzh9X3FfJNov7A93LLzmjj24EeZyfCZSqf3K/YYiO
ZZIRR5FQuzI9suBplajsNckLrkHDRF5vjGBD3f/tSJ8jTOD663FWcWTlaOMBCSFf
gnzNOJ+YpuuyVxcgWfOAf53I8CpPZ26Tc79XzZ3tHuaCz821EdgKMWeho34crXv0
OEGpcYwu+rYJNdiXdzY7ltPdsXlyY0HsgG0OuXd4FyJeYG5VWUAZ/xkvrxSbKkDT
WHM7cMB/Zgexkcjh5epaU3mvBEVKnXyMo6k1zCr0hi3zprlgXMCnKQyHulMfzwnb
inm8NQa7jtyHZItOxC4bFkHXNq0+sSViJOxrW2eteYCEp/c8FO9b5JeZvkx41AqN
vk9KtYUvhvDQi6jfcXHHFZ//Enm8XeA/WRrcx2kKCV7ppWo1mZB+RnnORSFGTcey
6p9jR1TFflatn2P2QeweDxufVWD55+UgOOTUD++FVKf9Xua8hSGd+AiHD8F1Zr0L
zSlnA3LX5+grBm7z2bkIH+WRUO/m5zwn+gx5Li9gZpDRfseNuPOwDstnyYqb/R4L
0CAE1Hej67SqBz3bj7Jso9UfuF555nkaOxGRrPJYVDGDtmSpnXZca2Gpibm6rUmt
Uz4vl5h3aQebduh+vr7Pz9KHIyEzjfzqY5vP3fzU9AZrlYmTSrTRf2CZvfDjGvJi
sTy3u50J2/VFY/euiBQJRumS+8kt5VwCnnPqt3sRr/LwhVB4/kIXXU7+PgDzDmzw
wo6U4fP65VINFFVtK9HKcNhvn1LtP/W1EkLnAMkMxVh2Wm1LenQIh+71IkO2XrPq
VIJMjrt0LUEcvTKeX1MWP0LJzJ8hAzs3z89E82Wb59RDcutlRmNcWEHwg9kbkGAl
W92Pqnz+Z6CBv0RnlXNdxQIth5IwPNL7hfMhQoaIrOQFEButMHrs5tA22R01XU9d
vPMbpJUTVvnMNBySyaLhC7U6tOGkGXYr1FRVY0GP1qGtLwhkrCV2vXsg3iauAwJz
XgbZXdF1YoX1nzqt9iPvlWXkjfDlZC6PL7JGLVAKzBWQ9N7EBfrIAFT865PU5tO2
ukArzWYyEvJNYBxZRcw1rBA6HyrHpOkGbTIlyoYBlEopq5+p4JUpr8PBm50UccS/
0xyZ+sIE4kz/eK0cayTL3kSAjOrag79dHYwK4bvR5pXfqQ8Ph3KVxXdNSIGrqxah
Wz6la18C57Ac5EVgLcIYY0lGh2d8qd0BsPi/KQbvbZkPtbK4z1xLOHJAdy4/GTBx
d0oa8gqg+ND5MtK//3WiIVE7sUnwskXTQxQ0SSrNlXxBcL6CD75v0VXI22xXT+60
eOXaMKfHKWQ6FJmUOWxQYuGqCru5+68/+pGs9nNN7QW+KYPeDHWuqeEwjBwSdC/w
f0b4wDs+C4NuyEmv9zY/rOCOflmZZn1tdG1ZopL34dFzUSYwftMV0Ld42Yjp6lZK
11YoNAYDNsfXVQXkB4K1mHZS6514uhpjg/x+0DE+HJn3wBTZLMK1LJDM1YNRZd92
2l3xseJqSR4As/glhrH8AQQmCQsFo2x79Bw5oFafqOShPd2hASdKuhBABI7QI9SN
OUo8MfHkBVLWkf59aXFXNrf6oRrX+2cBvaPTvuiYJAJGTr79RJhQHhC9XNMFXjG0
5x1I/gVAuDIFZNeLphrIzAqpyyOplFd7eXmqB6NaGku4DgwJJoUDF2GyyHvIPgsg
UgpTzMTSWDkZ+YXd1bKCoLk8ywEv+IHvadHy5KvM/WENhYpuxjUFfPD+75LjHfnz
rn04rQVjJM6MZ83O5+J2om0c9XR9AgmcSsxlQK+/UcL/s3Fz9vXTeM1Y7/0kttmT
XLL0kz7NRbRSF7mFtgYzg0OF+ThfEh0ypRXhxHqs9+1wnkMdPQT9VTOPy2CPJsGi
NmYMrYigVkDkrgwWZ4rvFpNaAdBT9D5kolAyM3yg+dtgWeOdm2HmZehNuHFN6hPV
rolRU/WKBBlNr/G7vQD4OkqVpYD64twSDK4ydVkFl4fY24CSKrSwlaHkNHea5ge6
wvnWZmYnxKmYp22jtavdz7Z0Vck2rxo6DnLYmsKg7EmVG07rQJ6maRcD8p+K68Mi
MwgDk15140x+XWosVViU24K/DQhmika/nG67TZ6ucbiC6H96+w/7aPzBendlUClR
t1vmr1pZqtYMM1FJWGgZAsR7we7gx0/3eS/jDHi492PoVM0tmfkV+mYKwLvWEDeK
Pgb5F6pIa88z0wh7R/CnDj/LhaCUuc3bspdrafW/n8Kr5pNo1TOpyJI9MXqwd6b6
CXp04pMznSpJ+vLs3cL7BLOU1gQOcMIPwWn3leb9hDkStbCxSiagiEsUlwewmQgz
HiqmpgSTDebjaxY3payskYQnTXpwqc1qqSTUBKsAEeEPC6o4l69XjaUR4Mlut13D
/rGl0C7aVwBLucCaZyTlbhsNlxqfmRKVXCWahFx8Nn77DywHkXIlh/NRE9eppoBx
V76tXaqyxvByrvm65ysvKhTC1dw39n8YfA7PnxP3p+tTvujZWvu5pE5Xw6Jpska2
GV8dt7p8ZgHctqikLnRwjgFgvxTSkvq+6vjxxV+ITLhr2nvdl6DzzGKVygLZTKOq
Uo7LjFcN1Gl/FRb3VgKBbw6blIlJZUarhll68BcMZzNxyeZlFZsfHAmN5SjL2lC/
aB8x0jMmvqc94IubgZ6pR1P93FSFzkaJyb3/kCHIizt1+gjJGYX825LeB7XTw+vb
6d21JqflMrPnb9Oi9QxTnL0oSUgugMfSgcGxYRSyH+KCPbGCVjDslgcuyJ1Eqp5U
5/z7C4TJ0DTnMH9cP6FewoJvG2/t6hwESC3AKFK3TeJwYaZZLhCgZeMoIJzhqRAC
ECeyNGPKmRoQTXwbJ6e/6NAXfQewRqyebIW2kCSMiPow9NRfLmnfTs4/bj9jLxdP
R09QE567lNS++r1ZcoTUvVVFRfa3DaX+Ux263/6GmE60hhygxORwJ24WHGQkbHeg
KNAHGy3877JWDokXQt3g53KNBaZv6gOj0MPw8DGR4HRGxpDMSQY8pa+lsxxwtI6g
QCTNxsWQl9yfU/NbNc4AASPMSOKtubus8nsQ2Zak7bqGIOXEDJ7HYACT3ndZPT/N
6AEuQ++EmxlQKrnx6r6Qe1DHJMdEmJTGRF8tUuBgNAMGVZitk1eF9bSD88q4atAi
Maiwf4bs4PUfzjozP72oHT+4QOs7DixCHAIsmfvkWZNRRVAzePIhP4aSIqhOrM+z
9zMAN/6QJxUlai1EwmGN4TeCJNlKBZAt8KIuBiL+uWeMuxlK7yyMt5hKr32NTfUQ
+BOd2XGStELqwQ6kUg8Ku3hRjfUDUMopoHMu62lJBVwRjdJsFCGp/66D85Tkaecf
6YhDdsyHANPohNernCzS1dcHwv4cjBsLsjd14GuyE1lS0x/fhXd5Kn3sLzEb3h3x
uJ0RnYMlH9HJOMjOYfY6iRThfGSb0ieb+YWYzFd10VhoQ4t6PfHPr7Aj4Ia5hzkW
pUZywjQq3UOFG/ejwR511GsI7t/wSwwhvFu3BC3aQaJgpKDuBAttbmlEuhAj4ovJ
nIPalUv8XRMHZK5szRm5B04sN7dNGWygjc3+JjZWgaWC4ima46nyGqKg5OiMI73+
EU5XoRTXrs9MpniZy1ClXBUt/HOzMrvBBj/0UT6myknNR1icJiaqUaff98lT+g+E
b2bh7wxso74GAtDX+3rVWQDI4U4fkTnq2hDSeP4J7nDoDzhFy74kgnt8Ys0Bnrvc
hIfU9BxRw30PJdaA/wysY2i5vTrwPsXIg3ZsaZe5o422UyKJDhqoEMb0s+YokzZp
t4EZpxKlAUwdZJq6T1OeyE1hL8C0io1xJxfscXuoTmEZ+zA+gawOkTLrQObmXiNh
7sHRHazL0vS1JBh0cOcGNRJ00IvxFKQcgCreShGmERcjwjKueZ+6b/8vegd9YTeI
nsKfPT4MtsJ5hw03l/uscTr53FFWF38Cz+6dfNkxE7CTirGrZ1j/Wlio20FfjTMC
6agKp/9UUASbxxK01duYi3DJEE1BkKTdZMNvXnp218fztbKlL7afUmT0W/yd8vHV
IjdAhBYsmJgnUq3YEX99bhDRlN8fRLj+3hyrNOHAWqhZZBOzGzTOUfUtrk5sPKoZ
ojdRXJplr9O87Yn+r3TwqY+njrAGjUwQe9jTGm+EDAX7x3uJXxRDclFAc4NmcjgN
efr7UguRlEettGP00uTHOZnTGjrNb+gG4575lODTIiI3O/bqJFRgfgCGfEMRvn4h
6iujBcf0s4kz7SOeMjSBv2iC70vOjSe0ZJp/lcFhQAUd3XUT28SJweeuCtgvedr6
9d6DPdSVRyDNEO5jFCHpWpR//uiBKNUu0BTF/mBS3DHzCO1yPY6YsV70MaeLvGyE
T78GZOtFw2yPsy7QGO7GRe4yHpfYos8jAUwxlW6IwDnThQ4d4sDCMcJG1y90BQiW
FbKYzgy+eCRnBc6f408k2fMux/kH/m86nLN4RGMrn0qyUlKZpIm8H6GVyutTLL8X
iR9Y/XY7yh2oqvH0NxXQa+MLS1t88gw1mj4gI5S0eFlNcbminbiQaTHGTvOI5veW
z1JiijkEbpxkxtBK39zqXtpIxUZfkbysTnkcngdxTct6qPUtat4veL0+352po41d
PkWaMW9z788WK4/nPMFusSFw2dOhJuQjrkZIcxe029tu2poFH9N25Z39XzOGj7hX
Ln7PyiiGFjD1TGXj27qi+rWHRzYG4ZFxLYin7H7CfGe0FFdJ3MHyslg2ae/WtWno
yb14iPKJ7VZ7WqjwJM6wtRovLb+5zs6LvZojcQvqAzGFajizxiZLXoBsJIwHSvf6
OLHbCSmwYLTxzF5DLZx7WQYlwpql1IAMe2EriO9Gw3M1ThrfA9Sb+pv+atde+90F
QMBiihyEbABZ7OBr3iPdMUD0Dy+4aGO4CPLIOaYeAymQgCgASOiSxeUalHfJpsWL
zafdwAzlkpclIgaM40jkoWH3j2EsLvYCrFk8UuunCCn/PT0fnTPdmaEC1hi4pBCG
t836fZ1koqXJWrTUBdywrCPZLpUyK9+4TAN4gDBYjw6/5SmHRv6E2JFunHzkBZQA
w7ZCzZ/gXInNks5PvAL7guTlGoCzyWpxrMlt4ohRKHE6kXWFFCWI5aS2cxnojICy
muz4Lpt8n7M4m7xWtC296HSDbodr0QQ3Z6QqF7nvdK2j66jqQ0vk159ICfqvQwcw
zxWQHHYAU1kBkkqvWdTYyBcL3M7tpvSINlKHSLdb4Fn9U+B6O+455AkqfEKYu8D1
DLaFN4y9KmC61/CjYmLtbyen4QmSFBMiERpDSz8GeOKv7o3oK8jSGH1HDLWRGTxt
E8It++sqVgjlfuD1nPzRnxCmoe2Zu0QOw8H/rgWSABMcUdMap0SnRaRI5cS0K5CH
nvyZqgHaHh8rO0N9aLJxr4VIQaKfBF9d9kuAVS8O3yunYU2ZeLm2HU1fmX+xrFmM
UnzxH13K6Bl/sN6bafKykjXMVn5lkjklH7NR7BlqPd9omYAkXbovv82wCtI9+0np
kMogmZR0nPuVSOBNe48ZB8Nhf76Rsb/saNj8hDWVODdf//6kUC4IlGaIfbJCV8b1
9eoe/ILxbHPSnpEIQkeUfyIZkTkSRFBoWCm6i5vxcbIPDsdxGdpmTU1nCLFyKHoj
zCEL2q6PSjYeTpwftrY6FdsaO0p6jwQQZsCaycrezQUjp4+M2t0v1Yeax9MPBkJ0
8Ywrp8KqGJJAuUdX39osL2MnlivAyziQULpN0oZB+XvRveFOeG03glboakTmur20
RsK3bNlWh877i8znq1quaG7TWGTmnNlTuedxJAf0RRVRU/yRgrFKmvlScHHfUMBS
HAI9qtU4/haN8NHQd+U6GlmHh51W105vv5vB3rdxsmoXnxjLt9opmr1ZZaiDSFCJ
Zwcykmvmz9KgWZwd0AjeS+cy1BkFp0+acrdvQoPJq1408LeDaCcZgEHud7EpY+6/
WjISNF2JqRXrc3oWp4fM3/uAoe43yQWD+LfnVr6Ttjz8pP1SC48VGIiXxxsQFp6J
ZY97kisC3ApjBu/rG4jPBucu8WirVWDsFZx4UMkFQysTH92graRiBwV0H7Yo65sQ
rPrSYbfJbbplpqkanjVpOMk/BvQKOUqo7P8Ncun3mvOPDUHyr3JsVLsuhIRVOrR+
E4+0c8GDn93PnnP9yCG1dd3+bEyZcMrwgHLUeNqXnM+B3Cdxbl04p55WNPUU3J90
sJhhJJA07WBNlBY+tOuRpHlLRfzRAUzrKKcvX/4PhzuudbDmakunvwlamFB0Z2b1
vTQe7/azpzC+iia7Hk+72oqqKjO6YVyfZW+HKCNo9x0HuGxII1zmKJdWUaw0dQQF
1Faw+7ElcJXR4c4m6x+VgmkoDsEmlQbLaiAwQg/eu1J1Eog7hu1SQG40qbdAUkJF
STwARUc+Rfp5dYEvaZkqep+ibRiMr5/hGFcYQlP9uePVCiprmewUJAa9wuL+TXAe
dYfby9sSBD+XnNXjRiy9DjOEn4krWCLcJ0qOXyOJJ7P2R8llMgRg0XeihJCpqEzm
iTd3BqeIjk70JJR6mdV3+ZhbqJMzWsppxEagE01Hw2g90OzxZjwFYK8AyPh5Dx65
JAD0aCUM3Gx00kDk2wOJ0MHW1cfapV4VsApQ5Un2Mu6/1zvhOcKSR0JN2n6Aajec
HwJjwhBgU1CtMrtTa05XpExZlXVFWPsmENAJtrqlnAUPop6oOgu3bluXqO9k68/8
errNkRvS/Et7mZc8OfaqOgu2oygUKMyxDXAbARBsJW5tlhsgqrmOQV5w4oc3mJ6w
f3f5g9wQAai09V5dadCyWxOEG+0tPxeFxjEZwJcMwVQtmfDmWAadZgmsfGapVBkc
M7CDuJm1vi8cPVNc780NHsVUyayxq+L66x1i88bSy5hhhjvgE8IQ7JU7wXZOFFYI
Hdzev0i2I8QFazjjRw7LkBrcOGZO0AF0JJkq4Urd1UH+V/EBTK7UCUcxqq5iZtEO
uqPlPx7oXe3AlkQf9xfsgI5zLl7qXR3ukHGkTW3KM5Au+7U+cd61YRSXtNz7Rmh0
W/b/tk8Dk+hZ80mA4Gt9OjiEHP3Y9SDUWkLYe8oi0kmtohuyHJSesTsoBqO5sxX+
W2laIx2LxnAKli4hgMzwgYR+xOBql8PqbYE3CG9uH+3tmkt/25G5pwundmNtyx+i
v3zo2W0QX2TxglrHkk4QsTbmkxwZ4lyLrDB+4iNv5B/u38FHGQK+O7D8uCXQURoL
mkh6QKWy64x7wRBkflcdZfqLtd86jhbWDQLP8hIWGbc5hQkGsj5xmAqtT3xNElIe
3H+RGKPmmC6YfOk8rYfWyE5Fpm1BsA6DPybOCXOURCDk7QNuCVqc1sA2TP1DPKT6
OIB+vPCszzcjJk3iUMq6y73vvQU10mNyYAmlaoZExWkW/j4c+LUPjw/b/rRwHer6
jI+PF/My2mOQijPjzcJNkZEwEx5d8WIWYUQYgUym+o+FT41TL2Og6KAFs+Ra2/ma
l/Ts4WTjgSyC3Yqmjya6dipm95ZScSoY4f4F7rqrN22TSRK3qjCRadfvNvUteIvS
v+8dSAIwtNGnNsJqfrDd9rcGteVnvoGEOJXMDLU1+7C45pjRUwKweozxQiMEUYt8
Z/wag802sLNzdBfrJxr8oH8Z8CssxjPf6CsK5QJsYwSc9o5kwmU6NZFVe9qLGsVk
LYTLAD6Ry9MANTnT6JFC16oMh2iI6Yc1vdiT8nh+NFsaBKsBxOIuZEK35WGCrR1M
vOgQSXpF2G6HQo2AQaCRQAtdOae00Lopnp7Wh9NplVQDVibV3itg1MBH6r68PqHm
XgcZOyhtztW0hrH1xlqsabgCceIP9Zv8EHN7vBhC0+yh+BXetUFoGJhwTut3ScXB
34qjd3s2MmXi0iR8NZAgo2rPBdtVu0NwDap+q7maEu7wGjc5RcbRYXn325b4seV0
8kvjrTx8pripLY8vrX+fWYtNpZaJQCWWcJViEA4/jcS65Gva3bFuADGIHN8eFRgp
gwlWq7mKwoj4O72N3fAn1L1I+dxEKc+1zJYO3Rl+1vRTonQkMb5gJiFQY/acj3O+
VvSFzaCgufxWEdpVgddscnsZHc5bdIV532rWxnfCh7HdDvwWA2jt5rq5tNJm9Ng/
7IZhCz63zD1ggR8cOuDzTrhl+IKspezR7VOU9Suq7VGHxCVjAX+FWT/7ZOfiHrUh
Xd5cz/Q7JAF7cNDb4P1c7G5KKLxQZP13AYvCyj4L2ctUTUsRv7h5Au81KqtAzEOt
oCbY459ds2XS+nTEB0NJQeTPQlG4Fcwj9GUVRwzMAVHgKNnYQ60s190Qu7RaJ38k
FUOxrRmzT21eeqTnWHd33j3VxkPhB2hgqh9JEQVOIBuWTJy7L24b2nwLyOl+Gwhz
lYD6PuA9FtGCHYGHKf2THOH4mPaGYqP0ahHtHJuQXeBIHs/P6aXWUPNhrpVtpHtT
BG+8UT+rRmAQ3diK4DU1WxFIDcsCgmLdvpVfqB7Mp5KICMaXDLCePT6z3ijaT1+O
IDxDoE/NQ/Ov48LMhETnS43NVa3xclit+Z/ywlvwM68R0MLvBgE6R2V6rtbpO3Hl
Qc7Mek2zygKUMvtpNprL5lTX5nCYPh1i+FAE4UTbDIdL0Svh7QxoVL/4sABna1dp
bYtfmXVh0yQONTDpLDTu6PRBF6Z+vBQ30kZXzhqAHOnpUiWBdT5dndHeKskHRoFT
`protect END_PROTECTED
