`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ilAuNGfgyuvpawSH3d8o2yBNuRSnUUrF58GO7agh6E/nIKojlWeMOtGtbl6IS9k8
PK0l0oalPPCIwxZUdEhibm57fpbhLQIAcuPhYinBDf1WjKQkEEOReFybfRI50lyS
FzqtMBygLQaDjqlaDpgpEZN+a4IwpVt8jukV1IhBF/bu6RUe2kXXczFaBzsi1r/6
dczWxM1d+sdZ0+iLSxf6nSCCQKmdbi1druTt972qZnpP8AtXpBq05wHcprdpdd2S
ENAJUc6rq6FodB9zhEucC0kXXCk207ACwmgH7zyYfwH4IVEM4eTiSFrOZSN7vzDa
kjrS581k31od6wKdcrTUxIEdMiv90hEYApbwcl+WluMP5AyvWBOhAC09QEDGXH9T
k5TluX7tbCYiOUkqfqsAmJ1K0Mx4zlVYIGMWgRegJ6y+Y2Lo2RyR+9cb1U2/ELgj
y47vcCemFEhBdvcgbWeeQlKeQUCdeNZQNAefvJTiP1dKKv6o1b7WvX4FG6Wpdh09
9nPF/kTtlr2jYGsKqVvBr4MFJUAlN4XK5kiMnoS4EBJ/9/Uk6K96jLSeQYi5+75+
8AOy2XhHMI79KZjJiDI2ltpsk0WOwu1ZsseqThdkVqSl7tAFsaOe/n8CJSGZiLHq
do4lkofyXyC04Z86EI6b4QvKkvMKbHxPsJpujL92Tv9j1apt2K04IoS3pmYltYp2
Ej8lHpXcK4m/fuNQnaD7fZ8+2PdhSDBD0noJ/m6VXOGBK/6xjVtBWMAx+ghFJPbR
eIhmBYILL/6rarRJhQEvhVd5aBK7ZT4uxCpF3yH+Nh1j7hUWnqcVXasKDwBB7KR4
pftkJLXQGNkSg9A42TA5sNQNLRy3LY5gzAistTJKA8mjtK8gxRYRO/8gCrVrMFEF
4EjbwS4IY+4wUmUixmi7n8kWVzM4k36Vvcwgs16riFgLiaK+HKjJUWKFjDoA9+zV
WdUAN/d7sBGMEd0IhgKeZvr3FOAi/nuNnmxHOvD5lWAVIpSy029GC8cLy3TeVeHj
SLyCQL8df1NGjhCm92cI3XQ3JBEzydQ6L04HYpWYrVfJhtRhzZsc67UnGOQQulbv
EogBtPPi5e3Uj8l+u6jvxvrsVLTKYHUekAWNiBCU3Vmt3iWetQPQ1S9J3CZvUyRp
OH1j1GjNx/fz4F/D8StXEKw7gdNgIYAs9LowDn7usHS4dB0NiUxYbfNwzplLW4sM
`protect END_PROTECTED
