`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
X0h1lTkZshtj5aRTe2aTIKNYRnq6aDzYh6AnwyFfeKBYmBcZBYzjbbXUPgtDTm6+
9ZapMuhV49MaxkxoXidz1CRfaaayl6fSG16xDVBbtoeNlC4YGG1omFwn/bOlOdGX
tqCMmCVBd11hZsN97C4WcJr9XISdGdCM0JiO6efGduY2MFdJmCAagEva/Br/N1Ul
nOoOHuRaoTTKc6tA5PxZYN7XYMVlSn+Ar2CPcqT+QsaaSbNkx+TxETsn6PmkOz8H
Jab20qcxyDVkdFHUuA0BAFN4btR8JFyeqFnufjTJle1GmSdC77T3/a7Dr+4FGYIL
XDl0iIlF3LBviOYh8u/PjFt2Ln1hWBBWVQdtMDAJI++DidGinjpVw+QdDgONpZ1r
qjfn3VtXRa9DoXbL5nHwfvKdYxFMKFlV2BlabOHzpPa9Sh9yndDm46YolIxFYqiq
hLRLIPQr7mbipIZgcjCXYN0nwmspspu490OYVJl6z8uaHslj4UuoIr4ljFcHCsTM
Sxny4M+pkOQr+FxU+2yOBpfa9myn1PDUYn9EvzbZdjXr2UxOY63UMQ62L7Wv1zuZ
+m4j5PcQq0bKJ7Pe/7MDovBgqi5zgVKPf+stmqqy4IyaZ5xDyHMt8q9lll0/nyOU
7JnChPe6VU5/6etAfB5Wskeje5CSDn974B6rIN6+oGNr/pEciz+KxaF2iGI8Ohq+
EN5hyzpS5qq5q8Y29i/BgMSQB3ArTg6H4bO9r3//1DXNXfBgjCD5l4lM639Ur+Qx
qD9pAzxIPqO4U8LrqdetHPGsrH1xf/KuMGBLBvYNw0H0C1H/RA7WDk5nFXgXXVQp
QjxFWYPmB24bMk9cfH82/LDDJIEO7fugr+8wV6tDJw46ChQhnVCkFcCIT5ybE8j0
wwp6kLn5myv1jmi0f/EGwm6U3PCeqhODmUegFRbFt4+Au2WnzTpYxo2HbhdlWbTP
BVF+cKiyja0GxKnKiMMATmU7R1nduvAUBA4xZEa0rz3H06zuDHVvn/q+sZiVvvBu
j1MTZphF2bJUH8iM7/UKq1Gj44Dvw82vPptKg9HbWq/1EGgCskok/RuA7zN1vR2X
FIzzOLZzJzJ36o60DO75yHEL6Ti0qTNzNGCJ9hUb040UBgyKFJH6sNet5DvrrFjS
3/jf/7nntlCoBOMy8ntnZDmgGV04lVk5RPCUrkUdB+myAcCZI+vG77l+eJiSVXTd
jq3kaVFxBCuiPzzGXEsBkYWJaIEz7RJJF0FRtXQ4PNqBbWEvh9Mpuy8YpK/ltwVb
p0ua5EQkuyKzK8GC6tNK95RK4I+FUv4wA7nv8Hf54aTPJsw/ak327OP0w3o+SMEo
wYLJwlM0HEhfmswy7M+ZHnagOnQRSigVIhycGq8FaOaVWcvrJJKebACGEOMUFzfo
sM/OBP32M7zWVXOhGfgv3+t9ck9esYqzgaiwsHlbgHwXsrdovBHIbHLiDqd9sLTq
p8Qv5ZBZUBm8ADnN1JPqGHDA7zgXUAziXnkOgNNqIcR8+neXZHk7+3QHzTqxcB0H
QVEI1n14wwN19S9/U7HP76BdpHVWh4Fkc3Kyqzg4VTlEzU0N16eyMHWfPMPmobOW
S0niiN9EFtFDIhSln+5QNqtmx3vElfVFzt+l1QpO4rBKElhXECldVkzFRL5c+n5c
7aMMh8xAmzT2N2Q8pNUwAV0TGltzIX6LVub4UE4Gy47PGXZ/mzLo2Reb2IIjt8XL
MrHQVUSLXTfGzcSAPLOop69QeP6N3f82DMK/MaNuicuKqxZmtd5PJp07YEwrMrTb
2iMmMZgDLF4Wn/PBPBHpsaXnoNwNpNz18AbzAIKB8NYIZDFfg+6ugBLcuSKJ7/jo
Nk5IwKPYAkTWLm0s9LMsX2vAnjBl8RVaQYw/+2kjMiXHLmZHWKjg/eELLJgYLPoz
6hpcKuDBdisdmzHt7PrILIPgQWj3orAJd/5iW1vwlqyz9N61hOof1tBa67G1sCyC
zGU8ea5knAXBsw530OJ6CZdQqpC59WjCJcgU4imLt6rJBpCVf4Os/Vr7ZcUXHG+p
vV6kCGZ545BpNy1W0ED40OkAX9q6GKJRDMWk4WQ+NqjuogLIKIMK7Msu395G0SVm
k6rn72bIhtXRfABnr28X6ZcVWkaF9SoHVchgO8DWRoVS7STQyhU2TI9BHGPSxbDN
af9jiv8+GbrQUkKJPydhok684GnMYCSMvX2rK1+t0vL8xgrX0FhLDVZ4ynoTlRLK
1OzfrBPSbmdmKwglYKLbxcGRuqTEGvB//bGeADDAPKkmDPfe9QWNqIUq33sxwi7S
l2ASymuUPSlqyDaK89xCrxJSWlcmTg9ogpGXOgotJwry7yf30LKgcE14fwmvPINI
GT2NVT+i6PMRQZwb+hKPXVMx/kb8/ERzy+vJSF30q0xuUn5VyrQqiEtIkuUJUTBE
WZvMxN/yzfpwilgzBjPtdddPXs/TStGZcS+/Zy4BC50fPxyYGrhL9+WUiPklY5IJ
ohTgFdzKFV3JwjPfBbOGQV9UwL6KwtLgzkshWbnV1emCOmrPsu5bUjURVO4wpg5J
dp4rg5sV99qBVkgGXuCmKhsdiHP43R6U1PO7JwqGF1TOQ8zSqVbVP0XMXPLWe3Mj
qJWmClnpSjBHHSU31mfvpJ38x+Ckol/la7xUcFdywjPnu9JYcLAyczkC/YPnjih9
1atCElfvmkQEAwN07csPHL1jy+yBxeM5HDhSTTbQdw+2sMY5jApRs0Kgd9WEOJji
peeK3Vritvjpu4Lm5MxkBBum3DypLv3ezQhCxt1DVcStWzxOFJei6wV10593gCRM
9v8PkZk3QHd4wplBvrRwnINKvv4bYrLnnyGKDJk4Lyyhu9mAS4QmI95g7msG74rE
dprJSDPyYZujIOhl45p1vm9sMgGuryV6JeEWTUyH6YPXypBo+S0n4tNkf+N19vXq
w+5fzZ5u2YqcOjxbJ/hm93uX6M4GCdYT5mhyPw3FJ1ABP/yV5/pl5jSDVMwWzTsv
7KjtH006CTIBjuLPvUvc1/Mgbpjv8yHtEAPWwemkm6v1n364DKGEilcRH3XlZ8kd
gf/VeBhDT29TdJ44wF5Fn1LVGjH71mxK1whLwjnWWdqOfnq5edweWNKgIKLhCaFb
xbXOV9TfRL8cREWiQXYNTDiyNT83wrjcdGZugPMf2eoSRjkThE8UkQmIE+Sy5dMV
XJyQ8c9WWvOCAZ1g+mV6AEri0HBoIDDncC+0OHxc0b5s+5Fyj8rrKNQMmdRNKzpe
Wj6wv9IxzEMuv7GBqWPYHoCku7y8Wepj1vaX4v0UVJ4n0ORYx1OMlTv4bRHn2lA0
m2giTcYhcvBe+JaKM4Y7rsGoeNrtZ44svvQDK/3r7/lS4eEOhcippi8/qQ6JHF5N
9Gfnw5rR2+qw8873gHizWJfR2XbTWLAM9Tmf4J+4DFqJvvWBb5/LXtS2OKO2uj1E
UWUSeJ27CTYDieniTDvz1+ftLEP+AynyhX0aexBu7NaAKTF8Nc2hqMBP1MHpZV9a
vhECaTzVZ73ibTR+c+eXhguE6Z3Hm2czYLM6rHUg6E7YIHThj6AadxiiJY7TuPls
eNKcBVGn3EB/LETYu9DG3eYQwisLrgksvWqYHAtLlJArZeNmdm1OtWfNT21HIyPg
ApndggaexWfJ5YAgRps6LRPpgyOYJLkIdvKPOA1/KV1XcTgsKGf5k8LRSOsdp22V
MzJbv+pgfWgp7FpRgT6v48vGN52pJJhT9BPBqaSXaNnqlbSKcHN/mKQkk76v0iyf
ZI9NFyQHCSFqMVKMSFS5toMEpLvyxPWZwDzrK4/rwjJqcBGyAsq/H8agUYmhm3Sr
yRC2Je165XIjpmk8StZ9iqCNUt9d2yIAqrvqZIl5iIhfbXN7a7e+5cBGrMX+3Q/v
7UWJyvDcdHY7+FTyuUYcoV4WeYs+vLfauLdIrMh8GPsq49uwD7rRFyF5d75SZBJT
lXucFPseuU3DbbYfz+NPEtyjpEu467SThbuGaG8VGABREamEv+TNOh6RS83DY+th
5dgW291/nTuIZk+fKqD0fUljmMjgnr3mtRmTNp4eK5WK2zfh4wfNib0fFTgjBxsC
1rVJi/4gYqK2Eu1FhalMQ0xbNBRzevY70deSv11bFzxVwRqITjntUMeqKAO+FwE8
+sVyjvRB4JnxNwlBj2Dps7xiID21jdYuXFG8XV7v48jGXZmbc4FzWeMltdq0yKok
w+KEBcAJ/j6cQhfJcSHcc6i5Djg1wYEmuAAr11vs8J7DxAw/MLqU3/0hz9Z7B4HP
y/i2rCZPOER4cU0SdkfdTuqIgiTp+bl5UYTS3VaZechDQ394a8XEbycqxhPw3JHA
AbWZInDQ8mYW4c8GpQIKba5S08lOEGTan+odsriIqfMd9wQ7EtM6ioQeJAYU1FVe
udWfLUJkN1eRlX4ybDcBJ2fNkukniBCTv6mWnd6yTFuesRM+ZYbXOsC+Wgco8TJf
6xM+o+SezO2k7B8gnagif7f6KWwfM5FXU17UEPJ/+/kD3DggbHwTt0YCO1+oy9el
xcc5W1pehLN5URPM+Ef5wCyeBNCqR/06u3pyuqIJ3suUGUtkZMHlkiQLoY1JUuZ/
laGbB5M6mpkcMyD15tfv6snDIFcuUf6DyeZXcuDvT+shJaFjmM6oIQvF1/Blg/KM
TrTqmCw0dAYFdNsd5AbCmsBPIvvA0Xm6qaQCDANnAY7vzLgRRCucK4XAWYN0eI8i
A4ckeRyPJqOnYPr0gn5jZMex+E9sIVlUR0VwZv7KFTvPsUZe32gf1owK6jkvAr2q
3o7AoTAOuQG884c4NUWJxjxPn56v9bpXJDEbafs6ZTZLQByniTBkyYV9SAKseoCh
Jz1867KOUlqqXoHGAECd38V40NbNLWPP7akYY2A0DGsk5ECghTxZnDjn/fo+K1Kv
lr7cBK8qBMnXM4oT5AEqkKqrB0WycYqCXCY1o/8s0vf+HzxgFxM2BwzuVNOlaEf9
+3JZcdDWbDHZdnITEs7n1htiSEKWQ8GsonZu27xssz82bYA2uRrQXE4l9Qtwfvxx
0J3aCvJw7OZmznG6o9yWz+FC8qLFrQvrH6ncYZa2fU1/0n6IYkE3RlhXZyZI1GTu
QceShmbgLYej5nk7zgX1S796OP2YzNYLtuFfDDpXz7vSQ+2lAhk4dGB264q0Xt4o
6rliOgQxYgQKw+yihyulN+EGlUvPAZhquhiUvx8jyAIE5aPz6ivrjqTMJBdzEKdJ
6qmvL3PXd9mHtrpZ0a9HcKE6/zlqkQ9cWuhchqB+Ti90qWfipOG5v7Bo2GOvC5AY
UdN285ZDHzsKndkF5gxy/B85iV8Mce1iEkX4NaUQSpJRW/G2QUpaBpzQjrgAZoqO
1v2UOlzOkKKm+PxWZ3K+V25TVWwkk+9RJhSMNN58IOhUSi5Sx4lAyen2P1C2nkLB
ls8OUiyKHJcjoy+H5JhCCV2eZ19+2umSeeBp0ZQJUq+XM5Q9GYszf+4nON61R2w3
+HWTAN9Zng6h/bkt5wwvatuEcfBMr1J+BMaUksxmd58=
`protect END_PROTECTED
