`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
H4HKPiqOMPSDehFyB53nkRXmnfvp25KNy7xfQdt+r9Z0SFbyuv6H/ZUlRV17Kooj
whEIPE3qdURlx/txLNfOLJJvJtx8AMMNk2bLTBTP5sK5b711p2iU5zIywbKkp5n7
tT5Ek09hMbGvdFNCBpAiuCuLgftRsF1ZcQe8T8h72ybtBDNY6xV9DrNCOY4h2H8u
JrUIRl1deeVT9N89oKIVL2fmSefK+AiM/tusuosmv190tTkRx4DCMB9a2HHn6Xn4
SnXJmKqZwNcFBjRo5YRcSznv6PwjkuiMVpt7sipLwYerGUMFSRjWidLsxp0f6Ip/
rIgOVAtRcsQVt6xmhw0cupdZBU1Lf7HJp/lmbjhMGLZrAaxafzxrfAPRsSebF13K
gTQcGl3JRw/oxaaGkNRrfuNbUXX5FW3+BaKcN2l9jINwVSRN2KXnnQSUQYinl6v/
3J2sFVE3OTINRjLezyUjBi6iNTab2jPCmyX4h8OWJbwJF40WWv2mhg7SDYR9PQ5h
1fXXzOPKsiUjh92dRJY75u3dfjwokpHJpfVrUNdLBF8iQ8ImLsUvaklI6SGI4sUL
9SLsAeZev/R3de+MgNFMzIwIoZO+4zo3EYqKHpjfqYUWEiQ7XQ4mJjEZ2Pq/sSj8
vbXJWoWb3r1xJ6aMSiARIWkY/KhfOy797QrertljTuK4KS4fGkDLXh2umqDVw9w9
/8Vj+fiEEB2GSAammU4Q96NEnHgLW+dScyX7fYqwOAzEZuLHQMS6VZ3yfg8jWA7V
ZAdxZfO+7E2iW8oj3ujVrFkUyJ4L69LjmhmMaSPsS+zW/79E+0c0VFqqaHiEA5XX
eFb73vFaXes0UcQHPejhJvXZQOBqTllfV+nCa/Gna/byWZvuABojmYDKpUXrBI2N
FrhC6IHdcmwVe1YZ9zp4M6/n5K0YMD33ICAkkKC1aNUvFU+32daAhBHebmWieLU4
0LR36gMnBTOdLjxxdg2yq+SeY7LRf/Y+CZLUZk2WnmM6gaqrRzYbnYgvD1shlUPD
2F1zIbx8RTIY4rzo7rnB3J0+F1P+1resyKRBtiMZt7lj9qmXidmQW5fxPTldXZ5x
DxbFrQxPK6eAevl+TBXk3VZWB9SDJDQJMdJNgw0btX4x2IsBdmIoRob3pZaTkUZI
qxhkwG/WcclJYLgh6M25U/1+YyRpne6xZq3FhQMhibAfF4RFFbAUJW7pYKs7R2xg
ePku/YwQGqlhci7GfUF044gV+icy9lrt9c84ankQmd8MehTYl+9hJPLN4fq/DHXO
g0yAlSkS76t0dCy1QXvQdZi738eynZpgPnPaZNZJTOQfyZNHMBc7OYo3aqxsCDdb
boNPDd7DntuhE2/aN9340HEOcq/dHFeQZQIIkqSd7f6nZjpMMdTZW7aSy4wFAeGP
VhNYMosxJWvLWb8OwykOSYrtGQNu8SNrS+1JnYyZRh/GLbbJp7ILi2d/P04In2ZJ
Td9tM1pyROPHNRNDAyWj3DM5zx6A9aGNOmV3nLd892NXeDAhf9Rtp99tGmFSxysh
0FCEl23qc0Yv8HI7MRJVT7wNB3e6axbC4kdcH3nEshEKkGtcBW8aNWGfthMma4Qa
q/Ayfzgj3UQaF7MsGb1F5rXkCnz26o24ZrFhdnVhSvUG42eWula8AwqHVxDZglLj
olXY6NVvy94Lsm6a35ZrUHntxm01pjcsiKNscRMS9YUff4728V8jWYoQshGzlghq
7xmkss7jAUEXE+uvSF7hHYS383zj+xTk3atuX950yAlKNr5qkKt4wNbqiWUkDUIF
LEow/Ft4apsEWGilmOD24WviISbG+IQ+0Z6srndITBFLybbG9cJfRxxrpDFc9Tev
ecTNTV495eQOZrpwALTnzXY4SMdYSv9RYBAowTHkU0IdKnzBlWgJLELsB7UQOFs6
dXgIN/z23r726Ys2UaiiUxks3kJw4drjeuuDE2Wa193+WGkEFoW8iR3gVRVEEttT
9kS3dEHmZT5TV8wc/VIAbh77N8rRjHKgZHOyhMrk0fwswzqUvNyRzWO14DbHMfs6
WO86hYDDeqEunIVLhAHsy1U/pJVy6V5a2hRRoGdpdOosJcP6CZL5X9ivQ2+VhE4b
O299OWhYjgshUU5hSr2PPbQReigG+kQayUqF+hd+UDxx6koKzWI01JXe+eSpzJs4
xr5KldclLvIkLJSJVzH+WFJBABdYgKwcLR+HUZBd4UGUA19onZ/azD+qxQ9TeKJC
ZjFy4IW6pfsV2ChJPlCNqMc3mWSDf5qy0y140lpZPg+Dj6maxjRH+aRfVHCBp9de
ELg/Bgm0+1NdDTc5tC8MyvllGzlv0xpXzoHIr5ows3mGrZaUmPaEHpk8idBLcaQE
m85XWYe4jj2AV5oTLzxwms8vt0HTESsFVRcccDL1FeWz8NogMj/uOZJ/AcqkOPAF
8KdP06Se/PpLC231pcit6IVsNLlsCvmqhQXSYO8ywuC18jVb4H77F8LkwXaAtjYA
THXEImtobvsznudPnJCMpkVHW84aeYFFY3fw4IA3eL1YEliAslyWXOts6+1Cu+Jb
Ag2ZHk+MY0d/lveA886VLX15JpNQciDOPCcBp36d3sLgsgOuP0H3SQwmDfkzKMzF
FqOFl+NPwLcn36ADTXftSDR2HEFE1pzPguczpShwL1YeueCc2GTTGKTRoJEgJ1pc
erPNm63c4pRb0LRVNiXXqUihatbiIeMcUl06e7LuOwCdDr7//TAmst/iuljC/1Sl
J7bW538WI61Yii3j5z6HgLTyHvDSHnRktgQYJA21v7nDBC6UWYSYfS4LhWBI0NU+
wGgt1VL5rrk2hBLmBJ8E+erAJMxGUTVqnrGc3et0ZYoWBDYW0716+03mVXB92Aqc
Yb679FDbJBOc3IWThBuTDKRuFzhKkHjjt5sPTX4gCcFgJEgGjTjsAYqQJ8xi/lY4
iKYl+F4JRSLSpzULkDPf1jElh2Wsj4YCb/xYrmpcX1zybfI2hMQKJbq0dXcNAg1q
aqFr30Ija+h0dQVqugaHF0HLqpAda3nXBDLhV2GzUOWYj+hY3WhMM6xxJBXZZwG3
2607Kk2nYKjtPwGud2L/gYfKM+qRaFXejasu85Wb3xnQPKRRPPYR+DUeJLMX5RaW
lnKkTQbpaf7/dXePTZGLK0HwwubVhVuKk32YzFMPxIlDWRD7mf7UduMB14Mw5f3M
wKeggCzEmc1cW499AX/G66calzMe50GMcL41CUJbJoyrD3yKDtgDeXIJcCtuIih6
CdX0wXR3UoE+u2VVQYTtKS1V6VdDanOFtTPSx5PIfnvU4AFdRiMc1peewpvYNIhg
f+wNYh6RDEQP6ZGA/6Ze5N4dh0xsX8Y3A/qqri228lMX/N8++CogXMu0pobOJlAW
TN7aej/mHFWeZeTvahQGZHLzylkOfu4lkQHSRUrmL3/Og+AnRIuapLZ+fgOQwbJD
CQVtyENYRlPuevYvfQnptYjaowK3nG1AxFTnLfFcR7AHLmcvQ0Pb1ChdO+gnvu6N
Glui/NkcD7/0AqkqEgNjQMzW+iWtRpNKYNLi6N4ZL2YmPfCyCYpBRs+dJ5kOyZqV
Zj7qqGHFJOBxN7ir5bDmUWnWN3fhetNFWML4XZCjDkcBEIfUbFmXebQGWAhYJh9v
CqYmimMHfBVdcxt9pxl54aJ4ApDVHqj8w1NIL6up3B1FoUUQ5PQE2ijN2v51Wz68
Fk6R5vbqPAOzRMxPcPTuz156XJ+7iZxh49G9205xLaPMHLoQAfOHboruWXBPCDsD
wjy+KmN/GWDnLqRx2NujJhTyJ2n1Zlq0iCmXnzakNwMfPqN3u2ygDjNTV2ExkMf5
whmsGtu7wqhvCuuF0UjhTmmHK4kBjGcune+4824S8FpSpHJ9QsybAQjX0XCzjCIL
J4XEb2oCqC7ysabJrfWUpsrviv9RP7xyGlYjzCkU0nihqZQqV+kEbw5UgRbNSV+w
ijcNV8bMzZCKj6odNpTiS0LPSvpPyTyT/edg/vuRlSjFC1bko/nLWKGsYF4j4Ki5
uoHCSfbTzPazxfmfHj6TaLohfwJH7XX8ZVOaQy/LxqTcJPEDpf2UaoyCID0raEGr
pdkwTHGKQp2Aiv+EYUrfwu40d5EI6YepsM5pidgBmepUQqmN/vbtunV+/sguXSRC
lYts32yqQZUl9rzlFsreDUxuD/aakVItmwshu7XFKg4NUVe6Bj9CUEIBoLZ5oCEr
+qYZkpQzqMFyfnsKFS3JAkkRkhMUjZHc8wsSm1bhKq8o8e+DP8GU7lbBEpo0bu+x
Wgz55GvALsK/RgmIxsP0n25+cfkTp+C4Si9knCSTCldRA2IoUyT8zPTT6y3urdmj
X240TPoQaxbTP2mputin8WfV8WB+kKGcqxbUeyG3a2cFgmFwmru0F5nP3jmVPqIW
nUc/lulw11WFaPSZqMhlFvDzjy1XNalcDC3ZwQkb6tiMlugoTop38OW+bfyOQS4E
wwN0Aan/1Y+vSthVEMsmxCecblogE+Q6BHlp46wephMbng79rhfvWQRckPDWUsl+
qb0BF2HLtMdx0vzoqNcigir/yJKWRlu/qINIA4ZHs7a2yfrcG9F9mzud/jaRd+zp
MhqvovKxK5Fx8Na11RFxVPzayDZ5jSE6IioxvgRqK6xc6K0o1Hw7Mejxca73+znK
InAo9+Nnms3mDMObq/MAaNX3a8Qn4raMEpCnoLuC1zgcUxcz8/Oj+aZ3rnEUtwTk
DHW5sgqhFuHSS0hSRJN2vrAtcX3smvoY1EDNqNVneiuBWg4yRDVALvQIPL1TXwq7
Pzsx/rSkLRxkGMaZBJPnZws5ik+S++Rp1n88rGGPh4miKY576gQimAZ1JgSjlnSG
KImGU1MGXd/eey4qnwzmRxVaNS00KKS6RoG2ifxnmmooueuBmHAM+kbON8Q+E6Ms
0kzMvv/EQVftE4nzjZb3LQQDEshNiQ4ift+vzivP9NIT8onfohKdizwSh6zc7FYw
xfePQD0+O/l2J9aWdP/q6LD8EMGeIoK8BqfBLdfsMMtgUXUBZya3EhgQSE2M6/Cq
yqEnxn607s5EUa0Q6u+zeYZSv0dj+duBDYMn06CHg6JzFX5Jw7krct1NpTp15aCE
ibNTRobIagvHUJO7XTBbM6NkHnWhRj4fj+T/8KvG2MZN+gcbsEiNbOSaKpEk3Gs/
4pL+9Ez0MdW3jQSiK22Wtk36OwfE87bmMmACyGa21wn7BLM3QIwwnsykTWBdyoRh
iXiFgFz+ujRaRljjKgOriZy/e41bbcv3ZwoCFRgUP6C5hrOvwepSMDCle8f/Hmx1
+eCbVBtlbTiuwfUitZBNkfXjq8nPTeUHcPsffF2sUwR+1Uufug64TK/LbGiLg2SE
kMg7JL+ngCkkSybyiEAMj++cjdMfHRl33pC84+ikHkOn+MMBI+Ik66f4kTcT4os+
g8QJchT4YJ+o7hAG7zswVxthTBJSG4cjz++DMRVGmN7EffJwYeAPPmqJ3Ldut+fG
rmPnEWk6zNuj0lf8JVqnkZrUWxpBNSDd5yZdv0t7h6MEZgOfcnkbCLvR1vvYPiEJ
Gy3vyH1dfBRIoR0ufcpO5PwWo3T2zMZaerjJCSdOlA2rif/104P6iagwnYudzD2A
Upe8pHUtjPg93AdhRryWkg==
`protect END_PROTECTED
