`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
V9I8YJnurBgJp/vsdm9KCUd0PIFarrgBgt4hGJkCDGj4d0CqTdtG4XWsIqXSPuKi
RjnzOsRIfL87XIY8GK/MSvnlrRBaF+MqwtxQYaQgWGGZ31UPVEMPDXoT40qC9q9p
n1K2NvqeH6vNGi/XKkpbWt0s0r9OmXCvzUEdCb4ZbJEDyOk2trsfg2iiNxyzq4Q1
qTUhe+ABmaHbw//X711h+z7X5260VmBgbM6XHrMHPuAfE6QKbj6XWyg8xBs+KeNC
HFOVaJ24XbkJnr4Zbr2VfSvxZJVxWeSfXgPKvTCNeKA6URT/bIFCP/IGl+bx2Qu8
+42qXfD1GyPjh9r7FnFYFS6EFEbqWpGTTNn5blG4LWATL99zIix3ONutWkPMn6/O
`protect END_PROTECTED
