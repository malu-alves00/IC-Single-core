`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PfbVcZUUCLEhYg0ZWlerKx05pGBcOByQEhMQXzggnGw1GqfC97NIMmwwxM4H+oVp
4zSz9vhi1sIQvUS9YneE1USnX6eFioxevlo8ovUeI2KkrkVbby9ZRqYeMzoQGEuj
pPafW7cM5WQD12vvrZrWjXitTtJOT+PT8ORCb+Hy1J/6GiiN8w62X0QD5wuFhroz
/q+FEEV0QRJKA+4AFZaaQM2hW7nN2ofN+Tg2nAZp0oS3tWg9L3fCy1i33JRn72XC
cU+kIbdIObX0hI8ZdmmYSlvq7MXh3DFmYOv2M7OcDg2bc9TcZMVkFjhH1OFR5G4g
BXKqn0z1rVmLfnuGU8eEoYRI2FMTdj31xw8yPspLxibKnt+aAtW+EyK2oeg72Ms0
9FxXdWtZlCbCvtl55YsTcC3p0gsQeIFVwE8DTLpaRLM9RNuOIgUWTw23l/bog5Ge
IVrl6JhhYHERAKSq9gqSprz44OGmmwjTnxb7lQwLeWroPGKO+zb/eodtD01pLiaz
mauUq0/8l0RtC++xqPtCd2DAFL5E8wO0gEao3No7JsBtRdFysfQ7xYLq4bBWBG+q
nzxnvP7pg4e2nnAn5h5U8LwBszRDhdNXvdC7Q6Ve06z3MCxtt6WwYfXYygSp1QbN
QS01eabl61Sr7ex1Vu7toCVPrWWLPlTBZCqzVZwnUVPwjpM/0RJSrvFpgOGQ185V
skBT+Z6Lhq17yqV2MPPUhqi0FdVn5kM0WG/7Xz9QYHPwZnD/dy2gUEeq4RAV1kUS
b0M7qWsJ2mOcfYleK8ey5JAi65Jy8Jrl7j6GLW1hE8x8OM7JfI/v3pJgssHrfdOn
DOmx6pZ8COQOgZc8qF0nWiRgg0NF6T7KJt3fQai6QL5ZlvMXJbPETcqClsXG3GRN
`protect END_PROTECTED
