`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Dhq7oVDoXuGqavJNVPtu7WJDCeV4NOvFLjmx96tjkDIDOwfKxRzmQvjHSdpWQESP
PkPWjGDi0fdQlUHpR4Ep/Mn1/UYKT6PyagChqER8cyV1X0V3CC5u7s8vk6BsOVUF
PNqrCehxuFhNIRpBoupHqEJzUZogIP0dl55ARclaq/xpaQiXSXW0bNq/070/Yi2+
yPuX3aoAgQHn+V+98+EHi2x0Hfq9s+UoGDEyCJZqjcQI2Mo8f93hcFuThl7jpTAW
jKu82j94J0ClxwCe1sNy7aHMiFiyuGYrpj5SioxnIXf5BjeK7XVFh/pR3nCKIbyC
mFGqzYgOAu6lbqpaHtXWvkjRJev6mrqtdV7BEWHLt2mygEZ3agE8DwJlJDUiqeED
mP2qVimyhzqv6TrB8VSYnDbONxs295xop3EX0sOmDvU+VejUC9SBm2r6KB7Ssfsi
e0XBhm1caZIWLh5q4s63u94r1BuN5+Rj8hzA1u7IAe8qqtAi7s1h7x/bgxJy/sQz
/NGIQFgUw9dAHnhkaR5cDC/ZU17GjibjBG/XXJ2IF2TVWcMRIuUhbX4D+F1OmOS2
/1rQ/y9GfiltNoEPyd52aG3/YSMn05Iakf6byneBzsTdIfvEFTKZuA7o8MHuUhDM
sVJXlD7hsJMn5D1ug1RFvg9t7iw8dyeMJdyn7FgG/iLYiWq1MZ+CT/ww3TgPylpw
3kRMjf9BuGXi+lBB2NVu42cr8AwC/L/KMEbLll2P/5TAZz2ztHRqGFtxBho/gqal
Nt4907ZLmDCB18Oa00hxrq7rVGX3ZpymtzqsuXkiW41Dgpyqnr0Evf5YPygTjfjZ
kMxN4IZXdLzAAkY+13W2pihOjv9JBdrlCV1y0ACIxZJ24fMluLJoOAo95oIe7kBP
584xoubFK5K/J9t+ZyUvlLf4fMsUtZeCI+qvNczjz2kYQJaQvBGwLIwUu/mpHLCo
THAaFwWmQbTvJxiJTxiib4eX1HzdNiJumKTaGBMAn8SJCDGvPe52cRmiQbp2yDvC
wLIo7dtDo5Xd7uNoDqQzwQ==
`protect END_PROTECTED
