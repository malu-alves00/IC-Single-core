`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bD2l4Z1JWBpAI68lZWkzs9Gj+EMcwigG9cCiPd8Yfu4nINo2APkspe3o0h/QCMyB
J5mWBFVezYEUy7zZM8qDuL4LyJ37R6BGC3fLetb23Dt9kkiR8mRqAwsB+u+6jlK7
UCgzIcUsG1SVlKOHb/soaS3PMyv2zaqtBdy0ygnjMhebZVR3RldR8eRlBYaX4Z+y
awS51zDd/IiY9Huxr034/L5XaQsu5B6fC/qNug0aGLlD3kTHzCvSXu7oKjK7tDpf
Sb0AfAUyOigqFALhZyOhintDtdrbMlZJAaxEk7bChMs6RchBdt4MV5SOgBfo9o02
895K7VshE0zZ61JGGOpJJSO/jZqF782vW9lKlAcfQdgIzQYSFj7n5vDju2FV3UFy
5sLxcr6pzQUpQ69ZrYTjAA9yI/xlrSLmlf939QbR5GXwwA5ZHySeWNa4O7seygfU
ODg8Zs/TQ/aITUOdjBciAzpmF6SfTwI4af7JpmNCa6Gz13b1PdWeARNjXo93l2/n
TPbofwkOVVlSzHoe/Ip2WE7EzIJw7vmcXiuf1+aIyDb+uw5BrwylApYQJHRObHFA
RlLYWzy9Up8DINNRzooSQEYv68BQPKpSKmVxYRd91hYeVWX80H9+kZUQ4mCKa5ze
ND9GQ6hqPn78LCePj0eZga1xjOZnDemXplKXODXTBexl7IGGCDEK89aiBGTlzwgs
EXjGPqKouKMRC00VJ+uepLcEv6wM4+WiE7qERjSbEyEZExSNn3ahvwpR2sBA7FVU
X/nvT8/IHRF6SG86eeQM2x2/4a/IlyDxgREO4NH77dJSvQVtJRsRyAW7JNM3asbP
NlJMVFpuowbBwUQITQp7ekJCRTgcRt8/B/Vnp1rAkdogfwETCOiETqubj8Eafsst
Acqziraf1ezhLHVVpoWl0vsu8sTRfk6rg9+X7TSF+4qujAfP+2uktOgZeKKd3W7N
y88y/jlC8vsOdBCpW5Fe1TUQUEM1RrOs9onz6LjX61dY4Mh3TwWCS0wLqQYMU55I
SX2si2vagKe9zi04zsPVRnmwvwBQ0ymEuxFAFAU/MfB8f8R/hproG0d7QIEncoP8
QQJoJcrLJKIF3D8psZ+MB+WjqdKex0C4GDGea8LYh3T51yGMltG/m4ffShOjZ28e
464Cn02Bnxu3m5OsyPAOU0omE3oLZR6eZtcVlJ/3tgAuIXVNzrWNgNqu956xn2u8
HiF7GiLWyuKVjjH451ioXlhesUph44ibUV70XMJumTraDLUZSErucWR2yQsmLRgR
oAnPY6GGOdtOC0PhCH1znjHoSAmvH2QTzb8cXE9jBN6vfSQUiG57A6x7KclTB+8M
k1FluFuO7GrvpKCk9qgfOrKcsD0loTqBf5pKaMmXI79lZmdVY07v4Z+RgJWQ/sGS
pxSyfyk5vBi8xEU0n/GOag3WC5KQ02mEXbt50ZWV/Cz3hMGPRVyPLVHrjd5zPsge
w6Qr+uJ9OeWhf4BqsZY5PI0cLYrzqfmYNqLJVVSc95ajN92YrQWFN2oCOGgqN4bE
i5k8R0yTmdBF29Sc3tbk7dbQ2/aF2g8cZ8GyihBJVRIISGiWGW/DL26Yw0niUVc1
3RyaMmnB1u+INq4NV9eHN39g3ejNQznZc6D9Ai0olQPb5VKFmiB6kJzrHWCMwXYY
Poqo6s60Kggl1X8Xr24Cl7VGe3wA4gPylO3DKDruaYM1XBVE/WdHRo2YsL7Q4X8G
PasgDPMcteT/BuloHpS28Y0TRS3Tl03q7s4IDHmYhhalycT23A/Bzvgs8kXY05pB
wl90hTYvmlyeD2FCa6lcix6mS8KX08ordvs5Ib9hkPeR5YWfbuf/Ke+DQoKMd2Rz
1MEbZQB2tisyYVxVmM0S6bsEV7eHTWje1fbEaBldAg+wd5BJJgquZuUfzP/OtIBY
bJVR9SDwFiNfPdet+c+cqFxHcrjw0p1w2VoC8qRBgCTcShHwwfmqMNCmDOd4yqNu
0AF7w1yMVUpoNh9001q8uxHyQNIVzy+8+dSsI9QQ2pT9Jqy1woLvGyq3VRug8Asi
OVrDFTmyEKB2dTB/ke8sP8w2M8Q/0DDmXMouidPIwK2zfmjAxF4KxnGAnjLxrW6Q
CgH4AfoVUb6M8mc+zy2UXVbendibxlSLo1kiyW4YBtr7p457kCZX/hbbAQbyVwBI
UwPBpvcRCXjsOeQ89XKLle/H3aqz2C7HnhFRVxpB/9HO0yC/9DljfC3GeNIXGxl0
DnGcbyI3ZXpJfJ+IFax3OYCwQUROfuGuy7JwivC1B3dAr4l+OMZX4YRVup9E8t69
JCwuT49SK9zKxrSsnP3e8rxivUJTSf4LtlI8W4a9j1nAukQgAsILtKK6fdpwY+JJ
D6tPWILZoefWY2ebyBpVizxeNsnoSCCsFqYupB0PUOHVq5+XY/+dQ1esZOtj41mm
abtWqHpN4hcjlZFVJMHOVK8O8WdFE1CaUXcuJNhlbtjb378y1Bw9sOkrXevDZS1/
rwSv5mF1rldiX6ol3o34BozWnpI/qm3a/pSs6dxql1qTDYWaFFAmldEwmQIt9iHE
IIuOpW4nBtZozETxC52Rt3ro+CDiO5wh04aB5FmbtcZgi1s6W4sTOb7NxeFinX3q
A1NGyJwWKJd/BtdEeaseoTmTiFl///ZUORZPHIH/s46iMCIZLZ6kv1yXhzDzN6wt
Q23qGkGxAh/P6I/XFyVix9fnmNLSEintmfDgpa7bbX97adUBO80RaJVhrmgv/PRh
CvAvVQ4K6mpq7hyUWjE7IVD74mYISCFHjYtwDi/jyRSjZ45SlkEuDzNJ9+fcCZK3
pzDRCtt+lk1qd/HMr8i1/ivXCz2/+CJGYyyT6GFg0IrdO48GTGGSCFvPtqt8dLnL
xpvw7jnRnrnKbfi4bhlHAfW2JtBoJwl+WUPC8FovdPfYsD2Zw0PcbAGlGK8b3Abb
DBawtJFL25RgokKqz0szFImpvNxH3pG7rF+MEFidEarMCV1nlNd8RjCG8AKFxpm+
wlzsEMp99gsbsuIwe2e4B6TEI7J/rXC0KO0D68ZmOAjqj+agaeqSPWXgAiWix1Yj
Vm7QisckTwWvrKJ9jqM6i25G1dxKnRcXbJgruf1Ad43uFuRo1PJyspZfsxW607Dt
kJ7nHN7WlisGN5SCjP+iSlBzQHW60McieHVWoUotW3QnRXQuG1iVoPoqzVp6nf/9
gS9urmKqeoA1YjnUFL9K05wCYBeqltGzFe+S6hPTtUFfBh86Y7S101APNCdISjf2
NAPwEx8xj73gak022LDZZMr1rhJMcWkAwAbNEKr+YDK6hcDFvFK+GVBRLG706Aem
uPU4hGLFJLbH47r2IKaf8AxOL/8ehNG7wJjhpxU/EC8iPO721MHvkDQU1GalT7ri
QYB/0cgWZOB1YK5GTOtWo012X2ALxg0aJb/vZfDRstW6j/jH8qu6sDGh5jBSJ48P
z0iQM9kQP9iyVwhY9j1VB68IVLRENIAVrAjvQVXCjRG/48cikFkDLT1UM1wySooE
aHcz3WDoSM1chQvNRD7Er9ovWekHykTDkHUau/BNdImKc110T1l4a5Zkt9WhepdK
bD57zhSxvh8z0OobLX8GD5K5G5aHlxAqIXbH5s/kVJxYAEGDEzj2rFGgOKiYzdt3
xRcIn87f1dTnUmuG1O4qqSqWHWCHkUEvR1Qbod9vINez9mEsK1lltbmWkRHSd+Il
QXo+wKKw7l2MbBNyzyV4+1GzDYnOPX+TEORC68OZtJ2nzAt9OgIWWINWTj1aWfw9
zafwpafQF+CxVV4CsA1Ba09HIMzpYnGCEPfyzjWPBaUhwkjJgeVFSIjnyTQ5Cqed
gnzWNdOx4ClyvRDiWdThwu9Da11mE7sYL1qia69k+RewHsenJ7YBfmO44d6Kb5rZ
8AD1+9DE/UgQSscrRTX3FCamsXt7XEwnUQ66oOapMw3x9XCAK18fmSp+Piu8BKHs
P8k5LxE4rgn70dGzUDTQPAFnq/VcEQUaACkl3SksZgEQMuBLbd3axTzMgnMItauZ
bl/qS1E0eFGuBVBzo7OS0LcDPwVa5v0nYiZG/ix3JHUardtvaCPdpMVAbwC/9LVA
Td3zqpaU9nJuzK0Ty7auL4SdaSA7spEjBfL3wt0WeF0w8c2HjFscA85QWAfQtgyM
Dx+fNRwMjWCUGqZmK0iRUAoA4NIx2ZRmDPn9AXEs3J3roUWhB91NqIX4pWn3Welx
rb3IEIQoErclx5q/xspKdfgATmazlOoCrxlH8SyQk6126OQGFe4u49w2tGMiQu9F
8bm4NSz6FAvOFB7hlr2Q/ZKPFnO+h4Uo/jf1+ci3tjLZjhY3kxuX407ooOkLEQOE
ZET3iY+YEsjT3pLXf7ThIE0+wEvodwSKGG6WyylnwiWLnnGUnXt3h0eLGrhMtsa/
PPiH/+CTMXYzCHPrsdEkI9ZJgnfI2IayhL4H09zT212G16xe/K4+QqB0ByMvrXJB
wDo8PF2Y75pQRVzoLDRHThJ2lMsrMzZV2KdKI9UfDtgxHx4S8ug2radjn30chs9g
yXeIbN/MDyhZygRJGd+ilqrwPC2qLs75QXPT1vg96ilx06S6JBvcyYMzO5zbfEn2
4HtALzLBmf5ZPhBJ2accR4nUkVPpKVGKAop2WqqG4WWcP78ttSgYYRyT5hQNOoZw
pwQVcqD0ptFfjoFe6G6Ap0haUpN21xuQlgelToBKT2GKECO4uhxU0zoK+47E2Y68
hPwHBD4p7iglV98ImDawlwtLbQP2Bx7Iz/gvm7P6hu0psHpRal1SYIpifpXKijCi
HfztclUzRoh7cTnhBGRkaY8GRT1pvlThS8whrB0juVxF0lqZeArDM06wCblBqEIo
2wYoq3WF0srm1VGtZcxzaYofhTYljAukuaAWkixTk95vMdp1v15r8DeDA6a4IRbk
6cM4TIWfxbb0k9IgTvW4aOGHFUatqTsVPmaA3jNpDEvlAEJZdmriCxMS5Z2OI/1Y
+wnqX3+ZP0qPVkcZiEgtWBLyzvQFGqaUDFClKwhi9Im0ue+PmZLQrN9tWBSl1Y7C
pueEuQGzsW9+/HEVeCKBVG4raTuCj6CRc+8PbWW+Y2uFwGa7ETuFrOZML04NDXns
1pjNCIW2zdOmXwWiJ1dWjj54P6zqaKnIKrIpRxWw8IryV9Z/r8KmL32njyt14k4x
SsbC9E8IP0eEmc8eLQ54VOWfITcwK44yS9+vs3hcUyBFUb3O72h/ZnqbUgOK2Lyo
Umet7GzbYBoQywlIgNMyL38ggBEU4mgLwDHz5hxejqICCGjNB8gZXmTYRr1xWV1x
aobZIeV5f/lwIv820dmdjco52dnfydNPtU7OKPWgFP+ZO6UHI2S56baOqWl7OUR0
rUhI6hpjxsXRKsoBMZrQ5HpuwuJbz7svl26Ur+kwTJu047zu9xf6nBx+bXbsSSpU
Ogx3nb9gjeOXo7MdJQszOQ==
`protect END_PROTECTED
