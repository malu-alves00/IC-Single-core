`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BN/KwM1//znFmx86oALYqKBDqZHaWpib6UfknGkI31eTbWXdBW8WUV9IQi9A3w1p
CRrWtF5WmFAmj7oL4YUDZRbHlVMM9wn4kztz2vIuFj/hRiwCfsz5iW3DOzgg1ZoS
FdInnYIXhaaiNn/IIi8LXhtIlnkCZ+mxRzw6bUsjW1v0eys3aeDaUm51M8+8eL8m
a+VWoyMyFEWE7NHRpkYd8DHmLQGbJAUfDgfWc6dshMppTdoLD0vJjSccPqsgq/9u
6ZoyMb56dQCC0/LCGcv6CDPmtQarobbkQnVZDDyPMlogykbnuJTvbv8B0Re3k0Cb
66uSy2o4DgXx121kFWV+Ch8csQVkZgSn43a23Vpfr8iJ2rYjD5jEAh86lpU/7yXA
iRis19T8wTVdb1T1jmP2R361poV5nZpr7Mh6sRBAqYMdJLagNqR5y3jvjTFSAvAf
g3UnaC2tNhdzB9Rn8Op9VVxDi4rNdHa8lItvnXlSLIKtkm6z8zpE5CafOguHa+XG
EshRoW2vFMX9+paCzgXkKC7v17qDFsyyL6GzYkU9njEMCjmbs0PwZufB6EUfqgGO
mPU0J4Q3tFJZKaTENxMZOE7vB2N87peuM6DBa5BDUSxAZ16JzbxbegUwSofgNDd4
YR3pG8doPXRbLNJVOrE+Jv2tIiX9FrQ3jlkdqKJhlhpfDvWv5I2DjcEXQ7GYDgAm
QGnuke5dUBvG6S0JupbGopzTZuqOagjQGpDu3V0Doh9w4QuJHERkBfSpUH1X77kp
X0/0F1K8+85ahFMreqC5hpabfXWPFxmMteOJE3XE28t8BqLC1bgYzim6sVB0tmon
7PjZLt7uLdPR2ZW+ZW+d1LWudQuF8kEbcOcBw4AxN9+KqfaE+bnQJFS8e02J6Q6C
N6r24nThEC1XI5NqL23WzW1SmJ89lSvkVCHmzB92c4LG8qUeQwUoOelp3rite+0x
oZSnxYJdedRlJbBIJPCJxb+CEsXpfuqyAMA9AtNBj2kAKnCiRztm0f7289D8VnxD
0MI/+QjSmCMnuBxxL98hMpVAyp9Dk+ANldQwyroxWffaeKzRsb5bb28XSLqaMcZj
QYbSYp+Dbxzx0vu/7bJnyNj6nyMfx87wgRKBdfCUvdQuWtceGBEwqlFx+2ZKyiIw
YMoni8Nps/NPm63dW3Iv9ym5sCLbYEfe1zBoaWHdpeNbr9t9QcEyswuJPfXxzohh
mNmGHzyTtS8WtGieCEgSre2PQM4PJvbGPYHX+IqiATwmVkyUDiZ23vBtXSpkO951
W66YVUk3EvAfB+9/QXAXz81Q+DdwAAtnyt17VwEsxQPQX/bT4jtig/0ihjYHgQZC
T9dXEVKIex1XVjxlu0q7ZLfWLpN8kWWTUrxODAi14xLVQ7gx0temZeafrbSvHoNg
xXN3egbrZi6fZ/gMMTx3AhG0ZZPr2XQRDUHTALc1JTvneIrqPadsKLQu41UOSwHT
BCPCZMrGNhWNbl6DNV5ijFJRGStv8smEXxjaCfwuapWNaJQ2usv8ONdgi5562h96
jTnDQ9Qy9NQC/mivUZntm/yFHwZpcPmHGtn381gQ62/E3aVXwQSzNDQaK8XIejuv
glmkZB9dYEWk8LLjH6UfEl7uRERdbhCLUA6sgI+xR2LVBUEFmRBPKrh+Ic2Pv7sy
gvHLJasEB7z4qp50/2be1ErcnPZ42nlNhYvGSEHE11LAhE/AKby5O6hq8O6pDTmv
SmQD6/7ddf4nrsj1N4xs19ZzkY2oGNiqJhZzCavf19UWbxMh6X6Ap71xtL/HQW0r
KlgX8ndYBU7pk0iCJoZJ4Ozceh+qZSnEJZlhR6rPsfn/5PYgu9e16F+u07M0RtnA
70tvkmhdal/2fWdt5L/XprhXg7A5rZJmjHD1eBYj5RAuG8hSCgxL3oBURKtUxIiU
wh3LKN+CHc6dQFtXT7gAVZ8e036YyjHoXWl2J2aXhRG0sAKgothueePbzLFOza3q
rrdBRjyWYr6KOfXzxnEZHwH7orOUj53kknO5enrMKUKfEPq6moYC3sHW2bkbhZ/J
yiCOPSHIX7sqWzRCYUUU8q+z6Vw43P6CvPi0dfntfTwS8SIT4F9SVquK8t42jqpY
6CuGJVPvOL7QV7HaeQH9v7PlgHSWw7qxfpise3vgH+RU8E7mhXnhIgItzmoUoqXm
JNmor65JZErA/2OJ7guKbAjnJ19w0GJXNSXkhMDSrl6h2kYxiZ7T10G8Hs+ePC3W
k2PcgPtQ1COfHKwva9gPhR6ZGzrcSvea6BX/H+GpY1dh5aNHzVgqEHwx2eSSXV64
t7LF4dzK1wKb4zK6ZWV4cMJoCIB1O6PvbrAU7duUmdtHYgIxDmivBNKItEs0z7en
3JMEJTwNkF7POjcZhY3PFCo6JdCfH3q3aKYNfzje78Xz1uuuNP7xpc0hIkF+DvRI
4OFQvmLoib01o1J8s6euZWEGrbdceU0zVR0CP35+qYkr2nJT3xTTVkylHj9M3uJN
n+7vcuAxgJDYDaFcqEqYaVIn+O2kUUXCZq5NjTYPlA5lV5yz32O2TMD3oXqu/wBe
PO3V6RMDN68050AOyJtYPoyBNYUal0/yKiVTbhcz0r8BOLhut5BIHjVhAhwUiTUN
FUmev5z+ctdawE7O4gBD+DadKO8SJhJimqgUxqEN4PSmjL9LyhjKuAK3pHxA3eK/
dn5fek1Lg/C1+M+PlBRPMckQx7P75xntM3EBbe4I/41l+RiJlE/J/n5+b0TFwHcl
Pkpf5U3CSr1ifhgb84bZkvudqTMywAuLrTEkfJo0L8czOirWUyLCu49Ws3e+PwHP
FxF7dO9z9qcbPxx0Zh0Wx95bF5cBFVUh319l5fMy1hJ+w3sRlNHPBv3nqEVV6RkW
PkuZ+Sf5whtJDerh5EQneApqs+whjUBptXHSKy5ACaXHYk4UVlsOv5VHQY1DmNPi
UYq9RH6X2QVgbqeDH8iaGAnPyOt3W1f07GH/23WfYJo=
`protect END_PROTECTED
