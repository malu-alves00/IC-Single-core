`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
76q3dQZLWTsCD8mh+fVqYLnzgwEe+klFHQzaQS8f4G2szsbqZYHwaSVhovz7cjvH
cXpQl1MTlqGwiplW1jEN+aBjqfNT2hPH2C66kOezq0ZQ4I+b1P0OoutbT3iXfRKt
ITfL6ky+sS8uOwkxGQa3+uPQTw/KPTRfthIsY1881cBwgnXlG5k27/Cn48Uwx5m2
h4AEPx75V4PlIxwJCaaTzQZY0KIEf3HDfzGy73gWwLeAwdKznsveQG3AkB8myEub
5VL62XxX0+WjfADC4AShGb0pAu5f8/6+BW2pGnrZkR4VziJl5VE4NIZUArrntG5c
ULMwuupoxwoSQ7l+0yiYIgybHJjRnInx9JHR674LHRk/QRfspVDVCBFCqn3lP8wZ
eG78HIYjZBuME+KNr8vaTkVY4sV3EZkArrmNkUe9+P7Wpt+5ewrrDS3O5E60QqGk
PfFgr9XjSUOg1ma1AsWC2016J7Jj+y849QRnechssiM9yLvgMCtGwyGVUbn1pIef
AzXHi+cHeZ6NZFWHHg0sVfhU+8G9WMHxvFSsnHIlh2TF5xa1feWGLmpGWKwOVZEO
KC2n/tam/yBSXNQuhkVOimCD2eGYga2rZ2AG1BuDQr+1gjSiZjJEA/knLXNH/YwG
+IKYV9jdoiYkjGRGN5Fr1JH94Kt8Z5O4pf4YKWPiTk6YNT1ROwVF5mEciJ3X5HUh
xtd22SESRweP6a9SSShqqcNr2Tr99SkRBOvtnlYWDs8=
`protect END_PROTECTED
