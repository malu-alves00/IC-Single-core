`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
adU3h/janbbhKHURCpBYEawQyNljPTGKyOIRaaa2HIBzE7V4WCbObo8KFkHGHKgw
vwbG2lR7F26kmtFdENngmWi6VwV2YmBrlG5hPz31pw0An6yDmVrucX+bYqpEnNSA
rGL3BwzZz0UcyF4uRZNPcsvv8bfmwxr7tuv/Ye0twXFrjjAQa3D+9dQLUiYJl84A
`protect END_PROTECTED
