`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YNkH8CalMELzXXCTu6soJrxs0nqcGrwH1axwJ1vd9ulO6vFkEyxJucxLfu81F8YT
DzzobtxOudhXqizzJ4LVC5va4nvqUzrR/bDBwRYIwBOxDfuxy5HD6pJGY1KcAxsk
LFd0g6IbXIN49YsD9rUmufh8ZNOO0dSu23Y4wvldweC1+RXwsfJ5Lb1OHQv1PSEw
Kk47uQL3jhOknuj5UhEFrM+nHgF+D0blrT4ixt7dgwUcNjidnUatVc5mzslqiexZ
1Hf/bh41UJrguFRW/sukDwWcVWMJDGIQ4f/QxW8oEEhxtAO2DGQ3h5DEChmjbWlZ
EFUaItYrnXjZFEsOqL8bXECmP0IxVAfD4go0Cexj8fRDIrFztJentmimqtYziyHz
Sb74oRw1l0naauXyQriM+O30hZp5Y/XZLJs/E50TsiG4K2/W3dELp0vAqCIkIj+W
M2AlRZ9Cohqv21dlyeiYa7OfyZwGGKleo8iiZAnQSatBmkvOuvHL4K31+HwEnptp
MUxd1Qmkqll56LKcJ3mVT7o2DD7FvepdQJ9Htc5Pdl8kXr0kGWoAv5IKYMYRGxNA
5+EAKxNzTCT43Wuu3KARu+udvCJ1jEShvItm2lvbq5NEN9mKDEOFjlfL+6FbrVUo
jvgyD+Tj5xHHyEV/pYT4IngTax1XNTuONQ/lFHD3aK+9P2ulnLw3qsyTinfhdIUD
stSDkFXeElr7QWxQ6cbiEFa/QbZNtAvpxZ54YHZOb9KwamBRjPRFtHTh77zxdODp
FV0YfDyES9qjVH9oatLEwNdzOKQfj1a19+DRoHBp+F1ar8xpxyrl2m0FC4GK9VNj
vMBtUlDz2zLBsfTS9biUE+HbbPSS+g4hUfwtFi4owmUxtlkb3N+5fsgVOIUtb1gv
d06VgoYXp5o2nRXJj/TLb/fRK7lZuqbg93TVczaTU45Q5hcuISBKnn2i70HcMr9/
+BRr437avVELEm09jYK00xCURfbjQBpW6/+PXBQ59P3O5hfzJmCw4vWFDQJpGfWz
9OzQV8yBB0e6qbQgtdxgYhw3fM4SIHJqA5vs6x9TVEx9IHb0XinLQtzSo9rWrlW/
wXiLgeejYRgH7mLEsoGJBjhwt19cfF/vIyoGfRTrVQANNP0waB+MBKINVNHHVGD8
ZitD6dlZIrmWRo1Jt1qAeWlHfanM+NnPBN5RrsJq8MYFzOo0FCXxWTnVWJi3hmV2
kyb68/wCeAJ/3VpXdc5Y9jUAssn4cP/9Sv/1UHPhcBlL8l1xsP65Joedfgk07lZX
m9dBBxPdhQ/mQTsv21lIfztWwGWpPMZnKvbqVAoWr0voLwsN06s5zcETps1Z3hkz
vDgSD6M+viQdox2zZAtaX6/zBAK4Hy33nKiscKTs7IQnlZLJSQaJuDCbcwG1ON9P
Kdzmx3CrrdH//PylsfzVcMncNZH/jHzqcUru8GvQce+GYwVoRURwhRmabaZ8Eq2s
H/8N2Q18XM6GDclwBkKClnCDtkvZC5ATYYgMoEbPzKmE8lGarculLg6BK99OgNJq
QCLOJzKtXHF8I6+v90c9rqFHiXn3A4ghrCi0LAmm0b7lvXcmjxYyvqkZjQRMyTCH
5JnrlioJQuUSibzAoHusNsWQFhbeLEfgK3S617hlJWRnnnrFrLaSfUiJGhKpNVtF
xJo1Y+tw31UVSWbmfRbdHA==
`protect END_PROTECTED
