`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nFHiW5EHJ5kp2V2auZ9W804zJ/FlDOOD1z4/NCHklMcfU/riCVAIruty1zMMSvDH
LmvtfqbRksERAQtH9TQNRheIEfNbS8FLqYNbSkyl8N96X2dNn/a1t6+C1/p+p1hm
b+NroTS+dT129nDMOYnEsMh/pJLpLFRcd2oF/PRlA3thl/K5N2BaaiZIA8JbXme5
Dfp42038smw8XzdMRrr1V0jwq9zeiDPuA8tkeT2b8MteOCdiFkTgzE7TbEgzMlfP
iCnDZMPsCeAVkl/ypKaxSWFm1zmpvRwsY2hSMDOoCeOuWam5O9UoXlPQIjEFZXqa
inN7xxX1HpAnla4eC46ALAo+WQRSWZFC6Boj9Z+VxdyyO5mfpftjDnrkyaadaS95
AoltXN77CWNJ1huF62OOZJ+jxKTsl2NfmsCgtm8wp6qF9zbKju+n72gMnLcNzCfR
0vHnaLtxE/XBWvd+nB5FcdGUy7hE1ZZ6tf5xr8yvRdjoB/DNfMAS7wyHfuNI54Nk
i0RIs6NkgOYAWE9j9IxSaELz4qeSny7lCsUxcmSmV+O1GW6/ftZrw0W4t2qfOyaO
6CkXIFdMsLultnsEHgjn0C0iT3znufpCphg2fdRdw4cYcea04iTaXtgWmhpjW319
kE/p84gpxLRufNwFtyzmzLtk0paWSEClrkhIK8+sZjU7Dg3Ek+XfN+eKSm4p7xI/
`protect END_PROTECTED
