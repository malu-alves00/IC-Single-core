`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6rrgUmPfJYnEtc+iMUo882Va8i0yhXqR3y0y3iIVbFKT9bS28jDrPqxLq/DkgQ1s
wgUczzG/lq0bFK76trvLsKys/d1UKDw0HdsZZjTD6ZwZNXM/LIQkLdrYO6zxW3PD
TC8BbI8VTa/ZuET+ucv9HsrHmmeU+OjQcVw8lCi0cPpSmMT9aWk2H/74zq9FSNor
PL2dOJ3HFBS9LusJYxq1yMVeYn2GLgRoLZ1/LSBf6g+Mx6OLu3Ya/OGGktzIekND
RoiaWVL20VqeZkp0sv7IMP4F7Oqyq6AGyDopsBMXC3WTUqpoXkPVcqiaH73Wm2Hk
YNuARppg/PmppGqiyfaXVaAj4nfNI9zgTGFdN6MLiumkXOXuq93+ZvrS398XG/jc
faeo4kl4OFMgwZfoj9Y6xlzSeh82xF6peQt+TSORY4afRncUO6o1aLRTyc15Lodi
Lw2wdZvkdfiS2K0pAxw2ej5n+EdBoQ7JQDRIz9X3r18eFZb3plGs8SskIaRqKIXY
IQdE6ui5LRGvJIbuuDnKyBNBRgDGXe/DtHjWHQ4+sJNsxCIeauQ2xbp8bD//x/ze
B5xIAuIm+rHQkez/4IYb/KQQRppX5cGkttFN2nVqinj95qqPM0irMlkjIZjzw1YF
bjfWjMnBYFlA6E5u8doLwN+oCTL5RKJ0FZtg0NVp1Ru1J3s5/vGycmKO7cZLBMHP
/4WLKm6OzzzlqSl0XLPspCgrx8WGAwoazKfRCtuzMFScGiGrHHnnXnivlQXjh3ce
QK3DRd+dO6YoXpzav46roVpbZVd44kOzXy8UQK6ArsyqCX5owWftE6Y+D1amXz+E
pNYcm6AcRwgGFDZ2CE++kaTcxdV0p/3C64Gfu3C5BGXlmqHhvIu61XWGHJBp/52z
0666RXMVjfUcMfnmlbAOPzEA9Blj5SPMTcpv8Zv2OQa0YUOqKPbgvUTjMuPk7v9b
b1nG9vu29p78jpuGSjPo4/6+7cHWZmFKAMx+9dMyglxnvMXPhc2sHrMwPLU6u4jK
czfPKOKKkGAfQFdUI6E0iFAUumemToPTdEiD1EVGjeUH7H/tu+noRyu78nqaLshX
51N7NA1sQ0ToyYkaevYwEbmO0hYS8qEO4a5HAfuZ/zqxZkEtKis+b0A88oLaQuZt
SWmR3h0q/lb8jiDKeIZFE0wSsMCyyn7LvjP65kJhvsGSr9MhyRDyw4o2vZSGoaxp
A0LZGl44T2xKv5m3+TKq6gLRyIn1SM7StwXMJNxMNa9U3fTcGp24DMhxWjoeCG2d
wAX9F+RFlba5ItFX+aRYZ6Ng5fqc7KeuPWywqsdPaCU4N0PsOMJ5qbcMupeim+ro
KPEIRUcN1JeTzxZtE1pUA0y5md+TNsJXbG42effj6zkjlEuQR+VK5QZWe7Q/6tFZ
e8o0TszbgKJwOQ1Lqi1ngfZSl5kLEORWXcTSpsOQlTChWY8NBWfJWN75XI9hlyLJ
In65+HFt53sOyIJIkEbMfUCN724aPvdMIJ7INmxh04oljg4wVuWb4Mss8tWkhuvN
koGltPF+NwnKpSThweUSHlpKorvqTdCTDI/CSPSub5OWnry749T1/UO/bH+6SuKa
9VhrULY69DiCJ/r9LPL3GUTJdhaIv2pIosiBiJEnf32eOwY5X3LNckWsAtSyp/O0
CJkFrL1OoOFVMVx1kOsTRDs9Lr+gxL8XSdfytY0CtG1PxzcjEQgitJ9T1C8jrtPT
jjC8sWXtUXjdPlOQycJR+jggUn0jV1enNyJT50UpoDlJOv1C4MSAhg9zcGPchewh
XdOEpAw3pbnOUngx6aVkuDnv0eAI28P3L4WiH4DxkOqwP5VFLAD1wKBvoSWbCeMu
LIJBRS6Ell+yleI7cXvCmunDfO80ECiOengNkEvKgyxal/8Eyo007emiviY0da+V
djILBpcSCqpPfJyK+DdEsdpn7l3YRV/glawpMweGrTfd6GFVTBksWJKTfDAuqCT7
HvGAjngs5xiP3uD5Ytt1aCDbGWbbE5p4RbhXbhrMNab7jO/M3mAGAE2TIM3KQgBJ
hJLwTKJ+k+hXYFJ7BRbi8KbDtGZnLn4j+/nDzc4JIK5hgkTkNPMSzxIcsUFe5DJn
/jzxAIwyKw5AO8njd6ttDRJHgLEoAhADO9Au95z+ZfrdlmbgOmEggYaw3kzRTy0t
/BftuFiiR5U1jnFud+IG8wxh6+MQvmtbWWD0MHAVTjyGRY5mKWsEpV1erdHT63+r
1gtkNqgeZgEpoOA+AkhNbs+VJTVMD2nKHJMFgkWfAbsEqkuacLikRP5L9k8KbY0M
W77I0GMCyPgSyZqkF+KO1xXjTKCoXvFyyU0ujETPP2KHY7ebwqYt7RtPJUv3QrXs
FnYKIUWmkoIuPTx6Rx9ZA0aXJWwdO/UkDENIiBGJvhG4nU8NhqZML6TdLCFVTBoa
R+Q7qZ0AOQ8VsSF3m7lmn9zJLOHx810XltyiMd3X3LXSbqNCTJEbLbtdBjZbwzHB
2iQb+6hDUMj3KkWOPFBo744dInXt7S3yVlTIAUGW2D3rX6ejG9zN5+WwDG307gmv
E5BpS1Sau66Wkc4E6A0vjmbnS6WYR1Igqhk7Tu/DA1GPBr5Yt75nkMDtZ0mlsNKC
+Mk8Q5G3gj2nUFOveBj4dfCieRo8jJnRG73y5aDilbCzeZpGyxluJNObvP7cvxd3
bGFNdN/Qc09Nmo45RUYNN1VHWQ5j/alanb/xP+w8Ragbd3ujNhb9qMUHfNvf/F/O
CDtkBIXd6tVQbUTuwO592nuvbjC8aVlBDRgsLnGsAvFMPSTTuxyOD6Kw0SuyAEFJ
Z7nKdSbBKxuOnzE139W01A8FD0q9+cAovTXMGiSGTlwYBo3lrxrVpx9eeAC6P6J+
dCuL0rFHss3Pf7ab66VvKwUI5FULfv5wqKkzJe1OwYuHwvKaSIT5mvuP1PxdMjuC
bBkAgiOilG8cxBMTnbzb2+7KJQFVTT1dV1I04UpmrU2aN8O2jDNom2aVT0a16zqR
I4eSN15QdexU+aujwL0uIR49NJpJqyU85T3WSGPtYegylXURNY8K8j0K46XTyQWT
k54CqKu26hpjOvtMG5VZjY7ZgVhMGW48LKhgDR4m9HCWwKffHUGPFkCcq3fvY29F
FpuemsmedQaOCfHWvvAe45UgoFLIf2frGgJ7ZTIWveiP43B8i2sYw9TJQ2f5wohx
cbUPbMK7kyYC+GBdQe25wmoU07Q1r5OMGZ3Vcjw36qvPKdBmsvBoMT9jOWmUk5B3
lGrYxYHGTkeIEpT8DVckJ1uXFCuQSM8qVDdRT3S7L79XFL4uoXQNWAyerT8NI0n8
lbvwhE/OwqPIGaHsK7NrmAshE2VubIOZz5ZOx7vpXuVF28E3o7h1RFGRhJLnja6n
8qeF44sEanKhwr79agjkO+oOzAUComs7OazYHhM2WlffKxumgO4v5LeQfYDxsv9m
sZUm/Qv0l2JAyBfL+M760ssGfXXVwQWWdNvFUdOqGOUPV4lkudGtH+91u+4r+8Ts
PNUKIDu/gxOKPaJAUASZ3FIWujJwG90ghFClidYrK5lLqahbGWbSyHDoxoEqx116
WLSuYUzYBxsxRjKZpydrMPy9+OPFKUXJbf/LQS8MtGAa9SNpwjqN4dd8drhCEbts
A33irpxUW1Y7rdidw9YnxU18Z30V/BfQcJIxAuet3QeKCvGtK7Fa4TsRIfe7Ejzi
0mRf4vFj7AQyaIJYAZ/Z8wSbxLy+X+nbZYnBxW1VNzvC95N1r6czg+neNYwtFtaA
CKuk6fUS94MHbr0jNMtRkVBCNgjAWPdoPWRg9PDK7xZcEdCusieUVFspgKysQas4
eMdPcMDWy6tRn9XOT8L7G7pb5bi71YccJ/WDo2wYYWdI/ePoeXFtk9TD0MVoTeW2
Erdq5g9VgrxI8ZY4hvc7wVUI4RImPOt+Ux9kl9ZCXw6jefkMC5dNWGMC8D9KQmB/
2nef9ExQYVZyapAIZJHQpvODt9vMI4IUGNx7kKlF79pQRGpMS2kRyOpLfjgREet2
/sY6B/gIWHa3t0tw/qE68WAlbaUjwMHbgF3mw5sQ8Aix2UkIM8guxnQML4JNFGG3
h/R4dXAQK46NFwo3+SmmqtHLBtY6Eat4VZJSlJdD/nAYWwjt5p9d2BQOTg32QUxY
446Uqx8b5CwJlEWZMsEn/hv27nQNaVtt5DKBusGR/dAIF7aQiceoPUpCzFeFNBYB
oQxPLXW/SFoUqBS2bQj6waVTAMlHjEDHSjb+5NAYjHrVtbf8CulgVdi6mo/j9ycI
suwg7kXkpBu7ERpNexDfHJUXcahKaFXUJZMdSe8uQRtl9/fImc+HEWo4RVBDhBQk
ohWl4n8HP0/8hXRe/QTxUycyXqLfX48S0V0w5QVyYP5Lnllsb73IofZhYg6JPDZA
zvO45c4A95krZcwUSylWSin/4D1u1/X74FrQ+CHOb5PFdPbTwaYar+OaBZ6GpOC5
VXDYe07kQ+7ZCbXVS5e3A+VsrZZJRWpyZhQZm6jGeuI/G9lDGVcqDK40pJlTlVUk
vPmWxTw007NZW98jriJRmlRmvBZ+h/SlPSl1Mm0jQTO308whyWIpPJj2pliIwWgQ
ekW2XKzkrvg1NbxmAoJFVk/6yEFwapBOB2HqW4zY5fHYqaEZF9a79wNmdcs/bP2V
qGp+cRgLR4Xw+anIWO7j09Gv7DE4hvEsBFCySJ9ZC0DzCZ4I4b3g8zqdAV/C+Nqp
rCxUDlyPbzqG4JLIMeu2EPmth/aG2goBNtzVKBOXvDrLX4jk8F4RDIbx0SXJyysB
4eIYqxSTpv+Q9yosuRk+Y3vn0a4PyQNfh5yBVnJHQY5b39Ueda5QikqPJDGHPc+W
ZgXYMtnE9sc/v0yUabjYjdouHhFfAQo/Hv1lYc5duqEnPDtW+qT2iOQCCwNazLSM
NI3XTYg4zxUipnLSs/T54bRsAaqEKEjWAGhx98VZ/FVgB24bEAuivv4WcMkjqWW6
2d5sJ/EtuSobIwp5ZAyOUNTYXjeZRDOa0c8h0tq4R1KOLnXEKTh2sg/cnilNBmPb
L7fRFdt2E5EYDTp1HPBeEUGrAERtcAoU3YChHtM/2tXiJPIibRZL3jpyf0nhnap2
OhKoM0klclqmiIGDghFT/JjnRLaPOUBJQ/iE9iDlf80T3co4EpEJDKj0dGyjaVIQ
P+b9q1NWWFqsoOsypGeJk1K6jPH6Jzkoz/0k1oZlKFeUjD1NNYrnpXuXK8m3PLl5
aRc2UHWCMc7tmj8FmX7Kxk0U1vfbyPpPPKS783nOmeOfy44S1dAu5rtN+HM6uESa
YD8gF7JszAeOJXVraOCMOqyDEhd/65QsZgpXP9+hJxf8h7xARb1OkJImFodZmtG8
gvpnrT4ZT/1g26QHm3i9NKSsZMCI0/q0iScFwfNyRCXmTrO1ZfElLBEHCFAqegwr
PGYlHhh5zrudYJrkU1SEtOF25UCq/537zgFI1HdO4u6TqFQlexXipT82AyXdnXLd
TyjXs2BTf7R5BP20M1OoqR8l1pGrqDbFnK3GxG+qqcr7UKQhiLnio9IICOSdfNQI
3uCub60iAERtxNNl4MUJT+5uXCdJUptn6/DEi23Pm5JkW1ffZdIhD4DvCytxriZU
YZJIVjgH9oR0AL/b0WUc3xU+ct32pBCHFmTDCtQmx2KsgZMjz4aO7RDOMHzI2PN7
aeaCvlcUCc3QGoTWo0Kyi6jTR1HFWkr77QGOpy62ny9wgpGUHmF62LsK0j/Jcvy+
0WEhQ3ZDjM26HG0ZOaKDCWtkmeiKXHSPJqepjnxYtacKciNvRts7B+/lIeJuS8Sa
WFUZHPB5CD2dB0fLONqo2Cs7GpKa+lybdLH9WlBOYX4zEaafmnTtTQGQEqXy4zd3
ZAnC3eY8EihGaMcjY4Skc8nxGPZtQNl1zUezyv6+MrB4FHpMmH5M+oSrZ7FSWg6B
5v5+/rP+hwWZwpidkXEVg1qdi1yfxnTfcuuTdCWq0bdmccWRe5Z9F3UksYmqKy5P
zOxGQmHi0TectLL56TUFTPPDcfndkbWyAEqLgeir8r+9JAKUviBeIjWdpGhqYyLR
yu/XUsJN/t+T3dYHw687GO6vz0EtQGRNlCovy1GiXUwJDFE3qdAIwcOXPeEBm5j8
8r+Ke1ttWizM0AFSyYfTZEBdyjfTMo0DSL2gz2tuj6GmmXDoh0QXHyxnavCKRvUR
QYA0V82mvLZGu8yd6gsrFaZG+14KCwjc9yrHzv4NtwlL7ENr9HbpsESaVf/gAujt
z/GaOK1mwFXJU6Y5eWeaGRYgB0nTCVz0j8wq6bpQOqPutIX+qLOANwz4oea1fv5C
ApbsZ4P/y8zCTQ85Ns1kLe7pxRJ+5MWKfum0Pwg218s=
`protect END_PROTECTED
