`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tIWVfYxvUtIpOcJvcvJG9XjS9SZnW4gkAPzNjCetv8p9WoVEzv9mIDE+b+ZFM2j+
lari2/+r90m7yEU3yhbZJAgeT6km1OOlYesPxaveuDNyG9bu8KqnrI6mxT6HmeNg
Fh/HsYQYMQ82VBSGj7bWpJm5SvD+i/GpN64ZsoygW1uWEWgDMNUlOWrfMDBjdl/r
vNPf4WRSnHkHyJipH8LCld/3dL89WewmC7f496uPcIFRiov2nSo3JULycDONvFPF
TZMPq7EkgUrjL32IhsrN6sqIj2McvLbR8YUhdCWwd/iYRMiNYYJpW+57cIBNme05
zSD/ezy99I45dmVK9ER5axp4f9tnRvP1B6Ha50+WqX7Tpiz70ElOFbNJipKYDEPS
2hBgRlDA6aKmCMQhdhA73L2MLi2xYKHxie9sliWFq4/wKTKlsHC2EbyZPnfPn2bv
xOS+45BSkUrnB4DNR4JZHXoMeLqm0YOBH4rY/pqhh5Y/jQkxWVKdiqBNZcYh8HAo
nAH70PY4zY85sGdU8Z2zjGjkXF6lbHMx0Ep1DFnNLI4=
`protect END_PROTECTED
