`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kWVhIiUiK/wn+s6DIj6P68a1zgXjay+Gq2R8ijjgwHd/laMwK75+/3K9c3O9If1s
fWGihVa5/sCeNxNW8jnyNBBnaQkgJoY0B/CusrKBZom/qSusDL218c/GM+qpIsWF
YolsRC2+8nrK/TY/dRszdFxQTV1jl+nqL81ZnlhGSaskME/MiSlYRv+XvZdKGxaK
iy4D70Sml3G1qGIsR1Mz3mvkCrceLx1TMf5bSoB//p9SEKhmYSGxtIXMCIO/lTfy
gqWCBFvpc4kMppUMSKKp9N++2z1VzHyRcfclS4eOqNXApIUJ1pThQ2apATUsiPq6
NwtA0BqBt9IZI5MoNBaSkt9gfcxAXQOIXVoWgzuXqIoWVHzRMgNTYwRv1bezrfNV
L2SMw+B2GznFwueNqiGHKc5j9Dm6p+woguo4yfhOvXwiFHxl6Xo06u11vP/WbMlM
e7AP6AtUbHYafboK+YS3qs2vSV1RD1fg7G5fVKSlZp4IADqxqyp813IKfkQa6oWC
GuEk8r1owBMjTfCduhddiMnncTiOkwr3NVMAL9FSpV1uZPBvnK3OZnAgb6ToIEBw
NLqPo7Sja655T3qSEoQkAbBXHw/IvadrcBtiIEKmpIJNhEvgGoaaWdGAwKPnk0XR
HbMWFA3CtCkFX6YtuRPEvULjaoNriE7/S3TqpkH+P6jmLaRRe0G7AAyQVQPgM58a
mf7uXfwVHQFYRmBIZDuZIt2NdR8e2WmLYGruGHY7Jf3LumjQty5Kj9uBmtxDXL5w
sr1h97aryitjkp+im2oFGaqJ6EvDQgtl4BYtnKNSYip71B4lMuTjiGpPjO4ZlTbE
pAhvZ32xFOEdz3ZNZihLuumOkdCRQPs4NEl9lYWdtMSQZOtbDn8/LPEBto2sFik9
FHuzFVQqh4T3oPQ2mPA+NRjc5Ncs6D0O8dNmZikxBzPbTWPzM9c0qgQR9OZ1AL3C
h6YDw8wEimudHjS2yvREfIDQkl1GLmieWDBWPKMKdGtYA+UFQ/HtqD5SnqrjB+ur
x89XY3/m4swK6Coz6CqLX+3mWoJKWsm2gzizatC8bUVrAqW6daBeysvRMNYPW18D
0/2K/kHW0m737UXARE0bQ1Dkq7LJH3PLuAVrACcNM71kb4yXHmuYcUgvp54gVlv1
zJxWtMHmIFS9glROfQ/2D7eaAOuJ50Xd319A7vTThn7I6BK3VPutYC6F0NnAULzZ
t00bNvbfgQnhiVM9FHHfHzWRpTwzWMv7qJG9UQQKp2EVOmr6VN6pNGA+cSD0sEyL
Yo4mdjqI5cu2kSxwVhQ2a6yurFaTQvIskPu4j6V5mL0GVusFc9xUIXO0Oq6nCxcq
Qco/7aQUHi5F3QVABA81phKv2giqxs3II6a/1mrbt5lxZbIud9pCqdM5U0n5o0Bq
8/FgMEnOcV7mP6AvttnLh0LFtOnX1Dk1TsCLBs1TfcVLxnMsGjL0q6d4QPKVaqPU
`protect END_PROTECTED
