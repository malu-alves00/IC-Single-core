`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JtcTw5hvJFb0oy4Iag+pDGbzPIRTbK/lvltrlXlv7gebJRVkiq4twAwE2J5pjXUb
F84GMAMySZYoq1+Y3vbXT6W6z2CDD3RROYhdSdx8byF5eZPgRnK+SmXcM3fOI3zo
UhnQl2tMuGT6DQsthYpqH9SH/ttsYbZnZuOjVABScb4s60vHfm18IpzHILdK8QdJ
i2CekihNRAZ/xgfSYWf/+URI7ubf0d9ycUSinxB1Kj1KicmWZo49sa7/lfSszTPB
H3xVgpnsVefs+KcVy0vxzwn1jZVvlsxZkxQbqee0nIUSfh311r7UsfeXs7P66JoZ
HYeu6rv+UKkphdC7uXYVoasg33sP17BBSWvhbTzO8JPYXqTt62vNLaPZf9wartma
DH29Kh9TNC1RJhu1YOayZIG7N9mldKSv3u20cSl+x3z7LE2LyZ3JLq1CAZa6mYUr
X7GpU9TdVglnZkpQofmpa0wXsGSEX/SdktvNrfvvlZwrU7a39sToFSorLDz3c2c2
Fuo1DHE+oVarRG6Hr4KvAV2u1JQLa3mU0aeKyjZoFxIJA06jT0fhjqFzLNwHawjL
oe/tXpooHzzCUBeETKjqcprfIHtZiZrDQYSt5mF5qnJ+8PSUbELN254hxlfE7xWT
kgm7XKvgX+wsw2uo9M/LAROm05hvoqGzVutMKj6niSs+A/U5aThGn8ZEhx1QjZmW
86J2sb0zKrLgUyG213vX4I7Rw2l328zvjYdJvkYh1hcOHAnusZP2XAybyGjfvtrL
v9f4J4YdN7+Lid6LHcP83fcielis4Cqe+XyqSQ/WNvGtowPd/NRRMypnKFnw08e5
o7ELziPKzv7xVPytUMvO5g==
`protect END_PROTECTED
