`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VLM390mHIdQq+DK18YmtWu1wdKPiIHJ2sF0/uw5FD85k4BprXm724dv59XCNKNIM
tAjxfPGuLAF3/Ri0sfLkYhHMB3YnCutSa0jwsm4YCUOtV2HPOfFH9r9fUXWczcNE
EzSl4xBfGeJ5ErNUKyX5V7N7q5clQC9xze9PiJVud82gFPlbDSQRuXAfebYvLGcU
C2Ctik+14Ncf4bOzvL1KvqwvvvdWz+JVG+wxCZQcqm5mz3ekGUK4d6MFd4ekx5Wj
bt9DeiD3xrVvXJV+Akm5HcntRO8Gr/II0isR4KvC7A5hp5tG9MTYrld3ZtHc8kka
s/Ynv1Jw4i5oDc2RmnSeoF0dSaLJc3DAHV7BmcXU/ZKCjEQnvj1LPUutk0zHMNGC
ry3wiRy7TGHezL8SVEOF+FRGw9HjaBHbcrTPEgXTaD1z4v7QBd4bHE7D7mqK8U3i
X5NLEzlUq0SxgpwKdVN4EDT0ihv6LY0kuemjoPJ+UcZJ9F3VmI/o0Tt000gavYf9
CF+SmR2uiWUac1i97/9Q/3rW/0NLClmfhYdyKl2KldQ9aSZX+BFwKYP8CKXWZMXc
3Pd1V1ADaaL0GTWEHdan1XL0BIBn4prqIzqnqKBqz7gkJEXkqxMO4kivODBfQR8k
TFto7s/acKOuK9IEFytPbYYbO++/QreUxqx52j3l6Vb69ExCi2HOuSolJ2Nvr92I
kQDKIRw/T1Um1cgN1vMz8l+GNAoWYhcPwIpva2eTf9YhehJ0CjVukw+aIZKbSJHl
e14NHEIpQIEkS+yEVB9etir9pE2ZjEzffh7KmjYBUfYj1E9l/tVu4T++WW02qo03
h2l57f/ku+JgoHWPJgPGG8C6dl5L4R3LcH97BzHhf/WviWaQBJD1o4oHzmw4q+rb
+8nO1FBKgfzr0JQPvLaQGCo6cunnq55kX8R3DQYczFbLDPk9I8mba6rhflYrYB5s
o++itjcC2cDmjAcTKdStf2gMt3jw/5FNhuiAO8riTZUEsrj5cmpR0ZmaqzmpxJQz
LqZf8/kR9I/p/tTyqLVVR0wcdCbhiisitjVSPoBYttk+ZxU6Tddc2EoI4bp579Pi
8Li9fICTsnp+BiYeIlKpit876Z+8DQz4YxtFnGx7AMit/2DC75IPf/1WMgs2Xvyr
fK4yBXAoSQRnhRsx1qv8x2u6Pe+2Ue1M0wHkKHbsOGg+8C9aquLSlvjT+yVJayok
xWJweNlLhZty+nVafHhBh/IklRdO6dnd3a+X4inDyJCjzTf9kp2ivJYY/IS2ILzQ
UOB7mfF3pI31z4Dpz0tdudWqNTIMiCY2IeVMyWfMiTRekRijV//kLt79kwWHoAx3
Bj6fiHJH0eXo0lV2HCgHjngy6MLiJyg/tQQcqVLG9iz3jq/iK3E23EWCFd1kuNUJ
REVsO7T9S79wd+ds9Q8QmZxYKzrS1t0/6UqSMTFiw1AZVLgR5+AEGKPF/u9okiQs
`protect END_PROTECTED
