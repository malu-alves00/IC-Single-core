`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EuHatXSkG/zojzpktdYg4CzmFoYfmUShyh+DOdUZmqxM6UDH2aoxRZYEol32RySO
auWnCI8Mxkvpv15ziPOkcI1pJM6lXn0eRSF5Y4ZszdDI86DNLid05NqwFiaVyo3K
Y1Is3pXtVaRoOQkROFJMLMo0uzpRx0t14tjeiZK80G0h1M5sdlToa1yvFIcXddyR
fMnEnkd0NpEvt6y8iZvYwX53Dq+GCRY304QsMdNGU1cxYZtd2nl320Xd2tqsa1vb
e2tYuCjcKda5oHoEIRWlk9dniF9dXzwRJr+UlWWOhW3C8JaGlL9Q0lSNzBgyO4PJ
WuCBiMUaWVzwrT9Oey/nClBWEYuewHPjoaZZCJvgd11wxkK57FCxWyDHrLp6Iepx
yO+WpgpuIwslvUmyRYJhZ2hJYhte1FJcvRJ6YZNoDGOcrscAlk0I0TRPTX62VaTS
WgSXL8vt2IiiuZkkKslCVm+zXvzZFjnkxUkp8vt9YTNZK4XlNtKE+i6vWg46kY7V
CuBOFmNL+545I57K+dzQ3VVzN9kF54+e3oFVm+fGYIU1OL6cd8XID620m6t3YcUd
/4sDQDi+53LqVuB1fbmokEA47IA3vj8fgXNN7f5hj5Mykg+xWcL5onlClzSQckhQ
CduhGdH1Xb4emH3D85myASSbccxX8NGV9hQT67N7yr3cuqyQGCJA1xHhyEZbSEVZ
njutwuwfHRXNLjaYW5dOyv5PpeRHeDd+ehFPiKGzUd3h313o0ARuR4oUlf5d817G
VRJoQmzoTuWmdt2q7JFBwpiH5B2yqfyNiNu2Wo5XlH9qOzvpxRjXY9EFlg5E8ws+
dZLWdklzGtgZRbac6PwklnvMvO6tcyjGaWbnRARe3Oxw1Pxdjr+d1PPMnhW9pglH
oqDQ/ixD7ubfgEJRquJgU2MpV5NG47tf8lXjAtddkUpGW/9GjSYQOT34GMT2Hov/
lwzpZ4vYxp/EuiqHCv9mB4SDQRDaZ5MJL9+3Fwtv9N76l2qGaauhzq5TPwXsEKaH
Gyx1gkCpMfq/TnOfctjIcWqPGiE/WnyJMVEKzF/K+9DSEBBPSU4S22ehWelkuUaE
Mkj61IQE5d+Oe0NjM27gU0Fl96Gu2G519f2IJ609bf4raTUqela31UD3Am0m07fr
8RCZWOR8VVogdzHcSrcqonbHyC/7pGb/N992hjgjonCp1jLZdug8Sr4dDo92Ozig
4VFLCxSqKaQX+lXNr0z50xuZisXM16gXok605WYfUsajNkO884+yipioMyrcItvq
ygLbc58KpcCcW0hqGT3G2ea7rYEH1V5SAOQIus4+lHdpeGOwOWM64ppDvbpf9sw0
+L1XMrGKLyOUVTYRSpu044AI2L4haZAVSX1PEbcQhQnllIiqVUB/fmwymfW+3hNx
IA7fH1BjP/riMHEyz2JCJh3/73xEjOQpY95wz+UyVWMLI97LvRFdtDrE4yJc2WnR
Kve3GzbncJvWkfiyNn0kcKGqvqo4MwPu6hx6/l6QE3Q1FTBqH+vR1YXDBxeb7An0
AqRp7eZLUSCzsh2ZtpCalSZOqMCWokl9ToAWkZm7Da8SXeeA50uBF4qip1NDreBL
RLqcDpvxDa0MYSKJN/zoPjBJtTFCJ2X9bdEqVPXy54hs48tb6aKLtWWN4990Vv2Y
6C686x2b2mPF0kDnrbo3r7nHHkUqEASwVlvBERczQ4JVM33qQcNI1aer811q7iwJ
dlhBs+y7hPQVXefTrRpJxIsB2W8/cbAvxScsCgrWbe969dYMVBfOteYjI9oZpEP2
y4cjp1F+/u0azz/Bqm0CJnv0Akkqx9LR76FlLHP8EAKIUvUk5fp8flOy+4navMRE
W3OFeTIrD9J8pZvOLbmwU9GOs5ExqEFmOiUwZEYjR2Z+aEbnjPdbonCMYrQi/TGC
oSToSCoya1b8ju8nXyVMjw39GYNXwZfEwFDbDbMJcH85Z3L6a7hu9jDPEY2yIf35
tEgDIkbqeSWLIX+Y4mkhA64UFxVGvQT+F3/jkczjUeHtQQMWDb6YJ9lgsfc+o7CG
jUbZetdULn+hG2DjAj93u5a51bfxALoW4XeFFnyFZz36QkhCH1lpZSoL+bS0UFsc
MTriksK9zm0/IlCBwvbxuxsCg/zHYcFLlcmrbXy6b4bYbCWBNH8AGzWh6vHNl83X
Uq/bpclsrhkLBmTDKfbi6MTQSv34TOlGsn6sEUULA9z4ZWI2DJzUKaCIAsFK0+Hi
dW5NfOTJOmF8fzF7i3ZAQeJf7rQjTbPBhxPQ5iI1G4IkDTynPIjcV/miANOE94H6
RKcKWKzcurkVEBv3ABaC84Tq8c9DFIsgHAFftAVZIbmDJjvxZzp3MBq9pdp7Dhh7
hWMrnC1nw2p9miH4PTPQaLblqzoil6NoSMKsF7JV4evyYSMkCcV6Fq9oHO2coz/U
jExQ08Fv6TbLyz8yyqJDPwP6wSThN9cpg8YAaNYaghiGl/i32zRPIgXYhuxgHa0h
xkwc2jJoNkrKMyqr7e78FRghxER9LSawLcGZWHIjzT8OUNeCgTETW5eQ6RhtmCJY
JgaHJSS7TIbhAaF7kJvvD7cN4V6S9wD43Ck2RDZ3n3U5Ed3Jr+gTZfwjHAGp5XG+
oTX6BxlP4wC6LpupGJG9cN1JPppiPbsaygLeaXFPF5A9EA7Hb2CnJCiDV03FECPZ
oSZDcbJfitUZjteEQXxqwQyp7lWdIjJHKTE7PhKJzfFwhzqYVLkQWIh2uyW48cBg
rqjJGyq+uxraOg6c+O5+J1ala+M54Q0qY7Zx+Wyo8QG5E/9UR4QsmO+W1oZycwYV
2FQZiBKaq2ZgIDWhOKVWNQAP4Vm1uabd/MK7RllALSDXnWVjSQUtwCNPDl2eUcWa
VNo2CTt+kZIwCPiToS90NJee150fkGpdYJ3crbn4/8I3fUUrL5V7XXsm+Fb5th1U
njSuH28RHGyiWcesmhoOoe3vf/PC1jPsxDItvNP7yQe5L5DH/Mz7bZywjggpJRZJ
I0JcueQm7qwZBOcS/Id8hVmhNzh13QteX88oIY3+E/e/UvAJpxZBqm2XGR2j7FC4
DuJpreg37ExMLyES8A4IwsPUnDg7yHo+7KLq4LaSOW3Exnfl7xb5UqKjKh+i/0OE
m47jNDq7oyoIDCfvv7zsrajqM3JvMjVTvzRYM8VzC8WYtNq8u0z5pKLB5HLAlddB
HpBiHQO35krVFMBfObWRuNbgGkVjQGEfrsemDZevD0D+7FlStO02x63lvYkiPCuO
8faK8yJ+Lge3raxc/SPyY4p0g2Kd/4J2YQF8q+pARxHuULCeCDVwo2Aps/3QJVXA
mnfOQT1I5EMnD21NPwdKQTeZ9fH5d9f6JnvW92qeIdu/5eOgs9szqBaE9vdUwoou
9ZR0hKPt3rDP3BkTnWjHNoUAuQ7HU5AUxQfOYt5pJhhW+Icyrv+TjbMA9ewUm7ZT
iQ+ltlfHby0It6h6bgARAzm5rqbXv9mhrzvm5SsM+ryOFzZlr6nZUe0aldga4ZZ2
yZ6iVvae0FbTWute5fY4eHQ0bpWx2y5ZN4BzMTpxmoOH29QmObr93kz5tA3QY1rL
Qzyaq19/38boanPLUyhzWMOEC0X1me45lOuZ9LQg7AVEVos7ngMNJQKKvmhqipaV
ncSG6yhUOA6wxmBFlESJIqpuqguuIeZkaYYq1W6uvQTQGxZOyEdYNlo4JbVITP89
ukPMKIgyFnHH1YHlSZtn+l/TAIuaPPnTgclNKZk4U10jyDQE3HraWRADS0DBc+dt
zhwF1VjsVeNdGhHDZ0uBXD79WwauhmpzBNkz00sTgmelUvlPcR8VTGdR0bpZPe60
3J07qCev70GySl/PGmjtrqPKPjCIqYl3hRO/X7o48A8NprVY9yS3Va7f5eAgW7R/
0mQOhOLtlyXULKtjRjexh5cXxQBvATlIv+XeVGZ7KLGX5eqNDzN7LtRxnKvXcZUs
7z/+XGVjnw3epUQ9uJBxhvU6xPeWOmT3qO67SJKQPd1Np2a/eAI66YJuPxf48EL5
qPv1CQ4CK845A31TSPfmHdBlWoceWtsGIAnyo+2qZF+c+UeLLl+A1Uxsa+bZw8a6
Q3JbdZ0ZhfsPspiIVdUy/BzTFACGjCudP081k1h7dmOqcxELFB19a5OQO+EvIFas
IrSZO2MBa3sYfo9ZansJbx99KkX2ZVdPzjBmcQGqyJD5ETWkIst4G1FIY2TjmpTg
q/fl6PHKd8GepPEIwrKE2a/I+JN+vxPaT40vasGHxCCyAqJMmBwmPnVEhi3Xkk4s
oGJ9184SlVuOGypH9h6r/6ozKZkyzAh3Oa7xkOd1IzHeYBup7+2+mk/2NCJPVOsV
FB0qZAWlpDcP3mNrrTbFDJ8zNLoGExODn/B1cW/M42KcghkRCwSypMRIdqnyiE6N
DbxNBMy7P+QjodS5FcLKqkCXCI7X4v71pPO+bzFvCUrD8fdiYKvI+DXdnc92O+IW
AKaa/hn8RUVHYIjwOAPtONP7tLIlWrzCcgIKtoQxY9aWg++lurua9KU8xXqW7333
uehOgsTKVy0YaEjeVmYByed5dklwjzgBktT61GNkMogityygx2+HiuoAB4QLliRa
xS1UqDKeoOBvUf56/2/Q18aioDFDTZinM5EfUoS5EkwbqtUNObHTc5zgcqgpMC33
Cg/l17CuYAm8pmQktIcgshPNDAGBdJbmhOyrJUquSrYHAgoAowkdnalIDkuu0+ar
jzjrlpS7epmT3nEJcZb0kpncNTiKPPRgOaMC5z0G9sFfXB2+PF9IWJeQKFDOrdwR
Oy9ijgsojbhWJJN7k46Q9eY2Asku3jUKkrkQf6urOvRxnLxdGPM0SYM6AgAPJdFT
R8Ds04xa5vnAoSc70PC5ywLLFg9vWELeIDFJyO88QQLCuRq3TP6aONXUmsqgB2zI
I3ZQygflWwxtsqCYOLSVyEIgCFetcrspzoRlP3ySOf4nPrXcM/NR4kPSpkLR7nhB
89vB5hQzvMIt8rWgkVITJqJ74L8ugFg6uX3ItfVPh0KY6QWAwUlMkKtH65sxteJA
akq1hi3HLtfkgtLd2GEfZU05wid6bILqCpCp9ShLwIaIWSTIX9NIOGa1lzkG6VjK
UHK7lkcyepF17eFbWKIOcyNjplWPGEvIUBvjjmvcCeTxIRh6czAEdah4q5JHjZlb
MvizEhP63+y1fSf4lspXWLpxJUy78jWMGqfs9SsjPgDv8xJAHpbCrI8avDV3isjT
QjsmTBv/vo9HBMseV9xhJdR1brvym1bN9k+zbP7vS44v/BlKkU1ouhh2r7N2l9L/
aJJdf03ItcAbbIxlHN2cKcQ9sEJy5NsCRlRtUwAOPYWcVXcDepUUJe1pZapnuXDi
/2hF0z2dkHodGzUEOhP5JpGvtumzs4uWoEYrh9hd6Ws9OWtNjXnTsMq7cG8F4b+R
EgIqEY3PNph543VHLxh+S1Ra+XWTr7yeboJBiJlhs3QIAHBKsoFc5Hq5jFg//hun
b1oMIVsbzhVl2y/eX2+qLBMvs0i8PWwvPfHXscM72vWvLK+HhDbmP+pFAi78nFFQ
QIavtswhO0rUIrja4Va/Ldb8yQg5o3urnPPpIdcT85S5OmKHZJwf6elPW8BQJZ7z
qp3CjxnPuzlAQtE2ctEPtreNAP1kiihPlSHI7eBLe6Nf10iXlYWl8lBvqmtSJIKE
J5KRrMGhvpJn0cnbvkr+eJ5DdH1Q0V6xSyZHo1yEyblzs5FyKoWTv0/xrh/XISjF
N1KXbhdwLbpOzJvQpBT4dqnaa9UC+NShxDf2Nb0wMcq8VTNg0wJw/4NW6G6QCNgz
A+N+bd6Wg8gVy0WqDQ9LH8p40n+y21T48sfyUPrp9R7X86y5hE0061wbtqdsNfbi
7cRlzVSGqluMJm408MyB/q3SMcBSHBYwDVh7EkqTjCB9mjwMI3eZiT3zxjx98rKy
eECUZGpgunH3VohkGaqf0ueBMbkat75z529iGud3YlZjyjsdPiNn9TfG2kfZK4+6
1kuKERTKy0tbp72ZD2iHP00aqbw02BpesvDMsnB2mQDvM55ByZkVmGC5S8t7mArp
j6TLaDQ3z8M3v9FfGHVlhFcGwGiM++MDSuxkrWr+oJLW8iOnrg8lh6KAVbQRO+CP
mfpN7GxPWUranIuh7eSg9v313/L2E4NVWbbi6kTmVx6+kGOhplvguZhpSR8ryZzd
ryZ1iBl2HsJG3nzctCzsTd/FvLmNl6I+uHMnF1ABX+6bRvS7bZhNBp+2ACnQjjo7
3dFKiRt9QAMx/nbbjKYQ20Pvs3IrMi5XK6RVZIFZ5bg8P7UWe+SNxlyLoOecgCtW
swAN0uj5KVnrJ+K3c1yzrB2sWzCJGevy8n0iiO1GJWzECzwrMagWfMOpBN+GhwZu
oQeBgMlm/iD9dUL7JxXlV373PdyKdpe4CQNBat+Uts6MTG7fi2PGtnDNSFUgC8k9
R6WBPC4qvimw5pWSj060436xqfb9DJKt1/xyHC9lF8gYtebjy6iIu/AlnbB+JqE7
ynbxl2xhdpgR0+C2ZK4oPMvW87RPq6syLuUtDsJ8ajHt9sKjTQH1o70ZG0G0qC7L
78d0tHSzFfYO3BO+TmjlSBwn/knZ2IbdFwHKp/NBAzgJOj7Znhlzs9TdHi/nRcVT
GGbJTb0a1xY++enBfbviiA8PkgRNmZ5QNTFN5vsBVkMvc0DkrSO4HmQbs48YPdZC
y4UVkNWbUm88VIdZNgsGUVsdfkw5bSdaiymMv7gpBa/Xno2B27iGDtNQWLtdCrf5
5/F4kZDp7MZyeyny6kVM6hCGMR3kzl41xhdc/i/Mtjugs3xgmdwQR+zF21xze5YR
MZEaNeruQHHWPHfq2siB9eiEmqY15WQ5B0zO0WaGnIqR6wMmdGCwyHz3WxLGUe+w
gllGg4p9zbhUMcpMIUCmNt6Eu6QPfHBwOsVtg2pnWvUjyPkmS+jBE+ctDc+YB3WC
lSN6E4VJ5l7lsAPFuUat3Qll8Y6yPPcwZejlNlIZWMgBwTKcfiQtWcPVLCL7ILmE
VNyzYPxuJOseCvdM54qSJbxN7wBklGbgYRKCI+AYDGRGGOIrywJRf1VZXKYyvSKJ
0zwi+s5ZFtjGljUj1uutF383njryDvA5pJpdxc1SJgK8Y54cVoizEVeRaZdQtXY8
8euBfK3E6cZ6BTBD8bvaII/MNLOl2Rbbep4rMe38f0weE/agDMDF7ldAI6l/gp5B
eJ59iYG9BKqvx8q6KN4XEXgvI84lv82w69gO9okoh8ASoxUQJiGlPJWa8LXgJeqt
oZZ1Dq5w1wJoAHETGxPJXZpxQ4t6BQR6VfqcO6eBuoliWCVGK/OHy05O2mZmvUui
Y1EKGuEWiFFpkVbD9Ak+aM11AAjguxaUCwWy+htWs/XU0s8yoHQ2qgcUUksPw+CL
ZIxb4wKOnELShFbY/eXbQMO2BpIMsBr/t0FsuQ7JTOsGEOlcKTJz4mBYsfC3M9if
0bBHGcIO1EdfaIaTMav/yMvIYvaE3Tiu6LL4x+sCWFBfVnnodXPDhsVWlqWU9+dW
aN/87tEypyEnquqgpCO6C2wqag5DXfGRAXAMukXQVNxN9emPDd0ymhMmrshKd73p
1r4LPIU5hGidAONqhhpjOMfxk4U1nsIQR/lz+vSTn9WExKATNShQ1d1lGnfPeD5b
Ld8xeCzI13z/rZ6U4uCqnHd18pn3+3x45aqXaQ3dU1u7PE3EclPS0i5THpGd6Ytb
BsLABYybXLsaEJoLwMCTVvNW2r2KEuPElZKAa4kfJjfT+hlqgTQfslBBPojMzUjd
cGKh9xVj1k6lLjXQmRBZ3k831TeZGNPvRKzXjgSV2swRuUJHGAvUliS4e+rSnvMa
/lJRE80Niqy1MGVA0DAcXd8AvAAaqyWszUW4AR+nZfJW+11QaOUBk1jHxcHc52K1
ou9ISeUsHNX/uwGnKR5Nzv/X5leEtU/cG7/mqaz0iF8zabItCGS+HAmUQKe06O81
1G4kgOeSi+aC6IttBUkSx4y4RiiV1KyaXvsObB3UvIMGKy8rlq3Bqkv2bTBZTd/a
8+fRm6QlEsHwneMvbZItU1kOf8Be6euzNHWyNpNNs9igTsRBrfs4B8sgyENScTEn
49RWInmAD0edHIgS47IzDumziV2fSMYuilq7K43qso23Z1mXXHmJ1NhNTD35n46S
iTatNpcvfwN8o1LFeof1t+9qNAjBrgV49QU/tVhbz62S4MTZc4MLVI/ZWOajC0cg
mz+fwGdMrn8sVMOWdgmJwrnsy//KV+M2zF+0wOQ4TaTgZ5VrCcC1F4MXW+/8oRPC
CTM3oc0FZaf9MK/5uGOp4WKbTrTQgYScLGHz8qz/ojyPJYcz0L7VnEjHVkk5iXny
ywpnCJBaVdNa8pnz0P0V8KsWm2qo7q3Rxe5+o+yW2x/hODM9QaBtAZayTTErWuKV
1nxiz6LftO4b9Hzkx9sFPgL2mRnUPbthUAWDEysbMJ3sq1rF/WClKvdcsUH8hqFv
1mZHEClyUS7iCSmptD+HLh4X2epJpyDuGGlZRTIDngrjoiQwJKv5bVSwJpY1Uuin
TA1aQC8spur/n2EluegVPwzxgvbw3kgruqi1EJsJI+DjTXdcn8RUFwFc2ayDa5Ln
p/TEAWuENCRttAaxbmRwe6Y5gO2j8eG8qBrg1OU/Vxstj0eguLWBzSk2O87XMKFQ
X5Zf0s09W7lnXXdMguufQMvu5LK/nBYsxsUbdYuwg4WPgFO8E0CHi/W/OdwOCabf
G1O4T2zJ35WNpufJTkSHhFBYx772AvxMmVKWOUlRy4yFh1ojwIRdtOP1o97ORLkv
ZozXFE/S4rvwSRfS5N3pDkMQbn9r+UAZPr2RZ3cUtJqwFFIj7V7aYKVOFpOZlGYr
Jzq7QAZ6/opukVGNJfjt/WZGaAiA6++njPN6NyBcUI3Do38TbeAWnvL9wi4g2Gnz
AWSHpSOmAtU0EGhe38XMxVGE13f3N337NoTpqQM543/MdmJ5KMVI0wHRyEYfDG3G
izsdp3q4hUSJEiZky8CIlJwkN0l1ocL9Upci2TWPLGak6rkcVF2VyyquHdgzevAI
LFugmlYoQP8JCPcOlekNxEMi3en1N1/Cf1UhT0yUKCG4E4eM2OmfAl8nt55vgzhy
fKw7PdY0BYR2fkXDkJQ9+oKhK/PgSUDcAD4DzJOFgVNr4x7xS6reVO229a7D2JC5
KK0QrJ3yc3YKceEYxZAY/CMjwCG4DglQGunWLB45LsWIROdRRh0wmB+U4flZRv0A
x4qdobKWpLXj6eLLeh3/HMx5Q8eTcneqw4YpcapgZUQqpu91kbF3+QMfCEyuoPJU
HsyWNiLcwlLyE4h6+VKRIidJP9ofdpH0+4dF9+rzdEDrjhuEEk1c6A8BtEquU8IC
YkGSxtQhJti8iBMmWaZ47UeEwnJgVE5cDMN1+PZRLR926vNFroX87XJS0m6tho7Q
6srGStmXm/a8po1pIOsdIZ9fdwmgkEsppNxX0wQupmUabGDaFh/C1HT6NIXRykTZ
XkmafqyCSwjTVzK7bY0x096A0xp2H3P9yzIbzkD83G5uLAijrzGjJ8CfJCwF/ek8
+W9tXK76uEpudVhBvJfsHR4wes5ELNwRCGSaudNpLx8LkQKUHncckLOyAxMthKon
ys5SKtmN+2ZMUpz88Z+ce3s2LmzmKailbIZCVv+LC31Gy8dFnOPWNPCLMocBEFq3
r+PNnFkcKJHALWthuIwVBmCI6b7PsPdHWZCvQvygOhqVMUvxqawtCvoWSHxZsK3s
+F5pfi4OyiKAEsJ/aS6TVYXL/94e7az+PCjfsjfQlhe85/F9+5LhT4ywNTUED/DT
o0mcabtv3VrBqvu4gexTRsng+ubWaG0rWBdAIwBG6mt6/RtQW1/OPpX2GbAwrB9P
IHGSTKU60YowrjdLOrBX8eo9s5B5ELKP+i/cgg00+7P6ZyQCUwCZxTbkCWSbxcfK
X9pMwKaI3NTzhZX+6C/JBFvqRxuRkOhTyeyK1YEvXS5hKPPR2SSq2N4bjq8uQHlT
/u3MkPRgS3vG4gchYrzARi+OX1pDBYddH0w9Y5RN9EdcmuthsKp65rRcYJzPIpA2
ldhe+LJDgjpTae81ewhgL+YmPBndpIOQQ2TbyL7HDaW7IF1JFPVBzH484W8o0wz+
lOVXblE3TEW8ESp0tJhkzX0Ng5UvyP8Vp7FGi/UbIrbXnT30Ze15siHjyzAwN9FQ
B0ivZAXkQUaOuYCRWUYrf95kx6LNK5iVuXTWD1ht8+t5PkQxLUhx4kNrR5gnFL89
uPVBwArf0RFYx2ZZN/R0HlnJU0WzrsZAD92WYpq21jiGSQhJJ08sJWwx1q5tqCOE
gFs5q8Z3WxDadItCUEIPcDZdJ21FEcCntQLMuyJjeoK22TU+jJ5wSvUW5+WQk2py
7EzqzcKJk/37B0SU6mfwnK53GS8r9A95int9C3nGR/ELSDq3H/uQDXzxsgCaQ1ys
wYEzzuG88eNbGt0HNXoxYEuG4pdWG3Db1PdWINRhi/H7jBEPNystTLkZTEcGH8Eb
H0axeGHTfFHAKCUCtvXKNsb0oBwS+m56DMWbZdmFRLG37cvI5idcCGvrUihweajq
/+7qpYpsNKz8kWhbGZufI7A7mPl6owN9fxvylq9zmYQQ9XLnUBDzAm8FaQHAZQiX
/yljINVvXJasvcVwTxNq4yDgpMxmagT0THkxazAvas7uf0D8qOUg7nAXeLmlkMlK
Sghi3uXnl1IasEbcRE4opmQV9lZpXt7/0/HFIPviHSzDZmunYGy8toyb4FWpAIb2
+v3p9l5to5wimJnl6DV+OFJJIGrpFDaGcJy6XNozqVyl1WI6yRt/4eUNqDAvE10Y
Bu6DMAxnG3wFWzwx95BJl9YwbpFw1Tc3OjKXg+PqvfnxfmvyC0ewjvhPE4kQvpJO
aX0NFS5Bu9aoxQ/GRTriZMQ64g4GqB3Un3CR/nV78hpUL0MLI1QsXNgCFDW/w7vJ
oU84VpZfksgrIW1WD33SGI7kkZBOihuWeKCKc2eycBqxhB63qupkQHEWh5KOBQzI
5YmZMF/ZPV3ISTseRy5yCILUc2nOHi3sZDLYXZIvjorc2fgJ5xX3qRSH/8QHRhLl
1KZhR8+QR/vCflg01Ho52ESH5gjJlqbwLEelt6hbUDKykWLEib+oeUzCyNsTZJGK
tbU/UbUeLf3S4Zp9XxB3ZbtbmoI8TNLQmTsJG4JTDhJIFJvpHA0cOm8OrdXWQG8H
NN2CuMg8px5LRuTEgOqLv9ykN5fBCGnmmPn6Lc1PlH97FQackxygEwg8xZEBfEB3
vbmiw/OZNkiiEi9/qbUVuv/HnmOBbAVE1flDgwayp7wl6CP4ePphemRReQpExu2h
ZebHiVEUA5+lu9oAyohzWDMCWvkE8gEDQqylR48YKwFA7mkUNHBTrR2mCvClU+ub
X++Hu4kA9ONs9rge2j2BoFVpU3Yk1KR5qVWu54RNip+a7BtLtYqVwcDvJyIn/96j
hEZmqHllBAe5GPM4kiqm8/NQAZZurgQTqvoIidlA3Ev2IskSyt1lUhQ7dwrNZxsG
ktiYRQHCpOMPF2IwEGywNMs42YzYjIuxPVpeilDKauJkLldFM9whmETVMSFLKB+0
AMlHSMrQmpxNYA/bqab6fhinMB2nT7CxK4ePZJyy70dyEsVEXo68PsenosL5FBEs
9xq2LcNT4G5h0D9Ao79Xy7Qt9uyzIonXWY9Uihq4S5O68Md6XZH9lMnd4nG0cofK
72brrgYazujwvmcx0VYFOMK8C+/2dmlX5VLm3Wo0L6FWJR9B1eaniRVxY+RELMbd
qOD6VcP5kDRR4JFRyBiznMhzaCrb1CR17/5KkCX8KOx/e6G/sEIzv+xkJ+QucFi9
77b8ryljqVU5CjMgPLFm8dsC3dDUr1IVehla34/ma8YMzQEubgL8buAFcxvXZwSM
XU3ctduGlktSVD4SBN7THDoh+0gfE8p0dwEzZxUG9Bidqgk2LUmTrv3UocpP0fuU
7pj1VKoZSxunkr8v3I7mjv5hl6wq8whiAv7G4iUuST6NnFWhzkYDal9cG+aO6ULN
HFsfSf7/5JmbHX4n8KYn8l9h1/VOZHLX/mRfNyvkHQfE1aoA9f+RK06Ylzsh+w93
+QvWDWwR7S7mhpNH5YbC9jm+yTuOjGnlLskHHXHL9vuzfC5Tq+fnhSEZ7Q3EcIj2
3xgviOfKqp/9l5kLv7anT3OyFL15A17efkvrMjtQ0dY9kPePjstDFxCBYMgWrgtT
T4gMpy488SXF5bqDbJBBj4sov1uemT6rvYSEfvHfL6kAYefgRMXn+jrPVwCfJUGF
rXFVEXyq9yblLBnFEoZLTUPTqJ9N4jaYVCIcfQ0PrIwp0OOmLBHJa8NhBxsvj4+J
1m3YmIN1QQ8GKLky4cXpfZPl9Dpa79aFaHB0q6OrmRAnHqMNQElXozKcSWhdXjab
fNMFAmrVXcY9AlKeu848g7JlMDA4VR+pirMuZorLr1RhlzSDl+YbI2wUCLKKvUem
PYmw4lNje5Fckg8RZHQq34Tm6PZlE/7NTYbjHYykrA4roDA36D0MBJ7IHRXw4d0t
Nkz/jzxd0nKtcIYusQRMfGwqNUPFMQHmK1nxhWGqijOnGrNRpshiRLtSxTnrg7AT
QJ1gVw6l9hFOBMZFqqiBQXGsLu+VpqWH7ilNqPcqUJGTnOMTICbr4BrbSNdXRB0T
mJIYR7FMz0wNKs+ZUHKgzGJ3qu/l0HBzbJeMuXi0qM1BowDb+Dg3MjbhNiJw9uQE
KaHYFp2NLBT75ogjvxDu3iWon9UH9XVq6q2XeV0LrjQoC8FirPCV6zhRJK+vlT4x
NFsUgyHsHdnA+I0EhcCQPAGujjClGv9HqbmHt5RSgniulkc9sraAIRwCZFxtXDCm
K1+0cesgGnYq/nXLGPVEBzhuZwooLQjrOpGMhC9Gy6qLgCuv9BF8/rK1SxW6K4KS
Lsmz9iFxRpkhYmeMXK7+q79UfvlgysSd6/kGLlb3Rsho36xwtktB9cBvYAm0oMlK
FsYRB8U5lH/tnUTo5JZt5X2hwaCXiGPwhw76N8QH5IGIy7ZM5NBXbwu17Fe9zT0L
dgbNpBBgi6up5S9pqcZ9AuEgo09cTBnmZTHMud+s4rkRqEM9yt/oLKfd+u/o2949
VzN3qBt3hr8ci7EDoc8xam7TZC3cQ8inOTZfiaol28MSTZHwkEL0OIVpJUuEVU8p
TIvbTZtxkuaE+5KFAvKNsNIiKd4IyTlg13hqZHohnkwV1tR6wjWernubDeDudj+k
KTfItbMF1rqnlIqJQny5mM7cGv3IuJdM0+EpCVf8sK5GCB4928IZb29pbBv0Sqo3
4WBfcGVqY7Owv866zrqdBCrm4WxCMl1GibEgeV84KThUZkWSarxFKbr6/7jQFB52
5okHL9TrAKCR7GvR6L2zu5PpLNMVaW4vBid4eLn1fOHlHH8MkO93CcESZkUhhQmK
wKOl9chSYMlcuBXUqMef0FhB/f0cnlzCWpS13pLd8A6gjzBVcsWuypbL5V1uLnn+
iyedKOfCXRiaLxbb2jPwUcGHfynu/RTwesGowlB822aLouer82GmOcSEe7pYVGPu
voIoP44t9Rk6U0kot41+wt7hI8SY+OxgxW1ChHXgn8otsZG3vmHGtgIUr3Rpf3V9
Cjkp8IrDmu+Vacq2f5jVSCyaBtskcMTitaVJ2w2dtRdgc/vfqARnirlUtJpXUJX3
X+bNHWF7kE8X76rKxgPo0hWRAAVLQ3xAMqOubNU/CuCfhB6jJW0vW/WmKlX00c9h
xleDPTTUhXjwZIL/wiDz+tdVv9fbWhx2stQQNgGgb+UuHyfHF9qJcyX8rAP8MU1X
E0GY7fWZqTzcn9mnVnsFpE667l63jOFpPLNpfP+OCbImboZs6kAReYdNPZcMXDLk
wBKWJq1dzPf81UB41oubnbWL1GzMFb6cz/21VQEnxXe0IYTD0QLxEBDwlUc/ZyjI
22GcS1lTq3N9gGa9qCe4oOcwWQEEZ5NUkg5N7qP9N7AnAjb3tcIlYeKtzsCP3skS
UQAfwI1dYXiNvhEYi54rAnbTk/9yocTIT70UTz6QcJqbx1HadkgC0U4tMq3NksnE
6nSw06jknY76H9g6lDaXosjqtLnf5fS9zmBvDGX6bg4two1sGuR8C6ZLyYMcYpOX
BUHtbysEf1AweYegkAVSpXlMRgFecvTfUMBXgURGDxER4rwuOfARrNVWV3MATWz/
w87CzqT5MUeDi1GTD6xqzjkAwQA6v4uIVLHAS9KS9x8RDj8NziLSUwpCo2xDZbFV
5L4hSTYVrYFQ7A8nCH7nLgCgeR2aW9yD5H4RlbdLTaKlpHm2kNpP187HgcuGvRID
WrOxtpomQ7PqtOfT/R0k2Quu4hqz3eNVgdNWBQwtgPwY90zBDwRJbcFs1UGIsD6o
3IInbQQtnJfh1W3uJOCqeWOreNBDyK4xMguzm716DU2ubQvZgwcgltG9zicvYgwM
ns0Z2DoPoxay7HuUyDAVCb8/8rPPVUBgT704EZxRGMesKLDjcpgew6hap+HJmdlJ
wQGl7qZXGHi3UQrUiJt4TLAbhrJBqXs3oXzakR+gnmnBN0Z8+7G+zai2eO56L772
SNEsBwrxbkkA99J1JfqUpkkWd59ezmk0YIQRfYY1BbVLd02YBHBM9TdWn98uzARd
vRiW/Kt2SsRe9xdM1ZoFH/esgF8g5bcT2sft9wJgrpLa32MZxp80xd2N3uldLvmV
P0eZI/s1uw5YVPPF+ckxxllxMP2ZjUT5VcbnE+DlR+gcpOec7h6IwspeFAsfRhmt
SRkrxQrh0bqikDtH57zDeSEn+RRPdcTsTwtS2fo90drmVjqrov6OfKc93rjq9XMJ
TOYXjvv+vtSSM1xj3x1VS3wo2TJu7EoQyPDgfVrLCQVDjaJRRcPV1SmXldESMtut
NhpzJd65zzkge03johF7ICaeuKER4dqGTBNLg+4xVpBdeQ1TRHa4y3TqQVGSZhgf
qponezT9T6B9FD+LFJ6LwXyOQZ9zX4wIFrF0svTsJJIfdbSPqHREMJCsesNMV3jo
g+lkbCqm4fxjsv7ubfsKzLk1N9/AibKtxDhXBrg8lTtxkFhCbj0ddRrHBdRqZgMc
pEyBvutaYlGXev1XqeA4V/GmODfiQERTzMlVc0Nm5urZ5HTqJJBwrdxZmQhJ9p0w
s4qav9X5DlRXsV/4Tyz8CUCxpIsChEJ2sOOuBtyTS5GCMJ+Oef9xKmXe+SXFrdZz
Av5jbPG42p848McKMF0jg5te7zNXZFlHva1Viivcfhy9KIvnK6lJ8e2CS4Z4HUi5
q1WA+rx7YG/fkEbG8jPrwzLzCqdpivwS1ONEKQddlRmivYbUh8o1R65pc8SjQ994
cmz5VffApC2sFW4Pe36LvQ==
`protect END_PROTECTED
