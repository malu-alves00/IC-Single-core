`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ncLJn+iruZfz1qJITYpgRr1Gy9xE2g344R+JQzQ4JgvrOI38CO1YavSOzlKywzxL
eknR90NQhWYZMtbK8h3tNeEEEkNKzCjEpNfXnH4DFM1I3YjgqlSlBtPO1z7YcZEA
BkA5DHSvkmMDjj3CzbD3Tggm4JhzGTGElQXDn8dwy1VBjs90QCeKpeChNdWuh18o
1J1/WE7ca8yJvc8fXhWBSRB1nUrrs7jgrjTCX57eonEJS1FQDc+xwxsD2suatERu
tn8IKWEzJMvxQU+kLQe7fO3fF5qHWx4p4IfcilFxSB9aXNd3ZSZwl9l7hay9WMIT
XFUbwdAlEL+9GUoUFO/VyFekfO96OWsdJbZN3PjSCH4NXO0x4qRIP0pKdTFUEl9c
E3UQH+SNT2lY9Vmp9YEzisQZGJTksrju9EwzvQg6+3WkoGxWOB75JhqTj4yuJ9XP
SgZZGNSsQzlCuFaAdC8c9yZlQ4YpjLiYZpffEx3N7VvVtfMtgoYlq/tW2EIcGKRU
pqiuvhfRc0SN/WRkuHuKT/uUTnOxRNHfR2pMgso6VFJrvGx0Msj36WJwyIE8Budd
e1lr8HZlgRz0TAXWGbdMlEhr2Zg5oQ5BK//WekpEPJtq5Kfgls+pQkp0CIZFBF3b
XHPMJsWor5lpr9bx8CsOj8M1gegyoFHdOvk78ncs0O4osvHuuxc8xbnB/3S11ZVQ
AjQdwTXaM08wH5WU4SX9dxJH69mrQdyO6xVtJC1mvFv9wgwWK6n/YjIGRyOBQNBX
qyx4odlPmFucLPu88GMJEC19uf8O+GtNLXWkUH9GjFH0ePKq4l4grtwdU6bcIeIE
vJOOXlFcSL0w2HOWGph/3zKneLlaXakaQO5yw4fHyyQVN6kMYBfA42TtDcZV604g
qb9turelvTfe+t9TcokhWzc4g/EwDqACp6J/HyUZW8JwwDnCIMcNEf4ETls5/iEb
nIcx8ErhKANid0aO+E5zSjVkNZrfDQAhUS1cyIwWybbEIUkxShQ8eFgMG//KERU4
Ueu5UrWNr1J55Wr7xHlM5wbFDMfSVDilT5UQMpOS2RN+Fpwb6enWWubjUrXBGg8G
Z0bv8NNGnykBPknnm2XEbfYMPJPa6+FIsA/5Q5wwIhv3s6M5BmJynjdZw3DYziIj
6RVTrGmMqMM2pSpyYFjxb61mtlvDc2OYCqkstj5b1m9UfkN/jguXzEvZUETyiA3C
9elsz2p4QKszcj72gU+IvXheiIrj7GluN3KKdD01JFwSRuSLuBug60KL+8bBR5bB
64dJRIfRGfjtRxiARBVrT7XVbv6D/vZ6p6eoQIi7wmEx80zHudN7qwY/7sdOM2x3
767FYgefNb021tJeClQDgqRF7slX4Y2gGpQlE5B6LgVIQQEkBonvjzw8QxI6XoXx
J49KW31vPH72HFmT85KoAlpcIup3qxph966erAUBPUbpxsxwk+xGyea/VrpJDAJM
ZBFriukog517e7fhUKNbzMXp6og5KHQk+H9m6IUC+gk1RkAKpaEhp7OVVn6/RohY
OqPDULk3Oh14u0UllFu/cIyuuH1fLpgsaana/TYQ5c+juwsg5K/nwpVSFSJTmZok
ikX0dnBhjIbcVy6e85d/nNrhBDydHcZ4PVGify1A66D4RW2JZ2Y5UWvJeFcsrxwU
iB0qZ06MbjFLRU5oVtdVT9SbvvPyyxh8qCYgEI4pkvXmCdLfO+30p+04nvvjMZqe
f920xGMZRAB0rSJUwwLzLBuvk7mqd3EkbaNDhpZmVvEdQzKC/skv8LQCqMOc3IjC
bNSBt6UE5VX4LDlaD1YUU9018M4RJo7P7zr2cVi3NRrVcE0HvZn2tURdqnfHx5GN
HS4RLcBvZ3m8OLXkaE4xMnb2gaDTdptIsXnpnQjMQ12/J7JspCYVVI96WnCwTPGB
6t32KCzPlWIlU1edU0pZLBeNqWYHPdFs1lthljpfdfX+7yAZQlC9zmBulrZXHGec
Y/UnbkjTZzfn6iWXFGSEzRSZD8Z2we2i6iCmayXn2lQucKFPtgLJXYSi8IW+ksp2
iMfS192yhnfOQHg5ykbG7g5frUUhl66obimFlPYaiMvzqoGg5ufqf8BmbbddXvyo
C7v0lh9LttsEFGxWn0gBjWiTc4lH1agADR1AeKMjbgHPhE30GE4N/MXUmsfiVU7n
+lP8C+XvEM1GSGclnl6Br0FiBwe3QGjqj61kpIwx1pCHR6OmWf6s+pB/5L4Szqsw
3gIaX9zkkzlxcDylZBdQ09KY/nwwfl0ohfzq8+13tIAHeFvDT4B6Iot2o2w+RIZx
sPu8Gm/gI1drSlNrqfLYOH/vzEnC6AFiQ4Fszu7kQsIfx2IrZTTKNAfLIVHo4DIA
+rjc+3dxpaywck9pdcjv0oI0905e8dTF0CMmNgfrDLUobkFSCKKXhEcabboKPFuT
Bajyud/jxHD2RsqmfBfnf1bKKJQKnnfmrJwIKL0BYgzfHw9rFMs02BjKz19bRm3x
FhA0Y1PgqhG6jxHr9vMFTtThGgNo9F7JxWRfZgrVAME=
`protect END_PROTECTED
