`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hSqSlByhz31zQewyagKfOrfNzHEAv6mPt6sxPLb5ZGbfBlkRF+Wgdy3Eh4feACLJ
/k8ryGMjNKGcT1n7Aq0lBrxGWz4TNOOYG8BgQwiF+RBX+p4IS2usOXi6oWbhkuJj
kp1TtUvvV6IH9Rhq4hiWHuzAF1+rWaCjXlKq7Up9ziL9n4OMKMHtCh6KM2OkQ5eK
iiLGdg10G5e3f4TqXb+X9BBdxb/+whLoWgPhdpQBXbv2D4ueIUpiBTdnkAjR6vvt
XJVN6DeAyfHYLfbqbtbZmnE6qpVUKiMX+dfeTWqhvemgllqrwzKDcJg02p2X3f7V
JyXIoQ9uUh1Ckmf5amJfuo1e3fqrGlMo8/AAHJBvvZ03/hEhNbcy0Smre5phEeH8
r2UeaCYHfvgAY6v7FJXEP1KtGsSKq2IVAdRIRVVClmHwILLt1HRZFX0w2Ym/+LMu
K0i7pOva7sdKkgtF+icTSi7gY6rgeXDUQlP1Coyr7JAoZV0cQZz5+3PiUQ6fygHV
q8CwpRJejpnyN05kCm/y2IA+fHnBjqPaN3+YIGQqJ5ja7ReSJRRJ+UhX3qQKVij1
/zJwiTCjLFjSazYJv4gPGOM9p0O+kL17JtEcMEWaZFK9W/0zAInyooAZ+WzIiPNG
zSjOI/RPAz7QTD7EUpP/6IwZEk8LkQwRfiuU+7dApAYLa6mXVmWeWlRdY3acJVcS
h2aglPCRyT7kO0zJCxr433dB/yxsJ96GkQMIe/yeasudMBgqEcr4qd//ZWTzN1Xy
oFcdlcwuIG+8eIeN1xE0gxsKC9xfhn+5TR0+wYRB4C2Z3h0nSlTwKYFVqZYDmhhc
S9dPhRH2qhEQoYzEGcgiLyps6ve3UeTISj8yGrIqMR5y7o3+ksyj3XC1Ta2py+hq
RCuAVgZFztqrcofgFCDkM94yEU1rnHHdv1GknqX6LRFzQPxusWj+gRLp0WPQwzIt
j05JHwGdnhGm/27sUacO0+4SkTLjHdf08mOAMH+FgEqWCpPWYKVB1/xIHOshpxxM
sAe3NQDsB/iodOsa4LBl4SISDJwcMCbmlra5G2NwIxcWsCRTFDwEMGxuYjY3kWyZ
xnfCEJoUmwVcIvLGpus6sZXLfyS5d2/D3w+LbqtibqbVHo83ZvaFzkV5dzT5dGdO
6zeK6ehMtcIV1gTiZQx1vAKEqrUqhLQzEuftTpINFMx2JIlDgvBsBTSi9a5lQjgS
8MJ322/EKd0r4LgbjlaqhOXuybtOvEqiwLG7XlRTYmD0oE9Nhc8DMwQ6Mo7Z3M1U
Q25JTqufO3Djy7SIWOM1aSBqB1QuiAhVz7oxxE3hBE9Th133QsIUlrmHuWpZ+Dtn
kDNk8vjP3K8ZPr9REI676OwnRepQDsWh2RWJvv6YECVBPIqej1v/2RLUiTKoGEok
EG1tQsinQeBTdCaIP5js5vDoiptbj5rI8g/P7jDS+RQvxeHdyUEU2hkJPkElYzQg
T9EOGsVjXwHrm9ojMg8RbUHANmndWh1zNvFMyZMzrtDy4RrI5/2Gxcg4LgeAGUki
FSUN3aXpQtBxQU+p0f8SxUUz8NZze6hUR03FA3EFq2Fo18Ua0FJc3e2o/1qG19XM
H5l7HyRW04RYBmsm2+jdGMXids4+mBppz/PJ1IDQ+Kb3t5FUIAPMebU5LmxzkFvs
cU7o33onXUPY7isjuGz93+kqdiuqm5RUp4RefOfjgEOrtv9+eJtWKCJJ5pGxfKR6
9QXUBZVvZlJwnyqRQZCxXsf30eYSzjGMSQeH31gUsHovRGkwFndt76+G+btKP9vB
DtqyYJmgUhF0g4uwzR6PHsNXRqrdA7e0RBugEYe1bIFySlNmrFtuTgHNjMl23MjM
Fju3QV0GTGbbRjBfZLxyGtYm+pE1pD2TUHSBIH8VWQwrLyQ63/d9kgAIKpcxWsC1
kutog/iGlLDMINQQZCRp644WhgzSG82yyWkvmTgGjOSH1pHnOIZdgRYATfS7tCjS
kjEBxkWqQDKFaczP36+uY+HL02V4UI0yhAJKeU2gyMM/BezARd7fi0MO+4ylg3le
lgFiso4ikaazX88aBtoTjYiBrgKCC5AQUFc8YbPLCc9EC3tRRat9epqJhgaEPySK
3TwyKuQ8hypEXJ74QooYwRXhCVoIJ+9QD1wUWKYGIUOHg+Z6ceqIKvguuGwD3efQ
ERkGAcrW82lvMTgfPiujIYfDsKy2icbV460REnCR+827HSNmiypn8gRjUpFRGf2y
TYqJne5QCF+Ozh36HLZk+uB7U2EY5TO5o3erv1n4Q1UqOp+qT9V4GHgBqt4SBTdA
YXwDwNdefPTyy2snvcR7PP0Y9WMXt80JyqDuY35kN05QLR9WnW709XWZngaDqqic
55rjGv6XOEJAcbo8N7bI3VKwTVjzFQqyo2bs9DUrVOOF3en6i9DjsnkLrlJZiagl
fZCfYoTED3TTPmaE/UrqT8+B9QpUad3mKGIDvkZ5QZzgdG6EYXbqLac42YYP168P
AQTUy8bUGnzep5WvJYclRFTUhxp2VzWNdaeoFSWIodyuyS9TsxIjSCEAK+ujdxSz
H3ufHoGHTCz3Ecxc2ozMsvJTk++ngTi0Z485W5NsqkL5/n+A1zgGXGkdjbzrfgG6
P3C6yi1jhpsUSl1TWfX1r7Fw/RwVmeMznCJ7Q+qO6Hgk1Z2TGOCSOlf+AafqYXTL
61tEdoRA3T171bI0G/h2lVf/qh8Sz1dzWrIGneKtRom7knvHuMdSjD0gwHPgReMJ
r+8ulGq0XxCwYzOLoxKBorAwj5IqdkmAtO8TGyF0h5uo6+VFIzGUD7Xd6eKnJpwO
J+snuHkLijU+S3gU3OpFaCADXHAVcuvYj6ndJCa5b1Yai8szs5qEgUiraEpTQoMy
RPMmuaO2RFbbPuEf6DaAxDw8EkZtIHCViOhDVOVjIqiRkxQ/2fksgjY9Im4LVinb
OPJpoHnleIlj38CArxwhk9naZXKaFNm5cw/4R/UiHLVPAG7j3lYROoKuPxj8mFCH
xQs8q1v39ZW5XvYuqOc2+9n/ariwuGB9X2rbjMxHuGB7lNLJjY+048uEUMHjWonK
EMrW1RHEXOiSgsR97Jx5hfvkof7+1TpIHLn/40G6ba5e2Z/zTNUjiKQfo9B4dLdZ
HOqNYV6QRuP1P+A8xADa4qKb9FC3rkECyF/x67hYQ3Jqw1H6/tNNjKO2i7MBpEyF
YQZcTgJjkPXpqOkji8IwoFd1VrWmPNRngSbyFnLsLWnreGbR+GQpL0Nzemnx59ec
Tgqwf3NsF9QpZLeIDG/4F1hj6DhxcevAs625LSyFaj/MmhOAZa3H1lH05QcI4R0S
G/Ts8+bBbIp0e8CsT+cKs1UzUCHYJI8mgtdwWBoRXNFp2Nyuu6muIJs7anr7Ac13
6QyU9wTh6SniQaTnuaGm4MLFcwqgbPisIVNQlzeh++3mCsvAPcGMNaso7q75awPs
dYkyHNcoCQF3BelG/LeQzAWQWiLSTe8e0rXLmwzyebTJcVacEOcVDiqGxtqlMc+V
Kk72lSvUIUGTxjWspIqQTKcBFreGIaaEP/8hT5Xo8itwr50UJ+paX8mUSx3Zusy3
E2rLB3aSOhczvf5vH44GyjXxcelSytGBZxL0DeK/cT7W9vxmFUnr3iYr/POB+huU
clZsSUO+V7ZFliK1QLMyAN1xY9UQOezAAQxAwrgftxbz6cV2rF0sCHiQ++clq1oX
`protect END_PROTECTED
