`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6UW6bGn5cQSd1WgcChyP0RpHlClMGU7mkk6kByg9f5zghqlrx7KxV8NkY334QWSa
A0bO9adrGU0Qk+j5xyTIkOho3Pq89Fz35pW4iHQxo8m6HfBIJu/+EcZRzqsmaENb
ji2IYxJvgH09Fp6gHOm76E/MFxeAAv/cIKU2DTfkyLX3CT7tr69arie94/hqJ4Ev
UBCd7isJkOqrk5rCcJzsRK9dMvl+eXCK94jri+DPG/+KTuPwwc3qbpbWbLgq7SnX
aiDmzqAvnO7fSpvS7HTRih02GQoEMNetRc46sZ1Q3gzW4I8jYEczJ7c5kABbjmJ5
MzBnIKwSKTukS0msaifpZdkCDGZI/+AZQgXayYudnV9TazXMKTQ69GWdNsg33m7i
jPRzncsDDvvWpeMfVL0I7lMX3ql7MIMW5bOdb1clNHw=
`protect END_PROTECTED
