`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5/0mPZuDozRc8BZjhm4TfID0pnDuGeWZ1wk/z5nWSIJrR9f2JmRdumKbpJKFnOMB
D2DpJ+KYjZbv85kflpArMqaTl5uWH+b4dTBEvedG92DGGxHtFPRPsz9jzJJTwSZX
eXW3XP8fJxpEx9H9i20TsRoe5FBGeanbnyoQ3qjnSNunbsN4GKgWebrHh6nyO4BT
O8rpLTdndTdKAuCRszQvb7di9kkodisyzxYc8RxzzkTAoft4jhyLJqalw2Wm0YuM
/ucenL1eUuNSWlH8sGBxd0OBuRBPIfu99mvN1Wj9MtxO6vBK+yKiN3eI53gAv/CX
2JXhcvZWMcuJ0s1Pe8ttRUNNAL+9Ll1iB1fZ/ZV3hMYLj7xZt7yUV8LqhvKoTUvG
B1VRX87EHj5/bTVgOp57jN//MqzvKDzu7Qo3IEWzFMTvcDPaDNGYVXxTRWEWLMYz
1LvkK8sLzIAMoUHODk+DahSk6RIDn2JxS7JfhjImh0zUgfoKdiGVVSLp8rQDGsd2
g7U1jp64QauTqO+7xUVkOmbcpDkiL9zOOQCfMpHHmYRZ8K9Rx+88iGap7Gs1F7pH
GNtqNUMSai1PgP6qmxz1pR9Mcxbu3B7H8lwBPGL8d463q04WChIeuOYpWIQYnClj
dV7lO6YMkG3sdnQ7Vfuiy7pO6jAheK3sWd+Id+nsKFtctCX8E6rBTTYhOIMqXlie
HGOu+huMDxOWXqZk7gGKsvtCAhSAQbmtXlvTzA5seEI=
`protect END_PROTECTED
