`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7letFZfws0Bsyf+ynp1wCBqNUqI3EkEea/SqhwBkns5hsmKroJYhy3gt4ehnWhwk
C+3vZfB/M9xCrOP63WAbVauf+HIvZgZQjAZb1Q41lXHQjHjEkNB4vPUXsM276pfI
39VDzXVYXYagDYkOs9U2+bXc1LHGxSYl69XwaY5th6H0Cz6OwV1cFftuou9FyOrc
Ds2hReQkrdOu1nVUsL0owl9Xuv4mTC+rra23WcH2XPEl7UsKIvkZmJQNLZ2IAKq+
1ITOk1GPbbIgnDU640kLNcYYIY0VtjUvFQTiOzNmRDFu7/nfFVI5Kxg32vxT8tKk
gC2BaiE6VoA9II+ke2QvNOSQkxK6gDuvvcSjyI22nQIWghrEKW5i7/uxbr/CghQH
1OD+uA2jLzWDnus7IWP250AxVQHZ4wtrYghUeE0Qud/MSf16rDm0TBqM18grNpyA
eZvMtpbUuU9PVLYJg5Vjp1DOYbQqMQHR9WFG7vNZnSEtXB3VMfvHZMmnCCHtqiaY
v4Kq9og+iRkO5ekCeWhD9cLl9TaRVEuBiYZeLUbXLWJUUUMBmfP1hWieE4NmTPZQ
BlDY4EJxieHE6gE0uZIBxdUmG6C5PJmHS0mhcfuO2kxzcEvIz9phz6FggIL8qzqE
EdHxu/Iwi7ML8qWYjQ/gWZGCkmnyg83HfdlPn7NLVzQ8izwZEKqitxB+pG4hPfDb
pHFjg1EwfQzc7P3UWq8nFwsYebQJOdMMbCflAwKl1b70HyWTJ7xPatz/jRlOAzIS
NIsodwVVymP7zRiAkaMFzL/ePvt9oVIac0+DkkCEY8jc+4ad+GVCcE5TOISfnrXO
qL2FZLYJEndxlEgaBMlrEYpUAt4k4Cex7DT3a8rwm/U=
`protect END_PROTECTED
