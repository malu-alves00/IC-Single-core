`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zZHuyXpmeLQ8tUXdJEYNKWEjJCuRJw4kiyb/yVaxZjxjlR9FkQhv7+eUN327dVdF
DJ/N9JG+mqI0peblKai6pQ7Wl5zsetDZFEOLQqCYPN7ipfSNjNkdKd4z5vcKp0Iu
CyWuTmLWyI2zTLUEXlAdW9fYSKK3VG4psnkHz+7wEqxtw82QOTuX2SRuX3dPpakm
vcM82SFTvGRmfynKhK3V++taf/pf5f+bx5D59acEf55zB0z64XC3OO6Db0gq+pn/
3qvRGIYNmUegefJW1o8CxA8iMEVDLAIs+3bOF6qVZnnYBq/E5TIahJW5K+BrRVqm
JKHQdn2ZQMxuh3cehfkg3+59nTzjKS0eRP/JNg/f9JLiB1yuiqstLPx77tpuBp86
MrMLCydryGEOuOND8tM/4r6e/pwOVcZG4BL9Uk38j7FHP0blk6lBWvDY02rqJiL7
JhqtWL5DYPuVZQuw4d7NN0S8UH4FpYNK5OgTvCOdEl+Y85MZpVq8myf3Kr2KIhst
LSg7N59rFQ+oQa3o/Y1kmA4V2HjwiNJ+M5GvXC5+mi45ciLoVQIsBImoVrtl3F0p
Dr7i/rQPGtYH3V7a6PWFR/vIEHq3FTtVYPfTEeGkeSXvkyZDQDXPgCfNJESOGbkj
14e8M5y4LsKB7LMBqVpnAuqElrOKUtHyi7LVsmc+Ysu0R5Ve6RNvhsvTE5XuR4od
y4FSEd6A0evIVNEikT8B4HqzJHZ7+PVCRnjgmUbR5UgcN1FIJOTCFThte375yEGt
OyYsLH/45PwiDSu9V2K4Wv/bjG2voK8TfcbMZliMSjrySfN84oQAKL2PNnKVzJIN
LADB6HE3Slh2SldcXXHJmGliF+bNVe1dfYzn4YMsxB9Ku9Lyb4BAXMnl1JE5gZqy
b/XwsLzYMF8tgehrLVsD4RJ8JuyhtahC08Ys2mn0EXQU0ThxEocqheI03C/5wPcV
pndw+3MEkGfH8rmOlGaZ+Ug17F3CN8r/CGKZdAWpXJJ6digrfvZRFdEMALOu1PHr
fx+CfWyhV/ZpNoFEN+VxKwNPx4EyjvVFPsywS7CoFEC9qQXs61lOskXlCiCt9lDk
NOxe+To3qRAN6+PaEpzC2rWLzduZJynnQH4Zh8aMADgrwTZMWx3NBBKrqc8CLtUY
QPbTQEGlJ9xsoO7qo5m+nnXr8TYMB+sAz9Law3E0+7D5ayN8Nh29iO/mRPlf2x2R
4t3GMM2r+6yotDd2ELNDm2lYfb+yxIXZukPUcJzrgN8PlJBoonbUlg7QiFu/Kn/F
mj6SUFtg2lpTYGcFfPCvwIPZpqYQMHcbcAbTUM6eNVbAEf4wPmVSuv5x0KkTNhVt
PCGRTX925o+yAAUrnaQ/2Pia7nCjw0bxw5oLOcg/dXYULzGfAcdFjUz7gv8RbT8p
vwk0RVZeksOWKNDLS2ruvIvlwzFAiXcGE01gE19KbK/wq6iL8CXXvnO1sJc75Eh+
KV3rEr0t0yMryMtAJ38bkvcLCp3pAexElszkHSytUsLeQc8q0QlvO5YcSvHiTd4y
zmLnwvlTsLs+AC6qgC3PUS2dbqWjpTIvxURW09s1aQ69bxY9cj34LRvVyVd0C0Mr
IZqlwhQcJH5oMRecOcLX0wnhUpvmuidMOBKMJgOVSpHN2vxGbYSQorp03TMamf4i
OanflqcxYQg7xYiTXDZSAhqUgca5dyesP31oli2b5BhF18OA01MnZGb5ENCLX93j
Hc7U/8OvYp7sKWAAepxT4O1VkGgEoPJiiuSGsoiYY2vdsLBhk/Pa2exw7Ic4XwKg
BlvkdwA6ByasPAmxzo7zetqQQcJnFFm/Vqg34+ItMqsC/l87OtsghAXQdX+6ir1Q
XNTuhk+6930xEb0wW1f3cxjj4C8N+vF6E5GRX7HYJPu9ktZMMNKVnm1GxrrTomyG
8ymeo+Nnt0CmXkCLKlGHsl5AfYgBZUFGITEEO0ZztWQEYopuqXDXTrbu/YIkTULF
u5EwYTA/vgUmJnPr/4MWqCZ/oxn4N0AViajh0vzrokw+2harhEydTmHwOTkEuQxU
5a0zXu1UZ38OibnGbmC2jl2jOuI35S8o65h15iDXOQiwS8FBGfIZ/pt8PHjRQSMQ
2jfi0ngS3dYrL1ZfIaU2Rg==
`protect END_PROTECTED
