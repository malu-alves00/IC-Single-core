`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BOy4U5MBUI3rZLL17W8jSFghmxY06w0hxjcEe6ZvL5nPVJgOzvlBT3tA1fVUCphY
482ZAEvJLH4txLvippSw5lDrxbAqcIiGmxajPpx/qctnVQbTDknjNrGLBQ420bAd
kOd+HfcFKLFZBxEHvMOHU3lM5B59mSyTkG96lQKKQRh01k7kVDo4xbebpvm7Q62W
MjbDSGvTJA2pVmdjBsHHm1Z1fln814IX9BGtPGUBEE1L6eGalU0tDNo4S2nighAO
7DyZOE2EvmLLFvwL21Yehnj3B+4h1CbJkFp8HhpgbAtVaiF4qgQ8ihNabcQgPhY0
/QXVWRpkIuCG7tJ45pqh45aX2UWYDRbqG6X0DCuRPTnJW+x1yQqljQMK31LW2HSs
7B1SXU8o+6txBSHQOT2dimcwYmiicUINAe2bMfhvp7Hal5H+woBAReDm5AJmG7Qu
jl3ZGyUMvTZimyki/NCvV98UJ27h3r90umpdXxItwht2red0GQFXlf4kJyPdMhlT
GZpkc2SlIu6QyX7Vnd03CfI+DEAzIHW/AJJ3jKlJx/KZsVuiycY7ShLbjmdztVy3
L+R7cjvPbd/Vtc0egmmeLKie+aIE9apWp9DV6jRJFL0fDjWme0gE8/JeC/mEpv9f
`protect END_PROTECTED
