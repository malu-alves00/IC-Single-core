`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
q7t/pPgjOEc+nu9A93vNPCFAE/aLI9kaIRBoChzLDktMEVKab1nwocxqq8Jk3enq
aVLdR1aHXQVpox2dVOlD2Eppv1/TFrJzxRKoVw7cl9bGs8W69dClWuOBE1VM5B71
TWLvPfnSSZXQZj3Xa9rLUDFAEk3pbXb1cCUpXJzgbXbKxh9/acnHj/bfs1IbYzJ8
R2Aqc/I0RVdng/LsGa5PnvcPiCxjX6ExrMMNq6NO3GLe3RIgTFTbaU1hzzBB7sBi
HPST5sLp4ltSbxFXa12/Lz+qMd4urQm0dlepmNV0tjeKKgQEMcF+siQMweOL+VyC
MNqfrf3Tep4is1bjBNdqv46ZqNJ5/QTw2wyMjirnzPivxOvvt7TvOblHS0yjRgAD
X+0yUaXdBFSvz+XGtj8tAi2cRmxBY4gKCiVARY2btjhF2BJR0m++M8CtQ/xjhCHR
8zg/S2CHbHSuyMDfYD6xmasp53a5GMuHZqk6iyhYPJTy6HQve5JQGwW70MbH2yHv
XBr/dC4P+H2yw4hYf/Hd1DKvQrkN5a6gwl7woFo8bh+yY6FBVUwUTBS+FaxlgoXd
1o0eeTq1hwjCe0nC2r/YojgFHOjglD9q9YpokgIfFgjs4zfCqUaGo9QIpcmojlRW
6eL/1q//jhvqwfx0Tuny04ReWbJRmCc/+CfWnySlYiiRj0UCDoseaccoWeJ/yQEc
BcyOKmwBUcWPC0igm3on9TXqL7sXu36vuGqA+Z17S1YMsC8xdgH7kb9cGNM0+Vr+
+avyB0iMsWgC7syF0vEVO2XYoC9NKS+Izrm47pO9Bhdk8UspQN28Qo5XyL1OaeqZ
f2VmALuIDioMzCdTTKuUdw1jJ4Zg7Fb7CtFMt+GWUTKIzeZ0IlXbtF0voa/ro9tH
nS4yz33r5ABMECnEYUFahGgBPxprEjjcAfRC7agXqcAg6wcbyjAGWXsWQ+hfUHi5
9+dTlamkGrTDGCXEon1e86kENst5zugySxKy7AckA5E1g/sF8KSRvx2EF4IINmQk
G6Oc93TZEBFmqOCYupeCzhkdOM9lB8sY1/HERRElogFhIRwja+bNnW9qQP1Iv5Tt
y8naOX3UbCbJnVEZqlonPrLINPSolRKWk77bG5rK4K4OX7i2c/YQXXGgrudkpwdZ
44ERRhtX3zsqbvGC/dKbWnSXJ1XfZQA+m9qwTp1feSZXzjIq8fA9h9WbA1b4Hbos
f9s65mdk0NRmPu6NoXvwk/pF1xmSansEp7eDr0VEvR9TZwn9teQXDLTOmgc8KXD9
bRv8c9tNMSY0joVbuyfl2Sd62d6ZF49IzWmre9yYHGjc9ZT4XIj4rqHQonde5IC8
q1JdRbGaJhpI/FPV3W+Rc0uJ/I17uU/x0xKzkY+eWk3lGp4OXwObvuc0zphlD1R3
Xw1+y4Tcc7bzaLNdRAUJypcUR1dJ41wZSsLToKRkzrMYfUfWGDmA7aAcPZYJki3Y
2nebRJIrvU+PEuBzpKs1/DJ/Hc98sjCkBVEgUqQFN9jRXK4OBcexfZx+EGfjaGDJ
WiRp58IPD6/M06Lq6lU5XYk1AU1A4nsdCuY8aIaiRtoHpi0eLyvhgkYORuc0r4Qo
asAeHZZaUspuHiw8Omhnp773WU1377rHGUQUA/OLD09pmgyp2cy2fdMqfcDNDUWm
IeDxDhXZy+WJYVgEcl90tKLL4w+M7OJ4KOBykHaNxkYDEHou0Qkj4yF379aZdzZW
7eKxococb6AQw4knx3lGH/Jty7ctcmh4pYLkMTd74eUC+02++rjgIssJopG+Thnz
8WlaLxDI4ajbODclAHdxEgS1IOfRLudhnR5D2D+TVMVOUj+OQbhnGPvefyMkoVyg
A/R2p4LILQy57ZZbaxXCy9oHsbXsM75W9vwGqQi2/4Nn5Jv/qIE3ISHSHAYL1TEU
tobmRao0Mm8rXdepwSjYPRvZWTpS5oO8VogZD7p3QP9la6I/SrcNcCnwKzSKXsHu
VIbwhs+/DeAmAhPSzQ+twxx01fbKxTESAzgIg9i347OVd4b6VdpXBamXslQTbUwd
sbf2GP4jwZI2wa3V8huqCdwr1zfrERB51Qjq28FUov//JQpgspIPPJUqeaz2mFSG
a112g+Gxgy94LgCCjstCUcvSVs1KY+zaFKTHK3idH2XZaYZe9Ulb7psBceNjO9pk
yd+D84gG5kNKT7yVIpdzjeK4vkP7aC/Y/UFgrGmwocJbpP780wgAQhv0r0EMIP5H
ySSo1sVccA+xVZCWVeO1zYiwiXwzifqMjZ36Rz2kyY264Cz2yMvb4DX84tfv7ftO
1+unEkwdi4PuITt/VrBLhQ1MdUvr3BfXE6nsuHwYJXcPLpVa/TKWzTZffTd6qpI+
55lGXwCCEg4OFLZWtQUAo5c9yjzkqozWe7drmNhQHzlHN5X/Ewf66i3Cg/XnYKsL
EBrEC6PX5QByu1l9QzfF3sBRkplQY4qcfkqPZskSrrLtfy+tcCrPm6ZUW6a7aEjh
ICjo75aXcVlGSzkQ3SKMIw==
`protect END_PROTECTED
