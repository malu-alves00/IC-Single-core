`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+13iODk3rI+kuVM2CszHqgjefWcmSJSuO8QIdcLh1yW3w1TgkOcsGNDVtDviAt0N
to94dhXZVGxN/FP5T0DlUt/dNOOvt+miTwEdyAfGOKDf55hd248uOuq2qnMXRjrI
ghn1yd8iaT6lyGkhMyzr4NEQdpP/12RsM3Vg34i0fDRyPLp8gU1qumekgS7LRFUS
2AgB3URsGHzNdnyBk03aBlu1j3FSA+scaR1iMexJtNqvmX+/eUX4tWl3MiMeX6De
NCzL+ERomvJ4ebHUwLCVJDoRsP4OgM21M4JYAfIxxAfds8oeH5O0JO4OUHI1fEhS
O4FuLUDedBcmC+8X9dv5EzR30a5FjJt2kC8LK3DeWbpqY9iqV3cmPiAtaHwo8fDV
JAmb0XTlbCWr11dZ+2UP0oNH9sc6SW5GiS5FfTNp6ZtOq6tP7EwuFQW9a1YqBtt9
w+SjFR/r9EMidnGFjOpTmRJkWNwvO/VTf5Jeh4EpAESdWTu5a1ZZdnxUeMuDvs/w
KYaPu7eR6LmoL/TnpQ3UcEt+CqBofQTqA4k8UVZHUxyRmi9/DU8TiPJCh2fKbuBJ
PGuy9+Cea5e06OyeSF9I5CtPzP30V3dHyglX0O526A4bQ5qVG8mcNoNlkavzCuRJ
gSLIRM0Qvf0+UZ4U+HW+gfktySrGwmfBc3nmlFiV6fnS7vi8Fxmen1hW6rb5+GJn
u7X3rYoC3S6uTVWTZktZqBTH6+mOdJqYMICqt/j8+bFJ0hQvi+0VOk36tm16P7/z
eQAFaDf4R0eLTXT0wpZNnHaRX25p6+AIFkZCKezodpl0gFZo8qXIXYzNux+aCTHG
pwK2W2A+m7UV/DVUDtSr3w==
`protect END_PROTECTED
