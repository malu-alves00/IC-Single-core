`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rAI4P5v8MmmXxPdWcVy+VYOwbp4YXMh+iPOflv2ZPkrfyDpOP34R4iVAAwVBchM2
yp9ye3xBYzWWXtS0oS+DDnLD/2bj6zu2/pUkYGO1z7gPv7vJNTA9hmiAZ8YTCgOy
5qI07SlPUdSvnQzXfumQ/wnzOtGRoVamKAH4uLYfb1x7VVggWTCv8eYL1z5OxZDf
0wt+CJ55ORCCGmTdWYzJLe3Ah7G99nFEsvntmKDGjNV2PsYzTgcAXwa+OWHribM+
V77ZItE5rFtKLoHIyHoJdKW/iYzmQ9yJsqTJKSFP3DcHp9FPJSS5/tMiCZFaoOvN
/Fp5NdkaTznqQaqTasnojRzUrLL7vIEZXleZtOdVHmokxymSvBJg0+esRqTvrg43
m3jKdLrSMHfrZvufRS5ifYLxkJmVdSRssnZjBOLjyfTVh0Hu0f86yXw8F+TxqEQX
1cPaTLCvQx203uRG0CpJ/O4yxTFdlfPXE3eIbw1zzUpMJlysDPSWaeqJzdCESlJf
xOFE4I9X67zQBu16mKdp3CSdc0iGQXlCkG466LQtPTaOAU/uLeGGh3C/SQqTO9BE
4iP847OrDWC6fGPmjdv2PtJWPxWK3ktU6JuiKo+GP9YAYiqrP5SP9pH20sNFayEd
BVx+lrd6o2JgKtLvEf8sVqvVum8Zr0AAQUW82G8+He6pywJcIbh1rmaNItv7GjDI
aqp5q+IoNGRKwVpDZ8chUfX/myqyQogEqHxvaz+r77ExOsFkBExYEJznBYhog62D
79zbKZtFhMYzsuxUe32MvXI5je680bBywxEkxNornWHf9k6+C0SbJbCm6muhp3yM
1n78aaObtFEf3rwefTYOawptVprekSlcoI6KV5LZyQ6w6PEkVCG9kDhmKq1qmtEC
kCCYsR++A+qSHH9cl9xUucdrYB5rxB4LL0P4QP1NlY7l+11W/mGr+HHEoEhePtAT
h878odDg3ZD7J7dyX51rGHB5W4XjL2DDS8nxUFgDpIZamJ6qef+wdnub8oFs3sgu
vlpN493mdCxA+Nug9knzVv8fp9uf4xtYeWZOs2jFLPdxYdxt/F4FMuV/fIXpM33S
cSFQFn9TXmkpPRVS1N2Z5lAUu+dHPOke03FOEMsWSishd1WTAtPYE/v4HLx1Y5J0
Jb0qiKaUgjUoa+zadA/fet14ZjoaM4thLBICV4OGmR0paqS3HMaqObQP69JPOGgD
1pBeWJwg78oiruzpM8IgBYlDvW0FgV4WVCwcgB7F2r+n6Db13OKPnDSzli1NZs6l
3cJZwhcA4fLunaXg3PFvQBunAuNn0KBsYtpTWnPiUKeH1XVVAh3Q6JIYkHm0UGV7
Eqxpqq4nlJzspntQimj6eNDApDHn2mNewqARd2uLbItvZZpwbZDYvT4nYuFDGHmY
pW6AavtccnVpbPjy9IXBE6cSu2BC4SQCHaQLNTY2ln/zeU7njtNtUAkglST3EeuE
vS0Cpj8m/qx61T4WQGkDv0Z0VstruaVPv/EwLJLmYt9WyATwLkP50jUVL03Q9k2t
1CMQ0lavpWUB6aqtgNbLNgsG82/C8XEw7HMENDMoVFfS7aVK5drkXXmBRlTxWS9h
6QBA+7DJ7eKpfwji84U/KER7kASTHN7ND+k8HxuIZucWQ4XX2AoEOKWGR8ySCDcl
VyB9p4EBvCXl3SpMhrp8UZjBUPRj4cdda2e5/JXUC7ckvAlhMSX00L+WbjFV34hO
esyIjwyxR5K/7cxiDzszT4Mv7oRIp93OIJyz2I4yr83GLpXmLWhVhziWDNgahQNM
DP9B9XfD8n3/LGMpS4FLk3KpBngPlPwzuOkkeEJY6waX8yTZHAqruVwSzw/OMQdq
pQXu/TBg06S9dsGpPcspFAdDqgwzymrLKu3vm83tbnQQUlRyGczbJ7TpFHyVnL7f
XI1991RgkzZncuBa+x9Ofz9KW2Y8tij4X6MGKKUSy9Xnc7rtMQeqpBlR4bH8d4Xq
oyQspwb0Qa6o6NubqNIOYyIOsJ3zHTXgEF/BaK9t2q49lhEdo/OguoHDoU86Ypzj
cHpWBKiGDuym7681bTlg1nwFjgU6hEoe1l/Qu3ip6x4jJmSGd+jtTeYHDEnij7gB
OeDUPId41Yv8Q+MTWYvKtbiyTs5VdILOnXlZ1kCmIJjuJ7CzHUIn1jcbZDSXkcDr
So9VvcS0kpPhKRFbvHOQnog06XkVNQWlhEIexxc/hVLYJbSIwwCAInNdvjsupv2i
CJYs6LkDxAKnWJ5SHte6VAwoe7Q5WTJTISnMyZ0HbhN0O8hUM1oPEVn0WUr4faKW
BiWxPM2p7AvbPRl4LOUkR8p5oeUFQ17qTVIpLzLbkuD+YuMrCE9hchal8/2M5DHe
CB7h4MicjsQnrr1gJUZ991Gce15Jh844VDMVmvyPsndI9OKtwbvsoh+yv3Z4n4wI
fAs409ZUDRPsalqahf/3wt65RHuxrOjA9mIoUkrGtI/bGdsM16vYTfu7AcnEFdGC
MtuhlxdV5cMpivMFHf8bBct7w3mqz++OuorWmE7D8x2L2Q8dw5hcQtTp4du72osb
aG6Q5V0LWgZMA8EXsJfpeniqtbIYf70uIaINJXXH6TYL3TzX5wn68YrK3Yztcpdv
oKGHiwMTTB6hDad6ZJd5aT6EjpQWMRNWOLXDtoh6LxXFVpG2hedJOukcx5Tti+N2
DOINf/61fiHRcScuO/UOhLWn4VZ2LddS9By9gtbPVBmzCcZHRZR6DSMvfrdyPZpS
YVmNN0CbciTbG08TKahzymFW0SjvAAPBkWrFTz9zzvR+P2x2CfmSDawLuB9/23rf
SJPEeyHktfCGWKUSCDFrOxJTOyzzNd8yM/hnNdwWbExeoiqq6HQ2FfTJRPyAwGeX
Cqn11k6ikuoouW0e0yuoBDnrcb4wqv9DBs9x/eISV/aNRGM8KXmFbOmgPVrOFKH4
ewOl/AM3kmfQiO4NpZ9SA4tDFpTvSj7DslUdU1+5NeUlqWVSzJRfcrkV46i9BPnZ
p82h5yPpXMT46Y471ng7bZlqZUFVz1w8xG1ijZBsqunYQ09kNpWfhz81C79MfSUI
BAIlnhwaTI0KbbkzfQOei05kFQxdEjoy1yTff2rBJjch+inWMfqmdqQAxrOxVnf0
0pvR2hF72uJpsTWrUThFX10fMvy7C+Z1Dj099qEekBXcUj/U2sIVru2KZMdY8x4J
x1YVy50gcDova0aE8+bkM7pqIPpiijYpDehGc9PMs2QrzbRwI5rkj8gmFS3rP5p6
mIqihfeDfK5QBmRBT8GyHcTxokHxnRyZ02jRfbUPhOXUQlotImTO+Qijew2isSyp
fSVkZfZjPywp95TdKwbMuAVoKdMyZLVfhdJPb1xXuY68QRIhfuXM83Tcagmzo87M
AYoy2BHPYItr5SnC6RY4hj4/sGyQ2st3o2VZHUegI2o=
`protect END_PROTECTED
