`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9cCp6n/8DqL3dVN8cv80qC+EBqDmYDC7EtrWUD/8zMitz5oAnTwfVA4yFR+qiH68
tDgVDZNyeUUphYgHmmVXRgTAYdxxBNEQW49x5t4L9DtLIa8ARvqfczjUOMvaNcJu
EmRqgZRH7RGQxxGct/7uvh7YztdQxLrnFYOVk0TL571D1qKy4Ypln2R+PilwYNzq
n2Q1b3khGj9xUDQyq1ogkcd2cct+iQw7CBUs1s5pC2R07JnngHU2fZ5jGk3eYfAt
OxOmsBlBaPawCgjpauSg/lZum49OKdgeF8bBaMF88GI9DW71UPyv1+oNKqBSFMfv
No3dlM2CfjEXxM6dkIxO0a4MKZPKPQClUtudnRq5ySgMLXjovwA3qGP65SZVJOZp
c7SpoS/n7jtVY2SF0xRk2Lsg0+w5HfBuzqGGMfJBq0DTYyK4kPs46C6/rPCR7mmz
SO7NNN+phuAtRtrkQL4ROARKx3VvKsdHP8QblVWnp2dIbWc9vIut0mqPQL7khSII
fENpwSp3awzZpgUMoYUV5lfTq0zuVkqN4YOXKnrDgI1064zwj7Pgt/D4QpTHuUdE
IOK6MVEddW3DH1a1iKvkVpYhxQj6tYIpp3XqlvQE8sbRf1eC9mooK5tw1sv/iAy2
72vWvz/emJIXEe3DMxO6UDvS+ELDqSzcgtexLdmmVIgumGr57+G+XZBcegFPaR7p
J4HJkGb4Ra207UYVvnSh13P2MekRCpN3eT1keHCgezDDHVQP0tNSdVq7ReRJQffV
yMaACiCNgnhJAgHg+7aG5XK9URYSo88DGJN6e9PLIWGl6M6IKjcfAAFIrG7WNkA7
BpUsL/ns8xPSJ+E+/+q+A5xKFPtsO0W6vyPxNNrt/gXWKicsDSx6hQXFbAIJeY8K
KGlQmcFgosDKXekh3+Kd59rnIntX+IBxLsNdfnyIBVqaF5EN6HjIXaig3o/xgCLq
TS+9a/WIFK9xZYU9/vqGlzCYkqkgKaJVBrSftjWFnMa17IU44z0UKuJBGaSgcQMS
ufJc4RBJo6/5Co4zUxbeczoREsGo9j75Cgw6vgYiO578bggdJSq7DT5S6winlXpa
doWGiJWaR7PdHQbv3eOHr9J1GBGFx0vgzKGzU83kmMT/cPEcWAnaK8PiBbLBzxN6
wcg8ldjP43KtN/UV7QyC5MNg53bhS8YNi4s9KZx5+q9dtoJEoXBLmO4L0CnbiM45
+5+gabHlOd404SgdwQF3BndZTufsHefBSG0KVXitYcod1ZzlopbZFIpFU+c3TK6+
G/lzpplB8tazoh0kIK2aaoYuqudDNF/wTwfk53TlAKQm5lMdAuIDIObJDt5tt6hz
fxsIBFMZxwjuazMvSNC52zmZIzAiIvU/d0+9RfjLNdD2o7cKTujIjsqfEnyZUbPF
v6ceTNoEXbN9sbdVEycCib7dETVbEs4PI8kaErvZawzcwjqampUk2h4LWY96ufBi
8cedT9U68r+B0/WVHPrxYapTC6fta06kKRAjABUEgOV1ItTKlK7B3WuMY98HYGg8
5z81YKKP8yJYULTN02JB02uITS6qaE4IFCTEa3V7t38u+0Ed2980uHTSEp4tl//A
B+g96mQ/XLtCr5s2/Gf014ONzfj//IUPGFyDvN1JRnpxAUhzvNnRt2EUz9cDiVmi
ZrzN4zVvJ2y2wRRli6aSXZsJOQRQC/o402FcdOkwNS5EnHBbzcvBNlpK4ZfAn8ac
uaxtlEw5ZmQu0xyu+d/3jqpqybfUXAY+JuhBlVKHtDNMDVg/UQL5W1A7Y8rCuwBr
Qmo/bMNFEOA6LxHcs7KH+ye8hfUbkvOFPZePnHKtLQic591QZ8mPH1uPztaiOauQ
if7bHY15xIqwI0V8RnMPiqhj3imxdK6jtg7hzUBb5ONliwWUVhMOkZsKv747wwgX
YAHbnypuAXytzX22uts8gchuWW45uO9xwkByiG/iJFysSiiDJFPK6nUZ3x4T1Bdt
ojWT082rL1pM770CJaDoz7h+NDJPNtKYEvpuGqDpfV7uEJW020scGfs97tjYS61w
VqDHgg/dkgk3VmaNy+Cj8Hw5JSgjmrzDjyGKoUhExRZ4JOPEbhxVZA3TlkBNObsZ
z/c5L3oovULgzGJ8IVg163e5N+epegwncXmNfHtdNPC69l7UjrpWUL6K0/tDPKz7
OWPQ38O8hmxbe0kQK6ehXk/vX2lRTvjgJlV7tcqiO2yuSwmXkLL0q3SU0HEVOOT1
Ys7C1oWccs3IYqi4oO+M7tpCFnIWkHkkQ2/ZRVFlg3L0AhLu6otOCL+DHHem1EWD
bz3UeRE6Et4G3seTWuT+COxHZnGDqK4Ae6fdazcEpp1LyIsV1Br12yalpTgwfas7
avXTkIbp9B31/3gCfTLFv7U+MxKFUtCe5AAqRzHbkXduW0sDIkEdMTiLBenK3Ogr
PlI/82z7BLfdqk9gYkE9+e1JRbCfzG0gFEFDw4PIJYq06vnnxwGGLRRsq5AwS2Xi
2XjcbDeMnz8Vr3HuyIUtvdu2zfc3Z2M2CtVhrsf7nn4dBI1doVXOzzDMAACdBn32
wDaXXPt2mh9uZP5U567gTjpXArtvMDMnKwMXiJQR7W/JdtkqRzS6/rL0iSMEvL3G
SmHHBqWTNDCI5XVuQV0NfZxw3iu+qlXRV9Q9MzawURcpbY1Y9T6EuJYmucebX4ux
k+wBIPLmsOIEyGAzLxWQsa2aIrjV2F7gat0IkgQH8rYzmD9XkNIGJqgDq7HNYQnl
DRAXJdOqby/bppTmnL0yJNRmw6eaen/H256P867MPZ2+KS4Pafjb+ny52SWbVd8f
SarmOtjsMEif8PHlms4Upcu5GJRguCh+0aS2FTkgrn7eFee97AIK3VBkcgHlrlRm
2sMeRzHSLch8pqJ3boHHI7p1QxCFlIRaMe5ePko6RuvNu2w0b2JYS8x4gGXSciAJ
TEFCpz/ZWxqSn80Fec+lcWdDFlBo9r8mJoDPekokwWU695gQv9fkgkm5jLs/m7P8
GVu3XASq1fg0VuevRMPwUQtu7Ue5QEsMR1FrQPsZGpR8KNB48DudLtESLBgprHgY
xSvI4ZI38mdHBgzWjpe38l1lUCpHWxlnO2156Bnt07itDoGpCWqRzVeyDLzlgf5v
bvgpUy7DEpSsiZKxAUqLrq6z5fE0mN0ntYokb7mlVAbZli7B1uFBOWQwj5APNdnn
Mlt+z+4H/aBcDLvpe2an1dLkQ/9yp18m9Tb4o7vIBPsusnEtpsnHABswYhF0Tnfz
8oC6dyDa506mqLEE0qVI8wK8tojTEfV89WhQIUe7ByC6cIMQW6rcQNgr0a3L0hqS
PcIlH0y582eO1B1zZ9G3m2fb2BFKzK2eVl3NCOcPBUe9dKgMpGjyhO66/nfCjeP5
u/qJ0nQshayuHsCmasxLpG7JTWAkM2dMcNps8+NAvfrWsh8OKcq2oVa9qvqRGOCC
ESqKPbTUPhji8ZI3j2V8TvTt76Aw2qi458/MesFlEf0VXaadZGEHtn8KU8O2nxjb
3snfZmRP95sUE+1QTDIrBN933jFya+ne2hsdiKRDJ500W9QzsJN1tfCsTgR8KL1P
H+28k0rXRPum/63BWoIlAbQ7i0J2Ra7ySI4UdmoVpKLUILwWqZQNxiDrsmGqTt/5
ZXf0R2D7/fBuuc5H+bqCoCQteBjCMvhxGwKUrZ1bpoBGRM8goHcEKc+vR9P2tFEo
UdTYHRCfbe5QABBbTR4EyiT+ocD7zYOsu2e8NkSRTHJMEEp+ZY9GIDYzl0tV4Pup
iF7e3trm3nnZoURNKRwcfuJwfBl1xLM9eiqxpPd0VePtx9psD1nFD9hr6H2W9gMe
+cDaR1168whRQr317ABB2GW3Z/v/JJnE0Q8tvEkJDVPW4d0FrgKNZJV0ZO9a+7Ul
NICr4hB2aB4wZ23STat6B1rqPj6Mq9RMPlMQN7UlVDj8swJvBDzTu0h3mlxZc5Qw
7z2NF6XRKZp8+/gzVfDZ8U9wHxtM6Uc7tTLXeiuBn/ita4lTK52b1ggUMuom2F2P
51u5rho9t/4uwEW7FAoB1RJiC8ftjnh9MgoYyAu8dhT9PXUozD/6zG8x7W3HeUf2
1BEcltbj6ukysvP1J9QQS1DKsVLjlMAte+xzDNPvqGhPUQ7YaSEaabarMDFGHV4b
MZn+fzCSk+Z/juW1SH01Kg9+DbN60BYhxTed76BXVi6HzE5a16A36J9sReVbdT+J
Jzw8agT5rsk/BNsurdYQLPTWQPSpcyhVARqR7GHfgmE3Y/svTJ+WDXdRi3wQc7fW
h4aR73Ttwl/AvSv8mx/Da4Xet6fVvxrhDw7ZZbtXmRbenvZwrNqIm/6+w6ZqZVC1
c0L9ilWFFIFlFxU2mhQ/NXJkpMjHVNe7OrUgblF7QnBLWdPJeYS+2sivLiEOgzUh
YUFBEuRgbAlNz714KM8CsWyoIAwsV+adj2p63RLTH/mG5CuXh8olmVb+/0LhDc9s
rr9eHOy6kte5DlBxXkMDBx3EHpQQh6c6nJcia3QxrSIJsMukbHO0RbZ/ipwqH93n
LvIxHut17WywLD+a1SRPRJp7/E5SgT/4wgJGxEWc/z9I2UVMDcspCB7OqaAI7qqV
eSsOnN67t3//EZ/+lvcqJrrMYa128RkMiG21iyeSaYVZoIyd8LQl2eOQfzAWrLRo
gy0w9gxAFxaontCBt1I6ZkKcxfVwP+8d8bQbgXhdLv1d9rHwVf1r+fVQg78hawGf
TvUKBFe03QZR5Gglf1BRmRus0DIU/fqBM0ZNkLOg6MG9FZyE9L5bPFp6kangNXQH
pkdJBCYF0LY81bsFdL+2/aJ6B5C6uCGM1nJHSmvP/Mgxxemu4eOrSSM9e9jhbTHU
7JKEWw/le4deWMn1LlyuMqeKxnoOTh9zsrP2V1m1yunbU5xcbB1rmSGEeY8Qqss5
eNnuV4RuHWjDF8W3nRG3TQZmrkx8GNGiVGlGgxx/UD2uwgNr2nAoX8mhVmHEInsZ
L37jTZMYtvGlOGO/fAQTmOW876KWTxuZ1YxYMpr6WyQxRP5WprygRzw/nFuQXvJl
U7mUWtmaN3kSEEQnwuvFTufzBYcyQQO9ycY3pTW8NHSjgTAPPkVU89YWNYBrEX5h
OFX+1XxgO9I9xU6JztyWkMhOYcFie+7nAzrIE4uWjkg2BHJVql3tIABvcDUp2r83
sQRmwRHYyZSvk5ZHIaJQMwKfSI/7gdNtmCI/YxWA0yFi5qnzSQu+FWqSp3c83Bqv
QPcVNtyJOQ15yUNYGyhxqs09oI/amWL6AxYAMeNAi85/HSheeruilrKb2ZMVyAFR
A6t85dKYvd0nhXMj0q29mlAY5/XqkBi0ycccHN+qhdbD/OrnyT+MvC87hvqFMwJp
c6DJdEpN2JrUdXoxJyodZzro1M2HppZKa056jug4kad37y2CP4yQ6iKgNOKKQ50t
ccnQCa4N8uT4qVyP0UyztCSVNV7GaaN51xtROEYUeHFlZjgA2cfhi3QbE36x/rv2
X5CyExZVBD+XXOnaHaQQqFLvxyd6AHanDvZzU20BIN0GitHEP5w6w7Zxwom3Tj8X
dIbT/q6WdAhxOwf+NMHlY3pqWbSzGM9aIkRZESLceqN18rfu5R4hXxlOowEwnK9y
vsj36xfTOwdN5YuqdRPdKl204pVF01CI8Bonz/vDN0qUv9bfRFgNYnu1eJLuHOyw
rzXE1ID4i1gyqfF5OltzivrIBOq+peiiOc/8W/4DwdkFRSTkknCBzucjVec7nHCL
N9Pdys46JnrG0gbxJYV3NcpxVNJAj2vszgbLQMsnz7Wyn/PrNlTsY5CHmWbinE7b
H3Ug4jMtIzH2ApIGzIQJ6MdbkgoxOASbbeb55hZdnQgBq7Jz5AO4X3/tfq8Z9T5S
8wy64FZwnlXtTCm8nx/E6lsn3XtVe3BNSt09R5QG6ddHZhffN01QukhLfW6iNQjl
5UDrq5oXNCzbubWLWCWadBGNjkfiO5d5ZlzeLbpOcy9iLt2u6HEYEi1uKa7+msAY
9KnnEf4PnszELqVKIfs/kLl9LF8JF+Vi62TnsyFE/As4nuVdJyqI4e143/BgukbL
UlvwFQS51H5yzm5aFeddIfd1Jj7FL/9zDGInNS/bTL5sH/kZmWym1HSdAn2KlEcG
LxupiNmhk2XObbqGhlHrUf6ObEPtxK4C+St8h0lVFJVo6zqONex+rfBfuHmQ2gYL
DGchnFBQ3sL8j+MqF321zWoChMz33BWyyCEgU8FZz53HErjYWl4mgJ3v4Xb76DIa
NLbDZccXSAGzjFtj7hEAx5BDVBgjlByONrnOIK++uKMjDB4O09ApmNXEI3FGxyFm
YztAFwwZ2zcJK7s942ZBBcVFqqhQt1Skn1c52figaMUp8gjOmqxJsJbjXH1M3Bbh
NtjiLOLtEMV7+X07HBlG4+Q6Kxk3hmBRiPrKs7Fp2wx2qW1JSQo0vdmZC3Ej05gE
lSw55GVqUIpSYWlHylnKaeOE16Xkgt0+75CDhjurdci23mlTsTdK0PuBrWYVJT9z
EihvXAxg+tVZpcozdZ9yYwXU7ORMM66UP/jVBKyQMu1vMetGrQgDvBuQb1w0HFjK
wiz2LxR8MxqTKdZiJgfIg40C8DD+am1YyA9rEwgCpA5jYPFONFoH6MXmixAxRMgt
oar8M9pwlIsOaFYgjxKXIs9xqA1rD8KQCJUGDO31nC1Hwj9qHUWyBF+GyTalmhXK
8JC9RtzLcieQu3NgsSDPOhdrmvDD14FEoLDLY3BP9mA1dOuNARhOTx68hmOyA0VD
O6124ywz4PdiLh82mai6nt5vajvbnVq0+pZIAKBT1Y1Ebi4+bfhfj4brGoQ9alAm
HqbPAHwx2/jQ1JjJr+SEQnJj0lyV16cMVvPlTkxfFjv6tat92zZDP6rTnPS5bip6
6i/aKiJEPuPZ/mAPHBS5+S6IO2IHkmNvJWCaaVwyRpcjKRmD+/lms2ZvKz8gn/xJ
Fg9ZwyJO5HSNmSCFesG8LLOV2CYL/yvCtt6+Uo2n8OMpTjRsYCVTK8+2zY2Q2bQ4
o40hPF7WXEittM7VaI69Cv19quinkGcl46mKPETeTx7nBYTwEGkFMGzR+vlvbpzi
ahN24uf1oLtFvmCGKkTnmT3quAiFGagE7ePao3UaPbvKOnlCh5Ao3piK8V49UTpV
N0WLlCLT72Lh58AlcOB57rAzZbqY5Shs8MsydFqGMSpJTzIuqV3CFZv5ET89Njuu
Z/7hNrZGGYYL9GYGJpPP3d+98PSgVRhrM6o+U/qPQ08aMCGEilHifkYG8wQLJTOX
DGEj2i1NxdYqteP4JTDWK8vJbL9e5faMyXZZsrnYAEDESVL2Ta/vz2caIHtG9fdw
gsJPRcGfOo1bVsc9qbQUgA3sGsx+IS01tamzRXJwSM/IUzv5IZZ2tD94eGSnxEzK
UaJYhCk/6VdkP1azJ5fXLoR0R/UfoLBj9rbLD5Fy2p56AVY5Ynqk41Yv4gBf8LMF
cqeZB6QUDUOATbPOcwVTvs1/Y8Mlc4AqLztTjLPNG9RrwWKJ4HMcUY0Om3Cnzkpr
04HmTwAnqKPO+9VJ83Vdp+VVfNLKUj05HlPVZQeTwJBEsc0cK/MzBuFRFzZaAdWq
ahnjBNlD6kj4QzuZSoW3iN83CGEac5vDe8qsyNA8VDbvYfkODY7BEJrxYVsQVtQC
Z8TR8Lq0kdp4q7ahO5AWs8ijVclw0+iYI1y8845ESE5eoAzhTkuT2YeQgoq4xbS3
3Oap84icmzpt+SMkzeO38ZbeBojGpagUQLZV4b9rooZ48IQ/slKN9+/hwMZ4HA/F
fcF1rKlR/yH3LQHbkI2EnJnF0EGx7+39sEtoRTXI5dVFmihP0t5GzKBM4zjhpViC
7DntR/f6t7CZfws25Q0X1JWbtZShQc2jsrjeWqsjQnQn6zu/oeet4colaOb26HYH
siSRvUsrfzPsH4TNnaFaKRdAuVnyu2SD3iXh9oia4DOq/WdBp5E3M7k8aP5Vv0Cc
IhcL3WS8xZmdMJLHEH60yj3iogLmuc4Q8y7peRCQIucVHPIjiMwKH5vBHuD5MFip
h8o3po7ADYIwtiPrM04SnKvCrub8MZ7t1BIOCyukxO5AWlJi3LV3krOphJjRTZ69
QhLgIjs/x3gyLvMbO03kJwEP27DRALV70+DUlthxqWzVH/CDFXveHEbss2/gSb9I
wLZ4qzrqSgAQNxX0Yx7F8w8IoYLNWZkCfq8mWYeJTSNa+VeyeQct1eNa30R+OOob
BE4BmZp7tpX4PfsKcxDTtjw8h4KMG6cmyneRgwtYGsy83ozV/Xiw4I0LYgy9L/6B
bRPwRjTBiUyHJTjPIcobOvBQY5RFQ02Y7NyvPM0U6JgvT417QIMY2G4ECGVfgThF
dge58q19qdSd3+h1DdfGztBxQ55f9J1uUi4fsyLt1cpp2Vp2euxkFaqjhYGUDivM
cNkNUm+NdCYPW/elr3jzv9EuxqNJAuoM+Esvb50m8w75ML8agep2HtC1oaTzL49Y
FvfnAqEaSwH03VOAEZHp50NiCxyjtjUZ6fUKO7lFMYnnHUCudrsVLkKph2h9e/7O
hK1p6NOR0/l51LNGyl0aeh40uuOrCX7PVtjbNqnX7D4M5eF0ZiUBuNjEPFpr+mMQ
pRI/RBECmCJ6p44sAMxIepUqwPjXJfkY7gLmr5NFSXQ/AdsaJ17Q7zOW/rItivLU
7LfxynfQf2aJ6q4xID1qhM8WGCpOmH9ufg0ngQAGn/YIEkUj9r2wuYlNaiegzz8C
FYAREypwj6OVvaGYDPkd29fzlb4MK0yNiqNmQX2PDxb0l8JD/w2xJixgWL7sLaxN
YN+OJiFHE33pPORNArxykdpGOkrgD6udAtxYO7VepYPSSETxT/Kmz1anTutx+WS5
wj3vgdMCLzEqK3LBq+Xzt8NBwOqaz6cB8v02MXLTV28kb5JH2StqgDuzn1ZnpnSQ
PPx9NZRzEUa3pYqRZ4nDhaYEYcugts6ofN92fv/DySZ7lVOv8Td8XZr4iXRHFbTi
X9LXtVabRMfVXiOW4+5c1L6lB78d0ryBi01vmnC3ZEBcojzkpoGCNkTgvHQRllHb
BjbePd2LNxChcdlmVvMu0izUmLePEomWtsBUGDiJ88g9P4VzJ4SaTGkd09AP2Sn8
vFMVnF+aiqXiuNpgEvVFpvQVqXubsA1shRbMk/x7LX9uewLAc4Lgg9NAaL4kj87G
5zTH3assyKzzjMHuqD8xiiJzL7E84SwYlbw+smb3tiKi8q6vK1lyQOX2ncH8wzam
l46BYjThakXpUlWYUkofPWMfXGWw0m0C8SbJB1nP9lwd75WOm+3d7blFsKe558V+
peiD5DF57R4xHi8zeZCh4QxcR5Wy8o0Ad1BjJXWCFWLLWIydo6fUIEq9uyCTJ5il
44J+7FaYePxNOJnswhtWPYk6VYBYgO5BXWTS5yrtG+dsuZVPoRKZ/pekOODdP0/n
0+CVMW3CRwkwjlMcJxVmEnRAdvBAC4d1arXE9DmvAeKIUAoipX8QC4bomz2nfoE2
syPNlJE/bSw5jkgJC66QjoLiGKBleDv2RtGT0GeEtowEWJXNDfvy7fVV5kVdbrOt
7ylatfWp/Z3qopCvKOmrPrlA1j9Z2efLprKGfTRkbvB5qZn0WJu0dMF2lSIbmgxA
`protect END_PROTECTED
