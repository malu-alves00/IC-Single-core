`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MP3RTZSDc36xf5jexeyDBX7V1Cf/JnHr7FXoQVh3Ci+9FG0rLqnITBTwzs/aWyvH
4S2YUeCBaidd+++/zuw9eSbMxPHFdr5S7XE0CP1tXavjTnwJRiDFiJMhZHQjwVDZ
qATQVlQ2nvkDQrhPP2/CP+h7nk8jsQIxt5G742iFjhtMPu9JseulhJ/P7aTIMkTL
DAMRj/P56EcpR9NokOAnbeyEYr05Jho+xzYW4pNFoj0U/DHAhabeW4xAHvM3+iRx
779rM7qWWoaGimfpElFPKdZwXWOjYLa1bJ9I4VRbaJC3TG0OAPZBv2M8hS0neg26
6HUHGgUvjqOU72ooFszaMwuDHtNwOFM51hj5oetjx/AGpUjiYKydzFJojJh7Akfw
DnMvFU/s4GI473CcLfzs5wEO6IHiAvKeQm1iucfVA/VlHxzuQk2pH4QXWJsj9qHd
jcRNHMasVKzGAQbHxEc5nE4aUBShfTG8vIFxDki2Tq31BbC5m5M0PW22h7VoCI/g
LSeRq8bGQsLJP5zTqEqj6Is/34ij2/oPqjXl95aMVMm33ZoJBeJt/ZVFt2Tm8ZQj
iD/UW29HgOAtigA69LR+sZhjbkj8BwEJPPyN5VnLpkXOKpyY/Y3lK7n1zq/YB0wF
xTVYezlS5ErmLqrQ8457HCVFjqcZ2TB6+07POidwPhr1xKkMTWeYDym/1RkpPLP4
X+2jk5emCn3IusjNiQk2aPo3wrn28G1LDqnfuySfV6GoauuehLgvnB55FPAuwEGa
z7ET2TYNpHtsLU7JMyo5Vk/AvfBwCFJRZY6Hl7AdrEuZjbumbKzYx2LaGCuB3H5e
U//y2KzDzGiO2TzGWZdzgUmMEzempc+gSHV9VCcK6e7ERqrjMR1PFUVH4zSft9rU
1bl3gfuIlx/V+EdRmFM97q5LvTuDKx7uArCe8ha0yNWjMwotWhX63f+TuTb0Ux6Z
GjvMqsBSH4wK8pA+BpNc+LpJdTrc+bt1TaFwk9nkAVjIytYT0UcF/WWCdKhWc2rQ
gEQSTL0GKcGm99E+wX9yB3kYxXr9nWciw7fByJVUZJmTsXo1FuEr+rgClJb/tN2p
KwA5OgChNFHoPmE9bj+aj2xh8aAW8EFOarw+YLghWXxicz9+Ouf6s4xIFafWoxba
d4GMc/t5Mdq9C0VumlmynICgJ0ntocvtAMNfGmBjOKX2q/zZIIEeZoN1DqB00ani
fZ0wG3sGPZjeb652Nhyg5dQji7TwCNAjMcHsd/K9oqHNCNIl41SU7dRudI9Q9VEa
/3Axap8VwN30p3rNspnfSuOqdxX21g/R3FwoBzswsW1rmXIHS6M5mwVtBj0RZzNK
e5ijh3cMm8n65Lvr436Ww/FFRvPDX+m/xRO9uGSo9EGCD2TnFPZDGyhD3twOqhfu
KgnWcKIhiA0BZBuXdYIf/DAGO8gU4n7akRZYI/sojnxiRGpm409Rb0HW8OD1HEKb
th7oswmx1cznFzI8PHvHM2i5ctw2YbVBOvI6tr6QMoPKZpplgomc0KG4taeTNsAA
eqf7CosBb/9KCWoy9f1/1GzffYfve3ApHV7h6Mn0hZ3skexS3Amw3qp4kOX2fuI+
cd3t/3Pv0CcvwvIQzsgck9hJbd+5TWwEAFWmJkc2O5aosdOGx/61U6P0yqMBNj9g
DVnqnGC1FZDtfKwDQdzNAjHjcp/DJcHjJ9fUUBS9v4M2sn2/3qoZI3BOXU21HSvm
eiMlBhXvxUMY9BHdazcC3vZjRFY2HsEZpd2ZUfJvX6riBZIgNsBdc9C5XhrNqQRM
rfvA8EcIdwbTYfic+0B4sg4RIQ+dLGFWy42Rnu4+r7h/6ODgxNh+5c9ipOZ1wMZu
vK/X7+nBEGpUoT1EXJKlUHkabnn4ZQ6pm4pcZuK6q9bYVrorrtR0Tv5dbIf6Hy+u
pOj/b/hYqvS2YnDP7g3ysYjxX7+DvE9iQZbjnjnBszSWueqNZpqQbHa9QC7EMQng
fSiQ7KhFmjWLBjd1r3pJgBDH39eMFdd2BIsigSK44dOjaJNDYVBJXJ0vgUpTopLW
z5cTLSMd19O6ZIT23qX13xoCA92iqZ2TZj5LFGasOrlP0h7DR7SRn7W6Ao3VYmfA
pPSU527B3TumAlCe6oELHvZT/ko5C86raIIBQBWvhwd4wpI3g3sZQm7FG7xyS61V
xBNAKrfH0VH3YamJgfHN8Vdd3WSQ9V6zeoworJmqU0hgf0pwi6mb6eGfrr6Eeo86
2VTTX0JINmuZfdgDgpdRMOk6WMUy5v6NwiYAhdV3y7eFIzf32KM1RYMk5O2GwHuJ
3G+Z2BzFgCzSYcGr7W1XjfkJJnJ0wfOaiVzY7LGKWduo2lQ4c3riYiomz7k2IAkr
nsmF2ibdqkLZQaryLuc5VhUSLZFkAuUBBp/n7dYm/JVh84HfP7uHqZtxWthT7ECD
OGJmaRnEufJ5DR1JPA6JIqCZZ7bQtQS87U7lf+bf+y6s+2rm5nPepn2fOmESBWf9
pkikGd+Ou/vVVSRLm28VqCfG12fC2y98VOXrI6wRtGuyoml+AWe6JigtI65f9gXP
8h2gnT18cI5jqPiTOLyH1GYcO5bkDycnZY+biJbrgfpJWK7yLmZNS8sQ3Sw2YyIM
09b5jIsGhaaI2M2N04G27XRbeVZ8P8hUm/BbN+3cpl0RtSFE3ssi2s9IH2X2BHox
BOX1/DpAS6NQpGfDSMqCB4jUK+ZFGILmwHqyTNX5ADu/dhPqOdmTx7PQxBMASSAA
ZdfuyIVhRB64ceHHQokowyULs3F33/hccMnkZtvJFvoIr8GqFYYKx+RTG88oXp7h
x7cLlGrofUsl5M7jUM7qHreEyiEkWSRCOK+WSuM4YLYdv/43+6lFEgGf5YRUCYWN
yBOgbcSVXhvDc+OHP2oFENKWyw1DMuBqwuGTSS0LTZXN4QpAPHe1x2kEWtrCEAIz
IBIT5rSK/Hiv5d037cl7AYwlQNNQkIyJJfDTJPKnIh+8nJx2v5qgGkFh9ZBucNuO
dpT0VPhDMA44ydk7Y9zgv5iUHaB0MZfdW6yW+IOma7tQJSla2XgvTHuzDMMg5SSZ
1VWIoaYCSU9eXsCm2xKp/rcr2M/YgsVYIdvikbyfjfX+JGW1O2GE3U8S5Jhb+fDV
SV2vZxWHAKTX1gO6YmeA2MuRv1TOcWXURnvKJX6IWuhASbh9TPuiR1IYigPHEW0b
vpaguJGSDA7Kt1uwQCy1TUbJ6ZuIQT1H11u5gDuE2bIQpSMeN+Y2OqMGEx3KWux5
ulHGmbWE4vua03HnD9pFlEs9zheZXGZH2f5WZwZotnjTUTpmKyn3vk5qmJCsQh/N
7QS9bFmcAMiNNLFNmEeDJ4RsE1kiTkgprMNvZkGVk7CeGXcL10e9RxcZQdXj4MfN
2eSSJnnU8qRZ2/IyY6G8d8evt9TYZ7Z7JE/BoVzG3eQ80YbtlFq5SVda9zQAwW/g
z11HqDcDMVg+33vNHFY8jec7U6FaYnoFGBhf+NWSd2BsiFY6kYro/y1J3/nIq04K
nONeZApgkgb59ZdUWyW9R6fr5EpxxhXjxMxWeMhs+d4T4IbwJURfj+C8um0t9s2G
JFFnhXoecergAXKBD6mScW0yTnTcLT+rdB6Lrnr0Zr77+8y8yEmIQsMbF84XFCc0
wtt5zsKevYQ2d+G9d2bbxC1X8OK4QNOVMqn2ql0BBqBzw235UCgpC1GitvUHdst0
OIkoTYFTk/H4yaCaTl8f1vErZ52FM0XDm0nmFewhPz0pAYRUnmkyElvcAQEa3B7d
Asfp86gtUH7V0zw3bA9Ro4u2IwvNDqt75sUHJEt9CsPbCexDriWGVg9Xbr3DVVFc
b7YVj7T8ayw7FZHVlmpsyc1vbm/bfjx5E4QlQ2ZdjdmIuq+M+qHLB30j9azTFL0X
zHYUuRP87hC8S+LqY0z0GN3+NCdaIeRg9Cb/StAvTD4nl3NjcwEltxj24Ik3z5yR
cdpmh8gd7GBzjV2K98hNUWOfkp/Nw707FmhvPAdeuHcoDFxBerG60aZCqo1f1Rm/
0aLGtxTGT0sqMqpqQiuScWkizaixuNqgvVk23sXJnMHDhuoYpQ7dLe1TUCO6so/r
YSnR40FPqibFHyFd9K/IJCNdSTuc24VcOsvDmijTjw1pdB5eVt57bQ/ujxkBOwra
lLLFMhoP8a7Ak5PqTqyMi8+bu3EUT24zyUqCvqZ9TDTaIhMKTUEC2KbGfdrPid5c
/7Vo8J1HyUoTaNHb7p12phtjjJk6ukY8sd/q5IFyyGXhFzOdEnVmn0drKVaqLF36
amECjI50Kva+IFR9Wd1+45eFHi1OJIN4zH37liV1di37u1u1QdcKS4aDkzPoeFzh
KmS6Bm6bEEt+3fC1O96X0tDWkZ66fHJs+8rWrP0M4kjgu2Qu4/nPcJaDd6fqNzd5
AaCQQ+f1HkFGcsn6LnVhFAQ7oj6w6MApDiH08S2imLk0wq52G/WFtHgY6IAjSjRp
lcMhBaZL/oJzzjMOG7nqWvJWqLl3zMHZH/AIrGIop/y1kzsAsPYAmjaKAZp5Ouia
cURFdJQT5PMVnH4+A8rxAKkg/JDyhtvsPpn8sThiuHYXmmrVAnSSCb0fCkHv4ZcC
bkt9OYuaOHR8e73UN+5qO/zz4cBl78Gnmag/j/1d4ByhcRBOrnzQiUy4O/X4XlNZ
bM7CvsSazUKK0+YWsegO53iZKQrQ5/MoGm2zeW42Zap1XsKAlTSoSwuPdArBHPSC
FKBRDsdjwebP+88kS8LzDIRJiCTaS1jPonTCeJmO06wH1YZxVj5Wfl2NbvThEosw
Q53j8BaquB7tLJyZ/OncdHvboRMx57E8njCKIoAKM7vSHY8SCinh4qa4xTAziwuC
xHF9EEoECoWdJGCuttexd+a/nurA8iGn74OYQcNeCMKES3AzMKSL3WWjsjmXpewp
To8cvn+0/6cvl41eS0Z+lQCdJ10S9cY86sLzDAq53YP1z8WKv2+rPhCgNcXTsmy+
bzIDQyZ1m+2UQNCbdERoRcsU887mVvpQmnA1IPTDHGw0Q92z+3YroReCW/p+KzEe
sX+JS9CpWl5XCCo5LbHD0mx6ISfiAe5mADBXTBgxOMAEFrOv0YxxhCVLY4PoTPEJ
q3nERI/dR/Mywwe+wdd+HZ2Kk73I4mLgQPe4jh4p/6a8A6+dMtZipBfN0PN3D030
dnC8jPb3cjbytFWcMDIitfllLa9I4eboafydfbGs8lOu9nxT2CDdIvs6lKG3bBZk
rYWgTftQCrTbpILnnBNvcKC6jBeVy7UYrfemSdL1VXkZh5MzcN4stWU78uY4lOjO
GgHYJNKn9kNPhKHTXcMdWT+CR8Cl3+e16eAi1KnqwQqUT1Rlhwd2KyhdpEuUybdM
PDPALQfxoV9OP6atBvKf/oriuB+b/T+7Os5jMazhteMVRr72vcPxvY+EbdYq7EGx
G3mpNzd0fAWjkdANuNg3cqEK8IhtL6ARGUqzzS6USwCbLD00o+r4sj0E6NvHohVE
SN2NbCL0DAf9ACifcb7xIQ+jA5p9nvSxYKdLUFEUzM5qdDRpyajuaNhJubj+UPOT
eSJdnx02pEYhWcFoTIhTsJtbJeZW1yzdrtp3cM63gVVqUhx+fFOMrI27QeghRUwU
NP27e05nsvglLg3udJKubkHWurdqe+RdKb/C95KwhXud0s+N++CFLYVTMH7Sn/tV
mqT7BLPThx0VoZruyGghkxCALcgMfk2HJMcGTluhp6yR3NjkrCLqBpXprtgwul5w
A2pofRGPz1U6PFXiJ/5+w077TkdtGWBWwIYsoIc6lfo=
`protect END_PROTECTED
