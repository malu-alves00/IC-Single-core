`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EF1qzd8xmKUjP/bYAD1fQ/crsmd+24JKYyu24v3j51KK9+PiDioaKgo8CXLRA61y
ax2v+egRG8UjAMAgQWDBQzqxiZkajvcxvmvg/Dj8VRCThNo/J44WRkEdhMh/utL4
w8cB3KpTueHxBnbpQcIHPr63DmMxnliVVK2lHkSU+81IT1aN8bxEyevUzzbK7R4g
M2FWr53FZaFaBvkNgavOQffYgdrTvNLZzBOsnS+ps4zW2JVviKBgNk662Cq5hbMI
nVyxslf5M4z8Dr/yJozcbRytAcp9LfM7IBqOiAAFboJw+23YRiItOczFwQUrFrdu
6ykhm2gK26j/cvDxWPtx4D5NwIebg1o67chqSELATWDFmQ3WMfpdMQAU+EYIWnFI
sQPceAI91Bpn1R85uSTPXucBmNPujQugwo6y7FwUB3sP73J69Qpc0Jsw4nPHvCyf
ZiYeGjeJ2RGcQGbbxzRmDIkuJNKWmb5BP/WJw5n1J+QXqKMzouwykbDVwskfHJm7
HNpQAQdglOLVPoVPkzQ1/PxEHsIVitzAf02D+5Np7Oc=
`protect END_PROTECTED
