`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CDn0S+ekRpDdgcetQXYTqKnN+6Tj5jfYCQb3Zg2P3fTgVUcoM032JemwFzh7N2Kq
StDYKmHnFexE7OeAoIWj5cl8dmWqFAlXFqjKyQdUU8aVLNDFy1hPyfbJI0uDuXz4
zUrNEldFAbTSjW188YX+Nn8lLtLKroK8f8HGfNbhrA2uCY5xxOiDyRMCwcQnYcO6
Yi9qJh0S05h5CHr7ZnfqgR/mf/3ODEYa2PND2LrrjMwIKiX5FN93SShln48T/UWA
PytpCfFxsUCwwRNELoMyl1bqDmVL/VnvwXWSR9xdvZHacdAC0A22/AYFN8tRE7S7
HW8dxoIu99yqdMUAoPxxHzyBvtSOWZDGplU+jmil40RpHluiPINyD5ISvVlq2Cmn
Dv/UEMNZB7rXZ8QIYRNJNtmOwKKm3ljYO5E+DAGCNPnThOmmJkjiabw73OLbRye5
9ozI6XJQvZyRrZr3f/vYE0FP5/Fd2YNAtJI9q/7CcrShE1oY/PMsCTWlJEe+yLI9
SfsPMYZLaYYWt/ySpE8pWJtwqFFr/75UAO+qM/e81N8CNoXOY/9iNBix7GVjkPVq
`protect END_PROTECTED
