`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fj/gKhozhl+oWuEW1K/QSI4iW7AYw2VMHiy6SooKi0jqzF93onznsmVAGYGz8NEY
3Sdu5CR12khv3xNPysaM93c8EInke/mP9J0lqf8G/5S+59Z1kc8hJggNhJTK/Os7
3n6krZ/+//i9f7Okc5pIdzP5WaKGnEmPa1R4btgFLcVtywUkhM4Srgfj5CngRtXB
4Q0mxTCK06wCNt8XwglNdE+7IFeWzHD2QPGrRS3KFvPWq3hCsgxut/8g2wKfjx2V
KpsebkYShs+6iSKpFMU7HTWMbNPaJkcv9Pgr16T0uCUe+rAnTr+X1Et8WgaU7bvQ
teK360cxIDT0Usbk/dCgXVWZrNpqP1UXrpDUeM2lDIMIzuYDy88OCGVIqQ9a7VUw
cvM4zWvi7kwr3a42xrwEGK8ePN04xy5F94TnVX6rPj6trsDagHwGBcfIK6AfKfso
xqbGYny+9tDpI0h+D9ZkyygqNZrhB+q6jJHni2PdycQ+9ikIKTxxR6QDAU22ntF/
AcFRwySSjbnaw3gP0wFK4Fdh3EDpPEbeti7lrVum+913yOWG/FWINUVVSWWWDqqx
6vUiILPc9RDYn8SNeiF+V68bPMY0UkLbrpmk87mIJn8D4R3hFYRZARXqZrYdPqV9
mCbGK6EbHlIuA7nEEbXrmzIPn+WGwFr9GVjJ67u4TdHbYgKVkLAYupQzsy4eO0jF
dANcBEsq5TTTJANbYGpLFX6NTq46MKU1ytCHOg3G9pb00hkupbFjwyFlbTyuQFhK
fORRI/4/4II0sVfhlUoUbhuZxJhOTSx0oum0h5tSY3BMb20UQ9uAc5pSfyVwsl83
vK6Q4h/HD67gQ5aUJXPes0ffOJtVscFXom1AO1yKxEB8F8wUaUkFysF5ZyxYCEMT
/fgE5nVqx+fLXTpLyW06Gm19W7tL1bEeV9vwq4+5i7ccC+onbDTL+sCFWdrhDZHB
/4myfeR3Hm0JkXmiY+uBCztTsmvcwiA+1l6kvaTKKN3z0S0ZFHtRK1DjDZX35G0K
AdQkXmxk/uH4KbTqUvwiT5+jnoKkW+v4kEatIKrNVvygV5ymD86+YNh9ekoDV2/7
EzUZdYzPmSk6ku4uiuzahJOvR0Ehfalw+hp20C9TboZhwF4LNojpLDvNo+SNNui0
BvLz6kfLajGjj2j0SWwtLL3PmjDS1agAihd2XEJB45xhE3ljaW7p0oWpZ5RNvppQ
4MDB50/f7H9DkSDW0HMCm8Xyott8m+O2g+Vbu9uNBkEhV5+jh817F+K9Ndotp1K0
3yOseuQFU9OQRVXmD1OLYZKNa7zHwcosRa13+KnDbWRp5E8eAitHJePzkuKLJtw9
bYkRmMqm2lIXXHSNYQZ+3ii/4QvMh83sY7iKVBsD4G5Qq1dQoKwHuqpCrtef27JS
FabuG/rvrhkXLcFuYp7v29emNWtB+H7i79Pxq0kS+YoxTWU5ZwREJ0tsKqfWBpwz
rO8zk434do1zTy7+hfGvPBUz2hiBWjT9HzFxyF1S9al5B0ZU9wYepvXoYRY2sO4G
1M3gtbMDyBzVMHEFsvGoCN+5APoL91HIwFa8EsD4R9POZL6gy7wefPhchjmcX6fV
4Fb/ZT4vcUn5RvjI98l/H55jV3AFX2ivrIl613Ft3VKCrPHMLvHZYGk4Yv7gx+VP
bku7jvoD5tINAUX4CVCN/rU7xTy2V8HDdFd5ZzuUFeiTQL4mDldnKJ2pcJEsx0tW
0gTk30nL4eKo+IJczDVOUo0HmSNLFIXosu7XtcsgC40sQlpAp4TgaSzMQCHUuaVv
oXLMctMcaysdYOmERDbFSHLPXPJKnOk5qPn2JHAB1ZWyQSRjAEdiblP+RRFEWUBf
8KN2iSUb6pj8ijKZNMzH/vp2WLm1z+PHb9GPKexaMZy7FmRQAGDtWmbatW26HoM/
d/3rqTnEHQSxIlGrl2pV96argXntOStWUzvCchk74dN0v/18DpyEHJg2D0FBwV4Y
hfFy/1xZuog1AhBsylNirDsqficR6BOrXuWtIx7xk7MHWG399zfABSPw0emEP+/w
TKmYXmFL9DQzRJGFMKcHragR/Bq+l0tUC7I//W3MVT9780XcgRg0Ia8UiYXl1k9b
lzKpna3Cy8CVpvi0yBX2M5Ea0wnNTFk9MfSMx/1MhG+57gT0RKDnVoGP2rdr+yIN
7s3qFD0W4xJxVHLTwNkIm0R5hgqOaKcXlCMLooNlspJ1uCiaWQAqu4tEMwwuro7g
kMKlV7Ls3YI9njJI/T1NUrhfJtDDIYsH2vHzfzAfzgpREedSW3IIMTseYwTwNsgR
uknNys81xlCtBL864PSpql+2VPh8gPdwVsHokWHUR9KG3fwYgGMjI2gggCn/N5um
/5c1yQzPiywv7TF20FPAU5sLsPlJXzdw7gU3f4NGAFGA75SDn8GH9h7Q2Lx1yA3x
OmpPljNgjweDzf8yJ4PUJk9d+eD/UYiQ69DpH1PxYigyQFfcTwoUE4qq4x9qNqE1
ztCcdslpujoF0of6TbkAh5ewVpONNVj4MffyhBsdPWJ0bPYfXvATbVypfafKy75B
30FvdIB+TxWtAVbH+Nor3k3WMVldTthvbdxBPm9HxirGeT714pebPXnFDh/FLF3z
AspPlRHxVxcRUUWaR6r2/bvrR3LL6Ttm93koTPj1IENk5XbStyUcxUYPXxFwiSXk
XrN5F1mA/X1aKdsxLzF56y7ZSEJayLnqmnq33Ht488UVPdLMstudBktcvNAaOQCz
2aaTNMZrHAUO/z9bj/7BjNfrdNVgUxF2bEg/IoeO7CRehkp3ByvWpP+SwytJxhLB
y5e5EbYSfSJiTu+qLK1MNo4QYaqPIG+4axNPsa/udrE6oO4oI3Jdt1gcP1XW1ggx
aIeD6UzLyDreNKCDpYP2PGNzOciKuFD4Kxnix1me05pVc4mcDda7uZRBz6ddMGbH
uFEU/6d90bCvcZzdCqr4Bb4RSMUGRTVZUIV96NO3fHLQK1ppZPApU4IzPPXquSFZ
ApQyBbiG96oEDTml8gEmS8rMKRaNZeDY70etjPwRIhneBznbRa04g7MhzJgvheeK
f61OeUjBO1hcObCp6HFqbBEq9qatsiItcXZMPX3L7f7NZoUuO7/0lPUZ5vs1WIuR
yarmErIjAjLsOcsHBNIAHGH6gK0amceJ9c8dJ9ofE80V9dMxcP8A3b897dMvEDUb
xmV/FPRiGFmrXmSKTOxSoOfMXUo/q+mZgufdXbTVHfeMwJgoXDg+0jMLaiadHMHu
6K30QSgjyXhEUz202dqzlEc09ketxOG3jRKVpXwROR3nwNQHXpt4SOea4sFdxS7W
EweU3UsKCuHzZaG10fRqOduJs6rOljLCO0EV4VSDkXbcZ0RnYZ/ERaZBFc4OTI5Y
Bhr4rsCH9uEW5ZZ9x7YlD0Y2oNfqVTLYtMylJA3WYZRmvZEtWtVxqF5xfPiRLja6
/vp5CqY2QJhMYt2go0p7CwB3AT8Ns0+X/IM0fVlX3lIA02dfkNb2xfjAG7jTMNm2
Y8djZfmkL3+a0Y6Zz7Ghl8tvHWx5MdUxlutu3Gqf5qOsaU+1BuXqooQ++l6WAG3S
NQz0kMlfHfHJBbRrxpOjOG89rYwZ5QnjvHGD09R7dlD5bZDGT2+WTCMxeIqPUBFg
p0w+ue0LPXAcUARs/2onSzrlvj+60g1Oc1vwAlKDJ91ZB/4kdd4xqi8i0ogDPY1L
VPGtStP45PhBuXh2SuuoYvs6m87z4GfYH4TivUNaVUVF1Zh1VV3M236nzO0st1cB
ABK+gtdf/jhSG5df24gcy1MrCPyfiXKrP2N416/kaeK/zGz1cGg/YzUhiWehGFRX
5hbaxxg3oh0j6DO5qdIwGKnJAgzgPAzUmjFT1hnTzrvlh4IN0QHqFndBKHGGRSZQ
istdNFS4skuEJwgYwGn8o2CPD+Qxxm32GRA6cfXG4m0ADGZeWqLAges14iMBFBXB
55TP6jkVYsbthSp+TfyWAz9eWkpsx9Jr1rtwzD42fYVgZx++Eol+Lw7Wyq1JI56k
TEyPEav4q+3HuvjJAw21JU64ufqgaU8pUUSA+f3ZTqecxFyLgqqVOStGPs/Ll3ds
xffQVlghXf46Vx4kVpRElyBRvqXTwuOi6ZJGn5NJj30N0UaLayW1/BZaufVzUd6L
o0GgJQY4oiqwoJMXVYfkd0T/HhmDhqWXw/sBc5oTI52pxhiHb52wZOZi9GJGaHh/
p7TRbAL746W61WStgsF65CeTP76dWdrCwhj1SO8Pi5kx6ZB/bQBkZ042tERr9FKi
z/s3t2mRESJK+zwQuR0gskqjFjxYAaPIP9NJ4cQIAPSLq7UFG7kg2yJgiNvfuUYM
VasG+tOQ67F3eNmRTviQqa2I4ChgT8/QJ3TbQny0POpH6PAdYmqi3O62HXkKBAXr
SS3O9bBfwppC4RU2oQH3ig6+moc/OcN4SanW9niIO1YanXdgyeDEGGyR+RGupx4p
diX6BtvElgwdRijDeSV8JrEotW9S4e2/Ad39Vjl7bWAPGlaFr4yxRW0kgE3OUUSR
07KpMMowO5OC5LqZ5/bGHNv/OVQC0zxG1XZC9A36KtTIGm7CqfBz/Ti34aWEOCeK
R7JK4ajiuKRccFl2GVNPOiO5kIZgVSAOLAo+YFBWWpDcK9eZ72L4aMy5nH4GvDW9
AndIDMiGhG2YA9EE7OWghRwdRbm1yqd3sSQhLxh+H7maGtYaDhsagw94r5Gsl0Bd
SRqLCGIDLqehEEJCKpsdH6zZrOL7rb8bctuKIw3O3iYI/HQC0iNxwZ7jLCgFsKkU
KaaQNVtaMMsfS2SnkKEsTQlt0FRw5ZzytaidcpKgbtUCqzLqD8UJ5+gAYuJuxCAc
LSAYaLQZUThzc+VjflNPjcdxJVlnDYC3Y4FWtsqEj6Ez+RlL8L4asHR0G1l1KOyh
vNL/8sFNsJehP33rlF7+5aL3EB/GrFbRA/92ygECxG7A7kMZ7xsXuy5nWJvzljPr
EL+U7sBiokEXae0lOtiD4X6p7+N67fkYJ5Y5YMM6TxCWQqZdsrsDeLVa+bj7iHKx
CMOhWTrOQnw4c9vWwea1459pDNHT9AqGhrLa6AVgdrihZFeb+EMpwKOlLJuOlZYm
tI00qheQUwx7gwnwHTkIYwvQkDqwYqPcNOqNL7j34jMAWy4T72suQ6am+FrTC+jL
M7vfUTBdfncCCbKJTUtkBk8WbtEWn7nQE6zlPl5LdijXIH3sPciV9bp2weFONA7z
osqkZezWjaFznwVgn8JXqdx7zm3p+LgQnTi9dXa3ielnKnzKHhS0irlolbf4Y8ST
40Pe1CU5PmSX7OAgpPvpibm7VHmJxylpoHSjtSRyGgCpDXVVp/UAa9gPB3ak7PqS
vAq6PuLQzpgHECMjSSIZ/F5TpqlXtgZP1mjFkMMfnZuL4f09Er3T1QJrTu6o0WIR
yJRijislJ/fOE7srZLZsSrdDQfGhLU+LHcTaWmP801tLm0W3BG+4V2s9GjEqnV4a
pfWkjYpAnUFgMCbKSDi+5wKKWB5e559hpSa68tyylKCvx3HuyvqvVP7joWXgE4iM
L5yTPacRus+zwswJ87HKkYcN25mNPJoNmEu2+xffdyWelP2l9oXn/vlfGzAByWHP
Xud6bHkmea47AflPKAMhjwVO93tBhFHek1ocJgJZO3PaZeC3QtSgNfn+z4Ce0nk+
Gy47FmP05B0tBKQzo4UYefjECL9SjBGaXdwNhLfz7pForZjuz0GX/l/gtbGUqJLU
ATsOk7RAeTxwmKz8/+EXoMkFtAT3nJENZRYOh1GVjhBJkckj3eCvY7ScouGPg1z0
UrOMW1YqQZ6Wo5jcrZyKZIGm4T+EdSYxwfxpvk2bAwAIMN5Vs7VaggoNzB3ghIJT
IIr8L/oNIcGpEusI46KqHkDa5ZlDPdCsuxIHwHQPeKTO124P6q15rdvfFy7PU2c+
YB73xY30+8Ee2ita+uNfs5qeYeGwbn75uXl2aMgvp5R5NtixTrIA30/Q4KjhFlDa
eTy2D0P4qTtK2d4siISedagt7QCyeGdBe1qPnY3eMGTnBiHfzP9HlrkNId92xQlF
FG6wC/O4laW42FksHtQZBL/MRXMbXN3EIOXEaT9AyoTdfgXYHXLNilIk1fYr771i
VdkmiOoY4Ov8CLno7OnYpxn4whlDqc0TuVzatsItx5qXiO+sViu1fk5F1G6FijKT
JfoDsTCQb/GnVkPSJ2rDKWhwenpkoHnrMZK/in5xv6PFOhmL841OjVqfUBglCgmN
mEyhMAS2lVFWSpkhm7b9Wm31TWVmNGOrD2TC0BBLIbmxeEHxDfk2Gjulgu/6JuK/
4pCgPsKdNYiPJFIBP4F7tq3rdtwoXXISpXLcZx1BZ3A4PCLYaRKtKgyCyp8QcTya
m3/iB4ajLuOHEdcYJTbpVnCDd5+0R4oHyqJETMP7k9W+sANbdzo+yrqnZguijf5B
Ec19dK3UOEP/BZMfpHjHQuvaA8CsIB5JF4YQmIDD3XrP+g7/ubhm0GA6swpildM6
b0Wxid0EKVkP4FmR8qimgkB4ti+DZJh89SD58rwwD0apu1BZ4cgi0x/nlDTyJJ0g
FYbEOx6Bx7Mgfi9AcrqUJuvOjOXMDjG1RzRlm5iQ7Q+FNQa5SRnINGFQhc4dgjI+
gJJzIhu+Kv57O5iU9KXfZvWf/yCsycNWvyldjxShfL9ISCscPydPBV1ot+kTbwIw
GIvU0UMy7BUhJjwsyrJA3l4dlNl2PRhRgcqVCyqlY2SEV8wXNhVqy0PxmZo1x+aN
fwKx0m57Ld49rQ6xFm55vawcDjxzgE3ZZrqPtCzyp+8LDExhGq/I0oH5o02h3zdw
/dKQIJj6uf8kFH97M/PV4Zo8/xD1TuO+9F+jpRl1ch67CLelPezDhR7fCNcsm4y8
Q3BtSxjMmL7cEcLOBJaQ2b4Bp5lBdKlj41/mzNzvbJ14RfRMYWg2KMXOVw5Ghh4f
k2oodvjn6I5k4a2iV9DRedOA3oU/LOBxwuOhavISHiifM0aBKipQ//3x8nlScTNJ
MUTyaKwsX0/1cXMeRqkUpzFDDQAH76raYtHPf3c1Qqpc+TUUEXheBwecpftwH+P6
rzXqRZShThvuhisIWHcA96qdR6k+/BWlDPdTJNZDZ9GGc9WcnUGbzphikLGwi1Jk
fNtoC8Tm3w0rCKogJQwACyHFrmOajvwTgZLICC0fh20PqGyIUKOdoH1NGP7wyFLL
KoLhBSCkfCn+9023Ek2fGxj3hua38fRcXNtmrMwBCeQHxz4Is22+MVfKTHDYgzGB
rwCksBctQ6r/ya/9VYoMTi+gj7DanP4+i/cARDZ/ZXoTBJZ816QU6uk1eURhvAb0
iG+E4DwGT/UirHEeP09+9m/3jMOoXhRvGhkwE7TgHSR5is2SQaRYpdXQ2htO/3Sb
luMYM/0oVK8zb++eeAITWk29wSZwUzwXrkclYum/Xfgb5b9Z38Xz5kMM531NGZ49
wgAwnkBE++uuqLJCBkoIi641XlCRKWBxEA4i5PzjGXJP+pKjFRXqWnX+MLrtOW7j
xQtTGrPrYonCVM4TBPsGBsIc93fY/jPvOY/TWtc89MK7Mtl6Jfu32EylysczgO86
ZxBUeBvxy3OYNaYWugwLnIQ39sYq3jFJfe83z2hvfxvcdMXAwIZ6I9oa/nKma+k1
CD29gXAgg4+YidctUi+l2NHAk8BrcL/iL1CyySjabVk24xQxVhczL4+VBaUhdhRB
EfHpy5zV83WjT6lEwwel70qUu0ZfmsKuSlN1bKG6nMHWW7dYx6+ij+FMwbmd91JX
p2nfcL2n7vdsSalaEthCzrGyk4ZnluHHr3ZEMzeXo8xbgmweaL1sHSg/bkJjKG4E
v6Qpig06SAQ8QpvnzBsduF6Y0K8OkgfZoUuNAS9DutL/t4pvnyNpkl5FCqKCjj7s
02XsO4TAa8CGAx4luklM7zheU+WzDnLdXH6jO3kiZ+R7umqSb8HGZMn7r2mbNqpT
BlgJTQ1B2o3Vb3N3M1RyVc/hsy4rD8prQMA4fi/QXgt+biK02JIhhHVOpLMv2twZ
fIWYopOcflvQ9TsQrg7/R8UvA9meJZ5/vTLsXUadkpdBRPcrDOpr+29pfrddfI+n
UZ4w/cFN/Sp2heSQUMk0YoB8z25M+fGsGbf2ava4JpFT22oUPX3VbMopxnwg84+o
mwQ59zwRILZjMlhI+UV5yXhFum+c9IwJjJgNtxOUhYUtuHUf8rvfOFbM2CHHNte7
HO4t8CyHfOmvmAGXLu3bTikg8Ru4TGujTjIN9Dg5T4pbzd/rgBngwqHjQfD8rQLi
jbbIYiY/yrzpWvvF46dMCsg2mEx7e60vYy1avljHknIagXXZkuuhtp+wW5HoiaWY
yOX3dAdIpe84v6DU0raRN1aTqxVIukhPsCAmRrkcwthBdbDHjBBfuOJhZUsQgcvn
WR6Gqdn2OBq0MdaE0omQGvegfRGBniKq1FmxqzRG77Vwt7HnSr6Sl6HRom3VrGxb
dtj5g8B4fuyAyU0m0po7AUSWtoCs786DNGhveBQZ0PDrw9ylYBgU51QwfWmFyzsp
kWX2ooeN+Bfn1l1/QHdrIkQttwpODOGBBS+HnGumfFXVR+yI/gkOjBogaRyLdvcW
DncSUsQZRKJfmI0DogDqK1QXRftehXuGO3hFZ0h4eVY1dG9cbZRbzP+9cXfDCBxh
mjmH/+ZWNDu2y0HBkqcDJW90RQcLFaFGmj++9Bv5oTJJ4WgeYGjki9kTwZZp42kM
/vAgXFgvhOk0CQiIeFpjV1gFuUz8TOJN01qUXKYyRYxbJgFK5taa1qMaGtlPl+KG
uxFfn4a2NfavCtVoQl9ZJ92haxX87PVPsU0iminGsIhm4+24ROgkiEr47QjKViNl
/gMFfHWDrxNuu56fdMgClhs+z/5FPRK+6P7VJvNiqe5kAgKKq77W0sMwN6l83LT+
a+GlDgl1QqSf7W6aVEgcmLmbqS4z3AO0MoWcyZrwxdLeL+LUsvOWUUwUft7lUyHu
zeeyyKXefsgq83KCaJFEo4s2XYDDxusRYQniNX0QPZ2awCvWZWEOojWsnB7hapHO
Uvh3SptDztElxNb4u3xJLUajDr+4QDa5vz/GhK6ay6Vk2i5of7Rla5+fV4qt2uBu
iEC9FPaRnPy0JjqMHWVIA1tX6KVJc2H0QnqtLCLFGD01oNc6jp+LWsO0mln7l5z5
s4FhkMFthkV7cEsi7CwLlIwb6DyeQYpfdyPH9XroQYGyMVh8GLErO7KPEy4zKKJs
N90PRbtPnjSia8G4ISTyL00SV/RC7yaf6OQQEGeKW8qR3bARRdwVQI4XEOsRrT4K
DOcSFLCqIVjr514BKgkbkF8RCFf2NVAs/O6mQZWymblJQ/t/d5UtVVZrbPVCQIBC
mN/0cTXnhMcPT4Roukeyw4GHw7TKPuc5JpgJfRUY4KNLZT6OEN2gaGDH2iMhsA0+
YzzByS9fhviu8rGuQv6JtAaJHfF6tsFlnPpTuunWCP/Lt1PURhRrj2N4kjLBnYTW
7catee5ZX6uMMY9PdgS23OInNhmhlKBjoUIaiUsbU4CZQjrH6vAxLY4sgL86F9hl
RfZky4G3jFbzgTyqf5xTVi2iQ9rDlX+2raNN7UM2GSlLUOUwVXaDDh6FsnBgnO2+
spF9VguH4s6DRCbXpxExMUmSGG8T/l+ZA47nto3taTm1sWHbpMVkE4Afm/IKF6gO
1dvQI/vo8XgdDeDl1zFyIap90ln0lWqyDJ/OO3ef/cfu9TubrPcuY8P7LxfQ2YNC
ZHvc5F4ligdxqMAdd02YUrcMQ3moWhYDOS9itk9wv+8OX3ceO5ZiKA08+dTk8rME
PnKG01UWknXvNVdKUxuWFDrf6/zFPM5qpl57icFlCLlo/5HHPEue3zZPIPMBmPkS
GxhjcQY3TG5+q7Ww+0UwqVP5kXVsLX9O9RA4V0fVAnFbri3tRngav+M6ciZZfEad
aZgL608WEvpGqdHW9durZnSG+2uf4T/8RnOy5ABDHicai6Y6wTg0MTyLAiAg7NKD
OhNOvbubVg6LcjaFKhoCCirt7yeQbIKab5HrxYCRJo0stKM2kjRbLObwFc4AwY+V
UBdsZNjoXvdItzXLk/XX3+MyulGFmpx4sppBKqDfj8J5uDP3bsjDvg5XTWk3pVdo
9IQRvKL+CTlx11kGN2kXtIoov1aMnNWwWYUzItVJAOcTWPy/Jq9r2onxN33S01PA
yiCcPbbFLebMitcYuNpxH40N8kyBhGBeajgCd9GfoioAqzGQ+67L/Zr0f6apTo0C
PS5eGB2/VghhXZ+4Xpm8rlZOTkvO5Iqyfdka71ZqwhHBlIhw6AUVeLHCm4Uo2/Wf
UflJ7NawDCRIctNLm8f1WKMcfK5F5xs4XqsUudivnUaGV+d/yXdfnHQQnA7mvJ/4
l0+QD3R01khCn6p49zjs/CWUplHGc5dgg9yR3Wmk0+eHybTH1MWnzVlby1M2BG7K
/RXYhQB0CngQWkLFoTcwRTlsYg6E7B5iG8wZjQnliCfakjGreSeKpmongcfg4XW1
JoycGhSW531Yuh4g/A0XYAa1MrfE1vo3mO1dilnfYVYLONEW4JApm60BdlPJI0PA
bLjjl6ZNLhiTwlBpqfYZMvrn9/3QooLVaKDGA2lA7bi0bhG+Gk7MTv0lLko172VM
oSkZn6HB+AgvRUZQidU6QQ+81kvZ+XfsRRae0F12g7SdsIJ0jHaldu5y0g45sLxH
L1ADSOMhXVYfNoNyhzYOCHMbJJV7Wlj5BgK8db8B571l+K8sHr72v/e/gtMFY5CL
z8HfO8k/3tP6K0DQsfzs9LsMOxrXhr1mxf4EECnBHYTmXrb6Q7a5H80nJcvrhN/V
qxpoKS1oAnm2ZZE8ree9Aev2ca9AI5BEnG0VNR7CS0keVGRe+PlwYDFiRP4Vffk4
ZbxhQb+oJjuRYXCUARqXd4iQzJP/K9pEj+PcXgmOHQMNK5ZpFBZp2eDJHjLnmCIx
/iIWapAUcIK0UxkOlfgYmSRudE9zjsQO3s1yuMxxvkEJ+6Ey5xj/jbdXi4bvXk8C
8H/HFTO9jGALpQJRScspjZtwhjwbaU7oj+SmEu/+6sAG03iAMFY4JBMRhSK7094r
9XcUv3xZXHeyKwXZGjRAK2n5A4DLQ+z2dCq8kSGvAQvABeJ4plrk29smWaUsKCE/
axv4XnMtNPHJSHZVXW0htJme45X0u38peIUN+3gCz1wxgu2m96iLP04c018v0zrN
lL5ZnrMuGiJzT15Az/lJdRIvIU0xi0orhRr1oaxCGH8Carm2A1GQCaa+D9cX8qaT
d6vVKyMFcyq2XnkJs3mruRuVr86YVt2wO87Rrwv0CwvtSGWhlnR9+FiU0Ph7s6LJ
dGmSFa7s4gGWgi29Jki0HuGJ5wGKbIm5xqsMPPUpmcw3jS0KGjEhnJs/pr1I/Ps9
ZHlOFAjqh11iwWrQbmEdkzzrj9utn6Im/G6LjIN2qhSuOLKeK1HqDj9q9k9AGTpX
bV7flBpQLv3iatgn+DRofIHOw2/aIs1oqVBdom4UH/Sgv+Fg7HE3CtSgOqbeCR74
i95M5x1coGpliFq9W/m0ElSHDoq1PPEYUEKgEpbjOIGCOhJZuY6qPHlz6XCl/tk7
Jn+AM0juA+tWQdMi3VmOO+fF4tCX53pwH1tEwctTEX55wP8gc1p5iw65blFYz/rq
Fl4q196wdQMa5XveQOoR19vnHxEYCAOcxtRXEajznkgXtozk9O+E4vjxByFXV3ML
ISwWqJrPvjB6nkTcMDUh6s9QexTK9sivcWbS3l2KKGYxUWYlmHNgqLQ19ui7uR8K
87U5AyFfZt8qwoSpyxshGKPs3FzLYfukrxTlnmSlAsUrgw2en+jwHMAIpb8uQW/C
bnwNzQC3OWA3K443wmpCcq2eo0BI2OlFHdcGxoqooPFDvga92LpqyHL2TimAadC4
TE9gOViBoKNr4QP5n1bOCfBfZoNxKZ1O5E1a+gvHww1srILz+WrLrXgHLcnl9L6p
sZexNBYCy3WZZ6mubUvT2sqqSHYkiti+6xQBW3/DBIVy1eMx8FIi2S7tWQ2VjQhg
H7vb6wP9jHsjJGbO+7km44vG6hfF3pcRKoF6XBn2gUi8hMoEVFfAmkGVEleGKZUk
wQo3KeCYlwz8dYsxPKHX9pDyd5mToXpiH2FLhhUzNkumcU0JUSKbM+iUTcv2m0Hn
lhj3qEi1W4Xm6gzv6QMPyZDNrkk6ti10INtFtWgpqvjFsauLrSDjQgqf5wc79S0H
foS1ujeSwFP9/977bb0cyk0ZCu9PHS0RsD8gsasuuk6PZI75Ipb1/h6p7yZSfMEz
rpphhTc262HwnBKqMrhtYAgNOi+26+jweOmdG/wS2Mhwm6Hc5Pxlkw3wW3/GkKz5
uIc39xwOSiESRgMJVsQOJfjupuw3hMNarlXvyPXslHFvDh26y1MohILYpBogJZQV
c7iigW6QrC//jtm9tGYO51hjsMSlGR2dTno8kpTlyVcWDy+D96aM4es/2o4+/GPH
kmNW3e/VsJJuQoEp5q1y4xjZivrmmu8SGesf+HnFk2hVg0i8d12YLZfgUyzdVWNa
EFTDIC6HMgWD2XClmsVBCjFIgJYBQIzGR0Tf7MCeMk2PDAhGWk809qz3qVnpWVvV
DfyKTGGCBkH+IhFylCFbN6LG8K8VP7DBynaGKCdaX3E5gA4+V6+OJXiCTwwheopf
oj11V/FYXKyefZc9zJUt96wKTY77m4L/UQz3I14ecg2HweqYlH5JJZ1YWZyogr1r
8KAnJeVU516dsOxrXe4ATOqPN9zPR9rHOvnHa589n20WvuVurCs4Ru8vdwV3E9Dz
g07qiPcO8SEkB3zlN8K/+B2ZxuPUmQ12eeAUwXQ0N2VuI+A564M2SQc3P25RIg3T
tmxarxe7jsNU93R3AVZ/owi3C5LfCqt5spkIeiOQmdZbWBA4raznCOhRxNwWVv4a
DqDI35C/bC3wocjpd1Rj0PD5vFReLB6oCD/61re5OmgO+Ll35M4zH5bwl4n1ofDm
cagkD8mTzs41EhlMsOOEpvWHWvf0gpAGGeGtasdaEbHq0JaikYbUeAKCr+X4BMIv
NjoQfGDqcdgNTqWCrMUVuL34/ytYM0YYje2VPpSIWuxGayAsomMySW8n8Lm/ag+F
T/XaOvgQCwy52kRiTkswy5qSu5naYaxG0vv1lXTXVXMqsHF6RTDTZpSUck3+lA82
jNp7hDIC758D4KWZVho1DiTUAODPWcUfOOYwq13eddti6zqIP7RgcjQDpN+Hhowa
CW/c6xt7l4i5VRxACrszQplNb14k90LXSxjKZrleeO/TB/I11uny1m1CdS9hIY4O
Y1zFfeqYzosHSKOdoJR6uH4yMKfljxRq5I6ww9YWCbD+Mfkt686ZdTIfOyySacO9
B7fWgd2r7hvDcvgWrE3rzfwtGxa0/MRlWZFJlRajO460yU0enQK9tMbiKsibfUVf
IeWe3DeUpoXmiG4OrIlafFGDpIL/uWaGJ8tramPJ4syqkLN9ON4329Wub7PoFpP9
Zb9lyiTbdin6NxOsLY/N8iMXmudB//MVvOeQBodQaT9hU5cxF82JkAPnkhJF85FJ
Jqnz1m+nLv/1REmq5OddVnyQ0Q7uHU3+MuuBsfhxOohKg1riU++v2G3cnffJ0SyF
yrYuPESJBm5I6OWmQ1BgO8jo1LYORrJw//W0xKCNWTWnvPbfGexPoi7mdio+E/hs
SEgKI1KrSVU/PcAziJXfpUFfyQf6fC8ZPp8c62qJsL3dm/1yt52rLtB1pTaR098O
vk/Ed8atQfLrxr6FbK+dRVFDZioqerxpDlr4kzHEyAunfEl+4kKuS4fnMwqcrI/W
O9x7xPgYF5g7BRD0BCzj74lNmk6PqVS6r2arV6gWK8FPxpK6IVd0RE6boEhLQrQl
9/ceS7lkQ8loYXrPMdfRvUnRUuV7GWMTr1/4F0kwgHy6b1YfcVB3+EKPkBaWnStX
78u9uZNPRo1mEFOIC1NoZDWZ43RWfexL2bvEDYFnJXk0BPhLp5c3N4MJSWzzap7k
Wa5r1YNkTBrxRimG1RkUIy1SxMKrHEqxO7jqo03vp155+2dmB8O4rmiEaQQRN4z2
LKPIyX3VDsnSn036P/3blNHyOTdVK9GBIxVahLIQxA9r6djgpxcQYQ5+MUrrp2E5
n7Rw0xgrWfzKtQ5adt5K0VPQZtcsnQ22r/1bTnybM79ERDzlp/6BTmVnxdxDth4d
KPc/hC1d7r0br9x4o9NLcEIIEr0pg6DsgNcskB8gStbO4jDaEeFsm2Ly1XppCD5R
J2XLl6aV3lnEpZ8EWtsz6WRrhoXdVmANHqlQG4tQde6X+wskpkJnzf/hYtsCP/Uw
cOikGp/SGwp05oXbN1CejoE4vN3wGpNCEAA7F9Rll4Emn4VfSDcPcab/VK4gnxZp
DvVwerejcC5LBjSHiKjHx5DJ0uvwUFVYnUYZ4OQFgVbns60Hl2E29r+etqLANUFc
vm7od3CCI10SqC2kbSUrXyUts4TMT6XxumZGEAuHLjXe0NAj3qULIbSTKX3gDvOk
fDeQG6g2LvkDgeQG3Kl92RWFhJt9cd+oZ2Wz1A8MRn0hxtZN/stg+7MPqUtWaWMT
6mRuuyTdh6aLJa3j764hwTFh051UdtKLSwN1YG21tU841F1HH+wqsoHx/BL7qQ13
uOE0kQ+o3y//QweE6b1zouDKIF2YX/q8YtKW8tkayrieWHxMjifBz7Wt/KVIH2yV
xULZH0AkuWcfaSYyPa7HdMF3fCBc6JZHyCBG0htSdb0HXj4t7pxnNQv4YltFBX/b
unlK+5IR1LJzjFVJ1lzzLatB6BQLMQvcyTgHwlZSwCenZXqw0MMaTZ9rc0O6iCSH
Y97ZWfMS7T1YjvKciuoLhNKL9QI3O1az8Maa2ZlMJVAPBMrZq3MHDho0pQ4bcDo+
DYlbr6odXHG4XMsEjWKjIjJGh1IdVYat7IVJWaUaJi8B9S/RmR6Qp87zNAtKnzia
f0W2yTlYa1ukJD+kPqzf6/Hc20NqJ43XihiA0HIrqDfxScZijYMg/2MJR7Tf6eoN
qdY7jlGWx2mA16+8kKSQAEDvIJfsCG8HOGwEGG45WWc35sMxi8O3LNeVTVvGtQhp
trIDweEPfWqXzwNeT5D0VcnPfGHnn9z1YB/GT8M5fJFPEv678mMlhz5T/XlcMx/e
20BvOt4sySopLFRnMb4DLT4nl/B7v/pglVHhwuF3DGSr2dSLH/wiKByPLCOnbUqR
cgjRc+BGYrrquc3U3RJZ44zEoxfKl5D+VRVsd+VnBLuBYqGqMAkIucW5RiAu6PZc
Mwx9uxim4tBDcOXrRUtzX4Es9ZbyQ6SbN+YwXoEcA5H8XJIQhMucMgaUhEPMpzIw
IRPRYZSXD21JLYlmje7nW+JZtIuxJ7/st8N2ugUv+LU=
`protect END_PROTECTED
