`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bwt220c/634DCGSbn0/pYgZ6WN2qd5j2N/sspQjHGeA/iTbEGhr6mBTeICMiNy05
sydTEqkDSTDw5MCdequYTfyad4rbAb+0a21zKC0OsIJ8oCsMZBTCFR/o6QJ9gAqE
xlYcMxufbw1B3QidG97I0nTzxOL98K0++JjGG2mrbskQuzpJVGSPRbIcCNXFTy00
s4V7jqeCIaoTVnlKl1XnQdUny+8LSAkhcJxvmew7DXEjfEmmUr5NYVwll/Y9yxbQ
h6pgO6jy+BinRhFex4hmZ+oNCodlePHh/nU2wSIzRzMNn5CaafaQTfC+y/3zgcG0
0c5D3WbVlV4OfdawCS7SIS5GR0ezfbdyNYXcoFd20oXgptvA2CKRXb4H5Rj/PVWA
Ywg27Ciw+2QRrD4KqrCKqm9gaUH9xw2DSVSeIjNJbpmLjGPahXimsnM8UjxflkmL
IfCQaz9Pi+c9B6O1Aw4C/gRBTSyuBGfUIGcQk3vJ6gnGtl5+mN2gz5B4h1BfVSln
PiKSRF9zZLDYCO1mQLlA8XS//vbGHCadquA3c/3G3wpuIGVObOcRnK8RPrFtx1Ci
AAvJL8jnqXmnehZ34dQ8e7HsgqSzjlkHmrOYnuZDCdmgM+NnILaMNF/peUZ3lpIt
lGVd8JuCcKqceEy7z1YRgsbN7Qd/VJpjB5hFYBv51iNn9ol+SAwLiZ31PCiKopdX
dJzotsZAUiaMJzs4LritoWG2Dsc2w6mm1PF7Vj0ZaKXBdUGKmjcJ1c/Ry1jtPzD1
+YcMlRklqq2rKYOc4kdeKKzyfGBpRH9axM2NjSfH/aFipC70aGezIJuRHYUhEZd/
YEz/JHb/ajOkKmBoaSNuIfOuFai5AEvgKM8M5XncXlH1NJORvSGBL1INPdGOAd+5
0XSiTc+EUlGnsD6ZdDDZZqau6QGuvGQAScHO8FmYDzb0L3rltYRygTk+qaXWVOse
HurTgPHgNuhBISVt5bxep78PJBpoeQV2Vie78myCpj9zo7KkbfC7KKo+jGH/IrZy
zIZTaQ5940OP1BBOc+tVB13YaKzBVEcjGgcp+gbw/jL1fzY0dIwVNSzJBhRZAco+
9imtwOw6YPlSGLZfv7w0P1eglpsHtBBEbIDntVwUdaDnjoerXSk3+is0JdXI5YTI
AG2DCfgX9HxMjGV4IUI1bkWmHAe3iip8nF61uz9/CWAP/xkAW1WobfW67tjcGDDY
hCTRSWStdgoQg/ToiWm/fmPQckXnz3IzcCetDZQXS4P0di9JDCPJjmD96vFwRBuA
9GhH1KHCRJUgP+E9GR4pHQLgw4nV0+cSP4HMVg5+lr5Ps+2+eyM0v/ggD493NLUO
tyQ8W4JIq/ZVKGjksMCai2aPC2fpk1r35KM+gFynwa+Xza2cJ3/oSMCPDsHwyS5r
uaLdwtxiMWH3eWEXfH1bMAuS0zo5DQLP5iDaxKIu9oD6FI5eqK4aYMzEuCD2T9No
4SqqxRWtIm6PheAvHV045GW+0l6G6V99MwXKPPcL+Yu3CkrCQ2ZD5fHgBJ1bKvqt
JrNP2qTfkycoS19LEMOiXGYkt5+kIcfVu5Qazk9ADS063urOmhDV5OZs+S532/KT
CRWAp39QhnuTZE4GsLC6L2G7U7oTuje+sZfTUKTQfcwqbPW7ODusRLW1gQYKSYzg
o/lnH8UUpbu8FiimIqMD3/yr52v05BUS975o4j/aLJt4s+IptinlbO0NfskOPoUi
2BVRXC77/ja4GWTx0nhGuoJ0F2pXXgCDqhfyTWcEllEd4MMUtX39cJ+hC1c7llwG
2y/rLgQejLhmMST5IRDzoO7qkd4aT6lwaTv3pV9WxojAYZjbsoh3AANmOhLIDuad
9pJh6xyoH0R+n1b0ORAL3sWHxHax1JMtmYfQ0V653z5y8Cgx9IZlPJozrq4YfRzV
kvYUpgURNBP+wOFnKBFEL0qFVuDUeLoxke07BT3yvbeHHFdLz8AUwYnM07REVGUp
`protect END_PROTECTED
