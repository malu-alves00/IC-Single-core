`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PiaYcavgzS2fQ5CXpWL+QEGvMc6yR+yKDigd+sDhJWbdydeUA8ibdU/wyF+xAgkd
DLAYtsKuypol2dmk0nH98CPdGQc8A33bbipqPJzdZiY4uoXRWoK/fTxveU5hYnLw
HrJRhs+lztheWiJiPFvc5zDtezPkgCIXvNxlJz0EdfauzbzGMahYHDfq7lUKjWkP
iqpp+rk5IkqYnso8TTTrzOaq2SHzAO5TIRIs5IqaTAfimuwzxrvsgEUVGQkh/t43
n4JZDkl05f4v1mZje6etxVWELDXkafoM5cSq9Bd7/m9Mnkc+I0G0qhYEvJ8E01Iq
kJfgxVMs2K7tsMKDfGs9mHFz25gQCCqiJMaXkDboYV4tyXjKrSo6Tog0MRGIdzwF
YQuz6aj9EhHecIl7AkU7LDtSpwDil9KM98s9lPAS6NYV/WVk1OjBSod0+P8pqzmM
VmgpzjrYLekHIt6W+2C78oi4PTXWs14T47qvyMb++lKz/Ji88FEcic4dYemoIs2X
vmf53Tzyy1DFc35qpO3mIbdZTPs3iF4maFJbNi67JX3tp3P3A1l3q5Wpc+zJnvPC
Be7G+V+upVdH9QAuYDoeWKshCMH43MZwaZ6k+SdXlpH/kZNrQYKZ4FhthJpxgIT0
MQHFZuIyMXTIpuoJVzCGSZ8wXBYgyj96r3PD3zWYQ06MWb7ukG+P27Xccs3LKX9t
aq/nF17b9nMeeq3OwXAV9SIA9fCTZGIvvEgMB+Cthb7ABHGZLb+m2369hQjuWOmk
6qryF21Vk+hFIxVsBhGpPrICKGLjLHHaWeclJpa8IR+Ozs/HEMvmPq4OPjwXwKgB
N4hL5+CZHNrjVunhckeuYZh6UuB0GW9Jla9afGH7mABEb2z6w0YSHEOUYOF1JlcR
8dgxeOzis46JHCAFL22INMxeDmhsMUTisJMqgmPzuzxT13dkRE+bTkibsM9BsM7n
+fFb1OLYY8JEqdv/uQbNWLtQ3rCfZQ2rjpZlESWg+qoajHDzjwojW3zlzDT368Nd
i+9CM+DrNQ9xB74tQj65tYWlJMzC2pqPyOhziZx5y0A0qXvxXQHgp/61VD1tjibz
ZeolAL7jISvmf/UhRleJgqr6COsP8USWMuliF/rfKxZ8E3qa28npHKSKmsapw6Lq
v/nuhIE35iBcEC/bnSLtzg7Bt9Y4BnJ3E1oTto/3wUUDHDYFtMaWrFQZhdj4j2xE
AIQ0yCSvpRsUjs5pHidXmVbxucOiY+S12qUDzsjwIE88Gdh1rUrEAr+Ff+ewX5c4
S3aUH0xEj9HDDWmRGG6B9qkJyo0/qoVmDU8ScIsf308A+dDOuhyKFrOzdNkL/hqz
HdQWOloPxeLMUxTco7U5BoeS1zCESJlCHOIXuiJLuMGdcAR5DUY4BJesUg0WhiEr
agjLHvDcOAZ+xCun2g4iGZCDsMVzAOVJOzhZnqevGPh5cynAG+e40BnsstR5g3XB
//ie1Ou501n7ectPF5H1VFD0Nf6qFsVmzDsZuSE7Dpy9CS+wNxXEh7+/bepkT7VJ
xc7iInkcICdRH6t5Z8JVpsPuhdZ61Sm+OxU8iH5G2zsRWTGjMdoMzgwzdvqSxE/M
ty7YbHKTEKzM4KY5fe/yU23+aGZ7pnGn+61rYi4mTEmdKXEgo5u616TvEAwsIDC5
n+0Mqj9oCOvSkTV0HsosC+HfU6ESTipTY8uUIcEnCIaONa1PWd2/m9LGVZBzgZGi
dYwWFbfvaz1il6xlbCAkmfrZQtgHSA3vcSm7euqmCJepX7coApVDtGegwq2SrnTE
zx2ixMBNgVpzGJYc0bloMbtIEMrCNoIl3vIL8WML2TcFZAA8HK38Uf+o4EO9BHaC
VPUas0nlKtK1TUR1ROaC887cbhD+lU28wwyAKLo2vnwh+kJiSOFIeHBfLZu1N48F
Pm05OUDXBWYK1WUnRUFOTV/oqbRLnqD51Xn8JvlLu8GEkOO1IZAF4HIvtKPby+m7
7APCZcVfiBjROpmRcf2vSBQrKk/xOk1Wyk4bXTzZOfPY+wGkp4GLGrYPAbyhFgxQ
iEKn6YqGa8+pNAR5AjqjMwgRJg3oLVNtaLrh7FpI4CYavEJcgtRj5UYafjxfvBbl
A3KxW9xxv2U4x7N6fEtL7bpHjUypumIQSW0+XUS/aGpCzIoEoAEAetUPCoSVtGmE
6vfyy2CdqWgv7SVrgMuQ7RekL9SKLA9YmJrj1rOAMdN0zlua7yWruXWFHUQ40hFO
lxGjAdYts1ijdYYqROefp8aSNNaQhOhyTv+H7EIA/b+9kv247lwox4Cm8IIQjug6
fIbFvaAQY5uRAxpwnxbdcN2u2qkZ/pZ4P8ZtFKhS15FYqsOApt5U9KFRRbBYt8mq
CxvF5oQ2uQkFuIudXaHzkWrAWOMCGcGgScMAdUfPQMTntm2A1kQmVcQxjTqb0qX5
kj4owG7U1xEjjRPtxx34CODLf8t0EvkTnaITqGFl9KDiKbTLF0olVsA070o0nAgc
c4lA8c11rQC/guElN/KdWxNPF5Xfaqtm91ooenZKUwO9pLkFZaqq6oSjiC3/OVIn
bolYJ/3OgqI+sBEhOML+t7cXiwn5UXRetCiXujd+7iuLDTenmlaCfa1UyoODUoSY
rb4mAJGeRi+KNCMB3FsuO87sCyv2zRZ/xLB6ZsBkaBvwBB1uS6tW9eGKEIkpDvEW
+7q5/whUQIB5VEIh7e8Neof5P9eRPKiMuSOaMwSXIpE3dsZbxGV+smymJV1CX/TI
c22+Zb0RJT4gJa078Zz3E1wWxJ5grGQOyg3tx909GY48J6EJ41AGgA3HCk6BPsnl
Air2xbTFJnyqdXIZg/tYvCO5126gQYtcOtWyjJg5FtOsvoPa80Md3wOO2FRpDvdT
fQa2dqCABBely3Pi4ZWx6veqZ6rWvyZ+6WNsnbqZ+gpbSQD2jwHgc7nQ8r5UU4Jf
gpg8AHnl02BYXS97A/SScgsWRYXGjbe/ZKgYf9OQHwRD6vQnyD2aKecj6xHUse+u
3k7R8mJLMVMEqDBr7cOcKquJ46bqLb3CiEJi19IQSGQFGSo6M/OE0zu5NKKADnzb
5YwjU57zp8f2ZemXGYLsCc2oPtA6qLBP5eoB9xTPQGe4uo3PO6PIA8fAfIenAj/A
lIdz45yPbixp2KnBXjICE67gip+NJGBWY7qg6POtAPWeYWNaJb//3BYqeZ4XFvh5
S/tq4+HjgoOefRIxL2PRL+fcQjUS0fomyIG5GdsFacGpQJjvwb66M5ogFHtJv6NU
koJfMFg1V4SH8Y4XOL1EmHICAdopqHU/QoXywARqteIVxVxRDi2ApYY69Gm6xO1i
ldVVl99ez21d4XpPAa7I5fCGl49JD/v38SSxXrc46N79BdBNLn9W85JBp0HGcLgp
o73l7OYit1zvD1k/gwEYZIq4VBxSTRX7H146eFH+VNMIjmItH4rUaeja0FHgGx+J
NbQ1Da0yReOXY5ERfvfl4Z7B80k6MVEY7IAYW5CNCbTmah0qaCiHPRQv/N6UEwyR
+ighVv9xnpxd0SBqPGEBhyrI8FdzIS8Uol8bOqPH+WnLg0n/1QI1Wh6G19NgZ5e/
zqnxKDjwTdTT+AP6bIjZ0GkuoteTUEmEyT1t/j7AAGWnuvgi6MXT4wtvPtW/x80O
o/H4d7eP9BpCa3kZrPZXvdhQTurZ1k3Po9khpi21XZQxnpoDsTT3WVYpSWjHeyv/
8Ph7n4Bu1O4Er5BZ0V2G/mAo3uWj4mfBpskJVCPj2FF4paWGO4o0QIY7ZGH8/mJ/
O8xGVElHOy5uwOLkM0LWO8yfn/cZrms0O7IyvN4kwmHKOSoCgSzBpFLsAK23ZNmD
Oz7SUk3Ca1lVhGmYUG3iETQdz0YHHhKYNNHfm7NZr91EIps+yHBydlskUMToQYCe
+yvuOGx9W1HWiOObj+6i8prLT+0vVoXslV7s7O29zUYhJs82YAOCKTp7W8pES4KI
ZyIF1nkNoF/SJS3sInft9N12bRI9+4MfdHLH8vOcUSIeiU+bl8MHwl0PlZ+LsnqZ
hR67uyGKzLgsCTxlibnJ/X0NWpw7ye/Z0O7vs8SBBvFAjVirWhw5k+69dOYMhEAO
vjpbhtvacplSN0ZyP/mzcRVEJTmTtdbG7DSlQiTPTOlpkhP3hcmnS/fhz8nfd3cZ
FzMEuDI4IzZ/oCmeE3V9UTwII71859dhwwAnoxxtEwciiXXhK6GE1f9hr1mJQejI
jKGMbV7ywTtqo9XPi0DoEGiIZkhc3uFqagHPRPsYpSYb/K5KUw9Wo1uWQKD9meRT
cCTOG4l3xR0TCMyc9gKi3sVbv+b7g/Rpdy8QcKOlQgcCjO/frXVrLoUCN8uWwLeA
xOZXOQiqs0o09ga5YrQ1OoFVDM0zrMcnozAiEt7hn1Rw/mirTfADpjHeI6Mpb+3m
NqXnvbtPS9hckMrU1sn0SF265iRHLo1htb+IOdMjM60vWhGvlxZb0HLsAlA0rUyn
jBQu+PxMr3eJGR71xScqr6kO8QmWopabwdJ7FAx7dEr5mv1QJ6hOrt4EBqkwIq3G
l/NEMU46ihQH0ynKZBmIDEbZYWlwAC1tn9diaWj5MwRBNXinFwVTsdjArG4Wvg7X
9VA21K/12PvmUM4ZK0GZab0MujPuCNcNrpmv+D/ver8WvtpoLsnf287FuKct3vtm
uvCNWxxKi/1FTygBGnQsd6PMcMPs1hFMYACRdzAFZm9ggSmyGd2hPVTLSVD5QkhU
vTfAuTSu1pMoCFHyWWtYgywFCZCt0s2+MQKniur8klPbDX8TrvfZeQo111eWxRI2
5oF/UOPHCMeXLxfZ6JNYu1shvLBmfGB6Z6Ocy2RzhQWt9mmMIhes91kS5HEl2GXO
CwqLwZY2kbK/HVg78sRrRt+IgUK4Ok6iCW85wfYcD7YlJBfvcCG2wbzABJNVPztR
TzcgwBBHvEaLxmP3wHvEOmkjfCpzwaA3U1bfoUwu3WA0Rqs+d6dSkfOXSen8Ph75
I8TcehX/+jDJ2uVgMdIhQJIpfNAcl+tjSrH6AXUSxSPI1Kw/ITEPZFef/J57SLEd
52YXPCd4mEg/X1jBOy/v8Z/p/UdFViKysrHrIKdSzxwmhgILVp079oswGAAFs+bW
JwVz1JW2nUG2O81IW9bOY8RPhQwClUYXylvKghahwYDCaZZXg+wG42DzmmmyASDe
jqX4IRz+enb6+JU8vdzuqqIUDOqGLTA4hLOXYlUlJ49J8etUo0REpXLZf3vmw5fY
jD6RjRtKcH8EvOGk89qJzdTdbDztMJIGinaFFkjp9dNcpGHpdkfgCk/QYaw5tOvr
hMGpMXzCmJuXDhYVzDuo4FZM7+siDgqLSfzfsjjR4XcpV1O2vOHNwlYE7l2hiVLj
cmQC4lVajRLjt6qkobxd/TUb/jN/jXtpezhuDie+czHq9zst1hNkDmLyu7XffGYG
TAcx1OXiRM/1rQQ8eveR2kGPzwB51EacfPaRXoeitSuk8z5nCubu7fngUyY5AG/r
itEsBR7sxfeeLfHclebTBmO848W65oRYz054wWBzZc7+obXNcHVgeFgNZibmCjgj
EHNfvX5vTqGqvxIrl/vziMcu/e6zdGmm6A7waFatI5qXjaVxuhtRWAGzohC2QlsL
7my/UlKTMnaPAzE3FsVrnMdth4QJOxq+mwF2ZIclQu0wFjQx9UZlBb4jSuwcdSUB
1j2bdQKaE3XExsvYkqJqVmY4993GFNTn0pE3+jmgWDz+sG6BAOtNX/T3uOll6XEY
EEX5xHqILynFh+34cuJOvB2Z9mfjLKnWI+U8gEWY1j5xB9sW+hbbkoCdEyROBiNW
UcgWlxdl3sIkEBO3BZxihPqZdjjzDM5yy8Pd0Yl/zwfC4oQEgATFLxII1ixnorVR
O/MQYFYrISO4xXAGdrCzDTxH+d7EYTqQjSX+z06nV5us6ZvV/EapHo1MQZHDTk2F
BZaUhPwn/BAgabmrMjJ/2rzI5Hgtj+u6RuqClt0uHj3K/mPBpv446V7r89EV9X2Z
ckTTGGnCff8tXEcBH9OlgbZnGBXmjbOefmWjv0ZkB7F+jt/BNY5qRNxaN+GtYCn5
X5+IvT94rHfwEoTWxAhc74BrY1VV9OWk4u+r0+lVLO8gul3MyuWBjy9vJhDATCjb
BTvdxLCEa24+GIqbGQHaTSdpgzO/dKP+2c4aaKGEwVnYJ2fZRQ+uCTUeGaAOAeNK
/N/ae1EKSTei2wh4DhMUZbvvpcwhZhEzJDlIZQ3lR0wenQVSaIJUJCEvqmlszTtS
Zr3Ovv1/BgZJPaalwwf/NkSSvyqknNEhxbn0T0FjgaYO64WEA+P1J3NvXYCUPUt7
LFLrA9vKaeg0ns74kib6WSbJhCEFFYGJyEiTrXysN0L6et3JCatMti2wgc8GAuNB
3b8PqRvdXt7TOXhvIEp8MUvvoiRsfi6aawc2SPhGaihJMB0fUXo5RpjgZ7KK2zJQ
DxMToeCLQqhw0bY59WBPhACFTD0C66FXPdn+Dv+YpscyHZmTWIP233UnFgIgPdnX
MJfPZokhvckzkm3mhHyzD45A9LXRZulADPvKIeFkxRxaUk8+U1sY0SWF/0w90HSw
xOtiv0pl+XmNWI6YO7GRGFpmyKFEd/l01FKw3PH8K9ipkgjlkpAkIIXAiuvg0MBX
WUV4UG/+FZyWBEVF8Y+MJwGglPwyZhZa9IjIY1ScP4AH85HMYcqWCrCkk3BVI49+
4BnNvP8k/I+c6LOoQSnd/MFZCDVBm73XXR0nTnvGsrUemTiZD/KgqMprjcCa8ah2
Xfkh+U/Nb8wmv7ZN8biKY2ejWEnXknnDNgpZvIA3cHMEXYhEmEBNsXzg5ZhfcVhs
ojYdyX85GuhuxgydQyoYEVhLbS4zZzuVKqdKu43EXxau0y4ZROl02EcIgqaJsplo
eOM4G3FX4dtVthvdjQLxWSUmxTwYI9RdhzQdtbGtjY7dff5wRVUD9la3kAa3+O8b
WjGIt799p+g9jJ5Ywgeo/4gFOPMvgfHbtb9P95leoAJ5pcY5CAyvNvSMtwhe6gkx
5ogdzMhYBAeyfnD27HSA2F8tJ8IbuupcvlIaXU8Ob2y6xxAlSlE83KR/rUKMehXf
B6CbEcMkEbSJFsO74IkoltU9cxiawYFBJCR5vyt6mW0j0/VFjv0Co4JoWRj5QQRF
7hMehoSwpvoWbwB1BC/M7B9aT3DGd7ZBdaybTIM+DtOVT7NVKcgH29sRGZI67kxA
QcadqSUYR5iRyzJRRPAWDZwD8mkMvdq2M4IHO7qxoq8+coiqyahN+m5kCiXPBr/n
yTIHpqH4qEF9W6ucmIbIjBTqyI6Fs13r6J/bKKdxeTaAA2RG4qiP1pXGf8hzNHgX
S3NsCfVVKEARYoyVnb2+jW4cvhVbZxms+HWPLO292a3r57qazFMht/2unMjB2sqQ
piWJ0wDM1geEgNZyBF8feT7dxXrkdh7Ou0hEYaAM2R8TjI6UvgiNqyf0Krn+bg11
J9QFxh5PWS1weGEqqrhrdm3HssPbD5r0ukgAGK719oUCYV1Qeo1KyGnj/dnchT1r
VWct0ZA4XJVd12QsjVSK7lP+b9iPU7MNLql45+MkC5pZd8Z840C5ycKYNjrcOrIj
4pXM6WiLdLp2JxVfEHxUVOInZ/idcJxeufGbdtwWIu4qHlhvMQRC4Q+ODUkGE7S2
UNgnFxRjpcugSyJupmoxYLD+Udmzfu7NQ4LyEGOJXpduft7JXIaQ7jgtn/FgZfjC
/+LkKiVeTIVySDmPXZPMFEHJ3FX8hFREzALHdUMVXvsuEKL30dVblOefeBcNPSWy
SmbEJMlaAeE/jiC8k1DfWo/2xBhD5bFe5rPqXSIAw7SEPnm2vPj+Dh72lT14pAN3
pUDhoNzcIXYiR6u2wUENpGoqWyi7OM2To38HveKOQzurju1gx0YLpGIGioEcf65x
Z/46lTk91maf6IqWsm1JeD6YQ8UVdJnzRuY72FKlZZs4ks1R2ckI4GOvzxVdsAdh
AeXcWXVBJzbbaIe2ipMPowz4JhjtzfeGWLOyCltSYno=
`protect END_PROTECTED
