`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vaLbNyYtm8me7n9lpjC7nGQZkt4FSCWFDb2AE8d3HZ523FuSuUY+lJr4E7rW9eKd
W62xDKiZdUGhAhp0dVCkYxa+TZERavHNjSPtru8gvufBQN2tQ/0VfukIsYWNduul
Utc6I4LrDgXMP/fYIqASk0noVo6zanjG3t85tuIg1f0zFiyvXUdvA/R/su5x21AA
EB5rDkME09oOQdUiPulQIo+XsYxx9uhRCtDrd7Y48vI+GlQpao75s0Fimo/L1GWs
VTB4PCQqY91jQqWeYa+I7qC3ldAiEKkto1qkrxV3EjvLwUePtzRgxLFStu4j/tjn
NcckX0+vTJfZb/UuknoY3I2rgaWirWq+RYUj+4mVqgX7jgzmR19GPkzSu8HQZvZi
vycvMutzYxrHhODqk3hscBdxgYFWKHjqDOcr0s8tE+W5RHcGplNWsbgeMlilNjFr
fmJKSqmezNv8enhyHbaGqodZD3qGSGBeoLczBX5t17efwDrABiZJ078NmmdQiOuN
cbzEg+bSAZXPfFVlmWHg8vgB/FjL5+fvNEbCFXPYNohS+12LYw4EAn7RhC1QWcnJ
gaG5RW2mgA7sQtks+Hxc5GExX77bmuLLq+bY1pKAtdXHnOAHT7Z561tz4eMaF5tk
94DStYeuS29ghCD+APWfgGDrMeJUD+oBRylWjXUbEE/MbHG50cwEKaGORyYnaOUz
pSF9pczF9oH/6KEKplMLTlS4H9kHXZPSK5XiR4+/0A35xd0LCACeetU5FMBWdBvW
Z125MgATVwIpRzC4pI8YscE7Q3AK+ucWPeh2tZCYQWKbDhjsZdmrsHtgcGRmr1mn
gwAcLcdFJSGrUwRQbcT83WzJN+jASaYDPD4o+AixCkEY7ZnCV+CEgMYr8W37X0mh
rqzwdUmz7hQPgEPRpcDBDuS+LcwuOfK81TY0su1NLHl99UTNA87F1GjBswXdYC6W
VK9vWCJ2tS77B1n8NCPPgd7PSTbJacQeNAYQpgwCnCtELeWwXkLugXMNhk8p809N
tuwgJ6oth94bgval2xcdDssgvQ6VxlaAWy4NhQ94IAep0NtP8Wa23RymfKJa0qHL
FnNLT/zMCIXbhti+AXXhl+Huy8JMcAWHx+OTSBfQVTWw2T2kzAhaBn/48zHpzTre
cYSuY+QdX1p1ZOcrBZ+61otrmRPYnp7biZyJw42wAd8Zoi8mzmow897KABgF2d6I
LKuktwfJxqiyjLGsvmsPsNTN5JjMT4VWdEXcXf01BI0=
`protect END_PROTECTED
