`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Fs5RIw1fKora6M+Zz3NFS4fzLp8jSC9ayulfB/SJyN50mVlfTahuwWfVXTs9Hbr8
pNo+7bGNPCaMlVvwZcrh94x3H8MJ6p87jpTseVuCzZXH5JmBxiNvLn8QRsg1mXtr
/+5NYXzL64//OFrsJntNGqdbSgYcrf9HCDRAEVCcwQjGDAGBneqXpfJUiipJKnHj
tt+3y1xTdH07kemIyq/7M33RvmkpAa9oTmiyMQT5liUQOSrO92EAJLRbWFR+rXl5
lpE8Eyv94MxlemfwYDh0l1xKzP8zrlb05iKQczglLbPtJnBoUVJzZlWA5kQwsD7i
6s8avZEQAk4Cz3+boNiDYk5jIJeAmILnj/r9jTVTMmfPnqRGaAkNTq+hhCHqjKr1
nznJxswydQVQ6InJcUlQtuLW/numzRjI4JKNzt5kAgSNDAItDAvahNN8BOcnA+ww
e8QihD5rZT1iahY7PmKvqzV6nmdyWRAka1aL8EJOe/E+4ZwNDgumHVGOvf3ADMA3
idp35Eq8sS2EovEGhuNDIindCuxhUg4hsT6Uh++uqxv94yWlbFc9NRaPDOKHtmb3
tBrJRWAiC5e1YwQieaKv54RWqebJOHV6LB7/Rh1uoTqo1UvZpKfSW0EGYYjPCOem
oH35ouprXk+ngXtOu0wOMkyVl1d71XOC9fXrx1CJe4IClUchLRkWekW7wYuB10Sf
FOIZavxYS7rMYtnI/v5A9w/iWqK2eyifaKZz0K+x9ROg2b8KDcq24sVJshrwm/Zl
BT7Z8oi7CLeA/+oC1G7dcBtLjAjaftLzamPfSytSVvMg/BuLOQuurWaAX/XYJTCl
UsUcvjNe6kmDPWjk1FXQf5NRkzkUueFGVJAOCnhT16Jn77OWGocj7HmdItH8fDss
Z/Xc82KALcC7vIvWXhmmpqzxdS+epRktlUaKYKq35snXh9cwvvl+tXgKkNOZDQaG
`protect END_PROTECTED
