`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Sx+UpFqxcG5cM1Us3WEesG5vr2zF7YNFtCHVYjCR+yXH/lam6kukLr67xtpyw1J8
o0upMf6am73E0vbT3v2/I6wTbmw+ZP8YO/UOXU5MC7GNhk4VXGR1Am7uHAKu4o41
mUQQowbnK8LT3B6QQJNZsGkwxQETsA/znmbCnJH0YZWXoprcD/GPGBX7h6LsZpD6
nwANb5TYWztJKWJY6gbtDt2yZug7u7qgjWhx4SM8iEOdJiWX3iOkQEyoaQnecQPE
CrLNViszQsmdFzKKec1xUFVFtXkwQ5wLIv9He1uzN6a95p1ZjS3HeGD6EYfPUtAE
yurVpFvlalHQf6Fs/h6oTefGc5z5omoC8Yil9wHmIR/JDZqiyx94Y5m6PZBR3S3F
B/T9LUCzztE/xULt/Rcjr/UNhof270dpoX0GhRsanhDOFghYXqiOvao9ykY9MVAE
KX26290M8Bxs2/zk5sFUX+m6v59WAKtwTwgD838O3EY6MNhXiQ/+KAAL8nFw/Rnj
SESZ2DDT/JP1ZdoLD1/33OrqQHfnl0LcYSBSehtomFfKyHNoTyFZBkFRBPM6R8Xu
ThK59fA61tww6QvSNv+f/CdA/R1chRZQv0MpG/56jvKtvXPKho4lL82cSdc+UFhX
ImLewWojtNEkGRt09wFNmT+oLGKqAcVWHapqdr6bMEhYeRDjaF+C2Lg84B9iqsFV
DcaAnI1a/pBeYt622X7MdCi+rPl+f1Whxpb/7pF5YcUhEAuaqsuiKsMZrbJceFbf
0L18YOJMq4XhviOcAvSd42MWZg3T1CIOJgcVY+3vF87bweq3yTnUXDapPL2VBPbV
yRjS6gyLQi8r6ev1CsLn5FY93UkCLbAfw8wXQJUw6ZtNBqZklO33Mc08rktqC9ij
PqGjuaTk95nsfGF0GO5a4c5XCEl88JMrdTzJabaptia4hv3xCRQjcD52Zlxr2U8R
xN9CLCfI/B9udd/eRpTfL7bijwrnkCQcL634eBcRrVneI2UUwrmqtjYYzTTtn0Ng
6XlhOBgYXpIbhL6HQeyF7ssCaXsQ1qmXlfKT60HkIKCnVJONoQ0YXwP0+SUFSHI0
lamEBZyhbzfP+avwTiQpY3KqBGvKnZwbHK1HLhXPGzPxgKI22HM2VTJyKM9pIz+m
2HIx0J9JyZ7k5WrhpuQwIo+bN/iNmP3GmInpQjC3C9wrE7J8+lquwbIrxlFS3PAG
I/UEC84jexFtUAsnhZBbALJuwcrGgskbab613FnCfiTiEZ7PXaJnOeMkam0kHstf
/N5WGw1ZF4ZwR2MwvMjRE1gjyIFPCSiv+gNc9MzgZ9ifxGhZiciNdZ8RrGN5cPUJ
r5XaGRvy+f7oG30vICYT1NUUZmuUS5GTc4MDxeKZ1nO53q7frc0LIpKTOTF2S7jE
JuH8ghAkc2B3pORetj7uSnyuIMW3b62mu/OvrLGHYZ1MjfwTHhpcqTvmOhYHD/MB
Jo7RJjdAuOnuCuXQYIAJ8w/SAoSxsGQjCeLOGOpSJomc7NMT97dIWm4OSOAve91h
3AOiFkUUg8y5HMH+geONsm5yTaZCHtFVZoWdUkKdB+hE4A4fknifgOO/zNSazfoe
P+Y9ZsBLrUMVjpgObrmL/JMbBDJcGfGlXG40UzfI8imFvWw861Xgmgd4NDpjUKVw
Dg+R0d4OPt+iIu9sJh2d7c+PUwkW2tP7tP+1Uq29G8CAwfZ8vIOJau/m4G4f2OuS
NsnoU2qpHhbgWvIQfU/4PMrCrzLNoSX5mFVdkaGMYp549ipaCIC2RTTMRfJZLzOM
oYpe0+/kHfm8NDNQphq5LOnH7zq3EfINMUtxbWD6752m2w9dxr2RHWhEGJZtJSia
pG0Qda07rgQLRMk+oFTDUXe8Ft1h86WsWe2kR96HAUCWcvtrsEES+/ZGQCTStEyK
WngEjWcmTIZHH9FivLtn+PYJVp2tMdyFMPlGoY8FkrHyBaKJj82oj6Ngbw+vNzyg
HJUoMmBIy9NbUIIxWsyNmP0RdqFJF9LcmQV3XY6gk+zXT9EFSvO3RudsAFFmV161
85Kb4Ty70p876ddnldaiYOIyjUZtLEAwKS3zIhBUGhUpaYGBB9emU7b6H88M9Aa7
BjOWNVD2ZI/NS0jhl7VQwyOhNtmQQ1HWQmABXZp0BCV0vJy8T3CXA3gbvniWcpTb
6mZnnWop2H7s56RFYg2CBxNGSduv8OJBJSKVbW0Hvp3XwCgEbRupZzd4J5yTB8R1
5RDVNs1Qt9QKl9RA3BHiSDl4qjXFnCTni8VbDXkszw1dBkIJfhmyNK2s/DoMU0Q1
btJPRHCpZCTFNKAK2+MF5kCi5Ii7qnhWf3xhhbKbJ2v4jNW+2vZoBCALXVwm4ya0
GY4Gg7hw1C5zYKQmUr9h/lezxw+ph47fJlgRlsKNQ2uZIbSuxMPu/dC3Y+6XE2CG
y331FPNTha1CxgIjGMAmiscHzuWV98R3Xn0n00zvlHL2aDjQSo30tC6wuqp7A33j
L72S/S6fHklpsYgfc2gGcFTrl/6uY1eZcqzedpl/liXDx+4LB2761XFZfsKTebZz
rqykMQDiCXtA0UphSTgLrltt4b4FF1N5UbdHi+i1QsolsFR0rtQ/Q3AMjJjKyGPt
D4DWEl3DmOA/9izm2s+fWl61kUMGwNyyGpeIwRA0vtT1Lp7yCvP7NoHP/NglKY+3
c678uOuGhZyZY0aBBd/xBKOLvD67bYJy7Y2QywqweiJdd5UtUrxX3dasqpSBiwHb
56yB0fi1WXfUt60swndZnKIQCzt2Ep9fyaVcaqZM9RECWapFF0UTQmSvsa1D/iQT
uuhGMYvRNi6HFsszG5lwfdikOcLKgaZzBDJvYGl9eLlGh9Ux6CF0IQir0zGNyaHX
VHqyiI266gcTnLv2NRzNShvRPgikvqkkyB5ZhvxdB3O94AGAUXc7LGgf5j0BB9aI
dq0UknSa+QOpfV39G16uZAgO5/skD9AzLTNtNIBkiDJvbZq5YgUfodQJjsRAO7po
N99zgMVH6im4g/qdFZustvczTDiEXlRW2qMYVKECwg/6rnNcp9Ectoteyuf0aNvS
aeX40ocA5fc8bAH8XC7Mh8BmcuCtMm+sSeeeLLJWdXXu6NoGwFtdMGD7fw9H5LKt
bDsnwxQrMd5mnMIsuZtpA+6UbeH++OQG7ms83qTDK2SjEnZdflFjwEiFprnqWU1u
rvoFosdmPi0Y2IhXKX37LZ07t9XYIE/d/HDbHgvd2Z6sjpFILNsKjskoNXNM5UVf
RsJmEkugz4L5/fg9P1d4V679t6jR/qsbSZ6PPyR522AqGZIFlYJCJ9rduqqr/vCn
aIC7+eNOZsa467VuVZnW+gTRzLh9pbsgaEuw30X4rtIGDCZrkB1mBlyy5buA/wPi
TfNSPffbQwazV2NK7jNmpNNaKWsD2VoyKtgU8/+wUGeT6dx1NlCqVxrOpglOG6WU
vzIbPh115IgtJ6/xHVAf4RIsvwwJIWTuMYQNXzxdyNbIAS/76pPHswS2a+/o0Hwv
g0oJnYy6Alue5JuxTNHUwsHVvZ4M++6oYKHm3KpBr2RkSNG5bxEMQNHadySbigcj
BlGW3niQOM62tSLiTKNYWWmysQiDJqubnOXq+GAG3qB6rHnt59xaAjXX02DUliy7
g4kUm9oqJcJ7I21CfOR3CNMKzd5c4nkJYB2/BB2/MVO3BjnkmbP4rMp2I/RYrNy0
AqDMenUpizzmsvs8OFErda+yhp2pBZS76JNat7V4kQ9way1sy+tdVJDb56ivNHl0
Xd0QtVX9HNff9/jEGffdrhWeeNVTQEMqAwAs1GDR48ECWIHs6nnVJh6QRl/aoE9n
188tXXcem/Ci70D4DLsEWu08ztmlo75/ECxb7pNOc2qIb+rH7jbQJNFEvQ2NHoro
DzfXlKBkLa3hbVW3/bPgF6ZyMPgEyUCOmt8MxJ6qTHDGWiei0MkBX+Iv7Nq+ZZ1k
issH//YhXEOo9NWr/RjQzEDDcFPm8goOdcw3FwdhhLzbacojf9enpLubycQe+Ug1
n6wgPzQiHI/mOw/9R7a05KEy8cGixOU1zW/1xwooEYrLvct3OX7qvEyJ7nsGZl8w
G6H1C8E59tSRcWl+6xR1SASH7KLC87wzcEeglKwEuT50ieqey77yVj90jvPS1rS/
9eSRIhpZl9IqNjxOu95NMR9CNmsnaiGT6wVOF3PqcJRpEp04Jn2YGvbJTa5js6Nw
H6+GIPymPhL83MmEM/xvGiFkL7jk4FzHpsAViCaz342vJOXwVxmhbP+xaW92RIx0
n4hqjhtNd/OmnxuCOXByZ240DiHqUrHzHTWg+/MfICPZcKM5Zb32dmQcIC6t6i8e
YjPLes1BvyzgJ4gLr2/8NyAuIclGWJg3GT2HzqRmCFpLBcn6yoivlvss55LkoiwY
mNPEevVpgY3spbUYoBbui/ZTLjOSSelULDSbuLJlqVHnJg5yI4JA8WCRQcuHGmLw
6Z9bf1IAKigWBxJ5gKuxnAmmUXzlYYA1Cn3yhwHubQxS8lVRTyfSREWyuOw8QcX6
40t+mNObEGDbEYeWsN9LRDX7x6FtbW9n3M4SVq5LOsacMudLk6ViHvMpXrlcjqcP
aCgCwJCA2/ZkIiYJ4lbIFWfF1dXXkEDL2/TUy71kc1TfS1C/Gf4SEsvxhBcSBxNj
CcCuP6jeYO8ketKj4x6YEUyPYUSpIuOFsgq/OAcjQ4ThT8fKvgE1OHmvFyyslHj3
rT3GknM9gzTI6zyr/dE211D+vssidmf3YfypNRQtRbN95OlftG/Y6sFu39FItcLY
h9dNJgRtRqgqa8hYYuzeCb3k9mI4YklUhHNglqkvSRxJwXmN4MJbl9hPCGITvcOF
ZybEgKAzIjJfKKQEdixBnO7X7ozQAg2lLeVwCMpoJeNOVTKPWmyV+dSk+BTjg2b5
spuL1MlNrPB+Yu2ZinG88Nh9gtpxJLaRltgdc0gz+yW3FQ9BIstg6y6JS4t6qemw
m508AV7neOlH/Xk4Eu9eV+rVhKRUoNOmAVn6Xph+incH8YjBlSeqJ3CfWoYP+X5p
xy6bei0zessZisRsmMy+odZiT2wzTGQWKC98nNxopCsJoQGC7Fu1fWdblQ5tCesP
1hv+/jYbEhcqRcfj2raFn8Y6KbUskDk2DXnDfA4ECkvZxMBS2INfbP+duElNdDSm
g1jZ6eJrzzW+FqR5JGVNaAwmSZN9lLJDEmNGkU31bPQNFtI9iqWOMoo18HywdWTq
6RDAoOiHVH06SuNyGmOpwJ4bQzMhmZJqI5Gybgp6DEqdZOQsbRVl79YNDQEhCilC
ZYsxlT5wb/979rVH+zTHAWnceVnjfVPrtImVnV+bsdLG+FfLuVUZoJFpZfSJ9N0D
PaXuIU3+vpOTub/jHVPgP3ABupszm4mjCcqz1VK2OAxRnoabUyiDZ+b8U9OrceBz
1DLQxPOZtM+BE0HgAttk6lnZQ1ByFpZivkz0P03XaGVXrK+iBktqrkfo+NaQuLj8
plL7QwvFHtnDoGlLl4aZljYDjzRiDlVceX+PiwH1NSVo7EZRTtol3ygYnksN3zd8
EkcIbOaPwof5rlscTABrwpd/p2/qrtGh5DU6BZjuMlLuwNCxKnj8K7qEfJuZZjts
SNs7xHhB78U1V4VAvrRsbQiE1UCwraQjR/thmpjH0YtGoH5cFIoJygplpcnxQ9e4
2H4crsSJbjf8oY+bU5rjwgto5+3dLAvo6hRv7JwjQnAPAA0hn5Yuoj2vJ84M0flY
ws/8aOjD3PqyEfbBk4AUJJ8yWt9+hAJEe6qTaHbA02dJZqwg1q7OG7PNmOlFHF6r
hRFjIxpI58r1U427K/fDh8urXwuEQaKoC3RgAp+9wbm+TCAIqxpcNNhdYAX/nDvc
2aslqmXnehQwAz6ylXaG4/XolGhUZ/XSTAUOOvFqbr3U7XixkCdV41u3uj/Z9ImJ
9Y0tAx/V1yzNyQFTkpvy0FTUkd3YEgacuKc0u8Bsvbv2SJx7QV1HGyOTZqhNEJSk
YWdEtXpaH06Q9MH0RTMbDFC1t7nZrM0BblGCgMzVAtdD3+gMKQC1lRfPBddGBifs
Rt2iqct5h9arBSrSR48/Zug9Zn7H57iaoo3jiJIv5hQPEQ5aZiYEF0eIbgr+xGE7
HK7RJpM3u6ZCWZeWu5wKiL9PNjtmDbcGlP+wpL9Dq8Jdfoee8ghXt8ChaT9sCBPk
3Rdrh6XlLrBg+BEbIWUvzgpRMUup5kaCQ3n3CnPuN9OYEudiBovK7zQlsGnQ0x22
1hIr55Uobi03IW7osAbVN2DD2rNWzaKkpJ4sSrje1GuWefshbVWCeA1fuOElPEAC
W7j+84+Se9ly53F4EbUewzQZQDRsmNWZD8La32aB47UQIvEXOiii3wVzSCpkCn8p
AR2Q6PKVYQ40+3ayoq6t89PYozRkeHTOd361RkaUG0w2RJEPyBBBMYrpf7Aolow/
/KDf3aay08JWoqgzZjdC8BAUF06Dy9LdFH+2fkMmQvDR6QNie7+f1GsdeonqQ0WA
`protect END_PROTECTED
