`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kojxdrnsl1Dkf6NFTbZ4CD9eozCi0JVpBdlZDR6reH+jVhmHjrpmRmQ76P7C8psA
cnBSuGJayn5ryHcwAwL0s4t50XGuTybERvHR9Xc9US/BK2t6rVCMEy19WPKfxwes
JP7tE4h14OqdqkR/5pwevwt7BP3sBG4W0JhP3lsV183zbi6Tl8XpozKxB+K/2lws
tfGHNpIOWfjQ8fWCTKhHoZLP17ZLIIT3yNnIMr+joaYPNTomhNV0TMuNCIzsqhxu
pyIJpxihL4E2xsAXFVXkGmeq5kDK2CFNrTve4qxSXHFZ9ZyOEO2XZDR8ipFaAcqc
Uz4L32ZRi4V3vp/88eUZaVze6MlkRmLL/nOwsr/TImIdqvX6SewVsikb6q1LFgn8
4tqi7EFVERt8SPqsXmIJjL75iKrWm9cBCofHnzeJ/Aapn8YcpCP5QN2BE+WS1Te3
JPpaXpwUWtWdD3wHy6LReCQOMEvCqmFZBAXQpK1jVDOgYEv4CMyM5kCmtg0S5afz
K5R7+HN/yxqRD6aSuZFM2g==
`protect END_PROTECTED
