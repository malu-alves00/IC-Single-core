`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Gyz1gpRPouJQ+gQeYKfnbspmztdnF29j+VsDx89Ef7zCIxNO2fWqiVqylLZYEzcZ
/9LscH39Thp9gNtTcjRn7HSZE1z9VGJkPncDpWdlWAAUwv0XFEeru6DDpYcVty0T
m34pqLrYZNTmi/mzjT2t05+9qJbTge+Z+jOQ1ueXv2nEoA7EFvoT/H6wN2SXa4/t
Nzm090gIARfXCkOelWIejSsg+TuCx5nuWM31zScAhzbzDk3rqAeR4PtkX6c5m/dq
OTrImovAJrLaP2ATUOJkrifs/xveHV9heur8TcRxJGnulj8+ns3RV5idaRne2M3M
unOECWpEBIkDAptuwYuM2tojDq6oyPcSiKj9f+bSuPN1SICmCQijYcP5Fa90v4wv
mgmpDRZ1chyG/IPZN4XJifCnyuE2dgTMVm2+zQLyNdJ6AQ4l5c8wgdPsyGVKXqDj
dkWtpYejKYSLzN58x6hIV3RWT0r09IpEOvii7+UqCvv+Z0Q2kvBjurXgwrKGe00g
T+xliOPFF66dERpu3HF3B0b3b64d6vNHe3vi5TnKFMe1YCU28ArnJEWon06tWc6V
qpmI+FAEZ5kp+zaxyPzv9siSDE7LSz7a2eOkqvhb8YD4I/jzpW0vGjmFbGvWxbID
EUbEPcBtTI6huQRG96mTafPDNddb4F50ik+sQv5bf54RxgzHFaJhiCIOgVZaZfs4
OpJmRWje/7SD0kQ024vPb077itGVGEP2gd9R5zP+sCgovJZp/4L6CqTQWTdd7hdD
MfB/k8wUbc8EVGn0wW0nWvjvngamRiTJud7LaxobvSlkfQs4zqXYgXg+ypYehqhQ
NpjFzpadE9UHrUa/JAorW7BI2W6T8VlnE6MOXv3o5WhgmC8DFah9xjP8oOrze9ev
uui/sS7qnnNGUECMnDU/D0UcUkvxeH1qIRdArzaoKr/v95wNkKqwOCXmc8X75uzn
rTQgvHjwLQolVSCWV5xiZRbvCqY36/STWAQFn8Cxu7zx7p7WZpvfcYwcMzOBPH0d
VcW8qOlu5Csaxhyb3Iyw8mHwKH7jJu4yGwsUm3jHCBpBvbyhu2Tjtn2zmnZvNhs5
3azgEOl5Yg33F7HEXbGfI9Qzjr0+oGnlk2VN9kKAbfY9fe9/Yv3FGFZuOvgAg6nA
/Fj7zm0yI7qEcUhfDXe5aiWNHnOKPvQkY4Fa9oENsZdK+znsyf/y9eruoOwmKU4p
zclhVt/zWXadEu2NmwYC4kxfTZOpoXl1s7p0CW09/PTvP7gt4oV/oyz75wy36pts
e8mFFXTLWfrYFvvofsvG97dqOHMQSktB4t4Fc77+DUC4LI+0kxHbpdH3ZPwJwR/C
mkuzKTxc3Rb0iQRvP0/QxQhVExIy69usQqJoXoRrRWobxx1thZ5ktX8Y5PhbXEKT
2ADJPzG7g5jbo0MHAOpaOxn1JZlIZ5iSr+EQnxeUq3EIvG+6oDJuuL/paomcis+w
1QZf8fav9Pr8UtFkS/HCSKDhnc67GGB4S2M0WYD0/0NMSYTnpYRBJLOPY6d5keB3
UMuXkWMpOLFJ74phmDxZ4wlV6UGGMxCdYjIHw+Ae29KDynAmtu36nsi73XyGq/pk
y0fQnMhm8fX/x2vGszxE38RDICMwFLFK0S/+l5DSQ3SUqzSJB9moi/Sf1yJ9zSXq
NCnJKVz6aZ2KmhHA0cF7xf12WRzxpvRJMRfBey8UQy4+2b9Ik/oxuRh/v66x3y3J
16ZTktjzevW0iie/Q4fSjFBs4yNABS+V3Y4VkEaNuM9ibz9kiPp341tTZrqmBOrI
tUT5NNcqfoA5x/WEIYlgXjaC0YWECaT+YifyZTzUGELpQWPzcQpIiuUtl0lk8Skl
69HeTqYV7/bR1DtGPCyVCw==
`protect END_PROTECTED
