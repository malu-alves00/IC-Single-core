`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
r+s1AkibFeiIAGhoFRo7fjpU2YiFJIC26biVCTK5x5nI46utzb5Yo6ajs3X5hHB5
H2mL4z7bJw1TzaTCBhFIJNFvlU8x1BZzUXBE5KcITCJ+y7xbp87gAhEdoiW+uruS
xixNWNjbi7FB4trVsvPaHOkj0KTeD4nw34KlF39ELHSejIfQBquuefWeeC2PBTBq
rvhSVREvsX/MHScqnyDrWKlavUw7jOMhXltiw75KuRxCRJaaObearKm+2RQ1fD/R
qD9ZSHYrQU7cvwFxgNuZ3jeFQznUxQO4lMx8gHWZay4n8K/ag9LA+KfakG95lFPo
G9G1lMlQjnkEttPLfQ6kN/RpUOCgrO0aZ1oosR2pk92cUumsyg9rd/wE5F+4pnhn
5QIFWxTaa7aJaNCESrHuG5eo0WyvSID/hLsUj65d+XeBq8lLN7lTnnn15XsdiA0B
TU0pwGigN2Mb3rb6vwpv0ScTdfYmbownHBcvuu+DsRAiX0WWg1IJhms6bwat3RWc
pwyVRE0OVjfCVPxDTFVfSlq7iNfsIMBEA3Y6dvCZ0aQxGaiIxNYNyjyP2zhpV3JW
dazPg4GqNUOy8CFkVeCG1Enarxf0nfA5w0xElC0lSC1oIVo/LwRyhP/Zk0t5azIp
SdupNM69Snizg4ysmub/5h4skCOd4MHnPGhxO4sdimKR0Ve6EOTzIHhBn+3DUrXl
HuDPcac9Pie1l2QL9xqxt+f96cHp7g3xSAqE8vkr6MLyoG49JoLD1L0xiYp2d9gQ
FEjpJp5jL/n9dFLtfgIQEmWgjCxL7Tc7wI7AfHxNbq3nKrQrTMw7OqlW28FhCQ91
ASdQj4EDhfgbONDfKh8zroLizls98cxY9QOla05e1wIAU9RXkRc4aw7qB9kS8ERv
X0wqm6SOvF3SNnOO0opfA8J8yHqxVQKDGmlPWGX5+WIeSeDXg3+yF5WGg1bMLQ1H
fHj3wtoPmmrh8D4DlVnwh0UUlRQWWvdq4B2KxMbm4SwtB62DQ1EeOflib/nGC/D0
IkViWICcs5j7r402DwciguG+cPzESxwopzrqToC2DHMKFPjsgXHCtbMvqspHGQ/P
znrAPcapnteClV3XenUtLNHR8JAUHyR7G8sMCR9fuEprMsR0uGhzNWIT+S/hFPWn
2H1eC6qRhncdjceTcWuuZEWCciv1lHNM/1e3eIDrXE09RoPUma+Dy0DehylLwir1
6ql4LBxLVpWQ48KsXCzZoN7SInmzaxHKz+WGmGblKzt+erHkr4CeSG8bDysxFFQu
eU6uizX49r64F1lYkiJaICXyGITIB5TtaGQ69F/5t+6/zu/zByEiryw7AqqNCIcI
lamN/Xr8tQKc7aSXAFtzj4jnp6VZ5HhRLj0YI5KjRIEvqclPRvBhXTL4usQHaQQ4
X+oyql8/ZbGlEWC3vzGN63U2sCnUU6G72yw8loOWFaIAw9P06Fto6Jzohx2yMUJg
`protect END_PROTECTED
