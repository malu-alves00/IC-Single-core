`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BSfrgcQ1M4GYU+DX+61CYrcnjoZdkNTqulqTEx9gw2+TvDJZ/bOkqAMBQRfTFVaV
fof/KnhTz0YsDLv2er8er6jstsSnG2Uc6t+qTNICTvaU5pUHxQjUPsC08qmx9ZpJ
fNf+eUzNVOmzoglvbPqo8YL2N1nwAkCvZzaJ8aCWfvrdjIJ0awp4asGCmThKtn3w
Cip5mSZIyupeyjmnKF0yU0t/FMamiBd7de4GkNsqNb9KztV12HaG5MQC9W4wsy5w
bJix9vFeQ5LOdwDU2Nw26qiq72sF4Mw/sX/65GnWCZqIeMZLHpnYUVWjtfsTpmqw
AxO7iy0vZnx4PXvJCWq9RxQ0hpLgTUmtXH7YOgveIJ2LmVLDnqzvZSgzyrL0X++j
X8r2NQlcAluAzCrhxRvTpxDxlKfq7VwA2XXTPSMuQ3rQ9+sx85elSJxaMv45zI8p
MQKSN6N4sOXvyHwUylwBjzR6sRfz/8QMi97iWAlSmS78SGK9lEmM8qPc9jR0SPbA
2goipkWWVp8uzt188+7eaRnRCMbTa4hOAv45TevB41CW8dNo90Ni16bvalw3+N+0
NmnmsZDsg5KnwfyfxVB2hdwhUM5WU5ZC4CgnfspH7grWeSyQdoqy4Sgdn2TOprbh
Ih4vcxoMIRSXZQfyIb/+XGzkUODxliVSCRhy18cpY6yxDkJrPDkE5rguvhGEidlP
qw5qCcz10Sl7BLLPorJkSi9R50YINEWGEeo5aJvQokZR3qM37nBIF8ScKyU15gXn
OWU2KDdFuXGsCzAurprH2q2iZmxkQ54blur5oZ6RXRF0QxWCQibl1gLC9FFPYbZI
0POhd0l695oXnPOwWPJxflM2Tctw44hdtfNhxMHUk6gWVxWrjJm6+2b1L/ugwTKx
XRkPXyfY/oS4XRmeBdGR3IkSFbXD7VwTN7UBTalHjd9MvuIEqndV7GeeSNnKVkG0
We6nZvVq2zhoe/roa0pW4EynuT7QgUt+XI/rmlsG31qTf7TMcKwsaLYdR+mNM/zE
mLvnl0mW38hXff1gGtAXlnWq2AmUQpy3qEXfSV6Ucb3tpbRE4BHdx2PqJwQKUjM8
vM9QO4XtTOoDh5OrGlLQ1RU2E4hEaPtqOKMeHodIhv5/yubcMQFGRnotZkn4GaoC
M5oCx5xy8XX2RuISKbPTNXeasRU3aaM6c40AmtlJ0gE1ZCA97x0XjxWfh9UlrVJH
I0HW6wP5tWbRSPaDfZZWTm3yKwaNAMWQmhAstVn35cAOqFGRRtEOB8xyVngLTpMy
t/N+iF07gmY6qx8cwpbG5muuOVOxWtQx9d8a/mGZ5sbXRbJ/9WZhvk4yibO/3F+J
AV8pUWN6OH0KjSO+knqj64PEqieJxenZ9WSI5Nj+28qsWBRW7fFuI7gwuZxZDSY5
1d+JDlmxJutur7l340oVKpgJwVrFkSUoXcLMkZA+NwqTFd7k04IPUoU8gTrfebmM
Oz/PwVIRWwzx75SiewXvbBqJ0UHUA3e5iXG3L294NLmLATgzFASiHTdUP5J3Nyxz
dZOQfYlZiDFxg0Et2LKBfGjzK/c7FvFVW/W+3KcKCd695P7qZoaq0G96TImF1xnZ
zsJq0WHpIb9kjE6FEXmC9AuKosy32FNqNU8b3Wg99ZhvdOfe/5uL8f1s0l4+aADs
u+DreZgfeMo9lnZgHP5HoI57cynYZXfNuW5Qv59u8akaIWumIBAGzzJrX/I0wa0U
wDJrks1aU+pSP7b6Lm78siLgK3mmG6Ic06EcgmOUfi03FjZ5WnyVt3gNIQPfoSP4
2kdy+T1MpHmwNP7C1ef2NUPabD6B+Jc/egziVcUXGl5shSxOTzynePc0ghqzCpC0
mvwV779oDA8q1SpbJsS2T6HYtygEnLcVBb8IsrIVN2L68YZJAXA0/QHJtlr9iwUF
SsyLnbsUAGHRfkArc9LZ133ndRgT7YlLSHDe1Bsnj1XKi0c9LFwD+ESuQGFo1xuh
zkXsa0VHyFTQTeA3E7Hpi8Wags6Hjo30q8lHPjbUmsRoiwSu2dHAI045kD0dk1No
07ABwXLjKfdCYCIGnLVMtqLGRtIbNAuQHqHAfcXiCcIsEMBmLx0Ykq84CmLGULsh
Gf6YQTkx20oTffmSJEBTqdlNZi7/IvukhffDhWg2B5OGYsR0bUXODS++UdJiWWks
CEvbC4xOkl2D5oS9sDb9QzBOrRRldCYs7VTjcZr6MYMm0uC1m5znF4Z+LebFfuMg
Rme1PVonk38hGb9/49d3ithvCg/0zWagQ4nY0U76FCgrWzUaoKwmVr6DfKWU5yEf
iDxk8pfjo8ZvrdVjEPAwyfa7LgzpBIsmXtqqC/ZO1prr3sPuaWnVLUPNv3LXjnt5
DQlM8PjZvJf4VtLrdU80f+lrXPm4sKTenn8YIISdO1Grux3qMQkGMUXJvc7RQoZ1
cFjO7qG0vKPv+BlF0xdcfC64P6lKpnClq0shZhOby3EgXTgBAlxSklxzx2znO5p2
FM1AB2pVJ9rzyTbtZAfRhcak16JAija4yjGw9ZbK4W89c/wgwSunkYJWaNmK1vLF
r4hVc97mQmkrxTBP2t5e/08x+BTmNod7kDQXXI0Du8ZELOXOqvxkAHC1l3NhwHB7
GQo3KaWnSN4aEu19mmEJvxNX3EZeCsS4MR3griP0gr7oZ39z1H2EdTakBluarTnw
AnMHMNRo9PHhbgC41LhuGRghfB9XU3OtFb+CsHM2KWNNWBIYf/j2YwlY5kHixal5
Myx2I/WuHtG0DADXLoWSa0aHrZTzqYs28G1S8OMHJ9VuzNx1/hLVNY4PizhcGbVs
EgsVvE5Pvj7gqnxgndiwF7XAZXjHJv+jLG8eZ77EMGBjOHFNB8TB0U4H0Yim9Oft
eTbpsiIMl6u+qB5L1lqn2s8Cv+pEcqx+LtEr3X0WTK63Mx6LgfGpN52sM1DzxrnU
J7vCWcc0uY/tb+M7VW0xDqoyNhJgPrhiz0XKgk4B8Bxn1fS/aNZjZtehlCdHjGGv
4VRWn0G1yxVqgIpNnCnH1fb4z+pU1JqelNB+teLs30oCHwRYZbyRXuYjrAQtf2OK
Ek4TPvDT5QHRvv3gyO5YL8+VWtgrJNkCXJ8cZoR9jHRZxF6SNXB80M4Br20XD/fl
YuA71UByEzgHOV2KuMNa92msfiYLhRczXa1N6WIYk/q3XaPoddMRPJXIVr6XriR8
R0yWoKV9nj5XENXzfQOJFK7kxUmvj/QYDERJHBhOC0972DeaR8CRhpqx+aNOvcVk
3QhLfSEbz3S/xHtyaDkZ3O82FO6FY5hy29uXdB+cZ5tmHMecL9gaUrK/CRtOCEw0
WzqliJkEJuDpxGCSXCKWOj74mEEczjFbu4ujUKOtRU30/Pytn73NB/an9heTxjmB
JGUVruGX46sqIyRQc16luIv1OGa2cJf2Z3ImEkt1mTHucIYXc3Uum+lcDDOFHz43
Q8UC2vrDf/rvSU6vTTDV8lRrICtDDhkMKhdz/FkD6kjg0KL4t4vG9MCR/VCJxjHB
WgZ+D+SrI3SVCbw23CvlHAjvYOm42b5EpRWZHmn1qBOnm26ob7ZFmgsR9laBIA2y
dGOOg1Oxh7gAv5UQEJpQT4dbtLTdQ2i4e1VtmVK8DdQBx/U2kLEPVgdAdDt+cjxx
RroBUVHaidDwZmTnrdxRVx04Zx0LrozdkLbcebc0jXPkqPDt9h9+uu1YAJqYE4VC
nkw6Z/Rp5wHYHgPb07bKuvunTRfkUiPnC41zeWk2nB+K7H5Etd2GD48ew/6x+UeX
iHBa069FEik0y+cdYk1WJ5+mfxcR4bCOm8V/iulu1IyXsAJaLoRz/ZMXJ6Zm0leR
x+tJp8NZ7BBHeCK7MLXsFNKE0uf+2083kCcW5h4LKgKDDlEtaiWx5iJqIEj+dnuh
qpQR0dMd3wPUZioxGNDNQYWVSNfNmW9YFBOo4sDElPUB8ncfKuxwxNdq/CI3W0ya
hAmhxDcGUZXbV39m/e06M53/t2zfcAqyA22Pc/YSxElKXmkqbIz0c1sYHf9cxuI0
U2eCgYxX7OO4ijn8oYFME/rwpKR29P2XMVL2l25wmvGZ7vEkFhTaqlArXytgm7tB
OQ+HobyNPJKiw5hQt8Ez1sE9Mj1cdUdIzac2X1UWZ7/4NXNrmeeTG44mEaOgH8QU
+xtnFDkOcxZ0V2NUIQ3ZxXC1kAGvAgGaZHCC5qMhhJy5NFYQqRMLFggPRI9598RJ
66AFrjYxtVCYz8tj6CQnxHc9RUzPTdwzum7GI9WYoNqac5mgVoq9iO2MOYWHyaqr
omD9pAoXtAGlsSPuH13BzoiWhRZvfwVWAH/8zlxtOMpmEOJu1cXbVJdUsIIlAUUJ
/RMfkxZB4yo3KKzcqy8DVD31qRST32m21ZIgYuiS4NV/Wjn/v5Ald/pdxcyy5peG
14mu4K7l3khj79X1T+n5ie600FzqGm8nvLnV8GhME2fUeJV0oe3/uvA9E5J+Gopw
aD4XX8i+6ORB/cr4bzvd3xe+fF+8hObs3yQoEIiizLIP4Om2iyG9J8itWE6vwvOv
SfYlpchqXPrVWiymmimLBfxdF+MzMVT0AbGoy2e9PfuCviYm7X6oMCRx8DwEHUtD
nMrDXNqxeCfGU+QYaRRfWsVXlzmutzBRBRiVo9wJpo6Siu9isoTqzQPhv64skAj4
yEMu1z4XfB8o6n1KZFPRjYbSwihkpbO7JJH9Q0MeLHmDPr63JQGEwvELIvwmrie5
IeD6KFbLRr79OLwO6B1INpA3LkikNgGHFwXwSy2oHRRUCy7T5y3inLbJDzhvMVcU
PokZ/YRsA9rPEA8Qqz4m2J/4J+2pjIrL4tu+QgrUadgV5AMIh8hPL2Xxcj+O+kSH
gePCJ2Ll6cghzYR41MCJi9DWIEsYt9GCOcl1UEF+VI5bMiVfKs6Awzw7dJe1PZZQ
LuEikITK6/bbEPPL0dgqS1sufZWJ70H7uvROyTJ7R0+vRCHR08sDv4o/r6xDpJa6
GSpE8dGgO0punM8/A7DjRjtRRHsa07WyoGW/iEmLxjYzY4ZOhnp19raSa4A9eqNt
VkPcOXsaBxgDW855S+D4gw7YQiHZbq7qax1t8hJZCXRmhasgvQJlRR7ADNtA+650
aIy+GGmlL6LMcIDWgydD3RPF5ExjvwC+kyZdvZsRQSDJ000Omj4sha3spoe6JVWM
UBlBigS+2yflcg/BChqz2+UCNb8Y3DNlmRhNH04dKfeD1XGJbzD66menUC/rA7Dr
v0PsHbKc96ncJmM4ZfIA22UT/BD6642SNaMC0mScpCAjNZ2tTWhDwjaICOkycKc+
yZY6rynMiPhYQc1DsfRLFmEd7pw8EItYFFZWs0cvQ93/c5iJM2Ccc2prLoGuR+il
/02HdCgAdj/0CsUDCxBFGo8eVu020Ki3iy3h5+cUqtXFF8mYdb/rae1kdjcGpxCn
KETVo8jhuY2ySSDOVIcjlvdjK8y7rINLjIghOh72fT52vYr4f6Dy9K2n6yWplDES
A/D0hW1ZnPK7F/3O0n+6lACBs/haJn85l92aIlpPM6ld+/SDd007LjqI2bDBu8Bu
EBZmULGTRpTGQcd7TZLA1bOHnxi5v+QSrFx0IhuBXI5S7kBY83AKoPpb2F8lriEf
eNn+LZ3aJSBAI6Y9m33CgF95H3m8GANwY+yhu1iNm3fb96ocVb1V/whzF7oG8h/c
4LlOQo6L1ns8HQu9KV5zI+X75rHC069MKFIe2GSbhmTXQBSk4haEy227BDiEyRmH
HA8ZybLLTKZ9tocEsOB9UyGD1lMBK9gS7QYzUAtXonFe/h8PdO2sbm5hA9ZA6tZQ
V6ytAkCA0fP21dO1jcuLy2KlKnJmxcFV9FVvA5/bflfBYwcNd8b4QcgemH3FuhvX
Tc82pXI4Fj9Iu7CxnNDQzpVhJ3txZjj92cHE5+aD1c+JANHVsk3TYEXDRYacZK95
kHnMgKdUkfRaW77l3PlhPir+dkJycxNKWa9lFQCPKh6OU12+Tfr5hMyV5ei/xDh1
onvzG8Jsd5MBO+SAGyFHYSVeVI53jSrOvRJsSTHCE4UbOG9/Zt3SQs8GuaMhxg7c
`protect END_PROTECTED
