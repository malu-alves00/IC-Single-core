`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
h12JTzmv13KsPcLvEmDXpl5NstljCkhH1i3zCpocVkiXipzG/HE8TAoJ7IBwK5Xv
nOUvHiMNGonnkFNftpY26lAqboyZRIirfa5R4UCf3rfhVwr5Y2/CfPqt4HF+WPPt
GlQK0y6d4y2um34F5XabJS+g6exgbmD3s896xTJ0skZiek8XzJQ7y7kTXBvpxMfY
H1bkCK3pFcVHAF8/w0YPfn2c6y6RIILGNYNihn4RhbjaLnpFjYXj5mqrAZKsaXfe
zDwz6cP9+gqb23taKIAJBzRMObS56xSKFg0H2duyjDVtB7xLSZdywZ4nqTxPwcG/
jRTcUEXjdaON5kOtuWDWQ6gnxxlzsYgKtuL/FUoo/+nKjHSych5+k1L5kOncRr8l
swcSWMR/PC/JRrTVy14/xzZA86GsmGhIi2/iFn4Fvm61/PIqVQvQG2hxzJTxllEc
TRW/nnSMxdnZQFRJDoEIgxiM0NeTU9PBC9duOuPQlmSLlEjwrbR7QTFLMXYBS/14
P7YMBShSJieP6TOdhe8sb5VbdgvdZcAmb9Hb+9hwpXrguhbxSmtG47UAzDm9ZeRv
yT5DibUV9inj9uOIAZf+X/oi8brpB5D2Py/TzfII5TJ8J8W4PCttuEso7E0Ug6aS
`protect END_PROTECTED
