`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Cahx5SJ7u8vFDfRa9+zl57LL32WXusWKxdVW72MIDTUCBHZkB+q7z7UMjuN4+lwp
U/xgrs6hylqcBGuHJgiaA+WwD4UZraVzyy2YwuBjQXqHuqdY8aJR840GcM2tEYQ2
SJKjDRDs0cOwSFR3hWDXXbmhNVpLlotHhlSp1p9uwGHcvl51whWqttMJxfx0TdYm
0i6ZWlwT8+VEJI28qfdRiZUS5QeDE2Xrqrdk6ekBp9ISCf8BCRK5tYeL/z6GbSSa
d+mmKS89RVVwFw/oEL2qe45NJs7d/104/9sB22IJjWUCjP0np9vyuMc5ixI/UhND
ME6jU7LVdFTkm9THz/UGQdx+dG6UFt2nnqiUxy2v314jrQghUnso+MrI2R8EUdu9
jJRvV5qeMpF4hxuSf71O2tWxcc6ZTiV7ScZWhme6m+QB0vnqpAMwClWUO8GDrmEn
e+dqOMIrBK9uq8txkng05jPuVjvZJoz3bxP8vv1E5F6lnYXtPfTxrPg0ZGvqAMYq
i37YBapPsYaRQ/xphiSr9WhX0OWdO4jWz288IWphfQ7h7OLdlhRNZYSIhY8t/ymB
Qw5SFsn0ciNJLWOzGrJF1h35kQS3GRAKcN7oZaD6d0R+FN+GlPfcS7cvy9YEP2ym
nHGJUQneN0buMLpcclxpscjmjP4dMu9fn3MQUcfRFuPvPCy/SeaJEB6udNY0Cl7D
8BZndZ8eKugNnGnwT+vFX2zcRO+z+y0tAmAy8U5nF1tjYf9p710Hchzc+H05ZiyH
PS7JWADpMes51IZ+l8kS2AjOIkhagcqV6RILHIiadvHN/gLElHIYsKInr0ppKNbE
XuoLJXuUeogTOfvOfBxds2X3cgdMEIuFT/pOJ1i1vgESP/W/0arjFZjURlsMv/1r
nC9Cz8AM+xm5MrXvlP7OWFhoIlq3kF8/O3G1MKDSQzVuH9094pppu9YDLqS9voHi
w58I3inNmkP3H79l2BanpPxXDCH/bdozifo8R+5dHa3CkdQ2zKAWVMt9XNbsKQAL
cXoaXuJSrmbVFmrWKwkC2ePYoxiA7oCePcmdz3THwXMRmke5vIwKZLEqy6STYHzX
exp/DKx6dSCnJBRmU2O3oFxmlhEFBANLTbrnAPr8U1VLzMG5l3BjOpaltw1gNPzs
4TuRpwpCXXzs+EYIfO/Zg72iwH0Gwz6CpuNZVOXEp5xd0SxVICdXlawFYzvLpggn
IIkUyY3TLz6zgJElJpLU5cT7GDqIFUudyljaXbmyNRLfNrD4/Wn/lE3A22UvXIt4
A2k+W+SyY9mvntNiViPAAm9KRF/AbQpJsP725TQKWeMvpkeYeypttfHgsS1L8WK1
QmxF0o2WR2TxaGqHszKmoKW/Pvdg5lE0IRIeT/kd4P/Faw3qMmV3HKQnOWtAtrju
/lznNHcorSt9S0wCC7GL5IRXntU0GKoWFOLhVbZDY96fdKlBBySVHgE6H0eGnaJb
lMPqSoH8SKqw41sUS0sRsu1VprU3KaOGiBi94EXuejuM0S29m6B4YxmPrOrRBkwf
C6qxephcHR93PT3VNc1eQfvv+oPgr8PrV92LpmQbk+r6tKdDo92WRIgK3TgMBrJn
ImeVb68FmKYTqFOw2a8eYZW29ln5LGL7VoOGCCRvqLRLp2luZ6yw4J1xo3Nvm/+h
b9Ub7vDAWyNan+rN9uuGCrQ0CM5UvrcVaCB4chhMnIxWXoPpzEJFJIZ+nPZ+eRwd
vFVmawWkHpJ1f/fHrK7FMTYl3/u136SLSzbk/5ag3EDAxXKJqgiqI42wCvR1vPlD
3bCkp8jWsu/MnyMHF+vr3FnTs21AuQm05j5NgQKjqy22Gpjxz0V6dJKPpfhSFbBE
MpH2CK+w8mpzMpkNGMli54vUyd9TphZmY3qEDaASxAjSLhPuQEI52CyAZuSCalhY
pWU3pO8UnrTnL32fLwy5oeAFyZ2dtKA7D4NhRP6Cyo2kdIETyfi1OLjImpnsNwUb
mhHMj4VAfFAZ7I/qwDpK2YKY60LecGRtNQEW+2OXwgrQ8/ByHXssL8wtC/VU6iKM
gHYCqEHKBHg7Q3LjhXk2QePf3BFTBHQCe5PbOc6UN6ZyX2Z7SP08JV+KQEKSSTHF
I2xC1wDh6D50LkRj98spCSOLInFDcJk2cmN4EllxvAPeIF8AM3dRfIxGFvIFDvgS
hNqGxXRNyH7d36CEo1cssIRWKF3PvpQru8lQiUD3UzMHS2aP7LQhChAQKGsdeBar
bA68CLJFz391mvXc2H9VoFtzTn9mx3Z5rMnwKGT3mwmY2BLW/qk/pDzlltIS6lj9
NyyPmTddiTrphzvHi0abIrbo2bYP5JhxQVibGWqAKAu1eBD/+YLRMP7LzjzMMPQ5
9cLA6vefWUiPfb7AHwXd+fTDlgzZH0pOHLpX/XCz/9xBRI6iAnJBarO2jmOOO2mk
2rSQURFBch/WpwaHVmurQS5zTwKC9acr4YoShTARkom+jvMzXVnFMSF1kY5u52vW
Qlzm70ydKV3W2d2u3kK3WbzlG9bo0Jyv1qVhRVA4Kvsp5ZU22YuqXiWXin6kSg6t
5tEqeQEirfZlDNlm94jRiJaQfdFyKAeEIeSCUeYeiGxDxFxYxo8x+UrOKP2Eq5AB
lRo9kUG/gPn3jr8OnAtuggU0DDWIKFrLPCWf4+HHXCNLd1lBziIIXIV6kmGBHk11
zw5tHAci6Z1lBmq5ON/i8/xrMrw8BmmaqWZ6lzAs6XQY6xzziIpy9PCsZ0tVr3Gh
Jn7JjuFqkzVJSu4h8bWY/59V+31da0Hx4lcVI7rz54mH5qd155PFy9jlzYxGnxKz
O1UX9FpM/S1CN5ARBhIaLvSKc9oGC6jWOq8JkiByQiWzHub0Vx2MEV++insgyCpV
Fck11fVDDWQkkQ5uR9IH63ZoRbgu6rqgiV3+2fkBRZHBXPgA/hkUg5nK2k2QQlbj
lDdShICi1w4D05OQ3vHlBGloWQ5zh3NfFE1uJ86s2u5LLrg0cBStB+RAucoGlSF5
Aktycrz3HvG9FNF/5jLxQKgNBijrXp3iIdTred/YPrJ5Zd/bFFleCSFTDPTol1JK
qENnQ+b8Ng6STGYd5HOpJv1GTlsVeaVN8YafPM3gXPlU8jKtFsztEeSDqnelHxRY
C8X/xs74nsRoXvrB5tsyKRnGyqnAalWm74Vvgy2D5/IT7gvdSQ7ODBiS5Z05zIC1
K0ATx9YuT3ylbu6oQkjByrA3yH26NrxEG7gWpUpHX6MjiCBMr7qIgBHAiqIGggVP
eGTjiGcettzmBNCGSD9DmDxLnPTOopXiOhEDKWW64knjF8XalJ+9Q6wcxKbIzXny
V/zNpwlbyrP5dz0/0G+0mTUv69JFc7oH5KBEuFgpIVRzVXEFamlT8LnIxv0njJ7o
uTrT4fJk7OkPJEIR9NuYoeIUeJklgl1nr01zPfimKTzbOsaX3XGhbZ8SP2QtB77V
aBIeArwytaw5QmgD6jxjmSFlpB3653Ru/jRiWeFJwj7C+gut1Eu9LrsWJWu7ap2W
ns2zo6q11BKJ6wt8g44hh7zLSiaXPSbSXXhEkr/TYyTUOBcFcRD785E1B4SckjJs
Ew3mrJzcdKfNfnvFg5tJpiafdMZXPL/HBjBIK2b675CC4w7lIBMd0n+D7ZZXjx9x
yDwsxSE0uqQGFvij0Wbl+LgCDrzb0ZtAcPi2aVNfwKXkh+NkWITdbnCJZ5wuxwuu
A5/U/jljQekwYYsfdr6ufbGKBNzVEdEwvXqPbS0ngpaGP1anIWrSKw2FvFmTKEgy
DTnNSWWpmmnefRz4UT0zUkuFzlrqRzvUsflOcI29PubylYpIPOj4ZP2KCmvsNSzd
hIDm37n3uB/PUMVRRJarqb3UPRgV/wUhWqRX1jwKN0H1ZE4tBe7fImnTrQkI7KPn
Hy/awDjtOU6ekfYI74rDyonid4KNr8rwm8V7me5T3KkOnywOj9q5xG5Hs7Vwtf/V
wg5SAwtc5/w4oIr+vukshE2KLSBIbouE/z/ja2f+CqK/ImNd7jl8QC3s/YD0dy8K
OVz9E84gJuTbMnaK1CMkilUpyYA/Yvez9kdqupWwKsKcsEObRU0IeFHNfngzwCPS
EkKBzdvIQk9HZT64+LjP6XWXMoghP+sdM5wWu8QdwToDwu4m4dfQhbr6BZX5vD2u
M35WiAMzM9kcuOBaCGWeZkCp0e/SiKqOZ9Sbjema4A8kXADCv/Hq4Vto9ZInp+qw
yiSRfJNmQf2F/w7H0he5bDswUzifOjecNGRz+86pIBjaaVbAlN1QrSRfPkeQVID7
NAfX/oZMAvEXiXUE5nf/ECRTh228RvErPYR0OQGeOuqOdrSSst+u75xKTPIlm7Jk
zEptjXujp+JGsvDyNoAPXtSdWItn6JW5SKOaCTLZG+LxW33PwAknfu8An4P5TTB3
W6QERIdsNsskVfIVv3SN33N5v2BBBLAbC/r58V9FT6dvErHBGqFteEkBGOHodnRt
VvjofDM9dqKGdTrK2ixb5DzWQavETniVX0qt3skpQy4T118f/zE3mSbMLV4q/3F2
yV0PjD4aBKTaYrvre44pKo8g1wczqsRp/DD6QycBtnY4KQvYR4wZaDl4/A4YiDCL
Djj6P4NhVVpX/oo9lGLb8MVtaaSn/UeeZHHlK8CiPvQoi8mdClvI4ECjohjevr98
Q77pBBWRymCSL5TVyNMkMnCWJ4Ea386IpL0/Nhki1f/y+HZRZp0l84zIGrb5Am6R
ghsEjUvjUU5gb+T5ZAbL8ApvBscallL8qMX2WVQPKjWws1FNci5Inxlpt95EPDKT
e+GXgsyWyYmgSB9fRTvqBH1Ly4Y+5s8ycqWgbQ2IW+gmv9aMolwXzW24NKgr6kjg
RQy88prghRFI9bfSrfuaLWW5Wdq7dS3UfQ2DRCOXQGYc9TFBb8a4G8nTHlFLON+0
ls7mhCsk7suZOD1Ct6ZtnAaCtMYTl3HXkNPm3BrZsNaxVcZuQPhu3hqX89O7jDsH
DJHVgAESNXGHndKTQKMlVgoZrvtqhvGY0y7/+ZMNBwLMUR/9dJXQJn+BIzp4arej
94tSFPDjKDP2yGPaekONi4OgszfIM93EhkBTAHf067jdULGZFiNwlY7TudiJW3qv
VPi9ijmWd2vD/EAJ8A0Yvwv880kAFsybzybIeue0CDomolq4yLwisDMNjq/BBD5j
DwPoJLSyEpQXBEtcrFU1Qc3VOYhtLNgJmdn2V8XyN+50PRnxaeOojSQhbh/pReCb
tEpCMuymtWLKSDrCQWBmjTe0Z21zMn82amcy53YklXt7TfeQwP7k0kv0sqHm/IZy
9UckmVJWw59NpuClYESG4QWHs4as7iDo19wQJPhlcKf8D80SB43P4Gq0AKTpKAWw
GiHDRI0liksOAtEz9ZM1Cjwem7aro+h0+IskV/LRRRB0qPFxSFE2lAstGzGM/bMo
Hs0JFYaAPHQDJAX+RhnxKCWzP0TUNL9fsgQzoLzF1PVcODD326EyKil9U6SLqjBA
hYGrfohEswsNWDV2q13+gm2j1AWKnv7dB5SHc3jBwe3PEpZbtVrxXNkXC4Oz/mXz
KZ+bSnLx+C5bFZWkgiX7xhC5cnp4znzZTZTFT0kUkHVB9V7tPt1Xh/MpZ1fB505W
6CDBs/VImVWBbpfXU3t8aIg6cdeEzWlmKb6yLPybtvdU98n/cNYwa881mpzPEvr8
ZfCVPnmUr8TIJ3bSfnOH4wOPIflD6+EL8oKblfEvEotdTvSsxYkNZSzSygXjG0B4
SWKDcQ7D1iT8Ourxgu0AaOvzkocAbiLyoxlKzdtaapcQe5ODffA5XsTTIS+X6Sci
HmhCkXcDAkc7l6Bjynx5HytWxHCgwDqzgSoE0jP0ZoKyC7xXoZVe4ku2oIyW2Jav
rEbGDg3EENCF7XNC4QtnbqfceyaKNW03ILw2TOFv1uwVTwyea9d/bbN+yd3PXgER
BnOGhGjIhoRipW/mCWVYl2udVzPgEAA5IkPyL9OYm54Qcz8+G6BdxaOHVoRn+GjE
E3v/SNocw72A07CRJH/HWvE1Xar5gHbfZtDxX+a4vZA34klZ2ZcHzx+mjgKh3xr+
rW/gtKDJVDGuhN+/pzg8Z7BobW9uKiSMdD0TVKCqRszDcdQPCuyA7OrSUGYK1s96
j0uHylfBKhNw/kltNAHCFHZwtLoQKscCIVYTukqJQM8ywtBbxMU+JWCHVI9JAAnV
LIjF+1kPLqZKXW5Ppdp9Xz/aA9ssQSrL5D9bES/ygqR9SCtmfhtJWcZO3+gClB3o
vRoGMANFjY8L2eq1THrS7+SQu4LGqegnOMUsl9CWEx0B8O3QHz70EX5xLaBgS8tg
G6kV73ZVJqxMNGBkoEt6kyc2Ld+cFOdrns4VdkEq5E7W7i2ujhb7a7qjhzmGEGLi
fnCjpRFS1h/XxM1j4FwUVlBuiXSS4QFPKS7dypuo22mxV9cmi0S7vADHa3ln8rIi
Dv4LDLFNrkDcuqxKnNt4DEILtTT9YJaCb7T+etY73FTgrMf7l05v3j2sLE0cxWH6
kTv5q56x7NIjH/nE3dTYOidQgjUfMT6qQ/FpiInPRXU1g3Ec2BwDmd20Pyxs4gz/
nIQY2qPMtPzDELQfzCKrC9yBV5COxLLoP8JsUF944oSUURHadUFn5DXver0zRiCE
thOrPLNUgtheyHhBurZcpgWl9i3t6bQ7itTE0P8HE/pdRYxLXA7VIf0AqQyCmij9
UvuxWk0f966qpKZNmMgwOtClh1ML0/2kBDsNMCmwFbvV+W60jgwTI3Vj4dwMvdiA
vgSKRlDSvx9MweeG8R0KoUoKbPNURfwXz/uYy/C/QphyEKW1Swp6rfXAmTSmXKyg
fKwVc7Uv74zMjpXZApPTr0Yo6zCR13ArH+vucb1lTGpYEgHEkFZPB+4SaGQ3Fc02
mkejxNhZIbXXgdTt5Vi9GH7MRAWMEtAcO5kymUVtGDR4t0Ydh+IhRBOV7RtJXoh3
kYxfbaelL45ITD646/KUbANoYU2D+BsvfICddsA1jr/szc7Pwx+3q/hKQcY4k0rL
spSc74zyo8meHi2v5ZZX7PKxOZU0MB3qNAbgCVnG5Fby3fabo497+GrnLGl+c0h/
khWAb1EIv+XQFdkMCOfSIVIm6VTRtsA8bApoqarQeRMvHiLhqpnwfZEfqwfKFf9D
JhaOrSRYeamnPd5UIT97uH8RCIM7s6p8LaWOwKTWqH91wpChCTCuSYaOeZOQWFCJ
oyi+nsUYifxTpvW9FfpZ/w5tjae4Y5sruSEwEHHidqwqXl8P8Pt86+OllgZOaPI/
gYdRK64nrQV17sAV3Y8JeaaYVd7x6GXblPgrtC9tpKay4R78I8vlO7dsGRJ8Zp1h
1hBsWGA8ppxgLH9V0FZnk1zca7l5TgsUOokWx7c/ackK6QsfsGGohw2hSpf6CSPH
ZJ4bzPC4CrJ2qQHDoahFmE/6/2alICzzPVmDYqIOf6NvwonUGyrYF5wcIl6Ll2a2
3NUC67etM65Gye8aDfTHlaUyxc+aUmAzicnZK02Fj2MOkLBYhXRFJkGmVOxlKlpk
ecDA5/0WrYhHTRmZ64Rf7ZtF/648gR3IP937aa6CbYGfzFkArGQUU5BNQB2mn5fc
cVtsMnOk+ykHqX/bjDbOTyyJN1nUl+vredOVn8SfvM/jKT6ZH/79jhJheqUgDg1m
0/BdE0U+iMImxt3y/Lfl8ONRm2LowSQIk7DVZV7JHuIzus9uumtdLCMsmCUHETNy
FMGmBKGwQXKPpx12jYlPEZ/iZbloVF5R5bV66nbkGIeyEhDLhhmfFxFLZ7T3sTn1
PNp6wr3a045zSWH5Cp3jV/cP5Ff+WNaZnzR5GqY/2rj0tW7wsncHsYRIfJzsh/V7
ldJCFLclT4GkLIyc+slUUHld7O9QaOxwtuao/kj5Gy2u8CWTDWQWWDprSTa7CPKA
8MF+s5MpXXhjUoeu7RDSlaaOieEIsdnct2hP2pnnrMVuKzptM439dYq6chiVKKL+
wutfdtUgnbkqtUqBqXEp1QyvZsiZ4GsdoDuV5aLPpOAhWcR8oWLMoS3sbnPjDT8x
5QI8Kkjk5qGYaF5rfwEIssuYecdXEWqcOsYdp9mEibeiRcJTFTxl3bTCwFNWBjfE
60D2X3mlfDGY7Zoc0s1UHqsYXSSumdQkQjXgeTb8ph/+Hzjw7cHoFjZL+jo8YCWl
Ba2guvciO5Nnz/BIPUOfalkmr4XAWYBgO75ukOFHU5QXOt3j2iOgmd4XO+YG2XBm
opo5w9KvpiwRKq0g5HBkbOlciqcnqYiu17wC2R7dr9rMF9kc2K6sH7Hj6qJ8mO1m
0yeJHoA0QD3gf1zkKDg4IFNUIK2wv8edZ8n8OL3aZLu5J5Sk62UMSfyxtGxaow2l
atnFLMKughVcBiK7fN5jj152S8YF9Tr9nKKAHc0WfJaF5Et8scuLFF5PeZtTmFIi
ZIe5dNGuqGKH6499fHPCad2A06ZUuH5JogNCZTKwy/+C0YL2DaGNcdIG1jz7Dxad
kcsuL/WZVaiS0Wza7orJ5gq8zNrh7hzoSQI3vlLzyBWJ9IFSZw8gmtoco0Hr2Gcp
1c+izP//S4ytL7L0GBjw4GZVG0E/sBjHqqYTUwrZm/O1jYFXcModIdxk2wJ2xbI9
aqDVkzNeZFwPnm7G6xkkRCCoG9ZemZcsMoDrKPCLu6b6cCSi0a/qBU113f2tP9b5
hdgoq1fdJf4GtAyPoEADImcvbrchJWL7N3AEIaox7wdCFZSYtngniMlYsExDT9UU
vmdtTyEJih2H3tOPRmRw4XZzTQNwa3/WL8P+QOWxoCDmP+ZTg3A0ruSwhNWHJeMG
CmNUBzdVpF2yfs8m+TrdI9MsDQ0Gtz9wYg/0ODZ1YINDF+jcyArWSG79kQy81VTB
P5MS2ZkEyyI79Ls9JdsjAR1NfZ1SMQaXC8XJg6ojgGDOLT6/fqyEe+/hCafJBHkF
gSiQNxTo2lBxIdRgQnO4es8bj8wwNBTFWhF52MLh7vULFJCpuIzVczVnkb48GJYr
dOJruNyQXxsgMB4ZYGajuSjNCLHl6MOgqaftXeEIm6ZEMa+7z+NrRYyhfg4yzvbh
yO59r01ByHrjMw2scv4dVtx5FDUSniO32+3vnc0lvVD/ZwVY3akDLYV4uuuHdh4w
7Gjcur4XHEXBvOUtjXfFeqr2vc3iC61UZM/3gb1cQ+8w5xMY8Ws9ygFQBlnCPlWr
EA8Wj/UwXfItjPYIf/617szj8WIiKFjVAXtr3uMZKg26ZgXFMZ9rvVeUBwRGymcf
RNb/vK+bPWzff8wTD3usuk2XKiFwcy6Taz6W0mALcAJVCZGauLLdgTWjfZKmEb7j
tzS3KOs/iRE6SwRjooMujza5LGRdm3DrTxmH8a+m9RXeoSPD6iX029HGdxBoxFJ/
HmdtrvVW0x8KfJllkS6S5lkjfBthmj0F5Js2SxpUvUvVKaCrSuIsVMYVpKUua6QB
Ttmq0zyG+GB8kTOap4mclDzWis5v+TUmpxIZmPKbl3mO++60yd3O9mSp78gesLW5
dVLPefSXPoBVCS+acRrzTk1kzbM2uu+ZGrUnDTZWPzqrC/1w6rCDXHczAhoSzL8X
3Y68a/uaJ/W8l+1bAYIm3Z7oUa0J6l16LuNfZpfzy7cKqib8Zz1rXJjqubb6E64F
hfdNfH2UItUo5F/YGL/0N/JTII7gOyhZL6hS1v+bkgZNezZRiBEjeIDmMHBup9Rs
mf5ghx4ZfZMeeaQPZajRN/3KRRrAZcHelIpvUodxJTiZ13HBZEsO793vSyGmY0Cw
oKc+rsYrvmOUy6PmVy1uODoxjQZorj2c2X3Vtmuq1sEdSAM+aGei7fKThZwfKqPr
bAhwbm2yibIUgvdzEM4qm7rfCMpuKtW4B+CjoE3EfZnHyN/6pOO+uD3pOSK8SNSQ
88ijnM4wc51d4Gjb+lErkgMYGCQ7P3qmPiC7gexyJseKwZsZ6Yyh4J9e/3MSz8bK
ZZGO0lDY1xhjXcPk6tDBrVT9a0V8At9k6kFS5X6yWjQmXOqkrMRd41tCMH853flJ
eOqLuCBMX33RjBFCOeibIVrNgG/5hO9XlWlxE8/JTidEGyRgQj3MZ957b3GDFNdt
4O666jQxZS9Ufmu6hyzByDYZlNFI43x+dmZBRADFI02qQFrCJtwaZWm8QxXX79dq
t8e3fAeUWfmYKSfnQpVKOpFtZcWCDn1SLmvbFqJBlw61XO3/ZExJG6YgD7Crp+Hr
QY+NQ8Vkbp65G5GD63omcKGTJLUW0liEx2vt+9yr2SLguGtRJx12RFT8yBdvG11S
H/U54Qm2E/9T1+2azRQWj8QkUOOQnnOC6JxGbPKsKE/owgDwtreBe5ksaRHcBEqq
D7L5MjLAVoBYr+6XQbz0BraeXGrsX8EC3gduYTZWnQTBsIzU7SfwaKihmApjQjL+
Ytj+orNozGdXPfINX79poCBJbKcbbPjqNWP9YfagzToWUpIoGjS5Lct2aJOZLQVN
5SvCBuWBWBWOOKGugf83yKoqROTtsQk3lcZd5IrsKlbfrTXDfAQ1tk08ZIjHPl7y
UvBSd68uy+xXt6/60MA+kQAU/gisIVZjnlXHUQepCLEqZXWhDGaHyClmtwUE9NoE
lH91LtrrI0U/otXEDdvTp+ZpfcxG312CSrbRx8KTv9qxh2Rvl6ESdJocfD1VGP06
r8qR7azmn4mrGDYDQmikAGWTXdBP8aaDGZirsbksMvkYaXsH8aiH+w9HKhm5V9ue
aUAWk2SIbmrTjSmviF5sA27efBdTatWdVS+8A7PCq0jq4VqBUKErlUsJYC2yUeN/
eWw+X3eatb93aOhufDabrgnn8PZtDS7LjlBsw3FunviAYggTk0R7XXgWpXcEmmrW
f2+Iu15mWY1cuq/mUam1Fn0W1+vZQDUiblByOTu7oi9rehDe27LY+97HFRPSR1qw
/crMjsn+I0mCTs/Pl4kBri12FmG8h0TPEejctMVvSMa8xYJ/6qxeKFJ0C4+WgtYF
35iodIqQMK7u+pNDRsvWD31ixcL5hzOL9nXhZVysecbw793Erpd/Bz35As4fyNME
6G8EW+SF+QF1bLpH5RDQlChdE4owbE3mijQpxjAXxiPIjcn/SRR3W4ROTABv4fvK
jyCN/koPA3c8VfUR7QQsAwLmnN52iBvzVayvE4dxaeCp17lQzyFOHnDtNMBJA2TT
msABkSSgKjGu5uDAIQ+GVhyXyZ5qiRev7w0j1P6zYvjehUjSSNza7ttkRYg1DQsr
imGAlh1nMMF6gT1M9wAVHEXA2SW1N5vIGRPJGDDoZ7DDXrr6M3Q8nkRXGSzjZh4P
q48gu3y8aR8Cr9VW5VRH5ikd/PmxJC33dE7EmgqvYaurYCxgquiVkrZRuo9SRJuZ
Oz1pRC5pxD1bJguObp8KVYlnzdIGERGoLZ23j7RDCY3gbfHoAUIl4fRl54Q4Athi
DVhq9oz51hAg/O4vBY/6UoYo0ufV/hG6IFRhJhJNEv0ddY1sGwgvaukt6aLc3OhG
fjKzp0Uto4GrKz+1zGmGXWtvPRiBZi0FHU86H7Gm3nT9fWs0SBCW/aqnhdgu1Kqk
G9kzX0TAmeqe4Cuam0vnEYvXnXSKcvreDi+AlVG8ZXyHyg8smGGGHGRXpkqV7uBp
/ntC067bpZ3cSNdMkLghPV8iK74rKrnln/kYtZgoG1m1vTiDZ6wTt2/b1F98IOGj
6gO0O1zdmNKBbaG7uucbnfsbM+c0NUZaRQpg9Cry8neq19iUuZeIqfzeRwl+wnJ2
kMr81uzwY06ZQWH+ZSkoh5zduPMnISAw57+SWeCTQrtlyCZKl8IkIjenvcl5K9Wy
3HwurWQs6VCtXnppajqZWSbnjxpsOpmOkxooq/WkBlICt3yAOAiOG3S+A3fEF/Om
4q22vc6ommLcVr0f+7aTh58ODruvzLe6XHRU7pljklI+yGKGoUaBrnaauPhu9H88
GMKQz3LzHfi0RV7HoL+4lojHGfYl6XYuqe2ZQst5IpaAufeSxll/+fpxVv4YdZIk
xspdJEnpMK07M76ELoUo8l5Gjmdd2HuvQIBHigbIIQpTHbwuL2Ph81+iopsHqfeo
/uHRxG2YYDZQaoM41D6Pm38K2+5w8Kfdq5acO0GnNPhmzTwRH7L9ZurbJu0K7A4R
skVE5TU7NdH94HhSQYM6EMeazzRcJIraEWeFpRjX5A883N74OrkVHL3D6Ns8u1o8
VZzjkzvZxvu7i7Q54ebXeu0sO973Ftq3k7KcJVu0ErsaLH60YhBOVYIoj0Esy97S
/bEK0KzdGSYKzETZp5Vi2Douc59Pp7j1eiAMysw29v4lanhQ5cbJC4gVKi+IXczs
UAx48Zh/teOf2AdlFAvivp2R0p+19FqTY8cOi4quh7zPVt7Yy9ggR+F5HRrV24bs
F046SjgSl2VF4p3Id49/DEg8+gewUPOsPBFr9hKd4x+fwxDDjFqVTbiCYQ5yo7pk
+8/qvm6JwjJjem6kEzS/mrd9xFzQkZuMZ5KoQP37iFYjd23prk3+qmz/w0W02t4G
bVEkph5KsZJ1kSAniKLQI8nRfOa2sjv7gEE2lm7EhEuQmp14OB+xEcFYJydwXdtg
5qmRakH9kEkLhiFtMzw+Ej5kkkFn5JoPcbBINRuqiXYUZJX3gTN5LHONyX6BEBEy
gPMw7rW2a6zuzm4RgfkfCU8BhGwlssXFNzGTZgfkkLbk8DKTkgNUd42MNyeOABoK
ZD4XNJ9fyJLl5UKJTjUKCRZh/gR71U1rJp/jjwNe2zhwj29mEv1krdamrXL6xnWo
mpBTjHdoaDTzS9SVxVDLKNu+ARl4TlPGjmDUKhMCVymDOq+D3VmsZN+m0WTc6s86
ymskzy0qb+NqIQ/Tv1iW781wueMU4FfflZJ1mF0I7KgNiNhVOvyEA65Sv8CuqgPt
xU9YYaHbJckRay/kw6jHZ0BJ6r60ZuiM7EaRgNM5M9nMMYU54ahP4SR26oi/Ip7y
SWufql49gkCuM0XfV3AsHnju55YqEjBVLnLrDiF3Kp7bPIJhvZRk2bHxMqNuTu98
EeA3QTyk6dHIjR+7yhuACb/LCpRN57UgleZdXQo0NGE0wZJ0wqnzkY9gZ0rWlzmO
CK9KL9pdiQoGYnOBukuAxPFCu2mzkQlYoUxV9OKRmQ3C6PqQyjSOXnw0oaJgjqpQ
WTaj+W1vC8/DNkabcMlQJW+3/4wiZGMEfoYhjV2SzX1ut48QjBhMiq+0Sgig8NvY
rbUa12IfAlTNlFyL8+xJznDm5SMLPq6+iabXYS35j+G+hkKb9z9X6EA4gDAdDsvp
G5yPJroEYp4jpGdGhanmLTmMswY5Rm/4cBe/UtN3UE7BwG2y01iWzXchO0raoFtD
oeVyBe/yUyvUEOoeliUkC8OLYaQH4e+iZsQpoZqAWsf+yFOoF1ZwANdzKnW8xDIE
1nqABptQ+rZIxvDGvXgPcAkkYzTdPna6r6JFWmHScahnNwdyt6QSvdKhH1YSPWf+
L3pqI3umwd9Jy3OCVU9ZlozcBYyaPegRM9XoPp/umr/duFU6dWSZUYfbO/K0DTNL
U7g+RUa9qByyfzn1dDRHsJvZIbhZg/3BMII94VE4orvZS1qfwnLuL5XTCJ9C6HT0
WbRed+ECyXURaKiXZG2wTypx1+G0Z9n9GoOndR9ZzOBYiM6shlhsE9OUdKVkk/ef
PLje3rOgR7jdkaV/31Z31Rt3xl68abxQ8B3idVLddYUProDiYKRxV0l4H90Ov4kh
JWc6dxx0sE+kgPR620zs7bFP8KkI5gUq/7Oil0YM4KXAaJ0vLvm87w5NAKFgVIk2
IPdO7ZJwt9mARN2JOIQsTyb1LRAoFlH8sT8G/8VDDDWX69gbcpf34cXAa25qT7WX
0Q9YRw10GgFevD+OxboPnT1yceo61hDCvU7w+oR2S89Dp95vI62OMXbMAEJXGB9R
QGJuBRBR58Wv9ANVBJ3+NC4uvQxUPdRYfrp7//RQQ5Pl4f7M+4uSLaTvM470Usn9
yKjHOeT+moxFs31R4ovi9aeNWkEBfrbPsdJHf3lIO5XWIzEOZRkROTMGZ/KxJHnZ
ZfvcE/QY+rC5sI57I8YLXGhEr4BiZVfpVBP1Hsmj13Ff0VGuZrHiUUIKFSVZsJ5o
8Ezdft2DFNAW0aRBmFIR8LM3DRHoLMuAXF8DVQnuZog90Rq1mFIOoduz4JHbi2RU
qeXkZS2HPaexl2zBf9CSnPl0bN25AhcZ5cBXxXT0xk7ptQ4LQWTJB0mXP0B1AhGC
cCQ1UNPloAZaHSaexjkB+6FA2SyAEQLxWK6wPg8fbpijKZAQMVbQTqbdMr5dbRyN
euhw3Qv0pXAQYaYmKWH9jcT7b/vQFrTET9HZZkQWKz3BpvspQva68ryuca2aliEb
1KBJ+RKxK55EAR/b/suQWHLHFPKWkTlmCuZMEL4FeqSUQOAdR2brGTBP/WCAhL4c
Y7OYeZIQ8GU4PO7cI5KEFz8E0w1MSyLW862K2S5SRIw5k13vVkMd7UU2sR517Ria
GjQzri2Crnz8EeIkAiHFLfG1FtDC87GeIP7xIOzJOjjNeO6n5rTqFT5gM2ppeKbs
w9bnLr4LHp5I0VF0i/S5HmckGbf9XyzKxkblJHWbHl4Y83TseHD765RbmJFLsvVn
bsZu5RFB3zy2Lrua8iF6/PczVjhNcENycuv2U7HEO4sLxu0QKpbjIFQ9ifg/bVZP
N95BRNCmQinGsNnPz1R7N5Sk5PIWbwGcsEsvsgEIPtoQYmUBU5NNp6eYaCHrB/H0
bSWtm0LIZ7bR99pvd7US838FGuzS7sjg5V8+PFPFzjRVUsHHsSwqmyNm9RAgrG5x
DVu/hZEsDDBCqODJO67ynW5x6hyoD0rAh2MkcuiItQWPkV4RXhR21FjXOcVtaHN+
pSVFly/GOFZ1qUIxp7njsao1lkuGgFYpN77lr2J31+Ssw1T1rehIZTY2qpjRtbOL
h6jsCheqRGRVGz4oFq6E7fUJKpqXvfR2OOmibxgdGtk/zQM8fWgcDZQmGymHgbEX
Ng3gIa3axt+igI84e2rsWW/I2F6slTljgxjTv0GXMFYQoESfTfT6iOUwdIhrls/V
tHk+S3LZf41l9A2fYtW+b+t3+ePkRu0aQy67N2I/NFC3F2D15c9diohUEqq7B+Oy
jYDWhJDUMYse+jV9HYk1YbttLQCqvCq+ENINbJE4g6AL6xn/fOMUcCYYvP5EMV3i
e2B7PMx5lK+ITEFMB0Fb27Vmgyulo4usLCoo74TZjwJJxBySR0Pw0kIY+5vEpRSB
jHrK5RPw5WRN3/QIOdsXkF/lcyJloG3kEe/23bO+tNMmeX7Yu+W+7fjSYcpWWXFD
9Qt2Hr0WOrcdsPZykkaOXt9IeuFkDiZEJPe4LBKTvXiaCk3ULwElHA2FM9mFfwo3
rBP04yvO04hviautWFRz6Fw16EIEV6yqWS5PNdnqN5tr3/s8WXV/NdIG8GsMWs2r
M3QhNluNUCf2OhVS72axLHkLEFMboXAvqMAc33KVs2vqhARJWlZPDbLGDomg7Wia
c+i7suK6NTJmPVxyXROnFBwz8xgRDNioTofpEXz6Ob+V2YTxhxqfo23FT/9EOXQo
pUyTWYG+D5iY4urakIz2pKifyUJLQzRJD1PA2mSIf6j1XUv+AxTWLNHlat+BmAR/
jBicAAvkv8yU0+766ZifsjtstPB8hKjAfsK4nu4LpWXe7LOowjTuj1ZzHhJ8VuB8
cU1VwQbHFM91yUrVaQn8lnDvjcLkHwWyg4WomeEMDjZGpZ4FHK6n7ybSyRMQsgjK
owOG2fr/jlfkn++awOOyQO+LX8eTCMWUC5DAuk3DbL22KImcaunKPebwfUD/M56p
gaDDXlua8VU1EQUAmScRMB+WcgLIe/fcYW6E5pF0oZgWTZHOd8uXVqJvOfkQmDMo
MwoKVWB7ZUxKCa/QYr/u32SIPm6gD657nceRtNvVeHLpaFpuY4Cl4MxXSF4bhf55
3C2n218DCP47LlNzmNSW1wu0qPHOQ4S7+3ybB7CJ2WCBLyegwy8unlbosoUstTzv
2t1bsp/tqmbQF+3+fb3+kwxKVqVHkD9diQpIVz1CjlM88ZocTeyRSF3Vqt8UhW+4
Pv622cYHav8bwb0fmKgpA5vSPZY+lsyDsSQErIkXD8gJoIFivhZB/rcO2G7V9gmD
N9dyYR1NO+pAlrGF27f+nvcH3CclquuboKTTm5mdTvxeeubOMUO1GZHBxcNjr+Di
pPCYHHBATXfS7DN6HYQ+kOdzQUDuNE8lZv52jlxC/ftYRq3zq28c++Lpcii1BwWy
Q5Zo4as02FKFimqBhMwoDPPlA9xhzYiSx1PXLFgck+dGPKmSrLFtPiC2xI91NYsE
oL9li7wcJtL3fDmfyRPotrHmDyeLc0/lr8gUg2T/TWWXRRMnmMEP7+C0fUKZ4soT
Vet5ebrowGuWAfDFNgZmXqbl0BGYpvCe89u+44AywZsnDRxgfJwYwrjhCH8Pa0nZ
DN8c5xMfVPxPjWzz3NFSnmatgmGkU5mA6Mv/wByDkfEll/BTRcgO5T07DND2TI9U
/gDwCvzQDXSbcgkDlwODILI1HvQ+z6I5E/9ZekPX2ap7f5IOnB1ytPgdZMCHeYKL
mIJLlgxSiv0mgmrCOHvjUStU+ss8y+aUAGDhIyH8B4jxJSUInwaduXiM0+FoX4Ow
aJVIsyilkuoMqNk6oDdxbDCKAEvOIfOz1PZ8Zt7wbelIZcgZvV+Oqp797KhfA2fo
c04J/R1CWS2Ef+PDv0LFj/jXb8DsdFiQRWLaxCdz8zJXy610zn78EcyuCzptSc6t
E9zWeHWJmJuB6kBFHjSuHfZ2lBC6JULs1LpV+iv3dLFUAr6YMU0R1mIsgzzs1fQO
k96T8K1PLUmUEbC6fpk2gMsujzca4zvXa4gVIlSnCo8o5RoKdoCMprp1yLs2T5F2
ptVl3WHPAZVNaMQ8MGtMrwTTqxhdkby6rVzh+54gFlEkESEuQkvFVpFvvbXnqVQ4
eRbQiVmd5v17iAt3Pe/mjZ3JXKaAJoOi4zumtqVow40A2g01hNsZByZmEXdwMO25
v24idqpcubA8rKd2lzOwU4PgKwiXxtBH7EASX5q5gjW6FX1drmTVCoFEdwFNmBcV
194YGIWtF7bKg967UGUfF3k29RqGcY61twSqJOXUCVhqkX5tT+5+nCFSXCfXAA34
TLSoYu9+OeiLMaEDxKcNL+c7kiHKSciKAwzZ0C0A2qxVJDW3ksk/3LjowJf7yH8B
aG6A9hh2puVWTu0GJtoXfYgKy8rQJb+ux9lKaOffAIzjOQ4e3RuUlSknEOOsBv5X
AvheeJyqbRaQlqJ60kA9J8JY0hwqaHxDywvw3hDS8o577xcvEddI/Z+zo8KQ7WeD
kURasHTswhB4qngXK8uu2quGxQILzSA8BiVwpRFM37F6NI2R60v1y1/Ku+sq2mTr
RoQUQ70nlBrpi/vC7qhVdP5250nLxtyD+mRV4YGOBKoLy5do4vGx5Vxq9GDxCvkb
YE6YTm7z90/LEy5Y+kCjvoaMtRcOQsn0/XJ0pX8hgMI1WC0vrU9ExXMMSZYXNCC2
3cj0rLPB+9q0QjNuqYfSWHM92WC8aECs5l/vhjVe3lmS3uPzmlhh6LfrDavVZBq8
p1C8wxuLrVjFf37jInsdS7p6jjB3j59Av+84Iel9Ne4x3ZXmfxtvLSxfXEabGJlm
LxzQNT1Bjm8dmPe2XEEH5Pgs9hGA5ZsVfbH3oqr/pnPifFRBG9yjgLmD6TdmjUG4
bc3DhY5l5GhZbGtgdxOAQex6JdDXb+uyZKtTVfpRVwJmz1rzm2NFqywHMaw+Yq6H
k6fqhYoFxjVXQGZWhO0/NJcm8sCrk9tWo4Q2q8ag09uiqBKlxV73nbVYrMeyRm3D
gqyaYvNm/kKHCj1CgDGYK91v/AesSJ9YU7BjIxBUhbGPz9xTaUplgUEW5ROpoM9S
Za1aXDJIWD9ZynLa1VC7hxn/iLZymvbggHQxyWXMzjccs1BVxOzouQj9dY/X0Fph
Fcg0XZt9CFUzX0xKWc3HP49mjOL8i01cWqbivw+Ot+Y0tVD6Aqx3YjE8kxztjiNn
Abw+7KKTsXFMVHcNXQiGHRt+uS+8TOKF+oKs3EEavD+vhpkqZK9M4im/PRTXltKh
8UeRmwgaSkEJR3fj+a4vPb2Kx+V1Qk9Im/H1aRU4yl2XgT0XhCEc3Z1pyjoioJUU
zX636TBaC9P/M40THIE0OJYrTVcO5Eo4HFdil+WwO2LLlb3RB/gxTkVpPMJ2KbrS
xf94uQXyJYilCkOPSA5ep6DhAI2d+fXwukpDDEGNoOh7YxkspNZSRLIq88Ve4pkK
chbjiXgrg3K/ifsnnxSutVxsNuNsORzGyDFiz2L01i0zr33cAxAw73MC8AHuXFkB
LepazZl8JguxdF8XI7L2iRGi4/OloQVhjZ/Y4g/EUmueEK0uAlp46pxLvperTngu
94bFgtYK2peLS2tenMIl92n9ZgP4u1fJAK5kzGbFfB7kz2Cc728SzcFzkdFMSuqY
jBsgEeI8064rmccF1QrT80/eNwUMn8eJHuMqCmea+ElTmj0zB9qfYV7GxgV+8RIn
aIABeduzKGPH72DcuejPwMZixPRMQNlxe1wEbKItM6CgcQzu8mO9bwjmIMPc76nJ
nKSs8tBOl+utlqdqhzK/6H+Im8nsonISv8wGEoLCw+dV4py3LLInw/7Cx6h/QHU0
N6ONXzngvn+IknMIGn99VdSQRPP3fxxw8rYVx6UfL4XCiTwEyFAN+y7I2YjlQXzu
DghCvruRJ7mmhWFAL2BL7zXUqtxvPYLd5U/AOf5r/fEKElQuifoA7F6SISrrGQIA
RDw0iIuCiy4osfunHNeSRHSlKdgDW5azWGUPllYGajZmInCpmy2xC5Kgqd9HhJxO
56jknvItI/20s7abMwj3ZSf895QAijMogfpcPqcIJOkOipwj+pQjRJEa3HwHgxxb
U5IPiCXf0cOOXsbzWT0OiSl8zYQcmfuAw4z2UN+Cqk3C8T8MRK89U1K8tAIvpWPf
82ZDR2fOaxIcFs3JPduLneDBzbD3gGwUMGK29UjKQsbZ+BteOtkwc7Ym/D2+MKR3
fdcqkzBh7hWxZfzKLmSmeAmO1iyEZPvtAxo+vP2BYgo1ibW4nrRQIVmCEa5I2xwY
W3wfrV1LiYcPA8odl7whMPbZKu20UItHKRZRV1/yePBDC62eyiFqwzdnvyorif9M
L1JxSd+65eN68sIcb5lYylFLTPqcGxaTgB6oe2CNTNAWws+lrwvrHIehFaozI9JF
8zvQFwx/mA1wqRTZR+NUC+rDuiFnHX8Wz1+6gaFjXjRL6mgy7h2KG9eEpaeEwipU
7kv3CNBj32IUW6ssfVdWZv60z2UHzZ71MrjdPdgSErQT+VvhD+WRtx/u/NpN/aOF
QW3bgfnjFa9T+p1v05R/ZforOlIKJ6BYInUq9zh1wGjknu9bPUD+qZuapYNIQ0Sd
9xh4GNjt/dj5GSgcwo7ZNTcSj0BPhf2BO06E2AmEx04YclYFh2pV0AVtZmMXXMcb
Z/OT373OGWqNmExm65X5VpmJSz/f8BDQZnnDqb0yiTNYEZuLrQ5OdkoBzeLzJL5J
l3UD9E3Xz8fpzViLtkdbe+KoDK/tcvZU2/Y8qIAhY2Q0uvUQzh/e+JA1Kqsypzkw
7x1Gg/TpmRpt+dokjWjI8z3nHZ5sbDqWLNK3OafbPJGplNHIFHjdVB5k90tHLnWw
rkQBnpXIx+f2PBqeT6T4v9BTbOUNBR5er3A1BQW0axXfn7racpbXlcimf8erqH63
D1IPHOEb3D7eGEGr4UOmUp3T2vYqba2N4oTCjFMK2pm7ZXMm54OmAj3uYDmKs56G
mT82SWkELZ1Zx7HmhKUQchUycG9hjDOhG9s7zKIaIeRG8Mq3VAmk8iAOc625mPUz
7RRXBnisIrWrLNp9W9zEVYCL2lZ3A7gsq6OFHIEfgDzkQZzJxnR0H5DKcKKk3mbM
Xqa7Ah4zSf/Gefez8AcF5Neqhed0gK+Kbx89qx7cLTDDHiErLURSLw4hAVQ+GaGc
rHgeI4SwyyiascmduYVAhh4mGVw4SChk+FPOGHOM89xNn9yKWJqJMVwDNcOAA4lb
8sA6w1ahEt4zc7+Oc2hRTqyO0Gm38MQfiUNKJD2Sass07cO9wejWHmiEszCZg6e0
Lm0gKhcC3VjucPaAg02m+nnCzGlhMJXwDXjWgMhxjpzHE+JqV2nnnVI/MPMV9FIk
ix6jmeWy1UTMfV3rLMNLdoPYB3dYOoGCoUaEKjAHevqe8MvICzbzHv4oZhDH/dB6
kqRCVESwF3kIAExgV/fF4uEOMNj7PIEyXjTFjDrgW5S+8umu4rbkfvCjcEqOVjaL
yQHqV9v+pBncmWBlRbRtrpEMWrk/bm0gUxO2niy4l0EIaSvdX11mMtIfX/5p+WDW
in6iW1HmumgVvact1TgCoLTGJQcGKRfYdpQZ0Q6ewi3tC7OEoyqhBXd5hr9N+ctm
60+grt0Lg58k0MIlGsvEqg75iStEeCvlhYn7KkU2tB3dvgcxz/8dJMGfcTI7H/W5
qWf9aykirBfQWNnBYCsAnEs3dP5W0WgsCBTOgST5uwQMRLh+IR1jUjhARsdSE6o9
7yJS178fEcFMspCYz2E9dEWKcmfA9FPcK032qM3xfh035oRvq6I26Y/jYGuA0Ob9
aUGto/mf16c/kwMhBrazhcVQ+DJI+8zHLWB5gV4gxp7acLsJda5uRvORN5d+XDQQ
GLfZ2YlJpbaAUmpFGrXnsWzF46jCjvuDtdAMplzVcmn+Jy1BKBsLkAJeFpqU6CtX
m218ExPURDvL0f2nfDQBljuPAWq9RCkk+0JRq+BW+wjwkAUbX27fu10SMKAjsiBx
4AfCl50IMqKJXCROeedeC0oadW7Oq2R7cRyqieJRYRQzcsqbGFJ5FZdJbj5kAJIf
Mrutbw7JusDCGFIXXeHvWRnYFy86Eyy1iISqfYmS68jf9vC4PNwpJ13t0L9E8e/4
B+1goyl2Huqlozr9ibtVhA4MYUuaa4p9z2+1JrMoz6afzWsc4DmgMips1uqFv/0E
Tw/C7EdVdAFwi0t9L3gJNG6ze9IPfyWWE6w3x2tadYTDuLNzf+Vfq7f+dwbLHV3k
TZJG5/JGsvD9etGLvK3+UxQ8faCkdKPywnpxfU8P7QWBG011XSenQjr7Cg9EQL1h
XklDGo2ZrrDlEynaDnv4M0YfyNUSDmUFjsE11JMA2QA92Z3VuGLMjYYWeqF95CkB
URvuK02VFDsoP2TXGxC7b7fZEXWz9F7nVh+TmwSkSOiCYhXK2RqPQMx9NIpFAtjL
+HIXH9/aRIPW1LlKBT5vVqPam0tZgfafHGmu0P/NAWygiLikcaLiZmQ0pwJaynZX
pzy6KMsvQ55KQOni1Pyg1g9rwHhKRQrRCOHBdunI/xPXq0cs/l4GSkpRSy2iUuRj
+eiE36LGwu9QB9yTQv6J0yveY1XLZAJb6L2QBgAAZaMgRZSBWIXPiefhZdrctOp7
`protect END_PROTECTED
