`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ILgVAylycpBG8Ig08ieztMoBJRyfMbNfESWVK2aSpUCOmlBmFVvx7saoLYb2/3Bb
qHQyEE5CoFJvnNpOQjNDgaDHQZOhBHhH9l0OAYIlT9ZoeZafoHkMV9pHxF56eqkm
QcnjIlJHfVfT7M/L4jooKKF3IZ41iPP471K2YhPs0Jhmtzu4OOs2v3+FFTOXqBl3
Z+e89n4Z/V+PyTPOMdgiTXcnk/xRdJQ2nryvMarNX8ZNV624glyle5xRgyTU9UUk
1+LQcqKmkbm6kktoKtX1nAwl/pO87z7C8h2glzwm9IGhaeFDmIfAKTJ92yPMDtQ6
Rnk9NDm6AeqKcJliELviHi9ZnQLLxE9I8H1DK199hLIEQZxvE9NZ5K/LbbLodmS0
F8wZR3s6IHbZEeHL8vUqaZ2IbxSveDuQowq4DojyRiqvz94QvlixyDMDPTq78NUn
DGNpJ4XiH0AiV37bi89IffRVQw5E3wsfzDrtsd9IR3PCC6/cqGJF/hSDQMuETUwb
XqARsMW1TOWAYIbK80IbpohKEl4XPr6mus4i2fJFvfHOFw2vbtFdazkAsdPz1d3H
hE/wwyvdt2cNm6iH5akfnA/p/3vqHKfzWjUd5niPIl2DQXdKKM1/Ex5+tqyeKsE0
xupY1839JYrKGIIADdIcQxDvoSlCax0jQFW6youXNucz7RFqPjVsI8RzdOQaK1hM
Xu7KSxAhl6JoH3djCklSr5WaDRhaLacgbZSIeaObsmYtcACm59Tfb4PBGB7tbSZu
jnphi/3IzQimcXAyJPL6etn7Y1eiOJJFnjj8+4MZGY79FDzchjzmMsnP0r7f9plC
x5IClqpze3lYaPWyPrkIgSUy/EQ8w/WgiAvqzr17+ZgsZCR9xoPBPyL/MOTn+Zq7
zqI2CAZhkB6THmwLZ6tKZTTKdt6jFRlxEEkrJ6XtwV4=
`protect END_PROTECTED
