`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5nzwFG/n29SOaX7h46tYD/TsvdwXrm4/scjE2YEfAcaEecmicbu0z57ffs5Qa+E7
oGZ30sAtDU1niKRbXel+L67FPrXs8UIohFi91xPzJ2ITTeRBIbRu4RZ/QAF/ov7Z
WUHEFZCqzy6lOU59tfphx7EV0Aclun9n5c+1ae5rKiGKmdfIzRquWwkFhSsGWa/X
DNx5Q8FNSyuWgqle3HiZIymz1xrZ05hHabDMHjNGWcu+FMHNXTbZLkrOvI9WeNSQ
V3EMWaZ+7HHDfOlyi0lnQdtrVfGjN1zndkO8B4ovnGVtY/W7DKoWBuB/KKTcuBuE
ShjOlZiuG0euc7aY6/+xmwm0PGtRuBMCnzlof/RN6oR/fapMM6TxkaV37CxP1gSO
dsbYcYJT6ohxy+e/gqQW5vgRMEVE3uJWH5MhrPNHSDWzCKWGGUOX+TB65f0aDwBj
UGlNeKWhHJsEz6u7GZnmoZyGl9QQW+KRH5P5qkzsxInCYF29a69lSDhZWjZ+pleM
GVnyYzN57LrP+PAwWwBjPRWkJd9MXOg2g8Mn2v6jGcRm5WipXtcBVienA1LhBenI
1eK8AmzGQTQ8TOQqAY8dflqDmMgU6CX00eMtKOns2V3p0JjN7q6VBQD63xq3wxMI
bx4AGpVNe0pSL2u9ktQJgGcVzPWEikhz0XsGLNn1ib1cegN8mkwnMUKEdIMqSW4G
YrSRTwylvVDKkFQxEHc0eNa5+vAD9BlzjplhSZQYgPPATazrBZC+LcI1ZZ8etX33
qSiTremGAHyLSj63zwPzidGSzjVn9A2ItFQSOawrRfI4VNN8o+xERYqTNnpppZ0q
cPjH+SP4Uu75Z8LiIe7pho2NOLZY0LVIvcLTtaq7vys=
`protect END_PROTECTED
