`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JzcEut6n5jyIlThAdKgQs2UZE04TCK4PJ8MPk4FfmDwAfF/Tp60ZwRAWTuvnIxmq
B/mW4z+AVxewy3+6MTBGzsO4td2HYxMIaekdUJ7PnC+lEVjAxpBsCBIEXO1kB+Sf
lkbyRvgoSGtnVqrnyHGtzQvoDZ3UilVhUTEWc32uspd2gLNnPsC1GZEl2MGhaxsU
e5kqFACzJ3zf9WqKwtQornRQNfTavNMxWA313Budt0QhiYDsPhDCzc6amYfNeiLQ
JGsQGI8aQBgo45Gn/VHsbx1SuX+OT+FItw3I62mSfPw8iRSn8OHwcFIffEWvGhDD
SIHHF6uMy3XsP73X5ACUzlPikm1B8vjquokN1LVj4EjPEuXvHzrPFQXKjkimYdo3
IHCqB5xsOVxUtsgrPvMdAoa8JlBOhKrIOCD3w+YhE6wH8Vb6iE0ZfyDJXkD2lAyq
mYDyaXx5V9TdksUpfbVhtg+ox6HgB5bqyZDA2ZfJaKKfHae3gc+vVxuN/wHeFe0P
Rf1O4QhaGOuQzc0aPzIaUkBh+OG1bXZt2XI5+5HeHU8+U39yPXdr29HPf2KPgUQ9
kPPUuN13ozQcyDb0kdOKDG3zUoKAeNFPNOK+YocAd2BPyeqwMT0luG8/k/guQaAb
i4X3YcEq0ZU0AXfH+fv8tUkQjmZ24E/abh9EaQ/3l+Vn95xHSXQ5udZNz/b87bso
KQscgELoI61g5PLZjXfrx1R01sA/KSYYyYrEhRU4gbT4k452eRiu1o4FINFITcQh
J2hQ/NF/v8mDb4HfBRax9Kw1vldQ5VBYveqfa0YF9cc+fdtrEd+V+QhzHkRCD/6v
r+b6kYGBgVjvPwQWrFBCCnwPJtxXXkWUGyusvdh95+LAWGPjKIfhoGlU5XduyvXR
qEyw4rw97ITpyV3oS2Ns/Ocw/fMRgBBsFjd9t444XaDhhpcicV/2YxyWSVCUVJWD
P4MVxDuta2RhRtZNTyJojQ3FRtvKzaLlYTmZxFcNo21IHRvzFFtSpu90o6c4CLgx
9nYRFzfQP/phMjtJdr4mjuMKoE48QYnxCR9AWsbWbFlQH+TqYNHjTxDvrIs1i/0F
nW2y7VlvrHSzhrULeWhfQwJ4JS5VfmTB0+dM/ebiWiSFXj0kWF5sYneRkyhRZNO0
c2zDNDKUL9DwMsytufOIC3sw+wNMRBWGeSJAaRUSjzGrW1aQM8HcysDULmQc2IAs
ktDw6aY//7Y1iSFuG4ElOtsEd27WF41I+akxQ7c+D77FOBQpUUcJbofavAJQgs4b
hpD7OIqKpcAbKCyVJWwil+u1SLm9z/Rr1OKMg3W2dxODwBJBKkONN44HZp437MOU
oQp6PWcwtSpHZUJYRQdcHgrO+9mBmYxmgANZYzguSjKRWJV2egFosh1xZaX4Zqlf
hNK+nz3RVMa9pGn9vwxm6OeSwTGuG2oBuzjc5oYO8ieiNvn/mn5yLavSuHZa8iXC
GwQesw4SYshL96rt7yHro+zx2aUwBfuZMVvlL73viE7p/6zDF91lxu9jeU/bBTEh
IWTfM/xcqr/xskVb7kfleiCHooh62Qgv7xmD1sWo8aBpI4G0A8e0mfE35ZUdOfcX
2rRoVfXNETBO51mhbkVqjPETjvGY6Pc608nT+lg5K6VEKO5Qm+Kab0PBxlJUl9WY
wwS+7NasavC0PSfuav4YhZl12tkPiwO1bIH7II6O0TjA0Ea5VZ4+7LdxvGrM4Ek6
+5J2AqJ5AJA3KIDQmSnAxMcL+PnODeHaHLOfESGTH1oNH13PhCsAw4NuwGBT/af6
rXev75oDu7UkAsyxEYar/Du6x6HeojI/RSDaNnJMOV64EC/WTMgNnYgh1o6y1cPU
Pt3tcxGQq5INRcaTLod67lc7i/Zy/51qO6odX2asH2gBXM1SUoHvaKZ34h2YBElR
QN/ntVFSAk3CEdVKIsiksDqmo7UycKbiuKwO25tLaBtkWlo4AybUzF2qudcbY2Ng
CUvp3R+5qe7Tb+WGqwHYRTViSH4F+Tiy+79MgJ1Ea3hBlWrZvIiNgP1MVBQpgrk+
M5dR8lI5EOdJLysvHd9G/v3Cih2mGLQAd4Nl4Vsuql9NMEgnwXbCfPPGkheQTuTR
4pd0a56r4j4XTYwjTQgOkjCrn+U55mGii36ySZzBNLbeX5cwpPM6AhzTc/t831pE
T7eaLWoUFNJm8BqlpncHhcrazGlCNB3fCO1l5gTKNtkzzk12TOkpRQudLwcu2Bd5
o251kEV5oP7qp+rcdxPUf7hxUIaqHc93Icvz49zoqcc6yBjuUZccC/vM1QWSwAa7
l3u5TY7cNIbYicNwHMfr1YbZk2fHmIqcg+vLCpTvyQRWwhPpSpPIT84WSKrIPV1v
GuQFSG0N06NTO/N22mqWDnYnyU08r/blUVWfQN39GqsT5OdUXis1SSjmS+rHu5BL
WBUynZAr5W5v5Zt4+k2ZoaILSrfUq38PtQ9K9BCibfM3KtK0hFR9zlAKCKY+dqIq
T2H0TCqHDCy1IwmbAmqe4Kt5glVYzV6C+q4i3N0rga1eNSGJl97veE2LyNBjgypg
Q/ArW5LMA2ZGl97oJ/DVgyi1BZPKojEcw0+EPrlb5/YV8TBp3a0uZoQpk7B+4/kF
5fOQcIjarKIpnwSRewNArPpsMpx5SuW0n7tKwGh+YPC5b7kichM4Gg1uvs3Vcn4W
Uc84ZSWdGkDQUlnrO3FXRaQUfO+SydWRGNzg8a3zHLSzJMO3hrm4RlJGWdxLnUKw
pc6wQtG9tzuMW8LrtA3xr4LMAgZk6h/x/xEJJA2zgfHEZHlpjHH2ZWAAvb886vJl
q12Yu2HXeIGTIB7nnlSe8V3BhuF1HF+MWt2gMgaOHGHipIU8+6VPVrwihImhtK2z
/xUaaCo6vZv36c/Ou3RPuQam032nRPH1/SPf59ey+Pf6wt/Q2qmPHD1CoOqzjIil
pbirU0MPD9oB2SW3fG5N6v7ijY7zSmpBE2UAqkpobEQgiv38YIid5DCwCVYeb+Lz
bq/kBeBPJLCpCfvkyvRc1duCMMJxmShCSUXDJCGfq8kfphHGzHIgS247YMfFRjxz
IAICt/5+uPUqcBQZjHXsY/qhnmt77fwG1N6AkCXuEq+84NtqZmwsmgHglD2ZUSjE
yPNJ2+K0ByKIQwVDnJJRZA8rme96i6tr/ojtSL3aR7/Hz86vsGA5DRYiT3OHFT0c
eZqdDb9HflpkGwbEEnBM2wxizQiDgE+GEWqj5OozlsW5TCK5eyq7V9SPjgP4Xdzc
bhbblQcRD6GnbBb9XOPw3HTNl7hetSZG+w3z8XLiN9rnkhFg0HsbFvW5/strNKvJ
U2tVse0y4HNDMFk5rL99c8NGPxXY8DnmiLfpysSW95xC8iUPdWR9IHqTpfUM8b0p
JJ+Z8E+xtMCM0Je2sBupMeuFec+WQTzxBswPJmMSglRLzUiVaFPZvQ7gHh8tNcv4
IFfPH1TQdyBKZMoR0zMERC7NEuHDJg+iepzR/SUp0trRUWJ61rS06cedntN1u9jd
HWo6CnsDVD6e3pKxKYsyLpnWjBplv4cfEIu5iNaGZNb7H9Kws0Az6mDQ5EHjF6hd
h+MRyL7MYwFAjAPZ6yzH7Q3wbyPkK77KUS2d4L2D0+MSe+IJJK4A4lV9A8Jz+rk8
3/2QKuxxggxY0RAwGW4XkriPX9qzPIHkXaeh0v7IYV9z3u7LuqaXRGibGhidb1o1
OQFq66leQtThARvh4wKZMupwDg8Tlo5GHza08IF5NrGdOUMPeQjAx6E0XgaTC4XJ
4SI08OYpZhSHndS1tJ8SoXGJl+i5Acwt7/8bdPs3VRxU4G2x6Gu69ZAOIIA9kanG
3hqH5O0oeyAIsuNqHNFr7hrIO+i/WJlteEURVkrpIpzXabpO4ku0Ic/PqmyDbD4k
VbTms8bbtK2qUQQ8nlvrnoci0rRsB/eeiSAJchpBoboxc0/W01rwtS29xnFwYD1O
yPDWzkcfieBqNIshry3vT4ChxS9RSaFhFk1KGbBs+ckgqTErVbbUBztDygWt7QrC
io4FHPK8JMzm2Zeriunu9u8UmCQ6FIt/e9rF3cY9pYFzNM1vCOa9ZC05eNvlHDFT
vNChsnBETpOkQreFpjSTuKyKSCWOWNpK5+GH1TO44eUOkCyIZz1Owz3BFO/b4Dt/
ljx7MT3PdkNwMMoWPnfhIBzg4vg9CqddQoc964zkCZAq66Sbk8uHu/5iJSHpNTjJ
5lkGrlaoFXsbYVHFZdky56Vrk4n4Y1WJQXrDQmTog8faXO/nQQ0dfa3ZfCfHZ8jF
SnqIAVCgpSAO6eLB+WTpwCoqRL/hMQ70qFmtAjbKq66/X7FX7oIo+4NFXvHjhPiA
Un/NQHN29f9rsM8mziwOtCgYjtcYL6S+Aa3VopUJQ4U0j8FSZ/RV5QDU6geVsXnj
JFKWTYfByafGEwFp4b1w3eNy7I5UfzAspg2edYcNKf4cZtZBGcko8d9pykkhNweH
O5MOGvdV8ZUhjDea/mL5QNKzp+PV4at3iZLweeN7tJ5gcLQHkmguJFINge/A48j5
zxUhp2H4t3qngAYvZyWUUOB/QC9aVsIqR2zIZgk5u+M24JudZVTKoCU59dpTcHXA
7Kv9jQ2H5+WUIuNIKEMq4/wDOqLwe6Gr/04JKuKzSV/zaK61JMZtDIaF591Q3oeZ
sfbA1rS9VwSJG+9ul1n5uAicDE68bLb7RdGlgLnh9aC0kaXYwuwfbOOOxObAHjSG
hhV11Bn6LTuyz/XOZuJR8UsCWyjQO/XqCpsKjMjUXiCH5V1JBCQFXQG7Urgd97Ro
LVo31QBGK4umgo2ftKNFQVjtH7XnJFJy/KLa5rJV1K3b/1h3eXGUW0daMrr7hvRd
3b4yghFe26yA+o4Cb2jnbEP5KqMTT8OfYr5NixIicWOOPnCYwwBt7z5+5k93UxgR
AnwP0IM+qWOeW11CZ7mxsMQeT73AI1kNQ3C3PtG46cIDwUInZObsLpyxPZHpERfI
d+Q1ycsNvcpHBw6zv1Ho1lOzHr74iDqB8lusAV9b29q5xQkzEj+DKZLry4IW99/R
Z47flvafehaxxiREKC8a033GcJsTm/7aG8RLtGx9gTMFeC+z7Upsg87XcA/g2yOI
Ktbnb2lLAfzDk5OUI0wRMCUrQxQrLxt9dRfJjeL7tSVApbIDlTsQMFwxA35e/jl9
cuygdWgom/TA2YVo19CB8UbO5UdM6Md7AI2ffjIrQdiRTI2UO0zwaGDP2njJRJrR
OfhWyFSqE9NnSp/AW03E1443KhqqWnt6MjiX7bX9FuWVISeWmdydWEH2XIIdas4K
+q+7bvcL3f7Z9t1xSmuAgKmqijYoQ1cl/IR+yNE2DRnceHQgXoru3EavUpKrG47m
e//T+IOAR3B7ArUK4udJzhD2GB2xiz9ziIKDWTlkENu1iN4oo0qjTC1hgm8DYzkU
XFbzj0gkAdmJ9k3YP9K5eGa0rrRV4caKr/cqkp2DJIuUjcetY4xyXrOqexv5bZV8
WEA/lurvmKFRTo1afalsX53KIELYXfpsNiH5+ueFO9Rj8FrEGs+AFcqMFkE7F7h+
ap+NLfAWtD/OcUX5eBYbNb/58O3JeaaFnPtD/cRyb4HUgjH3tGEU2pfxLrwYRh0Q
c3NM3vU7bmHWxVoWqvjjQWWJIZFvlJvoRGTKbLCKgQwaJpDOujaYwFrJYoqAbbGI
UkGrVhNinpBMa5pqFy8ykiFBze3Y5Odl5TaVoaXWLkRcOz7QMLfdyNHG0caztVhn
zz6kl5nJ+BBjq8zudDj4MC39WAfSl76kuI8djz0o9m4oCnqN/Pmt5dcP+oMH47MM
2t1Is6+P0S+9cKxG4zDPVQUBQN26SfQtQcj7eAou3QHFOh3ay0omn+TDZFr2Gmxj
I/slK0CQ+IUlYt0nBgow6AszeHLSRNTuUjm2doQRMDM8l70LLrt8zfildbK0vRpu
5kac7ug+7aErpPVO1EQSCHwUoFsH6bYv1nPyvnyr+BA7wY3Euh/jvNrxYg22KTOM
ChKXfZIEnwIZRZLChQFhsNaMkPPtUivfsAsyJz2J/t2HVbyyUoSPMb0UHdwe2IaZ
ddpp9+XYNhpxcV7Ln9d8B3Etg0cOR3AiO0VRStHvw2rXRWepNAMyhnD7x5N+9/U9
lSDy+dkdi25+pxIWvzbQRYR9ny6qD/267kVKtaWBWq2OEC/Wbz9EhrGs+lp21yRp
XmMKePB/FGwN4u1LjJAacjnZCvDU4mO1LhTdNRCOPfU4JX+ysKjiMIz34aNJh3Gl
QgAi2gXuEmfpQ6KnohKQupHnI0XwAOLNI+mSXYRuCNb+1R4aDW7d7D/BiId9tofE
mQBEnNFWQDs2iRnnQ+yATwTYw4/Fn8pPwXIU5UsUfQ5aYNI31Nh+cfJlChiUw9vX
hffqsz6mqCFZ0BEoePGm6jcdAFIQGCLZPEOatqXQMIy13PBrNBw4SeVyTLeft+vY
hcJs1Ygh7kmusBHzAnQLY6010I10ztwdC6jYToD1/D8WOLB7S4NpP4e2PROOxXBN
OSWJWxaJ80aVtTfd3HcGuBOHlPIS7ZCdIhkhB16prEFGQ8of7MwLuplaiBIRWdEG
NxYubnhDBag0O21afpBQkM83P03T8pIQzjNp+BuF52QPUD/RfQKd8a4Skx8Lo778
lcGU5rtDsy6Z+OPzeNv0xI6jbHY3Isuk1hWpzqHhc6mH0OZAwhsJR8WKeBO+qcVy
H8CXOnFuDR+fk/KMlutj26v8JSdg7AZRwZdNan6oWK+NullHoKxNbzjulLL7t4fd
bhvj1owX01v/Ng4RxINWUQFsuKnP1ziDu7euiyoTN/NnZFN5T0M8YZP1bWL5jfQB
tsiENoSHdKLsPYljZpLkTjqWk7qwZo7fcN6h+Y9emPu95n1bPZA29RChs7T/6GKq
U8emT04247L8lherO2AwINqJtJtLwTY23nJUMAUlZJ+5dUtbTwRzy7Mk7ApH61X0
yMIyCdNxPnvJBiXxsuhaF+ZkfbzlK0lhc6xxYCEGUcZAJweVpxWcKLYru47KXXeN
tSG1o0VBRZHAMEOzF5nJ3tR4ZyzL1u9v02AyLdulOizLdvR8mdRnkE6+YPk0tXB+
N7UJPsF8F/QBCYE7rEPzCgDsXhvnVtm2eM6ZSSLExjr2o3Ky+tGuvs7JxpsssBxX
wZNgWTcfkUb0QH/THClhdTiA860mtF5PtLxAmyeV4Z5/KDu/Tyqb9Lc6r9oM7Uwc
huWED5+pWqPZKu4h3Y1IcNtpMltIlOzlKUKSr81MKqiqcthXTa9sk6P3sIbttGh3
suR2OPz/CQyAbGfNN2L8lpAqTYwkMd3kUowR0dhlCgjSYdj/aYqmeIzh5HVzw2+I
fCfesrRKtlrHW5Y09pMO0lSJdHWOhIDHVh4y6eKbAvXW0ZlAO8fU1NdrXkeMenLM
zIAmvUTO49vmBwvQ2R1eza/LylvR1tCSZP4snI17r2z0RIh5RUOJhba0ue3AAoax
Af5ufqhECDQaC1jkbuTWMPzO9/Rg2CD/fChgcVW5HBQFRf3SSVhHalWIY8emD1Gt
xtY820YltJCssjWGP/v88452od6Bvd6mdQ5gwAkXy+MtiIsZRhc1GlED9dkjECZp
Xyq0Mvhi4S7UMPF9nvtMUBYeVpCg1SHbWG7rurkebrfTbk2cB2N88ZIFDnH1njDF
libE2SB6b/R+te4zc4hsbAMChpWKzoIKv/5Vb22rj05FX06ZzTdfC0erDV3MlUX6
ifnIGMIoB+nSlRfU+n1Qhe5p+XO/n/pOKg6yzDO7oASNjyC/BTT9K70GcghLxrnd
qFnmDcVTA1lZDsIoSu5ej2cL0KNV1zCaCs+ICKxjYoJIyQ/GB3nZIN2xtMeLPkRn
ueH2zifNfM0/uIifu+scSnSNH7ebJgChPyGp5/XoCvp3fgYo/rOg2eq9mVCiawoR
55uLLIjSY1aQH9JFayK1h/Zv7wPjM2cmUS9xEyyYN7xRx0hAIntjcW/qEi3c8a3J
+IeQY/t72U8L5+nYLkVx1tGBDGzCl37g6wMNOBz7AcUJE0Fpg6aj/ZvVFPQSxo6m
0xws+Qis0vuTM9ruGK0hvLI6caV+FJvx2Q/J6+lYGCEAqmgPeCdn8r6xUgLAqoAj
GVXA1s0ZbxFcuSZGukJrhyP2WEXhkQbrWcN+VRm3q6W+3a+jFmx12zyAN2WM45kG
hLMKxCfMCsd7IWxZ+5fGML+lQRaFhr8xKfX4ykHlaJ8fnCIyua0e0WSmY9qxU5Xl
M4d2LKL3Vaxx3QnP2MIh1WIFlwGlVzxcOiPLnryOOHZHyGdW1LQrmXG1VYLEnloB
xk9p9my/bFbKLnww2Daw/i34PT4aLakczcVF5PB8Apz4m04mvWo+SCXE+rtk0JHi
GVnNC5//Zu8/d1CIgTs5C7WjFhUtuSi26ORkcfELQWA1YB7PLMMJQFNmhqaj7KuF
7whHMOlnyd9AQdWDVybUDXTIcRGQByZTHUarTpB8KR05/B89E1NoRueeJEV2U+Eg
s1INgZBy2yDH2vh1aQ7j7Y5t4SMws4AtJFumVEA/kGvTXPgxa+kkuUsxBa8zqmyy
8Ds/LkO7kRGhl8CypCsmOwVJoSF5zGHl11mTjqyPCms4qgj6ovm1uu+pMuFaSVb/
qzAkKdnTLM7F8XzBKE4xFOAYy4hSXx7007aBvJSD5XOhWL5CeVZbXktG6Q/tlRCg
vf3PWlqVmC0dafNvIPGdsgrg+lFd1+QS4MFfaa9f2zF+EuOEyCWDWN7QtYX6WFwT
5uYEPysZ0VPwJGQ84S/evIodn3s48+o7oQ7lOVdRP6ZYV2YtrPk8A/CQvmnQ6OtV
9oyips4ZFfRF6dtBub+BKLoHvFQITiRAGp+9wdm0RCGtAs+uaCY1X7M9UEEgyV5l
lrTpX80yYFhOznbQx708cT9Ff7EaliUqqyu1/8zGepV89Od8AZPHcYQd1uVj9fog
rFZwFnNmDJtrAuGqKFlu7I9XTHVj9LIWZBGnKtTd6veN7ygtqCzTXpIMlAi8t/Hd
/pTAEE64NEK9rCB3ZYjXRRw5X7dT4TVdI8MrvjOoLSvRpuZUdxTSYyl1Cp9jX8q2
ZxvW7paclSdf0dzbdXzg2i4eTi6qkmsDdPXesW4Biazq8o2tbQiqIcIbbsQLA08H
SLJ/AxFZ2Qste9enzLKQ5BphRXnC0gQbI7YFsqncHWHRXSfEA0o9zj21x65a1tHI
tvaR50JiPeKkFE6oqEftD8o0IGe1laW0QNZE7B3CT4nRiTU4nV/xLdAtv94PnHkR
muGIhUi5ycobG6ycTMwcCZaOmziWCxGR24sKUcDCUzCcqQadLHOme0uE0C4QG3dp
CjcALs30pPRXRUIbr8v4zu1fLdkpXtdXmOmhqC/z536ilVKBzJMvFHAfbgWPZoOT
AuGcQzJAx6SK4hQVk6jz5UBkb5Kej6HwKKGM4MGIEsNtMIS1VCheu4NblkqB3uzA
eKj0el9ORUEgKUgEqe+kFTjEplmXzNWniRU64FByII2uhrW0zvQK83hKDKJLCMRE
495iuWD9lfVYZqoZ48zujMGtE7S8sIR7hNmJzchTlRLlwbsWu7NQ0aWb+ZE2V/vh
4Yt59BFjJ+Uh0NaxUD1Vo8Cnfsjurk+IR5Gl0twEycs7GNaOh+f4I+2NbUzXihp0
LE/JSCl6DDuVK81QRIBoKjgSEHigRjLo0xQAAtZu82lF2zH7Dj1rA27ik4na+6bW
kyW/E/Vb8+K3yRDQMqH93Jz4tqOZpk1yd9C2WdExWarr81/zQUcgqYAFB7TzCyBb
Ut70RPIuTtugJdWzBUZ37aSYq2MKBHcjyJbPn9k0hDlwXpdyGtuJyx13BXRa4f4O
uetgxHXVIHCtcWJAjxZCVa0SWinoSK5L8E1Wf6f3oYsalvtcSbFPFp3tPMGkYAFN
KzWVVFGYn7yJxqqZXDI7eI8bkRD4+72Q3u595tg3IFHpbW0u45ArBBRCVxx+beY/
3bFFp3on9FacL6Ehx7f8gNSQN8KxQYo5v8K3b+VSTxheSrWHEoGPBCPDdctTzl/c
sf7ImqO+7z6UyRxYiohuzfotQfYjj6Eam+ko36sTzQ61ccm0D+XdATqd6hXycpa1
N93+AJ/r6NyWfPQVoPBRiGw7HGxdwdwXv7sNqn79bM4hcgc+BnOdBMDBg4WQpGiv
LnvIr4G3aXzgV2L7FYmuWqBIxUpDee8Fb/aZo4sdKEFrPIiFQel1v3ocrzUuhHzO
E0lGJ5vloUyPDS/pFYhBEmYyyprvTXA8MCdLtqh2mDW9BkQOGjkbHNr1kBucmvrC
xtMXV6mM/c0XS9VVy0WH258Y7oSDgl595EBRvdjtnYA+tNePyU/76ycO5y1eU29y
nTUslerUSPs8KyifqEfb0MHCelHbFJLzLPJ/ForFw0dmYKs/m0kPuBnN0Sp6of1F
C6b4M9K3n9gElmMAPYHzEVVc+Yq1A0FUv7ExuBizZhRTGoMG+VdvvhxAjE3NcVkc
2gjaBQC/H23/hr6PmTZJSwAqxtxdUCtE/Gj0tm9eANyZIfUj9wEuf779vn8DAHVP
oq05SvGom0XHPjYKRbze4sJcxWPXs5K+aYaacWqodcd+v1cRV+SXLbLKRfe0dHXB
4uMkfYzK7fPP11QaVdKxsaXSIiUd5K3ZTIkxAaRu1OO14cwlk1NTBlB7ssUNPzOR
4UyMHd3xRBOF4Xya48/cLGr4oT8S6e/Rs5wnruBaZ6ECwWjLeqfWjmscamslOM7Q
QPOO3OiWKymocWB1NrhYYfA5Ha5G3f2Z2Td8XQiIiG9SvkfJ2z2uzi78IzkFFF1+
NMnOeA2OYyeJg18TH/M6LCoMXKTVV7yjkrvS+/c9od1pOJ7+fTlZIy10NOqueJ3S
asKJSd2aQP8oqYRermCtVVaWLY6oH5xBSpAWz0gVHc21hpLjF+mxaqEU0/FiL2ej
VtS6Yku0yn4LfWyjYLwtYlcRy8Yai0caw/luywPPVwwIrmbkCS2jv6BUNAy4qNtO
J+Uissdo8xDKGka1WhtgyGCfIxH/iDSWi5EioTPErN95lXdgqCd8ysZaIlg1W1xQ
6LNlQSr23Z9JzJnx0z4VmkZUUkF0WP1SggYbJwGL1Ik+ujEE34yZkUS00fu3Yvm3
+asKdY2C1auUqYMQVtj7bzyjbU14fKHKXMykN7qbIposb1MC7IaLf0vaf3RUO4rN
atg8UQyF849pqm4zi/TMYVlpASJiiY+Y3wT1WyPWIsR66+XMpKv1xjalovrc0wg9
eaQWWyoXkAv7LyYXxcRlsR0A/bOHiYLK0xMoBY+hwenX61/2hDRbJaDGbn8HDhoN
phlva1TWm3qU2PGKHCUNljZkzX8zBqDsbJhOjFMxg3z0ALjuGgYjafQjpLGLGYwn
nh77mCqGpUDMIuFu0ouIablYyrgPUY8m3Di+rEXeexjl/ekoEpb0HN+Ohy2JJ62m
IDDGngPa9XVW/rIWnvjOUVoxFwGRjKVOoeHj4sS79Tzb9gWfqxt39UdMDz3zj9Ry
Eu0lICMjGRJUthN0hoaRW5gND7S0e/ewxxuYu0PrzrYj2EvYBOA5t/lk3/mIdFYj
uB8srbHDoQiYuh3Y7vXn8aK7LDG8aXV9YSEm6uqiLxFhyIYS1IbuUJ0Mjv9BJS6B
pDxIzODyx+HrtDccZ35Pakg3exxoZl7meEtF11ZJGVN2sVrOdViVCoxqbeuhnOg0
OPaP1pGOPDKnbP/V3yMsusdVWw4HQdfZ+QoRAwJVMaCEDc0PcRbfMC4CcqiBL0v6
sX0dlxHtULsuUeq7wcpGfFx/T+VQmSOagw59ri7hDIFv52DWJbkp7wOkA2/gkDJ1
9DYFBGHdrS7RXvk9JhqnXjhu1kL+Z77YNDka/TgfDvdkB6+XEOkpsRepQKmkCkBW
1yRF5gxgNuTe5JZtoLCSRlY2GdgT3QeZQBXgoRI9wEH55GeA+aLCerLniY1Dv2R0
5W8NGFd/i/zrv+SqB6Ik4RiY7OKdHSkI/JPRc6N5FBXnJ5QEEmev2sZGTbzUz5D6
Rr2w9h+VVDOaIzjFVdwOwTM6hNrr5xYph+X84wx2VAVq0mdhmybXSPI/kOJTkPCh
2hhAI2HLACtc/zh8KkfCny9KmsC6kR1PLQVCQVCCmDqmbTDu14gok3RnBR6Q2eBF
vZ39ZBseruXukhJTE73Wc9FUMz5CUMY5X4a8sHvNuaxEbAr6sdQIBWZKWUKN2luK
UJNhuzfzfCD3ontpswREr+I+tDVV7FNKa0nz3w/J1TA+YxpZhc4JpJjwFOWgGxFj
L0g8ouHUgJPfymwNZpk7tysp4KgHzbLJ+taPtp5vcMGSJnOWy9y6Jhijf4O8+6Kh
265jx+LDMGQUqsez0qiHWI39y7YR+xG/ijPNlJeSBsletmmJLZZuHMUkEs1r67tz
RGmyW34cazB6Rt2iQP9vln6jyHvnrghaFGpEM+XEu9KLBJuzZqzQ8iD/K9gQy0hG
as1kmTI6/iOfGweQif/wNr6PprgmqhcavF+T3PdeJlBkl9kUC3Xk6AI1rj4FoeKu
ECNWhVGi1tPsqi82Iob8zlWvrBp/rVjWps2T1cDB9DyGEkWpEbU0lHdHhpPUjOdE
LCPjJJdBxKu6KB1O2VlnEGL+NK7402AM9/kuO9nyTHp689Kw0qvImPeVT7QLZuxw
EmM42x67yi/MsdZsG3b0535sVSFtNxClVdItueJsWFuxwDq2uW0DLOF+iIoVCQcj
RfV2NxUHMHbXfiW9OXoSbVpdLS89XMX6qk+z91Oa9ny5gOF5D2q0a8Ra99YgoyAG
Mj1T/kmuJaIoQ+hsvxXanXXCBWFY4o1zeIIUPzNYQO3UBq5HZphrjizpdd/zzjqz
NFjHoReLZnd6CeR4MSWurftRa4VRuN9nuG7PJIIvdBDBdP5Fn4MPyP01Y/YVlt9+
`protect END_PROTECTED
