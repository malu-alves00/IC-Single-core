`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BNA5OTYao/jelNxyOXRTO1yhIgDwlFmq8xdXY8kEI0dFNr3lqouX5yLtlZC7+hz8
pHgBMzuqRjWjHXyOJB5cafwNudSyY3nYU/hw0E5il4INZOkrSwGsxR5/gosLpU/f
WVn5qIq9MSnWYKkB45fQ16QXEnWq6IrP2y2cB+Cz3Js9gY6p5RkJA/yooHX6CBzh
4TUAGL6gPreAovqMKhSGc7wMNT3wk5LSfWnxu65S3mNsxYjuJD0BxlZnMN/Fw0hy
2X7u479SM5GImC4rJbQdabHPVjtwcJj0NyREiM0nZSs2At1W1S1VnO7vEQmtscwv
Bn9CjDiwFE5b7MWdu7Lo714hcfUpoBOkQ5tLdc2+0u9Op4MtwS4w66l5JhcgdBlX
M4wlu0BpFUNmlQh8Ffvkdeu9OBrsGNq3CgzjmMCJwlqFWHFPJ9N8pKIE7TCoWuj0
3z43DO/uHvfu/Mp07X/lqSmu1jjrVNigim196fnHiPcw7FvRHQH3q4bCZbxSgp6y
IfQHRAn+gV9Dbu93M2/CPLDkncyWr5MCYule3FYNNA1Dzfv6VBPu09X8UZu/MntK
usvzodNG6kG+NiHXjfx4tfbWNQsVZD7xzpcxNkT6QiNrx+gNFAWkSZlDWLEvoa5Q
mXR1GxLMPBVFCuRD7N1hsDEHF/4c3HC6pwgQI45csfhX8ho4gmT2e0gP8Z7RdmBm
RiySgqjbVfiPWBMjH/1oPCC7SIDlMerRmoGaafkU6dC5N3OQeVjWqP6i4KMzLR+7
aCuRn/okcsqfBiIMnM0tvQ==
`protect END_PROTECTED
