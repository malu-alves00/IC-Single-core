`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
e3lkFJHeTaUMynzXhyj7D8AxXJ5PoMk547CZFf3L4piheXK1+ILmAzL/UN2XcA8v
jwNrXEXtBW1s8A20EL/UdlPj4S9Ui5M+JD3eJQp/A7NmxbPD5VGJ+AoFivDpvGTy
XCY4nbCmEMbXYX1MydJgh+o/jjNRPGKYWa+PBplpB5a0STJVXYwuNZPTtXxmeIde
bYaEj5/aaGwCdgB/rjbaqQALTWaEf3xpygTyOZhl50W0kMPTwdKxS8Yah1D13Zph
WVI37kjqOZsC/l9CI3IANqAHyk7eaJgn9ziSYrRIJ25yi6zGmHCPnmjUsSGpwuaa
8jANE7f8JMNXVEjOvSfL1eh6B61U2Y/K3DMFeXCLx3WhKgYJ2ZikZR+jrJVuD7Nz
42rkbNrNWyeCbjBtDacLjeR6tEZKYUBuK/QxyfGVLu+e7wuENzQFcE+sbd9XeKml
xQ2tjE6DsXyetpO9/8d6omzheSU3vL+/5lBLsfi2I/NVdD6zMUdgduXdiLb404hS
XcqwIzS5IvofUKADEVek6Ng9caExW9xdHrtzJsxWoC3JqEy8mqVNYYVHbW3jxNrL
tPV6mD1Ytq8rduaHQF4sbt70q18341JabFsVRg8s3i1E6aFejebODOF7K1sGb9G/
Nm1jgYNn71gv28yICfsgynq0RR/v2Jh6xr+w1QqY/6wanNtMM3PD9uKFNQ1F1iQY
Ox9vCLW5T8t0WL+OBAsIIjb6Cqrz4Jh5vdPQ8rleLbpwFPiAJaQXs8vRv6/AeJtF
/m+vJrhO0RQ1QIbq3qguO6kg+BxCUBGFHQtem/Kn/52PuWs4+Y/t6cnDrxzR54nt
OkmkIIKPokfbAB+ZIvbarhhG44mBrge9oc78+rHDtnkMItZtCDhePcVBo/W6w0Yg
eG6wPlj7OLW1XQRrm+hTfzFmnGRphCxGhGkra4Ry8ag0iKA3ApoTfOxbAGzHOaSr
qQTSNax5UIgfsKhHcDVxB93NtDVllV0Wk9Ym2lp9airCxBCFbjHKKrjjz0324heY
qFqrxeRXM9DbQOJBwvGfvCLxt/t4lsXP9hYWosMOTNn+t5UFeUMW8NYn4BGGth4l
SUrm0HN66i0g57vRkLrBowQfvdb7tGUtq1ook8XrRERyTqZUYyOzwTCeIMPTFDLP
vv5ktZGPSFkWSmk1Qo39bkP6eOWFYAyGAu58TnSWrNp2kZ93HSxj22qwrBzns+vO
ZHOFiYT0SK0SnTs7nI1Udq9081hQ2Fpgm/Lws52V1noiIsvJECnhd5RC90kMKYrz
C81euz3EFaU7i+2+QdN3CcswGc7pY/VKZIYKx/ys0W495xkelEsrjdLWTq2uOOEP
P1AQKONGQSCZ6Jyw/YU67nqp2rUs9uqmvZq89PkgfQXyls9wuvRKcfPGe9Mf2ie9
tyU+6jtSA31lQNavPMu163yNdpl6PAPzGqCYtbmv/+HI5WcmOjXbJJmKDYweCkfL
s1Nj0j7IWgDBW8y+xiJVN40qqOTRgUtD21hVSirhg5Y=
`protect END_PROTECTED
