`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QGMTZI44F0wRwWKSo5QMUN03v5ZT5lrmsNTLFrEsCZ+nC+XFY84/Sd1HyjTLyhsE
Zf4x7qci4l/6bHaPARSPrpvJ/cEcM8hIRKRUWbp8Ca3ZfXRFU6L7CNpNoFH0KeLn
17sYZpbSe4Xan/WgiioTvEN2ja7hfFCO5C+zoCEb3LY0ONzM5w+Ww9bF/RPs4z3U
p8qhlaibOPs2uMzSbexvokT0hiVFkoo7QtNUw8g5xhgQ1S0AM7AVKRvx9JroBSeb
zC01TFMBY6fBSVlvY40sHKV3UV4Umy51KgGGTyiGOvnxcLvRMo9VpOs9ucyYFcqD
l6xUg6GEZ7uliSDN/tHQLJtHZ+1Yy+Wv4OgCXFN9XWQqQu97K6pr38C2PwyNCS/+
r14xZ3sx6NKsSMLMvFBlsxAevh3TWbsQh+lcOR4e9ND3KY4xoBo/Ub7tWWH3MxTT
dRQbArcLWOHAoZrbzpmHuEVTJSvEFp09MpYEG44WXsQ9E+nISniHFzlbC6PKChRV
YOx43cf7nXtvjXJPWO0HUwsMknyiRMUZ9EhovJW3DphvnUJyimoHzFH2ln1fKuYj
K8DJDm/hoq3Zp2ScxFfq3g==
`protect END_PROTECTED
