`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ql+NvCwQPX1qPlQ3LLQjQ/PPJyCtQ5SRcqRgEHicQ9jygolik6Jy3aiDA1dMAp9B
aHdT9oYIxnikVDPTekwHOs4SI6kRjlrbC4NEYYxI80tFGJJBru0rC9PDHuFMP+ab
j0zIMrVQDA5bVKmoYJvM2jBcHCS0XzaChHs80ds1jHOM7gj1aAwR3W1UwSdHOWoC
ywmOKHQOd++DKjKHGwAJR7fyKwE8KV7POyiqo7fJkfnCtD707OieEnHww92znv34
F52ygIWXxtHQOj5axRFgEeT21ysvPYhUvbPynvgG9CWN5rbQOKmJ6qByPREYB0o4
3BUAWItAATJ6BVEA8GEviDYHViPOyekIBq5DXvcgCCOxy26sil4sf7rRZpTskqbx
XR8hCXqQkhrGS2tFibXm4sKBey5nY9QTBrwr7XTk6uOULMwz6hD6QTnDweKVYHyQ
VQtM3dtJrQ0J+LzODWhrWZIwB9BDMca5txq8bder/dyayhD4dwuFKXOsn684v5rQ
aZ2j7f8qtYIH6GZdfEi/JMw7LsSEUrShCIHIF3O7CXeGGswtJhLnSxPiOjYEiK4V
84aT3ltnJca42lziuYtvsWU28ScIzylpkPZ/AaMeiOSR2Xuz6BIYk4TFB9abha6i
HYaQ8F9z8rQSCX9DKYZZ/FfH1m5MSGrkgPyfeE50ndwymwiABYR7rrW7mjoBNmKw
4eFpCqxO6/tGyF/1UC/Naahk0K/ZEKefV9RKArUFoS1rDPZAuNWukA1sqAArB2jT
HOwINS2HLDWtWJm9CrX6YC0rrzRpMw+TMrjw3nRgHgLGuUuvpaTx7AlcJbsG5mpF
7mDTYn3QJCkGQWQqW6bCFUtv6CtwDklyLNjb6bI83rAj6Z9/CayK2O1Lb3SqBRVZ
e16b4HswTREhZIqt5vd7gbJlaW0/RhUCjPq/BNPK7VpvsXTkITMxS8cj25W8r0PS
iBKvk7GUYQyS0FzHzDXo6As5L6IKMkVQy1stmpU9u4ICm/rdf5cFg7GCU2nYcHtq
KbjuaW9m1Ps6cHgAH/1t6pTW3v1FumfSe58vAasZE6rdrFcuxnSfGqhl3R2OEI12
7/wkzKBtEQynr9zT1XS2OFFGH98oz87JWrC8TMWvHJx1R9iBcetstAdU6HYgTnKQ
EhIa6BM4ogbdFpnsvqj88bkaM0wavnmteZpIbOpY3bNqcmknnB9aWnTxak5jg5P2
dR9/5q3lnEpU7RqMGhn7JKLCL9HA3XwMsMBCEapysj2nIkFc6SL9nwJMptgN+3P6
rR78wM+DX5ktb08XCcSHYaBpquAC8FPndacBMCWtRIGpxfboxEAWk63EJJWs2fzP
MGsmZt1LQ+SjboXSU1ivR2gqTY6s+ktYKdJpNBq7kA06kSGUVYy0YKL/TCDMXoua
OBYuWeX7NAPvS9Ed0/9v5vwJM+lJ7+vUBp8hmXwgHQIXQyKh1uIJk9wF6jT4gF8t
jgVy6i9E6qLL+3FPNrk55gXLHfaJcSbVdxaccnaTkTm5s7JDLA7JTKm3ZnyciTWJ
K353TpirYmD4/vAZE63gOE5IR6YUuyAW3Q9IR9qfEToXpdEECDPuFnQ7tHG2z9Sm
9Qv5qtlpOOrsOSY6mVubaCr+le/PvM2J1XcSxwjPSQTl3r7EtXMRHnO6SHp+RHFK
VwDnHgKs5QXfPDZPqBoTgoQw1VIf9adj6XpGvqeG18buCq6cr3AHtbqm/r2AkxVW
mq8n7BeqED7KAH7T1Jtrr6bKAhcMiIb7a8oeDMoDhqRjr6+a1v665xzYn1Wwe/Yj
8dnocx5/5Ed76abUZWX1X5qPMUuhuki1jLU8x7icDhJRU4cWLamXv9AX4cS43qa6
Ch2S3xEJm563rP56kMnNR93wzPQCCbeqyiXqf5HBQI8Zys6HptjAHtC8mLQ08eqz
ShgjPZMhDHqNiY/rCx4FfHZrbeFDSzQsX9T7HFUT15GVsAHtsmBbmToV9z2bC9OX
pCJjp+HxuxbXzK/V0EpYNTF1b4xlCbHBliqwLOEzUgIfdpqEc5poOALmmnagMHOY
VUwUTVXy85f8xc/iNiRWtnoyZw3A038MA0Wo+H1YrhrZjsROsvoRrtNYtZZ/bJfv
CxA6FsO1/W488qrUfaRGezb98+P1KuUKiG7iCiDXU+h4UEpPOxR4v1mZz43hXcaK
jRHNbAVMakhprVNeMPnwAoTHRCtgCmFz6MzSl5F7fwuX9GXbax+W/LZuMBnrYvTr
xyKpasBFF8WAgFF/QmMhXHeinl7lzDRhcayfjXKmay9hOE9JZJL2O2BYl12QN7b2
JgoPXd96oeySBiUIfYBbBjFM6S1S+c+ICefGAt5xsyz6dWlfifv5+EosSyO/mF/y
eBSsDPdN9kdx+yhSR6+PZ8CgcN5PsF1YewEvbuoirlxRoLsnjloTam+ddWOPta8T
lGYp59A/qJqOjF3FZ/gonuJKLRWAmxQ0x2rWPn4TOKT81fj3ubjaj8HjvPW2zzI2
AMO/CEd71ddq/BxuUvnCeBCoAAv7j6gsEGQbV2HR+YD/EmDYqZquPZU/lgaALxZo
NgH5NgHo2/pO5nyNZY3oDuHrtgPXfLpRnrqx4kaEkGt0JXwu7bznGbXanwSA3mgE
xz/z7/DUiBWOJbIheSuVxq/uiejyyVCp38YW7G5DnMQ=
`protect END_PROTECTED
