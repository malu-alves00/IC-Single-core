`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6WHgTGIdkLvufjTT692ITykK1wXjn+JiE61KIuxZrlRWh8nxGlN8PI/ltvk8PQFN
S9Ohb5wjMoePl6g18m4O+ZzhZI/1qTZUQdUk8Mxh9WIfSA7gUFlwZROp72fLbbHT
+8TeCZ3r/R0hc5SYSZbBhAJEgT66KzKgdUd0SiJ1RC2uCSEsgxrqDlFy54OJuCHC
WM8b9TURcToSStxlaBy5PcjNUaAZYiSjNsh0hoj8fe3WYrDE0JURvk7bw8spkZti
gIa/i4Ho3RMtHWUB/BG+rUIinz7TeHS6rbWV61sZ0X0wvvbCVgDsUQCu+cKd/e4j
dHKfZDxz6wmowiy6TW0/yfHDD5G3lmxMO02WcSapjFUaTX70lv1w/KFbbk1GnV0O
qrlJvmHh5y3L5rPD/EEkpn32O2bKmC60QaEREBWb0MOlQITQMqX0ecsWtcWoR3cG
dLVctZDP1+tMf57QoEhYHh8CkUn1cbE/3pMmU9K/86oWXnUe+Hnj1TqHoJdUYSnU
tYSgpASc7V7nWw32PQ+jZEOc9hgWIsPhl9gWN4x9YYIGmLYmZy/S4AMCsM0gJBgh
7ymVENX1LKemSrMfpuzAhdIMvCcB+B1qknqKBwxp4WHL6636e4Ar2HwjOjEPJREi
uWBt3hsSMYxZbghA4f7UO0cKx/bcx/l5jpZ9NurTgRtJiU6sMbqqDKnvuT1FWkz9
rBIVDUkZIFpuVVlLd0BQv8T331/MVMDnGHgasWQ1vSglnMBoxWsiGBjghkTubIzs
Cff45pAON+Ed8iTS86LwqnSxxzAnYmlmh2Qbl705MWb9cTFPwgosFd2qS4EGib5e
mzqzqbrRuYIphcS9G5BBtk6T6K4iX+/jg2D5CsQuMec83XhIb8fIcZ2YID4U/qt8
h8UwUvPAS4emi38VCttJ/66S32BOQGndd9TGXhjblyw/4HSNCv0qgflGN2VOk2K2
Qr6x4yoUk+XpZhdpmPcA1Lm1g/D+NutAN/VL7RcJxpSaWBS7Wz34VBEtpj+RMNZG
yDlMZzOst4ivcpNRLXzfCH6GVynuYEBKjdyRIEXEwLeb7xJ9nHAirBf2NHUq6A9C
4B/G8pQy0rjJTt7MkxW6YGzhtpw4XI6CDG27w4zUs/btlxiBR2ElQoRdEFb0uXyw
YhSQNDwRHfZSxy33sR9yLK5vmkbrucCWYBtAh3At5Bp0qK2pzwgZQbFz1nBZSopP
7bM6VkBZBHttMgDpBaGuvVO+y+SHRlI2CwkLOHxvrnpHQ20Wgz8LHxgXlx+a9ZMM
JrKsYFUHNXorLVqjHDHxIihVxCibZXETOGPNbP9VR0pJEve9wmz6s6yEyFtPNL6G
nUhn5KV48xuWjfYAdfxTiys1e9VPHvVuWyAddgTj440ISyCbK4l9egy2mXParzKb
6p1XCe7OLHKWyUwCC8/DmW3U4zAOq3xpSdgZ8NP/O8EYUyYtI0VmNr6b02erZohv
7AI1nMIc2dS8KeYL9rdeUfsD7GgtA/5x+SmRIfGs4ZLtVowlJtXY0ewLBXv/xHF9
8Q1fHqLZQV+iu7Sq35f7nkT0qehQptOGT/jddictq+sFXxxi0n7mgQPPbQJaxUo7
LZy/3n7JAwcbOf/t3AxC/xjhAeRwPE/VKQrjbcexnB2U3zRofSpFTXKe0riWonuk
68tSws9gAu+doyDy9mAdcd8cCxQdHMWDH/E1piAUqFnGH22S9TTPgS8IURvndcx3
UTtpd8etMbCRITrNNh42vGWg2cZ7aFx+YyZpVhG5pIcevrmr0+TqMvysW9S0OU4t
SCBU1iynVoCUQAiYN78Zy97Rh491a0hddf2FhqmxM4iJho9OHDkVzMGy+hzLU9eL
xtWSKtIu0aHUtElws5goHpnY69Bk7lGVTq5t/5+yW/7kI5nZt8/2cvAjoC448+3y
pynPd7EV3AtmPngU2OZx/zgDz8VR3VzzzdMtt2wa4zO1CQIkH4E0AZDh6amL82oc
uvbSVRdmXXC97BZJXFch68284vpppKCCSgp4Z5/0mQ8HapfS6ZDfYicM4NoFZvms
ed80LNRJSqIwmicu40blbP3MvNftOPS7U1aCN2bsEAUg840t12Y/ejCeI/VjGsPv
pqHsw9jPwARCyjKShBujVbKlxxNACU7FGJ0Hb1TtlBRrQZPCoCu80gBADoxLpcWL
ykSI9o1cttnGrZ0oeh2/4wn255zUWsCLyZpImwHbEVOheBgZJV5Y5OpNz85vg05c
FQFB86mYJH+L7ZL93veMpMf5bJ7jCBhpW5Mc7+qujD2ucpT+eMTkOc2SimrfqEk5
ZYm7vAqNG+7KHBtBIoN06uaowjVxVdWQjJqFy3Xxk3S+pzmVajZ5fZpa5KyrFrS7
HPMGzgocHzzIESAG47zQEhO2rBM9RhmkkJ4jwDehyp/9wj8cFtg1h/6d/NzNanUG
TqYuIYfFgg6G7yt5r4yzxRs5xRT3BBjJg4zZ1Y5S1NhzRU8/PQcI0UN3/n+XUauw
QF5nzEu7xkrgw5Pzwz6Xyyy034tZ3zLwrSP2WXixDt4jRqiBezlKXkpFKZ2GNeBo
7g51U3pmEzvh5MGcPJ8EszrAIV/a583nkygDtF+rJ3AGvNlc7P/o9ul1DBGFbI/u
o/Nfs63Yn1o8Ej2IEQiy9cR3nVjR1f11SfGQQSTDtHaMoYN0M5u/iV4Hh9IW45yk
/3+5cUM2R7tquluT8sBZicUibDiUWUfxW9L+2yqqyFuiW0yV9fNzIrSmMQrAxG4y
5IAGLH26AdcSASrCbG+Gz8c77drnp8lmIm5O6gKSVOGRMMgZgo/q93fljfGelf/O
N9969/PctbkkUhJ9UEefoqIqhxGyMRiMfHrzQU8GttNQgrMkyTPYq0UU2hhSNQp/
h/VZSHGS1yf0obhiTYgkytHRyFUWohGpXjwpJeA5PszW97jmDtw/eFLoD8tnM5bD
9q+u9yDPs30PWInpQlEHuRf67UM9/RO4pHW1/oe+gPjjioVL/tym6Qp5ZAudqn50
CpaVyNOtemqUuG7kTZSXYb0kaLrrBfG5hC9M9p9yH6iqsPAwbKuOuLrY7T4fSGUR
CMu/bBWJLPS9aHEyeIy9tbCx8XULHMi2OJAZtuHY1J5yM2zo/B9m2im8oH3j+B8T
Q4AlvcboSQHRcwm4VpzMHbFsG4eWUYb+wP/cyYpoud3ui3/+dqTisZtTGSluNxbf
TFuhboHifq/JkE7dGFepkXqIssoa3gB5Ob+Swgt8tKIIiNXsB7dLIgQQE6tvvlfP
YonatL2JlZhDAZKMJANIS2BttLrprotKNeEhe9Pl3+yK3CNZlfZsBimSU5EtlEcC
Li+Y9b5lWTeGQLinE0DOc6EsLEzjS1kzDjSFaEGpsOErKBfyRZiNqTHH1MgoaccC
o1L7u/CB7fS7g0nBto4UjsWm6+CLy4VvRX+qYe18Zzk7a3Vw8rOhoH7RZMh+wCIh
qaM7nRhC+iCw1yV29foxuNZSbUInwk0YbH0dmwAtzjtdORi7ObbbVUj1hOX6MRMG
XLgYWCwD3kERycUUUFIfj1BnO6rv7lxeBjKecQsXTohWwFzsLiyIMU7btErdzRfs
GFUThqKDClYrW+PsKRznOD57NVfb3tUvna4POeo/MGccf9IO1b7gEZyiVoSzOhCR
3vJVQMynxuBkmZfh935/vtykPejdPgtwz1MiqzWqDYoQ4JR0NmWntlS39g3+NEAg
muRiX+/O5YTBDXHHV04xUiIi8sQhKHQLUsRGkuYDeUK/vmWmB8Q1Afaab9LgfdQ5
rXiAieoEcOeHPmxT3QoCtaiVCLp/qsKJzlrYAyHHos1WDD/6EK/DMHILnQslhU6i
lW4fxjajtb4gj6NNchMB1BM/N05nyLo5re9AcW+N/WNkF4POZ6Q3tfRRuQNH/6lr
NXWlAl+O4cQA7fY+7pqI9MMlgvqqGxepjnEDCZc7q360XwtngY4UL/lO9vBjQnQH
40chGLGhBQ+20ptVcMYqyLi+ZMjpogjyVz0OWwepM8ZURFBNffPsDSO+oF/ET/mZ
Y+DegGB6PafYzAn8jlNdv7N/NEt72G4aZUUSeDjMrvv18+q4F5pM31+eEy+mJGEZ
fz7Ay8N5pKWth/v1bpPiUh2XoWJlkQhGpCYlqowTVV+WgTd0y2VtRWCnJtCfnVG4
ZM08GWTdtfA/vqK2+EAr88qFGdG0wdZLjgJJ5TREAgJ1OfK5HC0LcDXImNOsDWTS
eneWliFT0qRj9Ex0g/5YqnZGQ5JfMuzh5gqDnmbexuPous1RRXozfmC3veIndPY/
xn36DnINOB8my7CBnasBy283bl16+tOEybkbQZEbCfQ28hyQekeQbI1eVjGPZQrG
3s9VSIArxhPlzMXSRVfxFzmUFAKuFWT5wOUo/mLveXDsihJg4cPww3jueajyqQAn
cNw35LKSj5SQBj4ulN2iWnEfaUeQSE647rpMV6s/JbOFPSxVH5tcKpkE4RNyNaVP
7XecvtZYY+esD/l4nUiSJz0QATht0MweqeUZCdL55m7hrvUzd7hrBO6OiFuK05BO
J8oBucbgWCQGoafldM0RK6WcE9pgjWl8vpjG5l+BD/yUn7UDu1Gtj1meCAllPQ/m
TkZXUHXVrxaCJfgyi/Z7F4Qu5Xm86pgRONbOQXnFKpCOvU7/ftDWutJ3bUuL0Bqu
JZuwvOs9c4+3AJZDIGzX0NeenFafojQATxrSFEB8D7aBLLpcJQdc1K7x+7g2eL/8
HrAfs76yNFgDkRjJhjbjWAlTaQ3Ammee+IazNRckA6gDPEhrsq0ii/YchALDJaHm
8IQMI93TtJwqD38HrrM4E2rMQ8Sq4tz/UofFu7us4TNAdf7X9+ZgM7C8NyB3WUps
A7mMVpRv2h08HkWgkYjpFKBApbIo1xLsZZRXApN1D/QKMA7jztrY0hY9vDsLuMQ4
9FZxZC+W3UL/H3P6TgPPegro4iZ9vLBXmxb32nWhkBzNa4JYXEqP29Mo/Cch27yy
E547S72zKu6ldTkYPZR77BG9eOt/Tb6+ovjprXD/BYK2HeI4jf2Bb4O6ANvJQQTx
vAXEdIeTNJP9s9F2zVygSk2Njodg8tQAOaXQFjZE5yWg9Y++gZSxJIgeXT6qelyW
UnsgwxmesMrRFmYHCj22M1xBv0H7aq9Sn2eFve92p3N1iUolQMPlccEx/YihDVVC
IGwGxVe0PkTR97QX7O7YHUfpUeuNo4nVpJNEOhQetJZZK3Bq8yyHXhhnttAmlhwS
+6VjkO/kmtdPM7CY1VZWohVGNVCPw70G34THDXaG/P1exEe5TEFV9WSuV4CbmOgR
zqPwdz86og7UXdJVePgfPU0myY8LT+jaHneCIpxp/VjSPSQEPLanK95gfKL73eSw
GrJi/+hSTSbnKP+H07MTFEFbnsTcAZ/LQR1Kqjto4goaWQ/WPKs4OXUBJcpF+EPc
yvmz6IOdnxl1YS/lJBj7gHjDwF9bkYsWpEounrJmjTu4/5aR+ju2VbMbrbb/mbYT
DqJ57pC5neEhMn+Oz0MLeARJDJW96foRuSHjNPbw06fwY4e2+HPhzgIf3jJruFtW
GWvMR2yl+vVdzNf+uLLnDsqRUwtSs2dWmg2nSqBIC2g1C1d279/iewWeWPKAS8FC
KXHXi5ZcUVxMsAVXTLbzY9clJdCLW+CFN+vMVIZYBruuKsq1No7T5HuS7UTjGf4x
YOXFqf4yUkOI9XwvaTpSeoiURhROFbaFwJU+OURoSKF/l9A0WG4XO5o2UScLqmJW
vis8aJGj4lqu4CdJckVe21C/wY4/dfxK4VjG5TZrpLGd9/wF1mmUmywmWynz/da/
OHQABlQwaRQ1w1hn8KkkgaKTXmwNzBtiljgg2uVs2KxZqbU69wbdz6KGcSrb2qpB
sJ+jyObm+u3VwXTYhgHIRB18UmlCXeVzqBLXIwsS/DOBCW3okc3OkmEAF/t1WsK/
muKZuGxFF3yyI2nef73Jmxvsk0IgqOkw6jdT+rq+G1HKmc/+P/EYnUO/aRG18AFa
dFEfUpZvHq5Ht1HaLUxuz7mnFQrgVOVD5CP104efNBWPbehzQEhHU1uQ5b7pvx/Y
mj8b3qh4tO/QSwEV5pM0evwEK+QXNI1BFoEMpl7/16z8miQ6wIhivKRoRUm4lvMC
uT6wy430gPvmLOqW8g6kZBr4aE5VHwrgUT2HKUjX5g2JThagjNp7NL124cRB3tL9
73EiZxRCpBm8AF5pgf0WNc+1WMKkz188+sb9LlRJGHqhbR8ujMwy1pPqg+FKqJAS
P2dqzZxbiUmoyarVchqO0z3AGROmTcqV+ugieXG7t39vg1lpDvj3fLy5cOuer9H9
5SWjruAFdXW66QPG8+Q7XtTZnJJQy7eYLnMeu1l5SSN2K2yYvpu3VwTSI4rfy/JX
C0Tc+1v30jHTP+1/8eemHC5nEOZ4VffJkDQHA2YFYDwXNYz4jDtfKdLfcq/6ipCN
aSnIvjcw7Qq/Qgad1OAa7W77G+odZYlxuhnq8zL+tsOt9mXFjiBW5I6FIls5FnkJ
WFxxnDuiSEfcwO5ji371wV1rWb0O1LFmqOeAtfberde9EtQOjfVBPHWxG7OFLOLu
567WLCMa4m3cttcVoVr5J04hnV9pIb8gXSruDf4pCd7erwyh4uCo6CyMEYzz3lha
TXDkEppJj96gN2/vE0zDWUSf1nHcxuWSeyMOL30qpxLAUtlrwHChn8Pdj5YVnfVk
ERdVh2nXOWMVkTL96RrHPD8a2Ij3ncNG9uUJQ1y9sTh3AeMW0/oeIQlsG2AJ1WXJ
01d9Wuo0tSQq3iMFk9jGzbDN5Bg9yS/kaF6gSoZ3IEJ1EcyGoK7yL/+6jojb3iG+
tRBONL9R/EF/0nyayaffvx+GRpNGgnpt12UDBI0u30+gvBqQT8cEun6BpQzYVCkA
dEQjrF75r7cC5+Y+XcoojVltp5VzzuAC7oCBKr2GKdzIaGTnT9/pxF2ABkBKcspX
N/3Wl3nMq8ZI2ZidQls/2spJ7gd8yL7iS5LmKSvCZfH6qrsKQqYjIXIKYcF39Or3
goyZzX37TpVBQXxSf0lVgDFwBvuf4Q2V9LHayCAEmSd0F3ja0PEksoL++erYuVPc
pUh2Q64iUVDIwmtIA8MKN4CoEZmJC/84FHA0fZyTX3WnCter/hVVLH5IEWToCxmm
ZIK8+XK9HH8u5eQFyecUG3sOBxfGM94S24YKFqVKvSDaA67gKxGLhrnXSdAkf53f
HP/6eKKfzZIpC1lnD2cRILhrXPFDinUw+SmiRCIHStDBSD6CDRFVk8R6L7DDK+BI
UN9OSxTxW9sNyyhvRxfeiuqKHFTbbwktsFfelnTe/Z4sFiqlke5ZYLnSpKBUPaVW
ke2Jp6kmz/9sF/dZGuPBO0cYIMK+LQ+UZ2ebL1RDGiQf26+WpmhGuCkk2MzLuQFQ
9HR6At0XVNLAXxMmJkBgD80w/e6/VGeqfCd+D+2slmwklT4ZQ5a/1XQB+8MlkW9o
pdKBOks9pE4SPqBw/gCtHserhOHl6ZI64A5/ivPVZt8uZuTd6d2HHRtI6qUvV04u
eKYhwQ+ul/dvPOXaca0Y5w==
`protect END_PROTECTED
