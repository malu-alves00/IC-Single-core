`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8yD5a/X87MvKMU5Eq2yJ5MmTuVhVguTwJlc8tGCUdhR7bGcBwGAASbDBWKFfqgMn
iKM25CQCWs055MPzwPmD5XEh0thLmFbtE1Ec+6fUYchxuKaCZ5BBAxbqLqktlLeK
RXbZFOq1wWl3FuPbpVY/4nS9LBIMTLpwW/xC10BHileLv2C0mJmX0jViJdHI1CPP
qXdGzAmcoBu3UG45LRbqkw0akrmxBrCRwM2mXbuGqtKCr6SMrzY7S4PvefjSNmtZ
ksjEd0VEiUOgSp5PtgGuTsomFvdylZqgMjNXha81bzka6yyzTd0YQnMlSIGae7Te
J2IAqe3QH0AbxgnJ8qQa0RzIX33rRnxLAHhlzx5uHtG2NhsS2ATWg6V8BylC4ZtU
5yA4dVBbqvWZ756RdfmuHGAaJ0YA9jHQMoqEOrIVOAHn3bgb0aIoRT9Wpvl0f2He
6WZekEf/0bMYP13zO78Sc5JjT+1OU3ETjj5y5pgFYbh2DqOj+VstlzODTGsXX84m
qYwDx4WdjUUIqlGW58ygz5n8p/dbsC7lDmuBq8mXw8hyOe6tHidytqvhXzAmUnnE
p2U4nw1z7/C/FLobp+s3gF1XKwnpXmcrkAO2FILsTn9My4CkVHfydfEcxBDHC4dv
zudp4UHGeDMxbRzk3+wh3e9+zc6Jydt+k2ooelT772KFUkvxuoJ6ZcRM6B/G+Yes
0FD9Ki8trrGxCzCLCny5zSmi9KQxfG0g4x+ztObdRohCVavwcGK0lBzNgiWl+KvT
g3tf1h/Bce2S6OcbIwpaL3UaurIgsN+HxxfcwkdQ/9zeOeABPWxWA89vyQLYfwro
bCDoJX78xaS8+2l+vpufvw==
`protect END_PROTECTED
