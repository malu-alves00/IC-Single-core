`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Jlyg9LJua57/TTWh2VhyWUz2v8VDeqFkHGb0Ds0/Pchpa80qPWTYVOItj7sdBMi1
VqdeHaYMTl/779pMmTwnEsWNsH1v3sebmFBlQ/5bPV/ceULG6owRNuEyfMAKluUd
TFUOqES4x2ITVAS3PgsaE29K4uxlZd3wKZgu/09VqhCaErCf0JtqNgGsx4vAzgUS
v9ZX3R0sAppiFXt8pwlFdoRCxqxyoUDkT8OsYzOQxKMZ5oyQ1SxZLuQrobO24trU
xoODbKHhjTtzVin2CYbIYiSihtvO0mzO7A2wACo3PmJtLw3M2aC2C5AE83Xb7NnQ
cv/0SgrCXxSEcsXMqir4aa4WovvDxJYBlo+LN9noFub5IyP7jqBLjhUEp0PkJOeE
PQFuKd48yz+wRgaUpcm14T59/ApiAUJzXImUAiBpQsDcV+w5VuBrcovaIFdqtmM0
Q9QTUC0UZTOwYJMude25L3pVFXXylImzAYJED6M3TeGUiN6/VSrh2g26vI7ZHyqp
EWidxnOv3WO02SvAVLxm2nmYrSQEnZ0ghxJTKAfdpuuYh2FD3MlNXfJTuEIAKJZD
hhtHLhWlPinVUfpRsPuximaHqPOLFMciKPEGMzrBW2cNGzW6lkSymA4kDa/JkAaN
LygiPIlj1kVlOoHnzz8VpqRqYtyxeomSN3rfBx/q0mndgf4oUa8K9Jn4QO0Wj0Fw
Uw/YXbWxcCbpIn9y6WCw0O1iANXSECC/3wot5F8PCxynJjQSvIoaG967hunvd5Hn
Ymu1L3d1sEE+cUiHWUiyVbtgS4uLdo4U0spx9RCySHyNsscFsYhsFSmLN4p4c7jS
vkNmCMGb1EyLp0SYrufsBTp8P8HvE67ha5hB5h1UWrYf02rP5HfZtGNItOA1Q3Ca
ZGG2UMZE0PaMUsG6r2+/0jKisYhEwxiRF+crZWwNPKvX2aGJg4eOhf16iVWqVg9J
CA2RtbGjD6WJCIOcZ2TQDnJxbv8rgPJI1X3f21JpGU8exU1RqD0dyf5zBxRcQYRn
Rtk9o9wrtiFvixAFRKf0ffCfMLR2ZoRtRhc5kfd49XxQrK27Pl7kTs/stv9yPKyw
DQHEcq0VtB66qI8C2YZtJVidZ/qW8Dr8yE7IqBiZd1/exq2cFJqy4CQJ/B3qMUdZ
D2miHcxrk++C2rf+VLqKCjb6ENTJbE7sKk7LTKTy42clwxGpg5/fOGzX9NupO1RO
Im4V2KzbK5X3iQCmqCEAeuRr1wkMVhiIRtV8l3mFd6rMua35MIyXsQRaPPfM61V0
RXCLbX49+V/vtrJYdzeycygOnmJTzodbJcy6R/EGP5URSspqPLR+c7LE6Sj9UJ5R
3FKbvXtRGfLkrNSvfRqvx/00LdgTy+L3MHZpB9tz32/qWoy+GpME7i42xMupo+tV
fGsuCvt/48+KAM2yRBFre1k5PmNiyvqALY97OcG51UlqmoVRrQNnK50ztUYi9UKs
kNmu+rrTj6e9ImL/zIoWFV64+rytceLV/eEpX40e81TgKi3hcJJkowysdJo0wpTT
16em02Ua+6EAt7i+b+ae3sZyk6tVJp0HOnPflpvOfPXCJ0JUPaHvLG29UuM+h/uS
/7HoUacN/B0YN8HE/zMUc9KIVIl4TUiWFZPkiu3yVm8dZq0pw1CPUkOzad35gXrY
Na53bJMeEpYXaUjuAeNiEgoG70zH2IGVdMDt+5NwAyXt9lUVUK64NbiuVPL6AUkX
BWKLmEFMy6peUsY4+4UcIDA80wL4gJgJEBE13lQgSPjljY3TvE/PHmvJSqtY2cH8
QHoLLlIymYcHDpW3FeZNnPfe6GlPNfQZ9fepcSC7eyoOD0sfPKKg9ARhvDr5a480
SZJ9DIHlh9W67SdiQ4bADbD0lt0UM//FwMQ5NwEr8m4egK6JgYKNFIwM2aM5SFYH
i8yCRN2UGg2GPfd6RE9RMN9+/EXpYwdUq5sUIcCYiS2FLbu1WPmOEmsPGO7BmGY6
2l38VT1h3NJ7xWwBV9CgIcDHgDoIXMKB40FZQ32KLRvuxypCfPEa/ZLLZuePRPqy
R3zyDkJ6Ro2xiyeXhXSGR/khDoZx7cztgLv4t4bgL5+INEoCEETPVUy84mTI0XSK
97eUMHycU0oVNUNtrlGzlFYQGjQBSvNYWdR2gVLecJ730jnPjWHkvod7QmV+7AS1
x0GQ2yhD18p60kxrF/GQqmDjCzmGIdFeLRru8Fi3snjJYPRTnaGDBX8d18ic1MGP
UxM4kJ8070cVEM138EUC3d+L1VzcZAIi96nJicHTB4lgxrEiNbpHSW7y+Ue3bOfF
Y5mWSaJqdYFbOWWCFDo2VqYu9qvSDCS3myWTCbqMi33vUCGTuBpHYdQT3f5eJ+Tm
emG38kFg6K4XA2QqtMYFxJ6Ki7vcwnhG3MghpQ8ckIyGf+u3QOKIw4iek4JpnmlT
GRwxjEzJeTQdv8xHpwoXdfqBO24MvG0dsABqr+dfj5Do7YBWP22NZtHvS0gxIXwm
1Unajd4+7HzMuLie6hymrgre50JnVfw1x3B3R4k726D6yJTOOEoM5OohQLW1h43p
SryjnGKhU85QS2/FD5lSo5s8yuZr8QJ1BF9sfvYZDWqO/94X1LjfXg1A+4co79i9
uiuYWxdkpzNnJxIhTzvAKnTCbvlS+mXsnIHYmAv1myZ9JheaWrrQQlkQlHiyB+4c
1+F4yXoA4BssOIRw1TMuT21EGmehvY3E7UYiQOCwJuQX6LCvXtS7Gh83U8QxTHT8
O4O5Vi18I118buF0PuALSrACy3Xe0IrBOZKvQsGIJzBqpEyw5JMIELGSDXVpOTon
6r6KqzlYBC9CaLV8ne+Id3xXGKuoYLFApgtEIS9qQ0JJmpkbv0daKSoRoMctMR5K
GfK+48HPVOzeWIKp7tuhJ+28R0QRZ1V819RufFLMcBz6jmqYVc07nV7r7dL2r4p2
Ky43Y0WvF/dDAwat2La5ehPcU9e0PVu90aeyZ+91aRAOOLX4TBP9DLvanOn0Hqvk
FvCZIEuSqlE1pgZbBmeXJxGB8YzqRycUvHAZNowB2KjghG/OyRAIRHiu0SndCnCI
EowI0NpIE4i57dLoPOl+5d6CsMjJxAIJyZ/HZCeCvCCIpVL0n2X22Y2AtpU2znXB
WZr1J3qW1uOPJRphH4EgbkQ1mQDsGLbwyOCLA2B/dLaDORWgpBb5oImHJEPsxL0d
gRKT+jkFOy9FlRBsKpL0quF0dS0K8bNFD+vcat2BdH0uSwKkGRzCAlRveE4sAiCw
r1YvzLen9aANawK87GeufOmxe4WhmPxmas+cO7lHsQbhNjIpkF5bETTNbm/AOEwA
8aJ9LtVs2MAoCNnTc4nnXGrjCBFoOFqwV17JC74boy5R8BSNcw5nT0DEjjV+gte8
YWKnPq8jw9miCGXUdiA40I55BqhChDY8v30DVQHlPp6pOAJxlCbBWkkWTP8wld0r
m680A+1mfy+H64hLa7/MeReBXxodtOxWLdqGhEFUDVWA78K0C7lxZQWhn+QBRKbD
Gcmi5LbJmpzriKtPmQL1a5qJqZd4T8qCcEyjR0BmKMGXgTMQ5ZlYXkMc7FFciddb
4pNNWeQcK9CZLLpHFaNLdPyV+J8jIuX1YMLofHJBuHMDNI0L4XPHUSLashJA4aNX
dA9yQICKmpcctUHjVic1sslQlEzeEasZfjUiYTHkuEKBGlbdYx20oZeki9v1nA3Q
feHrizOAgGDwFCyegzqtxEfEDS+F2pmcLnOHSU8vP1TGGoNrCm1GvXqufoq8bRSR
VRCWVztf7s2QOmq3AHi1Kie0JBFUCA7am4Z72eT6m45VSXEoSRHs0eDNp78TC4tz
4iD7eS9hiP5GB4PJFrnBBJkG+6Ln83TzBH99l2EO7FL5lC43g/xSONt3NxIGG4zm
lDL7QF7IYZTzWwSsqmX1ZVHLyYGpDkJcGJsnt1Ta/S/l7cSWAEPO+IOFcNUASRXK
JMlO8S2+GONDl7N1ake9gWeni+AJJv9Y0v5YzxoFFCQTH7ZmMAoZYqaRj3VIZEZO
CgFL0+tyrMJ3iqTbmL/cngEA7SWhgky/1Y6iH/M2dLXsdeuG0ulJPjuCIeo29hZ8
7poi/+wQejcuVgKi5jlLL3Vt8rbKRNuYk7ZaQdCBsTyiqTAm2YcNNICk28H4n2mN
9yw4Axldyj2zznoWXU3x7Knv5icwzcHMjh9x3ca0yBVlobMX7X+c3o59KXX6sER7
SPNHHpHtxQCmyZkreUOqKldjNMun0TjBj+iQpMI4W8c2nGDA9A4AF5D26ZIx7Lh8
inr0Nkwu9+hSqL9biYToOwmtoookHUDppA1SM5Y6mOqRwrQ5HAL82yEV4Jhd4F3e
rL2Qj7kF6N0SwKWPFOZgsj5Z3pQRCbkFxhuC3iYNYc8lwQVUzUX53yTiGBc2kiBB
VDM++fjwVdNE7BHu9TT1LnOOcILlQ1sJdBqEphNMdNj3Nkc05kYAwUTtPv8kywrx
8/VLnU7xfzzFb71OFubrKso8UjH5HtyfMMc2RiCsIh0P1pvdjnTUkfQ2wm1gK2tM
vTDD0zIGXOZ6rGO4xHGGLD7VX0h/Z01m5Qz9zxg80WINmhWaBdi88YUMEXTR6z9W
yuyjnNAFDuhJAw3au/cYBzIq+s42ZzAGYXNmCCaFds98Cv/s8jfwQNcuQiLMOOC9
Ykz1i+w81ftw1G/pY8sRijygtAX0xLKTMIK+g0OoW7ZtvnAGp+bO/JHHUlc72ytp
OmXTTcl1gf9rnYTerci2+qXCsVhencVedyvrMaJjGgPyPo9VjwjeppPYtvKXwtSb
Lt/V8033ucBoxlqCoiI8YqkMcJ57kKHHvNA7OiAkjCnDUlm97NYMWlK209MSmXWF
zCk+6/ZIStrUKyWIW90/eYjeQ4MSrmbwTb0hwVUa9Uq6nAcISh86V6qjeezlP0D3
2TGZHeVE4cEcOCjWx5hfXP4KQ/Hdo3pzpAHEgAIuH83bm0j8rUAuNOU5F/vvpmTU
kqOBas8X1iWQ/Qc7/2sy/O/zoQB0yy/y96gf2kekMBurIJOUWdHq1XRDb16ePf6t
W8nclumnWuagnte1S8epCDb+b+yO6yqXdVzCmnwTilEHjz0BG7M6FXOc8qnzjQ6C
87KeftNSvdEycRLWyP8ItC5lH7cUOhG/TFwLq0ArHEbdz+DW9TB+q78GnovQUbet
KTYPBsQocB4aUo+MqiesP0gl/HLEmkPKxUDSsNdOb2bHt+rTajAPobCLWn3U6q0l
GFWms0glyI3mRWho2V96wC9KEQPhy/YJAq3XvNCUshkxsmhZgXcQmCcX9dbFeMTX
Xah2QL9U5Kj2otQ1U1e5ux04Ws+c/WrlCMLj5H18gK0vWD5jRmpcR8UKym4i2U+z
qGKrxrvhkYGYepuGssVpQg68abJ6TouN0ocEqXwxpxPc3STApjsJuzFAg5SUb5et
1b414BC4kkbPzUtjQuRwiu7t6MvcljRVMf4oCMBmzEv2pgzjNU+urd+ypwZ0fHFQ
uxEN23dyGCdapUvutXU2bCwkzHZsVlgWacyjj3V0KSSA53RM8JHegD1TxeKf5v3b
Z/zrYC78zKlNeFQE27IoLz3TP5H6f0gbySSQhuv9yLrfoJzyXP9iduMqaccOCJH9
ou0WHB046P2v65cdLVWwM9MCDCDE3WTZUcdjVKvsAFiQKM0aVbf0gHvXr+lsZXBN
T5WMMC5vBE7xwpEsaVpJ2wyQxeEVwTof4RhUKpLlZ14LYODnyNlYFK7KzqC3fUEf
ikBUitm7QW8/3ivY6EoQNPxx+nMlpXH1UlckunsQvcG1i89cCagOD69FOkTiv0kB
tOHAJ2Ul9qq+rtSjUxxa5uUp119G2QaU/Pp2LTXSkdt/bEaQ1vKXJKk2dzgx7y70
9VdUOnFgwqb7mxhfNM0cYICvfq+iFQKgGDsJBYF7V5DUNayzn9a0vXtU4/LgIXtR
/4HZ+2cHg6Ak8Wa9pX3ZzhBFdFTXa+aDeifBpl+Dh+fm9AtDtFFoE+R+c0lVyvPO
3IfEcEH0E8xIx2tCauWYPwHtnFy0NfYsldWzgpJIBNCDj8Y9Gbi3dJyGW78b7ieh
K5Sk8CUfDUyoRzMbDixY8dkhk31ubUmE2ICgN89je7tx/azzt+8bjHDt+fdDWogf
EJzmhGSb++IB7UtQdOZqaSeiVODUDVP5p8NFogmtI8uaGrqQa2Mc/bfB+pCjQXsd
Q+cf5Duoenak8cv9Gwb845FC00MTCPIDWqDlzgTWG7TGCwbyqziTiY8PyH1jV7Ta
DBqwMMPe1rpr33sb1nLtj+dyRhIOYArApt5chtf0trQ50PCNDfPLk7fuZQPQI4UL
TSrJGVaRKKV7AA5OO5IgkYtjIo3NoST0hEcsCbgumLJJQmrfzj4GNqFP0Xovcf2f
3/jYvIPTNj9KGJtJ9b9BISp4d9SaZEmCgq/G+8lE2lLIvCV22+6dsARFxZeUuq8Q
jE7J64JngIj0pJRg3xp3ZLZM5VZ/0cGrrM+K7La4uFwvpBtGM2u8bOGmhH/rJHQZ
QxBaxf0WOwUbix882kFpMAWLCeTPozKUtF3Z52RK/10vSiJKFqGCw4pRQc5K0S+j
siFFT0pNOqZgbPTRcZiQdmOe9P+bQ5GF79GQQh5qBRnK3Bym5ME9PC6tvj4TSMmm
1w14k29aXe9jOO6C9+d9z+jWIYr9iVtI/cUqusy2gBC6zdV2VpV/Bw/mAOQrGOSL
TnNZV84gabA+qLhZmefJ0mcIZ/EPhTjTOGzH9pOt/FJNTt359LdzwGSG1XsCv5Y2
/l6+K0C6JP1tmVEWLr4S0m5OLFZF+PVJkTOSF0wmfA9Dw1tnZqtFl1vZyJXFEPax
/JfrPv1hqRhuv1sSDAjx/l+rWbgflAQxOyM4QGIHSQzz1G+qY3pkBloHDvgXs+RO
RI1RIH7ZpOcQQcnWkZBe1+r2A8s/vI5zxfS2Wf+JD9ILh4nxGnyq65gzJja2KUu7
ac8TW215CVYvg/dekEK1UsKksgYv9sEIiUOtcmamcU4/XeEb35JcSsnnxcEQGbEe
mGqolZjErGq2htK4IBoHcnPo9cyBRQjJ4FeBaVPr7Vbm53eE3IgerDP3UFB+vG0+
s6sG7bLBakJ5hKhC7VPHqPj07iFepR8cbSuAVmJYncyAaBo5+5i7BblEPZNDm7gs
7MvDwATM+3RhB3r9qbB2rEIBPfREgCtHIkocpsoaBxFOt7mWJwEB2xLjxVnh9H+0
c0XVLYTU5f+axQjxa+1Adq9wfKNK/NxxMd18h+D9WHAlR7D4q016wThuga0smR56
BWQB5KvMfVkgSHKezQ7oRhzwjmGOQhMXFG46a/DU5CFq71TN8xpmN77RwWOu2kyN
heiOKb7SIh1YCUePxtGe63Y+hUdhPJoiKHGWuBAWploKns4UQIjpUD0HDuo+oyqh
37Qx8AClalxot5TqdH4/Oq6+HTzlhN2PPg7yMN1xkqP1wNcDC4Ao8ApuVmYuF2eG
KIiO1f553kdaXF0osfhapr5xehJ6COOtyuhnPnUGbZXy85iWRGq57r+wNwcfbFHD
lY5NRVSkM3uD8b3RhRvotNUvF04XnPJKGVW09/6g5WKAJcRM0tFuk/9Pi9NmQCZT
KW6xJJb6LwrozRbDSot5dXNLvnro3tqzbppqpBVhrVypggXfONUtwT4hvJcUpSsD
PnklAOAW16Vk27RphU55sVaMLTJffNaatusQaoZ21Md4RIIEZJNKdEP0meBkDX9H
mUXIGMICdzFXOH6awKUpyvx9Lu/0vs02V9zRwKk1MGR73uInQ3b51P0bzhBSU7Z0
B25pOkkhOYwl49qj8xqPOOinuVo5E692tkwQGcrGhvQ6HDbxyO/kXtnFF65Fz7k6
2CPHeta4bZw6Xztl03lpUjYYmmLyzhoP7I+k4NobaYNTxGJM7Ybm1/yHjSbgkfJB
VP05rNU+xBsZJTWhraCtSvnm4+FGBtjvUZXIVCSeqDQsN5sWVhKZMYRw9nUQVkpn
YADtbVDzc9OZpCF83h9J2xkyO2T9ZqsRet8BTTLentLEy684iGFUzsCML/YbxGkF
hvrFsCqIPUs9+jz8G3vOnxTOOM2HL0UmioUq3v/a5z8pyueVKxTuBUMkhYgFpvqj
V6iEVwzK0Vx2ghiHEEbdTLGlDvCpiMJoDAxU5yI2J4YZS6ZVPmkIGmUPvP065XWW
Sf2Zhe2GaPlIGh6OSKZ/y/Hbz43zqw4dQarCuvp1GOIXWF5iYB2cCNMJhczyuxMC
TyerK9HJrlTFSnZ6k7ma3uSNgi0PcS7DgLjk+Y0XeqA5lvn98KZgnfKTcJGFwODh
AeTf2JDUnrIj98Qm2y39wPAhclcXEGq7hUdzrk0PQhnXDAp8fLk9ZN+aXWjZ2oG/
jzL499kZQcFe68dyDw/6fwRA+/9e0xT5tQTL1/STYKtzx74Wyv4aupSpdMbaENoo
vMBiBEJlAiXr9JAtEh8QquHX7tLb2KhlQgg/Nhour7/qkCroCej5LmSSG/LJWu6z
0afZlfaIQT6ubUdRzfDtP1Uw4xAtsYe823OTbp9Gsk6VT9dGqeKSdeYncilLxtP8
/1+9FYSLnXrNljnHlrkF/dsW42HMwUqTN/9wqMOCygDxgZCBYpouGParLta8GtqD
qZkGojx1im/R+YTH5Ob6nHU+AMSo1x9PqRlucKQMZ0sMQT0UQqD0aR/AT5/OKGbw
95S7a2Fayw5APfnJxk1hGXBXh2rQz5lN040V49it0nlvDyCopFLxlfi8LX7CmfJ4
lC4IclYwzx2NQWeSA9b8cfr8Fi15t9XrGSVeuo+hi4lmckNW6yrRGX6sYVhjCrb/
l354aI4uSTxgu5qIhe4budgMZv5hzxE6aFg8+1GSO93S4CCpDwYBgqV4afVpwYrT
Rzl5/mxUmNspHEOhZ5bhZkQ44XYNNq4vbJepmilPmIcYFy6J0kfzUglxk/rp/8hQ
DlJSqQKF3dbN5T04/Zb72+o8NfAQy7YSRWclXJmvRASaErIHQvcAwMqEbEcstleN
ehcqV1Ro+Ax5IX6r7MrVBQ+AdPJQ0RDdyko/VRiK23GCLV0agyQ0URhJTyj4nL61
0mynxo9Om0zrF162FVj4UZI8ZezyT7LF0Cuj3gHY59DAhKAICeMZQk9zYfjjjHR8
hoUxIvY+X8yig4EuLrIj7e8QIhxUcBQTLN68kwhvtt4J/nJoeXOqmKULGIAEFyYp
qtENGTdJbBfEQyNnW2AgR8qh9jXimeSrn8jqB9gbB4d5XBn5+HGszDRkOgQFovdq
zhBFb55QZe0Vzr3BRBgtFrfjvbtj3yJFoJQUbu2BgrZd7Qf7g1By9wpZkwy3qfiv
QhLE08lLbjvp1tv58bSqujurwL76Q/w9B0GnFFgLB6ZuBHo6RyVfA9j6HD30WSdI
YbJjo6w9CcrE3svtpvukEI2gayaRpxZ+zpRgHWR8Lk8e1m++rEeyFdE4iGGY0FCQ
TBdRuqLKb5kw6ZgBfT7j5c/NrUUUVIWfHxvs/nDys+iIXiEkwa7IHmjDuxN+IMkF
cBrSaJ0FYA8xqCqGprb9y7s7vK7Wggpg19bqZg6Z9Xr9FaGaIy6WtWvMQFen4yeS
OmypoP3+yEOO7XBKwCW21tzBjhmC/eU8W4Wzt/MdtJDlZUG9MwQSwSI/A+GumKHY
7JxTshwjEaNIZSO44ehShn7TjCwTVFzP0PuhC+0aBB9vJkXiMP+8oZDaCkT1SBR+
`protect END_PROTECTED
