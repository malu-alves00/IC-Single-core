`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
H/zc7owYijo8w15fn3m60aYilcb9XcfeKt8lqME23jS6LL1URLB7NxFw9KxIEkcj
XDaY31k+lEvMmuvwUyr/cyKSaTiaFLP970FK1fxDBMSiiJgGoaNHcwR3nigX7fvW
Rz5xCwCigiFtzFO/JzAekE8r6vmv5KHvgiqU+FLFRJcf7AS7D8RBo/eODAC7wTK4
+bKpOjr5CQvpHT06mBz+cti7yNLwd6ukWtDlG+bteYEQkdagr9gQSmqn9BgNI5Yc
wqfH4Etn+QFu0JuYms51aEpXVM1u4psDm0JFzYBzBW2Wtk5OvXBLqaKVK0tXuzvH
2eHmu3ojQtPPRlt+vKSEG8iQUJdbqL/OsooRVKX5UwHXDHoOOA+dvgPUnc5c18r3
uAGl7Zrw3Bd3u8xVdsbJTQGiljqHYl/M5jyZfTa+ASc19sPRNYGhrRvyhRtuz5dJ
W4vlJt46rcW5Fn665sQht4oftYRNcROyfy3UIqVu1nQ7TWGJsuo7QAkgmCwco9iP
zKG3FoRBVM5tEmFjuuheWz/Z1+xf1IkI7uI2y4HzS1eeOjatd6W8eRgRvZzB0kwP
XIsef61C+fF+h6ntM67Zg2pufREeGzEKUvfNubQFqRWN9x/TxneLsXZPA/y4txUC
KUbNZWhikYhZgTn2Z5Qw/P+Eb58+T5BLeUjFsoLcRGZITnMfkT6BkKsPXY1qioFi
MPFwFYx84PbZazxy+WKdEvxLhfLmMJbth5LWMItfx4VGSt1AREUA3XD7gp7pxNHH
a/06aAoCcFxbZW9MWLxckRODucoOXTJn00zqWzIhHF21lAx9xRiboC+Ds1cHlU+F
LHuy8cUqjAl8DzId2XD4riJg5MrgenE7OoxXqAMY0SHxWK0ebyqw5BIvzlUyD1bE
+QnMGMXNr5azEYFiyoIZRar5c6ZzF+stBj7UvaveZop7YLzPaGCxDCeSVu2f0W/4
5DxE/+wcnSWIe06CxE40t/ZI1c64vWkk9VkCX+yC/4A963HypgWtGYjizk2viWuR
9ShZ9Z7FhcsOCAR/mqNibVq1ksgpL4ak1scWjuEoEHNdduRPZy7WCe5twUaaSH57
+NeoEIPJf9saKPEPivSxGYCnfaofK7abWmTqR3UnPAT0v1MHrNLj7cn0sBoGucMJ
MeOs451o3pNxsKWDfA+yhrjpeh4SnOhL0J5qHiN6JnYrZh4X+6mLtwy07oL0Lq6s
tazObfu4YFi0UTysPqM+gUEB3n6z4JTw+Iymw2LMOVcPLepw95+m37WGulylCllD
KSmgcZzv7tarJMBjVt/ANiNWwEDyjNY/yxoTTzGpFQMTw8VJSJ0pq2inbEFx9teA
HvkKJz5Dyu2JmJHNf/sKVgtBbcNHchf2Ro9lL4LvvlM5g6CqU5GyuBTDJ63gjMFY
zBvaVdLrp/usFJq9EdE9nuRd1mPXSmJ2QgGf6pH8LDgDrU10h/dDqJ+FivyCBNYU
90IdOQ7Kz5YBOv7l5hLDaX14A94c/ZKoS1BtDOKJgz6cQVjo8lM2XXCaFEFHIcg0
1qLBV4Hef2o/StXxfz7QQDD1T5HiQD+OHQ2M8ccj53hRab9Eec7L5YorvbqLQMSX
dCxmFVK+sd7tNtdMKakZuhOv3bRtHTeTZHJK0TGA2Szfaisxf9rdHVswlav05AUb
J3MvzHi3opnKIPCfgKUBCxtaWY94yaSb4ZaP34dK5JIBMkT9R0brwZmm4DHOWS2G
KB8MtJb2+VSKrH0RGwSKmekV+Jrdt+x6nSRHp25+5lsTPU2ZMvPFozG6QlkLh/do
DNKgR4/E02yQNAncNx/4lSSErcQVwOlHzRCSgb10kjiZQxsf2y0asA83vFaP6SUq
eOD9MbrbOX9FwoDzo8VUCji4Aw6NWZEyqFNPz2Hi6dfanrLx40UQ/UvXeht5LfJA
WWbplcXIT76W1ksyzoTRksSk20gQXrMLnYANrVYHysnJ+WI67Rbnf82l263vDiuR
2w+oeyvSakXtDdQT3PlZ8nvvRRoSKdZV1/juLmHxqYvFCtYskVYsddUseX0d9zdb
Tu3smO8dvF+PEjqYVV/mzW/PIKU5g6mjcWMtjKEgxk0xTooHHpNEvMfy7pEf27Gb
wi94zr4e5uT9GWtD/BuhXDcSidhcoZysNWTM/+YU44Z/VJTb+zYJ1wrTEifQHsFk
UeQOjgckdLLt2oGuV5Y1xo6nouZ98RP2btFiLE8T345Zgsu/l30c0fzq8HSf5G4S
oH8pVNy0pIlbl97fXThQBASZlFJPvIkM3NuPgnYIamk0s+5rtCaRlxY0PiHLdZdn
fTfMh/PNyeTFY14DSjBT5LPxxfohNevrz6X/D7YVMfiIPyQwFG8QgYvoOuHR8EmL
nF8PiwsxE6cgU5cflwTd6vsrL42zd6uWHCTpN3RSFOtNQQJq0Uw4Qil3yqJID9tE
kC+qHcthkrEo/xy4K8cgZY9GmfsyRf6GxXg1eGpFgczSrPLzm9k/ccLGw+i8OMKk
tWT9dmlp5wVVfHaHFnP/KTyrLwpiQZrn2uWMlj0QTyqft5lcHeJGM8sfxpZFnHnG
EmbFTfrKgk2ZnRN3OYAf+W1uaAcRNasted+6k6WwiwEsIRGuf0CXyuhOgmnbF2bN
YUIGI6v16SdY4phtpI0cQ6jJSwEpyndYWt9wqP/0cdAI+XAdEOaifVZup1K829Fy
mFx6dSVytTBbMLTsyOK76spjY/lkQsQRNj9YVSrkjLxy8JTkO/5XzPgMmIrcknoS
xVrMMIxuQW5jg+cfkjfCVCwOvmxt3os9pV6SU9nUmbIjZJLwbfX6gD6et2UFzovQ
Eg1Rd147rJ7R34iWLKpnamYudf9nXuFi+WaAyX7yMePMT3yTKdAzt5OQVjUHwqz3
qR+7jhpTRFzoi5B6TD83cZhUpLUuotuygtGBalbHww2n1+8OwmzKHGT7M0Ruf1Z8
zWpCGsOFAELyRuks9IrP8g==
`protect END_PROTECTED
