`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5DWOctfsdkLba1Ip1TPPPCz/U3gmyQO/BXJhSMhSoNSijl5hMqv7LRpNiYBZ7/AH
jUdEjlZnhKM7/bl5U1ichtxXQvzxbcis/TZS7qfDjzT8FZ+RIvIAAsXscpDwHuXl
6lfhz/uqd3PHaY+aLOyCcPSCe3NGeC0N2Wxaz/Kq0okT6ukxIhivBZQ6cUZtBOEw
4BUGCtCl5wBP4rYv/fzVFrJs0MmBndVOB1MG/BPzH+KyPwbLNh/1KZfaajLwB7oS
+5CJN/8Tncl3b39C1CSpb8PiYGlRNRusohsJJu3gHZG7iRb8ASvjvT7wFedGdIus
IY7fg4wtjb0i4XdydaVJYk3/jNbiMCGk9uWbB5FDjPXd+Wc8csYSrpmFMy4J/8Bv
xS0eK6W8gcLPtlte4EfhbG2OuHcIx4XI5dRoRPV+EYCtuhb6vDRjAht/ND6seV4s
IQm1AwsMEracomVX+W8ai1rzOtrK8QSGhuzNXwWxAeXKNMPaE0LcA9GVo4zfUyou
y2jaDbGDBZolNLXEfw+w8ZJh4BxyuUSmdIV80+f2sG470+jljsk4WgBjIoD34YuJ
EwrfqjCblM61nnOFmlFFlToBWaYcmNHnRRHLA2PMo5Ykj6hVU77QF1juqd3cIHyH
84MOIdLq98AKfhm74uWFASuhBRzvFlTyAGAGJF2/V8g++jaZTUzeD5nUJjHPWNI2
tkqJZltMBBDm0qP7zkiLQsfaCk8V2T/34bFPT5RKH9pSTI3mVLRVN3ntQhtpwlp1
YszDRSIH0gLGSSiReDKvy3hjpdaTFGE7sj1/Yg52d35eJ5FZ2SNLJoBQrZTGDs5J
gQgoslgx/jMgBnmyXKZJQAZK+jGeHacl6Ry3MoJxdQQ1y6RuFoDpH17TLIiktwkI
aa3k/isK1FXGMenJHDZWI6Nh2U7jiQuf5iGjpiidf8GVnEp24TZDeXI6pKJ+li3g
nE4gZkMt7jAhC8nUxTp33W++300U99Egon1ENn+7fwfbm3UX9ivMSALDIr7Mp+0k
m4idkFcofi1vkMfTimXP/4HMXqz/WW46M0CnvLv+nYP/vgkME0ZAaEYT+qzScld9
YKsoETgyi99GZvchOHnuyo0Xar51+GRlyjJbOaHvLttVWO6J2HTDcFGKTYCjnM0Q
T3Su8pESjkFAcemt1GzhtYiE1KLm0g4yOv/oraFLYdbAfZYJ6/ba3+vbXlI0BVmp
Pkzq0Ms61MPyrHyiMU465D57or8Heh3P4wuZgtGZgSSONowNWUTooC+ENksDgY93
mI6Ar+7sNUWEUSteCeKz6fMoBlAMMBfpxtk8bVKqT2Q6EQLUzJSZw+oVFu3PJ2Ns
Xpavx4ne88DMrSYJrDvdx5gOk9Wi+6U1xEof9SJPIf4uMSiXzn2QTwRILYlsZ6rK
66JqQFeUKcrYgr3YfUEM75CcFT1dBvxZfvldEGqfPstMHw+yA4xDB23hthHLlegV
OTXHpUpNCCGGDowVaJTjKteUCurj/++mfluZ3K4Qrp/RJussxbBE625U1A4pc8jC
o91U9LGqv7wH7hvMHAJr6T6L55Hp7gN5u61QxB7icG+FKl2B2vAipFQ8LVlZIgqi
08wZrO/2L0+oGKoo81EEIU7URxIp8afoNBYuQ9Dzwmi+5xsyODS4SJUDlniVbqD6
9xjJi7ekB7uTYBNDJmj8tqvcqvNpeQnJJK8vT8dBTaqdQ7Q5a/6Ttgn6sRmnnVoS
4aiu/5DHxUKdBpojaFhqLizWqB9LpGhIuOEvN39m3aVr4A/6d4mFTn/jNjFgsRwx
dZmJR14OHOFc68kYbgvjIOTlCn4TT50zPRRRehdvCoY6QkLN6usEuhswxjqBD0Hc
ZHH8C5DcbxGc9sAxwNLMNMN90FCWcSEcLgrSfl2zAZ6Prix3bQU6oTyebh5V1ZjD
AnKBX/F/p2yPYzFqnvxDa7XTQdxR09cYNc3ibbeU99tsdqnCkV2cMB0xtP2sgRqQ
`protect END_PROTECTED
