`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
u7Y7CayWqBWlvBI2rkCx51syHmL/KsmIx4Cm5SXBSttvOVYlzMYDJ0IZO6gzsUYJ
BepIKXdlO4yycPejltNQJIpqnrTh6v3BzwLgQtbhyBXdqdDGSjJbbkXxM+KNlgGM
jcdBXZLMOKVGgUWVfI91JbubgBltrv3kldlk9/KgMF0pIGHQhkJpRR24CEx8ecaw
QAkTYkE4MR8ZTW3UJjH9mqjSVwaLWnCFVOcadC+0RhsoYc5ZY2zg10ifT62ncmJT
XMKXM7kG5CBjAH3iu1kTbFuGJoMKm4oJlfbj6hnf0Fe02tdBn1fZIw986YDklUNI
sBNRuxmBqd5+QnKV32TbW/qOXWPqKy3GZ04LufDvm/U4/LDnBtBMan+QqApy7uXj
W6j+WhDTq/vFAvg0Rj6RmII1PWLKdWaOYh/Mnv0X1fc6fc6L9MeRl+ejhXfwIwEm
EEtednYnP5uDI2jgLxJ15Y6MbvHUKSYcqwir5DukCC6MCpfuvaEzhhN3YVrU9VpM
EFIBk/OSCB6a5EmHWkW+sHqwQ6CCBUvnso2W1KxFxTF0eOw/Exf2znjdkD3vCTus
PzjJW3LiXnsvnE76ENhrpwFh5yD2Gt+wuTlPaZBmecuxJN9pZTy2f0/SLPkYNxHx
6J7h1l+LP50BmFq2xMIOE8hz/lriqxcdFr0btHcwMFsnC+eZ599OHT72xZf/2Nqw
njb5O2g1UoixvRtwEnbF1NRb5WjVftVKAqV7w8O9ZVRqLrlTqqXOr63mfStPKR6d
FE98qAnKD2gFtIkvEuyGNT9xUGl23lquSnTtDEnvZ+INUMcDgWinKcudg5L/yQRl
lKr9DaaLM5schTTtAq1DyKKAHLQL0lCPfGn2vtR6wSl1b0Mr9GOd4lOJNaJ7lZtI
fD5ZkFnsNZmcEdtXq1Tg11lurzU5eOmyuBdmX0ft0P6WrIkg15q7hZcYVyfszZ8j
O8MA1V3h+qRHq2YRWgYsX5A1B9ezxEKUoyvUiTGrqXJKpq12CQE6HVH9k3J0NzWU
jkk19+BjD5PB2M0U5Ycu6J+LTGyaXkdmBw4g35Lho4M1PDaNvKZWunVwsOuQVEbl
9rl7VEYBNh/XYSMkMzQF49IUErZJVbBx6ComFRn6XVT5W1U/BuEOBBAQJEo1YWFp
pzf7ayFuZdoNH3nhizii9A==
`protect END_PROTECTED
