`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
24547Fula3tE+3r9R7TT4e6FZIOnZKa4UwsjygS23v4kLI2gUyPUBF/l8x4XDr/v
xC6Kh9R16FURDUMTsO9ba+iiYhs1zN7oMOsxgAF+6MWbDbZ7IAL925YcE0Eb2gmQ
XDUY9Bkbzwwo/Bv+Hidsi1yv6DXUMBkuZwq/tLHdNxHlehACodGji0QnSmYOF5LM
hryCoFu+YUpvx1+NiUnHUi0uXl3fKhH1B6YKusuLg1xmqBb8ZPdKW9vSmnJxPd0t
IB6cHER3hrM4q7qAAUweMg4Ycoy4NZlFqewGgTOhcSdl2mQP7V16fs3abGhxz5Qk
yNlUHTMTUIYjvbO6PHNjexuS1SCZCQvcdbMK/HMmFxIhKMhUwrlggJU/t6jR9KOf
399USwhS32ySDGOgeAFkJEQ3R2VjegCp4P8Y6vVNtKXdcNaEYaWPJhWwxrRYj60b
W1jhy3X9ilmhFZI5sjzuzUQCkZrpJN4coSEyWaO43OfGjbRHEfDlt7bN77mjprEK
xI3/vR9UBea2EsJ8rv+MgOW7k0OTWmKbz/N5cL/KWOyQlbDDNb8Lunt/JRdAS42i
zcFYtx/EWJij1V3Xz6RTk3bdKj5pDEJ75e7JjMd2esxrk63I+zT0TTbZwr4Q1Nc4
5MvrulXlsbVAxSN0IfTVYyROIN1kF2NhvppwIIcukE79b0oEZ911fbpB+zuc0KxB
xWOINFviEXNpeLSh6OHaa1RRwXeNpWWG/HVoX2/hrizc1AGCwL/u7sgvlUJHkmGy
aYrAq7b1njEUnaLfAVb43QKONAFekOjMXY2Lka1BU0aUU5vUKxsYnDxCS1AM0SMS
37opzmKadKKnER4rAV6duLDtuMTcKtGnyCEIezpdv1zmNUG7cYOh5rmvbp2LvsC4
+LV5qftTKGabhrkawNnDPFycNbHCbqabouvaNYGtH3vOgtBor0f/9FGa9Pb8wflO
Qtv7avzLCMoJsVWu9hOgDzEtXbxhNX7Rz81RQ0niYCBgsTjH49mKost1zA9Tl6dL
oE6wTb4CvXzcj1iXRsC4iPoi4/jdLkBTxwsKAU11jQX6YZeKeQnHjAmW/t4WyKBU
`protect END_PROTECTED
