`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2eOtQawZdvyP/Y/cHZIKhpbQh1UgR3HApR44v94HT9P9mz+gdkU8kUuQ4LCyUJIX
lEIKbkQ+X7AGyZw74LgM9cTQyei5znOe6X1CCgdY/U/ydBbqjmzN26GZm62E9sSs
6KvWdL96ZgMBKcwbMblnx/h67qf1GpdxsdfNChLP3JsZaxE36GCsreV64RR3J9Yv
fH19dlNWy/rGD+bJ47mFPRYzxM3fUx8i1Y31/knuCGjVcB3poStWVX8YmvU6snHt
0+Ef9gPJIM3IVdGYnsnGTQXBUAUkSoVvyJyOUXEIlKLra70YHcVTNgO7qNECgppe
WlV4e6BtQM6LDnihQlijmWjqm8v3FWSX5z5/eiubgmJ+rgQeijJmdgatZ+IPe2Jy
WNDSTYE5lSGdF8XfeyUOvDE0uiOEZv+0gbpD7h0Pqv5bfn7drwaY/MKI+afriVtP
xyccJ8uB6hrygwQgEABpcCYFEtiXwZCGpVEf/X6TPAw9EYNwlW0nZkVdRzPjJ208
bqGxeAxxrlMO/LWbYEHAYJp1DSvYo5269XuHTrGm2V0N3sk7/N4hZecpUzVJgGqi
wFTnhupe0UWz+T3ArB9JMIZ9q8q1Tmh3R/A/2sRsjYmRVqRvXRUSIM++ElXBhU0N
FBEDkTulesUis6+GIYFIgKMjxAKnaLQKZgTdPF/SHICI8bLoA0hBXWZtcweXAhtN
/gFbgSk9f72EDPDQtQoRBE4F8hUcZqre1Wu5p+6xPXSoa5R0EL7A6Z/1TxQKJe2B
EtHZh4AtjpRtidJtODfyhV5vH1lwUachHMIM1/mB31O2g5XoMA08fQPOS+Se2Rdm
cWV5kpaPeCv13tLwhVX7Hf39WniNGFzTVFlwZLiDVtqaWoAQu5upRtmzmONfKUjP
UrdpuA6An2Gxq9v+diF8+qRbUQ4gFc6uwny9aExtICG/OHTQpuSawlGMvwD7y7H2
8l5PTv/9wSxOlKKZ8y3rSTn/U0/YTaKmPnsE4ZoygaoLUYovaUyYbLtIW4BSe/t3
c4KYGtr5eUNGama4pwmiTo8QkoQTxw938Tr7YJ+U3kFLrgi2oxbOBn8RbK8VEQE9
NDhnTs57AyyLMidd/85UxINy67TDTjmuhQOuXdVSKKqMDXSiU1tBY12j35igRhAp
syH1oKH5qAXAdfzOXXm7fDUqqzJL8VlUt7jNN+Eg//ePis608BKYY8b0x3LzqnVS
GLTo0LRib1uSyj+hrrAjFhqUz3bTLY7HO3z/AvkOousz7DKC5G6V01puFSSIB5fg
jApH3Q8zPxBwI1YTo0W1Xg2sFz5SzsqnWVDaqhD+ytqJo+Pyl9U2xH0h/kFFHyMg
XNhsqDaK5M0lNfhUJaN8QyvNFxgchN6FAPQb0SJ3byw=
`protect END_PROTECTED
