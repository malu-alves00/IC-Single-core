`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mY2B2B+rCYK0zS2CYNZzIWeYME3K80a74ztFpaXA7IjjdSBo54aCkSNV2qsdkZjk
7lUS0PUUAP8Rn3BKGQ3X0dtbH5dLYunsJ3iHvlXm9o3grMaT8QQaS8af+C+crYC2
Ko07L4o+CKAQcHDRAGFeNTha0Al2UVsXZONgOPv2rH0dmSBlyeVcg/JqAhH4+ttt
BSaSXKmuosfuTU6cvdnkQiHHpHFer/ZTIKCEPuojdCgYR6Z352lD364vVsOY/MT1
DNzDMszTTyiPQDhi5BvJT1i8NfZwztKzLH9IRlPMwhrHXuvlLRj5YyHdvz0L/ej5
mWF3NcogqrJ5jrtnGHptAakkJZizpYG13vWD1fYVpQuJWp4iMq2A/FTTAb5SSE6j
Mdymp2tna0j5xkqPFLDPtJ0kIQjFPeCUvfZrRSCrM8S9g+yD34uVV3TAX5RMkS1s
uOw8SPujUcyyo546jzDUmcmU6n6SmTnyrwuEVWTscXNGGaWeI9kuTwzj/u4RinMY
G201xfNthhyMlGfF4sUZuFiPmv2ssRJUTrIq1qSTKRjgQo0IKlsglVpikoEPWjGK
kS8kn3gnjWTxDJ2aWo+VkSxqYy9Kcy5qw0z+9oOs6+e7Rw07wFc57Wv3nVGpfPr3
vXuwvRfC+oAe1q1uiqNTFx6gcigdOQlhiGohLPDMHin9+BUQeb42Or9aUvDvpu+v
dASVEzB77v3vKGWbxywGlbcV4ZnzJBKGiBVIqJMaEPOssJTKXvhaNdr4QQVR5Mcb
pLTFZtsYNi9rykIBXDkwKbq6uKmvDIkQSfhxnhrqJViTMWMUMq3BIAFy0MS5M8Al
eL3Z0iGVsJUbCSEAqx9FEfcJMXEwSynQMcWWdYyrYbh6Dej37q0DnQ31sKcDbfhX
/fZnrum+Atm4TPqxXLCIRUVMvgQ/Lr69KzYelKnVEakhcIFJR924vyIlS65ZbEL+
k2sTJreWyEbSfl1qt+Pzd9dMezrhOC7SPPvaPWZloAhn6GgnrxQ3OuLEIlO1wEm7
Dsw62UMP0xxRZA9LaHgQCwvcHU0CU5QN2QTXdSCZtvtQphQk2ZCLnQiDOxeyZP5u
XoI/YtFDk5VuvuscrJn00Pi2IyVYfVwfExHvcm5wc5Si4NvbnGyXMwwML6tx1bqc
lpGAftmrWTMkes6ZAae7Kj3QwZd0CsBe02sOW1xPBi932XpsH0XhW34b3bUzL5h3
4Li8BtLjn+OT8W/TIwMCzF9+WVLBr/hkwR4uQBrenj0mG1ytnYfo7ZFVT2obcqto
QIY77ttwnwvAyCuhhozaT9p/gHH4U1Od1EJRl81QuvcSNK9ZCds31+6iCWT+CP6C
Mb7N56jMjefemvvKwBbtjb+gw/DPjI6/8C50FremZ129hckZG/AbBeYf3DGwymIT
1yC7t46SPl1ASt37rvn/Gf6x46NlJ3Nry5MJRepovJ8d9ExzN4CsWqcYArdoTyqq
zlvGkO8Cic1MaPbsDfcBn5Aq86iqACOHclUQKklQLon8JyEXxqTA4/Y6tlZ3fz4q
0Kc6GkqyadynyUs0IIZll0eowh3oaCKwDWDx16jASM3MSFFs7qKJA06VJOYPZ8du
XeVtsPlO/lTM6z9C7dFsVlZkugYvev0QG3GIaQU4Mnz155BO9zi3ZTfWRo/U1xvo
FruVugkRg773/Xvj6OWMhiEQ+8ZyC639y3JpOFgksH4eegnHf3UCaMm9BjsDLpNH
1UBZ+IuQBsAHVXd9hvKhv0bcI6yZ1L7RsgCm+GUc+/TdRXaG0rIHpByGKF46wcuh
i9duTypKJJIbLQR5wuyf6jlw5YhSOEeHVaAL5+uizZvKhOEiSPARLUyyrkObINor
bF4U0TpbgjBAxTWOEsJgMUvSmjwWx8w2QCkFpFyGl39oNSIgQTBV+ec4remMYhnT
eKXXoTfp9Mp1cfmuDStQOt1aWh6NN/8BVpzpevDLhmlvwr+ywvXNwEoomM/Z+ZjN
lEKVGIGHtQ4bzr78cexU9W33Di0KPskA3sz+C0mxMcqrp7iCfV7NFYdr9wHrwgRq
Jj6rmQu66aJgCOiY+h5EOxNgbvra/V20FRZKjKaPlIrMCqT6aa2H5VUSODoEjhUz
D5USPAkhm4R2ECnS83pyVaj9dwa0CxQqJJEuyqp29tMQj1l1ervCJceoCNEl5mh7
WzW3otcPvNrLRnoX/+GKBNUrvxfLceIzpjsu7tvNJWvYh+J+j3GIB3eC4z6gtNxl
LlwpLSuifRZ6vvtHjF1W9HVPjDSdr1z4jLaegj1M0hBYi/EcroRTNeCmRimowXRx
+++M/xIbxc7rKt0UInMppNs0JyqrDjpkljMOxRdEr0/Q/nokSJqWWW45mgyWEnX1
2zgfxnhtIot6QzTfDm+FSqUL3ctm2neYOtWNiZyyaggnEk54v7LvuK+Xa1iO+JEL
NBQIoc4xsVDaLLfDaLJO2U6TiR8io/MEVpP5lYG6mreOjOqnKBsSMFseMWkeVyj8
39V33yxGKbk0cujWf1LyoGT5mM61uuSWUH284wj/5wm+TbLuBjLmfqO8AxJon3TH
cl9C+ixqLulNX+U4LPpDkhLW6hZGZ5nZubxePpdSyXjpDhNFl0D5Y7DelQW7MJQP
dIjsX0HuVxbq7fvUeIxTjFXAquT4ortTjAsNzmjTzS/fKTq1VEfLhCmNu/ZYvQ/r
d49AHXuM/2ap5yND8NvN7RdKC5+vnTsulyUgStETy5awg+pb3qkWYn1PEiMWMlNV
z9hdslTPj5Rhy0ZXkQd5z5GTbw+XwlNHjKECmrAUrE546j2j418rkB0mfeFC2uED
DYvynjOiLP8SjjQ3Tdr895J+mUGXTl0cI36k9lnsajMtrGBvCeqcrYxoLpDAb3qZ
rGrs+VI2+gN/oke7m/d72S6kJAmrQa/DvKm16qNRIqKG2zwOkZONY/8KLuuYdS3c
KlsAdtceyMaOyqECG+8R5T6HSS1yYChd6K501FzcAbIHj7ZSTb1I9+jirhVrzEJV
o/NUj4q/VE+9sWpv5XLcm4c6FlvVeZUGe1FEH/B1U5lNrrjhVTwYZc6HtM1/ppEh
dgP5S7PnVqkYPsjm8oEMb7bYEqN5C/OfTpmNNySJpOU3G2ZrQKWu1c5ChuO+lBWe
Y7Tdkv8gnfV7iWEO/U6ifqZm1rFtysPqR7R6HsElQpSnImyX9KbLFjzhTrI65Eiy
UtzQeFao9290yb0kwFXy1npM0OgtEGFcqJ7XjAIj8arQG38zxObYeBzl/lF7AIZ4
1cxqImY6bvmf2BZ+zJGMZgKeUfly0Vrv7qHTsQhdwLd9ZsT66bBhpPYwZy9GAjUo
unuAEAHuUJ4NA+B7Q8MWx022bW8YFyiUtzq/44H0jir5qr71w0T1P4UPBGzYmQLo
vqCdQxQ+uFIq56lV/yOlGGw9OWrTcDeUU8Pjsi8X2qAur6MD/uyWaTH3YxQFbXQe
OpUwAgg/tQTfco0qUTKDpl8lFrh5A6Rq5FKoPSSf0C8ipfBFif8F97Ieof1Bhf/O
KCJpICmk0Lih1VAJt0aslQfMCxQdgGKQ8gBG7odKYQGg6ZAH5j0VDUap5TU0PFOl
2ab39IAs1xQD6AoeGVTTml+X7JngvOuvb1/ARYsxdTqHIsNhadHMlD8v5AM1tABM
41NaNnY9Fu1Y2ZXYJ+UNWpemvkYZv+aY+G1EFuqKkaCqfKczWnloyvyQ70u0jtsl
Dk8jjOtYjpysyw8Bnh2nbeqt2/VBTaeOLo+SIfghN1o1OW3TXCKPOY0A7dP+GGeN
0y9omopitgvyhPO2jzOvXOWYZYPNB3Rlfa2mVTkabPH8Ob7fc02ORP4VJrOCWuNk
dEW/TZ92xDHyve6F3xqLyQ==
`protect END_PROTECTED
