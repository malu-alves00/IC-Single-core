`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
c8R4mSbsWjEAsGFHYsqUzR96AM8Yt1qUuCLLmSNib8eDZGth5E1qkugJM4Znd41t
7g4JZYe43NLmt5cLz2MUcU8WktWuHyJL3SLGe/fGbQrcj+fDeEkx2rUzMiOkTBFv
1HarSHrFv6hnUngO+jf+eGuVM96b2iObY8wOVe4t3aawTuuynhe2GMGIo1bd9Z2R
ei+yw5u2DT82p2Rlkkllm74UebBaE8ZqzB+cZuhjnsezd7FztqfCdquivoG4aj8e
YeJtbE/IqHFJGAQU95XM/DQvY/4JbWPP6sExGOy6S+DlWkc/FPBs3/tj+qZFsboT
t1G+tCDdkr7KpEvY7z/rSUhrGfqHwxAY/DXF4w0RECNAU1gDIZSQ7JounD04eBJP
0rRWTTnewCYdog82uNwfrxLhSXbaN2fvPG3sqlirzaColYp89nRDdDXfWHTd8Wbv
N6UFAMdMXkBtYBVy2mmc7VO1qPzINPvLFa+D69lbgRmczC7gUsKxqBwo4F5etaXT
I8MHY8/l7XePWTvUhfHTW3/cS3DdO6wg5Joe2ZT7tfI5QPfetk9hSD5waoI7/caM
j0337Juby7p7MaxxH60jG/DwEXDs2pwSf2QfU2wx1TCfidjlzeJVW9cHhB2lpPD7
hoZ8naZ0/29UEt4Qcx3OVcEC9RT+QlpYqDJOLgCZC8d9cYtbA2r6jRvS5qN6Fs7Z
21DxIluxC34uOgIaaMfSOZHUYLEFxGnq+qCd4oJPnKj37OnZ7l0ZiDxACO3Ev5kj
lxIKd9U8sjHHRG6KiEh0qF+uoLqbV/xCizPCOEOxqkhhTDo2i4uLWmsiVMSt8e+w
hFhzwCISQ/xzfITkljFMUg==
`protect END_PROTECTED
