`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ucxGxLNPhFeDMnG3lPX2wyz3ppF22MqeJ7Mowho2kqNmEQdsU1vKMuiBVR7HGn36
ckFr0VwdOIcJvtUArPtRi+SkW0uHREQDJ2xZdzSTlO11KJxKW+LLyCuizILcz29D
BKQjmRL3s6J8yFER1RvzOuAkbzA7EgBLO6gwTD/NEjeVVdGjw00gWPPO4RyY7wHH
c8kQizGONIxuMy3jy4u/8JxsN4ycn+cZaKOMPlzcxFi6pBDGy4w8kOcwdNWW/bhh
231o0sYYBttVa90VPGwh29YW2ui/r6rrU4+gLL24R7pslwVgOr8jJlS6fprNcbc2
UoXGG9YEi27zV8+EueoOq4nLjKjfVRvAUmwx83peJ8i+AnVWvmHmmlZQjd9/e1Ya
M08qqmzP+xgbrONyjqlsTEUk2yaIPcye/HZQidfC4CjLd6kVTgVaPSwxDYeHnf2Q
puvvNoEfFhnBVtQIWWhzFIT7FdAvKcKEaOtO6/zRKAX84QLlABCsB7zg0LdT545y
1VhYGbxrh8dPHiw9KmZEI6sWIWVNiee1OjGE3YUkGWYi9U+oPGR7pDEliBB7V6e3
kRgtCeD+W5pDLIzLDXMNp/QtrJDOowP+H3NtKfL+zG8QqRgEufB7jsJ80uTRVBRD
2UzIO9aYAWsZ5MEKRdxOXflf2T/pZ4uLtHCuuEGtw5YC7EdDOkXbORm8MBtGlyW3
8ON12Je9DCVVaNt8csqqb/uz8oqwx7YVpNaKzLslKJ5wiQTXILLUJvZt5S7MEIF5
/ZDWT+tr0JwA0F8eU6Gb1ibXfLqphtOiPyB9hlKen5CsvcpR/KR7MXtDSCmQVSoN
lWT6EGFVMlMDjIMPB2NslObjDXAkmgGhfV925Md6LM17h1O9G1Rc/Wfy21G1XilM
CxyNG5+t/qtprhDTaY7mIh9Pl9JQUl8uIwCZYVo4+u5OT9xQanPe8wuuvDVSRdKo
Vc3V2vL0OKkSZ5wNkN44m5e8L+atyRhSujnljIMeKzVUNAcbaQSUmZ6HHEYkkn+H
9Fu5i1DgvwHp8fvcJxK81jLYn8B/vXn3nZfoMgYTY3ocMxcB3iu1pOK1qfx4aad2
sjvAEfcPzNut4UjKcwd/3SU3f33d7NXnpCwRF+/NlLeR5q0EWzSOg2hMGgynfJVp
5Yon09+rgQhCfPL+s+a3uA9TCpQPoVLT/Y26629SPTDHDJj0GDacFPZBevWQN2jx
smPg6yD14kEUJGeXWPMSvg==
`protect END_PROTECTED
