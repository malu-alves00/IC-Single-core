`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UiiQmb/OCQgkg90zTg7AJCkfChh6v3edB30cCubctJKYt1U0gvFqZs6xoozo0bnP
3Djr9Q7aG4KPTrlyOu1SeGTiCQBeQvnmeZ8eqwN9y+EauUZmZKY0XQDiNBEyfphw
f0e68dhFNmec9KWRr+7OZ7CpyIEeUCkyUT5+o9WG91lZkLG1KGjnOkORSxSUuZh2
jhsgotx5DlN7uBBAq/WoFDX8HfSR8lvcECn46dhBofaeiI+M0i+FuHMqPjkcX0Hv
flrb3eNidqq6LIcrZYOiF1jmEdj/E9xHX1QHLcWfDJZCv+wYb9exgteJP3fEvKzD
MU22YitbF9Zp7iJjOdsXp4SNPe/N7CCyauC/us2go7Suf5eKGPtTtPk3gBsPi1yg
wroJKou+UJwY9KOTMiCse55KJQU2YPkvRggvvCOIujX8rTHYQp0c+BVkHwv9HXAW
I6GF/gCte48GHED+0v4DDlT4Y96kP3QvFGiQ/64z2k2mD9l4DH3cR63NhFn2m8yF
Az+F9cKn05a3CYnMzhAASQMh6RT53fv19iK87fuNJytayLZ+CEbOB5nAEOQTRSI9
W0vuAkGu/NcyJAnRmiCGCpxn5f9XJbSBT6Hr7VEc2c4JxgS0oqLonr99Kxnb3LxD
d/mb4sslm1+AlxUgwDe0cwwURQNZmrmhgT/cVhtUdt8uYwDBAuikDTTIrIC6niKh
pM9pbWwQXO8q5vRDUxP4ALG5kslvWtxcYz53SRgU7kzn2WL8yu6EtWAsrfkZuJI1
A7cAhq6or+9czXo3nOqMSmSazsCtAWfytkYXXYjz3o5KwBJqNtiSIaz3Q5+y2S64
HNlRWLcd+W3rkY3PGO4XrGqNj1LK0IDiGdjVTSyDUWkk5QGMM0nqdPmv1oM2/t5p
dkyNWLhSjGDWcByHUgefwbN1XkUqW8v4wJXsfHF72aijPHOsdk7WRB9AGrHtdlqr
A3292c/J6ob1G3O+L1T//9btnXERgLKTIATRvmWtHnlImRX5J3OTXbVDloMUOmGj
LH1WxQBEgYNg194sqHgNaAkAEYLjgGSfC6/9F5Q9FB4aLtUib0y9Zp9cJd4YZwWa
D/zwW2ymc4tnQRtz8xbsKDZG2wcN9eJaO/cAUyqJViNyI7UbaKqMcSHSmWWJH6eE
Ip22He3N6NflqUigVuNQNw3ytd8nx2vc04wjZtCqCiLpnd54zCLbjm7uyAOMEvhk
BCC3am17hw3vQ1d5fGAcrGuSsr02G/i1LlC8VBZANELBar0Rek6uKs7bpYHhi+V0
hCIs+tFnoQN0Lz2u5Nn6TZshImRNTl6g3Oxn39utbDtXdQ13u9cPJDe/YyeqHvQa
4dIIQmsJs3A+IcrWZ+NM4l4peQJHU3EE7u7xTrdDlQ7xyB9FezkYZ2JVMT94UI9Z
u3Mfj4CnP5BtwxBj2rnwWWzuMr2c5GTBnY+ELzvyDyrEb2kwf4ihWxg9G6fw8xmx
0AA5o+V4tKSWIJx1jGutl9tjoJ1URq/Yd9iU6WTFtP15TU8QvN4+Yn+z+SbMOFZg
vMkfuyH5XGSb20XN7yAy1AluB3seLG4jctPQIWCI93v8n+ZHBfquHvnJvFcHTTWS
AxkXVm8j+j3t0ISFy1BpHP0RM+NftjceOUpJGqYWLl9dJuMAn2t3FhLihRO7S2V0
i/lcPL3H0HsSDVW4HMnBogdeom+0goiaUSijsw+dACczVL3wy8oBQtmojZY/Oa8A
q5i2jSGSkFRJeJfWLyP0HRfzPquz6S+bJ7NOfP6ZCW0LKW6pyCEAOA/W3AxlutT0
4Ucf5UXf6i5vqTonk5AD9Pe/BirZw8hBx4DcR1wXXTeIa+9k9aCQm14RQgaGHx59
i807BQst1OXH7SnDbOmiKUnJC23VrJ9FKz9fv/5gK+BiaJWt6gzVzhqnq+hlz4RX
CMu9Np6NCevLFMAQ7xkHvUXiXX+IurLZ4+PIaThZwmx0ZvJNTOewlzRp/YFRX8US
Lt/5NQXIPe9HZ+3WErUZfTzGpdh0x3UBeGuB5C0Fg/+ET3k0FHE9ggyN+2G/IgXV
kbGKfyclaautMr0/ppv/ft16tLWQAVV18dZSphGZmcigqzcRIHIY0EXVCVYMpsiZ
edrwn4x2jb6KMMS139fgOtK1PHfgOD0WjD3SdC3XcUQyX96+gpL07Jy4WmmML/IC
HI8T5TXCbR+Pec9UQK8XD4felC+WSfzUx61R30beYcWvQOxWrxVNv9IzZXRUz7GD
UABvZGc3UxLpirVBp2nukMC85cBCmVUaR+5tc2FYu6s0ms6GUJLOXLZpp+9qjVmZ
fCd5mHOzKQUWm36EhmiVWhbGUKHEX+H1b3CotSpZYsoaMKfSw9nPEToCph6dlB5D
U/0TGbDz3wqq7Az9dvMNrwkF4yNwwMDSUAx0FCyqbsEKZmbI75iK/6IdA4FaIXxK
F0Un6E+B0H+H7t1Z4gJkjYBj+a3e1+6UzSm3J9RXQof3dD6ZJDE+ycn1rSPgPyDC
gxHS0ZSOu1ZtXO9Tdnv9VwV4jVY5owIh3k0ItCD+YV2PMJ42bD2yaL4Yp4lnzBBO
gP1QcwFXsq171sG3C1XXlIS6V2KbQmBcaUmdVEJ8LSVohlEkwHmvKUuCwyulJbo4
Wg1A8pIpq9CEhKsjlBorsA9suYO6e7Ypnyyxz67uniXMTzDQ9cpog332xVmMFNnj
MyzKk3NH6ILyAcAEXfvrsI6EMNJk8CKgssK0qWmaEoOSBqsBY34ZkKM7l6YeiiI1
/TItw1ib3f0ON406n2c5vcjwYqwgHvmWrlshkodYIar1uVjN7qXAdC2eWKbU2ROL
iPB3W71jLfJpXs7sgIN4ozlHhkTQjWzMamlLvyNf3mNCskTsnS+vUcHMV2y6cIFV
pHORDrlm2PdpoBvVdvmGZ/98Ccr1ShVaQjqN/Qb7fn6em9CqYPYXfJtMutz+BU5K
plSFKI3gmVyQTU9xBLL9y28WwRzzbr3ON9HsjyQL/7NvhDtbO6semFU4S3OXBk3m
ARYNSW8tMOdrJCUstv0zxS+8oECZiym2gK/o4j9KCzrkVF0A9RpQm6F7CYdn6S9e
8evaZWbVKDQ3FSmqhAWzh1Pevabmp8aD+1F0J4nWEiTZhRr3jaqPISubtuCdhEnC
WEPom5D5DZbU+3Qoutpjbgq/DFVvGgALMaOpY+qSVud+6Df8wfk5HYY4/YdZpklO
5AkUV+oFO5VgMAunpnZyUry3m3OtNURv0yIccLuBICaGMPmTc6I5S9sWqsjnoNVI
gTs/22OOb9YM4XTrntiuwVxcZvE+GB0URaPsetc6SyWzrE4rgpA1xtjcA4IhYnZ+
2mCbzWMa8d+G/4EXzihSVTPpF8lVLotfmo/YvFaWwiURUCJxAMr+w3HLlo3sNwBU
3zszrnGVslNxEMBEZa6bGWrlb6+Uq8Lk5yJ3mF8/p+/IFlteIFoXsZNNWG9Giwf9
E332ld+nhYsleA/Rc3Rt82BvlpaGLPVTWvL6QddUv7u2eou/X8RmjP2eEAtWlw+K
wlIfGIijQ4YcQQTj2a/cwp8iR9ubP8SmKTko2sGGrB1ikU9lcW855B0IBs7nSzZd
UnyeRsWbOGhSuHQ50/OkWZO7NBBT9oLz0iYM2UJmgQ2OwfJFeQ6VThhjGgrxBNz9
HULkcDmCId3tT5lNrv+hi7kG1yFEB3n5n11Fj6gJx8WUi1/lH8VTO80BfGOL99Zg
eFEtQUeVHQz6Tfx6mOUXb98ofFsIokvez2cRPzeNrhJEtpoAoDidUVCLAR/CxQKp
teqCanhX+94llcskoCMZ8Nyp8v5thYqjIin0LIyjlA/mruuhj2osd7SbuFeBXWuG
PQClqOVF6r2P8KHnb0idHFBVYV8A7zFvv8LwVuHmeLplfNTDMuFbtluCGdR5+Q2L
tJxHvKmrah/EVxpeHSIjuaoAjAxR7DzaWzAFwZd08N8jusmexQJtiKRS8vi6/zeg
kzhKK6TqJxY7AyuxextsQGnJZnB3an5qoE9Z4J6EmqzMJHShzSEIxMdcGsKC1Qaq
YK+VQhomdV4I52/SNqA9nYMrRyrC46iI1TpiUeco7Be0IfnNi1IWh3zsD6qWP18+
kTkpHLWIwBK7hHz1sFq93RQzrmupVdl4wFqgoV8xYtfyhFscyx7KewjaV7FwHiLD
JG9zYuAo9xGTSl2tFOBMC/jVIXUj5PgNaxZD8favMeDvOIe18Sm2tFEsjxbW9xwf
OAFRTpot7oU6TFtG2mq9K6a9bRVXfL1Vyv74qL2wmqXe9WECaMsPNKnHqKH6yLqZ
RcQEBlux4JoohJeUnlB30frl3GeTPiMk4WOsDOGg1eoQakqrBhenE8NUZy+kchtx
KHZlFMz+X2pELw+ATlaNuYK1JGP3/rHFmQ4JN7p6QZn9B2pVCvBOEnPUpOiK7kyh
RnJjUNWUTXfB8eQ3w1BWXl7WwvAE2I6pPYIJkC04CdVojMzfothjH7C3VMK2RE40
/GXVsFcpNgiOrktCkzZ8q3+Rt43Vxpjtg5sWg2LCuk/1u6Bid/wbJz1psSrJXnKL
mMmAxfBbI5dhQyKNGnMsPS4EQXPX1yW1u59gwnqJHewd28lTsly+Hc4Cx+0XMkb4
4ng3tk8ID+5Ph4HH8IFhEE2SsAyRPobmvWEgnRJYpcVWy/H6Jlg4IW/SOc7kuzmI
u+m6Sf55O8toFQjVyvLVCjVs0Axc1REscArsn3i9gG7Bf4FP7l4JIRtYfVm4raUs
D+Tj6RrD1WMWLknR3Ipsfl11urtxrYaaCBqiRICpQYFMnDWKe7pFfnWnz/A+21BW
ej6c/fDalE0OKGr5TyYEGK0Vz3xq8zq7lGt3+vImwo91ekwktrxebu/Vf5NG9d15
smEALcbo9C/wBLhd20+idAjIMN0n2xqTws5MTXHtAvehGFqaGOZ1Vc4ejY6hSl0q
RDdCNmmoGHd6tuNToR8k3/VdVCkw+BegyhQhn4QUIwEupx2WymwPwgSH9wSNvyYX
JG7+m92Z4V9mzsLN74BOdNaTr03W021sYLwvwO3pmQkP9+pAusRjRv20uXttoygr
NtTbeUJybI1vQI9Q7eSZygff5Y8x7taqXCe81eaMD3PonjqIFxIsa6pe7rtRBwSZ
UpNqqUPM2nviIACcM0vxOpD6QGWzSX9eu8Yf58/Qk5K25RGZDLXh/p9IF/ZYTN2x
FYKgT10p4Eq8nij2Y51rQn0MVZ5M8K2VnqysIxlFaWxqscjbL018gc6+l/9/KuaK
CsnXuVIT8+P4FIsvNDQCtLYQ8hYnevikv3MvvR5nHcsrVSpEJGYwPrh7zFNUsUXJ
mT8748lYrFn8gPZvoQTIxPbrb16i1qTt7RPY+6d7TGuIuyWVt8es2Sh8plh/fUrg
VMtLoGzHqBg70pPKy9Vw85YE8Ghgd6SXkvUkN4rR9afdy8vOPKb5wYwF3HGoDE5A
jjjQwSxSuVKy7qpkKUqa/vZx2lKt62V+wNA/w1NKEp09Ch94TtCsElX1aTxMrQnu
gDQFeFrPLR/I3LmwI1r/UQOB5ltC+9qhmaTNGuVm5B9FMkvQofA905ESTjLwPd7k
E/L4YhRRf6cRq7Z6LIvosUdR5+hib2tvuyq0uUhW777dRNLW7rV0nXw1An74gooL
nkNRU4TbC1ncMtHAhq8bteojPDJlFa2E73CVVep2HQ2rHlhcXM5nhhPSuzvRW+H/
q9WiwBEAFpgkFLh7INBeLfg1ZifnCUjJAhWNdjVgn1291j0SUaQXs9RgApEQzTkK
xnVO3epN5262Q9e/y7YWe36W9jZb8EHAObDj1CpL3DcRCeGC9qrhRFv+Gir6nbF/
y72qpdyGPrb7qBoiUp/SC1TdjKNov8oGVA2V/oJXB3Z7tsqZuddmDkQ0HK4TSPsj
MaCUcnRalA3HcCVP2Kjt+5tAWSFlnKNz2lrivzmdztK5I0kd1nWxNk7wT6/lSwTC
0mIGA7Tnokc5UjXcO7RArkmdifsHGnE6NjPmdw4K35lEQeTs7PXFuA1LAfIwX0Ip
PaMuDmiYXXMGRFZEpUbiYN2kL6hB1cMcHKhZLgukRf9uIhl58QAq1RSHi8c2/G+I
tySf/i0C7QPdfvTPbg9DXLrbtgSIxUvmLjBckaWHkkKPfjxywCj9O+WIDrinX8vn
kDxfqY3e1pUKuUAmdjsO7S6RXCKcqJ7j2GtOlJDEAiqmGrG607PincQ/zFRLn88U
t8ANV0DEYxBL81sr6TB4naQFi5j1QWTZRHzcDQFGpwJSpRCWGDYxUx98rO+HBZZk
micUEsWZaOMmHhJlFvst7icZMfyLvk6z/jMtsez6SZT2idLrJMMjr4FfdsNyeISx
itbdwk2+HkLz0Nbet3z/4Za9MSRMJjRN3gsfXVolEzJn1rSVcrdjZ7oXv6NfewZX
yHhBRxBvvG6h9qODoiQV+CaajecfP+B/+408Uf2bksbllPTYVRx30Mj0PgMHltf1
q13O9UNb122YbD+QtZQz3w3x40SQw25qmOYvrzwK8weT/f8UfEO+sOLlwIO4EdNr
i+m9/A1VAtFVFV15SS3L19GiEyXWP3qDlXDu8IyeWWDbAKDOQKh4wN8UW7l92RWx
ZlUCaO3APOUjliZtNqutkF7BUnt7F6kopRNX1n8AIu8gJcVB+PXe/2iawYsAGFAj
i0ujyXBMh5WTUCkDomBWZqiqpd0/7q8qA7ZnKmFRlJenaf1ygNVga9EWSxoQZ5Fx
W5tLCkugfBVjVqd+gOySHjuF/3ghlXwUFU2KWxwULmHNg4uh2o1WpUG3LjPW1Xu4
Bd+TuXxeHonHM/uHvzn6pgtSq9EFjh/5DguZ/1zQWxlbmXsjONFLSxc57B35dekK
zIgzKlM3TuLW6q0nh9Rt8a9+YRwP9yeAyQ6df9pT2/7zxQ3XWgWXCWw7l+o0C4SH
JGe7PP54/7VCvAl/wTeEC2+Y5qtjg8U8AkjzatzJ4Zi4rCBl3NTxIOPKopEeWa7u
uLhz9DFgE4B0RvpIWykKbVEnRLjH9AY6ZWSHdiubLgiN6NVDCD5LI7MvGs9FPYCJ
4wIGrvzu8WPSiIf5ol9dnvMM8b20gMVwVBsK36sJgBuEKGaDx1hkW6hI7fHbKCkq
kxVxjtdmjITcVKmggzHeJvL21B0stBqhHHdW7+KO7vjHBqhyy2vnSb2gDhzmmyJ4
dZfNmi9aKrzDj/QfJzxu6O8Gc3Mu8fTovw/9CfMuKNJ7f8IWH0g+rTeg1IefgxbL
CZqC0pqaWwyNx67j9O8U98uU7/NWKpMhmjJF/0A8hug7QBI2I6s4IyJDzrGtQSWB
GcyVRBbUr3+jzyjTHaXfdofX0IQT8KOQ8J92zk2jmM0wEufVVA63bELOUeRCwMCX
5zP5svP2EL14DPmHkXah2KAknXWZ+zHujywK+YoQGZOntqMj1tLSfl6UyslG6T4O
XJeIMLUHNUKdOQqQiMO65zBpbWGVfr3Tki0ICRcC+ivZCA6N8jb7zs0fLBJfnbCn
QHpNg6n6zV7wV1rxDwIykPaOCNMJjCv6/vcrDNFdlJtYG0PZkXB37Vtw2+YKtI+b
+nTN+AFKxOADeNcladnarxqEwCDxEJ7P7uSJNZSQDsMsEENIpTlQdIe+JZOFuCsB
T80vSb3UybFoAn4hRTM693nDhWgkE2/H5tqMt6qkblobRQvX8ndHLIYs50RcVFbW
uN/XORjI1RX3kqmgHmgZqaM33crjRbLr5OCio3DCDvj1ngDpXJXNvEDRvPyFQTWg
sFhJsVP7xfxioDXVEOfUZ0OkaqUkK3HfOa+lJjiwQf9akVZqsV7kA1QPDUyLMcQj
rqjcvCXEUmDrWEgybksRC2djznuvdI+c6naNcRKs5TVv/zd4cEpoxJTMtoSy+tgZ
dSuYdauEg15wTX231iCNBUiISQ37OLKuXeDD8/n2d2tEkVOnvf8jzuoiG/VKOzk6
mmZ0A9fuWwy5nPblvUQtS7H0qxEUBL/O+a4VWo8B3ZYv/5HW5OHuZjeCgNrFVwCP
h6crLlHV1dVsGR4Jq210IsMYhK3lTMr1M2P13+Fa9QmuyfvR2rdAyXAXY34kaytJ
tIyCGzza96rn1iBK38po4G6aF6mGcTZ7c9yFkR3we8EsZ7RfhcxXUb1LElnqJxBp
O35dSEoaJqy4Ez7q0NcyYMYaC/N2FnHaQWxql+eaK+JrxLcmdWEyj8QF9zWli98l
KdTopyCbvr0KR6VWGPVCT3MiKT9o1mWvkAy4x2Fxz3V6n+iPCJ93D+kSg5vQhDa4
SPzTXtgJ4nlvvBPZElOYminPw62R4+SrvmZG8c47JoTeefc3GrOp/qMmKEoTwXn/
u6vKUB5+UwSt1G125Z4mqzRv9yfnxzNazwg4xzcQVlLKHCQQIKDrinkRoyMd4N5k
Q/hvjUkeprGHq6GZJLGycr40bla6CQcTIrJWjrlAoM3Xcm6VJxzoLkqBkC5MjUFe
KJzobsLo7xw2oEWCtQ6GEu/6MdzX7HCcrT6muEnNOfAc8N/+CFufPhXnk7rivNSK
+3s5nIuadyv9IpuriNBnAogZQZ5PcIRuvpk4OeL1T3SgsPa7jNPAxDxpM6zvzHhk
BS8aiKkhOROr1Y2Mk4J5/SIX2vLBkDZ8belCH2GSbes8FynJwLgs/POgHpe3WDdD
uKwSnaXQb96InFpsPyY0q06KBpHwRQkJbNnbz44pnhOTwQ25JbduUCywNbzdpck1
nYYmKY6xeClUGUtJhn49Epi834fkgi/7D3UzR7i06Bhtimj9ti/8JIFYICgrrJiS
Ucnr4EQgcKL7MPCtOwc3bagaYki1WPNTMwBfpiKnTrKnFbpszCv+z5N/ORPPoBcW
7HSKJBfw+XkkOmiWdfl+upKZ8cutupkWxgowTg7X8aMJyRxzcBoajxpmAC5yzzyC
M+HcCJhvh7FPU7DhBQx8/V2PX/VFHc4hi5VhMGwWujfZjGaNLPbjfHApO7mXj4h2
gv5+bvrqSeSe7Sm4YcVirIRuSvxBDTlwKNUPafH2xxRF/YEriDWmAgQ4HLSYG34I
NW+e08JlByzeR6g57dA2t3rik4tK42TdLA5WRb4qyIP7+1VDH1vd6W/K7sCfoJ6c
WtiiAJxm0yjrBX/TrJCQjzjM67XH1f8VieUEL2tVUjiXn9w996Adu6A55oV+tQgD
2BgppYFCm9lBezf3liBwhKFbFZ0wJ3JJhRI0iOAsBFl+rVQjtlV+XaRTQiu5qvXc
Z1xi8QwUY7O1noIRJ1VXeiQgduP3CQtOrzsoCEa6xr7abGLOSHGtQWAjMqkfdfKL
5cc9JrhKzZivSwxt3o97MyC+i4/z3nd9ZokM2Uziyc7pzJbhbVIzMQR4njBoLjN4
sIgBsEJRzGaapPoWqN7IE5zHBQ+c3cvZzTEUhvtG2vAFRfZJkkkF0RGT8uid5zHv
SstFAHHFv58RvGiRk/28n7aIuqaNG3xbMzpNgch/mkRPKGQAfnoZjclIKoNW1HJi
qgiGo8HX30sxeuUM1oA0kQNcnvXrqkoC0+2ytCz7ZdL2QSxkBOlch2/+tXNkJIO1
G8kgXmJoMoq1BE47ytOT1iqdHzOMrH5PGyJtP/yaIEOnhtagBxOvjnnrky2KXrwL
6bwt+aZkLtuSwUQrtDS0JdUkczFufTkUqdGQuEDc4e3+XmxktoUdnNaxBGm1adJb
R5cFnX2ebj7fuO2EtMlezvMeL2dDYfxSn9LNCGcljLvkWCAdyz8DRCFvdMbbxqgp
x1GxkHBOFrQ47JLTRGa3oycOg4alVdfk/CyjUB9fx0XjFiaEy3qg95cgBrFzo1eZ
lOIjMKbbwSutUjypi6qmrgesTqzWPn0vUsafrFd7ZjCFUCobn1yHfc5OWYTd9eza
27R3sjHqw3G8yL5g/l6MHmmca01hvZb9idlntLevyhI6WaS2hszxWx1tf5EMzegl
gV23aqjYpdcIjHon2evr/oWN8O+N3v/iKjb6shBAqz1oKAPOF462YvJJbb1mEruj
0egnkJHAaJ3/jVheq1+nKquk/knO7jHy2fskXjSRjIgFf7uAZPhV7BrQ/3pKxFxy
lpfo+YYCjbAV2JFGJ5uk8TCYiQ/pNjoveDhmZWuW3qGHMUbUGRgi+Ob/woD9At75
n/pri7J1eQHqJC3mD6bXZ787ovCGF3u5wM8CfRMQdyunjPaC/GvRc4gZq4jNuCZj
AUYIF+BdH87JCRVGIglN0GZKAZBMunanpEBZ/oh7pj1y1Evxs8EzM39BUN7jj5qU
7ygt2goAVODpl0fpE1Oazmcq50jx5HLB1Q4QuUwzk6fOT2EcMgGuPtjHVUyWCupA
BUL4Z+g7vxccKYSakQc1L1rfM/lslhr1MpzKgJPDjUPTHzKWMm+XM+QkQMsO5AKE
3zGLW1aouSlI3b8rZmrpVE2B2NXsrMhPQGi4dcKJKI+T3YHT0gcEv1K3D4vPHz7F
Ppm/hJXeBvr//0kzNRWZeRkgo8Wgx6zdFYnnMrdu2+znM6rQrxipQUFQbzSpe+1E
qQFqly6keEmBAUd5Wefj1M/jCVhAq9WW2CgU6jqfIXa0i2Ta8E/0g1PlFCM5Yw38
nH2sNisXolfjTEoowmtIC7lZ/kpUUzejvy7y4/NSJuxg+r7ge9ats2sfUucUURdF
7WGL6w85j6NfVIQDrrHdz9u/bPsoWzeelyjhF+i6rxR68quU5q0yUBIApO0a3hjO
Sq+KmPYA+tAXxFKt8qqttxdtnpYSKRZtJJKzX6b+atQjPoj24yyhBq1QUb063gDg
/hN0iSaehmQd43D96jkEW3/n498MHocsTIPPEarc2YLXFtMl47wDglkDxakKsoUo
T5ANpSleiJU2Aqy9VJe8YuDQ/jPtFtarwIiFeNj5PPtDPa+dQFJ34dWjp3vbm0Nj
WPmW/M6ooSsRkRmx6ushypiNxJ/uYmkhbAFFJJRo+YJ5heEu8jpUClbHG21HQfEC
b3HTmrz9NRf8kbDVhyj7QgW2+EbeivFRkgBvuEUbsvHOzQT/hhL3Dyo92b33osRn
lbFUF2zMIA4msTyA02+/Nz/GIf/MvNZTHQ8oBR/drdSdNkw36xbrrkg04SxYr89+
+uRFx8by0uMeAZoSZ1HcQVsx0c+MJe/qSg0h9g9M+O85xVArhjKIRYHp6B9b0A9j
MZG3HHw5XKHh4SSHSz5L22pOHCIEieOzj039lKh2LOCrbrfEC8ZJHvq4bqldG2A0
rGv8FFABsZFej5h0DYf+3YNQR1JuEwjpQpEIfGM5na2CTZTwpDPvGljqcKdxoPLB
tB3DV3+wkni39rdea2pVZqJGjdtHCPqBrosS2cGjazuMdu+P7pFxhQ85aYAWySjU
ZtLLdIk+u5Ahhguqef8VXlW1hHsSbYjdURbMII5lIQ46CbUqGoJg5jbporX4a+RY
rQPOeft7NdZ02wVenCKVqGRJcQbOFRbHHXaX0QOe7r7rTIjZ/qj223D4pNQYYZQH
BcvcDEk52nZa5cAt0qVhYpy19vxF9U1BImfhUpgm6MdHsbZGExiLm6VAsYGxg30h
LY+M76yKF04XVO8fnrwM06DEjo2xGQ1/HAINbvF/Gt9OjpzsQv6eYUE3AhbvZuJB
7PlrAN7L3F9PYd7z0mSqylu6/mLRX+916vCkST+R0qwdNEwBst6AuRzJ33Iph+Vc
az5KS/CMessvud2JuBeqdoGwnXV5lvKEKyVYcdnTpUNYdMxTvS8hd35xM9jzZLqY
5eH7O56mILQVFPAtUixBSrAgd9Wj/bLlb6RTWs0jTjRX+GUcuWea120qXEJXICx1
xqS1OHES4/HegMBr+tEtmqveL2/BkQDC+sesgvpnpg2vmeqWFQS0px76G4bzh6SH
UyX5H16LoC+K9Pyx/n6k0jRuCbCWGJSRQSpCCHjKsQ59dpytUNV8UmTveyxeXiZ1
Q0D77kibZCC19RgOkFpgxL2087Cbb8pNjRQdB4MFKl9EFmq0IWCTYe0HgYjtSXzE
x36LcKNyApDVK5Y3EvIyZxc7sxiKZC038FHPdeJwEuS7g1nkBe2miy07QSWCVjIr
2RZMTNMan+VDdMEbmQWmGcIrzhrDKZrAh2lQrEKqQq9V7rNbtKgfuD7v0p3URDf3
wtMftIetanlUPPyz8JfRvZdDteXtvtJVxAZV4hDbWZvFT+jI/7Ych+yNByP5vvs0
hXvkJOhLu1OTV5BjJQMdmhBEYu1Hz1GtsgQ/V//Ar6ZvTafahe0dwk3JAOQdKXbQ
Y1BQ/yhpJb8lolHCGLhvAQDSW6JGVe8QrKPOfkV3y9uFjbalDJq3AY7AqssI93rC
FwJ2dAr//GUM7Tsjf1QAIs4xh72cmgpXyIAFQ7UetJQ+wY1mKfZMyz6bCV+6ahfZ
mo+yyEwPz0QLi7wmmshvT5ucPqo9biVBy5GX0O4hrg3Utx+tN197NizaHMgqidWW
lF1W72T82m0LU5tLlMiwPbXRpQLIjOXRvUiefzBSZgmxcTPGpy4fmLa5X9gZmTXt
h7K91TqEYwbvZwhj+HLz82HmGXx8RaNoRtwtqfWitouMp9ruktEWdL5j3aeAsUGX
F+5H7fG2PRdgraB17EFxdfhP5M5kP8mVzALFU+DUIoxJBLDBszqlx/Uf4xoZUOVj
lNTotPSxVB/hH6ec+5Owh9l0qdYe2QkXktpsJDGIvSZZhJr2OXou89Gn9yldN+F4
0gwmPvLwhvXIOPT7zw4j5RMN7q0owQyZdFuYbbvhrI0KvvbvfZofVrwpjEaecZcN
3T8uZOFWh4sTOYo+xNNiL8O8AGJlCcOhjsPfrMFK6iXXUjcEk0zFWCALu6rwXfoS
ON8NRBc6rMaJZv+hQcyxE7xwZgkQlF2Az1/FLm3AInOmBGYolavOKbYMDSNt68+T
ImsT65xb1snY25BRvUwS64FGx/1k39662DgvhZJEBEVnbTQchd8yGIOgEU6BDFfE
wefgeWHxmiib3no9z0jFApjvhg+EW22+vjAYLJO+k9SKhZtigw6bypoQ5bVo+KHu
VmZqNhH39LxY51SsWuh7PzKZwzFIewSgUGFZ9K9k6yd+8Ori5JHNe/ztKj16SvXA
LFkshRn5AwfTXUBH8uJm8VNIV4Kl+hX4Pv3cw5mIM33EeXMdV5morkDjn3o+Mc7n
KBUvtUk2gefuNX9nw94nk4XdR8U4fLRbU+D86+fXRGQ5Kr/daS2bIRw8/EB7u9Wb
L2rPSIFzWA6dbrlBq2Bb5u7xMosOMWZ8sqFExZliNZtcyz9h3mtZz4n7Tt5o+FYE
YnofaohEU/ccLsZw0F1vOAjU1Lgvuqj4QRT57hFK5F0RUa3b+8rZffUVL9dkMbX6
ilPbAYiMPQGbh2yxbsLXKM+xi+qmZMkKj4eSITsg3Ma2B9O5rlBtBlVU3Uh58H+J
LCS6f/pQq/7LoGUNXyhbhGrLm9NbVfrjrMZ0sLeQ+yqbDx78UhtrZm1WNFA15wvy
YeZ7J2H9I+T046gEEwFox3LVqVH2RxJxjOozGMGXIznSrnP4btBnyeHy7iDygVCO
W10fY4G3fP9JAzkyd9JzaYwfTAn1SthozDVfSdWI5kWMfjhvVQO7x3jkkOSZineR
tEzSTLXHtsjqFo0xO2loGEdsPt1HSRlsx09RxQSuY49KxZMbCg85SnFu57yUlOal
95nt5UvdQBBpwpAOpJHViBBhauQPqfVgdOs9cAt/FUUiUzMOLtevOFbI68UeaNmq
lVRHq4MwQ7ZZFYhKAMD/vVqT+s2MiLuEhCcLZjaEInx/dyb7NG23PNAN9OEwxITT
+63Cg7f3yRjGh5UyW+bRL/HxEJgtfUJWiNCLr+K9feak9s0FC0z2VNaayN2+EK6V
a8lgbVC/1Z54KZmto8RlkCWK75pTpUDgXYJ3qrZPPi+vVJP4lkIoKZZ7t6smhphU
60WFJQ/P+jnAfCe/J5VuFck6UDAeK1s4E8UZ36I9SOb7B0KO2Ji4diu54wi9jM+d
rW7xXmWpQhUI3b1Mb0kzTK0qrKmeZ2EHyf8RueiBLKW9gK6ZHwAbg1Z8mhtklyVm
aa+qArQIdiic62UxZKdch0gLXp9GwglOFa6M4sx50LefmaAtf25nJfhG04CCUkz+
BS5J4E/OAFx4sseMIDjjJKU0phFTOUtgZaVg8Nv4+jVpOl7jSIp/QZZ2USGUhfG7
eBK1+QDMxfVdCfsSZ6SHZcjK37PdD1Fy1n4N334iTDdWyLIcjriXgKnian93PMYa
UColdio8eER4EOSPShi8sigrxGiUNmlLdx2Ku7u/9cx4K2icOXZ1tM7KF+UH5fS9
/o/CnMMzUUtMyor7sQDq2sbKOPobz7e4R8kQnhjy9LWt8KgH42QMIk6CD7iN0ZH7
U9s0koMLd2cPEB9sUE3qujPXjXC5Jnyr0ajOS34lVgtLV5KGYncPaFjQs0hNqzI1
wE13TlhDhVGY99iERapcIu5x2mOPlT/Zcj6id3OB5nB9yzMNTWyx/IGQd/+Ay0OJ
TLtKQFSrJA7CLnLTxfzt5zjAU0IIItV4WjHAeykZeHNW5UL0/1C/bZ7uvsy7CxSz
b0uN1SvKnOPfjmzNCYlmntqfE1pA8SfdSrt4DjeQ1jW5i0ndE2dLVzIThLYCX1U0
LDC4Pd3oR1eCl+KMkKc67lbODrEKLDH+U0MdqXiHGWq2qUCFBsgZPG5jRv0MeXxv
+6xuP2EWRCd163GeMSr/9ad4aTFGgwi+m7L9bdGCTBxFvLp4/2ik842HU16BAHP2
LMDV2MLVOSKkUaXjAGJiLgKBMZI6KCCiyhwfJRrR7osV0k3miwF5DzxrAv9ipqIC
YhyucqxgaZgbrbJQnWLLnLnTggy7vyc0U+ML1FCjlMeCdwwk5UQh9e4x1RAotBCz
SxkDX7cLAcTmnsDrHFGdCQz3GS5w98i53Mym83FLtGmxfzZZPfvt9iSSdMChDAzH
kn2ChMXc9FGcBu9/BKkY+2B14WxPEOjF6hLMmp6RKcll8M+VPBCSWYqd0Xk6Cb15
3rEQHvuMmn2ItuIjYoQ1Phk2QmLSE+UXrUlg5WQVIHUOOzGeZFyH1UAzOzsstlxf
wOlrQbMRwbVpuIQTaRoVA+gl0jgRw85PVDneIYJQu9iPWzutnRSJwjX+PnY4N5ko
yxDHKzSHeGneeEaCXMPc/pc7+TrBRHM9RKvdcgFgxXGET+L0vdMvIjhyhJP9XY+U
74oUUeUW7mLDAl6G4lL5y0Dhz3smvefdbaMj55zswj5zp+FpAuIp/6cIGh264dK1
fJSJ6dLBVxPlrdYLwKkD5Q+tQofj1fd0cZca86T5veW5NSNWJ2wkC7ih/Zh8mT24
Ds7MjIf7u7CMwXnwdq2NtzbQDZ0GWo1f6OBShFye9GQUfwoK8qau6GicUvJLL/Dg
SIlCZh8G0pstZUrwgEyzQr8Gz7EZm2dG2bMYw1jUfPh1/At7bo+4pkyKar3pbJHM
xPr8AuB1uohp+WHKiU03IdO/2Q3VzCk3s4rKdboJz3EM4MwoV0EFBURUikUDSmF3
3bhmHr7n74hRGXyPMDD36yXibo/o4FaE8srKs6yOIhGLtQI8Az941v4fJ3HP4t7k
XZ6vMqruaGPJ4DqbJfWP+SHFtZp36WYSoNJcOfjdV0YnSz9K59T4dHzSRMuNnu2z
3xB2KGDSOj/AND23jYWf/29apQ8mgt7TjI2kwijYn+eqZrXHiHNStXuy5mDSzd3f
HQMqQoQlt4SctgKDrwuAEY451nKNMIBm6CCrmpKH2poJgafIk2SAAmoWuvFAQq7J
CZfqPDRLOPXkyfPZglAuKQDyBYYwO1zJVAY6J8pz4UjvLMTa+2Cb3epEvTnqFj/f
8aWgzaM/4T1EeJDnKpvIs8rwKm5x6a83sapp5GKI0sBjGhw6GqHHBPlih6qUoxUB
FpC3d8ZVEku58mqLPIHbh86Zo1zBC6CaCWQEdA/4i14DawHkKgsvS4RXOneICqkg
F6E+v2EWm4e1N2bHkdA80IZ+RDGwFyoBYKDQzGaAgteCjqawGcOiwvuTk3MR+kW1
mpG2U+7YbjZAvd6nFhypkys29Vc8hQIpY8B62mYJggQOgMHvkikgx4s7o01lmh5G
kWn+n9sNWQvFDttNmXbh4Ub0W0NT+lpl84Z9u3h3dYh2GV1jXM/7rnR++CqvUVbX
V0G/UhFcejQSr123xlxFZpY6yMM/uu7Nivk251m/L+/ZAccN/byoJSeaj7tzL88w
nSvBsiDYe32zgDUbDW3a7AIfRwVbSlOvqwygi6+Z2B/I5ut9YBENOadTuMFXpB0k
1JKVOTYUTZaeYI6SYGSCXq7zYhLKzlcy7wnZFJ2p3KphQp94MuFTxO25tBDYHDs5
HPPyBQO6ipCiREL33YUOHjTRxbKZN0QbE/Ix2ihkDtmTk8S+hgjLoRtVGtNzORuC
ahn2W6cV77Cw9+5mx6gYErmMgw1zo3FZG+OrMK80o5qXxg32SgHnAQUO3k+ncsUr
pJekEndS+KjrSqEZf+ZoCDTspobQzzCetvO6bbAinwYPO/osjyXuAmP5p4oVV0uS
eRv2w+YwXB7s0FIdB5jzbRifxWYu8GI37DEEC/y07KUdYgEwZ5T1tek0CCbNuXGn
R6Ex+UfI0Y1sIhFBgPgSF5/Gl14BMXD/rwygvWsTr05yX8F88ynUTBe9VFhCbjCw
d2z/9TLGxA9W/EjVtWD6NG2mQjXenAj/7qalyVas6adXZaMWoWuGcIa3u+TVlZdQ
SpBnUaA+pS2CzaYlNh2/SheZW3LRAmsGAxP7y8+P9XhkblpSwkkPMkDppaHkEy8Q
fNGLg9oY0HJ3TWe8wTjiI57IflnVQWgEeOaN7tUNitV2ph86yDbBDngeQmaCR6da
ZZp2fnwawidY1m3914dy1odsb6PL6i6+1S+QTKZMXJFeDwjSODfCexBI6j+T5hR+
QG8z3JuhI/EHeD6v+7SJDJbE3q03MRXPJKTc7gwPofMeCOfR9fA+D9mCPB7L3c+r
JSqReifXot4CU8PVwhEIyEMNBTL8S3kUpYrQl+M2rQYwMZeQ7VgxEoy6bSGMyQIl
6ImWuG1rHeIag+DcLMiFoBIHPnEX73k5PnTyHWBUZnNbYbfQ3V6dfPlrh59GgqDq
pZtGvEz6MN7pGwrsVRj7iPiRAJ427DC1rzUf5vYGZTJ4Xxuh0KNb7phsqP3VeOVJ
XuC+vB2eYlqmKQ6ZUJGPpPjVa7yA0d9xNJZSkmTZaRIxZ1X8tPThs/UTEatkpkje
GhqrxBeX9D50SHHUAsnqE5H9wXoI0P3lncXhUP7SnKKYosAOLS678vUGJLy+wCcM
j7R32UsU33MXpw+YfOGAc4KHfvYqOTlggKfZKuPsinI7kL0DbYaniY0SefToLEGb
yaacdFVQ9DD3DXnLKMTwA+lqZVleeGg3NjauiCigrTunX1Ax4pILx3raRJzL8yP7
IV5UmaZoIRdqHH/u5asnG9clcoHT4YxyWCz0X4rnvchH5p9LGhmUgDqN3kwqmjkM
lilMW2QgjwL42Mfxz6zdEnxK7ncHgOsYh5tR7FOJpBE/w8JzlNlAXi8AKJoj71Mq
rQc1rofBW0tKxwAJ/YCBuPNF9QJTC5jjzrKhUbej+SH05hmnQAQi0AKpD8Xe9SDS
VbXqY2kllsxoAUlHsR9lAFoXOfmk5pTfhXyULfrVIBnR+jO+xzlxEBenhd3cqem9
sbsJRjIbwt1s8SydfNIzyIzWdNlb8Do1ELQSoGVWnB2W+MVViTK4vFPiKaQP/+FI
kk6cs81rMUrXcbT2YTA328Pje+/rLO0ARUqkQvrQ7hIwh+ce4CHJZyuFUTA6jEOO
tS3smdDi/vfz5+DXj+c0wqEgxYAAq2BXBjxbil89vWIa/LDNPcX2Nkh8YA/DoBBC
7l9szA4azPae+5CIsqtQXZHxPYSzkRxaHmXRmYq5ApM2F2Nxkyi2gAMzD3w9Z3sT
554uxFePgAkzWL0iAo1blrXVLgp14m+3iYEOXB6As/mQ43kWULwTaQZLAc7FTAlC
EwY5nNh6AZWnP0RNTyBzNduJvkGF+MCPJdaq9zY7TLWYYaKBSh6ach1Fg/8DKVOI
yw5jzfGCOqtfYYNfhZYIXFLT1glPKhZK0F2vxHStp6ww+HflXTBHcPqHEP48Xcbd
clqNMd0qQvQJVw+ZGtUzzOnt1ZFGWGkofVYLIjhcTsJ8jrRaqjOQ1/vmIPWnPHGU
cj4GiiDuu1MMx5wslxfgG1yPBEPqU7YScKVMfg6/Il6JBrH5iVByVkI56VyeQePv
jLf+7iC5fc1ppjbWo3oZUYA+6La2wTBMNLjvno4/7AXHq1k+UVm2SXb0glGZ2QZj
9kTbZ8WhiY4MhXfRSIfv1zmAPFKBJ7gdmgoqPTCguqCM0I6b+WgyOHy+APFWHNer
qj9WZEetAiIFl1seiPDRYjCXsnKg1tjbiU3yJvDDO2ZPYXlM8J0vaub2lqvrXgNq
+gh1g57JSXUlgWkVk26bkQ47vm3xaSM2aNzwZ99dJYFmSbUAgrTGdkRGXJCNNAg6
LYqGujHaPgNlGC5dfPGO3S82gvWA/2auoyrwoocCYz/1bQGg+4Ez+Q05ltMgSwuy
3mhpJEKsZ/Jjk4+djcLv+Wta/ewJ5g7KuQcLHdZDufCbZIf0zbNXvUcQ6wqPM8Km
+DD7QBHnTbJ4/S7ciHl5fy9C7qZkaNqjezVBY6RN3DjKkY0/dD22uSi8WtwDSWf1
3343HF54lRMWtSxttq0f/AJQ381nZT0PGeN360oM77spCSfKxq9NsBKFUhYX7Nlz
XtjNCbFpvxKizCmZPdpz5yutrDT329lWtlkYxisN8N+B3hYt/qBf1OW8ZdiwuNqc
yJoYA3Yafd7QTNIX1yzVVItylmSRc1gC/NN+n+ooH3OZafmcbF+cNtWtyFQUh64b
cePB2KJU663ZipJ4KzwoSMCVVdSn6M6wPG/FiQ/YTjKGqKb6x+5TWOF0GrQ1fRpG
RYvSYa+2mUX4FyRcE8Hmkr1rsftSXPWI6Yh/Y2vCqLufTUv+kMFkg53P192tj36v
ZNu07ZBh4hgI2liMt1PHxjMJvWrgHCYRem5QiZHCZ0dJ7PXcfAOI3QDm4jLWu+3D
l42vA26OgVvh2SlK3hFcwY+ZWbpQNMnp1etTzWqMq/ihJQsxYLDtAIlDPx08nFJh
pef1zfr8H9O/gu8e5+lZcGOwNe4eRVadVhwtn57ZZFv0RHYCFixwjLXUV/niQ+5h
A1cG4jd3goExgTAaHfnVLTVacyozdvZ1RGZ7T/8Xv/2atzzJqd9ZiBkp2NX+sKwY
z13KnKu4tnGm7cbvo7HRPIDQDJVEnlmX7l1+XkaWwG5/L0cRIErFwZ0rOZkk5jYn
jTrPUqedQ3J9rTwS9dCxARcAzaT/zpLvP5Y1S+K6qREtdxxR29Jbb6rwxM6pATUW
04qfwQAtoyBHiUC6AW2RN7tD3Wo7uoAP1+2iUyFLBVmY43WCtTFP07B7uc26SioV
9T/HLMqeK30gDUesUSfDGJDkj/iizQSSF25RjWw5fxnTgcVbHPEfL+nq2Ii/ohf/
hWZ9OqE7tsMdvK91OZaL102p7Mt5SVDE9OtxlrQ2ZBSE3UTaePwdbmO/38RNmC0V
4VoNCII9Pp8XaL6p50Bzyx1USt0LRJrhgGqbgl7LRVgSvL4ScJBGm4Ysl+JbreBp
+PWA0HX58Dfx3DOurmmHm0n8fhjT2scUky05Og5ow8Q6TTsePDrC/iT/uDkmaHxc
rLxei+r6KS44AVZSjq82oGkHvqocyefrsJf9Je+VS2Lzm9vpOKqYXez2GhCenWC0
sDYsC6+6HDVBfYj4ZG0oRQZ/EkiaxUjutBtio9NmyqYQPvziS5RCV+jBu6EmjIoT
9hSYVqISq/aiQU4V7bhCKiNclNBm0seFYsGJ5fBO4MJfKWcWU9aZajfpSXwVUyH/
CnB6wHkl2wacZ4QXRPKEdbJPMArUGLmUvXC+/drpLv4+ESV4obFYwmRreJE7LoFY
M6fcw8Dax5ey0RxXXGT//mu7R9BIEJA/qSexrGG9T2hb1dSBF5ZGjl45T2X+foOp
hx9HAMXjADlA7sKOG1qhGClrPpl2G15Lwxw4+NXXxSrALIoGVAQM0mWIR4DpNOeq
zktyPcYyCI+R+MXFst3OjmD/gtF+BM24kvoNJsW+gSXJz9vH/uw2FeprWpAgU4bh
y4cf0gCTdNyz+SUkl0Yu0k/hx7FmMsaEJ3m1A+kXUtsgUWgNN8yzjdO/ZyE9gQsQ
WNJU9uaVv6Amp154EtBzNk0tcSUGT7B8b4pgj27rzX27Uvjwe1WvLU1gbY8vhJjs
lhmYLSP7k18jmJ/eWAoYS4PXeDdHfIOUHW5tzmcMdODzTqKFLcpYagycODpbI37+
ab/s4xjRJv6MxznGKuppAcAS58EIft1ezuw5qnGDfAB873ua7Ea9s+haDz2hCA9R
dcgRur21GoVc+F3Xk1OrBxIbEQrKc0VMt5Cz8PxKpsXyGWUaEIXwcvOO6J1w8UxF
bVQ2LHVgcctgX3xmna4Ldf95+Rr3qdYloaJgF46JXBuSQmPlaQqovm22X170CWHP
Z+UgsBEhUxuGPX43eNnYFFbESk9SXHQfzE2H/lBgaU0tLl+6euz6thJltk8rt/uJ
PWUiufOffir08r2alPvCbp0r7E0VmLjKM35T07IwsxyF1RF9rF+AwvMtcRpKd2Fx
DbdYUyiNwTi5Kq4SmwJ+394Le9ETeaPyRXhPVhXF7n/LHS/AtYA+vSxvHDkvUmMk
1XYa8R+l+59E8HwLJd77MHV5xXhuFiMzpsC6Bi5g8BzJgYyEWBtL9x8rgXGQzn/g
lkTdaBxuj5eNdJoK8MR0HqIap1MR+WrN/8kYE+E6SRPbbK+3Ib8fiPsOllbP2S3G
tjvfBYWSypjN7+CkEnf4GV1z3vzmKJ+1DqRpeoaR7ADnLQgFj3Tpp2mYkf2LMFBM
aKcbgxBqCuXF1pCzFBj89pNa1FEDvsZ/44BCQ1znt1IfpUKn2Bt5OvuV2ZxyIzAl
OYdVEuV6pHXI9ZN6NBQMJbAPLSjd2EJJ1nm3VBVxSA1U4WEDk22U78oum39ozQgJ
PIVJjJk59dV2NdgEXQdbVRUkDLvEyGq9TDYdgnEqwaMJ1qui2/VFFAd8+hLU6hsj
55EpcCz3vM2sWQi/G6VrvPwXH10F2slNvbygf0k97ogDKEHD4jMbASuPmt2oBpae
Qjy23LUpw7PtItPQy3rwbDDmA2jGMgDI662Rlpgp9XkJKdsvATVLbcv4u+wRCvVm
Ga/P6OEzJPuOHfk+miPkWNLynIsbgiQqgattRPj+c2YVPIbKz5LdpaICA61f4xL8
fCyUacfzOSQ6zqgSTBlPGP3j3Ww5U9yldZvVFhPd0ViQSfVkTZGcTAQj1SoLgj5U
y6wI7IjXODD7mDRxcoObIGkWVJ0/4cIj2qj7HPPGyQ1yCA0AMqfLqyDfWWDXBg9B
GSnsWyRgPqySBrkPtflG4OBC3OIqc2kvxLriUPP7OEHnafARTE2MkgDVHJBTyAvp
/db8DV6eab73McbadSHcLiw2HyscTEucbp2vx8OyZo7OHKASuxSOVvsFJC3/dwcm
OL+bHrPojf1PVZQm4QDUiMy9KICcuJ8UmFZsePGfq5gJ2vu8Fm31ADNk/kJ0Mi9n
yv16r9Zb24VIb4ytbHyh8PvzbdWgzZzNVQd7RSBjMou1O/Uzp4jsTA8PWcABUR44
KmfnXFqYO/21VLkHvRV5TAJBBMsA5WMp44aYv9H1OBl6ol4bWrHZpdpxe0tjvboO
+YHT1U6L9gtrJX8r/yaDNKFpfSgwDBBpgHAXFQhoRKmpKc8vT0gF9nslH+2kXYlc
Up93c0hX9H6uvJ7YoML7ikZ86NTyosw5prVnz9V6SZIpfuurNGzZdj0vwIsgHdxm
94+VMlX5uvOgyF0zPoP6nu9vG7tgxUuyezqR1gfX3e0+QX7qbOCXoLlfoVZ08P9C
wf0pQ2mpTBh2eZY7CBA4Ze28b3K5u/i0rDDv1Qc1HAWwQvS+47srxScP2s5hM1pF
7FOyIXuNy81mTRtFVecmuDlg0AE1nfwbFKSzGSZgPYSaXaMdpVrP0gZr3l0gsxXk
BsGvMncjHRj7BAorxsQdV/Ct0vIHyGRO8xU6s+9X6oDNYVyE2y379EQx47VjISy6
p9RFMihAKdC220tvLTaUW2Y7B727o/5ATYLVklBHkjngcmtPMOMn5cGbENsnBf6n
buxU7siixgMDVBOKiNSHJxa9UdM3pgZWIYWlqhKLWb+KKvr1LqHtBd4o5yTsSBvM
9jGtGGdrDuaPD3IQV2jFUFsZEFOPkaeycahCvYZqIvQGgqD3Jr4X27X+s1rnXqt8
AV7m9iSIfTGK0B246VkzCp32UmMOOci12UWBwQlYi/q7jQPhltmlG9dUP1+O+7OQ
btVrnsHAFcXACFDBxJr2S8YNvxgmEUqrt27ejup4d2JpK1GUsgdUzZYXeZ+hSEXv
oPRjo7TFVCHfC/xGwIdskWuK2Xyen1Rg1KgnL0JeFbXseWSE9BDCkawBgXuLZvGL
Ckvukw3fPBHqVpDQ+m8e768BtTAKqMDvxIf8Iyjk2Vr1vDGpXyTbJ0eEfk1NiJBj
MiwG5+zFGzMOl9UQVMz5Oz1/+mLXm/4bLgp+Yc8KSucnEZKIkvFG43zbQ4WxPp5v
n8YiUVJF9xpbDSwNUBAJzGd6s+EWZzQLt89MRUofoly5DSLmau3+eCoC70Mho7g0
7Fvk2DlVp+gks3sZuH/n9JMjP1vRMGQsrEl/QU+LMPQwCZqQ9GAhhlmoDe6iMh1N
ZKGLiu3QnBXT0cYNw9goSnVyoTb7HaeFSk+W15Cl7eMSLc6NjB0ZgBrBWeVEf3yb
0n5s2tAOw7rNeK9aVQyg5XlCeLqz0WFvhhG2mFwWc/Z1nJ2QwhPTmE+jzEue5M3i
aXOvQx1YAWWOe8EIfggCqpzO5ge6J+N6O9Iu/r65FbGSn021nLaLcFcUf4MSxUmd
al3lTOrjgSfyexq18ILUenCTpA4X4fCzX/Z61klJNcCtccPBE4VokWTon19JOgBf
RDUDuppP71fchVmhj3hegX9bVZd5WCOoLP5YdVuGYzXMocfWiUPsLTSyGtfViaKA
MojkJeP5Hrf8rB8dapju9fZ074kF8OEC8fGxzI6XiyS2o36NkXCWOHOd+kS89j+s
BRmCNQ6kmvnp8I/4hClytEYNNSPz+yZ2vSv90UxUDqEBIij3Ym3xyN/xa/C/sOEk
dcN5v0yKFcuD2rmfFgXU+plqfnu5glnm9A875iin/VJCPUwgNsZsPh/zmK1kudmS
Y53vF7fMuKHv2S/KRLt2q7gjr++zwgqhfUoHkJOv0nWKNBciP/etyPEJRwRroRTq
VrkmjWbfC+g+qkaZn/XyQaFlGgh+zFgkddl+ocTNS7gyX2C4vAQB9CSQPEcrdX41
Gz9NiER44Jal89HEL6cHs4d4oC2Gh/a8QfW2LdTBPMJyzlolBTQkLXfeVdK31/Wz
4Z70pAiHq12xLLUf2EMYN0YUpVgp6marNoYmopky6yphXa+qHilomuLYwnpIHH5Q
9nEAD9LKP3ejBKzWiK/4yh54lWzs1Hz8HFP9vKJ8zbvGpQGsZMrde0p65Pn+ivLu
OlA7ITYBXhKUuu4KZOH6G2b/OCHhNcF76uSmIKbTV0D1rmRBDsA96o4M937o5dJk
hiZLwMvytWFww6kpEA657i8wKkxBbjsCD0jwyUeozvkThhIgxygA6iHqKePZLbMT
MloCdq7JoXSheS1LHsd+vNrMX7rehu83uZvM/T66WyZZEsf27MdjWyRKZSX9qsyM
CFKEIzz0gDo60DVCWQpFdzHcsEtgJWCk63sSh5mHW/sWYMnArbNLVNM35Gi0Vp6r
JoXzM4W/t4pmLG8pG7GXuaM/v+1e17bdwFYnwdAWHJphIeCzf6SWckHh7WClo4AQ
6LuZWGQCauuLrarKgVy4NNkX76yT6IeTdYUUq/b7VVZCfhKJzEUxKjtW+erj0tYl
sbolu7tHOllgQXKs65Hyeyocxr70YeiKvvL6vnuHxKSlfKLE5dUYZcq3TUYe7wIb
CS2ES4FTb+wLfGHx6cqQggygH7MQjgWQkDit3mbpo4o3WaX1GYp7Aop4zj3mH+WK
42FVaw+v+Jw9Yeag56IQfqFzBVxc99G9Qe31eAXkn5GlsWlqWBPERmMeeHo61JZC
m2RfHviClGFAEMjXIFNT+HmtNQFo1bam1RpldDtb/n3drrW+QK8lvDRa1g37wkdj
rBoJa9G0rqLqZk0FJK9VzaOM+B8OCV7uftnXI6F+ldgnXWpnU3jSqM1vFOftLJM8
ULaIyeggr/86lIMx4NXBYVnVjAz7xsOGBVTqnMYV/GNU9JGt4/JASP0Z9HAhsEsq
CMbn3af0ys3pFItPGKk/n7IZPFWkB3IW/DSbVLrYyCvi6rn/t3kxeHzZwlG9MY5g
Vg/aIhXqHuPQH/MCRg4bC+8amIFQlCdHcp8ZoqHVX2L5iy+pbMHlnZ2lfBw6oOEq
vaxBJCuOWyG11VP2Y/nWP6YEiK603SkadxGZY67gY6GNFdnUw1QtKajNkJWpbfGn
j1+PYSwC4dThxLhzQt919YDjG5fD3O96bRhSloBzJjhyQNr7QZgwqENnjKEx1sjs
TmuwcKgkdjOgsd74kadg8G/NqV4fJzaDsOvrhkJRfhGBWl2L5WU/yV/ZRZXi/Y4A
29wszASPO1jaVD2MQOyBuiJ49rMzjw8wjTd0ADUJUiVTOum4o/ED/HqIsnj9Gogy
yU9L7AZ6AvHl0jE3YPgLDoyknfepyH06o6mokiZDaBoTNNapOj6taYwb4G1T7S6a
9rsmqeIEeK++VSzF1z/Q/vDPft9j1mlnbcsDasdy3aTwFpVIok3iMSkqi88u7Nuq
eDLMCmHibGVvI/D8WHg/ukAf4HmTdsWZQvosE1uaExGeAJ1IIWvbLupEwO5ACLKF
VeTD7/kMMU21sIUJoWeQBG7mypdN4+NTmrBzQlTROxUoFVU31fb78Pa8iRKwn6Ik
1kVuvcLniCdJNrkM38davGiumxriWgqcXfghuwvZI9N+pZRLoC3RtUXKDsJ4PYkA
xfIBUugRPGDizqz9LA6pCXn9+4AuRMrFLB4vT4ub/342GiHwozdGy1J58fDWmdfT
pwfJLPOO58OsRNS9uA9MqkpZAcIQnsXRXwJk/j8a3HT2MPrTYGu65DMPzb73n1xP
iAjAhuOGwNwLfJGXzhtmOYLDs49g6x+FT5GSHmedD6k/+thAhQe+qTGSC/03Gb94
Tc7JibsyH5aC7MsGR52pHLRsLP9uv+rNbGD8XgncWyMf4VydqtU5zb/DZiZ94X6o
2nWVTSsbVhGAbGUnE3pta1wQOJZdUbvKwSGTlJVHCgPd1sVASpT3lQGRQVBrHDZ2
Tx/aAoty5VlJHlS/vlB+84xUaISsP2wnkCJBL6P2M3dz32gjrqOaYCqRcNwXl3cz
dvYQF15GcIw13VNEpDz2basLvNdG0rgWQEIbqnbePYRglKSs//KZU6xZMHsVC3h7
+tRWrAe5CZ0I67Yt90Lt/DKW5hsy9rQlEwHH7+hiwB8qbdfjKN51noX1/XMVjmSi
Nfrt2t6QZtfvRTL8xrfpPYvHp/cKz60xjqZZXqe5zf/8XOnT4ttwVbhPjaqbf710
a1Q2RPXOQGcfddxwXdvBCS25M+22QoKUsQZ2A3wBCKNwyLmOSad1Bs+L5sBLCvmi
pMhQ4ZGEmwktaulFdAQ38mSKavdsB3rllN7aF0YfSdDGN1rZm8crm+DK25ry7qDr
hbymV+OsdEADxRtP3KHj+B2QAoLQyMfq8ODmnEBpVj3bckao9kI5xUHVsGfq8IC5
FMk2w3VmYU0MTJPRUEVgPDh2p1EhfKmYffY3PTt64BpH1bQis17f+IuARxGI5Iux
7IwNK2O/nwvYqnyX/nRB3yUeXX9P9ZNC3BF8DNwMD4UbqaZvF0zdzjXFrCGVTEVG
TLCKUX2hP++2xB7rtuUYl8GYhmB9lCD+M5ew0y6PgBA5rWeIjzttlLq9R7VumaSZ
gFtBDaLVIZBZVpfacwjTB4uMFbnL5mCtD3GMSN93Zr+96IE9e6JfOXOznAXDRMML
YvIcbd9mT8ZBFMxk/cKi2scArhQHOzt/fkbf4VTtdG3lxBSQ4joK7hHJJsaAbjqd
6SOBojCyjzMk8PrqXVPA6Nc5zaZ/1lXkT+XcoviywqRazBCOKG3WdOgi/w4q+OUH
S1T8QvX/p1Wgz6JcLLP19grIeRa2k05+ELcKBdqULW2UNiJsekw0XcBnu3FtZKCP
y8FM1pNqn5QOLoECxf1/HGsPoLWkqCXzvJNYt60fRjpUfdk9ykfjsvBTsOy88UKU
cuaA/Abbmo8NIdbNoeREod2C/ZWUkq/bpnRIMCb04u2EX1oiX5Sdu0K1tFqEMo62
0kno/5kYs0B+Z9mUNM/qNus4RgJ+/NoigIlJ2djpo/lsUurG7SE4SIwE2RLTN7+f
8FkaLS5HuI9Ns2RSb0a53jN3Ngpz2kLe4RypUocl0NF5giUiFE+5dFDrTQuWC+lq
NfH3o8AHQlp2eBfA2kVShgviJWePy+r9d3pLoBA7983UMaE/Pbg5Y/iewho7I5mX
ZhjtZMcaZvIUGZY85FjUJKxJEUzy/GdNRNUUgmC7cJXcJ9FG5mpJhUC7nowb1b/N
cA+CWg2y74nMrb4zt1vadmry3hi8y5kCvGKvDLLqrPF8p7jznBtAWLv27ra4SJXh
d1ls81ObTRT5/vMp+EQjM5kQiqzVMVEFHmIphvQ1cx9EririfxtTZssUU/9i/521
YS2KJccODunYeXtYXyF45WlyRWvpzISy9n0TMNiNvBkQX3CYjSNl+adag/JCjmQo
kqGHAJR4IRCr85TtVEciLGJ6oC+FZn6b7VHYnz2/AD1YGK06DWmFonK/l8mhU6sj
iFgsU5BY0PKCiqq8XXx+pk5LicdiArJ8xMdxkqgQXTHZZERmEEiX9y07Fd8I9Suv
ajzE8Ji61Tshb975gYt1c45jjwVsM1KFKL7D29KcsJuVFAG2+t52ItwgOAQo3usL
HmCYPcNwguISTPs/1Ux3A1BJKVoZx1B+m+00etShb97fuCApol3U5uwWPb0nb0fK
BzNjYYPCV3X+7CKmfOqhvIbbJf0mgPFqytv3lVMOjVIgqvg1cIhVkHQGLdqgp16n
MCPyrdmjJKn7Up6f+l86cPrNbzZRH5hHh9IlRaoQilBSaSBaPUFPBmBqFpcNyK9Z
b8Ora02mz+mIR+RrN3UTfBO8pwKwgx+ZSy5GBto4BbW1sueIRBHJt4JlnEnSLB2J
qhEzxgcyNehzmauaYdBu3ilFDaEh9uNbXdqolwUsVryPWjETFcb7Xs6HVzgL08P4
eGypQ+3yubbsXrynVFiWWuesWBJf6uxr2XEPqda3pvryKTMC7zQjmj1FdqlIm9hY
GTMJRgT9nZXNAleW9TPaSJ7nkh6hERbv8OqzUUJfkASI1w06PSAubScsjtggfwdM
sYcLvS6A9+ZXwLgG/PzmLKzJGTaoaaZ79ObkR1+deuGP7c9QvnNkUGBjQC8E/wgP
BqBJY7tcGSusygJGQn+g6VN8lgknEGd70mvWWPV26mLjk0L1uM2tGYpj0hr5sz8M
orCCvJBiHejBjZfMLbVgFIw6BSrhakGgNTz7zl3/2+yB8lZlQk5XF8RYQ85eShwX
RAPh6bec+j2WgkhJLA/t2vXNpfYx9Jf9ZJ/4dry8ACirO4RUB0P0zMc2w+BUOGHX
/y7c+8vYWgUMMlQPbkpYXLqlibAUCX0iPXKqzbVPL+jE1YWssTtN/T5VDcgC9kVg
FQ6m3Zf/9PP24+xFM8tYt2ahujnO14V/mYOSoJul+0Z5WX83thbtymYuQ+wLm8Z9
5PySHJF7+oYX9qKje1f/5KIDpPolCV+omKXrMlErGFxycqkf1DrkCzWoqMwDIrlO
0o+DGH9DEUTXsgzyHvwU/Bx/p7z7oZOOV5sXGFSzA8qbiOhNB/jtJ0jMA2u1jQxP
mKehH6YcUTUZN4rShOiTQEAHqyxGg3B3nev45hwCYeoP5Y7u9g4Smtaei4WqxQXf
d06vx+63itJZVQgnJxrZ1W0421K2e6bSrYXxBmizkc6Pj3wKfxPATTnbi0Brkm0t
fghKHtAwxmu0tcwhxwMrkfj5m3NjnNyGturH4PupgBEVAwucW8OX3KrT2adprwHE
YucJnIlsJwmx51fa22dTLvaia5vhN4Aqkb6BU53GOKhdKZDpzBHPPo3uqXTXDTk5
UXkwQ9F/2uCONv5GeGuZQ3i0Lm7nChLp+t4qlY4UyQXxHB1d6wISGKTNYLa24qeW
x3Q+5LVG7ndvplrNKDCaRkk+lX78OBxBVBbjMO/FNVt1bEdyNuFO1Aon1k410VKv
vBV7QcqEhsv1Gr4Rf+Wpqf4TnW/T7XKE7SkzyMzEuO4VA+3ZiaPgppDgi5+5r3Z7
XapVQtdJ6jjEpRpmXOjGZcMNv0hWLoSTK3dyR6uAJan9lbWZ4gurIMl1/t1Gm/6d
ZN1cRQZnjKmTgxzUoOWlxOAhY1oxsHZZnTul7xoiAG3TrJEkneiSOTPmhgEK5ewX
p893ZLc6VHG0b+1x5vW5JATlKWT9SVDhZ6qx9YeekANhJKmKfFvjStwhCwRS3jVj
vVARrQyPDTIDm91TfkHGGQZJRVO0aThLRMIGC/TNDE2L3vKXvx4II2CQljtN++0U
RvJMvxoMcTxnNAaTyfpNLqAN+7wFGT8DDv+KHIDIgIq6lIiLg1QP/81ev5BYNcyp
UufgS7ryIh/mhL2F632PajZmhfVtKKhK4v79ywi+gS1uCoHOvKRpOqYgAYV1pequ
ydIQa1Q3PFOQSTthyj3gMkvm9f90JJnQQxyV2X1NIsfxWYQKsfubm61FPpqxZPNk
dXyK0tnWczPdH1eOmwUBcctQNOVbRQah7PUB7pTHsBdTYWyacouYgeQ+mczi5vj6
XcTe+iX+AW3uQ8kQ7jJAGM45oK3cjp86ADwYdNqvgA38+3fu9T0SSRbttr7gtVFb
n9BRp3GrfMOHB7+7+QHIF0Jpsvuia6PKjc9IW1008SznuFeTwF+O5CSB2lg4gl+b
b3mhoWoSyuhUReNUZ0Ixd3jotl9J/6H+rATf/BrObEP7/0TxikWoss43oAu5KX3A
rbkZ+S0PSrq/o3NMx++a6/Op3arViStXd/xpYJAjIqnSi9/qlOJXAfcBRSJInX+V
ECGL7KLN/Xt7tEaquadOivgA6XRjz1eQGUYDLKgh26OnCvrDl1aUos6bsPBE9cqe
MLRXwWzp3DfaWVTcNQy0vBLmiMR8JCjIGVkj1O8Wsx7UfDdq9+GYLCFEsliPVTk/
r4ba7lMQB0We6dC8BUieTQvh4LdD8UUffZE+ltnsuMtg9T47CeuTwEjU3IrvrbhR
mKSsdLsIXNkJZhRIgpFFpx7u8hNROCz0gzgV/u7hp0d31pUeNIb0Qm9cEn9AzFFH
OatNCSGlqK0UIvl2amY+n8vp2BoJrbrgsx8n4tlQ5Cqpqu7t6qyki2vjJFcFuVLj
5GPLM/Kc6r4tKwlu0+OXgp2EQbPLba2uZ+22iC2JpPNlUs7xSYz9PjA6PAlZYcYS
V9tKM1L3+96rsZNKw5faVhVW2QU81vwgMd0EhSHrMzj1Qy48OBmuzfOJ6MR0CB2Q
x7fRbgcRq7+xPbK5WyL7/0Ag6EzADK0DUUCxVr0PsSP5Ki9Y9QT3h8bflcv2RfWs
2XuWGajSzaxDadQs7njFBdII1Wixw8bS9EqmwgaBcYguqn2jy3IzOIWeLYpjF5Ly
UoM+CMxms4fHgqxpDp3VInMgXGmAYepe20oev4x46Jb/izAJzF8OpELKcLjelT0N
QH/esZBbuF9FtYkCmIwnOLGyzNWKld/yzmanrG7cNJQ8k0qbb3d9LbNZhCp2Qt0E
892WK5CWISA5yyLc3QFbWZm4ZnILexBY34B5QMvWmbTKzMyouj5B+ZoGhLUeVuag
ImawVgOKhLulfMwJ8bJBjd+8htXt6ZhrjWUKKnffGDx+w4+AdwPAeyvjJQ0cKNKr
Tam3wzXgBpW7B3D874mEltxpHdWcJ1ylrTgigdOpkLnzi6g3ptt/LUJ0C5bWl0U4
NBMWmjTRzbNKVZiZjugjKGaTDR1R12p84oC72ddMwCN0ZYqP7/A4qartbW5++vKH
AThfp/sUr/r7Yf/8ySdTF8RiZLGZVInD0l/uWD+GuCnUl/jJlze2QaUF5g+3k5Ug
EjyqsaQco1TR34g6OiEelO2K69vc+IinmOPrPUmJWk6YpeKh5jc4pghzEIenTrHY
qF0tiKV/EEczlG5mHmisRa/DUVRy8XEFgvVdg/QLP9JYsIBXezVWX6FQ9lCJ45e8
1GUlYAGUMoFgQKxo0ZZvgrnR3CmL9W8UfUsjJTkVim4F8jHY0GxEl2Krfpl1S6wD
ohPSaaFcQe8AOUk+o1GxXrGWpJB5E2gafFUQo7iYiJK6lKdLjkvOC5KqGsd/mnca
U/mo+2T5yLi6UOQL9N0Lhmug3OvBNp4OOsX0MCZL3bfAPNW47zFQrGNLA9bq7spN
1P9v1pq1IsT6TEyqEU2kcY9g68ew5b1YYMIGm+IsqOfvHVwTmAVv7NprDsvekKFC
b9/D6CMWmKS3MoRXR6zFqc56Ws2Ackn8C26HAk6+/yXkruf+eEh05s+w80ZdNR9o
XEJusRPwnqYlPg9/vCH54cgvT/iD8IjPxZ6X9FzBMpjO2LDnO6QgHAngIVlPOyzq
zmNRkLGfgNHOsiux7vSgCXAZ+OfhRE4RNC8CseYlYAiG8NRkSt/+zPYhyak3a0PH
scAKO87Sn4xgaZGm71N4xbkCE4Zl/Qclm9M4kDnqrMcaIac/0HVED8LUV4+j74hZ
Fe1IRxN4X8dlrJhH5q9t5vuY8G5F8dwCWoWVCdmpsmjIRUCz0m41qx23eglL22Qn
9Lvnylm9X3/ymGiNee+Wz3fxrlWKCKlseJvPMWMUr6ONi+cTswDcagN0V+pRmrun
138WzVlTdxfwaSeEqyTmLEIPxZ5jgTZu0UndNcCs7jREFgvjKeIc79jPfc1PGYs4
v5cdBTk6nc/J3mpzpBLfu5YxD3PjPmuONbJoDXi4vkZzyU0oC+uYJbriuHE2l/7X
VljrBaad/DTgV/vTChOp7Eydp+FlUMrKi5N7f8RJ0hay0bdifcbRLLsQnjwSt5xd
KQ0iMbtAhpAv1jxraS75QyY30zBacdwVEjpmTzxtjhozOoCin1i4q1AdJ2+diDC0
G+vIKJAE0QsC21kaDqQqMA2WHTF952tI7RrwwK1l7vfZCZaZxZvNAv7n8B8wGzEq
GUX2KcSoWasBP+iydyKFqvOXReD1yRm66ezJAZUqLA6YtmZvQck3BLT8MXlIMPYm
CxZySKWA1XTRRNMTbNistPOgvjjR1bX+9QP7VOjS8btt2mX7vYoLij7zQCj/a7aH
8PY7rSEPxeEIPpQ0YG9TRMHtIbcGq6t4COCy4vwXzBO1yK4aU3eseqHAsqaZCFJy
F2wQAJAd7I5bxwSyTTfjcirgMBNSnUtpke9E245G5pWV+mTYLiMpGuP0LtK7DlvV
2vTeUZ7KkcDxfWvD7l3HxjVAlpLU5RTWem2wGj8G7al6M7fa1vMHTdwl6DvAd2Og
Oul2fjl3IBw6UDMFAko4njZfYfBnvMTW/itR3H1ZMd/H4GSAKTFlcUpAfzexYFTy
eFUJIKjN8TXK+j8nTYJNcWxuuzSc0tz4TPETO7xfvnBheni7SLz36UoC46xZn2fb
Y+wsYlLs/B4CdMWUGlYUZiZjt6juaplLs5bs5KPZPn9NGKl7O7ydVSkRgPjImJyE
iwz3FHVgC17UM0au9Nm0KUEu/BkbAcJ+iEKc1eNHsbnnjt2LV5p6GDva1Ng2aht7
QvOrBMWpOyUkxIuhWzBh9XYa+94n99JInlxWdBIk2LeHEmsZ9p1VQmjADL7cV3NV
oglKC66Awc3PXMuWSbY48ODUVmXXE9yppD5ZnliXnime3+KIbwnvFC62dEZ/TS+4
czTJPP3wpNuPXec3L6ALEevXmn/ta9+1dLjeuc5Z/V/VC1H0Ku/MVqWrn2IIt9yZ
56d/OBjT++q3IPMi3r2m+h8yz12SlLdkC2XAf2tdStfXT0kMSx+x9zgFaEYU1BI6
qn19C8gfg4eKJemk56BdpjeJpG1xkPR6oV57gnW2hmBQTs0qsp+osbstQ4YWD8Um
LkxZ9b9ncduoZrRzObVaTybBiCoivxsAMK9PGO+MN6/24w2zvAAAKpsDWTJ87yLA
Y9HHv+ag0FHGbtYyL93KtWfAauE97iiSN9AvEKuAWAawMmPH5s6mlP4ortiA9KM2
8+IlpPzg1qtT+WL2h9O9/Wmt1kuQbQ/Sl2roPGYoF9ybC/zbeqES3DGrh3jNpsKT
ITDSm8EqLKwvxsFFtW4evxBLYnVMKnWpePx3OYve0jBbghEGcNDd6KvQUpm6aSXx
c+5knRlcUFsyVGEBAtdjt4DeDB07fe1KKb4an3lkDi6FhVms+JX6ukyeE2uoz5s4
+d8NKVHVBauxCq9u/5dDcyAFGlbAKD7PB0WfmKeuSGIgXXsAKsR/dbKA4J73HE79
uyJWlGsvZqqi1sOA/xQju54ZIevvkCdwGw825mPHh3/4BK21qVEqpFbvq7idyUdF
fCWjXUW8f+8XkMlYMjj7rOhAmrtHf7uLsxapMAPDhgK8/QxHeIPm46p2JMkkRg2E
oPTXxFiO1CdOzRjAw3cBe2+QXtuJl/96yMy1Nso26F2QcSadHtSD82NeC8vvTu6N
aLMuZiFgPZuH1QIuR1oaSAZBwfArvPIpVylh/c7QzvcIwybG1mTHk2ZXELEzuB+P
WmO95bZ7G8izNnxMCu8s55JUhsZk5HvFtpnPcj4OihPa008LwSZLtl9rBnKlvwKX
8FPj2LEHLNf0cV0t4V4Fo65EJ8yYUP6DbaBhfimqAtHsexpEroTSS+cCgr3gQnHu
5hukGeM6Sl5nSuJRWSrZgh6kz/gOip8DytHebZ1vpPJdyeTBgs5rXXbADLuqpLd3
u/TZ4gqQP1lwLAhyOorIdsigOLIznO2hkQabBdWvm/o77qfRKrwSHusNxr8crnj8
xQkhOpgneZpCfNHBRLCPmjRO8T0puzdueVohB3P3ai7Hl3AumQ/HtSAbdy6+mxYc
crNDaqZHkRxuSPtJCMTWN8RajWHhfVmIhq71NXFPbljFwzDPIkyE7YvtVKGumKiw
DuIY1UD3//Qs9E1WD8hlT8WsyqCHG4m4hGwX/LP68SMxlbvsaXkZ3j0tulrAvLpO
9CcR7CkQyklfE08nYt4c9hBz/plTxYBdgUErZSX7EZ4NRM8+IcrB1ADL9oNgxB7C
iBp9XxQwrBhD6Hnd5kEKU3ebaKSPGoLfJOiwfnuAY4lcG/WxX+GQQ0GCaennta8i
uygu4kD4M7e9nUUmMZZY1el9ldPt/JiYOrbElAskm5UEdRHWJ/qR6YkwHxuDpNpv
E1Orp9eT0FL2wCgb6JMNz5qWH4ZN/CaTRoXGa/e7gIpB/FHDafS4XoqceAqIOfOg
HGjy2h4KGpOJcJRjWEu8ETjvL4eSNUmeS6FkjtTZiheqHk9znQkhfAqRlkzznwob
Q8HXsPPVJxQs2M+FYIsT+gRnrf6vcpIeSpVJovXz4P6/VByrWCFSkcYPKaTjQZf6
giDWASn+EcC/qAESHeYa3GQFGIeDydAn9f0x/758BI5YAG346x88smta+O5O2RJn
cuNspdDYP2n2wDkCMMH9kB1PGij/qevJeXpU648ddLZhwgRCCvz06Eatz9q0gwNV
uiCttzXS5SeefpPOZWPQhCPFHyjaZKQHznC2W2il7uEiWgMAMkPpX1HRc5i1x4Q8
94mMOotPGiHFj2gXG7E0yuHLyDrdiWUoMPRmeqONGxKFElwtinc7z9txV51ZBJAd
xBXNX9DQvHwMPzS6fxwyPZJfJVIlYu9+s0i78rBYKYgHoKvhKUBWxXiAgZDft/NA
73NFRytyEA+nnxh6aJSLyTyszDxYzRhcQSU6o+FpRDlBXADyV96xAz6OxCLgFK3z
FNu0cz/s3VDYb4VsG6lXDQLAcyNGsF/WHqsu3tC3H+cpLkq+Mz5FWMTn860ytkj5
exhF3TSzTqqlROJoItAc9Hpi0JaEkiQuuJXM5ZKWSHPRBOleeNill7cFiD2BKxyh
IZuJW6QNYPePeyueZwfAsc1QHFABA5o/Dfnr+1JjT4D22PWZjllHbiz9aW76/CQ7
wJL6yvURVNNVhu64mE7vQUADBDhtzCgqKZfiSkA3kcw6vm752XmD8M4zbbRQswSO
73b5J4EubbDx04B1GC/yxvTssx3h7KaqMx4P6SnnPd2JeEab8rkV24cjuS9VqhsF
z4bxs/m9hlwMdsnq5jDtnm2y7LyhVZR3esOacCSznOR6Xbk902KZ+dV+3lt1cZrt
73S9oyE8zqrCEsmffoAc2p1VPYfAd2tURIRXsmBWXHWDbVIGmcCMBsp3sIdSRgUe
33A6o12L9dqZEk1WqAbtWUl5WhGjGIblOYmOQTj/9Skm8inX62IN1kUVQllJ6gza
b0ZtwFvU4lb/m16LyFLGe/0zXpbhH7pcziOQTfZ07wCYQ67ySqVL91+R0gICMNn4
IhscXrfbm+LtpLBtZ3EWOZ3Zw/K9pVFVfmdQVJdFMw+cCMI+JVnCUOKZgQ/xcXh8
D5UjBD9LFYbpgcc6Oc/24/NPgd21T2/DbDz3YUgam4V91JaqLReSETeWHCB/OeOM
DHo2f1+HsL0+CbiKWhGve9HJKkdtUbkqlptexqGbbTzmzd1dm3emFm4J0HCtSThs
u9YDPtAoWM4gHbBUkjzg7PEKPl4yn3EgNoYn14NTcl//drIXbkK6TB7cbvsvtOGr
/67y9WPeqnueuBItQ5vg9HdNwJCK3U0vx1e8Qk1M59dUb/+6vKWnpdlvp+zknVWU
XzWQMDsVzv2Yre8vueF12pwQDxjqOE8MRoU2KYKYjrOqiLD4mBIaQbRUHpddQ6ZK
qULMYpCFlm5jqwYA6VNmarPczQIk0cEL06JZ8A24FFPTW2DnmYy3PpRJu15ZEOT0
7UxumacsT24dm4LbaPp3sbCQcEwF60NK8dVk2/egpL5W0NIX4e5AQODRr9md1NOZ
qdJk4XtNq21eVQ41AGVdveJvUujn4khVwlNfj1ziZ+J1sd0OCeRzUImqg6frAcTU
dJKVr1Tabb/TisZ7Um4a6HyXIrSs6VzfN1KdsmQQMNEfg0X/dhJIaFJcsyhyu1o5
cMC1VtBHG3XiPrTi5B1mUbFvRtHNe+MWpaIV6+HChZG+3+e+7nElq7VoSEXOGAEH
uT4VdUdV0bpZq+iC7rQ34hSlGN/C8mSpK7JrnozHXG18TmR9YBmUS7RSZ73scFaP
Uo3CZwvErw4Jo6cH1xhEEfxfBVaoZaRPp8CvKpekVq8CwQ+CKu4T5SRucsjxCi8b
C3AmvwBdzzJf2seJc/Lqw2RFv6zpniL7fQMTaxgCKEYV5+VwAmEIMSKV7lmqGlt4
njJd74pVjsvENmNoyg1CYBk6j8cU6Cn0nQNIPqd2/7qwlYSMKaQVW2vWigBBwHZz
DjJAeQ/WwtYqyOHN4aNi9wNZcKhyU4RDu5Uci2fbU+lg3YNnH1n+6CiNYr24SYEO
Z4yfQZrEMLK+bUgDopK+7MQftXDwLpHKOYBRkr17k81BFoZYB73bF4ja4FL9/RZ9
QJjPr/d359dd/LQUXhrtFNnfFjNwC3lxToCq3/RUUshSl8oeT09R+tVONu31Zx/d
oKmQlWCnzO0bPKv2BsNptZIqYuKCL9jW0psn3rzjOPEEA6Hsm+qAsCz+PSzegoii
ip7WqkRiiqpZYNxJ4VNFYJ5vSimBersqsjrlSVgfHnt2oUa5klBEtEvhy7w3BW1/
aG1RGRzFIF/wB387i7QlKW0nFdZd/Yh7+EeVFeQYM2D+RLKxv1KzA/wxHoXT2fD6
GRYIz605BfD5OnU/SyuGJ2PIhpb9BvWQVz9/nQrosGrAXJxx4JdH4EbJVutZl1lN
zm+lha/3MOensFPtyfBjWZXcttOY8Mrd6bmkZjZr9U2KUKCmA0ysWKxChcVfVy4b
MFlbTKjtFuRj8CJdVu57lW45UJggW9ZitJxTp6MZQdpD3JLPiImE7Sb8qQrXl4vQ
0DzsCvrfYuhZ4rLhYvTInPNa6/CVY37HXDKRqqTf+yfkKeyVzXVxEyW2xVS/6M+e
xnVpy/ArKvM+roldZunPcPGoYEYpdxR+KVRop8RuY8DS4bSKmCwRmmVjOsBn23N+
ygKJblxWGVZ1/m4gax7kICxF37skz8TEV3yVY7F1kSfkiZfD40gX6kplgXIo3sfM
JQhmBEqEC+NgQzZW71pTbEVEO2MTdd9o7kFLwF9atNMTieoHCm4maYEthCYoeZ/3
bQ7D4iH+bLDe/sTdWggXActOoWQbkCM0PCPPx/5Jw++xrJbUKnwpqQuUs/GD+XAl
rGkeBIJ74crbddgKHHeaLxfRJgdx3hvjNQhNEuuEpZj98tLahMGC1AAlsZa2CHef
UoZopPgOI8WVzUyXhU8+cTuukNpf7C5sHSEjldBQPm4kmSelzHCCLB1wRmDy6/qX
tk+wZPvMM4wAjW5/fiCQQVcwgy6fDPn4VQj2N9h6B7+HzqVJpAlt3zVIkL72DwNm
3cC2w1ImOH+e63jPpirWD996wxG6P7P80Emgw64ESNp4EiLKt24Yrpzf4NmpIviB
IXSlBBakU8NUEd7ZO2lHQL/odqPoiKIeOqlKUmTxr8nbsh9/EWDmGb3R8JEw/je1
k366uFGb4wRYE9G2SwqYEwyyf/LO/oBuAH/8yaN8S4tFjG40rE/Z1sBPxK3WJK5v
Ku4hoVsFs+MlXi56oE8fmV605ofvVXyEO8ayXpRPLMFu67z217n66Sr7wWZpWEZX
XF75n2B0ul8+wO0iI1823EWY1rTaJNZw/4yfu9uLT5P2jjZJKFBME20gPToQZ6BC
/ru07zysiZPTU/OJxOBt40HG2s6DG5yNwKY8DZoSgVk4SEKFDuFG1lPchLNdb3Zj
FQyWeE0ON9LIPh+TBraG0X6c9//kU/H0cuO/nYiy5qkCibEv7CyGkxTPEvouecgF
or+ZWReoV3nNtgQ0Aa4XkJWnjuc4VeENctru4+jD7WrH+TOaW96FRgcM9OenUqsb
aIdlSA0JdNpjuyjYZYbZiAgXDip6+0t92HtUDMEGXX4nlYznMLXcH7SdAEQ04quy
yAU0Qbojjy70UiNKz3xyO/pNCoUeB//vG/ZDW7hvqyRBxpPiKBlIs79oYa2wXaAG
xZeiZIOvtuRKwQj4SRim1eMC65a4VQDBz8z6z2BCM4Ap1o7SCjWVJfwHbM70oYNy
Y87tnaiXn0V+PtHRyXqWEDYwU1Kxh8720nuhBaABjSxybfTKje3CcqncLH6BNPHP
tfWWJxj1L7PN6d2BQgkGQKOZoM56sjhDEBFLuT9F3Maz3FjynnnvbsJZoklCuFBs
Oypp/91xjyrakgZZx0WE2BD8PWHyRzlSHpy1vVfXQyRM8w8e6hTg16DkJsXZlcKn
PS99pgi7pdZ9YxTBrGOG39R9O0OK+VbthaVVzgEjOZ8ezuDkFleFnldSZgqnAq4W
LVNvWHl6kHZ8YoJfLrdSdiYL3OdkmBoWqNnSZVk4rugJlf6DYcPWdvP2/6ljDoCk
Wx7XsnQ2n8SyEz9k3Q2myQUbEBEgfuQb9McpfINwejFqyZOEdIPorumJhK0v6OWF
WlK7O24eqys20nXRRyAMYJPedQSqoo0coFV7qAkwJoG1xtEJXgTZiZUYoHiEbudY
+qdU4oGtDsaWz22fF2tbyQFP3CZOi3lsoB3zNWXlrTJn5aQlKlWaqW62TBssZvGD
iH6hnzb95T0RQ3t1kXYa45qoKfM6YljUsu96vPZNYLdkQ7tNWVhYcaYHIRcdQxft
UFquuDSi7xeAevbiiwKLDJwadfLdVElqDEQYZ2YAEDIh/0qXWupyIWVMOmyiGlNd
KPdXFnzON00zRXo7dxWNuES6zsyWvEBRFT4z1Go33ffeGhyFNF0gFTW8FRxjyfEc
O6RkkreoAAJJ+qHuSevAGgEF8XXYKHu6guPCzzBGpL05A3nxe3soyCmyH2JWLG8d
+RNMQwk/8CxotqMseoFePHoQStXsxSuq9/tN2awx/XSSGZbaH7CzEbCyZdXU1/Lm
WXm6YtE0nnk7hCV5MY/kxTb17L7/R7j6YvhRcLm9k+JWtNcf0k5r77JGepmIWjfk
3OMmTxuJr+EW6v535acDntcV3gLe4zHnQQpSJRPjAtNg6PwOjr2eLuSbkPIiDlye
KEVfgAiZjepyeTFKUT2gpnFxaJ4eWXoKUDzsbXlI/kGQ5SwfHwl39OcFDyyfJtO2
IpmxHp3CXfOPR/nT3fb9b/VImkVlrSOyItpC5ea5ivNxass5fJFldSQ4gUXp/uwY
llhhPIuvNQ2vU0a7/bkwovynoeDXBdeROaui3FYiesx+/Mp29mW5ozk/XA5cZgY2
5qmEIK1vicj+TTyRFPPEgSl6ECJtXp8lCpvAGWHDFAvWxA6BtLr/g9WyxKXoXbnY
yXkC2JVZX+hI2SuWBTalsYnpbsQuNiGs9EHbvm1g/nBh/z/aY8OGwn8Y936/tFvg
SE5zZUbL4KS4ecB67nFHWmW5x4IFYEGvNox33q4GiiBFxbBCKEudgOrIiXQ45+FJ
ZnXiPhwIFquJLhJYwW2ctpO7puhDxjxiuFVq8SsJIeAN4+wjwq+FvvN7MQgz9/C5
gyHHynajuWQmMgYORx0utRJ/y3fRRLK+dzIakQoDSNl3yUJmbIMJciG4pTaQPrkf
9DKQiPMd1PMxR1NqrS0s2i8wMm2VXXlE7RplnNJWXmaNBArpQb9v0OcOIm7nPAFA
5JFcP6mJtudbhIGpMw/MGP/6UprV1/ez2yyS2TqJUlILvy8PUOA8pEyr79dE6gxY
nDsQ9Kr4IeDMZ0IRL0eMHKOEYA+7aB4FnBgV4PXBfD6KdR76iwjSXrfDSPILfZo+
Z8c5Vn0joxsRW01+2L4jMxp4TY+GF1v3xoikmSVanLzFAdW3U8G7MBwZWYtnVPiY
W2mcJuM9F0DaaWQfivTf1oDmWOXLSkvUAqyeD4eOcZWSaGOiKpZkSfr4gUcUBnJH
p7096jAkwhD8cB1SN8VKiugzX8WR+a8fz+ZzvepVfeWgSwK4vnC0WEWt6kNaRqkz
zznYWwLI5BZgDrh4R7yAXKlHjEc98fq7ibqkEdqn95/IGrYa003IIQpKLCkAzylx
T5ZJSfLkNchsfcMKFVmirbvDealPwbdAmytmcSBhG1uvsmv4uVlWOttOW/Br41fq
NgYruWeRYOvODkPl0VxDV2UQ/E4eFAA8cluGz7wjCIgBgGKDVpaXxwz9Kw0gBPvH
0sfXiVKI2etk7Ok0Tzy6BHrpSGzQgbmWu7LJ/o2GpBCUX34Jws/0PfBI8Hn17/lt
2Mo133nzvh/z3zagSQ4fO0ZGxsjk/o1TwhtA0dk6RYx0bzIHOH+/z6DM93my0HTk
HAgl0gsJ5ZqJuHT5OziokYlWgZYZHGeTV/TuMSrPzObMqDWCSTvAZL3vqma5nzZk
MnvJnsAtHN/aXsJ8WSAZldI7CleXq+a8nelH4Ew5neVX2edcjjoZJgF46YS42LPy
lqzslgnKX8jM6VS0g4Z+7NY8z/FhAj1SSyDuM9c2XR1yADlTeapf1gFfOr3k56jY
+jfjm2sGXStfX8IcX2Nw1uYhC6dGUy5Jv22r9IIUKCYXpp1oNv7H5Zl52OuM2lHE
Sqwbe9Jbgpc7WYxQKrRFUN3lQvdEqOMuV9fPHwG+F9xFyLc3Ry9DkjaH+FzU7TvQ
CsuAJcMCWSTO9LvOcCw5DfegkAJuvHv8gUWw3uZa4l7DtKY2ScJSf6mZAOw7ORp9
LFgebF6XhOMkOjlHS9lSMofZ83JvcyCrh/gkJXBHAbl/CgLZP+Wa5xo0g7DdBdsB
QevX8EVAnX+j8OiNWVdd7fzOrShkccojG5p2oQspwj8b9YpACbIcy/JkfFjIFPvt
cH1sWEKQqr6vSaionv7neatSo3YdBFnxGSzmh/et6lkRS06Y6C1RGJhRXcfTMDxz
BpMoP8m9l5Y0BCKX5w2TAiztWaScQc5TddGVmGLhYBaJmgbnb8DodRA7BR7odqpW
XbSnlXHMYIVmpaoP4XAuyoDaeTrD3uu5OPcz5hKmY3cqindCkGoaNRmbJxLHd1WY
ZORp1qVUhxYjk/Q7T/Mg2rkbH7IFU+11GdwDK5y4r2bS/TOvlpJJ5ufw9+l3i4Hu
4JxQS+U+2STcCT6WI40hyDjzA6htTDT06F3vehpomDcQXPIqrB2p/hsx/3L30uRO
gok0plpl4IFVA+ThYZGbU/TLVyxEfdCpFQ5RO1SJ7d06CZikGSP3YpUupl2ka0rJ
Uvmjmidw24odTeCOluTsCCMlUB3PBlm3tAo7uUDp2GOHxAi9PtbZMhYEX1a+tWlV
Y5iw7FZiNUKXAx6ijfXvDPMfeQMw5E0q0r6X9x1jCxjTS9pEM1erbpdrYRg5g3/4
X+UUQfDa9do+N2Yo8lfbbnj4WAMjNYslLuV/XSm/8Q+tYY584uiWzZemo5vPPdWf
26Ixzoo7+5K07QlpqRFYEdIxLz3DoJCJ3Xbrgutrwwh3mqiRJo/6azHHrjzYCDfL
Vasl5j5I8qo4i444dzfDwZlxB+yAy/510T4+QHBjL8vUQnbusoMF2Ry7lGsMRvXS
0uWCqm3/uwHADZsKbRebc12d13LbJwmP3gyNapWz/lpAUrvwrkovsMcjjb9ySWJL
0RR2vvKjB91GP5nxeD6MIWA6CMH+kj8WIuOuoMAn47u+Z4H0NYr10AmbzzX2xEmr
bVYJierbDpjjZa2gRm5lI7wqoSyhbwHKXJnX0zQM5fNp077m0O76qiXxkBPRioYg
jA9uoV22o/4ql556S9uo+eWjvlhfOswv9Usllkd2mXh+M4kMIWc+5LTupR9ast/C
tS1khIRaujtsn/z2i0GwvmPh0QBH14i4sMZ6J8EB9Y32SDNLH0sw9/k7IyeE/Y6k
Ktyh3jhPWoL6jB5q1ce3EpTAimuWr+kII5cMzarjFF9vMN9kT4j9aUZbuJCgcrbb
SKhbvWA2EmX+3hWDGlO+eg22SG8KfPHIQHDwEWqGnc2mWxrfzb/AJaLpWGVTnzR5
6yNlIUESC+j3nK8fAvs7E8aiZuPrDP2oCNAYeeBrS+YP1tV2Z1XPuncSZ/WmLhYT
DCHOu/EI26i+S12h4YKcKMTcxbzEG6aAw7XEPaHZ5K1PpA4gXXXMp1rzD8TizrKF
L3QLJwdF/7ChYBAQY1Kl80ByLqJmpa5BI7rHxUnOjCdq+/wJbtKs5qJKIrM/TJZb
MWK9BoFygrQ2NnhHkqcpeaTSPxEqt7Uwyf3a8QX9uENpWfUVDVVxzGkkR1IEonWX
JOEqdNksLh4ZOZxrAw9VJcLvFAvJMQo+C/efnlIu5Lt7b1Th3Z0K7QyrZBCUpqsN
qcR+jTgaGOVgHTHh24gU7M46roeHKj144lw8nEgriZ/4p/GcA29j5NBiewtM43+k
voFUmQgW4wfX4HxBiPhk7UGQwVXhLgTV/E+Et17GHdIsP582eBvxTDqivp++3dxJ
DTaHmSyu4PM69zL842k5LiV1ZQQcjZndU5cDTHLC/v1L1hVNxmRWAr/PzqxXkkqN
FtYeYMVuUuPUWHpnfWdIc8mMp1BBJF4V7txJXdC1RN4XkD68295kC6icPzvBTHzR
DfUwHWV4FjbaX1MXIXtITXPRIlV/MIOZQp7esN2XRjmm9bHiWotMxNMvNFq6LqHR
68kJaOBFe/43A0VtXGqPC2TlOT8xBPxBQTHViApLiWi+76qIhBDKvzdmVH7S0Wx/
d3kHYe1Ysp0tMWAKiu+ra7kDwfRRkj3ETK5rOzzp0L0a9UsmbfDJIV/kTVEbk6g+
4GZW5yoKXGbe8V5KkYwj0bm5jC0+rTxoyWBtSTvoUagmsAIe0i92kZlcdsOEWj/l
mhOI4VymLHxP9Vj8jtHgGE+OveU1EDvwoWIvg9gYgfaBPR0eedSpjLuu9NK9Zwm5
h+2fTFGKk+Argl+CD4qAeDDsNj9pYN5QL3Cj4oFJrXy/HTkT4w2ZrfPX/62P0q5A
kJWVor6wiVzt30n2h5OhzpC2JrCqn62aUUwlIE36ET4PzNE8LC0F/McjtkwYMM8t
G7Y/r7MZn+hv30MnqAV3nMpouUH/PNtPvPYS37b7O44l04csafz+8ThOeErxMWr7
77fkZd7GHild9UmJW0qEuR/coTfYJXz0zWA713+4ttjgkFExfv7sZodyY4UTZbBh
E7ORacnN2ML1cnoChzZlQLSamLhMncfmhdP22wCY6HJ3h+ZaXZmZog7ZkPLvQISA
DKMOWwl8pkI/8daHIE3MDFLjKb48Akgr5zGzQhLtQYp0TQ/7Oxh/9tTVySV5SGOl
PHyAy1N7BgWUl67Xo7hCxjLDTrWZpJZycU2waBKZXNyv7Nw3F0NpKmPWbXgQ4UOg
LpUGOSXAMx+u4KOG76L1vDqiOJJP8fcxrQ4Y/DEzb/pZULmMWMdKJRr8nqlbv4Wr
PV2mMEHrzFFPQV1geCwm7cqlnUYOxSQGzarqyoyLilB3W08yAIUCE/5DGdF+JGgH
0x4RMnZtEumh9dQI1sioTiqt02pcxY9QnW31k8FgHGWGELvMcpfZ/9Ecqw0LqKjn
S/29NX5AHZR12un1AWaoDrxwLofg3sZ6q9O3gAhf/Vu4xZ0SJlUqSRnafgDIgWrx
VWhspuAmoBI9jXNG5c9G6zQ64q9k9WzzOqey0xwEJXvMD8+Fl1SNTr8qZ2d4+UfQ
bWZ2KlLbUhSa5b5b/j1wCejIiCcN/DL1Djbv9U8qtRTBXgF+kuk6dRBCf1hiMcJH
x4RrUfcaRmngUL/h5czFMR5ID/Y6wMqQ9JtwRvf92l4rJ9Xyo9Ye+l7Ci8RtmyL2
wBmjLycZ8p/Em4eQ/8PG6aBbfPcRcicnRtm8fLrQ7x51DMrCswBvyRR2ItWA+DyU
DFSMN7c4SClMzxMYnU4+ScAGRzae8FpLKzRHWjl5cEJ9y2YZjPZ4KONKJvhRMnXa
p+hzj34KA4WfIR0w5RTBsUbc4vnzdi3dgzo+UsrDCa4yf6Hk2cwOhRSx1HsUngxz
Sctjra2VC2T7u+fQW0gPKC40apUkFknh8RU2WIUQIqn/+MK+7NJoIBaNl/Mx+WkQ
IqcqwahX8ovt/a8r85Cf41iXJzusCwOLczbDNqsyqs1gPZONQjJE/WL3eHZy/4jN
zy7V74336aBvjGCvmdeFNXuHSUnK98c6VnlNM5r9WhSnI8MQXUmxVSepRQmN+S94
djefUe5AlmiM3e8DDPnISQ87LjsHyfBtX3KbNgn9w6YT0sspxR40+LCjTGxWONN9
MD12FSB/MVgy5WtjPae9oQ1PLqcc1MNQ30o5DxUPrmNYqXWTAi0eaNGIqPvkXSAt
61gi5xvsWgqA+s9+nSsYDFw+qavnpAwUuD4c2yjx2nJdPWUK9FoDJc5uIdN9zY6d
/vYOgYcEClXmQRqR9LrgbZfX7VOG53IOjaA17gJw/k8ZM7O1gxVkJ57j4UsvA/I+
apY1FN5fRTNdjum9SxnnWUys4HEU5AOs3lmyK6cmQmfen3GXrJ5iMncmjUqTbi1D
sh2CAMhZbF4WY0SewRPApcrOYHjx4OToxpbM4xOD0dyIhB08Bd4ogV0qrE9SWK2F
Publ38qJ9Kv4P0nlu7RTBATIMpD/6Jrv7Zx0k4ZFmMBBpYN1OjV+V+JOWHFyVETy
DzPKhO95SxKtmGjxrgxW1g3s38Nqi8DwaFErHX6gsXb6k8/Oh8/OES9oKmM31bHB
oZbkIR4di0lqQCBnXtV8Gc5+yzKT+vddcRnBpWKBrlwVV3o1BLlojscjC4/h9jiv
c7WJEwpZnxB9aQPaqcdNoGXcbAbts9BTEvEAnOHCYHiObKSB5PGMEAeJVp5NyWya
yq4pktQ8to4yxUshVLDrD8MOejJwymb/FZe8Kqxn6mWmDTa6qz/mjmJ1i0t9UhzU
rwgGd3pJB4w5FthuizT0tXVrPxq4w/uu0pwAxJ42eMaueB4eTyVXBI8KZSyLpyM5
zpQIR8x65uYb+9wVy1gd/XjaC2tYVDsBeFAhGiQcXdS5HcoVL2erUgKTgeXW6S5v
4e+5viIzAXwrsPIkXoH2wIRKPQ6oEBsPXaulIgOe3kXZgeusEe5YGbkblQSyjOFu
yn5Yh+jSiqOpEkbJySKZeIH7tUZV1PTsxwmgNiO/OkEG+QrdTG1gRXKCiwyVLahf
/52oIUxFUWiNvNwVS16JaX1+N/9v54Z/vsoTsQ55JG95ltgUKpmumQxw5z+6GedU
zIXgxh5Nlr2/yQkAJsD6v2jotAIpM7mmTU/7Ih3v9fj81zX9QGpeOnOefQHFhuPy
d+GxgEayJ/2LswVoIC3TbT0ldFD5/Hey0vDZ98pqO4CmNM/Z6kWkJXpl7K9qgEQn
e5AOhGpKhDG41SZ0K3VXxEavYmojfOeKlo+af6uLzA1pY3CSgztxCu05syCukxN4
eMP7YFYpsRAWCLJzPtqoOiEv1SOq1oySxIw1Y/CNsqHnJ+l2uKR4i99IEBa0Ej1A
HKjH75VYgOXYLmL8ZYuSX70YGjZunwdYh7g22V3CK3q271MHg9/3MiZ7QkWkqeCu
ejeC1w9Au7VEXpxxPWdfZY/J/yY6I3jUD8+zNUgVKzNGNXEYL6/G4NRptoM2LRPX
WOhKuh2YxxeOOtRvIR3AClJrCNPcn2tSAlgW5mlE6J9X5SiFeQEAjFnySKmxXnys
ZCwuKbWBvMGw85hLd4NCvuYr04qjhNIOesl/YnGv9XNVw8sfIMjsWhkam3qtiqXE
aJQsMh8xWkv1WeJq93ls25AfLr7aGjhO4EUHfgUH8QFZPP6TJH7x3M30ohRXzO+q
UDRK0cboDHHQj4Uv79B5MvY3TWLrCmU8pcMi0yhFdFCesOAl2YOWpxt0lLaYy0Uc
SMZMpxhCOlpSypzvFMWCRw/IV8Wqp8ScUtjbQehD2RQ0FMJcb29Esqqyg6amPi1U
2OlpQLYUobyCjZCLI/yDgvJ5V59At3hsp1MYeG0PIqZT2aogNnk7KJUwxkIeWuQe
X5nihz6SaBW+h+D5Jlg46hUqCdG7NY/wVQJdqYnT8r+z45PH0BVmexT1A9clvA/e
YX7p8mJYXh0OJLqVuTwXQIiOQGryxNTNtAGhxhXc4iQ2OD3cnwnqtMhti8eEl5Tc
snjZptSaQBf5xIRHCbT1v+Nnku1sm9wJxiYRDaS3TQ+PEjTqedcMGcStcyBOPcHF
krV6+58S0419k/55NvD5HDg6N028wjkgiY1DB0o1vj2UJ43oObBxdHqBsk+FkOC+
mIbd6YWjL2H2DaX/B+FS7TdRYwBf+OAmyMzzG2EdpvpE+MisbwBi88MK4rNiaisM
Hnq14GozkFRgbXqkS9YZTBDaOVBCj7fJIVddcAn6xRTW2BWPzRJPnMkKyFxmuP4f
Xp5ZrFAUSl5Wc64m6ZyovP8HhkNuB1hTjzcVL7QIMFsnskUn/ZhM0+d8xhocp0WT
3BQ+OJjxel+JO1tvYxCRdNKjyig7bd7IeP3m1Ay1rVoLkdv+CEqCUSW5WVQJSdRr
RDvNMrGob2plhl0HtppvJUJY0wSPTNAMbexPYVJMdI8xZ8NMGGePgKRVPa2K5Sad
iBluJ5WBSqizDWNXlDkTcGyBx6FX/wNivLfdWRVVxtcsH4TN3FxlMlMAALIamMlA
Eua3vdqYQu6yyUHQ4GP5hovdkMZtG2kT3FLRWWQyUnrLbt6kem6VGKu18IAl47Y9
MswQHaC6D0Oxafse9ZJUckJ7JMDeeP8cm86g9o8usxUlhdoqFgtSp4KNPumuATMZ
h+IAxBNKpTv2p+DavOlNpD8TR8dqfLl9uxrtaaulwMrXwXeM4l0bi2IBY1B0ndAv
yz1d9gU3o1Qqoi4gH8xXhkuqa1EtYua2xOsqfyN1r7GBXHqJU7Yk3vjGS7uW+mfh
3fFOXef71szpFCRxnqmRFvMfYvzSbmAM4YqZOV1WNnZWYB7yqYGvsKiaAeb3O8bn
gVNkHGIoDUapAMBKPKzukU90t9wur4AqJ8u+INpzw5JbZsjt8COIhgX6Sa/MACif
qyjTj2dPOmj4Iqs2uDpQEfztvFAv1HSex/7i6eQbfvks6F3gEy7BqvI2O/7vuz4q
TclntttxqE5WpjJMPabfp0J+olFnbs9bPpwh8yTXF5R69iYIzU2TnJuG2I8uPyth
lCxaHcnc+tyMc7l7YElQHhBzAF1h6l8aInd+XvBBHkQAsthr57HV7jOqx1/akdbL
qYthLbkeEQc+YuXEbl7cz9JNFjqIreEjD9YtAuedHwY9w6AN7ZurzA/2ojqhaFV+
2QLtov85Di0cT9TOgZd9q30aEeQglnEOam8lwv4MpNUmEVfg87EaPT8RsMsTmTZd
euL5IDgkbn1acfUjI5LyB9q6+kEnxwxLW1QpJdy2cQ1oTGyXzOzyGjQiqRF9Bqvz
X2DasxahhpPbAkI/GAYkJtSeJUMCrnOnxxquOn2Lti+wS7RltTtSquuiy0v2Ew0W
Vx7JaSqMN/XWL1Xh6/iI5aR7vSx/p50X0OifxQHzZeEhsPbRlmeofYkTZ3JVceo3
DdjSgzOkONE9DQwVoMpw+h6IdSDeyMTFcjob52/C4vXqEM7Lv5Iwijh0a4hujI+p
3DjAN2/hecycVxd6dSg+/Mwus507A5L75zgyi6hNX0vOBUzS7v0rJj7zoEBvblpu
DF9gEqGLcljlJacVobU67OQ8ldH7Jz3lNI5oyi7/9EsqUdhdfbOXxSmyEJ8SFuw1
1QUexcBDgvL2P8ZsKkwFAn4pdL0EzPCOU/AtOmtIp4aTXOa8L8ApWN6pijXQsUjg
3hIUPw4Ki5zmZWf7pwuEv3vpDnGXsXxqmnHKly4aV56WYMQzELhs6/zLo5ktosrf
fxel5Lsbo45F73KpFuRJ9REtMdublTDJzqOTaPI6UyNvJ6ZN5BbniFekoFOwfh1a
eRiPpMaK/U6Y7msmWenIHYCGeknwv4B9YzsitUdSgoH18JXww80J0ma5R0DpFg13
CGYIM7mJFpMa82MtT98BY12JS5fIwvZ1YWVOigpYrPQ7EYPWQzc0h/y1rJc6ZlB8
oUx1l40K77oL3olT6bY+2p42V6l7WAko0vuNv0NbyIy2I96x8RYEUhTq+5803zHN
1hoS6RYedAJX4Uon5vgmp+smG5oljGWnuIZhvlRj3dj9ZIij1jPaHSGV32Mp0Pq2
Mc34brWRDJC7oCuLXH/gfVV3UyywVP+aJVsfWwJTVKnj5PZNKjTWPLRmHL+A2cKB
43YPyrSIdT4QHZlvF2YbgTas24wGqxjn8bVjBou6v7bzCByWSyhbBYXK81WcquR1
7Y7/6TEixyUaxxe4oRB4ygVkZxeQJK7VuKliQi/kmAPqnEoDi+tPoVJ1xHYqeiDE
NnqCjQadv1Zb73jSGgdUVRhX1NylwCWVACCcH7wLZOvcpuQYST2AHsuB6Of7GNpo
Vm76A+to6qKcUw+VMjkCfwjJ39pOedD0bJ/AowQwyfKt+H9hEUiBbyhlKJ3Ycbd4
PAzqM9+UcmhxPJ646oLT72dKLnZlHGYC0Oip6eEtKoqGEMyK4WyHEe/8DSb7W6ht
IY+qFG+gNwdmeG4Cl3m/r9BFNTqvotfVDrpGCDH+kA6X2E5qoe4O4tYL3dLnaGtF
i862PQFETeE53Azl6JaRHZH2PcL/h3ODZHOuu2A46efS6B7MX4rdvsziWyxizPj5
xuwZQwVrze5Y1ORWyUUIAgCwfaacD49hYCXZUxyx18TlRwVLo2AhNKx+IxPmWJjc
+8J0tMnTEUWJPE23ieJoJeJxyewvGynLX1JLJr6IhWqC4mfPGbfhmrxScEX5wL0g
bzWhbYzcYpLKw82SGGzGSe5GA84ZA86yYRneMAEt4MKFbJuiTx00qPkp42jyJtjS
TWjvbQ6sLbjBS8vsFrnvAvkHlDRr3E/kRuQxA8P8UOPa41kWGHYAn0APuQB6Ktdj
ZJ1s/C8mMWTNWPpAgwhILoQcOkk8O5fwm1eYfWsXn4+c4s7eEXY5of0XVczDHkQV
Nq40YIdAsh76C9dmAGhS/bsPt1ZY8IN/+wyzJLXxSWb4D1mpk98d3PbfGknEygGS
sl6xoIVmLbbxaBwaw1jYFe+fi9J6B/xUWBiHAk3ph267HemQua3dK4a3Htm4el0/
hqyvgRVKlFrjMvzMYXluT6JB6F/vqaoy6/YZiinIQzQdE03C9WPfekq2mSo6b6Ke
sEB5zjyGRpoxUq/myMuNu/hzhrtoD416r2vDAHKcNeZqnNj9V5ejLg5mAa/odSX5
IJBHrfNPDvsaRdesPC/LNKm0fMXXTzmxQ7jc+PDPaLPYviA0arrATJ+TDbecNOUb
uvmPNelGO425HhqOedXcbewF6ySeZLB97tLDMC6PXnTgfoK9OX/O5ogfLlzyI8d7
eSVP4i+Qsiv2eBuql0CgOwhpun2yc9Thp8wexvXnE7bOyY5K1RK2tkrZvej51Yh6
xI6xjPD9v9rgBGA/CZL+n3Bop1hh84t/Mua9DurU66g0befRwC8Q6DNFEsyNlSuD
xmK+CklhaIf831Wl/8wrB8Ekv0OLYEJY9B6ib8ntdmC641sP9RZOM2KURLPbzerW
teZBtmHUzylhcMo+j+9LaZRa1MPlOOv47r3dLvaivoG1RlmFxuxVRCegATl7yYmO
wLJt5vbhgw9vkeXdEGLsnn9483gMdhM+5MODqtuovkOTsoea9SuD/HzgivF9jGzA
f/OV0QrU83Qyv3a/yhzu2Pi5wxTOQOQCAc4t9kHLPGstxLLDTohPThsiSajB2xB4
FMdnk0ldP6iZWC5fBPQgFbuc0MC9q2AOeu5BEqE5VlQZZDCIsEbLq6CpaQD0UGSJ
wMa5gbK+Jsj4CyJ0yXa7bkk1Sdb8VoXUYyTufrjr/G38nVRq9QErmlAmLwbEJebW
gE9BuF+7ODB6/YVDFrwawNcbTdi1SQHQXOarXOXh5ZyNuTC09fU8FpXPbmlwbwcp
VuQTGeG2Ff274UwkpFMlQLFpoaAND4CG+5YZwohhJnW258JJ53wARNIQzkhP4s/U
79PLFZ7eUkOpLv+C9udgpBzvhEUtqIovpI/E/w3EGSmWyKPkU00yddXWjtMdSCbC
AvDo50yvK6j9Lo21K3h9IaXqFz5NehII8Fho81OEWPNSE1pUTRMO8ts3hh+7Ds+J
3Kb5K3I4FrA3nWUoId2xUSn9otXEH/qCGGzQrwcki6VmmZqZ0DRFn8Oi9vqDBgRZ
alu3tpVfhpAE6kLwDS/iaMoyfQ+Uk0Mbcn5rAcNzBhyc3i9AFnOSBEcfS+6PscKN
Bj5hD9AYxBkSlufXaV6gXhsClK9BGcAVfmFHv3nA7Hl//QEOO4uK8gyyXslJz3LC
w2j7uVsVZ2AdphwpMzAvLPxcyrxKWWWDNuTKtoTj7wtvZOSuhHnz/oZt/i7Lst4X
fceWxDdfR602vDdP79P1tekq1Jfsc8unZ0OZEGhJdNpIQgPzQDRsCJJQ+2QvK4BW
LBDKgxtU/tSNbfvfz8V7aM/PR5uvnBigiSCse5j/agpnRAiXiwX8WYeYNGafe+qE
wxPD7JtAi55XeK5fnju4vW+UnJCb8eJ3s48ofSYqZA9kf/ZwfPUyxQwpEw99AujP
SCHBks8aBaDJrun98LGuEkGnro5wWoEcFs/XC/kjIRW3wn2yIThFoOe8ebS5S0Ry
UvHduA2P4BwLoWZSiJT/iINw8z0MnUEFx8GvxKt5dbym5xXLlphZplsOLoRl7kBx
UOtR8gXLXv1FawDw4hHWKHxnP0bybtO3tDGlxV9rXIuB7yBv2oLitqTE/g9+fAOL
qQS7fTN4pZEM/bH0IX4AZU463MFcq79/dx3LRkmkj24XX8c/WWPdY0KiHIM3YEdA
3MJlOnPVwEFIpp00yklLxt2maAg26Tm+rHHQxmcvxfjVzHLBk4G1zu0C0f/96JfV
WFViTqK/l2vHi0wIN2gzytKaD+PjWFKUoar2lE/NRmJoOTysCWyaWwNYwJIOEN2d
pXKfxkZxefTondsDzyp8zS7bcVF4KvZKbIKisgWC6QhtLYNxc/hdZ97tqwrmCQ6Q
pNzH6FlVvh4rOmNI55wAci+BRkVjaRWIe5Bo6MizddeGQ9/EWG+yfr6Itzdr93kx
5QfhX/1O4sB9lwua1jB3vCezZGew3skPTD+I0uQf1AWQkuLbpG2AUEJXya2ame9u
VyeAnWZy9eggod59XHbszaw+2dkNpSdyj+hicCnk6gWMls4YloXpSZwGrsJNSwgq
mz9jFiGLCdE1mEvqnjXyvUELW7t4bvkhVHaj6X+nPeSgFugOSfVjM/ose3qcmX2P
v29p4D0afanike0J+HMmCIEXJ99vgcNevcPwuKTF7EvPgsM+QMUkdJZGmYo0XAx7
NBJBg/9bzZdKD2ZTkW8T0ZJI9DYuGfLHg2IAPxJR3YGsQS+ZtFupPMtUkklLiun9
NSgcc2Ss6D0+ATZJI6v7bCB+wn6eBvgCYhbDGXJMlRaErMIq5hj+wHn6mKfjCKSS
8PFpIeX1SdotNvSXUjF1zFZMcJSuCD0gXk6ie1+K8AtWM3IlXoDi0M6W/UKY7tiG
J1rQzkg4Z4nyjrEhDDv4aa7VY8Slb/WqiRTQkguaYuIuZBm4078Jr/LRdlz8NmYH
P5xkfGD0Ne3FC5/XQ31m0kcjMh6s862mp2mIeVI/e5VMNMCq9i+lubGoEjQOsbLe
2zzWPRNP7uDTm5nhL6MMlJXyrFnHvqrjAS47NbDzt2tirRnB0Y6wnmfuPOiEA6/w
X9dPY+S9A9Fl1wyLUhDyRNZDVdcz3QJMyYrbYU4RPjqcRT3lNkg8xRnJ7nzcJA6L
G5La0chDOQOuomvUfqAMoWpCHHGa0UAHOVVPLqRYR9+8nNGycBeRLW9luY4cnzhl
+MU4w+6+G0jlx3O4Ieq8vqSo0N0DoLntOXnIt81GdlF0sbcW6UhlVEE0PMFm48l6
QCszmLfIpWwzgn07fPa5QozzoWaKgBT+DnWXmkYsaA/qGAu2EQjlRXwufk0iSejS
PPmrfsxRo6XKkdCIZyHXyU5NasynsJRnAlOA9obKMHoP2wzWIRkvn1tNx7NsHPP/
vKLCb8o8aLmXLczJwhNYUuWLhswFq41h2/6qQzNDuooeEGI9SU9TT3rh/8OXbnMv
sqTN7nvtvZX0isJceiN/GJcOVrVGvkj8rAWBmGdquuH206d3zWs5AA+xl7WAjPlD
aSfmb6IgWW990wUf4GqNHWuxlgTN9y+PL/ML5yDhdu4nMWmydWOvOD7HGjxOKvNF
YH3nZS0XqfPAysM23fXZFHpNV10vIn7ofnVzw4u+dZ9dw33KG1wqWHFnDYG7xUia
FxOBwo2Ap0Gb1tMaoU7csz9O5gMPo9bn84Q225xObSz77tmnmRw6iz7oH1MupNrD
Ve6JdZOgxvY6Z4MYZ+5sgE8D39J11utjfYCElMfe4DhVBa37Qg9CNNSUPIRsYNhg
AEdn9ivOf6uudCFeddsRElQUDHttxaKSrVaio1CHsagKIA2arIRSzMCO8OM9eG5l
93ZJJbbaTgnlRJwxzc51/zlOy13Rfju5clCinxmMdpezez2FkbC8EgY41V34Kh1l
iZlsjliSP0rIi9k1tp9wGRR15nSBBXmkjDhFT2n45KrqVa+b4FNiGY+H0tT69fmr
LG73y9Q/k4D1gUsTYBvvTh/YKePKAIt5IVz2MnYBgSpn8XZPdi/C8+UQlpEt9nb5
u+FSpYYAaSJQzGO44yWM6beQ4nyyxySw+X6FnVT2Oz0JaOnBdNFLHfH8zZDsXp9S
jPEISDCIXwhkuPNeKoJugft968dnpE4zwp/lg3Y3cdQReWGG2TmXG2bvHP4SMZ8T
J9EiwS9qFk43tME9DJg2qCl6KvNMYsmyfokwgSuorJzAePOFTgziJohryxGBf901
StPabhC3+xSicG2oL34c/XBQetjtZwZyPz8+hrNsxZ6LJl4u6dWKJlHS2SJobWgr
hWbqnVRsQqBr1x/32cHBtynReSSIhgiSmbFWRlBskl60/vYUW8V9wRzcbMHClVeR
g74KjYOoEzuHrkh2a63Rg40vt8lmCwpFi0/F9uHitibBXIDCAWFIqO/tNhk1a0IO
h+EH9yHmw1zBvglEk6swdNds/6sGQVuAMXNb9orHtDEfSa/35otuphNiuYrFXogI
lvXp+7xe2sZzJq/Zx2OX/tCN7C3oKCg2pKsjTGGJ28R8S7s3/V5wOW5TWY5Kjn8q
eY0elcC+0eU9oyVoCQLghlX1lrsIvlwyxZYRhNoCLKhtRnuiMMkZEUjCWTuzTNbV
LHUXtGTMWwOid9viAW6A7MxngupawcoHxLkTuu0b13P3+flrNAQ/7r67XF174G5/
uH7QXOyP0OjDzRuJjFEwy10FQrWCltEWcQE9eIyCLU2Xoy4BMMtYvfH21xxw056v
0+MajqG7e3tFt1PR1j74IxiM1du5X+ixXB7rvDt3tuGS3wV8SNbLFFoZJehrxLNQ
5ybUMOJ0WZK7uFnx+8U80mQdpnHseskQSVNaWbEIneQxX7+absSH4n7URVeFtXng
+aVFZwX4vIr86GloNAZf7qV9MaOj8RZEGM9eXwmkltIUKApWh/Y5eW+qLvrpV1Xc
AWYiH79by7RZFZtwLl1M8ve2Ms1wpzN76EhfJAbVcAuES739YGHC5LmTjd/HGZg+
CuvvZ6jjrlNnP9Lx/JJsz/xdViZW3/WqEXI+S2crD+b2KXJhykgevSjICPnlS0WK
8mwor0pXadqlFgInjdB+WelhX36F6ubni52xnr1jLUQJRAw1UIt5mu27NLiOAfik
nkXk3vAUQr2s2hlkXuDhLgwQhQuM/hLXD9rja+AL2priSbq6zPsdbfnvOmbV/Z7V
7zQV0pmq5eQ21cM2T92EIZfvQajB7DrB0uDjgWPnjiPFYJuMHM1NV1xuc37q1d2O
dF3aLniOS3w4clbPlahWaWevPnbx92Aw/UV7YblVL0l0S6ZMddQ3AEHp0H93VtA/
tZMNGKylxXcJXTj6tKLis1W7l2QbwI73RwwlxchJWuRgW0qtOkD3iHdunBr6m1Oh
yNe4WBLg4DDl3/MFcRRf6hljgd2Rck/aU/I/KkclRFB5thmHDTn6LYkswqyuLp+y
LvamE0SabzTCNg1hJ4phlmWZCcaK468AOWvubC9oVQdPrLVkuNUoOCk3ETbUoFl1
myJiafaCTt3HSbK3YSq4i4E1joel6XSndxltMV7mCWozxWnfyxqfD9jUF8ZYXUtF
y0Y7/YEo0u3X9Y6jNkd8Yno/UycLJ0vbRPMyARV/mInwlTDd9htfXV5KNqHPk4Gj
KoEoKdOUx3V5K2MW+Qxiph+WJy/AeShR5gykVGHTFTV7EHCRDPCNA6bfL7xe0M3W
hMLb93bHdAF4z0Dv6M1kxZa6Jy6yTADKCLvWL65MeAFCQ23C/3V2TmifaVWb9je6
kE9urVXrkG+H/qq2zwbtekFHxNObXZPRdZhAiqySbLMYv2papkxG00birXOfjF9+
uq9wqk2ktYm6GiHWi4HZcF6f/F7nMGEGGr4nvBqHeave87QfUoEksByJQAotPkId
UrbJtJWxiqUVydmsAj8WqIhvUFolOAdno9lNhhCDwrOLoX3D1+tKjgLdK0AIngUO
BC05Mz6Aa359uNWFvDgGbPP6WMMo12ZtfeoV+Vc8dsUbeF6FBdy8ie9BedvemDYf
WPBIgSPZzaTVEnN/akDLGplVNhX9f/W8tgn5IQ7ohc4Zm/SBYRVh8fKSdudBqpPy
tuhSq/hNEbso+9qNW06KDOIagw+2D2UnCzPNRajIrWcUKtXMDIF9JqhcCnAv2eWR
KadjIXM977/lRq6IfTuRbkHYwfGYOk4cSxXYMhqCHPwi0O23hPBGwc7lUZzRHgBN
XEZ0mMVSCeUHmCpqaaL1SOzGd6mv2NoAtlxzFP4nT15BBxxSCGpBZNsPG1DVnTA5
XsBI0wHhgi3hg6wR+s9SXq6Y7jWzTzxGg7FzJPdwD1e7aFuQxrQHTTr4Ho1H+iGm
bVo1tdInuN9kT1JiFKf2PNY/ewkZjoXeqjzEADFbwbdncTxxD6TUCNz0MSPnYV/+
+NhVrF1Q66qV6MQ6Va0iAEEpi9ma7ARAynPdGCK2e0ATMtTUz4d0Fe7ddI428b+O
qAD/XSrPbQAQUHjGdvbZyo0WHPa1w50fliUOFHzHjHSS3s9juVar80hS1HZOyKJy
hzXeUqvV60qdTcIPws5LgLMndUvJn9ur/zQDIoGpGzc5YOeIzSGvACOi4/cVSKZh
rfv8nQn9SshlnyL1ix3/+KXqTxmuTLNYDQU76RH7e4VYWvhyRc6mbGTVvGysE6dO
o5J9Aj6ZL/CqP2igh3/OAp9RbKyj6MQX6+YicWdYJQuHhc03GYXduDgc+l3QFCCQ
yhYNecMn5Tb3LpYZSOChZm7XGpGWck0Ln8OX9L/WoCdFuoE1mI5kAO43VQA2BVBt
BG/l06FlQ/ZP9ueSKaoSQYSoEULIOdU5N24h9WLVdqzbqph0gfz/axE6NMb2sh74
RaPn1UginpMz/MGiz2ePVUd9Ho76QdBUT6mC0NLpKq/F6y77JBAWO+06WqSbfN7a
XoRLST9hIjhhDI3CQSjJlXDIndF7O7FckUNsrKh7kBFenlgAVvUR91R9Bu7XH/Wc
0AlSBnZcL1LDT7ddefOpOIf3z+j80sTEg1OWAdnYXKQnGMwDgnWPvJIN4EWnbxlV
KmD4P1AI1l+awncZOKDzTsKy46ZT7hH76EZ3W6q9fU0Zt75Bfr947H1XIc8nGSvr
J8tMtUmS2yH5tzQF3BaQWMQNlC18ae68PPrV0/XCCngFO5F7HvlvjqJOfp8DaTay
RF7gXpVFGLWDSQIC+yi1AABg+gSDVqQaJCAPBsNRXuD4B27gM1o+InfDhQwBvCzu
YC/YlcXgxzwP9Rlm8KXttPEfLNCnnpwA1pKSc8pL8mi4AmBXONvhmLPXaQgfk18r
hPzLSz3U+4pcGRst9BBt//1yS7RIBC7hsO9oh1axEoU25kTQ0zmB+Qjn/IoZSuGh
csHLlkVs7ecm0gq5VKiuMmtsScxoeHyAnJiZuy1bJny17jqmj+XoUsrpg7aTUr8r
PhYlZ76gS8qMGRI8sRY/562jW/0x/Y1Ens3utqlt5UbyWhmq9vEpD406ggoiXs+Z
6scwHxi+6IB8IISN2dDf+Y6VLDiM49GO+sw7KaiyqJkbxN1eXNmVWycSXJYl/3Tl
0FnszStv5bMCHOuo4p6EfihKOOaZ4dXdhSwFEFbx9dXV1PGxAcwQuUUEBhD4rtvi
iR9rGC4AZj2z6Alpt8v3SPGPRAPMqSTmRH4epdUip8HlpAqJplHHE4ayzIVU5J+y
uxNlTeU/eQwwecfZBHk8AuKeA5Cq8EqIxj/c/qkFAJKS7jsUYhWsTPbPDk2OnxPD
TKKNBe5es1AnTmziNEKt3nuunrwCGe5iW9n6pfAjMKz9NdHSvf47PFuYHdWmm8QD
MUURW8oeoCjBivVmmsUIAlHQxFgwzb+jXT4Zwk0DZvQgVPoOrjQCx07rdRfzfbFs
cN/exMzKOoFTlWgzIQaPdKVheyW8nUlCyhmEHmTaAxKHzg6ZYJsXTittu8rWRoOA
jS+eRK6O6HjACAlSR42EQDmQMdx2dDmYZNaINxnmbhGtSGSgRVUwVi9Yvecrj2Hf
aJzieO3P+r9THVifa128fFi9b1NeEM3pK8fkWkHWnn7d/H/JFlpn7o+1BD/321ga
IGQItnP7Niz4m3XYD/uni6XLROsjBkRuNJocAAstnSxKQZBcQtkDj2b/xAf47CcI
n7frsob3NrsMSczYSWxOcQRyHsv0JkbHAuuYPLfhHppraq2ohZsWEIeE174SgzpF
FmbMVtRdwqRac6ug8kfUPSi00rXtkilaltMxVvVlWNnDBMxXa2K53CXtbdoNvcSA
wgDY2Z3mgyoXBcRe7djLb2Vrm7+L48Bwf954yRoj+k8IR91/sozF/ffvxrEWwvp1
2lCwK7jmoweZ/jyHO8Pcvm5gIh/whgfBHHg9sdThMIX5rbKh6V+A4PDiIReF3RPs
YXnknsw7jChoOOBgOZ9u9fpwD+ym0lntLEhcISO5mfUcOOrq2syYjJSZWl++HXkX
0ied74qXe9Fvbm2rCPCoWLDBGCV2aFCDXk9AacrYK6xXQU1cy7SlPRFyUXDQYQln
wT4K40dOgAry1qtccEuy7ZJVMXvyKtZqLReFnrcYB8Bi08qiTze8vsDm0tUDYuDj
UtTaWpg44Kavyd+a7+R8zkt+8Fx7o1NzU7v2WTOOkbra/I2wWIlgExvXubyW7nvU
xyXQTY2DiKMcM8wr9iWcxxOwcVWXJdlRmkk8WqNBIA0mnq4ZGzhi5Oi2kng3AjrU
sNAHTNRQugsLX+P8SMLFwp8ScGfDgnktkiC8BaizFt2SIpyta7edx6dJRuYI9Twb
G/7M8Z7rWehYbcA0I15QWr+0L2APlvoO1ulacuJa9U59nIbiehQuqA8taKU1NTnU
FDKlyskVASJqiL1ORTinZwgP8JvfjOiJ6DZF2XueID33IzT0dM9amsawdNJooA7C
StPaSkEFHdqWyEQu6J+BTDlreDfUBGUCp4wUh9mgC84ozItHiscXHDYnmgVt3zDo
YyotROv+zRFutGU06D3Fo29wowuZR6BJTsX5oEnY5dBLFDi6/bqJagqjONmdT6aB
8cURGC3F0nj9SSQQz0ERAved1IR8hot+zr2zf9kbKLwaUTX6npGvBGXywoFI8HsQ
xJnCXTxQya2p/ZQH97qwyrSiNhw4+xjRfU3Klokk4H5dC7V7J5dDyFyCFn42iRTN
gbEmSuGimjaRMaPGi4eb1EoHygvmKJjDMC5pJlyYhh+AeBQhbjChGfwFUQpRBWLc
0gLzsCTFz09fC5nzD2BgFG2Gc8b+69Ohw4W66w3rTdmVv2RM6bp4laVoqWUIRp9U
D42GyKk+htOM+6PjN4c4z4WlhhdGHlJdU3eJSDd4jlzp2peMW8LkGOpTsxUF2AAE
zAgNpok2/Ph0RCR8MuSlDxg87+yTBVE5QHypB1fJO2Icb49Ok+YbMocgJuUIexk1
0o/U6GZrkUHHCeFSdLrml1wNZrEuTPlvd1BZKVydo4dT8Bm51jBc9hy2cOqT2Loq
VL02ezM6Euf/GfnHdByUnQuumfiv5rz2YEV4xTR9iGjaeE9VWYRwCo7HfUQvqhCL
N5OtXtciu7Ads/lBOpHmoAohJJiABBJLwKuUMH98wBrE+zgUPK+Q9L+8ShqNTFA7
K4CwoqsrdHyUSxpN0d3RwP+yeHcdwUrwpMndSxI90dlxzLrul2P9BGA+8pHvTIYv
br2p1zZJUSUOUldPvyQJ8O8+x7USjBlLVjdWwvJ0qorJUMpGBZGV/jgiKfivxg0H
9ritI/kQk7Mf1GI4YHsh+7irlMwALDpmb81QlEDPeYXLUBxW1GJiEMF43U9xg2Pw
mq1B/azGVrgfHo1qsDXgIj7qRCLoIqqeEe2Fa/LUZ4QFoWVOCXXRPiyRpXZoim7z
Eyj8UL0MNdhUpNABSbb8IDiscp4o1lcbzrQoCtDPzXZ/+ThcHOlPuO3kb2YMLnDT
H+hihGctAPuW+SdqwHKsUkd87DSL0dCWKDMrMWSHPV6qbkvlRTcD+5DWh7nEU1RO
VVRSJTYjYGUH+QbspX+82LcOeI8WfdRbh0Xhqearnng6086QJ5bw/u/nsZGV6kKK
/O4nUtvsKkdPemrrzNGoPS7OibG05yZjT1TktG2Kz18aQ4zvSYoRPpYHHJrDNr1r
CoEF6kdE07cL8WyQy+rmpo8CQOG3CzpgRtLDfV+4f31Evdgcq5Useh3BKBnuDTzf
9SYZrd11dG6b2S3BTVIDglqmzwTYcl7pvOwHDFU0tkbEuh1oHkR//rsc84XDQsIO
KCkCIUoqRZv61wORb36DJCBkHgZQmDVZIKo4vzsws7ZCfEco2uz5pJT3jiDqpIev
jpUU29AEzsWcMrpggVehk3toxfmTpjEGahEyp9+Vf+vAndzJTbd1DlzzsYj/mrWS
K+j8bLxpxZ0MHIfIHRDlGEZ/3yB5mLVY/meKdpB8ssVoei/xlweKBV3EDwufEPMo
BZoxHaQlNeRylgh7Ut0Aae3oBuej9w/uKN+DlwWvpjZ5VG/hbqg2MrxRzNXlw9wR
P541XtcSczsjCvQXbrXwhKFYKTusQbiI1Oxu74/vpbCZLxoZXJkJKeeoJApDCCcQ
9F2UE15l5RDFnmLoNx6S6lKtMSe1I7WQYolDKDzTGG1soEwR5Af6ZO/qrQ3jg9zs
poHwHZMp7vjUrB62XkgvD6gpQs/ib/n6wjRveilWCRsboGteAi0wz4cJMqqei3NN
QMyzWIJnZVBFgyZsv27mUlxNEY3av5+YI+ZZXso8Imomis+u4E/XQNvqHlGX+rOU
fstcvG73lhsd7fvYobLICdh8qfdZ1QF7+iCEwiXeC1TIdPKcRZv0anvWr1s6zWX5
T6TzJvy5t0LRM3NX2mud/+n/4Ea4b3w0SGPq4ezJyR6jtwVRt2EW+sMdg3LZeffG
eyfjhQS4hVY2JUMOKfJMXHJ9+Y3uDFxcQU6zc96kHaMdO7mAoiYtuhB8CukPIJ03
OLShuFi1biGxT+TjE2s2whb9qBheS1QiWrgDszatM3o0ob7T7CIM1ysyAYaJD8cO
YAubnxvKibZS26AIAThUjDE3BoLCIpy8HTEOwtOVF2rtHD/97Gate8BttsXf94DN
LLpc5u/IUJoL27/v/HD8+3QZg0+3WkT8WqynCov/yY1MXBqh3sJXE/ClxethncMv
5ludFsEf4o1GG0iLkSIvW3NXbLN2thbuicDsHnWK7fQvJRqGqYoPN8ZyAqlEeKjt
zrJvabr7dVBN/u6usQQeFex/qn7wRVZK4LywMWg8QkI7nZngt77J8CNvcrmPembN
rGxE2B6YRSAAyJt3BU1g0ze1tEMbaHI18D5smCZjocUVgVsPVmgcegMv2gw0nHhT
W1mogXBq4XTxxynvX44fgSjFikV44eduUb4xE3ztoZxQskjMF0JRWGqbZEWeC/Hl
0ixT6lmVatQX4/7OLuv2eBRlxheO5aTokmrRPMPWLtJODRYI857gK3VOB2TB1hMb
uh5mGUzfpbdQXS01MOp6MgvwpZVcBNsLx3pZl+RtPxw4h5OVQK1U2G9oQ8uK/qM9
devF951YD+C8BB4s+M3ZHVPurEd1EZ3I1PSVM2Aa7ZoMCsNSWEjr+3u0pF+HSlYk
q1qNP6QvnBlnIuqil91UiKL9N8G6q+8GZJgX9JRY+4BNFdIY6Lc9TmeBAnzBr9Fb
zKJNko1z8bmySmcmtPDoON+WrDSZ3IEYeC4/ZuSObsGiK2RRT6lfwZ+Ym+LtGJHP
SbWzYWbgS83RHgqDeXCeIQWZ+Jux5tntwKPk2TJqI5mkx67nMR8q1dL1NVNFJL9B
5MUVQ7V0rlZOAi2+P0q253QJ3RoKWsW8MQE3UdmmxyT5KYhjkzxcjTbVSFIc/qJ7
Cbrcxx2mEsZqeO2y70lFI+mmvVFkitFxzpXK93lUAXnFMOnhJril1DAaxdUM8xVg
aiNbdMsTtZOafWbwsRj/T5nUmW8CFjy9aA3EZ9MdRfNp4ki/NA4bKUa9K+sX5y8R
VvYOHDdX4qJEeqmb7IS4eFPjZtNM3pRnQ+zQTAvxD5h10IsOv5rvoFr5P4L77Yz1
w8ZXDoVKgXTIYJGUqtNBhsLVOeJ43DBFxrBwExM+1nVvm166qeN64PeVnnW6BOi2
3nUvVRj3ZbHEKkMQtUR26u8PGsAInJl0+T9ApuV1l+ZsozkYl7X4OUsY7FQU+n0G
XwVINSLTlPyUOt9HYyBEVpCyBRKI62ItBAc/Z96BKyxiB9/PQmFuUxYoTV75N6im
eeIAbYvVYo0ZFYPVEsvGVx/n2qzvSf/1Nd2+J0PjAhlW6ZDPQuklfMSjg5DAGVcW
NcjTO5rxM84G3Gdwtu0hTq8dkKeYWVIYT7lUcKfROkKTzrdE7QCwMbx2xovimE5U
SckubecFuHJy6ODYNOqhRtTFnd9AdH9lNu7ekXxbllY08afRmsCqLTVXn+xVUvH9
Yhxc0RKdB9ZsxIvaMqwDoJy1SfsvVvncsj+yUlRGF9MG2dqTG5s4nyv3b7mcltxF
4/u0xqD6XCgsT7SPBjTc0K/GrsW6TW4+r9DGe/gQz+OnXL2mHffndxEn+jjmhu/0
CH33g5JNa7ffzCN+CZyuZi9zSXiLbhSqDjDZ+WbtKmnl29OBqhQjeL1HlN8PUnOL
gDrrBJ2U2oz+kp7JvaY+u2HG6L7thL2NjIP/XykvRqTAibJ7QS6slgs43EiCtq7+
Uil+fXIe3dKk/s7NueSAkEq81ysupbIKcMEfTMBbu2New2Sk0g4w+NSTkIhq32ZT
URM8Wdlbm+F7cVQKgJshojb9T0bIK+eSuv96t9whDncOgS1KdTON4/jynKW6ae8V
6Y4dkInDxsWloG1QH0VMdURTDUm2aoQ7T3T5/VIUk4E1c5EnwkXLhad5ZJnqnSun
FSmTznqmAM993ctozHcfrJzcn1ScmXT+UqQuSk5JrXUPG8lx9vdWj1BlbC8EqiK8
75V5CTMmnE7IgEJq/uKUYbnfLhIRzQYWZoo4JtcX0cXY2mEGwIjR5vWCzgnAdBMg
4ZgCYNeMQbWDBQPXtop+amNkEevLH9coU02O//6HRz5cIQ95fkAGPo5yzKPjY82C
b45diQo01zMwkAE+FAtaQLjyUOA79JRIlwIOz2VTR2m8x1c81dMl49jDIRkuX3Fv
BoZ8p/feI+ZGS1HddfB1Ok38dcXo33GV27fCmnf2ngnDXKVE4aqb9kcc89Qf+Lg4
QbkW8Bdwz+hff88vTtyQMkQMYVlWHSjgEj6ztqgg/RQfN15+fPE8eFCqkbvT/H6w
S9vXpcL3IWeRh3oUPRGNzbCn3FmlWWL9BOvR+yLq4HhoYNOqkqTg3ZAaxFdgLWzP
OC+8+eUjxSK7lcmUrEyjkkfxyTYznclHVboF+2lSEoDd5yMZ6Wg7UvWtASpupVaf
k3jf/n931n9hNq5Wmht+hhPjzFydc+tasVKH4x3VfNSVVrV6sPdTP1vxGgqXGz5m
vD9FwPsdUzsxKbd7TwzH+6QtfspAU1o6/Ce0nEW9atmriKtqVKZD6A+ibIpIkhj8
IYxq8C5t7dWO8t4R69RQukmrtV0rL4lPc/2NWCLa56ffUOH5p1Qke/du5iAl8ZFQ
R4cBIKA5j0q3RXeyJuYH/8Obbrpj5NxUrKXuevnfVwJMXxHujOzqbVs/EzKDDrDO
8LGTWMAJgk343q6AKOY7ZsXSyNJ3n1tUD/lvp1Ty7S6n/PIIwN9bckUXoe7jKrqO
DEwTpkO26vurtZnWjaLL3phG+bouBmG9xJV9Z7zYqxEWan0PDKXu/2SyYrzhKrMO
tXC9jkds5UbDlscrn23vs4cFcCUlJLW7qWSI9DPIUQjTjarTwuW7u2grj2EgJh49
Q8fgYgnR/fQ8jkx22YOwckc5EAB5H47DYUNDiwZWgBTHhVzgMGcvyaZAItDQHQyP
JgnoYFlVvY0a5s0I8vZbxE2OwqXmk2WGe2HLOBx5yk+LtJFXxNi2FczvlrxYJjbM
6bveob2uW6N5AAqm6/TOc0VnSeeFHi0YehoS19Dw5Xuxha2Z81KcjzQtfjiZz6lX
j6reCVaLv7FW9c7NU2U/MJXRu8yp56hcGE4US8X7PlgvyCn0GFc8RiYRncmqSHQe
e1j3+RfqVGTbFOMqYMZF1oGqXzOLi65PHm4e2QYb5odFyzM+BvUORDt4x409//jJ
indTUXbynsR3c2e3BcY6e8v1180X0LhoFznZcxmaTsnXgc3PSr1fPDPTQaS3z+SE
RWON9Tn1MRL/h733XNWNOqJ7LjiTsGEkhruneBNf7EVUQJck3QQq6aUDJPBd4EbB
XVz8B85PkbaPZ1YzjSqtshkYCxbJEtPcjHym454t3AGZHAadt9QvmKm2F/7+GFc8
iEXjitLv+G5P+iEYHfhrknXeglmUZpDfjtJ8JCmVrGuOwZTsR1hjZC03x68guAg3
E6iKbqINZNI8tEe0PJ3iX0Z6pUQHxDZAjm+URYESL6WPJBX8kG3jbpNscdaO9JYH
T5S9CvQPm2+YAWtRzy22/ytD8eXJWQUYU/Cjm09Ipz6tZBjPaInqyvXEvXLqJJAi
jwAeqrDnhfRu1vJ47uv7BbXsgjHFA7rAfRUhazu0oziAwrASqPRYNj8ot+CbFXkz
niPac9L3QPq2EhJetZWVdp6cuivUG5rmf77rVbst35UvMbr3QyyootmnneFerMWk
QX91fKDMWIphDNRXP2RntpU75OhCtJsiGVb8cmOReO6TarCCfjnu0phf4o+qIod6
ejvm3D7Nr3njtXSgdmNk8bdoMsHPLyR91p9/9PoetZxLy23dxfCxKSd2Qglu9iXr
iNRXFC9bGz8lhxl3EQN8EQWrQnrjAmpqI4R2VBB5LJi1Fjen3Te40bzPDp0WAPmF
2U4WLPV/AfyKef5kjuLjMP5nAbUX5UQ/6RAQmK3h4yAegp4+hZHb4BumsyOfJVFG
qgcFrSBRS09X+kjT79MncATyO1XjcDwi1FZ/5gb5PMITcKYwCg4bekrMVjhFgZK8
jj0fvW9Zp2nt4KbcsJaj3RoxWePGFtrzpZ28lNuUsfjaMxqU7Hr4+kIGire9lq48
/m06Xw0+2py/v3vfKzIq24jK0Ggpo+cZxSbAzeVMUvhecYbD+7V7bMKhjyxuHxht
OR8MfHD/dcNyGCg9KKoBlf0dbQV/Z14UwSCZ5mfDDLD1d8NAqQWmdfeZXDMTDXiX
AWEPNfwW5tWp5gNfyFU5Gh66pZEHpAhuO4RerGCLLVAK6pSYG7mSczc+Mq4dcNq4
sxngQ9xfeG9pbm5Snhk5WmBCnuoKw3GKS1a4jIU22RplF+azjW20TTPjXligjQA0
JISddMYCLryRw9zrAKrw5jir5nXSxtrcS7LnwWjHHDQdLokk5HUVzFJM0b5UERdK
V11XNnU/VfVoIAw3bJAa2UxmqLcnmtowde/z8hrpq4CXw6O9DVGZZK+IzGouJWAD
WbbZBK2Yi+Ri0qoyeQ1znemdJbwuoTFpNnPo+ZrIeqf/RVWrw1lwpNE1jWMihsqs
eZKVjK4rLwnlLvTjEIRlyhMMcDTgOTDh3y+3FviZxmPmFA3vp83k6zA2syLIk8ic
GYIwFLEPZ6mT8+B0tocrV+0OeN5/cg0TxtfuxxYROr4TO8bjHe9vf2QO2gIftz01
1OPEpZUotjV9GNym2yfhndN0GuY/8XvSG9kokJS3VOmka2LbsiCqkQIqjYXvhdUS
cajBsMSJQk3UDDanZT/0HOAD/h8E6XgpwqIRDrZ493Wwr4uUznixMX2lx75NKiDB
LcD0O2AsjB+Ehg4jQ63y+xZyf0HXYaHFWiE3aLP4xu9cSx31RFCzGXdo7abZLe/J
oJlSMEes2sjRnXPJKl1rWlIDOhjdfI4uBoLU5mV7KRd0Y2tNA7aGutYSGn3vXGfe
0SeqwIgxyRbHjNwrEdtHRgCrHpmIfL2CNBEideQ/oHvC8YJ4xlFWiBOPAaI4Hhyk
Lxilk3uBbnhuLII+hmbIxbonwsocFhTUvvDp8ufj1WiotAUzvKM13dyROAP4kgQR
K6xccU/Ln0c94mIpGpHgfa8lOocZ9s4iYQhGxkw2Zvym4pbT9qtelR3dpfGCFkXZ
iJDZDlqfXsyiIKLllk48EoI7qHImoVusI3GxNq1d9+vogolWHvphanFtqtJzOLSl
tX2K9yLD7+A+6q96slobwdTSGz/ic6t5kBTt7EXXNCZgwbc4W/jkU36tsgcY3P7N
D9htwV0hERLbJC63KuBYY4if0fPC+b4bWWipBUxKPajxkiWYyecbw3GHec20aZP6
RVtCmfE6bx7x6U4ok6hNzR3NELWgEMycXvkymOebJMuQCDNqJyHLqnljZpmdSMQI
BTvqIxinMncCE78b7TPn6D8oIRMoWQIR3FPICq4xWCRNzDpSu+bv8FKdiKQvKQ1h
Y2anWdC2XGwZe0UAN2+R4J795R/cYaaCnk/tMj4tM64BzUB92Qc2aXvwOJmHM2q0
jcoME56aMfN9dsg1A3+hzmU2dPw1tNQQ7GZ6FmFpUUAA2fv4Qx+A8kWhZv5/v79W
GgwdwdLpG8syuUE7gPXky1tGXRXWekAXxZuLNSWV8IqLBpWtapTulwv3EFppjd8I
L2oUkn9wtS6YrW1b6z46HFsiJEtziWLzMaTYXJMxFdYMqnuYDZqSlaFFjnRurdQB
m9L5Z7+cnyHzkmxu7ooyRjqwo6ZO6otVP4fyvGVqJ4Dgg9f+Hw1R1o7u6OuR0ZIW
GB0nfB1NVzEUOUcSeVYaQ3DG0eMNP+qra9dyWnWLJvrT2fphKk/oP1YHMuW2qcGq
1A9HktvXRKUeC5TS/dDjTo6B0Z/k45+W4iC9bkpwdAxp7z1NhyPbNvFhzkqI9K+z
F+UytEDOeBHv/gHSkyvbK79how8jpWHiDI/EVLLMi0od42CyHCkgDDi1kZgkRT45
MI84RmOfIac/4UDlnc5l67Dyc/sq36QUF7YOGPb9x31jTAOOJiO/7WU/NfoqvUfG
If8EDPfsIShB1cvYRwN6oxe3ztUWwKI/DWEfdbl9dJ9mR6Lv+H02g4yf0DZjHgB+
dv2v7GOwJBEzeKkdnGbJ0VBU3o8DLAqIyp6bq+9Io34HlhxQrFLtO8eJygD3MdpX
pCOOEi2+7Eq+lvZ4h/ymEKrvyN78LKGAsqYYrBJeGqFcNdBH3qPzh6qe1/EQ4GVO
F1twbFyKtheHrtO3WTEcjLnerwViiDHkcAdGhIILFsuKAYoeQ/1goKuiapdPvxsY
FBDKYIpHoC3UsdTKQXrFD/DXD6K1d4QbktmW8Q3H99p0rw/z+XI1Zoedk7ZnLHN+
BPn9a0Mg1QTTHIOzi0SDN/aRLW+bIPIYcSulhLtd8awDYeYi7ywHw20tw5yIzQW4
24G06vKPktXthTkuPdU4Jb+AjN3mUIawKJ2ZkVWxDWkK57QQ5G5YXgbS3UrkiwmK
DY9O6V+PQTyr0wGGagg5IA/1eeLVBdQWJFzBNlLxIn29GVs2d7s9KzYsZlQ7CB5F
BNJMc+uaJwKT8bpOqZXUx+2LcKhr087eGxwPTBWRKPRfqWIcsbSZvUoC3/CxZuQ0
vqTM4cp4Rc2vvRnGzNZZcrHQXOhcvILByxv1EIJj+8irjMW8n3KSESplNokpMI6G
4TRzKzoC1WVEMT7pxwU+uC3xQMOhoSoVujUr94g9ABhdOmun+4QGcDGa1WiFfXsL
pxEU27NWCB+TSHauNUreBLgal4K6MzxxqDciHHj1C2tnrgL0f2RMONFbhS0hXVay
z2fN3esxujhTay2TNKuLykCTrfWN9LvsW5+Ft7qJEmkV+9wL1HtV8g5PNnkCqhsX
6UIFKfqtty1MjFylOjLKTmRfo7oJNbUNJPOS4jwvGs0G3lbwZL3NeX3AAqAojVkA
W3JYCnhEJzHe5Zn8m4u/lnsbw6EtLGpVFI29oY+9O9uxy6nQsD7xrEYTQvdotkcN
NAf/vLGbuDAUimQ4QKso4LWNGOLbcif/TfiX3YPieu1qiF5ERx7NeRyiWMvm0vKd
tjZ9mYq0aB29XrYE+S6xOEFihInpfk49bxCBSfxusUUdTncljsBitUFY/8mSJwHD
Tdm3BufiV/+t0in1TEtjICevlYNA3l4M+dkRIzxD6ZmU11QIM146UFlFCx8Ltteb
zR1SSddlZqKv5tyTIWiVgNZSpltYUGi0CzqP2f8k9iUma+Nn6OYE7U9n5Z1YVQoL
PXu1oEmOL4bEg08GiD4TwpIki6AuVFkjf86k0Z+eBBpoY4zd7Pyz8N4HOPmYAllk
uxvqcs6PtOBHVdt6dhVwT9nTXrC10zHH/4JVpCV63umDehb33h6VhTpIrmC3mvyD
blwuLGlvTRgw2aZGvp7+3M4mx/8OsDB/s/9UYHj/YtQRDDecClgczNWUSbqVWZpj
zjtRUV1CJYM9kfnKLJelXkYslP2YM7z6EY5xWVLAbyUxtRgBKD8DwrEhE2Xncohe
FTaB6w2BCzMtBYQuc25CLJIBKxvTvYuVuIi2OYK/hdZt+97wAdYTlpfp52fkduXq
5IgSGoZSlg0j8j9ex0cB4mT7JSb9AJ5QR1CmT8ATFPr5o+fjsFAyM9lUwtT7L9SD
69JS9SIvBwMX3udB9Ucd20clD1fEj914/3dHSet8T0x2bbh46eSVRBC8LK+FsJaL
cukzRD5QM7hFrn0zXcirST8ZCUu+PXbbHPR0tgruw9yZmuR06byYZhOazgNsCQ/1
L3WjUQ7Bmfdo123/FFA/mR+BlR7UFesrfEFp48WFQfdqghf+qx4q1BtxoWPtmBOa
xfTVSfPqqWcQbaUcjCakIFVGE80Np2TPHc0ZLzVpRem9tK6JVmpC2FoNJ5CgIH9n
nfxXOokm+G8HUOulEhjmQ1f13bQWstL31ZmxWavt9gqtgdd33F9iFEnywMw/deak
H+NMlOMlVOpJMcnIrBXj055qn72uDe8PzM6fv5Bp3gjZXH6QU2hRdg+dmIUPKui0
tAwgH/hjXvRgQzWnUaYhTPcdOpPF4w4ZmknBeC9RSuyPzuCbneABrhmGV4lp6RKt
OAzGNskfZvnQexBg4n7ny6HAOFhTeM9BW4fbs2WAQfHHRDGHe3Thm9TYUdIi+u1d
1Az95eb3JnItfNeLJcIFOTbJ3eHKXb/Y7o8XEeAJXg8lMoMndrHx7HYd9GuaQTjP
XGsLsf5FuawEdV7YJYPygBonIfGXsb5DQaLCmAgN9552hYX/lTRVBHhDa/igE5Pf
dzEcY6OQybprZT36bnlE89XurvPX8Z7w1W24Aey6sAqVWvftcOAd/RnoA42Rdtwc
Y2hu/1fErspGg0p2D/EN3AwCuDJgVe3JGo9H7A4GYiH+UFM1SepT6ua7GYW74J20
CRSW7NWtZJbdyWPkP7kuV7LLIOmgbGUCNtL8o/P3083gh2kjVX6BTgS8//bby2U2
FIAKlFA1M5xqpS1RNQ4mVBeZAOtdv4k2pncQH9PR5FJPNq9h7YPrmqNKpgnfXCE9
zmP+vI2I3y1QVb3SK+HWXqMWQYPni6xbkrZA8X1WXJCOBud2OaQyfrCnnqflJ2Yz
lw6LLuqld2wMY53rV9CxO6yDchOgx0oNdBfj/tOWQJgiXLIerOqiEGNBfZzkKj4a
s3hQJOtQWHfru72b4WZP8p6jRo7TwEwOoAEjxE0UU05+VqoOtjgMgznb4ntkaww0
UpGiqsGNz6aGCpAMQW/d2NSfZjPk5bNxqnayqoUuGMO1i8ZtyCu0gaxZZzynGTX4
S6MT1BJIMZUEcYebeMJ1XXl6n90sdqn2yM5BAY3VmsTulqv4WbkLGaL29lkpqmy/
oBG9o+WXDgVulRGc46B4GrJ2r/u8YydWzZMMpVWtTW7DTKkyLHwhytehPMZstKNj
wOYeDWX+Ebb6SFitKBbO91GF6C+1pGr6N1EmxR5mj3i5J4iJbhxbzx++MUQdSQTL
l3bAUy5pgjc8rqXZz125AJjPrg0Z07MOuC8tUtSD7KR1PUTCtRIHXvUvT9Q8Sj4S
7bQwLwSQupa2OzxVwwG6CYsoiNIUxj3Kux+kvV7839VtKJ3g+QKdamIHm6LASQ94
AzGXB3f6jIugz7lkhYTvm0RCsrl7bwox/rcdnNIodznz1ziV/bw+ZD0EEZYBspZS
LKcRO7zpX+RHGnoj0txRFTMXr/zAUw3EZ5MrpFIpdQytmbflTXfpky9DuHIQe+qf
5OdhW8xUtE13X8XPrpgOt8K6YQ4U/GSDEnBl6I0egfTkTLeXThott4KrgeLKqQCi
1hVpoMRmUlHw33blNYONK9k8gMgzDPb5ttja39YSOfRTKLsvrMj1FomISL816Ijo
GHUkoFBGGfFqGmhZFr1njK5Ny24TI6qr/Q+WO5GQ0xlcwsWSH5JT+tzV+mQPunSM
mkFTQ/x7hlrt/vR57unFN+5L4GOdrrByZcewfA4Cm2D7RCBIMP4eX3R72nWOXp/x
iocimzkVHxq/MNotE1j7rmkq+HrLT24dd9c5wSQB1GVgCF2A/2LJ8fTlMX0mEKvm
PDPxcSRNzWFfBoLdu3O8VHO8xZL3vs5PkZrBlV4TkaDbYHHb+wnCpZ5IgoPMi1jv
mcJmsQY1d6o6QEIH6ZRI2dWMxLfazEU5jX3/Sa8r1C/XUaDpKa5nCXp97C8iYciC
R1DWDoPGETQUlGhGqae9ZZOWO6kwDNKrKPGGnpQ4iGgJr49DTOlp4iWjduoWjXAJ
H1rSX4vE+jtBEwd+FkqkKYeu26hbcP6TR/qxZJqBP6fHE9TfQjMJJKYp1MDkn0cv
9MJQCG7OCY6+cr+/6x6HXhQysKvXv7ToGrNR5jbNZAymhCT59ytqxhOk7rr7TiEN
fi2Jf7Xz4A1M9PdH8gI4O1ss4BLmWKrT5TXSVZBQmmPCyA00MDw7tRIHjimktsoo
8u+RvNQrEO3ubEPurM2LLYzKKm/Z+G+NpVrt1p+Simm9PphDmPScI6M6/skcn0wS
LzVeaYNs6trCrjHwNdy+ZdD77euPPIC13liJSic2rucvIADQTf+b/bThaQ+tf9iP
DudN9+OMsxDeceX4nHjY10/QpWHnVzT+p4qylQVOrDsiH3tCV5swGzO7AYhrJukJ
M+1PCH3jYtNpMZF+mmYTrMFEZaToQnrGCwgv6b0WQiBKTqeY8XIsKCUxzh8CDSWB
Ujlg56MDO72aPDZUWWJlwpsYni8U82wZOe0T/Iu7W/RhPP8i9eeZyRjhDQTclv2z
VV+OFhlaCjjOYeUjw9oTcyGYJXcqx7LyC9lKxxjkrWUrs1Oo9J700uwDXMucY8YR
rLaz6yLr83G33gA2g/PG7MCJjAJM5Qcg4bA0HE6rszgW3KB3bJ809Za+vR754quE
EaSJmycSlgmKD4ZSiyNEzDhvPr3GxR4qdriMsyru3+E0Hqc5roqho3K7DouqI6kY
/UYtXt930kKQrqgmitW0iMPFwf/ZMrhGCoC99BsYZ+bW6ZlCqwgY5LUw2cYR3Vyw
/wXKcYz/jQNFyoWEYae/m6X5t0Yq38ijuhRsr38f8nKwzaLJFyiAJjMxG8LCVGOr
Yv3J2NtuJ9SYF2qMepEl4torQg1Qe48yEV8F1GFMTt7k/IKShbhW7YsiRYecOSoN
8ZwN6VzERynDnBJaq0ZZUYUN9Xkm6ECHu3ju/oiWrnMeZMVz5TKB3PybS240LSMM
aH1b6hcXDVl89/nC0JQrvYNpDK3c7wCsmypwVGZD7g243NI3dD0/UdlCq2yjMLcZ
/xjOSAm4uneFM74KBCjp0uJiZjG1GZ0rBFMDOOYiFo42nomW57ZqifE9OkOi1bLi
y5MJa4AJ1H/jYDX4uMD6aGj69iEdx4V26gyiFcaG+3Sg+02WZlEtXO9Dqmbr6mZb
00tkl7g4I7qZvvpRPbAPjy+rssqFL5rX3GBzkfxMsbhKbymil3ofNXh7RmwzVF/V
VPavhdpnNYEvgMmo50p1qvzNlC4JM4lkBghwmSKTQFy4W7oo55qbuopL4kN6CKO/
FeQ1x+QowD0wZ5F77G5n6xig1udPCHzLbhzWRO25bXtX1gd9nRjmIRDWbR1Nu3d+
a+KcFCUMbf3HPN+ZIpvx7iGl4IhjYFhPmXeQ3FsMqeEPnYi+7mKs8CRuJAro/mHL
6nGnq9rmw5XxzWNcmh/0p3s0U4OrZgMqz2qfdSO04AMemPjq5bByBTxtEmh7XrDH
Ga+vrvqzaL116rIP5av5tsaLMAzXNENUkExyft5n3cEx/9umDbC1Vy3PhG3Nmx7e
sCWogw90bzgObI+I2/wEQGJVG46fzBFJ4+nMRmPsQGPS4GfytHIxC2I/o9iHejpx
p8S6B9D+JfCLc17ejT9dbXkqFfkXvYAVNBC6rTITXxuwK6yQdRj+GngVg1QEJU5q
IltgJyy/21Zsu8MxPiKETG5xHDdtjNuCD81vxMmxBQOPdu4ydut2stOmq/Ve5PWm
4s1YTdnG4gxL7iCfV5KDwCW44J12DxX4Bj3T+PLgGhgZf05QYOi8ik5pexUCSCk2
DyKfxl6B6gnQwgNvXZI9fjJV3/1H9HNmFscokIB4zr27r5LeS9erlWg0qrgkxJ/f
YPnVbQ8+tZwcC1oD5PLkc1P6c7+p8rdQbxEh3K7Riv2aS3BIpU0/avg7iskBMx+K
c7nPI2HHyRmLxbF9b6uTTb9EKGHxvXwqh9jjb5ZoAZMCprsmvsjTadvwX408Tddh
AEAJY/YXcBkNB1pZN9yCwthiR5xWeGFuzHWfUbRZphD9kl9qpzEmOuaGkguNPei5
FOlZx+wMQrq95QtwjQ2r+0rb7eGTMZ/IouEmL+/a7igX1tkkVpT1yXoMS/fl07Aw
gJDR0J3IzRkLSotKkXkIygB7wQCKRcfXPtKQ3TimNWq9YfWtnVMhr6f5aMdquOx1
DsursDUwKWhsVuDTUghB4tdk3XDUXgE+jy3UdAj8505e9EaqIuLAljWRIunzhy9V
EO9lc9yp0lWmFjtBvO8ZVZw/+QS3t9S3Vn0NUEmygjcoxN7b6x+T8aWeAFwPB1VB
3JL0EF8XYwfKj4n3RNLCanAYeVuMsnIezbFvTcuHQ3vzsMk3gaOYUii4ZzrLV8jQ
oEqOn9EKz/UP/Ldj2KaENrmj9FigloHiO7H1Nu5RNXMr0PM4v8DvFMuTm4q5OSWS
eVFjR+B9DX38cwJme/5/BCej3pejlFlHeCbClJpN+ASc/NXnLEZvWAYf2TKcjGbY
dBjlWdRnLmPUC9f8LCj+mh0aUcF7EPAOXrNrNBdB5RvlNj0N5LgGRLb/dzeRao2G
DPvOuJd+scKufTS1dCkS3w2patL4tV2l6OozRqtbpi5WG/oMQQjpKj/AY0soyZbI
yxbOgp2NXjZ6NDPOZC8JpiBg0UY0zCRwBNcyh6T5rjxcriJgXUe9/R4qor9quOtV
hjD6O/f7pPlCLIOAt6c65f2uKp3Nzh2qJcLRMKy4xp6Y10onc+Jq/Sdo9nndAGro
AIP/2FoXop8SCWxtEdIskmNHFcvkk5J0AKGlxBIRWwiw1u04Zpkyv29CtvfsunsM
Uq2pF4frfQQg9AlK/dXl/rPiqW/fr+bjIrxbU7aqQFyOL/RaDUcoMRcjO5fPcFaw
HpiKQ3y6oGpo26V/apHY0qkv06rE9j+gy4pE3f54pXIQDjoPv+tFukA8+c+92ftM
kAXVOD5oDEkE6vUIriwUtnLSQ5epiaJBXvNh+SpmnTlgARsg2Hme+VIUju27IgLy
RvRAgXHIfEhslEvaw8v5OoX2h05DNKV5+D1QdeC3PIBqgTuT/b6zJmteQ7h4k5qu
KODZzz04jFDef9+qbDGElHPRIkP69chNxmPM0QhQUTlQAd4CxulQArwhFCjYI8F/
a3bsIrs+FcNsoSlH+IqHPwQHuIHzaTWADbZMH2+gpO5ZiN8f1/LF6Wj7Tgu9xfwW
KMIVFDgIqbHi9RiLBRuPLEGa0NMBT4obi/noDHsUZ/UUcvPDgCOpf5BMWrFdHg+e
HhawNwrqWaynGFWv3aSz0i9fSNS+nyUUyJ15HMuEh7xmaUMVW7n5MrLysikT8f0U
vpQYckoS827KihpT4jTjuEE1TsXpgb5Ew3fFHM2kLg1r9gGH1nVPtKVqj/r3xFcS
ogzt47Z8381cCjFjDvKkwF8oKhg0Otin1ikMl8/4o/sQbP86x7a5U/sHA8MyHdId
jp+3t1+E+84sTqEVB8SBsyC8CdbF0jq7JIKn4SMRMR3XUd3kgsLfFennHX34J0b8
RqF7SKemgcyAG+cisPM2AvLwo6suPEZL8aVeaXhhrZZdP4vws+HlPXLA1mSYHryv
wA/tn17tx7lRlEVPyIJMnQarwuHyMOLE/Gr45lKE84Xm+f+LLliAmZBqvVN6UxcM
HGjMLtrkH0u8QHsxQspohukKH2g3fC6n/CSuV8WO5uZ4jfg8rzbyq+zZGh97U6kn
uajU2pwj13zQ3HPzHYFN6bxHlAlq5QFLR2KZM/TIozA00ND9WbOGSKiXkaqL5uvh
C1yh/30CPVy3ux8vkL16DDV8CVDs3DiNZj1loNwTVTg5zjkByKhAXFF0HEfO1ara
6BYhqBn7W8bHn+2Nub655CQ/Lh64KDmqAXPZx3Nddj3fcRoQB4bjw1Vzauv67sUn
wDSndz9s1d3dGpPgeXxlIBGmXHyfdOBpedV5C1F+uMPFoc025HxuLkEUf4FePA9+
pOZ18y2DLGWUAPw7KG/jD9VcTqpkyHY0jvK0hpBKvRy/Sc2TJMBWUnt45qVNUP8Y
nUZT7Na4rWjNQ1+Cq+HzmobNs1YaDnhbuzOOlwV8nFFWkeF3NOLdxrOFhoysWRDH
ljkF2TgH0R+9cjlT2t/N2M1y/qSafWBftH6Vdjv+slsM7AJjfT6aTqDUtSojIcnz
5H/1xpIVO0ugoyM+cUASBFgs29ee80Iwm6i38uqRk7SVvepnpOAyDRuFqnaJ1L6R
bLmxZDaF+XE6NNxI+QVHXSsoiCGNaXI3O642rQwpwbG8lzM4ssX7HGgzSSOq55Ve
zOAHL9T86KJYKIQId9vMYX4inU1Mo5xYWe2ErNqDobf7vhdm7NB4DVlNVvID7+aV
RTUHx/zwdxjXUdC0kbFxCTidUl2HStk5SWnylxqNMGtLpL9xEDf12Vsjb6p4U/yO
SqRf6IjEESymoVxT5zx+/u1V2cO3ZBdPSPP44I7cZbtZmm8rvAVbiAkKLVYidYXd
fKG/kKaN7QauSQa/upiV/PEyOLr6XY5WaZc7kIZR7IIDlJOQu7Q/g7a72vSIBZGz
7/AUxn2MhDyqauB+4xQt1yIW0D9N6Jfx+1cUwY3Imau2D1USAIfUI5L16k2jEzhv
XSM+rb8pd6t9keIIKPjchLb3gMOCjm4ErP+Od990qhkWzY6kOExRwP2wDhqff1cc
RsMQ+4h4p9JzD00+NfLNt47sq8A/p5qUwD6MhnNeZHlVMHKp8OlVzOsg1nm3gVLS
Rnhn0DzDbARe6tXPQIvd7DmVWNeEtEAIsHEK2SjyoXtujxcySAbGTtsr0pOkiQVC
Mhb4Bhl6xIWTw54HLlbvttSQ4bwElWg+0Jm2GzkXVeaMDCxuAK6Y/t625Lx5Sh35
midMXybdNWg20CvuhjAkFth43MyX+Ve+84r6JenYFXsDkhM2XConfN1n5KEL20at
OQ/JlvJ4HGK5H9boi+2s0qUlYRqp3REGcge0evUPChdsuEmFHnmvI+U2SPOFUfiH
keA+L+YO0GmOBq3DApI829zOppP0sD5sbA+oT/622qQ4SW5hKLZ135Swh9jb0NsE
JVlBAuzLEwEI66+i1+bwB94dt/1G2hB5xQZdF0C90M97hnMfTbcZFYf6lLK4pGJf
4JvOYZnwx/dOoSv+ePdPiD6cUwXCZ2m5AuVuVSmRetmpi/9FNK0lFjZnBBGVphYJ
iyx22VQfhiGeBx38kDM9zmzKJbx3Dw1mQGeKVqxvey1Vt1RvLiTbVUXF7hGmk/Xu
V4eBKPhewo+IzhIRHL/YgI1yrPf0jYADh4elVdR2mGksCFoZZ+xyG0ZwUEkjbtfZ
DHwXX/nH9uq/iAbMuGAp1p9XfzzRV69HilsgQxgIWDl+uSwWnydhqqqMSQvLwnoF
3BCzJc6A/lxOix6KGLWQKJF2oCUtKMyr/mBhpQHfHMQJFanAtPWz5C3Lh6LN4RTW
nLL7bxguiZKCIYdAvEsD/Eogm09AiObjgenyEYgIKFsB7XEqhsFNMaZK3oKN/R8w
r6UCxSbhvrn1T0TgsgI+PJQnn6RnGpHq5PSrjKBorjdWsp9Rth4/uKbiQPtVFdsu
2cE1yY+TOvqiJY/3DDDctZgejslvL+legExMbllnr1ArcyUePSnvLKLWtqocEXjV
iHRiLYpHpVLB7V6IqbyKaHvTVeJSgvTH+dKIxeVlDfE4qni0eQ+LGW3KyiyNzyPK
0afu2roSDYb0vZEHqO8C2dv7TePUkZIHsEpBJ7gEllNBm1iyGc+r9vUr35Z+zqi0
s8H1lRra2uSGVGS5pEjdfr99YJ9Bxb6XcZEegQkaBctGbbROxGRYeOKyEViiBZdD
Khz5jiO5scrz5EloBdTvCKDG1TkI3kCL5E/oXelr4ST3HZ1OACsntPNtCPrYx584
thw6hHV8PnMe98Ie3XV+FPu2+On47FezPi91YeOP/lvKQp2hEIIFQhrl1lBpuFG2
4DizIWsl4ioKZgabHJnK2b4Resm2xCBtbmyj3F/zw8BQaXs8E6rc8zupzhGf4iYN
MpF7unyJUOB7f8TDuekS8usiTQHDKQo8NTEqXqBCiHQyH93zgIF/741ASNc03CX0
nPwKM+uDTVNBiBF+LwtrX8Klksrn3M0DG/Xiz9LEtdgNsCvxsLdESR/orR1oTXyO
MQtc+1mPfwQ/VSBQmp73W5W/9c2AJS/Cg/JiAfK+4ECPdueqVr+UVCBSQJoSWxZ+
RMQOHDttl5W400+ov3fRty66zkkPCcFkgBWroRJBGbuhRuFHYD4wK3UO/r6MtSho
IWTu1UrMMcVRCMiVUVRtzixOtvTiaK9NhvwlgbqtUW+VTpwfjTnRYz3dgZnpI2Lc
SKEHb5U3toIBroxvHwGY8dxaoKc8pUxmGVkOwU/I41vb1v2/izYOJGrXcYsTwPWS
GY/Lb9t7JE5InHwuVDv2UsqtcUDHl7P9dwzmm7F8TSe00lUuqQQC+QV6tgMxY5cq
Hz8iEDI4EdFupR+UBPfabMw+SuWxwk3lZ3ULb02HqthTMmop0oMTeTck+ywLxWXA
QXCu11ezQd9RAo0q+qD9GO4Iww3HwwfVLxsEpNNpRygYvaqXgSa3UrNxoxSvhSKj
QLPLphcYiZS1zhIfUU3E/BDTzhxUN6IncucMnxfcwGEF0IDcyzVjmr5FZV1rh5hp
+A75OVFLyMa22mpjNTjj/MJorcnsrtGHUv+sbT0BMPQRx/hd2gUiP3o2N83YZCpl
nafsOlMiP45X0fXFwqjYOlEE/0pA7Oo7LyMCz/vnFiJCB1bk5ZM9j7tX3ubLBqoS
zz9o98yCJeinys7UQmJxsWZmQ972kyORIYEuElLvv/xS8sos2YruWgf/kmtJzFoB
GFbL8PLQ4lw0e0Y1UfFzpVAlrx5vo5PuNEz7kJB3Q01WOM9Uk8/xKorgVWOrOara
L1CqtTtGAQW33NCuX/QgUN9vIr6kiA8c6KIEBJ6t4sPEIxx2b+WjHjVZiwGKrHXg
Hkj1dMfQru14pll49MIg5A4+vinMpRBTUJ9zJ8xAL85ezEgZ2vNQQszXIxgDVcy5
nXinnH5ds6zxuue7Y+JkPIQOOkInIqEyc++PdnKtcBMrol+FV4kITOzXe19jSq4H
bBsDyYP8/5SJ5mg5cBS6GcprlWPgH8xXMldWhzw0yb0hrRBt0BZLLhjetLAlgJAA
SSiRJ9p699AtGhzX1xGddOtZfcRTl74Y89bmfXlehavEKIF9w+WpwEEmAuH19JHv
14LIW/2ONruqGRMUlbhDGYTpIQ1aLL7+ExspWdh0x/VZiBjpagNydpE5LHV2Em5o
V6eHKHvuW/QG+SUPLhoMBf2xENUz7blqD9CbV9vAvbMYnWh7+E1k2ZlKfe9AaCL6
6ZoE0J0NE6MIxZnx02XRPS1E1EzKgURJX4oW+K/UYfSIEx1dwprBwW8a4/kcDuaN
A2GmBUMBUxDYC9ZH/72GUTYnUNY6+sBbeEQ/IiMxlP1fBosz3QyV2H1h/orpkBAX
dDr0Duzo7c2lVJCPKlK+4Ifj+8jVxbmXdgrut9WLKnYEYhpRKJFcHGHZJGP0K/7O
EwXACE6RD7foTYYMoJ1PY1Pk+0QT8rGrh+/+bTJFSUPWccSPlYKfCJl7J6r7659p
cb3sTlacSFjdzRBVBdHU10Qnkx/1ohMzFpfU+NDfpi4Z5PP5Qu7IbFs83Vuudi7y
JMgmmvoYGOJ3lfF8wQpkWftl7vlHI/fl/rhSRGP3uimAw2+z3u3gPAG0PItu83LV
ZFoYOWfleHfQHO+iwWOA0jjUzX88+n4OStw2QOBRNNh6T4iYBVkduJ7QaE/Foupr
EITqOL747rOVhqITiLrE/GUmesbldRjJtRDp+T42Dmc=
`protect END_PROTECTED
