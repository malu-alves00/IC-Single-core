`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
e6XW0t2edKbIAkmuaORrFnghHikgqHeWH9z7TYgnhPpxJHpUMbU5mejk44jpjeyf
gAurzKxQhfpfuZp8t69ZrHsI5y8cSLtDzU0+ZUMjV0WrRxJGnF6Qw4DNdl/t+Nb7
CaKTnHkk9qfZlrBmS9Nwtr3RuWpZ5ElKlD5KROoJpXlxF5Med5WjqpXmDuNalnA2
LSWY117Jyr1j3qi0yEmtMlGd4E75eG3ugd4ygvOcbPY5b4oaXjSelGwUH95CD2/W
7jtv8rnfd3J4U4Pukbimwc2On9sRnM/UO91oLwvi8pcit/Za77LBuKaZI8AgpEQN
RamUbIGuF0Q6nF0Iif1eaJgT9l97dyNa9jlw4cS2zj+nJj1M67ymUR4dd+C9Fiax
3SaTnz3Ko0wLup7s5h/P1GRb1RVUVFxsdpzdy6/JoU0EbFCohM5O+yLP9NuSXhmD
WEpmtvpvBvX/u3OEtxfA2UeWiFDZ2uZxaLyFoNFc/2bOT8cqSkxTyR/nt9oBqC0n
kZvdcKiH3KNVPPZ49ubuZv/S+xvI5bzny3W4J77NZas=
`protect END_PROTECTED
