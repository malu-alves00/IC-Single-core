`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Mm4kt95Jvb37Ctc1oaiyaHofNThrhrx7R6q/9NfOvCPPweseegkbOQXDq8CS86VE
+glUVAzrCq0NXRCV+3Bjab6VhOi6O/8wepHAsVTsNh2LNTahwo8lz0GRjrFmnASr
8aUFb++HsP9e19CrJsIp+WyKQRr0QPFdcbL1/iDtFx8QQKox88If5ND9tAdtLZ01
tIoTCbjP/4ejLqEzgUxizJvul5JGawpd865zxBLPuFGgyx8xSFGUkkp0mYmWHT8v
2sWhH9zHgQLi9ivU6IkulKjGe6TcOXWPGu5vnYnaVdi3qGPpVI9JXgl6HZphe8Tp
6belBZuHgLuYN7QtMQ44eX3TXMN0eiJ0Okn2PYsdQFQM8UJjuzRMU3E81wV8FdN3
mVQn84ZxU8Ake/F6D2OjrYoW89Af3yhJfthgoTmBgNdou4wcpFeHrbt9CahPsPV9
qb84Gur3TbVMJF22pZGSJng7xYpfeUKbit/gbmbaGd4JuZH+AnvBh2E6j/tkqKB8
b/6gPilr0vGpW+7XIaoKs1SttDcQlyhv5O9d9o3zPLJdn61iDNa7mD0yr7p6qNR/
mky7T/Vn9+l5msc3S9SqyZcX18RX137A2WTol5wXwwbp7zCJ0uAfcliH6fz37f5/
Au86yB76KZmgG1FztGHgyox9upPbC0obZ3ewySoHiEslIm8AVmQZH1vzHRj/VY/V
LawriajMZMm2oOqdjBWt8oI+k0TQlffFsHIxdfi5ka7gnL3l9eqXh7GEHhoDIwBq
IYCid/0CdIUI8jaVt5Sr+w==
`protect END_PROTECTED
