`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uuGZpxw3idk9SyaXCTMT7crCcEcs/w4vP2qLctTz6AkT1SZTzc5vU1pgO+SaAxm1
VL3wgrgAMwvMq3bd2W02+l00VzP8JKHrYbckP/DSZ9D3ELDp+VzA8r5HECH9HIwC
844cMhHDKz1JxjwCm0W+vmWkzCqJlsnP8tdfNcVJNMIKexYPqk8/10LTOgeIVvqF
czWkUeJaiJpe0SxZ1xfyqrrBaFSTNyIQj6ql1vzqBpz1H6+YcWNjSM0qwFLiEIGb
XoLx7QU07Fz5yxLWWIKbCRyjZX1UNnUY07hSuMqdOfFIhUArsuNf7p0KSdWCSnte
P2Da5vYJq0qU5KNMuKsNQqTtk+zAcco/DQ/RlnXbdNtmeQLhhhJavA/aq+AXghyE
nWnCPCt5qLS+C+8MUrE+jBOqasVkMZed1WKRhA6HjavmsnnRIdOg3CFmaEqlM9b3
npBmG+pa11u/eVIRMofQGBn38Z2ypT+r8ehSS2DTJyJogH+T0k4V9AGmyLhkuLJw
yAPqIUQ9UWttATArYiljlvknkD/P1CM5oeyl0j6jaDyG7BuIpklQvZDBN+XjuDcI
/lE+PqEMq1/3IX0+6pDLDfvKbg/orK3MZiUcX3NeXYqhdDZbSrkLO2cxRdIBxdTG
7o2zpx11lQGlIyevX5hulUBnaFqbLbf6fffXuzU9k8iXPcXhLBCKF8o4ldnRjuS7
FuivRpDGr1VYCHGckZlhWjFnJ2LZzYpvhkalkdzT9Sd/KeyMu4p6jKQVlhbUsgGs
Eu0zp6DeyIW4k3J3sGRHZLVMSntch/DD8iDXxdUd9QT2/C6eTglrvi4wLIp7wdiy
soBeHnl3guHOYfUhZNnPLAFGTZYvxaXwFhlnxNnbqFnCQGshC7WrM56aXUsaN/Ge
IUOaOIATi+QNh1lCR8Gq+G4C24cOHzLpy8IAZsv53jMNu1jIHxz4yihJCbSmF9T/
1eXtujBRCyjzFsi+vOuQLZLZiZM+mF37HPw449mtzXU6Dz3MLt9i+zSG9K3YKWpI
Ysc0M0prSGtR4rsECRt0vUigCxFKqfY2HV0keiZ9QMBfbkw2stz9j3BkmWUYXH2r
rMdXVgguoZXabrZlB3I/5cVHctw1zj2Fr/s7oksmLEqkWyT6V2JqwNOkqHcEWYY8
mc/S1QS6QFm7tP0ZJrHqqmL9WtiQFSnLXWrWfaRAWF+KsRW79j3MWhiOV3lzOJPE
u3c3G9cGAdC3x1Qv+XprQ5dd+DYtZWuq9TTeY0ekxJ92sTlUnVQATmSfWoLUzouK
RUHLoqpFJ9rrlL3k5J/X0JzboJcBValLCCw7DScpeMji/W7hir3wRbKaoYJXy9wW
CE644FE1runFH2TSoA1clLSv3UEyu272K67YxP+tInwL7HzHTVsh+m+p6Lf4hqKK
BOimKaaD5aJfIrwQyxa+jbqrmzuvt7MC1lIzNwy3af0P5cW7yAvs+pU3RemKelmn
QhOovNtH/g7Mp3p/OzwPc4hMSR7Q5TcYnYkAWW311I7kAgRm1hQ5HrOcsbSKeZRi
2buQFCEVcNSbVCLqpQ912g1V8+7BptLxn/qfVln8szun4f5nBOLM8gXxZZIi1lel
GkrES/c4SFsqbao3hUy39YlydBPLr3qIYCLaDr9TaYQF1mr3BvCKYA64w9uaAXO5
dhm3qTrjtV5wr6VnWfRaR3UWjI3tgwvZaobt++aY0yc=
`protect END_PROTECTED
