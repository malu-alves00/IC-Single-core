`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Q8hW7zwpsNYi8Pmw3NrXAvHGm2lZTHrAUq4XhiuoyLM8baTnVhQXvaxa14WnAiaN
n7XDetxL4gwblcLliC9/3AI1kjOBZOQ9o1Cmo2NnvXp/43uXAs0S79AYX28Ig/3w
NRbMsgoWsdDG4QoUfRBeMtjinCnJdCsMFVZLKdpB63y0sh+D6OXK3riz6mtRP1uJ
46SAqxh+pCOd6Z+AkX7+W8yHuh65lWc05wTWCrASC37MrFjpnnNqUgYDD6CK2wfV
mdtUNKUPEPZLwp1kgMe4x9krNk5sWgOQXaRFaI187g6fYR54Y0QiLDSKzKarTac1
0xpmOTNWkq1jEdKjLxjExYg+YxJGdmJmvCaefMYjdl0zgJZivJ4bUcy5EcKRMQB5
OSD6OI2nYrzfe/aynidi8q6upDn/YJcmB87CwfLwlkZXxR+Wqpdwohj+FSKrK3eu
T+ITPTfClRjd4GUF/Yz5IWsTRuxLAnmHBa9NESS2wBZnceYVO1AqL4rdoS5XhrG7
bM4pcLgH+N35bZvhMs3+VPKpuFCgfrQVS7oK7ZNsiLg+4ZtIAMOFFDztjHcbjhvz
x5RevsfQITX6+P+1FwTOCZRI8qGikvA3VctLiAWSF/HmaOF2pWn9LPHJGiHWlCA+
PDM7EiF9w/ctZNDjuTPZYwO+kIgYj5Pt6U0k6t8rH4ifwWoQ46/Tzzcy9jo0NnVl
riFoxlXNPh2w6btm2TU/QHUdtD86luB6l7At8+D4Sv+mAwctKAHFUQTd8XgsvjBH
4winUAq/+EAGV1Dfcg3n3EHmcKca6WNGL/NGoDIm7GifYc3alBI3/HLHQ7UvBTVg
t9yPj45eGCwMM52JfHI7XkZ0tmlkrpQmIOdISvOwzc6JZgqCWpwxqV3SYuX8WoXZ
NQ2mAztrvXW6nCttFX+urT/P3/RU+lNSqRVhURBUIDLjVHDUdhmY93KIMibq88aZ
/D4rh1CPXLibZOFJK8F6Cf861MwbA3TEkKipHnHinJmDfMlUQeua4oCQ+ifSpI0p
krHH5LoCbb4TmD0/dDTWGhtojrn+PrOHnK1DKDV2eugQYpKc3FaUc8JRGYjbHXfZ
7lVx4bBYTsmRiAmE5RjXDVkq0QdVkfSw/llmliLsUZASo9VgD/aHBuZ58OZAe9tw
IM76nNdd28ydctzNgs5xJ9qYVAk2NtuHC05aA0IiPkkppe9z513oX2YjorXLH5e5
2bLUcKCdzCeH2wXfCDKWx7rQTq0wf9qoW028e2rWduf//P6R8eM1rIuEzINoPgxL
xHDWyaPCkjCO54LDiI7dcD4JJeHKLrARZ9B35Ns/t3IU4YjZtprhZD0wp1HWD6jx
aAU5dVZiYsN+sY4oftd2ieoZMFN9y+QyH+q3eWyPfbSEkXKgcCJSADiSn/qALg/0
dAezFKuxyN2KfacQ8cro5Nv0ZfyxH4FqKuYxVLh9f/p1BSylyvk33RF+eDZCsxb5
dmoWwa3Dch/IKv5GV1hf/xbeJsrfjjq5wU1llFThAt/Z9nm5zZaMVU6ZjiiV1qkl
ymekWIYroGyjF7EioKMokrpYJIOQi+cWTmAfTLJmHXTitMaZutdngGt4tR/Pp8Mq
C2Yld3clekxHFz8j3rWr93RlpZO4EtYGGrXkMKrMs+Jvnop/dg4AjL/sL2RjoJhh
1RyoZ8Pzuzjf7FoWNDxf/UGLauwI8RJ3plNz1OKOyEMm1cSvQMGRpU5OkBR7TrIL
1glb0zYRLB/8g4sepEte0/eBueUbzgZ+jmllT6J+wbkgI1cL3CjqJWswI5bmN4lL
h8eaLQ/7mpAGJUaQaiCv9LSP7flMSI1LYiydp0mhBMdnIFNS3PXPFJBRrEKB7t/0
/8QejLvWd0dVMaLaTAeRtsnYuEQNCrgVw5SIePfr8ZDqvfYesC2OsS+iEdXdMNkG
5n1FPFeSgHEGbWfErFoH+l1OL8arRjUjnu6dOR6SizqIGQutZ5zJjOLSHHcr3t/C
WkGDIWauPyz8GF9P+geOdJOe+aIFPCFd4Cix8CRVtpSUl3BpYM/KYjriP6V1y17Y
PO3Z2G0A7HegtYfEiWSOnqP5d1NMBvR8CQT0cENWdorak9D8C0j1oklHR2gzVJyA
WkGC67mXAWWZOLbVTDPzoEhkFk2ERbOlUn02mWKwJwTDEXRaZeKxPeAmlvbA8lj1
qi+hCkosmQP5h4T6U79gTDUs5o+4vxwKgzswgFX2kgTLr33IdeWDBDhK3UaCSzPp
h1KztNROAjP5gh5Z05oQf9dmxGS9MP5rJewts4y0UeUKv1Hstjid3TjHML3z6oQ7
T83NvjlAeenki7GPOcKp5rYIzAbjP6vhusRGymG34vYQ9yaLkleRfl05M26Tif1+
xl73NI02uT5Ihky+Sx1xoEMAhMedCNTD4Vmz+j+AHlh+LvNnRoNWkuG9Lw41VVnL
O33v2nlkal0hY7yeVaT7e8PhBXi5G4k+KKx9M1nHHJfhS98+wFXosL2oRmntsy1/
DXeH5TC4QxarKCaISpWkkFrG51kX6hh5RJUEexonAW9zboJQaeUwdgNh8N1keleP
tGKAApR9uTjhrqZnJ63KrH1lxb0p17wTkH47incdmlbV/Lqm4DfeOzgC0FG7KpxQ
33TGGN8qxAst9AgxaoteQHv3+Mj1XIqpKn7BODIDMZ3oP1WIPyL2Je3bIBiyJR+5
O7bulpBK5ZrV005ddivJJuRBx/ajphOvXUKbyhfBqv9C3d/xccCiwTwMT4hORoNO
5eMZDOepMBUXrQEbx5tiGskhORTLX1LYKqbd27O3EI8f6QCJWs52+wVS38Z6+8Ky
WIcraqGeusXiKay+pg4W8pbjSDufZYQwIVthZFVTfJuZ4UkawSnZZH0gALWMcAKF
CRBgJBoc30GaSXceZrE0AZ2Vyn37R4q/6RCPbXHD9kk/AMeCtk4NJi1E2hkkTlxK
+bpotkWq9MSHwD0lYfY3UVtaGFivGSE+cOUeeWLlnm9wt5Vic526hnj8C9xIpCdV
AxusgHZzn162hj7SBpFDQA3xIECPPeqr9/BTf7kIiCvzfxgA/ocR+MI9PkhBOx6V
K8q57x0yP7U4kbdTFkGwm38oRAj7bHQo/PeQ4dJgIcTSMIp/Mg+PaSLXKDkmCY1B
kMkkxnerT0bCDZZq8Pu4rTlrqlkQANIeAF91Rz3ua82ALeN/jCOjQKS4cckzheVG
vadqesOPA05/azQeasTrGFykTq1V3GEmjGRDcuYKUlHt5XjKbRvN9amrqBwBctub
UvfpaytN02EGLAmtkd2aVjnPEIAKtd+tonlAkzWBRQToxgYsbmytctd2Pry5VOn7
NTYNNgrNLdJi4vDOj+JvU+IYAQ+tPLpEjTnnTLYmeqyWylvmb4TknquYcjC0Ytxv
fT6KSQ6gWsXOrL/IXn4I/opDFbPQVVJvlvmaoAhgOQBOg7LLJm9y/RgyGOpzEEEC
ghHzCTMaHkBkl3r9VjLdx38gLQ/+vbP2Glvl5LG7Nd/r7rFIrVONQPW/pbVUjXdh
X2XCi5BsWqt/fH6HI33UD/yrrAjtWeJq37QhmO9RkGB7qwTaYu7mALoIGQ9qEkAP
zsN0BS4kCavpFzT2BvZ41o6g0vh05Eo6TVlcxoTvy6gY6uTaCuckvXMc8/pYB9fb
cqYbI3y/9jDalA3xvncGjvaVy9vLO11SfjlIxXv8SANE+86Z7GS/aiZ8u0PGNt85
vXajxjFIXZAck0s5CSjF8vOiAwy5enxJGixpYj5RU/FD9ad3pNcn0TpwtydDJViN
6Ots4HpJcxXkEgs43PVUc83d2fDtJP13XbI95tYiHIr3dQg5NVL13W043ZNYFCVC
fzn9t/FeRpzYO+tGLbQGc5QKS9YUzZIYBYzLjz9qBIWdTfCPFHyiF7kqR7FiNNJr
kgLNE/znwzDP8SGDuZTJ6NYJJu0bfzQdX6pkvvFCrfeY51Dgx4vGj/Wo2oocBzrn
BWDS+pGPmMnax6grdg6cWo8M+3AGoACpzvzhkem1C5NOnpZ1LgoEvWq9VwYgsQNq
Upo6a5r4cmgx3sLyWw+K5oc0D572vK/XvcYFwgmkKzQ+TMZy1WWCaAu07eRoKtDM
OoeHWFCu076iVzPP5OHIgv4jHk0TU/kFImkJjdHnV5+p2XktgNq3+VTpfWetJWsG
y+qESmUo6mjHYq92SMG4pFvcQB4DwmTcOOScXstFYO+Z1TxVGav/7jCC/ADna8Ka
E/tJGqKR4bG3q5YPmkWVQvjt8qz+LeF1SgRHMum/4hKrv2bm7zcPH0+Hght+V+5D
Oq6OqeA1lW2JyWdX5GPWCvgnOvFWhF6f0B4f45pGi/JZW7wMgGj2Zr8fp3sX5+Qo
zCnG2YvMHFdTPDBeoQTfAeqrqevlg0FtJZreU+jt5NjiEnHo609rO2Ehj5pDAhrM
A/qcV+2901vZyklSF3VvpUJqn7afh9ZWWT/wUu669Nkm1Rh2uC+5BKlAGaNZld+B
N4Rg5MUSy5Q67xe9yrSy+/IXLS/IVoAx7xhYeef45iaVokVxJM8YdOuEaobQusMv
+Sia1wm9t4LKNAObkz175mDw+qiPQTM97L+xiUdBP+HQry7kK0f0p48TE1bEx/8F
i2IXOaFEfO5yPxNeXzd1V9CeK1V8ChiXYLyoDHAoN85sfCMfdHfrKZg9AXWB3DMe
ckig+oKUhasFTnAzXJ+eRZs/P8zIGb1e6i4CKJPWKSwfJ1O1C6PJiQfYWoddi8It
M6Aw79ApdPvK5lUlceYskVRyeKCCI/AlTjl3B1+FxSC4gwhTksJsgSCshymuRRiz
sanBQ8f6wGom/Llu471jT+mIiMgHE9HzrR4IQ52FIwZ9w1jQRv/wmv23ZL+B+J4+
yFqVz559SwKkRMedIy0zjCjR6F2Vxc2grh11q+WYOM2WeHf84HOsfddTvq+1Km49
CUw168T75XfIyjOGium7F7hZ24mKEAExLjYTqCjeKB+2DkZKdQnwSrcHLUw777fB
`protect END_PROTECTED
