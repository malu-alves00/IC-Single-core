`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Qtcb3Rct6Ca5MRl7ZLHNoyl89/8bNHweMo6sFarlOGUD0i+gx1dBoJQ7zOyyR687
MQAcmASFrASmpDyFQpw66zrGts2a++xTJnvj0h9v0P9dmZRtG7eK3WXwo7S9WNo1
mInH1d5/7X1QJ2VigJZWYe9CYqn7AXap6vZqOmyrmiJqD4l6inUVgGRHUybI1CmM
lm/8D4Vl0J5Gk04XyWgHDHh3JG5HSGKVw027mBY1tpBivelmIR/dSTzi9tsr6N5T
JtLw2A4y4NOmnehOP/4jNqlLKJKtG9E1Ae7YvClhbPSsgjR1j1DLsppqD5Eajq1D
5Ztn8+4OoaL+AKinHurXIGmt22vUWKoPIMYE5u/u2rImWXmfcBF8ZYldW5Pc6e/c
YI/CWxsk7pXZbzjX9lewdp16wiXkNfVE2/dguTPd0t9V2zv9PsPtbuOuKmnj9llF
9LYyIaJjKOqbQwxAn2rFl40fyccwhTupKY4DQwxAW6cbQ7CvCe35GX2tQohJ4gMf
xuVF3WhevoIYy6Rm/V7E1vJXI82XcTg5ZWs1212a2r1kk1x1Q4D00ItX1ea//29W
6fEwkOWXwdVuMN2sw7fkUM6ETWYGPQKw60ppzvxhsCVn+BuvArzXtnOjXFGoSkmw
gR4MTHKIsZGUGe/X4+/R+ZLRSacF9BkbfRvuB047iqgrXkxBu5ATGu/Lpspjhe5v
Dbvt4R8pMBiC2hGSfly+l2SjBjSz2szpxzOPsXGyrpflvsCaKhYBfrmpU2JNmVuy
4RBsZUf5f436SQn1ekTs72BIO8Pg2XZYMSKK2R9jbJ+QRjjcchq/oe4lrH2993uk
pNM+SLo2Mt9PfSDv5vngwhlUYe7f8zOMFJC3+wmW50/UQNUPD6vVbVjw5aGd8ebr
9UFPkDcawWiKRP4MC7kBkXoGFAnIF1lQbfZrxlvLwd70TCM4lMLGYThxqCvsxIkL
xfhKIPqrUONHzV8sDTsDTGTzxyfL5PVbtdVio1vcJJUgTMoqT2lnXnSv/doIwnnp
MrqTD2mi3MJ4O7qE8z++nd2scsl1DMGZwHolV1dt7T/tq48yIDzgQag1ITjOkC86
GL6bQb+lTfID3CxWl3+1GSkD6LM9ZsWEqY5DdYCkRRlh7zS20dAJ1LqVKJBOu00w
xMMnLMkndjk3YnvgocPq2IOupKp6R+5/9vRH0U5kR+p9nkmGGw6VSPuioc9Gse/H
7LbHmhJhJI9R0gfyHYNqhbxLVZTZB4hboA2s17t6CK5bwxWdTYpRAegSWCF87/7p
rN1ZXWbph9cGce5KeaIKc6FMOCuHvY39Pwl5IEKZi/2/AGv29PQesj7fCIcNrdzp
UVyfTTaMm4H3T+mAMGM4fvQUQ/aMlQB+CMdVMazMrOK8oJIkzOIDpiuqRcX6AcEl
dpjMRMdNlp6jGGhq+1geWQF+qesYsC7SqAo/OdREIKrj6nEBLlWX3xaDtVq1yDmA
fnoJI8en5V6DK1zBtj/MJHRWoHbjCP7uoVnGWmMrJMVN6p2QBW5UcuRWLYIuk7GL
viuDl3StFvvV1wBvf8r7mFwv2Va6YUe84wOnOcu5vn8+9o6SzABBE++BOnVFWlTY
JnlJ+gM5ATaqkIrS6DBMeE50EE3LcegLaBgnOQqRd30GzM2oZPp++rWuHf97xb9j
2y/MZDDWNoSaRMRAwmOx9r0Ftbm4r6XiZJgtQQk1+hu/FGTMml8dnozzMq0/amuz
bzr3+JlUyERZ2cQcHj1bMST1sbqLELAwQ6Ps/i8mG1+nLP57A7BL4Hi1liSIWhvK
UBVErewFVZwbmctohh7MAYT4qS31HQ9FnRnin9XzJWHZix6xevAA0O9PNoPUiBcb
shXojbnkjKdK5GFNbt9mlOZrdbzjZflkCYUF2utLMxfujkjpzARPrYVOrIomaM6r
Wd1OFDPmvHkjInYw3mwJk77XWCFRxGcna6XIYB5oOytnEY/yOrliuhm+xNzVImBq
MwxcriYVbliV+YUUNJOHyIsqwJKexv+wjbpP60YCO/dPWs7oBRJX3xLPCVEqyDAr
tK4rnNkeq3OLAoaR7zcp4YIlp1gyyAGeG/hPg0yB96LT+HU5WDMrS8uVTjyVEI9o
ElWB4XuuxQUR9tW4o/l/gSQmXwUbEtIrBxFXsmIL1DT+30wL1YFKU9q44/L7msmS
3v7Hb2UGDNHq4//BtB/sNA+9ufhQEXaIkIzdnYXpgJ7swzlY3a9p0/KgXgBDIdH5
G2LBdMNeZNwY9pkQCdZp95cfWTY8j7oJVjYI9u0NcGCbfq5p+r/5uBnh5N2j6DkH
zcYVgp6fb8uIwSMdTLHMm/gdExk7y30TYgh2oj9n3uz1lmF6z4/BfX31RIpEX2cl
7BiuSV4yQbinxofHN9E1sBRB1XFBRE5sDjGQ3d8K8gsIcQu769Iwl5LCLzq6dPTF
i4Wd1lM9MESzMsc2K5EYIdE1znwVTu8P4KlsMy6fHDlObT1hGNMwqQZJ3ntl7HXC
t8GKA9nBbF5IrDMJeshu+y3JqZFSuIovT8a1jr0/dNTFGB1AMb9D6wgYjGGKzsKq
ONuvtl01wyIgC75uV83LZUA1qSaiS50LcHSIJdTx2GaI24IuuZ+c4xbs2jMrf7Nq
e9ORaXuAIMXtfeDFsj1lUYp41AYmZV5eahClTCQpP4vGWQ5BqE8a4jEYQvyFezzr
sPo5v6DZTBgFBisV4PZWiWlUNUC1/ZWY5m8CcI2pB5H4MdyeSE1E3HkfX3o6a8gi
vaV+KkO+sjbR6LjnjIPrvbQuVZqmdaXgz8V5Tm1b7ROtMMrUQnE9Ysk4hltxGJGV
2bxdMFeRmbV5fRT1TyAlsfShVJluGtNiiVX6Ky2Aw1Lily5bULe+UPOjXed9vwEd
+93BOyGMfNsFqpukxdVZ2whBEkTswBGMrmYa6tCOwBGxnG3oXq+O+uhouLkpI+M/
zucP8wDJZl4yYkr37RFLRvw2OR+HawsOsdNS2p6Iz2LqZRoSDqUo7IeL4wl2n56t
u/lE7KisxAgGCgVHIAB9wSte2yvGpMncD6Niu8Ug3qEOEaRwRD5VVi8oyqU9YVD+
6Z+i3cyc7lusBPxbRgSMH9qYK83DmtuPGECt5tx7urPNne00jP3MTgf7pqLTC42p
7UhTrEW93iaIWLtjMk+e2ARAlC30KgJMRTMizkFIL0byGSBI7JBOvliEjMWyozd9
laRM51lbNdnFwGlRHImtKqt5JGE2ELCiHiptIOPd8BBTb9fCZVlKE1VW4Ly5+r1e
nwiDXDC2I7rCGHFSUhK0a/a5g+MrIXP6Yvxfc8iFjRZywpCpTZVGStcucoUr15TJ
pwFcDM+vxzJ50UE6OZTpwwm9ytgPqCHJeinJ+OOzZ4M7RDDCnV7rF0nc8bgdt4Vq
CtYHLecrqh7Q8/mrgqni2nO2mFSME1ynF0aYHCaCzxT2tvXHd2mXDRJvCMbmhLRU
SZOD2t9nNkVWnYEuhXZYLVZEe6s61uO7MTpyZ21aSIc5qsx6+4ZvNsW7F/B4K5Ya
hdrPKAsBOL5kjuxg9s9ajf99IpKXp/a6qCMSmzi0QI9uXV1tQ0WgnJaBv0zL+zCN
ts0+qlt0KRmQQWJZCMGOMl3RgQqgkfqbAX/GX8jYi5nQzL1lmVxvRjcfx/nAO61J
9whwjm1KANX4M8wep0o/hke2BHDilmLTp8ndez561Is5VPUnlTR/aA/lB8jzAqKO
3qC9RUykZV/u0Yq4I63r/aH8C5PfVvBDUsUXqx0KdU/TrAPQWnZlbaNI4p2DOwdm
izCDKCFQxeErpJ8v6UWV1GhJQ8xlHV1PBVfa8Ypmm3QIwtDhAHF6t+ve+dedRQOR
pEz/3q74LT4vUJVS9rqEjL/q85Dv6lXIy3MYkDM3qI5rE0qjlV8bPJZJL7d2kcjb
mYpJByExIB0SatZG/bSukp+rvpnh7bfN3o5iud88/GtRUADjPWZYCWpI1suRKftF
nfxMJkDl5hLyOclhE1QYbJCDH41oeerJroJTKrolXB2qk+uONqR5gtaz07REr+4S
W9KPa2Iue4uuTj2VaphHQXC3vOa4FxKznS1C/eIqoVeQqLpMUzXRUGRJsdQOqavY
F3Je6Y+3oxCdD8MwIegiyeTWu5ShZfAB4KEGkCSn0fJnH4eGoOW00ZEpChbktDS3
qO37Hi9Qfx1q1Ht4qWUJRdqtO0fIIqs5bGwcL5ahN4kmXCL3HP8147RMArpjJssM
Ezhbsi5Cza4c9sCv2aTjc0fWHEPbDHoPqNnZHPrcTp0=
`protect END_PROTECTED
