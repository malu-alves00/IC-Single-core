`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EaPGY9ALdDYSomhsKZpYdBb4PRRdKTt8bK1QUWZXdAuVnRJ74V60r1Ea7WX+mKyB
9SvIzC8NSIdEgZY1PAexgvTLXIYvkvkTssKB27ae5AHMywKCgoLe7aLzQUN/RMxg
zDDHnj5hILywprg5Qdat5zOeAr2/PXqKRh/eU9VOjGJpjBEMUnU7KtWe4ymB88e0
s5+uHLTxQC0OVz6U9k1KT5ZWDrgeKu+Meg9D3VuVM5fn3x9PDxfvcn8l6sFtgKHz
E99jBFgMH3NBBRrderv84G+ckUpDQwD07OFDBUAhFtcTwxB4t8kVKYqjaHWJpkQL
RmW70F2tBA/qfQsUb6QOUjiK2/yBZN/7mjsf72hwy2oKjhXW3ZphngseBV7XLrw6
yUMt7eohJfLjpHe5Z7wo5BisNGrPY0WwRZB3j5XFR8rm0ZXl1ZGIGLic7LW8EFl2
tb2UuVi7XMegZG1dpzOj5Q==
`protect END_PROTECTED
