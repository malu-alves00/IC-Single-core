`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rcjOWZnAN1lrD33hBnbLMyVEPc8+60t5foCNtIRYFx4nxvMSo7izHVA4xqw4ZDrT
h+NkkLh/xb0KD+YRKzbbDYaJ4zoa0VtWRs1Vfbn/9kEk4pHhSmXap6k9nUfpyPY0
85IkcGm/qYItg2mSU2TNyhqePX/F5cqa7W4C4/dWH8uBlsShiO4DwPe9bG000G1V
lNi1vSJBkWW6Xn+qbxojN9ypcJhNQtqPfbBR/dH15Ox3FyMoKmHLqHN39GfJYhiK
+3A3mEjUh6XtKfSZAdIYKmsKjk4Tfh0vR6irdrAkvaQGSuYbeXIGuNkFCmaWNZVt
HtcD5nzRGKCA7UVsRDO0ihhoSJ8Li5MiZrDVDrklQWTfURJcJuDi1j3J8oatpIvU
ZQSu9ROSx8jhWIf8TSXaTHVJ6eaL7jfoDjLwIF5ajxzaWiz1OAblpREvLXLKOkL8
Y8yp/ORf8xp43/TlIN/lfj6rR0ZF8FIMX4FN34TqRBMd1KWifSNxNEK7+CJnijP1
Ed1ZTBDEHj2XVpCzMePwv+dCoFvajKa/1VdqcCE0ngJUg2rzp8eubrBkgPGwSQlO
qJ+yOEUkXMqDy9zLfYwbRMb9PuemenIs+KohRFjxDGWcyJ4SkwGr7WW7Uo7UYmbO
GcImOs6hsw93AG8NpPb485JYI28mbKq0CdTe8D5uHWmrCRkj+JCqgwv8o4DRqk+E
jjCBoFrCkkMqLSgKDlZWp7TNo0x4no31r83zDrLMTAV2hjtt+gh7BcaK8OZaMK2S
QuJ63i6Ui0I394C8Ki1p5T3AaIwSP3ww/yRvDRaUQW8rAha4k70jFnp90ibkkow1
VIYwmcYrD0V3LgRk1hvrxA==
`protect END_PROTECTED
