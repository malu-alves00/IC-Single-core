`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
S+KKYK1SxUM7cEi1qivfyUuj1ZaIQID2A+zaJXuAtHvBHqsCB/5aPKXqSc8feFa1
IFECJ/lYEGU4MiaTG70hqAf791PF8U+7rBm1NdrXwngA6wI/fv6qQchs2c+XLw24
AswBnMYpvHnRnaMhM7YUeXPckDRTzHowZmxLmT0QxJuexd91olP0Wm1juNvLOrhW
v6GIbhAnhuKZtIi6j42GOM3pGTohvJ6XxCykJjCmmFUQvbKIORsjMzd/wFz6BQPB
b6Z703s9rVB4BpkZMrJ3QLpKqlJY3y5/ca5M2q3AI8r9ywtQe66iCFI9u1q56aJJ
Tawv7EVdspjW0d/MIqBsf2Mygpesup1vNZ4A5xlqXR/fJM0M8HtXPXd/0mf/QC3P
ODUyvCS5YuZ5qmTcCNAy2gVZfGNvAeTp02D/Cnl4S3dRrL2TfB/o9lEIy1wXyMv+
HVPc3qMbdtaTnSkaCzj0OaFpLmjPryy/X0Dnare3Ws8aNJZ6tCmpYp7bDdsMP9s/
gg2ZWNgqHmd9p5NxOXw2ziO4jA7wPfgtIiakXB2L5tNbJvW5BDwxdEvlad3I9vOo
a4t3oEbH3joKtFsZtXIfeJmDCKNN+oXM/vDEAanXRWOAd0cUaQZ2gRVN2f3w8aSe
gzIzk0neIhwA2EnyQYpTTekPkHqQ9C09khwf5Uzzkfwm7cPiSKKQHmrLVBTeA7uq
IwPu9c3hZop1xBLkkOmupl7Pnx4ejTt0HK1885Fvjj0y/wceXr4+C/BXC+mBDkbD
2I1n/+e6gOSiV/c6aim4NsspVX3y+BV1Ebu0K/uaiIe202RAlh+k/ZlJmT7nZ67n
OjjqlT9fcznJ0M/QFDBqOfMuyNP6kOUMgQfrUO9xLfCaC0VKBKzgH+U0w/eu0FJc
InUPBUgE8cjq3XYxSz7uTgQ1xKOGkRBUwcdWPTI5aXKbFUnfvrRv2CoYj8FxHIf7
DxzT2UAhlJ5YKq/fBQkb/aBpSW8BMtw+ztJQ2i0K2WQl1t6t60rYPmrOmCo708AN
1xodyebLt/GtBtwwMhvpuXCMGjR9znjSN52qsPRfpz+fYz6pQHySyjIdAGTNLMpY
8eUvXHAYKgZIoUHeltiiHqZs/4v+AxupNtYVPJYClVPhAjrse1O973zrPKY+Zhca
+DjtJy7wWSf+FHr0xJCa3BKa5gvEsqAV3NlZ16ssgg2j85XF6nYX5xPmpN9A8N6D
SFStzVcWgi8NcSW6HOKa8cO9PPAEsCeroqKw3jVNOvu43ouJnn24SV7y7CreCSYs
owm955fjtrvkNeqVPBj2zhNgzrRipjRuOUlPDDWPyIFjt0BN/GuiTeLq0h1+cCex
uusa0/IV4pZC7sZNKdiL+avOsFIhNxb/qPl8vszpmwtfmuCREnS1nX/adrheUx+J
ZiwXr0r4kF4JI8Mkq4kx7/dtLMJ2WkwP+wCl/Fgr4dnBQVmzm7foAJ/c5yD98AhO
4vBSkxTE++wKxqI1F6zTMzBnQglEfR4NvNi+vN3JWEpG+VUwhWD6ksN7X/dZOCJz
a70of22qTmaHKTIgVgLcACLs92f3WcYdTObxkSBIx1QXcRadEON1F9cOUkgrTI38
GCDvgaqOU6X/yXJ1oec7piRABjBj8gxHC6FD/GPKn0v6JsYrqmWGUe/B/odR0KPr
VOtTifJr2NOxsRk4rZTNeDgXrcCoZJkF65+L6DDlQWIuajpkbQgOMoclkAoAV8WB
zr3Z9VO79A2hAdTAeJKHAlGoPy+uG+79RFkqRahM7rkdOOnEdtUsKv3vPumSlnC+
z4QOKRIyy2q3e/QTaIIq+4u84gtOEwtlFdptg6h18lVjdaQYXANZYgoz9IqxXGbp
HEVvvCUoMZ0oZsiHG1eIzjnkNiq6ZURuDS671zsI+KA3zkqDxTjBnx7SqwvRBwcz
SyBiULcflifcR96qjsdRS89V2r2IhJO9bWHG+4ywCweFy5j+rPKGYdMe5DiwHzG3
E7gF00H3FSTt+chxfsKamlzjHi2nwbW5lETampwga1MnjasRg1mOb/rubTCaz7H9
xkFBJp6tfhO0j+BNTa96Bd2hjAOw9bUMm/D2xJO5+eYlNVoxQoOHoqq/tkg92vcX
rRnYxmTvxPi9vOFTiFQfJ1xpH4rkUQssaG9y68hoIuKp4ofMEPbIJtbOxBJLLt0K
+cnCtmCWU+hZwteCVY2blKgEtCgmtmOqcr+qBWWTQkxd54rVgCmJCyjGQCe+AtT0
P7Lywh8gYUVRzHIzS/h9q1f/myUdJak+cPaZw3Dx3VafM6LEbganYA5D0nQe9bUV
creiWvGuQIE82uLxcImgIYkkMxXKtSS4WJaHlaY+wmiXLRCYicbrfex52DmshzN5
fEiZx4QgHtYvCxrW9P/x2AUkOvvDAU78VfW7ZKxltAnJy7FLJGbfs3Zok0tJ4kW6
3MQ9kq+U1KrImIkTeU8nCHjG35IdmPaVSck8AOQcOIkWFARdBUAQIWFFH7z5KdtX
GvviuCpjnP7mvh8sftL6baqCdsOux1zXZNR/cAFk3XEkpMjOLLFhATDBXmWeU2E0
Yn45HGGz/LBQU2EZyLGWfpoVXQxyQ70+4HfuF/cjOxkV+0q3yFmgO67V4x/AFqRg
y+1j+kLY8D6p2TgOAREuQBZvxpLKtk7Dmtlrs4VtmVIyf3+XRzOH4YNekNoLHmWu
+Qf3wEP+Oa/dVsqWcw6kd/qAq25OhHqE7OALEefubPVzi6wuxrYXorwbAN9K7HYz
y9057Fih/7yCDrbZyFVV9W9BLIJjWIiOPpI3XizYARk4RDVtvyaZ275lNgcHrkTr
hpAwFnq5iHH4EQN+Zqy3k2/g8dv013ROK7OSnKhXGmdbxfOOnE1rlqCPzwafcEuK
3eMmjDa0Hq0MBtzTaKv0m2g2jVxwu2ZcMWgvxDAoOJI+lXrcg7CRJ4d1qVZsgTUL
8xvEa0J7N+RpDBf1+tt1wYrVQwcfH50ETgbNhTRu8jOHODHayOrLMjT6QvgFkV7u
E6EIyXaNeKYuRMgqD0LO1Tg3gvy8Zde5RcjABhSOaM6ReUMDQcxdevBx12QgrYqG
XWb58yOTWLMEbOXbQCPXyK+Nb7W1zvKbJCa/zCyv2KodZIdiaOmbSbV5yMWYokFh
gTv9llSgMgzz9SElag4M+8PzZhgmsH/b7wxPx0s8AczDunZATf0Ap9VDZ4OqvPmG
tnRDU0uPhIx43P1LXZ0vSpqqePluPmUYxR/hgg0sbkyNHOEhwstEgHIEppA6vRXJ
U7SMqJd3lxQftPZYb3RkZcp7ElXd00XTyANpCKaYFJ1mZHzuld+9GWh1x73JOrXX
wmSZWDQ2ffHBjA6uWEibJeLDgb60gV/Y1np2k6CIWxo2aphufpUuOyR5EYG8vekw
k8lRD+u7HgbEgKLrcijFE4tGgNSbQt6JIvIEncx+fNL41J5K3KVN+ONmVWWOO8Sx
06tTR6qPPDlCd4auvfKXVs+ND5AxMuUtOiq1GhE8nx//cSo2oDREGZwZVa34RnWg
o2LBpbRzC0Bx/Jjs/a1Wj8ihm/PrgcPRtxsvALyzCvQk1g5aek0j3vmllLJQI/LZ
MOJo4L+U99pOSm4iM/a3/OAFMkfDr/g3jZgcZmKsTKVN9FZq5JHEN8N+O3rTLWMY
g69jIwe5cjqX6dMGl3/EwWnypOSrZGOfGkkGp86bf/IcfqG5H4Yhb7E1m7Bz2McQ
DuTPhZc0c8XhMH6JyLSvwWSV7Br4Te5cpUIHPZQ5PCJxp7G6qYYtV0zzPqgXOyRP
xCAu/sLNdHyKyHfOR5C99AR/3kTNxdaQ/wfuHAnRJBAN5scCkiUQOvAjlilETFlF
8682nylgV29o75a/ytS7xgrxiJ8rdbZ++Gsy++ELyjXEX15rfMsuFmxI8Lcviaa+
LTEzrigMB3zC7b3C99Rwhu60VF4eDoPecZtfrO+OymKsdilblUg2YE/a/JN1L06e
4hmEmdf7AMqInf3haNM7WG/J5FP+0tPbGyDSLSB6VibnsBoNgdVBKBPYo6HF1UmB
T5EjcjmbNOqb15dfEYRBWvZeX2mgDvJ6gQjbJKF1RQeAkgdiLFaIM0kFnpRI1wXP
grCg3P5Nv/9q4xBMkm/IvdnzVWfQ0bTvWsdEOsPlXP9JeKHiFB84L4eRuNj0x39y
`protect END_PROTECTED
