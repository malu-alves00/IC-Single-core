`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OKE4T0EnaN5TFo8PtTxEaiLi1yl+k77Xd0obf3lThfFFiyCFcHjQxlVBal2uW6M8
D0ZykBt4TlNflo+zaMZoaJ+jRvyHdkhcvyEXmVhpZAJ0eUfHYmuzwsAFr6wj6SZJ
tPfBBpRsLk9LmEHlSjDJF++ESc/zKFBmf9NOPJcBH08rnXMxbFNHSFnzmC8gFuzO
rUvFHgCX3D6z+yMto5HGk+9NMkJC2KwISQ0LiDHlCSw5Q6if2nsRex8YMbF/v0hy
JfloVyMfBfcDEzm3MWwqIJWWBg42RYE0JC/l7lpCGLWog9rm1MdDb8o24UJxRLl6
2HHdeY9L1zDmBPS9+1JRXgMG45TxC3/bv78rjI/YUhjTWBcn78lok/BtTCSZV6fW
HiIIa2beKWBMBIH+Z8jCELNALBrzZ1tjdB8cFYHPUk8SslDQAj19VpO/plAz3BIe
svJnG7foG9evj2SBAz9jH7rMS8/7wCylYexSynBqng/FN76sIFnHxlPEfx0/wRfF
9NvIt621wYanlZHrYiV5ld0meKiHn3xUO728obh10UHff12dV9FyMORs25/UeDB5
JlXp9nlz95g+6ItLOlIXTTqfO8xQYlBD9KoVBCRpShUPU2vAbIIp87vqpcTSoAWx
9cBEKMKgloCx1txUjXHL8eGNTgY46/RnSW4xXESIls8=
`protect END_PROTECTED
