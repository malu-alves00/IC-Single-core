`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
W/FQ5UfFjV5DAM6DwWbAie+6HdNSsd0oCfvu+0Fv6nYxDKE35b7RVs/s9SSCbpfF
DNhn5+GUgvlkZLg4k3JwOm9Cvss8SbbpvUvwWFnVRBD1Zgjw2iqMgGMuLoPdv67v
Ucfgyd/L7ntG0iiGH129NdVKpuBN0gQbA7GvArgkH7Y6f5oGJsJkPgSkGLkZ5TCa
whPljfE6PsZ45MuYXhlTkCB3VbiSq/atu1bRfp0iXYw6EwmNtoUAuBFL4uQ+LrET
bXLzeyiw4TdKjwTMBOAjtu0l5gPor6ZHPK1Vm8B7r9hbpYOluzrSnW1CEEdHGmXK
iKZQ0aEYBssdt58ofNCFGx5J45CyQz62JZMJvAZr2k2YGSQtTi12phVbfUcQlQCm
Q7YK5mb7YXkMy9THAhmaozSMU1b63cP1/yW8axDXUaEuDwtuoh9aCBtz2fs/ggF5
8SvKGDNZN36zIaol2drdUv/qiHAh+qmcdcRyWY0fBcsRILyz1zlxVu9Yxch/rjIv
lVgKLUSXXMOGdB+SaW0AO78WtU3eY76sFQgN4YozaCstw78e4JwsoX8Wwju10qoM
lh4C/lOKgEGjzHRzKR3SWlieJp3ix+F0vxJIbsw3pfFP41Eo/xUEa9VAedZaJM/l
Pmv8e+XXL9VlP79YAX6fzNulO3w8QgqYSwUALT4xBcggJ3f/CaksHPsN/eIdlzC2
CNZFzW2amjHEI14sR6uJxYvlELXeXoW7h52hJYLz9+ml3Ec1CQy0y/Nd0w87732V
ipPuKxIw99zJJZ2SERXc7f5X0l9EgBy1ug34wOzOPgbaaGh9c1cZFtOgbs3qU76P
DIuuQHMzPWlciEWjOwQJwC6ioRF6rcRLxcdN4FGTvdCSvj2r7DbElbArfae1Or8c
yNfShdoyDHGsBvDsj8tKuqDebvAgFXZwxxDk7bAwQUqi4gwpNM4FWIlzyJe+NalZ
9aQJEKF7F6AWlOF72+zBjNUGSojZWkzMuzlP8ntSu1b0m5/iAXoMBHy6uKFWhOfR
lzcMPzkR5/xzMxgP4w+Q/gAecmcTreJOZaPswzmihNp7LR+FZEL2WCbsPV2ory5Q
P/6cbHHuQ/+ue8iO7yAULL/W7zmltGYcAHvGzeiB6MStErfsoPTJZ6l0AR14z1zL
M1OYhmy3CniJHTgln18vCb6bm0yc3wSJ+Kor0ZFZqiFcQrFiR9JoNu+UBu2LSx83
yeAqOIn3iAvsxUb74vI5Vtc9Z73TnSgUKcN7Nv4YvaomgRpbj3PAnprddMKyDpEi
Hjuq0cDnStIr+EOZ6nxxuBrG3+Wno3esmRwq5THE6hv93Hv1J7e1sNRLd2uItGLq
sd0DhPtq/qCQ6myI3RtKIMhrNzyslP5p/wzNTcO92IbABgitaAdEj6Mkj+HcqD90
XEF81YT/IEQkWEca356PxANjOiTDYmUR54QaBK+p4xvPLgBt9XiVtnQDjzFsVBE7
HhnX0kefEobPj1WSUxxaa/D9YrHJZbMOsc0nkpVMffMdM5193aG4B+SCYAPFlKvk
gIV+DonQnYfT1emfQv1JHS92rW990Ht6I0Bx9GliSgI6zdxWOGfx+YniGtG5BkH/
W1T/Analv/YpSQR5ANgSqHpvtAMxemml8j2hy1CrKaopYlkfYiC+qYR51c4YgnTk
CgRms3BgHDQaKFmFap5J0kjD3BlCmu8jqGetCAhs7f8LWPJ0Ca/ZIbgQopiF0ibG
995k79sbYTzVznzoT5ti41K6FHTXEufUptVq5l/7dnNeoiAxEngOZgK6FlOhJrkA
ibzmcnrgPEaSBTeU0oqDpynYUFkGTIdCDzM6dS9DS/PXlgp1MEjOZd6xXOmIDRqQ
Riey1AVKxVCMZUTOQ35D4IsbYxWnd9+3aLWMnN/W59QTTiaa4jSjozMy9OFYK63G
G4wpJgCgKKYMK0iDfC8p31qCmx+O2b26AVd0nZgvPuxAudLdM4OH/CcSPjGaIjCd
WKApukZSwjYjXTJ3MK4ebOJclmtuQXzz63dyswEoukEksP2JFtcgIqWGyq335xSK
7Z5V20vrjlFINe1RIk0DONEUu2Q5G7SWyRmF2oanluCfKR7kNmlE2uLkSyWn9B29
6Bv6k5lzygAv5ZNMdJtZTRlfNLdRA7MxqO5VPgxMc5ZlXE6MsWd19IIAXIkYGnlm
+Go4qqJVs0gH9WFyxvjczbqz0xswNn9ONZcbypJMjasbD4pzldFcvXG3Kp7hEL70
W0rxBpDvH0FFYwp+LQpHI/2XSJJW/trM1BnJ+0N+ymcDO9dUaZCokUR9GkW5ghR2
73v03aagcV9WNQ55DcZTW/CdyeJxJkygB34VkoTRUpr4opI5S31W4kOySOj1If0e
aTHUQGCc6rex6NA2mrDf0zvf7Asyc8T13gjuji359VTUD8SoWFIz5hdE2kiu3zaC
ueymwmPhlPFIFgHV3PGyNhrg3kCJQwOb9HL7BhAVGQxQJInV8HexBzATRTXOhRn7
GPyjhONokTGYzfU4kgRV6eqVKt5uGrDCTDKPbcKKGoM/DpuWAnJscW34xH4UysgX
zY89TuYbXDyBnKTdoJuVC/41mnEKOsuGaxM/GDeug2Wkp/0VI0pyqUR9X4mq6KXm
IJN7g/rVi66N2itCZ5qUCQcjf+WWZIFDLGju+fysp+6Omgq0t6l+mq9t32knZmcJ
+yw57hdgCkp8mMoDJnvZc/ontt2tVlSPft56BveslwSGCo6dBJZIKEdtw+N6bbpd
3srDqAbOc38EChgPoywRwA==
`protect END_PROTECTED
