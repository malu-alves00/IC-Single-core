`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OMfTEXN6+OrEnowat2E5l3HxwEpe/5rCaFMDHGANuuO4qoDiLG2XVjDyP+bexJnZ
d9VFNEXZ63wIcy2p3/o0RwTNeJHMDY28VGhd3PKX1/mexDIxACLgHMZaF1D/yfBG
mWZUEQhxsYVb1PRrPPM4L4TC3Cz1uV188OUu/vPCzzxIPOPt9qFiIfKcCdA1AC9M
32mxoLQT9ecba2jpvV0HjxURGISsbBDbPRAIy8k5netz8WNDh02O44bIMt+gI7Uw
bjjojbmgyaJbSeSgohaAazgmv+fIbdZMNHYnAsmHqxrVX4CNu7LVV/pqMHXlskUk
M7ZwRsOMhaPUv4QOW9iLU1RwpAgeG3z2s8r8phCZ71WS5UJdVbkL4+EbPRzAsWrH
uhW4wZ/5ZloD4oGfENLgH/0pwLorG811FVrEEuUacOIbGJFG29j/KB3c3sbxCuRH
GZanfY2vTXDTBpWqYzsXx+1cSx6BbE0bww4VjnglAE2Lp4TAPaJq6Y8EXUZrut7y
Y0rdNoebkPA3GXf4Nier8FioUtVZGmU22SdrkVrjS9/H9mrVgf9wFP/awd8py4rC
njCbTYDWmDBUutrggRDorsH41l3csRXEWDIQFXfas5PS1pTCygQIGe4a4O53rwwN
k2nfhj3Xyre+gT3XVdUoe2bqoER4HZbpp5xQhEQho+SbLuwOSD+hHstj09RLzpy+
g6cdpAKqEdS3NTY8l5zGBrq5JSkYe3ExXuwEWosTtYnhf8wPztjc+KfLSQihMs+b
96aeZHsSrJO4Za7P/ipInE+iehnjdKuG50hRYQrf4CZLE2ACFzv6vTJdLOsLq7CT
JeHv7la0FY5JANLSo/L00CxsucWP28wF+u2gia2bl4QvA1boRHRty/dlRN5Js382
zMGakCjx/9RNHqrHDXYkWbL6MetgLhOFdcrSdo+cwh4zfqW+xSli6QIjiY8vNr33
aLCax/Xfp8gp5SNVKh80UE6zybqBbqgqozKrstmzJ3R0VnVHRnQIHgVD55vGdW8X
ez2DToahXHxITHm7ad7oz5yleYDynSncdXJje0tnLlyHZhz3t3nTmo6Td1y709AV
sTOXpATSMF7sQg5gZEh50Mt9PPAaLd61JHmP9SYXlG7azVCpPnOC6/LbMZcDtigQ
MV0VwMtmo1UV0UpcMf8z/hrVCmAkAjh8DYY3/vH0lGkkBz7VjfBdoM1OKzJ4LFW1
+ESseoZYiQw41DmSwU1qTgGTasg9KLLaSUxc6JYBtHJ4JSw2Y432e6momsukT2tA
pMZ4VldHn84x/bVTmBJYdQ==
`protect END_PROTECTED
