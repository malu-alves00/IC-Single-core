`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
u5zj0E10WpVHssyxJCM2/O3ILCAveXnamRB4JfGyGExtQI2h1j3uPzHVdQu4lnHJ
BXwGwqeQrhQX33uEMGg0cqUJGHwzZ1VW76Evzkn4tVSyjCYgUJWOvaXZzmt1iNgO
fXLVZ1DDDfohBnUr5cabISdPkQzB0c/Qye5MQWMJ0NDl6WWWv6phYIoL5uZL0nHH
ilVVL55+fDMrclCZ19mnJc/6XwF0nUTEYGJLMO/AgZNFeNTvq0KdYBCLTNy2Y9GD
n0ObnlAZIopdkTgYU8vtstrQZYSvTouY8B5WfcmuSfCHeG2mjRA4KBjz12OeQDU6
9gnCk1pDS4jMEMowBLE9y5/7wtoe8R2koW2ZftCwKitDVOlFOMT8TkOnJzgoNUrT
wiq0EIeG6e0GUX/hCzJG6UYQrrXg+mrBcAKG5PUZHj1cbV/Yc8yagJTb0w2RMnaN
p7QQDKbNxSWOMWoiUuWO3wDPUjwgzCcsvZj05Pqz3uzvjLChV5zcnauBZlmzaKxL
UK6UeoVu0wozDAK9rJn9OkhJuPuK26/gigfQ21uDer+CTjSfNntksixCTd0EHjSQ
3gLc06LMpOrhdiQM0wuS2Hq2dtfHJHLhZ0qy9RqtvtM3Ir0I7DUn9+uR1FcYo73B
sxInXr7qSSZmhFTdTkh32kWFOEqNQuOFVMzszp7idOOlNE8JH9BE8bCM5nhkaau/
L/+K3G1ErTsogHV09WHUNpZTqgMxFtcFABd98+0KjNdQCAbOVs1zuM2B1a/kgBUa
DR+E0Ogom6DxInR7ngqTHzRt3wxOvyH2HIsGTmG8OUKeh4S9XTFPArgTA3YbFcUL
7ELHNz+3rhADDUbbvpZILZ8tUAcGZ7IS8VeZOT3hvPsL5TXWert/FWSArFsCpuv5
+GtFcT2Z631rrGnubgB75+GAt3gKJZ4h5977VPmQsAcJuHDEdv7HKrqz+65CzysC
`protect END_PROTECTED
