`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0J096WnLzcZNPuFMVc9DYfK5ptRLyNa3WRuML8ljrLMnw50saI1fqSZT/PfNEfV3
Cnb/lqzgz7s/2qsJ3/sezjfqONHMHOG5jITvsiuvIY+WeTfyxLXN3inD+xZ2QPOz
gVLseYmWAu8eimhN4s2GBaYmChJ4neIZolZj2kIFI+8wZiOYQDhISbbIwSEmoB0/
YXSHcPR2XjaWOyGQpO5r5EtWXci6rtE/dQ/wlpMzoP2drONMnHg99ZCyq4vzxhUQ
ASQZrx2w+pXw09e+eZGw/qRoVQ3AUIFuBr7Mi2seCambnH8FNDzai/2pQUZNR4p5
qBxThuJzuoEyylri4NGww1HllKtRxzp8sqXdnTAwoZ9YGYd097KtZlRXF7KuLgP9
4Klok/52VjDoWT2pkYn3ZuBKRZ0OJQwAhkzMrFvkskyWskt329ompX9mMigBRRe1
Ebs5uK2t5QC8rslLz5YujK1A/5GWE11hTyYHABuagLDFA5tT/xv34BiL29E4ULX9
kb+UPVhtcRrkFZZjPaBGIv4X0NTjtXOh3w+T1ENiTzVjS4RMnygCKWZjZ9WJ5XAM
K1aa1Ho0xbCKfxBnXtoq/Sz4YvreRrSO5a0tgQBMccpq74Dm3w5GDtHnsooFY5jZ
83ClIaS7/YtyQ+ISHKJCjqUsC6YlQzZGu+ne3lAaVb3mpYU3zVTxvkBy8UYS664w
ED3RmU48ieJgW2TqNi5UqGMtR04m1pXuVpNOftS92vKi2zX2H33iG6aZf8d/WHxT
FKe7DCJv7gPXfQ629odhcVSb8OkKHjucUpcfnvFOtuGayjT2uTDRi4QGtQGbZ0bG
3Qqh5jexKXrdnb6ZvELJNUX35F8wGKR49CNTWFGOGllCwyzI+ulDMMibLYFLg2dC
NOVG+kDP1N//vsHTV1JT+9QqmV4MNtGYEldmba3F5wpaGROpmDslRZ96DoF3UIlz
M90538DuaMgdBW+3eSPs0tquRNUClHJiaMu+KhKT++xzQ4AR9C2sDu6CI+IMu40q
wP7LEfRzbqhWDJH6fkgc/sdRpmEdnl2PSZ3qPCzaUoxtQP7X56gPQyoRdcJ328rK
XaLWGjubf1UXWl49o1O2S1y4Hq4+FEtDvXwIrlCzTGwWGUi500YoDQyXbtG2S44d
RmSe7H+0owSsQPN2mw6vLnniUgmUgNs5zflSjHQfl0l2QtIAPfKDnIy15l7lQ7T3
dHwhrvXAroNAzOXhhTUiSV8/GiNxHZebtusUrDFpqmHjuMw9c5SHRspbFsJcKH3u
02M1TmsraHNT84QKqPcJEjydpijmqXRXzVWeL9QkiXZozA7k0XGFKaj6mAcB7/SD
lZuIHPtvuObaghVHHVvjp/NvRr+VQCbv7usyMne5gt8CPWYRAod5c3c6H664nygd
EcYzpVENlCA/lOJMnZZC6t8wleKI3Xj0NXuwOVsNFjG5vSYLPMpeNaiGtLisItOk
a7JXuhUv7KB2V12qGLn0F4n/J9KWZ+pLD4v084BpyM9jI/msCQCnYtthleivAcqD
oSjVTwddzOoMQfdHOS3+gvi8+jwzsm2MACO764N9ltS+e0vS/8/K0qWlcqlztAZv
cmhB2sklA9TFKKgYjskU0Q9j+RRKweiMer06EJuFWeQ2FEqdDYtuWpOuUAp/3IG4
gOizz3Wn3sVQWMyaGUTyeylsCPGJPNpTQXzGGezpAat5x/IymaCEYxtZShK6pzvF
e7AyO4VQjHMTZQ7I8UYHfBGcH7lM1i6+NcTJvOn/zZvGA5zmg4NlBcCEuIlkjugN
tgw50va8YPgOzzzM9GDPY4oNdv19Dh8KjLNJIJubdUVDOCJpLpUFebdL5U8BuGj5
XgFtF5xSrxtaxPysBu/66pTlipeEFfXTdBMxvvgaJzNgPSmmXY7HHrzws8TUPonp
j9t5Nd9oylvlBYJnPuLGaYYNd/H/6doHULK8zuU/t3W4OBHUvi8boN5+5WMd5fAj
XSsPrYf70RZ1jkc9ykr3Ah8a7UgOd5m7JxlXdg20oLAvVXjwYjL4OieW/fA4jxbT
wVOqy4GIcLE2uloCI7RQQjLcbaAhQ5Q++IPkpyWWk4lftrvUSwdQt0TsW96PdzPD
0+2vumKRpNm8+v5WeSqHYeXGR9nLEPWHvf5hkFHcrqLouGz2INkP4Jzrmjexhx3Q
CYWVlvl8043XK/caFC3icvb99AkPOHk5vgjfoD9+oyi7d7+neU7OzLSkD/xSIdrJ
/7RNpnirr+lO+W86UtFIVr0Ghey3hLyL2N8Styz+tGx2bgixuamxTRzTF/qjooLt
dfLZcyLc2yKmsK0CKjOxDto5H2nVfkeW3eXLj7a++ckwsylI6bbA3GQjuawnEPnJ
4bM1U0HACi/2XpqgB5t/DF5PjUpUhl+9kjI+p9iykQbezB6fFNySEmRD4Wm5DPFT
Z102bz7v/vQXpp4D2Y8qG89Q0Wj35TxYljLDgQLQN5fqjv3mRaL/TeV6XjYImnOr
VGiOi62u1pzY0yK78+tINOS4SyMH+Ac4+cPoFo3HvOypTYsUvUUlUEuqE0TEo/GE
c2soJK4RASo+j2T76IAAztH3HS3Y/WKETWWXcz65+CNIJAIsVTKK8PMeal5WxWGa
nbPOFEp4a4ZxNM4Jw0dSweR4F7MXZtrhJuQ/v0mM3i0p/ZRv5jvwUkafw4YnhEhD
xD5YWaVIr11nqtDACzylmV56lKqeirezXqOqQGnHCvBS2Z06gT6RKckOQBPX1UT0
1TxwP8PYa2aE4zmXSWOMLqnkj1z1WuWuw1wUdAnv2Ls/YeHYLGvgCJHPZC5yIiZc
UWwTFQ5wRYiXzJ0gVnRuZheUznnTGOb18+Dd/Krw5TwGNBB6gAHWAzDBXeCMfXoT
EhwhhJs1tCTWAWRc3cgEawWvW25au0Zw/pYnrq0YwvHIKI6SYnNPRI0E6S1+zlD+
VEaUG+2AvuCBfyQGbYlJrm9T9lZIKMKfy+q6Fpny46dTsRz++9jcVgutVCUUBW88
qjDr5GuVfZl90w8dujpFWAxguVka4EQQUUl+6PimDImK3KtMW4TXUAQAUmOl2uXP
kFWErj7fdcJzRxNe6A5H1cxKsTOZxMneVxrqj10B6iivV+LtdPgb0IzahMCRKC/q
+9NeGIKpijf2kLkWdDkPGjxeox1beJKuU/9xRkPp+mFLiIimSIWXUOVWxowjwvJY
JwLDCAswpRMWn9r5H7VJFFBU1Xuhs9kZXSvTQCnAvfYZag/CR9qKocQM/s6g0Pz4
MnM2UpEgn0TlwhuTNcfq95v8RPdSBmSyCrxPB5L3i/kk8xlzX0CBjsZEHNLCgu9G
3Sb0eHvlpL5gmR5WPeOmKvJd6XhyIR7+lMr7o+QDn7JX2yrt8B069EOrVP1Eq/Ec
0aOj4eeg6GwIGBHK0j1iIY22umnsIN6x0uTB1aYTWBJJT1fs1Loelv2ylQ02Hu6J
73Ycr8h+kDURSSlezIDhsGyodiEJUTG/kfxXea83HicomU5xtJMgHSRA/BMXOfgl
HmXF+xJu1CFAiQyYtF4ECLzqJFs5v77QjG2QmH/RckxZcSyzNvhJ26dlymBzYOZO
STw1PemGd7q/vRyzOK3jjw911XJMYSRBI2Lyzzld7Sv79Vzs1ntVGXRChqkkEM8E
xXRsKgGfyx5y9qFeBKI4B1AffOnEWHTnkKOOsC+wxQsdsZtbnfyDAy9pWgBhNAtY
70nOoXnbBGb0MCGKDEeiO2kjiOtPvsXi6cQTOGZ3u5bfnVv4nvvv/mwsp78OhRpK
aMybXD73XtloB0zdhirTrB5CB83/Gt2ANfBNmiot0MblU5+37vrF5xPVKe38XcDm
xsNcv34AEGnh200cxjCTPrRPm03E3LV4YVZVUs4FQkaNV7+ARgMU7jn8s+//XjLv
lcBP16Bd84XSla8AWToXww1XfURZdKazcmREChJcZGDe0A7On0mHI4RflsTJnkde
DxD9vwzgBNez546uX1SvjfBC2YmO2Tplw5BAmJK7YQlKLPWoMZYWW2maVhjAuuSE
E8VozupFGFFC6a3xgvepyYpiyjwQoF/RyLgdiY18UjL2eR/oILOuIrZcAZVJZkAv
Q2JTgQE8Gt3YlJprq9MopPP4IYigzBvyYcSM0CiKJk9o8R1wpmf9MbdNVwtXk2tK
0AloVgeW5UFVqTBrg+e66qdLKFLW+mS7eUFW/jYm7OhQhl1zQAcGyY8EnRhmdP2B
onvXXXJHCIxo6T5JN7e0K7xNR1RZ6vIMKy29Vo8+nbJR+IJUJWtpuBw+OhjgTe5R
6jLUsBu1qVDA3Bhd2Lj3ri2NUcUDIJhAdGKgOa4sbyqO4cLUA9EwmrBA87SiUWGo
GSigY8+jQxXfN7uctZMB8jw/gvjFurwHbLhtl6sonFgQLt8HglBKdsi8dwicfumh
KDtd5r8DWWgcP8UT57jpab1S9swxCiW7r/aDGll/faufkJ30r8GGO/zioqBa7I7P
GQ+NeyLfUI8NEZ9PibLBKyagtoM+/wB6pbGbLgJqxj1etBHeC+NT+pFFBhYQmmch
4wTegYENCVxAnBn4SCW8cMD6zAJc9ckU4hZ5+nPqcyh36A4lshmVrBcDIHoouEqB
CKm3Eh8fgn9ISaRzKmDLZOXP/s5J9qL/y9SH9NHCbL99kSrKoyWoU4UOxNSeZbCy
IM7x4psu8b/+LuQeza9/64Daj2oESxDPTa/Fvo0VEjf1Q+/0zJ1om1Zt+hoVgY95
W4n9NzoY9Dgsvep9l6l675BOnvfNwtGRZyKIj5mWHVsEzhiIOBrrUo7sJ51C7z9e
egrjKXXSder6EYPAIrxJJRA0/AxnpX5mIyi9MmoPLevSQP1uObH+Px95AjWUs1Lu
E4Ezw+PTzWrsJxmcypzJVyWYwPYZ0AzOst01ptE1+cNKv07K6uiz/1moFRpTMegU
LWAtXWO0+15n2DBjS0U9i+0MoX6sE3Gaapj+CS9a+pq6Mi0+51exzkdjfEdOmztP
puVBgktPivm45AIHRLNq2SKKMaaR+eRyk/YAf82WOa6OwqomCcKBCXZuUBEIcEGd
UsXoFVZzeLKC/7kUee8z9Qw3BxQ3QhRB7c2kw4LxRlCc3XX9X/DhMrNjo3GAkWKH
aj1u7iHpiY+YI4WPsunJPuQXJ6m5snGrypFWEWSemgaifDMgZ2q08ohdbYs0Z3G0
HBI8KvCUhFt4IsmDBbowSWvfRK+CDlWBhqzOVqPmAbqRDv/lyD+6Nz2s+Dxd/jrE
Ye9gxANoTB0ot1lD695CcZb2/B+x9EE9GBLrxRj1KjOwTulo9dkPdCkvgheQbRsj
cO+p0ea4ZAFx2QSw7YRiUfHG4RQsumrIQQURb71IWMWfAMs9k1Yn/DQQrN22xlRI
GQ+mRZtG7P/FqWfoGQ9LWb6zapJ5o8fGwFMYbxzd0QCHWYXksGDZkKVH2gpY2EkF
RnjrLQI6eTbugSqbPjKSz37BKdSJgcfGjetjoY+AD8ijvq3iVp/2a5eqs6XjTATl
sQQAYz5zWnKj9n6bj2n1jdKGWbX42Jh+pkwSN6KtAQxO9ZE9szbr7J+tBZR/clb0
yvpLpvxpqvxZ2MZoLo2v5QqGWsZEv6AFLBVgV12i5PjkTbg5/Z7iQrEI2xtjwKR1
AoYf2oZXpPRbxcrwxmyQ8d7ZVgJeqh8tVfZlSCdQrt7KhHzp6xelnTkGONH/2o5l
QWd+BES16DITIQB8qmv3E4RIN/ZJMfy8erpX8UH5NAog6Sn9w5pDMDryIvDS4lT/
Z3b4jxSTn9wCm8dhtxcWb9/Xti+YZAqiUJg6JHRClJ6JGbKz063dZbplOs6So5hW
7ER0J1yyK+HmSffMUbQYQgDxj3YAqvUa2e5sxnShMa8o2r1t3rRwZr5tYoVKHt1N
fP97N+JQxDgeMZggXw50rkjmd1hwYoS/WbUw2dWrpmryrAdpSyTGWnP2g44U4pSi
l2XiH5Fz9f/6j/ADvSF+4iyBLrFsmKuhNPoHTjh/A/bgUG6wNTdHJdoUqllQv7If
2FVyClKbBWJQX2vNKeQjTn5nvdqY+d/ynQyI3Jx8VHWoCtRm27/ddegaN0S11vM9
hlumpBPfQH4vwQoilx2+uYrXVweYX61WB3HW1fnFsxg2RCp0wrCxM97Ltp/Xb99+
VT7duE9NB6ZO/CGIDXVT4exQYR3WOo9ZAlK3zp6AuiE94hkrCk+UrHaCEgSuIOWE
ArRLDOnMLmtWHOPCycve2uui6yFuay3zlX0VQv1NiHfF3+LApNbEYvRfbWyfLe85
056vFWF3mP8s5LVvq76+rXLtwsrkuwuEcvGmT4obTvULyMk+hjSfNXhPtoDHqoyZ
YHXkKqkq3MruI176ptlXIBS6AKQ2zwuiUYMZfLn2EGFte8Qjb3L3Ojq+c5s9MrZb
E0t3/4Q5DdRKWiD3udCDhRLp440KjstUWyQkyssHHpTLUly9KzDe/cUtYiDngGBS
jxGDo8iVTAgukythiENu4hwyGfmxCg2oG4l5IZlEjHxJvSnPyhRXhJ7oP4PSnXwq
he0bDwbFHKPkenTj1s+utSWl7BD5vUFIQ8UN5SSux69HgkdLX+D+CJrjIVtCPiYK
ecNA99OOqum1oZlcJFHX+CfWFauzlLD8OL9+vHZRLQsn66BHKyNWU8nsMrfDg7/p
YEdNsHNXu7nhWXoqApE6JcScdPl5EA2OQ+t9gVXxgP3G6mMRZPMqxuqBUM0D22W3
Jcns9Yd/D01RMBOLiISwMh70VaY03UBNtH1MfJyLNgkBJoX4eSVtzG5Su6CmVXSL
PC8L3ddBBBor1i/22iEl4ncyKplyhsYHLBeA/bI0ZKh2HFvU2ES+N/tFcu35x2cn
Y5uKuHq8d4XVJLsa/ZkeGplgKKatFFuenKIGCTFVSh02j8UKWoU7rMewSj1iFnj4
y6P1QYPP/IkHKbSA2US+UOAItBhIz2hSavxB8Fp8Hr5DtE4CeRvRAzPsw6wn5kF5
p1dqrOGXtJJHrSXqQmM896ZHEVcz5vTeOwtHomWrTvYYelfRYQdcOYcn3bLluYz0
AShV+DNxF7zu8qEDA2Mpi3ERcN4kYBEaaXOsKba38NHKVKuQmWBGpaC5J/h6sYCt
5devq4bjJFmjn36x2LbzHDms64HapWwjeiqKuL84lY6O7X0pJyEE9JuptaRvMYNn
U6gMg0ho9gvdUTknPbPoKfpNfac70KK7nYx6P0JR+hXhWLdnxqMnZ346im63jA+g
I/fLH/Jb4OqA9n+u/1Y3krWvRzGCUTNNrrbDcPvD0WPuyXM3gwJSMJrDZIdP8I7X
VoI+gncpwyuur9iFM4glu/HcievKC6Cp3IljqhdLzK8wLOU2DrV8+f5AKmLpuKGq
kChwtyfqS7m0Fh8bcf9AvUFxuSgBFt8AaiELHszRZoKG2HJwr17EkI8y3zOPRv4Q
mqAZDiD33aguzdRp3NAQ47sZ1L7Q58WVYPSWq49/Vt4lACo9IyHGPqqqy7dE5Jiv
TiICXpIZ4wr8iQzzRRYVuC5SJ9/q1q35VH+bIBNkjjeRxqEXPtUkj/5gtNluiaT+
FzIBxZrQ3NGOTgKOZ3DtVGSKu1ujXeD5/8wMuSa4nP0W4tINsoD0R5YrEUjCNPgy
hX6RX4kuxCBogq3JjNrEzR8zHI4a/6tFGWf6fFH5q7OJxaqYUCCyMYKYxDtTZ6BY
DnrZ9uzYasGzgWm+1Cd4QDRPuBNEN8zW47ah6E6E3CpsFco6x1hlIgrEMY5BM1r2
UW/ZBkyInSuhR4swS7i1izxHHOouLaCUl47b0aTxk3xQ7Y5fOTyws4xeIq9Hv3vv
gaEs93VTm86V3jxBS5BEaiJFqPDnsiJxeHx55H5vWTG7aTWy0P2QSH06mDXh03cB
nXRcExAiaU2K/YpZKowLZ5LCJtQZsW8nlBP0Z60T89Aj0SNDCC6qyVt/HN3jBhec
AyPraSsBgByHnwFGV/PqP64l4yzIyFT9FpBHtHvCqE/yE8Uu5orzkg9osc7lENf9
jl1p92GfTwxuOdojzXexxlIzqv4A7tRSgg1wC3zN+PR9wsTAd8AlGYPCeGVOzs7U
XCo22zWDNxuB6SuLYrD0+5Wla4VBPmEo1Gyc1CCHCm+KCL+Cnt8JuVwFc2SyTKf2
7w0kQBESZPBBtdyJyqY9dgRkKt9O6lPSJbwaQS8H+Z1q+ZwMGTA5IVQzfuWsX+nl
0W6u20iS3WjxxYd7v0Q3mLvoY/iPDKi7xE0rrrJA6RTN7tCeBg3IJ5Ww+G25vahB
kjm7qtUhm+y5FhiqRPZ6acJgf5nb77d+JmIvlpR0PE/gAW8rW3q4lxuWItS+uocA
s2YYuULTqYwl7SiUABoFpwkgNF3sQAC/Z0W+HkkisB80joPNx0l9cBYpI1G92iRN
oDbiETECqIs8TuNmIhawSHbgu+QEtjUS+Jiabp6zKZ95dLB6lvbhYReWU1Gi68+C
clRtUFWet7tj8Pun9eVCPh59vg1v32/pseNqo46NwV4/HqNaYbpRIVt6n8+J2kbz
OdnW3uUj2o0pwq4E3N02xUTDTrmaz8qaankdIwMbFJHcur2hIbikvWJKw3LRNEpR
cmRRQsZsmMApSZ67LT+cs3R7KV0TeMzMow8dAX07UwUItCziol0+xHz+Kar0UQWb
iGQ6CD1+fecucFnIOrarWjzhh0o+BGFN0JFjD22ArFbJffI6boWDVRDC8ocFE5A3
l/K9uWLtbr46F3Dd/pNw2mpmo0Iw8f+WXnJn/GjP4Sgg8jSjY+V/rQwhtSOg6boK
cll5gRVF4BEwcu1CrOYE+Vj6bnJwwbgX8D7+GpxOVQO5N+Pqp9odDWxpRJqz/fdJ
ll18m+q+e79pU9v800rZLzkUnaQusFZdxt+HBgjxW0jgQkgX4z0EUzhmWo+GZGJE
o19QNt9/7n80fii7EHhsbd1AyNKArmm9UdCoqMO45uXLUuzmqzXGBRz3uzosTKly
PPYSlHpxbULPrr3HgfRWHcne4tzz0+/QRkDjskr0lN57mHIja3viDn/n4XCtAyOV
BCaf+y9STarpVvxv+lOFRVR6N0vZM9NiwllalIn+TpacJTCN9ylxJxCAe3ldMYVp
YxDZ+wIBS3t2R61IcMhdoRaaZayDYSMZSn4d/OmSZpmgjxwVOiWDLJPaANdfppEl
YRfTEF7UPbGgt7lcF+Xsv4TBAGawM7B7LbB+8KCXys7Lj8xuXxYcirbv57AeazT+
shVLhI2PqaBrOOIzLxn5sB729tYorQRT0P5cFHNJ3KLeDc5lofs7gPaDM3M7Noki
/Q5vikTCqaEApuULN/SKliObHnCtnmKeEIroeNhLn0pSxcTkLxXVhV5wXh0IYvza
TzBrri9pI0+ixLFaJubKxtRu4ImiN+yXBPZ6qMObzT4jkeK/FHn46qJw4ByTWJHO
UDwfmdBm8FO8/n8nFxaEYetTkEH0M+xCl6HtL1ThyXAARhK7mHv0ZCg8f6dro6pU
kSdYDAh8LWvX+HcPSNHu9/ru7Pr1xPiYQubzY26bbnwuraaOezATjZlSTy5IY9/X
3sdLJK5f0gObQ7xbc3sEknQzKSYqe7c8ito5MKkm8lU1KE7wSiUfH+3y34oVyB3i
TFFPE8s3tUZqhbQo6bnWThekd/9Q8BRlXvB9oqMBGo6p2mShh+nOkbE4KpLz4WfM
ltCjbnk35/uVMxGuPqrXkfQJpVrsc6yVvy1muNkQk8L7MgBZjeiBcxJB9IvF0jp6
Y4QxbuOG89L7W8iJGSpYd4JXAkEaUf6QXZIRGag8mKnm5drl+JDLDbwD9v57mOX7
9K6OLg4qzzW95wLb7sgQhkHzuNusxQr9lk6/L1WRlzEJj+bjxuZDxN/KT9o7ik9r
MKX//nw3cWeJl9AMJAa+r6KTHEFjn0MvbcLM1XdFk2mKNsqLlKOZ4a/CmCKpEI5+
Wr6z/msJxV38ee7810xvf0B5ftVLsmxtHhKBmUX7JF0oEDk6NUeCp8pt8sM6HUtG
g4spk60fRJ7iby9fFGmkUwFdqyjHLmgBTkYsQ96cjvye1z/UnUFFM/ZIk7kPak1R
9rL5Q4YT5X5N4UZoEpsbwIqn2L379M+DLqdV4tG8nhEfXgA9Zdj+UmtnyZdHUHf3
krP+bezMI7n0SIswixwI59q+HZsd+qPZAGNzSRVgzHlnLTzMIfyQXRxAaRorz4oZ
ZAh5ZlLJkUt1li6LeB8VMk4EFlsplFC284n9x2qApyk+tK6eV9zm80u721BRFu+/
EAYijI4dOPz1SOjxWvWI7YUChMsj2qdh/0FVCCEoDKX4NKC/tnUWk+qab9eCA0+a
G+daNPmpNuEn62ZwZGoSoDTOAmM/UlkAgaS3G/XSWjMuzbDQFZYim/wH9RRMBtOv
CRQMMt4SnIyYBWWnI4V4Az1G7TYCRA4k8p+mBweFVirtBOQaNAye+I2qVrenQEfo
UAu3V3pahWG8dgDfTUe5Hvc0Z7aY53SzPaGhKalIybvt5UBlJ7IXgaXXPaVqJzlA
QT7GMgaqJMja6rb+DczvDWgzJSjouQmgYS2c1l8/ilLUq7SOaSlDBtalqGdQP49k
EkyKNDBPO666p4r2FZlYaYKR/B0OCUeXeOSHulUkUryR/qn+WXuPcqehn/Y45yEE
Dow5pY1/tI239hhT9Qt5se3gdGl1RymcmZKWHC1lp4ZVCNDekwBp5TjlW7Q/OYvQ
MqWvaXbKo4v/jKkmFs0DGzFCt5ZOwuZW9esA+Z7oQ9z9+gEcKE63GXgd2qDjdHPg
eLfiSAdHaftrcy7/klPIrYNBQCxU0rrKykMVgkB6JPMLWT0MT2tX8lq0epQZb5cS
iuLU4FTFxwW9BMEzgDl2tA1Vv1nl7l36FIb5Rr4qi6HQOO0ZLxdvJ8EkuMcrciVM
ht4e02CDM0aPiccmjYsTxHToiDBWDJCIjtg7583rj9keANkHS/5wHQaSjL3gwcQU
wu56sXCcs+JiL88OlSHKsvWj1pvhsVTgoLu7SlmT9c3LIlRzzDHo5wGLCtqw1B0R
RXZUyMr3wtYTGZozaTcj2uyk67VPRSN9oG6t9nWKRMzKjnkzNiTKawXgB0xmLPP1
w0da9YpDYU2urapCY/TnpeuvfjUZ2HfT8WGKZUUu0pAPYI4eDPI6BX2GvxhWTA3e
H9e8CBP8dcUZD+PTj9plRdt8SHOs1up3UqDP5TSg5W16iEx+o4KSAnmmPdbCcSRb
UKNtxq/JTPq7bXwjdZunKkj6la0TWY3Al7aT+qjQ8naz8GyTQMcUyufQbZiweX/7
J42ks4Shec3ZoQp6xkt7wVTUxGmW71jWrc76M7n6l8BzMPvVu8G/hbBsOZWl2erR
EKjmC8GPe2Uldt9dw6MyOsAs6NogG9iz2XGyj8+vO2q3Qwm6kXHM/lTHELdTgtrl
tkeRVqn8xdFu/pWHi92XYWL40AQ73Y86On+rbjJg6WgwdhJ3IaxcwkLlAiLrI/3S
Fj9Q1tj+yi9t9FO1Jn+xsw1abVx1k+sQ4BilsfGqaucy/lQp5Y/eTMlw8pUyESgC
BZg59R0uuWQbgJZBIG3iQoch6lAim1DKHJfjBawwyDfah8hmcSZz42KmVhwgWHKz
EhCglSUzCcC1+aF+hXC1awYjGKcyOjWUNwLzFq3CTJ6TfOvSW0nFN9FqhkLq2nyt
kRvKujygECUqlcDuLuol2gEBK6DqmRyEbeN3DdqrYSrmYbe+WHKsIUWjilV9SVLR
2e5RXvhrSO0zMJBdOnaSWgO5qiCjIIYnLbt/8b+HDmYW7xmeD2ZFpOP8l6i3l2WM
W2fRCasKawJXyaj9OP9CpqQ3pcdmEaaEsmbBy9eargM57QCNdHYAZbia1gYBUMfT
k1NkChjro0CgoMKDLXv4YLjMHqyRLEFfDCzE3zQDAtl9jmG9JHf7Vvf3Fn/B7HWS
mvNhXu/oc3haEetts/iqRXOlDS8buQyw+Bhtus1X07lYS9M868n6xL8b54Qhf/Y9
9vRhyevbIbqjD6X9boqFF8IeA98QBCwKtO0rWIUb3a4+/0wxFwqnpKvLSKkV70DW
Eo1HWTndrh9veeQjwbK7ogsHk018uysIvtSbjyvhdbrWLUaMVx+qwv+L0qauJWpI
kMEm0ngzC6UnW9qctaXNcp62abVI4oZMsHoNaat5s7g6Xv75hIx9DbPx5T3i/v+M
BzcWFnYYsNITfAvbVk82Q7Zpc8CY3uhtDcS2GNElvJ/jU9e1SHyOgUrQT48cRF67
YRCUoqvtGv60NgMGk/EzJBepdL1ckT5JHkbd73MJO1kpz09PluoVA0jSwXvf3Je2
LZTmdTRBt5LKteAuNLTVvvbqpI8k54fgehRbAYwsXu25TJkNGCR+vcavtstooVQ6
8qmDXcO9c8eXKtUJYym8IJ3s6vaUypJGqvplj7VQtaPFRIFFDX6fhzPnJ2RPIVuB
YDzSyRYt7iZWFrQIeeKvsvI7FpddBU50CHqxje6E5qzZqAupNL5vOwd0luwUQi1R
MSG9BBQwgGeaecwmSYDci/w14Das/Lvk1qu5pojvBv9bYXgqsaDePvnsuQCi83oN
3lIIOF95IvlOPXGDfD+/pqwkXAF0re0zURx8L+X7e9GqSU+VxjGv6DwRoQmULeXU
uluUdOFi+YXGkwlBWkXA3lQjAemrr6j+fXowqs/qg3uIleLI9ni1oPJIrAB3zWO9
h84s8pOKD98M4k8ZJS53HH8FxHswXvw6tAco0TkMK4i8glvcgItLr6jIIeGyIyBC
YuXxLMfQh6JCEWmdPdq9XVFcSbZmclyeNLWUrNAbkEahKeMSoSE4xmEDvdtYB1ul
W4l6meGVAqgsazTDtQRwNihUKXrU2QVaiOmDbqUAY2CsCQK/Fzyj4dVe676GWbG3
+zNel2TsKEyMgiaA3ECmlS3UyBx2gKEwPh7D5hpxD0PUBWs9noiWMzX2gHpQYzfP
ChUsLF+HG85YiF0+b+kvK6WvUweC278c8HU8uUM/omM0xPeOEMih9qKSDJuk2k+Z
UVB2XUlQWMHPYYgkMyeUPh6LF6IB+mGnT02AcC5pYIRgr4f+6hVE3WPh00O8JJoc
hKR2dPNPdrPG671w3R+byGV838Y7Ek/JNGYGdOUg/Oiv9C+2ImQEDMSJZ+bAEHIm
wmEPgwkG5FP9tQYtBtJy9lrdHljGpQJ55hB6nHvGFXRB19U8cpT3bQFefudaSwRR
HA8K5IZrAag8XjV9qmkV6QWH0DN53WVcEB4RweponBKO1vpmF0OPyfgJJnugbeic
ROFKCTqoUWKJ2Ka5us9aBY0Tr5N5NNC6AxrOUeAZZm8Qtuz/nPc0bK0f780bqy1g
sskQR3BgR0uVajGFcuQ8l8Nolq4zum+vx+J/GlJj/a/mz9dRy2Xahh1bCJAttHBz
pcWNL7oBC55wDInck06vkRZVOIWnXwHo22Y2qLO8+6vwoBy6W9Bm9356RUGZ27Fg
7uWXjhCbJJBapnOEvJWU1wc52cJyJ4H2yVAWbq8H1Exy8F3cYWrrrkEy1ipSR8qI
dusDH7ULIqAhZJw8KrV+UlMLIXb4xYI8JjN7ILeNEY+sTwS1B2unz1gqN6R6xWBP
DMNF9P7yOZBehrs3KCeITOqJOK4R2yGyq/meMUCt/01jHiNJwPoExa2znDQIZDgS
VVldcMwvJrpTKTSAYQBJzspeyg/Iw9IwMVinsWDqStNcG2tJifXOZStk2zO5eXO/
hEaALkfcUsS0UN7Jq6rFFqfkUaQ9/JvHxbkcb0nbAcVVe83MpVTFdjAoWgFmaQ+6
RJqTYtSRRmWPOtjOQQ3Qf5WRFD9fcImtMGKd9CH99ZuDCuh+sv5AwHekOLelIfVi
3nbhzRsVHFZm4EMoeBVv65oGqJrXP+eO659vXoB2ineIyvyGhHenAi2Oko0t9Kf6
Fxx0v2b8yl0f1Wqm8+/1X5Aq83JzKUdrf1k0Pr0nOQluKT1jSvMNIbpRg1KIrOKr
b97MwonG4qpFW62ykv66hUKEBwetHm8KUffoCOgNk6AOGP8LO9m6ezacKg0Vs5Gc
n6M7CyoU9q/qfyElDhgjAWhxpB1NLoAv8gYxdyNjSEbZwD22K0GEi/RnweSrNg5V
CseRddgfEcNOFcVDkKvg+y+SvKDuowFHaBc0tjvKz+DS7REX9VEjYlzCKZ5Sr3ab
GADXBt+hXv/bNTxnGW1uSm6e1qCm7RCO4lz8qACEgINcGFVworliqTD/QUjn/3Ny
4xb9lOWApe/VXBjbBMyiq8M3/DSs3/ilzqcq4XhXSw+H5/J90PLMV8vsVutzKf6D
6v18VLXR7P4gkBVvxpz8kuP8DGnYZV7CC+X48V09DzfVzuWehkdySjmkkUZ04vVH
zO4UAGCogs6qxmuTPfGywvZNT9DAf+D409T9y8blPAajnsxThcjymqwrnZpgCCI0
4W2ysAFFMdB5unhDUYCTl6dS3fx4dirJSFmO3/BUg4Rlz08TrYHP5cxuJrpLLxSp
L8O98Mb18pNK/ftYPFHoJ2EZuQ4Td6H2sNn9LcmwreZ/Rz0N3FOcPTYUAkmJjoQj
/Mc0zku6jmyJYii9vy8VQaln+jxdOIg8cbwuWxOpHO+Li/1Z71WiZB4MK87mfkby
whoQPBDa0992Zjn61MyoizG3FB+USDAygsx6/CwzTGUy+nhqlmtz1EHzyrd2/LMl
7l14gtS2TeUxgQ+vxYp2Hxr3vAF9hvwYDbr0WVFMAJzcGMKHcEWvsCEpZK8s2Vvz
c/aoFVZHW/8xGQuUAsO9g7x+tGLkdH3s6edjM1ehqQtvrnPBWW2FttzsCPMi/ui1
wFtqmLu1fEBpAlX0sKWS3FA8+5erfWjhClf3IzMuKdsFCQySutpDB1aKuEdGqPVJ
7mo9TJ/9/GRXF7hZCf0iEAqMa60TPSvAbLSo9ZoXcDfKkg2+eyOtcZzSb8Iw42FA
pmnn01IChzztJDNxxoUXSa9fAMg0pXI1IXGq7NqrePtDqyNyTp6rTET8ICSqnpvf
mn2vE/4BYCYmsbGDLnnZvIu7EwNCoPGWY3F45I5KV3A5PmBAewqT8bQXW8ADQz7Y
jooHyD0VlDu/gHZUnN3oXF9YaKmsDrzblcFtlyyxv0WOZn14WpGj63rj5KyVnA8F
g6ue+9bShlj3eltCtN5GUydm+264pZiA2uyCvZqVTWIM9DpGT10oc/Q2NZEnxd8/
ogVikijAxSfD5FR0KziLGTryiROEmsVcdy6sXAXcjrF+vQj27Rn9s3at6FPsz3/9
wzkYicdfgijsKkBmxUGev7KB0ha4dhtEp4FUvJS5uLPpx+Zl8vywkX2fpmoio00q
PWnuIJipjgY7u5Z+ZIfcxfxeVEH3HRwHYBij/NTIX1ygw6l3V1eOCFfVVZ4TTjpQ
r88zRabxGNcXqK7JwnlbxD5WMu44VvhT6LVXSceXxM6CCegrmmNnnJDUfJoeO4G0
lba/pYvdsKRbTWEsad8Xb567XKxnq2fmUqC2yMypPzii8z6jA8/6mamUFNVbh4Zh
xUz4LeceI4KluX1VGjwX58v++/nHNIwu7kE/XZHXNmSEozPGmawOXz4RTjYAwnkj
IF2VRzOPOxsUZh3KLXdgk9GSBOnGbrTnMmgIMUdc+luPl5kJ7mBn9capvdHpim7P
ZBwg+InofIuEAe9RNdC+pbjL8E3vwKsUH45RbWFYcBjU9YG2xmd0D5SJH8JMH8xQ
ajoTSGMipizRr2Er25PUIFePj7JV7BTMQsP3BdRIVQxFKXyftFyOXQ+6GIJC/dgl
fKbBAJLp9vKGVgw60MbvG1sy5p4E5ZK5pME1oMe4JUg2hE4tYNHjlsHoIK7mrpas
8WTJIkwVqFdvu0SiukZepyRJ5ImTLRxbOiVfd4ruvqUHRWlQ2dXlgknb4ar1YHO7
Np8H9morRTAeYx1qQZoTPamwuqCH5BQo2CiiWNhSWY1ne0/XFKjDYlQ3DO0tGxTT
BXknjWp+rw9WDprjHIFPvZG518pqUp2yDR7VEEFSoXqqEaKdXGtB3LrzEbAHW4IC
ThkQsopgRuH35fntNNMId3aeloY43sDlt55f+mAquA2aY7lwa5Wh30/prmZdy8Y6
/2itiHwqkmxIuTz/Qz11RAZ0c2JOSXjSArHtcFj6JnrmVNXsBy9buemWdvhJKygY
LQX5GKFAdImYwRe3yWXpxREepANF34E8HrIH34R3rhXgTILS0nx452yog4GEeYka
oVb/GiIPwh+HUHwkGNl6CRDO6C4ChpUicgtmZtXdJSyg7kQCtNUCYFdgZrk4Vd7B
EFODWgiSSxZh5GpbKeitBUXPdgrzaypncgS5gzxj5kBTt9J1u09kd1vf5cPFU8TX
UVC6jTuW8idku663daM69VV1+khQRCwrad2tZ8zLomtr4AXb6RtDDSuMjPXdU8v2
d876kai5NGQeGe/rkX/Na772cIuRWvc54eCgBZ0yB/taEjdQfChIndtMQIkipWxW
ZzwVMxIVkotKyOVbzvu5jzAqdu7fGsyZNjM//7TAPY7M3VtlUjfh9uyeV25HtiOR
eba3SrCmhQwIteWhKTh7XMUTNQJCTqNXfH+Ef5YPY6zZzshYkEfeJftp/afe+9B0
+zAL0xWJmC8wRWX5rP//h+VBncg2vumTqBElIHsgSLDZI/F6k63y8k0eXPeHvgqD
qSIW/GuNIPZ1ncst/99hW9VTfWPxIweFuNaymnN+jOYN2DsfsYfplA4URyEkXZtl
XIqeB6VHcuqISpyOVj4QY0zUojgtO+LBAfAcfiMjheTrnwAkVDacbpijzcfLqcRX
gagACVkW6kL0TsFVo7lQ43uE26jLRveiy6e59A5mwL4IDqWOvNcKordOXk06PcYP
PRvqdVNewGDWgag5lFQTfWbBaHsIDwUfGhBJviYOLHFYAmWw+byhvH+1CI3taZgp
r4ngLSlJ9djnTpt+A7CmX5WGBdr/5Y0l033KwW6cqa/FvoqinqMj8Czxn/PXvTln
leFOs2WA6P+ObPX8Mw7myZrb38FQ2A7sl2xI6Ola8psuk2u/N+3B+4pNUPUBPndw
5WBUFTs9FgVoHD+vzDdbxxG6UzPptM2w7Q5yr7mLoPNclbPYODhTQvRacUGY514q
EJaoEb7Q/uz5oH7aoAyteHoLe5QWHTWb4Qg6LrfqQgfx57yKKKGmVEQEyhOcpEHB
iBYHPifxAQZcafQOljqeWaKPmsY46c8TToQ7gWJlrXZmXcLrSaY1UjVBeIiHxjJf
xh4gyVOMHRI0mpVIHXE6NA+TF889RIfYF4lJ35eDdiuFkUeAba4FZUDv/KdJkA+E
ZsDBCjtACQ6I2j2K0KSlqMEE3iZlUsL7Pdt+RRxPe4gHXM3404ROTVtZMsw+H8qb
nAvNDqiUa1Rz/ssR2XLl8C0iW+/L+IEnWr3UQT7f1WggMzNqMApseBgX/BMKJGPi
5wm34iUXqdos4aKghE+PZNfwRlXnsZIsUslh0wu4zrWlg2zqXVwTX3FH8U6KUFHs
22EDyH3bytwn3z6RptmxGv7r4KrZuCDfR+nXYMZACqwcfGh9cVxPmCq0Clh+iGmm
BQiEpmxRQ2ieM21Vhn8HKWzN2jBZpt5n0+asRlpmrfb5NebozEMH/Jo0BYSCMvyW
nN9+yj2Yq24H1N3OdAfi6W73Uipa9cRicQe7GUiRCFrhutjchGM7rRdTCwHiQHdD
bf2xJaRgwBFmomSrTmfqwC8esl3s4f7eor/QyFzV0R8bzFJi92NuJ3OjjRevOxNZ
wExSFOaqXwoIlSevRtXYIcWehv2mrLXIWBIdc05KtnM7UmurOE6HlsO2ycjibyQM
ZOswxwC87jHMbKEJ+cTUkOMHKB8rCr8jLMvfIf/2xl/7vfBR1WpFe4KKohBWHUPs
nxfXBcQhG1LsO7tVp7H9KrHFwf7I5G0Vy4CBm2gidX00LE0znF8ijX9m8X9gKTon
8BK54wpBYBSnG6ejjXA16nueK/XQHPTvzPgQ85x/NLbGHkMuTufSHARzYiprZ310
dzrwZkFsDjnWSXC2DMsoNvfu/lF3al9qK4TJO5I8Px+RtBeiU3IKdIsCjta2ypRZ
xFuyLCXgg+CNOV6Od4p/I76hiugmWy066JfrtDm8U356krErde0xQbZlB3Mp2yJr
qBll+qlg0SnDK52QtEcijJWKji9JOnylSADHUEH/hpxioUERWGKAaW/S6JY96qlP
i/wus12zWbZ7AzWoSzmmEFn8Abq8S3MkPgsqB6k9I8cl4kcCvApxedqJwwc0OW2Y
+KC9dViydGx787C/vpHz8OSLvNmO2rodTcs0JOzaifoClcj1RksTr2kCX15lYK36
tj6SFrrjXnTs+NVcir8HeZEYqQ3SEKplWXGbjlJ+hsvye7Zkd7OluWqI/qZANN6D
8VT1/133XL9Xxbnx5i3CaOFgnhPn98p9bWJzbf3KHPrdpeAhfkncHiO6TadfY0E/
Wh18urRmOGsMRo1Tn+IjAjXMCd+Bgdrc4gPHvWW6v0QLGL1Sef615Oi5sl5w87aH
kwT+JxEwF8YUxkmJawFkL1BbeNUEXhM5/Zr7gFVG9LRt5oFmXziFjMFr6ob9jRmv
9RtoaTVtMu5LTiPjEWHAau2IQNyIUzncbQzH8TcdQpE38LKoX9ttqf19BM+lmaZe
Y6JMW1CubVAldPixR7ecwYkC1yCV9L7zd/k6MlmzMKpnPGD1pwbFVTktZa0oeles
mYWM72sYVQgbiU9wBGdWa01m8IRqPP8dS4dDKb7fdX7Q6xL0m2tjAdZH2Aa8qJTW
5vio8hs8qIkJOuuAot4EurVEmTsXEd1Adxpy05caUYOIan89HQRanugKc+I8+3lq
i4E9JWDRbeeXAAeOBiN3CzF7B8KbLxi027KjC3LPctvWMGPqB0d423PnuTRM+X8n
/9ISDBY+d3iaRcxpi3r+p0eSfXTr4Pw0kS/kEhLzJ/jK0qshOgy8g5e80KUf7psG
06OPemhLI0CUREMiB6OrzsYbwmioMpsh5CfzA2NJUeRHmq/JDP3C7e7jOHOTjbNd
zUvRKK/FdG4Z+l2AKgnwffGVQDoWAKNUO6WyTXpQ8zGhGX7fgrzRcQVrnF62bL2/
cKr34owi9Q/bGjKi9Fc+hzz689hvfxU9mlYLzZ7xIkCZtVHrB7KVervVE35xVAlB
fJjupED4dP0+3iqVvH0YEQQ0euxiAJxDxcVre7DTzcPC/jIzZjrjA01eby3JtMFT
Sfq6bhy3L1Gw8yMpfvCt7MfqFvAQA1XoDb2UIFu01f3jXwlSseY8cc97iTVOi7mT
8qwE3r+W0I/eC7LQcndsyPVjs+Y5Ct4uK9hK8h3IxUD8fX9R4fTvpFzYvl8CG231
y/tYahFrE1oM66FPFB5OaOAb87fKJFwCB30OXI95jJlDcQRJnqMpsU/lbfeFRtZN
ALnsb4WyN4xGeFqZvt86z06O9gVrPYhHkSn3eDDrecsvz1AGWr9PxhB+hzV9i/yk
bnfCqzM9RWcapcdsYXmW3kSCHqQa7mXcvVUbaRNuANBWuqN3dKiiee90rGnHRj/5
xFzsdeRtPI9Y5yq88wBhfuW4D8Z00yqkCVvB98eyWeYeNyj9r6YTnS065q3f9pqa
b0EVTS98KRzUKxPOJqlZo73WEc9i0fApdYPy8p/Lg5zds2RIkd64j3rJJ9lNRTth
6uF6HIB0obSn3C/uuDpMjcTTElw+4bn+gM4fgEydkkH+1QxqQIow7hPLtMhgh+2h
EupRwfX+kr1vICci3D1AM4exVDJRcB5QHQWPxdKGvsSazV/+awaOGmMoeYLwSmlN
McyrjuL6VWo2IFcynAcaoJZagyDYS90F1Qe8ueyiPHCT7KIhr4vFzYp5cCaWxDya
qK+eAdn8LbD0ROqVTOc7SVm3UBAcYnlPKcM7NWkihvspmv0Z539n396NqZAo/OlX
by5zhbYVh4V8xFV708sCllImP5zt6tKEIpi2NtsfFMoSJaipBYGBfhzYbCvsm4XZ
7PoRfi2ktE1wAF5HnttX9TS+9oBW1o9IRahOmaQ1g6e98/QncOHLnwZS7WXPGg79
Jr4HcJykX+uJ7otpt0hErxWiSxW8w19J1l4q2P6tv6AWUOmjBnFTasETWNvMbPfR
4QHKFtLs4Bg93NlHl2SoC/8E/x+zWifKobUUY/d0oLO/MP19Kutl8GiPQWGBJ3Fn
6mE8FBg9Or3kUqI9Ii6nE99tMhRz0S7NklvG4+xECDEBERhdWXkpRN1/f2AqfnMl
86C2icxxRHvQZ1hXKV9TTSt/z1g2IVexnK20gm1YqO2bWFpRa/mjyxFbGJ0st2vS
IjlcgCYXFI2CR1+UtkbmJF50/7N4lEnLinszV8mnxh73Wb8K/1qacw8I33c3qrVF
q/Ncr4rLzpK5St+XWTibasfpvGLHXkKVPXwDbYyPfaHwV2SMpZBXlB+zqifBdTZ0
0ln+XgfSZoHeijdBNpZvfYY/1L1VGJCJYZ2EqG46++jiR6HimIhLGNTiYKbZ2umU
RHAYoQfRFzjoI4nCcgDSpXIsGZqQqfZHbdy5Y4rX2pafzlLIitxMBQYb5Sw7NYC9
fmLMpXu16pCKty7LvLFem2kc9JWv0MH6ZkS2O4k+L+rMrvFxOtZ6/ut26XFcDyNJ
motnep5APt+to7P8UkpZRwEOvpyGk223lHK+HZlWyc3TSFQz0vzzINeC89Fla2NM
sGkEBnx4sZVA6B+SGAHe+L7CWFyzZuXk9OhyFSl29m+PcnVNpEnXo7vcrfJxQ/d1
pTSHbmG0jw+CilzXyz3yC+ITYzL+87B+Hnn4xAuUSKAwaaJJEHYaIWx8QOpHlvcM
jurAFmvprh26xtsGBeCJcVtmk/H4DipW4cKaZp49xL59nrv0jAGKlvHq+rS76B8J
d3+o5ppjZF5tpOHSUetJlfig2/nk5qbRl2yD8k0B02du/ivnvyloJGUapxoTRvRC
XDYQLmHAGp1SK2ZlFfdeee+PlbzCec5a+GVKBKjhyP21DdQrUOVQoq2bCKViIwau
+EwewSaGChamQEUHs8HceQnX4ynI47lNSJNR69f1/LfGGaE3HGOU6VHMOe2h5u1d
PMJ+V8rrUNsppSglQlR0qR9uEUh5ujQA8+DHE7fsgHc3cM2Klh8LMAhfvdOfQlWm
cstPqzwiWgUsqK85wRxHEz8YXaHS8EtMm5X7wHXZmt7AwScjohQwVwxHA/hvFu0q
jeH8VrrpKLZXSfvlbk5IQBJLJA2hjX2GMCA7bd6BHXD9R5HMIbWBxvqegzH/b8l1
bxVX0Zb900c/LN6oIir02DzlslH7ai24lznKhIoaStBTpBtXPTlZ7jadvKuZm8ya
f9xc6k8SrL+r4Xj/T6ylhR0upY4pdTe+IyCJd2+ZHB45+6bg/TmByN5d/YZ3olV5
mZXfN93Th8h8Ij1lCQylOQ6xsZLPlVW3ttDO2TuB1gd1jJe3ePqOpIb9gRbCESng
f+hs1YFbh8HWIGeZQgHfkPHp4Og8I3z0q+GD2Z36sDIkpLkDEUt4FICGj3wwwAfD
WSXZxLtxfa4FLCSA1H4AZ7vkj9Weivjp6vx6vpNlve8xpKysf1PMtxsPWKbV/BVr
o0DE5rm6LKtPZ+3m0ar1TNONafQcQQYLLUY74orf2e02LR+IJd+nELa8xmvI9iHp
YVcvN6bhDJsi4Xnd2qlSXou1ChImeF5S30WhTuxkAmNw4ix+eTydXR7OVGvPW+LC
2dCm1gr+Huq2gJ5FgM/H4A5RFcJmzdM8F5D7eVQuBVVCd1m+OeycfavoPkw/bo8Z
zbs40ABVKypjb0/yusk5N5BT3aiMOKEW2+7ohW/q4tkuCqmjI5nLQgccZxwWA/w2
mRnoibAQAq5/JBjeOjx29r5S2aYhCxoSxOT9mTEIUju7JaFe/YN72O1iS2nHEzgr
sbAX3D6omekZFP1RCxm+TnaYlNugoR7phtbScvL557Ph27sc22TSyyhFSzJMdvo4
wgxzAf7R184+63ggWSidLh+8sUNAoadw2Db2MxlCRKmQ7fbK3UgTljGyIlNCjHnF
2s3nHTc3nhr7SeLajLFdXBZtINHHAtSvnG+wK4tTyvFJAhtX5bQTpnhj3PHPupBL
/BI94/l6UT/zB6cIOse8vypmQHBAfS35ixx29PHWX/5f6uM9BnBjTgYMhH8Tovow
ir+vrJDRYj6qGR9jY3UVBl0i5Z1jyYqchW75PkxL7qbII0Y7xhxwLnugnX0ix9g2
4Ag1V2DUfl8hnbQdEOJOTzN31d2Ujo48X8btMzNqYOSCBp2nshwEdrFSQKSGpXI1
uJbqQi21O0ti84Ner1oi9dXtzD2cikwPUKRV4eQrotftYtXhgjkLCJTmT2W7oHDQ
ECKLSBNB4qu2wKe4pQcFhHxZHiunKWyRqrVsvDui5nsimqDxoYUCImIlsCwNWenI
6nRJoVUUeoOUe6nGxGmVUZim4kMKg76PSlMGGyrWUns6EDB8yNQoRpQYBOn/TpXB
xsnwyaALVHig58gm/QEzrwyMHYsq1U21vazsVcdsS90Ijlbh7Bj7rY9rzu3U77Ee
53+Gt8XPbWi6IvHP/21R/Lllbisn+0qSymlveykegXvY3vL8NK6MZhPFPUCP0dWY
TFU2TzOMViP9Gy9YZ19EGy2psqzQoo34+fHGhDYpV/XYlQE3VDPwkK/CPxmyokJr
c4gjkAtO9PAZvVjsuNsUMFIT59y6D4hISzBVfS6+AQZgRImZpEnKpUxEjwub7Li5
lRgD412RmWPHTFi3O9+vt+2Drf5C70mWfkKB4I+KssXKmr49EY7yiURu+1EnYM4O
DIxNEDDhUOqMf2YAQGA9h17LaJqDRTwqHwZMo8Z8vCLE3mbGPj9h6so/+5cFV53l
nNMBzpq7Sf66FTEep8hZJ7DC0eENkb2UWOPiI9SCaSTGWeqIMeCECpY1SMonJ6wc
GJLCd3E69nEtPsVEzD2XCNDqrAgKdOUGh+rPUx/OYlaNbFM9TOsx/e6epi4WpvlS
Z60mCTeUAwtxEqHF30HK5acnLXMzNZOIewWB4SVdJET65taD0RG83MUiQ8Px00NC
wiU0Zixqb3LgugjQOSQbJim53nir+JxTvMR/BTKQCsrhKNrxTwfOj1iVt6Smervj
7WneHFlUAMDh1ZXRWpFGXGkKpgH1Fa4Uhmn8zNCsn5po1zSx0eoZz/vLvizlXmyI
AyrAu4KxBhJvvzGMk+ph1c+BD1ddqNd/1RA3ODtWbz9YllJ5cLk3FKqDtWhWfWf1
tnMTSQZ2Nwm8JrRI5Dz45h6e8YcWb3hrcgXd65w4i5yVvWSWRj0rhQrpFGt6U33s
ZGREoYyv4EYAW6ARpKt3eskOvW/souDOdyKChubSM7Ly+gGKPl5XiYBC/FWeLR+m
y3FslfiNpxIcwWRlKJTyGGS8YiZl1Bi5vPkgBRr94oGOxZiBhMhcuNjWOQu/xupz
AE2QWgoiNpRBElODbWrsGY6y9/SDw7x6OYy3b2C9Tu74RKLZ2+BpRVz7bZFgeVot
Vf/2asRcXa0g05PKCWuZJolOBKfEfIKljnhWMDnlTDHzDodo1AqA8uTs0HdiPwWH
MwEJYm9PCajyODiIW25Ye6QGM6ghsPE0O94ebgdLdG4ZOmu6oqu/kWnAu1dVrJTp
x1CC2WcI5OYgB0xv4uzOsCwZHpi/8qB42Jkr+ZYn33ZqNau4on2795s+z3upZmXh
y2qVBLvutNfENpL09yTNjkRgw5i92egWknON/l0NbAgmGtKTcHVL1fPRIPqcIvcj
7qBTKeVQYyI+jhCz3cwRRfgbQMw21e/zBylRQ4y83m7kq5SCZIj74HWzPP7TYdm+
8t+B9r8hfk/YSlXS1Rk17ebAwsVe3c+SYRsBLLD03yrvfsMRb37GNz1GXltKSm93
vMV9k7DSUZ+b71GIqY/OGzpvn1NhzIeoReb9LUzsB4/jo0F19YnCncxei722neJm
lZNORWR2755br+XkBGJoTv8cxewOV4OlW3d1A0VLBfL/4EGPYbM3XZHOeP85+UWi
eDDCuIf8F01pprmHNZCE0Rv1uj7X8KT4BThjvvyENI64kuGsvy1cwQuvaH++uWWr
Y1pPZApMzAboq70Bdk88cnHTD9FmmqoEu9xcAZ95Ozwxh/jccEee9++pkanuj5SI
YDVSJEF8I1NPPEsS6cywVhz6zDm/Woh+RY82f4uKuYFIpqptxwSsB9y8DNF8+17o
sdE1ctxcSy/swjHSBE1DCzG2biO2e4sg5nMbNrk0FdVUr16Fi6/IQofPDdORC/9O
x4+ZXuJhbTlGvVmnF1yPv3N41eL4fUUZXS+X46DUwv+U6ww5FMZakuirVp7q8+N5
UGRMZOpdIrw4CnMmzNyakPyGm2o0ltY8HVVDxazrBNmmIOdACeE4Ln2Gb6l+24wA
Oc6ZmsELQvkpuzACXFwKDXR+HJweLuqw3l7WbcHOiHtKGSCwU2Tez+jvBrDvBDVa
ukri0L5e50iUZHKwVhEcK6P0PYO5K+4nFLZ2e0Z2rpbozL5pwOvEQWcHsoruFLHT
TyYbh0rWHp1QGoaqsQIR0wDMxYG5KfxbQA9fDbTm6Rz4oPudbgrz9+QkNHkjeMru
oP1lNvXeSeQcfv5IqbqLDVTJSDvWkjRKlG6GqkuVj0VKKgvG/NhS6G03T0lckl2E
x/ZcwmBt87k+dZB3SX1RJJSOjSMAnjyqs4jHEb+/4FBj5znTGcX6M9L88WVZ43gr
4h2gpiNGMvbDsHzgzCsg5bypngqoC8/hZYPkfUXtoT0SFV6jdlcGgO61FrScB2ds
vUMfFyID4Kl27qyh7jxv8/ZRUA4RREKFjfwyP4uG8LtUdkOilFdNnSsUxCrL96RU
VwvIK+MUfnXxJ9viZhWsGEpi+KEUhh4WO7vQEFE3WC4vVmok2XYmzu1AYO5jB6tW
MsuzJqZlBDG8SGxINYBo6kT6r7FqanIf8FDpzfZ4OpHKORbdrprVPdkoi/9qAnr4
AiyPifE+Gz7b2DqeS1z+KXwp57gFHpJo0rikVQX/cXOCeiiuZjWdqPl7CXmonBSO
+RzkoytWK4vszxWjJkujjkoOfKFJyuOkVj0lvRF0Ym9X1cwuyqMbp0pigCb9XUM8
yqzT6I+FSc+u+1DLxuK1mqEo3IxB5uXYOifTELtKVR+trjmkme/tmzPL0lar6lb/
waSKUUoj4d/hi/2DhohpyKBJI7JQE0lluCUYouTKlUxjAdXOAJmMXrVqMQZJmMqG
pdbe3O8+Vc0fv+Azk+//KMbK1yUpIpDrclmCoru1Gh1XvOsbE4ppOgrSg2mM6eFo
q8khe11WUyl2bUSL/CUhVQ19N/qX8TxG8cQes0v7L47tsEwKob4D4tqOlAUSf14+
6nup/pYcnblriWv5Gqz4mWU4vBwI9hFEqyJRSImD4ALZ735awAZaiKxfEbI+1np+
nBPg4TbhADC0vkucakPrRQN1/UTomtr6Z/pJfdJ3Y86nwaXnWZGYGzL6P2gEZmmN
QouA6wG0QW3Hh/KOEsDpJ6hrARVL0cXfwhk9km9o+XPHPNCAlADoYAEVmI3w6eeY
V6qnYhTg/z+aILd6wV6PT6gOQ6ABsNIMHfHyzCPIjMPXss5fdf4ddRj9xUQxLcsk
np5w+zPCpyhZCKjaZUa3V7tUOPERSCDMIzyL4d4HNWCHD8awq9ubsxPDKLeAGlbL
5pja6AMogO3tl7vgcPrx9F0oy95QU40YHKdQwgLKuCWSU5uReF34ak0NlNWJXFPJ
HeYQQIKP2R8D08LHg1afnaDElxsijWGNNs42qiUEs3PhMbWS7K4fRbLI+mMQUz2k
kv7Efl0Ge0+xT4S672sMCeiugbQInLaVwI6UEhnGmCFVUk5wFmyTymyxdfkZU1X7
CsZYiDVbFGV9XQZCBwG5tgI++o2Ke61iCry4X2lWXzVWrE4SJeSVDwTZFcd+g2+B
K3b1UcUMcV2Z1CieLtrahCabnO06P2/roKn5mOHFdLuj9/BKkj8WiPS2k1HODPrY
G8jnX8KCsk0UDvDJMzJPkmKr4xPRWGF+QP2x5EuoO/Z5FD9Kp4ieR3b8BbNg08Wf
tL0qgtkm2g1SGtnHnPJVf+9qSi5nvMSke3BHLuyptqRQMEYY3j3DerV3EnGpNji1
vM2woWcMHwSfXdEokXf9QGzAUGWSAR20lJLuknrV4YC4v9SarzRW49Hr10viXsKQ
DJgbSWOjvPZoz1IlCnz4PVJcDsjsoqBQ1Hu9DPL/xzxBl00XHEmuORcy6WeMXyeb
1nP5sA1f6/wRxfB6WKCtx4+vDyhYycCOShMbaXpdMVbjh/ZX1UTXkuuwgPZjTMJO
6Vk+1EpDLJWZhR1IHnD1d2avcqTwYDuBONAu8N55BsKjMndV8EOhmoM2gomli5sM
IzbyauYlkhBG6YF0e9cjAnXFs+11nS0BowVHKasQWvXSckW+Fu3JVxDaQlxdqkgj
b+Vs3xmte1KO4oR6gldM9GyfyY6QVxUrWP4WdOhISGvDMcVNpGGD5/YODNUrmdRh
CKnLz4is2cyXLzLAs3MSwwraE7kBaucOlUT0/+9lAeamruw83q9hRc7SrrSIb20J
OSK0NB4cyPPLBHwhxqhd8Le0hNsXW7+jyh6UBZA5yPO7HZNWX/368NNPoNuc1wuV
Dj6eIX02EWsUbjRqG12ygZ5PWTBW9KtA3K0ouTv4NZAgzpfmso9DMak1FLvqerhB
ZCJvCwzyAz+wB3eZ+HBaYDygVyvwmpA79kd1hjiVnwQalpmwBq3DJe2npqxPF3pj
KcMqnfBgUEtKDRrodS8ThH2IK91TdAgmsF6tQ7N19u8qSp6ge0V/jqH+D75r6goT
EncypXDrVPNNIyaohe2qbpMoFMWDNiM5isal9WEObg4izMT12l5PG1yl1px9Q0ZA
75Nyvt2CkxgiKQNT8EZFQaoLf2i2SlMCjTL2XGFw3FIrJq8V70KpKmhJr/0c+iBu
COFnTyRvm7qXz37iF7YDCZSi1U7O70L3mm0c2FJNyU3sMr8LJfZ/i4LA4sFu1lBP
WUnAIx6cRhvEn7tQ4oMHJ3mnxFhejsiiBqN6biIPg4HY1yb76czoY2vYeSwgzds3
tcqV1ZIsMsf7LQak8Wfc2bgcKe46/ZlRau87fGJyhBFn4KZ/BvINc0RoXVspwc48
2+d5NQmGhethhyMH5wPuXrQbKtOTE/oFoJOvUvK1FpBC/31OPw4XmU778V2sH9Yi
NOpUsOCPX4dgTtsRHnWCRXvCEssTiRTUjz8BX2Ymj/makYUr9AxCHS2JwyHb+i5l
+oIO00IS8q/fSS3UgHF1MzvdtHUPSeE6Yg2vfv6PUQHNgNZzs6PfE6xFsROojx9h
La9dT+hnbt40uJAN20sjffg7R3Lc4Fr1YkycQRyl8J1cROR79Mj8kjXCPioB/+ee
YgBBC64oeoJZ3ycLggDBnCueI3JiT461UyUWN7nt/5byjxNMLKTIE4PSf4hll1+L
tXKT9xMhz0CjTRn9eW7hi++ssw25RqMTF+IwiUfmPqTtVbun1oUZp2DJLb20GtNj
MO8swlYhxJ2gMHeztQE5mQK74M+2TXeYqneFltECY5QALdHJzwM/IK04/WfVIGE0
cEakhR9cC7tAKbaLNnmYOxiYt3BqwWN9c0p4qt016xtsQ2wm1+N1tNMYXBxwpgF/
rgovjVbrEpS8LBH8CRLWsu2wElvkQgqe9+2v48qvsFVezfY5Arosn+PYT361k/Ja
VC5AuVGz26Cd5bn2ki0sQT0Fu1SzAZtdvX1j7Q2D8EXS89RFZzoj2svfsmxgJ+Kh
TCCWRS0Th9vX68aOhzVEPGRd3xlvSVIVTsn0CBlbWz2uBl+ARDX4kuxP6LFL17Xp
pU8SNCj0CR1odi7XPsR/BtS21o7z/da08+9ZKkpoRhessbtKr74elndG6dDzTL7u
48OlrRgWKpVif9cOPri1H/eEjRh3E4BpDii1RUV63UkILVvOshluxhEg+WnbXG7E
LQV5PisRPukVkkVkhaKWR2qCYUMxa3z6xB8nBXT5iPgrP77tzthblERI9zkdBrqC
AT6JerP6GMqiCklV7mc6EgTHc2x27XuVIo4+DZBi+7bqP17OHciX6l7GrS0S4YMb
61faqkdMlb7YRd/ig511IEJiypI8qE6AJLxQtI0BgpABnA7ZT9YSmLomCjhEvi9C
xmxlE/MjHQdUXQOOYe7H4tghMlr2zcHr4p/jVw4E3p/2A2qoNkiWGpx4Vd0w/8wY
MS0pM/PGWWVFeWMCjgQNOFG9pKieG2Lx+Kwyv6BNHhF6bi/dkro6FLXJOW+EuMzZ
EaJEVMxhBv1cBMEYAfZeZzJdxHmDgkYarVGU3OWSgzpDmttzvub+gKHxWBPJ9NCu
dygsvXjw1GC7GqC9Q4GBOJzd5IQpcf0j3o68/wy0zY9myz2LuPu8zrf3sAGYLvsX
Y9FQ9kaV2Uj7BrfrRzHILWuqdLm9VidBRs1q7n4iXf0s1FKv/wuTMW0uCX56wB8y
1DiPqVDNZWHiavYpB0FsH6bwyxC6dMOTikB+rbvscEmwhAs9AF3W1nxBZyfkznzk
9maTpGROoFSCGNuOY62WhwOsK3V4wqPfItE1DmxwMqzXbdu+R+9T94rsAfhxhn0L
IU+xuER+GcL5yuuvKepCCDQCY3dg+l/YHFDTlTnmVjFDcJDMcjL11XUVgeGI2M4L
6OUQCt9ioTaFgTXQ59zq6P7fAfIk/FdMNsQLd8EbEpCJh7tA0KUQNQrwKGM8hzRq
ffKodgRLk+aXobIY4EDg0/UGck763cAPxuzZChEzjTjRVz6i06fCCw2zcs6SAG2P
ijgSAOsPmZ0GCOrcLlO6cdapW5iWslbxvpvbqtUUlosw8Hyde6PQ0b1huYWCkfoB
UqA0CMXE1lGVdOR/QsNsWGFkjOG7ylVLkULLCzzNLo2cGsmoiT8/6D6PtlsT44fw
xEDC9j1TYvDcu1lxlFDB4Ks/RghXyq5Xl8vobyUmtZhjX+5W1L2y2CrF9IXzlI/J
GLkT12lYswt2OA9d9Wvz6HAbLPFH794vmkp6WvT4dAdCqpVgRPyczacF5NhaufEF
Io11IBwiWZVxsNwwuHn4uMveaU7UUnynIOyyYpjFSFH5BEkvgdgiWjEHf1RRfg5H
wuz2hGWWSZ9Mf/9YsSiHFySYc7e+QOMQuPejTu4ePgzgsFcZb7kX298WsykS4ke/
1+UsmTEAQfCCZ1OIPVZiTeGY9dROlg27cmxZr7ilWyAPQ+izCnZGZ8pYujp1cNxL
PyEbXcplDnSex0v6tWBCUeTWe9JxgXwKJMlMj3apa+cPFPXVGMStHYVWeY/Mr+EH
/j/gLl8XmlYM+PCIm7MTXd8a2HCP053PVa3mv/B7tVDxK/NIiqWCCelf2dHBCFX4
yJMJmBCAKcP/IIMLXUpCqPFgi3RXbAVKB/zWDPueqNJ8J/o0HZF88r7OzcCdPy31
UaIGsi1VRt3fyb28VX2ZT4fqHMoK8h3IMc84/Flpckq549JVNJHuA6RTKlYGzjed
DBvLYJjr+qQDX4zlBt++/T+bPo71Ofa/wV8pilG7YdvxqvZC9dvnhBD0pwaybY93
IQ//L67mnmX/tsQlxwrqRdrr8HukS8AHm+qcTXU+lyzpxm6yUuR8ztgpntLPRlU6
OgTJGhBKMriMRYPGUEz3qXhGVue2hvSe1hXpMN77cwaKp24Agl5cpO0feOBClTWY
wPHReK57jZxtkpoHxigGONaTFd/A3ZjI9zO/BmtoeZ9mTk3PdbaQ+WQwfABb6oWf
9gFs0D/IwuaoZn6h9mTS6PU0Fx9AMqzNOGLCQT8W+SHy2Bu5dFNfdPHDOzc0kdJg
1+QjMdNCY9RyTb0jrhNrx2oRy8faWSxFlBTKKxVfnMQ7SIU4WI9qv86UT66DJc6r
qemX6Ts8NfCsQOBx+1yqA5pK69PT3XfB3se5idpAggOIWPwnR2Sty9pOfhOYtTNe
7bjqWcAkyCJs9qQMs8uypVa6vn33OxYMyqya+u4BhADrDBUeDo7wbqima8vbz528
F7EXNcmZwblE7bv3iU1ifA4znHUzuhf+7go2thZxyzhQBUqb3OOgc+P+6AOPfhXj
rUyNWLGNVgNmHeTsvBrXLBZN5jBvFb+7LJDKJt3icuHtA4OwWyp1H+T0XiHpAiJ/
vipm2jb9jgsZ/Ptix0WHXB0Hq7Tvd8ZFfzt/ur25SgmsXVbBOPsvvArsZZyXaalv
wv8YzOvmzejJJwUwLk21obMmY7ZPsRo3B/yhbojKySIyO1PR/hRT60GPQyWO61wT
zHRsIN8r3g8rsji/sfGf2oejdKh/GPkfyk6aDEwmj6W+98idNrcsaIsAC6h/iigO
Xg+Os+ku0cljWuwOCbSFmmV8fzA8wEQlUAAzoZ+9Lm+aQWaajeo+lJlu8xjjtRuc
oov3qoCqrn5ACB0686eeSEtyWRS1WyefWSWwYLv1KFEolHK/KKPPtsHFCJWEYpkj
6u7XNWzh2SSh0TzdY1ky7yl0E0xORmeheArFT65EALs54Jvz5KTI8M6VD+d4WXHi
vYpdg/57+dscQjpkPMP0qKTUkWXl3H8parwErYZSl15xUwNGGVyxpTtL+zmlDpGK
295aiaBYGU13MM2DHmmwtwC2doSnD0UhiRSB5gEdg1Eu9mnYYog9iUHJbRYlvFeh
rPtaNeoHf9Rirg26sq8hRKtnLcKliBupcTH/La4lZ1o5zuPJJ8aG4JYhMZUgQp09
1SOFW+v1K5qDUoj3AEaVFcSX39je3WX9fNfvnx8LtqGiqptUZBkOp+deTI73otTo
yFDjXpxQglG29o7MCFQzPylOLUFC4BHLeQNEPkqW+STFc/dcjuu6rwgtJQDwpald
vcKRaKIliMcA7CnxQJT1JlzsOp6XTxTtAfvykDh5PE5CAYzvaQnV0JrfIXWUG4at
CqOxO5KqWNhqSNxGt9UuDsFNC8tx5JYHggzwDF5C+6dgndjud73EIij4EiDuVpIf
AYSGnUAN871L4uRIKuzZxOChtmEa3JN2ocPvNFPITh0hfyOb+EvmViJythCJgNps
MoyGt+TFlXcAZ2GkQ2R07k/DI5BQ9mOdTIV8dgDzk4kHgO2yD/F8CvFfhLn15G5P
gQvprvHoAjGAcr1v0foj9lxu3vi0w2Q8n4+6Zvcyoi8n4YfNa5clqJ6pkbX9qyfW
W91VA5VMdnH5hZSFFCc51oGkBa+LF4gvF29v+vUt71sBPHRJz026EACIHOw+IYF/
Rt4fRfgpTP002bEQ7aMkx551dWnEp1GJsB75114YqQfHDqeD44LjU3YxFQGDk3Y1
nrW3uK5yAkgzSP5AnhbXyUF1JKpx0ffo9eulYFBYoDG7y5DSyqiUP0bs4BXMaIGC
KZ7uzrNNpkVwliD548VlGLaHFgYYsh2q3vAAzdWxDZCiKQopTR4iLrOJG7iw582l
ZysVK+X8rM5mXhVcEl2Acvvyma1jNhQygOejQy/QSltOQsJQfXFaEGuY8rWdmBDQ
5IlyqWH/i5X9lOhKmgADOexp9kXNRE4yWdG2YAurQcwVKvYoddCfCbgjfYgCIU71
FnI/jNkGBcLKTKotIvA3rkX+yKMMLsiF87M5hVpx5hKoYLPJIAgKgosfzdkwJF8m
PxZMEQsxNZRbchEwefySZtMaPCL5vxehnZzLBjPHiMXSJ4yeGWHjfLZqKfYbLIvv
NR+n9S6HXZMi3z2H0gYYblso+aWjnTV2NTHQVNwGwYlIqDbdH/6yZVNMtc/TYaA2
4uCcpN62zVjnGVTCiF+zovc0d2TFb06xKMkCTNivnn2pI4C/yMKfoANQlQhZ4/6a
yKF4ThxiBHaT5U1n/eA7R0Rktxjo3L2MSiomOJDhTK6vVn1B/r+M37TJmyHif81x
5CVjssYmyX4c9AsnuUtmJT91BaU+iMXThf2UWbv8ugmJvP4U+B/hSI3ILjS7JsGO
1Wa/HQMQ3bZVOcFL9qFU57LKJzGvS55lPZ/QWTjwrJokVFJo6lo4ucSCX0lcGTRB
5ZpBZliJBXa2C3njpWCcG3O4/0HmTu+GvnEPqnbb/aC/NJZOdG+2o2UobEp9WwRY
t9ddKs8RTh6sBOXjgw0ES+YoA9UE2gF/tP8RwMqq7s9EsRT+cS3WT0fSs+5+SoWb
BS9s1t0UBNPhzjxYpZPt3GHXXYtBYusy3EnQESWc3MhA0i0kb0gwsV6HdAZzbcjL
FwMx665OacxvKQ6emUF3CMAvl/tKs1yOz1AV1iY/gb0pCil/Z7MtLp5nxowLZZsj
ZRrR1fg0xj4YQcDyHSVFqKi2dOTTglcOoCLprhSsE4qa6n2DEfLeldYGJLFj23n9
/z91KORp1Ven+6gq5YUYmCwD/lRpONkI3q2Qq4P616R3NH/kpG2uFnJ3gg+gxWrF
58l/ov4KK9OOUoyMQ0uUxE879HwklgTo2z3QwP6Oz3EfJDXhIPEvh5QwSm0OEOVL
9Vx9iUMtvBoYm928Xve/itxycmDpCU9TXUEhb1IJJpJHxLKNqa4WQkOiev7eqpLc
4AourZWggZzFgmxopwEseksEssZ9of2b9vY6wOAZEUf7RCsrFcnqZkf+PJuZdjRo
yXXHDgdREh1xRbuT0+5B9xGuC8w9ju2jbVWhwBhY8iBmz5HGR5asvc0Tj4TRgj3G
IRrWisCWNnd1vIlzfmhVGaNJFVYOGDwL8CCkOaN2NBALiubPTa7kbceTRlYcpwwK
WsJWYHnw0bPxvqP1i5oovs6k6lM0nUJTNHEQk8p1M4xpUTPafsEfB+8Ju9fiBp9f
kqnRKCaYBhA27GsguEpnY7YrNVBKQXxqlTi2MMDA2mEt6i54wI86FStlXEfTciYD
lU9gskCdyWon2q/Q8yeoTAVmFqUNtRemw6beUoX6PgSgCHhAPlKhpGar7ZFxf65R
jJclH0wUHnnFDE9P4Dt+1h5ixAMzm/Qa89CCJHnLPDdnWP9FZV3818NoO3DRRBQQ
igmGNkkS4HhTipBlzGvP2QCU7kGABVO1Ob6p58ktowMlmrxO8JlSVdPD7k70Tob4
VAYZjOwZQlthq50JU4Aski44sXUGb3ePdTjHzE/NH6m6tTyj9wk5oKT+o2hhX8gJ
Sl2D+NmtODlZz1jTMxA/PDqOmq5+gFr/Aynk9Gh3fWWU0pLVfFEuCy0JyTX/5lp3
/DgwLBvhG2Z4UuY7bqag88++LuPUNNNM07gVkhSE9j3qOkP0l8XSqttbLdus7p+D
x9r69Cmw2D8F3QOMrz7EMDXwAJow3pLoXDvc6l10xFKlACeSY1GlyCxp3X337De3
DiUxsdymnzJ82xPm9c6bmvhPfjfMX1PV2zUTHx6t9GFm3Zq9MIq+78D6v2j5F5pF
P+CpRneE2i8SFZEuGknLDCB7avQKh1WRlVG+QOPOwjqK18R/y9awcRO7I7ZJT/y7
jyusg+e6LCsVUS11sBXGGCyqmrdxbmUiLmZpYclD41NPqUSYzehtSe6BSIqbYejL
yLj4T79OFpriwdE8B9uSNTbIOOt1nhCbj6vRHjS1NKPzFZ7N3P+CvlZfSGoKGYRW
L2Rp8ze6IyieSKeNgFrTUO9MuURIMJb7wWCsM5Wni3ng2nDbj4NiSp4Vm1ejZ03L
mJZDRBEGc00LcOeNN93UEa5nl9B9/g/PKth1hn/fG+SdbG0DV3GDhwDwTI47pq2t
cQUWmTu8qhmhOmcAol3D4RDHqpyzS9p43b3BDcljxKhoYinAc3udPQQ92yy7RNvl
Nx+52N1ePqwGzth+SMoab2jZl6ThPXdZYVzZXBJ513GXVn0lsHaJjeyCk+yL2Iws
GUuCsqcpLXv0N5D9uO4fzE08+ws4az0HnoHjeiF7mwrEYIvVvpoKFZ+rw8kxxpYS
vx2OU2EjTPChlKe3VXTiCwUDiSV8VAiHGRLACkA/xZemosIIbSXxMak2bbKEkOsX
t27EjPkmOo9u6OEIpy0SSZp/ZQdxHz63CFTU/Ki6xu3kxwzi0anu2dTYYeZllX+x
9rha/R5+sagu4MkTsYl0VytRDR3h5i7BGHyVyoBbIgHSBwoEInBvYPXX/Vtr9X8Z
XgOvBg8I/Z1wsdZk3YX1JIWrcoSO+FzFIc7BJ3hqI8TU+s1ibCadbJosIrBFqTNq
VWvlERJfuPlkN7WvZsRcrD4Ioo51nFLWwfggygNxHzqYqMJg6TRwjxsjkNov18Qm
ZZx661bn0/KIkucTSsBBWLM27TxXx79eQBvx9hnELTCuXz4D7lbUEtbnYgaLpR08
I2/g3N1VwKA98tiv6abOceFGZx/TmLdLmFZLyHyd6qHSH2wR/7jje5ppZV5LOhiA
+v+lTYiqW0V9qYIFiEe2j8Sts0zPbkj3ssWQQj9KeJ1Jl9GRZnDPp3LRJvGHyJWI
Po9eR088EGVSb5Sn9/WQwlNR2KNOCsCiFW+sPXpxbbz+NZ0i6YqqjM8uBVrtEPdG
bG3dOQ/GH38IptN1jkX/r9f8MlXB/pgIO+CnaKDBoDH2igh/1cvslLLwOjpzgkEi
reunY3/y2na1fStAAiuoZBvKJ2ULesiRDKJTpSaUU3mCVrg5wYN1hR+h2cNGWBbJ
XBzuxoQBT6Hpt5bc/9dadriz4OtuFp0dTOnY5wJUH3PQBlkfXdn9e+9BWp5MNSJw
rVm5bVG/ZRw64PFC6cukAf4K7Xg9GxUsab3tCGRalRQ3XPTvnUD894Sf4FWVoft4
hOj3YP14KT6ZqC8j8To63bqOI2/I60xFi+Z2eCDHFIdRL7Cz4eA59gwrM5CLdCPR
BMoTab4t1DMAqXJ5ktE3nDk7ahUQGmWQNSmvlRYV3wUUSLvVLVVYNf6uA+WsBUFD
/jca2eruKee8Mah8Xa4T3QZQqTXQ1qO8uDpcpjnFXCDhQ+Gydi/flrlejSK99sf9
uTixz91Pw2KLM7sQCEq/Hvars1k3DInV3mkDjHuhDnV0KjxPr2ZVsyoqQ/Bp9PCc
VyVt4iUypcuyeClnRuawTVe79iCPztPj608rMde3m6ar8P8712GPKazBgG5fLcIf
7M05UpATlS7K5GpKMsVPtdtSSucJ244V8GBTOEf0GU6yVY0pfZFuc7iHLt0l5smy
3f+NIfvOCLEnJoYJlUQWKr6kFWjCw4YqeM0tl4zds0J6Pog18R/znJM2O0zn/cCz
QUxdngM8DNFtgFBhv2NyV/mOBA47B3sRyn23+ePkj5iW9do1z5tEp+pWX+Iwom1Z
9A+DEEJRAHC2QT52qEmrDninyOzMAGmY3Nt/us04RhTLYoz8oB/hYDnfuPyCF9ZS
j5n/wNfYo9j7vWaPCBTnwmAyymwC+QiuL+3dhLkTrhl19028DR2qM5A/V99SnFNE
JSNBi2dV24GhSqn4mf2FTwVCAGjF+Wa80G0oXaMOqogTVa3IUHpsUKEfDZeZNke4
WV+SamLesrYxbRT74qXorUfiqGZxklqtx752Tvstoem3OfD2FW8FyFZ65lD6fUXz
y/ln63bsW4puUNmGH6eNsP8hprg+0r84dt521qDHvru1t3O0GMORJ8yWf0Fefhr5
1AWjkucOSWFGx3sbSnE1BSsN7bf0FOkNFW9kt58d/SfY5iHtZFhO23dUr9+czGRu
FpvnzQ+uA5hY51ssX8wVHH0u+g/WBs22UfrmEJoz+INFuvmqQh0+q4zGfoIPrzen
gNCY7dNVJ2zhK5TtZLbMQo/Jtuha11E8Q7TaQaOZjopBAEYh6YsFmY4xkTICT0/V
dxidsGf8yVU97HZTMh38Rv1xT08dvY+JSFgj++5nl8GYHB3xMg7Hw7/eWBPQYQos
uAsZ2kwkKsil5eAxc6Cmsg49K26CYFCkqNLc7WvV9Kcc3Q6/bTR5iFcrxhiEcFq/
0G0dTFdMQVmDXXWVeoEoSlMjYbDRIcL6FpByOFbkPej46DdtZsSLuaJsY4psmFCy
pqVP9zWXyivbvoj0XZE/crLQmJvCD2RqjfwlBbK2P8O/07A9ggkgdAvmSYEwYZgV
4XMx6Y/e8e/w5QqO//fFSS13PzNek/LiH1mvfKVYsAj6ughRl3q9bu4N4BNuu14A
QWuR8/34WXNK870VwzPxkrKCahYNELnMBDHdOPU1xPSuX5YUlGlqOU+s2K2L6oyZ
Cgr3mF1De0zQ7B2BgVV5iHxRkb6EZVrPUanN91cKHD5LS1AWxkK4Sm+JGVZ32m9a
8DyB053h7CPgqlLmnoNX75w+WOqPM3LxfO6X9pRXEC06743uTZrrga7lHmOCLgX9
DMhseOYDJxC7BtejG9yTB6SCC4ISDX68hM3zYkv3thCtVr97JWi56/mbmCqMz8OK
d/NpzEvWEdKZ849VAqwwkRifg4AfR/S7VV0QksEylsMEs0rmcuzqz2YGQrVfTUzD
6NCGKDOm3pdmNeaAnQCZhimhc6G6c+a/T1aHjs2TtfVIXlwsi65+xJCMkJHLFu9n
hwwVM6ssIWNDxJCE4W2Vx0/iJicJ8RCb+y0varCAqBeWZ+jUhZHxLHrjMCggGTyJ
Y0ApA4NqnPDvmFBznS9iGRAPswbfH6JOMLdsnwjUMgFVSR+u1dioMJKSlK4GwAl1
nsoeUQKGLezu/pO2p1GO2rKaD/GU17T35ct8G0tmw4NnES8PioHWKb9lpdT4Z0T4
Q0uLqxxCLWP9aCvt8cbSPs/lBg7pCZGnBL3sYQaqZErUrYiB6ijNfCzJ4lTx5SBi
xZt48qgyr/7bd7p1qK+CuYG/1lyrxd53sEwBCAWRBdqQMfzg472KeD8MCjh8vFwH
wci7M6w01V7ymKV88XLxKD7YRNjTLXtC31qQhnRY8onus/q+Dt2i/x5fFadSvI8h
LXIJbeQJ4jT/uPiV5GF7LdQOZGm6LSZGAmUhZviOQ9Gy1TkZExZMViFnH208V8/i
35+nlzvF9OPRIoIRUCXL/qZZSfeJPfhkFRCCtzy7H+K1jUfZI8A+N4E5f4Fd0oXS
EUZUsoJJ/ezSo8DY2ups9JkX0SJkQlZBm5TcAF9tfNMHk+ikLlpnCjChqJHzCdMU
2RO+BQuwRfqZ2R2KOLk0jla75V8loCN6wJKdlA3lswR9AQRDvJhNDuXP9M1Bcwt8
v7GQanu6K0c4vi89XAO1jRhZCW5SapoNvBaA6MfCxTP+p12RsoHP1SO9P4j/r+VY
abwCqZcoWrVssEyYwjRHdew4sSDF2ttnX6EtB6Vl87oyYBIZ68lwjsPYvL4Hg+zO
EReXBqQEM6TFvvJ859QASAcb8eiMdb+1+zUkigkpGUXtWbKN6MCFINJXRaOMBxNf
Srl/eWD+WvU0bkRW7XGlDZ+7q/xZuvZ2e6NxW8diB/WCM233cXJdHYFPnm8io/db
Q83ldHy1hR9HiZnBSEyUEBlHG8wz3UqzG/AGpX5KXBenBwNe9hW79t8KXAi4hBC7
gwJdSN3YRNYlBzbyt+4T3B1/uuaa/5NJ9WTXbl8SO9+EXzxl/mIo6dVpDBmOYZCz
rV3yawtp8PnxjkF+lx9sxiDL/fdBf7SSrFGx+yU0V7AA8mRO+e7t7ai0HgHJeXc5
AlQdFqHh7c0y5gnWEMX18x54pI3JajsBicI1/DTnSMBFURlYA2WYBgAFwgJTFavP
aHHkx6eDiUDxeku6QPoSyE6nWS6fBW6aZGuakcIDOe02DppsGYkR74aBq33ThmWZ
WVyFLGK9Vs/Lxnzov1Pvg+dxY+js04WsX9cCCpih0ZOv1tB8qBTg/owBQbK1UjBj
OqalTLWQsG8ku+cBoBIJk/Hx0rGZ7Bt/BqPA0Y2j8ZKWj/nWLYE0pURDLvyyiIdy
rpvTwcA+/smD0WXot22PRHV/1rEPq+76gP7RG00wAgDwzjAxoCr8JY4lYloMGSa5
hVmQVFhle/buypBu4ZgBLr1MCtgBFd61nvHZMYCx9b12dQa5H7g0NXoVWQhTfyc7
79c5/QCBO6ijiGAE7BVOq4+UdIUF6pjqqxsRV2nzBncvvky/xU6wIyaZh1lqOn2T
yjWsh0jd8N2u2z8/rSBI8dZDDnDyd6zSoAkX0PuAvFuaSaEnBiFOpfIxDbRPHkQP
zvhr1T0k8WpYAcxCF9qNOHg+4DQA8c0vNY6Jr1vi5kwh1NoUN776AGJZk1ycFKf2
lJr2pHYJ++mY4dOkBGZsy9NmI0fgosACbAWRMh7TTUd6L1S4AxxtDIGg7c6XWseP
p9Hh7HPecZ4kR1uQv0tZrPUZNbvJfO2csAyNtrXJN/W2+R7N7HkY+yw5Is//2pGp
+o5+QbJFtSTe3uZpkOg5BAhJOfnEAAtx7yy3h2+J6vHeUL0wacg+MapSD+BTejme
xSCZUscVlhLcfclwaeNp/WwLe3lPy8trlqUQZgCSPAXg2MztL5Ixpl1ytzFOcy6G
OLlsPrkG2KtrZ4DnYjKUM82ElIzfCYtp2dH+7epNUvH53ApsSVLgFo7ooRkuoOG0
qRmMm6gAF0bO3H95ZEHrjYf8/q9Jmhhn5PleoNBjTYsNLTKUICnKdtEoUYRFwbHt
1vcGpHMCVc1WhogyKqj+8fnIuQPFo8WLHjwTUorI4+GBWkwk5rnJwznhh3XAYP7m
IEab+YFGLJ23IruLXpBn4Uoj7+TRNRn9onVzH+fRS1NX0qgdJa751DOrXbjA//1i
F4t7D/zkrgQkFqUVBSKgBMgOyHQHAiUrJTHex3uPTuxga2tLbrNgWRbRHgy4F5ov
34HSTBaaUGbpnJjbYaaogtbhx4qPnTYL8Hwb8unU25Ur4F7hDPeGc6pjHig4yB0N
NPJ+MwnHyoZCyb5/Ie91kIfB4YFMyFbfPsYMeVS0PNi9ppZShyMv6T4lnyZU8vfT
iKOIp9Z5QWJO8ARPtXGrsrX2OcnNQBQlagrMGvZMxWUERFIKVMx9xIYPqT48JXJT
Cb2o5ylMY2M1EbjWWUq2upwWOB/6nsdpbxd0hpOr08MvljjCBoagkwcplqFkslJW
B1eUXmYHoosvGsbJvKpSYxfIp6yoq1+1RezHcP37Rp3pJ8VS1cEPSgkTU4XoxqpK
2/it2tFiVp1+DQ6V3elnJ1lewqyPyMGf0rFiqYMVwkEFzAhpDNm4uf6dnmoqBOZh
oASu3JJEnIPVmbJVGuCJA7AnMqYGiXo9QyAOgHXfZWv/hEYOLo5k7Ar8YEu9RJod
jQUrkyq7e7633NgZqQmhTZ32/Xc1Mn6xPQCpJb2UL70aV5k3a/Yx8JmNH2kxzUOF
dgQMkE9DeszgL2b9+17Hr8f+RCYzuVn3t6EPUrpWW1m1pFjfKVGB7hd17MTKwH7Y
t83N3hI16Y9s+nA4lNkpoOPeVVNCFaGmQMONYmptKfmFGuU2MVRjnwINhsalqpbV
Ow6vu86cRbEXxAVH5h6EVAGHzl9yJpfbCzw60q7mEiCQPINGZJftLQMbeL1MxzYc
7NIw3zjn1y+S18b6JhT7+1K3TDk1mWQ+x5wytwA07MBay16lv/rhITsr+3Xpgm+Z
pN918skQt+KIuBwKk+iytPzJ+fPQpVi6zRbzeadv5NaoPwMxh01uxQ8QcdB8AhGB
sJAF7aFFoooiH5jndg2/ZTMLfqNlxF34e3saGOEvOAznoXogxSd04UtQYfXQqtYH
O1L/l0CNywbTrkdgUdrEBCdwAOkUXBpFJjLh57Kj5v4D/pJmUpi4/qggfS/6bccP
gkRTuXEYL+F7KvYWtefOEXa/n0g/6qntVbGPkojUMfNlBN3wW60H3WUkFGw99Vvu
V+N86ZzKBwSmB/ARN9Q5+jlGqhWwER0Zs2BMxF4o+vboPOIJZxsWqP7duvDftd0H
88d/LE/8x0npwdH9ySGMrpVQtjKF26ahFjRM0qst/FjK0i7U4Mv0QEl+dH9egfs/
UzWK13PKG87E2q6Ha4z14zvUwji88lS0J/iMkJB1LE1KFJMZ8z0PXHsfpjPT4WP3
tSrNM89wGdEUpVyOKSe4wdgMHpSKEsxmLf7j7apHmPNhRQONGzmij6EvtOkJ91m9
ELO4cWWVKzAzgDJGPX2WD+VqJuFcobYdhsF36vpTjGrfFKGBYewgxj9KPkX6PI5Z
2cZqZ/HmojD0ztlPHmo3ZY6yfgmF8AwLc2YcgKTyLcAi7lL+43jlKT4cNAxxQMUJ
Ox2ggmm+vcbS6Fjv+M4FYGjbRiOMoDIIiYqwS78S5KyASWZac4jvxsR2TrUXn96B
Jhr2bNBPdt29HNga9YSudejACtgEqQeK2yO+nhaRhCgL5w7Y4sPYXZl6f/lVJYOp
/i5Ea+W+rdvqltBu3a5Gkx2yEYNtQqQvh8WYRKyEfTYwy6+tZ8Qo+lghePCUwDqy
gXl/5fIB3Fcjs/HbgcNoEHXdfb6BX9ngHkmKpU2o78mQsVWKaKgoz4YBVDvRRa9I
mYMeCvHvEsEsrPJg17iMAypi09bpBZXtH0bOBuDeBIaRyCBP771xliVFBBbHbwIC
ViyQcVh3Bg3ASpKyx492AugXCQy3xzpUfOfHdUsQYXOvggx9uGhfgDvoLWlYJSst
271knrEoPNKJqeNQQo1ofloMrWMBguQ5rPuHD4TJNbDynTJNnsgOzZosdJ3R2tXj
5UOUWfHMPHamyz1ZXVcptYb3aGaCeMmRERCPhZL9IheTmya7n0/XMvTc/fL98OGs
Tj9NMrZFo3iVP7tiaJYpyv+cJhfaTp5NlMNhZNbN/TxbkB54QOwaR6msrwmr8Ch+
Q6kiCOyMYzTy5Zh/d9eQX6csr8ZqPNcm4ZrYJFHF86iojqLnXatkl8esDDmURyw4
lz9KFp3VMlhJis/a2o5eOsP39WfuYaz6rGNfSiGm9Bs+ITbZGxRom/9KCuU8683z
96oJ6E9UWrkVHpqm6twcEeYX3QoJMFAyz+uTzbZB8fsP9kXBlX12r+zeOP9YgUXP
ny2nl7U5/T0xvHpeKcMQnM/cGN1owAvj/xqW+AiCPBOOLxvd1aQ0DJ7dZ/DJwc8j
kkepTbIgAePLeQkPdPkLMrrR/dFSdFaTC+OSs5lYLCdH+7gtxHKGa8MfcdttnJoA
z5MMWwdZv1LIl/PzkKS1a+uvhMrR+jiA9zrm6ERtvPHqY3wcJnGz4R1oS+CQ9niU
pHU5Pdr4QptQF/YbW0G337QoCQJpyiXfke73kUJSikzBl/kf6bgP3aIEswT8APF2
6M8YqJXnu4QBEIlYqxsO7l8W2LFPBsxIps8fK8apcV9TgmEJyKClGGFn1YLpAy0E
ttjrt6as4kbXNXOZDYuP/Aq7603SDtWTX6Crrxj3Kq6qD3afvEQhFV8pwIKG5jzY
aV+ptiGAkE+vFMG+DnR4j3KsY7Qlbwx13R0cTIKOxP82re6H1nAIYsatf8tWBENA
vKS6Q6kALCGi2U0yYDOcq0/eWCa22ATCXLonndyPvT7juVD30XmXErthjx46Chzi
PKvdwiTHxhA4JdsjKuJIwUYHbtuKCuxQYIkuUaV5lEbltTa+M1fkwx63nc8AsNjX
ZImvBZKhj8BYkrvHpnxpGtKq2ti18NFn/LFJZVyiHnjdsaI/JW0wsuRP9PdGNDiF
brZM8do1755iTrRl/bqBTBNL15ZJ/eBz6HVcvzmWbvFtvdo7SFAwFB9MeksGnj9J
3G03Jl3DPWAgXUOCLkk9K82sPNMl1OUKdsdIbHiQWw72bL9fJVuvFQCAxzX2+rPw
aQbqNBedLWSGmO5Su15QFo02Z3lcTXmLVrIaJ8STrG+GevRQQsx6LxBM+gd36OWk
+InMLGAFu4doen1MWvhjayg47QXn7GMTX5iawLcnSgqC3b0fQSXxjrA1FfLgf29p
HnQlqHvPl7aTLDoGb9fMC4ghev6Sgtuecg7W6ghnbYwwOFQBU48hPNgqZE4sS8pW
wPWQ25uepmIRlGgcn5iK5oNz8kZoa9ej4VR2OpwxQIyrKWD5OVzHgPKkAArOEbyp
023qnonLxhZuGDb1U1RIzkdlDyRLtqy7PpIbwUfgotEYGuWv4wEcvKC7BDHce2sC
DLekH6MmSIflnz89DiTES62zmRd31zoxsLBuZNK1S7KIviX59/g37zb9u605qGt/
m9n2g+4JAsGl3H2scDX3Um4BzAGJmgSCzhSog9Rf99MNGnmK+z19jnYR30JOCIZu
FLwsKBfThxgIvnInXpH2VYQCmUSE75/NshyYldLWbB5WuyVto5rrgENQmuS/JNgW
sh7e/xZtGE5nvroxvanZipUlCu46JI2wZF8ZfyaA+LmCAMY0wc17xysaTLz+1Bn7
wb/b2sVsHY+hpUtDeYIc068G6E1c+flkrA0OJZtVlzEV75luaLMDWU9U9ogZ80ih
1He0xApFiX4v22aHrn/ytsGQyD2a3epBUR4A5Z3+tiBbFeBqqbZQiQyxn8lZ6ngP
exfxaU11b6/SZs5uBxmxYhmCdFK0He8LeZ8B82Tmzp/ZqOyILxEEc+l5t3nY7D/8
ITp61zJ/DzlumwRgNmaU1b0ZP3qFcr8Ohpfdmw9IEhRFSV930NcWcLLxQ0N25NzY
My+KIfTGmnbMCNb7060Ac0NHOzme6C9A3yBZfNUSfkxMpRDAp+NgrA874pIBA5xk
FsYkf9lGop58uvYkUUwAbSi32jbEkNsU2NpIfpcmP8P1GDjbxpAOdtM7c0zu1rds
hV/CRJDManVCJlb0eEva9G5AdpJq0M/lrm4RViWQdjjlOeoTdWe9C5uxi6smTMtO
z6Li0/6ttdhyX2ArvtcSZxPhzNKwQIESJdaV0gJO+b4nQmwpoQE/7j786fg7Pz9S
ej/Uj7IiCYubYU2xBiPTYDNrY/0XPO+Vd10PmaZlb6Ht5jbyFBvp9JMPmFwIu1m0
Em7GmTOGKjyq2zEHCOMlwzzHY9Rp7hOBoujo6mQdv/EK4q43WsIvB9LtoM2LP5YD
lBHDQbeHkOEW02YvC0nWsp8nLFXrAer6/mJJycn9lWBOZA93evATUHSrh/iKSnyX
DWCM1nbTfKh8T8kWzaa78BShGMxh0m2vy7g4/ISGpVCZeDFgvLQpXjSTQnKxw3Ww
6vaOq/X0lpZYvcnF+dVBiYJvVINGP9HCptu3ZeJkez/yi4oYkLcESI4UbAO5wY2E
jfmUJPZWGeK3sbjAUySm4HY7B0/BwAsecgkeqgOXLXkVRXrryEQwJ/sMi5VMo3fy
nAzaK5SPNwAq/HrUqlNRk0kL+mMqP2rSfCefwhXFOxHmvyjefyTNwODMT2BE+geZ
PDCovcbIVQfGb2qIFdvXKtsZgZ5gcJG9x1++j04/gJkS7kJ7Mgzyb/N8ZN9QjVM/
tdZ9xk8NKOp6QDRjjzTXUkMYwzSPB30gZA9jngNKRqQBKVEUzpVhPs8Grpafz3tF
nkuMNUy/jI5SVhULFw9WtS0a0VYfo1GSJNRk95JTc4vWZvt/OjDcbyIBLtje31ok
WOHuu8kdorx+NaeQBWboZF3gb3dOQkXqlbmBjM+yb/L6cx66hFwOwiITKLgk9I0I
/a9tg0VkY0LC64AUt72/SIWOu4TEYXVtk0gyDC9sTgj8qfa+APG4iPFUkKDLXk1H
hISUp6/hOvAVe6DZrYsHI2XedHVtKCL7tYd94Hs78qiP4xqFXp8+2GtZqpuBeasc
nzL/nk55Q3UBf+HgL1cX5dlzuz52/6WWGgfXhcS5csRpuGtJLrRToopPT0aUebHc
gmwUyboNnr2XUFbYgcsFb6+EtIdKwargI085N9oxpHfDP5LYcrDT0gpZ9xkF8HfD
vaIa/zX+1/cazwCPH29s7W3LQnyuQV4kGVgQOH8KwDBOFKDVkhPA6u0Tr8d7dOaA
hXLanqaOSOL+H8+e6X5QmUvlxQTRu9bQwFpzw44irVKFUDbYsshBpqiFefiq6sjs
2Fo2VADRAU9DVzXdmQAPdrgkZJ6NMjOHUyioXb6ntSOUCuvliFuR4n86frWtHuFc
/4uulCdR0ceMf+etbYMps+j02OFsy7G9knGPX9xhQw3SMbh3A/lu7UoLRqKLmiaX
esI7ZTroSo79gSxrlpZUPZ81IpOtsQ3th5zjgTjTkKgHOscrw6C+5Rx9hD5lntHT
MEHzWywLP3Z+3QDz4auYRpYOhPLTgvoYlf6cm671B99coNcWB5VY8nXm0/b1mib8
K2KeHx85plGnfaQ1JiAgpywEr40aYlJmTFVrmMh2bWuok8n8f6dlgkl4gRkhOFYT
N1IhF181fQ8LCSSKLqS23sgubfHurXEckEoRwgnmjAfVAH7EelDmiHK/EBX2kU4W
tBasZFw3jdTqpFesCtyeIxPDrrADjlNell/mdcsJTL7KQMAxTDL9ZRCHbJuuVaoP
amxk6f+i9IXPeEL+GHiEdaOq1npNM9B2+H7uI1EdkaGaeGXxYal0lEtd/lhYVPC1
yQauf0pVIXhFjZIcnbo1966/w/g5Ov4dldSsTuh9B4BtJQXdwCH8z9kaD+3wbfwG
rIe87mb85PVXo4F8j6FN49XBS8X7Ul7LpHFgdxWwMvc8T5hQPPSPyii/uVuwfQoU
9bRecVfp+gCPAGp91QOvG7C6IEw3ncUmEeCkQ9u2+hqIh3RBxBf9OkZck1SInlaw
0ClNlReFt9Np3U9BowZCtyCmRIfir02bq/nvrOzr5nyOu/OJjfAclVGs6wq15hMW
aC0tQDryFvnp47VL3Fm4ATn/0puKtjk8ZHyj37ANe1+1mXjXY7SsmIjQctyMDr5h
gdkKXqCmUtECH8EKF1HDh3M7zXwCYlDkvWyOa4YwJ6aUOmk8FWxvNiRLZgCOFH5n
DueCuIOG/d6zKSSNFd540DfzrpnJjdtSXEmMCBqAyIAQx3RKMmJhjQeWT+VrclBs
zP6z7WPICSQuQi89UkTIYdhsRUz44TJoKh8hp1Y8hi0M13fdY2mKQETdi9aR48Ls
o//SphyiqlL2uki09g2J1OuEBqB1Ls5jdrMEilpzMHTdO7Y8FS+2dxCjeEkGiS+H
10pPi2exb2JwWhpfMMivPEf0mqxXrD4DjSUXD1IDvlkGX+XNrjTCaSxsy94do1r4
gZIZL1z0FGr7EFz5f3lxxDuw8253SfuJXWiM3XjQ7AVDLwtrNJMxN78mjBGKUleu
GALZ8gOqM/DEhKY3lQkicK7EV8vES03qbZQfgLrn7qCKPzJA1V7gVLnVuOasSMc6
NrkXkPE2lo4dHFvX3fO0ctrCBY8gZJbX0ywkrYGh/YqNIoTkJIYigXLXDMFaPG3m
jBwKrtmwg4PUbbhAjYEkZQtpju1fbft0N1Wnx/baXDm4Lxm8fui8I3/+I9bnCj4i
5jodrFgmUgtXaC++I7NTRzx4JrMtAV8HJBssZS/jEl/VcFfgH5JYBOIdSeVh9qtZ
AOo3HTWGdlO+3dVoTwcxhaX2GtvW8ymN7FPshXsGtU1iImfwP/9b4JeVM06KYggM
koQS+aKAUzWHH+TzxVULbLRyvw5MiiQLCGyVOHXD+WKERuNJHa9TnRGOGwRGf1g0
Vx/JhxZViaM4s4sa2i/GME0RyEiyUQaAeBXWWAATdEbMniB45jmHQ+DAPcZjIgJ7
IemANZgWDJElV3xJ5+mx9CVQm8ojsBN/5loTLffmfCKUmg5ugwkAQav147fBZV6V
fHE+QUYAYYzYeWIxNLB92FP7ucWjnZxfXnnPnb9qVU1Uj+kp5LPC2ObHMXSqvH/5
sTy1SOnW58QBV8umnurWOdQ223oqihtZ34KA63izu2RnIVxc+cL0PyGL0iEQGe0U
2ebTxfeOGZHPb4o6pricuY4CyZcfWx8gWv4gbI2rauVx6sqA/aOQGcNoXOO5Ii7u
m033G0a2NnaN2BLe0CbyzpD4t+KXqfKMan4CB91NoqxVlNHj6N0e2AaCc2QjOTXH
E3PbCnYb9l8Dv2cUHDsX8KbwOTMNG6gX5Cru9fDFW//sUp/jg6M2HxXs191xyzDB
4IoIuyQ309uaYA/+5eoEHo3boN4W0uWti/3HG/1ExOreC+0heIZ3x9JovwQMGOxo
z6LupoZVEeRhVjtgdKEiy7I5KLNhoe+z5BDF+RVtYpHHBO9N3ChsaYj/B1krt2YO
HZJUnMl7kgmcPtl1/YxQrYRRK0vFud9EwtCsHHL6E6BPwQXUQmkDFY79Kjud5U9U
CbDAcQcQo4tS6yEx985jBN3ALif1oHN1t1ldHw6BjmfMri07tQ22L67hRQHOsP1h
pa7D0DXeupAs6gkRvqlhqKMrPr8Y8BZZxqs0hDjF6AYpoLeSDCRBUjKRVi7cvaFU
Z+AoNmWRAO2+Y50QUlzexR30PEsomo22T05K03NVAnz3ke/rMOdLJ8tgXfoTbxH6
HBRDJay4trLFEFmcGQ9cmkgvOAMQQasqg1V4WbDNVSeIRXfh4rIHFRzDxqeu7wiZ
emmhjSbP+18XYiMDpzoXF7RAvOglNp67KDbJckTWphaL5ZlAQSTHMUuEmfeAA7aP
v6Sc3Xb5FiZA4JTEv/Ss7rFf0fpylfRfd1wd7/7hS17rEs+B5aa0qhBLxUeiftxp
tjtRMX4ZLSsK2bOqJhCLUOsk4Y4ARvfmY5bMdcCL1dtEW7Szp8xOEiciZHKNg9pW
tDm86iimbo75g0IV6S7j5MCvenWCMNqWQeJ01oC5nM8tH/YG0AnKeRe3RcoQWm3P
YbGw9TqwmOgjzG/bNM+mG8sLVgwKXzqdmHEHzLEzdAyeqZv7W/BLjsGp2ZjT0GuT
5ehApo2CDVDBLzhjFJ/4bmZAX7C/RAxhF/FnP7l4C1J7JH0a6+fT3kixhM5ZIhSS
oM3mj+iV39kwCZxybcjOtvmrhj2cdEE7IIipvIItpdE3ReHyEy091WfgRTIl3TJF
PhZW8UEONqLs5I88qNkpZcNE1Ncm0yUlpC4GYOglTB6KWGDN0pJYrEfnBG7H3WWS
3c10VgMWcsHx1FrQBm9Xr9tHfMxL2Q7Ec4+38+ieEmPsMkOGpdeJVoleFHCja5Yw
Imq0AkoyAxdtGhMVQMgB/y3Xf+PYM1VBqyoQS1ePdmCXeh5YCCTbqIqQ8Ku4MeSj
BavKccI65K89Tl+KjgNv23hSKc8PMOmMORWMu2hNbagp5nqdrijmG82BXlcQGfzL
ysyn+Q3aElA4mEMo6gHXnGUcQviCaCa/PVJ7pl6IHsXTnWo4q7gVw88jZtnV0vvI
GZLPzWY80CK5jQm7GExuYKI235vJALESfunQm//4jglqMqU81HX5GVEjfuQe2tBl
Kn/63SFRJKJHpyo33J6MUX9+8y+QuOVQURLU3P66lPwTOmf+uww2ryVIC3KvYM1Q
H1gZdVCv0FKEnGCaQPIIuXviZH4kerzNSu29OTCfPmENo6NWV550p6gIazxM/Fv8
bFjnZMvDmJUQRtZRhWjiF8fdPNW+Xxitr7qXAv/CCUuJXA55/bxB4KczbzoX6vrt
TwlP3yIIqtZ4TqUdy+cY3NzbCiHHSTn/irzbO/5LIgsHouKZdf/7Z6LKg8lcJvcU
iSt2a8SNjDCZ2N7YDR5Okj5k2FFOpJQ/ryq7J9tdNNnMJ8X4v3WZhuDV9mHvY09p
rOKL5OF2UDASWaib1xlhak6/p1EvhYOsUq5YF2y8WAGnxS1tfNBOR00ORwRSbh8X
owrGRq3NNHVnkm0iuAY2uT3fAQTuFtmLMuk587Tm9WuChztpw34/0+Mm2/CGAKse
sMNJwQh4VSrvSakZdhWqhlEYzQGKpw1aF1qCuecOifTGQR7730PbgLRA/qgt7swO
TJQnLyEcwmi3ovvptJTzP4EtTNoFYtDhykA9QSidfFfNdmODC0tShXiiRTehQxlM
jy7wK5OcgittL3Xs8jMXe2NEGhpG1iD8i6Cjup1VtOppWYvFqosAB1EmT6PXthcn
XufGoBtjM0x5mj1Q9BsE0QLyzYZxoEW9otCwmisi3LpIvqfsktC4xwvlXt496hIr
4XXi7M3SRblLb1y16kxxgoHz9x/BZZacKEbm6Atb8z/eX7nVXHHhEWGpH5xhruGd
de6eQwItxFdqwWT8RDvHDWiZNEj5VeBW09ssoVbKWW8oi9LPFQ9KllMCyiPMQdYh
UW98VoO1XxX1js2bdU1AzRPT3gJGiKy7f80Avd6xtt9vj2hEfhGOObM4T79I7AvK
UNBMNDGjDqVm0O6imFQWEU+BCbGxj35oOExuvkHbCuDW/kE8dDhkw2LHwdjAhakJ
+Rr3xXIC/hsz54rocQmUJMmMlFkCSfgMApSuCemAooQ=
`protect END_PROTECTED
