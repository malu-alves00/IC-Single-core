`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
elSEcIUnUTDyWUG/pkKikn3PRlzkk04CHrul2Mm4acP+h3rEItC4x0fYcEURERnC
ouOTZSwJ/U4YfTUcI1LCIjVlf5Yj1Mg7VINGURXD7UvRVBqpow1sE2nBMx9wjt/5
Ew1fDdN3CgMpDk+XculG7alsv9HqPQNDVVMecsvHH2DpFugyGkbuQO01nPymtWkn
Vj0nUIc7CnkHhuK6RDqD4HQyYLgn/DROoSYX2odQ3rI5GIP6vtHAMT0lw8vCaJo6
M5qNaLxtJq/GLl1QuS5nZMadCvPLieme68KgboUXW4OSoDwZJPwYiHVjvFU6gi5k
6OiciAX5WDggvFKn4If5vhx8WbEWE4K9FP2W4SAVbakrtLa4MiaIQ6b+uy2EVTVO
qakhsTOEN1XWoH4N/93TBnf9PmSiN/qM18SF//kkD0iVKYwcTZGiAS5hBCRtmSbU
E9dEHrzQAVmCCmwl635xU/73pitPbTygmYb+TQ8T7SztavkDDPPUN3Lg3hdi7RSC
WEJ11aG9qu/BtXvrwBrxQD83QJ0Z7bwpdwFd33rE0VW+4ppeCX6fgvXlrve4W37m
6H1w/BL1JC8Eoqpdew0Fe7D8IbDBXAsz+iprh2D3sOOFL5A+hDJmznf/kFX92WLF
rTMvNjXEqgHVTeukgpnDr1lLkIgJipeY9N37CkD3+PTfQnEr+TkEtlM/ZydTBe5a
efLVmnYDpbJWOgIqf6x2K/s9Z6b5Thmc/YLQV/XlvI4fHtzC6kjiLVhMBaXyMIdi
Xl8secq60XMWetEpvTldjPmAbARUKDn0XW+SAQpMgiodkOFN9u4xpijgZqLavwg3
`protect END_PROTECTED
