`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eg8CWyTN2QHccorsF7oyEGO0QHbYwEGV3Jaf+DRi/xmBiW7fQLG2TxoIDKDYdCWd
Gw3CVmXE56iqFUULOcsdv4/LSg+a6ceHwf8fDalr/f6ok85pVpLGPDvNkkMhOc81
dyvOrRDAidk1ZG49BEb9ASY23zNPmLIh8o/H+Kiqlxa2Z6nD3oVkLY0LGlMCBAJQ
3lNlnqLIpC7PKVwTsaCegm04+hvMfG4AZyoF0vNX3QS5n6o2NCujYqxrn4yvUsJa
4vZ6UVUlv94Yg3ste3w3ZA2CQkhGcQvtT1pzKruxniAxlK4zp0eVfLTY6K7ePkdC
pMe8tKrJKAdKlhR8Loz88rx0cFQNH+D3VfiWgi6vI0K5RI42I1VKskZFH6HFUWKf
jkRZok2Hl1/Kqv2RfAessbOqMko+Gccfcju11+HJROC9IUKRHwcEVnKNV+ZxEFHO
d0IMdww5MQ5r3Ode2FlP/sigirpGn59Xjw+TA9VjSHL2Jv2r6Lb8j+8TWoxQjjDY
HYkPBwRI1APHXXEu8aC51vwZRH88guOF3EvX9Ahzjp+DaeU7FCcwgb5D3i6pKdem
XeE7JWt8OZnvdFL8zmHBet13tVeKh5E5y4/DYv2FdnZpnbKH8OF+YSqXJjH0csFH
bHJ703AJjNz+rO51FPvoO5yu/bQsm4dRjvM/e9OuFLoOx7fPujqhSstsCWpHEt/k
6hbxNAQN9+vo3WevFqsomAQUfbBduhudmCwz9DO5Bf8rHaCrNXBQvzYY8AawV43B
zqSJxBYvEfHl6WcGmLNhGK8dvBgr30m8s5+ebca3nYJwji5OOVZgjgvURNPXcIU5
0u5I6qeFAscoTAUP7ZiWC+8lHVQkocXwTo9gKC5sUV+xENpvrIwQYHIxe8NL9C6h
uvPjyGJduedOc7Td5CoSTzb57rm0VEvQVN7HhM3fUoYBa6HmZdv2PnitgaCHZ0ny
Pgz9KdNtoY9wxhYyEZOClZER37vE+tqRsl8AZ1Z73Nbc8Y2wBFDwpi1RTuTc+tn8
4xUupzXq1YoRqkwiCMZKlJbtWBdWcKEkBhevtymtdjc+/pw1QvwUEcJaNDOIYktF
dCLriUNqQbr7W2O43x3YU2MD1YNtpWikrf6mowBAqSeYeHAh8n2as7DK5ZVJLomp
L68iYxQoP006k/cZTBotz8zZ+0h2tauE8hviE+fFmWPYni05YrJv1vNu+jZaWuTF
4vLD/FLRt6YZwWAeGj+5QFKUAnPUjqX7vJmtkIKvXeqlo8QQXoelSL6WFRmmy2cL
jbPX+voRfcu3B5BttC3uIqGKMW/xwAk/AASfDh00LH1A3an1xWa9QY2rEh3qnzl5
dyGS7lFoiegEQK0E9dYJ3Xw7yp1scA8kDlVf60xfvu6PwnoeLyjSyJd6PqQhMKq5
UpwjGR1DAVz0pNbSW16kk1Mi/rA7d0ZaOyaHzf67b/yT6qxLyV4sG+kUEfCjB5Ef
SpZLYIIkUc/V2z+pHhP4OqhLpo7qViZMJ7J6bML8f2Rn988oHEG4/5nqy2bnO7E/
9qKAvzaONflEbWlcmJrL/E9HD8sNVMIGUAuNM7YodmV81FhjbWQBmcvIqKe++DPD
UcNzSAygjxaPYC1ZtU40USqz+V68Db9xrSfsahWNT3NhaTNso7kzzBtLxzLvQxNZ
aN0dKcGaQ7SCfIrshG+J/XP5VU/fVRSZ3Why1BmAv5TKje8J5CbyEbMtdSf7e3NS
EOmhFlbgQNnIrbp3I9uJcVyPrjvVZB+KFQ0x3Isb8UhICmKR+5KhTYn7vWh639gU
QoxfYtC5WnxoKmBReOKniE2onIlsqQUlabG9+skHd2o521TgNodkUedy0GhChxhV
JM6qNXS0mzwHE/n0xQA69tyy150raQtrITiH+1+J3leLcZ0vQS/fD/wgAxZvYAHS
AXiyL8KwW/HKdpLHfKgU49aBCeDshvS09X+9iY4eajUUL8MdUrkNcgeIgLtzIb61
JM3S53scJqzsVapD1al9O0Lud/t+dQ12OC2fQbA6O9EUFa/lm+O0KPrwAw+IaFPD
tHyK6KHzueG2ac/vcqfipbNtEBQTpLTzrUQt+17r1PA39ans+SoS7XEHwlu3pvHn
WTHBJ9JO3HqpL7QjmrBLB0h1IrvY/EGm2iEG0Tk3I7ICXr28058jnHDonsLL+0nD
1A33HAwBzFCxRhfXQTfnA+yBVjg0fBDlcVAdBDTpfFhF8oTGfFcbTlP/gWuc0N69
SEfiyLwbO+QAt+fy+AlGWNsfcAeKGDqOk7cWz8US6vj9tHtII4J6R+5mOl7ueNGS
OmcRq3QMc+8ZLSjif1Wl8pb3OAlEUjxYk+8xcAUiQ+Kr6k8rhNj9OeUfTEDTnUiv
vARrJ+MU9iHCFmL7jofpXFHsmgZsTx++Xp/GRYqheUB513BBJyJTJRrA5MmeiNj1
P10vimvYI71pCKg5yflMb2TgxK3jmHfGW9gYjhhibpxbBfuTmAIxHH6AD07FoM3J
kc9Oh+7lY5Rc63d6RRTVBLOiWxkcFo8IdXeCKHkmD1LI3paLq0Bgzn8gtrfjeOCS
jM9uvYxg6WFZSBoRzFRmjFtEOGt/Y8jsipjJgj5lsTbDBarok3k/2hTSw0JNCOXm
ucDP1DGdIzIbTmuZ7dgx9W+SKVrtYpc+OtfPkyD+5LQOmbp301l1xPI73CAyOD4p
4wXrKpEsWKrufW3a7lMKnW3p4doXxNP+UTgbNydq7g65dCIIFn8yNgowiXr5YaMZ
94RVE66yYfmoPHHeCDjNhORGfTz19FszX75S2qkz8zYp6Ij5efhcM8ICZBliSn1w
b5dMQrXQL5sVijB8KWAJ+JLuzyqZYLmuTyW3PoDsl8g8x+/F+zXAGFcOtFDrYEEI
hGQ0uDBFVHeC8WvkOaPB3KIg66z9jTLVLAD5C4+FfqxM2SpFV9migkabJOAJf1bu
3Sp9PGEXqo8asK/qIatEduboz0naBsyCSriYDIgr8ZWXIPt0sk2QpZFBB+HsVnPC
MmTB9xc2N7HdTN6xqJNm7B2Oq+7M6LftbIWz7gQE3twRmfBnTv3D+uLk4DL9vdki
JzxB6PC8qMeIS5JilVC+PhOs+hyS1Cua0+fH1hOpIFzFRAJB+zWH1VXUtYhpTqg9
mqd8/DcE8dQeAnCWE13Khtby4OZ3CPkMT6ZTO1nNFEI6tN18pZX2fEBfP/MWMjgD
ZwWJNrr3CVYcFxK9EFwZdOCpadaXddFh404PqGINjk/m1pSMpH2FY9am3sYPAANP
b+VXx8UTj/rqfmDXensKbgGp+qxOuoFiIPgChUvKs1hczBMDncJ6tov8sub36Y/q
Cp8EkyXXozBrWXQwo18boYz7AVROFkTrSLZ9VSARHUdmyfSYBHG8g3A4BzBeIGZD
0YAK2+XgHG+xc7t2eiDGJH5bxWJqqyZgDPTt1wWHNAjpDoo/xstnMxO/zm/dx2qg
qCw0B/u0rTksO7RvYLn1FyZt7DswxxzkYB4UmNPY8PFPNkAjQGnAS3MGzEG3iP4p
7F0jKoPMKjTO8v2XH3VOCbYKvpBNfWSPjELs/qWvkD+s7B3k26IswyA+LhYnI8qz
2pd1lTUqRrdFymuY75w5NYILbeFOR+/plWYKEqv5TJ9zbbp05wvwsexh08aSOlB1
N5bxRT4vKfqsOKvXW2+l4oj0oVfidlWAuVj5xgfN5AFD347wXBBUwui3Yy9Gugtj
jVO+s30mC4TdYC5eUnoisF5mzMrHAlrAWKkX/EPMLEJ7oUYRD6IlKzUJgdsIQzxP
qz9pWi1Z3cM8nkhSrR/Rw1nkFbwPC0VJQyl4gFJGcK+0+bq3JJPIhbryAGCZGNvt
KH+KAw3SO5Geqdu3j2FpKj/0KYLwMpusAJO5J1dPGi6upCKgmp/bRxe3abdAtpzX
i4HloGeb1QIZ/KUL28z5uM0u2x6w3PSKsAQNHH1V8rnpBGLG5GdPAH9oBlF3ANIB
E/7IgnPR1NZj6z49iyMkWkPnSRsaL7Ig9rLrWcfa7+x+Y/Mthlk5ich+wF92grtE
lgEaBwvSPocumK1nTBpDwGCnxHx76qiai7HncXX5PKsv+L+dRvCpZoB2sRacuE04
9VqnQiMJkJFgZypRfd5t8SMRsaC1MRjO5ip2k61ZjISlPiqwOaX4iGmx3hjVg+Za
Nz3+RK/Bw6E9Z5g9NuwFx7FReSKoHG4k4/OkCnXrXNevCZORu7TZSWwFPXABe4ew
xuMYdpeS1MzZar3Y8XGT0DqczArjOjbeuiHoRvm4oesCgNnTfbGX1XJwUcTuIu2w
wCmLTCsPyLKnIkjqQk7fB8SWmAOkjaNcRqejZ7wnAAr+yKDhydsCV6p0kaNqgIrd
QI+xbUDyxM1PxHxivEgLuGLSr45ri2Xb7/h3B+s9RF5yl3WA60z+zkMov0AaJ4OG
ktU2aItE+YIgOmYfFlkkgbeZN53b1i71zHvn6PB/VTAuLaqbeymhp8mnYvrwFEhP
/vRmNbKR+F30S5h6/JlM66L6jc6gXZ0kD6C8H/J4hCcsPPO7/YSRNPZ8yt8QdRnZ
ug2DSxv9cHV1UUl+M/63Cn3IaxKhiD2f7T8QNXLItYoWIP/8UQgXneUxYtd2RqSf
qB5xSDHW0rNBzjS1CvmWq8+oKqs/lVdzQAeIb37sgx0OO4x9Zv3enB81SmGoib/7
gvJH0de2CAuvHSuTV4tgv7Jp9C2W144TI8/AqXdErRxIXUOde7vDsiJ0wRowM/Ko
oGmZTQdEPnCPnNl98RNeNrvy3TC1YII9OwnMp1zr+YY/X4vKnXHhxIydQBij2/WE
2RY4Rxh76gKbnuuemTJl9STlV5ZZZpUGouy4HMSPVBzFXXl1XcM1A3bEFfoLTdF7
+ZBTxu5GLJ9kWOTJ2lchQ+kZyCI4Bn+WlDC+r9LgBCZaty2BChIuhlGdacSy3b10
Fi9TKW5+PY0h8R/pL3bqndct5jRfn7i3GsQUV29YEcm4o6uTTpy7sDmyG1Lv62a4
nU86FoAZJw7MuyZepUPLeGnwkYY9yVpf0QQ9jjFA/6BtG4GYdkMQ5BZay9bDBc9D
IF3X70zQc7RKiqOrr8Hie2X0dCj2qfkYdA0QMgmIpcxs8Y1dwW+0SA2UF5VMKAHp
lf893Lisa0OA1QLQcLhM0NQTnUElqHVfL2gMP2KNTer4VP2FB4b8X/Mw3lr+Vrw5
WFJXUhvR2jAK7pY0MS5mMH/65jsrqDFvjWcacApL3cAir4pNUHnR+7rAZhp5Svns
OUjR4DMMivAcdBDwVfVRe/+wGirX809bm4qSLU0IFj1gCxecEiB2MygjX+u8Fs/v
aaxb3YsmfCMotUFNufkUnH5hxTR/P9e1zBMUSbST79gLsVO3YcEBr36vSsS6gJGC
g/3DYqonYAzvCqUmoTcxmYSGhqguR+GfYkHz2EiP9Yxjy5l0nzdIM9sblALp5a1k
dhF1YJHD8CgRtOOswVQgJxd/r5nSQJ6Y0uLGtR6YJu6EilL6VsX5bYzV/YJpvHr8
OJwhemqupM1uuNwnUsKVQfAg6LPySfOtlX+zij5nMcBZzGP4ZaZJOpeI60ahpk4q
NLHFtRlaiOoR1kutNoG79qGVUhPWAIQhyxMBrIX/E4jhdFlfpWe3JgYzIWnt0R5y
Z+18Xkd6nN9xBrV3nAyfkIbYu+RSVT1/Q87hjEG1zSXHHu+HU64tHRN61GQgbn8c
7Gs42uHAplAd6R+RfIRBcgx/YffdLvmbkEa+VThQxx0VyT5GeIEhzyDcjx5yVkwv
GzCEYotCskZPza4oU1+/sRvgU8PPi12b0/p8j858CvXVYcbRMxFPOqpEW0RidfjL
irqLSJZdJaI8bfTKdtVx+whjKsK+gEqzJyxjgrVdH6i+tJ5pdnqdUt3qSkJ7i/xg
v9F8aBAf0cZ793HswyMB0mmwQMn9fzmukAyDMtpPUwho8dRIk9VjS7Q4VtPYfO6e
JbUMrY/tSsTqSwMbfBFiOVPGK0wL34CycFTsAa1u2wV5EalRrhdwrx9sYSEPBNUU
YYpGFyIPXj8/1fX2jK1x4erzJqR+hojYTtQi9akjpt0Y+bJi5UzqgsmvhgvaQVtk
iq7ciHvEV0AOJEFz+4OteAdl4J1EBIO3SqnTlfaSJ2o6kTxo4NXQsd4AhXimsBG3
UETIQOu4AMdycg7DDZMqVNqO04321XhT9+p6ioCCMX9eZWUfg6jtOk4MCzpk5xOz
P1Q91TPnk7vCq3+FEjy4WM33Bpa5NbauMl7TyrUfh+k=
`protect END_PROTECTED
