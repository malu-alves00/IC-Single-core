`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
n+jjhNT8E45Iu7I1NxGkNffTbhLD5vrpi4WXxkbqabtCN7yGKla++8YJF7+BYi6S
agury1RJE6UVX8eL0jtzy4k6OepHbm/Plq9+Dk3br9tuDpOHN5d6nTYJ5Cls32y3
hEHfjXXU8ZevjxJOg7xdWLydP8UONhn+/wwj3Y9JFJx2oV4l9J//yA9RaB02cdCo
W2aDlt1oJbraTUN0YtuYqm3CtucU9r8hmKb8RWn6cr78pIAXBJa0B0Ed9FoZ9XqX
sMsGkOlerJ8NRBv9S0Ygd4GzW4LvtWeajR6ZFkKn4brycEDvkwlbb5Kl6IB71l8C
/9vpdfdY1JE4P5vcasZc4QgZE2HJLH+kxSz0mDjxRyGmcYKLU6PM+idN+gU2SeGk
Ipl7H60WjtH9KUshrBZnTFve5Q5bUWMaj+Tcq3rN77cGuU0JtRroqxI/mU2cLThp
0CPLMKNctJ/K13CAhXVf8XKnFOYYv6WLQoD30oxxKkbgRSNU66xrh0L6hvliTfSY
E+9YnwPBqN3zYl+SoQMmiBuQvYgK3hLSOZ2qCNgiR3HiZvXvS28BHD100xzBRrOk
34Ra7fcqZI6dhLaEkCfWVAoMncrTS5Hozt9G9i1BIwwKC4BykbNXETF6fz505GVa
iBax+iemFdRw/cYga4j6ZCF2HVtbPOGkc4EelPfTMKmZ0dXY/25vwrRotsKiLPZf
J7KIav83QMOwDfAd1Ote5GHh73dmW7341YBq56H/PzJdfZNk1gLm7sFlUWo2ZvHj
8eD3CdOpzX2ZGkFeotO6zMncO/bEvkWlclRM9PWBYR1zuxsnV1sjVj1EehVdzXNZ
/bUDdFVp0Sa5I4LRVfPcrih0y2H2o3wCd+tl8bnDM45z8YzhX1DOysJsZL4j5c2m
uKN0F9UzZMzkNVbqNGxWyZsXoDITPpnSktJat6rLmi/ok7vnWpWb1ofFafWRTT2f
jnvnqMn8eQmM1w3mQWCFYR9i32Pf1S5jXjETNy0XMWz1NdqKRPsjK3idNrRjcY98
z22rJinPir0BEOhKCxJQOQhE2q3330YRh1BJZUFSBY5ePNEON7ruoNeFboMtSDgb
wZGXHyR8pItTDVMvC87R9uI+zfucIAl3+TE1Df/ahZ8fgBlLlHiuDSSH7hulS4AP
twSH6Szw43vIUtyBTrhcihF3I/MgLA0kNhs3E7q9mpLNRRbdcskDNSZyGN6Y5O2+
dXU0aV32Ob7/Laz7q3SMuoadT613vWsaUdX3UVe4vbd2oe2A9ow4PrOtAleGHL8v
ReWIX7oYMoYCjWKaIw0OIgCNuyvwXRLmQzkmjKP4bYMchL83ygcwpx5lF/gKwu0i
wANmde3iuUsDWQm2LYLikKf7q9lqYPZw1kyKB8mHzE4mnVzqlTd22qvOK4GiT4bH
iawh8PaFmsODgFycpRuGu3znBJvCcFmx+IBhXXUqFfiuClxVUax+Dx9dEaj3Ow8l
MZWTT2nwiy5C7XmsQ0Hok2hTzzLfjWPwb/w7dYBJkSnjrepHxJ8uzbFX3+7wzVDU
jtj2tj1oeA1UI9LNuHGN0R9VTZTtSnPKAN/VPBWMLml9l8wo4Agn6WC8ftDX5X/P
Q7T+b8V2unjpBr4aqAm+puEZvHcf/hfkkk1fKFdIoeP+9D3OgZ+gY0VmwEI7Vdjn
Y/F+rW/kCo5HTWaUN3l7Efxm88qJkY3FCOjSHif5oF+MBUzgS/bjC9wLbdxekcpE
9GHKReTiNXgf1sI4S0JkuRqDatce+7fHUl/IIHrQJofTzmnLWRhRjBPtWDRcANRW
IIs21F6gtOfj7h+qNjxeLjXGALsjx6g2hKAE/emc0o/oAM3N39j9aSVmfmCaNJY9
un3vRJX4/3lkJrlphHix/bFxhCjRUlIUXg9LagGbDTYVfYvvfnU+1yKVQD2yL/24
GAJ+2k+UHxRKVdDNjOZma9w9vJshSD4T3EckFIza8WQmGOs8pXaKCNZPjxTJo1T0
m6c0Yovi9230aQ4L8UcyjRENMtd5+73zCM6bbRTXfL2J1/YEzEYEFnczKTeBaPmz
TvCj9hBOzu96fSdI8wh+9BQ2OM5X82QongJzVOsttRgN6yD5w3w4d+hhgvA6/YtQ
7OwTLfKeY61sA32Y6lPqsIzu60AZnPqVlFOMvlY3tU+ILochWZv1jf9xfPhqHD42
Ru2cdpT7+iH8UnaaxXCeHEPPc0danhcYX8k2A0CfYjVMm18VAWjAhCUPnjssO6v4
MLW6SI4o6bVLgWjrbKpLG8TDWiRhjia17SXBzHeLynuge1qCiM1qqLcNC11E1ug+
Bdz6PSNkguc9q5TyrSDxmngJEuqp01rf7spXImyUa0/50d9ZcsLF2yr8Asu5Lqtb
IfQGX567YIzOk3mEZVnVNNwroUtvrNo+oZ7aP30ukKZodB2Nx+mTEDB2xx9YivPl
WKimsB64aErjXCH8G5zjQWiWkyX8ueo5ZCEAmvxfNGedGKA5qblHG/cO86LlwWg3
pkBWqZX67ahqN3iclLg9euMrJ0h9XNIJ6znggu9GZlfDLy7qDMIYkoY3blPy2jeY
PoJuqy4b+b9W8pJl3YIiKmHChh6YVcvGAt2HH7cT42EZ0dAF43zEjSqhT2J2WQSC
i2OGQ9CE1VH695xjk6z6TA==
`protect END_PROTECTED
