`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Gync52oFpePFiPyK4l58wKuCHi/Ye9G/bRmIfL96VLwhHF3sDaOW3vyK5r1DnOMa
ZMxQNGMNng8Nu3Yvt5yqBIdwdSCnQNaWgiGS1AM+PnBl4U7uSUNNrWYsLJD9jkb0
p0+xiu781hHD2M0iRcrcGpHq/YnuiP50TfrkBZTxGY8tjK6KY3S3M6wN3HJIr16g
vxS3hsUh9j0jaz2Pu7+WuHdFxJOBHYJ9eQ5KRNwC5aMilDqcf2/jpr3hNx39p9tU
EoPqt0S2kMrL4O/fW1rjN1yC8SgDxLCDkqVZK6DU6ugCGIzya952zvGn4H3FL9L+
rpMSZVL0uf+U9QVwU1jQGYRA5nDMHLhGsJhW/aacepwoSZJ/z5Qg1kI/C96q0dl7
gNvmfMGjXf9GuZBh5O51EyepXkvdXfPapj1rHt684mb10F3jJvosYcDgIMX3MBRo
pFNA/0r2rXhomjElGhv7WeBXzs4NbC9b6OHmh3HdA7/XoC41zUHr4Gp01ZNgQNnX
DnOEDAPeJGnj5XgBdYJ9PdZ4ltvG1NOntbnGepln47PlLPUx6FRB8jMGeNLh28eq
In27/t/vVrVqUekwKGdiZ9fQ924rJnGnp5zeqGQSgnsdE2SO5cIDog1Wi03erAdD
UWNSeSNmCJK8J/gbREnr6grZ7/rNZos+iGHN8vuItP+j+9VRdZKGbxyCOZW+s5bK
H1sc+xI0KbIwzhV2O4i82TtpZaSqGB9Yn8xLCxSMCBYZ69USDY3odGu+F+OlG8Iw
q5DOzhPTgKKo5iBSge81zikUZyXdGFfz5DHhtdNJyg6KZEfTxiSyFdcvGGFuLCjb
BwHmE1N7oPRiiuiGHqurnSJ1DhPT61mmWIvUoEXJoeVjK48xKOemd/YJNtczky+W
59Ivri9k05vI5RDDB3yEnaKEAu9Dvkbb9oU2fNyt9NPzsgJPwxo+cL5qBF7TIDBQ
TS8JRwukDsrroiTyNDc2vyT3ro6I3+moogX36FTmpMTA46XI1hKhCq+EyLd30xHl
Ke3NN1NmR1ptEfAwonMV2EPfSt4A22HcxMPkS0U0lcTRZO46+dfZey0R6hfQiIzx
VsPCgYaFLsrDYg292ODmjqU/z5u5ffRg5LpmY1q1ZPqnO1YnkFx8oqB7cMDnMsOA
7CswDxAnYD89wmgRTYog9y6V5eWcQVGEg++DQ/+WWxroE0FhZ820dMe/svKATqXz
8QxILHTF7mEL1AqiWdG06Yhh9miIRZ1HS51/Xh9DHhCMfo6bU9L1L3bvCW3lItZw
rh8cTW3h3SOaPsVDgi3dX014V7E+Rt5rfUatqfn9zZFfcesVAEsHRfQhPnAK1ZPf
js3wixVuUUEZI7ZOXScVFgzfY9YEDdWELkyateh0rWuOJOSriQ5RbE2i8LkphIic
idbblDETWQR8Ows/PqNk4isI7UEg4/G8a6LI5q3HEYqm+9msB5tdttFfyAnpLtp9
G7w7xEvgFaqQzXsSR/g+8xWrZU3eZfBHjmsvAyZwESuznyXgG2Ey7NznC71RFhor
Z8IJqxYuK/Wcq6k7Bu5We7Mrkvk+A6SgfJANQ3bEBG1C0KDvaUpn9T2k45sPhATK
`protect END_PROTECTED
