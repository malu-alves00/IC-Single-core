`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VtDmo4xCdnuvuOIGu12GOuH0FjzO9289vPBo8euK37E5PS8ZG3QF/p+2ECzQ4WfN
uFZi+4pM0KivqXFEFTFGMHiGrE5Pyvzoqoeth25tvFz3JVtE+gYCnLcwhEg0/Vss
I0zSD5JbVbjXj5xhKimKv+ubn5qVBe/5W71XsuIsAClvtkHWiKGRGC9UTRVovxOL
WIGCy2+uiZY9VVcMV8TPf3zjWStqjRInvuq5LCGE1TnASTjBD+l3rN/eERkq+I36
vuhp1G736sYISDjqpWPF8ik3O/EF8EVNzLszyn0wTY8n7jyA9gtEOXMd7auC56p2
IdlpuXpwSXnK5X+CtVLQsZVjxUzMdnypoFoN3FcglaRxukHgqjGRhkrBUfNMg/Iw
Vkp4ZWi2NXIzcmScn4TgKbTov2OIqG6h+Y8tvgnNLmWy3THTI8IBZnly2wjnx09r
wlqf0rfMsY25MaKNcpmoVe3HLN1ya3DiQGfVJy7I0uq/bOY91Ag5D3HJZMgFg5YI
9zcU4Q2K1cr3GZg/ZdsorCIrF/JkNrNgTHFqiARcqfVCeXXQn46qaA3S8v0BMzDd
zQV/TrLqTsc/3PaqSD0KPCfoRyUQFyO+Fh06LnMh4Aej43BRTqgBMXNeTY5rNw5N
1v1mnOwbqaWHBhGbKxNOF1AIanv1TL16X5uS86vUJSqa4RJYk9p+gxrtSzUE4xVY
Xr9rA1PK5c12eM67jL1YVu8bt475XSGmnVz4p3mdgK7fxG3ouMAdtwY/Osg5dACz
rmsqNY4VpFSR3VjcJ/cNwKsIGzC3AbXcgrgsUtwnFj3eEXEWzANNLqUUjadevbFw
ip84f1ds9VH1dxATwpliakIfKoMBnDg8bpT3vG229CvcxiWV2w2U/yWItL/N+XUZ
lIj8HmUbu8Rj3b/DWMlTftUeq2aNAaj/5MdOGVRqcKjxR64QlLRBkwtPrIHaN5v6
bj5i2vZlavkQOFIz601IFbfasBV130eK2jTjtSDNCBD9lhv3KgUJjRDXplz8QyOX
yvmzEfo9UaRpo1dpln4GhxFZBD5t3Odj4MJapokGieEd0fSLUJa6RvyXi+aQzbje
b3J0LZS3bQOjuPs1/fV+AmpJX83ERqxHPZpjoMjkSL7tdFU3zmAP3v0O+uN8CANT
+JSdqDozWg1/e58TI69Nh+v1BgDuM4tH/zRK183R9+84JNCpeSH6HrR3BXcxSoTo
IMAhQ5X1cWOCeZ40qL8bzLlWlPdNKZB8mojg71bNQTsRa66lZtL+obS0yWimp3bp
Z/byWJ/oMmBqN2i5ZdCfJia0wJz/BcaAWk084SMXQwMg9Hvv5LTh6km+VggRZs9S
JJIMD+FNLhjxNMwO4Sj4Qut7XT+jgUSZ2z6U0DGNViNPEQ2sgkV2xGGk8j49cdRn
1ILfJatVm1o2wNxdCbAW1m494z1dwRDaDyM4b/msgS4DEr9pxVGUL3+F6LIiRKYg
0vp+lwhlvIGW11G5ieJkSKULSNdA+g8mgyQfPOKitAFL9HhhCEfNr2eFRzx18hYF
txANHJdw6+9lvn8gNgZXOL0K35hAQ8Kb7AU/njfqW2taTmGLsSz2IohDUm6QRxcE
r7TM9cfcol5csMZ8AQ+Zbqle7llqZ09grOgyzPkLKm24TlSTHBbmH7MYXmc+f5aO
ltRmLXKW9BC6Hg+AkZw3yqQ0YWtFtRv7GpuLgMCgmV15FskVPtG/I4bUUMTgTXhY
kU5aq13wjqUL/w+7hAXGxPzLNKhL+E0owgJWNVDhBWFIyOT/QM8d57Sg5omTfmDp
8nJH0iR2nYqcZtwm9xOFHpojFb1YXNuHDuWvOVjXE6vloXT4tF1AGpSBDff4SoPD
1WRteVK4QJ5WixPsAYmS1EOpGQOHPzSnLgYi0Rkfo4OCAdIfn/Pvkt9jvVrcQpD1
ZU+YZN5FdDpUg05e1vR1YCzU/qenrHIGR6PgSzBvRC/W+QrRygWch6e9e44fiJJG
hweg5dc76bu6uwHK1V4A2rh+5jYN7+UkCtm4O/jW4DG2O5DEWy89uO7ueURjXYSP
41H+O19aSLuFUdV4EDSSxigw1V32OONW0Q/44/ITmeQPJmuOYxzgiwZKdL0WsUk6
RYX7uPdr63Fr++fXW+4eQxZJZ/nwUiQfsiSL4lPuSh8g0oga4KdoGKOcaq3A9UCb
UeO2KriXieVBdKqJCENIJe881qBcFnQr02yTljiYZf4TocEo+4iypw3uACB/QifI
zL4iaUce/WqaAgSsd18G7GudjuAcyb9/wllKcPdohgR6rk5shC9J4E2/VrXs1ARc
jJD5G1nez9aXtusv9QUtULb2FFxT07vO2ruORerUUd9NtatjynTYOiqVUfRB7m67
vKJmR2cR1jd2IhEOWYKSY6FJMuhxWdxhY9Vzd6MBY3u9IeOS9xfZMPHQuPwen3gj
xsIxeJ4EX36HY+Q4Es4tS1aEMomIMti0fscMTdwxLr10BSTJQy8zaBuPoXI+p1n1
He+GDWCkqzf6+9eck9/iwuSIhbJCNYB9p3tc5bmy/C1GhQkeMYYKBe7XF0F7iwXj
ck9P/FuwPuCGL+4EaF7Y3ngmA4YybwhaINnogCUm7PvUno+g1k20Aa0fF5nNTC86
UGLscRB4itoGTevt8pdgzHTwKr5JN41+/FIZCto0GIpw6ugZGyuDLj8LCYLyqx3p
8uC1HiEQpvi5J7kNkbDWcxsiO9GkfZBMYhi/7Qfhfewgo5ESInnnyR7jdYqdhDWq
H+MKroyIUyd0CS/0dQogjf5qVYp8CZg8WH3tZus9USqHtGYPwJXRAg4pXi5Rp4vu
RrgLcXvbEENIi6174u86RmI2UG8Rc9NSpPhE61w0j1oC/szqJWU8ACAgKg1xq0Eq
mLqAzq+svJzsMoPzIXU6mf6PQXkA2qXzSg9BR4wMe0SFlGZ8t4MLzP89ZzMsm3Hy
Fvm3OIk/QpAb0+kQ3G1xKnFiNDKHt0xJaMLz5Bm4J3Q2eHzxC3LDGXuBv1h7kzrX
btRiOkjgWX6Z5T9yu9b5JuEWXsq/zsdnVR1gDiLky+X5kQczYsxUWRefuh+WdKhG
+pvmaUJgDjTckvIz91K5Yz+giPZYw0Pmg12QmTG16j+pbq0H4b7M+hz7GGG7OUWG
C4mFliuqYkCu4gqUGo7NB+4o0//dienD9BNrGNaEaldK+ery7YU4enBa8hRg6vQr
4cq7cdjyipnwwFwowQZjxVlUJ1QR3JafrdADLNiz8GesE1f6tgQTV6HV9Ww29b01
Vs76xQjIYm6FQj2bVdg/5oyiyXiCMyUNLAWv7k6KLX7Wskcf2X3JZXsRoIcJssth
WeP82TzKl1P4qEBHFdvFUc4I16kF/pgc6wEEhpEPTWt6dbLNRpojUcFA3ZeG+LRA
y7kd9qA9htysbmnxDnyX9uTMkLNMrI/5NttE8v7XELV9aR4FeWOmmUarkurq2xDJ
usDfDBw2DSAfFuBAtteL8AdODWNxdDqs+qJthlM7byt9t8cY95cPiik1UjbguGFT
PGMx3vsSjvslG9MjuctoH69EijrHHqr55buItnbeNqahyft/51vYgsJRrKxK3RV7
T4G8FtTH6VRzE3uenTNTBl/wOMbxw1ACK3zl+iokmhMo09C331JCpuZTdeZ2IGkz
ZNZUrp5WSPnSNBQgHrHze69XZTKDuIaZAKkiF7K5sXLwNfg5m/0kmfrGJ9ogZkxU
BQQEaQDjLv/W8jpvxHm9+FJzlkMrzCkpOZcO2IRTmVNbzaOcuMQ992TNFRZqi68z
VIdI/CBZqaTHOX4kSK0ECruJgX6vQ73PqEhemJgxVjq0mD5RVJ0khRiTGimqk8MF
30deOhHCdmBFWfuQpWry3ZEI0i06wzqgehptV0GdPKiDhY12zD7nAkdw3vyWaQ76
1/mFJm3zkEJcl4YY9KuTNOTPhoYsmbEaXUH0uJsxD8LQlL49mv9ATLcx1E4qqrG4
uRq5ob+lQbupE8IbVqEEccSD+hSYhL2ee3+jAb1er+GT/nKzyfiTl/8sMSEfJsga
ghoBiF+uCLWLHK9XbiP5xBhLDsQe3JxGHiJT5dId1XsEy3MGXs3B/A9cAQdM4ixV
XnQm85N5QhlQS35URfca0HMcTagvlJG3WCELaKfBL9ugqxhTlhQFgTyaunhwGboT
77ely2ClUulPDt0Qp6Y595l2puHl8Lg1fVx1UYSA4n2GcmNIHbteRYgVfLw79BRN
jZkJi8qmNMmnBlGbYYJrCROJJBbSlXl2NMkthIX0BuVWGLyhOamK1/KIho9iruUH
T1BqdpKT8756GSIb2ANdGXBfa2tHjdU5hR/xcoCOEcT4+e0tir2mgbwYzJD6yKVr
XROE9Ho/x7Jt74BOfXKHPvhoysDhPFwIi9Bdg9+TwPnEfpgUvJhRhURxMM7v6ECw
NPbCJr1GJKO4C+e6WQ5snhEAmUN2eDfyYhAOQrdiNznbmrCr2XbSY+5hB4iYPtxT
3Aplwrc+xKTOrIE1jHBNCQ5whcuESEVYe5VRKLLXgldgQMN0ga8sNBjuWWy8tfS2
pgT0sD2+7wwjEMCYPMUvvo/xHlt36KzlE4Pps5+ox8uqKeMinxd1swnhlWVUz5FT
QOupBHQGDZh86cAjACKkswXDGeHDj41YrME1Pa9eJCNTEIV6mQR1SdN62PFEEiYQ
qJB71yhXN+s6KzV+jAYJZnRtdesyzbQoUdp3wwaQKG0B23qN13h6LByp86b+iYKZ
slcRhQL91nv8VgCSiNWT++J8EQzICZtkrlxCAYimKsU+9eRRGp2ZfYSYBonLb9Dg
8BdlZ+bJmDUr+2Gqyh7YiCrvgTHbe0+tapeNNvdr/++tt4X2EWcuHuasPtEzJeVs
PgRms/qfhUAVvqbfYap6EPaN7AVGA2QtF2ZL4cgV5RMnOGE2pTH0rjJIzBPogstI
mSOU3qo2bSDFbxtGA4C4rxIjwc6LjB1K9NCswro6rs4bILDgnPwcCio8FHXX5KZE
IbakpXMGU6Mi3h5ZZlPvkEqPhWlGdjb4rlp63qsZ+5Td6NdUae9wnVzBlPcC5x2Y
8tC1HTM6b+4Wwe+0c3PQpPrXw/tpHFStuZnqITmp//UM0g+p19dRw2+cXwr/7ul+
iIHVLgoizZLPFLJ4z3+c60BF6kiYO2OrqpFH0QrVILMF7ic7TF9dmq9S6tzKZaim
YPkIG4yebqCfL9XJCl9MOBqzBcs8L17TCTvYpXZv3zp8saBf0TvjQ+uCD0rHVI7U
5sIHBzGGOi+Hzri8sIeK+r5zv1PIK11bp1Ai2xy4wYja7QRVUbYaZue4P+8G0uzJ
Ab25tX9FmcXj2Dv+W2JI0qB8Qds1hN6Ah9XBPrICJgmCrMpAjQ0jJ8KkA7Z+O0sF
uhZP1q8aXjWi8RFCbYYy7JqODskpLh8taXrETei9urL1cWRczqd7ww2+67GH+SJw
oPz6XQ2nHep+LSIXG67J0BpFRQoWTEAXBYvFQfARbl/rDhthhQUT616Jo8DbV4OC
e60H2Td4aYqpiNSuDz5bX/qV7llOKQcM0/y7i36sJpHy7dEA3JXVbhCZ3tpsyWFj
ZuAEG5fzwzV84Gcf4gewsnWeyHIN162v5B2bipxDNHe87sDNho27SjKzWwis0/l8
w0Nc56zqIkimnGqBsxDZh2XEX0T4eYAEV2Oe5CE2tq95CN9QSS5f7YyFVNFSJQ2Y
4Ek1lyVKIs2bZWw9ffoNgHGAX3kLJIiURY6AMJYRtIhCZA0fntW/esqG0mhE8LgG
Cmax8o9TLxQkZ4qqRXLriab5CG3V4bzY6HQBret86+1TMNkJGOyUxYQvkSQZGWVr
jp1/GfqOBHkhAazt3nzWVK2d04sjzKiYx9XCRI+KipZDY6+jgEEX/R1xZwSmsgst
XRjrng52oaa1fixKeJWVMmOOaQA1nbkwCPH3ZD0GA81MOdWcHRFQmvfpGQa5VlRD
9Q/zv5nYbwCHA9jge4aYfDo80i/ZYau8UehsgxY2KETkuKMpXiyPZiI2l6UJ4aBv
EvoORpoMfldDfyDRSxe4uF9YXoPSrMNejy+85CSJ3E8vL3n11q9IK/BzVJ3CNeeh
tGIWHhlTl6McNPqYfKQyhsLNqhH5YhMBr+xfGql1PmSNWJeotpV3J//RE3f0ulWD
W3lEDBdSvSqrr/qrzTzC6bGON17t89My7eeCG5WAx+jWu//ntgVRR2nE/LL40am2
JBYcDUln8CnsauEu8BGlUizEVkMUXUC4nVrbZUqGjRzWfwIB1IFGIXRf1Lu5cHKD
WyVlBpnhfSHn6ius7yq+RLvRhFwqgPdBIrLcxzge1/KSklWE5Q8Gftnptf5DOfVl
uvXDCIqx/bt1wDtJVrFgF56pIcPB2T8FlfP2pmiYFp1QpgD6tSpBG8Rquk14K38J
fJk87gkl15WugmCWllLMsJLP6OduPmxQZJngeEengcleSRswVMiREsYpTBiMBRk6
lQx0lkawu4THE/mAxiiCtuJJd4vMuyISngAgwpv9uBFZREpm0XpJHL3HZ5VdufFE
PWqi2uS1Sx8wcYcIKliFRDS5aDxqVwdd0bsf5kfKtlvvWNTgkl2zBcxCIgxDfp/h
UPAff5v/n+BzGtWozJ7FSnN3rRQs3MtIyN42eU/FkuW5TQ1F8023QAFuttMZSML8
VphDZXfIKmnKp4Wnub8Y7M5RpmIak/vFpP1sP80cw5j0lLwBuablKXwmFnvUYhgD
zF3CKK+VUiMt9XM1RqJ9W6NJC51npTT95MTm5Q9W8oBJiwo1yN8ifyDJbPYfFS1N
CeKaZ3tp8kHfS6bHoHi9oDWGq7G+R/svPoG9PGqBIOJdsYTncx8UakGArAk8ipyk
OYY3ibXOkwbLSIG/D+qJLr1QuT8O+7PmzZbzOBSZfho5DNIMs30kMM6Za4ioP1CW
jNDXx6J4E36FBNsHsTiAfoUnvTBiCTGlqljpG6uU+Y5qgM9JFoO0nc2JXl+nHmn1
NSg9SrO7ifDydhFYCqTpO4xqDE5QYPKxJU3xyDHvDpVmKuMAY4Lb7r71S6L2WJ3v
gixk0trA2MDKBimGqvzlJ+RqjxOqNoFX/zjQJCCd5TLucqw8KAX2xVCWi/5qeS47
uv5DzDpW2DdrUGNFihGG4KtGyk9SIir0qs9HcyU6GHFhhTCLeW+A4D2t2MDXdC+9
vBmYPBMIRmH9N3fzbzcGsu//0PluPQbaRQGIPmghrVEwaM9uxDKsZwC+YakBP35T
nRfAf1vNFpiOFyVtilfWQt+mfpKorP9Eu5wt6W1qEtDchCkrwdBnDqJmL0C7PxIW
feO0pnrD4tzk4BZU0gZCvC7Kq7PwB6Hs6YRCnetf8MCvG+kKwRx6OMf2GK3izG+C
KEDVzo25zssbUweDTwqo7vb1pGmb8bCCV9zPm6PcCfMyJb6T5hpGVL/F9Vfk1wJH
mLdJlE5I2V+210hT6RjZ/WB/ry4+ngVql24914WJ2CG/cS5fCtTsK3USvsSy12VW
jBblE25awh2hy4/NEEdAM4lyH2F0Pv+DzjZHgc8QupJmdE1+ENVXFzNSf/RZD0SP
R2A+9A09Rrs5/WHg6t7D7OnLuCvEnf/hhbeiqYmd9MHKzkkr5m0Ba+dIxdIPvm/Y
e+vyNWnveChIE7hLhhcshizOo82NHyhombNLdA8ECOBnouKPG2sq5Qvi8NzlXfgl
Lbo2QNouQrr6GH3hViCENmlV+KCiIq+rzz3710zrIrjkTtVrv+SRS/XMC9lwnD64
Bgt+QKSainnrk66w+8R7sYGfsbGr9llyB/6NQOhY9sXGZhPgO8H3xab4q7REeFj9
vOd7GoQwubUO9p9ILMDCp5B6GEJ76SiOTrT1uRp2LDeKX1S4BoMBGvCY1i4KnEry
M4bgr67ySyfsQhgjCymgx+ipKuyHNtaJgKBf/x91yLHGW40K4YVVaVQiejS3rO0x
C8lgs1s5KBZwAriXsjGIrq43511UFnvY6eDm/1B29csrO9MATl3R9lC4BsWO2/WU
KTrELzJofp73bGADTu0A9Rr59lvfQvLVsZLOlQi8YSyDVMVfC2XtOGjh/GPZcUor
OXcyzerjnyReXvxFS7Irt4CIqkhTa5GaYFyhnwnWmiuRhXPT2gZMX9LVmQGJ4oaa
CN720BfH2Xdt10w1bjNe0rI7YqOxat6zv2b4nmFOhIT3LeOb4jgZP7PIKlvmnj5j
ROE25tuz+QLk+OkzB8Zr4bQctDzbdAJ6Q6n7hkZXXl+wHMHYKTpf9E+Q2WMtV1CI
X1hQUTfV/ad+8ajtMd8iA7twNngcMJ+ldHLD24DyHOEforAZt06QMeKc+pkvl9LC
NucjbHE7pFe93612ECRVZAjfD6797YrMpZoYjF+hVfePCUEys6XKSZ/mF2JmuyrR
6X7ULYjVFFh25vI+X1E6uyfZ4u2zhRuShdS0myx4XyKtWSRt7jPMqXq4UIqNudVt
4h1a3GnD9fjrlrgjXRAb2gXkIUtLWYgb5bglBkFS3aqoGvEgQdacIWN73QJ18uL6
t7sQSZgDhYFDf1FNUXATobA5aIeVlvgq9jbD5PaHn0tw6gvEuCezk9Ch2/2OIPvL
HphW+WgksbKxrpl3VSTagcCisBF7lEjl0OcQHzM2fZQW3bW0vQWLyl68s4DHGhKr
GlQPdse7BEA2EavfirE/GIODnrkOndHvkGHpXnt/Zdz2mlLWZFA9Vc/RiF/s8jkG
Hy9cqy+1k7Ie7nHsaADOLZvi9288f4gScAvxjVX2JcpXzXzF98AFSvfI9V/wbhmp
TDgV8+OeaAhE1omncxgL4WjYUngBMlyYHhICiIgypEr3Pghe25tAXTSsERR7rXax
xnHrUl4hzdlPMHYIKth3eawsB8SVzQBDIuoHL6OedVTJcD0QT2NQtZOJWwxugRVX
GqMVtzgwmb1oHOphV22+UJtm9LPODrn2HigIv/2lnd5XndKarlAX87JFoeccALDZ
plkXmLVy2RjygS3lwGs+b874VAV2vUgi1xS4A1yugFvoteAlqlogFMXPtKLpK0AS
gS1wiQwfhMDebzOzl4lmp0vbFs2z94i1Ei9/2yNNFiKoul2MlXvc50bREblVuP7E
JhWJxUeqzk43VfBSzDuv4vZq0tFffSgYrTYZzkbI8zDa29ztJUc18fpO4FFzwgFW
pXbpORIyIV5mxqrdc4EzI+RvLtBjAeCVK5eLK0brY6a4yraBfrnYkMGTNWfliyyZ
ovmBArs0fXST26aDybOPWJxkLwPXAs9KENLfQAbinTlsUEiOe5yW7JW7IpzHR1xI
bwyPf1FZBFgr5wBdCkBpxr3qRcg6RWryWv4bGEnfMjoi+2YWA+dhCIfHZSRyxgYj
jMXzQ17z8HYNyNKojxHi9STB/QZxkkGX3fc7qg2tY5Vxnzibv2pW69jWTwNKRPn2
pNhAB2MZVAdCGDB0fl4N4HXHiKJ9T/rGfq9tfKzWAi+KSeFKbadZwa/YNMj4N6lz
lrW8tpNjJh+DomOaXGI4HiTV2o1an6HA+TBJt4HnNRYHW4IchURFdL+JOa6cpLaG
N3sWl77YG63vcB22mgh9E8PSqt3OPKxgQo1pY3iL27PLq6Oj7rMIZn0qe+2LcWgc
J3H1JpD8IS1ibvz7/pTIKcRbmOBeqVNVDV4r36NlbwlRil/YuwV0lQ26JIDC+TEw
hbdPvrAparRy51kXKAeA+/swzomkCnP1fyD6UPK8EdJL4MQleEoJnXWWECr/K5ia
fHjbq8aK0BrHLDxBxvjzLeRftQKMwb9WptwRsPbn0qvY4tgX4sEBg0YlV367TDWG
FMfzcCKGjkvKeYhFy+3yPNhdC33wsAH1ei2B/T0H+wBP8u3SnXV03NpEnCBr+Tk3
mwMTHr7NL/hDXFwPp8ICPMW0OEZ8bFU47CgpJMVIosOpCDzb+NW/i03eTpfvO6Vt
+xWQRlr0NYqPe3DAa82X3Cyf2E5G+ngWbp+ix+9vEbMcqsKshowrXT2/FdcmYhrf
VSYy5wxH26q/rnzhFcsibcORdy6ZLDUckuYen61nty5D8Qa9/SPWBkC3UkbCiEbm
vTNjQetunQ+SNi/kXoJ6ZoFOLkWEZk36/jJg1Vp9MEN7CcWa6jfpk1ekL6SO3b7g
ulnRGf/eTww4I3hH3sMcdQm45pHyx2tuaM0/t0hBxBKMDs94y6cT93kqRPmSuV+p
+mP3yfUAgVilwDj7B5SLqiVN2L4YmDEaRlelCKQIoBveYU4SlZPgFIgHrUE+lruX
TiuJOBJ5w9CUrJ445HM6FqYXVRAv7X9Z8nS853lURUfJ2ObnyNJrSEfIWpxu195Q
LhidGpB7Vc8MVoZlYJdGutUIpFo9ZK2JMi2vV6L1EFMvHxHn+lgX3Ko2CjOLUSC9
fuoAGfmhXl3sva2nO/T9xLq5yvZpbNUmc9EYKjOasmzFIJgwEgrvNUHnFWUqyRz2
5T9C8jzs713yApdeb7bJbLCoXbRKtDU/JmPShBarV51p0oezFI7YMIdGAgFZqTuW
xBLgfM5VSgbY/LrHJyrh6Ufz5sYEcVFOcUFZfAzOqAuiIjlZFOGlx9lBdz5K6AJL
Jheg/R9lwA3AgQYrERZrGb6gq6X4ML3KLlQcC8gAnTReQaa9jKgqqp40TQrqUIfy
piVA782s6+Td0zG1zqSpdQ6aGMcZB9dSh0Fb5muzfZo9Rpg84+Cp2Ef96ADGHFfp
YY7N6R4XaIbC3YsHQTPEw7RHpiwS64OnY8rg4baHBj0wUK0v6AFzYlvkHQhuoYjM
OMTjl7YBqNNoeGB8OmkiBWKOT9UxSzwP9WxM0Aoq2B0Qd95hfZfDKW9Y9wFaogh6
IWFSnRBab6tDYY15F9RnUowPQY922zDdMkMxc7h576hUL2X/8yTNkeIURWgbl4nn
uOEDpKEMm7U1YxmuJP4Hf2cQpdvf9LsIfAVQSDBF6avdfHer1CLyPzAlN0GibPrF
TiNiP7J6lqFfhZdKC/8SCx+r6reEWXnIn9z85EyDqxO2MOQtVkU+j/5jRtCZCOYt
NLR0P1oG3/5f7TWaX982CfL8zFuTRv09FQX/eISOwk6e++cMwxpyZ1IOdJuNrDqe
0t9IoPQSjS48fuDR602SjOzZV5U6bhal7taj639Y2uCSsEkPuuehWEtjOdsIWWUd
RgMy2FDgVpmskvPhKwNyotaZROc0NvY9tSCIBgeG4kDltjP1AZnPgqR5yo+SjN9M
tEFE7ptrt874ioBPsSe6UrPnOsq+5ROvTBBGBgVXkuEVIR/ALRSkTgWFEX9iEK5V
Kn7CS1yR60dI0sh6qrtjcfHJFjUumMyxheYgLPm2uL56fwyq0QvHP7yN12h/1QW4
Kr9SgB08a4NmXqVARrvOshf0uQJuKsGvGu92hDLcWC99xJNCg0OFCMBQZeEW/dGF
/LrA0J8NYo6XQcNx1NludDoM+bTuj+M0l9qvX7QQfMSGMS/Y2mmQ5rxv8tAEbJus
I/dAbHVr9gzvMKMNPYYFafhToauzxNxMff0jz598WLY0gVhE1loO8tevI4XgVCgh
NaN0cG6Nf6RDpbW8qXRiduCCcSOcF+itbI3+Aio+BQGVy8ngqNmiL+4vcZ7oLLFC
qDTTQws7yeyEASlvsx9VJTj6m08APuJ7GIQmj+Oes8Dr9drCDXsQrReaywNKOOFd
qbPiI+SchD+JcknvtyTdhgkryJZR32UzIxyluuEHNE6AZ5GVPrJS/Wu4DOmWpJ1F
aTgyt6JyEDfJtgQeWvHQo51R875dj6HLWsV4TcKfrnmgkGCjyOvQz1xB2TKiKRFT
JlAJ5qOk5CypCgWrki5H9gS6i9bm0EQh9rWhCHbprDygK0n0/SZC1cT0cps6HW2c
Vx20v3wD/Bax4/LbPv6lK9zgaJ5h7FiLixzmGM3IDR83H1U+SAqjSE7ooUaYrIUT
va0aMbDYM3XeEVbFGLhkbZDRut+9ToDYkQp8eyx16c4KoYDJZmHWg7GzRjRVfn0Q
D098C9kMVqfGggWl+UwTN7VG56SFhSkjMImKJ0pV/82lMhWSZcNEQc0S/WVQP4oC
OW5s6wDGArORjQAAFkObPOocJJzQZ12x+AiImPT6wMcbc1KF6RvcqBoM8IgB/Sqz
hcC7BpN7DNx5fVlnkTwCZf4hScjDOqIjiA26GBwWoDP7ZVcBln6e6RnaZ3aSpt4H
zAc8yZwl0YeWIZnjcnC3ru04cY1BNJ2YLqpQtayXUYNnRlOOHXfFuhHthsHXFa7U
OhwDiYz/uBNOBID8R0tueWGD/JRuNKCHtk9iHGBZGK9yNRYGLaW4gXj57qOpyHMz
XkNOXxxTKOjqFqqgs+0S/YBuvjpLTIydFoayg52yv26m+6h+ByishSYBsQg5+AZn
LZhIjHP+fNzg/2yl2xJbkRoXoSpB8QaIZdMO7j0phJR8wfd1iXjF53TD5iTmkuC7
jnbzX6E9ZBH+2UdO3ostJqYRAvH3P7GMX2rBUtyMxlLtp4HXwZf5Msj+D0zmMw4k
pSfLfwb13QeAmawh4B3G0uyylhhqJY6QCN1vhKmPiF+5wqC4TvsZndNPyrPi5a0G
t1Y3Si/ul8k0v6UHdukIkXpPDyvJiiL4qGXoBh/5IkZGCBk7aTDub0gTAzdvpdZJ
6jDrjGRVwrKyI9rc9yMrmZeQbLfcb8a9UbcJs07tbkIyw5pSppyzY+C0/JmyxgNs
pY8BptgIcREDTcatcPFo5klIVVWAUQ8FY/ueeUf2AVW94bVY3Hh0zIQUdjVKzD+y
9vnJcGh0uxOGlCE9yzuHGkzZPUBGDzItzEceiZLdgS/6rTqMAE8AL1t2GAXueZtd
Y5B1bCo2iK/qoFKm0V37ssNn2vo5T1arWFRVTAh9iTS7vckmHEghYblWgZHZbGNP
sGIK0x4Fntcu6oBq9UOQzTsHiFlh5Ckn07aOMa6lHnJuO4J4d8nujgp1SVRF9CoY
zunKsYvrCDLI8rrzhVkRVsDsTTFJ7+IIwPF9MIpPm4Hb9QLJaCyoqLQ4RoS8PT56
WC30E0a55AJoTxpDViUbb0AjXKcv/070jfnMdEpiWo2iHkq5DPMnDqoYSBfCyxKg
etfnE9npUGTSNnLwYugAyN097hwKtixdiHLwiR1LUctgESp5Hbzbj+wyU2sN4aiM
Y1T58BaLPTEE2VBfVSSnsPhT71Zr0cWq9zeyonBYtBHaLFuNPOAIt8iDZwk7rm5J
j2iq8QHpTerUZwHn6JSbNC4jfI2JDqH07jEYcgo3IzcoJgyMBKtTefF2FIjaaduZ
sIV/TcnubPfoJ3zckkwy8hidO2mZy1FKPFFoDy6ZseFYPEceJ8/jeHWb5e6b6k7K
VO/CdXFa8mXBST6WXLsWyGePABo3NTRnCVlUnLPbO1+QZQv5QZIc9nG+luCIMaN3
7rKJ5nz4nAFB6MVGG/hl1LfnOhpXbiWD0hz0mxbTyi36XlVJuDOrDmwjwZdxYFGN
ht0BZ4nZs0pjb90fEf6JabCrAFN8QICF0w7F0mL+QSLJntSxzbGgv3M8qZnMu1p4
tYn5fXx/iSOQwVTOn277Zg6Fk1h+SG47powlZv6tyOOGhUBjaQLIdhGlSb3X90Sk
zLQl46rUPz/+xaQKwHVgnCnhl+adha+RvoQYVoHvZv57/FfvOMfjarfQwSSw9xjX
DZU8ddntopi7rQwl1oIROoCeblQeSp4e4rr1frDKaEmhTXn42LwhlRK3Hyp0jwVm
3k/Znzmf56UomD4bEqTTZzUzUkwNZZ2XyqfA1/sCW5lozd9y48332DAyXYk8hPWu
TlyuGC+Ymqrag9u/davuuB+pTI9Zd+C/SIiy3/mJ7lDKl1aK5IlZnX3ijhaWVFLq
2kN7XNnRTZkC/6f366OM8IvH/usV6Jg4sy4FhSq0Oc1iO5h5ke1ioLzCY/wFX7Hs
UyDUv0/n+Xgl9Lj9aghehObMSTlsNSi+s/6TvyCWsv2g3fcU2TDJ1aMdUwKLctcp
H/KE9BAbHyon7cMuphDryxVTnZkj4gfRN0Y2/0RwLLC9cQJvaaEc8rjtLT52eUgY
LCQKNLzhIAeZHFgmuVQBSiLoGFNwzz7N/Yh3zkoljAQwAM4FmUFa0pCYVJnJSu3j
L8BGuP03xqRn77ClQpJjGbda+v2j/hnjjoXf/z+oUJlzzKMY8r+fh3RqnkzIKhYE
gShsNuuCAPszN+KOB0r8PPrTw8eQ8tp/vEfxX5sdaTjryVFaNiYPZjqgDcHBOvYC
qSlsLzNj0JQC0mUW8abQedQvA2wlA3iU+TFuo05nFhLYHyimEQvFQJGmxcMXp2QR
PO6XfQ6iLYmeTaoWfBrfSUjakOPDsLqKFgTjIjTFSbcxz8ZPwMlyolTZCZVS3vaQ
Tc4AVn4EIRPdYrdlNdaJiVzjxqBLXNAozcEvNG+pIwvuz7rTSt2LCOclMoH5fhmc
stpfPzDoX/zsc2FdjJvtz+HY+R75B1DABAXOWlaSx/my+BZ9JrUoGo18LDbe56np
fZCAf+pj2W7RXgbZn9rg4KfMEYxyKCFSPwlVaUbCwFONktlUEGkmuaNQ78NetdQ5
cpJhj2XA8C3DT8LI5Eiwgpe9bu9vYsnpj1Q53pQ5NvP9S4M33X5wF9KT6pKZv6E8
efvYYNgy+BCddmwhuCf3Qs5qsierznHNBonk7zUPCskoosRFaLAq98HmfXPHYYJ1
iGEe15pvKZQAlxA9i4pgWw4zCDCuf0JIJog0ve4C4pihjw8LpyF0ZmuG9xdoxodz
KUZPhSOFXFPAaKm1UjKA6THMSayIGBNVEYXr2aQCWpo5DxnshiqclPONuY1PLC+p
7LxvGzTBzI7DUPJ9rRwcBA/ivviOYdU62r6PdCUUKT5CGqO8eCJVA09GhOltO34a
G5HPCEWLjF/CWuMMYCE8BP2YB7Rsu1e34nddXoZyfnTFp+AZ1rgE7gttN7SnLpFV
DiBmz4AS8tIercC5AsnOGKAl7797Is+RJUu3gQn5t5X7pKaH3n7Q4KbQOBdC/i3N
+iOeQzKSluCyqYdtmJVQCzlM+PFrpJ+69jpowAaCB4Mtm2qlV08yZ03fZm3xOyPO
T6cZubMR21/fMTx9duPZaoCDW9mR1GEdSq+bLXhrR9upKvKSjuBnj9KT+bjWB0gR
VUy1RzvvUnJrQf4RTqCxVuh4lGJmUvYVkDSPBuQZpPw+4DfaYe15xDnJTy+Z5sCb
P6Kn7DBgFS/xJeVGAFsuTpYBRSl3F89Br7+LB8rcDaOe4DBmLrEursja91XB/zYg
bSgXfok5yWbyoMHJlpgDZdY23fbXbC81SpqC1nP1THExuUMLuuhD4v/1/9kgm7yx
A8EPtWzVhcxThtrB8K0HURKouZFmDEePtvVjYmyCFsZa1moNfl1nV9KtbfTAT1bj
QDfqkS4yORCzKnvbNzAKxBC6PMWQNzEFeHTmMOilS6Wmv/gl1ZeGUSBnB8oSLT/E
smavvNLJPu5oJvdak9d7rUO3bhT7SMQ4HsQonbB2JyUwbIwLJOw8lnxHoj1h07UX
FcrLcKNp4u8wpZWVzTPDmBvzWVj2cui60GMDBlN0Lh7Pdl7OcH/QE4rOg5QLQAyP
OivRZWQJLua0NtUY0v2lyBHUwr7luvH6vzQfFpxuLT2XSmH/u/0ijalh3Mn09u3K
mUuGRlpTB+gr8Ja8eAP+t5WLJQJEC985+3P+uG0xSZFhUVEMWZNnUZI6NOIN2SxR
x/oxHdc39n9onHxJDdsxIdT0qGZ/Iunle8T/7w6xaFdvMzr8OYRd2TJHsdmKY3hb
4jsugzN0VA7rCczc/MEdfKZcLGBuj559WJNtjgbA/gjnPkDhSHx+GxZ5pGY8cVMp
ZkjUHGLy1AKxSmfZlhfscH+T3zbdE59KxmYOlrCMrjZtSjluYsQvfLgiIoQRUs7i
gwvnlZcQurRoONdg6hMC963vhbO/Jix7QfCxIFO/eATMq2o6jEtmN3Xp/4Y4tryx
axr5J92S2CKq0G+yLMYyK9LMyY5pYC8XqfmGDgfktrt6ivFeuUWuoyH5UFHdCXtQ
svZRaGoB2RNzJ6/Th9hHOM/dIb617BjWn3W3hfnZZroGn80kiBrmbiEGSdpDfVCc
u6ixp0ElMZKph4+rtpe3YtHjW3ZQ9BJCA/Q/S0gwBQ7+RFK8sHeMC9nva8tkPhrT
XAo/qH7ljO2sXpdwzCYVQ2xrtv4YxiWZ1VZ9MSP13hxVanNBvNc7tVF1Te451x/a
D3ASQoBd51gWsIZ6lvGx/1Vp2SqogN7odl2eEW3W4VokE9ozPm2G8EWrvsDXEUwy
+rvuBskq21kGsvEHeHBaT5hGdm5zXXb1lUdSSpB18NdDA0HQ70nqzbXo9meXWuXs
2u1PLNfcYjZBRg+9pPzfB9Ox7t7ZCLDEn9kbwNDEi4pgTwGeEIeTzdLvTqS85e5v
S6BgtFJw5P3Jz4vjc5+nv5X3/987ggV1KiWrqNmGWaM4y7ld76fCaXUBBMQNktEa
asUDbLz+uo82qLjdt99YDv5DEG21Ps7VMwtkeUxPPsMfikhFuMTuGMPlFhhWgMkt
QkVATpoCuhkQIlSN47aTc6e1gIAPJE+sx4y/T8cYD0ak4JC3GKafLtOwC9Cs/SwN
0Yvx7Q7X+EpPhuKj9n3XwdkkJ4Uza1pX81Y5ep0eNa+HIoX/ZnObt86oszUYdi+t
zvDd5iwyKeAJd24qIcxx36EmYYQFecWuvMF08MUAyVLjKjknZaMK5NP+xr2G4Lp0
cheCqmivYQcN5lELdxTlLWQjixM1jJ1f/l9IIjmE9Zw4kN+ZTJsEGjix7lcCJG5k
QfLi9gebOyr/YeNdDwqULNKZvpM2bpnBWvzLHznLdLF7VgXp47vTVaxVWpy88OLW
WTbG2fRFEzVawnnocB/bt9zuJdagcCfxJ4BwoxauWPuKL+TUGxeEKhAk18cK/9vt
st94bUOhD8hlPNQDW0/Ro4i7rwQmhDyYara993NvIHG4002DpyRiEnIdjgp8f12N
iuzJdaUMYtpfvHlGgN+/Dnw5HE7XBfjFqeroDnfUt/4nKwE8UeJx5vKCxnx0+Rwq
vigL0dEgR1WShwePWdlgyoVxzkARJ6ETqT1gd8B3GiO/A3X8fZ0jMRlwXn8IGdUp
aFZeKTIBMxPaHmk2GJ0x/guf2I6nVy3RPeB+w8hKKDvnoLvxRzAVvlUvXLrkumyv
LWL57YczRMDeFBa58kT9U9pqg9GhVBnUP1jVA5AFuuiLnjSmDdTHkj2CYry51TDN
cXDjqiGyicU0+uA1Uwqvjgr5d7YhftHBz/DEmx24CULkIDXeOjmoVn3iMJDwmHbZ
rzW75QKugsAU03yleQKxsW72a5cbwPWpoTDael7ZnrtZWkbnMnwIuR4h9sSYz6La
VF5CaG5j0KT4vLJd7M4tjRE6wjBEt2B3yG1NnI/f2YQ+4OLOMPuB1+KsHp1Nivi0
CBCc+QiuEcOo6gasEHqpWYloBse5A9S7Q0vKhlGi/XWt4u/E/+JLrlZV+YxvmP6I
0Ko8uXce3pFgDHw1gfBGLSu1l9nz4oi8FIK/5cowuy6wLrht1bPvpI5vKDoJ21Xh
UOx6bJNZ+cVgLq1FuIrlvVl/3lazcFdD0ZijVh1yg7AO1y6DwO/fq5jA4SRWR9XU
g5eJMpn/FtOxk3a1wvv7VgVCqe82b1BjSuawzWThaZHVEAcUR9rxpzryCzzyaNT0
p3WA2R69091W2vYh+wLR+LM+KF0Oo2fWSmLLrBSLX3XFL+G+G1AYL9APzVKCozX2
Qv2WBScLwHsBxlpZZ7xq5vp7OjiR8e2j2T1it7EPVwOdglQds3TlMllrrFX5pW+Y
hULhgjnOMDQbhrikj9NDI+vxpmORiSeCRExqocbujrjYeeFpFRaEbFzuVe43CdTS
5crSKoWgx3CqgfB3yyN+k7XXinw9pzN2LC5W3L22ihrkgvtYwU9huce/T2YlrJvK
frS1DHBhL4CM5JSpuFaTJ13x46d/8xmfZF69AO1SBBUwy4XRmEMNdomfOY3H1WJl
RmE+elPwSKJ43mjdI3VQqd5iRx5Rjk/1DCKdmV47BUZXCOsG4oA9wAp0WldB3spM
6+IpfdQSYixppS/bp1GGtu1ernJKkYRtlaXuFBSVSNQDTTqVU3670Lu4cPu2cpz0
YMovDOFSn9K4PfwNn+/dWBSSiZI3qhyg3bxAojaAuAeoUtQgv3lysRPCUwUSOzYx
UbuXEwDQ3Zyy+Q8vpk5dn9XME0N9z71prXuXKiNy9edxB2VIgLO40/2xmNt79WNp
C41AN5tm1SiXm6dMTkNHsWSraEqs0x7uahKAzVIi2I89HNpZMBh6jqVwdA4qwxAY
ZPm7ET8eue29Q/1h9jv8uNAS3tOvCIc4AcHjCr5/Sj8Jq+od5A4/O4kErLoNVf4B
j5wzL3mYSCxWCXjcD15k2ZcQnbf2a68aQ6xHGeaErzC0reTtpZW8cG6qaKnwOwfm
5MsoI9/Vmau8Y47slorEGG9INnsavJNH48SynlFYWOh2uLGUkZK5uU68QW2GL4UW
W/xZeA7a7knvWwY2qyGUFCqtEtLqJipLUdttjez4UE+YgLMjBzNyHNV+Y70zlaeK
AaCeGTwchoODjs7WSOt15Qbqbf+bHkzGIQgShWU3xfRxLbA2vuh/LxrWprG9peuq
/LsdpY/PHVeDE621LBFI9HA+jN9N1t/6+JJ4X5d29SkSzKZih3911qyzXO8ULQqO
U1J8OLD8CYmvwUiRWgPY32pvL+aYsxhzgN27FYLIkbCfVRboZe3dSa1qTShmf8eQ
nZ2UuZANXEmvic/KLatIdtjnJOePly1JowkzXuRYA+mVJyEXnPool3ZxeCCyax1m
JYK+Md8UH32TQiLWzUantEL2/axQ9+5ZSo1ylB9EMby/F/i8bbespqjJ9nQFDXFr
s+vCMptQM5HCDv6DXBe2a88DKblGnOIM9iWkiYEMcw0fHQmtZAKp4Uuyc/ZXpHt5
BehhWS9DJtkLEUn6WwLXECeFl29PbTBQy22dG4RUrg3Rm1MQTaWpXAenfj2IPWDt
xbpZgzERbqCI23nFYbgNZxXbV37R9eBnTA9wAEodyyjwBLC2iDW2Azjor5Ftv9jZ
ZjlryeyQsV9InkCY2k+usqLkKzfK0IH2hmZpI0si2HH0XABORBUcLn3lrYSQz1AN
I1+0wBap0OkzsX/S5/56BfUzS/sBrIWpe25bLjeXTMtlQX7vigyeQgTBn8IIeYlW
cW1j3/bpC4Lg7hUxhgouPU0HzTLSKnXeTTcBq9a9R1U4FrdjAEVEDVGw7uyCgmzw
PrWREYXxQPdwUwM00VFPMFapXRpIpDDpXyruaTxE+cr3VDtbPUBKXmdm1GdB+H13
KrvuWwJSlUmTQXy1WjNiDQTRByyEiF9jMXxBaMi/8OOH79IUDdakxKfeXQKZaA2X
yVLPaeexcSL1OJmcDgavp3+V/X2AobBYSbFYOLB+x9ljQy4tUdMEm1EH+HoM8Euz
kzA9NxWed9AR8ABMddTXIV3z/ykC6SG4RNUc9CKqYOcmim6KO+xj+ya4t+8qEVIb
TeA2gMxNGnAG/hrhH7UNCwH9tBxFPOEdpeHQXNLstHxSE1SMA65O0XS3Aa/umuf9
eZ2wUPKDatlfk1ieTxyWM0tUQsA4KnqmzZl1jQlL/BoyL99eV8wiy7RadzoHFwLw
pyoLFC7C8i7ybDAaLoepsSFw4+48czgM4ljq1E/Oxm2vwHEP9ms9WoaLiTLvo6oN
488W43fkIIiOFASvnpwYIWipFhXzgMxToHJ5eD2yiFR+VEeijldpUjla7uMHWQR0
HZirapHgu2eeE2WQw4Qu+i/oUk7rj+ImBj6oyj9No4uXKEibLarhWisr1N1TwkPk
8lZpKH25XQJ5AWqmE4SFTJuC0sI4kl0DDR5epbCRbsaTS3o5vdRsGsRUUnLQxfgD
pS8lSdApTQfj4KSYkAhusDAk7KsBwP29Colvuu8BlZii83gS+mzXiIoA4J8Y1yCJ
v8eYrrtDoM5P9qjjyLddqjiu9jPdHlfngzd5QGlrFn8gaASP+NDKRNMnTBi8a86k
DxUpgqwyglPJKOT6a2bIXju/3+Ehxov3djbK6K1PL0YoxxSYcQ6lCwDG4deqHQTL
0hj1rAD/xs3JRy9uKr7Iceyy/fEnp+6UpsTPvIJPqDPhmb5d0Fl9hDuHvzu0ecUk
6CZ/kTmCGwUL+4UvGS6AI2NFDC82/N89hFxA5wJrFR7uiNTNxadNUcA0ZLve0E1v
DufqVIAT4oTXrgwei3xN3J6RMW3gceDb0XLNRscs5gDx4IZPVM8RVx7CIA361WyH
zMKFe8LKLL6uuKN95+evhGdblKVR7GI9NOcPaFvfwLpkwDm32p3ncN5/MpL0cYhL
+pXJzMihuoADA5k/hWT3OTGClKPrb9HPCbirC2kWYiAH+JP7Z0crePmFOgXC5mva
PPuGq0TLvR7Wd3dJaJcmsZuWueNvMCDerEShdOjUzJ793pPL5lleeKTe6t3JagWy
DG/uD8W9jBm4aNKXHLhxXs2u08uAwAxyXlkr20ZI0hbslGRY6W2n0vLO+E4OYMvx
XLqf2wKwQB0lMjV3bEVxe6atzM8soffnhXR5+N6xb8TLScxhaoHKds80l9GFQEyx
52IoHZrz5N3VJIvaBOdrnYTHR1LprKMpy6HigD1hcqFISv2QgXzvdRGNOKway/3V
BuUD070KknMCNdp8UYtLF3UKthI7QT0XkkrWn7+A+x9A8u1tKr8wo8qz/nq3q031
iCauQWHOYU3JWlSG993G1Q8CGhLHcGfeTaey+TmAVhRgI7/syLE/3SDZOjQtayB2
6FF0oUQ5a2yGx+bQj1aLzY/CL+mwMzzkrV06BlGWf9FjT+F9GoF1zjTzIYjJRrwS
+Qb060cG0nFXb4+yCG59zkExfEICSDqynKVeVsYAz/SxSPk8+RZOjNVcVW5hK8N9
JOVDRTtZGxneC8Kd5jErYk+5IhjHCEhbKMI6zjiq0TeJS542nCIF/tCqMkFG365u
B/DT+1aJcxbT0gcNmEFz2lvNtc9Jxd11wNm+jWrSJSPayYMf/s8GQmYz1Lrgys/L
Q46nVvQsNLEUvsQgsWOuxd4fn5Xs7SYq6f48zaHKFfNGR4tvsYvU3oCWV6HuJHUU
mfyRqydnn0C5ulFlRaQhehKT/dUCDiusAwue6HTq7Km296NA6QL1VzpyrmETRC/C
ozOQKmPLK4izwG5oB9JHW/s6x55NIrV1A+P84pBT98+SEQFJxYG/CMS4Z/y/b1g7
F9apYeQlwWw2URpbfEvJxcEVwl3mIjRhDcDfUhBz3Ak=
`protect END_PROTECTED
