`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PEDSh3JbsYyG3y8mNoi98En5+rH37BZY/197k1Y6GazdL0iynyuMOW0AUGoXUhy+
VgyVg0cf/4SgG8BhQUGJz3pX5KzBv4HtP1uig+dM56S5NTtlO7bYZBRANZaeFs5v
AeZ3Sx5sG8uWuH8nKTkeDm3FzFeq0z9ExU182hPOm9gJyTwyCUnpHu5OvCywkqCi
bjgMmKKzi0weDXWHYTwVGATTtMqCUeSNmBQdoKJ+EPKse5lPhVVkdgVXo7z1MqOp
ImV0YUuZGPm0Wd9xs5NE9g==
`protect END_PROTECTED
