`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oky6fyHaHQLpWpH0tt2ZWutyI6N1eDML5P2CxpuEnZeRvPavH/Jvt4MgdMt5DrRN
8ozTUPriG8fc8VIkVXQYg6TS1FSY4bSA1qhK7Pd7RaclRCjPgx44cjxzmyErafe2
XddLYkgNGZOrbDuuNm9sTSQFr0eEy+GgQeharQ8FO4cLMRtaxGSph7nRDOkaZK3M
/FzoaL1omH3cVf9SMUKuoX8WDg3Wmme8/wNkgFKQwl4yBtHSnITKsvZL8s4oFPLy
KQEgecV9oHd6aiWxGYaMtqheo5Y3cay/9sovGwksKEWEiSQgyu9Tn7/DJtNmOmja
S1XLvqz+t6CHI74FuulUuHxP7xX1V69K5TsdQySVuR2avZoTLP8pDZlRQrYB8GwU
SVhFj6z+4JuWf/ufBWztqQ+EhdXTENEjFV0OfOalvynd9rDPW85DG31anMLWdlc9
kiFC0zyWkFFl6GxTSgpQGROMxvCiNeAMCy5fjdafXhYDMR5xC3lJNbS5p7BVTBpP
OQZmoC30fHtoQbZI2PlWMCluUue5eGEf2L6KTk3OO/SWJgOZHWWa6pTRWgx00FyS
EuWrdNszcjt8uhrfd4pnZbKCdm9DENV39x8Gk0UN8yfWo8KSnzKisj5e+OQXX294
XtSqPdU0YKWEaWHhd2GQofheKtYvqHRuRrJt7oXKlScsFpFGnwWyjRsPwLxW4W03
yOEL/itIjJCRjnl1KKPKuGazjafICc7Skd7M6qkw9wQvkFx+gyGKIB4700XRKZZQ
bg1MGjk/6B7/6kR2MNlpgYMgiTyqOC5FHORvUdVhm+danspLhN8m5kaKce1BCXvV
HPvHgi4d2Bp0Xl/zXIlueGrcYMNmq7nVWheCUSiEOv3jzzV7PGrLSdtpLpNHIE8D
evCO6Scu0ZlxqStmpC+wwpQJAkW4ce+7g8TbBeVRGyOlavAlG4+PfC8veE32P73Q
WmIsTicWyxnj9aFtBQgdu+GO8yMz7WcNjYPfRsG4AI/541vusMLF4a64jkf/NMuC
6HHPn7X1Mgzp+dNq9dJ0w2TPdVbXVawrlgk7j3ae9dGwVMSZTbKc9blsEO5h4Zk+
q0ZFRIzR1A3JsToTYZtLLT/CA/bBtPuv7P1DEXVcUpDDtRyfMTLJnPtl+HQVgIvN
Cz07QUQbQA7pIOKvQtUHqClUW7ckqMd+CvmIjyWsG/LgwpXTGu4RmZ65xQT+37D1
KH8IvbT7WYlmZR2XVXF6/Irq8rpc6XwzGTT4PO6HvBmoKytYM+JAqX0EyrZ1ydVT
sKt/VaZmX5JU1AzkwR98YshaqDU1rjnJpUPHEwYzFQtwW9YP2/e/IIhe7lJaMq/n
pnkGwYxgg6T5sXa1WhbRqSyMzNZZMogJm5sQ+XpOUFWgqcriPHT28dtnfAqbfA2n
CZEWJDz4mydfB8WjR7Lfg58cUJhVw98WAa+4Q+di+zneoOnmvq1yAyLobGC2HbWr
lo7UoNunTb+t/ikfzjJXwfmDAj+Gm5HLtH6Fash6ALRIRXi+iLZBNSpqgVqdpcKS
YP+OFNAO9ciVBbn4QvLDe1EtZ30eKpPvueEGNwzMemA/iHpDPXSM/lHo35eP90id
xX/3g2JIrXoUA2EjsiQXH38acDf1uPCuzH/5Fj+pDHLdcFeoIpx1QqGqJhgqHH9Q
AJ1I11owFPgqoNanYwL6cdyLmEOO/Gj76iniVAI0B6VFus+2r/PAh5HzBhoFw7nl
XUJabjeMJ4yhG7B4Lh5QiEX9bOqLlxI0vByosKvj3MgFspD74UqA1j2DdziJ8HjT
x9jcn+1ZADH51rEFGIPpCEks9AkZznIV4GirSl1L3ygaGLNzI9AbaIuw/GcwQSsl
JMGA+Rg4CFLk6GwZKARRY42oi5VkRRNSgg2lC3P0zrs+xJyZjxTy5s1cES/0FSWx
a+7y9zd9WfTwCv24t/Tc5AqJjVyReB+qbq1vXmjeEx5xlUoezaPhRr6vVVp7eFDR
QH8p8AEDPbMejab1AJXIkevpWWV4aHDVqXErb09qxUUYHn1dLKoxqPIsYdkCv4+y
+5uylPmzdt5Skjg+NATDOeaLl2yRfNC72lA8e37D4BZ9aHBvGCNBnjDPnooV3I7F
dUz+yeAi8iKZ2ftdXDJbMbaaLRHeFN8ifi/fC4sTdXb4NlQAguH7+1fvZtg6/HL5
Z+c3eNSqIba3ckpTrHcpaVX5S4lUhmwQ1LFJadmaaHk=
`protect END_PROTECTED
