`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+YUlmZHZ8zUGXn44V50lHUgckJ4tqWGBUbnzMpsrdBY5rwgkx27ql/7xH7GxucuS
jd4hatunfTUKuXoZHxGkAaLWiD2lD2r13W2U8Yc67SYlSU5bUEyKO4vInvial95B
/xx5zw3YduikTaAs9YioBUfy+OZ5uLgmCMYlfPu3lz7UhUwtBEN8Qoz1aqVR6miD
VRJNQaSwHliff4CVsN4kr1LM12CK4mv2RDXLbPO3iElGZmZAN28EKnVvigQj791Q
Ur4LRdxJjLoB2QJj6obVRRdDv16i2qPMKYyEJUc0hIA5N2oZVRyFXCzPpMSZUuyh
zv4FtoumnfBTU9OH7oX9aM1rV1Rs+zeEp+Mgre2T6bs9ip+H701ZCqjVt66muBKf
aW7qUa/DCjipIpO8lj9XsEH+FdHH5jIEMD0AJTxe2lYhwUcTeE2o9uNg5Hzbf6a3
tj1rTC0ZKiTC/egc/WyiIfQZA6jyCiZnn5psMOSz/ubFAo3xUiL1MNLFPuyTQMic
Y91drmWOqR5FlK6ppY4ge8+9uMsg8IMW6hYjpsWhk4Gf9dwFZmZ3yMVYyn5J3NZX
gbtKQ2vAd2sk6o1wTn0YjuAysr3NJ7VbQuZdm/GCrX9TE/Q2NQqArErDspN/R9mp
RbcU46fLKBrSQlWAn4dH7N1ecmueKbyNp6IxEUtPZCFDpCc/hrNIxu95+MoKke3B
RdWgWqliVZJbq+/B2Td+mikPA41zVeXpb4bB6OlhAhrU43dejlI7AmI50jRkzmcj
KMnOA1K/QEVVry8P/4as88bs7htbu2j70tw3DNmyS5vQJT3jXv5kJNnP+Y0MCpZK
vLl1Oh38ztJp6Ab+p7dp7LzCU5Z8Xi3WD1FhiWVdWz+xgEhbtM/SnErmgEoJrT3k
wjkhS+pKSg3EPtezNtBrH7jN7mTVVT+kdk2itbFDVoEa074PwZUg9Mp/DMJpsk5z
`protect END_PROTECTED
