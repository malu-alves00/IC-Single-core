`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RyMwS9TcRdfOLEYerFXRfj15kwxGD6oOMXC8UT3zn4eS5sTNw2s07phyqs0OX7QQ
JHSgcCmBfm6ZgdheeOR0gVpCzCyCJoLF/JAFOa6RfLglNBEg022ZvqIJEsaXayZw
TzjLEoJHSBsdU80amZNXfsyVeBK5jo6VNp08X9+iQwQmHUikPmL0prbcPmEk4SWP
0506KrK0uJ2IygjZ+i1RMGcfvmyty+28EjM4Vg41woU/BXtxLc1E2le6faZWbVi0
4DYS5VCZEQNY9ABdpLWNCzqHtgMrFiYqCrM/fqqqlZLvQnzCv/4j7TQof4ryg5Kv
eg+6z9GdZoPHuMwkQaGLsPAt71PVEhPNGIFw1CcwA1GRG4cnmh5ZvCtT3LkAZaib
/JIxjRHUSuvNKNdrvlqMWKqj4QEmagtofiCsYzpnAwFEaDOOdzPk9i3b2WVQjk/y
WVzDpZbS95RHhEe1xQ+fxAkavHOXHuzRmQjIexopkl906IQvmy/Gkyq62Qt2fDfG
lUWR2Ng3WCnZcgiExTyNL+M2eQyCwzEFx6XkauuVFJUy7wsolYsRvm2RHRWkTrA5
`protect END_PROTECTED
