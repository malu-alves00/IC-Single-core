`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
g3y6EeXChNBhzqSQ3dOoPSYOb1QzC41uAXKqEAE+ms5RS1HMXlw65titsXArdPlQ
tcENSCBug4csi5PE3HUOigBtPKCA6WyDlr90VANdz7rEf1wKlF+Ul8f63+dzrn1N
5UxQs2lpg8J0bno1tvTNFPKsB3zw8OeoozdJFPzWGkTxpjXHlaoJzNTnydChfaFP
8QY1rtoerkDTzoEt2NZOO+w55jShUnHO6qW2Mf7ia7KuF+kXaDrhXnPsVg9m9j90
0EJ1zgTrWtOzuahijlHtHk4evxyNBb4EC7aCqU82MVEyV57xnvk0HrnyAg39ugri
OMFMQGxQ2/jbqwQqbAnCbm7W6J74e4a6+2Q+sYZIux8=
`protect END_PROTECTED
