`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MTAnJHlVNULH/t8enaJRK3eTqf7PZ7lJmobCBAoEHi4wZweFJxmY0uPzhZQhsusU
MDCUbeCD2Av7JZHQ53uWbpErHfu2JKN2jygwWlt814smZmgbGXsyDjuwQiuAavOy
D8iPlPndQeIfz381HytpSFaxYscy4F5gPVv4XL6Ob6XJLeJQPgyR/LLwiCZib7Tm
rOqJhIq5ODZilxchr8dFSwYemsEWlHu48W2jZi7t3WxslS/ulzJ5Z8r8W0z3iKAY
7ml/M6BWEb+gLf/OUKuwofLqjxhyv1VISr7JsnlESxp96Lyk72JlbASe9CArA45j
Nujqr+3nx/QzUrb0meavQwFlyE4kzNTcHm63Zl/a3JA00Y6+MFZK9nqHO3Y54eB8
DLPHe3c4KxvrmqgyF7+x1PGpAWUjB0t1DBYUNJZep5pGWILbWS56vNQw7S+h4Hg2
4t4lxFDkxqnu86KnSG6M4wJ7Jy+T4cx6l3RAZ7HLU5zWzY1tr814oa8B0Qg+VKjY
yeG/d4zncRosV/2mkGJJmkEU0FMiSQTuCv+m3Y7R10iDMJ0M/FpFYySnNGmJXRJ/
28eZ1HFW9dSut5cxmB6VEGW05SFPLX8Pcwe5DrfiqQ1Ur4RFBevu8S7QXmsOzgop
aCdguhxzH1VTlfYOFr4I6FD707qKt79j23JS7a7j4xb4S7yi9EZhisiKB8T11kBU
IfNCoLDRAay4WOp85Cw4bDoI5CKi8mZSQO9qiljUN8JqO6u2jAg8//K4bPfkyOWz
KkCIu70FUkeejA9n/HITd4tUDlhjC4Jfvzus3GY+Gf9suApYcYJX/mJ1drouHLgq
3eB7rYSkYdgHRu1CHNg+OY9moLQe16Y8caQZTym4pH73AiOqXze3LdgyIzBxiyNo
gCHrLw+EsXMF4bR4hbZnDqhlADx2y8gzGXTnHV/9BMWQ2K05r7IoNwbYbGm8RaGi
sSgHuUeWb7B+dIsp5dJnYG1E25MXrMzjmWikigdD5SDQRrfzoah33/db0ez3U7/y
SIHOGJ8hAgKEsSQAvuZoCHSpbKVr2Wup4k9KQN6FH+y5TNSMHcGOGiF0v9qD2zXT
zgLPuym0JXtDSZimtmuPbIl7tDz2R3LwMXEl3D5zWpcrZWl6gRW3OmIfJjQc2yQq
6o4uyo32Lg6sc5/kuepLIIOCSBKPmpdKLMCnqgpRZFI7BpCKYknnA4HW7jYudjfn
rBs2ppXikxdQyRGFIFxvRWlPcenJGVFRaS95TU3SX5LjJ8JOUGu0cqc7NMRYL1is
YzXuyxbRxo6sEJsWQ0q3hDIEqaTvIfVv0hkJq1baPePOp9RYszC7cbyfIg7UTIBI
Peqv0DHs9rshzQA5SQR9SevecIgDcT9X59dNGmcEjqmHPy8mV+scZgJREuVlt4zV
9/K2lgKCAdnVmG7KaQKk5O927t1ow9aEbKUS5jrPMhjjJtNNMcsrmrBnNkfTPapg
S008gCz1f51T1jxPOQm4dy/7llz4i40gC7mGRiV11rB7Jm6zvUygj2V6DBPSMkBy
Ic8d6UEvll7gFIuU+758JGVud9RR06y16swbzWw9dwU+RR1iyjg1EuUj3CA+FUVu
ytL2TV8bD2mz3kLQ4ezYyG2qb4McU3xugPxtSdCfWsCARekPZKPKX7ygzqlEyEiy
t01VczP9hUWpOBRdbCxtK9ONj2kW8mcvfBIhvTFUHsSJlQNWlg7UpucM6uTPTxhC
jQtRQzKlepJSuhF+5A49UBEy1cACZVA1KyeR9q7iMujjIfJgLJHJd0Jh3JJCV670
7oh3whuDyS3i7wp3jR34z1CAuNL1nugdrZ+LfoMZ1ARE4j00ea6+qDlfV7BJJrQy
T1ljoGjlJJ5Kd1Xb80jB6Q==
`protect END_PROTECTED
