`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nOmuFN4kiY3v3JZ5b5kRRIjYjogHTaz6CD/eBHisUkeiIJ2xDfGC4Pf4nYKOtKCp
ywJz+MUCAiYdWRizrzSr4MweIBwGpxpsA6f7jDMjm/ixzlHJ8trh6GbvLRCl3bPL
12Enra+ScDnoEX4hvfZaAOWoucxFpJlT+sWrBEi6gXOrk4Tv+mhhyIzfIXdaWbNu
VsUAZa399KgGc8vfXR1+mttKrmpK7lLIwaCcXAFAKxYIJ/IryOw5Nyve0dom0CGA
uxzFdGBSe3RYVxB5pI0DczxZvwsJrgj0CHn2RpJLBjxMJxcl9D3DTiYaIo99Mu2s
H+WsY6iMxYUnP9DhQSfSkWEOah8ShXIn8qicQs+6/gFzTu2lhBKTCeDTvBnNfftq
n9r2bgP71rzyRVobgVy+wSHDYI1TMo7VJId3QW7VpWmUjTYDnOrsLMt9RuAJkLBS
8gSxI1GhX+CldmMt8+ZbcX45yw5Mgsnn3/7ektWZJmTK/54jMgc4gRbrrqI+nTvI
8HfGoRXztZc/iY49PD1XaJOktO7dRH64q5iEf5ykFJUNRJqM3df3mcmFrnFF/daT
GjtChgNseeA7UIzAfQnbkkzUe8I2BHUAEdfEgXQWUqu2+0xNaV57H5qfyrawJJnL
fDx1rZhx2w7In0VkwD2mgnpQPy+N/r1kmnll32Np5LGhZw3Kww2RVK5aZVKZ/Zuj
lBIaWGuTXVe++Fbi+W2FrA==
`protect END_PROTECTED
