`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ut4FbB4pfmtevwkW9Hc2SmnfEE3ctz2RjzAenOCBkWiPs72YQzOOZ2/UtqE85+bI
22X8e4OXbDvV49oeZEOK2aLet42C2Z7a+uVXPZHP6nBCne2IeTk/kHH1m6Iqsw3A
ouxqY/ULq0xnNMtcaVYLR8qlRRM1SmDW4AsIasbADFVZPlbROUIn8LK4c7ZN9e5r
G+8zj86PFX6VwstB6V+/9ACPEeTjcn8Ga1aAILHi7vjJe6CZOuOirI2/nXxCfwek
0CAhwyvOV6TXsjWbhe7wWBzLvVC7gj3z8IPEmlZQUG982hYJ+6sY3S6m3s0y74Q4
EGTGtjjo4cUE4+FI0NH0RlcEwl99zESR7BRZoFv8Yx+a165ucISUGYPFHBYEvsMm
BABQIFMb07q5GtoGGnFiyKp5NF7l7vDyRawAxQKh1sxrA2DrjQWMQWoEDVr/gw5H
+aaoycF8Gixon0rH+ESlyDkXyKU4/1QREVQL4Yy0U+zuHMcVnT0UJ7Viaz/1ZG8Y
+BmPqnQPCnP+sTthTgqpxrLE6PA4YOTkeAElCSa7u8UZvMinY5d4WLLX+lEjXh3l
09gVwQFPpDJgZwym+FOIr+rNemLM2iMpA32EKP6TrRT+SkxAco2n6ZDCpdP/+pqA
LPhE5K2XBx4Q6aSNjI0EdAmuoOMr2n8a+CDNKyHToL0P8pC9B9iIRScgoEJi1dvV
h8fzsWHmzv5ct172hsXFQYRcpdbrwb4H1TKEtN6btdB/UZk7PWy8qWrJWHbOVyso
QaY5iO8L6IJL6kr9SdIXVHwBLmLUX2FXZ/8Vv7CcvW+jswc2RguYr5+yX14lc+t4
QJI6wL662jNbFczGEVPRBxQ8tRfd7ASuNyFKimzicCgSn/Lk4eRQx4ae4TnPx6VX
Yl3coIj69yzbmMwTGHrkwJmiIOhXvUEDdCKdd8dLHsKFfwNU1rvtkjpnGCBnl67O
nXtqDHuPD25wrsXUfZofxqoXW9zFlnMsCMsArRhYds9xGydeKR0DFoX6Jvbpdg44
qmnHcZ1j1mJQRF79lpS9GldnL/GSt9yAD59RqXzL/zWyEFIMl+a6Gv4Y9WW49Dfm
Zah4IWLiCmRBZyx0jmnC7t11CZjo9zAeF0faZQF4ww1cJY/RKzx6Li+/sZytiVJL
M6Y4++FcDom6+IztrbakIQ==
`protect END_PROTECTED
