`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UZW1iy/b3gaxvdzY91j1fMm5fb4xq3pxTIdl8ChGZmW5+70mbk6D3fQMFpVdB/Xl
FpDQQ2FrxN4718CzUd8viauIQ8/jBf55h2xBm6ZDaWefnjc5PdNS73L3kJ/iXAq3
paGbb7gx0JtjS8fsTlE5+BE/bmGb1emRNeGe8bZ2u/L+CDSeNAt7SxVi2eyMImRW
AAQ+oz/A0G3eTkjln+RvhF8ooqKMYNRytNXQDJv+KloYTzZ7c0S4jTVYhamJCO2K
6qbZjm8EMw/2jljUzCK+rIx/JMnYCeqdStGgyNXeR3pq7J/hfiXLVqcdl5wKwsRp
5uEh9RECkQzGVLWG0OkGHMi1utT2IRpXeFxT03jcX7FNKwpd5Hma6sO6/D2sHwiY
qUbEXvdL9SkE9ZrdSbQzewy2Q7FwHaRAuK5qcwxyo9OO23cDh+ckzJoU9oORU+7E
SOSkVe1DOcOXDbEKtHeD7aybkoNKb4Vxn5nCA8kCZPj3trugWUGzQsrJP3N0ECYL
pJrrKUW1NJatligiMJ189384QkMfk1mvAf0GZSEfNo0MmVC7Cl6PicQZOPhbzkt0
h4wLa8J/iPU2GfeSUR1L6QcBk0T+5aufMW6XPBOePTKM/bdQhJ6NnUmI/NpNsl5p
acRf3Tpd5Rnas1zUNs0FhEPQqV+PSEc3oluuBwnSFxlJwskOw0VCTJQrJllRnx+D
`protect END_PROTECTED
