`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uZ3+LHWb19DjAuR6NMBG0s6UNPERQDTf09toSRv9znmC0rs82K+Kbt3cbx6xciaC
3hpE6nv3KDadHVwmuTpHziZGevqvy4txt85ZR9DuNxAOGu0V156njZWEcDjioOfv
wxGpjMNvpdWIEwtX+vxNAj/f730kaF6pIcPMabXuZNoK31n3NmoX8gsAwQEZ660X
xSIsm6pMFnLZuNvKsacTxggrWRf5n6L71b3Y/Zw6MZBhSiULCquAgHxqC/189WU6
Bo73B5DT6oAjZxx4tXG450jz/RkEFDjVm9AWMezE3nY6hXMooc3/p8Rpn0hqO32o
sc2blMLBBbG23eBV3EnFaQnuWJgnz5J00LpEyi+Wlg+6Y4rSeHs3gPiwXe0epryl
Nvp3mapBWgkhq9f7cytChX+PZ+uRaF/MsXyTWrUevEuLM7nSAoRhu2TwyZunAZ5q
9zay0Xj5tnZW8E2B42uT7NGBxNBC/GFxhIpkEnZSvi8wgax6OZc6wpkArN/ks++K
a653jWkMDjsT0BTPc9z4KfAKRj1hHBzNeRvZuUiTF4GG9bryruAnKVD4jNlsion/
PpoCkCkou+PiUuF58Rt95r/68uQWFqEShAKJ3GJsREgWDPBEWa3lG0poG/JB0K0c
ty9A1nkkgKeF7BKCzKyYysV4FJloitsID34RNYOuF9+jEfepYckyhnRFuk/Fb5im
w8YSkBXF2sXCN5QPPoMAosQYVZ82IbZrIm7cWtD5m5gy+mao0HLaDQ7SrrnRcHmQ
F63Cb+rDYSsCbs5JvjxsdPfycoU8kPnnIHyjh9ltLXc8YzR3+lw6ejFaFu0S56zQ
lwxQUXsWj/SufeYem/29Fj9usLcO2VtINFwUFIvfxrcgzqJQ2z/14iMHfzS7aknZ
Gx6smeICBwBj6mzj22wbt8vqdWun1DFNVLSrXqOkRPH3lfGzVvKztkh0C5YoSuU4
mZcPjsTQoXnpVSWcUimTRVxdeu7gFQELJlwd2SfDAFZEqFnMqebku7OTuctJ5Rik
jWGz5QY1yFm73T5Wm9Vwykh/7f89YUXBxNXxlbNX/KkRZ2ZYWxs2gMGqrrUtARvf
kLxnyl76N6+MdzKDxJCdF+PABZ/APb18Ygq37lDVfMRJT/nuQ4qTZIxdUNbl4iHX
2gF22Re9suZW5rl5KCM0CgfZHQmj1ijpiImZwFl0LBr9ywbN91xTs1MtnQjAwRhP
XLNuseuHKc/h00jATKoGyA8E41snscX4CIRo7uAITHSwnTJt9Bnukhz+IhhZk3ax
2ddxe9YtrsO/MnmmEpQnLE6rnNLumz/95Dil1EhMb5xtT9B5Vk4Rv4MnNgk6IUC2
MaEhMcJcuMBwbilxdmwssOIHXUciVecXLJVBDx8dDPTNDTpzyhiQRjHzgLsr2ZFK
f3O/HrV1O997By8QXXDf5vIJ2/m0yVrKXjCBVF7iwDkzi4WtR5mIRuPUOFMTDuD3
PK0xqNzoJbbI/nNIvwW7QYqdlbG8eeSauO9sm/1iVgPKuF+BwRszJBZdevZEFKit
eugh7/3uxBlF9brprc2jgqcpWnnLnNZ15vTD8uDrY3dfSaNQZFGQUrpjjYe9kNH0
4fLGIR7LlnFY1ifuXeoY8BVxYkijRScuEcOjzU/z1oiRJ++ebyvErTHfoxUtsJhH
T7pmR5OeyXWB47Skp43toidDWsGbtGmHTx/J0YDcbC/EAbrc2GdhF2ebbrJQHeSE
9uO4jzm/z5AIrfVbK8Ju/+uTvC2qLbSwK2oiwAimIxsBJVIX8A7z7RQBRu/8huQc
v1/D5P8e2UrXOgHTHnpXc7B/IXnk07qWSOdksf/VSZR3DR/iKVdWWYp2GTiAZdt2
4ou6fDo+NwFZENjDDRDDF4+oe0pqTAQIjmg0IoXVQb/0o0WS79+BtrZR2E4lrkCq
NUqHsmBI3IC7nElhmaABnD5/SKzebBTv5LxiMso91JhSP8VFVVr7/cCaYYpd1cZG
F5VMW6T7fw2NCSciNPOyydq3twp99qifySe6EYkQShjzlx4BMw44COpU8oAsAceq
gImA+caOh9GJEMq/6CJxvsh144nEEJiSDIndk1DA6/+s3THN1zzyakPrj47jKtW8
Yv6UCYS6jziVzj9K83mOyJbXorochcwe5L9cmuchEfElGwwp4y8mFJHkzGU8Fd5H
17mHFdLylpmWjR6Tss9w/CXlry1WxMu7B8kB7XFCPzF0B6Y6JmF2T1qnyRpT0QIi
KccKvNDYiLowbN9Is0oqXz6/LfRdM1LQhlAdJ5vdlaolOpo+p1RRh8h7qOp4O6Ex
QtwCw8HkfGgx7AcjOOf2MkjhS4zZJkKsuawMtZ2B6eh1J0zXpLbl2vj8BUKtMzd4
56HvulTYJBPuLkE3xu31o+8YNTTFXxfVTpF4+NeRRvh0MnqYqQjK+iSo8Tt/2zmC
UhJv9juDnsdVM/TBjWUju/2Iss4bHcP69VPehqMQ43G3gI2JtJ4zhUtye2Q/49v7
rLJ0SHZo1WhxR+bwvEzcuxbzjfvg86Hd2Pdhzg9dq/9IwEdm+BIJYiNNiceSG6FZ
0bby61lHQhoj2H4+2OG6aNN+X1nTn0KRqVW+DcFe08Ab4Cy8/g+47VpJVVadOv7W
r+7cRO8NEjLDbyZo/Hk2eDtNgF9GmPG+Ex7NS7fXa1VX6JhvZlm83ygyYiqFRlLh
OpN+bZ6e49J4HDkNmgFEd/LLms6GoTtoSFEjE0+fYmMssd+7qVCMrCEQhUiCjtk1
yBvbxdVFlQw5DJ4w+wIIzPnvyvh+v2i1E2T3lPYrdYB8NAPi9XTwzB/galES4pbJ
NuzcMNybYpa1ScyzZpsAFfkbXJnntwAVRSAeE/gHF+R7TM3L6Kzu4IHHj/4kvS7P
JkLq301QvjNYkE8PKubvSq5ch2jJcgsqLeuhwWEaY7CeL5d5UwsVFsfnVE9DPAa3
w6o06qwMIG9xdtRUY2tTdnTgepflwzlo6fhXhQusHA73m78N6SVmKWJ5IE3DdaBv
JqgDsunmAp1Y0qxerf2T94C0x9XGMFrvnp+qmU4bqzuvTX+JjLohpAim0Ie8ns1r
pHfTFoiEb1C8FP0pRfUQwU5WYECJ0WkcR8o1UyxPW88m5N4fosIYuEV5gnllp0rr
2HPqU5F8Vrc9CIuiYj1AV47IH+iOqJ3tRwt9Bv3B4hblUPv33XFe1n8RfFLpkfZV
R4NAqmjw/pdvC7B3SE10lT+8/s+z4RlwvmgIzzOZcUP8vqzG9ySs/AWfkNL8lc+z
T+ahh3QagnnG88+z+WXBYJ56XhL5X4Muw0KQMag7Ry0np9tqnorfjCPvPQsPNXeU
l79fVL7WQLRqfzqyp1aQvggIlGN/3cyp+ju3SLSnsRjvCC7fDTbzdG2wVg6pbK/4
SpG7pJw/SNXPiWC6HDQkd8xfYZjHE+HYM/bgIkXq8wyQB/QzbIBzzD3NGT7TypYK
wcOotqQgGZL3GRO51U7c7U4nfBLm/RupWUbpAb2gOwBfQdpbG9bGhkHqSe5pvprr
GjH+r6JgcH4fv/t0u5AyKjRDHPajL8gbGyyzjOa4GOWr5e/BUIUhBO+SDrODX8yf
YcuSnK/efj512GSEmxQfyHnm0DJWls2dlafRRy9FKd8BXgFuUGtIX4cbsaBz284W
aWFApVPgtRXK6XoG+Mgq7KljTKZxLNhRnJsnidpEcCJsSzAKjQxMXEXzvFjdwNxC
tQ1la4n/ejnbcrvUInncpE74w12V1YxNwV6F6ls2ISUOnme3MtwIfKeynUSMmnXy
Niv5y9BdZ4M5DZbX+ZA5qd1XAHcJONOCLq66givFcETl5U3KaIqnIyGIlgFWA3/N
va4BtjgTiC1cB/SE7XthwQo5VX3GmzMEQ0UeijSoOe0=
`protect END_PROTECTED
