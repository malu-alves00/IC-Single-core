`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
frwlPctCbiiX+oyLXfIeKCoa7jw3pfcPRYvE/Qyjf5/ngHYs0iXeVbEGCoiHibEh
u086H6kneGZ7vlAij8gOpRCDCd83TwHLF/lrfFZM5r9y0Z/f761wacPj7UASyH1P
Sx0LBlnrz2/WxP23N+2t50yg2W1e1BY/W7++5M7mpci+v8Mu3Gdyp1n5ktYDB6B4
783kkYGQQCw0Y97gXPqBRtEzQKdc5LUl5P7H0w6G5xXtyD0Qg8vVRYeP9DEUi7Cc
OruhLWuknyoPmb/DORf0B/fESBH5DHGnZTNiCYXr/M5brjLMV3o2qNG4jzS77lHC
dw8pQGKTKRd6hQvh8FUVrQMHYGMf4t3yNGSPQIKL75wSzw+joFwXqCkKJn8k8v4/
5BMR+weUH91+dxia7SVxf95I/Fjy1NBWBe1mBA8l31LhwmpGJ5/emEHO7cR6mcLX
OkXw/q2wCZfw6RxQWbGKM+2lP6WSck7MskVBD5Sr0EhG47o64Xvg+eCzIi7ss4BJ
z0eb2zY9LQO1u6TDCrAk3RARD29olkiadmUWjU3kHynLXvOjwexPVODR/TfuePAB
tO214zQMT1waFuZePjXcbZdBUGgOfERrE+6K2k72iz4Fp4jPXHumyyv6KG3tgLl+
d8w9RbssSIvN0rvnwRqxErvi6N/iYgAr/k6JOSQoUMylZCXwHTBtNcJ+LjN89F8Z
rh4sGcOVYs73/BCPSr6AES7qQp5ZWfXydJcahlHxosGe8l7Zayj1yS5tP1wLQxvs
FfW6L0/2iepYS9yBO9/zub5+tqokLHcoNGQ1mbcLg/ra0+GzFzuEttOTDqEtI9UM
ASBrdoBIUPTd/sLfJk+Rm6FCajjSr8qv0Ou/kqF5Qm25la8jW4x1D0lnomhzU+57
nCWk5mFW96BmzJK4dp0JDghSpm34gfIinkWEWYF4Qp4CTjBGKDLXZ3UbxZgI9Z8s
UD/RpCpqp1RpdkzsraVPsp8FZNuRiCFI3ws0Ng3MjyI64lZQziXhyB82gEsf1wa+
MXBRxoguXD8KOtMX1z4jK95gOEeZHNyCjgtc9SxTUHIz5ARGfPz71VV2mwYRotwK
k50guXx10AaXIy6NiS80hxV/PnqaCPptjegoGPXJSEyTPHbMSdCPsx8BwIBlFf78
InkhCdVNBd+3WnjYwvI34kpcfbm74Z+4FnvBUauKhQHcIlHwFdVXwvNs6+N+Czus
NDBe4R5UMzbGuJ+1rA+ovH9dv8WuomYZbM6eV0t8eu2zH/T3TyzT7i66paiXtz9j
/xdKyAfvq9GPnFXmxr2SRmq3sfvdJ8ypkSfBk/KcMd02bF9R5taBAM5YA8UACAJr
7caotrVRpJ1YQbxL81X75MbTCvC6We1qqEZoTVxTGaV8pgAWYVYAcWIyQzAIZqJr
zmJGD+OK+opcn65Yqq7OK3tILiYDHySAcEETwhvgeHDWkOXhN2L3vg78vMHt5FUL
Qg6pZUVa5xImikiutsZApy1Y3xQ3aeSXGJDqwMiECgC7qdjEzdSZ6cgZm7nQuS/L
/YeKFlBjfCz6SS5z960npTNo6rkws2xny4rwBmjv52jscFdWobAt1UTNtEJreAGe
lf5rI9GNZxzGpGgvbMaKWKIjb57UtBW1P7XjW//FKU0cuF9aQ2jzWEoP3vzBXDKL
t7iAAzyx3FAP/SqoCxPIIjGDlSZU1hocvUV4YvqevpzI9UX7BnKewPGW3Ym8mbnk
69ViqPDQ3UjvYXD5f8vQ6vlBYfqL+2A8XMsqDgRIombNIEubyP8dvYTaqZgPxc8x
sV1o4nAP+ujra0BJh00LQrOMYIuMR5fYsUpgQvyV5aXf2Ui8zooWv/PG/Odo89ld
lq43VEE12Xdgte4HDIBQL76iQNx58AVoYJAAuRDMwq5CjZFgYN39qPNFtoG1HOXG
SCpFQUOw6z6IXi8GisnPLkVEvRVefN7VK/QqKGFJWh20ChU1FQcABfCBfBjAx80f
BFlHqSlJNQs6iKnbgzgPw6QIHHEbUI4Nm/A3sC4IC46okM+fXBxOaOps+FkYm34/
anE0usty/UBGj3r9BtuUFn2Yv+HoOwd1l/VIvM3eRpieTOIlB7cpMSE0A5afOlji
NL3sKv2AXHS4niI5vGmPrAxMCjntCHNVLG3XEylGD3/It59h6DUyba/vFeQ7ruyA
INlrkwG8CTm+ZOef0slZvhj0wGS2XulIyG5fqpZFeR1BA4NOi1E7urmyQDX2xsyF
h1f6ixvjHK9SRrAPGdcwlAOar3hl00W5HgkLIdVDSelav7rvR85ESf6Z83/PMETT
VtYIhusY5h3LG+7+Ho5Vu+Fa55fzh6B5b/8cP1/vAV2c1RtmKEE1jOi8gxOKtVnT
fzR2e0MYCLUaPnTQzFZSsbhz8y8Hg/gzgC0X6jzx3mQT3j4OCozurkGeTgKVmueU
a3tODA8gg4dAyTdd5zqLDJlnyibU+a2SO/mhB0LltllzggdV1EtkbSiYEFzF/Pdp
EFZ1fKtXcU1R2WGcti6YKN5W4xx3GJ5X8TtC34C26XjF9MXxnkx15qwvP9dc1DiT
kvL3W1tVCXq9EwlwATLXmNOV4o6jldVbZjKN9g+FXs21wZ9cxAAoW4IgRdDnXJdA
4xRdwDHlrgtD52kOA9nSoLHm5JCaHiT0LSwUHEHtkXDyyuOZTbHKqJSl3LpIcZQt
PhgN0l8Q6xF/K5XZFSZ5YFGKYFapoqkkY/Oe4s8lBFTFITwTrcFFOMdDWtZwURsK
2nL8PP3dzFgsrs67bsJGr7iuLgS4AuJ2JxrTncbu4W8guZQSeJ5kwN/oOBpqjny/
`protect END_PROTECTED
