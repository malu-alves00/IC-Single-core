`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3qqZL19UfV12Ge0e2XAJksmNOsStJyhIwUQSMumXgwzdXf9cprigD3j69wlr4jmF
B0n9tkcSc4h1pFsefQml9lRz2mscFcBC4FFGZ3uDIN4+4OB0FWmVxlcK/y6w3R70
iqlxZN59tMGNB6rpCeZQ6GRRA0Tt5t+i43UaDlAetEXALLiHT8Zz5lZEL1hpYsk8
qMBqLap0YJpNDuFCau0sQLZHQCbuJyp1ocRp4F1G2FqqPZz+qgyrxiOOFisJyqfo
dgQEKBAs+9oVFfnHkGMcQElz8VPVtHREiOcwopLMvrvGLe6jLjFBly16328BbPA8
hDUycRUs1W+teguMz79Jf7Rz97vj3bkKNj4W775cw6L2jwY9+6S2dAB76G05xTHQ
+zRezr3O3UC/V+s5NquQ98rrJJFHRAM56UvgY1nOaEv+Qqm3OejEitQ8xcdVsVKY
Tbkdi9YxAki7dq1DWwn8JoddllkD9xEFciYCEAm+thzlfNxNvmetdjd5qS/vu09K
tF/8vIo44hy/2p1U60+6+b0IN6Uh5O7F4D4gQzcuk5oqSAJ3LGPVBhAIpgxhmL6f
zRD6V2HltjYJjhWmTapU+gXtftu1LUlAIQ+FMw5d185M5LmLwxaHCwmWXFKWp+8R
nW2Fj6v2GUuH6qh/K3UM3HuC/UaBthDV9H3ejpFKp960kO57O9eughDJZzWOQBLf
ZQeZPlW6XOAiJbSjJP0J0bBUKFrwfsA4HNVTll8lQex5uajKWk+CRIQEa5g2Bc91
RP2gl/sv7Tu9trD1JXO0akJp/xtBcsI9eaxOHYrcNtyrrD69mzsg/T0nZH1u1oRt
XCXXRnKvpX8aHOi9CrT5HVnUxBFwFVshvqz8kzJ3ek0zaFM+q7UeM3zfON5Ec7RO
6iHSst8p5s7Ds7P57XhRACruLoa9H1aP2wOYfPjP68s8eCllI65HtKVLGl4mPppR
apxiofivxWgPk3I9e70ml11tqHLAUefPWbBll4AlxlfzTPvGeriKwI8E6FP9tN47
`protect END_PROTECTED
