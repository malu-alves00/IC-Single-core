`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sg6ZEKWcIx6u7bdKNgNVHOWGWKrp9jysM49C7HX8RFBnPfXM3nRV9OU4mUSgHceX
CKALofunZ6fcumwcBJ6chxI81RYauTzDQFkxMjlSnPU38uP4Df7VR4c3SAKOy610
IMcitx95EsR3HdG1q4pSt6PskzCiEK03y3ErYtI7MbzsVnw7NvZCCbCqVBAbismt
mUfcDB7dLrWGHKNPdSQvB/iCOtwJBGuuZpkrU2Edswq791dV6pwr1bFyd/m3oPsk
I+GMxG1wPtMH0mEJfpAG3OOeo57pLMO6McRrihYlJEIzWT3wz+auXtdblRhM5Tw6
mPGkN/U4KwLvFXRd7HVjaaQUoEa2So+2ZwSlq9Do4TjJFwriQHO5lIfOxMX1VIWI
tUVUte4lA9mIMUvz8JVURKAQOUN2p1EBCgNYNK/sOicI8pcNWUNPVPXs3yAVTeM9
sYRE11+hE3BZTqRwKnpBNpkpSa/LVAj+fTEAqfQaDrZxJKNFqkneSkuTqR7HSHfI
cbT8DZwK8CcMBHEBYLOohrATBb2V6zH7aDbiXqnq9V6mJOMXCfTDtFKCWW2jkrrt
5nDpXcJzw8I7vLiAYL8xz/S3MH9Rbt2xBZkH1ogcokooHcPWZz2WRS1foc5fHWCY
0iy6I+qJOlqW/3iFKl7ysWGmGBoaa3WXg/zPIN9HzfXeyMzpADmhO+k+fKt1U87Q
5uZjS2bcB4K0PJch/OHzdVAm88R2/TVf86j0UrHbJCNquprN9tx5hFfWY1Le3erR
BRgRQoe7F0NGlyhBk06Bu3HJV28no/Xc4o8FAdqRY6TbJ/5Wqh4XW33/0Rglk1v4
4S32NyxjiTIlQi5mSkihJ6iekLY8Ij/wuWpHEwFWl9klKBBPCCzWXZuVZc5nLkuF
TN5Dg5WJmRhGE+cQS0I6TaoF1Q8yaNFGz704Qji7tvmV4w4oClKpN6huz1BhDt0h
UuXuT1qPqPBUAzCHFL0wItco81r3VLrFHpXPs4uE+RUYlqqk+F3OiV8+2zx0QLuZ
X6uZpZKo+5xT3TCnpfsWOUzw0MqO/ondA99hPdtqv1x97EeG/mJgTCOj/o5YMZQy
lzqL5Wq91VyNHC5ENn8cwLEoEfpiWk9SdpeoAVpGL0vi0vi41bxia1ZHo4vZZjly
dU+asPfVRv4EwKRX85X2NzZ/mOzLaKtuioHgFOL731lSI2IgWOqQh7907uP9sJk1
xrveRs9/POPQ7z2XdvytuC9qpmb/cqGl3Ffy+/8uDWag8Nnvh2fkS2iHhHWnEOh3
WCoZTNvaYuh8h4AHsF0e5iPvu/PFmVuM7mLzcCB/pz2de60HejamHKagTpCXJMPy
anvpkDcz/fVf+HcglUDR5Cz9KI5wqUSgL04jeGasu+rdGuBdpaPFWyPkcG/DyeK3
UheCV+fW9UJ7B/6ZMrapQScXlNiM7nrIdrK/2+a7eyT//GEjUOS58h5LLqXHdfD5
Ml2cmlFgN9hlUfM70RygWZrbW2ohd07unMO6fIHRkfHAjOR7Gz1vX+smVCLtmgIR
2pUSmVaZEUD6GI7lC+g60+/G7OTEKt9Zzpmw3QKjkiYTdTO5lKVnssYd8XUsjK5a
bbjKI5SziyoZnULmzb23TtvkK1jZDjMgWEkz4OEp9VD/lKb3JZvlHZTFiBfYJ8yR
TPdmxRbhCAQulpiF92yIcxcaGJKMl015/+gCA7Yp+npTik9GB3D32Rd2VB8Jocxm
9KfRyoysiIM3bemTP7RPQX562FFyndkcqpGxTCJxDCBb1yp0Wob4veEhtBYDijSS
`protect END_PROTECTED
