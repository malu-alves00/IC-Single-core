`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
I6gp5leReQjXo+jwdkLzUnSmzYa+KgZR2yq/7Zkkm4avxDk3gO/9P/7cQ2QIQRf7
O32rOiin3cTWrtcEfdEwWj6gAPPKuk75bIKjhb6p5MDylD3dUkp1pvW9Qfi6qyTy
iOHSjEqEQoDwyC4zo5pjhCNAhKGrmBhgQFaKp8gac78ntwuPTKlu3tUj0Ft8OoRM
1XykWhHrbJ4I6y3mb7RmsMO6sFmkynKN8EL9rXlrHoyy4S5iu16wAofgKYYpexDn
ph50uQjSvlyCyhbIsFfPsriYVomI6EgpoAqmt2gdrcNOePT1WB9ViLJUwfXoLSiv
Oci+q8hkEA9Pds80oCD0DTh6w+j5AH/gFiKd8a2PKElwNUvaf43id44zJ+q63PQv
FPiW9vZ5xZH081auTCRnX5OObgXvlW/QXhBL8iUwhZOss1W8cJehPgK86Khxv+ZE
tPzNH4zQTleXJdCiTZND2rx1Fz3pF5rt6XOh2wF0Se0EVBeN57t+n00W2KUdJwdu
EUCCm8zi23pdHqf4BqdgeRFatJQeuQCaFGxou9wgbd9p2qjbAx1OFgnN4NHORc+W
HCgGNADwH52WwC7av2DRP2i6D8NnvCTNxyUgnkFJnNJ1pqdUbrrJQIYqOi3RpOvm
augSBayX8O98K06zhae1ogVHykguZ+r36zUIryUPK/M89iAzXxCMMZAnaoda9P3s
Nv6cCzYoOnq450xuWONcAbliud12e1dNf0hmskWevFvC6YcJBseos9ijr9PICmZv
8KEEc+4RyTb8DeSr99BvIQwJTBdX+6Iej4eZvFn84s6ygMR8cEWEXzl2Wcpr4I0z
H4qWsnvmh+j6Xbh9ticMjDwJLGWcFHo6/OjJEQ0ZqiU=
`protect END_PROTECTED
