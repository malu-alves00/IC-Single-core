`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
x1Csh5YPGBZhoqPi4KBFdKPzR3WYWNLUlakHEzmZOgPvMgaRHDH4G3voxBEBdWS1
DrqDZ4KR3m0M8sttrWpg3EOz/WwfV7Pe6uZ6d42p4b7hGacJPxGnCEDg6d8jNlcI
ti1ruuDBPTwTTxwrzkmfPYwtlLIQKx0jEb3x2jocyPgKd7ZOi0Tz9ImHCxJbnNWb
gSRtlU+kmRghZNR1cleghhRAAE7K3gRTbZo3AD7yLztx67OYyFVGTvx5bgO221QC
QGsC4x+K6nX/7DC1Jq6NqeZENxhUayhYF8njcse43rds8SjvZfnxrP8YlPDVyp7s
yA+NHkmW+yp6TWUCyvU4OD3zRK0N2P9eZqQZ7BMJ2YgI5pRuRbD2UEpTgUghuzJL
3vp1MjFtOrC8Hpas5EuXCLroiPVpdg7Ztqz3Gn1+eCpG0wbXUT2/NaLEVx29wxWs
pmo2PY3GQM5lyqiTn2H4Blba5J6NGIWNQlWcLboOwPg0K/nNiZPBSyTX6uoDlYgD
OpItMYpZ8CFN4wpH1jr6UffYDWpH28mLw57n3/HLV0I9xmQTozOzWJUdqx03GT3W
75s4GFe+47fJy2mTJZ/Rb6SlTywAK0XQtLk2nduj8oGfexfK/1vm+DaCFTVY5L9f
7Rh2MNgxb56T5P8VlgvuPKz+OFLV2lOtc7c3BLrtrQCsGCy4vIT2QBtdDBpyxDBU
e5f6NHkeD+kF1d+IJyeahKMS7EfPOAccyhgc0fh2sgQWNmUoaNfJoCwIqBxCaQBe
wUaQEb61cZ/PTAAF6YlEAR5iTJgxBXMXY/bshmpGMxc=
`protect END_PROTECTED
