`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kY5KW1p5/JPZmSn695lq4ImHe+G0lfQEpHoDLKdfHILAwa7olkssJz5X0VXJGJBH
4SEByQepcaFWV5J/oJ+bsEVzuCXv8FHKUfF1Yn74sqWR0ns/HcaxSrnLVzhTm9Ag
gXkIBr3hJRQUj321cMzZZ1TmMDSAnaXSVvLhdy36yohzdKpCYrFIbS/qIPGm0VJE
5wnfTWheUKDW0CPc3DmXm5rJOpiJ97ccRoQzLdrIYRteXWM5DxrgvxNrTNdHsN79
0CbkYOV5exbz1N+g6Pcbj5rTVoR/n1Ey7rWi/pI5GnamxEH43cepT0GvfeMeuyWP
Qp8R21TgsNCbimRSwscwdqIpcHKflF3fDxer9axVzu65K801pPsKXz/hCZEn9cx/
lg2GdMG6qHS2ivZ3ApeUQ6xq+BVFEbsgkeLu0OHRUhyGy2eaYSRqfz3blDB0XarO
z+bNJGmI22DIrQRVVCEYBDkDfb0jfFMn3GIe375QcahFHR2N3OkxMpG1EKxjaxvU
zDsVKCcNLO4cH/sMnL97qCfPrIVAlDl+v+2JoD8HLUcnZ/qwF30p4aSAzUZP25bP
GtgINdN8ZCk/ID5C+TGsTG51nGT1UaaAJ9+9JCJgBuUekVYbGBoVO4AMD815vjAf
TyFSIGMLIw8Z+YDFAlXlG7quLs8Rl6cY+vH4ChF1Bd9P2sKdzXuXlZQHHfcCvS2N
gb9hvhoWKlGZ0VVNZge3J2gr9vwxn4oYT51qjcxrOFyj+imTN2WiWlv/GGmJJEQi
toz2IKu8gEusROtncXedt8C0pK2IS3x5enVCeFm17uJI6Peq/MDV4jdyRdZlhsgX
Li0lf158Ld1hV+lsK93l7iPYt+ZtIV3GzKlOh7N+yQAWXpI8nCh5A1Hl8lqLOMWL
07AYceKjg8/kI3ckXene8Gzv5mY4ZECg3clq6UIUL3gMp4s6VsnsvDT7t688kVjU
643EsO7mzLdeCu7lL2zhy2ll8yPwCpNIv/d6xtFOHgOMruC3GcpHnf7m1Bue0dh7
gpb8pNzTy2QFwO2D+FB4P6VB5Iw6+mYM0s5e2UcBYq9+RJMC5VspyVvdAziT8Y0e
YwxjCGjwNd4BYsticFhj9RZWG2B9q216loRLBG8VtaIg/vH24wwnOaX6+BYvzd4Z
tU882z0UT4aCz7l9Ld97P5++7iKJc0vqF91M8WWV1dPcQbYEhbujHpeTKSGKJfHl
iVIoCT4Fb+BJ1VTPZBxmjeCMKj6wB46iri65LIW3Rlvc2wlN2IX/ae3Ag0HmboLV
A+HrkI2UxAmXc/3cvwNuHtyDAy0tZo8MVLyPEkkCRvUuJleq6CSYk3AW3I4c2Xmv
8W7C5vY6UmDsfnf14ozqG2YpTKK3zpoyR0JGExxwhxnu2TL3CTAfWj+LmuR/WatO
g9CxtDOZCDKFaJ0UC4iYHybF3xTZbbHzkNqUrrQu4QPwoEbvkesZfmUf6rg9KtAP
wtBzrgBUKqaZT4wamguSI6FvldWlQu7ZcM0ektQAYw/rZ7xNI556R/55WfONBfgx
ogA73UkByctyEfqzPbEAa8Q+gbwbbBZ4bXCysKLf+fZIMWJaKg5itUmjF2EHM22d
xxeGPyoIzDsTg7QkZvIhKysEZHFNLfGU44TrANTBlr6ua91eTHpveVZBtQM/eF5J
HWOPOKMO0Imo+svqi1fQcsRMRVc+9bvIFBD2VpEXI7Sck+W/Fj8y/UXzYC6Vvxmw
kmyRhGJ08/+XUIyO021V3Zaxe5zfJ6+U4m6fwtx9mKgHx6tnCQjKDdjitl4YGvdR
CbfXMnxh6nfNH1dl7PGF8Xmk92MvIo92pM0gGI15GTVnwisJWSS9AAwj+SpF+jir
0i5O8SQUcQQhRVGZ+RSRU2Q+f7slvJ2xVWs4hFqEmPyQL8xJaYY8Lh9kF0g41IHB
F/IuUxjCvJLNpLanDPrTXDe7LmLcxD4hNhC+8MHgiLtp0sblwRg17t3q2gqxcL/M
ycjWg99i2hmODlJSA2cVTAlNQ7IWv8f+6K98QV6ivLYDBoWBbfgYyCeIJslAk+s9
dLykQrZ2574rlVFzTnKQTg653IjRU1Ze9oHGSf7jf4IHvQPrd+C39dE1SPp2f65k
M+Qkt/QcyvMwwDpwXzEycPL2eYOHw5TP3rgjim9FCP1sURS6Ff7Yp7ZR7gHiJDUK
3QfdJ4hujv3rVz2E+lEstWvIXm1DsntzSvt4Qvzxdne4dt9pdLLm6PSXrRXyc6Zz
l6qXnU42aj/hvlWuuHHKDiywD7ZpxsVB1YXE/eBBsRI8iAmjW3F1LSnny49jqhLN
NSnxsu4HtdobFKXsQkpZ1inWtxodbzjRVz/fth+nfB/tKSzYbXg6qducy1dSX1Qy
jl3APePjOGxdKqJtl5Mu5Fym9zgpSDwPIaDIbGu9bmcWaKJuecq7or6bBGS5uOYf
E1G368s5UWIZ6RFbQfB7kVU6Pzjw8c+LBiF0bwy/BQ5hRD4E0fBCdtKTjmHXbwdZ
QJOoRuXW9PjCOcrzM6Op5E6b40kjCahDK0T26MN5cVYIoJX5KGuHrq+gM1BrXKzs
RwjqcxOoJxwLkpCeOTHa4XsPeq1v25RqRI5kQbdpyCeAP/AdDGpenoBs73d0RyiF
kbDYLUnE0tbiCfq5qtp5nsveC3Bs3tbM6EmynKp9snDFCFBGmCuEKxKWhal4ycLt
XGkfejZxRFP6ucqdVPYE+s8z1Hgp1ALnTi+I10lcDQX+icU442CC74P+MJNHlQwM
gYoH6b3Nq9JUpdottafvdfLEmvZ6pkVOxtRhgS5Awq4RFVrhVgPO9952ginALttO
M426A/hEh39wxw6EzFRa99IrzSo1JifyhceQffUgSCUYMv8E4s88MkJXEE764VO8
YcAIk1xUsIxH0RhhAG1CirFSjd27NjtXX+UxbhiLrF2duhHk7lPB6EGVTB3WHaGt
637iJvERvODqhAC13h1qGq04KW8T0qTU9w14n9+w1JyryCBfi7jTY4sjhoWkVg0H
`protect END_PROTECTED
