`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6Z9C/6a6LzpqdYHTG9AOEBxistedYZDTBjn6Kmi/AoQ5HM7pz8pMVVkpMuTJ6w6V
WFF2DynRO0comVavtiv2Xajk8ZcGCBLed2JqTgBkaoOYHXUYDIXzitLLIVm0iRf/
/b60u11QsKOAO07pKf79lg6yvwb9sKSQATtptFuE+0oQ409UTcTaIo7n5xf8zMzU
JnhmVTGt58raHsK3dA0vVj+o6JXEg1m1JFbsuZ9Oy8dMVlM1/9wCNZRbL+ksyTHK
9YOO1k3kogbYXAeJi8iJJcuh+paz/c9yHA9nFf4HaPjcEl0Rl4Ozv4ISCh7PQe24
8NjFEsY0qOE231twEEvNnEk8eujGLNaQGw7iTmh2yd+N7/Egud6IqLE+Q+gIRZS/
fvLS/pzexHC5z7yp2+mV7VfpCmy+Qp2cytwKdFhJ7tr0AB//IaFPBRHUZ54pGec/
+78deZ6SH4NAMN3l5E8dzcZV34Cr6ow/Cy62XbbkCIowFTrRD8t0TJp33XeKJjF+
2DKTJOiv9vv/RObisYm+frwawGZJ2v1ljcq8DWCAMBVWfHXKWJqoe61jAMTXjIA3
E1te6Q/VpFHy9eZOPF8D3XRjEJKlQGeIP9M65xZB96QWqn0ZkEXTfSfu0BNNJaS2
JTve/OGXrIip27GeiJ3qPcOz/O1l61zybo2kFaAlRcPuxOrq8jko3Bw0+Dn7FRup
3V6He+PcuVDLsu0bOCEEKUjuhZEXRBB1TtrY3vDcvH0ymbaAeq1riVNtJndCTeie
Gqk1aR5TcYzKsIU5nHaCvKAoyzNlHcSlM1ygu8dfdQZ2LjpctxWZh16Q0VQj4+z2
EfRTdohz2Ku0oEocwXc2/5oDQAs78TLMN5HerAB3ti0ivy7oJmQoqiEgmf10iz8i
YRNS41wer65nB/Rb9BAnKB2xw31689cFIeyki707FI6faiGnePe436rw6apsNzKm
gVfcfnzXbYL0cqqbGmEliexW+QnkQueN1X83eqjU5DYUQ6+cuw5rCBTzcv+IdDPo
S7+hk1ZDw2+Gm+s+5LcqoGNRVxGJalPtUgi6Cpwh+x8oCZol68yZV/4nHdnnHH28
BwIop1tC5ZZAqyKqAM94KPFMcw6szpwqMUVBDjHWtumXE/BCsr5mPHjDGIQf3dsA
VvqdrOZbDQ6/GJ0sbTIG4Iq3uHm3D5GHUIyAATG8LpGfjlsovwqM0w83QikDazK6
lQWIgIu5UDCgDsEhKFOy1xLbJJJIf6a4jiiycs2l8BGhwr7hC+m8bk2TwLqOLZYK
ePlpyooJZanA2vcz3x4ncML5rYKKtcZBRekYWrosMGSh+7hNO8rtV4hq9xDW/fGY
ov+mIthzyAFbgG0QPOiGKQsc887Hb1IuvsWz+SQTSlHvUea2INBrXp/P6/Ap61ip
4BTy0mA7a5BAiTsCnDE95lBP0aE3GkI1t8KLv3WfCuNDTtlgdjysBih8bYH8aMtQ
RVbvYEejmZvQYXP3X3jfvd4sJ2JNZzFyipFHhr0lNR295Ttb4Zt1FFyy1p2dThSK
FjYcpbFl/Di2YUGoPt97BLJeYL7pX7Fsy2mXonRCF+ZAOro2blM4mh9LFsZe6iIo
hgQjcPE26JcdY4BNPL8LxMiEGYRrA0vxUyi/TAoQh7g=
`protect END_PROTECTED
