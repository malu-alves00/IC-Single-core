`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0cVoxH+IhKCI/IfJXmvmXvhZ1kolzroR1iOdmdPux6dz1UZYyd1rVKQ56fcL2lS+
GuiASY3mBQdhW07C2S8jEyTq/MW4TABZJ2bfhBM2R3YMdG+FoiTJHASOybjl3d8y
2Wwr1u964aTaSlrao8WxvJYTvktfP3/y6/fzA/zeenssb8vH5b4U5ndkh38cJ0c2
RyQYDULCw6GGqsa9WwA7M13oV9UWWV2gGtwScE0scz+OiHLDgZOGBjulk4Pe771k
S0qypuUKe2oXnBfdFpLFobyd0rdyUOXz3+4QjS8bG4uIGzDmPhUWV7WBi4O3Jd+F
ItvffP/OMBRd7MuXTb7NLXQbe5Z2gMZCQQzGaUNVPn6v1ugKaqEngMNcaB4VwrEG
6182mWheJ9cJXcSXe8PTKMWDq+JLHREh+QeynbaAcP/R5Ow2axnqKSi5oLQfiKFA
OnartVMpmZDht+uDgS2lo3yHPB13gaUwbywM6fKLxOCukGM9Q6CX0RCAxMB/y1rS
3MAdDcQPCJNBMgH7G0c24Wyt8boLgPbbDPTeHhDocsOEzpG3RYJOhYqmXREZchvk
/MyJUiHvRuSbgkqzA5zszq5PhlfpmhRxoyeTeeFTvObhl+uvulyekm4ZqyN72yAs
VzOSWUWjFz5YVAVU00Twqs6wjlHKpk8J3kr5wS1KMDpa0Ms61m1S1tbLUZayiZ6B
kmVz858V2XjhNT5EGyl79NYr4B80iBQnrBLhstz0L1CHyMpcXmiix/apLQln8K5g
wwkFh3tkcPE6aEp/vZ+UNWd6bpt3Lwtpl2MXPVqrO85gx/u9v8l9MZfcYm7pYlpO
BSL6Od9u06eRCZKS1cOl5PGHL6pdBvYTxdp4JLv66/fyjbInPQqctVfMB1DSMH/V
qDu3aW8eHqLkn2q17STlPzjpSyQqCt3jDoSe8T81ShX82n9ieRUlin27kaWIh2mb
rKwrB5sfCRDw6RsYXa1ExEpIdn/IumGHwSmI1+CL7A/1t7QUR6dPQn7LNDDePBNS
WIZTF8I5oZelIaqrdEb9G6uFigjwG7Q0RyPWaYvy2StQCj+zSCyfangfLh2IVWA4
LCscURf8VULSiYqP6Ab8K5oVzjYTDZpIu9n7hycjoTqEsObs+CWmIWSBcda60V+p
9XnBdl25L2h60c5KcqBES/sYPScHJ+iCuvYMQuLHZjWpyj7K4JfDAkv4fD/7FM5O
hzyil7SvWNXWy8mxhl/TFQ5oEfu6S3Ip/To3duu8zt/+9fgSyfNtIpH2+o100v9X
i0bNUZD0SmUOoAdhU+SJAu9P68kQySV6icFs3zbIyBcefEWFZQBpXsA76X3kan6p
eMRXjRthoGQldhOKx0qQmXSC++z4M8CZAmHRk961GMe60V3oGASi1Tkn0bhskA/s
H5wXzVP/bMuw+ZcfhJs9Q5tjrRwCjA3Kl5YgdW7btxJceShyHNOQIQKF97XqDGxe
hcclarj8tBRv7/IYCfIdrhvckEXi26tbFFq+p4NF/lB2vB1BpeNVB+Evx+rfWD8x
vDjv0Jh4ZCMmWFSf7DkJtaHeYs2NMAjRDEBjFb78k+CON7ueqnUoy4yulCJ6yBCa
13S4yIxCBxtMyoeq6k9G8LGKYeapN8WINx/JO8XMBVg9lIA9bUj43b/BS89LUQZ7
Z5wgrv8C5r+XBcBjun5NClvTMfvDPDDKWShzW7WsCWNzyw5kJoQGG59GdflCjHlc
h/ibPhTsnadS2IEJmzhHVSugLYDdy6JwkJ2uT8CEya4yrHSEqn6b522lrf8muXrv
jMyLNF+w2j0VcPZCDTsnjucxLRHt9o7gZgCD8A5L6SW7xGbHIZ6XXkRUHXEXKrTE
FbaBAXWakIgPik60Wt1JDqt5AI5g17RmFAwWDsOYZDrWKz02WmGTqu+gJtEOHeQZ
+xFT6W10Holr2kVNOMchP4/AGTfAQgi/cLqfvJsIHP+ZolH3Az+qHmHEHz3b88NK
uZPwkY0lZzWuWeyhgPkkZn/XuqUmo9brxvGLcjNbaeRjQadPVZj+TTez6RzZlQ5m
Y+yfePdFurJqBYQfSx+nKem4MShO2B7+ugoIBznzlYlmux0RGUsAL7KoC+XZqPg6
Xkn6OI2rJZ9fGS/Q/gcY1QXQR2/MKDAjrkA2me4MIvq8xaD60ezgddLYwxKLSigF
VSXMQmBKMzRu2ZHCbBPkj08STh6jJ/8wcg/qP/aZ7RsSzplucEbX+IQLidVk97Vk
zRd3Pdgnc8ClFAehIFdN1hKpuT+QHpwREmS5nqFXbdV0+nxYu8ZRVEdM7ittOo5Z
avPVw7pOgIzluqoGR3XhM1mEhfq/p3TtKhbetqpMygTV77AL7wTL4fncPtOTMlC4
60Xqm74JllPiKabmBaSZbhTM8k3g9cN1gXMsJwD+aWc6uCIHCbhmvK8cLvoeVJN1
zgrWFo4rNVbeycqN9Z5NziPlc9WMIXwxcWTEv/L/xaG8DSVLjI4mB4KC0c5jVrlI
B8L9YCSZWHlvN0N/MFOx3+7AoOwaOWvWgyAdeHxPs1k3UJNYtkmEjsFmd6VsCGIw
T7TawM3x8H0xfT/2SpHhGD3jAZLgpEgymJRCfZ9WrKnDgw/DAStJZBUu+a4gPPaB
QUGy0nFVMOijLTNNzIjY+Frj6RnTkUc9wYcY49fcZFqNuss6h6fmoO3DNbuAYleW
bXY/Q7qWHi4zvdWlnbilBNpSyDvimiSjPRRfzgSGojhPzPJqCxkRZqljHL80/OG5
AIy2dSR/eRHPxQlExRlm0RGp0XIW3JnBBcoTOpD6rntsA9Z13RnFn4nvU1aTyjXI
mURfeovU3z0or+j87cK5V0l5pPykWRaYkxik7LGETo6sZqC1ukKtur5gltGcbLYH
Rsmdx+Gy3iGc5uhjBLpChZ4Jq4ysFNTuPCdaJnhbZFNFGei6pRKhH574c8XfmOx0
hYks75vwXGbzP/ibFjRGDbrR6puhHYz+tQbTFkUtZ5B9MUwB9W+HLTnzaOseh6ff
bRMZe3AqUZRWINArRjpRFnNuyq7Hv0ILaNOGDPvM81hrAS/5GoD/HFKZ8vGxbt0W
rKUgKB+xgggBFuPxz6Uq3sqIK+OQwrPYQ7CtRtRSGeSk6JznwauVzxcsXGpEvnZi
adA9pyXorZXWbyf459AHvSO9aJdBO7BVxKiVrcOuFxMt8n9S6tdkdjAGG/tAjE6H
CYuqGptgmdNmRoQW7aoAMFRgE8hffG6PhH69iTHGeAD9nsRpk88RAlDRh9H0mWd6
4mOnAl3BuVJAjtBVF/iyTcjUC9SbTGV/FN6nKa1ZzEFxAb5vK7oxSwgS29zZBwIU
cvg/QgYxVFQtntgwEfA10+vKjnCkh4leR9pCz+Rf00s=
`protect END_PROTECTED
