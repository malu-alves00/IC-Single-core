`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yNcKuQE++4+1SjB7B+ah4HOBO0M+uAu+06YzNVlbkO3owvtY8ENWzbgUjiZIbL57
t4H4RiAEtGsA1uuJKD7xcQ8GWfaX/xmcpBTtj58EavAW8XZFoexgpdyvOzsqXPRA
D1MTJwNJ9EJ9XcStRmbgVljJfgtkMrdQyf+pTU1tYQ520cW0R7SLjxKNLb0lMTag
z/O0nLnoc6G0F2wNimi0ixkoUeeRjDfUMWHeNlZJ/BeBC4SEAIKKGilwOhGPcWg/
X0cHsyChaSSn/WrXwlXae9+4KXkefPpV+33cvgOws8jOFtVNmXRJY3cMtxBSZbjs
WJk7LEbFRMSZ+HVU5yxszMu2xRfBVeFWV75hQYkTM+dOGbC2WrUxTNntKmhkqgUn
rMWvYTEoOSfOTr240uwO2YHODHol/yl6Gd9AOg9LQaShr43ZYZYYmwpOt38Va+UR
gPF4u1W/llDNMtVwyJ74Dlb6mhVvbj39fC/O4CiRVEYxHNnoKYGiUk77UMSn+woS
au6nKFjytzdwqyY/3aZdj+KDLgvDyo+sp/Be0ppq5zIf/x3OoDI4UDsANtNJC1/C
HcEUctwdu5B3UcA2I95Ng4HoPkvDA88pkc27kp4EQ/a8kNYck2QG7tFMCwXnCt9Z
blbO/tee6rtuJdFD+McJ08c6PmecqXiPbmlLLeSKTvpdyEM3JryKlXCAnYhYSbWM
56WwkEMdbdDSC0y02BO6BtsJ6TxmfAeqm7b51ozRW0mC88sjQJbApkXXyBnA0anG
kEC7FOB2PPau90tzIn/r6nK2JOoZn8y22IBv6Mi0nNHxg0zLiWuOJAKF0EMHuTaH
4PLIDs+2qYU9PWMZ4WwI9EG81A3on8sUFIpu0pPKIkHjV78ntMjIobxDhumzJ/px
f/+zrZsRJmP2Ndz9aXu68uBAKhmes438ccJhzyJKhHn5oTlmo1TPf6jAUBvliHNF
uwusPBt6nzlPX6f7Mr5hXxZIbQdLS8N2x0Nas2FY+ZA/CzBvejuUNRi/92KF/2Wf
iAG6fwzTo8Z2Jlp9EUiUHTfAK64bc+/3errAo5l0PpwFDz8+nhSBczElUWuomvX7
1fQl+SNjeQYaJ2h8BgQEJ2vchhD1uoVgCO/LxYwQAnVvGA+WcODfg4oMy/ruit2z
avJMVaZoSwEQlRKY3XOYZ5YZ6o/sLhRd5UWgEXSQ0UXBXX89zRrPDdUOutcx3ZEg
t4ANg3vT/9QaNCCO2xlRwAyR4OsIiHqjd7jVUG1pENc=
`protect END_PROTECTED
