`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
P2u1qdLRIR7GWu2dpAb5zbs5cIyf0Drzh2o8NIe9KZfuLYupPuZYqZvmPQ/u96gU
fr+TRJeQK9xTK9bDBEvFK70LSNPTM0Pq2rGfNXYai74fmvdG68hoBtl5biK581di
0zJbBUknE/R8C63L28/99etkz9wOq+b6DTA6z8Fuy/HwB2AHzzGcYdj3ayWg2uQH
8qEveDNaUnJrCXQxldkR+d/EE8Ya3jrp9281DptC36ZkLed0aP5k5h2EAxVxuuj1
93sjtSpYBK7avJaOSFIusHtXKcsPNLDNMlC+wHnLGY7pe+ZeWu3vKszp/R1UHbp3
RMmhLLHpWu5Xbz2EoC2i6t5aR/IQUDF2FaKq12WMyH4iMjM2J1gsjor/2AvzM+53
TiW1WNQIYNclAIN8balKG3KWWpbYf42w8b8t+somiQXxLVzDYacDFbi5Ts0LPslK
1CE75JYovwXyldpuY1rJch0arMlEdn5uf4CA7VuHqM1NzWbWY1jDGJZ7Dfh+HgIQ
3ynzXoeEPdpUL7OTwPj/LCdHocEXEhCeRVHbVC/6qwlaQx0psl4XYRlOjfQli3re
KVhDTG/RqZVy3GVebAOoY45bnAb6hUH7D/UlXHL3S8Q=
`protect END_PROTECTED
