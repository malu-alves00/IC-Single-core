`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lohdQuF1Q2GOvRn3Bcd6PIxDxh9FiEgAZs8dcPGsJLGv0cHNf/apNL7X5NohprG8
/ieGD1/F7YzSyGEez8z4+/rX1z00TGdwcH/AkVc/lqR5Jmbwj/oGFDDopRAaKlCT
7JX8TE3bUyKKXqLKdQbTNxypvXrlJjszm6GcfcS70lIHu83An6gHabgntsYpV4CL
dxxKnuaLcM3B742ligVsCZ9ajT5s7eNMzhx8PJrqRM5DcjCLIyxApvKYzLeXbL1E
zlYgSIfdOi75SEsU+ClHKIalvep3eStt0tC1CfeHkfmCCBc8Kawnu/iXrf1QTrfU
Fo51GI8UJe44C+HOZj+sgltJCyInYkbRQZEzcI/s3oXBMCFOCbUVAbFT2GqoVtNg
9fGvtbC4AumLh9SEEsMNzrHTAeylZ/0YUqP+gP99tZxYBDf+TYz4UW+2/0BKXKdf
FvSvzrrLp5uzerRvj5qAhIZ0khsZrS7HL6QqQaZJWZWP9K5E6Arg4mJB+7KLTp7m
1zIRPVwRJV2JMcvyJQaz+jEVlUFDPAe+570nk1eHuXdTNATDA3GBrnkNQHqgyL8R
7wPn3GXJUjnEtrrLDaS0tn5KcMN/92tH2AHm1gxDcCoMHarAC1937o54YhjbZR1w
k7wExcZgQor76iFchT6Z/uWPmh8+YqXzByUNs8MbnBM0srZ8YwqFiDQ57Ul5X5/a
dBGHsAsaDJ9p8D4+wUMZfMIAb+WxRdkMTti7kikpAxM3wZTohU7jCup41uCk9Xuv
n8q55NgmXFKqXv4Xz1XzkIeFwb64NWaajHjuaAmle0QYQuIvaTbFu9ITc5eiiv/T
+AmaArBT150zKUYDwMaiGjePSpewRTaGt05i/+stqznra1QygFG4tv5TWIDeUJqz
m4o8vRi3tghidl58HLNXQnIQ/4wMsCcv7C7PKWIv9MAEird8RHKyzG/ud21VFhOp
RDrQ3nOWmohvOEKimRnSURRMD8g5IGjqrUVRoGxOi9g37GA2CtQq2BF2JTUZ9Gd+
gIr4FVokkAmITO0qlJO/F5j/obzfMJihLm1+GgVlmgFKnc79Td1/OGqGrgRiFtkA
F1W6G3Q8qqiExe+7sckucwShq7GsGrOvHYyBevASww6cmjnflUDkgSMIWsIomxLI
YeXvLDx40CERxDmSidmqwOu99+Sx7TGyQv43Hv3XovFmXTuiw6DUfIMfI+A6Masx
Hf6g1LxLh+6KC8dcCqkDWQ==
`protect END_PROTECTED
