`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Z1TRSdyMIZFfKDAVNliDl0tWlVzk+1LELPokmg1nH6/WrFJ9EaC5fqO1uy7uzL2x
QgAIxIGPpnhWR4FnVlt5SC7i/y2SymuJguKo2h0tKQlXH94fLgI04nx00h1GUXDN
/40dTlKKWEZBWPrsHPPO13vn2fPZGJz5lNPO5Vy6QaxPDuHOnxCcnF/jfc8E3gKc
1dJ5nHlu4Kwe6l9nPscuBUsc7MX4UB/mc67DzWiY4QhUmY5TI+/hkAE0LdzRkCav
PNAg4qSgDSt7D6fGsRlOsOaVEAr+Kwv5gS/Ip3F9RARUc7nfMXz3qPa/m8uLUd0a
HWnSiYtOCT9cC2SjvLQs2Ouwft5f6nYXfx7ZyF3w5Er+aqzxpeKgeOdpSl3XL8Zh
iM+ixVFLs9mbAOvBY619q90Ph5jHkyk7G/id4LORIzkRisGRzpM2QhxvMNFKIoy+
jkOSyYBjbZWjWHP6fxeLf9thWzbs2Fj1La4tzxaYokV1pMmOnln0pgBNwTSn/0+a
eTu6aJzZC7Sxmhlp/lp2kV2KWOIzFwSC+2HwLT9WsWQdZcEydIQltfKBE8Sv6Agg
xh1s6uSM8AMuJ/ANShM9UqELpyT/92yhFQAicXeiZltlgmkzY+x1AQIhPthDV2yT
s3aqlUKXkNzhW5y446jjWagaYjtShAoxmpwqmH8gQtvj0hsOh7kROlADizaDM9CC
NbRbBaMGBIrkrj0E4SwG/qNdr7YK1ulyFeAOsx4tRnbPVaaw1VKJQq4PS7frUa3I
yE93+CNkJ6P3Um6ndEwNxPpABwKYVOvGC2of3lXvVpdx/Z1EMw71MO4ahkBKydDb
RF33CrvdoUvVMnZ5CNkmfxPGBzPDJkO4CLQrar6yFPqy7i66W35mhezBP5O2iVMN
NhSDAKZbXDe1NHOyL4nPXJLx2CVYlTuT0oRTG5h0tPQxD3sqHgCqRFs8wFzlm/4p
cqNs2VXSbjqnE7zN/6x6rKsSGbDqFtQlE7uA4uY5otc=
`protect END_PROTECTED
