`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ndbeCPeO6I4CfZrlHxkSw+oMZVvtotJRaN94D2SKgh0y3lje2NsFazBSvD80vB2c
2oxndGIFbraNhMR9GIAUPvsckNdOzppJ0nmC26e0aEDiFkLxt3p5qZwHGVwbBRxI
6QiENf/+OyTKvwIlxfu5OkF1fb78gGzhHq0lf8dcZjilFE0a65hhsrjZqkBy/jZx
2xNCGQt51ImwH4S5VHY3FCP7XI6OH8dlsSWAEvTXpWqSiSOcoAovOsu5/Q+iYCsQ
klPFWOVniwreENfIgZGJg3wyTegUONFCOHvdZauDvDa32ZKlta/PR09SKgVD4LqP
k2phYmZTveo1Xy1LH6bwBVPnYCQQOMaa0Aj2RUYlCHHvx1WvgS+DQZ336QL53sFp
0SjUqOQ8j/0oWgIpx2CrmGbCpEhnqhvhv5ibyNG3x4pC5144jyLDFxfdx0BKBWe2
lxGKftMkLn7uy9lpAB51H6xoSrlECdHAb3k3u+l0sZML3xH/nCooK4zQz9P/xTbR
NgLeuArF2RfLAcPughFUJTEdLgLBeMZhQp+IGLYmQhAIsr3XyEoRieiki2iQfKjJ
AJQ0nOaE12I85cxJ9zIkjtTArhaEO6wq/j7GYSriUYNR6ep5vQAuMypnjuqyqCU4
bh/uvLRsqsoeVvpQA4aX3eO+T1VJHTHehkjZTSWz7vBqHNHHUUZTIiJ19yCfYfDW
k8CUcp9VQuH/V3qDSs6TeacJiDZtRp+aUMYb3wRiHIb9PECDUO5et5LMgvbpHQ04
iB1GT7/z2FDIqfUvYTSX2x7aBetED0qYBFmAS9u/W/2I3jbC8PwNOvASl+ca6H6O
eaEUjaB9fAf5FMm9m3ZWdSw9qv7GuM5PJ/dus57n9enSk4MVm9kf+k1Uf4Pqd3gH
zsJM74qzIaPR0IolTSvUraYhhjel2lfTXw7VPLOLRuRAAGAD0T0ngiVcm+O+k30e
yRalQw/blq5HrVao34mnl3LfkKeHJaz9DaD/bD+mvVNW8ARtUx1R/sbx+NG8NcdL
H+mxdosbJ7mqjyYEBynr4HjsBTq+ybkdSJt9ly4v+WrSGkVJslqpVvvEXEq67FZN
9ZQJXybwV2MPxREnPNzVMiC3qZaIiEO73oKE0HulCzNiZMNJ947AznFqSydM8/T3
WjQgJryb8oUU5qNRDO2BjXAwkIh5MENYmH2ijXunr1qUQEkJRVNOzcUSaRHhrXxv
B1SiIyY/NxZFzSObMgwvGjyUDUZUzwpKjk6qmFCR3AcgDsGuelKlin2uQlYkQ3dJ
pAR53Nzh81mxUdXNcDWlRWMzMB+23zjyxJi47phSAVcE5onWKqY5FD9LLrRrE94M
zI50fMKOsyXQ3i6MER1W3vZK+oVVV/nLRhbDdOUEVcm/b85eATE8ksHGpj1eRXzh
LkPav2FfjY6JcqLOYTbVO/uNefV73LnS9eP2ZDL/xb+xo7kk/Hs8jiGvaiDlLQZ1
pwKnlwTTuyidCPxOOxlr7YFzj5Cd05NAQMHVusyrC9annvdQKJoKT0eu1s+x3SHN
90uy7aEfBaVKwU2ijBSh8JA4y3oEkxbRhz7sIPkq/1jWz580KZQN4N7EO8+U/K/B
1njO4UnK+jT3iAcX7g69LLq6OS3X6eaENLbVZop7rAiAU9ouij5kT2fPw9aO6j5q
gZ0OlZQX8I3ooJdkNoVEANzhmzJe1S0EITthNZ9q9d8XVswnJv8e1Iqr/1KhMyRK
gqBUjNbFrYhT/mHSLIRBqkotNPQv8bAMc7fy6x5/mg9Q9KZhlqE8cBvkQ89t/76d
e7MOZ0lvxudnTZzHhdskWX2+UXKJ6eDDPPVk3vNefD1ZBVjcdLgMhgPRZ9EaJ1zX
4cXV7gPivt/T+NiDQBFumIASpIRTjvBn8doppPVW1gfdtbsY+zVTqK1OS9TIFdZL
1nSgRgiN5kAo7iR4agOXcA48mZR7ks1MlcJnrOmRe9GsylzDc6Qjc2qEGWCjJmOC
D6/O+QTnPnhsFEzSbqVBB70lggvvfUBPjVVg+43aOKpC02rPCzDFsrPGWDfnAtmN
Ji3I6NuE/xqIBhvgcpOVMW902YoEJzer9Clld3TUfbSCoA7ialo7pSjae18ngKnW
i0qs0TpBWEmoho6ngn9ASgClAMMnOMlqDdfnjWdIaCoHaPN6yPxgumjEiJ4sVdxn
1stqh8tsI3qBgtbcoYmHC8pQEKXUI4wNekD5qIUfjJ2ohFAn1fpTK1tTC1xZaGt6
gvjkABuh22hLcd2GnIKFw7X7KmPrLuI0CSU4Uarb4HoACwQw1M/MmZ0r48QRrog7
1BKvL27RP/tsi8S7UoNd6ZX6IkSb0PHw1OjBXZ5F8BzS+Gyrpbm2c1chPYMHb8vt
GbHhal90JctmlX7o0vqFXSTU0kdYktByidVw3pdXeG7CVYRym9cCxAJPt6heNMwJ
A64TKpfxPLTVMA0pc5kyhl8GVc6E8pdHO3ra6bTXg6/0Df1ov4qrdiGnEB7a+Eiu
fx7WevOAPuTg4UkZWmm7bdcxqbASWeWLPTtbQeUBntkhc2MGJYTBpCzuf6y7KtTa
EexkrTu8+auXQUNdfzP1qfm1d62s6kKTvt02SWNBKS9zZltUaJLAKclwUp1uZ/01
95HaT8gbOLfr0SvghMb2HVFDPCYvfpdFp2VFkfO/BSYAMxa/ZImbMqSOjvg+JbZk
ZXGBcmTBmWx+2tzNUT13pXCt3jtkyhYVa5FXGA1B883crafMi8NApfotl2RI8ZtT
Sphu89ohT0WJIsq2dBIcC6forxqyyVRFTjpfJXdVvnuY3kr0PREOESrkNMYLyg/A
DGDTUWezE5dry9bw/MQ34z3n2+Hk5ZgkkIl1IZl0jlOeBhmeMcroiQv8EZ/mdVkq
NY6Bu1JtGDnLX99RbszF/tJpJu5yWs6gphiv4P5em+oG4FOH+sFKAxACja1TYYyL
bnXlqWQJDYS4dRovVv+XhnqmihJg6KQI6qNwKuqQbRdvCp4UezBTBRVSwEDQa1PS
07tmuq0HkZ/ErnJS1PBCd0ajEMNUTz24bz3rV4gQPPSRq8H/3umIc5ziHjDsqyNz
SYZ73+Xb/6R9OucCy3X/SKwTKi2D2ZgNdKk7I4kkAaTewMAej6CHE48qm60HHgUj
K/fIUSSRYQRVyCXpFyga574BsXzrppTFC1++y2WyddPCFUCcdtGQTXE5eskI7go9
IEIeTkAgaT2+mIy93LzqTf+9BB/W7poqW7s+fLhced/d9vwFXHWkvijW1ioYFdI4
+VCbO51zk4IyXjwobOfHWLF6M290/rIZqmlaouj7reZpw+CWIIHwU0yFKznuj/0m
+/uy/Sl24HhJ8WZdN4RlZama9FhPsCEccfdr1PybLnLwmwgQShrgddCCofHeRKaR
/T5GPyEK/yeXVYduq9DFooKTKFmFHnsd3UzMdT7zdwQSJZButAKr+poXV9ilmhf5
4abDMhJ7GTIrIPVYfH1IN1TxXwYkioBgVcTpdLaCh+fC/QqLGQbulJufYSLrNucQ
EL5mxEu9SPBVHSRTRUTwFqtUmQXr4MN+D6HJzFwDO1Jvw2bdi27vFZ3mQKtsS7wq
IKA5rU9+Sh25WflppA944z2gz1/GoSIZFKZH2YqaENB6B2C00pRWPMLsio3ccWdR
mAjyvPJcNOhKJej4JabIz6E5R/dTK3kLVUbEoZ6/nyr+HuJR3GJsLEf/nQy1iVfh
omTc3pzw3hh1I/aWsShSKogxpwH/YGCptaEAjZqjZa+RrHPbvfXLR+axF76Su9kS
uVWxI/0eJ+J74jrNRVfuXwkU+mEckHYVHsnc03FKlQQ8f7fWZLGJHs0gexQQpywR
17f9oLd9yhkeOYMbow4WbaVIaBS78aGwQnULRgquhf5f+ysEK+hawjHwiKf/Azm6
iYXYrhM5EGFEwicJdpP4ulITbD47t0Q5PBlokQP+jGZXsSSKfGL1Jykh3BsP9QIC
gW8IggL32zZB+3pGPSdmhP4gNWfI30+/lXwYZo9jlOG+KTSvUK8ptdq0BTA7GQrb
9idI75FmHlIjPaxorMGdq85Ja4tLN8ktnP+jKjQXJGSHBltLzuJy3YlzfLhKAKnd
txobR31bquQ/LK6QserXwZHXInhr1jK72KdhoLD1ckP0dEdmCgjXIktHz9mE3bXi
JLFdxa1dLK380XqCM4I6mPtd8yPMKsqab9EC0ywlAd6mJhiUx2wJsxWSN9GBc0c8
JU11YThNs0Uz8tUZwFOfmT2jLxIEjRQm8nSDlGjH4q3moQwCJcyy5Vy2mXJQvLTE
Jt7eXyNnwbPcuncQpbA5koawjReUTPxmWQ/7d7dUL0nIJ/FbJAQcaoc1pMc0niuD
M1bi0XUtVe04oUzCYk/y5vn6/R2DWNU7xgVrQhXdp3ga5FIGbgcpQJRY6feMOpDS
SE5OWrqCuv6n4mFPeAB+GDKZ9+nouDfzLfTY00eS6S5fco8yCN5T8AKTQAAWMfU2
e7QVcyFCJzMyqI6b4N7G7ByHzJqrp7jkxIAwim+wfNiI7aMKOiTPQNmu2vkKygV5
tf2f+uSWWVyHYgcvT9yDbHsn4g7M0roUx9qJxARTEhcYATUBaMnOpaPOv2/ITV6t
ss9X98HbNQuak7vHxY/oTGTVgoZB5nSJO+f3kyf6WnE6VWIFel2Wa3W3kgGl+6u8
c4KXrBxA7c2hnkcjRjgh93lhfDVKiKiwNZFgWcHuUfqJHrLFQXxSel6qIq9YmQ/g
e32Y+vnPvUx29IisXxPseUVoE4rgRk3zwzvaVMh/x1YZ3KfVl+yCX2lrbXO31t0O
AT6vDNjXDWXMOG1n1U8vwbMCseXTVri11V/TbJ7DJFRwJ0zmnILeb8pkSf5GMLT5
z8iDB1QykpP9nuB7zWHMwNULWQeHc7QgZPtBV6c1eLxsJ+11/36VuqUYKqRfF5O8
yvgVFIMU/IHooRS+qDiXdCcnAeiZduJIAxu2g6PmEvLPcASpwOIMCmQSFo/0UXm/
Lt9y2TTLreP6yH1XdEWKuMUnFx+qexRXPwtyaUAVOKNJxHtZl2OWI+NkfBCU8yUJ
pbmbOQP7Dk8NfiPJAQD8gV4cDu1NLh4FaZA4giRZZ59SMxMUSXne5P19geEFsj3b
VxNRGlnrigBaK6bmj0vB1BqZBBU8OHTih8VkxP/0W44K3NOGaUzM3MusfO1bQYDJ
ZHiphNzjLWD3VbUM+SI0RDg94grt21qkgfKhdBTIjRjV6yf4uY/Se1ujby6keuib
gM+y9/yNbiFUBLgnUrrnVYVZev21Fsm1HWMe0etyP5A/G5UoHLq/PYtqUV2qS3gb
5EzTwbZEqVWRAfnpJMCER9/yXsthTX5AgG06rXmINpp2qExX0tQMA5ss9j0OFF2V
hAIhf5UjKBVcnhBIwbSbsmUtgXaeyO0f8R/U+SCXczCVISUvzVolisHUbSYbZBTL
cjtrPfgwumybMmt7uEt4hcq5H49JRsGcfPFYhjwPhj8btAx8lyBqN/4CVpnWVH5d
gsDF4zOyeig7Ac3AxxSmDeBqaqd6oEe+aPCd6z+BxGj2KD4pJkZietJraXjbIzzJ
IUlTNafFMQ/PETWMf1dp8el/G2bL0lz9WBBex4B/f7AkmL6TajaNKtRDqNByzSZ+
yYA7LoMiJa+lLiJDgfwSXmKSaJgn8DRMhHHHZ7+6nkUpNdKCUoO9769maJHvYbnl
X+juYXdB6XApILe5sMsKhm0dVMfRsTuoNos576gvdQfNtFBcTQop28g0oC0zzzJ8
5MpnvvLYafpNAxpbc1jBptzaRjMYGeZZC0dl6XW7PhrohNVj3VCr2VIvJmtc4y3X
l7xQxvBNk52BTVM6xWcD8iDW152Z3y6ebEFSkljAjTHAvbYifW9tAoPnvXIEU0ef
WUnnTJd6zYocj/KmwXuo3m1vEf9KtMsyXoTXkZprXzQFwDOpYifhW8KdXDKKk7MM
Vb7L1XzvtXh11SmTP1YuFkH0D/I3iMGJPPgYukQXmKEz0Hr1DUfpJg/rQ0KX80kL
SJx9ZITZ7UDYUAr/WpfjgiEsg+9bFKtcAS9cvwqYqqd4L/QvAad6pxZ2sftyFHCR
l1sOg/vDLInMF7K7jMANY2qO7aO0n03/gBqPJwkfzF0IdEgcaP5kZeaqMd+/tJH9
wYOU+TVP69duKfHyQ3T6PmL/7ulrdl+waeZ9DdqjwfL0zMZTQeYQsyo8X9gLlgjp
2OAtjcZQ2UqDJA6ms/10C2guhJlE1qmFRNaImtCYc1mo9DZ6x22Qyt1sZeOPGmnZ
8yICVKKBrEQ7HL0FzXLMmBefqQ6BSrKDBCzskPHG035iBuiHfMBS1/hbVn56zOoy
b58Y3LA0KPJet7JPXMN4ZiVBa9dV9wXrSY2LoHEY6cPmi30KpSwKwsS/8/ABk2Eh
nUNzxUDtNvvBM9SlU+N5EEQ7DisIRAGkmNFvCczA0XXlbblNRLBuM+PvCgl7X7yG
ypzcyMgmzikHt9XtpxCSlTYhYc2p9TKiHjEcJLOAI0MVgIeXkUp90fZJBU3WgQJ0
K/atY7fVCD/MqFtKK3H0IjT4B0TOIA4eI7H9Eq7hu4mJcG3v1irPTVIOaISwe7qd
3ahPjZ587O/jd8//UHsdOa7Y+ipHCKM/Di2z9th7/71/9tzLX+fbc4UVijv45POb
KtkXHqtrDx9sPEITzzmulgiP1JuF8ojQuQRbSdQNd7dIa3ymAeYVl80qkCy9at1D
R+mM+0yieYmk2Su8w8+K3oXz3S931mr8TWrhf0l91h3O6AKp+3Dnv+0l4Un5m1na
Uej0RK+mP3bw/H/iew8s0c3uUqzqZgvSoCv7nRa3I2vjppHMX1wSBiLAO3gwAKFc
D6wSIbPu7KNOyZDIJXYJ65SDVVVjblYt/Sa/4CtH6oQzY1DFcueJZmiBUppSNean
zxEzgVVlwSi6oL1DREWbar6kaSqx1AOQiejAIQaKupPd2s7qMpnIwNT8qF/Ddyoc
7YK3CP9/Uy0sTYqFA9tPPgpdCpJlT7Ho8HmrbUNoJQpus257SLEPs59DY3ojFSh+
itLF+8+/KKdveEhQpHdHRki1UCYW2BYoQirqxA/oRMOUzLE10xQLaM942DcPw+GV
hUHKwOEq9LdS0NmFU9JN+9V+wDtIt7Z8FBGH+ZtZ+iIj5Bctvk/Jc8lm1qzXp1ZI
64rnbDBmNGKJC7PUcfoAEx3MLco7SmCkiBJCSCBoAy5BcSc+u6AJlCCPV/Zsi9Xd
s+n+pBZNP6CcfNY08jIGBLJVpWjHyD2svBo+pN5WHi9jYgxnOpTC0hTc0a5F6vBz
EIJaQro2ognScrP2gcuym3uyFpzwWhhdW4UVmSCk1gk1RegFbJaMkeKEXZJhOHNb
HXzGfFE6BX2jZrDM1BgK8vaCvOHfk5C77DGv+CkkMXFgP5YOEVJCIRFTRDoDjCoe
SfXSrK68DzgpooohmISpUg==
`protect END_PROTECTED
