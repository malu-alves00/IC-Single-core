`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nT8KAZjde7l2JK9EtDstDRrFmHjt7y0E5NpGvRCBcYTsusiIH2Rw87FaHDQeKyn1
SkWefcObzQPDQu99q6XWDzDkm8AXZC3MDe1eY2REyY79yyBdIG4zcQnklsIXhe7X
c8ttxbJ3aE9wbH+an/i/DeuW6fCIJNS3A9b5nM3bZNUD3rFDpyExFDpruKnwut7e
eO2+Dyd+awziJ4SYLnrWmZofb87fVsY0CiLbdMBqC1YXRvQBvZNPy0J0Frob65kA
33DC25Vrms4nagLhJWl0Jrxvt1XvW3rlW3f46yo7C8y7av4T7uHc3SKVvJOuHw5S
vj2hTDpghKkvdoiE2oSD39p2l/ujt4myz9s0FwpDh7azb72St8FmqP1uYhS97VAW
XXwJfzUe9Zf4uddXfbr1f+v4qPQ3lvk6aqz9vj48xB6G092Eq/sK/M+8PhRV+Rcv
SGCQsU5tgGVa0GEZfYIOPtjO/a9bvvBi4lfcrU3z5ODibtngSU85JG7UTqqiRw5c
arg5fFlCpEZJPnIpvHddMd7Qem1cm8erPfCS1Jr2DfR7y8ZtCeKoP/7c9c3lOER4
lqi8iraMsPruOUfDhxukKp4YBQeqBQ5GGBXwHQ+hkxm4Tuub64hBsS50SbwR8E2+
RV1St2MqZu/QE4xqxyigAYh22OkFlIz8GPTzgxHgdL3Ifyq2YqIB/pR3wsZ1pgXY
tdX1zsTbNwXvAQVt19EURtIbFZlPayXO/50QekeE6X01XuenhFDgwFr0+i5B9mbX
fROcAqFw2vnasVpD6mWB9llOTQW+LUgcbD8nmZWzbTOPt/qEVlM6hRElMckijZP8
arvrKkOq0v9V0Y1iZ15YxED2AVAu52Fu7j13zbXVC2NKPdLgGblkdaUqk4lTNeb0
FRwd3h7BD3EDOcTKuX5iJElZzUBofS+SxJ5zBuOzIdMtJlms7CkAb1WKJ6bRXCo4
qV/iOb1dGlIjjJaPF6fp52F3rkRVTnM20iifA84objZGpCwjPQw6tCQp1KxxELFq
UmlOJPtisobUM3fC9Qk50MgiZJeD63kEqQJYCLlKauGjjIjcz4YMtBqbpwUu2rYW
HjoILiLHVt7NiStTGpcJoaUxmHwofcbCqo9kUUo/gTEzSKcdfX0ULh/akHS/raFg
zSGKjDzGKpEETD9CV/aBDcJebeeoxiRejnRUIWN4+SZH06km4EuqYfiIY/p3M1xb
dHMokAip5w4nzTdNI6/aq0osGPqM9EsYcQpL6/2gsStPxgb+9aiRDujJDZT2MDWq
M37n9ySfTzBXIzIslvmPyAmp+zWlYZ7faB2mryFHjTt4j6x3kzOKG2f9aiKnp6gB
LoJWdBo2q2Uw/NoljRtNTMNZ9Nu1pn9byy+f0vYjsQXEg+CHRscvg5xo9nRXRRJw
mOgYEEu9D51h63fmsyDkzr+k+OCaYmAwkoW4NqViOvW+N7uYK8ublflocn5PdEfM
3P789gzgOwJY/Ft32gkm3ZZz3zT9pQ+LYLfg++bHS/L58SbMqc9dI6AobpwAaGOf
zPzMKCqgflehVq/IhJlw8oQBWd8rhw0mqIVmWjepWyEWolXhk90h6vSkHSYibaU1
dG+yxa5+NsTWJOfYmZhC5Ei82LArXi4JLmTeZeKMMyxhKROgUcnvJ3Ez40yoPppS
HhfzCJhgpwa6530CnNe/phRRb0YMhN2sR6TzvgGGCoNOtAszovrpnIpq9ZkLiQ5i
MzobPdjIa3i00FYiti/V39kGSgElwiJV/NCWVNXivF6Z2YdtlET7cz/1YbgjIWKq
fmkY/J8ubqZzz9y2OdJ/QinsGEDiJYlYxL7vP9xmzrdLAgs2kPLa1UjQIrZRBRDE
apQedEn7UxPd22rGHQBTc3oMDv2z8cqrA85BhxqT7CQB0NdeVqQbcP9813T+jSJW
Lmg6zbO+MYs+G/zYLepg2upEDR9Wdh8Vg/D5KBP8e1osC4w25nDuKbMudoPa01Yg
CJeEy1zSQoDPHtqwjparu3IUQxdULy6T6X+zWbDXXFQFaI1vS9SjcDoWP5EVs/hE
SU9AHMDt7yaKIQV9QVEIGRPnvi9wU9+2D0RTjYI4oE92KUEtOf2k+6Fiq2VTzPBE
1Bynom1i//qytQAFEccNFrtM4WiaEQfTf9ADd50ujZ4oa3VKxU6V+KTIKq1Mos/o
xXzyxegENP0a5TVT3GvnSWgHpWXUOmBaWTd+6qc2BeL8NKsEkK2l3BVGbkPcl+WL
AkZKhMiSx5A6mORgQ7sREGlPUschFG8hAqKy9llxDuvRUIZlMRK05iVB+jarQU/E
cYPrauDLp89eBbmeM3zfj5zEX4KudvAwbwg2209NessyHDVEREZExSVglcPpD9El
Kxp3pkSUV05p18x6NIZgdcoylK7au22QqIcFjK9xGdy3IveYfoH6mDvpdSElw2cK
zPqc3wLkLjogjKM50G+7eRKuA4v0z25ooQEk+C/ssESRdSHqs1rKzulalIICDxeq
oqg1zTQ5ghb+9/nW4XtXGQQSrrjpVvOefWorgqLQZpvMN0CFnvW3sHcZ3XTGXcMT
zG2Gxwt8R+MZBuq3/1CyL4B8IxQTCX95KVU5SKFQJDNGX3mNU5ycQoSs6vcy/RzH
pgcJV0iu2GVj4KogrDR1Yu66YI+iWjiB0zfrBpX31UVT4nqAetuqdhRkWNnUlfyf
0PYcPsxiy9UcyA5g4IjeWHENHj+nkvbR00U0DxiOHnNlMdb9W0mQSACsUOkDKFZn
ZOzFSmI/6CnRaWIs9ryayK6o/BycIzOjQP30i2aDESBpqOGJdzLYPr7WYuiP99yD
Y28CGA3vdZoiBtATt0gFOBoKIZ9ojr5bitDBnj7nssIWjy9+P+EHHyeX88LnIgDO
9OoMPRv8CFf1/UI2Jz1O2FmhE8V2uzx1TFEFHflwYvhgTAEyPunLHXlpSxZjxSsn
XagGsCLfnD6LuiFA/lGCEBWBBaw1G3yuCjUL8lQAMSiGNwnQDDdPwjEG/dlZrhoH
yrRqgfEK7UTBFxChDqgeO+LxOZfQmhJJ46tgfWANHHqSuBkoSg1cW4Tzl2WIRltv
ViPi4spH4R+Tl85ZILehH/JYL7bctazWe9Ad73fkaNWwV7Chse+/Sh6x3ZX40GUl
ZhshO2uvOrlHH6uc+x11qNXbfM9FXBgDv6PQnaVnWhNXz9ijsswV6kds83JVfAkY
PDxqFOnQZ4wGvyClTVyBJ9ed29jaGUcNnjU27ZXmdqj9gedw1hT9o52rp9YoTvrn
GGV66Iz+e6NRzjNch3XWx2tPicVZg9TKsf4UMNtiJI3GzF+Ue7lR9qj/xmM49OQ+
IqLBX/Ih4tzUBMntgCPs/5um3TzhGqU4t9FDIjEFkJmrMOi0ReMRXaUtv7tb4J2B
6LcGT4IKJo5nudQiob3ymGusthMI+WX3eBqOld2uCguS5FY725sKW45vi7Givw7G
Ru0+awSL/+7onI6yvARBhvpZKQwduiQ+n2K9/LXzHU24JcJ26f9QSDcvy6muGQvH
PMfYBrzKV9UqVyCECS4XKeAdEwUaANWNlnloCZWLuFSooxu7w1FawqL+paDwEoNM
3QxsOWFe5zDKM4gDDu/AGh6YuOTZ8oopzVd4sWVjlLSOGv1707EXRzQUPNNPg9wJ
uMXcp+9BGKu6gsr5o1E6u649tWSfWNju3+zqYDvZrXSpAfYd2celyxXetoMebfqL
e2DLf0XSGyi1O0UiUP2ZcrMSM2YW8DoPWJ9NeOVfzbd9IJSFHe/DSTN1xrntBXpY
hBCoXyhn0beOhfmkNgksKw8L5E2bweACi/9ehT8MAmOXhmJc8nvL4s/60mMjtRtS
cHU9KJ9yYznYWlcWbIdKU7I0QUqJy930BIex+nWwzAiT3vYEYJxaK/sOGjnOyLa2
AHO1k86a+tyi2XVKg7XXOoEYAMf3OeTg03jEEfMr4udzij4gRlNqkkb4pz7vYI2g
MwYRqexrMCZP51aYPgJgRmlesWRTTXK0wgfP7rRoIRQ7DYRG/iHetrQ5ull23m1i
6AVefBCl+qCE4JcwO6GBKF4XKcvgv6MpU/3TlGrnzG6WwDNlm97ZYt9t4IAkosxt
wcy3pqDzeXBmdTnSDbTaaX9VwJt+qb3gIpAA0WE2ZHIZpLkh8msxDN+3bUvN294B
gOJ+Vh0qgSwtpUAWviiQPmglqWHsKC+MoTBsgm2OPI2eU17U+e8l3h0alsnyMT4c
rI6XF6xoyKmTwnJg6qFbIj1ocyntz09G59iojNFIGky8R1eSRHFmZLYAZibeTARL
IpPa3/+cGTL+qQsAtsJ010Z4B9qlcfLfAtZTNAOJfPH3XVBUmVDTBelkUE4L1B6Y
r+ptS6Uz+1FMjHchdZDt2neNNqb+OMkmhAWEFkmcQOSJxkbibiygUsmA/XxYcDke
9cLVnMIgWXVvLBSsOVryQZHBMaYKe0roThIFjQFp29DwAW715PFwUXKmQdxsSncX
JFQM0I5MT9uVHqJIf8XRDLiKPc5W6IW468oWbf0Bx3cKoPSPCw0VFUy1yeXkZHm0
KZnJrPNMk3UTv+bjsESsB5fb7fkpJX5/C8XRs1tTvXrtdD+TDduf0c61qFxu9Yyz
pW2RGMLR8hhQHJSKU2az6czzY96hRLS0uvXRQxKySlSdMzM50QCVArsYcUVRMZbm
irOizYj6acPmJA/Pa4uN62JtHUt1t92B9fKX0U0+GlsT1R9bkA4K18EblpHu7oyh
rxeUEIGgAlHERNGGTE72mlJ65j8xOpMytwPovDAn0MXfmSWWG0grGFkVacsHAM/R
GfLUfqkzXc8eRdksHeo0czCDjQAFcERNuRtHzTGogDXs98pAL1sjSjChRN63fASG
GmUETlejfOQh0Wu/QiopEWD2L3/ViOPDOG/vxREcbq+ZvEzGBSXVLIkVsgz4lw+r
YDNczZbuyz7BJ5xxsJfr8uzMe5pISfTS6JTToJbBFdXzW5fkaleLGgWJ8d28ROTT
/xPSlyIJC1EoY9e5RSOwJw+xg2S9OnT9hYNiCiAyWjEtTs/mZ6jVVpNx6chIUsWR
y0PlTuJ4ufl57pkMa8KbfXx3tjqbcdX1BpoTPNcxCo/+hXdrgdS6vXs1my8Rs3t0
UYqMYSewbI6hvDfgzan1t6G8OIGQDhYn0tpsa9EwIhc8x4v62ZbbFbp2JRXQuaOr
RHE+DxdI+CJzy+uRYmHXK7Prs1z8NPY6TH42jE9HUMb0UZ/0xvX3CJHRmt4cfj5T
nEiiBzccp2GHLTQvJ9rzqMwL/3/ptbkOQJgZG+0ft/G+PT6b8bETUfYIODfzvChX
NBtZMbqlP0nN5fVtjDxF7Csi9lBBU/er+L0FUMb6/+ciLpZJCYGpewhRxeoGuW1K
qczFHSXxn6IfYer+AsWEf8nOZsvYa70+oeS5S+IYGXxogxvIYSpvKpg8L7xmhCVd
eDC2BxdUwNoxmgFW2NIX/ESjADuOHwy33+kFuP/1eOO/VgUkXUvoIslP9v+UYtzK
CmFIEO9sR6ejT7QQhk7x3e9EY+UzoHflE9DizpdZ5X6It5D1nh6S+yP80BGGIQe/
eT/IABqAP1UK11qyAdpkahyXb28SbVBZNs5Pv3IhuL0qE/fqSoVEo7to7vT3Cui6
2m9ZaGDAc1fQpGeNps1UBSlNDG7cHVAyGT6qyP8pMJgJ+4IsEvQkcgX1juNQzNGl
xZN8QO9J73d2qgGyfuryChm1OGBtyGvpmwWupztPRFNY+TXGsNYCY2BZ1SfGvNhu
Mjfuj3HxASkB9nJlRpKy7yDQ7vimEyEHtt9Qv5CY4ESDhvn85wv4YvsK1/znxjHL
L9CbrWM3w6duWnHqyM4sRIDYW49YZ0sqDMlqKvR0qLRPfigynXt7FR8e6Q/0/lCA
meE07M6uoVTbOkU+jRWsc8bkJPLYbg8sVmIcQdbu/OrGcBG6PA7X+eK6WFQP1t5g
kxG8wJv2YfU9oMGfiDflTJsuW2qW0Y8SPJko0oXdsW3HDEl1mi04J541V0Rb+Dhi
dcoOnNPGNK+i5RuYD7Y+t1gGP1w8wkcjK4git9Ta4cPHHzHGPeY8QixS+45Q8n7s
+yPm/FWyEGXp8WAXCmg1KDD5TbPigrXD0t6vlqI4+C0MhbPXeGsh6+llrPuDL/lC
TGxS0DRoIt9I3oFf9j7s+H/9hAV+8uTokxh1eQKQ1iXEHHlig7oPAzTtRDUPLUBK
5G/MXC5crCPP292eBd7+h+pzV6Xd4gvdpIVC9KOH3sVEVjqVGos2fGDjY5WYcScJ
sreJhQsrWYxakpcHf2/q4RE6SCBwnLcDTOP/od7Apjx4bNNQyzmIfcs7a3CWoCPr
aSu8AzRH/wL9c+407A0zSBsYZ67rtYL/5aMSH84CxRuKQGsFeP+FNlRw7nGXboKF
KGtbFHey3OorRseBz8FCCraLYEJdycOWgnjbDXEPjh03c1HHwIl/Fd7qKZtwRzKV
ErMcud8A+ZR/mzgyCHHgYMYN8acSEcDZaBUcJYpcvoMvQpHLEVaLX53uwLYkj83/
FCY/mvNI4Tw6rmZ72gjEYZYrmJnXeHJSqetb0afbHgmdns/StuYNLTXzlOnCWeOn
F52epOQ4pk0AHfB+Z5O8SiIcCOwGbAD2Xd/GjI/Mna2g5Q2GflcyVw+jqWtNJWSQ
tDnY+x0AO+G0yKWUAx1HvKgAnvtKj9lSlobAYhxmKup5rWVccMbWGELFUuBo/vQx
hKOx8ijYHqPloidcARqhFAlcnEzunh7/KL4u1sydkYhQSc9C8seW64W+v6yVDCti
bqAe1zW/p0/fNWiH3ewsxCmIMEt/Rcfmo0W9lcEc0gJtlpkLHX0BpZ3CLUk5fU4l
YzdZh5/3c06iimBzvNRibs5dXhVSxvd9xo8pht8XcP3NuABBc4pAd83Z3btTjF6O
CU0fOUWcuj1Wyp4m+RAfzHrRTKAmkwOoLmeFxG5R7opuyAVlotZyfVFAQ9LxEO8W
zlb1lzeQm7prhL21DjXDtE0NFCz9lFR5MfPzpv7VnU/K6Edl1N3fk7YQSgh3yoKj
KC7RXRTGLALrLwwcuCNyQ5ET+dPpSLXnXPzgRRGrXIZBtHz0GFSfj4+J/0I+UU2Y
WC6nZodBQ2uXAfmc1kg1e3tPpFiNL8P0xFuGAdupZ8vKFtjYHFAqd4SYRsgNCbIa
j/v79UL/VJpOtFaCg0YD185UoiGvbm/jjKwMTabnkHzHNW0Cv41K/8hDrgD2SLVo
TbTpQygN/uN8yUXWSvneTGlaAvve6JeZ7AFV2nj1XcXkymyrb4Rxr8E4yugv6bQe
py/UXtWqY4eMNZF5Mna7hI5Hf26+xE6WPYvx6yA5vkHAKES4qSiJBITCiOid3Ajb
UDfzj7f9BPQeYBMmkSkUzs/DnhxKYBjwWbvoc/i/EV+ByDKaXhXSlgQ0GUsJlRbn
c6AbzwrlE7szwPhCwfkjFpYRuZXsVPLvBgy9CiwPlh0lyL+o2Mo70yDJ6IMb8vUw
TcpjVaZDSP8ZQS6Wr95epIqZOuCiJ8yOIAknnWd1gsBNe+Q/BgigRUkEf055veJL
zYiJKNrKiZnfMOTWeRnOo1lJu9bJmtQhTsGXROX9cX9fWyZoakZjsJ/zlKCaum7b
ZtzfuNt0gwQh+S/VKUpSHtzfsYjYsjxlrxb14BmRfNZJwCPzoPNT7yBqVBiZDE/q
M0KPtWrzIWPgNAu2UoOFO2IcqhlIndJqitDPFy0TpwoWbajBQPOfKm24VFzCRQ0a
J9iMLlXHJCMD3FtekupJmax21aF3equXaRFbKiD54gC91g2uysMnuoWqAC1n90j8
e7TKSHy9QxDE/DufdxlasorgsAWj2AHmeYcvKZBcRrtlh5ns8MnVZe/kkWBuSezH
YCbiQoH9swHhRZs//ZSiHbj2gg+CPOGu80WrdkNKX0s7bvKUPTFsyqVva+GbzFbl
+ka9qPw0O08iorzD0txDzGdI08Iz4HT7TyXxgXpIkJSbxjuf8NG07oImzZG78AAj
Ei2y7RyTbB6r1F+eKqBULjazrIc7NGkKo+FPzq3DIfFtcT0JObe+JaaeBJONMOPS
mnxxbivfFYgRXbs03qYFuwEqwbRfxntl3Xs3hBSCAYrVE1krqlUH3g+acWfgGuNL
Sm0F0c8B5rR5W4YTMcOg1O3/Q3LEQc6eniDABKk/tcIbW9jVP8yUK+yQE1ukcN0c
X9qOsEQbp+ZfPpLW7UagSj24Ml/LhGN+qgqTrUp8b7B2oLprhyFnfeT+y5sYR4TI
cSrViIDnkIVklh+S+1dk4vFgS/6lv6Q+ekIsRUYs6NwHKb0uav/475sIr8pnlT3Q
2KWRWHHgc2F0pGB3ErYl63pVPqjlvJJc3+5vUkIA9/DtUk2FMEjDFGND690T8bgK
c9UGuCeHcL6mRlKwigXmzk995t98DWifUjM6KTy6xDEVf+Utpem0avzZJ9p9QTuK
FJmte9GEN3AxU/zxMRl4NH+rdEeZuQLmN1WhNaO1GO0X2VpKsOTJ4B36YUWsRYY5
IJi2hb2CDT7bIsduRmxgINTTc0A4mpNT+O7YZITqmVZrj8WuGy/uhEtJQ+/DYyGd
a2NTNonU3XxEX763VJrlctPc+D0oTjnSBvc/I8SiBqTqOqceJ8gA25TXXwYsAspT
JTU+WhwHWILNaDPxsmUKYsJQYUsaz6XSOQL5rGP5ZlcHKmCxbG3k4HvNfkiGTBzh
rNt5Sv8zup/C6QQumtqY3SMRFqYFrqD7zDCj4AA4VreVdwUjlkwRH9+U/3xUIDP5
GxbekPwMm4KnAb6oF7fAEW4xrkA01lKDVVbJOncZ38Tqt8yp51HaS/Md8dqhcfkl
LWMA0q3AgsnIwylRJLnkEWbqK5n46UGdy9e71R4t6XSNG6fNt/x4flsFW44QJWzW
K399G+Dc4LyyHQ5Y8ummAcmy+XaNz+WpfeSJbvjIG8yTzmJiYw4kMa4ge1K01n1w
GS59tEskcEdIj/FyLofwD+U3qzGAjrCl/xehpL2LlLaGTXvhqlhTyKfFgp4hq2I4
FquJLuo3nsKPItzDWwkWKT8gIsxraUzUE95yws1sKZC7ee/JPYJpgw7uFbmLxjUs
bzii0eyKuYMGkSKMgJRYxjlEye/TcqybXcr5OQOrDm29B4iUZrJsk8O9mm96C+J+
jI99jWt8YHaggh8cYwEB/QebeBed5Ooe8q3mOp0L/N7FZU/TSCEGWOvC1slJ/NUm
cRK/Bpx3kDDcdjg1FXKF2Br8+F7Oh0F5j9QmDORxDAdNghUr8UlWIPsvp1Ts2SQt
/fQksIiBqUt8VRl6PjtHlmV1Qr6p57qRaBDPkhyR7YtbWC5zLQdFoM9e0Azs6XLt
UrzniCK4aGtX9/5qkajOl+EABCe29Ce1MyOLWVr3rVy0vTcZvXlZyx3StC7hS6D8
+EoHWK7XafNGKDCc1puT5sxwn9lvfVbuuHI4hMrFxbSkej60UsT5EaPrpSy3HpcQ
XGBpIm1t8U1czovuy+yRvcSV36IsonrC2JgMrwz0msBPzozP7s08/a8ppR9t9FTn
PNVvJaUrbhQOzB7OkoiE87phNl3QIMxthhInyPy0D/foQEhnMp2QYLdqKeo4P2lq
PdbH44QxohyuQcBKj/HX6Tq6u/WFW/2bChk314bkmvI7Qs9/umtm6W7fdzN/eONO
Fi0dqoAwN7f7gbGYjGS/usO0oRFfil/0wzih1gIfEfWWdgorQm/YRwQ0j+vgvHeI
pUwT2t1fjQse7ZQMjFrg+9ZPFYRFjqQuLRqNGlV80siPBJ9XEOXnHtuU3dhadgBT
RJYy2bHDx0F2/RmKhC7GQaiJEedGgLbF9EiQAsjIpsLbY7Ene8YPtXyBvCdpt7Uv
ExaMsD+JAKH1WeqKtiYglzGOgTHiLqzdxbmKqo3fFoVlugpepuZhyFUW8D3oyXlk
B357r2nOIdn8+SiHFKhDn37M9TSyPKkx88YlpwKh1XY/oum3+51UG7z9y3Iu5xpC
h8hxiMaAbjLqvYo2OcO5wudIgcNs93V5hhAgGiZ6+yz3GFVoqYTss7+V0V3JGArP
cqcj2at0veXC6eoxwOZTelAlY3G00wx5XUmJGOZqE4xo3S8t/0SyXK190YwxNqGd
V6N41LgT7VxbcPeV9YH1EZZ6meJu3Xuzc/jeNsxS6hhOiMDLr/LVskdfYEp/W8YX
PQYPVdSVDzCvHAbh6OWGtuI6ZRXxEV+Jqj02Bt+txGaHtpnUxBpvdqdYVogyx7yu
549EgIIJFnvVsXMt1stWOiushfTkqbGMAWvRQM7VCCu2ZQyXP49l2oD1cCQc83Ja
pY+2vTNfrc4FwScYg1/9T/KN8XgoIbfwNE8Q2YilxN3tTP/SlYzHjJlL9p69o42o
bj+ESKpCZQpGG1v3V7i86td919syFmUl229A7Hnk8G4uppgXcKQMOfJtc9kEXRAJ
Ps8O+VNb0wkEenJ9fFhfWtrrrZuVe6EL9FxW+8NRX9wXbWFDg21hfqvVWargBkw+
gI0df1zVyzMQt60oW7Cz2eO1DDHUDDic//vwibbl5yj1U185lfF4SAHlbbBG3dha
ZGlmRb+9ZX3OgbTwzPErWmBAy7B7KyPeIbFk6P58RY3ejJ4ey/PWzBP95JffcqDd
QsuDIYb1tHG4Q/BEAcRyJRGYFO0sQ60rqV0Q6ADG562S4uHa5u3G//bd93ZCsZJx
lcQfKC7ixDsKF6Ty75A37MK7laXYtrIt2pS+Eocn6DonnM/V5LKvEOjWTS+8/7hJ
8pJ8HG2S6rf8LqJT5OnWvyDVCvw5KxGb6XQewIH43RGirdvmFws9KX5RUcn/OoG/
m5b0iF0cGR9LndhLmuGNITVysrxNHmyCzEzfFyzAe0b0FDmiwlUyfr9XT0BrjxSS
CVLnrLd0m6VaS0rQei0tXo0/3sjms9699PxwpDTtEK8nWtJk/J5WJelkYxhEqHdt
+dIfgQQWqnTVCjU7Dp0+sfI7QxRlNQLe7lKRP821k4DZ593LWCnj/mDQLcbSF6Eo
WzkHLi6bo3JSuDZw7AP26Tl9ZmpxShU3KXiXlTWuT9vuTR8zdaq8GE7Xl0kUIj9E
a3VmDT/Z2D74oU7EUrPKHY/upsTrbK7vTU6l9Ukj9qWLQfgBAjN3zzUL7wQ/Apob
ElSLLwy1PWX4fWTUAVj3h12LRF1J3z6Qi7gBXbRkLqPxKqqvtFfnCuiLyAc4lqs7
0EbBsBsTBlPRTmENw2OkEQ+7orjGt5u1uaOw+h8lSHG3TQJAEwonmTwea7bZjwI0
YLvnfvcn0D+SBO7pXKNMr6ikkItLQv09NskVv2LI0ItuKJFikceTcTj7efJgH3wx
S5yTu9+Raq1P5XvfbtLuBLeeLl3nqojEhxEHuBtFWReF/vignKV13GUb3uvnr+gc
xV5I/m5sS1NV68Jyq2GdhE5Fh02tPjRZttTt0c/t0DKXXFfv8EdF0pI1nBgt75PU
jTmSwGo1HfZP1SSdKcZFm6ZHlzQfaKZcD2A6cwpAiKN31GYloiomQ/BLbxVhjJm8
JUgEjX3do8j3vavnpoGsceHH7Q4v1lXygDn2OvtyYdJOCIaQ3Lpn+2WAgY8nOph7
L0fUkC1OJvOWoX03Fx7w2wpzozTkdEhciIEgQRD8FknP0eHYRAicZh0sPcGzU0wt
AUGsUx+YVKNt0YBcYJR/lbOM2tQynmSs2RgIs6OHX8ALsAQ5cEPQDo6dNgB49oa6
vta0dO3UIP3agw0jggFvALo2uLLq+42i3JXBIj1+PPrRzPODG7eRzH2WYtGmRsYo
QYJ0oX6v5nbwMZ8GqQgqyXvFCIvn9wvQKxTLu2aZmU9QbzuYsrerC4k60bO/4Wgd
6p/ANmpFq73pVNPslQK8d5MZKXTCVPdyp8+6TGfbPlYrO4GNHNTnfkK03qToApm9
w4w/MJ3gLMYO+gFtnxCnmMOmA6MO4q6PvremvGwlFk+Mnq+ghaRjeDlH7hgC6cy3
P+ykq6cH04XgcBUq6DKTe3tEGcS9TQIM5zBstf6fznCHQ3y06Qovp3WXWqtB4xwl
Nja9D90IBYkpXP/3AdqR9IOiMJ3AAlTuoZkto2hP8CYz9pjWk8GiEp2SIjeS88Vd
u54ThUK3U9SSlkSyQjvHWdsxjVX6QQgTi1ECcZCw7G23r95M80PjoSjrjbLr3WUT
ZtroZQGgp+AkeVrXGtdfH0VGz0Ph3IOBN+VTY4jzDK3XV4LbGM37CFj/MS7ymiRL
Wsg99YoTgQSSONA5UVYn4ZO6vp2jqpAFdF2gGQh2uQMxtAfr4lsMs7Letzgg/noJ
tBY6Qgk6HAi6rjivQstGUKiepMmbRiSC7abSLuQ2MjQaGRzRHv91I31dijt8hKCW
wHTdd/UPloS0W+KGlxtaqOvfKAgiFc8BW0zlx54EmKe8n1UAS4n6+bmdz3Xv2FBc
o4/6jX8xpEppHb4IHBcr+Jd3neIX7yns1LWOkrT5v5YEz98vojHxjIX8Sem4nMBn
ZQf7lGwF1AYBPUeotrEsWYa1G63p9QXp+tBu5JZBEcgAnXLtdt1HmORTIx03XMFo
DLQrhiJAu2BGm01dGDAHMLjhJp0iSAIQ90C2YPoyd2Qs+DuYzJW6dldrrt5tLxE2
Oo/ebzXTBSxlh/i2qNwyEAEiti++KG11mbKXumk/1vlTCKxoLWZNcd/JR8qVaver
bsL6KDF1gBjPkbsg5tKadWCO3zhWTN5JORhEjB68UrywYuV9Fjl9GQMRrhWc07n7
S1NmBxXj+0gS/LPSaLVczoLzL5teFO7VcjVvbczmi5V6ougpjQeSrSIutCLMjCVC
UzzqtW681C5fZ05Q6yC4oTmK43VZ5SqFhpg0+POUfWJO0ZlapIebSvGPpLUVOPon
doGR5k4lqGswa7A+nHKgvNCdGWUBkXzPO3B/eLW504X6K7Gm729Enr/d3J1ZxzGj
ekJOw22NBtfiQR/+9Vt8me994yJKY9v7YyNXlnjIAGmko3IZXRN+o3nX7Hi0v0gb
QqLPnXMUHFp9XU8qiumnref48lD0Gj42ooIKDhitpO/hCMdu45J5QF/XkH1OcaC6
crOB/48S6qB1jhAKcemDqXyQQH8+shJvDIMTP7vXPCrolG46YnOeQHoJrVQw7owc
zcroZ8YjI2mV76Y0Xe3/RHEbJGl8+m7RPETZYQ/db6TMDCgIAi4k5Od2p21FfldA
nmDKDKOZaN/FOR5T7GZIo5FpQn7FNYoZqRf3CD5C6gEhikpdqxxvQaRT/mn5FEay
Gsr2t+Qxf8x/GSTirxzKIJX4r/Nnu8+21n0zpKhor+gSHup/K/SAWjOy1FTGEgIK
G3q1CB0YSyLdB0yVgz1q5cjotfISoXyRd5DMKXIaHlscDMgAfnjQSCevOc7eHqSB
qtRqBdKhg/QmzDAGaeO9r0mryVtqYm5J8ng8qK4rHgoS9Hy8d4twAOQWwl96ZF3d
IxHPq5pRvhOP7bK1v3eTokvQ+Zrmcsv2zRt4H0CyigIOuoe4qAeJWd3b5R7d3Kp0
vEPACqaeKpnxdXIv0pI1mpYeUvFLk/eVVr2PRsyWHn7FoQa/EbLKJQc2GuCyWvZj
HURd4I8EdsnTZdIGYLx/YOsOxcgFX2phjB3vL3x03cq2/LKqGygp/+tK9mOgFbA/
QtV85nyLZsDBy9bpimR/yAI14q4vnuhQK0di7dlj9GorJo69hsQ8eMsDSRLOz2XD
z2t5b4YKXqF4b7rLr9V/30UCAh23zixpxUWjt8rta3puIrRf9Nylo6vWSOY87eMi
R9CfbsAOeDuTlay9k80tS9NwLuBypGamKDkHq+WN8dKhUyekh/TuMhc0H06UL5Bk
n7P5dWktF6/8GmzrF4OvqqCw9jr7PCnTpZwtzoVWmX4DcVt6oMeO8eNPqoHMvOkw
taj1/Gzch9wlC2n2ZTQIZcsFfV3iqpfqlZmcuE/D7eHf4IeqY0wriyazVu6UGSiA
26C1qzdDfJMMVjcOoFx+HJWGXI3BikBFV+vvzPtXlKQTSXtuJu6plwjOtvU5JG1/
Jzdvi9t1NOwTzQJJxERy0iC2J5CXfrR7KjvF7lcd7048d0iAY5xDt3Gt8hccnXY8
2IYdCYq/rKOiVFFinE1EhMGNDq0sbHpBeKlWSA92WD+BzUm4u+4cCK1yW/2lJEhW
k3vcNCGR2HI+h/I1FbYOHl3Y5zKvzlRw3Eaf75a4w/01gT2RvFTIH6ZxLxsMM1MF
Rb7Q5X/4+W90KwOIvN7SCazpGsCuXudSQ33Gee9AgmcJ8wHcJbHI/IZEh3Yu6yUf
aUrnBG6uY239Sw2OrXa9G8QMkXpkUr5vdETaEPaOdaLjvM7y7B2ktuwY8/ucAk0t
4YKCR9vC5tGKwrlIw/ALf7If6nKdDH2QwdaNq5mJum8ulE2u+y+sDa/IpSl3WPex
6XQHmWUoLyzlBzOyX+hV/aGniDUdsR8HXYDV9z2fEQ6lQOsQPecTKLRMgbDLZ7uP
1G6/bcItGR2/HhDipj73QtgqKRI/ezoLxf4/5FmY85reI0qEVd1O/2RZ33VBrTdf
9860e8rTBz6TrFF/PcVbG9n0kw7dwk6IQykaUVjms4lEI+VDw+NxsUIQWVB87iQF
oYRsBqX++YbV1SEp5nopBCDOAZw0UHqmKwe8K+Wh18OO1XR/odlQALW1YGkfbJ5s
8jZNTWeSSGFUYsE3Np21WZz+IGp0e6RQ1Z53SzlJabANniX8M6Uqgm/r90l+NMNB
/bGTfWnPWE3pzyUhBskZOi7gRaV/sIcmVxvHeK+VRfnaiUq08Y5NoV4io90OnaHp
gjrVLQY07ephQtIJcEC229/szNmXh6C9PlAorRNx9/UUKz1VlpZ4OeRcMAFRP8J8
leF1BjobEN+lX7kWnJ/SondR4n7JIEjODtaSbzirdcRw6XQilfBD+iRBHnYchU0W
BIEiz2+7lSiT4w4DBP/Mlm6oXJ+x7a4XYzmwywHHO5PS3oBzkeCzTpNYykQBnCvB
kiBd2p2RXLNQtMD0BezSAiT5ar/HmMMOMa8ixoDxVdBnhm5ZrGO5Z8ofrgE5DAPE
hheP85Q5sbdsb8VyfcrcAr4iaFpVjZrFsLF0EL8pLw8o7pvuIjYs4DY1N3gjo7Fb
jZTJZGH/ASIefO1IqIm2ZjE8pixpV32I0NYuuL/AwHSo2PQB5bY7UQ4yyPJTN/HJ
1n1NotLXRGkUoSP87uqU/hrtxfioGafIRQ4GZa/lNfJPHHesw027u8NpfGd3CSQL
P739QiGaPbZv8xTutQY4dj+jm3K7HSnktar5RMWh/w2gBBZ3D/jLKnYNBcx4Lq3b
ZR4e9CTKmj1jS4JRkSs3sMa2MAJEpwMt+J6xHwKhF0WHnBsUMCmMFbrKtpFen10i
VSN1LCRbblsEemQIXdbXyEq0RHl2MRrfN3l9hyyLyqc1G6wGtDxCRpre4WDB/XtC
HPSZLbEOqxsXM7vzzTWHC3cP2vVG53S+OfuHTy/xyLvSBxAi8U35FeaLeofmDnG7
nsZFCaIQ96FvHzZUjPd4x4CZ7j4qu+MYSS4bsClojER5ViSmbb68MVcvc9yvNiRy
d5rz+f6NMyy1s7YzOgozMVD/huUA4QICGCK/esHL5TflXZe32yKH2L7pYWq4G59E
8423tAnDleWB7Rf+aP/pHRSYWmKLmEbNFkK8syUe+pkHuuPWinR+/SfVlJTbCq2a
/XXQTK6OY2cup0V2QDLd5+aeeuj/KuO518VmXlraJVvwOgM8UaIxMEJe0gnSny9t
+caVY7OZdA6n6tiF6jnfDlqnuxjG2ZkOXUO5OiwyaPAsodbnqjp9epzpEw4/QZKU
dGPOo7nKucb4f0Xm4ItGyRQeYdbbGp0xxY23nxOAnez0hLRuooB6+8ixEMtr6eJn
qY8k1hKWJ4kaFC3rOEA9oEsQ6SuIZLlx2rsyMaqYSTwJLr2/enVre02hMDypW/Ca
Hjgkgrb9qwP5UFjXODP0ZcgfzWS1Lh+ABV2zXs5N8UhhO1yNePKu/Zm0Pt4xJwM0
W8IiGYnXbCD5igm2ru8ucj73MknTVYRLUFbi8+aEplTqr5R6Y/TyQ7yts8Vi1TpD
nQEhbLo42kfF791rGFJc5CKT+riiMsUF1qLU5P3fEjyLEV/UJKMA4wKK3HxtIk9p
PKwZb19amtoqB6mToUUJKMt5gz55vlbpillzixPTT4gXGOd6wQS2tTneUqwuBrhB
7M/tHk0qFrodQe4XfitsxLsJlDZA3qFBZ/Qeu/rQMZ3jGBk9X/r9xD5EnZ6fS2b2
4aOMN4fA2fOIdGYoSgp1RQTPl+feqFA2TKc3n2vKrhqWSz5ITdna3OyYpIilg0SX
f+C6X1A34U7QcVWTjuOnZgTk8392b/knW6iPEeZGqvrgbgyM2kJTRJniUI43ropx
CDjJCjvBK1/aTVm5mu62rHemYzB4jf2syG/bLgsmyrwNwzHgbgCLm0zqtI7wwNMm
nkMbChQhy95vfHRS0vobIrLruJTw2WiYvzj0FUU1BEjUEsryiXiNUZemXlAb+Y5p
mFnaEF9SdnT13McjsSCt4LzFx3UHUqHQV5+StoL/hPaOudPnf9IljvpvRgyG9Ac0
pgo6OFVnEK/xGugi7poodGMAiYffxkSUjUfsFVXxv6leNRxSf8dF7+1ZnRQEBTzO
ZaE5Rh0+wZmwyZph8dLStBa+/OxwCPbrcu6tRJ1AaZCeNwOWwcsuYFuDs6mi2ZUX
I13Qnh/mpbCLudak8aBaMxJ0rVGxzo3lM3JhaMv0tshO/4lkDZp/qQ+5d1eNF0bk
MgRM5O+NZ16+1m2h+ruFpZD+26pOJQarmnwfvQx+lv5PchQI9lrua1loi3GMO7wB
Te/GSxy9emDjfhA0sAPU0x9v8oq42EUKC6jO9yIp7FqrpnVuIv1TawkgjzLDIgxC
3uEk5j7oxvQsfkh3uBGVEKmhny4hllKD3XxQRvDXxnXnKyPSEPb/7EqxSODGurPv
8mW+q46fupmHSxGHMJiFHKNB6GwOpEJQWfMJ213S0/YUbcXS1Y5Jn26vaMK9Dq6r
NGl6WZVtgtwoYQrOz5ghFlba8x9eaVB6PYORYmNtKXuP6T7MIjQjG4wJvMU85JwG
Z22HqM1zrGuLmp/W2Id56R1m9ZWgBydvaPsL/RPg5z6371uwMFExqzEi9/oH1N+m
UrduOyYgybbS0mIKPkqY+2O3cwqc5wfmjOmu/PZ8co5gC/kfVrTEUeSpwQg45scp
X29BhxM3VOyrff3eo+Lu7oCabBE5uQsIRpb+ZtUwIj5idswkAf9GYwDo+Au0/XkL
LV3wi4uUim39i2XjzKSdMVurozFwy9Baoo8m/9N5qM/mGvcwEuqs+VH/cxLsAzGu
JTKDF+RWSlgJp4LeaL+FGh95rA10/TRr5xOOfOi6MLHBYtHyOsdBga0FY74TDE6O
TZjWuznrZpp5xO9BWKEoBRlGf14B6WqFjmduGEc3HiPz7LJhtrCjXLGT2VJlV/0u
G8EtOMVK4D2EBGBa1z4w11gZXgvR8ynjyMbPm9i8PV6yO4tJMN1kK7ISWpws5aXH
RMMnkZ6JK5irfNEe5oC6zc80rHhquwdbANPFGM1s4z0quQDpNkVdhmpKpC/usWDr
nq/EF5mXQ2Z4sxqRUuPHTieeJfhP3AVzekAhbG5FzORGgJh3hjBYMPi6epdObgLU
C2Gq5p33Frjxw48yNm0zM8Qn0KlAOPvn3IivFOPbcCwTrkRTbOyTQ167bjlcly7b
JxAAeQu5HkLxNvCkIvqXVioF7PxsrGbSLxGm1KylOuInUwn5/9SzUyIsp/Olpcf/
nvRmbGzSUEspgWnLnjRBkdDr46TJ3LwOBBLPI1MJmjajWzdOuyXuxV0Mncl9xv5R
fpOkm7qgQxs+6dgLxFhailYOcnzjBqawMVCX2WPMh2b0zngIFbWC325GbX1aG1vq
rrD4XvxUC40zUbg08M6o248l4p0UK5QetVDx9b+0rQKeZ1TqbdjNOvVA3B4sNscr
7eVWfiQsDwTpI82tvb1eX58wsKMh1//hGs+c4udNV/bBZab4guYZczEIsT7udBky
J89+3rdHeKHqDhpKfxlFxkdkp8mhWkNRdGiYcCQEaL60IT+IDPEtyG7pilA2muyw
985yykZ/wLrzsPGRN4SwkcLlfBBecU2em3uetY8OGL7hHFX9eCEIyXVIg507EGuX
+rN3SqbCtYi4FmLu5Gy2w2QQqoC96wkg955EsG3UdQ+SB1ARjf26u+H4aQmsXdEu
GFDirqElXAYoMnfgSnNr+SQfShCl24aNvdX6+QzBRAEnmnJyLXY4rucOSe7eyvjK
kGMOYWb38xUx4jgsisL+nibeSJGfInQmIVbJGBfunxL0UJIKoDT+sGX3x075JQ6s
5uSuN8GAV0NneYi5k/EppXhFXnlLsyFLji1gvZbjLkOHzz4QYVoRv69BnlKVZtXm
UOZhqawsQs2Ff8uGPr+Hfi7VGKN4vrD3gwuxs7mrDN5Og9FFX1Yy6iDySOVPFzD2
j61Hx78U1nVXBQjmAiTshTJH6ycNiXH2gR6cNX76VxxsodphCum61kw8tjvSOXRh
0BI6LI4N3EK72KH+jCJftWDQVQZGEmhPT++FK6MngbRgagAmca03PRagWAhWpOm2
mQ/mlfwvAn/xSAj/pvkSUkQxEUBaqHXnaDPFC3CaQsRM5aMD0Jag+QmoGPkgt39n
WHIgVnY9ecsc/E3MD7DnZrSAwHh9V7S9L3xgm4keQ0r06ews5dj23++dW8dOgCbe
sRek6GTikIqa7kXIX2aTwJep414Ow2kbCMg8ExaiBMjU5HzYahESQXsqgUBtN9RK
t5LP09/Vp/30ny1O4C+hpdgQth3HfQzpAPkKZ7pGrdVs4Sx+QbpDPdwo2U8F+Oz0
68WJ53ZglT88INU40ERg2oN6FC+UySjfMtEGGl5LcIg6t5eQl8M0NtEYecqlVsOu
sxM2loTr/0wz8ks/cpH6eWdXNdaWYCebseB+oTUgmF/S6030/xhAxwnPeus1lQkE
Aow5t5XH3JgXFeP+AkPN4uGyRliwKTV+a+j+pNpZhm/BdERLI1eecwL50eb4LHq8
zAYqJ4+LjFkh8KsKP7ABGc6rBgqh6T1UObLAtriZHY2kCRW4WMqBkA+I0sK0iie7
T/jIlq83QAlGghzfQFUpdebgNRem6TEl+zfM1/oN8K7+RTNvMQoXGhRz5EGiQjr7
8+YGMzYD/G1qJkINuGRZgcCRhIlN4aAerlMOU43qgGzc0s75dRYC8Ye90lwlFijX
AjiWdAE6k678Va27N5T0z5Z7UzCYHMr2CljXnpB1w4XjYTw9KCq3Wmk96VU6Y++F
u/8QK2PjfbNic8WJBzsIXeroOyk25TT1cGsWMtMYlYKmoSfbaNZNiBwrarS28sm9
jwsoh4XRtB+RJE9xzYojXDqvccJtjueKLfzvKbgQuyIgzJmvLcVpnGZWkSlj5VFE
hgprN2JwrRJ1/VcAhEr9++pK8x7N+K41tzWqfYer8++nwkdquJ+1h7WdDd/kLBGY
2Meyty8C5M4UOsMbcbVFy5P3tPw34bETeaGA6YFskosSsWFAj8cKcq6B/DJb0XtO
nkUlhiiZ3DVDcY5ceESWqXkvI2sORS8/UW3aNPUEyVFUDTLUR06G1pPh7UfqB/Wr
GCyspicz+hGDeyLAFxa2Ropvy3UgDoMFdwYZaIvTunBn6ia6OaweDap9jIeQFVhA
GXd6qPTFkRZPAJclEP3P2+cIg8H51O2701sAfcpsb0n27Ar+Hc6gKqxsmzT5UQS+
0Mq2hHAc+ORo3oG6Z+LwRzVmzgC8xP8yXcFeEuvjFzXLXs+8OppXbn910VSVwcez
asnNTw0EC8lO17bhV+NJRh7/wg5JBvHLr2mGBpOSb+A72ohC6uQasEGs1e143tcY
e+np0hYpyDexAHOiBSLcn3a1LBay3C6a/jYT9uDHAdNFskYxhzesWMWL5v36vkd1
Uw21SKfsVpSUFwxBlAE31i3Ou42UVNvz3PtDNJB1Hl359OQChvWIid67plvoGFIL
mZbshSQTuTDYaY2vxfZIXX9bkPOBTZOhmZb4U06G3PQ5nGsTIRdx2rRktxeZjGDf
2TQGzXKauHE86Hdm+05SysOuD/U8SHDO7rD+/WEdqgO+rmj5Txbp54nR8AUKGc8f
etQbRef0pVhr8q+AaWNS5E9pt7NfLC8XYno7LAFyb4m3pmYoP0EmJrRmHqi9ILmV
9gFm2dtWL8Zadc+9t6cyHyNh4QE+GaV8KuEemAoNEb78NwOH2x7dxZmuCe2/x90u
ojAbiILOVoF0GgLwwajrcr2qnQsUkMPIsm4kOfO70Nu2a8P99QFxnubRja0pdHUf
4LGAv8k6vjl9YgPmbnr3NwvclwEGAJU+HalsrWKV3vh3PgjvwgoB5Yzb9U2Rp7eJ
i+BftDY48P0b1SCwuMYezCcGkDKVEGHrE6RwSlP9uqOX0x1BG1BXMSoIg1XarOQM
ruWyhJ9PDpHaEMgyXvI08INLxVgGmPrdc4PVwy7uqXN3aUU2beaerjXmgluHO3Jc
Uug4ys42uLC2fE1T/kEACgXZRi5Sz8VFIQAsGeLX76FfAkXxLngiljBFQBzYN48K
pEAirCsBgcj9y+zsNEyp084/c7++JrnsiGgTC0zRbvBiP496KOIbbWhnMDaUEQFe
v85tyAEOIkhXEtmxBPMdSlg7s3aaUeDslyW8OFYGPxxsCwmBo0v8zABQ6/bx9aZ1
Cb4p0AmrEiq/V6qgOLrtvydO5sQ6csPAJ6+yx9PU5Uy6u1duRILqD1p+zmnXRHpc
YwNa9bCVQuCV8xQRHBBpegDjCCl5Rk06ew5dxEprPzkFt9eFtiyuRZpqQL1NdtDw
qapYuW8wfjtRX876KfoEQcjtIow1LIsS3PGpzvQav+oTe8llU9tIA8yMbenCDpjq
2R9vEaoMnBhvuxjSOQxYLBkG09DfChPzT98wOar7Q5CO3cSRiuBl5uTZVQ0qXHAW
VqaBosCu8uy+alqOt482DZvXhPJK6iyPsMC0QvdPRvG8JCz6JyZx0kBBUlKnrThn
IaUAWI54SLh3OvZMoogF7vWZKng49TquX89/IC7SkkfRIg4uNc+pgGFF2jpvoFq3
lO1AweClbIr7sXhXWOoHZhNOLx41YYwpdmGD++PZTpxM6X8tBQeYlOObnw2HL5AQ
3SzUeUjRkCLpbdMH/4ggkel+ChwKAUEADjV75ZbLng2eOY1IL7OvNhGtsebjr18n
jujda8R6BCwLCAc67wBBs+47FInLhuGH4bZ1Q/Cz+Y0j04yRXgL9b98sAtUDsKj+
/tLvGotf2pzhpSNwTf2JclxxSxHnpQ32b3PKhCVZ+zKYc6pgszcKQDTLImtN/01s
pHeBb4O1Ay1n6D782wepCSH2I4pL1NCc97un5Be4MIyb5+PvZ8x95372tHgKsL8X
lGuo3Wl/jW0jiNGfsJY2/nNVqdTalbHPKLhIjB7bMMpTadFwX07L76V9rsEo8Fr/
vEGkpPIDkOwQNo906ZAq3qzcptLqd4c/w2lbYVVpuK9OgmWsb3RYPaHcxTEokYum
BbjDAsdumoakUNNL+O/UWouT9LmFRGhOIC9sb0qAgpNGJJORZF5KopXvhpd/V6ev
fKL737ZBmeM/BgrjNew2pW9c65bWj1GwfeSAIrRg+wxrTV2jPT09HNXHNgfrlF15
dF3SzdEbM0PQ+QkAKxp7q6QzR60tcc/GfdFUDrbOqZ1pS/uiN0BAOQlBzk+ELuok
ZXA10TYp+FS2XTcEhQaMY7vfcfagh7q2yvpmlt4/WsWybtyQnwYIuGWpGhfUkTP4
8Nnn0ngV5GXpEAIcIXle3qFMSimHNcxnlioc3ymA0iG4gm3SB6OSUueXovwb8+Fx
exUx/mpZNwi+gPWWjf19jmKGqhsx1T9STRnzKF1XogaY/kiaTX8PLAfRqctqlke9
ihWo2qg9Dox3dTvBdzNvtGTFIVwZG7dqrDkWQq6d1Cu/aG9TJg0i9LTwHfuPmEuN
i0CWbQ/RCYTjMn2kXVNrZhlN1Yd4DGDBlOqKqA9uIhrVmv2JqSBu1ZQBSoIQCR8Z
a0HGTviMg8ZtFZhz/c7rUGlariKTbSsNRTCZ6wUlCKjje0LpxcuvhUXPMlS57Csn
+d92EI5mIarI1ukGMJLrfoMVGim2iy5T8VEczwGixyu5WSDkW2NlKyIOwGKrek+r
TgvUP7ibRlXvxmAnJOtmCaK1STuE7IilqMCDoU6flqiFOO6s9VMALogU345luGaB
diTC1mUBY65u3vKF9DNB8mt9RUrGQuskZsyeqwcp2JAtpzj6bgRioQkFOdTd2qkI
RVBzJ68RtmZKV0v2gShbqt3RGgDHms0NO2EyD6GYutsuRLqGEqDQj27bxp/JEQrN
Gm2WGnEubmO7V+f2K/m5CeVUo096NSQcKG3F+V5uuY0uXFSVnUS1vHLzgKrV2hnC
ZA7F3P5G7Mw7dtFeUbxqO85Lnd5GexArwPDXgw6/dRu0v6CqJ+18MdIDys/KEM5x
bhj/yS057mM/jRfThbSJrKwRcBaWmFJuetuUBSRi7w1lfsrCCvT9VDuTV+53FnVo
9Vo/1IiyeT1GAQIU5PUAvFF63zZf9FvsaqP8azPG9q9pivcDHdY1EEn1Lzabvc4z
ENS0Ifl9suTlmHHv76ldlwDWnWYqO72yelIerc3rREcCapaK9BYyk45/NCwMsjKK
zLMMprX3vYVm4XsIjNGb5YYMMpRXbZfPn76RVHhVngtcayc7wWl1Bc+An01POsCi
EbauU0MaWEM98PpXaljZ2ufv8Q8X9hEbqmf19k/7YpS491tulM92TQPo5hwbWwZJ
g7c19hVzfbcrO0v/xvmUAtvRLOGsluabVoYInuDyK/Tti5dF5BHBxmReCZGK2dHl
yqNZVAmZM8Fc7E8MFoOIp4elCophy92oExX/zz8pl0PIrVL+2aJx6Y0P0UDRNnLc
xDtwrpGkEXOxEDpWiJgMZfrDzVyF0vEiA03d5TMDVsrK5O+3IYTGzvyARlsjp9zs
vFq3xfbDB2BI5Ym3JEBWyYVA4HJZ48NbZY4MwZA99v3EAHuW5MY2jcUn7mtyXYYS
uy5e8FLORx6IpQUdTLYtxXiPLMWjXAglN6AGmuLSkcI55Fihn34x1j7QtmGCPvkB
6bxA97er3HcR/wU1xKc815cQ5e/xl+Soip8DQTzTAJMc19DuS9uYKqkHcnnSJcAX
qhl0tSeORWFjU88kQmSHUe5yVuxvy/Z6b0CemLSAMoervnYiwioUS++OC+WEA+zO
vTSVdDM14EYU1BAVSzt0bTBrg9OYq8/xXDYxPSbsvKeE3dtcjF3MQgt06i+KuGwu
4rzuLdW55cnY3CkHyxgphAiSG+M1bLfNGLhUwyJazFewNudBtj3DWUmtd2Lxr+Fi
USwqd90Nw/76HB6F3EsLmaL0tNjHN7xjGR2GWk5IB9hOYK+gZLut4PL+aCpeY40Q
0wfa1+NDt3k4J6t2qqfb1Yg+c/V4D0CjjFJxAHuSdmAI6OPIhs+8tkelAzTXe+Ye
sQHjppJgpAGxrTLS6+8gU2vpxxUXwI/tYUS8PcC4yb6QH26SbmqH8zlpaZHSYH8f
L62bYiygqtMqyBA+GAr5l6EZzu3Uc+DFzQbrYHg7Wd4IaqXHDSPA6Q2tar0+DVb4
mN3gVS6KilnPUvWTkj+wduJLfeqQhZWL3ntVZeZYlJ3InnML4ocbFHi6YcxufTfU
O9BwMJeQNhyxn09+p1uhQtEshBftqOFhu/e/nfZooT4pIdLYQ91uGSoMsmFtxypf
XdNwEWBTFGvlqOjbQa4FKwUdlK7R+EKCtHf53hgS+vu0zz7uf/wPP9+Np55vgTcw
d4sY7lK7GiQbhCRdETvzpswqIjyQ/LRhpJHqDuyQGZ/mwy91MXMxyHfccOoBFIpm
ZNx+vE6/cO0vN6T2NLFtekVUdFaeUTQbWUjPfLZN62HQ2Ov0p/7CK5eY5nAEWv9/
fKP0o5xj8PCn0abfu6SaqT+b5pqV4cyX3Hmk25J1D/FiS+4CvN+EHxcd0BscqpRG
Y60nKMITXvzWuZnHGeS8GLIT8F0U/pIfxHUQfVK387TJ+ZsRPlP1sEuhwE93OUyq
Xcy+61b7ESKlldopcct5NnsTwoKfZ/6MKoWAZQP/p6hqQaM8NVSEtB/myZkZG9E2
S7tt8Ni201qKUTVus8ca7ZIhf2iEj7cA19G+yVS5NkmPgPzn30JOp7vmmxCtipPx
QCINHfp3CkeNnHGG6slLDACwoJPSatL9athLwhOhMwtsXuJCEjm/miKc++yjPCuR
TtME4W7lhY+FN/ICU9IHO47SRpgp3ga09XHW2aAKyY9ezbmNgSQARVM8WqpGuXwA
wxlZXKJblZaC7e+x6kVpcz1DNlyKNnUrVUnqFDoTZuK9NaiPfs56jHy2GqsJZmS3
HVq1BqdvtrzcIWPd+Hr49C2nPRjRAhYa2OQLJZZMB1XU8vXYgOoQVJHbIw9VSvnf
AImZ/07m4BtGtCHrwKglMEgqAAix4ogxP4yg5rFCPM57ZONhcPyca28V1eMz14la
G9wwbFs5Fv9g3En8a8xslMiSUKJQEA+h6iMKtaKglW8GnNgIzi1VM2Z5SXQSFWSq
icJOW1TMCEJaCeb8YYDi4KCSQbZ0B2yMgb2+1/ck+cxJdkaylmnI9rZ/KuPC/+P9
AazTYW5OM45WbaN4f9oHKN9jMRtvAeZ5qbeZkdenZN/LMzbrL9yOCtWEpnZsvr0Z
U0VHxpDDhsbW4RxTleT/RFEKuoo5GWwygHgKfpG1pyScpiU8k7WANILYEhCVjGe+
ZoFxiwYEn3vQcrm8TO4BZEugwVUbge+31HBsHo5fOgeWJbr8ILwnxSRUvJpRdKF0
ua6h6MVr/Sk0f4wHJkB6781uPsjn3Cwlw+thsP5x7ViWc3CW/1v1TZ40ZW692swE
ht9hkQM3vL3ZmucnkdDosGdC4USGKqYrLzn1nDTG86vOXiBgl8VncmgPPbqwZ6e2
E85aNY8TxQUZV/2RWw67Y0yxmGzCYvuGqOfJHcRz1lgLniogDi9es4zETGCYoIx3
NUAO/Is1JMsusxGTW+NwH/41rnL1PEAaudsooFqXRirlUDtoP2tiYl8PMIbC5u7Y
rKTTcJut0kcUNHRejEgThTtPbFVc61w2ZXffT0xVU5KUQJX45I83PZdKytBzSU/s
fZysbkhK3gk/KBxXfNhbIrfWuXJb8xoSm+qZjDmaAbAvcIsKWGMkze+scvTkyULl
FyH9YCteo23z+NomGj0od5l7ziM5kzfUEEdP1wz+7uH3Kvy2OPFLFiXzEl3LJP+N
qEgcYz/PeIw+bZO4aZUpWIRs2LyO9jVbz0uKRikYAAFB4pM/lXtnzaIDR1+kmLH/
tzBqIUMss5e+D+kZOEKWlkrylWYARaDBECZi8Ng56XlkK4ftL6AbOw1uTSATfNBS
2BV/fy8j+hW4hGXG/KR41S/hXxFzPpOAnPciU++rRoMjuDueH/G9NEFlHFy2X2E/
gaKe0TkQ3b1WUTXRZa+TQ/OwLt2Brtxwn+ELUa53TumASd50tnQkbOwv+8CFBzUq
YgMc7n/NSZcpbziRGoxwEDM60qDIRFBuNd/Q1uCFvVoHJxKePcLIfaEcMaCthRng
vHKW1x/OEKegRrVawVw34Uf1gzAWFjF8x+vCeHIojp2VS4jQtQELaoWew+wUer3i
5Jy9OpsYtJxOcTYf/n/uR4lSUbXhXu+Ul7GDm727ZnK75kBiOOK1t4at4FfzBcgY
NFas6kv6zyNCJFGat/N92oXBaL0olQqre0kRJUZsU4Yoiaxj77t8kj6EpHr3fTxu
rA1brwdVY3v/i05pQByn8qZKZOrLuvIQrNRw0ZkhUtFN7SOkNB3PWHg5/QZPQDY/
NGHEOHynJemdeUUl5TSE3uWiU0Zam4hR8meeZPD+jc3+L9AcXOiyf6JDSyANZDhW
vj7a0JAmjJkGdAcrthp6wWVZ6ug4IthrO/tBwpGnjgtM7/uvKbO3J7HaDrvuRG1T
1ak254QIDmVaOmauxSIh+JGTHwi3XoSOHbTd0ztYRMr9f33x3Q17PfV+jDWSzxf/
fR2eNkyVj1WHcIHK+eUrRKNoOvQNc02vaYePV7sgKubBOvSMDOfrdZrN4obSQMnW
ST/kuho9S22exoIDDQ7fy8QuCZFJ3TIVDr8BQbvwJcT7trKj1oncqLSdzOKkCk/U
Y6sfQysraAS6SrLXJ1Aku9nhsGygBmtXcpgBR514lqeaNRcKMY68/Oe0i1wR41X2
/QSrgKCmDDPfEYQF6+h+/Pn2Y1hBIHKcoN9pE+LQYebFf3gpaZFySfr1xevxilfD
MxJJHtKxsw6ZWIuE988inqqdE4ycDNzPhw8jDiN2B1GaWklbw3o+w5WfDd1zoSdc
gcky3crbpjwTzlma7z5SrhlIlYdOyZAbpKkMbeE+CI/5Gac4b4dz6sberTjQsVAz
LuK3aLaXgSzJrPUZT+QO2iKFf/eWffYk4VQAO+2t6I6Sen3Jvd/GiCRoj/KePA/D
zzL3sIE/Wnxva91l3K5jpdyFqwjbeZbSWRcZhqXQV97IOIIb7Tu6W1GNQlJmAaY6
xHKeX+5sppTaDB09Y0QSqV765eGGvAXOSST4wa/IYQJBbML7CV+So7ZcBGBXiruR
WsR/cL+JQ8M+o5dRFvNOwKVxFvQv98mVoorOrGy7VMYSZCrXe8D12l1IWhmDz8/v
wWZTHNwAWQaReUOF8IL7ewhsjcSVpIjgQAX64Hv5sVUBA6xqsWD/zkDQwGkxMZ5E
oB6gbn9AMOQVn/WNcqnRa4KUrRsw4sgHDgDuzzOYCAHffEUZfcJ9Pz23UtQuFPWq
CmRlN8GMdiNnLDf24azkfvLLUjCarrrjl11PfaTEsfgpSrNljeLpBT+uthhdU7Sz
OByiBzUOF06X9oDVJIM1chzJZZi3sB54/YhH3lUFeYGaYbFmq8NyuJyhwjCOCNik
Hh5M8leyDIBwC9GivpkCm6mm/vRw8jMHK9hlyrKDip2tjX1TSJjeFXzN4bfH6wby
UbKw5KBXI5S7G54bpIXlGcR/to/MgXi7VGWunZR0FXDAO6lYxQYjMS9mhpeFrRKZ
2DnDv8741WLIehoknlKpwAsHbVDIB30E6N7FCQFcjBmGIzlyUmYm7rawJU9L9DeR
/ZuGbmOqvm1yOt4wtZvkjKnH7QKNSQ0scks4F1I6W+jtwbW/SnTKLFZ2dIRAfbzL
oyPIDJ6cw+qhRXSChEjRvKfM/ctv37uaAeAkQ5gUxbzxbI8Iwq4nKofB6iWNnXNF
R3Au0qhFJCfZKvxl34s8m9ronLzPCRjUB17FtFfh4tnPqr5FFicl/DitUlQJRVgc
Jt6ZNlnGD8eiswdf8DXbvSzfQB/1ECe1WJ8yX8mbyH8ZdiHINCraySiZtk3k3myT
iiNuIM91VpN7QPtVIbTqJFGJQfMXBICdLDZjRl+1agWhpHzP3H44HrhVqiulAjm1
t7y8btzylEA2MB4cbpQC07T3y/6WfUAYSM0tyNTxcRfP/4KFQpJckANgSoegF5Mg
OAwUAr0deLCfMDJCzs9vJd+fHUcqlDM3WtY1Vt3K0/DZtJAZr+gaZkHMwlwnS4KG
qOsn38Ig+cEDM5L7XYmdDyS+MxZMjFW3j80zS5gRKKbRFiD6wS23MaO55l+R4sKw
BwDgSDKirfxI6tVnGtd7o9Yq3FclTaYzZIJGHT7PGXP2EmAQ7Qn92tbYQZzuZwbw
poLX8VhDPCVRAbED//NlLP2oTTdZSqGk5G0VsslVYX5TkXgVV4ae/E26eezosAXy
+AneIaNRWu3xBCWyK4QBi2ITtJfAOiw1/SK/P8Kh0Ihd0RQjkn8vbtBDpdolhKTk
TPEMxoUhqYcdTN3YyNtn8z4YpGmXNLvBJrOU6oTEn+7BXj6EOOIemibJTJvLL6vs
YQLJq3o/yhiL0Ur9DurUF4HwkOGSl/yDSXgpuDs0RdfREanE8cfoHB9HEx5DdsD7
Nr1+XwPwwiNRiVrit/sjDp266zHT2TH33t/gRGhmXkC5i9O4ELNuLtvYvB2bO8Sw
bvjgVehCFbxzx1rAFCtEeueE1XsMQAANRuQu+eziww5rlMSChtb8uz+TVPbArI8B
GvBqncMAABqvUK3E3QkYPDIRBudcHSCLQ4fWG9cna+pe/pkGorYw6bQ62SX/juUu
w3fsNsfeZCMrwk6VybLjMC6R02UX/rZ++jxE9NnTJ1zQ4/zEyMQDnFEryu8EF1b0
1yLHygma2i24zygv9iysAvi/yFGPHJnhiJoLgKFJ5nKaGh6CxEoV0eHM6kIvk/IL
Ul/NTnCUKHJZMm1H9/K94pBwhAwnA7Jw/OTskVGHgI8C+Ds3iQWMleke4GqEFH4E
DJyEB6u/HF2E0wrfVRSmbyCKL2XIYx28O0ZbrRsEIdiScwP+yHvyz2uJ0zwRPnVx
DErC7Q4SNs9RkB7S7F4nJ3LlMVAYBfCWDLgAQ07+W6EDaaU/KfD7CgunT+pskpm2
wvQY7k3v2ByLK1paAOCh70HfRL/ZT2VWWy5eNfpVT4wA+Ot5/gAGpWsCn5Hvp936
32EMec+RiVi29z7MeMA5X1HuBXa8mfCrl3iLgpRtJgW1lKKtixerm1o3Th3qDc8I
PMszwyOWOZah0ruVACQWVqo25XT3eCANwhLUg/bADACr1WrWDbM11zxqFyNAZ/j1
C/8Mr4YbJ4ehQPqMDg7g0oexpOa+3QT7nb2EyUXi842wghdVUOWIe/t6YTFP9oG0
7xuIHgFlMujUqeu7Gj4OmNb0gP4VeZHXddUAzIQrozlZLoTghR6l3qkifkB2lg5t
nMopgo11kXj64fEJtBDQ9wNJ/Zsqc62KI+5Bsj8wWp9BHrjGRT+B6YbUOb0tiX1y
PRXQYXPep62tF2nhuoom9REkCvysDFXEOxrIy+9iVC9zg27iY6b/zc6faO121drW
DhstDm+6X/B+4UFvW8GGML+Q8pJpUHXSllqIyx3SMsBFb2+4ijr8rauseZqMr/Mc
21uo9XzohUConnj3awKu3l0+gMGmkCiOaQbsN3J9KlJ7P3st5L8D0doR5encf6GO
6cJrzHs4RRM83bbRprV6aj8BWFvIGgdR7sgcze4J8b4ZMpAM67t6c5sMH2omMBOA
5tdx1y6Uw2mNG3NZVfiTqm7RCw0RxOdc2yPhYOYwS6FBypyGk4d6QBijx2cP53QP
lMWbF5ZpPR2JvbtesfeGFIUNwOLfDSHnxg7QZ4CQKG/fUX7Nv8SP2F7CD1yw7WfU
TnNHR2BjmRdeYDKDi0ETDN2fayi1YGchsqiYP7seEuCQT8XsbBDQ0UOkhDNl8OgA
9ZT+votVhciglyKeQUgXJc+mLQf4RTmTssz7WB3xWBtIHb6c0Aqxtz3rWY4FwaVv
oVNSWOOeeE/fdF91wDb4W3uEq9MuJc312RcylR4tL+Q+FqkZcdJ9lAJvpBtuVnNB
kXlKKkTuBJ/+evKBm0zCHZDUHKJZP2XI5CH1ESHvcEyEcG9EWnvzCIACA1O4+ugx
sA9FcmY4nXoP1jRHSmW/OGPhZaEBJNf67TLYPn/+elZMWrPdlZ8AfnFyyKHAhMJ1
hSitEQgMwnnuah0v4lddddjMSCPzDR18L8wbB9597lyc+BOPWAxG0QA5jX1A4w0P
TDi6aaC6Ki6Q0aGwYdip+SBMc8LiFAcTR9RNaqgaR1PQJ0VdQhrhyy/syv/gqFM0
ymxRUDl9yseLGIsES04ufbTquaaEvcnZ/PfFWfkLAStgUzih+rOkaWowb/afbPup
IZMHWbb8Q/rrRFsBRYUigL2gYiIqRLhAjAdmvh1t43esnYtCfSKRMVxMhusrCufU
zuWtIs0sI5QE/JUZ3HxTC0+ditsQWqDHeagqBS7y/wx3kir1h46fWxTbRPQUw85i
3FAgmmVc079HnyJHY2dZHVOpazcowdyKPjP7LqGG+kqv8OQ5vnYRZ7y7n6BnIS38
bREMNQnFxJeR78NCGHnIBTlLG5E386Vo0VUzIMKfob2ISWKaVHvgdFVtMO3QpUbb
zGRM4xZF0AYR8sVYlA/Op+6kxhx6TgGc3CYpdOK4K0hcwKNawRh9rHAI08HZwwS/
tmKa1FL6hvP1uH0Eo1oKVCqHbXpxsqyERnvOjLJ90OkGZC1dmq/MrfikVg6Oy768
kf/UJVjyVdNJ9p2h3QCn+4+zGVuo7lHjjL7Lj8saC3eQyP0JXfE+WCGksHPpxKal
5McHFs5r8ZuU7x3uZyqxARREQK6pjH1HPtaCf+GbhottiUFKazKFoqOWiL29gKOQ
QVOr+2cB/TE50ESSgIKurSPmBpROetN8bPRHJyH7NsiVTn7rPqREnLuIfrfx8vWR
rqRbJ3QIRlWXjNHIvc+UlFdQlIK/55AIT8UFIkRtGJGfnF94kPis2XMecN/9Eh6i
7wt0OJf3PDJWehP0d7fOl9KYyAjl7qW1zJtGgUsk1H4dxk+lxdMsIEVhTvFFrqkW
GBV3/3/Ov8wJbI+AYbYdSA2jmkWDmppjTLQcR02opk9I5gR+8lbqpKTwjaAXc1mP
C/Fc0R6rVouC4EVKHeBh+Z2O3qKKHmx7PWaUf2xnhgy6iCGpBlq5X6ZTC8M2hX2y
O00C8WYr+5E1/YoyWNieAKMqLaEaDY9pfwPteG9vDbq0tMpU4ZAGKUXeNYNvrSMd
X+tQyarW8M8BjPYr1UCCCoFEcLOkEhOf2EvmNi/szqDCpoxgIPaKESQ6qz4FHeXC
UfpijYfpu98NGgjh1Bh/Xoo1THBU1tG0drwqzYJ0uzbvvIkNZBXgEWB/pzI/FUSE
qkcbwdaCIBbPQRqkDfQFhTGC0rw1TW5xo0OBNKARSj39CzCVwajpupr4qulO6f5k
53mVli4j8LrUvmtIku791F62ouwG8ZhvY+M3DpkXPF1R9qPBjm9b/oWaq+/fxD3K
iaZWAO56XNb3WBW2eGcQiDTdSlG8xHzwc/cOa85DBq5D0gP/RLbqweYTZoDqG4tb
S/H8B6tuj8flygdCswO5kFtCM37FkTA9IOQXMXSlganIrvEqk5gM3SQLOXAFWAac
8VUttYrGtgBRp5wRwB5ZiFTff+XAl2Z714gGFdxqiAyBv2DyfsA1VTTu1/USs4Y5
3Zim3JJ0mTiS7x6Zz7vQ6CU/L1XGh2awnmxgIpHM8SZ0DkFsi59Cv/lZrfemPsaN
r9XYf/bDjOAQZAuAQrmg6J9z71GVBjqUNvPK36IA5hYO4RyCILhsF3Yyw+mrR1Mp
R3NcNwDSueuVtK9H7ftwWJ9MuWf7lvk8AuUoWEGmZuW6x2gdj3bg5ZM2anla9O95
8jr13E1DeeImegaagR+nKIWhv1Pv0fh+wfVoSe9f6CSQqkGy86svIVvxGeRAIyMe
J7WdVXX1ssd3NygXKN8e7mHSi01biZVZHDp+55Ox7p3PrCkFHcs8qyP6rUK6Vxer
ZRBxp3EGxcquLViPHEpJ1Rd7PWzpIiJgcnmXSjsaISXqFwasyotlD0nbVH5OzKwj
mAUIq5+o7rfJsOlcfF1TAKPDhx+CZYBUTqtaQ6lJQKe+cIxqbwYN1xIPWjQX5rtg
+dNRYINlsJ8qrEcx0Ctn2tyE0CtsPKa/+hr2B7mm/tWKkOr2OhqPV3ISfCnxFETy
EoWY/rrGvl9/4NmdZGdT7SGwjs4e37VtiQl5HHqtE75Si6qHI16lOOGKU02SYzKq
9GF7R7Ybt9GYf77u/EwXdgvjBQUZvcEKfP3AdMX4r33bdSW7C0F9zV+BJ4SXW28V
wqFujOmg9rfXodNi3bhN8qFbbKMndsTpyKIFHmflKx/7Caau+wCp60oZIj4DpglZ
j/BxFXqm0nqIwZgf97SinWdBsCNxl32L7VI3fjhG8kwkrqSk0I51h2WBSbstwGsG
TmC12/fDj81+wlOhnwJ4Y2EmSdaq4j67dxTCqxh2mIqKwafCYs+KuKzpBeQkjkvQ
M5c7WWVPlMrbCc5aT/23ayrrPbcumfwQd4dWzcAHU3mD1XlwNJevVlmxAAWv2MOm
mpn1pIZARhsMolLXMmsISG2zwFtXjGS/aFnjQwW/86g6gdidPzH7TWXloBag8yxH
cQFAnqMqakBoex2WPHWXAnm88/I9ZvLkxnsp9l7yBf/t4w5kRxEY94InXBZ/yk1n
BRWSVRYERvsiIbTb1BGIRPuk+I8HSTX8FCSmqA11EbCYBggk5GQOszdv3Qt/hwew
cI/+P1OJrCyZAlxqU7AwdTRJZBMXkLUZiCaXWnG1ubb+tLXy2X+fs+L8q2MmQ6XV
tJYXNd9ovduETThFGN7kncL0mTZvW3P84RZdlhcKUCh/wKxmGXbgm2eJOUnWTjhk
SKJHhx/8S4/3N8oj2OJi5LVpcrJfno4J+1rB5XTCy5FCBvNcOnIl23CUFv7mt/oO
RLyfK9Yo8yR14lR5tMvhhIGC7FiDHzHb4ZkP3CzD1adpynpyUXFzhCwFWL+efAiZ
c6/1ZgofKujc1mWr49DZ8kFS4BQ6ey8fsJSaRUsNSuGxEoJKppPqM9fUFr5k7d3F
mC0/6e84FVW548Y9yZFvnRtQUky2QzyNSaen51sG9HNnhvzyWzk5tG3YmN3xLy5b
TtJZesSM1LNKMslAzvQfh81bxBNnwL6IrWWGDNDKOvP8VljOKFxCznbxeD8arZYU
VkRcUfIuUiPRB6B3EmkQZCt//KkHdfaZbGSSbZ9TsC7X0FdSRNcj42kUURFaH86j
RDlgbtoNLvgQi2bf4nRY0pZckt//RCXO7QFC3pIaUqlCKtA6z7qUkEvSk/NjzRv7
qD5OcnkQg9a8pLQLo7ZgprRJ+UlzDURF4FHAzduY5psPndGyNLtXkH4LvYaVegfE
PpErhpUxEO1z9nqaqptmz8oZgLeFlewkJqOJ9wDUW7lhQgptGAKjh0/8uCnY+NBZ
MfEvQ4qXgwWBjKn7f5z7jiNS+NBKBLw1MXZyAMfr2r4LZbs6qEmlhdpitRfZlqzT
XV33iEd0eGaA2ZgVIZ3bGZQiZFsNigygSUzDW8cjZ/wWwTPkYm4PcHEwTx9wiyAY
fTy25KeKc5U4zm2zY/6R/mnSaiKr6CaEMUf17Qxu+r72JnpDs6NX8OBWcAc8+dhp
1D6WYkWzCwxUB/Xk8JhBmG5DLD4w1ohlczgNwU6tBKJUccfHNdVXYRsmPzXaifCq
G88k/N0sqPjDymqqrHJuyCXXPILAFJMGuDwDohKGYPbjmRlC6cBpPV9X9Vpe7vlC
0BWhTUhdIKrjkRGYMASSHtQqdop5mu01Fnbh35NhOOyM4t1JIs+99U1I/1X/2q6b
3nroNzZ7PkFoGy6vAPF9CYivt5GkFNHa71b+TXyF3fHh/Z2vtAoLip26oNpyQ9UE
Gnqx22PfGO8Cp/Wh6HxCcSiWzwil4olZVt5wFQspcr/NZTTUtjnAaDCYvnEAkFPF
B0mNoDrZlhEoVLK+PnRNHbarX3wISkS2jB0AMff+rH49i50oRX+xQSU+hpoCvWwB
fPeUJCiyGkLoqqtQTk91GzcpruPNj2fYUS2ED/f4WB5/k69lUz7baKQjIIimMfHT
a2xy7vdkbqr2hgWrSwnwwluJ5MCY8HHGyiw81g/qS9XZ1SKeNryC+iQqgtMdwpp/
DrzGwYcaPvS6qa+KVhJEcSxYbS2ybLlVEbQwDTAnRnSR7VNWR4O5mDUyjPukmqkh
aZmYUEMAZ4QALACbegypBWDW7ATl00kk8TKLFPGvOmAamNFMv9Va/WS5gIYvs6Jz
L0fyNhxCKv1hIlsCaxnTDMuS8dqfC/XAL5qlsCpBd5nLdjeXcmrswp8dZrRqrc4R
qZRFJrFPSjyWARpJfuAK8zgi1tivd4NVFX08WcOnLa4cRE23GUB1In4vN89HVbxl
NM/agUiUv+OAP1oV++YKvJ5fQxtkHq6KubNWHEjvL9DWkCGLT9wEeT1/NFY8GBM3
1mLuI8cqZk6gPKRbEIo0lsTDMTOSgO44qZv/7mtKrhqBKCIlgO4uQLCwACQGGCb6
AU9GtRLVzhh4s6s0i9mgM+1StSUOeIN9rzxZTYexdA5BfK/HbOPE9ZZ/ZgyQn+5I
EOfNuXD8iRqsXZCjJ5WDOfJt0qOpGR6LdbaeTG2cjN7OYYiRqXcPjVPDk8RMPCBP
r4pE9rw8rHQbbLKYPtU+BRDs2HC67YIGHE7n8kqHvmwT918pZQwhzZljMy9wr6XV
bx80lJ2CJU7tYGZU7yGE4U0GqSkA9JOQxgyyM5E3P8G4XkVT769+pg1DDcbHcmBA
/ndDfdgBe14qszilueYQqEIuJ5+aj/Hj7Xnz8C2AsowJJ4+I2p/u06wcheeSTzTk
+8AcW8TJvAym8vrkRBNVcRm7MS10jZAGFE8xctygmy4iS2tK9oU360jArBG0nHTX
vHvFOqpK+1wGY3qGY47ySEoj/00qcLe2yyl+n3ufZNcpcgYg4H/B0JqsdVpF94jJ
n2TLAUG7D84qZfSHWxs+Sx1ePd3dYUC5uzwa3Lh7IcvWeRPMcWm4N4ZGmifDdwFd
Ur6tTTTFJG+aeCTRwWXlj68TzKKq5P85o4yV6z2FqPd0eBhVanLzfmknvim8GUna
FxFosE5zofoWNzo3ff3zYByOXp3EYyRTHJp9x/Ur7MW6ZB/uoUZ5ZfBACU0X0k2K
tl5cZkjTEeAy2k4gvJk+5AqwfIjRQ2dsXXEgaXp75NSwzxNwsENPiUpWdHUKh+ST
LuKXYSr/TNuKnqv0UGDooY/Cy3/d+GDkBJmopIHf9t3mqQHNbekSz1GOJkLJbXoG
MeCkIrWsqByG9CKObPMxDH3Su9jHT83dVdafTUcI+yAWlaKd0H7R70vZSmu23XZT
HY6aoHgzT+w0TjJLYp2rD4IQph51w+UaJiE2D6OeD5dVVcPHOUTGdLfWm2ZiwL4z
jEUs/1A7ukcKRhYayYFx0dFx5wtD8P4YYxE0iKeNnGL71GIuiKiGM+k+MqDj5t0q
QpTTVYLeHA/RM+u7u+rgQuugAwX9oG/VUFaomHDeSb4YgMjds+D6a9JWnulLqsP2
AmLEuYQjq57KascsZyOheFUmye2OUAXb4Za0KW5ebhvhIfg+mM/56MgaD6siuCpX
9v346KI/yxK3WxZYVque8IZanUZxiCucycyLnYFTcmtnSsyRyr7Fn7AFZuODqHW6
0f0ey3aWGKV2LZA3kVMUz4SIIMGEbNrl991IcYYom1aikAsS/ipwZgG6HB2cVG/x
kDNYY9Wuqw2mo1l3efso567a9blCe8pYD6SH3EO6leoPX7DOtybIxc5oLbaq4PT4
TPxLGF8SCW1GOCxUbEOc3AlfUyw8TUQniOTare4Q221bKJpLeDmtyNyHl8ibk2hi
OZfPnlmvGG3bzxcZxRlfkbJ5RQPNa75CddQsVr0YT+ZakQ9dHeclfq4/Kw2oDfau
WPQdKz6ouqZyMNArzsgLEmBGB4JDqcwWR+BayeydKQQUU2hd5px67z/OL2C+IMAZ
IwT+BDXCGRqq+95S6xD9ovE5H80UG776t+Yt1EGiB9MPV7Rdl3PNizC6+qXSyOfx
Z/t3eroqgduKn9CsnUfHtE+/oUKRO6sFada9sXmERujNJHHYgmWEVT4QkoUi2KIH
qmjc0C9KE8SOKIuHkrbEPxgHkeFr7gJ226TrMs2EHtRQdtmjkVWpRSb05BY7XRLs
0TAnmcW21kcM6n3tR6n2xDuCrdQPa8lSZ493tFkQy783XJv5le6ynVU5vwRR89Em
F7lVO4F+d3d6121jQ+yWz79fCw6fzgNPTKSSNtkHqwta+1a5cB23Tcm75r0kU/me
p+4xyVse0KHb2/8khDtDmihQqoL3Y5SajDNXzXmhJpRuyCJjayJaTS7KEKCmLQP6
TvS5glAyWXLFnL+FA9jVe358cQpKXbeV91nP0V6mKI0+Yv7bX9ilb6VzqPDI5o/i
iO8o4geSrI9Detu3A+VBLq76fuKC3eWm9C2oyQPXtL1liszH91N7Ag42B0ArKzA3
K0Tgy6D8XGlluutr/WoiwbXj8zm/dBswGYwL76bAQi440vYqMe+N3VHPbvHyBi4w
j1NzPXEJq6JIe4JYB4Xc13VPuoms/RiV81v+39nN5MJIVvez6drk9FD1oOL/RxNU
qxQKRTvPZFuZNtlzYeBvjcw7YLSXb6pY1wo5sy8IkHB8X3nzXmD0IxvZtiuieB+R
Sy/ZzhorEpjm9+yf4X/slb7SL1YQg36VkVapRdMfVsVrLzEbDIA1LbTRzEL26c8q
L7Lj72eUPrM4coCDXJxXwdi23GdCJRZcBaG3PMVoZNQSFuzfbNKxzwg20EPhFqgJ
X8rV8HcPZm9RkDa0lEZdswQkzsPx3ZTHSAJouIUTIPJ4ldW+qC/majl9iyEjPl0y
1quEi1sSSOpY6TpBSSjJqjvKF4EeY6cDJolLriKIEmSwYiUe7D7d08V896v3Numx
hy0O+6OL+uC4aPXZOvmAGZNHOLjm323hOrM7Nsx3ZLdth0RN05F1UXyBprmV0iku
I6DLB3YnJyPX9TRogBhbOkolG/pryUH3/ImCXrf7+5vmS5NBAAmLgixzuxSwIYYe
RIUR9vNCBvZFrgwgsxA8KzdHXub71Z8mitefCjz/E2R0KzwUEFLhX+jlTdoxEdnf
JejdznOPT2MBWMpAEMJjMpKXV0fpUdWTCx5p7NCWAET+OS5shPoQjHKR6kk3pqhE
ah1EYl7LuTKLB7Q1+1SqUvkmWXyE2mPgAI2XAE+YVxcp+6ClMprlufDEruVVNf3S
YjSlhxShFt+8nP5qsL0xcD28oeVeKs3QjDjDUtDFcoGXvgqzgKVx11fXZg+KkR5R
w92GVu0ZqN0cPtghZkSq6p+y1N1ChJdgoXDPkJPmeo6MRRE0GPnPhqnMxdYfGFDs
l0tfOaT37OhWl/h6KEvWNmSJyKgYsNsB0hj89CDVOpXCoW6tAl7STyrAVXqKt/wS
Co3ZO3RByaL5u2y6x0ruQ653gcfUPpKsKw58tZrhybXfDS4HigLAK+aP0l9ohUVI
XqQtAIRD2cdtvFlHkeTX4PvhYoyFhmoAlJaNweqa+WtWjjzVMsW1Ypu1FvX+tbfQ
cAQFEMUfugj6BZU9YTd53j2YYcCE97YymN1PM8ytzYBuCS5PLxK4H+UnDXIl5AHt
woo6WEaFL5xhMa21K6aByLcbFQVePP34OEOiptGpogliNyaoCkEr/etst+z+umt0
rb1K4g0PwPUVDdqHzBRBsGxgXywJT/T/tab3CjGw9AmmvIVFCOkShDtXlrKDLzbs
kSJE0VwR+UhRwIUT3VEICENDJ1duD38yIOeUM30eLYUvTxvd2MkhQYRe7w3gVVde
pYOCtehnbf/EnhlLXTy6fAyelvz5Voh9+5f9xQFOelB1sAn0KRtYsS59yl02sbny
4zJjD9XHp9dcDRmSjhTEzYTj3KEk8QrhckgRO8AwX1XBp86SToqoZxaNOtPWypll
5eeXKaYf+fi4eUnBethPDq+UMk7J/R418CyrEuaI/709BxGgoIAA2AkyYCa0ocqI
+36VmDoZFN4F+yJjZuJJQS1MCTspeZjlMyqTofDjzFtOJVv9exWAJ49XAqPMj1R7
Drg2LVERWb89Zr0CFKfjN/V6KJfPR9rOErOihyAUMC17BMnNR/w59CR+d2MdEvHR
`protect END_PROTECTED
