`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AQP1mT8o+cdBkWQ1JIGz/Gd0lEmkvVJWKgma9eOb/XLTheMsMOUYZ0TEJaziM37Z
Gog/wmBNnEDw/fj9S4h/6La4ysgS09+84z/LQ7IWSIl4EIIDnbf1j8ZPL9+y4XHK
/KeC+MdP4/SipcdJespdVaxEwgXM3iPDkiUvDT8KQE04PPqWSx/yczm1ix3pjc7q
TzoEpk1M7sdhp0rbHfyAdn9WbCw7FmswsS0UHh5K7OIezSCsfFx9Pg8QAUz6qHpM
RddrsdQikB6aKqNaD/hdd6izlFUUjt3bHvGt0kNFG2X3pWxbac/65tbziZK+HdR0
imq3Ke2rAQtJntantrEW7H3LfQklxnam+g9EtJd19S0uZKtgpKZUygGkiebs2ab4
h7jZJ95oChT6Ki0Btpdwfg7Mu2EM/O9Fkjqd4rVYTyByTIKcleYbhXRxWQybtfQ2
hl4wazvjL/aRi9fMA5sImrwmlHIydMPj2Uyn5OUcADMWJc/vQljkWC+6hUJBvdb6
nV4WPNdAGwFJq0IZvBiJGxZaXyHUfHHgYEJblQLyGYqKZ6kzdQID/8XnvSeuBPU3
fIjfJ11qRAiYf41E892pSJYc3lFcNSHJrtDJAY58mFVlqw3xaMqNlApwdw1jVGz/
`protect END_PROTECTED
