`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VOdHu7uba0/g+OiUpPq1aeN4bxgtn7UhCJVAZvGnHDAR/I4WpPeajU0MdRqtU8MQ
NhuMBEkRV4ydeKRtYpi8ftBhwwEWYOyl3bwfLUD+k1lRV/YW7Nm7vGiGvSb5JF/s
WUJOtlvKalZDfxKkpIIrdut4MLW/G+zZk6o4nAcEJUmJxUVbG5oplcJS1HzXcwQM
ZRpRmSclgT9YT1QmnyWgq737G9Fb8kB/+M+k54+aorjGImM0SNZ/pytylznTCtat
25IoLy5bMjJ290DgW5JpmmlIRelNAN/csa9MdCtLDXoU/vuu9/afqYl4DOiUXmg5
jYY0BRkz+ngJysXq0nxr5c9+2kS+dEACJnEExzYSpgTFqjP1bF47JrQNsrav4rUs
plGgeP6iC+/BT4/VCB1Xht1ts4Llo0lbO9pBoAtH7SejVlLivgdXu2u7TjnxHfaC
L6YC3K2jA/U0/i2NU1uPWvPEmYJp5Ly541z6EVd/rKOgfk2H5MZiReqBCq7ri+Ou
IFjI6S4tO/JoE4AXKawKFJViYHUqwival2NcNLY97wdqH4ubko+HKTmKEfc846EY
xvUofM1B3+iiBK4dHsTmUnOBOXyeb34lyYaBkIRlfMgFcj2iqqE/azIapwpZfWmu
ox+trLLlgGdzV8vASav3xkdh7TURb8xYiuWgX4Od9V9I4AVjoKAvzXjfsE89I091
eiLv8l+f0DzZBnUVcewfvDsbRGybm8m9H5GDilRmgoh7QrMjSqHQQdwUUdSE9gWi
Co75/EnS5/ybGuYKZfeNLz0GtAbCyxFvWZie84h4uxBMnq13R2NJT9J7uIiTpeWy
CjMmHrsOMpQHKTw5tjfO7w16rOXay6ijYtOq0bwuSUbm+ZC5eDDVSgEjY3QuXtRP
D5JdmIf0EFmU/LZ9g9xR0L4QZKqvZ5IMc0L/cvqNEBng66lu28lJNNy9rsEaF/oR
+ji6WPMpZx6oGw4r4ueO4JDXhabC2ARMx2p8PO9LC1PuBU55QW1xMTHxWQc2DEqc
ma1hq76+2hUwIQbNwAwkdBsbWoYOYxjEadNiBD3prL3LPehib/8yxpF9//MeAsZz
GJwnjQeTLktHjoDPypLgK2hfbQsIVx+0nnuG9uVmZAvzi6e2+kt8Gf/HkU8jQ7Pn
C8HsLmDu9Nl+dffF9Qzqsy1tZe2Yeo6tDtZ3UCFAH8CGAmTUJN7BDHBEh5HMM9//
mDtWExdo0+ddFlQuWYwLHiSDQm1y4tC2jXXY7bOmyrePyaflubkBqSR2fCBhU98i
B9d2zFgft+l4AZaOjefv+QDAVhACutEe++cJbkHKWksqqBjqSnw2jsT6kDQXxquX
VXIIMTkn0o5/y2xZYVJvvoC/dhXu1sdA3xJzO0nQG7XEKAyEaJ3HFt4myIYBaC9J
6i39ejotgqIQ7uI54PXOqIyW62j/GaIxh1T9tzoJbEJo8HDoKx5otP0E240xMtEq
VH+w3wvnw2p6gsHaU1ggkbwFGN7IDtV9dN13xutc8j4srYRUNHzIbMNKws6APSZ3
oerOspwIUydAET+VmKXk7jYd99iOSogfFj9EZcpf8AxVxNMDxERAywLX0n7qsJka
mHYCkpDIR+NcB4DnERi2gadQPh+uPwrJ2CxNvec/f9Q3hrr0BEA1UPYxyxn/Lmsp
AxMBKbAHZa1NBw8sbPJme5C7QERtuZIf9Zv5w/H91xEuQC99c+/bxlZLpkhdgdq9
nlcairRiLLexVdmZOXRSK9Dumuh+VQcrAXuTk72HjvDFalsEVY9gSGA+abtidYSF
jJ+A6Xkwahk60qhtXnLP+WiNwPOg2daPW/BYvvfDza1XDtbONJ9PFQpfL34Qyu2B
m/HTp1SNdVMx/7hxkZTDtVRg8iKJR2+++W55UTPoYpCB+Pf4UD7fUPfk8zL1XRUc
cTfaaII8fRz/V+aq49dQbIOhV0byjEVEgvSCsCM/AQhjGJY+X2tt9mOChptdHpE0
brV0gG27tbrbeJwsnQ3OL97Srh+Zk6eSzZy0DCvz9VDZU9ja67L85bQjMI2nhrZS
DAOZW2QjZt+SuYvRuBGnUseCy+QMrckxXwYreqvd4adoHzpHwdg+GcW5XZFbBmzf
HYjRiD8/Tjl3a6l2t40OxjyC/TImcqm04w3f+jq9pSLADGtwCjxmoR7BrL5Xq4+k
iI7L5mKBTm1xPvd37WYR4Zn6w2QgeKRcMP8MsfMFMtF4+h0/M1LBLzljEmXY4rl6
3J6iEgW38ZIVzsMduZ8WylF2H6NrUwYR+2CumZeWyL5k285BZLf85ErFqOugJgtt
c0vgSZXlZ2ek0zeDzKcUaHsZpM8RWFC0qFNuaWXA/f0C0tGiNQW86jqV3k3gFDnB
KEekmtzSHnfxIKRqDufcyLKUjPGC4AmTiLw9VNFHHR2QyQHYW9U1XMJcG5r06Isc
maCG4I8zk9+oBBdQTH51wYNJ0Qpl198bOGB1JNFA3mMb4GwKFAjJ5WGBE+jKvAdk
7Es1Ei2UT3UuhYVO7WkbgeeuAyXD8ZdraJHR/9kiAMMzAlHNi495uoebegF8rXhy
awV79tNEOrzMjk1Om/wljpaRtgx7pdpJarQb0v5VrGo5z+5bgYMgjAB7reXp3C1Q
tfM15Q1FVdulbblQaSAaJ81ua8Tem/nXGFkl4p3+vsmk43gFsP9+10h2dtd8viNO
MCcYvSTUhYX73WX4cnU9j3xC9QNIRFDo5zCqb3raLQS9k4wGAYPAdJw+/wzBLNDE
rPWXYITi/l+LSmAK2HThfFR05LKrBAoch2LLQK+qkhEtf0cSXGhZdeV1hnbnRnmj
k1mWaFwtjgtaq0tJOIFi6gEl9pA8llVx3Nt+1NO3bHVCCptGwSdfx5hdqi5jOPOk
Ev7+QM0Fjq/v9K2q2NY04Kym780oUc6dQmMLKUbk0eKpnapAP8RWQ02k5yUNLTbf
moY8K7uhNqqOIxYw3zqG9V4Eqd+b2hg7NIJ5mxlU7j96rhN7CCpHV0Z6sqvAi8gQ
6WZ+seXtisp4Kn2t/sttnC77PVhb0IQr1ecodrau1G5evgZ/1BCsMkxFofdMEtnA
tLqh4e8iq/DEI2qLP2TNkxq4NIQBlS1h5W/F+aCO6shiQMDhusOrXbhZ4J8AbJQW
ZQ9r63JswMV0GKJwHVYhiqzkI8e4Pi8OVGVuVkz6DVObd1NyZjDj2VpFcPz8crTS
q3bnUQU8VZjHHU2wIvCBwuYbogpqOBgYqAYJFziOR4Cldv4gwhgFvBXzgbZKlVox
uRHRod+T/hveY/BybMg3Wg==
`protect END_PROTECTED
