`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6e7Tn9ZmPknaA1S5FBJ96fM5ZQVAhB7OyS+tx6KwL/dl4I7uIKzPEXgXuQ+KYVFP
0M5HpBJ+uLoz0aGZECsqb9vMba4H4UuPAdA66Vh4E0OoXrCcObzpGfEkEpSH3mIE
iWH0a2q5S6BNdEq/yXubX7uP7ChPZ8NAQFvuXcxtH1Hk6nYdwJjkhtNTXxNHi7O7
QUfTQKY/M8d7162r/pXOD0T1mgUTkPRLuOI2diltmMvESrb7PCHsP/wqIjxYLLFH
fekBKJINHeqzw4MbW99aLaQkWUI7zpolEDyKEbnWQky9xaCMxCHvEQHTRahruI13
9t9AdFdDPpDBEBvW8j91lbL6a5NlrKiaHSeOURWouT52nNN2d6zYg7XaPFhCiFod
kv8jYUJjzPNTIigVMFvkuipBlxLKvufYkiT/G/TQdNuYaG+1OVwTiO4npZ7lq5aj
/T7se8bw+y4RT+uJGl3Xzb0hsOqpjBYAZUoumM+bAYOCTQGIHJkcLIL75WnI7rTV
SNRGg6+wv4C0hKE82mMRl8t4lalo2Eg2d1nz0Fa459l9g1O4JJ5MA192t84h+MwT
V0dfXVYFZGsGTbx5U1Mi8GvU7tll0RLMM3bsOPVwad/dgKxVjfv4qEVMrfkP2yAz
5Pa+3D0QVlTit3QTkDUDCPRcEbKCaN2uG7xVSRWSny+f7KXH5sHn4WK3SpNFZgIW
Exhd9e++bdwSDRmVAkuXxvy/UuTEs2O3ZnJQP43mAFPDPCGncQfV9+y9UfJCreEB
6UNXF7MoCkNUmCyhLYAHUDHgCmbLOfZB/0PSd9AgKTEJmBcwvRx24P4rP0EiwPa3
h6IljXwQCZjddkIv1hgzRzEQUK4MBGPuSgnsndidGfx4JyBv4oqR4lBuz0OsxA7o
yxNvl5+sm9rvdKMgdE43tSbgw7EMsmYZ+z/z5CjbTgGGaBurytgLl8+IqO5rLsNf
nST9wM/2k1OjLNOvaYsRq/0L3vyBlkURnaEFrQhxsua5ciGt7vk+MPg2cClKyX6L
ot2U0d7sFMVLUy1+lMDrJVKOmNLX4LNPV2O9u1PzM7t2xsTf64NHu5nOVZZn5JTZ
Pjweh5/UUJ9ErKlHQobihq/TVuZP8NJwf8oJNX/e8FrvDeIUGUMJbNmp5BYMAkbV
gBMCrN2c416RWIhFd4M2i5lTbqSDF3EAeUpy/tKGKbut2fkoIrXaQGhYB+O5dQnz
Ww4I/lR3y4lW8RKGTz8K+ZrijEi4ImerFVKrJQF09mAVfXkKj39EY83iLIUfJCGg
yD21WnJi187oaWEl8ZFq5kcgXXkTOdyLKsRfBmCIIo60lW49iBf9zz/HgpsTjZqg
IloXS9N5itaCk5kwAXOxDVUR0egiYObay0OrDwONLlcX4701kmoIQqaIfW0vlq4U
plh+2m1mBNqIG05jN/Nmsgjg2Jks1AxsgoZlklAGk/9ECgWz7a9D97ZvGKVFVN32
95OjUQ6cQW8KWi5dJ8myNMzKK/ZP/WukdNvClbZC/+l/vWKq9/NZ8cWapvuSKZJ3
dA7j8rHGWiqfzTiynprAAFcPdWs6zwCZ4Josq6AuSyr5HwlkHDsoYADaBjTWHDa9
ecAiZ8FYUsyR8v+IPekaTLoO9S8/iSLWOm4u6CbfwrNAi/B/llgpgIVjSxDsMdAB
Us9G5KNoQ5XomXJvbC51Kw==
`protect END_PROTECTED
