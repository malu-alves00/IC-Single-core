`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
N6rtOgFOaxXJOBgreAouVkYPc1KcSa9oMalvpML3p4gfM3v6ws9AFNH8tgcDrxLu
vZErBkYvIoAzk11SZdi4AUSxybdsBbGqn3x3/2VHAJpP+D/HnyBGLN4tbNhZSmlN
w/UhytwayTtrSeBM2TxqGaJIeo90iXoIZBr14JUQOsFo7xb73XIuolsD044Cd5kq
7u43LvIvmeH2QQrSgL+G6AEMtrvNBiatuwnGbE3peZVYs7tWapyTwPQulW2a/Bit
UpMuSb66FjV0iaZwEJib8uizfh4EWPFUVbqYgmMUpax911M1gi434sZfCAT4f0Tg
pExZ2pxgxjxpAscQTksTUDkde5Xen1lhgTR1JDWziOH9H3bozE+bKDR7EwZobDlJ
BRcZR7pMMcTUx2vNr6tGYLLYl2JUMY2jab+Ab31oGZGNp5obAL2BQmePQ6+eFVQ4
ood7phPa1iVY5qSYqT1zR2FrS9JtwQEbX5biaJuUMSc7PIMRzEWvRJvptDt4TV+U
hUUsxBfmfEuXi5mAapjYoBBKdN1KOQWGkAjHdcogXfRhWhkKFX0JNzry7IT+J0Wh
6NLenOGBGdkRN2r8TaDrnTDDtHNUDdqkA+Hi3Ng6lkU=
`protect END_PROTECTED
