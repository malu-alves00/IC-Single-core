`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IrS/7m9FNUbf+xpQBrBIEoICwhGAqa2Gn9LqEv0Vhs44q8WF9rsOZ17bEGjindOm
D3gEyTKMMIbKeBjexx23mC0oJBgJ0hHY4JTudGpy64sUuoRamYtufon3D/NJGw5v
T7XCCDdMmVNHhGZrN7oaSF92KyOAvYS5NvBIdCEDYZOF+AwtwWEtx4uvcYAYTvp8
f1J65l+RrmmpOMe7dPCLl3F8iTx1+W08PpDyRVOcsB7y22xJuKVH0IXC5jMRY5PF
Lk1qG8ToOnSw007rFH3VhKJcqi4bv1idsEPZ3enEX0W+5OTwPbueoDfafZ9jCmwv
vnJi3S01/0R4nFluCjQWwm7o7p74urCIdUQDIaxXTP6ZC3tkHEgYy/z83dYPSAeZ
`protect END_PROTECTED
