`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5AqMPsgFCzjVVUhoHidIS2fO9Z5GRGbkqBK8D/aqu2DKkRHGCzP2rOKUZSQ9/qPb
VnWZyIeE1hHut7HPgXPTBm+IVnFrHdhbvp6wlrmZXRFiQLjohpjMwyG+q8XRPWYf
ZzkzxdacP0b4rEEYlPHB0o8YUp0nO5PG8uew7wEnc+C8/lbs6Q0dQS0GJuByhd3+
CcfXlKVL3CNQeuaTZAyKRZYXOK+9JmuOTzBzQBTvGVPn3tgb5JlLsdRyO3Xd+hk9
DN6A4Y0Yhi/OE8s++jFkN5U0vjunoEHw2Febu2ViVp0GZydD0E6iGglxwffHMDVm
G6ImXcV9hem9ppKXurNUwD24W1uNREXxYShrFKrjpwlywZaEfluJjZDb8ZG6L8SU
ldMLTSBlqDg4TxRva2tcR1v9AlD8Hg9FDxeKnw1gCB2ROFifpE6EWnDhxj+TOU4I
k3sMM2/4rU5oVbELhYMVM2xReLEveN1h3ODHgOxzNKgv+4Vs62jBXwJveX3f6W7O
zsSsOeG218ySXjdjpbW0sbLQKNBdhHNtgJtZPQNAUhr+ELn/2n7r63bTtzMa0Q9F
/m0ghTZ5x0PnsIYZropdT7z8RtCHE4Fh8wbJwx9hWktt7I4a8KqLPTjIRVn+KPM5
3sIz9rCeX+MZb9Qz6g6tL8XZPj6YM0VA7xbMx+Vh6p3ooQlGFJRXLsXvI/iEbKWg
eGLwpCItekK7b2PMOcftovdB/HLfqPcGSzaYvi5lILexbOkUWNV0whZRcJCWL912
0LoVNXO30RreKYTc9Ozd41hJZgOPMfLomDZFBLy1EEGfVmJMGvdYijZU49VKFGiS
ld57ngB3wPUc95HJw78FKStpZpoyogX27g9hjFIS6uONKEnmXpVGJ61X+w8iURL4
bbZSe5uoVJHEtAtDC1mHk3E35Z9g91XLbuQuvup+g3uTSpM6Vr16E1kT/T/n3q8/
RGQXHTtcNopKTN5dwrU7w8GvGMsYqRx/kGR8wwLYcLXWP4jx46DlEDK87bT7WirH
KKKzsu/WzLv8b6BYG5mOir4anPaiCMuTF9uRFtnmpCAalokefpRDXU53mziQDPLQ
X/qptWs8YmWgRuHxw73tPR7G9pxzb7Am9i9ytVWTPiV26Bg/j9c753bYqWaRZgYg
6WRRKH6yqtTw9EuwcUpM1ufdm+GE0TmjyHOweAPzHeiLh2tYcewYX45/nlWbjfVM
RjNN6dwE2AQW9R9PaQOEG+AkmhnjN/OHzFVdrhI38pmfkP7pNt3U9Qer1WlfjEch
Aphxq0JBXuLaVpQc/WlcvmHg6yh4kyHokJES+IVTveGxbEBknvoUTknOhRAUeOVR
wYr3ooJwXcSRY9tU99GnN9VtUCs8oXhZMSNr2YRJZXsuDv4qNOvTNeiF1yk2Gj1f
VlNI+8Z7k2K91fAyFUeZRvtW/dpkH5Yazdn6QppmwyvfC22tXt8HdX1bBj6zxxEg
2eOdWHST+hxE+rzHVfrx7+PqAXqYQJjz1AI7QPvcCIbPJ41KvotK66qv5ehG4UZN
4Bn7dI5e7VA8mjMgmzePerZR2vPE5orTytXDmyCBh1DDPuB6Av9CVmwt7eLOB6ze
F7D7gawq8IzsVYkoyRrS9J06tO5Ilko6OsOBkqu/DuMGv26efIUi51UnqbTdAn0a
iUt8Nr7ZReFIovi1C7ewNmvJWJt0kdbh0V3MoXLHGLO3mynJT8spCc63c0Xy6N6R
twBBiEszW1f9k2xxStdoCMZ6pavU1R+v5OelJtbOn9YiEKoeMGgnqdskPsSF8GY2
iBa/Msevv4wB5g9U3W9UCA9hyaIwWrHdMiOhLLO0GJsHouTqjuSUqs1yknpsC1N5
cnAU1A5nTozxp7odKJZjfK+ilZrEqDt58Jbuh1h4zATQbIlVS7Q90yCL9/+9D/pT
/iiC6kiW3hFta7uxbBi807S4k1GaYW/yJnqwIe/3Kr4YMZjZhdQ4SJvlaTp0L+/1
hsopse0eVGxN06I1WVDLPELZgiMcqBK4sMXkC6NoBwguWWtoin6cIz9SrAsAL7Cf
kgu6pOoEamPJMkOEDGPfRzDVA/1+tc9F4PJ2v7DeVHCh9p58OHDZ+WUD8rdA5q3f
jtsvIsh1/85j502dpGgVhApEWcoC87KTI+RFIHyFT6emrxIA6C/Tt7DrAOXqJ+JA
AY8dEMyaicXFcapPEnfBjX17PaU/U0G/OctZPoAdJqj90ISNm7uvA1d9sLt9VXOs
sDqIEydnHPpRcN+5gnxaJYIaH+wFGMIpTFXcYjk4J4JBkFhjdZBQu9YWHjC1ipvK
DaABPqVW0ItUh8Q5vIPrFdDz+CESFaLnD+rM2UW/rMw6ZQPpCrvgf1mMOzV5/tGO
odv9wMrPk2X3oOHZOykbjldtyPap+reoVT5O5vdknqNQKbeqAhwt4j9G/lapj2eS
2LMehRhpcCMz+o/fCl882e0rAUGXfBPiowPaj0gGeibKFnLjM7fF408LFTdO5N5p
pbHexOTnqc/vAY+8EJyyA4/2WlMWu665DKwRvgBYtYE9ks8WrIzgkLbRlEg0xSyi
Vt8wm73uBGbBL/X+dhZfwz03VBYbCUSZ3BC2pAOs5XB7trdsjp3goYTnQhu+0hmy
G6rlKL1djY7kE4eWrb/S8wYtjlwz5TLKUFwMsTz8IhcDxBl9J+hisr/5k/1bnlmE
W+ZnZWtI9oshv0nBDhGWG9UaxFr2O2qqOAHkv1g3QfCTfyY2ESqY7TAhs2wtytE7
XMMjWD7XTchBrJrTH6Gx7gN08zjalvgklJuU0sT7jNGkahnoJrT55qXlwkT1IzBX
N/rf5NqtaS9MJCnlz+bloPvqWk/PkCPy1aDVR8Zlkb15LDDoJVMT1SgSc96CcWxJ
GHSLgwOyPp86ZuPmprt3ZD60ILZDwR4jacMZzlJhq0QeuXFqFuv7BBOipqPTErNX
SWqewgHLUw1ri3Em7oFwTy5xwetISAaXnuycA1aKC4QkKY5eAsT239WGDVvT6S+3
ehei2M1jqaGTUPeee87NJR16KvnjW+cpTM0MO7s8vb/zyBNB3KpXvzVhZ/j8BAtv
HJK/jSyfoln/MuzhvCBeqASWoeCz9v/PFwdQbCN9lAe5doc+5+Crd7jg7b4FzR99
Iy8vgs8aFozQcvJBNA3H9KDFOa6kXIYMBNlzsWdGeYHWPa/tBYUsIIZr+MDNAVIT
gdEFmn0JKzINzw1QFS4fkm0hnKailN1F0snoWiCkO9Tuh6U7iGgl52str+JMqTRd
KYJpLcCPS0VYV6JXHPVdTa1zxHStdvb0AcOl6Zl853aGQuY24n0w2qgtOgY5OLs1
4ZPuWt/L3RlQRaNWL7ce7cdVCqBVRbKQBNfsoHSLFXWr0FauHWST3NZGcGFqlYSd
TcebN2E4P2dDB5zY9idscX9a/bAMv/dLCBpWW3lX87CVOgHYt/JcpceVItFhwBEZ
jqJVTSBXeSBmte4ApAEqNbgvr4rsNHHnhUL+3LsHC2mjaMKuHAUqxrgX4q0YoaWw
dyE5KGYo6bZWg34ymmaSPc9HOJnXb7M7DFFOCzO87IyO152+Hi5jyc6rXzMsKj9S
o54x8u0wk3BEeg632Zly7+3Nx/sbwfDKTE5sRrRQ0/wpBwLUOaTtw/1byJZ9LUPz
tIr+jMbf7AMWkfdfPQvHkAk0N/WhrqIcQwBL+nOcBfd/Q8EVQMYy6inhmU44eNBC
ru8MEZTwNlXyiYzHIBDWOXJjZaft4BU+Hz28AfT+kuG9N3SPLX9Ge+eynwuoF3Ra
7yzIkm8WpOYMYSgS6O62/fm7VNCok+n3NaXDrLiIQHMwQQimYSrm1szdObWU4CuA
EmeWhLem32+nTbmUUtNtMdygVSFpY+e5FyZobYz4xkmUdHdXNY5N1MaDIINj4wax
t0FM+DzasR5PSYfef/xyySaiDBZtX5pENc7Tc+ozf5vN/az6oPVbLFWQL2FIt4J3
6Oc3pogPU+mrs/ckYQ67oIkVJemGz6IDBmMYz1Z/871h21tQS2NsXZ+s3HmfKGKS
a+OqN6dK3lTfZlbIrOX/i4N9AFSJ60FQuixOHRUSTOYs0zArWdxFhEHVqs+v1lFs
qwOfZOC9UXCLhjFIwUzliUzXNp8RlGbmUp7l1oeMO9YjDFQKhaM22fbF5+c003Mv
32+tpsdBXXGKzls6Klq9QglG72PlKwtxiDv4CyIP+YAqwF0xWKQwGdwmR/Wol8Yw
WkckoWMQs/g9gDldk/g+XVNM9VkRsPq1UmJiNb+jyyg6hKQIiYtXO3t5dyYP5zTj
xN6OizZjI20Wo8xiA8VJhDe0qAnHWSFqhqHL88t2k0n64Q3GOPjLeoyARiz37Re4
YONl7Td2PUKjErw/x0z1r9VyBYfgNeDf1dEf7nQa7tVnFJpj9+/vwEK1gF5g8kR9
5uZHhvQhwglllc5rCsvP6BxPtlX3B72Zo9UHzOfqw1CmUo8uzvXZQD9lU8T4lMmO
In+dogHH6NAOytN5607jGClgRi45lsvsvYc4EjmCW/zAOAD1EhwMFHlXEp62u/mG
T8JosMl7n7D3TkalicPzx9MIKDeSe56lvRuIMSUmhP1cUOq+vBwQ1YZB5dD1JDOF
htmDgh1mC/SAjMACCTxteW3GuNcsoXU1ygv1vQrBXC0kF3GNguWzIwEHewbABaPG
2mZvk14U7IYMYTuMAjO5MP61+cfcmUb2EYdAFVaUIeiaGHtOQfr2qri8CK5qctkT
XCJIc+1fALzSGJRtDwemgvzeOj5MNUXpgmFAHjrdBfaU85sgaMfSm2nRpeyo7r1u
xui3m19lee902LF2MErWcplfKBRa59UpXX933oAQVaQwSs+8GoOUrW74VydwYvzO
v5pwBBYVrmenn57YuzVCfns0jMhAAuaC/S3M3s9KuRqM7m7Dieue2MK11IgDehjk
uaf0/LymgPC/7ajJG7mhVBQaUoXi5MNtexiOXbAcS/1c7+tTwqKGVofBmaxO3Sfy
H36DIb0zRrh/S+zoTt3ezOZ779aDnB2PicKVb34MObyZPUelFo5pIhhrMhDzYEP0
ozKyCqR/O8SPjkeU17AoSMfe5GQJbNZ5Sr2zyrKNg1Lt5wC9IqzRCBru3tFc3Wad
ajDDbj0H50WrgYUY1D0nAS3WGsO958lCL3MQViShx472coNkAD43C1Sp7ZEthuNk
VZ62iNcWyf5/CoWJPBnD3u1Tk5LLOuZueyKMMwli9BiDTDxrHv4+uCGRbkqWtwwH
3KnrpxOpknaJ9SXzXx/eODDGo5Y4X0jwLsJ+VC23/wbXnqtiwJhWisAyXvBcpIq8
Ynt+5LKcDzU/8ONPYXwsj/EQdnJw5k/hi3ikmhu/BxEUbtMFSqZnnwTakLDw5iAI
QV+Li8XKraw3PlytdLlxKtjoaojK9rqu3R88K5KNQLEjk56ElYBvASEz8Zz/TkfK
LAqRdbD6FbFoGBe4HlYeBzm+jN/2vbPbpmjNOw8DxHB6k0+vn2Stia5qfLlmBFhK
nza/l4vCeehmHJ5rAtKDnD6RHetkNxGTGxv+Vz022fljjh+MtHJdY6vfD/y0+XHf
CCS7ja0YyjvQV/XzxzcS9nK83u0phMD0u0YHTTPgdVBLuL8MCHaxueed0kCytwqk
IqF0DD3h7wAhi/FhojGb/qIc+8KOVyj4UHGnw8d7wyvj3m824ISl2zelkme1TnIb
YC1MsO2Iu+ftWRbYN+C8zYbQBSYgwUOpSHzloQrfRD+mahkolzpFEUufETuNtqOf
edP9P2e5o2aZFOgCUwPVC6PG7wBiGLnR03hyoQsls5LzxIRzrf7VPOaZXcQvQnWa
7UgxR50RLoFG2fPPTvYJKwyd620l9sNE2mVd8hPb5Y10k+VWYhwArLh9cMsVSQr5
P1SqMYalZt8UWBl0ztbp0iaioLsFjv/+jmHrpnTC/c4/jlU9GU9O41Gejafh2+1m
BshtqtaanSitjpB8NZeJEF3G5RY8Lz03JI+R7AlEVs2BZrGAdDuiwhFwXcs/Cf+J
K+O724PMZMvvC/tWBLJP9N62/OqNt5e4OZZw68rKS50BPqIHTvwZXCTClGJb7A75
ucVOkaDCEv7Bvbo+LnqkSYkBpYxTFixLDDRsIBDO7mA0sMx9B3gupkSEdhROQnvr
vg2cnJtUx17jo8RUJky1+3NJ9dhWK4pgAfYcHuUXEfy1znxiqJ4oRynxd2nQb3BW
4CgKRnomvOFKGFx4B+K0sL8WpXlIUxNlOKvuDw0XxwJVbSgwAbFiXYKOgtcBq6p1
Kzjy0D4yOfOnLM4YQYIoFWSTgvuuhIQCtFI8bDyJ0pI/AIxz9OWyXjGZCBFhQKiE
mXi6LvFbPHGjDXxJYRKqOHR91DEEhvFNzihW2Lhd+/1laTiQxymzbWyYOPjpXQlQ
zclsQKPCPowpNXPlM6iGnucmHNjhBEFDfS8K43w5HXfbcqPvTBv2zt2pnlt+Y9jH
oo/VartkCOD3psdW08GZ4ac4mGCYZ2OvSBr6tAf2zfia+kG30PQwxzFyd6+d16Q9
DP9G70bvnnJmNtcFHnUSxForE7q6inOJo/xrYxf9PwPVapTSSCHe7YKg6Vk4njW7
wD0dlrv3TaBtsrol3SHp6c46tYeIQJURH4LsNTrEjMfXCr04rAwHtHPw02f0T+qF
2T8E0PqlQTjnnIzgUGzNiyk99ASF4Zhwadefyr9D5PojUXNhiTyPsVUPa3XIzMiG
cbmrsD2Kt5QMbMkvMkd7niZNECMNwwAqh3LDHH0nf6Z5IpjGfxUvITslQHPmqN1H
tIxHb3+oOtke61lExPfAHSyH5C9p+g+p1/Sy3zw9gWgCnDY7EO+jtjC+w0/nc+8x
jOx9dWH5scYANRjTmuY2f8SB6mOzQpZXsVrcCv8NhAa7z9f1cHz6omI+YtkBtgoF
H6dHAWIRe7nCGSjOjxLsc9no5Cn3ylRjsEZq2CNPYWpjz/wfG8DqRA25OMnLjmjn
LNuLGvAadwKagC7t5q5yjzc8Z+h9Ijt0PEWQ9+00lFepBo840CbBVr4GPPw4p2hS
u7LQzFqy8AkvpypNe9SWDwiFO5g018YlZGpNeCeMXwH8I5dSk292hJFVBpzL68t7
XSudRbzRKR+jnDxlN8GMU5cLwv06mJ9vXNLOQImboug2DDJll8YUEsqmv0jKnbov
MtaYRv2LnWQcjqZClD3qNs46JsJn9/GvF2e7x6QMT8MVH9ThAZ2bFLK1fWXPZ3lT
CpE2J5/pukMAC1YzP1WWl8daPUGLgqAkJrzKqHx0aF7ZSEaXP/N42ik7/UDNhT/W
8VH6e2r4X7gZUpkk6g7rQAWC3oTBm6XUwBwRz1HqFbUcvPE3nAcXPD1E8CDGYELa
989OCs2YA8x8XTCU01edcaIFlPcRzukjl69sGlioVx3yif8tnW4mORLWyTBPg0WD
ZtO4NdlUMwqNJJoiYECC3MLoOeSD2jgL3hWn84Nx9wChXiIk7fXRbepqPfSQlmhN
q2nRWlWfpwe5xA0NmgfZaTjMlmN6UIjkw5I9I93fzJv4d/67h+5Uc8FFpp1Y2Dpm
70MmW9DRJR/k+/vP3GYhX1xjaUgO0Hz+4INTT25mf7IrDgkytxbprYAMGYhkk8/v
S12AHsSstE0Cah23hZQ1iA9qPWuF7+wHUajzZuoSojKUkTk8cl+p/XPM2jZrTzO8
ZzODadGe6QjbYs56hmPbjHz59HbzoDCbFpwVGlKHfAjjfxq7hzqdnSdn1/KaFKdD
MNhCHRGNpWgiUME6NpMTfMaqvugvyht1/OkeuTVC2TXUmohBT/1f6dt+AJ7+JbV3
pglZUfkhfHvZrwaXUZxPEm+WJIqCtDM6oXKviuQDpRXknuD2rxLJJO8DHZE2yrHU
Xr4kOw80cH0rBIj/zkY+KIJbcOQz3mxExDp53790ChOVNOIS4v9pt0t55ZQgC3QD
d4r3k/3VNqFg0/YKdfaOeg9c6IEHcAVYpa0jsLYjuySMxgjMKQJhItsx4LsQJwvV
9kIBmpT0m90QiOSv+mvOsTqD9mii93EPqI4En2jTzXSgL87rm+LnHfGcWEGSrBbV
j0M1qL6QeJXsrUNMY5/Gd3LU7Ey/so0SAYorwTZMoMRmN1aNqTpPVoz7KAx/8Hpe
7HLHMho9lAOTYJhGm/1ueL0H7aufuPLfqmcWPnZQmCrGFopg0L5AEk+B5eujsjYA
D3Kp7yzEwnKEQCpGXJzbdbW8j0Ex8B3YZ/VQuwhFxtNwZWcrNs2EGpkYYgDU0jyO
G8sEISyUeIkpgkq0lsGsN3Q8nFEnLvQ7BqQbLSouC2hI9+TfieOrfAcAPePhebXL
78Kc3cvrHPLux03Td8OTGLCGfeo2z+JDF3nLAd8eIaJ9AtYmQ+vgkjT8o13GJ6cv
jTmzDyWUmn1HhNsIwb3UGPysJS0hcFyb0qQo9VQ3eGz+5nSqbv2022rqMfpZxb/r
SBhXSjAso56asW2ystKk99V08hYovydGrE84KUTyK3Lathg9X3IkSqtLbXHmXCBA
MRmFDaziSZQx+sD8Xv9g/Qk/sJW9RzgdUJx/MEVlIkyB3mn75xnzGmJGR2EFAnsI
FSr2xcDQQ+lby+qine6mHAX5GLHBvHYqPRc9DTRoeebx9o8iIUp5F9Pav9WEM3Wh
p11+LClRYIbF/lscXe+WH5WQdGl4hV5PzooxS5jRiZPUXDsd4MBuAvl4XoyMJLc5
WRen0b+Fz7N6SyFuk3KAlQi6HedHs5MUidh/ThzwCLrNw0WSUwPb69zwcZNLjT62
SBfu8YiOgimBRiOby0SlYYDMJ/znd6HyTIG+TUU9v+49OVGf5ZPO8TUVeTxCujxP
s+T+5TcbfpUj+zeGyto9sdxruq7+5tRQOwj8WwhlYRzhF5QW8tmlvpO/wHvi60x5
Egd+uk0q8uRtGx/MCAnLx/N2/VMNR5njuWiaPpXbFBAN9xHpO9HQE2W023YNOu2N
V+Vn7JGix6nnPB++2yWDlfxlWI/7gfYrq7vBqpISOHvmt8bQjL5H1a6i7gQDZLx2
SSQuO6U7Fyun2RhBVvgeofVus3S4YK7sstPDNbTuqwYqG+p0H5F/Ssz/hTNmGF+G
0ky1gBeUDact2JthawizEBgM+fJc6oybU1Ck2g/FDDYGN+dB7FUdCmjfritOlwVK
VZ/horY80h+onmhbSab/YvLRQbhah85TPf87el4RwMFkZPsRxIu/NrfwLvFIRsGS
mwRyr+JZjkgfFoz/MyWCPvxOHvdhFG8q53CxKHPPM1p0i038EWujpxBfp5lLHWPs
TJFETico0GuG2FtnD3Vc1gzessG2nVQz/325zl0J9XKX9VLv4l/P9pPnvMFlvvfy
lBoaRfD4eUXqVBNwS2DW9HzkHyhTEDbGN3Ah5RNZJ40x0NnCmI/ppaqqf4TUsKZO
xiG2o17G7UFcAe3RFJvkYWadAFJd67XiGq1hgKNuaropa3boZ+ZY8ar7gfc+p+u3
FkU3rhUHECThYnJ4ZdQKww==
`protect END_PROTECTED
