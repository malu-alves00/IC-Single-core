`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EuEcQhL9Bzp4E6O7YaEvPfXOcH523i7P8MT5u0fqXCrQw3AakFij7DG7bjq+pcFr
L11GhxcVy+Ig7OeLrVatDDqouQsmPLVRxxfcWcvmWH9SR4U4qkghsphV1VmAoSe/
aoyJ/oGdevM54+l1kxoVFGy4ZhQD83xvbT4TWMNw6eq0bwRbkS3tCjWcBYw4+six
hdhlWo+OoEhAmbjZTD5C3KUhUwKOUAeRqjCYMJhlhGhmYUDieMWKdZicAMixDgeG
pfR/6Evk9xbhe2VkTathomxl4WbxPAoWskZmeodeUpcLWCao0xy0t8/PKdMiy5+1
HZRcHhqakY77wfsfCbsA6Xsd99USy6CJ1P6XhMF48+PKlT2kK1+XnqoOijQFmxar
`protect END_PROTECTED
