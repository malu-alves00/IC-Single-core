`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ENQKTMtMHzkNbTq8113GDXuk/PNba4UsUWaT2U7JAKDbbQ0ZuKnQIS6Sfnz/eMC+
ED0NUJ/D87qZBsbjOAx4bo5Y65cTGTOQef9dd1raq2Djl5N8YFe49vdCuEBShIZR
I6VKucquZzyL5YfQ2GC/htn7NuTbey3Z4NqnwLSHei63p6X1r2DJrgQjANqQrKXy
O8c8ZdrVPm5jwkBqiCJWzgGWgVCdm/5t3ZfXbJZBp+MijHOdQDCZlK6KCLwktDMa
nQSmL6dfP7ycQ5WQ76MDk94hsJGh8hv+L340rkp+4VN0sud2v2lrkjmE6KIm4WTT
hVXOgA4+oauI6WAayDahC+NWuY6Sma2vXnCT2I43gvNT2TpNxYUhv5MgrelHIym7
7pztVp0cml7CCvmwB3FE4I8AUT66VXBTpbcSUCnL1r1sagRn3jtaPCTCW7PZsbZV
Vd6oueI4Ig9CekhIG2ywtwUZhlc9RkHraDn589ys9TgEhm0bz57h7uY/UqUu1QqB
SoDv9mFeKh7Xdz+V0c3PWQ==
`protect END_PROTECTED
