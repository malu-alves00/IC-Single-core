`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Lv/h39yAjr/RdGd2HRcp8FIimUKYFn1XE5HOLiTdiXg75apSnTP+M9P1itirn6l1
WM+Fyy34Eud+ruyXbcztzwuC2qclXQlOr7vx/GQYuFgbVwz9JLondl3OlaZeT8t/
SviykIHLC9pJpZxHvB2IxJDJZ0fIEptdrAo/QUH974DkFMFMSJV4+8Gkk03oqI9L
M+muIQ7iJ92DaDzLLPUT9K6oLdcSW+Blem1cp92yyyQnvHBSMHChpeVQzRK8hRs7
CviwbyuzI5BJFEXKxJVoG6WBIQTrkcCDLNgfPleiISBOJLGOq0eYd1W0ChJGe0vc
iU981ErcyEjUTDkc+j63YiVx+R/bWLpw/RG/Doo/tEabaxUIZ6nWQcAsAkqWbZZY
GQCfLHdS6jYTkANtEfg6DjKxhpkPPlN9iJX2Lj5FV9VM+2GNTXXhgTOGomMyjLCj
N3hJA4FFeJTNL2BurUdvJQ==
`protect END_PROTECTED
