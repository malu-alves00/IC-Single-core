`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uYKwRXk/y/lit8xJRSz1UxblwyAy9/57ZlisOHhZjE/8fQlUnMHzeKRccYFV6MxM
Vpwoi8g+wzU+zc6yO24LKfvdDZKGchvy2KFsvYi/mJpdSPGRD5LyFsyIIW0ZUsMJ
Xq2KC+WX3QfqQxV4hEvzRUrQAvVB+yu1KV4EZpL8lYm4iWJro10B6bqVNvIOA4U4
RrC5gd35vl0iOno7ct+lqiuZDWeCgecbcTjjV3d4jg2FQr0x/suboLz4MyHrNktG
LkXGEm+lrckV+Xz1B04/yC9b7I5jKDbCa/5oTiPo5T79aUAjoVWsQfd56L+QPtAD
rz552QaW3Orn50UDoErjB6jVyHlmrRBdbltPJIUszSdSWD6DU6vYq5ENi1c5I1a/
rAyYCfCoqWRbnXUpvJwE7Kw+yM2ba2RUdjGY+Y4bAwfVNN3xmlyJrVSUuQV3oFjb
wie5wiwRidLHBaTlLy5fitTHhi+GwwAU2tvwsFIK00+g6aSITN+9tqqsIgDyJio6
oeLSpdUweYpSW12afY8LeNm5MEM/QioMfLvGxyxFM8Ru7fZ8jkL8txAsyXzGcTcX
MSYddOJf+4EXzEmATS6tsgw83P+pKEEqJBukcpdwiteHIWfySs0Opsq2UDqhSE0/
L4ddRIgateiv9hEVt+mkY+4cWaVzA0L0KziHmVbs/Du7ISXqJAqvFY6bPVBBxf+e
RBNEnRaVSBHwOkmq7NV6XRVhKzmdapNDpy2w3j6lRLuXB13T6L+eZ/4XiOWdZrYT
Bp4eOjDcGwHOzN5gdPZzkP9xjb1/sLFagP8WtSHG/5gywv+xPxjoElAQqfbHIqj4
VXvX+LdTsv0DMNhF6rHCMSZfVf36//F4YQ4LV8KtNfThcGsX0xlNKCGTn97S9Eij
/IU2dG8XIRxcaiR9KAcChJwW3+ebLmVr4hMBI+tvFioURS3Hq8SO/AMWs0tBRKiG
A/Wgj+vIOW3+qCEcZS9MQCk3diuYfCVd3kqP5UALDsC6H36CS/cnvNb6/3on/mPp
US4C8nio5I9EFGK/Gg3Z7Fl4RTJX9PIb/742KNhKVUrMFAXYKVaUMdslezB6J5TX
AhZXE5DnBSxbwDuMnUkhkEcchhzsQdJgAWIlLRMPoofERm2WIQrEO73ZRZF5nAM5
cWY3KkJAwwKdhaxgUwg8Hjw/HRXdG0LlIFxkkjlNqtLEpDG792KFEcm48UxVt0Lg
HtrNEAGirgUWYw/RxjZgmg9kwKOuSFIcCkqu63uq1MRpE0alveSaBj8h17lZp/Tn
8MXb9S9jxufcSjeHs732DyeKgjyFz82+OYISWscVA+ODdoQegorotxD305RNPb/6
8DtRiz3H6o8tcwxnh6Z1GsPg5Qs/1513IM2te4xGut7z1yGdbWZNnWdTIcxDnmJb
sUuEl/Ob38I2qIAUdmMZHOe6VAEGjPD9C3JoPmqkVRqJsjKOJYzl3WRgLfCCxD8o
X9syJsLWWL/P9ZStn5Z4cI5mp2+2ZmIERQ9lopgs+uKrS7BQYOV+utv1VhJojsbo
Oe9sXNyOnDf8V39kOuaaeQ==
`protect END_PROTECTED
