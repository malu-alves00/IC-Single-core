`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ct0hmA3nBwHw9zgBEtbGRmxbK9ljEwQeAOJDs8i0sXiUKGtRltZD4+add4AyDe+O
weaMQDLs7Xv/TA3pBgcnKEQH4/Ky31sOmxUVj75Z/JbpXd9gJtyC80/JisxVVH8d
V2hOoMJljqnOg5sgQg9pfPYeIQP4c8kI8WOQzJvyqaONfIYxqY8zCi8IzA68/N8v
+IIx4xvJ7PIcq4ISwmxMsVYxHA0/LPTVwHVS/y+mmPoiJ34Rlq/fFsjj4Mc5Nk6x
TTMsV6RABrt5wbsFpSz9Yv564hH1RNRRzloef4iViCsmFoI+lWcTfmCVn9D3hDxn
L1BUgYB4Q3vClR1k0Yl1x9uCZj92VNg3BCrP3y/FSLg7FuszOMdkP0yxeYxsSBZ+
`protect END_PROTECTED
