`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8I86h3zUiLtBJX+vY/+lur/wc4lHh7gUgxwScC6l1clRboG0YHG+0SY4vmj1CGR2
DUiZmK6vZuHR7YP9mlQK/erZBGFU7O8CZSmQenFiNqRfMovvmNO0ylakxEFv+mcg
mR1TTqR3GVdSBAWnZ5DkGf8eh6P7ARLhX3tNvS6ULiIcmweUcKUVCqNPsE1UokEx
Doe3qB7zUDxtpE6Kw0joSCUSWhYKKh1EdJ4bPsXW9hH1wTyXlQPFE5/n75IYqmns
kMQkFGVljEKO/zNGiOgntC8aY7eexyFWFPlbcpSMN0x5b/iqY57OWzTWSXD5xRXI
tP1LQlZNoUQlA2wLqz55/LklmpUWvArNk5hT9GZmU+A/LqpPRHC0b5FyxJMNcMVj
qSSvlCV3Sjjaems7CrVkhzf8E5mWz4NrMzHxttjfmY0GSiAh/I8NxeUMVBbqIbA3
m3/EkeGeykAyNaZ4rj2yg5S50wJi82B4/m2oQiinYObIqb8ejrPB0svEfXNU2/1n
18FuhU6lojumt4xYHd9lowQfLJnBtyx4hrH8lIT67Y3DhncpP2SSplOi0duF0qg7
ADOuRZHQg81U2ztt8PnPth+pr/7rPK3wx/AJ3FAYdvdp9gaWy+UWoAXJDp4rWEE5
7TqcGslN3w4NK4eQyRlKRFv5sQym1YQoPmn5OMJPrFkpJGKwFwtQKBCHNsOpNnsB
/6EoOx6hawsfoFBWFvumV7SXH6kLnH6rZsnXQarP8LUA7km5q3X2k22zx4mPPw5B
QaxJyrtf9+SHuKJkbDhHHDuUnTSvtur30BsWhjrwoU+Z0T6fHqi0vVcbevqfPajt
EepLP/Y8Fg2WWAo1RaY4TtgkKErND2EJnoNUls9lLfiYX8282g8ThqOF9blBz9zQ
yolATLgYhnBdyC/8rTEYM8Lnimw3NeFKz91FOFWqMi06Qu2FzlIlJeqoz9gRPoU0
17JTV7w0WRVBt5Y8DEmBB6x3Uqe+p4oPlXeSuPNXLs57oF/fW8SNqdKsBoo6OiOe
13hp0yFsiVJLVEyPqcLx7zGVPXt6GxCMvt+/WNDhWHbEmGKlqW38RBeablMSk0Y9
LkDOEQbFy7pfby6rqzFdM+oIDmuo4bszGi66H/bXklOBcYWeS3vj03AfGAlne3yo
EPRZYnv5kLoXrs62grQ/Nv9dp1IecISNENaE2XI3pSe7Unj0MFxagWhx1YKPKEFm
fZ6MeJhwKQKYhofFWYL55yfHQ/AlZZO4J+maKE1NeT1GsZRUvWr5/HYL5ifpB10C
LAIuf7GIw9cTZntneP5QCX8lkbngSfZ0b2744O22AR+N9ggl3uJml32kQHnFrjpE
xyvjQk8wz4MYTWsrtbvU/5udXxW3KrjPs++Hnb+PHWRW1INEVf2sDgVYtv9Ik/h8
KmJ82/icJ2GkDaf428VEL0fs1lxChAWLG6Al0TIqCEq6fKSWr5MhsRkeodHsN7hQ
sEwLlTfr6oI8JwGLaVizWqNWX0YPwTT/T9rxs7bvKzEbkDvYam816+49qyPVtkNY
i4g+bqzUQUbKbEVUSAtDwyDsD+JpxJPaUbgTLpUGRU8QL+pkjjLiBUTU5lEpQMF+
fHEMUtGgCExgpAhzJeO8t94/TPUJ1Nr7ElNteu+COq3GxZlK8AKQ9ezPN1jBYMRP
4p1/2cV05xc3pnxPxQYOAhsXscj4MO33HFnvFbZADss74YAaVUxM3WHIALrRI+qY
T5/JlvPs2D05YltXVkP4HWdr6qOU+Uwqh19RzVAMYsn09Xv4QVnJbqNZyRgVFi2h
AL8aicZR8rZUu419zie5pRg6w3pQ1xLj1kN1P+dQISogObP1I+ROs2imB2ZebCnf
RTL2ETyKj+rNjkGbZgF5GVhVTYS/DAZCLaYzjqt3lTiLPxOMURw+7u1LgjWmOKnR
phedwq0dZfGGvry+l6IR0QTpJMIOAENObUjocJtNcpsVAxvS0Z16JGBPb/dvbT/l
M/dJjcnPB4fTdn5s5D9NlC5duqOmvMCzRrLYaqSW8DCymExoMmt308Gtk18V15dm
cwwR+YB+JG7HYtf5mEuAvubAJWZLqOlShJoXVDAz6c8iys/zBmsArb10SDWkqzZ+
BmAksgUOAHEK5b1SZG1KRb7mChMpPESw1/DnMIXvaj787BA8+2nLNcmdd9nLDXfz
NDweJwqQYqbYgOKjbCDLbtBcXPLSVDrLeS6F84YBHPQdb5sT2gxbp1GixFduI7Av
RMtwZeF4CqdKSLb8+Gl3q7bLEX6iJPcLVRAq7c5AnuV5zhdGWklJ0VIXaTTvUd9k
Xv5dQRM/0As0BRVV4Kn3e2p5ZI0nC6LjjNbZ7fqetIemJuslSlAAbHxL2QNh1Xv2
gxWOTCHGwVTdcK6z0WqT3oK8S6KTcdNhEwanUfTvFKVftWSvF95xliPuqxeRopOE
O0pHCY/o0V02TtqP/DJk/denJJTUX1dPbN4Y9b9NcfejMmGjm3IWbmkJ/BHUgEtK
jOnCdCRs3sV+Uv21wdkyDzaKbmsMHPXhqrtmfvJcw6H5YKb5mSZW9AfJjLIYJAmf
O6nxPZfnGY/Oa3iP1gcfsopvyL/afpXpXRuzCNC0wYd8CAvd15FfMomYySUQNOi/
oUqyLCSrAjwSKEHD2Y5KRfFTIyESWv2AchnVXPJu2paev17Q9t1mAs8EbmW1q0MD
L7mUUHtHWjNKNXY/wVmp26pSmra81lNfcoEbJp76+Ez1ve66Q1sOn6Rz4lUBIOvR
wOQb6TGrBEBDiKSV1QAMZ9cICaRBvXRVeNH8HyLWtsVJT1LlYkVbENfqWfM2K2HT
Uy76xwJbwCEF6mT56noYevXchrEH5ajZY25MNRzJ36Tup2SGBsno/GVm2mS6cHsd
t0naR5omD+xEJ4LX0jSJrF9qTTS4Mqd0pmCcfaGDhyROXm34A3VPgNkTK8I/Nm1Z
mHrM0b6afZHIdG4eUxJyFrXjOB23w0WVAz3bYUqoaPsN9Qa0pL3IPhEPlB26r7Ah
6P4i6NzYYaEZBGoesc6Ft8IkLOXfTSj45Km/0PPqdfYlbFs7v3/sHOciO0y4pK9i
hYpKQ2OkRD/WDAurkhi9ww6V1K5aEuTowDEG3wl6ZzGJEjdtVKpQbYt6PkgJR42/
qrjwNahovbIldGKxahiw9lGyoimA8jwD3/l60bGDXK4x5g4W1HpuL98dlGMm3BUF
VTlxvbT3g/zrWW/O4XZ52ZEmaZ7eXazuEDHp6Q8kiY7bLjeuv1AKj/GTv71n4bsK
OG+vW+cKSohoGLWwNZKq+gNNvfEIQk9saogRNSyxgGc1ZOMQMP8JDKdwEMsniuF7
gVuWzH6/igg0Axwy+fs+QWLqdXY1QSW1hYdvgXJw/ZiSKgD3MjJN2oOSNXzQNlIR
2SOrLEztzWl1AqJ2o5TG4YROmvN5Q/IMjL9/6GzaE03xONezTl2QFZSF5RYiowf+
SKa/4MIS9K0tk1F0feBqW5gilR2+6L/yjbelMFFE8kBGYVmX/oANiuIR8INu1e5o
sTgNJqQQvx/ImSKeX1lC7cwT3LAEN/PWUFe8iSvlOTVq6VhKCh4p6u4aASrhmNfS
BkFSnz4ybCPdkvNeBTu6uQFfg7LoHEpfiaGo1+DjjLZTWdB5ELheSYXhFc6ogMwT
UdPRrdYOpUKZuGSsqvXP40Jh308BJHevBhnZ15kjy9yGIgnzf0JlYfRFwk+N2ZzK
MiZWhY8cqj4jz88Qou8m5N80AV6m4TRDj+3NH4Ikv3K9wC+oJ/sWFIPKUWYPMImo
+TMQ7akLUwbaZ8bp2evKOt1t5RkDPzUMkHiI01EUcyNwdNUZ1W7Uvymx3nVeDPOI
8MMTM3EQR0oNXTTV4/BVX7XEUGhQ9Y8MfpLYxhMKslMY1/CpiqLit8/ULWe8vqdr
MMslNxiFLA+CTz7UlqAOIDOPpTmYP650zfInjphgdXm9Zrsy/qy3sIlpHyNwRv6X
B/lZDAEN+ZpqdS19UySdHpb61ZdGuMrRgA8XXmSgELFZ7Xt4kgkxGJi+padgcHuX
4+1gJwJB86C+RpgZgRpZHP4WyT1EcseS4d/zmjCbu9AmCU6oBmKNx7C3XSG0FDJI
yEZkfk4E8kyDpvEuI/iAik0DS+2R4X5IRgunrInPo6dpJTdQk4vsznr+zMsOyjYN
8HsT/nTSTGRjNTwwgEx9PZRcw3QnpLy0bp//eau8rLcLTWpj78JJqvKKGTtEaAad
wN2NM2G1x0K9tu7Fgzc0+ZKnvaZWSi7uVCg9vE8haYhKPtSpuHgEtz6I5mtYgKNL
`protect END_PROTECTED
