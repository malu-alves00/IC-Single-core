`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Jp8T4O94b3uRy+fHlYtjx+7g0wxgl5JFWWHj803L3+k6CD8xINZhRARPKi6/jI/F
/qHuqPJj+CroFTVtSkSCRFIIGtcFqpDtfdN0hoU0K5sZuRh0JG21MIF81/6qeRBw
zN0Q3m/bQ5PGzMB88BwIb1cPs82tWFCD/v2hKhRvlORxxRqUtawIa0JOKNARDoQY
VFOwR+8zxoyHWBq1JOoCy3K+YPpz2mcUjyRX+xjX9nKe8O6MAi0AMGN7TGNLg9Ne
7zfTM5P6G6yrXl/TS0pkmp0jd8uCfyqFKGF4LhsohvHi5rmc0cUwBD/iOE8cT3Vd
0LfPoo836nejS/MZzHIxysa907yjGCrmTs4AcUgBFRIB2xzVfX0VsQhQZvbAc4GN
pdv+pj1NeHhj14vwALYKzNBuf1gxT47o0i4XjQayi7UOSPYnKmvgFFSvgbsN2NCn
cQIot61g9ZDXcjEjGm7gTEmUQCAO4Jz6s14aQ5sMkT00pnAlKQwssnqHoZyV7zLt
NVz/biAMFjg7be19Q6OTHrRQ+LfpO3Jx6N4jP8xF71HalILFd5oz8JRzy3iARZ38
NAq+hpFVdxcR9HMvOCVSiz3FC3NKXRKjTvAss5cyA0+XREq8lwfPQAJz9Cc+7u+G
v89NzrU/JLoTXS1SYr03CNIE32+uhnT0QAm+3A0q+q50T8I5x/K5byr3qK9+dEYG
UX0W425xjrco07AutYPuMusbvHK85G1pkNxNjsaaqMbSIT1WwaVyFTBXH3EdK3pz
Bs3Un/OiW6ZTJHmp/fG6hadGs05rInlkPmxbLYMOi3VI6BpJcIxuqrrpCEKJAPNa
u/PfeU+zEodXQbGoVeE+KmrlUTN4L6C1MPTeCA8mj1z570zv+6XoInLOUTGhrVYG
ItY2KQHL9f4M1QUiQkklqQ==
`protect END_PROTECTED
