`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WoAYIbX0qmZCPg75iY8jVkHMXikZlmGMn3KQaifixGqFSY64VzmBgyIpUZyYDZ0R
NZYI2pWek9sGUVIkvJXmJlwU+KUAQiLL+ZNGObCnie8DBoZ09sLkaQw5rZCTeUMs
HLy6nO7269Io5LRk1DIC1hnVHxNrAlIBkQB6v2Vkd24eRBwfWJwQvbMnPeVVQ6Ro
Q5ulIaCRQZmnMH3kRl4WezZmeW6gdqeyR2m2cuATuSzXURdJuXsi+HsnCyQUzLtt
3v42wRX1tLcQ7Ho/KDkW2S1KlqLTxnD6RJZORiqJfGYKRun9BtaeMZj3yNevE0FK
Mc6lq4syKX4eok3RuxmxugoY07aqb4+uXViQ0EC8T+Q1uwwZYXuncSNI2YGh+E1q
7bz9GXFp/xyVSmkmFQfz0ciG41okTiWdROxE9HCTx8mXMb1cCgn4qc+cfGxfgg61
z2sVM+oRmzlGQudIGDw4FPY0KFDPt/LRcCZKVBHsH5txojwStGCvN7fcd3sRqW4r
l8hUKZWhqoYbREE8rL4mSigImd03CIlTJDl+yovJojji+E7PFXzKjSLVOnICfCL7
0EUFn0XEaBGGeyDGUC6ITZTnbgFANlWk8awl7gaLeJLQuvIyArYF7QxWgsQ7+xd4
BebltwY8LpjLMS6tISGLLX9lvf7UHkVn9jIROuYYmH18cMYTWTCsYAZ1mPZoZbOC
JArGdyhLHJQVFIbqA73Pqph+qHhNMEX/ctr5jUFY/tOdxLNUJHtxbkJkczot9uCW
fxqpsbaMs/VX2ixSiqJFaZR2zxKdZtYMX3ITuicAEARoyo3cf7yZTUcTwErRTW3i
PLzC/97J0WkP+EUpRXtRtwFIJ82RmxXtmkZk3ii9YPXJApDWDctlVag2MnCu8o6F
zi0/89nSDlNGMKgQ6bABu9H5NSk1sxNqhOcXxvwzPcQ0Y4/NNSOF51S8brK379Yc
1QUGhT5E6Xo6m/vRFXmenOmVNgQaDHoTfvgwiS5U2f2rZmrgiLl3uqjiRtRu9izJ
AF/sHXhRSLRSvZ2RUrIRF2hM1tlC9crYCAG66LM60ZsXvkCaVdXROSXVm7vB8mik
+YREgFZNu8XUh6qQjcERz0W977z2CoAErNwHPS5ctWRLiPWV2opG0YSeL+a6gZxg
KMtvnbu9qlLJfP1ALshy/w==
`protect END_PROTECTED
