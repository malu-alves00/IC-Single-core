`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iRlWqOZ5nVxkNTkaLnMzVaeiXaUyWPcypFrldajWNZWEiG08/4NvH4UmTwDXt5Rz
Uts/IbSJ9/3ZvZr+9EePs/QXGYa3J5hmVcbYS9tbeEjywclJ1gm5nrNtp4meueAO
ZwX3N3cVR2QHoshPn5GEaLRpK+N+wJdyF1uoJ05Vyhm9GbqLdIgQ1spWFDwP/Zse
RalArfuE9YWrpv5C5gyyheELg+Kd1ReEE3fjtSMYFy7qaEJlpAAKNFGoPKzmrFAE
adQMo6PWmSjtBJml6Op5FiLyArkdCV9jTx0Z4zrEbXReUiLSewRfMHXdKyiOjxD8
CSDnuu6XJ/QRMKCP2M67i3ERZqrVVq53Od9SFA18pk0kutVAcZb0jv7OLt7ucZQJ
eWV0+ZzUZ3Idv0MDwmszxH/PmeGNkSu1qLiLrpouY/+1buNs5mdo7K6L2sDzfSxp
StYaM6J6UinmhqTWd26oPwffW9fhe/oV69IaB68NWNhHD/zs2reY7Ocr7csECm3f
9k3MN9ZP/o7RWV6TIBjuOJn1cd82z9pNZpE6X0QDs7A6RgU4MkkxHmUYAVcNKx9M
2chtqRf+612ZJwX3sEEuyOec4dZtjKx/W41Hc5u1tb2uU3Wgabu6YtlC5yltX6Qx
lCd7fUCXQKeb6ckpyyqMPkZNF9ai9L4yWNsnj4GOy6blxgKNTr25Juxe+5eFeb1K
s8SME+TjyiOOd9rrvAyx+R2/Pb53+T5xXPoDzbNU2KeHCMQHy3zOC+kkkCTr+inA
j2shzrshAuuHOyTLSAaOC1/jlTnCt2SaMTKddHqeIFgpxamWUx0jh9Dr+qNzy98e
E1celsX2KACgj1/cAkKZAFBT3JoDOaxkD3H0v1spVnAHx4Io/ae0B+gQIZ/i0Gsb
ZWFRabckavpc3SuioS32MMRZqv91CH/mkqi6rS1MEd8QsmMUBTgdvsNb5hesSFN+
3R8ntvp5ypQGGqIL24gOQA/Spa2XoIoqSMZ6I0QpqBoENHdoGw6MttmXWJL/mT0d
UXyVeZA346/9zIuMa/zjruxjplN952GWcnX1jrhmtvW/F7w/k6g4WfPm2dlD7qeJ
irBucTXgUlCUO4GeL5qyhieOQbB6ApA1XJFBURZt3EyWpnzpAoZitT06v15byevP
aNmWRUmTZDXOJCVQblSj8g3HzhF4fiDyHf9CfYDpmGV27+CXCpW0WnSq091Pv0vD
/gZ78vxm/SADK1+Ypi0eywXJIPi1gYWd1Y47BxOrc5Zlj9HJYCwMc4a4NY39EeFa
1yWdc2vLTBDrjy1DENTpBSbkTz1zOimJ0fhzEb9Uns3ziaWkFo7bcQpGE2TwohiR
SuyRfTFxyuua/q1njSyK9jQEk7sQX6xZpqVhG+1XrDMqwffmOMweDB3biZJwJi9m
2kPgY9l5xWuyIc+UcmmBqycDUO6XkQ0ri+TEhCaLRDr/CXn5myjR4wXvfieRMS5v
`protect END_PROTECTED
