`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yi3P/cQWPC1Gnhraw6iF8RaRExw/NMxbG3EvEpQFtNoSyEhc5/d6942Lg0vTQ1sE
K1MqdylzqB3/qaJSnG3ulX7pB5y8cLJ+xg25PrAeV0NBCkhlO/wI7dsmWWBbW494
l/SO3XZ7BZGkslzaE2AGavgFYGTIp5vCBhW+Ixgk+D1d0FJUIhDtxXhRdeypSGOg
IOdk4JOr4RaU20GCyaO9RtlgOKyURb+QIOQ2cWnBVryoE3nGUiMi+vbIvV0aQg0L
UwivCq2Ll0w0xEkJURDckd8rx0yVJ2gy7lUtzGX7rAv05Vn/pvlyjLNCkTVTLkZ3
rHD2po/q1S8fFfcGZZeQo/jA5wADFiUUS7XUYdRXERlstSOk9Rr+YsZr2SSLv/U5
lz9bLhAeR9L/uo5dzHiJhK9HAffop8CtPx3iDLFahGmcfpci4kvAublhDVo1MpXJ
NX7sHqa0Q6vLy7zuF5dpfRQjY/Vv0Gfg0wL1JupV5iMlFq/wLltmz/uGTEXeqazn
92gGlk/GMLBm+7/N8nWr7oM6VF2Yp87/Na2YQ0HKw9GS4rw6y3qzJ/ozhjEM7t/q
xKyIuAYzgTIuhxCKYr4CruQVuIS1o1an/UBuqV6UclncE8SM5MuRqlAVyjmiKyeg
G+MbfRKkBb8oFki2fGeZIxSdGJ7RV9jy9oTANvPLMdrc+/uZ99bAxunZs92qYAHv
OmpOBGltmTaK4XoN+Y6vf1skKdbT6EK9njBPeAkVTBVZ9eOx4QejLz96JYAHXdZ2
J9WI8PAMKrID4WLyM0hYgW2s6X9/tL/aJq/4DGcJwjO3hycHjme46cxb/4igzWSh
xVzYjJR/sxgREv/wmmUIqyRpIIxer+T4bZWDkHkloYaF847P/Pq9YuiB4jsN7C7U
bUAP4ia/9TcjYLgzUShXBemgvRgsSpA34Yc0t676wd5tv7yE49t2Dyf0w6A11bUi
QtTLQcP1gdtTvv3OZsCIs6pTsJynOHhxt5A3+58kVVY16NrgFvCs2pYi3j+oTTyQ
MyWXJ1RCoe+xMm0Q+2Vq6HJHXZmCFAzvffoAluyvKQ03a9MKT/V1tQM9cWeET7GR
GN10bXUaLrqaGtSWR2+dUS/iDLm4G1f28epsr4fUmZAxDPtTP8oG1Da5a6iIXpRj
AhAyDLKH1nS+P9z3XNaGl9+Q/t5yQVMWO7Taiggli6YclB2YXfg6gqWvPdxvh0DG
3r770J1U9erW74/Bk3Qhgh6/OR6rXCKQAM7BEuRdJMdB2KJHBimW4OeHKUiUItXZ
aL7cJ9uLeg+FL59LkmDrRbI6o3nQfJo8zMLKXUR8scgzQLgfZfWTH92Zjkh++EZo
2iR/PpJYxVybcZGL9U3Q5qi+i7mDm+ILEbfAytP3yXySR/kUUm6n/M3WEPHEUrjB
lPtvwiFJoOfhRo81uHYT7ud71LRIDw+cB0blZw87HFvff6q9VAGDYxpoPSSv6V/p
4VcFHTmFkDGYTOcfsymbABDsljgUVreqcu6ubrOP5ZnyCaLv00NeerBawQwYRMGK
864eDnk/n5vfxisDEN7jFzo52qruWv9y0ku+cPDOLb7o6+P4Kwji872ygm3wC+8T
vzAumzzjjnP72Qo0Dc2k4HLeAQFiaTbjjEkxTgK6je6dUdj/9CSaCuurhB6oSxze
qPfgX9Nxgp5e+MB/oBukga+Qe7Cxx5AxfAVuMfmOLfkJYFHilnM7aCObW+zUZdgS
gXX4kNfUuMQC3/T3MzfyNeJnekpGqlIOsLqCKV+j5aRmLpU2gdoyDWVKQFv6ljjG
oZ2b+HNWwkafunTorLeMVVSx/pV9Ep893EklTQzlZor8ExrBIEVC7xC73SAMlU1R
LSnG4QdAATjGgMFQNucFXFXXcW6r1YA9BJIueMwVUdFu6HTbdN6Ajn7GYn4fXKCv
l9fWZ1n1ZwlBzQgNv6lGv3xOA5hzEpQ95wFZau0wdK0dyNQmli5c/ZsHXzugX8cC
PJGzXWWuOEO1iWj/CF6FmOmcQmieOlUl7sYP/0HYxRcrYu2deU5nVSxkAZnyez8O
JBAro+mfxLm+egA9aq3/IVDUvdWVDI9v+zvORb/9Sexztf04A+2RvIEF9W3oe+Lq
vH3Gk+cOsMeQBYm9EeJRAO8anzhVZx9egBumM1QtBYF8bhisItx46gtcuTiby+VM
Oqg148/BG69OVMxAq5vdqGiCQRCug62Sp/cwzWwBAjxNxcec5L4ZA2P1INTPH7ZQ
XxDMKECtLl6zv3c2v8ue0JoyTO83tvlAZJ8qgDyUm3S87b0TxZzC1pJr/5uU6fYC
1HFpag/nBMX0SrciLXagxetKckGS0sGo3bc7qwHY8EPmVOKtFA9O9N3eBco/h/Q4
njiutsLHiifG4NLKmcHMaIBf34ya33WtEZcBz9s/FkBMYEF6YelTm4UpdwA++A+Y
Zwedd6SwtXrSKFU7ehCFuHycbUd42m40iTot6fe520P7jOQyn+ZRmj6TodjSCSWL
DyloIlRAh0U4HllZ3h2plBumnkh4/Hgzax/LtE/1d5x1UqgVHOrgYWCDfx8pBGnL
BFwC81X3/+mgaOFvG4pnvbKEwrkuWubH8j0yn11NdkNHkUBC57dg3sWPy19+ks4G
64BL5MqHEXsh04ATyb2fi8xKP9oGLOcbTZO0UKJGpx91h9xViktmp+mDjMM3LguB
GOdFNwa3f3WWSYE9jsl2eMlnDO+N9TUWOdt+6hw16WsX0Sv1cXqjw5CMDviGoD0I
woKFq9TqVolnftFOiOIpaW1JaWPMRTYWal7tHek/gtFYziRuVKq+cStUxGvB+2/9
9p6enIKYphJ8afo0MzQHIAQvtwUo2knry8LnXcUTINZUza1doUEZXLjCq5AxId5/
SH2kVlVN5Eb4ocOOK0h5c1j0nSbgHKw1U2TMA8ZaSl6FfOYEnuLBajo/ak79086G
l+UCgMgzA2Pu7fr/o5ZCU5a9y+Fry7XaSAnoVE87cHNvSfrnF4eTdiizXSEIrttf
0+F50qeNXXQk5EX9AjJtYXUk2819HgSowtllOuJyGP/wo0iibm5juXJdDIm5lh/3
mCkhZ48s2WIES58A7Lk7TKy1ACyCME4GdsudfohM3ch2RKEFHG7xt2EOlGwfL3AF
gdUpndgCa7VSFmhGRu/CI0kAiD80R0VLBQ2RTeayORqosvlS8kPVO9K/HAA9MoXO
clY7Hec34xGLUpGbb3utoAVfIwAmy3ZsW1izqhoEvTG4NbVJkyNhIL4GMbnQnZiE
3sTGXaBAhkx9q96P9nTR70gYgUWokvkiSYWzN1cEZM1+W9kUQKTsLbz3YzJA7zx/
bGBcnoOKAwVqkkfpABX7KhZkUzfgVLlTktGkO7CsBj0UuEVp9xP8fq396QuZkVhP
1gzq06OdLagoe9iBWFGbKbTpGhg9+KxY6W2YkR0gDnod9xfLCFDzHbww6rgKBnYC
+0f6ZepAyYL2vSno/x1pWItAzyDWSFvpioDZYJk47Ta84wzoJ3X3jXbNpYjcldDs
xOryyrpAaalPYyIJqEIMsK6+J8A16sn4qdZOoRe5/XP3OL+nk+zY06tIvXMnjruA
nrikL5QnALy0j3j/BydEE70VHr1bdu2N/0vjmKrC80Z7EJ2usw/6hHzida6VXy2g
FiWP+d3B8sIcye/tCx59eaCY/+SFZXgAGNrGdtgmAquG7nUhDmIItbdXZ59V6slz
aO6SzU7ssnWbN/J8Vvboqmy6CUN6rt1R5NdUgRIKSiSYtbfXJLiT+33CE3eHQ/n7
Fz5A3ln9zIDtvTCoXcSN/9P3/CIHJHu0IJSMJNXfdwKR/Gd/52xnHaaRKggZ/y2o
Fz/4SnHNBzLKonsDbDBTYQDWNU7G7CWK7B5PLZ3SvZ6gMDDxmGEqtNOobiDZbhtV
K6VLHDj2OBb95Qj4GfIxUKWkObPhhdf3UXR09BL9NXikP1Y1cf3LlZ5TFaGte2JX
xlexbRPytiOc2/84HgqR38ilvmuOw/K3HP92XSrrU0R+g5W3v2zhEr+r6ugx9UH0
a4/QV9NMEtD75Eh7F60sE99n5XmV91oXLxa/JV+6IZrRPWHp76GFlc5MsllzoHYO
kXrLV8y4lsTnJ24iMSj6Fl3eoPEIh8fMv2L38yOG4/OPvasdFPiO+5/TOjxaW56P
TP1oH+BVx0X29FGOxa2jM4rqwnj5PG7lIgafxk0p2ElrCdF1OmPl5tgEOIaDcGgU
8KxJJo066mayp9zeu0mBxiWxEdeKS3PgywRzKW5TrALl0lGHP8c5Wn3pn76ldJPi
wiU/fETBWtxP+kdR+KV0HsA3mmnYb8VtYvjw8ltEKt/FuwIwt3JsiXq4GiCl4fzW
uKXXPkO2wvqBQ5D3EaZyH7VnkUUQLgh2iKJujFgFzvA=
`protect END_PROTECTED
