`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QbMOtydBcAvQFDFVlnSWqaya1Glf3o+HwlTpGklhCne0MXowC23/5Iiw7eQEn+Nj
VGcc6glHriyPzJq8F+0idY9QgPybJ3BdykH/XI61gWXxz4cxBWKvrIviUz0TEpkF
QyuTWFLzeERF+/YZS7vR9bTq9XXqsEWqEn+jBcKx2NqJKTJwpOiBD8O4ND0LnPlZ
x3zJIV+flHOdzZZ+iz2y7ejamfk/YF+m/+BwNGbSX4kaDSiPJGk+CxyI2q1Zqqup
gBMa0ZUEC/6TNuuWXKfv6NkOo5/XkgF3W+EOjbPJzmwPVenV/QAqVsiYJSAmfV5N
BaKrGYDpFso14auv8jGLaK/tmQb5j0uyOv0u8Nd06/+fB+r1tVeaBaF84fSYCvYZ
MqlPhL6moPt0zE2FjsRRpPbN9x/KJIUkiXArq0UXuoHvTg5AHFBoLoELW7zGTsdQ
4AYhlJCiQ5WDJ9n3d0sQPTzSlnubsNUxo/8rSESVWEvyFY9fB6S4Dj0v8ff9HFK6
NI2HSdhOQa7AuEgJDuTkreamHAhi6xtmZODB/5aDhln7q96Sk02OlVQ8Ks1oxq1t
J0na83gd2RTPLJuNCyfowwereYnCi/vL1D/2lGEG9xOj3/3pi01KkSlZNNBaSW9G
nG/j3CQwWSgZ9mQLWKeSM32LfGc43qdSL94p23GWzNZsa4RetRKbuuQSwza3Xugi
6CvqP7bNYIh8p/wkoOOwzGNwazKbzo6wQqNxVr+WN4m2GgSUJRQcMM8QrxN8Nl8N
lyIDaxRW01rjOVVO0KOCdAr1y2WJNte0GRfMfdP7sW8M2Witb4g1abNwH5+32MgN
20Vw1wW8AYMMpz7N6mV+vo+vTqEbm3XxsqSJOEjPGfUDt91Ir7cT088mcJvMtgFp
oZFsgT7Ajto1iHyAgFP9OOWNl+DPt22tMMxWYWaDI6dqRDQtPPJgQcO7qJO55W/d
S8I1UVJEd2VTqfbnlUmEwvWhBIQ6PZXZ4Fz+kzl3ZG5J1txY2Wj7cwFyZ8QGYqdd
0Zj90MEzERb7hu9RIJktyHAKeBvtHbM+UNxg9J6R63ziAr4cKK5e1HIvJq/FcJ0D
fWG/d0uYv1vZHNN3i5zeGznaOtMGeEAHfsOslJaEVgjVzXJLruZ4NnA/IEYnp47Q
eJrxmlDz3v880sEitt5CfrRRgfrIYHD1r1Gjr6BHbN7vS+v+RENVkrE4rVZvhtuJ
C+e+E1N8hff4PwUUZo1cEZBKRrD3Le/6wAiWA7KimjVywNqP0T4qLEYvbQvb+RL7
JwtsgYRB130AtIvzyrXlZKGAsWl3PNatI0LCFViA6Rl3tkBCtXOSRVQm0KznN5HW
UK5q7jHCmWZ1CFqG3L2+vsnz55+zhLaEldJ4fZfOiMVDGtoYm5CHupPFfdL1e6Mf
vYThfCTjAUVW86JeKB/4Uoddm3SckyYXxEHAQzXyC8a+Oqjp7Wyu4m04UkKVUny/
L8QoChZgOSqe+QceFNsYxsChig2wuSijg6e3PNWAMvok/lZu+UyD5dEm6PO27ncD
Mp3tC9Ms3d5kfRG1FxbZhFWYrRR6W3m8+99oOEoSRjC7Twl/q4rulcZduB69D5Zp
M39JOsf7NzEKIUbR0wFnHmWCgnyjWTFbWP31CPf1UXEoMNzgimhjEB8DqdVHK1d3
k0NSq54lq7Xa/5/DcKZFhPd1pf+oY3iuJPZZgo+5Unp4oC18LlUxE8sD8YJ4eXFr
ytcG38T9b+Amsuy6yzFti9c6SjkTcs+XsOlx0seNW30VP3/UE5B8bCInobsPFIe1
82+nVtqtzjZC3KAUXRSxS2rQH/PjEUqEbXtAAPMI6d+5o81YcDpifH4AV1MhT4O8
HJ4nOkJwAf9pcX2sHOwmfud+VH8Y/pBjEP2/tqAIYRx16saxYT9n27bfqLV5flMn
ImsQLSqEVMLXLgR6brTz/OhCrWyeK9qd7s4Mm9OGI1Vqyq9BMCt4p4/EhDFUG5iz
obUXSjvILL+2YpX3FDHIT7uHBNDVCRsoqIQv7ic3zsubNVdyPWB2UOplpXxi66fz
djiZRjAA0Ga3ZzDG8qOIO5ysLqr3HgYyl/Ov8vWyHpWKvOpWyoQTqOIO27+rXYoR
MJCwDaByBAawazDCAnNKOg1bIE0nsA8mImZCU3oi3r0NglBMfZjvQ1Tmvlo1mrxf
U2xAk///Xxlu32+XxxUrMCVaas672QmsDv2XCc7bzSWamEEyeuU8QZquUUFGpC4g
PqdesH1fdaHZko7F3A5wulbTHmA0T1Ppumpv12tkGlXYVP9a/DKXPND+94MrhQQ9
Lq/Rl1bWQv2Bps83CHIT22sTtbNqOWA2NOokNz+12PrSo2yzIvHvbtzGFl4tHkdK
F2KaPCSU96v97apMilET59VOsT2AfEYMCW5cOzY9CKDwLARfidhd1yCOJUwUSGje
KEKPGYdn8gJH+/kf+aqzmKVRu+BBygb4L4JcKT6LolIBV3grFjKbIuwjsM7X39qZ
Nsv7710nynhl8iixR5F1cOkc6av3MvIMRItQURmbY2/rqUVZUQAthxPmE6n6bARY
jjTJrfxTMQMVRbHza+TrscOH1xiRFzrQbg9X6fxkbGZjWCHDBlUvKCWJj/+XWy/Z
0gsExJ9Qp83yk9IjiVGd4zM5h6Qiv9uXqWIFgNLaa0pKuvWV/A9zZD6bTbXz3xPn
y/V4fVXSZy8RXAIzb9PAorj037O62bGYTu4Ag4HaKw/jwFFSBZfJi7N7YT0ZBRaw
cuhz1h5V2kRFr7LhriHTkY8WGnnx6DKcGkRk6foPFSIeeTYOJZEvvuDN7guoEKIa
5d2bDLwgZn90adZfrujXC95OIvxwV7lMQSVqIUpqlQBYwnkmsMGs6Tk2SRXlDPXU
khJFjSoChb71VGouqmQTk6laL3Cg1YdHtP/l02/CZCyDN6eTYfu65iXtl95ZBjXo
PBThbUdD7yGyzkF1YrG0NkqceWhSqS5c4fYlLZ02NVV7GStn/XkNFqariK2MoD31
+P3c6ck/WExz701Wnk1iPYxYTKBm0RyTYQag79mibAsS8gnsDF1eiAI1F3V6hwr9
RK8XIZW401VgAQIW9Zv7hpWnYdAfhcrFLO9LKPymzI4r9Ag9/eMpWPCSf8ZPxlE0
OlY4uq/f+z4Z43E90DNZYWv8HWcggnEMVGibPG134zZ1FJe0vch8sN8n5y9cCpWP
+DDHLfcavXj0hsij28580LfQmCVUFOFdjmBexCkqq35OqBg83hctHinoExHXovOC
4kRnoLfH4XLF7aixgiUib1ckfEpq3e64Ni2pzDJrTnhpFVdN8TGMGgfveDqlwZ6d
EPOltlRQO7cevv1mwZwEATTSPOs/FGnldsspIH+VQgrbEVUJZbDi70TDshKTf1QX
rXhN4HugaEtFa1Qr1SPgjn9xfUSaaZV9ZzBY1Phua+2sx94iXTIL+nvw8McWNsYo
qNovi2yzD82Y6z8XXf8eeYHaoHhAsWn/JHWj3ExGEoQBMkEsrknfphqqykrI0ffR
uprY0ezc6sJ+kHdwVgkf9GzQblAIpOR9FsLC7oFV54JJnVubzVJ0vcBq2Tud4tl6
eRxtniAotzM7v/u8oFmOaIP/N1AbiNXyrSgUEWtm3xO+zb6bHtzxJV1ki4qu7lvV
7IDANuldVK16JMKeyoiCS8y2DUQHoR9YHg5Nu+Ck3L6SUKW4Egs2Am8oO0oLzB6b
+68LJeHK1a3DF3D0RSEAN3hWpskAaFAL7Kx8ibNYjpyPD2Ive88EUaqmC67Z0T93
ubP8BYcQ6F0cjfC/Ml43Hl6bhkMMTKsEnz9X3kwLvkqOlQlS9mxmDjoT5qV1mJmF
Pbtt8eoF7JvcMWxYCl1RivnEXwhRoWkI7Ob1NFMVwXTY9i31/33wgnEjOpqcIYOS
wcl9fUIv5x/AXhf7+zEVJH8EALAYWBR67QktvAyUVx2RSoDKx8pcIJ5bnKKfFqvd
UTjZE4cr8Tm24xpEGYN63b7A3KeccULSfIl882s71eaAEs0eFI8zaI7NbOifQ0Xr
xLuBrKL7Dc5UcxGz31KBmUutiZttWaunBsSMJpd14GuAz/dzMZlP5MVtldlLnNSb
slJmF0HzpDbAtpvcsOJNMCUayQfOFEraprYW1yM9jgXRnZfXEOM+hFh9lDORScDG
pvC13udBScgMZJgp2+uxoDlw5sXoX8pN7e/Crbr3jROUlS66A457CdjcGQ1l2oNC
NCux2LSSZXNkEVZxZEKXSe4BLxgcpjR8ag0bBBuS5cCokaDQ/M/Op5KCGCNkTE4Y
qYC5DRKZ1TWTKrT/BFDdZwJZEPCr67DyUB4iX/OoVbS5KOCXsCNoKpy47nNhzf5c
II0zHemgvpB7VcV8ZaPyVXX58yEt9/wGMeil75nxn2MQMfF48PZ13hqCPmyiZqsX
ovJdnmzgebXpHggpiWR7DFY5papTyH+XHPYyTxzzQuvjYJvWRbWGMwOKyti0PJbF
y1ZVSByP+K4DlPflWKmldAmihqtQUXW+vCYO4pbGU2gW0x60Wl2rPnk+y+cpMbHy
2earjwzAC2Skje5voyUesc334P1d2IqzzymZU50D6HGlahfV5B1jCi2FZcYnPbYf
7r2EQmunF3wNEptpSg/XjajnAqbY6g5Bd/HXwY3q557Kx/kbMgomPA1L33PtM5Up
TkblfqfyH8zr3bo2oAX3ibRlY9dZX8uDJbnpIlt+ZL7PkX/YKuRk3s3Rml2B4GGi
zP2Xlamt5jzzjvvZ3GhNhcR+ONW/CWEtD62jADbWt9KS/mdDer6023dECrhiPTmp
wfrAmxmfV3t2nbXK9PijHXRdsJtXNrHi0oQRPf8bajRiDTcG3a/kuQOHWtLMj2bM
DimItg3LTSAe9KbDcmnLWnvn3BnKFWmyW5sarvDrdfOKz99se+XzHW3D0dDGXxoH
AXzKvVGWTSdiaQW7rFwcM1loPCHJpK/5+lcPqjMxHhNuGjTE35XWuiFlkCkgLdN/
gCWyob3viZ9hcufmeLbvRDuYTd0Zu6lkiMCMkBL9FzBTqNjYFPhJW2BS5UFSRZuX
Jacfz3FumkgeeQ2jALZfM1ltYnEynO70WTNYE9gSUSaBpQtVySsMNjtMl2j6Klj4
mgji3NKwXMZCop4uaZYrTVGkUX4piaFs1AbE53+0NlRpEnVvSapuRQl+woyVn5l+
CQEOxjTjY61pszf1Ts4of93LzeEP8bjgso4H+aMotOZXqREMajTygzVCOCVs0FAP
hnDU9NF3NJDazDLdKxk5y53LmhV8mzRkmerJAuk/kKuI/gSPcxFFNtRY6/gVNYqC
Y9youZcyBNnv2isgwG4KSkEnlhUOi39cMa0+LKp0IQtNyX7fULtmmQpjanzJfgrP
U3VaqJISlpYFY+0BmWuDnseBu7ZyNiwCBA9/pTv7tJ1ujSn3CoWehogdvy7fa4Dj
IoEDq9yYd/z8qSNgB7ak6Jd3gXz7ztdTSm/8Ve5175XZmCZ1NiN6wXzqxVFWdy5y
vDc+LeheDLUl4VCDShsoe2fh/ONrUNtUuExWlagDRxxqhkyQcy4Hh43DyCrh9V4R
N3oVj/5P597A5KXrPB2GzfGJU9np3WJNWiuCjdYBO4/ELDVawU4BAHNjarHZiQBR
JQY1MLLUSKwa1J9iNQZP6vGhMwYtw0PiCT55KpEBDu14YEplOcQS1gLzGJxgR2Tu
ei3HgVz2PmeXhpWLpKDpWV+E7DeW58cCBYgja2JiJOkBlPkRjSMTLggSQLQO/DEB
H/hyoEhkQpypm9N0jg7bqYU0FU3HK2TUM0GQMTpmJmMrTKR7/mQCDlh+BEPDP+Hy
Y56jlN3sf1snOUHisDFGsNbIzVYgQ3lsZh7vHcbReuiHssd0OOESxT46cjEoAimZ
egdpzl3/j+cDUZ4Rf3AL62mbvbooy9uCw52103EMntbx9SVePCiIpydfxUmviJXH
TiPR7A7BwiiIXTl5lSDLBT8QvuGUF8wVmYlcirM2Z2XwTIsNqIV3coHjM/vOk4UG
qA4ocTwB1s/qG9Dkn/cE9TpZKrbpyUvuw7zq9+glyRb4sUxWo9QC5sT7emb2skMy
iLg+gJ9XbN/7ZgwgnzImZLbdOONlJg6MdI7wbdXpscjEhVzYCiFhoiGRVTm5zXJW
HtPc3bbFm8ieJaIFk56zWYyWsKp0r+JS3kNGxsaF6U8iOkW41bkZCZckJ1mabynA
7PK83NrjkufJLx6q4en9Fmk21l3x3MjpCgHoylh+e1NZrZSDaeUcW88D4nGGh/qk
sCVVXfWdOAlmsmEXecBsWbBaOlJ5S/aul0k1z03hdcOC6BnEuFZGRGY8IKl/IRm6
STiUjDOP1chAhudKT7Lj9tv9TCf2o3h10gzsDsiOY1e5Q/6P74pX0xk4BQCU9OiA
lGq3LYkISiRuxs/vje4mhoH5q7Dp6+tEl0mXKEYbZYk3dJzugV07X1++C3/NuHnv
IzOmb9DiXTOo19/mTyWSY7LdwFXIoD5/9l6nONk6tcHgcxFeTR78t3IAW357CamM
tgaJOo6yKcQg6l9YsDSpgpFZ/wlA1UBe8R4YeJSQqsri+cmc/LkEIaTEA4upYSO3
jR5gptVrqCN8rIEIY8p/A5i+9rQOErGb9LV73rmBCrPep4c03yp2QDwHC1t2zeox
ShhAj0K4O3kL4KzzdExQ85r0HArQ9I6UNu97yWw+7yUEspSB0wv9Ux7mUdJ3CNML
Av25HBWFBHVXr+xHcABe2sIAtk1e+yG9D/5YrOaJ/F6vFHtj30UDNbQq/ZE3kSR0
MTTihHxPqvqSqTFfHgzG2QB9dEFQ9KdqeKhzXGlyGJD6+JJ7QlAOZfiCeeRpFtpE
pOpVs+FbmlYpC7VQLudCFLEnyPNzJiJ/25AvulIKjI4fq3pMVJCpzcEEgvusRGyo
KmpwSeJS4ErtlcJ+D/Dh86r/3DzbGKP+/aGNWwLij7nPjxJESNtSAMJcLV2aOXrc
YudiL58IEv0Uv00k6r8Scg9VyMNjUggCQ9xjTpcMOjjm0gXpHKld89Ju32heNTjz
Xo70cipEPj5RycDhUlReKCYOn/mbjVK/+Dy7m2hUpL9qU/i26nc+R9Ug5rsdR+7L
Za4Paj27z1VVagT1903ffJ5bnMgxLzZ0anNKS0CBN1UNlHGHuYtsd6pSce+y2CHN
Jol7xQCphttsVJI5LapAkeqffAEUwI3wxTtc3y0e9A3DZJwcm6qQrMrA5Oh72NXc
1kGeufs99Lm0KY5I8jf0iOEORfaQ7ZC2wPy33Pgwa0zfdOMTHl9t756y3+ALMcQO
gVaObjsoSfwcC6ZIEHTG0uDR5VY+zjUEbduL0FitoIDvizsSDWPMy3UCBFCiQd5H
hHek7JJM5+b/+VuMNVIv9b7tWkYEj+yzeHu5LPtn1zxMmS8SfKDdPtbGxPFAvkIC
KyuS6sWwotd7PSjQyBZTiolGQ5RRCs3PyXA55IqOv42vPiOOmNXIZyTbhiGPxlOJ
qK4bjIr7rCKoRJ620DZP0ILDUxl7Xb0c/zXgcQL8yDJdxRSLDDpsoZK8NRPPgbMo
g8f4Kc5mg0Px2BMKeuR7PUUdX6835ZgwYIzIt+6dqUWMUIbRR54rjj4FFG+GHN4H
NqiOCaoz8TLGpb8VhpHlWebwnRdS0sgGVTmEU7Zb5Jj/N7r4iM7NmIoOxqytCE3v
ZGFmVhREXjYWBq2bzIdqY+3gPqxNS83My2kbxP6KjcNkXSgRs7dMkh7njjESmX6o
U3Vrai5lNIP3806xHHTolA==
`protect END_PROTECTED
