`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TrRfe0lXoQeXVysiaf8YkLI5H/mTame23v1ezrk81o8lJIsaJkrhuzNmRI2QjUy+
vlO0DOA7S8aE/5nES+Vvfz3I8UXMb17VW9xkpcBO6J1W4e4vxG/l1cTm7IsBSOKV
e5qVLx5eZV3H7fZKWfqDLikODvm5aRUCvQh5eGaHLxyfo3LmjnUFY35MOPk9ivR7
H1JbsKczHcKLOfJk6JQpWr1uQm5gLEKedLSVxYNovp/wJv9yPRJhXsAwvfVm0ub8
6T94AEdcA9grwtzPTZzojEYYwY8TLjoypRBvnAMBc56EtKE6OCVLLH+ZkV/4Qg/8
6+ml/A59lzrAB/mEiyUSUqI/v+hzFUZMxNiNpvkbU99w/yITZHQ3yN5UAoNyTPlM
tZyoE//DpEgIn8owN0KVrAnARu409Xjryj6W3oIaQU3RotnCr0jjJjJKGEvf4Z5w
KbIxr66YFX7CYnPZrugDF/rftC2rtmyfzmOlU9B+hGhCOz2GHEdM5eYd3uMCiRy0
QqlY1t876in/SlSUnyJHhwTh7PuVYPGaVzeZK00smeO1jBeuEod79fourV4AjZy+
ZuaBfhUlDse6A1A7eqb10MUd4bI1WmzbzcYIBPGvVyi0Y1EOprLmJEAzo9tyJQz4
krMu4x3AFw9AuXQVQPcg3/8ELmRT8zyBLclyqVB5XT+yMh32E/3iJ4pDdp0zH4vL
M0QRD4aTgiWLZa8W298b89xgVXoEIIbRABnj7r3UTanYdVsVZNzGkPv/RChp8Ohs
NBCHT1OTlh2tZJbDS15Dm9QrmYvld+8qJJJj0ua9SKoZNfzCBBEzYqA34AcfqG0w
8OO4iYgg5AB0daCIajK6th5ixNoAYE1XIwLUZNPGw4ZDjwC2jTzL82H2s9Gy/4k1
JuJub4kNQtL8FPbsQTmuJye7hfiroOF9oMnqjEXMzsUxuxWj2E5qv2RTjbuowjPb
2rQGiDLjeSaAwMVpsVc3073Ia+PTQPLhZ0pONElhns/wDvSZgSfqKYg4JHAZvrnb
U97zNLZaOxtAbFNmaTU+u/zjdjAnq3oFAs2+fXlwGcq5a9lUEN2p7N0+obil0E8G
PUY7h8qUuJduhZbNtbFsAEQmCWZpwzb9iKMwUMeT7Xcl7RSmlumMUV+YJKb08dfW
0D0zIA5Ob11Z+nNtxThwhBpZsNlBtIJ9Ewz1hMH2tn7sLoGnt1nS21f4ZsKj1fnn
73LaGL/qvgQCbs9SOPqmewoyI/L9AJ0zmohAFQjdUsz+vRmeOi7xdwvOhtA5OugS
XXhI2I8ld+uBiD+FB6i/aPpCtwkm7QDTWsUZaLjyh6DrqBdN/Q5c81nl87m6szzy
LVa6hM/evtSL1ABWmYowBo0Sykn156CjWbU4H50XJUxHJDdFSK976z2T97cV1HOl
X3l4mvcrRdw8usYUSM8WBWulUvMZLQCH6uv0TRZNbS7qpVemrGnmFk/tJIi/rLxp
k/TH57nKu+JlEu1CUMF2LUIVeA89/RqbC3cSnGKzRurckxSIruXO9zscUBDuCnk1
iPkoOW7c85hjf1sCPNca03ttlN2re3ohfxsX1pWBKpHIAx4DTM2qYKSYSIDCLBQX
MYbGEkVrdILMT2F2Dpe66A+iOyozSCaEFlr94h976OXnxqssJMG2FMdpuPk4h8E9
PovNh9oxpaSr2p01x6ws9oHQAUTXrDJnjDs77w1AbKMRifdx4rZwbVGpS1CWyw+F
F8gui2DPvz0FcBiNTC9hUcPX20ZLWTU7wIkUsUTwohui+0YSDL8coV9iPbvgs2F7
kVZUXhqGoOoqTrbt+tToxvledAIto/bxmKzvWFbVMBnhV71GuJCDacUI8uBuT4RL
7oNX0ZyYLWFRk+e13oDMi8G3wpq5NweWsaRCHbx/6606cX4dKarMIOfOpNMBjnGN
7mbbbJMKh/FkLfnd21p/zyIZXyZJkFwabYQ62f4N33vVvaLg3/VCd7QvOR8QdOi/
QrGKa6jbYJfHSx+lSgRRhIeg3sE/IShm9INAxWTeGZc6sPZtqfbRI8LOh/4JSids
f8NsmjD979ftzBsIsNpha9MemOEy2I9GiigauHF4KjLoHo2miXJBX43rmx4LMrV9
pmVBfBwW+kha1DPUtgwPck3ZGq9VtjRhGet4aM8aWmHqS8a2K4ecBBsnfOL68lmx
0bO0gaylJ1ibctmIiyEZCB5wxapJ2C1sZy8gV8te94pnOUgOvOIIyj9BGOWnBGSL
Ixwup2MnBeHj1yYLG49WoPAtGAQsjiV1Z7RDMbnV24/zF0usMnVtPT9EGG6w1AfD
K8o4NPPDoblWg2VaLHJaVu1neYM5odYY/0VXEtq6xZ+aF60tnOnShG8Qn3/b55Yg
3RYA9i7FAsuPqvs8EyDSuaHVXn0iVAnsq+Ev6ke0bvH7nWAPmbTscp40bSrf6lGy
IqPXr6/HxDl/kOZC98RWBeCNgelBWVqRJQc/gGmCFc9X8rPwZe4du0bJpkcwK9We
heV1dNHl2Nt1aVA+PTSwkhVUhs6amwcETz8yfkx/SKs=
`protect END_PROTECTED
