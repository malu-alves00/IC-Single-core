`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TQptlU5uz/UQkfRv8c8+JCEubpKMX6mWa79XF5vE4cf217jVS8ybORy070A5bGB0
P1E/V7zxMqV9H65FzgE0cK3/6gCs3DXkEfIK24a/28QED5vEfAY5rEjnMjnyb+jo
4T/qCkbA05UiKCOTcrAjyhuyv0UW6lzUJ/FqnfGl0X7d0LF4243wqsgpR/d3T4nT
zbldD4bd4SlQszqozbVaF3lYIAJXNMre2hbwDraik2rCiD5OLyjHjlu9GzoJof3/
YHvjavLfcYN8JyoH6nq7t70SxWs5OsVaRk/DpW9Z0Z7ng/ug1funB6JnLr+7pC5+
X2+aA+mT9M7RkVNJU8vkXgMrUaJmmWW6WxEp6ssMx5K7/wNJgQhHMi48vFgwRXWq
kyumcvStNq9MytM7eGcXYDZEU3p+taRSJ+yxpGsix4ml4PwviTJ72LnzFMbKiWN8
eAo1b4ZxtXI7hCBM7SbFfeDAVeVyh27Eaomyu6Pn13gmHEfzk5ms9M5O1IexjbcQ
xFOWEsiUWWKeH6YJ+13rPmbSSLAanooKf/Uso8nOu3wIfzhz0DDY4LDYhFryFwu+
AxdvEWE5G9Baj3okxCmwXAnUFRF6Temx2N9EImu8PmO5IO/RBAh3ASrOOf+4z6St
5bsdfA8rzWGXGcwQUAs1s1eTfBbvgLF+Ds7G0iClz7JiMimVbFk0JwHbeuubpjds
3osv2Ci/6CXBKLPVG99KBmvJH/ZxVJmVNPvT2qaU67P/wn4+GbipVVSlLhwKVlIF
QvDyjqq1TRMIPeH1BluRRgN5vyTZweKQxxwWs5fDG7vc7tEOd+LEvkwRjG/+4OOA
T/IikiPLK5V/Bu5a8xiGtaaIAZfEBuRkFDtGNG7xMv0uuNk3l0qfpp2MnqGA4VAC
JjypE2tV/ha4MqWOWVUMLCO3gKxQE2+YXw7P0sZK14Jw2Rh7zpR60dr1C7FJcYC8
OG8Gd+NikjWr7g9tOR0JOpElW4lCQyTFyG40MZczf1Vw4xoGRCMmcwYqZwMHuCl3
Z66DSHtzz/tBwe3+pgX5bC2TSVyGYmMwuFZQwdIYSIz92et5S8Khdke+fmEshimx
8VtxAFVbqi3HlmTPvx6X9dqboA0eDjxpAHndUzSxfKemeVu3jSjyDch0c69J12Q9
YJELbZHDcFH60VSrUatrUDYHMNYGHz4EqSq8wyfsM/t1X38cQ5KBfI5K+uM6Ksmd
68KmADXJsmQ+v80dwCWHJFFHWRNsb4C6iLkgdKNXeBx4hFh1DuTmQN6SzYwroA0g
2AH6xKGoCYZGMUZx+erNxxurbEHZRcpn44mvBKnHUbdO3/a8Zz+LRD1MDJbo0HS0
yomWzMGNYxwfnY/IBQOda+iPoAZr0PGMIrtj25k3JCnEKOk/FhbWFkJfbqDrPNtK
kYI4C7kGOaFnJQJ1DV8wl0EvHvjLUorFeGqwmn70FhMIfbihNwZDoSQ15+YA4vnN
QmIG/q+rCBusPbt3TUfEY9YdfTBr45hSahOWC26D/7TFIPUd6Z/P9/t32M44p/xB
opJn8yo3r8bCD3l9QtUNjRxrUGnzuly8Ioo/aD/isKbQe3T1vKHxshCCdPNDr+TC
L/EjcYbVMTPd0G/CDnd4iNWZH92XS5tC44tsxyaDWhuFVNAVxUtZJSZoIOx9FMee
8bC65Owj/Jn14Y5v3vdFIggisW4/yUXEwo5MySrSeP98ly3PQQxrA9wmKQz2CC0Q
tGwkMS1gWHe7fVhqBpr5cDqmXOcPKInT+VPzB2ayHTxcq7PU91gh53W+98RuhXHM
nqea4hYqW9cIvdoU44a6gywvg2cKL0Vh7D4AO+OjaVc9L5FFhCnexFw+5VW7xGRU
ajc4wK8A1dpk9uUzc6Y6oQglkhf8noPfJipfKnArGOt8QIeMrPB0cRW3nUCMrifd
3Bg2b0y8NaTb5tfx40C1WZxzzIR9UlJ9b2CvOcaeKOf3lqeqgcXXKmD978g+yhM/
8VbhIY7+5PA/wrL2ga++oZql1UqD0Otu1pGYYt5zs7gwIrBiTUCnFrKoeEJOwgUa
qET8SGouH3PQXBkyfLAW4dVFj7MoqM/R/Od+c8J8sWwBFmLKjaZzurgrA2ZXAtAo
i0VhdH+nQrNrTr1rUUqamp9xJ5N/lmZlfq+EHjQP5m90SYfDXNr+M1tMOArdbcUb
0xHJlZHMklDTu/YcZ4ZMyrPhj6+9RSXQ48SzZ/omr455sel43NfaY6IW/WLokKdG
SqhAzMsf2soWXLREOhbP6EvZz5bd+PxoaEyO/TMxhqs93Jbk261DI2CaUqJmeD2z
qyt8IIuqoX11rSYuuCrvsQLt/3F5ff6jBK0CffTIZCsNMM1DU8Md7iUBQAVMg+3Z
XGfUxcXs+axIXe0GHppkHael0gl65LIGlnkzdurs3fi8EdHtvQcZ1aTE8Ft4k4A+
wfwsWDS6WHEKqTLSTkN2wylG2Zge3pNs+x1gljUbP3cb6NDNNprASZ4qwGcW/w9M
VZmCdPsuyAMbMGg9CrQ13/8v0pi0GVC2L7DxCPqqxpHrmZ2lTP1CPlo6JFgJUhyS
bQUKvyidDoKT1kCW+/sQEVIZ39BDoRLWaCdmF9h1y3LlZ6iuRW/q7KtQXmN21spW
/bxR7xeBlpfe4o3MSVoI7s6HtIme8HmpDpouCDLqOpGKsHVgxGD70y1zg1hfzr8v
s79Z9j8+2b2wMX3zszehHAVyHu0nPMQ0+xKOlt0o7WO557nfecC/ucCoa8nl3rz4
oGl6/3KPAOsf3KkXQcjrseIYtUH/UO5DIIbOJf8TKkDtYrSWrjBlZn/SC5obm7C3
KJiMcujaqufTYrn8L+zqjTZ4w5LV1rDJSDsALTCaFMXQIHtbZ6wpk4xbPtWv4+jE
Pzji3bddiyvFjQOUa2V5tEypskXFGxLKDWDQCUc1MVk95LC3+SVz7iWVTWa5dedU
3BDfhFeKIfS5JnEGG4+zE+TeOlXEfsILBMLm0KjzD4o7tRzvQw/JCfI3OC+kfYi/
K+CF5zfThCdy0W6jLEqa1bEZw+QVgo+enjUa6fY/PLK6CtgS5/YUSX0oyxXTST6l
EzxIhT2qxYhkS5kgxbmLGxhqQj0yE+HYQwrMK2QrDlzy2Hey7yB6smwjLyulLAqz
7IvlXkyTCJsP91udE+/wj1bemrxz35qidq0j2AUYOIbUC1dvRSl2knND572bPeTT
I2W2wfBgUZSV5yo9aEpftwbRbulnAqDMnLxMcS5XXy6eWdYhJxK38LKeXmG8sTl7
P0CK5+qEuzRGI1Z6AWuYfE7B8yPQWEd6zB1eYD8RbtreRA2MV4NhA6qLf6yaAaXt
MvkRiQFmw7n6CZGLbB2qVFcqtdFE3Gz03cxVN1shhh4m+OUSg7ys6RwgLa2OexZp
uiFTUhaFN67rXWkkr3bHd/Y1dtXVCZAxp18RS5+6PviC+mGfQtRx4JrXLjngaOwr
7xeTyJHf2/+2BUNxb5AVl/44LpHFNzNb9K2G6mkG1fOeGEuclGLN9Ix9Q65PJ5qT
jzeahMI+pc7QqaMDZHCW6NOdyeGF5oaNcjT3vlAlb2xi+48+zwC+jv2T/G4RTCQd
t+8I4amlR891c/YsBUpyYMqf2slAHIiVn+MEYRlc68jbylrUoj8ZVlLRh6naSdWh
cxIorlNSsXfoPA00ZY7nlcbkXkHeBvpapSfF3jdE4uCvGyHSJL34EBJ6PBkdyuQs
oOXnAhGrobPO4XqntNVcmdtdFf+oFomtFbS4JO/nsPDnKWWQ6XornYTsRMRgQ0F3
QnBh6cx0FTacE3tN5bnEAiMUgpIFmMF5EKDcYhBx3seUpujMd0h3P8EiGXoPSvbr
U87ODFMH/R+4cv4981EQxK9ipMwNEzEMcWAol2xF+vcufn1dHAJJSmLckbdbMCSd
FQQw/FTdNKKfs9tnTxzhmXy1sPEkzYX8mytuc3eLyhzZLSdNZz/tK1GRvAH1PCjf
lPFGGFdkjHCf60slgH7vRzRQleLEq+gAlC0T0II8a592by1ImMZ7Cswj6oQwnR2w
76M38h67tv6oHuyIqQ9yTDNXZ14VHvlIkfeE34YyMkanoZVC83addV+ej+I6qmTV
tZwDKyJKnwndu94hZk/ZBifLgAoAYJFce2MKEHBoCWlkfc9Hm/fUFen85TEArbNs
ba3Q5H44iJqJvmEpS4zzv6HuIBkC3ezbgF7NS+qt52goeZiu1G78gx2fej9cGm5p
BDMrvKAsWPJhsgp8nqhxMXh83emZib07Wyr7zQ6Avk9aYftIuh5tBvRygXCzzoAf
4fBuNxHnp9UYPgRBS7Xk9wlWa1SVi6NgzUDAAyuV+egu6sZ5tlQnVvlZlwU2LjAO
VgZcxzhyYOQ2pjoaL/Upxb4Hrzk3GWescBy9t5fAlQXYA+t9Cb4877DE6xm8TSxo
EjFfbfacuq63cQn2UqN7DzZReYOLGxevxU0jhs+1Yt2ttnE/beWfFulGoGZ0qQ6H
S9VRNUw1fAJtyvnm7m37rO9kdicnbQhsyHRTQLlb3iuKEDEb1HL0XGbid4AJYwdD
XizWtbkVTmP6IxQCjPwKKHH+/3H6HclLByZrnTkOISx9ICxPxN6ymJ1W+NmwEh4o
1Dch1tH+9X+cFi07Fdp7eY46UaKubqQvZ7B6HtEceRKubyj/7bmu6XtNwrn4Plcm
wvHQrsjTKqq5B4AKZU3J12hYE4B00zTbUjttuDlIsN6cWl9OY/XkeiVQqRUWSEke
tfcwtd7nkFVTJN7gxT7KKTwVUJ+KnfmCel8O0nUDcvANxgN85kWCdDDd3ZBvMn0E
ktBEKp5CMZTHqUAAchYCJWbrFESifAmUKaTeceHhJZPAJWpBZgkQFfwR+QokHV6H
5odGHXwOETpji/vX4jSZaBply9MXQoCVhcrBLb61ilVtGZ9W7ARo5KOhU5CBty+R
FDlCg+acx1tA46fe9XSNL8+i756SF+NWz6irKEhwRoRfjqN7qkgxcCMfbd7mPHyu
EyI6di2NCuBsa36DsXk5B7BOuOLj/PK5UiSRx1Ssn5mmt4MsWP1b9YcLqv2drsMt
LyyyU1N0+AOyJ8SVyGjtbQ==
`protect END_PROTECTED
