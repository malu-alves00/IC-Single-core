`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UkCR8BCpJvsgxQEOoyxHMdnPUvtbd4Ciag7KFXF5S/0k12T1WXCAO+NMx3JhO1bP
S56gvzdJEeI16uqlDABiYHP2J2yBcAPoFfSMNuOmgn4iT//RhslO0c/8Dx4/rBSU
3og0jVhuEQussVZytzejoKn6im1Lf+shRu6v/GTXtcqhPkp3UO6GmJXNvM0jIkvK
IR6HmXjyj71iJmrwLuUHYVq0PIYAX+TRKuI6A40L/KLxG15Na5/rvgkIhcxbgJ3U
0nfTxhi181MCzw/EAnlmrLkk5IY2us2tBnelZsaLe/2il3V/rG8V90ilgnUiQQvr
EEfBV5rWk9sYja+YVfta33F5XshfFRlIBOPGwX//AC1eV9M7/w2/FaJqxMX3phwC
PdE6NAcK2FE0+v6ysr0PRFif85h6PYlfyl44rEoAW2xhvlyu6DQ96W6A0vz7m12O
W7NWGdmfe18alH7Ec6ATEYPQlLE+ShP3NJ5TU82/oKP6dzyT+Yo+WHG5U0Qt7m5I
SI9exVCYQmOjhcetraXzjRidu6YPgKs+DXZBo2Z2WpACbJeKQ4wd2ocjM9zSyj8C
gWGPR3f+83VNSzRMhkFXwfqVa3vKVfbGNgUV43PTy2KUS62IGYFm+xivKPI2BM4P
boIm2Om8Y/nn0WSwk8P5fEav4zqL+q5BZxfdMrvWNsuORyvWlk0ABlvLKVcyjCFz
SEmmptGrASgx9SrL9Z9V1xR/89PxUH1X1aE1JZlcZF/rdppjFXLdyYYbosNbnp8F
onNz4/fRri5VKyOl++J3PhJvuTlQbmjY22rysA33Y0lNKqP9gAV+JkPqIFSCNS0C
XELEa6rFTD5yLnXbSmgg9xKGRT49kPPAt+05WolSXSHDZyRQsgMv86OAdxQsv52D
tic+7irs2LqdEjXNZsIwI9hieqN2TuYu8KtDW6DuFNXm7aoPCywBL+8zrvLhILm6
AV17XX4g8y7mHE82ErHp0sd7zR6uE3clP6kZpAONXpIwAaEeRa/vF0YS/cDaJ7Kt
Xdlj9YQofz7rYSf6cWSCT77xMdD0A2AEGmZJxLheIWRtujuQtNpTeCbAiai+kBS9
D9jJazIJBnZFaspIteoPwr5xVe9MNhR+HVpHO/4T3+wkNeMPtxj/q5P5YRk8+1Ox
+3Dnv63HNJMgVBiugKo8CxMWW47ETekt4IyOuHs5LLQ59TSiSJa2n9MeIrEBBBFm
wUBa+G7c7fnSy5DXThL/S6fHBBg0Z+jeDQN845H596JGi80gUjSr5RdMTSaJugL8
PnNmUJXN065kzAjgOYkq+wRA8tKo5wgggdMdbJ8IWoz9o1pSEEsV2uV6/cFReost
9rotNsED6TUKTtEMwnXb9TKfryl18fJRMKLfPrXW8j97L7cfQyd7AmQjOfFsBJOn
N0UG5O1I7G0zKfm24IIMqzoMELuZrjEO9ZKhlxD1HXEj+a5WCrDWNFRAUHxZDf/s
rD4AUbJQOPR0twljF1k64hVJMdyfzoVg9aajf9bF4QFf6oHpFnDcu/nBiHfdc1ex
ReotbmN7FRgxVnAXmrsXP89UntlnqeYthd9PyJDKL2fG4jFBeo04ijkWgRrWuO30
UODnBn0Gqle7DcZ9mQklwpIcejqIIyHdUB6JuEOvIOorJs1j/a90N3u9v91crH4X
dAYQ4awhnc+/Qht6alAi3LMKDZOj6HtNZN5Y7gwMins=
`protect END_PROTECTED
