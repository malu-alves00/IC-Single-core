`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7uaUp77FZevo5MnNmJaxtMWAzx+0ZokDJQr14QqekPpP8PaNYSwPgqr8G/KiB2z8
3RIVFOd1+VJb1nx8V3RWlVZMEwkMCDKCPgFHEm2ihuO6e7ILb6G7rWnjl4zjWqZ3
D0aRNBdPObFhBEt+yrzE/MpBEJKLbHkTXhiZdGufh2LzYHorn61WmXmRUTr5rTag
uJs5A7iFHHFwAFctPGPBnwJt063r2JFmH9Ime27r1qmHcDzc95g69cDITL4R/YsH
U8PWuwIwlX992gkOnTIKiRlMusvTIdEmW9wueFfElf6nfsT67mAyEv+6/WnGTPx/
g7vRRmJ7IdXydpRHCSVPtN2XlKk6tBiCz96CLQxQjiMvtwGsqSFvxmnViiq/y/Xs
LWCKuDhF5dBf6TsA/3rT5l0x9PSg00DJgxqYZbaHrNCCmH9/aIAnpSuCII7z2FfM
woKEx+X7EcEyMDpWP5xyqv7DuwyEF6xWP1IWo1+SPMVFCeWNG0QsXfYps03XAxGe
2F8hV8Fn4p/lFilfrAdqTsqujqQ+sEVmofYeUQZ/BVcrd0hyg2v8asIf56awM1/R
xDf2MnzdYelZIGS3DUEp+bC/3pIy0i3qIILpB74Zkn3BvJZ3zPyMir6nZF1Xg3LE
mSiy9cQiG1Q/VDi5ECggWhe9gU4hxNTy1/9kM7y82AubvR9CbaTVW5R8uFOO5Q1y
6QdE1Wyet8jzcwCfSFki8Tu4YVlyLn0j9zbbrtCHNq07wYVHNQjq4bkTeoLRI0kn
qwceyb7yUhqg/kVZ5dMSH/Hra2q9RCb1I8xbAKDO/aVS03n+QJMbTvGtvCPm4jGh
G85njm/oLhWP2IRMMndaaL5eyqhkE5H5uJzIW7gx0hxMXT5cs1tUISakVJt5dD1K
Ij7pVlBVd8rO4zsj2hK8Y7IQsDvkye9v37ERt852hvAHeEBm6pEFpUNgg4hBqHtV
Nx+TEW+RWFYlvNsUHfk6Lrnd8QQweTqCgl35dJdXUa71SQ5Ogcf3F7b2jCsTkAI3
dahJx48ggBts3XbJmzhJbdNxuuHVLqY5jbhh4jnglbaqXkNrXKLId7ybYvt1V0MQ
OVA2PV6e/TWyiRNirZAHC5qYBQ39VwRleqJ3Dy0EEXm8iwf07e+o2SXn1wvEHA5u
T0mfd2bt2IdWy28wnOTjM3w3/en/YB/xg4vilM680pzaXp9wRK7Mz3AUy0MAsfvl
3WQzqgzlW0U+ciszC1TUzSrGmxJTPpWNLVAkkiDvESHxVV4LdhH4v1APeuvdJuyL
4DmZMoweNJERbviujp/sXx+rB9bVceMMz5t/3Z7RRWj1kE62dJeo6HneafhDiizn
RBRYMFamXcASfRjs1uhofw7BYXbDTk1p3rB+p1ot7ZP44aWaX4VCnQRDfh/fX9Ys
H0Yk9MtIqABdvPwrGxTsrA==
`protect END_PROTECTED
