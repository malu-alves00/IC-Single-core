`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
W6Cpk8r60Jy3PDgOVG8M6je7nx20GoIs9n/WH5kn+tFtKEuBAbjmLzMaCfpNs07e
wvUvgr4D0uUzudPGYhrsBxskYBLUCDqndRUC4hWqLki7NQHDP9glXq8GNQcL5zQ0
Zi227lKRazIh7Or0r9UpTMLNgTzX8jl0xaOV2UpWclE+BQ+h9af1AkZy17pAJdrg
PWbtYjvK31+F6oaBLqS0hBmEqDCRb4dgC+qlE/Um8fAx+YwRkwt3oESSC9rbm4D9
gtUl10CFzO61MW32GtFq5xmrItbnlFoT5bRe6J9XatH6gVTWbXgX+lsb4WBgUYf5
bdjfhxz5lF7mwXk6pFw6yTxwAtpiq9Brswx0NUJIQFHcPTOFtF81y77tp8Ao/a+O
fdgp2nV1401m4q+D1uY0KkCBMWQIfBswckUvJVjq755ovCn0RIr+sTxg/VV+ZRN6
hHFJYe8yeIATr/S+ssW+EteuG80M60EFknVDHTW1AJZMuBWsnE9U3YwCGe9OPqVO
5UuYtHYiVXTyNdKj1TJ6IviLWYfWlk8WwiTogT6Ex2M0A3HJqyCeo8OtJtzNFGz9
rORyjhbGAk710udjPBfxwpte9wMTGPQ2btVCiUNBd5fjw+BLdsFbKCzdRDqkno0w
GxLZ1z1taUp1jfjS9WILhY4fXr3Z6fTN/sRGkZbNlR52Ktz3dZyHBcL9g/X1/xfB
O18+6TbdJRmGC+jKtkzzN10iZaesT/PeFDw3V4/oJuhWLHj5QL5CNiGivknTzezf
X5kp19HmTpjgxwC0cbxp2ZGvR80F9uwfpfdTUTOzT8mvPwLHtqyBj6KfLWHH5O2T
UhUsVJj0zugg/AJv4d6w6EJLo9ystpnsP595W77WHVXKOwo/rBuU/j4ywUGAXelH
qSvC0IPiKClRjS2GpwmNk9nNxk2iRNp7IttEM/Y2HJC7w876fzg461MtFM5THkMP
nxhkBCojm8uGfwde73cInlq3ZBKjLaNfCknqcsWHxsfMRWImcvSQG9UEu5u1gtq9
a/X+lIStPzC8QSFC7ehKv0Lbcdiy1Dht6/L4JlWHo2O4CCMJgVnMZKGDhnEo+uyG
Ok8+Fri26mVLd4k/wNCR2m13tQuNUM8JFgb7hKWtyZbvvauwDdrPlCWU7j6tY4qN
Vn2LCkAQE97RSQWKH1ERpfNI3f+307bCzZZLA7eOF4bEhc6yuM4OhZpUDw+U0EXz
Ynh35/u4vZ7/gdvOWXpj9PNAwIvU3VS8+vCljrogIFtYMV1vbPOtqAkoUJYBMof5
9wAQGU3Kfry9sm2IHoy5UiLx87UR9Jy9vhYPV4/mU+kjGM1k7iVDILpsQM67EWfr
Ym/qi/c5rRK/eadbvD8QEKuBahZBLkcsjsQrCQZWObdGmeGn814THUCdDciipta9
sOsm2JqLYYz3CfvFWwYv2Pi0e9qskDSGnrwBvJQm/RsSBIN7U5dVUsd+MJM1Kroo
V0amwtFyXnn/GLnubwwB388fRSncETx5yIO9wOfp4Y1BNygmbxHT93nd8H2u3kUq
MY9HA5N0p6uDhD4jRHz8lEAqMAzaCLxlhcgw3Z5B0rbOouMAMrd5vhdJVAXq81iY
lT36XgNwT24eRq3VNVc7PJ1U4kHfNOTu+OZKs84UGBzOrBPZEiONw1L/v+eF3z65
ikhW0R2+VnDiunEkXBHOALOiMeQ34aMvDR1urcyF8oMW8nyyJQ4cw5sDRdnYzaGZ
pmYw3Cmg0mVg/N0g0UPbhobUw7AlV89W2yKAM33sI3uxWx7LMVkDsmaEIf1nQgz6
GO/rSOxirydKBTIIVQ+V06BSctrwWDzG2B8JSZTcjDdU5Xgqf7pKRqorTo0k8rME
gbKLivI7cfzKye4WARU4nCL+FxBRveWOTNKP9RWXnBY7Mt/Gf7XDTHyRXYz9qZR/
1xGm/lq+DSTNP6gmuCf2E1BHG2qLrcmRPBJNVkxK1R3wK23kdTJffH0jj9z4qNcK
tgnpK60YuFyxRcODAzpjifaBXZsWfa1WkW9bQNn/CgHo5QwbEWe55LBL7aQjC1H8
kCKjvhCaUwTudqa1/LSBcuqMHGa5LgE5JubwkKAx82V0rsDu+R8PPPZjxbJw6ptk
pnxrvEueCRMAPL4sh1935TRVgfZjI9WuYB+/Lct+akOLN+xZ3lBnC4/gAX/oJJlI
x6giY2ZtfJui/M+lgCsugHZqjF1jPiR4DwmEbS7sHWXk/iM+ozJD+7IfDyO9rCYI
gHFctLe0Elt8mOSGphC8/VWg+YduT4dogPD2Tp+R1YH3e8jSBYuqg6XsXmWD7/m8
NA/p+8giu0X7q0NyN6v2xfzNkkptnXfKV8NWrmeZeEJpBFCqbvEJZp4yS55tbldo
fjyTBoJ3lRGtYFlrn9pJAh71qUBJjEKFn0eJnmlnFRn1FG9rm+KgO4d6V/a1juSc
4Fu8EFZCGvto5gk5FNItwHskK6acF7/8Q6CfAD/AmsJfPTDDqSWa02vU7wHt3Nfi
RwLvM9QySMLwFQps/37TOiRVRCQXQK7p83VP8PojatxCU0yOWCHs2UwT6vb/gmMV
`protect END_PROTECTED
