`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/OoOm8TaqN4rIrVbj/IAlYqkaOc32U2x4NJgvaeXig9qxUyolzbpGnioJInTuNOm
Ix+FLUjnScd4ZZbJpuV9qYlxW9/vFfNyrZ7cblQgDLjY0FiEztvyUN+pgEcA6qUN
3K3AEcSherLbgdgk4KKAHR8EkpM0njd7bYySXIK82ccMfVmIXamRi4L2j6DTtTaA
1axMPyQpa9PdAFHkO4Zrgfa1sAVkppJEy/JWBEfVDEru7tMOIrZuvzNEKwzcoIzE
c0Ow4OK22HFSRhOGyjUSiQFvIiuiA0hB2l4ZvMu+lyRiqH7ZGVuWM7gOOKHhTKYR
zvg08/beq9MKAnpGtaN3ZWG8kRqJauMpfs3bKA0SLWeUMDL8U5LXmyUzXI3/3LEt
9F0Ord4CHTt0bVZJ5XI5Eqap97zuWoS49QyeOh4py6ClU7om1N+sGv+h6iLcdCby
5D/HEJqYfnyDrQ33rov3MMErQjJqkljz0B1T95I7uQeERSD5DvLWXdHUgBB6c/6S
s+oi9ZsTBSzHj1YGA79JrUS4N4+4r8KzhKOtz438+n45rxiYLVoKFzre7Z49mgBQ
Z7aSBQcZbLL4b0IygPDw6wRZMXJcfFH+ily4rwNisiLp8f0TQhPzAqOHHJ8QC9UC
F92L04Pzg/zSi8ZWc3T89p87ZRIg4Zl8fKE/Zi9rHwprEzr6Jqxqvdbk7m/i6JMs
TCFaUEoMlx2Zr1UD3rcZjxi5ezlRffICnYFbnfVRsjiLzdvaACVsvVH6mzcp+inE
sMryCdMoX2sOZnBmmvgMegUEoJeQb+5KXZPXw1oPkiO5Ke39TcmDKloXC6q3egLm
zccK0Q3hvHn+w/hHYgFUxC0nCtAeXsnyRE8qlNQnY+ABoVZ1hjPzEur57Jh+DXNb
aqzD+JyRZNEuCRp7bg1pr5osRLXnXDb2asj+ulo3pBfK8czOw6wmGxe/U2glnFdP
rX0keS+RjZcnWiQP6CYl1UmAx7s4jY+X6SttFWDiXg2EqDFvHh3dE3HQckyM4uLb
yL6QH4KWINYmdrCwNRRVt97rHNWjX9CMKyUlhSHIhAsW4pclJnF+8Q4jDuDUMUEu
SDCY1N6i4i5rewFt4EbuBOhFQR1R9sWq3v1PyRUbcxWLm3Ru+qoIEy6z2IZxpJZh
CmFq0Trn/SaBj5CuzYYvm8lGeI5FeNJr8XYED1ku4NWrZQ3zXpdDHeR+VCQV18MV
1WR0mUme9wT4llyBfwPAQl/d6r1swx+fynm5tp+Xtj6W17YrhiVeLzqf0Ny+AICv
`protect END_PROTECTED
