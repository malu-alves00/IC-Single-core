`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SQ2e4shMuC3m23KWbx4B5dbv6DFsWyCNB5IEywxei7u74YyRvCyB+OPWxi+Wv1pV
I/hXqhegmk85VyEFjWIDmgVQYcWkUlecrEIEyhOA4OHY8FGlXCpukW3txRG9t/lu
esRO/ZYIDQZVsj3TQwjup0Nx5nQ4UC28slQHLArdu56VY1hpAcg/2553kN0hVnyp
gSaIxDieo1hd86+PcXhfcLvdT4JB5/q/9DOSEOPDLVYERo4GhIPqB+HIAN42UxV1
iHZoC50/B60rh9E3pbaiWg==
`protect END_PROTECTED
