`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qzjPMGS6UK/9qhOdcmNldyY8SO69qM6hiXQLop5mdLLdyVhcw26YNqMwmqFi3V8k
nRUGzhOskXh+/xzZWqP4/3Di2QzZEr/bSbftJI5YYDEBNZv6PN+h46hjQxaV8ZsA
NkkZblC3TeuUUdeCChCi8DugZ7ofp59tysonQzo+n49tf1bqIT3wEsMoT1hYzPjd
78mgaqZMHy9WxFFvxRJtR6MQux86LjMBbW8qRZDBVXEcmiu2glvWVGrhohpfuQwr
SWsKOKA/8kREXzPzRe/Ya8JiZwhRJQxkul7ryyrrQlOlSOI4uGCdlWpMnkYc3ORb
tEZB2XEKixj2+n8ZClQ/qEaRhl1WRFtmZ1s2HjeP1lcVT9e68CBqOUF1NE4huQg1
Yzydf5LaP8lawlex/1aWdpwl7MW5o/KpisARiOCVDsHm3XxKr4n5we7/Laf9XKWa
7DCedxenkhzo4qnBARST0W0utsKjCSih278240i1HC2DV3Ld48wIu8HgFzLhl1/x
ZZuETDXZbF7Oyhmh2RK3Enf2yu/iwsskQLioMlEXkoqDu9+XUbaMoPLhOupeW4Fs
WcrjDpD1qg+4IDvkWfd/z/7/aUVauszTxbu2LiKEMWTrT4FP5nfNXdbjzAixAbXI
RElFMH/6Sz7gCigSifo2bQIPMzGVt4zXPRfesTa3uRBqfuvVQRP5OO2ghtHqDy9J
nvnd+sJFNWjycBSFVi8EmD1wJJmLiIGXm3yxuZZjfBT9W5qx0k6W/CjV74Y6eIgv
vBm4fszRek9lhR2MLtn+kELj7uAX1jaLRkx/EOG1L9xNRPnLVWDNyx81TRs/erQu
b/i4dGP4uSrlM6rhq++k68UKMaaAZrbUFVakbNYzcD7AJ9nFJPn3j4hQk892uVLx
c/iwrj17w/cN3XIcRjJLvP6cdR4TG91Ej8TnU+6P3XPL2Fbzwtbf7BW9AD08ZO5B
l7foLNzRbxGXG8UsultmIuuwfRs4U7YRatVhj9nVaxebzEdmVkidA2ztEh2jWP1Q
R8inrUMaNZbvLNAqjuYgwTEBQWjhG3Ca17UdgNqoDZLzChH5zlns+ruwI20erARH
UahPcQDLpISO0D6+orLc6P1e5KI+MArprBILJ51767Ar+ic686lBv5OsJs9rbYKX
/6tFEr02/uC3h0FYasD73jl/PILoNjcJ5BSC+7p6W15SjboxMeAbrn8t9C3vDXU0
j5a/Cp3Vml9XvMqltTNGcgQkB5moIpfmBAxrB2SgBRQ+UbgsD/Nz7MfescBzcZmm
X67O+EfMe40Twcf2qRelbyQfmUgpP01ZxrpxiMqzpyNUaCRzdw/ik/MvyLj3mKQO
uoYxbUNQu0rtXTsuU8MPZqv93rqKjl1opBTdD0BY2mNRxurNlWaTCo8+sdNtGeVv
++xwyM8Egw8HK7TG+W5MMWopLf8uGv1XrOUTOyln1tBMu+xUIL+ZbKaI3cADRgbQ
`protect END_PROTECTED
