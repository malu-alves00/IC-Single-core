`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wNJZHrhN8KOQ8xzyCv49cVQQB8KSeKLPmFZ82oHsrWYL4BSEhydHtV6PgGfx5doC
1CQSAcrTmDTmOVzAuFgcECuonHWHey11ytVueoGeyk1yOiwSmoBT7crQltukJLMz
TrktlJC8YU7a63rn+IOd8hpMwOAspkYV95+Rf4EepORq+gUSA66jKL4kZRcDb2vQ
SLUIZfpCYKo5yyPzLPNb1XKAt0J9yyw7kJPwovkvg21AwNc6CRgdhLkDlWtESq4J
O3z1li4AEiOU6GhXJ8MvUqoz25Z75RZcicnGTtoD06/tlQ3BXMxUUOM3u3o7LXux
iQ1rKwydZ07MMdNDHs02clsQuyvcPQ1Ax2RJ2zlPJTcJH445jkd5/Ckz4o0GqHSa
3bSt/bmdz0d9K0x+j8RP6HVU4p13G1gbvbDPdFXGJRzmNtPdP67D/wajGlwXVFaC
wfYrG9oKfVShwEjxQNhANsDWb6s7Ym+QNZ9Z86nOU7NKVAPX4xp1O8ZsFHqdNDuh
u9hm0OYwhfpXwilIEMlLIR40ie0VQI7wa/A1RxlwfL5x+vtGs0DkQx/nKUe9JJgd
B/jreRAM89EcbZLtt9WLfU5MLz0U/SbomCSEQ2L84INrFS08hVccXOGfepUMDy6/
tGunzYg1DO3wZCr6a/GA+nH4VlY7FdBltVlpez0PsDlt6+nSfVvBE6AQgCVGXqmT
dEKXjMyU3ZTVeI/Enpk7Y8+GiZERLm+tJTonZhLBTcNJRsfpbmE6wZUOHjfyQfLN
iDMlrT8iZdriPh9kTso9agDN4vBJ9vMhTrVTFKbUKvcJcTeKvHPOmsKnhawQn5+8
VbFHrsaKIlIes67Ql00kHv0YOzYI2o1fMRW/+zO3QmAKooDB1xAYeavPn5wqmFrm
poQeuV3IrKt+gFijAHqdjB4fhUrxUeUe/ZtUPu4kDpSW9TQ7Z341mqypgg5Dha0k
cZ4/gkJ5v21lnwPADfKvTwLgrctM9V87ywAlUDCu8s8ex80tS+VBxUDn1lFce2bz
kk/RwJzzjPcWYzmc8HEi4LcyuUXdgEJJlVmv1KTHSmeUDNEidNXHJArz2IrTDYrI
1QbqP95K4sPXKVs9Av/mgw==
`protect END_PROTECTED
