`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rBV3PUCMWEvDZmK+WZlyH0gQhST7wKBXs+jP56+hkBbUEJ0lC/GiGrsPDRGZXBop
HVl7e/M6PvNqmoBVlg8fiTjxjZfp+vuoSIawYs/EY7r5vxNPkJ1l3lzPYE85GdFC
McBjUZxtGB46RlA9yMolSXDIO0yIlrKNdyzND7+Q8XwzXlRnCCvkHOVJznbmULOt
hJ3mJG83pLXABSELZXYuE92Au8dpy0dBF02hssk3nyelJXci4VIAb5KgwVTial5G
NEutcs7ROkasm9A7LgpYIaSkZxq9ghsSf6Yr/JvAYMAaOE36Gx1C4qGD2IYsnrpq
Vc2WyORZ0ny3hwlrSNTSAFIqj+uuisC9azqxsKzHhjbeCCFDM4k2LS3Gv4qXSlrh
8c4FP84cyfzPzfoBD1C8GgTHz10kKYgZxJYDLD1mNQpWB6nvEuAU9QslFPAC0I0R
wI8BZfnJtdIFK2/giraqoNNcN9ZVDsjROeoTEHYZws3B8ZDzD9Jp7KOGj4pcPiBp
6FB/cj8jOxZzYu1PzkKH8gM742ndhDdnCqZvxdzSgdUeguG9PkCav1RtihSMPtiq
uG58ypp7VqnRcEbE2f2Fg/368LY4aXyJzcV5kpko5xmQUlRIXCtQBLLuQXLtCtjW
I9n2mUmqTq7sOFBKkNEFJO2259NfTgZZLng1fKr1lElauYPQBRtpPriYhMyOwBNQ
IQDnJJwvzjOrHMv92Gn00QPt5jqGgxZamifGrXyd943AbuGYJsfqzT3Bw4dbcu4x
7ofw8ojZTQYr6elgjCO7H3Pnu3u8HgYwNChzj9A7WXvghwOX5E13yBYbh/RXddSR
UyhSJodkA5i5zQE4FdU4Jl1n1JUvUc+BbTTiF0EZ5yB+lbwpEZ0L6UlFusYDqkUD
wF2WWlE7qSzg3SOAmwofcRRJI6ZmQZbpC8HEePVuWJKx/mlp1pPprHfBAwEEQ7Rn
g76nvIz7UyJ7Z3CBPARUxqhOmYGk8vAZfM1jQvh37bor3BP6Pb9YW0y7e4B10EMa
MKBHtpnvZvwZUwO6EONR30w4xa+LgY42Et6dhyOWH01GJ+6T/Q8mNGIIXWUlFhBE
ZVnXWCkpnyy0E4rIAurAcW2mhv3hcKFkuwx8wPGKBZWx8WX1nBzdwwEmM/ZiD57r
aV22J8TryV/WI3gce7S2DoLYBzVPmvoL89ySJhATlYXOAbJgNrT947vu4PWcDARB
AWBBDf5isbZwTFtLTBlX0Iz1aEI+LhjdY64lFSaWO4YRHZVchQlKqvqzkQwzTLr8
Eh82IOFagU+FKgkY/4Z07Fu+Ig25jDFEy3gXXVzbS5hMFyKTAzo8VpyLM/pb5+Br
7ySB9FYy0L1Ug6pxcDu+iBGpWl3GVO5hJqReBZXSCsNpgVMKsAKbSuOABZhc1ijW
e65Tqgi8xTC+SJq0rwGrV4WnRle3T/8c1IXYajAm72O8ZJObVzISv7taXbRlBeCl
x4MxetP0wW9pl5EGwh25QBQ0/cuxkbS7waQsaUI0pnIVgQiwYYyQuzqs+9VR1xBn
ygYLnT0OHQYboHm/GJsMCaZrbqavkm7k1FbM+dQ3R3lYn3y7I/zV2JihWIdb5b2C
ADwvrQS7Aq7Y3n/nzq6IRWynyeUpW0hPblxRHbMfl77GhxNXJBTIMPYIPQTp9UYc
KyqWpvKx7vPUj2ne7i1S15K1k7GjuQQlhRQ+O7LbePWfHYbjvIDwKY4aO+FVH+uz
xHrV5lnPGv7kTEMjd9xtDb5I3zAhL4L87Pb7OKGNVsPtkmfQcvuc3r51gRaBzAX+
Dw/yt+jRidqyDmPnvb0wPiGKT9FH5EZq+wAwWQ+kJVr5avcg1KXpThM1D36i1+if
uGWL5joTwY5LFkJyr8x38gof9s0dU8n3u2pFO4RVNf8o53z4yyYq3rVlVF7HpGiX
TeIArz7YFa3GxeaQpUi2NRYG45igNglbVj8bGWWwfFsPKTkgAQ9yq289BugUSAoK
X3q+paJZZ7d5bOEjfraYIwsXkyBmbSxWOU2eKhX1W6PwCf/nlc2qSc6roItFiXnX
dA7C09dqZCEBPogm6dfxL10Ezg9SBlNF31jVQBGivXv3PuiU+jTRHqXYtTWKD2s7
WIMZ4EOsfohekoiw8LVRLq2f9w8F+ACsx+H1TgBmGyAuX7I8luzJuwFwngc4WpwR
vAjy21xpDOZDusCf3X52VH3KwF/jdShmS7us6/dUNyeAdkUG6tV8NM0MrcdnzBo3
/HcgcVxHLhUpIKLukMDTY6TaGq+EPzouTjG1F65VNoaR/ypTrIdexDKSCEyymLYI
LJIVuuvz2VPp//07d5zltPbD0opXig6OGIJCNyHplbFzc5ZLTdpZ4BNa7Xhs6t6W
qpeBxqg74jAQCVFMJL8HU+27TOkBxAaQIh+t8fAr5Cn1+UA2oG9fJERs9+ZYyHob
t3KMu1aGYVdB+KGdrADzaKNPlXbwVLai6N3FdKtl0ks2YmN7otKBHk6PI4kuBnSq
r1iQuNeeEDmlGLtCyQLj2mQihMdUWbbWmWKJrI8MKaPII+yTQOQ6OiGPGX3pbL9f
yqhdzKJKFBqU6zZfGIVTm52llCTcTFCggHDsCzAYQtp23DZBHpwMrhd79SJdrupJ
NnutvEPOLinPjk7a9M2tOfiN9DAHRqrKhSXTFPASLCSmz2rC7s5U4zibCBcFB07A
wpVeLFGsi2CDY4OmLUKWRpSnWmO2IyrBHc75XjBHRupFVLXAROaEVS5LtD6avjVU
cdW+YkfnZf60zNd0evSg3qYc5tnZEo/nuOjWmtIxipRUCh+nByhi8jus9pQ37Uoa
3Mjab3YWjEP8NnGi9TvIUKEV1kVpebnyj+1+i5FuLj0VPfEOcgctMJKAp+btP/CV
BG4VaYHasDTtULla0jZTFfsEjSbKkg7hpPg4JgrU6E2DvTnDPXYDSEeoUY4n+D3I
oJTfX2U+Z1lUi2UWyG4ouJReYh1fq9lrg9zDTnFr4r3UbL+cjmjS2gR2T8v/N04r
1ghNn8fukVA7vN5f/exo7+TjHcAUPf0eMbq84ZkUxN2cQ9JxdTgJ2ZTDDfzU3LI3
rCqxVvzR3fuymDYbnG6dz07bxMp9LqcB9lheCdTEv8Q+jLUPODVrT3/TrUWrcl+1
rzLB0lBieuKWD5khK+HneGey/jDIBN8DrkGwF95mPfv4KCilLmhKj7HTrQ+T2jAO
/OZfMdFB0hEP6Ihp4toAtPJ9vprGT6EGuBvYVhz+6rcYUAvXGmtOSZjZ0Em6GohD
Apjc2DY6CfebnRZZO6P895IrcEtiXW6IWtoXmRBEztvMW8qMVhJHf48iLKMPw9Y5
7vn/HbPCSZc1jep74Hkes95+S4Gvb893KRzOJOTxGe3dNviB2qEfxwgX1T2Y/qxB
nK3UbyleAXgCGJR2MMs/lASRf8G5KtWGeAkpyAnb2z1OPU/N2ru8Kjuj56P/5/VL
ANwx4KyotNXWEX6I9RsDR54ixgym8n+pVMirdYHMqhB2ny8yHiHgHg+1kiUq74vG
7rRN98K5dz0J2dRTEkepOH1YyNZVqmJQZYykzLCWXHFS11eJ615MRj43omv3Ue0Q
jweTutIz8A7hYDy8if0i/2YKeRQIgunCP4SbtQDAfz6Q0pNmH/bMDe0ldvHHkp9s
NOsCOns7zJv1WRXz44UoaoI63yCjPc8nNvXXzTOb8Xa1vgbC0sP9RrXdXWiO1U89
8pc0q9eHGLrdZoAmD5b8qJWQXFcyYbwq36rFxm6eUpGQg+IMiQPCQ/1yY+fKRq68
8PD3he7NqYsm0PSDpWuXeiCvFzhXL8bSJYtexnnLHvgEaUYTkm5M8MI3AAaeomCm
2MyreQHlKM9EvoyPunu4j4KAkqN5gu5Mkg6PguSMg0M2zJK4kcRf/GUBxGQSe7+T
eSp0uEXlf+WB/QjQf/jY/HH6DBoeC/qzQwoyX7a/rbF6UYCnF3YYgqWbheFYkpVo
Bu00vM2hWjKiS/eaVbhUA59inJPxisDEI86myDgopQYzZCUaArtfI+cWYi1UaOMY
GZt5irJEtIExRr+gLEL6VII9AZl5XI5P+4YrAuKiIl6wnAAXJarFv7Tco20XUvQ3
+DSuA+7oUoPxJMbiYNMwWjH0MWObVYpA9UKrDRoKKiryF4RyU1lVWbm62vV2QHWR
g6inHwkGc00Y+2DHyCLw8wP7YiSzLQ11ZnloZnRGRDw6mtSsKUqAALGfojvLeLE7
dwDsRoEeVdTN9vJBffFBulQiKLgUEINPkTJ/odP7pMFQQtQtjWzy2w0ZJRfZpoJe
31JpN4tzsV/HPFBVt8uibLR1cO84FJ1JK2jufjHnORR6thxhTJuGoGRcoO6UqNgD
48GNlGSMoNnUsc4lmN6IKsdX4gkiuPeKumd+a4/spiG5k+UIo0Cd0QMQVvoBypZI
GfdBcnu+PqJvBJpTDcdglbrJ2eX6xvdN8soaNAVVLA6keb1/dgcB9/blz3612kQx
RDT2bLLxydPhE/uft9KI32VM+WCzDcKM/Y/Ahe2A81Z/sXfJehFI3gFxnBGyvJCG
RswD+ssSBH4tdJnJAa9rV7D5ddENnonqp5rvEEFOm+AkliqvAeniWVO1aX2tofAn
PwkTDX+z8xqdFhvQIO7Vf/usJk/wf9GaC8Haq6HpY23Tct5WcEKhN5VDvi4qiGW+
7xww9XK0r+lRStb2J9SkOhQ2nxt2qXMckNakB+B5NiLWg4A8iReovj5lrorx8x6w
mS8jN3tQbFaAWQ7IFh2rMCSD4YzUETPkHMvg+tlcp1LF5F/RlvnXGIFEhP3zC700
fy68CGN4rw7wIc2PksD1worCV2K47+y0UpBCQBRlU4LzEvQUqtakqODMTZFR8hkd
r//W5+Bevfp9FBxwG1mHj3IwLl/hOxwnVLx6D0Ae2ABR34vtVjT2rg7VBb1wanuZ
iMwcMstIW+6UudOa2Cn5jCp4vXw/2rfzlB0UQEQm3cUizWlgl51DBeeEjbrwahxb
ySVji2h9kZqgDTeAY7y5ru2i/kLY1Egigzgtps9K81F5tfq89Zu/DzVia7mrmSV2
8kIas9gKBFbs8qFd3JBXg4Mf0Kp5Vz6gCjAzGjzSfvEZGPJ9CBVn/dCPucAAFBBV
h/6g2Ix8wya1VLKrAfTr01V7K6CrVgTBImq29Z6+gtbdKUdRih+WRdGt8IEDDshD
tIfOi+im80O0E3B2FsqioETh1J9Y45lWaXto8+WHD/faVvhs+SsC7dPJZ7XRHcg3
iviIaCXwQOte/mTjnEOPwra0SaGfvB90VKvSE+zqXDXM/xGzZaH1qPway6sushMW
foRH/eA6hPWSz5jvs1k6EoB333/dRW1iX8uWG4OB1BxyBrzo+d0HoAnNuOUfH2dc
j4hPHFvi5UnksU6DO+x6zhFJDpJU0HL6XQ6AdIuVbBdCIdXs+HrogG9Zq4xOiH3Z
OW70nfocpdFT0B7DFY6FtNjMYenQXiDXlm5r40X7XHsI3RdR3BO5WfT//BWMjCSB
gFYkDAth3Su7aemhZ/NAwFtqqJPy6we8dfG9tL1C+vGvCuc/LK4Fe7BfI8xocBnm
E+d2PVIORZAgOyvPnQsggtWMaHXNN5/GfagQdecpLk1FN0E8snZTmxd7je8xD81j
AjUmnOA9BRjxDkoqk5/LfxBmSMEU95+i/+Ara1TLfoX2/9ueiwE+OTnVbaS/zdFm
41ofLoYtba28SW9Q0ML7P5uVykzrrbsQ4WS2fX4QzTV3DLuEryOCX6ZZabjGPCDr
Ydd5WhqUXFQsjKXZ80VUTnS1AAZGPr9t2bYOTiQ631OccHdpA23Ph15O/RzfX1JO
Kz4B5wyZRv63MWj/5xvEzcm8rvaKySnnIaKRfhE8nnT6jbKreZoTP1Bsjd4ahyhF
VR0yiQVFJNhhS1Fr30ITc2Qc55Ss2Hu7SMEr5nHV3abNCNd95GNemipr3S6bAW7G
lZB8mkqQ9WIgSO8q3slBuqcLNH/m9RuXKNIZxweu1DZI3E6Up+vUf7tnpJuRnoyZ
XY5sShLxI4jJs44sHIk26bIMY89Pk4i9fMYXeOD4EQr08WIz6V8z5Db7M7ujrjie
jfOzsuiqIBRH7gCLOMLqtSm45VkdzRZV1L9cCGxAnS6OW5dtJ1td2/ZL6Xg/VDTC
mSRX0OVqTXFQwPZzqXQUcuyqMNMw2RtwXDH84L3CZbliL70jt4X+kp4odb77+OFJ
Sc11qqQ3W9kqjtjtKfZCT39Ltq55DgGvgOk+q9hIbFfvwRG9S/2tPJ9t+hAPOY/0
XL2xlly9sFvJw3/N69M9laBHiztbm+cbt7PobQbQp9z5ZQCRNpOVwYTjvVPPREaF
KJMgBey+AZ1mzTMgAWRRYjF82UW5ig6sNXTAw0VzrX6XbAP4d+nFU8uttxhhIH1i
rhhp3pvr2mGRM+XH3OXEuFu9oDRraiOh4ZtOneebgERkmESBwH/pH8AmQkFnzgdh
5hh7HriX20Hajes3oazA2X3QpjmT0jydmDoFkmuzM5TD/ERGNtUuuOcSmgMqym63
JU1r9x0nFIBKhjlbmCSOud1Z6lem0EGr5nTM+uNzK7vz7Dmfnism1lmKcR4bE5LD
TBAqHCGpdJnfeqDe2GD8V4nAiMkexqyI2Crtt+RoaPdLw2Ypy05f0b+mQnhI9YB4
S4VOdvisZBZ3fNFB+vHfS1sxyNOlDWJHQFMhqJhWZDOs64XGlLHJX6GBsSX/RwIi
zP1SMhjQd3+y9u7jqpolPJe5iUozxMDfNqd2+/+hRKXQd3fIqIKpcDroX20axfZW
xmTpP4Zqi790iS0aF8qROmJuqqSufMSSuIeJFM6iikfrur0qvybuZxHjko4heNiw
cTdA13IMu9ZMMryQHdkjwH4Tj+ePoHdEimUQ88nVaH8yE/zHhjWIQt5iL0X99mTT
cWBnCwHtRdAks3Pf7Xrwx0DJ5YjDnyuBS18RiGnydqLDQRd5+5Ggv/jz/zzG3LTo
730U10gEW1wEmcDUr5nqCHt6UjNwvhpDG19xArOLmQOwzjPFyPYPB0JtNmq2Qfpv
nJGzUM3MfuOBgYCmAZj2j2Yc67eDrJY2q29hyNCHk/NjVDwjadKb6mUbDNC07ZoM
u9E/QHJxd7nseOba3/og3G3S6MbYFjR6cT6aSt02Po12lnWWZRXaR6jpG5bEkjHd
B6uqiVyNbLPmg4/Vp7q8S+s4eeRmdLyjf+4P5MIylCHj6Yc6HWC3hAw2qisZU/gS
/wpOCYPHII++dN6n3PW5Fq1GFuXAhygNpnNqcqbL88ENRU+O7O45aYmc5/yKrsjY
3AIfRgMThQ7M7dy+bZ8733Njy22JrP3LWfkNYAvOaA1lyMYXc2cBifWttJQKPzO/
5d5XE244vLwmPqxaMWTP8R5npH4e5GjkXPFDfvXRUd7HHOUDfzwP4XRN1sdk6Q7v
B9muDIxlXnxFx8jXNWoHJc2sMUA+As6Ybc+pkNXqwLsMmPfF7OX6d6MtK6wKSl20
uLDCoGn1igtx6/f6U4HTXqJyY4z0aWybkr/O+Q9JQB3puAzaRzCUt4dq07GX0eqK
FISjfNCHwdEBnEJwwTgVkJFlsiy//9ZnQj3XjGR666p12hz9uV5euHQI2I5bpJKY
xkG7e1OAT5osvl+l5Z4nCrgrkAYcLS2wzzj+RHQIwNQ8ItE2oj15dtENP5V2D5y6
NhkRdMiUn68pMp5KwXlnfiFCQ2lbMWgW16aebaZvOIopqBueM0C9WxXYJCRASr2D
hTcxWCQrxFTl0c7Qa9WXLHiqPSCyEjyOxKZCQnhcCHImi/BYAeS1stU3UKaAn2Cg
U/Ui099sTCMu8n9R1I7VWGe4W58oQG4MnAt2yNj0zxPZ3JZoWhwLHJVfhnWow2oz
rJWsCxKJRWkH2qCDrIb3ruPYsXZJir/nr+EyWQRMSOww0xGvxwPIELeB/YCJxDNz
KqP0hZnvufYzATDVE/wBkvooeQ+0fYrfatmyfBe/gs0KhS8hx55lOIdNDdMxkg/V
+ydpPjMdgBjXFH6yiUHM5sVG+C00o3lD7RmVk6hW4r5gbd6QkfjOg3oXJN1N0GS5
1mten3cN1k2SSQrEmtLnZzWD5eiwLEkT5Wx+pRrHrNxlWcGOvCezRn2UjEGgLjtb
IQYYzEfaQ8jKK9ygOi+GtqupeE22pky44Z6VJ8ksTp50HG8JUMDtqX5JG2Z5qWLA
hM7xVb1B+m0dRJ2gK/nPZoVcwymI/uP7qe6b9Zj199+dePp0H9JqKD+m+GAJNt6x
D9WFgo1HhRDLopQABGKJmx32hsGpl0/frheVmpJAISVWBMFCSUxJM6ZNxY1yJtgi
Do9dNe52k2H2JacQ+ZyHlHkkwvhhfzNYKT1ebY7lZiXXxyxKspvKO1Ng2gI30jVK
5Q1s+Qhx/PVXg3vB2HKFSWv0usZqVlFyjTxz50dbcrfZ5xXuhu6J2N1cUKchSP7M
clSRFbrGkmlonFiunmnbWdY0alDOUsfXqLVc+6FyeUpmAKZfyCMx06mY25guzb7n
fzg60iY2kINBbuk1neKXT88dQKllhx7s0qq29YbZ4FJEVXRAI6uPIXdnvyNIqgvG
j72gUI6jZMJF28deWaVIQOkvQNXvAHM5/x894e1ZBKffna/17PFp5j4oCMhXGeLH
rPCWifTnMJOTbM2Nf9Cw6i6Ic9Z5pwrOi2MlSVqbtFVwA1x89ajfT9ypCQS2IgiM
Z3q25NYv+ozfmV9LClBT5w9EP73H/g9Mz0tSniMCRpRuaBN2Exm0x/ikuZ/HSUWj
kHHKECrBFVADdwWd3PcOY8GNiF7jissVYPGVmItsjpKTjbl5Soig6SXhA7B07r/Z
HRaEGrGSWKBSqgfD1bJ9WsI0M71N8jwdHEn0adBMY92vhSqFAyr9jtUhFhAe6NZr
OMJI8e9SVAWi7nwG94NP3kLosa3a/tKMkaDyuRm6xZ7neuqkLrIWlj/moRxf0yeN
fvOpXHQCJrTXfjp/ytD/y7Lsnf0gsy2sIJ35Hm76ZP/z3oR7kkjl5dKSYEgv6ml1
faOPch8F18Wp+70ehQC9OVLdCEL+1qYtIU0HzoQldKyS6XJuwA4eGakJ+WJp3Txv
nLN9s0twgfy81OKziuSHzWtBWywUndVdG+OCGcFsJ+yI6MHeMuBY/Y016v8VsU8C
EojAG1VFfq34XP2Kj91WXM2UTT1nA/xtFdoG3AE3jyzRVC2Ajj3WJGJiBw/c3cQw
grY26G+rtt9NqnXQxItmblT5SQ0KQvfALr/8jGP/Vt7p3QnEghn29UuiLSKUzA14
6c1r0RlJZ+juCm/h8cOJFB/znGzI6JFmfU5Tkzbk0U7LfeIjC0D5tiYckfe6rTld
5svALlS6YQv15tBVuhRFfMG3UUyf6IQAKw4KTjxWEVYg0aaB0paQZXsLmAn4KfiV
/HNfvq+hbUmzf++bGHlMDVYAULqhmsbhiFaVZ37bB6ITjWBku9l5OU/zqL6ax9aj
xGtKoRf3uFofs5sbcgeAoYvkr7sh8jWZ/Oo6JH/4TdBRfu4CFJ/hGBa7fNa9ihdF
ot1Vd6apKtlax3ZOr6L6hn7eURmvtkbhd7HGzgyrripMTgFsUoVEU5cSE4wkFEFo
UkvNv+MgOkyB+vwvZvctvbgZSPcXNPdLq8vNQJexRQik+Dfw56z04vGPJ4Rw4iU7
19qaqOROngSja7uBC16qSnIFdNaKr2VX9fSMButRaX2A9Z62xOj/m0jcHhmPE10f
uGZ4jOUdvOEauS6KRX8/3jkfERBKMvs4bPP7N2oXbViMAcCt29edkO5znFk8hRz/
pSuoNoq/4B1CGq0Nl+uBGXx5DLzkz2R0Teb7iWJyLi3wKOWq2n4mBUrOeOqRRWAT
0djwHQ3+JYR0kcTavIhpe3lCg5UbxQZcW0uIiuMD7FAPS3oGJsHplgTN4yWWe5+f
RDnVjVotHou/hFtNBiqaaqWUOvf+hveXGA5cM6F/uOqezLx2JAnE1tyNjC2lJBxY
JSI/43MTx/BzEidMv+hh8MbzkidJGmP/eYdV4MngkD1btBEN0dXs5/VGStsPvMF7
oFC4xnrqciMnerho3poJnJPu1AhXBgd7btbW4NvAJpQN6T+sSG31sn/qJ6EwEwG7
K2rT8QyOsX7u90In0hNKVDgMxDTsO9VpnkRibC6l4ixRcbsDSY/MvYvpHTk6h7ge
Mupdt47DdcQBV7EVun+f+xwhPI8FZeC5f4eDqkE7XuqzqycP1JBvtuCauIgZaq0N
Rq7r0tZ8WM/aaM4xa4KAv+5CGJo1B6kImGmPttN4o+InJCIpvcFArxjeU88J4570
y2ihH9J//tUDPgEkV5B49Mn8EgNwVVAVDCSrYGtbmgFEwBwhTfCHTdp92yHzr3sC
+TcueppEkjdrUVjzXqat+U4maWjbo47aOyF8sogqViPFDegQtKgfBf0OUUSqO9Wr
bfpx7/i1cojAiyz61RX5xdIfqVwd57N/wgxjc1U228+8B5AMTaf/hs9xOulhB5Tl
uoZ0tdJKYatlWIO095lXheDYgYiun7kJJQ71ElWK68VCqfSncy4YCCtpzHKqRAGO
KY67VYBXPdTVEojwkENq//QKm2t0zXRK9MrZurSiVus3aAhpQWiMf5D6NqytTinW
wmKD/L/rYvsIbiUE9nchEzkzWer8cf0DZ2oxKLNND47tH2ysDKrtu/4QgtAD+1Hv
I3RqDXewIf+P1FqcoG2z5Hc2B8QVEhgQcjtEGTxsW1Unv46v5F/R1vTM2gqe+Ggm
Zw8O6XVKcVP6sh+kgo+bI9yJy37YG3TUM0M3pOVhC8qwD7gTwOKpfTAuXZ3JmOQv
twiZxbaF2KkhOsFjFHUQYnEf5PpnIlEZZodkk2rtVczeLcuySeoAZXsV7CHsOW9y
neRK1g1W8JOJfXd/s6RHNYnkJWXvxkh6AzeUXNzpB62ORQBeSFJR9tzhIwzPZxlP
BsrG5+GjYNOoOQcPEgTdugb+cxuaY0LL0KXez6qfy4uYuZg/SL7gVayMf/NgFCAW
nXHo1VAPzF9+LDNATDHk866u1XGPzKDsElHN0ltEdKoZA+QW1Vyarb1NrZG/Z0uf
TWSIFi/5b/s87OJUaf5kMqNbMQ+kbmALikHzkGwVlpyS1ESoSPOrLl5XevlRBljM
NTS4qCQCBa/r5Dr2rB4u4kQB5avUS4hBpKr5NfU14tkD8+uO2daG9X+H67Aaq7Ir
VXHGBCTHaijqG0jmzc5b4aoQbHC7o8AD+AYzr2B0SYpYZQi/qcez0m+d3/XdnOSQ
ctKr4nLVEpd1gk/qlx2Riyx/uOAw+cPDrvsFpjdil0K3YHEzsz2uajVTEy563KbS
PPuSxuOQsFn4uZ6ZJEEUEOdVtUXoRvzW8eDEiyVfngnjG7xgeZAmiPJ0zng7pgbq
Ul9JGaX7Bu16ocAvLCTNDsim40jJYeLUIsJWmCodQJXHgj1OXvgAT5QsjkZYmjhb
SfVYWr9z2xEQRq59kyjpS4XHl6L/lNI5fqNfSPhm06kd2JfI5fiZhgsz91aRtyYF
20TrzQy0LtkdLMceGyV0L88pgdgaaxglvgAbazhbymtp+lE6chInMeU7fabtaIlh
E4rYy3w5NFSpE5qXUtH7EUgjJU8nBzfuOMDg1WnUm89akGcjQmGOYsqhMJHw2vyk
L210jWmCkrrtOfMdvMua8DubF2NsWL4LMCTxPfAuunrMcjzS5rTrevwmwRuFdqLC
T35/7vPj6HAq1XvcAP/AibKK3ok2+70UoV/9Vij62VkeF0MTe7GecN6Nodwe7dlK
NUnwbyE+xEiLL9ElSowxdMd0ESQiOvSlcSCj6w+VqHDcUVFNUmyQ9ne7LXUYZpaC
sEq5AbG+G4zqyP/aidBv32G2p+zrINANThdw56aA+9FwXXvPFMivdUGuyrlivk+U
cjJyIQw27iBufQlkyx8aJOLHfG9hclYda+9USXc5gjf7qrI5rdoiyNdIqyHCo0cK
yflrkX9CApoXlvoClDPaZR8JsLmVXD6PCl5YQiO+U6XvL/DxS64hb86TqeXqf+Pz
Bc4322nVcQFt+d8Rri/l4/aEjE5Vz0EjbqDit5VjtVAmW2iN25B65ODKfSRHO+x1
uTglqrKTC6yeCXnD0kxxn/atTg6rAQovdYg/Rzh/BM4vdM8ZP3IVsiuqyqX6i2Bt
4FEEBzMolydyVx2wsDooqXxTSmYEXBMZHHrz2GiKiIqhJR+kHbV1ceOTfM5Sm1n5
esI75m/hkk/n6bo3wSypRiW0MkKOdD8djr+Sc1jLARaAETOs15uqW+JNa/Yb5iFu
YYdDJdibtPVFYnWE9xY+Nt7jAJ0cmc0hQHk0142DwftkLC9UwXZcfT2UhIfImx29
lYq9CfmWufJefCGJVexWxzk8qwDOgf3eBPrGPNLEj8WaIZWowlS8mfVWmV2u7cYc
nIKmx4rKCm6jv4+Ah1ylprSxJfVrkm+Ms8vUdrarn9jZlDHfEDBvF0s4DXcYc3JB
X1L15mm5q090cD5IZG6RLun1U6JWRFpaXMkmw97umAp+zrjgttL8r5v57iDHEvCH
uYhB0hooZI0mPDP8O7bVzyD0D54MKf8xuP21AM5P5SpgNjGePIwgoL3IQs8d/K6L
CxvNz/iZGM11nkrEuA4YtY3u/vPJbhIwhQeX28Mr6VHR+zutWn/eHwe4Ob2sGY2E
pdxshiC5f0NnbOwHwQ+39zpaRRlL9v1iTIn3RQUmxPgE2VsweebZVUR2NeG4unjD
krpnl4eHUbxG0bt986mz9AjaJ28RQaO81c4eirWB3hJnnyoHMpeWr5me2PRPBZuH
K91ATgeYEAcuRWXEdSHpMJ5TTsSKwJyi+K3BC3OEqQ2aTmVzB1iDb7m3rpRgxua1
vuczPx/C32jknW4H0ZbdWMOMKTmCzlmChRgwWffqUYVk/YYvrHRapWsdzGDIO8j8
DrPClBWaQTkW3A4SYwGdd0PBK+EMUnvFBv9qwo1GC7yBPiaNgaTfhek0CWDT9kya
dq58KMgpl40Pehzku3N7yyYj4n4A8352zLU7V2rdLs9DZhu0UmdgeSxdliWIqg3/
5gWw1gA0fLQyBJIhwkepBgxIBcbHknUgETZP9w60v6K5xOTi2amzocNCgt5CUEB3
bohXaUSjKAZ6dRZe+sNbT+4V0bziDL54x/3XCBAIai0wGLrSaeVaqzNYUGsms99C
iKsvbkB5q4u4ZShT/06N6RCEsvzRsX/fJbyNJPO4ZuSQqTgId/l0aLy644St8U4g
Lxpe01DUSuN3RUh2Q1mf3SmMdpp/DDrxSQyhw6N2rWQB8qLvilnRgSQlCTKWjJFJ
rQqV/XpNWqLDzMG4A4Ufv5bozLqro2MAsK1eAdceMwtIh74zvjmGeNrHu3ZM04Yg
YE1x4cLHrgZm+o9Pv4D5mwOLo/GWn12ZqQWYjYIczuerhPWJT8skiNS5WRNUQp/J
gYXJvCEtqHyyLK26PrXRF252sfOs/7QEzfBFrLenUf9mk9/iITsrzeYkluci+gEw
MTNzAXO5lC2fjyrUSneT/H1o7tf2RfH1v2rMiWLLIX2RwWqi6YhgPwAQyWGwaIZH
O81J/LQuAqlm0dIybdZm9Dzn5N8YWAsyLwnsFHFr8JABXAN1FxG9FN6d8AbxUwiE
sKUE+o/44PULaN8DDIuyafGuIc9A20Ujal1y/YIrDSNe6USKKlxduig37j0TS8w+
8Efr4qSfLHauUjaQ9TeSW0ruqToo2reL91yKMdekzuwpxo6bTEVDKxEpJIAP0mk7
njIRG6ZqDYIGjK4/UT8ucxj4Tt0VpfVya0eeqqpr9dIkB4Ef3dY3lFyg0xB5A3pX
na4xiedklArNQR2ECg8DShyI31lw5Tyuqh2BFRGSoe9YeKF7Hq9X1jTs0wRtvoIs
KEU9pj2h3rz22NyttByjrKMcy1AZKR3ogHnSHGRoxbS5nZhHb5LPAa9QpssmQkXL
fmn0oXVKLeVQEIecaBJS3p6LgXbtceTHYschObOAd2xNQC6LVeUHOb6WCOhLf+V5
3dSWRiOQBS3P+heUNXx3N9s1HBMsMznk4M++x+AojTys+2q4VyhOlzvhqzwl0Upk
YA4pkyA3gBY5OZaPB/ev/6aePYnQ6cEJW0YvrRqUEpkC6wPj/iS4mZU6bvjPZBQS
1Orf3P+rodVe+eK6801nAC2MjBLWJ/2uL8rt/4VBBAOcR3TfRjyMozAECPqBVvoU
ZkoHmMeJ6SSbcuH/3vQYQPK2UXB+2M3pmkeqb/7RdXwTvx5gRxdxoWeH/gMWFyME
ZweYEKon71s1QPKLg0Hz2r+BWIfKsgPrTiakxDmqQHJjRQtDm1Sc/cbRkOpRawqE
xf2lCMqiEAroetmQVtVYHGpx//XquPkayw6X31qQ8k7ZztiMfJGqyAShm7fRYKC3
rjHaRkt/c0Q1+6GrO1nqOwBN+LJOUQ607j6936J2vy94+OEZ2h/kOc3aDKxGrM4i
g2M31tHwuwbb33QTxWJGZ2BvsNnnCWj/vfn7TuZjBpFmZAL/iMNMol8YhduzUWuo
dDLViq5NVwx56wqZM9jotYvZZWcCx/GbRBTDeaLwPPl+uxqzLHNT6U8Pd9FhA9U8
8lZHLVS3aY5tn+TIBMqHJneXqvMhakz64zMhA72kExLvi1DcLwKutQmqeJ2zOFk6
2eqx36rUnoNcupWBzhEOs9fLhv+Jw604FkVcdYNYdFqylhXVsnK3e8onOmNO3M/j
HKb+Y5ffHdizwoa1zajC/0rRYY3NHKw6+D3yQGqKidF4yowakGvvWH4o3R4wDX+x
Ybgwr+M4mxYVeJ5EnuK1xMv0LZQRq56JW8l5KpR3o+sMOz0k5DdAzH82ohYTKb5y
JdUnY3e+6CT5baOsKkzQb0NHTs+bhJDEukD60kGaR+xJvKy8H7wXNnkR9ltQ3F1H
QLmm9pRcPYX88SuO28MW7Rw/JcjKPn+iBAgtBDhDs88iHTSfGeDvl2nkHG+ZJEBg
9TycXjULbX5wclJ+5676hq17oNUTmdNpW3VC20qV5vMdss8O4T9KCGSDTuNDMyCS
83srJz+hNRBf6anMY2PDITDyD1DHSguijsN6yMNmm7BiApFTVZioQMiOST05JU3g
l0Jy2uBxz1niXgNsYUu24mgwtAxOYEsE/+gWMSTW9xhgU+Y/4unQonEDgPqEa0R9
R6jIeYNnjR+R0Wgp9a9UL+BihJsLVoUQ0ESXUnrOSBQ9cApx5vssOM4fxUCiGTbG
DmhQ8zxZB795R1d7DCIqOhbGMqMP0+gmq9utL1y5MF4uvLteIt+/78r+UpKQIN1j
Y9KDeyu9nLbS5slC0gzy7I+1iZmsyrvl2PdtVZH68kX++CKo2ThWkQ9x4n0Mlz6A
R98ApRy/S1WIC8H6rYZLITkpZAaQyOa2tXs+9iJWQNIOPjYjd5MWi+qeobULVixC
RQPPyHVQU1pig7aFd2IimwfXLRWiGRzd8oaHopg+LaEUU94Q3G+2jh2p7ZgrBUWw
wUkI8VOkRUeiS8dNXzyIW6RiqlKUulqFCFW3xvpeiKbJDRm6FV9FXdJI/dFzuu0W
p0MWCcBbit2bgS4hrcdhUK6dKKMklOOa6TprdaFcxgBTtPzqZPy4AQlFnEAk0hw3
idhox0ePlODcm7a+8zFKZNL3DOTx28JFPLMtI70tcfi97bOwY3Rv7tfk6SlFXmJq
jd/7lT1ozBrArzBbtXdVOCxBRQNlEHq6+KWeLdEOpgqjUYytk/rabA7GNoLUF7Q/
T6wtXfBGRaP7VeWY/8eHcYAclreNWe2CR62nx4wgdW8eqFcxK3Eki/yl+WZ3ensx
CI8NdBuv5h3NduxVBjFzDTOyegbcTQxJSbAJIo4EqeNK2axL86OnAOEOwN22MocC
UNQHtHaWWobqdzHZDt8sQOo6M+muLtrksXTtMwrCzP1hCfg7sffzeLTnrP91Xg1Q
B0mrPvCt0avZq4vVjQ51bQD+HMIhTgs+f6EX/QVCN5JtB/BGZcPGLHjpufL8eWWT
7t65aOvmkMy4EvvZ1RKv1rwv/mVzm6LUxeIUYxnTpKsSV2RYVoI5zTfypCMvUN26
dft0MavidLvLoG/kB4kWHaytF25qHfcr8ETG0y1aK+bQK1RSbdYGFdAnC90/oZDj
JHOA1nv3bOvXpr8xy3+VM2DCbtaDcwpV5L/5/AS4diJmRwUVhKH2CiyPX+KIGGjM
+N+Xq7zlFXktoSlxWMYQq+L5d22n9UsbW1jIXv9BRs4xKzcAlwBhrHdu0+q/jQwc
9XO50LUPIIkf7ib3YOGu6JyA/JxnKKIrhJra5mvWH67VybFPnkYCaMlm4bfhniD5
zWfQAixhfKeKlMeD3V6Wro/9Dg1vtyxfo/6TUjcckSi+spuq0uZ24jKQI1ZQcfZz
ET4XSutj+vhJhTyxaAKkM3VZK/e/YtVOzpcGQYtyosIJqZ0muFiIOw2MPHn19NTf
kh/m9j4kdrNKAN/Iv2goWuYNjDGb4rS8c7w0p54EW0y/Gep2y20+G8WQIT/fyVD2
UgLudhwye4ecUi0lDPI09Rtuk0pfhL8yWMZ7HnXWvDUGhdXfajj8oEoePWw1zm4k
LNmbgPZFwN97z0b1v86d3AvRPA/rCwGdtGoOc86UBww+iAoAdPsouYUavZiVKt8I
qPmwrS4+GhGgvWtlDd49ybdTXg35L95gVTuprvuro2NSFkHrbhunBLu9jykS7rxI
7/1wvIFpqSz3987gprUqTmqhSRSM8RyI34E8pl15jNLHVAUFIgFpYJyCGbCpBSfQ
vPNClI1W2nDpXaEsXZZA8HBWseuY4ujSX54HVkMwTwl+Deb16eBQIhqj7irPtLm4
t3hmS/tViUCgh0LN41x96QgAi641g1hIdIJ1Cm6jUMUHC+YLk/wqq6mbfN05uGGX
/W77IOUDE14Kx1nB1azESP70fKDQSlVGNTazUZV+S58zmQ3vIXeJDkpaZP8oFzb5
DdRtYgcGLzHYJaJdz4ntFna9U9xztPWNwVq7TLn2Tx9YXepObB9DhZ9u2g5aVXhX
F+56BKmn+sWQd3EkjR/USRBhPpOW4Ro3Ro3fVUNq4bZWqhdn7YuWM6Hnul7I7FCD
7X2ZJXX5Zhbg3C66A+L5NtWsgDGQmbr+aGg8HTyeGkjzeUGg4kWaLLsprd3URiP6
GMWntf+iK/qbl69HwKhaVgN5Bdx+e+B6Vbu/ciT+As3dW5W701CeYxX22iLLts2/
ecDgLCeQ1+zxJC86hCM1FJQy7/89XKIPFt8of5tkzfHcLcqMLrJYO637mcW065gj
Pe3NGcaIBUEPAcVgSHQ0L0/bFnzVXsUwtMnnG0qeYqK0LC4lNr/vV5fiFikOiInF
7+fmBw4KqFABtFDFSzwyXSpabiZyDgERbz2Kl+vsZ2526bvBEkavPT+fyS71u5js
3t7JfCLJqsGLadBRHAlC4nxlYuPQr7PM1LKebiKq6hae6gSxDkzeZFOk4L2wXjoe
FlsEHWN3UTfawHRadOKTotGXJQp3+A2w51Mmbd9CjJZlLkh+8SVS1pd2pEvdZ1Iv
PaLK9hIw1UWBPQPMmn0OTm73HlROeJESGbL/JGtYapLo7Y8sf9FaTI6RoNKNdAE/
ZbQoDbzTGIxPhas4PTPkMrEeJXQCUxyGPLCjv4SSRmA8EMAyobRWnU7Jbt2U2Y5F
bbOznToqeEaM8OyZUKdGjSBD4510JhOdWKKHKSijcqpBi7dfPApSBNwISlygQJtQ
SYO4sXkxhX1gL/0/4DoUFU+xfSxJHCmU6+co7spdVTx02pge8xNUej5itjmaNtTD
Ju9uCfy/W6L4xQtffxCO/Mbfau9s8hFGDfK8I0cTZF3IxwkhZ/VkQnLPUcZqDdTa
WjIkI3eLHCekTSkeqFEoguS5lp6zFp3smwsXHxp/PLP3rqk7AxkX6fEcUvnOM6IZ
6g3aHdzFl0GjLgL/73FDZG2TPEtSoeWSZXQsRAJjFiT6D+ZbRsCB6Ruznf/ltYXp
VUx5G3hb0lBh/Cswhe99DK4Eldhjr4aevh2JVdzF/wyp9kMbd5NT60Cezl1Q2RD3
IqIg6KNzwIJD6NI360GSAyn/ALucuWBJ9qV0NnWB/3UOmMsM2N7oQE5fcdFME8pg
FMhnio52M+k9mAsiBeVnAvZEtWzKZ7m1SY9LdsESpQiHEwT4ekWI1i2n28cF8NwV
+AZPEsZvVzKe1vg6BxYqz86Ec9Y9DHTooa01CGbob1OcaSClebsilBPLOUDvMlZE
l2PfO9KgFKT3Ra4bJdPzDILSw+RljWlhA8p8BR8S5LK0sO9xiNs3A757afjcgiHm
x2aA16bDhCH3nv4NhGMaBrTOAX7vL85iY1gT7tAIFEiWyqbeqb7U0Wfbtv/OwM0l
bBsJt5TQQGqdtbbBhSolk4y/gocjV200vhXL4eZOg1aU3Hs5D34tF/067EIUklQk
4yKG24oeCWTEWGvQLuLR82xJIQcIX/JC9DOxR9gsE/vrAC3zAAn0sZLJcGHrYprh
0AYFC/H4eNG0u6/j3uN33nhm0TAOt3reBIYk9M0d661x6Xs86IT41P5rMNCEKjAZ
KdEfswi+WMBfcvSPzgXStNOg1pDVRRmnYtMoJ/rW1375tdse4jECskRvmwbQaEAV
xrgyA8TV3INcnaiXBkMlxpZNbmODawGiDsUmIaFNKLngIaQ5AjRkd25FM/I7ye7T
frlsflsTnv0WDvr78U5p3qgch4uccngXPosymH4/001XpNz4IRlM0vcrmolvDryp
UTPUW2aoWxUnG468iDzxJ/tZ1J4GYDBZOiGXxbEd/lf5qv7TQJ3XPK2KLlH/aYx1
EQSVfjP5UAuFutJHcxZCDZTzkzdCa9xEejrYl8KgRnqnNPMBn+ytBkkjaNa92C+V
Cs6GSLcWqRoRIRXzTV93CyTSgm6iuAcQNnQEhy8lusSUI9rjXm7P2OZoTDlYTk6u
VIL5lGVF4eeM7gjnFRHgDtNGQTyi4KxGvsZsDnxjz9DV/2bm+PExPc9ChrS5owH2
h2J4sjzt9PJMQm3gW20wlIsmroLyGCi36QqEopuQIR653UqwD5r/ztXetynsjhKe
Cr1LGtZhcaV/MSqqH6HvacChezR0FOOv+FsEf7tFPFt5sDWHH3IoNoHtvCsSvoLd
29uylfC+qrSCFgYIKFKhqZFz8tcrTPea3Bsl/NeSm27ZRIYkReI42a0DQO0EPVg0
biIo+yOonAGIlJrdH1EVXcn/pFcaW4elISCD8REih1ONqBong59nQJA8x/8RN3dp
YoyIOx5HxANb9vpYOMIQweocjBuNyB5YnO/i0EhsKB7HMBtSXVT/rJop1nu51mF5
kkchf3Da9vNlM9sU1zXwKZHistfn8NCkgL0PCeJQEJHd4kvQi/9Hgf7Axtm8J339
gIi6kzYHQyI5fS2S4dCwQReyHEiNGEqJLla8Ckqx7STFKM1uB4tmLO3xM6GpoKog
4iVozhK2+ONXkaJ9UxNr03x/R6SfIZsGFvwCqP263Lc9DNu6isTB6K1qIywhfGqV
6w8TCmiaPDmm2FwA43wd7KpfZZl7oG3BqvXdHrleW5agbZvBk2WYbddAO5qFlExw
`protect END_PROTECTED
