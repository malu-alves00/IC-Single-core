`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yYQcnG+sRCzN99Kj2Lz2RFL4FgGuXyRM9LrferLcdu36Jka1L4yu+C3ab97uIuec
pkGy5EQTkJ0FqNRBfXAx0qOvWmrQrTeN03INb9/AlIIuTTmgK6oMDvMHd8TM6ECi
9jnZPX/RJj7y8OHwL8XajMDlJJ2f7b0DoN7TqcLcRsejjoPVDqJ5BUNhU7BJD9nc
fW1rH5kp0dcoDw/QWJ5LrDkRPjXsOXn6ZCpNdO1Lmded5GtMTC5R5N09Z3RCMawa
/BJlNC+BfRk//kCgK4FbtaAuS4OTKDgvUUI3l739Grcv7DGiwjQQEIuyfkgU1d0g
zH4WItNdnsxw8vUoROIR4hAGbYAXFP4o1oNyOFQ3pp9nNiHuUUnAReBaAuifkCuA
dh2+ddqUf7oJ59KIhxXaKiRTS9phENasCADiIz7PmerE9rYlBlNArcdECvHk0I4U
0gLo+ANrO7vMCDbzHTzyfexdG5oVtiMQIDNv4YYg3JgAqKJDqKjZtyZ8o66aprAa
/FgecjYZS8GZB8fe6lGraeIWZfot+6Qq3eHA09Gz4V1wDRE2BdUA57TcTUDNuE1k
eFmyf/w3KtkswRIg74efElmyzSqXMaAGXH0jlR4VSnl9Y99IuFk8bnjgxw3v2yUx
L50MDGYhYn6ygKnBhoPdC7uDdWH4ds/fX1NOE31lW846fklWNUvMoJuXGYtqOf8b
cMZ7LiTYQUqKBIfuMAvemkrufE+nhc+4zMOMWc3cAf9kC/+CjA06N5AhCnXFP4yh
Z7GNP0CmyqDCFsOEzZsjEr+tE+4dVoSC7JdednO77H/RoaQ0w1ZMDL3Kg+no6F0b
M0WqPwDLJtAH4dkjEXFk4L/Ep9DLm4ddaU/5BXfm96exdEKm68OLQCCZG/QuJwph
xNUqyywpKNmngCJ4Ptfg9uhbj4dv0RVVN4ckLr+aCtHizWFLV624qyzPGH4z7mBP
KGPoYP7k+ZhYJQkQWyuY3hBINyJLhpKxSsE2MF+Kmw9OHjEAekL3jZkNH7MiFdnI
ZNjemV8ew9+/utzeKusocNoKrjRlyJiCiSNQGSxOuX1K8e0+Ys2LlZftBBx7Ce5u
uu2eOfUQLa7WLqZ7dEd7yeL0ORTJ/VALdn82d0r4hzY6ffWCmysKueGjy+mEqqfS
LgguJDOKw07jEWShGm/i4ptpG6wkRI9x3U9+efXQ8GAlS6GrE+V6xDqHq99fHxJ/
WS5lTQm7TxMRAwGA4TKvfJ8NPzfnpRxdnDuV3k+4mGWaC22h1EyB9gB6rUzvvGyy
Jf3vvvfWAZ2soQB7Rcb9bvJS3dsaGA840/9s8Ef1do5b5VjLeMqzJy7pjPEppzG8
RfaYNL/oKDqZjglEhp20SxEAN3cA/0qln1h7TOm1f63p3hFbfuvUpauzYfnOqAxs
oxwHV8sZDPj4MEG/qXuo4D22vo6NuaSlEirCjU28I/v77qDooRAjfz3K0B29i8bP
v15zFktPuOrt3GWGGkfCmBBfGndO/PCxba+/JIMeAe7jzpEFVXmO+adFCFlYSmv+
iyBhmnCNXmZjCtWWjqhEtN5ZZZalOgkr90OoSCYVb9ZZcrQGGyfJKGguHChW+d9h
IBHUzv13sHl+MbOApzwGT95XyE9LH9zfaKuH30JMaOLovWSXAS7UEl3/aWER16H8
zozxmDovjLCW+g7r0Tl9Yw==
`protect END_PROTECTED
