`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
73biBCEM239AcGCG+D0pVXqxNASuHGMRVTh56+q7H+/ktfjxbIjlQ09RjDAD+78j
NRauVnYjkmyJNoJimLjIO2LVSPlon5PvTAsdck8g3MQts2FCl4xM1upTAlCSdWgr
9EBKPwoNiWwduThFv4ESA2MmzOOpBF5Q7kqQv/32+BEfzgDuOfllMQJAh8oUXqxf
x7C07eY9SRtJSvZXcgUmkmbddyG7e7S3lydekYeAetVV/F2+zrqGA1SWRP4TwBiX
e2qjO10wwcSoHAx55/iagr0ucFM9dsjLK7fnI+Ba+wF/Y4tf9+a7dfa6JxNToBBC
1rjLybvPkvLekJIxYqJESlSpZXP9hfKXBhnpIzOHPqsddhCNxv22L61GJm3UTm9T
wnLqndBy2Fyhn/ZHvLpg/yVwzM+tK98r7Mnt502GlrqQ1guikz9yqeEEdgTLKO6f
PX6n7P/ihvjPXTF3LG4I1Gnwi+SVAjEG+jtixPQ15x6SSRm/+oKJoHoYYJIa9sWN
qgy8n36qvhouvGJFTbrFVw9wojM/IfDSssZVhmLoJWwgtYYqoYNiUqVw25UVWcDf
vm+DDZgDEjhR6WRLVC0f2rrz7mO2bmd1yVxKyY79zWRV4gqFrNojh5dbjRkWz+Fx
`protect END_PROTECTED
