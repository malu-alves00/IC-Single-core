`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dDNfxFHXPr7jiTiVSVbPEu7e3fdb8Bxv5N8X+/5XHmLNfMpHRkyH/e456+LMnMU3
bz4i1vdDs3gIaJUcwuzhN3Er2iLv7t2o6kxjb0Rk/bo6dvJNfjjPTrn8dTQjb50Z
ndCNnh6AYwPBUvncDCgVSVpU+YeDERPRWW8li8NgZmsTEofp8hHycQiOp8pOtYHJ
+Vfskt9D7TMyWpbezpK8MPJWvUADhlAnLs2XT9EM1TOQhbZqnuZSOGVJURbMK/6U
5d+OPpWzGiFooDKomUeb4xTeHzqc9Z4dxtbdHGtbLUh3sMcZCyWLNAVoYzuOM5zD
ufx/nIbQGNBjXawmsoMws5//1PxrlMnMIu/iiU8ZmwNKe2hBe0Oj/d4vQm07wCO7
ljwe0vy0A63li3zgBdzi3/IPRztdgnHfNHkxmYWX7WnP4STKPV3gj+sWXnuY6Q68
PULelhzCxT8Qa10aglCVcxMSYjR0NETIWiWnKOGpjWc=
`protect END_PROTECTED
