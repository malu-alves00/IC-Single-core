`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Lit1TA1A8CnGw8tm0nhI3FgozXurMY8Ts6TxMjtBrZovLQnxRxLxNabOAj3+Nijk
fLoPCb/8eV/8peBc2kA0oQqugJCCeWlCgP6XTHSv7OZKgtPd+S4OPfM0sGH2icZH
dBrZ7aQzyAQRQSUpN4b5JhM+2nLMmXOyNd2NTYxEQcDm0xtQBXdTEzATX7I/eTp0
msyfumlwS2Qan8QU48OK4WsLSOUIOWFN/7sgQDSSogqgP2RaXUjVE1UByuSfvgeY
3v9aFavKmYixgLcLjA63E8yCBBcwnn6LXAW8GsmbfU4YoRteF4rfLBeb8bLywQvT
u/7Bg3TpJjtae4T8TOCaQ8zpPbq9gizeV/T1zOYW8DQx+fX9E6Mjuiqob0DaSuEm
1BWOU4btiWx67LTc0/+U+N25KgGxt0/Mwu+gXFoxeCFbc2rG+YEeguJHwqWgW0oB
VeRWXcyExOzyrVjtfE+2f4J/g2AQiiIhP/rGPfC2TuFtLMG237e484zaqiiFmAY0
DJcBFBmmAy1OKNdcmnJTiSs81nfzq4x7CCbjMOJf6RM/hFV/8rg6Yit9ddiZu9Oh
GRiVSQYSOPqvwpx7mOz32A==
`protect END_PROTECTED
