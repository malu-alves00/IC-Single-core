`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
f4dywFudkbeM5XscpzYxHWhSLk8Bc9FAIUYqP6/YtZu8JRODK9ESfXkQJLbfamWq
lgtUI7+0/4/TeuIDQgZGPhKqQKQ8cLb3/U5pgSWfHpCKmKvjOeNUJhh+vHWCB67D
HJlsnqQlmPL2B9NDJe10ymtPnsgrGX90EDDHYbPDVT2kdooo9b5jthsq07wEQZln
4X7BTr8LYwe/RIhn17i9x0CaaNvGErDNDQ04d6MELARiu+k/EVOroxU6jw4ulCtc
VLyLWNcN++myVnBXLvvdxNAN+ZkNSeG5dMMMq20Bsg09xzCyB9MWiEJa/Nxds8so
3JeblMVvdLwfmMBfMkU91v3n1fYMXCeTU/eba5dJbpns3nRXyPIeuOWlzoLEokqr
R4MkpXhYrmDwyfXLeCPYUSTUiZjV8NJ5wc4YJyNu2ZDW+JClMkEc4KOC5iN9i/Du
03OmXAayRL5fBqASmFEn3OV9Hss9OIsu6CJtbeqkKgCPkN/CEAJxD1nmUF5KnHVL
qJaOZYkZ6MOsFx6hgXvoy/rToV7AkgBrdGp3EH2d6UFVQyObO/vrVBlWWZ1qjnbs
iXFwxDHgy4j3Cvtnvi5T6oEuOYTgWGph0rl6n9dlc5c=
`protect END_PROTECTED
