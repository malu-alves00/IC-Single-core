`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GrRZ8bIbPK5FatCltHtbMF79i6fA3Vt7u9Ht7bw6c9/U/oD7/0otIC9E8DbiGcr6
E4RlQE0SKE47V0kvEzmyd59W06yiTDTshGV5nFSpGxymXNuPDibyREIbIYfmFUAM
gNh+0XjoDOiHHzimlBjYJEIJSUVKuZOlF9X4canXJ8kvhaKKJ+i3v+MNjpR9e2ne
c/hrwlLiXJDk+VEm/7vVLD8Ab2I35IwlQLtXOj5iOLrDMqM7tgYgrIR5gE/2Siv3
9EootSFgL4gWyebrv23JhQi8pAK9aOL70EKMv5JVEqkTjeNyMIEzD5/ILQGhuHV8
tNml5rBgDk5BsWh3f5PG0Wdr/usPvV1oXjbhLCDM/uMuEh89ZDk3cfH4kfzMslAX
j3nCIa94053LJ6bElF8WMtbjeTFmfR7jBgaciprAx44FKT55Fri2OOV1R+yjefhu
7FT5SCNh4filQrIIbXzf1G56c/gwgL1KVRQaPfaVuQdSXUqZk5tJ94D3SdC3Anfn
JcXf1j3Bw7VTD+Evxs0ABwwbmXZcNcnIQAMgc10hm7S8UVlaHPSlBmtCEwbk7cyK
+0mgDyv8ZBnwgOAjXixv8MUMjHIszzZ4nQ3yx/B6MztAPlEfh1wOo1AX6LFFfv3r
4fwIh65vvpk7lfTZCYR49gLI/7j7vcceJQriz4ZBumKZ4D2GtkDoFbliuovkyQ/Z
3QZHR/5V2Y30QCtCjU1RRiKSS+xYiS0/J/86JcTSsyVYhbGJnXJdRN/hqbabdHwj
`protect END_PROTECTED
