`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TdFHfJcVWhThf6jN5+y7lUNIBuk3uQXdDFwmeE21ahh2X5bD5huo9/U3KjrjAwOB
9Z2fMbZRNCh9gzRIbIv6futgaA9L5hdgCL19PIjsn3OT3GsUpQ/dkahypHxsmYpR
gOCNkJplDukn7tGku1mzI+dRsatPjAjSTjXstPJX5XhIZvaK5+YQpNZ9NwNRXJNL
ZwNiNfnoKEmGKNXXRKnEwYvYexfjL/J2XbUZf37ZE2mduWGVEqOlbdKIs4TFJ4+i
K6oX2v1yZQVDNm7jj7YNdyRwoGLCycc94VbcG5EoEnPLK6IVphSAquuEWETOcrBc
fF392m1uI2kjBOVdwNS2rMJl+8NsNXhzGL6q1IJvQQ1xdYJkHtl57ch80hSFl6Ff
NCpah+6Etq3YKgEJ66xOimfmvE2QlivAwvN0H213L+XudoRxYS76K9TXctmGofbS
Zg+nVCSk8oo6UyTSbJHA7s8NS2G4YLKlgpoOSwpNqnFWvdTJ0PYGgUqMDxYx7z4G
7bgyTqxviZqRo/5BnGbjVZs8UJ/+fX8YESockqwce2z3v9CBMN7c/Is1W6jXg3qf
6jgwrI6yWFKLKm/lKipPSAnFOTHH3h3n9fJJUdbnV7Lyjagmbk7hD9cVkXHzf1VI
vjJqQyM0MkNh+4KTYwy46GIpPhJT6SQ/dbNREs0jinOZa2p7FcBpvQXSC4cbVtZv
l7tGpTzAqSIG3oSQFF+gYi+/WfpwzXjyQd/n6JWPuW1RP+B8soWhJQj8sVc7vQG9
hFUI8XEAD+kawGf8aqS8xUYGgahtKhOhLTe+qWHPW6Vlzq9xUqDQPW/V6R9qll98
DHZJUJWO7m/+kY0MfMNlxY41lrp3FOw82FtgsPtZZo4ksI44xlLucmdb8w3kMgwg
LBjz9jUuTY403qYD6qCOgrdU4O/htAxUZ6YIhI0r76JLG9Ei7TF/coVGpUMXzvot
A5sPEkxJkGV06jLMWjsq6BcSC9pu5Gwip/lFHqd/pj+CfjUyxlNn/K8B7Zer34tv
gc1g/HrBfXL2v9CEOtY3Ahqg9XlyTUrM8k0/blMvCWkbXHkj1mr/bw4ReE4OuRAs
dnRViQBw8iZCSL0MTwywiAZhVSeREV1TIDBOMgY1pVw337cjzOuuzk8myZwphd2T
u35GaMdNDR2gUTSR9oaWbe//dNSl9QmJ9wcd39biJtQ0Ya3ihHLeNFwuzW4ZhYU9
D8/VI4DBFMSsiootuRJFc5l+alqkfTrWXCB0q++VzwC+b3a+sfAisL2i4eAXEyJa
ZgPvvFBBu110VEiKnoM/FsnzW6isWtFpw89nXWwyU28VEAfeDqAxM1137zwGtjpd
qae9x5Z/nfg4ngPPmJwBq6131Nln+e0upHt/z3oiUSS1Ubnqe4YyiT3SOo4PwI9e
O/htigB7OI+Zrok1v23BkA0gNFzWReJhd90vCR+AeCJ+F2WfqHjI+Jay6w0CaCx4
1xSZHN179f3+C7SMDDVpcO/ESv9nzPKlFNDQ+/jzGsxAAiV4d77sPAe9FXc1xjfj
Q/NI7t29BEoQsRR/QEsLWrENqocgIAMJAetRIME3unr7xpfnIaG1QU4WBefAxJCG
2SM2oZwoS2wcnxO49o374f8sOq13RfDeHekYBrq2TCT0dm2lvlrnloRYLvIAAsY7
yDTex+fHiBJvgqMuI7PYDYPewLNYo5nWV74wgXVmksE+Kwhy/r3y+mIC/II5yJ8v
Y1SB4LEgyuj/z0a9Iw5lVsN5A24rnGpt8wy0+KrcqsUd7s69DqfqGjHzl4glaQp3
/VeY9/ba5ZitXBUBDv65mJWTpQ+2bkKf3ooNCyBRc32MKwtgBDVgHBBw47rSpyMa
uD4QZtDDVG8GZ7TTM3R9t3nRfqXZRI9WcgdEMe1e3J1WaR8cIUEXpSbkVtmwbVvG
zemEhJExpdn66IxeZOhHRNOyyVaRuiQKbHIYFxecD9M3MUxsuPZfdTKpnxLEbBTo
hNnVnHfrlxNwNvnffd18kxuwQAsdCKhuAfyBkBcu0bxNGpB3i1JzCZ8DETbTfoCO
TpObLFtO0ks8oRXOJ9USh860RbT99R3gx5lR26/+Q4FLukHrs3D8ucUoNsTZCKcH
Fr9lWsfkc2kziJkkpDm4rXc/zdMkbYjudkVu0ixV1aexLWxamUp3fYZu62AP7GvW
2jVkQARlB9vObfUpJeUeZgE+sZQLgZdm11Qe8NRBPPPFnNBKyNmokBWrPWUZJgJJ
sdvEGBgvWxrzjhHyVecGojxsBthIpyN89tmGwNykV6s8npVwhd6ycBC1U6vizCBT
skf8CFyCKmnwFQW0Zwr89PyOCQ133EGaAtYQGF4yITnv7SEoUvoHeSJh/VXXeaZM
wwbmDwh6lqvlTee/deE4NZ85Y9vrcuIxaAvB1ed9XEd+6K//TZ3H86EEYisguguJ
85vIxxXAOHYcJLeeXhCykw==
`protect END_PROTECTED
