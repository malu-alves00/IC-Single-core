`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ix+HIFrIaA6yM7pIB70MpIBlUgk+WsN/ShQG8MRQZ4+tASLL0M9m3AGOMyMa2tHp
Qe8pOYaBiAaNFk0iz87IEDcl8HUeTZxvkm9VlHsc6FWTx1LBDj/Qx5KgjadE5qhw
Y+ZZTOkkEAGZkXfDpNJnv8jcKXNqgAi1xvNt+HTlEhDoW8wRfwZkwXGZkZ9GtDqc
b7Nv5U7KPZXYFaX8BSzcsANoJW+81rOFH/mIny5b8DXUvGdnJt6OffG9YXw3A7Kp
kj+8gr7q1ty4n0WImn8UDwaXZONFxVtBKAScikretjt0wzmVxV7v39FoiNvzsdqt
QFxY3Gz1exOKq7lf1MTObRHzev2fGf2fS2HnE9hAWp5hcDfBgNUBIw3drC7WhUq4
awiA7xxv1yzCVEhtte3SXjyn2tHh17mx9MkaXr9TZqxVn9R3S3fKcTzhuhTIO1xM
w7wiwid2JGwdxyCAd6JiCCdQS9mdgDBFhPYnuWCavVi4OiDsvw/3x+ivFpEIfBdV
zziCQvqvONu6WC5tmssqpIGUDoSJFqg+s4uwyHQqGfnFYHcVSnBULh6ZG/cpx3sm
Acm7VLlInVtzfMNpKAocBjWncCA5WEuv9X1YWxmS0asN9opMIB0WYNJqmbOb+/Fo
tSCkLXsXR81QjktqiOXq1vTPNVaV4eSY7GWez54XxUU18vZX45AOjI8AC3zsrwFf
Ne80eDlGDK25NuiYl/eMrF4HdqN0nh3JvQsK92efytIH43ACzR+updOfMGriBsuW
bxnvfi18FcdxRU7ppCbUpLvW8yDi363R6hHiAw+i9MXGf3hdgV/myQzg+VfVPi1s
FtzT17sAROIzjw19AOc1lsKqL2+VxD6/DroiK53NaRTzeQBVGweYUceDbqlEYtXC
rQP6yh5U4z+IjgaD6HWYaPDE3+XqQzauGsi1WcETZzrLq5JueKbpvgkScmD0idbA
MDV85/4aPQmudqNRiCZRk0ueVaVkEYWJ4442z9G+HR+mIPwQ8qbqTNyyU1oIw85e
POYr0zk7ZeO3Nusc4T6ElVM7KL6sBm7Daq2+SzPd6Sb4h9UYhZey03iItCj9uz4a
tQ/yNalPlywaIHYzmjE/HGV2t5XgIuvJf0q5OPj44NWVdjflJtiJALaS5xNu+QG2
YSTpDrR07P1WIv/mMi79TDHTuw0/DqTQ2eL/c8uwd5QgWozREzSUurIJg4Q6e/+D
I+vEUW7cL4eJ6q6Cz/lOc+Vg15Ulg6tpUzDtO6l2Xw63x7qycc4eW1gujp59wGNY
wDn/PevIGEgvGwtW094toI0E0vB58R6zFJAxT6S/dUSKmOhhoWcy85615WVuvfWj
SG+nZxXpA9B9CeYbn/P3asBGxGPz7s6/bc35is8SRSKXpAKxsZs47vwr8tCOFSO+
fk1gDJVoGc3X7tekNVhX6N7GlRqDzf8RKMRPfBB1OQCt/1CFl+u5Oh26LhumuKt+
f5u2iz6AXEE0OPgcRhP2yoPVggZtQ1rzL37K0eyiXEf+8b2rY1LZcTOtcT+v9Q4O
qPIC01obqpSV/kTjDNp+JNL28nuluRU3S3M/i1Pvwv4HfqrIzapX4JNK23sl3vO4
uqX2aQlJhr7tLWRlfiYrAuGt8yQyHVlsFGTCa1vV08jqiab3d531+oINhM5o9lsv
9ArqoxyEAQ87DUFWTTZLVosfeXAZIQXKq6fpivM3ybvdqMyhrIZ40n+cx9RhAu6E
CENHGjfthlTrojrF9iuFMEHUBg54zl338xG3Lz9maNivARnBtQkPMJ3Y6EZcPds9
Fai2n/OF/5pqCEuzPZswzQQB0YbiWgJIMDRD3RvC3YRtX7MxlE2kirDPUW9KhpDu
YPt63jtYP5o5x3b+BF4YS6sMKQJYdO8NUu2hqjrXx05knDUqbFHfUzEFL581g2Zn
ibpR9kxuMFEAYntlweVXGmgMs4Q+N1iNF0W+iMso68n+PDmjXElx0khPGrH1YmtL
bDKc7ysrStnoV3K+srMKPAYCFwciHRzajJ0EzGcRncg2AtuaHPHZpyRGYSXQe/QD
8RZ0Lu2xhufqlQdhtVx8LMYc3nYkQvFt9YyOGJ9jpop+OjklZXMRBBJHG7TlJM3T
H2KOfOqmqho/DBszf0PR68/SzOhzRoNsT4Z1OTbEdE5px8G4YdqQ/s6XCkiNGWUt
toqYGdZBU4XoHyObokLQXNBG6PHYLuN8wGc7Wwh+Us8tjpcM0IO8ebmh5VkCNQ1Q
0vDnZkY+GwW49xTbyS9Nyk7Dd5upRc0fzTmRQ7l427kmlHUhAI55R9iV+XtUmWoi
2Vjs+6l39E8o5RjliXIXNbkhcE25aBjT0WKG7CIhZgi/CqgqwVKfxCBiJGl+wXr0
qfMh1J7mp6OBuXCSEu9/d0TfBLxk9NJbdze3h0zgLF+XJuJYP3sZxD/grIDh/l+C
kDSJUWX8d+ZdnZzra0rKG7fBnfQ/EatJJjobj8CL8jZo6FaAyyngVyQDYAC+Xxp7
6wyKSAtaX2cxdGQeMsXYPEf6U+wIb7Zr41QVVzA3csH+OOXSlNHi6UW1iYDWNz8h
Xpm4p5+iUd5qVLDdHOs2HuUXDN/Iy+sk0AHEsVRmMxDLEwqrmmUeKEuuWDhvUncc
GAfSc8ykJB2kQghsh+yRNUQ47F6aTcMnjxIYb6pa3v09HWq8Wq9q52KqS3LYppGL
8KgzFXntw5dYOiCx+H3TMnieTnydpkT5HrlM5tyeO9wBmCgd+4skkgf/UfnhiYHy
jnpFu/4icvhS86C37zFVQWL8KGcL0LyDnanuWqeZ8VhY2vwrAxIpYVlRJogxDb5R
r36kMMVPvSig7zAaqruvwUlO9JAwLHJ3luBXQZ0Z7+ZBBgj7MJxzqr3RU6pkSnBu
WxWs7eJ8teI5LHzdZwk0b3Pzw5qL1kKOvlhGAdH4QxQNE4AeBevWmiLqEAEYPqHm
K4MYo19F+3WVy+LbbYHDK6I69fAMLczB4CiqS/fz952MSjTgWZF2fqUd7OBXCb0C
wLh5hIVzD+s9zloH4UuVysXKP4QsIoxai/9xEdoARm1TYLcqwVaMLoEGdi8hIAGl
R8ONLHbmp6uCg32W0W+tNNMQlc//UpuiAj2R7nxMJ3RTBaCLTQUYFjGn26pAjJ2M
yuupv1JVNr81q+EoO4EJER3UiCqICCB2l+8CV+/N4rsIuPho7AE+UzUXUAYOG+xr
bhkgxXboH+uYmDXubOWPvFDFf22FiTGIJjLXcgDWQiPjQzSM47N1GL0Z2+zrljio
wx/rcrIi3jPkAe8PtkyUvIpPb5ubNXWYlo/FHK/7pMrJCZJixCDwy445jzG0CIEa
HHS8188j3/ybrVfc5XC2jDzpSZ/FIuoAZar2lTsgIZ8I+M6lcN320TupEj/HeD4q
QJLZCxBPjbkxZZNtetVaMD1v3Hf5D+KPkO/YxrF2gSsqHyxfWNng2UFhXJFVh62t
ZeoIyxNajbDGb0+px28v/JrMmIqvVvQvN4kDY2jWKz7ihIFQGyPMY43MJDsa7zln
6WMq3q4WKoBfu/ZNO5G8ziaxK3fx+WfhhkaaXs2C26Q+fA97zvF6sC6BOUkqD2nG
2RlQSP6khCy7qNOQZAWixCVrM+kKHq5Hob3ft8fzoOO43ZDKqT4NhaiC8Vd7HipP
YNA6qwLgLXr1A8O94HSGtXZbzMRzlzr1xqAhY6wEixmNbn8BzhsAFo6j64ChV+9l
TFpn7vwjiu63YCuPLlSbF4ZopSBiDmsuTZVhn5iJDBX+GDmDKwbk8f/dFc5n46hO
QxylI86XfZ6JzFTqLzMMZbriZ41I2AbRQBi/01QAIkv9w7pBB92oQ+AU1y6CasJm
uarTz+yxtHw+51lP3lEQLqGgPdpN7btc7EFrCa1+Fv0a6iqazs9FyyGrqw7JEgYm
EByEzqCofZzXegqslHuf4o17bwZFOV9/oKYKBGo7AWLKGwbw/Amvf/yXyzf3Pz7Q
449wIXrK1HsBs4Bxa4m3QE/HWYG+dfGRbjNXdbgFZaXy0hCH7U712NIDUU253dse
tphidgStN9EyGM2jfxxlJHEu2Zhj7E1HY1LzLmxKf91r4MysVd8FAiNQqq+teQWy
Sv34Hd1Df1dz3Nym9LWBdB7HG0xqMD+gXYflhOsUexmh838ZGKmzSh/IVKRLCHcQ
fVd5V25xp9Wz9J/FFMYYAvfo2UnimWov5HPVq4DRQ9jKsdA1Z6vqXQpwp6RmKaIK
zx5qla6wdeRrqGgPDpw1nlF3yHN1D1MgRY72zzzkB+eV9tFtssVE/3n5UHMcgbn0
MLX3H8W3XEqcJuoAtQydxqa3sLscc14/NsBZDW96TSOPKidN1dy5WSowJczpDGpT
DF6O++m/vzu+OvzuZEMo+ie7COOPSZ/7GhMSHkPGS0Y=
`protect END_PROTECTED
