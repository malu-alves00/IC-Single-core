`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JbwhIGx6vtVZ/hXcnyvSG6wiXrgFiLpJ6Z/jLJ42Y7+o83qYx7yMvYQuy5KNzHAW
vto+ZOuzdYjao/qi7Gm+p2F+/VZ+GyPi42ZsR0M3AzIBxaS8PcWd61s7tx1XJvIM
NHWntIxHbS5lS1+zQYReQ+bxmu5bGxexaIWsDvlOFrTUF2xqdJ4TC24oRC/E5OJE
Ofnwmx9JMisrxIOj5hbVpC+HfpvLqUQMh3NaUk+XqJyYaAa8C17dMFL9N9sXU7wn
IseZz1IbBLrPJxhiB9sUuce7vnrO7HjnKYE+B0hU02nD0VgCpfA7DZaL/61+cZgj
hEL7nGRW41tHO+bSh5XbQPN7jCspHwzhoOw14XRBNEt84Hw2MvFgUHT1WkvVES/a
TDe7iefYdfJULuYU6YjEgZTfubv9+7DQnYkUyLTCuVO0qVjpL/3QNPnnPJfYaxkB
IUOVLy5/AtgmTkj1pj/iaI1102TB3h2je0OVW1aRqT5KwHtx9ZBjSaJhjk7eKnpS
+xli8xpyEsXicuQ2zWeZvx7hwA697bA/7gCONkXY11JoWPbpNrnaOwFFfp3CHWSN
AZHnGUP+czrGEUQWp2HstoBtA/W3Iqu0YGW0aoRUl0b0syedpX3TIqDXRI55y/5+
WewCjoFb0CUkj09bsjl4zDVxMw5Q/EPl3DP9yRZOcwsxJJ6lOPqG3g/aWS33zhOr
wZNICBGkhTh32MAQ83PXNausfG0EaNLK7arrbq/T5u7m5kTdYHLEvnRMtRVo0z61
uc32DAKyGRpt+nEsX3L9Tc1kglt/kcm7Lc3eBUWN14JvQBRdxh6J7PL7BsBa2M9m
3EB80seEEWdfCTEmAv5XvqXRnEvjZV5wp+NYgYl5cwq9PWWUgyZJhfuEcAaJkLUf
lUKQwQrT/2xH9roIfvJj3sKhs0+qHGkHGD4rPPsKciBcYQlxcmx1CNzz2MWqHpsE
xRBZjFZhijdxfWM0Pyb9yv03WRDU4Wv03IMWu9eI00RgeLLWerlwE4Tvo7cr5kJn
/pDWStxdGiDlh40+/s8OHiEOSxcIYNpCE6qoQbTv/6u8bV+UxaEmHp+yM1HX6K1a
tIz5bBJrUAYkiYGw3GgYOGlXRSk55jyR+adnvl1Z0hVV5vIc01S4usywShOs8M+Y
sFwV0qmTj1k7T3UXtWK9kIIegyutf5ZEwEs5ZrTanCAY83zFlMf0y6dC/Plmwd7H
OL3Omyw9pVArnJheYD9f/hW5xLxYTyJ4fTE2j3dJjhvA6p5DW3ALFi/biDLvINOX
Xi85CVgakXTvyO2dTighhMTwIp2k3w+zpjFz7EIz2hax8rXzZYFy/2hj23+D3rBR
sLxsD/MRkL1tRuUzNYzDeK05ipNSIAXVOcyqI/V40KqQRedMnVviXwVIa/ebUx2m
QVBFVNafkkP+zj+mM6yY/troSUshaGY0KjN2WVXAjVLKKDUUvb3hjTZFZTMZ1R9b
9+czjpED3NpvowVNtjAuY+Ca8e7JqIKpYaxrk5T0DLJ37V+yCLrQ9lnGGzfIE3bC
W+XfXrFYlb6yPDYtzAMOEoU8qZdX97Dxqz3+qlKBKg1gSfPr3YZ9YzIuPONOSZFV
QlQO0Px2XAZfz5luLc0f9CXD5b48eliDdDWpWSH8poO0jKqaGgao7YQXqzfNQfmF
stNesI6iPMyIXl+FJpvNNs80HV/bpvMsh4ivhBch8naHtCjnv1XEh/a9j6ztBkvl
xff0Gh9o81zSkBQOoWQdG0sLtD3/QdHJqU9/459Rf2FT36ERdlm02PYXtkIbCnWW
onVIZyfq9kNBODHMwaCEQJKyQI03tfqkXoXag7PUrF+1Gjecu21i1EHre9EShgQx
MDgG4pSIBtrBRCw73aKfuhmHuNTe2GJ/ZpH54sMHNbQcjKGlIya95CjLjvp5abS8
VvnIN3xIiLQid0+qmGCLDIzPHVm6oHPRQ6sJKKD+0j84zpjfsrDA4qB/wp6DuHbw
8SaaalBOQrzr80aRNjQznM9kSu7ecDZEwOU/P9GDXZWinTMh+W/Ly369KE0ky4Tf
pJgGa3hDhfJyqsl07ZbkBU3oniXxHxhjSAyz4NSiqPSSYN20xzpPgwJtQ48iBW+3
HCb6xi37GF/YvS35DnUqAPJQe0Sd/DJntKJ/QWLhy5KttlkeGi/B3+3vd/WQYsZb
nST2wXEuRFwAEQUVMfz3+ktdVMqdJHY95sFFaDcEg3r80FAOg4OphRUn/iA5CJCL
xmfMsK5Jbxl23TWSHouS2XwbsR65BVDCBCGUD3Vp+o7mlWv5q2EHwwYbbc8aZs55
S2daiB8emXf4DRTxvAy/mdHhd/8ZJcJKAJek/p+KVVi112yHTXiZvx/tfcPy7u3p
x5pP+iR30QLOyqOoU/Y8BGMjj/N47uJ6/wVy3phZNgcexKz6Soxi7m4gZ5UL/Xzv
+iVqhXtVGmvA775nO9bavE3IwwoMbWCGbomlsCmZwF3QUYn4P6QLERzPcnKbim3B
IiX+BnHZK0+4PqWh3QtKK6NlkHF7RVQtrH0W3DJbG4tZgGWGBx3kDSeMKI1i1uZo
jUivMVuCKEwpv/YPDr679BkvsM5GFAKVy8BrQzEa7jwv4fkLhGO88u6sb9VTlRiN
8pMsKx9KigEIu8+rXpyg5Ijylze7KCY+6NRDzxyrhICyacemRJJ3wruLyz7hIbke
jIoWEXbSwH8x+L4lZ+WVM5VgI47XLIvSKYtM2675jFeSEjgQjAy2ennWV7j3w8Gy
4M6ovqkcjiaZQLc5pR/N+qI6HJHM8phpnh7DD50HQFEC78LZJbXQvYJEA/lqgDpJ
cs3rg+Fd1Q4lIVh1u3JjVhFUQ1xgQJSZOCRoVfay7t6Odj/p3Ffw97bGz/LhZG+o
/2BS27QZogJg2t6sdjlTyGtxYEWKZGXrFb0Xx3avQ4OwcOBXtNUnfO+FxJXE0iS6
3YXGMF+GB1xMkZam9vfBK98EHriQ39RUmxCtnbYtVin6TpGQNI9TWYqhcnYOzwt/
moZKTGcxETZe/G/BjoOdFiy/mQj12YFMU77+1MAXSBl8+ZLLSd4bzjY7ukGIfZCU
b8SdU5XSwx+CbqcObXbXf5scyEmyhxod6R/it1Jmo8aRCa6P+EC9yFKEjLNK0kzH
hAeqa2Ggca+8PPwESVk/GLyE8nr9NFiLwbylnPMFLJ8pqQOEo8wNaKSrbEcD1TvV
tuyITsRVUCxbq7+QcKQt+6pXQyLCBUgcSFkA0b9BCslXEo0c3SoWekDMwbcH3JD0
cz/rFbTTvZnjFLec4p4fWZ7+LCf6mhT3ODw9JMa58w3V9IwUBOY2iLO70g7hT/NB
xWhUqv3SfZGyihFzy3qFKmyq9lUqpqR9J1rKysqfu1y5PRnmAl+9sfyOHjRkITlw
s/vD8xCPa++Tl98s7epUMZbMaiGaPQR/GtYRGtwgKYhTmZX1fLtQbApkeaSHlsex
us0gOg+5BdMr8hbVT0KLG/7xY5bnRJgwNjorINBqXJRdsOTnxVSJ0OZIIHg1Y07C
Bq/0lcL8T+XWA4zp1/NG+Hq4aAqKUq0tm9XFC/S23ojnfDbmK84fxZCkBqou8Wjr
XfNQ0UyHs5sQXtJgpBDjSVvGsxfraNIN2IF5yFrODd+a9EaDOuXLjEiQ/sPmB8oV
2nqfhdX0kMrCeiE3QGfrDNCOa271KmgudTU9LcQPj0CRzGQQyvy3f+W/4tTO8kCh
Sq0YiN8Mvizzr+uSBhYEwOFXxwV7iu2aaFTefJHSjpbbVExAA0cgGZ1IijG0Ti7P
0xo04iLeoKc4uasyWm1Klr0RNEUxdP5SMwOXggN9lo2/D1vQyNlXdoNyiQoVkKWO
npNvrt9x0nI/EOjS9sSztE5MlF+lBA3ekJ6+OMSd0xwhyZp6bJ9fQtnSQ3N2BV4J
MWtND7vHEDFEXR1flHNUlFh3TIqOrbR/n5FAaehOcr5F24mqv4Ey4beLgvFPzID5
S1AgFFlf6Mwrj9dTQqjlngVcXDvNmNyOxt5sCvsXfvdb7G1tJjGPm2AN03Qn9VTY
yJXEePOtxP8yTaciLfP5pRMeIs/zljIbLm4WFf8706aB9eZRRnD0bhy1d7klRY8c
lnDy56Fbunmot93W6BSeAf88ClVK9TY2hcTdYKST9M/cZ9S7OaGOCNL5tmX8QuPp
gfCkb9cTYFnGhxUBOmbQMTP3gqM7tGD15mIqHZUrvlZF45I3rgN5PJgFdJfw0MAJ
Ea6O0T5OjGHzzaYJDyk7+6efykxzPIItDg/B12/t8slaQGZEh99GueIJJTxnX84F
xXdCAVvvvCFJTDS9zZcd5ghFoMJgnM2kFPdE5zTGoI9prJWGawMEj3BqoyiqNdsR
8i1fj1LYBuCTpB8b4Rnv2rDP96qWzvni2Oph28DV+wEUpo+HTnAJy3gVhIiJwkhX
OtNjEA4wc7W8JL79OugiH3yyBfpDzF8JBN81/os2wRhH4Mjdmm35zjYNQ/7Ymy85
DL+LRsW5RvDtNgmTJZ8gUcaClCb27pOHbeIGcFCP3p1DbXIzgW/i5GrWmiEI5Gy7
hPVmEbXVYS+0AwK2HtC8kqxPlGEHsZnY2z1D7+oZgWZK8cKQc39c3EiBpTC3WEZS
Vf8wJljVvKc13t/oJIQmrRs339Ruw0m2b0fuf0JBma31zIQrk+KKiJ4o/gol8ZWe
SBV5aq6qAxe5jYxuNbKoIc5K00DwHXZKBiTgAVp/IQSxOZJGzpvxRLTDuptLEwLV
5NKfenpohfyXNLnIghkrMigjhGYjA7RuhPrkpcQV08nko7Z0bH2hBdK2rbGMsK9U
6Whhvj0HWEhSyByUwcZKA4Dy/WbmunHkaMi/Z95+n8iTAyvOZvnGBHpO+Wm9qrE1
iBS2sH/z4SwlJ/yDpTcoZv234gRtYAFc8MWgzpMp4E26rY9m6JZ/QKv954ARrxuS
ajAQqzEeRHZoeY+xQ7YGEVb0+Aie4MhyOgciNdSZTcIBD2aAVJLbpk2y0QOTqhB9
cpIOQLwpHzbVpKIV20yqmhL19g4OW6iaCuESnIySSz/jX5RUTqq1sjDyyWJzgp+e
YLy2c5fn1PmO4nMx7j/L52UqN6gVhyNrWgQVjR0GupwoPNeElcwWYHGzi7jScGxy
YfiWFzMnC7wh10zLDTYkHiQWSVX81my/a4N7hBXW46MpiSfpcacfMUu9bDtbgIkH
Rms3GDQJPf8szVdnxKKTcw6A/j8F994STFoifQmuLQZgfXaMTQXpMBrOMf73lkHR
beqiW4BzntL5/jy/9l47tFvvLfuw3iD/DKOX6Y1j0tBBSqs78fLsFZaOdBrK+Ycr
GEQykAnDOM1nM0Zr3TXSRbp/aunp/6I+xnioM2IfGKS9BvJa9uMoWmTj6oKeEUxQ
yXU13hjFTWHjaOK1E42d97boa/esvuLLkjT75tCnLENJ/uW6uVTzZHIGF1z6qlzP
Kd3Ds6tSs9VmdG4v1UeuJObRiJprO1cZ2N6ugux0fSx1oXGmEB9UFKslcLzBmcU5
MkrXD8jnhogeZ7LxJwtuF7YHJumUwptJLH+Fl0l75dvcd2kFVxQnA0Ht7ZNSZ9xS
YXYTRGDBIhUOMh85U3ItaYiU4jCuT2qLlR7EXQq7HcBqqWG4sumGIM8hbOLiS3De
ymkA/8m3S9JdXZh/Py9NvBxsuKsnO2zTHVvMpxIA24JthnvFit6qI3L+iqbUq6br
i6RdRe4QIHQ+yWmvRls/aaYP9C3nXD7eq7QnzkeK+6E8SQ5tbwgnPLW+vVvMMn1i
bG1p3SxWqajRUPoVUDtrm8R0W+JpYUEQIgs6dUy1HJu/IR0Bi1kE33AWI+VSe764
BRwrObMJtNbNPM+SRgM+5p5KhZ5IO6BSRNQrQ7oYY60VU96n8mbnhrVLYg9eaoxs
rJBfxO+AEQLi2vpVZdfacSf3Adcsqw8ibRCZg5fdErEpUayB3j9i62sTUkW8fECF
Rn9M0XCsSl/LfAvNCFb7VCanFjOLtgDX5m5mXUduxWfwxtqjQqdtfJKL7IsuNhLG
3LN0qb2uIq1PS+kVLylm03jJ0TskuLuHAnwaehRhVMZoPQY6roRLhD7YY1b5pBoV
ypKKZGkkx2QygW8V7qb9OWmqzXH9aYatrcJatlOHcoo2MH7ljPjiPxgONkgnSF3E
QTlXjxyhKEniNKEkFpO+r30sOQ5bMnWxqUS5zlmzxMxQgOKIEd3U4HD8sXK08n6i
VoBoEsxT1Rf85z6FG2pMgZvixPXH3Bp6bga/xYBaweeSydscVJ6s2QWm2ye8esqp
hsTBWyPcUy1scaTR356pL4gcfQjpXHfG1DpOBCpjESrLWNyZ/4mfLoOMuLwaZIh1
OmTbuZX3UvxGFYwTSGzgRDYEuawWfj1giFK91KzQ4ImJzAzz5TSwUYlILoOiSMIF
CUmWjLrybS0LqYNgemPpF3IKsupq9PS7ZT0+rRhsigNNF9lvCmZ9VksOlj6TaNlw
H4oHJ7ogn9ND36y922wRDpluVdbhqt1zw/u67FVg11Kia3RJoGcw09gG6pcTwhe+
zbxM5lBb8sQyXRdcEMjZsB8+yQmcYbOOeTuZ2kUeMv5rGx93oB42aITa+obBsI3O
aMtGN7Gmjl7lkFmFBtF6D+BBjOZcnGaut8OR3g2tCBHQbD/09AnmpeoVPF9v/W+A
9Zh0pWFPMKbDmebRjjlW5Cw5G1FsseJf1mcIvUxRG92mzn/CDbZCfUTLHqmBlH+4
auyP9EZUbiJucoQiqdvr3ec3vNQT/fmEBjhoDBbGs5InfSQK81Tk3tdpgaMNPU6C
d8pJB+DaKx/P/eCzd/9VFPlRG082cfTtiutxnH1PawDTlxkXX323c41R+hF/RFbJ
74nKOMInaSg90JyD01sd3utHiilmDzlNC4hGfHjRGmpB7BBc0dDB9xFgLfwKr/0o
JLaY7w6/3v0DEMYozs6Z2MEds8ASrQkoQFWXhDn5qEjeR34og7kpDwtlSJXQ7kJZ
Mzxb5hWEzhyU/M0n61+H8/9rYFkbVyVBrlldht0BRzKMaK8o4ntu10nY2SN777Kp
oYqL/Kf38onzbKJNSfzDeglbPIR3PA83WfOXYCQz5dfBlO0nA6yTLDAcVK7ZvhW/
A00SE+6ZqXiRqn3+QQOSHWHsESUcnP7ZqsOyfVkc0re6YIs+ciFb0sLap+l/Nmtp
FsUVYr++es6MtLqdlNUoUGmg9OImXKAkaHHeK41MXUJIOPOqh88ZlZ7mllHrwPoR
pRe3e6SHI25zujNiyzqSr/y6WCrP4tGeLr9Oe44F7xxAwzN4EgJu5eKTNBfKNNO9
Lr+R3D1g/dW4g7l+2R++pZjy0nUYPM+DStghuIrWBSu0/+tkLXmAdtt1Dcg1r9Gs
2kYaixBeZnRvxAWLCxWur0HfFCsO2IODQt+WPGtyGb/1/dDU8s43Cs+lFbQgl0y1
s09UeMrj3GGNgLnG4j8tkge7F4/MtWHb6f6aPJWloK0uxSFDpsRI6zlVRusIZ5Ar
6h9BGNcSrBwwbz313maldWyysN8Zw2xtACYpRH4pJc3LpDV8JTgUZKVI4a/NYGI6
Kmjrg6qT2pokjaHj0nfkFbcqOQOyXI+WhujfluTpfrvfnK1hP5IwWLnJols+xQ45
r6MFVGmGj144gyF/hz92DvSZjeYvXoGqG6sWVfRC38Mf/oJD9O+WBIJYLmugoy9i
48WqdFJYCT0qCiDJ2kQcON+DFBD+SLXplJ4fpartUSEYCUvbPCkHmJ4nQq/qxG6D
JGrTv4dy69lISfkMfIU7cieTpjRvogekLtTtqSaVDMPQRiqYDOeHjnSY4XneurTe
DmMZuprwFh2qVOnmlhkgSWOPT536+QkBtrl5bE886BHi0NUnEqHyUxc7LuEnTgGi
g8GszzRaa7eao88w9xWqfd381NJBV1zInD/4zEHLAPspZDBIqdBGqI0lhH12pM21
+3onJE7Ou/iGmavZegQtJx9wBHJt1KlpW2tJC9evRRJRuWwA4SOEqT5a8cyHCnhy
PSh0XVYrrPVl2RQIsebpr521jYXTTb2V8bRmr3Q2zRLLdw/8nIj1qMd3t/iP/xV3
lhbzKLs0hrwEWTeEl6jssuMjeXS5gfkA/H46GK57NlUBYtUeKuAfsIo4z80w3/HZ
97ww5M20wmSuGxNBD+x4enkRJrJUjSBC1ac7wQsWbBt9VU48kl/+yak880kAn9Kj
a2G8igSKkCNhgIWVde9hElIwXHgvh960p2Mfc7WPrQdR0ySej5LIPPxInhfDb8WO
P4FRjaBOuY77toHNLZOSbma1EGzLWQnMuVVBJLynq4yOjh2FXtlKuR7m/fSgrWXi
M4XJULVsqnNycBsYvFMryW4XLh8fwJWAxWHMFPGcdTcrSgxzhCpMb6fN6L9TbOpA
4SgWjiQjR+QOOjKhq58u3VdD9QmONjFLpx7I4u3G22H7rxSnkR3yIV7VOD+g9cd2
hFJd2ervFbTRnYgACvxfPc7uWYRKxyVNgRGtBl4FrK3iSe/WutEblksglxcaxtJM
e3waFN8UuyZh82ZJ3h9RRyh15dK/Yuh4jeQBHXskNgbPrtn/zhiGJeyWxxRN4dlN
Rn5WFebvfiQqJeLrO+Ar9B5hxNxL5Z7nmPniXqNal1+3FJHfxOCeMzyHqI3T2F/R
gz3gDPj+lYS20m2ClbXHzBRS3QnI3Ug3Gtv274nYCr6nFKIDwTSWWdfuyDmTVxiy
sbzc+7U8TmGK+rpXJTD3O/5Mdm8RZZwG3HAHJyfN7xu+3436f4ec5Mk+chYN1NHL
lXr3pl3KmJrT+BxbKfVu3ue6/8W1kMmWGKCLi/hI1IqejpnTBJ2gUXQhhF3khh3x
E+93rM7YwFb1FEZjpuHrVw/+ZTCOiMHHmlIQo3v3vr9oIw54WPyxgSJ375Tmhc+q
cGe7AmW4vF4f+onY6prXQOIw+E/59fjuGkdEZPSqde2gBeM7Bco7vZ3KDIrMyfSK
+hq035lXsF+NGEtwR3ybRjrSPCLKrZjcwTjPLCbAv4R+5hZlIIBrUDfIdTl32UuE
twJHFnscEyE3zTZLMrigZQN6VRbD+VpviAzJ+FtX2pUrQgoOYNNK8UCNgdofqYsz
z04Y2Vp10aEMtQsKLY5XVWoIC0O7f6OSMN4khuUITvkGiY48YwHBHJ9wf0181uPi
gG4KJGms+/2bics4vjtoAR/UZXPEJXDSsCPWHieKNJvAQhD6wlS4ij0j/6zUk/io
ZRmy1kvCPbkWuJuVf3Knw5nbm5Uq2qu47MK6rsqwAOiuQMuzHdOFyvgbpaA+OFig
9RR4+hiPmek8dfIkuAT86/pLTVmhMUWyjBKvNkhD3kxKzZZLAbBMYVvK79ZQuPHg
YrALK3+3Pja7At6XOHMWIni5+cluHD4DmexJJKc7JsDyxASGdyI4XnZYyPoqdXZR
F2L6XgqU2mmRjYUR1pORVVLRFB+ppc/NNvlhsCeK5KMESfE8m6aWFqEEpX/Wg1tC
j03tXDbkxmxPtbYOph1lMw+9zsecb/gxYd7n0ZdE4pGWO4eOMvYO+2ooNDCJW73j
kwyPuc6K5UD/C5mZ60uVn84JDNhQwqcTdjFJxOtylsUrDbetyar/Dgn5zFi4hdlk
Azt98BikQ2xePnG00fwAEPx/owCWzgaSjhZNl5e0VK4bQbq8qUDsAZ0DkdogG1xm
lhQcw028gyaGJ/3Owx6YOp5fiWW3tZ5G8y2r2UvusRf3Yx8e5WFb01+E/Jt9kQNn
YmbLafgBVgK6nNVMigGcnJQJ+6/cWlLQBL5KMcq7vGMMWwbiIY9I7QnFKLZax1xw
FIIZLQQc2rowj2HT/qcKb2KG8DWav8qPSdt69PZNaX0cZeKmRJBt0jl2bOXJf9mL
PIQR87nD6R/F68WxmndRCFXM2j0Eh6R5/6cm201IFvNmurbJGzqn4U0T0X7+a6LM
WCXYZzgrdPTvUEAIZIucHvgRW1621v4Hr1KGCegYHx/hSJF4Df27/tZRF/Nh9j48
czqbiwbt1C2On886GaBPQ9GZlvQQewoffGe7STIdHypTbsvXbFOwnkIV6nDnBVgq
w9OYDKo8XNfLOa1EZJIG81cvW1QY0bUrhW2pRwlXNPZQd0Zz1CJ/B70mCeuQLhzG
8YKAo15n9erYE8sJTt69uwNXRDfNDuuUjJsmiUGv/HJVqW8yM1/lgom+9xBdIfdH
WMX8Op9OcIRQppiQjAjGOWQSFocgm0kJkBdFQPzUSmShRxcqeA/BECY1/HY5XSKl
+a8KF+8aVPgmPb6gQ1PAIC/G2TLPiSaIqfm3Ms/31/L2OIuyVAhZTzu+ysEr+fKM
yXXPx8MWkk3EaZ/DvjkbzS/c4sqbqxXRUsYvjqeQZ5TX1OnPtG8kibrtZC0FZ/KY
wqFszAYmgQL/2mgXm68Lec/Ov3bFhnfH+y9QNISLyZcCrdf3+HhB22QpJW0Q5gS7
J9FAHKqrYH+gQgFwE5Qgqb0nNwd+gAX7Cl6wdUr9hKQ4RHxE4QYh1/f/58bIwTHs
Za1j3vMlh03B6F0H+tffxQ6MQI4VomHa+8+EIkAKmYwtvGQoWnRvIlGx9wDdEf8/
1koMyVIM55A+xLN5mJVqXT6c5HuZ5XkTxm/iFaPmqApurBQoW81l4IR4/9y1MDj1
BPTpha6qSuleC9OPilWsjrkV8wMlN4Cn9GtYvAs4P0XeDrjJGLedI0M5WfkzGXpX
JYc3Tl2fSd4JjO0B+eQARNu6nBfdquD6UiVLF30MKdCen2khGUw8HRg0szEb9cHv
iCxwIhrIl/xP4mEtCi+1mYQ3+5m9i6sqMbM0Qs+NK8LiCpJC/Kf4AL+9oXw3KoA9
49xv/VNhwgmnDyLX+38RSd6IN63EVFHPLZQitx6dNrZTlU+AUCA7c5sceSFZZGBq
UlJ+Ms9VP9n4GAY3mWgYZlIfB9jWPpABd1iqZ748virv/5yZG/TNcezY2VX95Vtk
Cj5uPyqd0NmDIwLzkKLL6Npf83jmOZTjWki+Bk2f4hMZME08yV1V3Q7EWVrJ7igI
Hf6RxChzXtMuNm6VhJzG0jN71j6ihW73qAyfmf5ySGYQoRU4jHq+gRyWp2rVlPMR
eo9qOd1QR6cZtRlkzja8znc+7ux+N2625zezTSOtPo+4r0tyeJRbjwrzAnasYaAm
KQn8dsP6oPSlPWCw6ixCxxkDD9e1Z7psbjwqP8tZSrbP18BqqbjTiy5scKRn4lfM
nieUv3iMYFmIDiXTUWxVYcJEkpo02QMyChz3A8kWCi3AncBBvUMhapH41Ryaed4e
CAiSVrgOxcbFj9s/dst2R8HwzOR6tYBriDbluXyExR6q+VG5rSXvqV5slb4nkI3G
aLzquZ9dD+V/vuwB6uy3UoFI3xV2b4ShxdAJICTmBZUnE9+8fgVxZz8+mMjX1Srr
uuL/yejyznGAeacd+vqn7bkKkoWPaaw/64UvUrgI1u5VTRCQQwWcJQN1guq7IyRX
SaSNDbAGbWlgcdxu7vk9d5PeJITDvqeySoqq7opcPCQslXwu9aGy5uWS/9wZwq5q
ll1ymr86IzIDOxdKSwpL4aAtYa1espOB1zpkRereNE7idfLXS7L6Aork320Kp0TP
jHi9NmusfWtHkgqIz7JbtE+NepXNEKeNQAY3I1fIxb1hg2wTHKmRFHo8NMqjlPNA
bI69E6Kcl9fiJaAarTpC8upCNAgV+bSxnZ1x9OjUyuBvqBcEcV/bREDBUZy7zdms
PWgNIYRE0Ab6/rMST/YtTLDt7PrgjNq47tBXCLIzGg0PZepXwnOCqkZTCvARwQU0
bTTgZNMHbuoLLRiTdGfrGoZyHnIwh8iCggw1pBG69bl21LS4A4w8JNux7Z2opBmt
EAzbBzRj+d6cTs0HBQTAVfm1fHK7LZeYV9IzLfYIHrjsBzWRqPMzSfLrveRxr7Xm
QQ9qAPjTp+E4ea+Lx7+YJV7/L0oP/gdL8hshpHV8RrQW0ZdnUIsqo8peeHjTaUXR
H428Xo/0/q+/ASf0IP3eEkmHxAWjlJ18SSknpjDAMbe2oOAeqkD9KCUPo6juaqmR
7Yj4HNG2hmPO1TwaYsrJXysADTE5fUfc49+SnfEwvqg2vmwr9rUXMeDbYZ4i3xMB
1MgU42/7JUCdgJOUadfEeOFzgW+3Hwpua+WlkDK8kaXJQWbWpnqhFgrYZyF1z/v9
YR+8UDZRQlhZ5Gxxf0+iI1s35f0ihbVF8SshMVu425eRvqB0l8grM2REWd55dbnC
iw0se5nXvuAIEAH6k45G+Hf77edSbdoWCaktKgwkFOQ8Xh1vprhjKWZXb5US7sf3
J4Q/DyE5n6ATePOpFOhipmxQUEfwOU5kRUjHvUdqWxYdez8kovs+WbwGOBrTYbBF
p6dTx/6PNqRyHKLJMJXiML6uS53Vz94voNIzd8ArbHxM7rThWJWdKATEl6LVakgX
wGzF3/EXEpo1c2MneNnENEc4mlKyqGtiGZmAuzer+3X58HFpxFxjhzJfZo8+4ImC
PUkiE2ySITw14GUeqXmaO21c3ugOlNi+zSaoCSOffFnIOuk6FsSHB1Gp0ekgkD2D
RITpjrh2urXVvk+spS73wKuUEogJhadCKPCS73fJVQDMLFzQOkgTNWCtuozlrhUp
bLohTKVt6/BUfZsAnyCaDKfgBGCos3G86NB07eEQb8sQ3dbiOUDmxk0W4MishlGa
a++AMrS6Iu56se0hJo358vcO7CO2LxoJ8hItKOOQMZkq/RCYZfKYxQOFrToO4V1Q
iIaBs6ynJinZCI8oXJA+VyYdpXcSe3x8Cij3RA0SnDvDUJMdkGWSLGJRz8TxsyWn
7P7HHoht06VkTy6wVL9cA6gymGOmV5UMwM3vf3e3YexUZLGv5bwOr6rHKe4EKsKg
YzN9rlJN03RN03uzmoF2bdXgr5yoX2DXDcfd82/ab6UoXpji0adHlUDIseg5dhki
i6l5U/3SJmilUBuETDO1RP3ecOWJZU1JmlXUc4IAsPWhMWzIEldDwufZB4V74UUk
GaspDHg8/7b9QNSRdTNtceRB8QbUdQSmndmtp7+6FS4N5425M/nBsK9/xvyqzWZG
5z+MMLnk1d7Oa0PsMm5UcJoCNHd6vadGKqathKE1cGAONr544eP1DzMXZgInPnYe
QKjvqFJaf9CrkVLlqTvQ57WmwkCm8QxVumgzidHCRZ4MgLFCTVxyWbriEaQqqQ0V
AxAB7t7KunmzKB0qrtQ5KJZMq1hQfjZf5fGK8KqYJpd985UKHIMsIBkKsafXq9qE
u8YPCKukumLV2GEdZqtqjseJwKJj2t9+ykzs0D7YR7wrqU4+LGuEOHnDcS0VEd+G
bAlvttVrrRDbCvFm1fO2YChczB/FpqtpLYCdFOhZYCXrIZF7c4ABUIZYCo3d4lRt
LuXcbNyckSpP1aMLO3Vsa7vzGEEkhcgWrEAYQPel+yULEnvbgriuBS50yBhnT3K6
txo3gDHHfEnZnw8RlH2vfefaoJdQWvNTxoUKEQPfjbuvOf/a24oQ/j5UwLEmFTUo
JA74HUEOwvghKTSkF0tIqK9CzwQS5F5EBbqIjeNljFu4E7F2yLWRc+TR+NijjGso
giNNwbIbw9z6hJw5Xcb9laFBq3txSJCdYuAeP1jUJSPmzN7A1nNi3vkd4ThNI6SN
348QbFWq3IE4E5SBW2RXmffSIgMVFLZRH2Enw9HsKRU4YovzqyHCBw/0Bc357PNn
46sWSL0k1OVFJIENxCJIzdJ/0fBQGkvFpg+Da3eV5oAwAfW+rsSV3IJFB4uun5TM
0Ux7U4OzGc/fhFQARG4ikT9OXR1UChE0gGo0CXvgx3VTrVdZMvyqz+3nV3Uzv93l
HSjfJXwi3SfOVxaQ8r2iPw==
`protect END_PROTECTED
