`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xcv4oswvPjaoJZ1lJOj0L+TYyGXtIaQjurgaII9TlDGzbKctrrHA/Hcbph9IlyLz
j3Q7rZgnzXcVFckODZkeoZhehmZEj7WkoNU9Iulnx7T6MZ0jKe/7pG/kkBVRWHPE
Lt91zT3OjQcEhpIk6h9XHM82W3UvBtn2+EGDN2UL5N2uWxNnKa0tcL9S/hH4E3td
ILtKYlQ+KObjYFkr/0oTMmNOG1Z1v2TRqfaW74XM5qZANpYxCRFsAoDmfaymK5De
p3P1TaHorKmv6yL+U+gpm8fflMuSfiNo5LhNWKGeoY2AsraUYPKePvLgFrcGM88s
JRFQDFJhCU+98c08FFJhgaChH4wIiCKNZhno8yjTlt5KwgNYQT43ki3sBEamjuWE
goqplP/kbJO0DcuAjxMiSMRaBp/A4ulsW7mJKnYQXVQu2CRdIUYx1w19E63qOoeW
MwgKTCBf3gvYCoOsKI2ITtCXu83mZsV3DwsWLtkq3pvOrpYAPNWSg8dVSB7hjdTz
DEn96ObcKTiEWORDHSv5fSBA7Gi6YLUSSMQ9Qs2D0kr0Yp9BiD8lOIH11J78KZKm
lepTxRJui/CWSDXnYBZRaXntR+S3dydZDp9o9E+nCgGNLu1RClUbFDZOHhA3qaUJ
gg/qkBG1Zyv2QDdDx9RDFXLuqLtJ8i+XswJFubs5YP0vlHMyzJfsIm0cHWfYOjKY
NPeb1btGDqIgalW/nv5T6Kb0XBQCysQ/HT8SOvLYbOT4dap/qc+3kjXdXS9NxZbu
DCMDCCHn12fRMVkbpDMJcj/6ddAQ2teUbXBiC2P9MLolT6jEkBaUB9BfRHFJjE8k
+K1taKTZ09UE4oR4gyUo12clyQ2g2ZCDVwWPCozLjiKf9UJnwJhDSDD5HVqASYA2
1rBCMSZI/Uz2tf2mxaL788qm2EwNQBg6Lz3MxVxVPQfvVy0h7MX1fTYhMooXNSit
jN3XF1oFEsCnTUUFoB9oz0lWiFMzck/JVZ2wCN1XhpRxFKOG1j8qRDJzus+rqm5g
a6e0zKI4PKFJLRufMLm+rYvgr0fEtN/KKoNh44c3by7LeBvryX+rj5y6z3JSo292
V5/Ew77h9Zgt31E9czfCcbB/vI4g9iZdJ1qfDwbGmjdbufktfFP5i3l+UcnytGij
l54LDa5srBlrqxIHEStl13srno/m1ABKadqJTuDevEONm/CF6uV2hZJkpeQbJHZF
rsinrioHuj9udHn0PggZ4grwrOvYR5bxLiZrX5dYmccFaKKyyknDIikTpSl43yC8
`protect END_PROTECTED
