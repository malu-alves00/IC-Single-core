`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UC+iov/fvpZYDv8T7sJZNVPojjtHVMY/pTWcXiNG3aFqC1TA/Vkl/kDilCvxJJzb
+yOE+E/V9h9BiQwDpp0kEMsvNOQKDOQ4/tXp8nFU023nPNBOGet4Y888r+JJiVrh
tERa64rbmmeYUhXKzkvA9pfw21sw/cb0MZq9mVmExAcbks/NVRtIZxgDKxcF4ryr
jfRNNs6KIxLCuvemo4v8is67OvTyZISzAgVnK47UzIru6mUZCy9V24jfX3jKhx9f
W8AzgTc3WKLq67zCl8+uY53AfgNcOrVm2t8WfVn2S/hdpBqTAipkDatyl+GDvknu
cnVylY/DTnwrUKZPvDMeYLSDPsit4XPH1tVkoXaIKiMiXBuuBBoV2vDtkskAvDJc
`protect END_PROTECTED
