`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DdFMT9GKaBytil47rCV1mybW4LgPfKjWMnrYKaqSGtPb+yIV50YrnbbRjPWqOrV6
BVNH54dTYSLZ3CbkkFJq3OmrkKWo3J1D2B4knXXvqmPCc07gEZ98v4t4wuLjZz3V
6HGEFuEOAL2a2xyIiMWscMWWbMl2COm1HUDHeejQKhrQoYlUHqWR6dLOXgxqFI2C
R1cKa9Erky8dbWW3BgFlIkMPeqFDuGPnKlSLJ3gMiNVp+1XIiphnNb6PMwL4H/Nv
bJs5CJQidOfrrcjj/wEYR/z9zQQ6Yz0P+pAoejyf/vP+TXbCSk3OJXyznPgXQUYl
ZY2R7iqsdcxIqwZOWZRC39ftuzkN/knhWQTmTIsm5soWw6zkyfBu2QGUMdWE3I73
F3QppSgHWzDWKWA56g/2gG7SR5Z4jp1VAIfSAprdDcLWUAtjQzNb0D3jhE6VHhcy
U3ewBJuqKEmpG07bWNfv6o6uQDzD7d7AEdXpPM0ezMsywH6R/KriCkke88QI7Kl/
aZkEoRxWJvj8gGRJuW0pbVbM3XM/4YZZlb35asMmgvM=
`protect END_PROTECTED
