`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
q9xFs5ylruUbs3gZjEyQtM9pCPCu0hQ0Sda640ht6fgZuX/aowmaNxGIjTqGdFqc
qIxAjC0alIaYL45TI/yhqhRSWvxVZJh/pXjdtwxcxGOtnMptgtLLCEca4XMuf14s
xqtVBQC62byFRhsi9YxgIGUDNN7M+mYCvH8udL6G4TXORgoWy1lx4ECriELZUUGj
nxVf03kLNYALedbrPU1XKPpPr1PTp4whrcS9QbtoKpXGOnDh0Nnx2vpRK25MWho5
M1da/I42+Nec5oyCFvNEtrwxCQiFyTLAmiOGJJj2/WwjwN5fqWujSED6Sj5ZnBEi
CZy+momsSLmxeq/kC4swfmnJNfMdto6vo8QgmVPOecGxG1FRKnAkF33Td7W/Bdoo
Sh/LYb36TWVod1pQIAKRDK+uKIKA4zuKO10GPzd2Nfe0jUyR5qGmi6iOHRrFi0ev
8IwD0guExel5fpWB153rQTz+KoxplsQQnNEreDhS6NOzIZeQP2f8wmcsokFeOFsj
WsjnRfr0GVy/ywE5ODyIm8uuPEt5SWdDHWKCzpcNvg+Z9syN5HfTdW2t1MLXsYTF
8QZE4t3OzEmoBlIcBc8uS/8fHiTNTVlAze+RgufjkKUlcBfG1wUtYdueqfZ7L1s8
tKGR26HsRQ135o7GiqU79sfYbfMRqDDdMCjHzoH+5y75Wd8jiiB+sPqArTcyHu4k
ArD6j7XeUdOfu0jf2CdaKxs63JK864FRpGtl01wWT/L5USAbcGuU4JqSjPwDpQkv
`protect END_PROTECTED
