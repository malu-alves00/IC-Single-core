`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Frxxfyqjv5ZYQ91Zd0l75lTOTKAVqgRrEs/yhA9ck5Or6AstgdpPYX8KNbzk2JDW
iNMgOA/mssMN3I3caZlxmyvw2JDmQjsgtW8OaSpG0umDeGD12lBp0ivIwKNBWRP+
dQH0hSfK4C8J7ee1sy0rkhm1XhZYEajIkIddHQR65PHjjd2UswFJctwb2Rc9oIvx
GtUgS8K1H/v7YkpdlJ/uyoVuQlSwaJQ1qFtjOiske3lXd2+TPXmmhsK0kYtBKlVZ
XnmBIlNTbsakzv4ZcjY1GrBwfcQvSaDULQHAFE4XKr9LZChPLSeWu7Jd0xkv7+FW
mOtIs3nk5R/Pe1UxaK2IfEyKVi6xfgj4tYGpx57frVRz3L5b3wxwmU1wDhvK/OqK
hM8Z/nN0AiImguRJCm4oNG9LDNcxhNP1zxSXjUHr7mtOovIZlMPc4lNjB8soy2vb
Fkc+XHN8ww+erXhWUINJe0CtlcwlkmVzWJ71BLl/ehwiaRlyR88PgCKu4pibNBZC
eqfwfFtsBfdr2cLoGxf4dq0jP25Awig328F0zOQ4Z3X++vvBjpF72iCCXQHJwnKx
/qSha7cWwftz1EVMU+WGJJBf7k6UMMWPSvIXwA3R4E8bbN6IJgCML204f3uPnZle
ePUP/zhn0vU+YalkIOZB4XcV1VwadY30/an2pwOptK5MkI3VM5JgOXBO/tqaVRVn
assoCcMeBlFP7OYFo3IBn4eTqVnaYSKQeCOdwixina/t7x3ts66chLIojOLypdPM
iHTKTBvt+04DjcossB0zzYMdhfV7KS7NJ7JZxvlZfv2ohvpOdJWwezENrkzOZ01B
XGbhxqHxmQA+RmlmypU3QeNur2mYkVlBLOvF06UfgwpNHtvYEyOQCmqeeyNMFAr6
zrUsNXHwpgJHB1l+BDPu1prl2sIeE5NhjwWlhz6VcFFI1I7TLEgW90Wu9gGActQn
DPQ2D+Uvg73IaqgkzCrU/b7ZyrkJw2YXBrFvCIWp9zk3UhWlnmMCXFaP0lTxRZfY
S9/C0Rspmt+X6ZsMqkzAh6srMEOBFvDZJOevFluUEYOlNWpLQ//khGmpxJYwMVok
MsW704X/ArF1kC6nYKmTdpNPnJrrl2NvlHZCDy3OGRgz73o/so1q4vXwMOlN63QP
qThA/ybR+ULgsEK8QapHLO8TvH1TYc8KmeaGVitRa3UIo7F/ut4yfcYmFiWn96lO
hkcPI9VD/ubFMs8aUxEGdxMqS+bcH2WcOzQ4+yBB/AAFikNxNLUIyVpNhKAFEuxs
MnsMPHKRUGyUsF+6x75Yrqzpkl72RT/cTscbex2CFOmtzHWgKAh6jsLV25CC02an
qAr3WDuUOJaqLDkc/dZPdarqb209rl6Zw/qF3UeROkr6xtbXR+ZssCgjab13ISI6
25TI5CZcw333XezV/OzKeijwdiaVCn4G/uJClq1zguePcDlHPOt4HXY3wpjO6MEL
tPOHI73hSuB5ZGllPijYOFEKV926skVF22uijAk5GQD6w+yHFcACZmZ9tvIs8qHR
IDnMYBYEorb3slVHELRBoA==
`protect END_PROTECTED
