`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
g42wey4+pF/2ty+OQ7aa0Wa2mzEl/O75yB2GS8QnNNotUMGd3jWo8WW0L1AIPFLa
nC/8kqO+cxd4FLvjE9Fv0gSeTE30S4mEIIPRsmcy/F8GAK0vAOSG/X/1n/+8oylB
fUcQ0DEdONS7AYkZIkL0GkmWjkv5bRWAFtAt639Q/Ebo4ViyBL/Rz9h1H8oYWlVv
sDtEfp3Y1sRa93FNg62xloAOfz45LCS3qjYMiZD6yngzV+VBklTrkGiTwlsFVT1z
Gy5KmbSsppA+Th5VX/lB9krmzR7aQAPkx1jyI/GfJS98Tl45IbX8sar02iV+AjmQ
fGDDlqRR0aOcyOQuHDO9FLSxRPOe2Pc1wJZH8oLd/o37tt6xEFar1aiv5GbLxiib
SiDpFw7+v8WYlUdLcqhQRxkTjufaF2DepD4+YR20PutsTB5JbB9wNN39qFYBwdN8
KJCQNRLIQcKHwjkLqm9DEO7gwvnc6KPnjEFqUyUcrXdomo6oZlq83F9zdOhYK9Rn
eCAnikljxcj37l25dcaB2RoOa5auNM8Xzmza/gR2QoJm9HJ+mn0HnCPH48jJjTuY
w1W4epVrKotUffOXGsyi4yXeqrtUECbApQeQnAiwW1ypUb2GBwIPLcyYfuwGrEhh
uWYprsKJkO8hjK2Y8Gw7GNuU+g4GWbZx8toggA+0rbLFAe95jSEwG0JkL7hHC1jZ
ShGEb5vs8/+iqNfLPbVUzuhVhuruRFnbFb7glz99sIprfd7mFjDXdxQxWvYU/UYO
/GqNAWBdQoiKQ2MNgfVXUc4wyPq9dazFBm1YaZDxHyCCXZ6LsSn0+RjZKupGrV0O
0cZtyOlZTOmbNMqqqGzQaAgZc4ePGV2+2WttYlxE/cdDKdgIZn5lCtg0+6PfFahw
7PoOGit+yYlD4MCo0TvKA368id7mT05OykCMuXinh4kVPNo0Lu1mUHhpkXDOuEd/
l2Ar1r/flA2eeSRQ2v71S9pbEY8C8xVmq1O0EHtxqYXGOuoPW8skJ0gZUrJughS5
JSBWJeWo3pxTrYoq0uHtO0/RClDS4cmPiYvAkzAxOuwa4X1Sw1EbpiVCA30rOfj/
2LRU3p41cV19nxt4rQf6hFUXA6h6DDGZXW6epaxPyokK0+an8jvI+q+K3Pd0bhHv
sNtzVb7kGHBfznSITV/gcOK9wfu4dmshSYYOgzG/gnNqrAYkrWAgORwYin80mr6/
AuYE5fRZNP6m2wCEhvwa46aCzzFBb4Wrh9BPxK5h+Vrx0QnruFvRyrTal7GthlJz
llf6h4524IAITx/BaPNSxkjGIHJD8DsDdH4YhI4gI4PUYaSNOMTe6KfmZ0vofJ2V
JT2OC+T4n6+0+S6pHHJCXivoeAJnWNWtXb83shRwOcE0B3PNvRi/Fbx++CHbmBEW
VWI2p1eh2dS3GUx2OqwfeV/6mKnJp4hk1P63+XwgfuPlv1nlmruDgDqN7NpCUDDz
b29qpmnCM/3Bx/WqfkI4L+dL3TZxWNDNWyeV7txDkOR42qE/2nzBNF+DfEd+rlji
aDssAKaP1XjDaaD2fmaKoKYMbIj+zmL4pXjQJwd6mLKBrsWG8KpEvaIHJwwb5YlT
PAF3d/LB74YuCFBR2RGkRkvuMsBf7mBjg9cAJGzSm2E9ft7rN8z6ptcJZ40gILAH
84to/sMK8+zE4cEruY9mX9OrNTwp1lhdzACi9zT2TydQDf0R+niJOdeqqTQerxJw
ce4xPAPRN7Iz/t/mMZT2GNHbswU0h9Sxy+uln/VcxzEkEHlEAPUOBj1HsTT+eirz
2CKDyq5w65Hyi/mgAobLWp6mJxSynzzsMXOnTxKl0OwBq9YuqV/HXInbxf1FIo/I
bFn92eZAprFO+SAKWvLXrKkakUANzjqOkrRevAAqQ+m99ScXbMUX6I22jDWbhg6G
ztCKDY/HKdZ03QMRykR2EhOrbndqyHCTeP6kPQGjI7RS6B+sEf2Yi0RbCREdvyoM
RVJE1T3U7AD1co4HhiQEgAEzT8PRcb+Qd5wJY8o96+YuBanbOt1wxOYeAIwSTUzf
f8P5n9FPqejyuEROrUB8PEepNDahKWRQjH8LolhdRSUpDXzMBFVIlVJL/Utxxw28
8piYbkUzxOsbMU2QlSld9fTFAPYWL0A+OVmZoczYRAX+r0Q3jjWyMT4oKgF6rPkn
Y5vl0USV+Pclb3zVHdEu0nN6rxaRshwd+opGYa10T+jlPAYl62ZXCiKU07MCSqyu
iekfiuHQG9MlhuStiQ9fluTy5BrM4N5bfmDs23LJPbMPYHE3PDdE+5TuB5O6UwaK
QJ9kDRtwotWzUYFStzx5x0Lb1J++iGrIEl6kz9EUqnVddWPnGunODUlKOgDyQCBm
zA06/keU8QRa8zx7/43/PJS6Mui9/jf1JVS9oKP4Ew8n2La+tlqcFSe+bjuUDL5q
5X81aEz1K6bFyslb1YIv4jHWhuVa2VperkVswd4MYNhyzk1hTQX+n6LuNijMgiTH
5YZB23GXAqZFZF4molZ6fQotZhL2EyGK11AbgDZptbf26rWRCNPtH4d2bb4ogqGy
adbsIEvd04SYQQ3HCRQAfn15FueNGFTfn0vMP1Iob2ezOW+F/6CJzGVI/AY/G9n0
1jvrbrovdaRKIwgMzOMyeKry8OpLCfS3i3xSusrQL7CY8rnJsXO2OiApmmD8Rhpq
oXs//F1QQ09fPdqoH4AmcLfQl6+DkhXaGvewgFil8tlavrrRdP3itoVzCktS1ryn
AdZrWRCtdKQa2Yn4Ou9Zf1bqSneftF16P6FeZVfuaHgbG1jKk3AA5nxbMFxZM0TM
yxTD551lNWi/K6Kb3Hsn50niBKgdIFyUHA7NJItA4ijpBHQjfMAIMansDQk9UVzf
V+Sri5l8PLxIVbmyuoW5isgKitRKhc8ngQaToNkky0HQV4pS3kfLBY74XeZxIFI7
3R5DNtM4GO9x8h7/iNtKsjK+g5t/FOfgoxgkZTATojSnfB6SmK9KV+ojAe/7phq8
R70/fh+2KXVDaXZonLPsvQOX8PNTfcH7Oula2YTEP9eEFtbjQvZ/q0Y8j9HGlE/8
j+kdyWtvja+oxm4/q4ivoSXEXj9Ef9JIcRVCXG16w4mNXIarQebd20qDUg8RSl8k
OOwKLLHVn5mcyrlIid88uzjCHTEW5EzhpVSO7ENMYPCAi4mJ/9QRGORtMI3LHOXK
q7CPte/RI9cqNjeNt/84N4X6scLN1LFs95p10TZLrEFHLoiUjMx4WMAOdT5J1P9x
7HmEjxhWsxcWiu5kpfZO2fdQDf+GF8tWmvAmoET/9Iz1cHeAqru0oBEL1ssgiDIC
ifqgyToUP5Hxt4ZXLG38l1QOOL7OU4Sl2gY11RM91PsMnn5AbWWw4HylKPT+lLYJ
cFlyBhEAoShtd+uj/J4eLxPTX0vuuYDDNRu30a0eWCFXyKGbG9nSr9NiekHgd+zA
97TrMB8CzJ3iPDm+fi42w0UYXs0sOG+fuimSXFM368PPQN7VNbizCwsRBH1wUMIT
f6TLYbGeuSzDhkK7HF/oDDo2Bn34q2nEBlLF6KsJOjIE2YQxnvQobLDhPyQCbE6h
L1SZ2BbL5YtmypYOLFD3yueh5QGvR0nkeR+rbmXmJc+NNkMbrmRBeRxggwXHUPRf
wi8toYhnCy/e5VNVZwJ6jZ0TaI98bqSV3P7uiR+G8PVzNeGdI+y0BK2O4jfJT/YB
`protect END_PROTECTED
