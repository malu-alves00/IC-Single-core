`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mRx8TKXTwRqLgnDH9JdZ23jwG6F888H2MVC3x34wyrR+wdsQyGKtGKcWWS6L2A0R
UK8svkA+tmkn4JromlnnvUdqMaiCNuYvT5BWuWYHbe64bi8S1AEqkhs7C+JYL7rn
8ALdnwqL2u164ILmJApxKTx21sBrMyFvaFHvms+sK+EZ/Ij70xbi2u9m8mn3Agje
b9cgE70O3Mt6v97uGg4piHPERGFTpLDV/Vp9WUJ9ncwZVAUFspaXUbI5Xp8fZJB8
4cGAufUqkzjobCPUZSkAn2zfm5remk9N/udBTp7G/Hhj5gjdLHOLcOjc4QU01RfZ
19sBg+v8hRSidGD6fGVlAHP81/hSVxOHo8t8jYiFNw91BSL8Ty19JHv4Lr3MoVI+
OJxxZN5rMTXTOBtAvd49+QAn4JWmLVmGkaU9zaTniGHeYHHaexLIl2N2/fdvVVca
5d1ubsOIaPMkjABoK/A37G8G91QB/psrcEU0bMNMOYAvy+4YaparWDz5xQkGbTLy
TMCvSwwcqDtdXLK/j0RK/lSykD/cWvC+ajuIYPheSkcDKWWlWdufx4FfyXYiH3Sw
nf8T3nwGL5x/Gf9Ds2DdVl9i6V17QmNzfBwCRqv7NbpoOAugw4jb3GmIxtxqbIsD
CMNmG4CL9Pr4niCgZNEQPoEKvG40dv5zJqoBkoaroPUBgTIbWWEWySg4ZKYIWRQ9
1PDuCbUDFQaTkywl79//zzZXWwmQ6lluhfqeZ6mVTgs9b8bTQkiq3uet9fZ9YCbt
Rr8ZwcDVq8jji8w7IzJ3y+PEY0iYB4cGNGplDdvJvkB4pQZbxm2CqwlsKTpjHMeH
aaj+6Ob+dDzLJ1ZQPqkDPHIuGln0fHDnVoOw9btHL944dGEqTeBunGy3LZcXaJex
M5+pvTLYWoHf9PeFzWGjtW3fraYLrs97aRQHzzWzDOWnVQ3hiQ34PEzzWvP6FpHB
lrG/vEeDLh07JwphoS1uvEeTxw5BwVjDgysnv+vqqU6H+u6jc2n4RSav7e5EF2hH
`protect END_PROTECTED
