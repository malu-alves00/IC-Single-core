`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
abRrd/d092PTv9Mrff1bQUBqz/u3ROAymSiUnDKDPBYR4TP91IvZbawFYtdZYeoC
36xiD35q/uQCeN1KDmq7Wc8XaTmnI27ZyybBt91eYyA7vd/mNbSpVRZGmSb7vNEO
7GZ8KtcAzEuVLf3MB9wohXpMgLGs3fS3A+lgttOQ6rNcOzAAO/fgLJPElTnkltY/
VpBjA6CfodHQCGiDrS/GAmlemnEiJUQ+FofvH7tkfBYmBubHdcLTBhH3VlkalbKI
neAxb7ruZGobOGExc2esZ+n2TB+yGXk23nOGONFlE4Ypk2eFMmZE7jKwEtfto9kg
l9rQa9wDkKo6QD8tXrUDKYaLmtvUptWS3scB9f5T0eT7kZHXGv0yIo6FLJt4m5iH
5aikIiQZS758hEUAzKyJV/TuHfx8uKmY5qIrF1ku5DsNr3yt90HFZ4wNPge1g4cj
t7VcK7PML/1JdI/0jS62ZI5FxvG7uQB+EnjAlNp+mINzhsi17GBZAVdFoESpTH/U
MIIqk0RGb98zzWGq96rxLQ5N6lJ6Iz81uX9sfnvMQuhEjPaneyqwuK6/c7W5BHLA
FxzJbRWZ3LVlMTKyRv6mMghXHYXqrq3lvl6nsMG9nXrl587AqCLZlaw1u+Q2xnf5
MPt+6e67IP+fi/nyzb8HvMVCauFvN9cgaJ2ScrnhlS548YBxMynNpgZD8s4FFpPo
JLlqzeb4QuIlr9eK5yUdtlIvq8LVVe/7JRTpzWiryo2MWw2XkJ/xbfnbjyfyJmgK
Tr9Jh1ehs/sIPv6Q1yFkkpMh4HnU1+icL+zW3FAyDBMuTeRNa8Dc5Rb67kwVgPfE
4UzbNC9DgrLTR1Hzuz/AH6E7eDhpWCpqbEwKNbDolslKa2vkU3Ve9J6O0pGdIVin
NL6z9dTW5Z1tc4cdlgXksm6fLDhK/Oe4bsO53tkLe2Hgel6USa23aPZWanVN7go0
urc96RnPC6N/DWqYCzimUoK8igeAQ/VnnhZOy6Pf5w6y+8qcOdd/rpeglzCGQ38O
bDgs5sEygWshaKvzEOe+JlB+XGt8F7vcHHpzR6JDj7HZ3Em7W0bo0NwIeDiS0P4+
ytrflqXqCXKpqAkpptS6S+12ZF1RyVLqChh6O77j7jXtJ5TPsE/5EMpv7LB+T8ad
WR+E5TCIEG8G4on8nHuLx80LbIve71o93yZZSUdEE85+vCGy1Y1SFSnJyQA0rUbj
Xl2wkxpvlZ8NwsYLHLpxZXCvz701rTQIvWZINalDsuHx4jSuCDcgcAIElbqaXeLs
dXzxhXN5TZuvfTVzFmZ7ig4eV7WWBaOgZEsKxRGB8SGMNZgIckgYCOib3tPDFJ9I
`protect END_PROTECTED
