`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Y5/KitkFUTQP6BmUqMMQqZQzVPnBX99wws3Jffx5P3WoaIoWBkEK5SGIWa1ChW7x
7ZS46Ce66h+jin0vBOuaEAvfpPMK6jJp7JT2a92tv6lbX/UxRDEsLKdI8hM+6C+A
4cJM5fD33Pij1VPlTZ6AMEY2A7wwyBiefTeime8QQiFiHXK5TXAJFa4yePf7Wet7
svRDtmwUuZYuHuhq/tETUVDXIze1g5aCFPcn8+Hc2dnFJHlST8717lvtkE/86PzY
8viWLKh/S5xcteJ0XV2WCSRVHa0ts4796xJRu2sWrWeTpI0c3s04xDcYiwRYCV2H
sjpbjNpflKq0kp4Qrkcg7yTCT894jREkp/LR7a2rnJUxNXWP4Xghi1UtqlgEdOSY
IrA61WM7O1Wm2UaeOZE2SDdEumnPdxE3KyCU889rVChVG1GBPqgHGNkc0okocyib
rJSvun1B1ErRNxHDdRrUdPH9FhRS7OXnkedH1oHaiQ8NrNjUZpL8fz0HxX8Ao6bL
kz2eQyM/0DHHZvIG1DIOOE656Bih+mUieq0Ka3Famxzu/KF7JJub1ATmMimnocOU
Tz9U08BqeRW941xTwloLCY1ymXZ1n8U+i23eIm3vece2kKMEnUm0loIFuWm8bG7Y
4+fV/dqdozHISpI4I3JCS2SaZ0H3cBE3qD2LXngsrdW/s3QgA/qGNkhJAgJWXyHE
htJlim5WSwXZlduq5WZKgnhAiE2dRlIU2QOlpzw2PEv5p0VKtFP6bRyxEzYzVO5T
NTuilFzGvxZdgI144UVLrXhuj9p0NZoS68nDb+i+iaAuCc6jpfaeM1Xo3cRH8XI1
3Ep54NtFFX9yDj+va1p712wDVXahs7+MIDd6J3WEYd91tk9GUPesj+Zb+1EtQZAC
b4uXf4T3oI1JeC1HlmEiEqLSFLl+jL08SNRJnGNPiIZRG5e15vfFmJ2L1Ex6yRUq
0te4aLtIxnJg/tVTa/OVxz2OTyy0hcOHq5ZSDwm+m818mChORkKy0Q56GrzLPOxg
OzvNKIT/NkfXunEEY9hnfl2RukdH9N0ngqWuILRoRusc1EnMYx28jyYd4rEuUuVk
Lhdcy4Ok7NnUk/zJfHHEHbAF558jvVTOVIRqt6U0x7hNPauRX8H/DLxeKpb5Ffq1
idIXrsz1fxPX57fHCYYPjm1Fsydcyr2KFVmI9h2QNdN5vz1hzY6obXsm/OE+DWD1
KmSNOIZjTOIFgG0GG5PEJSf1azCmx4UJ181P0+7unqx8gdENUSc0Qksue3R0sDXh
HLIjdsnzyJlpryz0KHkOOGsTrgLmn5OYrJd/9mTWiWzzUcKy9D0afhJiOlZdi5k+
MK0tInqILBydFunLgH3yv3dhgNpnGwUxR3r9A0DBL5LOW+8GB5GnYcAZRmtAKgGO
9psi4XTAFrGZMogbRDvcuknukrZdTYgIe01MgchwWlWUE0VgvECHdvKz6BuvOQ+o
ngYKJ3lcTcrEVxlt5iDe55bPN3KRtKFv5emQe4Ts1Zc=
`protect END_PROTECTED
