`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RG3vtgRxME/02mmb2ImfzCFRHCCAQjSCJJ1fmOz+5I3HPcBRWeLcX5cCzdntDDG7
ypxGyu0MnBFvVWGuazL7X6+n9G9canx0ayWDScySkojPMUbWfdqLoaq74stzKcoJ
47IRYSQm1zcatiyleLMxfvktRh9sGA2AATC1bF0gEQm7JAx5skXIjkje1hK/r6kA
SI67ai1DSu4fP6375CIRXf7AoIDiYdWjgGi8kmBALLCeVuRqKnpr3Du87UtIHPfA
xide6QheAwKn7Mpyn3KGRWQmZe/Vre520Q1zVVf5ynFMM3N2ma0DSmnSDUXtvBZo
GohKvix6aytnoXA71LSoeg==
`protect END_PROTECTED
