`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Nu9TnTrDQe+IYQSK5+XYUlobg23o7xC7oewTWl82CkQu601p2DH4CUFOm//zzlak
q2bnwamSmWtPtgiWuT/G5hm7F0sQzS+y4aKfNimpRnHeeX9IrsywXpbs4IXtNW+e
O8Jef1SgH/g5NTrabAo8FdTflSHUH0yDO0QHSfaHlIVZXsJSGCqnq2H7d4cT3uyr
A3T8aZwQUt//kTHxGX9tbekZDqw2qGLv0fUdMe+rZ4D4+XKCyn0vpSRbyG+6TsOx
UaiEslTEUOWxq+NXXp1gY9w+6dhYiFwLoCBPxjq3OxinZJnxYuhTKaFXoUnfVDcH
aOZ924FroETj8PvraiBuvHd3x2CEQ0v4+CNaERaSHzjwVFDYfu2UCyu99HK8cYTL
73J6vijkk6O0HPsSRRbyfvaKqtIEDOTUuCWfoJzdI8KOl88ikDRPVBTblLKsGdMI
xx4CzrEgZDU0p2wbUuRyA3olWlUEQtrTvgFmi9p7vLXl+WrqWzcsR6uP8XsTuIfs
YzsifxHyFVHxV6jHk15IM46J5n6CB1ACZ/v3m6b5X11cPoc6rJU/UWqpWQGoh9Cd
PjzoC9CYoSE9sU3WSkJ8NtxuMVbTaZOTTcSL1GpwIfUZrIek6YMqqcmR3t2CbvVV
hpZUrpYnyx14ToZXYThkdiITcoBlRf6Ep9jE3CIrxmIRuAs+RhS7zS9OFbPrZQ91
6BzYA/U5q7LeghQOWUQBK+SO060A7QCxEDghodfVEbfU7KA6o1vRGTMuCljYdlFG
YKa9a14mttY6J1pO0/HmUxdGoRKsVd8xHHMyYfzIa9g5KRp2GX4PvB+o1mHdTamU
hKfuVK2YBpV8mtgvaxckhFVQ+62KknJuq5BTx3K4O+yT9HgBJyW2fjMMgmAX9WYo
4dvqbxZtkWzdC6CpYvFXZ7QLjj0f3QxsuECbrlSR4i5w1biHmcfqA7jGOrT6KjEP
QmEnbd8S/3nxon7P4zAgwYjMuws53JsE2pA7EueF/8lBr0KBx2dZ+fQS39HlVZhy
7eRIPRyRgFPxI8yKt8JPtajcRKQIhLpcmae+g0dlId6nwBkhjnUSfVpqYc39uK3g
E6bFAGWnaQXTqqxZN1VOdOEIAOBg6hdckk46NBRnGIkX3Q/dPlLfOoJADBUusjJI
/K6d9enYPD9NQAu87akihurw0/yywUsUXMOz2KjE6XXQ4HRzDBIMp06EyXKDPEj/
mY1f2vozJYx0jGIaS4FkjAHlqHSDZIlWMVl+peJA8vac6/XRhNMZFm3YwZBMlPgn
VlxNtBrpZ3ee/Hlsvko3EpRRrMLS1TFDWWdRHDbfxNl9PPDARXey2uwAkBzi5kkP
jew8b5anJTVd9McFjB5itZYRVifKYHljK8BM3TJpd8YznmZ1aCZPk+nzlJChhQGi
v9EoBztFqTNK2fuEQdG/c7XPwtSwuHBFGDa2A8diILqE8MAAeMRhukq3AR2LQXg8
jSBGPwEtpi6C8HO1BdDPkEAc0ogNsP3lUv/sTrQ14KYl+NAbEG0/TulWcc8vBpog
d9Y7NExwEUegvSET5dC3sFuYVQwbXM/y2f9P+CDlDpnuIO5RdrR9xnVMBvMK99z0
fZi9Pl9ccMGySInFlCBw0iGo6V32wSehDz7T/EMcW/OcFFAGxz+fpJX1PzYOOnxH
B+rvmzFiPDqV72BXLrvS2zFxhpL+tnGpFOEYjNuR8jit6FwLkodtbWgn+Q3NZ976
xHc2e31kB6NdkP9JD8ncLgqkHgvUvAemuQVrlvWyXq0h0aXmSjbD6mZwn1dlrkFp
yMx1mSy0Qkrjtl7tcerWsxCHwKZ3oshY0iv/QXZDhirh1SVj+1QClcJRnDepw3jA
L75neLmPgz/TmxD8hHowzEl3T1w79EL6nshxz90748/EQ4CnTd3TY5v71/wpekv2
sxdArX+aUYkrtFK/P+dDwTuJ7wN8o3se+JyPuVqHlsb7bB59s6/nl5i7SpUIj8Vh
0yJctlNAK7AllSD2x5Nk2bSADeuZV2RuFFtn+B9pDC0GAjbxynO4e9B+idRRpt1T
zByiX0NscLaeGFclDUl4rjLS674CQZDIFGKUYzknogw2tuTt5A1wcjWymsABOVcJ
S38FhuzRKjcEPnbz8+LuPvCmePGDzUHur5L1MzP9apiVoKsRl1kbS2Dwpkpl/94B
WCmssIDx6x4uFsC0wOSyetk6shqf2mNAfCQ42BfjNXEYLyjFRVDDuFmKMbHAvyer
GdxxbQEX3myh9ibeByzIHruOtUEhrFYkrVtQPyCjwtHQzjBvih17O95FHgsjuzRn
eOGbDxQu8HJSGSvOsH8k98YcPWrmXzXKdWB/noSllRxVTIwIW1chi0PDujyjCYZ9
YJTmMU9uKBPV4SRx9+mQV42/acPxBf6klIR78d+6YnqELv8sOHp0R+izbriwc85y
R21QCqP/NZk4NUcxr668cOa5+UG1BvT8jHduUz0lEnaamHrh/b5SSt/mUoylCopY
hCJWPTDEpNgRa6h5e5mwZE4EzwAFSYw+w2OnLl03inQp/tBO1dH3U8hq2UAwHKBp
nZkQumZjX0LYxzerL0Nt5NHnG79qDA25w0hq+K5pAwlD4csiub2BWJv1py8XN4sJ
/ZcEknh7J0uHZWiBdDgBrYdxxLFmWDtr3sWbemVtT/HU81geArP28Rxn1Ktyjh9C
tisHir9ZSygzitwwOTW7iphAa4fEP5n+GBycOD8uDfCjrkSOu1LJ8t2eZXvVC2op
VYGm52+jxmqeFVjX8jfWQwyh7z9bFqumrsnlesJ9SiEKUkQOngnT0e+ihHhPwwCS
1J5VeaHII0Gc++GJOj+Mr9HXob1WFEefC273hEnzgxrEx2IjHLgdUZf2Xr7WegHq
L4DS6xaP8eHHndYboNY1xiaB6dxzs5o8dlQ2KZTKxdmDPk8hql9Zy7jmrcK/x4z/
hygVBl5kcrerrfXFXgoWzDAbFmz8e2H24UqGV1AJWubkUDmcSojhhV58wuvhBaMl
lgCtZPHjUiKjIIuG42fNy8CJyfS2BJgxMYQ8mCNN1h/SOw48EidZZhFJa6bgyrNK
8+B5VJNwXGh3KUpKKTk/d0D0yI48KhzBr62PU+7lx+jdVbHBLWAdA/mxM4sSItBm
Lif0tzt1ioRAGgrfb8lzOm7ugVaQfz48QEkWGHkjm4bPOtKwwH7+2tOou0/EzyVR
5M5XGj2gPy6CIgwhgAxGV36X8r/XL7L3E7veRQ4JUvmFyvMXNi2/Btbsdz4xAYpN
RxZft46yj5eGap0LDFwy1v0dVJP39h6XXpOAE88G+aju9r+5Y8Gxpsq2fH8NmumC
Nw61xtEWw+imzoKOaT+4MP5tlsnGI7fYVKmsMZHOdqhpOQ5jIpmS+OtiGx6zkEUO
51+oAbkzdJzbL9S3U+PH2VjaCX6XRqd+zfLpdiwkZBV0njThDbV5tJS9IcnnF1xB
pJsDaBxgK2boe5101Rc4FJrOOyZUFyY6PXyL5C5kmKMwQ+yfNMGYdGuNDTopZE8t
1J/LbhFN4ocvf424F2mOlhd1/Vls0U5dRo6e5Oo5HkyQFX9wuhzg6fa3sNr6HmS4
r68XE6A5lNJZyridVGU1XONFH4RyL3T74/z7qiq8v5hs3x7Aw4LTeC5wL6u9UloU
czBKIXfSvoIomqmeybO+RSk1WYKMCPUS/A3sKBgRRRe2Nuw65/7a6HfLK6vx+H1I
gOMkMqzDPXwJz4ytjolDMe7q/K7wtfi3u5O4lJkwwhLbDnyJeJh6wP2rLN+uOIGN
yHtgzOXLH7SRWlSBiz+05q/Z9q87zKu5NKtIkoUqI2skHps281YhW/sPKtxdmyJX
J02FdxWlBBmB62RuLY7Hqd+LAc2tVnJ8gpOTNA2m+URvplLcsLFWYo5Kj5viEDLV
Nzuj/0gNq7n/0NiFBGwfB4Oe1MSkIz9ObPY+CywYqE+52CLsrGF2WxyO0O2/ChSW
tTa1kKm50aAgCZh6VcA7wcW7wH112dfiXzDrabAnWB2H2WK8fwAMeLY7jzZV4vEk
JW+aQOxhGB76ttBeDWmlZLUtqWWSnT7PR7Xe1tTbYBLOoUrCT8pd/MBesk2U+z4T
QFTfphrcAK6GKs5Qfuui1gdwfSkdWN7xQz8tBHiLsGG1HfcS3/6nAmNEc+PuKnU3
i2IvjnjlbV1yOkHFIxkYVLwRKtWvtGrtwUG6cHy/1OtvuMV0nscRLf4BLF4BHhB1
e1BHs+0KE+fdoeuZ0Wt459KPLOGQl/BPBmSRuQo1BFxV3ccdcqfUtXhO3MpYopEx
TB5l12RAcWsAL9nIQpwuP/QGun+biTui6/aR7WImYn0j5KAPm7ki6R+3LSb2Qyxt
Klx1tiYUL/oILzIZLGbvtVawsl4zO4ijCnXNSu8AcWIuEzKiYLAVVGt4e5QBWxXE
MRWSBkI9Kgj3N9JhXo8LpzzdSUKonK7SoSUOp39KJ9Xkml9m8iYQxHh7rFd3pAQA
HvjHkDkmx657CMnQe4Et8t9mn4DgmO8rSw4cGYX3cPutgL+J8zHMrJm0J62dTbyJ
cngVOu15GBsQnrt8DcT/3zMHoODlc558N800AfXZJc41CZLeu/lTsXzgNaQdKF0n
hMttFJ5MQlkTkc5kfDxqHiv4VLL7ya+8MnFo7om0WoqPZ4B6R2N85o4hfOSk1Zxr
UumJwqjUknFEO6hz1IF5L1AWHG7TLvTUoVC41vGpCgjNKXogkvxKDWg3byrsVXd9
Mc9ZrejhWIjqL79+ZLFVsUGiUn7hucSFN578k9Q9UjBVBT40rUtU2uO90EHOtr8m
ui6fAka1sdcJx9fferD8ge3fSnSTKQgM8OPEN7Jg7hJo7FcZv231C121luT8gfsq
7tzcUX4ytDovd95G1igO7mhkm0Ox09vk/aA7VnMmqyGmn1nN9wWbpe4SbeUFk+Yp
Ro2zLbtgCtObl/95Uj9w4nCDfmLHvSco+GbTKgWrfB5Zrr4gwgg92u/xvQUsqdrR
ON/frV2RLOgeWYMoAMrQqHe+vh3NybQz2KyqREekTp7B9aKzOHkybDO5ywRz0zc/
i5IuiEZeTYfWxq4yQ8N09+K67WhU7PAaWJVCC6YJXPLseQfmv4nAM2yMzHS0190V
DB3NrObSKzVoUAO0+4Y3GA9xwmRxwowv9zhshLT83hGkJFm5qBYjoRduagh9LKFF
mxQ9EefBZWthDkzk50FZCR/h/xPeyk7QCRc/ewXCfq3iX4R54jeBxohOqNrrAlx6
vLHJ8CQ9RaCVjyfwDgrkmw75d5W33CDGCpcxDqzdP5NEKNLjzAz5mRbDVRQPE3ZK
mJ8qzEcqfEC2PSqYNiyg45Uge7eIp+24/I8eJIPsneiJ2PlXyV9704PBMT/GOUZH
JGMve2gA+o164JxrKI2HKC1Sb+NQwebydr7cy8RCsxEzNIV6itpSOELws9pO4gW7
zt33d5hXXyztKBzh0bVqNQ==
`protect END_PROTECTED
