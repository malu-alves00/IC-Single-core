`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uLJzCByRzDnxI7IhVFxjzRBnj/GyKA8Jh3gTkCavTtOMgmBDjfutnFtWV8TCOoz9
RWhIua88YsQ8rMdgkJFLF02u6AQOxq3Tk9Ognr61Sz+/Q6xOm7j6aKP5+RgufwAI
YKkoM7tb2F/vUewQKW8SR5jNW5mKExuM3rnh+oxUXum3ilN6oWFZM0Gn06WGd/QF
rBHgD7jOChK/taC3iFVfaVTANDQ3sFNbYX5qIZf2TtCpXK6BHo8gXgCz7BpxCrAN
w8wUi0cqhjkJcCnbc69nuFnmqP+2p2CB/br41J2Eq6Mnnkekj2K/2Yej9E9ztUu/
QYQLgEtOGouZ/OvtKvsGAn2z9PoYWZV8slNPtoMYYZalzPG7CsVssRYBeld9rW0s
c7CGxfAoEIDnUTft9MDUJ2pXHsgkvf//MnSPR4M7ZcSObZhU9kU9zbpaS8+pKT9m
OqcWz4SXWrHWyu0MjCg8FCdhpm2z1DmOAuoeFCtgzHupVZc9S0Cc7vuTZOWNJlVc
ibkAFwJGD303gfT66Bx/olPGLpy5jxUSf9Re7nL5U++o2hDvMzC14u1u8adOYEbA
YE5zEjdqVdZw+5SAWtJwoM0HnMOpbA9GxGPcLwHNoTvPF6mWaL1GivhHvBpItanz
fL7pw6hiOdqWdvEhedilxIpb/JA+VMpt6uYkfSwfZ0VYb59UPsdv4cAjB8RQi3WM
nmt+tMZJn4kY6AkEIqtwu5GU8ZlLYiOsulf6cuJeKg+XbAi0WSpffPtxXbPPRRAw
mfduXAoWPNppN+tg93IWTA+LKvLPJzyb5IrxRr6duaujkivKIG6H9b/fNu/M4C6y
DM67joMmKQ7UuGs+Jg4sZGRjGlWepdogFrj7QgUBl3kYc30KOQ1VwEfz5FA4IP9y
PaAl7PoBQWHnXZHdlrm/EVF0BvU45KuyKKp86gQzG9Au43JWIwgJUloExA6pd8Yd
UXpN8fmnkgtv1PTQJCJJO2bR6yhH0vqUAg2gkVjGZ7vBB1nQVyD2P6Jtf4jn8mtc
Hawgp9aC5nfjU3fnlE82ZCzr59WHj/NlWO+ZQI4Kx79GBXMxLSVup2NN2VmmuCK5
9Zz8ubkHAWLaZ/DAJF5sdTshbCwjBbtzNItgJDrTepd2tYz6bpewCqS99Ltbbko4
Txja6fDcJS7OjElqAdbfFz8JBXWYp1TS8rvvkSOTNWpwfPGA4tOV5CJYtvhtt/x+
420ifrR+oEH9bRUtX8XnuOXIx151VTC+NBC9QHB1NOdnlWXu05wVJp2XGVH/Oax0
TXgOrKdayvcw9XRgNTO4K3U2i2EzX35jl3eBdMMmJMzoYG9qxK0QYN+PFV5PlGKR
bN9E39WWxNuIT3UUZq1exLpDdBhwRs0lawPVA9R4trzRd2Tkmvh7Y02yul/i67/D
zX0hJj6sCg8T1nvN5XTu9cLcW0c8Tzt/hkOreOwEcqZzLwSKmHwSButcdlasnAMd
7zE4pe1ct8N8wb+8N6kIvU0yk/ohym8xH1DwhT5ylklWqOg2HSFyouxk2HupSh+u
powTRrj/9oBGx3VE9H1JtGnnhU+wDDmGsuipCiwFcH8kdOqKXGhHiV0FwVhp+rsK
0MtKZn0ZC4jNJWupQPSzO0bGqVmq/z0rub8EwB+8LLd/+QeTSC0HaMVvF1gabu2D
0FZZ8wtGRloXrMn2d6RyGXWvvim17d3E4IeWJ5PYwmKg2bddeKiCpef6TaXOubAw
/FQajMZAmsL77mV0wDAMnC2r6wzJgf74YpLPE8EJWDtJmro9EeHVyMrXk7lY1hir
HwhPU6jKDG3QUWqCvSEyC9hXA67iIWc3RQehFJUbv6ho388LW6ikeYy+ZWGuQxcI
Qk9Mp9fGxdBspYakBT6LpUSPjGdBK7mH94eJtFJ594op+1akr941cXv7dU2sV00e
WZGP92WDal0sByUqWY1+BJnH//L5pC7IXN+N0ir9eFPghDtQASyK82lKSK+8lqD9
23EB5DnYkebC6PtT+FJ6xFyDt/3Rk8rkidiuEdxtYNpkeZ9zWUR0KOUbKC4nURl9
vZkrLb8lhNL+JVHNrKwBEKaDN8SL1Z2GvwqKlGh78yCJ6RGVuTIWqKL47yRTvJZb
U8bAhB3MRkpz/HzcoYkDE86UBNteheP55fvPI5M0SrEDC1jgzmur8DhmHnB71evQ
nf4DGn7bDwvc9RcxLMfR0IChz+69TcoilDDz9Kda8+D35+3MYHV4HSJBJp76Iv9C
NePNUAqC9sw4+jtgzb+oxfcHCcyVnVeE8mTFq5IWxWRRIAjXMHQh8TBXoT+FE2vZ
1PfTP+cjfEKnn/4WWO761WCBG1z7U2ykGDSZAVd+c3kBPSCudkKbPz9Hc83LG1eN
fSttMuABbtDmM+5DZqI2fdj/G8UJRn0zPm0j7RHerjzSMekq/zlE7dyzj6knGbL2
tl2PyoDTtjnDH1zpjicfeNamts491PctRzyvVTMoCVuRU0SmhXHhSWz22oZywFw0
aQGKD5+Atlp6G5LHuovtgM5LZURMgjqQcnqblkoSjam2yi8cLHihjBa1vF2FGdG2
rpryNu0GgsI+7Axkwo9FGm62USpeZ0MzZshgLubEQr7Eqkza7rjgerEYZeLi5GBM
ngCC2BWYsX3XTV6goCuDj8ueH8lwFUs5uy6DDi1ko8yvfHuPf+WwFFBLxbxC5zCs
UCrbqsA+C+Rbnq8MCYmKS1A0wnniFP2XyknNPeHOwKXZU4qtAl8tJ83+v2Xhb4qv
WTVDBNXjPMQWUQ4PxrbP7gPq6IHk8fgFZY4NGKwD7rLnI7G+LcKuUvAv/CX+GIWh
TylBgWyOYv/rfAIpRFMmVPmjRtX7ez2E99ohwOJMoKy+HzowPix2sA7qLOvKBlyg
iD9zfRpS6CEfokJTBse7CwHtyc+7Ey+Wwpb/DqrbTu5712DgWP2OnTaUPzVJ+C7d
lBr6Am1+WPw3gWsQhfS0E4I+vOQ6MJPvWbgZSqErkQ//8r+X+4gFSFwHDcYlJK1F
gEp+S31TcqnKyEWTqQHzIsjWaI717ltO0JdLvtO+Vv+BQMa9nTkHlRkAT52zWFLz
Eq4SVI/niLDbFqlEvxU9gmYWheS3qGekrwNn7XR1grj4utm6oK2iLvyOmB3hEpvm
RTyWetoZbq0TzZJzmW5zmx9NP+NBLXQobjqfTX//eCZWYzv2kBU5P0/KAMNLYxI9
wpVZ6lmmz6626LuOmsrFt3drS9kL1s7ZkuZU05qiqrS8f3NZKEVoBXNpDCndLtKb
vSP2lTM2Pl7bUNFjZEBzgl5p+ZtEH0Fi8CCME5lEslbYAIHxbW4w1Km0uBtc1eC8
5nowfFN1LIH+BCjr40X1Pclv7uqWJmUAhMknlhyubntxAH/Y8veZvcoOvH3GXRHb
81dKIil13/GDpnzIShWEDPVcK4dyik5gaBB+QubWcEYHpNlYWdtoXmgNHX2DbQlM
AjZfuH6j64jDnUmR2/bJdznx4hEzyQlMLmfom7mPp/WueEeSShprPXfBPtQFvJZ3
bMFYcmQVB7EALxcEyZk5hqAshXOUNzZOoEijF+W7pVyGW0pfIFWOuT24aoQ48nRV
Shx6cf81qgnxg+PGlss7ClREjV6JxDmhlmTwm/Rma6+kf+bqATkdorhkCd80aJkO
1OSNjCz0A2/xPvVMyjUkwBtV/r+ayj2qEe3jmwiIs59v+sdh9znJ8E0uAAr+cMvC
5hJJZaBqd63zc9mwx2qPP1y7tIgJqxr8gqPWePr7lLivWuhNpxUASMeEdATnsRPm
uwkU95h31GzdWsG5+69m5S4TCEuPEMjvWVTkTQ8ohfsLS5mx3WYO1zUWIdShqLTO
WzAHg3yVNUQ28h+1oQIBw4kLqUT9zJ73AqbpAvTNO3KrqvTJrpGwo5MbpkuvkDXX
fmkN/JAR0ZuUkz+CZEhsDAyHcMeancb6vrzAgDXv8S0lP98O5/Lg+W8EwV4eK35C
4ahHBo1p/QmPU+m8Jtr3pyjXAxqgucwj7R7Vahb2VpwD1xDNBKQG9IIq6uYHe94I
UPHDpuTLwQBUQAvLv5VisghkayFJA2gQuNRFLEdsTr48lniGt+KCAgjRKX38oYOK
oPcjDEi9fzMrJQ6nbGIpHEXPHS5RnZNptCZPUk1zQCE4XX+yc1XX4x6dn9K0xL8E
f9S83YsZTogBStp0Jj+kI4hN4CSGu8mCQ6D8DGCABC6SN6HprFJV65M653kuebkD
MSFwJ4jBXpQ8eqSm6Vl6Nhm43WJgArpr3oaUi3VvLcZylfECpi912qa3ctZdS+P5
`protect END_PROTECTED
