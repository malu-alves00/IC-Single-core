`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
s3eRaBhRaoLIAn25cbfevx+2jFLbxKsO4i5WcbAk8fM5BYLY2IuMTksrw025QOvp
Rgcwcb5z4/YH2QRfoZNwWAdBfeuniO3f404TJWjqBUZMyNyPXbIyV3gEZ7gulUsI
4zk0dw/MSZLctrbHhB0J7kTNQgXQs3b1AG7scd5PS1ua/ccg4QC4gvk6zyEdNUL7
KZX89ELJhOeI60YP28dSzW8bolszeLepa56d4n3Gfn6C0B/FgUHSWCMWIGg3eQBm
PDF1TRnypKuVoLzgbSBfieQHwOyQFAn/jyvLr/HDfjbCV4NfL18D3uYnpVv/9NM6
gTTk3M7L4AXK0E5MmjMNNWqTXYo9zaknOlbkFRICS5wDcaPAxYKcPAecDHQAkFBv
KYfheSpZwkonibVl3Ka0HBcBMf51DuWPuD1RBqmLDbyFdf1o4jm1ywYK3GorUZI+
q3XlwIVXevOlYoMgmxtK97t4Xvno0eFRQjhrSOS/UHzv/4gVdaSL3tvG8NXaKlkZ
bBk0Bs3RQSqlMul2B/4E8RnybMyXTMCVsa1JdIbGumWtZWniPIpeCY2nzoPYex7L
ccfuMNiHyKg0ssAo1C4V9QmNmXphyC7Z/R0YwzumhQBTJInpHED7nPwhGLImmcM5
VjHqV1JRB+XkZ+S+ugS0hhNzr/lShrV00bi/n3LvDVdAEuw+i+Fi3zFshPONIF8e
c2120EF9Ae8A18L/eew95NKWJ/KM2PdLPJ0hUcYJ39d9lvqVsKu9Gc/sCKp1iocm
O3b/h2W2mBIh5xRgcA3u0PWJ2FtO5xmquYTmdU0q93M+y+nftw3p0KBR21UlePo6
YauBG78A7xYdxo3qVJfAUObEBAKqNN/nwrnzYumnprN5NfjHXyu1oNeW+45qbCHW
rWx2PNUS/p+HLKrDkvk8kg3FYfAuWMp+bl/L+uTY81ZZeLkmxO/V9B+v9IKV4Bc+
ic2KRCsLDnH6/HmmHysxpWQhTGdb7vDkzXPeQGD1em7Ra6xhogNAB02TezcbXfFN
azpSvdiBY82GFG0UVt1UPuiXE0p5oGg7lQRxxdqNmUfYMGDvSO35mTB0eU2beFAJ
BwczW+syCdq+FqhsvhWVOqZm7fpnOl2WPozP8QtcDJJKD6VpXe3QhOJG6weyvpxR
zgXR7nNEXYbBIMmQNTXyCsGCNeNM0Kl/oRqEb01YRYnDxSbHR+PY0vo5/P3KPxmt
2ZAVsxutzzxGgIMALFYWJoS7LcimMdTKwxnvhKxtmzfrTIIhgoBa8lQYUBvBE3DU
W4kz1rhci3vU+ICIrvvaskjSoA18YSBdOOmyqfCam79ON4+TSM+NWuFDzIUx04VA
7Ou8YZDtlle2hbSUiyouszWR3pOLWiwQoOVvUTMP24abs2Kq95W9fZ0Qhvb50eLB
Z1xJCII5js3pu4R7CfO6VyLVQat5uyUnleTEcXSJco+amX7qeWeh5RMtnYnZ/gDH
FlS3YC15e4f+8EfbioW3sM8CteBAZnt05ExUX/i3KPImtmGADcYkID0rog0Ox1pw
G2wfmU+Fha9syPT9p8sjg+Laq7oeR1t/IXMdXyqiBJqzq/41NS6hWUqzVMQp8uN9
KN0KhagHquxwN0P7su1gBJ7UAGYYzsKgudlfqBT1ec1r+g54dMQgheC1b7i4O+uT
q8swJcdbqFYm4PP23R828MzdQ/iD05N4cVkxmNAnfIDmemn4gJfUc8ycbDS5B6RB
3q+gXGJTnBJqeqkrz8zLJK7wg/EWk3adkGXY5R0thlcZUo5o9x8smaCF26kCNhSu
U5Ana0DWJUQLnOfPcvASRWwt+l/d6ixiDjGf8oI38+VxoAxAxYuMRHDglEaifwt3
Cr9ANR3nUavJOO4t+TsjUdWzNyX8gCFLJHuAdhl9jtqQGDYGxRwHs3w287zZnHm4
1Dnwh/imeUuCthpfLrc+EBfytPH9G2hGuVIBWGyH2jbuNuNqmQGr37knmK5KVSXI
HGh8lNsQ8xR5aRl7wsn0tSefiJjduhFNmD5Z4rJ6fNeTaxfsZq8bzFMJZoi1TH0e
FbiIuquJn8Aw9rS+XtPWqFBgsHe+xrEiXxfy2+/TAOvYDz+fgxf8bOPfojtw+3/p
4Ks9q4GPTw6654NmBuN8vcl8MAo21hX1HUgV509NwEUbnB1flZmUEWEE2kAvUU5+
Vt5psUu+jhdI5gZ9VXeu1j2DcrEW7976YPIGju+UvESUq/A4QiROEa5CMGvdBTjA
Htrc8rTfTbJnZAl1UCaVLD0DyJ7MJcMrkG0Aqw+59m4Ntak+l0kzbGCyeILYmeJy
RQLhrWM87x46L5AykY87EGtuRooZcFy5zDXeNIbJpkLw5PTBTI+Io3y9UtpmECEf
vfFVzmZSWMyT5iV+H9rkfzAqRAUOuSRkW/w3uO9Kj64q0o6NyhaZxI0bN58EJPrk
RRFT9CwnBAt8NzGOfmTfvxWGdePtc/UHjSTBHQl8YfHF/rkRVrXfsjINTaWB3+1W
E6GYW98AvDpkffdkem0DhjOz6hogUJtf1b3aBny3rQ0h2r48R0OgyOXjYIdXld6I
XrK3oAVMukswI3Pe3p9wXqCpe/zzFGaEGLP+PMIyjRcitBwVBGa/xliop/afaEU7
pd2tlnGnOY5Q1XB5Dh8aFjN+8VGRS6i0j04vnK3Xu86QVKds8cS1gKHBOu+8492G
6mEHe2yfcXFyPjHf6Amae9m0r3H01+12xUdyxjSz2c3TBhiQWDmicbn4yx3LESPw
2pbqqo1q3FfieeFMSToRy1Yb9AweBD7MBUPOEr2W5gjO+NqU0Km5sgyeWsdkUcGr
tpLcjFCMDSD+90AXRt+s2+Xjjc2iaqXXLjMWf+opye7kSnK9d0Jc0b0qMrFlFIsa
oCYeRhhTKURC1ZSX0cMr0Q3CK1EPi73EohTSWQrcMfCbrygftofIwNKngxejRG3L
Yh0XnOPTjpCckmXOfRvdoMVPLBv/dAa8AaDDA8DglkGMjVPlxwFtpakLpK6xCzNZ
3YUqBcaspwq07jZDK0sLQW2jcxvrCzoNuqCUYGqpfF6CBC5xoeZ3zC4wXIX+vGD5
JWwjVE1hReoJxxazXYisH1zqjDxDKH5dTngZflJ8q357rhCL+TuzqjKYnW5OwtJP
VTMdZY/Kjy97/s4qGI30Zs86MeCYuJg/w/ufBYDroOnF0vabnxpP9f//JHk5SEQm
LAnm7zrFG6jAzGbH0HOlJIrEOTKCB4hbkG6gJsQBuPRfi4kD0LxkVCKllQAzKi31
LsVyYvXmzZP5ylKD6Pxp0vB3oyJk4IM9FWc2ffeANPFhw053ih6GDWIqAUvb0GLR
bEpHzzBx+sJcXEMkWcYsSF9Ut3mv4ml9lNc147FoG5g28o48XMthnpvI6hYp9DfT
q9U4cBjiTTWMyScOrrsav0o2r2ss3kofbeXDj8nECbO2B9oCYwX9e70YyxnbW9r7
P+q9nDFYriHGZwdynALw8MTfjv1k02AQZf6MWjChms9awmFdqrOqGENs23BA1PCP
2qXCnvMt/LGckNbi+6Qp9PvQ/xvoAJFWo8Ns+3+6cvF9v62IcL+XjdPO2ClCY+Iu
nVWWptglijXAN0FLUaUEg0vBSlEE7aMcDoYY1uVmOLCFt8lwgWJf/e8qgbcjhShy
htaeCWNfbbPMOoy6Jbu1xqNdecKCWurWLJDH0MF9os0NPbKnPToPP6PdONJLPGWx
BrNpkmZXfJXk2OkQf/MyTOrpxbdq+uQKRQeMJABBylAxaAztBOUq27iYxWBvu4Qg
ax0ToiRluv8M6mHlJfIEHfH+yhNdCHDCaVAmRtUUSf6WocLb3NucfnPr2l/n0s5A
js2wyMtRPkRY/UOlN3wIpiH1aesZSeusK7C4gpAF6quYi3lBf7EPHvyy2WQXw/Gz
AMKaA8SdwUeI9BOju2EqcOwIMzfJhEgU4Bz8yLcWGGQqyZ7psidjT20K27djUrHw
Rz0VMemgxhyXlYMPSw+YhNi+ck6TjKyIVwfFVLgEAzrl5ZgdLjMKMpFLS8GH7oOY
pnSMX1ndOlVMO5I2BPtG2eZXVCR7wL1jxyqZKqFFDok16fCHZqpGPag5hIBHL4IM
XsNP5cKbKNtyq6+6LdLkRRnSM/xqz5dyzYpuLL2WToKYvY1tGdReaipLkosJ9tsu
h7orwSm1O4EseslxVbUhJw9KYC5heDRkghX9zIa5kq4qhSkgnEJJ9GMfVXAaukdi
pRxKy5rHrj5vDLZXbGzIL/bg2JFPuGUHbTBQFaCXE4EKx/utRekwVThJzRRJSrAJ
bLQ+CUMMfwMhWvkgjIv8+robA9VnWr43SO+4fip4lK69q+K4zWCFNQiVjI8tflsl
1KCKtB7HPceJaYtCXk8AJVRVOAKnKzt5kjfd0YnUx5QSStF5vUZDiK9POyGYAFHR
kXOlE/af+XdXYO93ZswknwFyML/YXvLqsZ2un+Z+u6ANds9FJT06DKX3AaykrDoe
Ls0ojKRWRKpeIFBX5mdh5HIFwA+c+5jhzdy1FGc25hMWdnneZVDnaDQkNheTCi65
dSmvf1NZgaOEw/2ejZQJIF6PibT6EFU5GAl6SH2Hu1L8BIE5vORIcUDX/F58OvdI
3KIBoTg4TfgdIw78KWvrj92E/D+00dD8LUfcsgLeQaoy+8zeU8XNSagl+uG0qu44
gG4HP3ld1sEF0a0i1Ps6EbNuvWhXjokFfTovw9Ub6tsXpZDUyEUdLgQOJ94ASR6o
HyJ1qe6jPytnnc2Sn7ke5LQYqAfye0Ede04ARaw/JAJ8Vvw4iVEJMk+TDMaGqFQU
H7GUNrWGIKQ165ghbCOHGQ9ChjW20ow4NWqI2e6LPHPC+jVNrO2edFAJY740tcgK
GzkV0qeaFIPyqx2uUJ40wc9mLNsoJXVd/oyYN4eUbfCaHR1QjehNF+NCDedfGvQc
O1Of9psPzgT4UZPHEHcZrLOM4fpbrScVH4lBuYWZ3SVZZe9wjy1b9mkeI28HS26W
4WyFuO7f1CwFm2ie6tUKYgT7ZTSmgi0pDCRlFtF6S+3n0mQmx3UpUOjG0VqyPpyS
boLAowWBCjIceAQcGsErOqpBe8WWnomYv+hDBNZfC8oeqGAC9eP7ZX9UtckN6EG0
HGwqwqTBpWIgnJTosfcgDpd+kbc3V2CNANx1d5+CZrU64qub3savIc7nWpb5ixoP
f5JxKzdVI/WPOTADYR+swyUrJt8wYshT0rO/WKMO34nRf/60fZ6fVUucLfwJhfV/
3kRVjIvdGAiYvbdJ42RLhhAHPLWhgX/HS8pY21zUELcWH1vW6VW5tNEnH0jcKcIM
`protect END_PROTECTED
