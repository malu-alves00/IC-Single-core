`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XpD9hmDll6YiZnLLwqTk6cQaSLOFdxmZSeTDRn2TQQXjQKsfHjY+pBty6UpKibxb
NW5clYkl5xQtnTRxgqa6BgeexwNehIPCsFQImgy2WPhcCAgBCWLnGUiGzCqcZ0ru
sMY/SW6HGrodLQWxcP7W1V85i1fvEngeQp/T9MtJmpdNZw0v4p+Ef8xT3c6vWrAc
sd5tczJK32UM6fCMtM6Ag858KAOwzJMskSJ0/6yqORZSB+IeeCwoalkdWe0YBoCw
eWnFyvwdG3X8w2UcSGh1E/yWOW7hxrbKntFAc5jLbD1t4INYCcztkWa3LgegchpV
7IvGIO2n7kpULT5QNF2eGoeI8lwMlgkkOQ/ZH2/O2tsaCKwFXa/ReXjafq+xgvmu
+60IVyqxxRE0SqmZ0zUCCWUKfYVX0gQnfpX0B2SmLIUgTpeEAl9XMSEGI5xF5rat
4GLQHCNfEMwn+Asp5a5vvdvHVj4s/iDbK1eS4+220o9/Jz8xrFph8P467vMkn7hV
ljOIyd9JEX1jI8SYVunmebaZK5v8l1r8lSifuvyc4hapUmmvG5iV93gTKvsdRn5z
M1BRVH8nDyU5XVXqJt+kDncbi3VRhSo19Tk4T8niHRDtRDd71W9cgCn6WM1sPkFi
vQ657aZi9LcM9iswqDo1cc7B9mqRHv9T4GrND4fdH9HNlHuVMQELgOCNqdnzA/xI
Li79ccMRSCBvXQmqm4idQEu/y7/G5av3zQHK/15jb+W+Y0WQAfx9IEkOFp4ZTm6q
h4e+gAsacCSMnyj4liB+C1xkUAcN9DkpFvk2aOTVkRxL8Aja+AtqIfkoBeEHWQCo
l98t3yhSfXfjuY0hWbO77TCDcG8FSvvrJiGCpB3kRNma3uHRW5lYB+eKsjLCkYKu
FBfeJIxwKYGTpz3JRwVZ9DA/QPA6AWXUlOzwm5I5EGTRJVvPB/sVhOf8QxEiFeZp
pDoajkJVV5uEi1v8jpuxFMohyvC/qBsijFeQ9iA711wOvA1lECndWr10wPTre1JF
YFs94+RGIqZWGgT5F4/g8CgghPa6kWIlh4tGv6GVrBGpS2TyGU/ULSXDFyeW+hII
kMmIEs3GZCTtvpAs5KPRyarHnR5mYZI1FU/b/emURQ9u4TxPiAccDsoTN3mBHlyz
hJDvRflmiXqEVHTt9SqbdaYJfverzHw14U90nrtEPks1BzYRZ4xggDhZbx9TAq+r
/mgibljbhMkeWY/K79RvXZ94Z7UhwiIy691zMpQcxd3HU5mY0sOTydF+lwVSA8Ch
SZgi69MEYrNIxneHRFqZd/1igONpNAQk36gZb5HaRIKrA5kcXh8IixpoCSvpFDUw
IRi04g5b+WGRlXJow+ZkvY6nWsCEuJgL772KniuQiZqxGL0kNcGfD06876KXI5qW
So34kfzEpLZmvZTWZ6G8HfaMb1MxR2dymaEYubKIJ+SqcGxIQXDObstH35Dg97I/
L/esBLY/Cj/KjbH931G+blLt6tGsbOl/JGRMUUuzNlma00Wp37p34eiFHRk6SgmI
ldL6sy49Tbs4VpeZFwnM2yy3XlUJkiftYH988oZ8aX/VGx8Ajs5o4MsjameGY73T
msahsRr7ULBdrGZIWuZ3YI/HQLvMYoD5SzWXhq9XyT5dpp/GR2DycisZPHRUbbxZ
M2doqAenOF4ISPFGt6ZNAjiY5ujH+wjWcJRdwXM3u5ot5nVqGTSSiTVjhaxgORHv
7B6nbYyBQvk9kxeXwLLdcvpNKQh9/WOX0TUBKNBVdjfe6g9+3s+yRm71bGUXzOA9
ZSo33Q1npUf8PF7hTQWJYlmPu9VbN0ef/gHyPsczs1FlVzJJJBMBHTWSebe4v71F
8Kma3bXxJ8y3hFX6ouvQryfch4V6Tgf0nsnDv1GLHRh8JrgpXPMtxicz/iqDOHo7
ZQ31cg4twVsFbZzGhbepMxwbk53x3kPAmWOq2tkmlYkVXXZaMVZBnzs9UP4ucUnQ
YWGi6C0wwruxObdQ95XONgEVCI5Ppnloomk/Ni51cW/n0EyZT+Wei4Ai1N5F7Vgr
EnBDjPO9l+dlaFl5/KxPq59aHGgqFzGbkiaRzDSK1We7q/QKm4oHv3iL7RHAu63g
STifHTczXmL4T7Z4NiRonlIwxqQ9IxEi56eZ08aIAdzuLnjLS6jsLgrsWlPIe93Y
ZyXdjiPZQ/+ssUW4o5Ba+i6eX88+Ed63xe9c8/cWNJs8UJOvJzNHFCQtTVCwcd9V
EvEu5CBO9Ye7X91k0c7VRqvOhYBCMXG6o67WdI80JqAph3rX5ncSFV0rYSF3tmky
dvJ/63QZkx0N8IuYUo4SJMLlGW0tB8AANAL3w///yPB4Bw08KXslHYMhwwe84yUi
cW6tOXozNEWQwEsEdXE2Eos1odwMUXYXbRLtz45uMEHdaOMxM5H0YPahq6GNye9j
yBANSYz9BYeV26LSQ+dovDl5ZKkeTr53tKU7G+K97gJf4iLDxjHmEHUemOS5hX0j
Xawii6ilgS5GSfVXl7lqxTtBRqcvwHj/29fTY/FBf+1vwbtVNLVXNoE3lx5+cHzd
JHyu41BdGv5gCzfI2bG8Qbeyn38fBPjJRTnlaDoYp/e0grhkEs+wu54nlUC4cdA2
wxYn26A8VHBN50kEGl90fNTwQFYZTErQOW99pzwGHnSb6FobBptde0wiBNUhzoi1
ZURhLIjdbSxFwGNmvkF4/kLuReDfpFcYO7vJ8wmPI0hCAYmOgyfYrO6u9pts0c4Z
+kYZwGZc8MxZ9EcQnRov/m9Y9YfCFLa7z+C3APCvTUc1D6UoIiOwIwFgqVn2V5/k
zEEGtJ+T6YrevxYsbknHiZvk9hPTqFEA1rvCrdMFHVrPazarg6AMyCxCRMfZKsEt
W3Lo4HgIPaTc7LhhHaaarUi7mE8wjKkTzq4iE+ATb1n3FalklD2nycnruETwvAAM
hHWnqtVpf15PKTLmJDZ5EyA8XD35oQHm+wxLhteSCSBs1DGditT1u1cOatlJ1r8t
Ozmtv40dcrhXzp+add63zEWQqsw+GRRIhS3EouARb4rR1+VM4pSSEPF+O97tNVDr
fmIeufOSlsIAxpjdUEbT+MKXKeEvCSUGRk8UhsTEBdnHsXkalNkeLvrpPahukbN/
8MO/ws5C6tlcYH/RHISZOZ+FK3mxoecYSbwXTsHdtwjGaJG2YpaGEGXL21fXxNqk
qYHcwlrO4zc4E8q6JZ48u+3aSUbk3ETELbLqQO1D669ZHsX6D1r/bp3cMEkvs+O8
VOFg5qiDxOeqyg8cacnIPuY7CkPbvgcGm6PaP9GD/35y7eAlYd6ThdcwAIfZ+/1C
BA1ffJwHuW5t4UtuBpLdDsvg0Iew9dDgUVhS8dHeAgY9BMA5hyXngD3mNjH4ZPSF
1Mlq+XcgihWUa9Fc+9QyKDG36/Y5YUcp6uYaRwFEHllUOqPN95JADlZlkh5B1qMG
NGGSUXyhCP7W3r3P3e+QN6yrZxNViMjl4wWOYQpKDv5075l2bUZCCBx6dOlsI/9u
vH9aslStzzQ6Qdv9NH86Z61ExFdcigul5hpwzCcALAKw0OFdlQy6/a9xqkdqZIJT
TCdLh8PmpFKpc2Y6qvsfRnnjSYzzy0QgTAlGThFBX5Vhy+IQ2t84moGSLxZasUfR
ehOPNrJ6WykR7TNkQcc3R73rLDA6R6vLvYYc6Hj6NCCqouQk8nHKfTSNF9yDlsu5
RjKG75n8ejU1SYR7qsKUop7x9FbG2iEc7yLl2Aj7I3rTJ6nyheC7iTagLrj3mTN/
Ybgf1bqE/h1NbLvIGuw/lCgb7dPJiYbD4lkPXKoNNXag0v2axMYM1CZqfGJ8HXv0
giuOAscGFg4tg4VVO/FmdJpLwbHoAyWKMyku+gvof1wmdb5l8Fyq2itCIAxD9dWo
MhSty3dd/lqTHVguHY197X6AHPugNyjrEFjInbXT3f6OTDQ5qhmQHRjPxyBW9a9J
10+sjrR1/+kZB4iLUIu82m1fq8uCKs8TVu3WgWyiHVKlYyhVOox+XkV2nJwe1ICr
i98EE+xCl2DHvO2afurVRfNJj0VcbGgINZfEqzvkX49dWRuZ+zI3zNFMolQp9trb
vpd3SU1J1n3m7jq/vLKLcTxonZjzxh4s+AgOHShNsxdgZHSCdZM6wTxF1xcqOwZ0
GlvnP4ki4fXoFbE/ALTFlpZlmUAfy/FRndzwv6z2XED/fufTqvbOi0Ek+qxEoVnO
HotzPP0hzU1oMALRJqDCifeBzELJr6sgQCwBB2D27vBaePJKsjqgQ6NCMy0Xd28i
cx9vNkFLDmTzT6PGoQ3nmD1WXnpctc4hK3xXDzsr5WsHVYf1c+w4Iii11n3d9N1l
0f1BCViMu88gX0EoLT5r4fcPGnjU0gudIeV9l2irr/6w/FVs7i1o3f5tHqDU+eqf
ykVAd+Y7WYKTHH8VuVAGZ4JeAgGaHJUz1sSHvepUQ65kFp1JyzvZBiDeK7tsPQnp
ZphBExbJQmrgSIgKc67w9MpLq+xApzCtkSQ53HFqA4FpLJLoPsjwB9QZYv4ebINs
1ylZ5NW2x6XXKiWJS0Gl6BGE8GirigxzfFXtp7jZ9UdRPwxzUZ2qWoJhNovRzj/P
SCTsv+DvJZjjgxqohf0qm17GtyH6V8I3Sp/YuHCDLMJhTdfhUAkxDvzvZcpoXIL/
G144jEUkTpk8vZ+bIKz/xD01WK8LECd3+Cza2ApxkYj7qihRs0i8CtC9dHtMiHlD
CElhhRnxA3urdvb1CYL3bt/cIy7/0EU6emKQO5++f0Pk1GO/zrkK8BHR5AZHnYCL
Lt8u+5dtpTQZhWGOzIOoYHXpZg7vkBcXy8RLvsYBZ5+GZsRO3GQ7W3SwORagg0yl
YO+6bZ3c0wWQOZrQSKBpJM0iqVp/j8I5flfjfT0RHwpwM8mcfHVXnHh0Lvo7WxmC
LhCrJr2XFiZMqMHj99ZHDFIPooDPo2Reyct7/BgwOGWoZnH/MubtqJx3RNSQYi8H
3szO/S3e7edrlEFCvoWMduXdDlTegQn5w7iZxZioNzL1W2DBZ9gES75caGPRDSRW
CTOcS7UdVj9JQ0dzle6gl9ko6iRcsbuRv80ywzhwDbNDo5qlFjeAHud/dCi+KgDy
sJWaB0KyNrCqJ9EDJQ0gtJec2mlWZe3vCt+2IYjZzWrwfcmzMPDI6UXtwiwZhnfZ
Nf1sl36l6H4H7/At/ocQCmu21CBl8r6sRhPpNP0TesgEFyyth3Nwcpq69GETaWXv
7BlZc/lbEoT6SpDpWj3Gg5OUT82/z8FD2zQQSkjT4PmtdyjyfkiYsQedlhBYTbK0
znzkgigcvU085ybdCRbpBFiL5CLnM9J+6xfz7jf98F8QN0kVP/zNoO6mto0AuywP
rwClLo4gUtFYmIq7PXUkJgbToHW4XQqVwt6je/UmF64SpZAKaGLhBw5Pm+5j5uck
rhy1XI7lLQ2mEpPSCec1RZrcWUWv3Rp4c5qo5aAuiVo1WNIPOdZX7N1yPAPSzbPp
n03VExEPA6uGtAbUgmjTNPAM9p1taU1MkdM+0v804uUBOEwe9O57cYGzg8IKnfCx
KyBxo+kqPXcEtYgSE6MEyBwjtGTbDVjvvL26y1qthSecuMN5xHuovh7T0ThvWINi
Yy+Ap1ocdZ6+YNxrmZLQxTgKl1msaB6UVeOve99ilAX6sJq9BanUSagxJeMqeXDA
qsUOLVhEz5CjjZ10cy1f4Bd1Ywe8sfGCr5hK9NCnSJtIaf+krClhaC9oh/z7iVTH
u/Hc6CURLznPLPj6hn5EWqDmoJoQ4pYzvaO9F1mNbXXYraIkgWdJxRwlJIElbW9x
GyF5WJ80JZ0JHgdHiqFmQHavR/hHp4F8pLL5HrKYaLug0dmONRmgtYysw57LjQUL
WltJlfQpBQ90mHM8wSfd3+sLgNthFImVpZUpBYW3FaAfI3ifYw4pOxVpLgADebT0
s6rOIUTuvnx4S4BdB3QSnZ5UtE8QDAakxkkHT9b9cjX34XDjqlNNVF6XvRGSWHQr
GoSsJOJZWniA+5sBFmiDjShRV4Ihu6cop6CO4fWO5DN5snLWErN48lZlfZIaeDW1
cBfCSjNx7gvqp38LJWZWNX4cqWO7uD9EkW48TVCYXqh3wi4A3lwhUtu0Pqus7lfh
PzEmDeANO86XJbqfSXSNN/p+EEttmHjau5dwp2GKrbRRucqyORXry02vuwduBGFw
sL+Afwrk7W74IwVsnlSZE3n7eZzdlL4PV0hbXL62NlVx0jaTtzwf9xMeZQNOIL5F
Gtj3qoTd2QBQV/MK3WpIPbVFK7gFwQoAHWGh3qHenXi47hfyxGp77SWcFIHtsKCu
vptwTEKnaO2FiW0b6SclHDUDGmgIEGNPeKqKiJQkc1bHxb11ebn7CJBtCFJPMEsm
qRUGdbc4dgXr0p76wORtBnZMC9JGKkbFnTdh1vDoKF75Dp8DPr8zipP/3GKay7R9
AyT9rZFOc0B7r4e9ooIGi531LAVUAaLQBUPVmccAOnn2e6cvS5r+wDd3SVkWaQO1
E9SQHqAxPMnw+VhMONMVJhLwCP9K39skPoxeKtsYoJkLplgThb/k2vt/YOWUUTeT
FzDyF38/rdiZQRbKjS38IkAQFd2h/69KZkn4DSTEJbBLCIcZL5aMxchoObeYk4Qw
pi4i9xxLjMc4NMPJ67Rp882ModuSvR0MUE/fCPY92Y/MHtsEkE+aF4PVc4+ypDaU
xVIjPB4/zTm8UrJzmzX2AA==
`protect END_PROTECTED
