`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5VVZAmyv0brdK8lYZdyP6ecjPa4vNejAAkVfClDKp/Iuwquvugl4z3NKu6ycK1xP
ej5FFD5MVuqf4hIUzlitu+bE2OkE70nTTj81peA/2MVVUD2JTgwTUbYXIFFoKEds
havwuC43yneBAossukOeZjRarksjCkQ/gzSVChlrT10VY0E+eu/PHFqIkb0zj8oC
yIRWwwS+uF+2XaNjCJgVsOXzKYt0dS8avuLovfRDfU8q0WYkx2FsWqp49jnNSkDA
y1On7vQTmwSfYK/aLV2O+j7EVd98iwz7sPhgi2PFZNd1xZjIthifRwQSUyGEyfQ7
jAPJBDnMSR5vWuaRXhZWZ/+oFQ4i2OigDx5XdVhCQBxW9uPyrxKFACJBiHGubtBq
dbmh+hOD6R5GptB7dStADsF4gnGaclQNyz/J9E3XmdcHc31gdfeDAGJW1l/BfRRC
Fe7J/Af4tSS4hYKya2BGsBmNRrGSzCpaMRMqqHuxTz4=
`protect END_PROTECTED
