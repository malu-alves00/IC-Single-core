`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7nGKeBDx12hXJfq85AEDdnht4bAqLQ8bZmDpAb9f19mkGVOrFbLRuoM0fQ1q4YTz
n3vB9xJuQqApQK7BF93u3ZQleZtLSLIg2vYncYIOhJw0OO5SgaZs9cHoMcU8kpAX
skDZYs7cK70hwWvM03SS83iSugd2+DIL5Bo6WlAlLRUOrJDQw+Thj+ZG9o5cm6Md
ZMHoi9QvCzF/lMNAKKQbv1Zw8iJqTKzD0kIzPdzHqZ4e+WNEs56y7AvWxwjayOaP
rWkGD2h77Eh9jnBGFexG53uoLNbYHs83iMIwmO2Jc/r7reyS1QCwyvafCjNiQ3IA
Ucbvfm4pmiQx6/D875awl/1Tl3i2xkcBSuN43UCPgNfLcfBAGgdpS05WcHRzNXxt
`protect END_PROTECTED
