`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DC9JKHZ2BMpeqyO/paaMoywG01s6QPmtPngKOZOFuCg2++MfqeGcqGczagl1iHHO
Iwv2NJGFTP/4if+hUTplhkpRX0LZ0nMVBGZmdDRwT/GFQCfdK+neRW5SjhupE6os
uCsqsznTtaVXTGrPLf5BF9rrZhsXX8cOyXpj9mNpst/O/jQjx6omFD+x81okFUQz
NSizx27oCTjJ2WgnkSHN0jtCKo4eWgzPrajOX+e8fvMMRcyaPOtMZk09bm7Y6XZf
DBZ1BGJNycG9b5gD4FWuj6U5C2QYxzAm7whDC8mBD2cC1YLWx3efePjRJKobOcCk
moeWWTtr0esI6xPLxB73NK1wJGT0ekX95df1mwKst4MCnPymQwKlJN8D/0ig9TeV
oSjxEwHYkRgA9uBd8i+7zD9pMKikyEtr1cB+ypVMYXv5Rj9Eqy7ihrdce0t3QCaG
B15z5FT/dy3mFtgZB5r4VvgL+VvXwfTnB7wbezYecDx9DsRmUFzG2iNC5+9cbHFu
xul27eD39ofh1vp95g27pQLkQWBHbHK/ggh2y7+3qzMBs/uuLkY0gcTXxdsivni7
tU3IKKbbqv418VmftP3Izb74Pphgdw09Lv8Ma94hb//zkNi1a3f5XUlWWXO+FAPR
cYX7YTXZeJLRUEDB2befMQtMX5yGEDSD9UlbNGt+66kVGpFZIr1M7z4kjxYFb7GT
xXuPC3/0Kk4KSOKml8wT4NwIG4U4HfLer5gjxuN38j9U7E+uTiYOij2oj6RgL0I/
lj3fTcOzJylrvnHe4Mf0vUYUwyFk1BBwVA6bDqiD9502a19GiF7fmeBHfjalCeqB
KKmZKoTSf4IM+lnkiMfYmaqULxl0TYtxidte6CcxSwXuAHmD16erFJ++BXdG4d9J
7E1IjRiQzYEbYpgtLTmsfrPfo4IVv1tAh6L6YSd/KzZeXPUV9UvCoVCiF1Ck61qO
UdOUhs2ypciT0RUWH+hM0I3FWBLlv9XerCBH2wNKb7Stau9nO6KpiWIbtI9z6gU8
eISqtSPsR5oAIeGhFiKqeoMd6Gdc00KA8cHCNJslkBaG63C0cSMNqdKIGrx4euH6
R/4A0t5es7R8Tw+zMHVByj4voua1Ejvl06lieQvnOvWssEx8VqqspEeA+Zc0GwgU
ymxmnoHbVzgtYR5xaiX+dAjXbTb+01Vd+mlkk3Und/OsuI19kO9JkQHzxi52XD3l
6YhytvkKouKqp87u5ekhmoQUN1p+OZ1GXFbyU/Nn2RHSVh8sap/WZZeay757Bhv7
leT746WwHYSxJu6hfUPM+kRzhjzbg8MU7pjZaXFe2OkyVulgWV7X0Ju3DSFSmxjx
VIrBAxMy8jfkRH+8qyUzFnVfWYTdqKeGsFG5Yp8aX2GlK5mPA75Wn3DXQVtscmjo
tRntAqRiWWd0ak4zYlzUXn3IaW50c1JtmfGXQfzSFKt10hdNYs7VaFHidmpa0E22
cH+/oqJ+dn+oK3LDIBq+6tZfLBCp8vhFEA9rBskffkh41wUQtbuHaAihPaTAtRJ1
`protect END_PROTECTED
