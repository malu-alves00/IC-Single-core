`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ASe6KZ3JBw+RVgOeQdGLk/TG/QHq8AvF+oEXSHTwWGOqnWJxKmOHzDXlLVqa1D7A
mV795NdD+9Q+UTabQMVDl5+MGYaPpZoXUSNwKvb9uN2MZaL59U1ijf7hk4C8jU+9
nfurbavDuyQmLMperuwV/hvZetrd8ft6sAcNV9phcVTXLaTBWTlqgglvfo3rRVZ+
Ycufj5wrcUwDHRRdWtFMbT2APpcizwdYccHzbWTWQD261jgZFOLIf8jJyEYi3pN7
4D9uHfibAuQtPmiaqas5+FZ5JgjcTr8aVb7KFVd/OOHX4S92+7fymAM9CKF+5a1h
m7eF6JOmgHnaTh3EgJCXfhU1QD/37arRHU6qokNNowhulHTXPhPqcy6iOppLJ0oU
+7uOFPJrSNhAuVKFNMYQZcdrknPWDjoFZnUuE9ZB036alAkJXVcei7qb09luV7cj
MviKj2cfGzea0eWNKcuVRoKEu7Z08laTt+xTc1FvxK9/MZV8AQ1oDzcJ5pkUjxsP
srVsA864+B5zCVlnY5LPhqcihUqWrXySTfZFkgjzHjovYZ77c/U0pC8RMwbTUQu8
itfMLghbBlOlo5ETyt9mFArWDHWe39jGo/bRWJjnEojH/T9lTnzjjlAnkAgZbmow
fLrUZ+GSpuL+xALbPrXVlFvPTXH/majYYOTU76t16Oqibb9oRnpId6dUTMWY/Q/y
FBeP9nWnGXg5lqNgA9Qk4f7g3yyNUgXnfhM0mnZzhJJyymnu/KMZsGR42Gktn37W
ITHrFeimzxX37TD7jvKX5d74t2Hm611O9ngezTgTGi5Jcl25+8p3/tW8zBorsDwF
1nXT+Yf+BbD9pjfOiJS8uRnwCU4qvf4bymnGdDy04hDoUrJ4bNlSeMWmV7Day8/X
ebSrInPKstClMBQViMcA3R4i1nnqxAj58im2BanOJ+9jzF947Y56bd01hqxFQdkL
L9cPn0AtVwe6odvnTUy//79e1dYL+kHQ6+Ayo2wxAy7aUiX5rHtGjwndI55jzsZW
RLQlGMpUXiqI+wnUAzbDNd2x/3fKlorwjsuFTitSNRMUu8swGY2aEjHjVx0hGSa0
HjowSsrYx6BTKlYUIYw3QxZe9RUpx+tAn9VkZvUUr4xlAo+MuNSdeByXVUM6VFEZ
j5SIv/MjyIMc18wnsPhq4Nsx4uYjqJlI6yx0ZxT81SFOm2cZoyremuscVTyaac0u
JGiaq4YKt4YXa0jm1NbXjpITFGcqXY8BFvDnFfkQ2t2z6OK9K8s6nnqO5UC9oM3a
`protect END_PROTECTED
