`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
G4GIGvhDeeBRoxjp3vrthskpEAdt7zhbQ+D4ReThzOHQnSWABajR8M5Eqp2blA0M
RnjvRc1CA5c7dsTWtpfpZxpoJhoUbIun/mBOlx6FT7aHF/C+q22kouws8kdKj7hh
0fCP9FLOcvXpFYck+/DztNxlQY+qOKquIMeHeHMazzE9bohc6HgxOYnNoEAUMmga
ogjFH86o0JqVaVQ0+XQobezE5jAsDW4Fov74sEiq5mRQcYrNXdOIcrOyyWLnWia8
A+GPd/Nz78WzchEzqn2iQAJHbyUFlwiV/duRH3twH9OcBkGPX780Wb35UG+XoEbV
a76PeEYDjd2OXWi9D7CT6Qe64bh4tXyRP+uCsXg9YJAVFSTSrqZM/fxxitwrGE7H
m9DRcbgq9JiQqb4VdSL8pKWIE/OYC/vJW0+wH70CkU+DsaaWOG6uWAXdoDAcThqT
hXLNPNOSrvtguq4Re73BvXoSCsVQv1hhy4RJ0UH/h/WrGkIBVdb4DI3WA59Ll9m8
KMEjmpVeYE0A5ERB8CdvRldZQOq6rFcQRImWH9N84nUIROPM5m61+dcpw+yFVtnC
JPL9/Zf5owI5871cnWHjROn31Nf5lX74Pd6DNt2GzpnQvjIpCa8LN+l905WySUD5
mcXK2WByWAbLzmXRf5vm2n3iTsrOGU1dBBA4ixQ/vO0BVJ5N785sfFOEygHQPxd5
zWUfmNctxFn6xdEi5S8GYKSefGPIVq+JfYtaWi7IhDph/4Tc25mlNRD8QPRE8WRB
8cLzQW/TcRFMOImu4Q31oEUMpiuu14aqJ6ciGrWR1wZuWVpVVBfUiGRmhOH7gGeC
YkfBxVr3CucajIfiafcY13tvXafpRLt/PLIi7mvY0hpJQoWc/6EzRV01+FuYYHni
IvyKc8FXfHsVAZGRe0UgypGI2UC1TkCxWu0YgpKpP04JvMr2wXFNTo4mNAWy1f3b
mSKg4LojHp2B0rffk4r3gZ0Ha8I8lTEZ8EenJqotItqO7Ye5qFUyQIqtBjCL18dX
MGC2LO4/3rOgnTTR56QASpNK5BK0h3ZM9EACX+EyRtVijwG/Ens00knzO5+RYodl
Bhf8L4cxlK7d8mYe/hOBymUlIRd4GZv7R9EvDX5KgskooQLTaAAwTgOknnHBu8px
Ijo8Xur+eyqObbtuz1XOfumxyt/J+xTFYE3SRL6JOiJUV6hTkDP53OcB0c4rVqYt
lXZicORwkmKcqbxqLyZKsoIs4THMnLYA5GqlaR6gYHWKWbqZylT90in5W+pGcfyN
ts08TOgsdJaWebp2DIKiP2DQdnpgdaGKOmDCCZFTyNaazI2gMWnzrVVJFJXQIS7q
QVUl2j0TzpN73lhLklaBpiRNqJvjeR7GnXCET+/WCLJ1dMv+dYeoCynBwhcADMcC
EwiHGHll2JLxkpXN3LF4GaEbB5WBBUV5K1a/xpDsOU9sCkDAqQYQP3vXj5kM8D1Y
Dx7AXwW7KsG/zFLxpo1FlukoQCg/NLimqdGwgcSf5Le0O+42QiUtmX9qq2tBB8Ga
XmMyvnSqpaJSmu9NJ+g3s1dpkgVzGq8/2a/vw0TxbnE5+xYwe8i+jFJIddUxiYma
NFpiqax2klRPBBucThURUSWJoFJDo7a9NO//8JY4uC2G/Nycvae5mXf2K7uET98g
GiJWdWEhtRub5WC2bQQwu+Dif1/A7jZt0HZC7gHzmek+r8Uw5vbMk+awxZjPq3xs
MUoyjyO4AGCxWgqttsXVsRwvxrnAshZ4rIEVQNE/V8QMrNHtPu57gsACSyfwvka1
t+gfxNp72dePf+dcdGahYOwt8f3zDIpO336gDhHQeZPp9MKUyPeX7ht76755XMvk
Qon1PeJT4uUGvKiCpk2OxuCrcacjgVYUIXcG0G/sOUFrv0hMLjYJuailfqA4tI6C
UVED39hu/qi6QH9srmzrNbGjzU2OC6YPJptvR037Ken1EWqjsExG108oPD8DPb/l
c45bpjJoA52I76gdjdyHQpZco2Jb9NQn9GF1M7nmQt2fpa3jhDlM3SUQK3Bq6lD4
GZYQH+oyeJO1Bbq8L9NWSlqKv0vgoJlSgVOQIoMoVz9695Xhiguim8joOOthRPBj
hon2rJlFqBuzBVBQUv2zWvPTD4RR2tXBXRLasK2S6HTzrpK6l0demKDKNT0KJRUS
yPubDe70yfq77x+aSUNsToMX+LnCdTRNo0C8ucHnTlP4he4KGREly3V9HiOt5PgQ
KaBgncqKlu+bljH0UtxhWL/VRAYMREgLMhHgMSolB11I58H+xhvIfjMxQO78A6rz
IF0hPt4MnvTqqlzorCqtV5Bm7LNKo9zWxgyEDF6CmkjmPHPCQG16fUpLRPmxBJ1V
wGwxTPxid1DrAMqvelUsedr8ij/Uahhmjl7uzQVywslEq2/OphKyYppcPq8yJOdB
N5c+cxaY33JE7+F/R2Ml80AWB9mbZXFckmql2HE5tpkhbXgnLWRZaD/CTcQonmWf
W9gEl2MZ1mocqD8Sjks/Gc32So0DmXseIK/+DmHA6Lducvl5PthXaPzkeQJ6CHtg
LvFxo0VrAeV2Bii9IYu/Zt3nNlOH4uYwYRhEeOI1lEjkNQzwPY4pJOP+pIeoUkDE
gv9/YzAVNNaIf/ufEeOZStYNQqllYqe3SufOE28v0fz08ZiFY/PpS58WKXKqG9vW
cc6vp+KaXHhAD9SwjI8DHWW6ez9T/GeYlwQjWG4BTDDjuJAO4nz6k4e9ifvSUFP/
2TaUDM6/bwThZVcV7dsOip7UqPQYLYOXMpmg9QjDEwp4UejlUfGsq7HqtH6AoPLf
0zi/mcCQ3TgOlOh3ry4VlNmgejIlgd1X1zvhlxtyUNMY14ouYRhLsSW6ZUo8wu3S
DoZtude/f1uQlnxy1glfu344yCDJBw20Vx0ahHaEDkqk0tC0xp9bOcddeM02TaQK
nw3UtVrCLe+x4LpyNFYz320kKviEGmPy30xTPbymot7JZIe1+1sEVk6PUduXyfOm
K9ft4g/fURB11oLnJB5u/bkmzEhypR1PCZ7CuY9ibdgmmNzjQB02pEKflUPBuR/T
PTGsrOiVLqd1cQuoEkg5Flar1wsckvqZQUmOwrjFq9+y9rFAU5UNmtT7e4jwoVlU
AqfBL2X9JNn77hZf9ttMnv00XVmla+7D/4ldGBpr1m7hgOC+kab5NXfAW88o9Wrm
EqtzGBKSFJpZVQ2ZREOwRaD0GYfiM0KuNIX7ysF5S5rFgmoPJFI4m9KuY4lLElFh
zQzqzSPaDBGO0KEbIHLYf5gNNc+q/tpuPkrE8U7uBwpx/pKnRORNYRoYDwUDh6Fi
q4waTVvUUfTipp3Iws03JXjHz+4iNDChez+UQBP0VPA4pJsDd/iXaaucM9gOTfcb
c9E9XMlaq5nEBVVRXPANiduLs2TTOLouEUUc8TlVk0/XCEJjnTs/QjAHWp74HxJW
/La2qF1OOZzQkt2eYYATHFQBDvrmaeK4BpAQzh9C/CvnCDHgIV9tcJjIuwsAQ/vd
Z00pGqcL8U/sTUmgfwp1iQ2bUBqMoL7Pz/jX2v7O5/j8aweMbNXnJjHLxbQ9WQS2
TUqEmDtVvIX9qnIdUaUryyDR05BVHwHTo4u1mzKvfQbzi0FYeMM2CAwHuoSZVK4Z
GuLgM4hX3jS+yU8asSpYwOWfpRPcyFwjVSX+qA2EcjOws6w+dFrEMdMYJHNzLcs3
DVH5zKrt+21IgREd1mhBkn3GKTJZu3j90W1qQyjQQ0FAb/LYOLuc6BY8K3An4lCw
9hhwyPeSMd4GevdmpKgjdjCRAikzDBXB20qjai3krgSxEvxdqE43yShs4MCdXo3J
DaTbTSkme59rSeUceFvDi6oOprGW7Q6udq7VjKyq2ZalbRAUQJQOSnu9xf6+dn0v
Mcf/FJGqR7Cq3ZrbI+k5yXKvtGH+iyRpfVuZTq4PoobE33qd0RaPIVoTZN/ix1Dc
h7D9wzT8vTH2SnTTZr9dr/o8C+Z/mregXC5VhmTzc3zjA4nXU27H7p/sJRnpHjaT
Ny5kBuBqzWXECchHtDGkIYOPnstnuGCxQlCnLqwXwQJzO0693eWF4K9pq/hH0CKZ
5QGQixTd6cdYWN7zql2qVwbmn2pdcf5kbELErFBArWdxlEXbsP5+s7fG4KuSvNXe
BEzTR74IW/8eToEVWLc6rnQI62fwpI8iY5iflJ3wFDrm8Uufwb5qL7n/iKfIPeMT
xkCCWykw5L7EHsylfSt8RZs/pGazcHKvgTOd4Z757QL2gKm45yoyArpsyecArI3P
PV2fUA2Dwzqo9j8flHh5YCRH9OMbF6Pc59ZgAoiYov1HhCekCfTE/n83+14iXNVf
GvcdLfAmnLTwY65njioRa4kPE5V35x44iz/O+UUuq9IGJ04LnQej30Va7wq35n2h
zGLQaw3mX7Zue9AtpW9SGzUiqNNEddaLZVaBdTUzOySoHopIHpbZzqs5Ja8LoqPC
`protect END_PROTECTED
