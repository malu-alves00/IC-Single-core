`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Rd5GxukYbi4tltUzTeICnwn6U+ILKZISBq+bUD9eLoLseUI0QxiCwuw+wpSu35q5
q6H03hFi6TkyBWcww/euW5KrMZQlNLN1ODBSrq6yEHAlcXKwRaBrvg1Txy48OnU4
jA7p4rNLMw/c6yVekvCCrrb8qNbLZU+KfpMMGq7e2YR6aQQtGtv4z4awBdsOUT3s
URpqCRi5AT1kw6xgBBXd1X1K20D6G9rkbcO+dGlBzWqewPlUOBlDCSkMCM1r10jn
0RxHO6iXSEM8ziJABX20bu5985oSazaX5NSC1rBqAoVMPAcD2eZ5kemkfbJqB88H
GfPI/U08SMcVgRIO/Uwbu3Vcpo3eRpbMQ6R2MxreoBFOIj5Ax0n6CclqETV2iD3T
cPjSVmBHsY8sgEn/g/dFtjUww6QnDNKGFA9arY3/1CViDXXu7TAoxph/gUz+Y+Hj
WFTduXNCVF6MIISc19VgBnZkf2Sr6DsRBjv9ljlV0lh1Kx6jq43+jCVI6Y3CKVCx
9iNjxD5+Ya92RYT5LCRzFIo2MwsJASyZs4umCv3bBFSx3RDJSiPmHtFPIyPr9aAR
EWoCBN/QpWjArXvc4e7jDYFXWaJo8ykhXPM5jtdv28mSuQ9iPgzs1psbcN6zum05
jeZStIzV/T9qOnCXgUFp3kplw5fOMMu8Osig5TPGu4mtW4fS5dxG8j+h9E9ex5s/
qu9QDOOkWfjT3CrAERo2BDH7/hXQ1v/yG4+fUfgRamIUDDCBJqwjBxrHoApQ84wP
2a2aKgcxJhnvdKSgg4OLpvMsbqGDdW1PO4RfNV05IXCSV6ie6sFar3jtDEpixJvc
0bczKEGF1XqojgYkPvGE2QXHVSqZFRP1FTwg6ogapDnjhDMCpWBsFjGG/1ykDHEE
EIHoPdSzDjgfLcadflKWjPepdZQb+Ww78MucnahJNFLu+5j2yYP+ahjnflZYNNlA
/RmEz7lZwUB7nUvJ1x4g+Foli/nukav7/XG3r7gmpuq9Pu51KJ5sRJAQ9366UxSU
gnQ269R5oi8HbnevG72HqTeRnOxpgZ9YcfNIyzdzIWKGny6nDq/XDfsxZzEO87En
SwGCGeQwMSrH7JS31ismiW2FXtOo1kydOBSGNMgcO0ydbHju56TRxQu8ZB7wrDpJ
6sMXjjNFctgTVqeSQPn+httqiy94oC58OKTfCoRSMJciGn9Sxr29yFruzXgLDwX2
pGZB8LcVmmwvOtWLipCmXV+wzrR39GrQJ5zX9h0wk0Dh92GPHX9rsPzvam55wjv8
nPcn5bDWvrFOY9fGsmsI1DT+UeGopoQSfXSRK2snq6DQlaxUGHP2pOOvEbdakKSy
ttWM6pkEzwPNGH/AfnxHMR8yeYpgGLTaPHTva162Og/npiTLd60GzkBOsI0Hn2ny
C3XQOVmbDko4T8hj/i/alB8iHh88eNHxPw12wkvpQYmCXQzRLHb3uTVRcRNjgVpk
gpa08YuPh/UA7zYSzBQ5QzDNhvosSVRAcx/ADZPuzXc5hnjze3XTtx1PHTSM2eye
WiRKUIXpOTRmuzbDW5dUBXeyGE8RHC/DCr/3gzcEbHCkQAlVbP6ysUdIYYRj0HAh
ZI2PYmBgHFaK0EIrowNNiYSMvW4uwNaA2nj2KVrgLtqQ037zjMRlai858X9HpVok
Qo08ba7Jb3BoZfo7Q66LifyDWpuMf++5FECnyNudILyPsRoNaBNo5M2NWdYZEvH0
fPuFNd3CsR4eNjWV88zaHFs385V5wNqzfjNxlj/GDOr6rIeOm3hb/AD2WIF92s+4
VSQE0ROCHcJoadUIzUDJNEkFJTlJDYnBLAl/6jC/DMFvSaLVVE+PT6k7CJhTneEP
0EYZLGbDWmjau8H6YLZSj0E0gI7dnR4oL2ja2TD+MDg6QCnHGobBu8uZopKqZCvt
ud4QajV82cT00qYNJQqk89NzXeWYS26bsRpxg/KyHmlafoQFb+TcpCQOdJKK5EY0
BboquboRtanRZUf+tk4dZNHVeuKw4eosq56HlDibqJEzil9hRM4eiSZSCMH0+wHe
yNtHkbeVQVRC9DzC87hJUom3wuGzTM7x9MCB31up90CtxPH5OD3Px7VUAEQ/u7ZA
6SYsR50JszSGRkDZP7zAoI8dWnQlrgL7P66pC3YHv5le8Vr3BzCBiZjjB4qRAmZd
2ehSolzV8eIgYvdoivatsVfK720DwhmEGPrrFiaJS4KmrhC94rPtwdCQaQ9KF313
e8ztANJPigRQXkZMsWRZDzdwZEO49VlvlLo5LqZrBaTpL97vs9N56lD7YPmxDZZu
8wexlmQCp+VAzO0z9q/1siNCSJ+y520Ka9Tya5kq0ZA1ieABtd/deIyQcrLQCpc2
cOoy6xEUcaLccEsOlXuo1QWStqXxx5sZjB7vSL4sl4jsa+BTyUJ4ckn2R6DaiTBy
Cyu7YPJfCs9cDSGqIJtgU2QDw09w0jrRo/g6vxfO3h4Msc4aLSi+m44+IiRmYgQg
FK4sKpx0hzZmcZpTwe7cjdJITLpK0zFsWf8tBosRjeZLZxv7auQhY2qmrrR805bS
09VutstlE5dGgowjFC745Qvn4wsgPvqHbyURIQ3hFcok9jZIBhsJVFWD/YlTw+Tf
PaAL6dEYclhdAmIQ2nGq3wcbU1iqOHLCDPadULeI8hEAVtJibdpz2sDOKZLuod4i
2406uj6YF+Cy8Hn6OgQHWfQx/Vb/0W1ngTBvkrZVtmQQ8uaivmQAap5IoHn2hmth
TYskPXXHBMh81yiOzyGYfsgtIv3//PrYFwf+YlSydZC1NqPizr8NA6b4CSox70OY
M59M7gZx5/KREw2e2cA7T2Z3Cw6AW/Iy4Ju3JP8XMUtKctp+ALcMKIwQsIv3svk/
8eQx86gO7d3MJrk2molixBo2VPPlOn/euLsCvYwftSVkCth5RRw/z+i+C+XXdKAJ
wc99++qWsn3n7ibnrYHPFpa2b65g2l4GQA1or7cm1DLeHA9LTTY9wHQ2MrlHXbTD
lng2t3J7N1t/Z8QQ+ZMFoUiCsh7a7BnkzHUFuN8mb8oYSuV8AgS1cspTMVXeSyRR
Sn5wqQFuhp6VHrCG5xtvYGKOG3ekT6eDHXEHWa1rOC0FOZ9cOBmatdJgVOEPe4hk
/ILyVEV711R+GSERICOH02I5mLQ40pQy6ZCZVb3Nn1EGgt7HDUgO5ECVq60mFxxV
dhYaSBJxGP5gmN3NwZrhpj8+fZLa++s4C1zNPe8rfiphFDSVbe2xuM3zEJKSoCSW
Z0HYZD3x3AjZOZEFrrvmf2WT0DO+bGLZaz9j5fu3yGzXpencHTc8Ja0mZBYkTe0f
8vw72NfEX6eOZzfj8gaMxjsFcbaYqnadyb8VOW9Mkzk35IumEJ9cRa62eSuxTx5k
H5eo1UmvHdffaSs1jZnW8nDDm7D8IeZ2skhmUJSnyuZAUMsnpT4QSXdxXNAmaMDA
PDP2eor+MprCMpyKY+6i4Yoj8FbZ8koZ8maSZuMUIf5v9Fawb1ilmzvHSsm6dIkt
an2ThpStGsgoDPDfqi4K9+wb0c76xlh9dWRq1gTqulm/+U5CR6sYa0m14BX2ZzOy
NPosUwdf9Ey2a9OaBGY8PxUFNYHzWlyzauluQyi5fT2h8CJ4qOK0CeMi0Lp8GP6j
WULiiEeZVOW+AAITUVZCXI1EgwG581Ks/NFo/z7h4nc1sbiUCZxi+p5CJ/29KMwK
qMPt+YNeRwE9jL8jCYsIWA==
`protect END_PROTECTED
