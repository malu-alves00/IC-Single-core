`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Sc5+oGN6a2HxU68smSk6xobjsf0wZx2zuKZ3Vsat52+9f11fgMEyy9+914pVNpQk
BkYYNsI3PWmiSuxCH45VzXrD5FYa24NbvQ9CL/pF/CQjPGA/gfYamB5JLkZjPP37
HYGSiLb4o0dgkL4wejdYe+ChpGmXgNpEpoiXtYHQji4hncZwEPn0Sui39cJaR/Nq
Xj3sPpHDbLgw8EWYjtKc/d25FU9eEBX8OXe5lPzQdJ4v99bNeJiHW38A71egl9ML
GXKrv3nW7kF1JUv90w+aA3NGniiZEkg+gN/i83I4UBD6sMbqoLXFNhBA/x0y+Rk7
tDxni9J5BWIrZBloDVmy5DLlT22Ev6Sh4hLZXxb5C+6+V3fnJKRhUeUlFkZjweN4
8za2NPuYarweiD4f8owd684s2yC5LsaUs3BLhZ3Ji3u1mQ6c794ETAIW7okCZwl1
CqTHlxT0LuVEMnsfpP8UUqAqPBVdRgTwnpW15a4uq/d3rDNbP+7YaH+YtAMEjGK0
dCqIeu5jeDl16LZaGPQia9KswJmfTsAlxBjznuPv5toshHBjQmS53eGOajHzfrED
TI56qeyqolwMp7o7wo0HM4d8fDLl3ZOxf30Gs5l/uyRIo9FKJ37MCBINLlrOuEi7
8M/VS0sik+YEgQpVFRGz4zAmrFt6Dx/X/CkWgVO4pRgtw7SE/J3196M1saWi++NC
8It9o4YSGUsapE1VHnu8zwG7IxGzKjyc5ZZYuO53TD7kVlS2LYiGhJTdO0F8bfDA
NbfuCS1rny/dztgsX9655u21Hk0Lre7gbb/kTDzkO2C3TSy2NTEmwJcZH/WM0CAU
9Cs6E7L6uFnZmwrFdGV60eTEKXeOq30T5CvjKtk8suMzQxFoI3JU5c9ZXSyogHxn
i9qSQ1QB5d4hZTqa46e76YiOSnvc+EdbCYP+5tL4tV8FjWAJrQn0gHo0np2sYZCt
7hoVN7t0gVi676LTZNAPP+AKg9zhCGD6O88E/mhOrVSLzCDCQoCjy9MQ64X0Bm1y
1LP5sbJvsqh3f8xpVN9CAqlki2xqOk3wGnUa/P/PxHKwhkddFhUJoCkgZdfqtcVf
1Luj/vlSMhId1n2t/OPJ6TTqRwg1Rqq55SY3uVDgodMD5vD65zZk4y8dSSF9G6Bq
eqXDGDu9SbAGR9M30rQSBJKU5u1bLMXWZML+/bqed7PdKFzT8tXWvTIwY8ESbFG/
m9xUoApV8ISn/41Dx15lfUaTqtEV8/6hRkH3Wg4Yne+RP/OkYqo5aOG8+w6ay/zp
e/mECemTHUikZPRuYltm9kb/btXeZSqa/qVw4SVF9fXgBm/PxNQ08PsB6LXIw9qa
mRqr2S0tiH4kdleXpNb47GrohBUbjYoXaH65cjJgS9M1Su0iiHVTpUrf8PaFKbef
N609tgC8y39p605GCDOClAKHcQ9WS1Vg75feJ4Di6BV2savLl3gXsULMc72qhE9l
DA8RAHrdasa7nyaJiaGi83Knvv1MGg/WaHF7Hnx8zBtQE/amveIMA6rMbk8+kuqV
SIraVdPENPmxa97OKZQx+GDP2ygKUDHsylaiOpGtgv6TM1rMfXSGfHig6TIVHOMv
o0cZiTQmht3Edy3uL9jPawoszlhej2wNaVHemmff00e0fmm0iLNfO6tozHgrxgi9
tkVzg0naWCuQzXloP0WiF2W5NKF3fodf7+hgRGZdExdcVKVPMwcGs9ztNu1dPlNn
p9m/kUygkmPGjbkxh4Fp3slIABjaA2+eCbGm71uBIYdUCCMyeeXS6C7W3w7gLjRD
LCaDNKaAemOPEzfx18UTGAh4Mmqj4f1T5+W1jKFyDG5xRNY8s/jF7xVZRY67wxDR
z9vuOuhyxapuucNgtpsA3x6yAdRvDG2VlkZZMPxW2E9WLH7dja/BNI/w6CjYgfL8
TWcZfWxXElZIX8+NRzITJEM0/ykIHPOBfeAhEAVqKQ83fflGKLQtCX7rlmAStNjl
iRjA3tDROqljhR375h3DPe/0yAYQIIYJXgpVDGvujPPb6M4KezRh1V4NcGosSTuW
gbymwcAX5kULdKUu+YO3i49L3aPy+ytTSkZya+xfI4BjjShCcR2lXQqPs1r3jnCn
m+ybYMjicsti4YC/1x6ILY+/ykVK3jdw6I+c7ONSNmJ7vl+rDpxNxDxdajCQXc9g
Z+iHik428bioq663hfVqKTDDYkY+0UTErsptap6qyRG8We7prpI5xK8j11m93teu
eSbtrXciCHiiHHMp5g9Xm3Qairz/JjNJAIIyNjgwJSYGuy4yY4ZuHivbCzYyLv3j
mnEosA2voXf3Nu/KIlgZM3nQvwPu9hML6nykGhkrqYnzgYzQ5FShq47gV8qwsY1+
SX3g5NUQAPlHcUyrY6G7vMszWtaH8kIpQXvjscc6I0gPRHw6JrAxLJj+TPc3tRtI
TkuFmPhAkjiUthOMF72EqAwDmhHFrTZsi4HW5XFWxKnSos8ar6DSvRrXbzGWdG0K
fLY1Ou6+HL2rByfagRFhcDKB+5f5b3JdqRvoZbrbNYpfMLINBNpIYPTnDWnyrtA/
zIQVQYw8q5JRb0kuuAS/yGqxV0OVKDqk5YGTxntwo1GVyS25MJ0VDzBnCp268hQL
4t/mGbRnt1eJfspubZCdV4ZXpvrXz1L7IG3KQg5i0nMhTz6arqDEZ28rodFZDZl0
LGDNXZFnDsQ886BRg9/CFxnYltr2/ERjLsT2/0zgm2vT40hGihukoY4yHWYmvRik
9yHYus28itcIkXnAsD2v+uPBBBp448Rb4pPs154961/PMkMK+a7Sja9vzPVLch6q
xD0ErZtbj/aG6ZBsBrmARMvjiUURD1jLg1btA3IlotQH+xJgA2+6C40dy9LSpcBr
k7xcvH4fWMUM0Hp9q7dr3GYecCNWbLtBhvjgqpZU6KLkn6+1IENes0lBZgAa8/EI
1QCJCHw0RHF1Mot5Q0JfHeTDFPXcg9/2i8BL+zJfTCnTQ6gszqd6fDiLMCqKULVR
lWd1fcDNpRNjGCys1W/SS1Fgs0TKq81Jr59XsxuhwHYMz1qp1J8o6Uyh0DV5uV98
uF358tEZnedZMx4lK3NygrYVTejOfpi03CEa8k5RI5/v5fpvmBvMxbmS9o9vnJQE
WUYptc06GEgxB4QxuW3OaqNk6j/AwBbzio8nDzbFbFLXaccoY5D0YZEbw7XVb+Lo
eZUz9v98iBWRQOfzqHip3+ckoc4x4BJj0xhNDAxnD5NRjdfqcMlVHgO4WRJNpPq9
93iuEFNrLHUTB2dzbsRXdV+bjFCPr6dugFKI648en5VU3tqIK6jjF/Nm3LAV30iW
FklyJXQ8sZOokTB1mIFDf8rzab181/GVvhCKzxpX70KZmx+SXgwGwIFhXuu16YtG
EH2vErkUyXqyiyTc0BIkYuLsF+PsQ2RYnhxjflcNaSLOIj3Q4qnJDwK3W1vAzlMQ
HkPh24azewReiO6yjychmt6o1DE79IoNCYnl5trcrrENih9T+RIImuXPI5Zcw2IG
/tCuplPTNcyU3Vu8e3CDctTeYnJaMOllX4Ub/r1klq22XOu1mmvqxShZS1ir/2MF
2iRo6/NkwxVq3fP8TmDlgZ0Ya/XZgg0h8Kg+6P9B5rh2KLgeJ0K3q9/hSunhhBiy
j2SQM95EcUYs1HR10oBzrXeZ7lIYTpIt3CKeSZaRTY9y9ZIQvXXvo6G/QfJwNuEW
R8ipKC3unxgVFfrsXCvT8oFymWx7sB6uIWA6/SHfcBQPSNM6N+61cqhgtNou1i3s
tQAZmlVUwd0Lh/ghqQAgHJ27ksMXuWZSlTxwaGhrTDWJoYaiTiyoM7UO2fvn21tp
PtGl/ygoLwPGbijnZggNtMgBtxxJXslWvRx6WmMWmnvxF8VqbBgonGrcGKrSgNrQ
ot+rh7HBWVuBDC+kTleWXxFPLRAp+LZe4iHebPQx9CN7MQFLMQDPmumIdUCtCDow
y2XkNNrIKnZN+Z3wZ0+lfa3BFYbvJ+cXzkk09wwnAwjyU4upvhwTIG+wKt1IKOF/
qrI0uQup/dT67qTlhP3b9nqBz7S+WR0QPlJN4/xf7CHGiGmXP1JPFZFtmNDIsWj5
TlGeZ2sPUw7sWtsNXi1vJVowSoYVCHr1+n8S2+3YFXUmXKoziMK+PBTc1Lq22Qh2
8OTSiGYpxIkiieHdmR6Xl/fhoJGQYZdh4JinShQVv11IQxctBGFB2YknIeRbR/sr
nPf7dFcLqM0OI1QX4R3HI/HaLF3M2wiz3fjsOWzy4dDDhtxDikT+m8WhYM/Cof+5
CnKxoKAdqzuxyuNrtQSmcmK5Lupkd06ojEHfZ8ZxXuozRherZbJZwc8RoX3DU6zK
VufxQmOXCVsTGxLpKI8kwWr4a9whuLq1YlFtPFI9D30nOfVaiZbCXaELwKFipVjt
wMIAK4Y7ra6VTP7f1MJReYs9Ko8mTEXvfdo/aYikXn9wjSICwbVcf1gnopxKf3Fd
kYWHdDAZKIPNcBPyCMCn54qz1+04Fp7q04GrdJPqU/fKbb13r/kuWzyqNXg00Fl3
QFt4UFNQ8W1aZJXe8asQ+pLBi11sXGES232OXKWzteEAnZrRFEFqz7ZaDYklZ1k8
DYHZmPK5JEszuiuRIl/lQnzeyG53JiD8D6jmP/3oC5yHSz/afbqAQhhdNXYmt08V
+jmssm8jErFcLhJ1oNA+T3zM8/PllhRXMz5oq5mk+BcwBLgB6yRpe9weW+Z/C01U
fcuT95eNK6BYqM8Z4cDn4h6bGlh7fD94Kl4WUBQBQyW443Xk+Olk2VaDMKVt9Q4D
Utc4ibTokzLbBzxr05GSrswFpGdcs6Y4AzPSRdWlDnpuN0Ey6rUtQq7DNCmoxYkW
WLz6KP1FH2W5epliDHGznfC4LbLl5pRO7uhXjbrGr64JUGmlzeTGl0eY1GLrOSRR
JMzg0CaAioYCMQLb4TSKEz+FkqPmR+VJYC0GQM+3G1Sie7T712wpXLDdF4yRgWgN
R1xi67SC7NMD0h9vGGwfKdR47HllwYGAitQen9x2sB7s0kaklQLxXVGX7DJHSv5N
Fn7V5Bo2bCLUCa/mnlAkfXmUc/2sO5UWr/r1TjwvOfk9MpWmJefYTWEgtRQyWPv5
9nWZSHL3NsTRxoxnPA5I9uDwW1CfilcXaXCtq8gm+4gYQ4BCHltbLGqzOsdkbbap
5Dh4XztV2zS2vaXadF5mm+ljp25ktsFX8fNy87LYTl+vdscVk0VcCnAKXyWzcmkc
+76OgboHsqxpEdx1Zhtia2dl91q+H50sI56MtPYHVOgfMqZiLU8NEh9TuZOvOhe6
Z5c7o/bLaUA7jqQHRnjY0ycrXQS/LXdTrbjGJcGaFBq08LpE7zNw0X3G0UNmemco
CBAPcyzWTfDPKfQfbuH5KPNG0ZhuVzbwY807EGuVU47buGnhZwO1ctLT17lEy4hb
c0KAK8m46SaoBaJVQxzGFsJvpOXGBM20aijzeBe4pTWCZ7NYMlgYTzExG3J2vhxd
yEwxNi9dgbutfiCyH5PpEN6gunow7THzayFBhDF7h6/78tzRVe4+vBO1KkeA1e2R
JubeKCWRYcbob7oX6PBPLBbq1qrZMXW9wBJTXlnkX/PwM8Wg2vrCQ1LuSsy92kr5
oy5VHS68zKmnbj2MWKXJpmrPDY2fl7WFBu61YC9D+XGvPhs6nR0SKaXV5Cjcct9O
DITGF7/YeBfEfNSmm+HTyYPJZN3nOF6Qxu4Tsa1Nm2Y0r1AJLqXleVNBrFuXHy1j
ht5LDfbZsmfCZhpWFCcMxEVLBuAZKKOAo0GlcKHGmUsaoIjWNZIPMlSTk2tufriq
WYjCRisd6f6DwT3U7z2VgVton+U6cnl38D6q+5/s7uup/xYIJVIyW7WQHRwPm5xa
kWzOMupdSm9olYuniTxubh5Jnsx3N3QK9jmiGxSb++DQugr5+1PgG0Qjg6hyXbwy
r25y4Hc4Zs8uHeAvZT8rRfrEiRHHks5lhCfebuSezJKJwN1vLRTX2fHGCWS/ipk3
I0X31XD++YMavFiDj+OOI7zhFcvI5QeFRkCozcvpmXNqO/sT0J/vcqAguR/Ur6XH
RgyPv/iaVVhnHGZe99Yeuru+DcMbIviZWI8pf7dRYysxQBvCOi0r/p0VIpqCwXEj
TAjdk25EvxdP0/abkSwpBd5joTU6SrNmrb+mZJfohNQe6gqkOmgIPwWr4YYbSAMw
OH4KmoOdpEroIPWY+lbh5PHGY1jKUPDyorQE2VQUfqGMrSplw5UYPGxqiJMlisf6
HRKhajh7zdbA4tU2pWEX8Kw5N3WZ0Fk4Qg4xKicweubmGdGb+zzk/9C4xHnXyNro
6TTeRV5yLYUg8fhOAzCTL1BqPrZmEC+3NGIGqE14Gd+2hDGk4Bljm2ScdEPvN9SO
LWgUaZPpbaUc6RAQE+SAPR18jaEkewMNnBfk+HlYiwCk9Fd8LFFbDS68H2/3PRYC
bljkO2fLDJuJUA+iu2oh0hxX11c6T1wQXPgLAFItbH2yhxePPLyl9L90Ii0eAFei
VLjFKjXwAAlzzN/Mcr2zltJ/1mLNJluXV+JIuKZD+Yan7533xOdadx2q8y26k2Ed
7nRkzBe1Wj5h8baCvL2whvmqA1Lgyp6w18scD9f5Yy42D3ZKAVLyPddvSKrYjNGL
QiFeVO310Du2yFCpzO9XdkJrmUGUYyNcSTVJzU/2HNTHe854lMjUUTuEtqEhzFo4
bLXEeHz/4ErLQWPCK5PLz5HsEaJIdMfidUfKvd84JrkLqD7oVP53/FIixfmnCIMK
QNsKbD3UBC/+zfBUp8JiL9OceXNRdwYm5miFemb8arrleEAPAZZZ7/brWBdPi3P+
WIeCV66VS2JM4rLkc60mUWqy4QiKnDQqJ+VvXhlotb8OhNoxK0AkVtDsV7u1XcVK
ReTzIK2GZMTsUVS2Wc+yi+nPGfX2+byBD1+VzWFouj62srV1E7CGxNfvgB+ELEel
3p+Av26UcE6vb9vSW8j9Q77OJektVcwHbOVeC752AxmFDAsDm9BV8nQanMI6j7o8
S7HjCSxxEUh8jrR0AEOPVVaVekhHhZWM2BqVwwCCXMTK+COgnvp9NcLgSBeFZ25I
19bXcqnHll7WA4XniqK/M024ZfZLwYYW+qQLHFg3hFvlpzU9P7XB7ImDpg2AbBl9
ZxhvolwwBhpwJceU1tXJyDLD4C6+HN/L3Jid5iG3/vuNkWbY80iPPDIqZnXuF/6F
PJQrFdGlFp0FkjSLMPduJbwA3TCbiykwL1wTCaKHEQM=
`protect END_PROTECTED
