`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mvLfDK7nu9bJWqDNKznoTZVoEmQeXZvKA6Ux+/1ss2EqjaA2EJXEZ+YL7oim7tbP
hFrlwkXKI1wdJlpPjgBRwsY79d8TQuQ62RF46mHmCgj2xZv6yWhumF2NnSqgeqm2
Zl5rQUtRw3TfDunExydds0KRfQ85vEEwMbAVnPAzpdi+dJK1YneVyH1Y7/acWksz
zC9rpLZidjHurneCkIjU5/+kqFFNOFUnT8st2/H5VHZG8noWzx2VWzCYK6rw09oI
h9PN3EyhdO7WnIyowCfkGA4Erl++brQ2pDy1XOAc7y8z9IsLL/8zRYCov9wF9dTu
q/5rZXCX3n27CNWDpJSCl+OsiYAdPI9ay1pp9G7J5mGo2658ZuU3peFmOPX05Fss
PJWTzsL+aewqetGEf/wRcWacvLNoMyJyLao941+PzCJwpRvdFUlV3yKF65qIMGiw
pjbsFuO0t3WJHBVujPk9Rj+Yp/kTH2yWXUVD/GwXBBjnpZUuqj6og2HEhGmFwyEI
jehtwxTKY4ewBISFevB6ATNhhb4+gbTD2GLOIZUD/oL/RnAG+SJzwTFdehd4aTIh
n2s9D56zjDHXHDA3ug5VE6lqgn35QCTRac+I+8bT6CmUFY5xoBplzGK9e5xs6Uw4
EN7DPIe69ctkbFXAYcPwXXIvUv19NKv26CCjcbY31kh4PwBGWYpmDmy3TBfOVcT5
7tAhs6KGAxUCXjx/U1nH8xge68kvvyIH1sKn0ImFHXh5nIyKed5Mff46b6o6R1Gb
1JLCBb7aUyvZqtETplFkDSvoj5Khcu/iuX/7INwMh0Me3QtgWjPCyhzy98YgUId+
EB7Nru14+EHIlVwD2CsJBVX81ZrNEVKk6RuxSDJL0GykFfJMCJmFaniHOGQwfdOx
XJ+dQDnJChuiZKlVGEpGWTj7ewYmgbI7SjOnXdTpjD72rD6bkyKg/FThSzfAYGTl
9BxG1eBKBQFSzForUeAN7i2rWaJGWe0vTD1AKDSKBBFM9USXzaX8s0PEU+QeHk0b
H8jh8xKCJdByG5d2Xx9iCulCAPLPnN3YcOz9sGRJcSTayCy9+bhh/67Yen58nI+b
IL/rmnZbejD/UC1Rlfi2jQ00U9aDOelbiF7EQs+nrPKPR082+P1+SDb4Of+t+CsM
j4JEorg335XbZxcCDdZY9bV2IxmwiBQDtFXLBZS6VJU9tiRdCP08MRYzG6arjZYD
6JeHYm0Whg+Z/rIQM8w4D/h+qpqGBKtnN8vKGGSJNJOSV/tJywDBndPupErNODIN
HUAYk9+BE2xUYR5NcHnvfz8ed6DuPbZ5EuKmr9p+nNTbz4zsCkSdzPeE9UIjuw86
tWPvZRUPgBRp8gLIx2hGSjdWCqRWMnVQ/G2lCj5fVQKvUC2RDG1Hd7aiLOucP4fP
U8a56unrUsA05gX38TUBq/gbViwFxrfd4YZlyFSucaAQbR09tu035gnhIPgziVjL
TtOANYqNKjiRbtjBvD/58ams9+SVd6hdE0Kaali6B+Mac1b/MJkIyfsKdkJWGQZL
rzWUJyAujLNaQvtfud/InFRJ8wed+u6kUKB2U5sPcW83Mbtq5jqxJQMkuG7HuGz8
6Cxl1ZQ5cSosO+wbLurF41oZklHCIzAFrf4eW9d1neIfxGLfZshvzcXMDXIm9FhB
uKMdkFpdauuU2pXtbpcq3xmAjP6SF/q03UECfJeDv0RYy5d3BQsspcfzWE40g6Mf
7/FCj0YhK9Dg8PpDwRzw5Ep1atrv57NzLrVyR5vT6l6qTwgSNmm5UF3zmn69bxo7
+3h2vDkLVH3VFqMomSW9pbJvnZ0myJ33B1U6cvc9iKDA76qIA68ciNNLZBfOxnOo
spEg0L8YBCn+7SMFLg1XH2Gp1EV9kiXNb1QVjsslGhHNpWPDI3mf62NE+kQDh8Ah
iJa4tMVW6UuWqtak6GAcIGnW42ZD16jjb9mh0rteDZFsSmQeh+TXNGNWcDbw6qFX
fZhHSj0XIcb0YscSl2nQMjV2kRDaTS+CHG1KCPTG+DyFe0W/yQOe91eME0pP/zV2
2h67XbfLbEfyqEyPjyGHluSr9aMW6msazS9DSM7QwLjZYbGJpZE1MteJxwkUlK56
4uFhxagghFNjqt6tPi+AngF8MoTaPIo1ykNR7hIK9JjsiAtOs8E4rhnF3rFVzUsW
ef6WMuSntQ8xQOoEzcBJjD4BRVsFR/ba030F57LheoSTydvBVc9E2Ytw6BJDrLcv
czoDwgY8uL55wB30LrJcOlXmr837t/LALSboq5JZUAUwqLNGfOGFVygUVf0yCvMW
OkgIruqYbhmWPbjRVlPh0MknLorRZ6qVBt0uc7NGQint8wgnYhvgiBuCQPVCGTQ4
7xz4sa9ZO2UGX63UASCO6HMIZLgRZ+gLIZdHEBuvZ489oUVhgH1+DcMS4NoBNV/y
6x5mnXlU4OR6ymrWGFcmilFAgwT/5V/H0OOriAlS0K+2MTMWGmTvMm7J9AxjLc9/
ClxpzFmt1bxCyx1oV50k0wTilwEQkEDTnUPjcW8AJoNS38lSPkUJi1PDaLZyzokK
DRveXEnvfPwyU0Uqn8pTQZTOd2dr5VDiCntV29TnSR9CvJYO2JzR+ijW+JFtRvfE
3oujub6rCEL77gwq4spB76ClVIu9NQiC6zHUVuMr0XHdgRMNKnAxKg1FMdegt0Hb
cZezx46O/9PQ9yZxlLB6noAC+AV/xkNcRCj5lD8Cr1qKY5+DOnKaToDRNdziUkqL
C3pckBiS85xJOzBPC9Xc3Ouzpus7f2SR12eGahtux6JfV72kj0HFX8YLy3AVao0T
r1n4kjyHnxOvYLvGdllP38Pr1eDMA72xoedeoaQ+zBbQ3KqFZZTQgF1vWh9Y3A5L
mmDesC+E4qKxvXGxSN1y3hVoCKxwO50JDmmA1LjzEN4t3RSObUDOgLuvpaeUGCpz
4XGVTIzCJaT657PPZGhmrPiKngTLiC2Aahr4QRWMO3aIv3B/DrVdf6FPZConn8pV
aZkxdmwRq8Bzcyg5cp1gDILPFe3NAvn8Kdo96aU16bYPGJQm6nbJEPDQQ6vqTKn8
KaTMD6sPBFCwlaKxQVBW4YkGBCQ3ubtHSMWf7AtybHinrVOSkxAqn0P6rMnu+VIk
YXEUXxEcos5yTGQjjCBs0PTvevEZFtCzFpkAE+lugIhxGX59gfNxOZ4FF+QCr2me
JtadF/0viefbV9jI5FqShkRGOzpaZJfCXylt0fhYI4qfnBQc28+vcQgKv9vxUIcf
y1BzrBZvq1vX6CbikTzDbu6xE17+dLbfoojFs7c2SX278viK2GUZ0RcYxoAi3ubZ
RYn5X/hfpNRGeOLlqRwxwP04XC8yqHzSfqHqV0bslcVVLWaeH6e5w6KFwF6MaYXn
YLmZkJaSJlOM9s27VKqb9FGZkQxv7hCihpSQMqHpS1gBmo0p+7X/FlNh6AY9NjJ5
Kf40suoKbJD2aZN8FBhyiriiKF/Xt9e/8egmlHYGMfXMBKXFEOXdQtZ3ZgvRY40B
Joq1tUfQV4SjANkj8vDE96aO00qEs/PVzfjMpqdVS8Ux7QYtv4XjVRAvy1Y1MvKZ
TqW8HhFa6JBUpKVdn+L1B2F5qdO1hTlwofrTJ5cqF0VAYEdQNIlFbhxHrOuUQEt5
YB09RMGLHKepbFNYi9ze3d/aj59noi/6SYdj89SbD9rtrJXFyzTvh2zPbujJWA5X
GDT1HqSbsJIBzdiRWwftSSBI+ukY6YPmY7LsPypOiciwHUTgOK6T5qBbX/6ZHw91
pE5tAI4sl6awwnif0o0f3aTmFIeUhTx0RrH53uWy59SYJVVG4xFRnbLV7ooLpYCx
AYQIFIXpqUjHf+vaQZk/J9tThUNwQmyBCNn9wRklOXdP/FWSvSBKiBtrFrpA4QUR
re2Z5QY97RUcKOiZ1zKbZWL8bcfCy4yOf3/7qjcmeqEh96CCtuMdNn9T2lBzHzPo
Xyqxw4BqihzFKd/t8K6W/JSYmc0oNFo7F5m3Tp0zOkJ6fzdoABj0kLrQzQPDpl6p
ZCHI4E3Uyb3KMPy0F5B8MlP7r368NFS+Xzc3qzPbWAAuUUgoBHWHsSkeykqxCYAV
1mbYLsuEvXI7sUsqJCqneIuYAuApWufXQV38MU2iSvISVeQBvFnE/08lrejWbmiM
4oaiI6nDb57A1V+tSADevegKh70waukLN29QHI7MM+3Lmq1zGIvDLNrsBEi2eX8T
7RDq0SckpVpk9EAtXqE2M9zrw9vajjtdtWhqLfB7V3iGskUWmrxIpN4JhG6xye/c
AuqjDTbAqwgg1ciIWgeq4ESkU4IbGs6xBOYpVS5n+HKkDfatBD3fBog7vk52O0Ph
chAoFTfNDRwxjHNN/nsdYgBT6xRLempCitREkv2rOWfeWRsNeRFTw++UtqxvjQOL
dyIfZEfNFL23bnmaMNzLXGe4yaFdmPZutPte8s4/1xia7dCLlelBf19/j+dYibXf
mFdVM6hR+s+x8Z4shhOO6/57o/+Oey+fFXSHq3QQ9hmc6fja8W2VdsmMRj0uIbXH
uutc6o5Q42WIWvykS+AlpoMP8TjbzTDyX/dHBJQGYp3TGSs2fuDBg1U+nvl6iCWt
65QQ1q6FyGqOUFeDxo363iUf0kSm1dB7sgr9apvAhvZDJqslo/4DFlmBKTxahSDQ
m1PwLK06vcfOrO/bi6eiAX5mq0GWoFLC66koJeXyR88llDwvqk2bksAQugWInRa5
2JFQ8JZ+1lp5VjUQyMOl1FS+VCZLrTs9kuo4jLvmAeoKkpxn7uFnD+Q5AHY6C7Se
Z0YqTqXwJX7VZ1rWSoUMoFSws2cqRb3PK7DooffLKp6GLe0rdTNuWSFaLXAsAqzi
z9GyAyxKW4etW6MyRFXl+f+w7v+cwUjpig2pb2P4vqs5JUrWajCPcGX9CGmR0m2i
ydYJhZx4hUOaAzJifBAoG6ajzPU/hWMc8fintqIWYWmy7wIXKPSkfzYS2cWrVIb8
KvyC9bckdViHKARYBuGSarXMqdQNqrfg6FH6YIBlxzSwKeM+3bu0m49XQh83v3/3
CkBt0QMf9B2fznk77XeSjbIjg2fiqiWOF+D2RbTTaSMENEPHGJ83R58KGKCvJ30U
f/Hhz2XwrHhqma1P1HcVwMWBXuLlT76gY5o7s5bZOb4J1op9RQQ+N/CvXCjltbu3
neoYQHvUNXoL5hxL9IdS/SawunJG7cuEuSpx8jTzWoLyiLh3hBNKkMUoCT0z77bM
eEVF6bh1glHa33MQGW7cNg0Ee6vJiHBKcYLi7CBCzf5VqecHDu1yZxHRKRKWCBbW
LhVCAHzMrJ2uSYSbP6MMK+h9hol2F9H97uU/zCF0/SlyrG1Y/WM4+MTnK/hvaEuq
tB2plFpOVuPn3JI5ikU1w5Dg+jZOAzqyB8wDf2V3TZo6Ymj3vBMVi1TPo5BACYIE
1AToucXTc+WNYAr8a2OlpcKi3bU0ak58DLx8J3WwxymNb5S4p4/n1JkH68cXd4NW
ogDWUWvyeSR07hmM5C6W+2enTiZjBp2dOPS9BOmHWDt2McdnlfAg4P7jajX07v8O
0DCyAz7+KO7eEEnPXx6KhPm910N+q1dTRmeryJZjk0uftmC4PGz8y0QJ0l4z76Iq
PEG+hAYRx7JqB2mMG3vDatC0lsnhSRF3ri9JR92DLGK43c3WV6DNtUCBOMKuNtEi
lfxfUUpnplKQHUAhAopwnaQDk5eYmZ8VsQxh1xRD8E1ODazqSxLzazBUfmEHSSOb
bFU2KoHYqAZMWew1ED3as8l87MUIqsvgCp1+1If6mwQX/1RG6pGWLmvxzk4wzugC
ZFmY/bIYipNNdrQ0Ucr5cVV0otgI40j1p31TWafTvJbSFZKL+bznQ7BOvKhuU/lS
w8fh24Y/9uazpjoa/OFZDufEjUnAlOYfUPAjkjRjBAoCdG7QGQHmLT84C1KsdCpa
g1PQOW2lo1KaeTrSlt5BGHtIyNWnvhmvexQD8OJU/zJDYHYzQOsnZpCBUCytRU++
w3Uzj30WPkQJUqP49LoWMBJ4h2ndLzXwwX3NLalC1htz+sMcjZ2ujhKxbThwSIqZ
3UvxNKMece/JOfumN+g0CzPsLb2umOj/l81p6ZgbishIqUSWRCV8mRYwJGdm/vjN
OTfGzRowju18A3hB+eryNFHKG/9d8XCyXX5ZKjt5T9h4qXiGarn9mypAIDbBoL+h
jJYn3itU6X+adecIQ3CBuhejrorern5CQiJTkGDCYwwNH1JIu4BLhQbMv6NZ0yfd
k9ipOKLqczQKiO5mx34NGl/1WPyOVGlBfIesHpIiEWys1UQviQjCGlQfxKCXsgbI
`protect END_PROTECTED
