`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OCdXA636hfkE5giS2VVWrcm3ojEAhJkxCgyhHe8+CBu6ihUFtskAADdx2DEAEIXi
xNp9XsNKd9opO7szMPK3LIqQU7jGEYEOFJPH+IMNiVT1kSfmqK9KTZRR9xroeIg9
Y/R8SS0Btuf8sQsZwZkb6+v0AcuNeP6WZinotjK+PAOYEeJaejde0hFb+bMckO4R
CoXia4b7WBdvDySgQygyUAkI5D3d786BzWs72BNzHBCfwhF7b+jDzSqpVMv0Qg7U
YevCnFJv5iKV6tKjq04U349X8hZdaKF+JITSPXpXwTbQuBMMtQFC9Fh1YQvQ8gkm
bnXuSk7wA4VZzloUg7XN2fSTr4E2/wtYljR8NnJ3drGNGpK9M9j0bCG6+GxFRFpA
Ye42njVhjqCk+bQHNJnUL1AqVdKfm1znS1lI4bzET6iwnJ8X8eEsFZnYE46NKMiq
GwYygRHfTybjXTZ+YeRSgrJV1bg/GeiypZv66eOAj9vRP8GPZblI+OXoJLIKJ20+
pp6sLv09/kkSD2TliKmZM5Izvlk1HCcc66/YRxLCFWEBjbrbSaurj21b6ybooCc1
IamSsSCgZGbN+FD1UIQhAUif+D8OapPNoz/D98Lam2xinPd5IHlBbQMJeDCCnmMI
Kr+9JvRKvfeDhsnIdrnBYF8Xmt2TnFYjcGkwTA5CUGUoI6SvbglE0LFb8dCtc2OQ
nrVJFH9UwNrcHYHb1YGcQb+3lqE/CtRR1ZZKOmxl5h11Gu/GL6EUiLJYiOoaGqpg
pnl07suNR1BEc40bVNjm3WO4sul0inKEH9AjtGY7CqYJRaXKHZ8juz0VCZKxkzTr
9mzlULyq1mVPgXYcyen5ZJn92J5zD8t77wdnTuJFRRMBdVLMyo7t81MR7gTyYlqC
0GcXXoW6uUbOORxsJWa3ZRu/QaHTF+zcNbPf7IGX6xfRCUGISVGyGSxx179dV7zy
hXsgebACLyIQUN1IeFjca+C/E8HLstSFDJJ4jr3LJBOVWupTkoBU8NRbS5nAiOHS
RnA0KC8b38mkt1qUZ+dKDpPToW+6JGTk/13xQa7Bf0b6RBNTDHXgPIOzBvOU7tfY
`protect END_PROTECTED
