`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tIL3d8iqonG2IiDn+EFdQoxBv+v30rUfU2v3HuvoZpHpcIhGnHlP9l39hDh5nj4d
dVb8vWyGfjSQL+bHL6BmwtL01nnC8If+4jVcSMWbEMRHD40pzT3sRwmvg47lQ/4R
ZrQ7aBlvDqJ2lpIttZuvVvj0n7Hv09L2bBpGAS2+aPBjvKrE/u/DbZx/14xhTq8q
gPqwTf+aG3+aSd+7uFoKAte+gyWHRQ38LD0BnTBhhquvOLWiNpEt0UWGV1KPEKwb
/auH6giP4BrViVv3RkOJL7vgPhcfUwjhpiok+K2+J7vyCyFYyTO3THdtfsTquJUq
LP4w0eqn8fISSrbXis2tKx01FORONH/2S9Kw8isUDHH0VAKPLO30SIU8lthhilxG
iZg0Yrz6vM30lzGD0fliu1Qxguz2XdkndzW5ekbpCjl6AiMvZ6cwtB3kBKWL7Wtj
2q92foSwOVHbpFKR4i/HHWuNBwA/jf5pa+I3D0Jx1zc=
`protect END_PROTECTED
