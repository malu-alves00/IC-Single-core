`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BEyf3SqVZdEPUnlZO/ODBCzmoLIyAr3cea6TFuAO0fw+hjnDGSPNbBH/68vObUda
UxMHRlZVCkuXExBQnHL9qfVT9E05I1/Y4CfMhl5pB8GVh9xO9cQEZa9/UuR73NAv
g9E+Cfzf9VP8ALMyPxUtfltcRyPM4hoDVFalQCr+FHzfE3IwhRhp+lthYf+idk3M
75xl2YWnd9KsrTpN9nMv0svJ+ab76baA5uWPzdXAkvc2vmEZy/DmEMFguyiOmmIk
q80ReBK9K3uz337/9yHKKALdPinZTrJq0l2VD/YnDvo7Ek7UJx3mO05KQOKFVo0O
CZ4qOVOQ0PYBvQhTbtF9tr2gD9492AMwXUy5+sCQ2aBZ1aYWIc2AywPIa20JJiL6
UHGWc4sYCnoqnYa6/ssWpg==
`protect END_PROTECTED
