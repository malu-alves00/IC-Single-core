`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ViEIvB/s641Z0SUmTZFElWD6YLXOPVvISZhJB927+7efVGTSsDzQPXPN2Nlpg38K
8NzF+9HuWxTEY6H7M2laJIQnaBtUlMq2APT6oUjPyml5BSeZKO0+oRsUPl25C93f
ZRw5SBMhj2mwuwPoryHkOsh/7oki9yHw1fsTUkWBf2nOIik6opCsdA1lSit5ouRg
LMcHFy9397nsRjvR6KjrJQKOAgiJoTrVgGiUWyCNevstR37MpxERzCKyCyJSfyCN
BvNh1hMWL2UF4TBXVHy594QCoqEaTVbcAeAFsclwn+xslUi6v8TfTvg44YuKR4+n
2XQZQoEAL/SlV5BdDt0KtC1iceV1LpktPkd85uT9FaNZghk1v1tYXcsDjdE7mt0L
NSu6sbWzcZ96pjK2hH3OEEwvb0UwLNmJ/+kNB/PQaDYYDgQO1FkjTW/D0rApo3x0
gjFxomCwlq6ChXI7kXv+bod5gvPrs6LmIouj8aDxJHlCLjrdB1/uNZIffaWtg66D
/58DFMHTs5MBQM1FvZVnOLFk58nxLdkdTb/hJ2MdAze8tbadDtt1V8ie4BT71Mo8
hQGspQjtjzDO4tf4fF70dT0JRBXNIbneR156+gdVVAI9xBU8NWn1u9ot+lNZzoVX
69m3fvd38eQAMA1/7Kz+VWyiFjwQOosh2k2APuT8FsPgbLGQVBTRVlXjRDrSFDoQ
dDO7TbwN58RFytDJ3ns15psdjrVndEZrEzytpZLDGN80FHFugGwcRmg/vOY4kwmr
ykB9P1FlYHdVcuT9/OP72u6uYGbRyWNVq0PmUSBx6HH/TrIBtkTcoI8VpNRVGZ/8
6oUYbVEy7znw5FZUKz+rug3drrbMAWYFr3R0mXU5Ml7V/L7X+bPI70m7MaTodzUb
8EDpHurTQT954PDmz5y2mxFiUy5mee18uLMB9fTe0gXQtrhBKMgZ1rsNO0AkYqwS
q4Wvov2JxOxhZ51agnUPZFkBshUD6uZIh/3fFD1LqD8Fe+e4zkQpaDIre9VXKzUo
EC/DyG6QQXWyM9tTT+zKsE0n8hfU7c1GKdG0qReyMXGRRk/Xd/JjFw5SpdoogSI1
ejzNqbLtfRHZ1+JyjpW6wfCfchAbzkxPmCyiFQcl3R7hsElGpUnoWWzv/5FhdY0w
foisSRzC61ehv9/qD/9FSQM5VwcwoHRSB0L5hVcJWY3vsSn3AxHrqSnAUpxfGO2y
Jl3yyQzMUNVi6tSMFCSb9WoeRw9W29CfCx9IQNV5vfDU0rDmICYNeL02HauKEnVC
egYiAgcR5vz4H2sqiW/bkrWocswVtPna6ljk4toam72OaFgVeHKA7FqDcV6nCoL7
o1eE9Ii48ex5ymzLCt371XlMfqGRMJozv5JzeS40L1QchADGQRxLQaLCTAVcKEja
Kh5mwXUZhR8kNOmmipkx2x2REgjJ/goBKnOXCV5EB8C0jcQKcVXs4/QE5aJoaAY2
ZoPMpX8GlLVmMlyZf3BgtDkg6TIbWwvjEbH0RzCTyRVkEp/ljAPt61uuC0ugLW76
Kr+nIVx/RYXq3EPYtTW3pQDBPhXtfaxBI1JeyHTQ3mXmMckExPPJbSmQjL4LlgS+
IYbdzIgyiGtcE4OBuYb10xLpZ4dn2yMxvLvDEiJfPxLE1OiDrEoLQ1YqiDFZLtap
de4Kx5w9tCGlz1Ry4ZDVMW5BwNkIEJNWDnOYmtAtxC+3UQCW+t7v8ij6M0IajMOk
KIozVE2K2sJe+ufUZFvAgCjfVS0QgOYYDT+FBJtwMH7t8A1YcFziE3fMaEUcRMZD
fQAEb6L/4CZjLKNNjTE3S4edgxnfLCtPJtqwfvSPgOwS1XIeFTNF74ZP3yBSkk7A
S4vJPTp+bpn1sFwW//wDWh6T534kGAc+7VTPb1I8fvAOWTbDDM64Lw7E9UrfEzE+
VMyaV/XhUg6EL7ewsoxyu61rBfXGkpHd0iE9gT2TjQqe404BRFwok9K51ocbEKmg
Gmqq70JM4ocCmoE0/sXOPJT1J972uXwugvu6KUMRkeeIztSlo4uaV8F08H7dCSiz
9rBe9dOFL0ArUbU2pSu1jtGmJaPI5jVRm2pFoRw75HhOBnkL7usrguxe/wfAQ4Xu
Ryj3RGhT3LHSts+5CkDIQY8Cwtg1gveMwbCYfEEWUbqPiS+Wng+g6KeKmy6TbxXt
j8vZl0GgoR3hOgOUlam7v/SIUKmPihyXYrhsQKEGLdynwor/8lwvHrGaMgNCmLKJ
/5LUJJgBCkmm1I2qelQyh0KcyYvN87zuR0GpwUELiyux6zhBtPnh4Zf0zoR6eZGD
eI6Uds4rxW7uv7IrqkaYWiUnJZHCb7AV7qxBjhICKgoxpdB8ewKpNO8IOebJ5mwe
JpEc0JQGWl9TRHTh4eRdfxmoAAx841cetAh3VIFFJaH2YCczcvZ81nmNBGYGIlrK
HKBm4p+706lyZwkpZ29qHjXHbCQXaY9jTOtZR7mk1zeL1e/gNUqy9MxyTj6lYd2V
I2ZiH7VBGAlJy9JafXepfjB54gtsfR+x2cv8rZfkiTJtJNzRYPJvgD7sND8uejn7
DrZ/Dolr04eS2yWMTa4hzOe8ONGtupYPWtFPMqVcvLk=
`protect END_PROTECTED
