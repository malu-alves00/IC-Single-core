`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Or83nTWm6sS7VYeeIzx7tXswEZ5q1vKAI8Xgtr81So0mEXkYIL3fAaTYYJtpz1D8
dHkUjBahA+FG5XF6SQOa2f8110taY6ElCZXfiv5jY8oKgVjluXBUit7Kanh5Qwxj
S+k9XTRNGBaBL0y3fdcmVDJL9UgUQ5PXyD3nbwkENbd3WWOu+XRNCY+pZo3v0Lvc
ze3usShLbWPH0ZWgS8QXNeA9qHtuTnRR5FASmXhNnRdDbDRZ97z2Rg4ROZlXRT8S
4Hlz0HrY3pqxMUiuiN+6llsewSWq2duxfCB+K9aDHdALNCpffazYvSmmi+ZlN2aN
DjgXmuYWhF2/PheFrjP9MjLnkzRW2qzjPSi2RsEnfdQmAUjIJdz32x0l+WNUKs4k
cAULYPR1sD2EKw7Mj6CQZ2ryWxPl229zU8uAKf3y+aJe3lOWmXr9EvluN7oYFXZc
7pyQLzcnPTxpdE377rbLmIG9hPqXnxsAmwbwdy0ATM8SHrF8HVu3b4bJnT9WWP4R
CIEiUwak46AmcnXmZteP00wtIDM75a9ee8DdAMhNRk0NSBDI225ufhKJAi0D/ilC
jLLa7Ma8jFIoXUoNKDFYLS3f737toUWPY1OhtbGBhbLvyOBWoT/vnbWdEhORZWTW
DE80ud2P+U4/VdyUEHS7XDNs7kyb0Hz9Vz03hB/9xaZZD6Q6lw7xX80Q3ZVaBkw4
XjEm3dxN3hNj2FOZFVGEUJ3jxzAZ4rLcZX6BZWwKBfc=
`protect END_PROTECTED
