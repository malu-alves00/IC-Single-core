`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
k8NOItO2JY4OIuwIhy8X+1va/b6BCXcwhV/9BpU27jJrBh0xaIar1HuP1ITx5GKy
aId9L1YekNoCubgUCr+cYtL3LPI8qXBRsU0PyE1CdPnc8xtGzaPDtQim1fX2ysro
Gc6pt/SHcbVxluNoh7SzdOMszXAMd8MEVG5AYqox1Ig8r0BgwlmRIwIxNXNnWdu0
ebbncbSkcCIEmuZhmp4arDJNZsPCC/139+1NSOWwMc+CdUOz2W7E6GtZVNqw+MoU
lCRB6Jo4YjRb5HLaPqkzuUvHzy32cGCSDCFnlDGjdnhLcJXHk3GQiUosIOjyBso8
cBvohYzmgHmwec7OeOOBif8LU1mUSQLG6vxB2te3ofCPtrMmNH2lN+JH/0OcBt65
hCLFSX4es77oNzFu+5DA544cYzIbATJ4LBGd3c8M8VkAauMt7ECAAjZjsWDy8irB
BEyzCKVHIr7EIChX6geXHMRI3ru92gXPlt4xXscQZYiL8MkbIg3/9IhS467tlKHT
t/xTgHXXdqH3E/hxuEPeSADN2tKCXnKhFB77l2/ho7XnlzPKaWzhdn1Tt6rnjUtc
tjzcwCA5HU+8McNfpkFEX45maPb6KY0iY3Uj2nBPU6iU8f6YCXBGJhw52Uwb0/Ox
HHc4TqnArb5vicUyOIpI4B9apUTtQb3ZFGdr+elh3NDL54gEb3D0bf0qGWHUo8tF
qzOBk/m+1dSYty+hx2Ey7MjdIFtAiQWC2Hi4cCdDYKEZIv84z1PxdiKD04AeGqRY
mg/ajxA7l/bPCG74JgmrHnGMRbjixX2PjnkLSZV9FrpAbJ2rr2zWtMyI3Rr3hDiq
XYg3RPxNJAZWnDSDMLAVW1IJoiV9ICBXbB197C5QcFaJEzx79a45WLRL85eFaBQo
pYfpyQhKmThLbS1FJ0m2p0Ye7R1/hDVJstaVtWfqA45ALWdkyQOOK7M/BKTBe085
5NmFNrLAANl/9bvliv40xdQzGvVcmr0BBtQad5bGr0ageqAdg8esjOmPv5xcX90b
LWq9xj6gdAZz+zKGKmO1VUu/4ur4X00LokXWIiCSHQFKS73nIK6HSi9OZx7aWSyx
6Qkqe6qiI2yuxygbuNUL9e8IYA77ofO1Ts9FyOxTNSR/11vCXI2ecdzvrRRulLf/
q6Dapu8VZwsQopJgucbAX+F9RmiFaZ9/vOKHmO0T2JHPzY53n7pIiSS5VxITL/6P
vShlrU6x5gXGJBXfUksWu6mhW/UmTL3T6MNGwIibI6V2v0VdDeXTqNreD9oF2tm2
aPyBR7J4VGG8NmxOGCsEEk2Ec2z/kGsRh8LEyisEEUg060yVCsRY8hpRn9W0jzWz
zrbWPOToYkRaYvGsUxFmyjo91Jqjm3+iCL3PCiNwbbB8bp/RoXtCBsm67Yv+4UIB
G0MUAuim66thejvHh2gXw++iC+qztLhVGzS7cgbeHpkdlmX2JMhvkIROFvJzEUoQ
m5vglRd4113GHR2Nh9AjL1PyJ4Ii15iU8y2tjSJrjqg2ixwD07RtMVgm2ER0D1Oz
2z4yNvIYfR1UtpHpOy8CWd/yrO8uatnVmBfKAS/V38wUm7WubZLl6HsMBOeP2sd0
fPPn2/s/Ngi+aRPr6KJevt6NzokI3TjkMpCU6J9SQzbjrVdAgtLkyMa6Y4v24GXX
ithiXui25FmQLurnnPDw+AmmfHgYHMxSflI8TyzPByv+uRybQSAl2bDFVD2wwip4
6dbosuAh/O+8GrhiPPIgWLN4NT/9LXo+KisqyCgrA5MeRudWy2Xvjx9rYH7Uapoq
PtXZlpy4oF/KuYdv0c9BUcjNcqh+JmZ14Pr1P+HG34jyd+c3JqohA8n8+AcqOcRX
4va8rrdUeJW1QdQosF+Df147WnMblVY9WI90ixmsVJgsvmsKijua6Jj1AI2aV9qk
jCYyW1phlKxM+ShwABv/6mFGAFMBPTEzRXCfmJw0Vln80r5zyQjdCIZIBm6o2nG6
aANn5+yMROk0ihM7bdcetMbhOKo9Rulsn4AQV/tZYI1t5XIlUmos+RjAVsWSp9cf
F8jCvn80G7WyYsK9Rs0k1mPigrQMw1UQMyiUDKtTXPedODQ5ZE94yvgp1BZUrssj
AGl8wj0lRbC1bvgi0fUjRCRFXHaKI/nezOt92aFNtVnbUmosigFhrX6NoKILe34f
mTownQF14TLJGIfKOzVx5RJlpWFjTi4cR4swUmnO+tUhtiFTIX61pt0Sv5WggbAX
OPSP1LrPwhazK9YX7bc5AUXUkyK3+EygbBLVG+8bNmVKVGLfHm8Pl3O5kSK9mysS
QUU5yNNRqskO2zBIPnKqXXWjODP0zAA2EwC2o8PDRiX6OHF4fgI1Y1rUtUAAZzHd
9uQtUjoLXuKiWzOs8bXdOZqQbiw5BT7PIZeUyFi1GqN5780eMH0ORCe2PyD5GGXe
KZ2rPzHL0ReJUNjmrVgOJsn6DvfeeWMcx4Qmcgx2a6B4klnEh+JkHPpLQu/Xq0EX
qwNWjCMDY2NJPovtOY/8WpPU8wPoiPoqDOtWnM+WuCFg+Hh3aiuBMFOqtC5mxzYO
k/KP9/eIoQxZOfNwckfCWTAyZxwZJqWOEXINN0AV9zNSE7dVz3+Qjbk3nlzC4y+W
PjXiJ7fe2p5Fy1iRHbsc2aMmnKq4piQA/odjXynL4RmfTUTfqJAG7ORuGrZZ/Ye0
o38UllgbFBZSarKwR5VYRZiXTBOKQtifoaxyZAl2J1KlwLqi4MrDzuqIhc14l9tw
xecPkWKmHpB1V+jPSt1q5UV3ZHuwWZUUnp0PdGFbjYMJ6DBfMWy8B/gWPFPDIgsL
FtywZipZKn1h/Z0U76VptJ5FnuCl07CTobp+BrVniSGUFS298HdcURh6UM5xituY
ky0HP5Lys202L3HFpoL9osr0j7mQlCppKC/5+Vn6PxkJ8cWE9jWDqqBdZ9nyQWiL
swK5nZThbRtUQCHXcrNQRL4HoLXldgQx8LIQ8/RYTvpjxf1CPaY978Lu8SLuT8cb
cEs64tefa+nuIrEZuDjZpqgAWNTdmF7IZtys/aBk/C5LhMR1SPQ4f8PQVCMjD+tE
Poyyobf8QQM4/Wy5grwuUH9ZEY3VoNZfiTdcoTW6KKQk4SiMI8hzwOjrtmyjNSyA
QUvW8Ey/RrrCq41ht29wPpgPPEut0ogxIFJrzlrFNNnTtSEJwLgtEelGj31qJ17N
xjye86i6ptujVvxw7fcfk4ydQFx/w830QPoJ29hP+705F+Mh7IibmEcQlTpPfFoC
08eOrNZ4gxbgNhz8eKfQyXZWlCzgXFxA858s0utavwi3vnafbBGVUFJvHfPmoKaV
hT8htavGA1Cd5srEe26dKMRGx4GBRzOcTl+h0EgVSOP3cWOTHjduFiFLkIV4eWrr
qPPtByWOoPo+BK5A/VHfeWRCmcVOStO2zbvDJ5YMkDuqEkpyatlWuVxr5lUIwM4x
IpFEte3N5mhy8oTMP3oJSU9nHHbllKyZFmQTanpKghXRRL4F7jF1RdxckU2mMBp1
GHANDM9mJnrew1K1m/YAkzySAjVVmCZHzDmy5O68WY0LXO9RLJcH5Q3zxt+OcIQI
UYf5SiBreFPOMZnLTetxPIooUU15TK3Ne1bOigQpqnCoYWoGe7UTQbghlxyFJ81c
GWK12S+NKJzSFx/K7prt0ZdqLwrWozChHgHcdO9Qru8ezMr7hLq2OEp41xtZZqwp
AHTomYsGLmMFD6stDkVvFVXBWvVmc3YnevEMUNaw4Q1gFPrdNCx4Czhnmto2CeVV
T7J8fpqpNRSduWvvdjOc43Sgr1Nglbl1AbYpZl8bcWoqgWikML6gARB4iGXc0G6l
EcpyPJLz8qS6Q/g4whJ8G+V/Lo+3ewqCeFWfizBwpvGob+d6Q2RbkKmuIymAZIpe
x09YbyxOXSwv2tdgSj3MBnaRLSaSf81uyAf2GvU8oixrkYcF5To073t9KT19bgWF
Zxt9oyoILpQZc2umYxNPmIyCLNAwp7cVOxbOTaYX4lTdmcI3H/49pBHMx8Pxga3g
39Ed6VfJUVEhPmW86r+piQpSzEKmQqCVe0+QpJ8OC3Q5fHy/cHlLk6xoXdEjfSp2
4kl1Xg2xJqkynjMqpheJeOIagvod2oY0uocxOzn1SUIPat5KLnDxCJ2mVjw68A54
6Er6h/8Mgak4+u+1nKAwpIT+gLaSOLxqL69jPnNLX4SNkwPY7NJRiRaUKu7HNkKA
+6E+GxgZ7z7BNQD7NVOw+Csd420bML5/KR4EuJkLo/D595VKQeq0YEAx7El7uZ/J
zONkHrWVfa1Y6pJB0WZKMJmoVvTgj/n1Bgrb2BknwSuI9F5+8NpPGwinSKndqAlf
TBI+hLscwaRLkmJQAjrlpmfmEm8KNDAUV/4eAOlaoeJZHIrdiWOD/r4H9o3s+Ylp
HSuf534sS6W1MwBsXGjDym0+cNCrCW3MWTyMc9XquPNFib9OibkLY3JkmaE/JUSH
VCfmqCKcSAn2uHpI+MMXRMtyEfe7N8DEkzm3ICX13MCdhx1CAfejeHhrMitn3jpn
LeQz+FKBIUkWlWgjdhiHBihS72A7GHqgDoxckRuJtivjxgg/WnEt66SHfWqU2NLc
rvid5MwQl1TA749zc8s7ut/TOGGdHnb6TytTegnfFA0zQr6UvYpwlodKzi8OYoIk
5O2RwK6rjFzsMrkVvhSkKUKOPuwBf2RzrMzyCETb2loUOqujgb9jU/uG6KIjNBiK
C9Go6XIgAt+bsP9fSKzXdPu6PfbirfiyyMDIWJxMOsFUmnF0h/SzflqPpR6QX09p
vVxPpcHCMzzvSo9Um316pKtskDHOPcFJ0undP8Q3rR0j3N/g9OTJOsls/uL7aVED
4y2aPziIypZyKVw2hOC/pILkaYgNNQdpInr4u7TT+JIjQ8DT1NaAWWPI849fWV7H
8LCANNnHj0E/rp9J17MBSioEX3sxkOG+PaDfozDuXeXqsk2/zeSmmMVQ7s1ieQvc
HEC1bPpqhFvv5UAV7P1BvOysOCWgtqko6Mj//B/TuIL3Y5DOr3do5X2hkH7dZeD9
3Flh2q2C1u7GucLbASZKauppVMXmm0BpIuCFinKaGR805hivGZ6sVhAHnq1NvaPA
h06urGr55CsdGZVAI4ImZoux+jd5/IwHHB0ZKr4AlNAyRlFPbL7jAaw2TSGzcm0p
Fz+rNkvbI4/7iRumSseAaIEsCPzD91M4wt+fCN2/sOW0K7nNaA9+y2HoHexResPH
sKeClUQ10eJ26mdX57LfzvKsbh1Lb2F648coQucKAlT5Pw79buemNBsxwvKFDeC1
w3ZEbCQZ+fw0RtZmfLbhIaUvyyaSNgbv+wb232MXv+moRCR1pjixHdGabAaZ2/E2
0Z5wArojlVKxU+4yC2Qwb4rU0vaZiClvbues8TAk52x7bCKFxihROupj63H+mHJH
+677kZA/3obyalGohGsRqTPg4UeHavR3ba5ivjZ4jyWMqoJCqcXAWUtBZzdUls/B
hXCYS//ZmjGcmnF/KhfCWyyIK+iTWhWyJrrujX+fm949KtY5HmrQt8q9PvLWRQnI
1YD5ym1EzKarFWTbZOJPwjg4jB3aIDX1YizldQFU68UzNiZQl0HDslGjZKU0jT9u
2FtHu0W/Lj8PdT4Rp/sxiMjA6Hz43qk3+m65CdbSWnBKT6WWMXV+ImCneD2BMLSi
yQ976b4ZteODHvofdQRlvJXObivsff0whwdjW9OT6wgptEwdGw6EDGCEaG++JXst
rD384lFYQV3XN6+yg0TD7cjxlDxxZ8DmfWX3ihvNkYMQKu620Ar1MURZsEET5T64
PKK6NUULA2cx71qmrSn5JP8cJjHAoZqP4gkk0XccfWZYNHzS4BzNSs9Teu0W2Kbl
J2xcz6+O32KSVhzkC8ak0bl2YghRsKZEPf4ZcrpuWSQyT48Ks1UTw6x0kgyxo9f3
rgJuOCYMf7tkYdqNTjggS+fGEyjso7cuB7FgLciFhIMvFalCpuLidjy/0WQR0AlR
dwrGmQP9sIZm98IJRHb8uiaG/kS7Ggz8Ldp4ezsGxUe6flnp4HKBj1qOz/+/Wl1D
otiPinsjyrqJVMS+nqEB/kDFgMpYAyYqnN8rIEZT8raAV36GHFLGAOFUHggxBHxO
1JmzgHY9pt8/fttoZURIGMuh1YcjoOnb4g9MqcKUfmn3A7YI9wXfUqICJetoUbFR
lYIrv97bivq5rLpbPjMGxLVtmpe09yAPkU4Wo1NcrGqr0t2Eb4tAJ1RYT3CBX+1u
spgJu5fH3OlXPruaO4fo7BEnXEXOC/foGhrmtgZdlX2sxpd2sM51hhKBKFInP2K1
aW4PBaD3OA7n1kHrl7/UsX+xl/mVaayzjTJp2E7pbrzUrFEWbrgPSjPGAY/u97+/
xiVEeFhVDuoOjQD4bvb7N2pH1glPSMWEFOyxgL8bUz6cSeBJsr4SPRVXqfPUDR/F
/pAJspxKulbgnbHU5fNnUIcZoulT9fTRnf6ju9PElgnh+krHjHqMvIiICGFHsgHU
Yr2Q7rZPSOFtuaewPjg3mOVw1FcVMJttpYrGFOzrIvy1EtHD1ynES2JNOPG1Tqg1
gNZxRVrjZslsqxBYs7LmHJmMMa2FSPDoXHy2P/kHR3JD6SY2cu9TEJNrnxJ8s5Zc
v85HVZR2ZLkma259NOfb887yq/l6l+tGRZ+IMYmxLafBjFkeCaSqftlg9FiVkTGF
06y97E53vBkOk1Aoe7PXFFZQ5dY7X6D5fLtSreXrLhp+bwCfpKF6N1pVBE3CPzEs
xxyO4Q1S8PUOqekGIf2EGECoaeN7CZwu5Khlz7LRAkTLCekiVBXu2JtUDe7jsZsa
n9nsqdXFIs2mhP0dHlRF9HvLxSTIcgZxBvQanQ88dkOQk8A8IpPbVy/yIFJG+aWm
FUEYBxU2K+iAfBrjdUmC38QrvyO7DAVjbmq9FB0Xm3txiPlKjYCmWJqHV0//dg3V
RkeZegGwEkuL9Ny/HHuRnatIje/3YhMLz0WirTjb2LC7jNfHFEEmD7HnKT3AjZBx
Gfij2Lu3mNH635WrdICpGUlI93SRW+GvCutjHdWD4CWOxlrmiDKIX+8WVtVRQP15
FNtJDLySWkvz2r9wIVMYh1aPmVAuJtS0pFqzp56ACb9Q3jpQ+dhnxFxRI4jhpPMK
5bGfNjUJTjrGKHzG+21/73r7pQteEAgVUhplvazP0OOk/4WTnGtkK5Cfefk2PXyM
Jw6kFxixV+r/mzXwASKEyWJhhkZ536Ssn1Zvi2DyFawzbuadRBw0HL4xBycZzhC0
qeivaHGp8NT88Mae8Oq1OHUHvAmGZZnpkvdM/SEndIlc8LEJ6n2D9W/qsYw++gI3
cMaPnsFnxvDQHgG3AJT7PABLUwbbumAJ9UCGczxBLN5hqFHVlklLco7KANSKs8h5
ZO0GLYMtxMBIhRVpHCKDtEXnqWLnlXym2Y/VTPaRwuJzh6c3LB5XYFsqUy3O6Mq9
3BK2gYM9Ln6Ercy5Goi4EC8EPBIRw+NKSplNBMk0hP29eR1ATgOcVU3WF4Tocvmm
/vZOaYpEhJvyu2ZX0EuLkkBBBZbOEnq8n6RxID7Quf0+GYMlP4hlfSeqTgw+wTO+
3ioaPXf4j1jmjF8ooTS9iTEJ0kqVkHT7XLOmuGpZZXQop9ZJeflkeoHX3pJZNLQO
wARn0AKYKRxqAIb/YqsCyus88iRnC6ArfxrbLA7oJV/kzr4jvAV8IkFSiyXERL0p
GwBlngI++kK2O8lwLux7bP/L5U7Ajy9eGy1w3qFZdZhQc+PHamZuKJMvWkGc07E8
BIK/99uFovEmXvpwrHbVInBtakKDn4rpFoBY5Ai07AVlo9cL80j55kDl0GyB8WDd
A3G9NGKMlqNHMS0nNKMwl0udwugq/38NQJVCEEosM93gapPoVp/FUBz+KPQh+nEW
eECTxRIEjsACw6z0WgUyEy6jwRNtt2hVBeGrbbb26Uq37YzItUehAiQ5grC6T5MO
FPVYUJKsKvYk1qS1AW/I8oKoyl+PsmBeV3dnOYId2Aozlfa8bxFSacT9rUBNsHg9
Kh+MI4j4Tcyf2DpglF6TpkVWE5oGu72aAQIOh6d9HjlYrn5+qy2VrvUamGW0z82i
QX3OKIXdlwW9lW2jRzAYBWLGxQzIlT0dT51gLSwWr20Ow/SFYitCa9jp4KNt90JW
aJNV92HJ9tXV4xcCvFfgfwA3+GNvkBZuLfvr7rUNYwzYDUo5slVufErxVIyuvbH6
C3yi0L7KFMyw2mYGJ48PSi14oLjkXGjkwJRm0XsLQShSkFhlVtF3dgdTgTi3irPR
ffw14qk9uBNqS7pudaq1hfqP3LxuRT1k4uY9EoZZi5W+UH1EBZl04tiYtg0w3H0w
c9ifmoCTCBqUwPtGedBFRCnZ8U+Gl5CQI8wqIvZN5H0uf8+zRW7sbomNsLpk6sI7
SeEGWuwHvWn4Mc/YjAtv3jD28NlN1P+T0ZBNi+elX2k7zzSu8sBiO4ouFCmUeZNx
u2LzxdIhjTzF5fQjpRb63FeQ8sPJLAZKTUrH7NJNUlK/rfTCgqPhn4vTlqURHohH
I0PEU5tKaOarg89rkrP0vCzrTx7s9s+hP5sKNghQTAErLCUPxncKxE85p9JvNi2O
DS2R1d2dyADtRMNboUaztHwUknChpWpDE9eKM1qadXRRKP4Ihh9HIZdyZtlQ4I6H
iz9FjzVtNCwkyGPHDp4nLPRczzqm4abE2vJ199Q5p42G3MTrUFya9I41hyfqmLTt
P4yCa3FFve5Us1TvZjlUtcdJtmGcmAfoHXGg3xAQ31A1ZYOuIBnjysxt5J6+1Xcg
yyK+m7eDeTWo141bdoV1gJ4TQ6XeDVmlHNJXqhhcokBEcAlToQkNmG22vDuG0Wh3
QRLTj7ONjOjMK97XDAQRywcWsZhHIRVeuexaK2Y8QCje5QxALxJzOUd6DGw/6Zpg
uSdnsrLAwvt+pkXUXYu24Pdsb77oTCN9ID/f1ilqsvOaNFs2E+pxk+XeD6whEllV
PFFYIM8X+GXZuqnT81Ue89Y0UiSXCwFhPmsl0+8qM4+E3QLhjNuxjkR9/7xu0CkX
21TfSOq/3HNvD9/vQxwgJXiK8L+WVaOEuNFEMMbwRT780NgrAc+NOvjAx9uu5QFT
ty/yVHWhnZNHhNXogm8CSC8asXr+hyQ40zMs7m9HeIzdQksC0StLUaexFNaHVOck
RRNKg5CmjoJT/oIgC3vd9OrbpmUTrVcjRPn9cYgVzCWP+FSreACJH9BEyRkstB5n
y2dw6R6FlHat2Rj50GggvfyzK5keAb4ZiPMpy8L31joXwCPxnq7ppsPDSPjgYcCT
XeuyEVJ/hlcLrBtoAD2uFnCCGAesjXaFVd54ZGxOW5rWwSmfNoaltBkoEQHv1OUP
BOMxKEWIUdVqY521vEHgzZ0Eae1N1b4Xa5128D0o+7Da50wh5mJ4vFQSHJ/GBKEP
A6XDT9FGkD8Iz7f9rqgd7kmrIDTewZEV7v82Rm9ocXYKkqrT6cLBBfulm2uGxys3
b/MWUeK+co0dPcoOsI/f4hIHNE+ED9trIuxHHjDIDg6YIfdyEBalRz7cX3pAZrgv
O/5w/haq4WC07ML5SWgXt3B3GlePztsxc2Ahp+39j4bxi5NZbwr2JmF70d0KO9Y0
vGOVPpe0T9Qcy3Renl5G7WDD8Pm2dFjQ36n1lknrcP1EQzl8QeVsOqiMD3yrk3ao
J00BJqDgMJU+4YV3ezecPdM9IfIyF+2OIrSuUr/H2VWRyp1jq0s7Pf33iBet1Z1L
i/sHB92ZqeuHOoz5S5Z6dP5qx6SgSEc2LdUbkSJdzAVYUEke7p07yowe5EoX5Dh0
MxXv8mlIaHvKz+JVmXrgwHzOtVoP9DdqkdjzMeJIl7/PHwdS4tYyvdvzgBHCW79K
qPEzkH5MDCJx5eiyCtUoJhxhPcL4rCCy/NF/xMDm2bad4nNWhYn/eU6xM3sPGkup
R94aNdZi0Ye/sQLONce1ilIRQAADWQMWAklOJjiSgGbOpPzgunIqYwKDzib0Q9ra
hOYute+fkRxJ2IFZxGEaDrAwNlDD2LPWcv91nNdcV6m97WEnKSMiqwVfgRz6x01f
jQzio9CZb5wKeZac//QEZiIkcXPGqZGOtD4cWki66TomoUsCkkzpFtyW8zMNt9SH
tGOXx2Y4iVopY8iQJgWg7GKcannkyHTFUezrIubmkjOA6igPmH88Wt+eJfeB+UqA
fXgiQb6it+u+uVJCoeTwUEw+mrL5UVv2kV18Jm1k1Vh/odg9EdjI0HINX4bIsLng
6Lava5SCjRJoFDjT5DW6x6NVt/hENQp/olVIlTi4Kz/fCZzoKTL6xCMs3IDx9dyF
6YW2XNt+8La3W9+6wdCkPjQkadKA90f3dAccnKhJVqu5McBSoB6GoTbb+lw+9js1
KFg8gM+noUArb72w/iov3CSZL70TWEvNMzm2dr215EOfHYdaRnPCgOS6+Uav+LRu
VY65ByBqKAjk0Ix+3CP6igiZ89S+v3dqLUwqIj6SeMKAOPdr4gfkjrADxNWPVbI/
/Tvs05JKmQnMip+xLg78KRWI5c+jSirMO0oS+fvwZg2YapWRODXoTI4wFTS7i2GE
aGsEJmXEqfBdaUuiJMIubSrnC4PpXh2igbaTJDAOl61AJhaCkgamwp5xjPcRxe5p
PVspoUoOUk7v6pqOMwmnca/OVlX8NEGVoOvCrFuEDYjb+qzn2WgyfKg5/qAs2HzF
5QT2eMMgWTnb4PfE3AMZ1YSG2LFuTchyvWKtK758BD8Ztgi2SyIBZUiFp5JVPetC
mRHJQVQKJJWCY2sWVD/rOA6bq4SRjUeEAcnTa7+L21gcXg0Sf79QTwyFCB01/fir
AaPiXMft/4Mwfth1CAm5lpPvS8kN5ooYAOMF3DqEspygYKADznE8w65l87F2KYx4
xAOtsvziF7l73A45twkkv6YCrWjSNl90Jpr0eCXnbLfaOHAhgbRl1OWt76oppHp0
rEU1IvCkObbwPRcmidxexjVzDy0HV2Z3JrPmAEkRsR7mRvX/dxdBs7224TCdCu4m
kSR/gAbn61sAtfzrJjcg28fkxhgUwJpUhIn/GpwrJ84sQejVHOPo8yx2vQ+KHW5d
JKPUu3XYRx/dsnVEONU0BugpevUaat8ItNEmxWFZDEJsTfbqAivzgGEW676KTk0O
CEMhL8Givaul++i3fi2FLE3PL7ySLm9W9FAiNg1V6o3zP7tQ9uzWbakBAHMbIwx/
eJuHX7Wb0s0muPcD0NfpWr1U6Ud3esJ3YRmQomYtrO2FzpTEeHXw7kvHhU287wZE
uIk3Tpe9RTlwQHdpQ244SuSUrzsJAMjS6J+hCHQMZOmUz7Y4cKDgoW8udVKjrokL
4ameHQ6+mQCjtbZLtNfKpBi09M29v3XJConxrw4tD/iWZLCqqJ4F5Q7xDmcnXNuU
hs+k8hSiZcmBdCJdaB+1bd2S9nxOyKHgQ2aNWma0jxUJGiWYNShxtyNn0iIXXMXM
6s69BNp1iPvPHj5H+dCDJdpdrAy/+iwsug+aeekDJAkhgK69bmti8FuulhZ2WoEh
ZM1ZYzI3ojc+cq0cyU48ycjgVgSWTXGCAYOvu+YsvEfQPO75uLkvNvQ+Ui9JlHyw
lqKV4LiwKujYlbENOmUzO3y2M4fVuwFxeB2//mdYMpCblotvhsnwFr/+PfQ0agCa
Gjaw9mtstyd5JrOpSjUst05TpURRNHnT39f0/+DbcjCOIzfadsCdWFEYoyVfX4Ku
hMsSMcAAWuaJWx4akZpzWbI0SXGAzwQrpQArX1n6mE6sKoVc81+EPwJBC00uYFFp
7GbbjDhE6OoTFbLMzHNvigrAKY9OIEy0eiQB9yvs4+PY3b9Adds/qfDvb4BY+LRd
Q++xtqI0NO9uq6jY5Q7vd3QnjX9hALeYUisjdGxNSEQOEtgtkMcatIEj47iFW8Sd
eDIKm8OQV8gxMlXQrMSQvTp2+NtIdDA+Za0feVNNn92oOvEvrKrV2zBhC6gZKmCd
d3BOMfBBH4XqGRj1/aBviC2gl++5Stk6rtrlS1EPDFR96W4vSCLFLmZPT8YL3aeJ
5O/hxu+vVFyio+8D31hIB9MII/vLI1tKPfXMsbFgZmNKH4wnlmlsgmB653cocyay
gkWFFz8tXEfDYKmp0JnUpgcQaVPaZBa3pQTG2nNHdgeub2zr5EBjAShA3yhf0kro
XoEgpmsLxnNn1SIFPoNTy77vqT5TkBGTThhrKrFG5sEdxN9wM8prHPkeuV2CjRIO
MeYQbGZpaN1LEkqOmTRU1+I2CcQ1eYDQwORB14RbKeaDWU8HTX452BWjRbFwU74O
9ssU/uFMKKbNdrzdT/S2BNh25/j1SWKEKX2p4hreR+TbTRu2mr8Z6jnHio/8eZXm
jlSp12/zLWMPPx5YsBaOUOvJndhe4YNf65VVT3AsqzR2fD5oFxM/LCc0IizQdfEu
tQsfm7JuB5TZ7p6VsmJgYwp8Azo8m17y5+K3ibHb2KywzQUYLocseZKqJ7yy0S5D
MyI42gzam6/jhY6oU2P4oezyQCRtN0OBhMFZpnhm7x/aQoRPVfv1tMsjgU8XUwYT
8xSj5H/5tQo6fsvjnhaBOwMKv8cvACRtMvwDb48AymeQ+WqIdiTrU7lCdW1ol8Wl
af3P5XtoAAsT2kL2zb4vjmbfBNZh5YT4KQU5OM+i0FthPe4J19UbUYgS7eaYn4/R
IX0gBpkphdvo1ClELnw1c6mPCjCeTpAjLcxBJSI50/E3jL+zeT+awScJbVeifk+c
+F0hL6PU7PpNL0AsyHcIwHykceJL3c+ifpD0RYggvuN73R8EWoNczqjI3B8ytEGW
uDiEWpIGFxvhqnSSzN7IrRqwCFoHd2P+Wrlh62aY3Ew2/mkND36HEedG1U6R3aA4
EZosULr5h4XQD2chT8m22MM16Lsm7Wg4JZB6rsFey8DLyFQjRjUiCC37mTcOL/Qj
sV7+wX3tL+8F0n1xP2ZulL2UTYrwz7EC8dV5hUVDnMJwJSIq6uR4W0qFSZ+/mI8U
UtGu+IdJkPUWc/cxu7MrJo+7sSCfyDTEWIJ9elHaoW7G6hxbYzooaiAyFbXHXTnF
1kX6NWlDh+nOvy9gjWL/5SAbrVaOnQnUQFrwXk3mrRO4gknL6SNYfNRXotOLLh5b
Q1YYZSo8Si/+9AXwPzArEY0k06MX/DW3AlpVhy/nCJrpAsCIWKA5xbQOgLVhgg6E
+HxfLGsZmOXuABhr/HUQVMO1DuT98c47wjeAoQDShV5AZw7sI2/8xt+gntf76rep
77dGWAATOC/bJtGt2s7jCMjWRNM22mwkrsODSRsQojEPiQQHLa5KkOblV5/+VxM2
JvvYcXkyH4FXYtvmPU7zC2T3dEYFglIJuCPWTsGAzqEihQepd8iIeMALs/16MjXY
7YR/76nIDKdLMTIWsPbM0c4mMKdIIH9S42VPqjSltxsTISGOxL4MB0h5MfWaEP3p
wcErrvU1Rn8hpSJcPk9Mk+fnIzEP+gUF0EwnaAf6y5jxQhNUS8u1k3t2NP6U9r0W
d1Hp3MRqQA8zqLsQPvNzMfRZARgGMzT4SfAkai2TzlXngUhfmp0wuQN1Wm+VbtL3
WocFAxJT/mHqbqYoyl0HE5eXq+8JVo3JyYFpP1A40VPtPKpi8Yfbw1BMlu1LRaXq
xAWay/zj6B5CIIrispo46F+FxdbQ4rTpJvS5KBuE8lQCQqCxgvLXn1ahvwQjPRL8
hZ9xT/CZYjO3vDp/yeSufBcT8BcfdpCwPz8dswO4AiX+3fGNd7S6SVB/6MvA3yEW
nja+FQHnZNHHuOVHzHd0uLvIGZxPGstncBcaOaEDapZQ7BqMZTc6PW2Sv8mphR32
iPSf+4YHjCWMc/RkOFuF/YUzJbaHUSa8YFhbbQp6hRpmbFIIZmdTa6mJZPYdTQFv
FcD2uHC3sNbooBOZCxT4TNwoLonCaXUqTMQMwGtKbHDu5wbBxmkZT0L3pOxoFdg2
ptVN/gpKeBV+bM2e4VDf7SQGrZ5bSo90BqVoV5wM2TkT7SVRToN4WhN76QzFequb
mjquoE1awF/rJWe6kyjzxw5AqmAH6wHC2inilP0sojX5xTdByDjZQZNs2+w5sqjJ
wdSrFTxfgJqWc9iFT/S4tCIXBa9QvAcEwyFLC7egDt7i8QTqWK0jLI73vK/NOhEK
vfMfXHitbnqM7zsI19q9BHfjgJcalsJ1Nlvn5wBhyxk29MfEXmM4sR2x9nVt8Md3
VWHJnDqEm86Z07wEivkWo/lcDxnoF666PWa6Z5cXgUOh8bucJo7w6Uk4N0+LFy3q
YbyZOrzRyyud3oG+5EDubgYZKxpx1el6NWSnn4FZYMOuiwkX++Mht6E0W9UoGZaO
zPu/fMrS+79fZTCAk8dC2iS7H1rAfdkOMCrR7VKjZn89+TFwNG1IPlZ/LwOXV4F5
GNI1CkyqTdLl4u4i12PYwNDq+BQTdXsCZlNU8UMGQMoawd+DxOC9ztwuw/ustfeY
5F4uKttU4kOgQx1NquxRAck1MpnLQBQhLeSX5ELTZMufPPJDk0zr6L2GL2It+fH6
0aFP2UjzTiZ4UeM7GuH48xKsaHAa8/XyppflM/+dPoqpxPKmmTc7B6ArZWkREdP4
Mtffr7cMKYnt973ehBbp0yQl9UUNvCB8w2iKFafRW/IA4ELQK+f6RO1ucML0Zt/Y
MKDlGwPRsLfPTSUMjyi87GuOLN48gq8h4f/nYQEVOcHV3gLYrMv7gjtUYveaFbn3
IwS2vqwvCDvh9akk10FHfOqS0h3n2M3Rr4ZHVJAGqTB58rEk4vn7WE4+YBTqK2fJ
B3jtqt6AaWr3JOEHN82hv3YtiwWhykrf7gssm38QpP4q3T2h2W+y8RnIVsZdI2Zo
7Jme4GgdAnOZllgq7ss50lFllIes2hpN13Q03HlR9eWgohNGEU7fRqyVZon0c9cK
117zaUDnRcsZp1b3oOgCwSB7LSgGD0CrZEqj2Gn6lwrG70lfSwN9jwfsKU0L0jVs
TAYilxcRb6eFrScYWOYCIB/kthyyBImZLnR0ax7kwseRImKLjqZMIIh2dqbQqTOo
4vSQ8oKgG+MULccvt4SsQ3cfwcK7sOnxUhLNkR06XJnXe1xTwM7PuHVKOhEyhXsW
qRvrxnBCy5Ayb+JW3iNO1/8sBBnn4BbwYmQDsoOm66uEZAkcT1sRilmoOm8TO0SH
CM+R4lEnPzWS2+Id6lJkv9CKzz5m6IxNugBnOVdcLIlFE11v6NLqDuUFkE1vD+Qc
DoMzswlFxv2g/n5dCglA9czAKULD4VK/hZpzLDbtP4FLPy0iudfrv99gj8OHQoZ9
B1g/9lWdDUjqt42iE87SdrWLqKekCq4sew7/5ImVcHKH9sepTivqt6qdTuYD9JxJ
PE2THfJSLceQi5qynN98p9iCFLYc7zlQKFefFXExDRGfAc8vAL+kE3xyT8lD1BfQ
V71Ew6Wv6SW0axDYwWw9vKs4LoU48jFkq7fr/c/GzW8hv1BY4IvTf3op/T/27bnf
RUSGqOqwkStLyl60YH2bAhzSUwkxSo3tiD66nm9fOZB9fsve/7a9TLsNVNKklTrY
Z2npqYbl5TuZNZnMHMIYpuBfBFNUhFy/5UFFBAo32dHZ7PJe1dXcx57PICeoEaZP
z0mv3x5EJBNy3Km89zotG1fGEEcs3mHuyDYCYJrAKOgWLH7MAjlYSnLogtfjWuhO
ufPmBhefiF2mkq3KnKlai9RtLBXutzZmueeKUgeSy9lEoH0Ry9m1ohXQbqZfS79k
lcXrMxDvuPJkK5CbH943YsWMPubuoqec8GBQQgKzVVlhcOf29vO0I3v0sOaZCWU9
jiBWGmSu2eKdIop8NDOn0JKsnxfo0GD5RnZbK5w7g7Fa7fgcsQJiU280h2e8jFzN
XyxVUTwzKo51eJ7KPKGhJjIghx60eoRdq0atr+zXWYRFVFpzjVLs1hk7/NXaFXZR
NC+VBbRDAKnXTNA5CkW/f53TBUQHH9ZbAKEnow0EsJfZLn432hjRiRjDiOUZryy2
AuoUnX3ibxErH3IKZySuoI2XK0x+AFsLOMEdJKjQITgO1RRivTriYX8jmXPyOOQR
6h45suF4TQ8jAGBmbJthXBBnhtPD51UNEbkn78iDHD6uBHbka3tXFAA2m5t0VG+5
NBGgABkMb3By0VHc9To7qhe33SPywBdntBsRIZUAw+z2hQrnEJU+NN+ouN10cmB4
zOy7/YFZe4KOnu9EdF1bxq5+X3KhI7HhVSEl24pUACNUoLwSRw6H/zhEzg1BA9SJ
wFAPk0I5h5JO7eDT2JYRvtZC5+3j/d5C62oRAo3pwIsuPLci+EtFhlHuechOmCu7
ROAgkLAec60HNjespNpyWlIL55MxUuCXVxC6OyEGikGa+tyLoezPYevu8D2geL5Z
iII7KcFVChJUf2aDxRf9FWtKMkXpsPZfMf8Buk00rT3AwYtai7FAypwGbRSLVGA4
tLEVilDlWS9CsITcbUNlfoZ5y6EMsgsVpfKkWcKAeLhT8VCvgwvv5s9ZqKQ7BOjV
rVchZH51l9IhUIwPtiU0SgmEn72sPFEyNRnmtGGG/d6VJA+j0T0gxR+YHl4J0XfL
MeNmDoXFqp/uUek/zF5OaSu/ULvyjEve5nPwBbPOk18EBBU3d/kfadZ+ZsGoxW2L
Z/oy+nk1ZFiu1eXkpXGHuBfsrxbt8/bxhuJbMnEn5wHwBJS5EQ/tp2rrzjubu+nx
MA2Um087/cbZEocD/SlCwF3PHHTbO8t5yt+FvOic9nf/8W6nEAm9twS8KYj+AvU8
g4zj8kdGs/Cmndk+iXCpU++bRPr7y+b1RCqhyO3dzlcwpgttV0JrrwVczYXiholb
Fx5fkQbHyVZ/TFMomLPdmJvuLDZb2jYwinZsftTvglN9Wf6cfhrPb2YpVjr+ag9u
Xk04z+woMEX3MHLf0lj0B2V8GbMKh6PUfSHNynxNv1X0vYS03NncPA68yXlJ55Jb
O1fSZnkLL9fvx46m91Wj7yP1nymqmUYNU1+B7EvPg0yF1IHrizDH/JUxIy8gHNuW
xC9uK38g+JFyor6Amb3D592cO42sdZt3zQ/GTf/bjKIl9eWDwQXDiKgV5ShQiYKk
RmkR5SEJTCKRFl8erCZNimNXegWlrcbHKlcXd+v/amh8Isrwr0/3ESja/ErgrPaA
Q69RrLHY4uFJCg8kl47CHG+ASoerF/b828WvcTro2rMsBUuSgG9z7g1nP7yTgvCG
PnZkRL5RbwJu0xRWLLw6Y1XasyP9pNOPmSQFMK3r0d4LXrvkEZFILL4xxJ5CQySW
VX9qzSTxGKsZAewaZLWqsWTmYx4rXIwtpF9/b4ffOG/5Le12cdRqNj1qXem/QoNN
0bvngbNR+lpl8PceOsIPUnpO4U7WhK4mNLB/IHJheYgHuBJ7sadl2ARU4fDEeARQ
xU9Xm5lTIpOqTA8n1wViZHfLrJmAxy6nqMeWOGzosbx3r7JeXdsOwi0lsOpQtUdD
a+J3BkPPO9AR+s7GqF0FurPcXIUi/cm5Iqlg3Vx6G2momN5It9AvJMIxmJJuo7Vl
BpZnNp03bedKPC9pnJ5NqhZEcHF8uf235zHm9IPRLZMrSZdZgmHZD0uxdBIuX/Ca
8LAfAPZIZ3V4EZZpgxguYmEUfYcgE4H7kuIvwI2jUC+bbBM+uPlrEm7Fcur+ED2H
4t9mmL5REx3sfiMtW6flAbYiB5lgu6i1OHgserlZ35rvfJ7BlkdjG14N3+AMQJ+f
gDpamT+ix9Gw4/GoH5C3KWJaAFATJZbWgZ7HHS3fLO26xGBQnYl+U/qODJqfaxEG
t7xdG6CP4ImWmmyMc7Ny0IBFsFVS+1REVP0DBkFRIMigpJNlpFRYScw4D2bwrpjG
xJo0mcoeljyC45NUcUJWyuiMlOfF4hObCZQS6g/y0oDr+Mesx/2QxMFoNg149K0/
heNlkKF9g95CpuORKJefIoyExz/0GY76XZeQs7NY1S27onxZkUBVPQo369KrgajV
Qn5+f0O2o5ZsPe+XIczzzochgFg+cEFzw2l9GDuGQb/0MyGMXB0J2uxq0JmH2tg8
b4JPBKnsP+AxwpyKovysboIW0wnPQHCyym7opkc8QQ6QGeTOZuTLnX9WajBYPFiL
qRzG3kQ8NsGomY8R/8qEZrYrplajcMIcbn0fcRNMQz6j9xbfSkHdsBAKZ3QNBg3B
uJp+obQKW3PYdNXtugk9suLFab3h1jRhly1FAmOOmAb3k66o0EheNlIsLk3lkSJu
MmHrCrX4xfaIyoq6CqlHBu9Wg/0wz88aK9tY04nBZvb+anuBpNPpt3+Q5XhsdTgx
PGJKRTY1vocEPPu6z9vHbGbwCfBuLg145fdMMuUpLlU+swOSv6VzvxVzn+BPW66q
Vvwb9RsmK6DBZVvcE2VyyJaI8LmUfzlOVBUObmHPT6LzeGv8JoBZNVkjE/KkbS5j
te+I5Vn1Uo9efXaWb8yF9O/R/IKa5lQ6BCv93ZQYFTsqMPAuDxC/gHPspVyM5s60
qF1wsjkssdCfJafXzk7DbcmTGA3tqed+LvQgAAsoD+0eYgH13omyAAMFL1q1Uq/u
chQn2ErLs6Q7mMpWayTTnNNP3TwS31orTrGxarhXZ17PC59AhkHuuiEdnIjL3ixY
e2iruCfutqXVCqOTZzsP3BTALY+wXYo9KhB+V7ORHiNV9Qr32au4imtoT1yvjonI
O54EZgNRea7aWTdqahqwPb6r1ejGxfh1a1P8XPJYjiWwTy2xJ8z6HP1wLHe1c3CY
eDbT6mqo5NTfEgw40X3sQIkLBYvb0LepFAppR4ovRbj+fHzn/LTyhEw2+H1KlMzl
PUwKLtyOB23mqii5S28hCee5rwVnBsY9QdvwThG6HWLFN5gc2zqvJNNwD/skiRJh
WY3k3P0JUAsDMtZnKKxUKkMNiljr5B5LyZby/Tdqn+hWf5k2YjjIanbLSlFUqfAu
Psax8r7eI7n9U7iXCfi/7DO1etNsF//xak/86Wbuwz3M0sVZ9054kFmE1OuhUdEB
kQs1DNYUkUALiEXtIXUR2YArgy6DwQ2tHBxSUO8+rXUNv9Xn+vA4bNt8hOEWkZmM
FenB1g19Ot2zNjQlNm+Q95aKa/wOBWNbwiY1jmZ5g1u6oKgLmzfnsnS/Sp+V30mP
x67NrzhWhCC5F22fHv+rZUpLlzG4cVIdaHEMxH2EN3IMBhwjaeJetCtpsL9DEIRd
sHL3iYnUSGScvWX76iEHOZd2vjAC91bsfDqaw3k1jwOd+DrtAm3qvgj7LcDqw22Q
0Iivl445tD65NFKxMpUJTD0ft2KF2Az2Krn4RqJsej3pj9TdQSMNRUFTRxjRvw/V
GruPxPZGRXlZkpmTGtp4jodlkQxKKrZO0PLp5MXD0bnHDIRnf4O2CA2Id36Ds8oB
VlVDSIos3jJ/A5+rIDHcAkBuKtaP5RxTjh6+7IQllWhwKWCGPrX7RB5oBCTGpeIy
JNQ2T4h93TP9vyT7fOzvSBX5Qbf4rF0A6iyZmdWz9XadpnJd+0ee8a/CnD5F5Zce
RZVe57aRMqHf0bjmhb135hGR1+cPdZ4E59Leewurgp3ZDX787GsrgmvvZSo/pD2Y
6WruWmEM7R/x/gDYL8nxxAQYCCD3GACF1xKiOZoohDONxxsM6K5+ymQIxc6M/nyU
e3ds31Mg0t4dS7GwT4K+BkUm/uTRj4PG34uZi8BKoanX5qdSejy/DlK3EzIQIkeA
N3aixAs0+J8SN+AgxPdnYZtOHltVGxLz6umni2XJAozVE7an8od0f8AhDn7oHkID
r3p4YBRVCWEFzhpgM6Qrmhua+c9Ica7OhMQTA7frVCWxfL78LvFjAxZoOFmaDw5k
wZt7p0fkrMVklJcWd2WXneg+zWle9arGmLqTy07y+IAnm8qHCr4Zs0sQI9y0SvxK
BP5Dsc0a90ziGv9h6zJcn/sP+mBwWORsN3NJ1XhpDYyLGdup//S0i7RfDrYd77qL
SXY3cPonSyPNiwhz8QXb8mApwN8mOlWCi2FBOlAr6FZw8HQl0ktxn23HXlN/gUCu
RiFPUdtCAsfWgTjkCnP7083XShJ1w9ml7aQiC8adardoNjzA+MpOvMtiP6rh3QmK
U29j6fMGBfdVzWmzeVN0/BxnJmZEpZgLta9dz8PdIVg6sQKaF6GvGIw/TLEr21b5
nkkgLpmlFoPpgCF/l+rZn7+JbBaVC/ncPLX8ffgFNA/i3nJHIzp0XLxDIBRhIr5T
tiR2eWQjaBODd3C2e48KjZSYm8gy/Ui2oBs4mQjJ/h7pimSm4zVLsqPYZjW7SBvl
kCkO38DTUK43H8BAOSz5csRi3fO3bAvkwSsOxGjlwKsTW947WSDMFY/nybOuS8E8
dhA2yOv52zTFLsbacPmXlocCUcTOfuI1QHBLMOLorUzABBzFahXNnrkdbt/mHmdW
ovIjDzJNuc30BTnQKNOWbojPfK69w1XJnolND9lDFBDY+SHOcKX+TzNOElIxPuii
/4/r47QQ70tegAk5Ab7k4FdO/V/g/Oci82EAauFURviLRHQLuDOS8sZEhvOgM+sT
HP8S6Jt9BzQEuGYIgiWkqCLi2gf6NFfdRfdAoMQNlaCB3XzxEK9K7nPOI9jpqspk
c63wvSK3+G77keNLHPkRFLK1Lhe6kJDhLZx86Juv7boMkbOUq3ZCrb5f/35OnoVY
46I3TiwBWoc8U67vk2wAQIIo/jutyT0DLwt/CoU7Mqw/SFUh+USXX5CnZuuQShDC
6fqxLDAAsSf4neOlJbMPkXXzudIjmwW10NmXLSQWNMCmln1HULGrvXSBls2m+O8I
b7Ctox07SyNxJ0QxaRqiPsveY2D2eYX6thiFtFsqWzodwMKZkUgA5Sq2fz+sZH2K
DAi3lxNC5avqjwwGYLazPcZQr01xwBPlRzJEGoJruF+11skGdC6SDbQybn0yLug2
kmxLX96pGhBcj275KFaY2m+siT58D34X4BR8Q4KCLY4egcPC0OMieaVPkLSsulIb
4+BsXudZCVhbrS/Das+wuPvjlHnAaNV3ZVe2suoDWI6ouNp8A245J3L1C6VWQFEq
o68tFuhw0jMSSev5JeGCe208stpiU3NRiJhOF5OsNGi52oCCqo9LAxbuNabAq5Bz
0aAzllQEERg0MHUqBTq8l4t24mS14I5VnY0f8qb3CJGmCaaiovXFOmJ+JGgtkf2Z
NOTl/SCePrH6S0DAz/+NFMdl5r2VfqTS7jRK+GENdjsHvA0lrtrBbNNBUIwPbCSe
0NhoN+U6Vok/4ywEamnC0JlDyp2RC78ziaq2tduDISKnHVGgARf+Ku7cU2LP1OEy
/bONx9Nfe5gL8+bD2Hiy0qt9pf6Abbi1uc+JCMq1pvLno3VruGM0mzksbHUtH42P
1ss3+ySOE9IBGyYoTA//tjpzVauoBW7/VzImjz7ZF4uexz02ZexhYGqTF75k1kPM
h1VMCTmlnJvxi6n5UMx5rFb6iNXi7Z9zpz/9AGsvkHBMSiA3bClre0HpDqWnvl1T
COe2VxrRIOwHJStYpeEPHG8DMBpgYqTc21EuPUWozvg7f+UfA+gnW2/Pd0a7V7sZ
9gFKT9fOJmzJd/LX3Je2spmndSco03kttR+PUBdhwnBbubYwB55iXb/8i0d4RJ7p
0VMAu+HsZaI3UduMPk8SlZE26bqpiSCOwtByok4sgXrLCeyemG8/ePFujvgbpMKH
BamkOx6sXYUU1pdN+ndGPogxKl4nx3A48OwdIW9apHrWofrtJDJohwFv2OSknm9c
wL9Lz4rIro/hn2B8ci8sCPQ9Txx8RjDnzfhRDltLibBvKXbgYF++eoKKnVdI9M3K
uYbOdEF8s9imhpyzbCdJHJ/8yAok0uC4RBnHtI5gCWZxRVzqzyqIU0WuBUKPD3uE
vphEep2RVAJCait6fcqIxYYdUJm3MtPlSosgkQWmiWL8sNeu9nxRPeca3L9vKFJs
oxFevx18nfbX0M/yyECb/PGhyFGXCFW1b1joiLQM9L2JTBz2VqR6AeeDRuSaLEOS
fe65XGLAM6XSLdBpQ6pqUlBPKOTxtg/kcTfaiv5TbYuTJRm8wQVuOKdzZikrBVFz
vrZL1M2i4cADdgHQj8KLrQpNx0m0sB/PbI2VyNlgPlZKNoeEfvzrVrRoYxobv38J
oqj7yhf3YQ8+NwJGsyJcX4IPu7qe+sb/xOfvVumYidEzI5YMzTwyhpWO5YsPwIm3
/MPFYZRTl5hgnwJOY0WYG/QeTFilyfil34FrHzdNDXxnBDaS4+IXE8YC9P9jQP93
2uCUOVAooHKDBAaDvR07K4nCxmfSAYAQU4U70FMtYGFXNCUjunlMoRSoTIpcO5QM
Rra+w3r6SsL4gFPo/ec4m45sUCgxppu8+d016fx6UFkCyPy82gazc/4H5CAtDXH1
9OjKMXBuO8cngqKOtuqkdveDKeTIou88cTaLMqZf3yMWQyLNosYffqYSTRJUJtlV
h2TE6Rde2kBy9QSDXpKQnue/n+a3UR2NYq7/S3VCV53a7iskc6uU5b3+fGeoLwEG
l65F0as8zgE9K3/5f80ab9n5MbfPxE7mdrLp1wPD0rb4PcoGUnisSmrC+zTGmuAG
8bXdTo25d+gUprosA6r6AD9SvkZ3yjGMatH4/ryuqJKZDbJolF5l5pSE22Cb3oHz
Tv9UXmw6MgjLuYCTLuJml0BtottIPPswmydDNknhwblgfIl6NTxjJFPs8umgcXd8
dY11gNX/tXY8aWZDiINiw+2IWq8eHdtcguYl6DepWlyByL490tbBxNy/Yuhwt8GA
NW65aB2o9zYtgl/Dizw3EdpCLrlAFlSmOFGMVyJiwiE3qpdw2Zlr2Y0TBXe0fF9I
yhEXdxADjmP5dSzX1OtM22C+4iwqPxkqnqrhj84BDMU7T4Jby79wh/jfBeOXVF6r
i87zueYFjSXJYnUBMr07aWS7DPO69QONkzDAvHd0Bp9odGqzKHxz1Uogy2ozw6vR
ZTIkwmoBbH+wn4++gHBMv1Cang1jmPgmi3yYSTi9H+NWpUyfNOF62vWcDVMX47G2
uChb36cf9Xr0ecNIV4ELCFnHqZYEi3UYTEXySyvHWoL3waAFS084lmrLtrs4PvrD
+M+WcCvNjVkavg63J8sg+9ODM/4KMbF15Qp/rComC4ToUT7mlJvu7dTeougT58+D
L/pCnU/i4DTCoFKMF61ZWUh88QUW3lpZEHYc95WybaZ9KHB8jQ6qwCZWREb0YwmJ
7p3zQB6eSfUWHVLeb9cuuF5U54gGOMac1KO8I4kttffpSMqXHg8kVOQpNCgqhZbL
+11n7zNp0zhU+fjQrxYrqt08Ygt2zvh4vCtSiILYQBNckkYxX2KdG3NmiuFaCDQP
a8hiWvS7Lj/CpvxYKhrOvtV+NI1vqjjbfuvSXaYuC49Sz1tTu6DxhIXxIA1G30t6
hlq4QNOtOrMOICcGAs3YdaPIuJpzNAk97PrIlZv8WvZw55FclH7YR+F6b9LnyRih
SBlx2RAxsl/c3jlO8/7CuaAfP5ca26Tf5Bz/HAlyORaJCPtuxbfP8gpjsXX2DCKh
URKUsNB5w8EQ4b3f48cvKX6l+YnMtn4a8wXEh8kAF+yyj5Vm0hyqD/Gx3RSjM8nU
ekm8h2ct93yl/tfDFuB5vpts/mBY2Ktak7mC9I6WE620ziVeMb0+P32khV/UzYUT
XudidArrWbYoGXLNk3V/j3v6LHhsme4QN5jFBJclFS+/cBeZC0MqApB0fAlEnD0V
axKuTOytSMGKehJiDzmHxzTrWgagOJgPoIavljv5fVaRx6SZKILBwONiOkGGJ6KO
gEaPhn90FCE59FPGO50Fo7S4qXbaPOB9S4ZG0s1cz0fskNKnTIqFDUf+qhAk8tvX
CoeXwZOebOwa3cS7wEtS4Do/va14cE/dDKBB5nMoViU1t7FGBbVE70gZJ6GV7eD7
koFqOZBwpAnf1kBebuFHwiy2YwAydwzS+390wBjxQluLVjHj/evFmdpMYxFwHyHs
97ntmSAfZR+VBVbl4veZfOTsUFjKoa/VjIWdhbC22orsUJNE3mK1JT8xomL8o+CR
hM0RmZuT1oMY2P811fDAxflJPJBBEdSm/lXNoGS93q6/u2CMBLL+fFja7H7qGhIh
auzVJ5QbEqsb8MyKes3agzikhdEJSXzjHYOTqD0Gj5I/f9IZ0N4ptFXK0bbt5nS2
Z6swNmpzT1WAlvpfq1LF/k19h/bGFP4DB/9ttC3DA8gcb/JtJoo1cIwbV4/ohaHf
/l5bfZlnfn9fJS9q6eWKGs/5M221i/8bERx3LFAcDsZc0xAfn9L9vRotewymeAcW
MoVKj9eqgyIXyaxIAtDUfQd6uA9O6IR54LLTCb1yNPwTFTkAucEhOsm78XHXTdHO
E3GQjSQgqfhTYJ8vCcRArRRXkW9v57EWJUX+TFCB56/fbeaXz7I5zcElGeRhFjoG
rXmiAbpBzIDGPkkI227t3a7mjqEzzNF2UySdndxKHqLeuVkyPdo6UgfSrqwQZ/Za
OQQF783QARRV6pe43Jn9PIpwaiUFsowUIYX5sFuuDxQ5kv2EYPdpM0ZdWBUM8mGL
UVbIr9NU3sWzdy6AmttGftcaP6VTM72cy+tYzVoAeoSAKS/AJfr3gA1bUbpG81M7
0NarEWjmeBw8eydvBR8YOVk3ENWA53h/+qw/cjKh+SVrb89P+cRu23igdhIeRP+v
wXCtX11K8yV0+Ggt67xcDswIp/NtpSPosnxwtbW2la80mGC3GPFq5EjpztWRMr0N
uApJzcSMFJYILOOQPsTrFA9nPMd4Hgas/yC3sdSyVlMLgL/uQc1dm1XW4DhVBcis
m7gCMQ+5s7RvlZkDqi3VoDqb5rUODn/jpFnyZdVcHcIDYSbyLBC8BeU79H7qKZ5U
UdpHVnyBMN0F+E1RHp1keAWkwAabKen+fe7Q0wlzuInQCUPToyFaX66hVZh7m+Et
hGXuznGQKXFb/IRBLLno3yc6mlReNjZuql+xc3re2TW0PgTZ+EGRDTky3aCA2AOO
l6uBZF72gvkuQZ1Vw5Xem4CMTIYP0rODB+GefRALuPVOHylO4z7eLiSgYTgzXMYR
6hubx/bGbSE0RzS264DpD7p0FVCnJKSpVkOHCWXJLffVv3uVgMxj7ApyshZF1Cxm
eqbjBsZO/vTAgFZ29vKcDmAtc5aXm5quujDdQzzKyKBM+f34pD6agP9vDKr7yw7L
MKgMWvEqnJu67jQj5T1my79VOQlVnQtNaQJST4ru7BykXAf9U3vuwZUe1quws2h0
YRsPtv0mYbF0+lS/qU2Crhoyux0eOZjU0YVBh8vHuowFlvFxgxGdlFcJr5116il/
tmWFJo+Y5FF3g5QXQu7UsgRWXqOfDpfviEUCVqK4r7ZIcbqL9l/zWcdGWCSgYBW1
EFZOTAFy3ypu8czzoPqMblf/EL7gAQeTkAARTXI43oApsE8heZBmCmTRUYiRWgev
8J85ko+Fc3cRF68C9BoxVCKfBqALeqldAoV7bsuq0mPG4lznQeXCXfyVgEXFb5nE
MIWDVr1dvA+mwuW8/7fjoOZ7K1mQvAP+VckC+34+k2RLX6MZsUAB6NxjPK+7VNTh
STGMBzzKFVQbbbiqwCNe1IlXQneRswv/7gZhrVR7a8/qxPMSQ5YWzE80oLP8kp7s
5bIKVWwziw9aZaOBwR12MYefqGMWs6fOKqP1kOxXJvAUVnT+8+7jvkgY3F06jhjl
nfBQ0dGflpmX5WUze7PCsml1ttw7Om8E42wIr46UN09b7mLooTpdNce06bcOubBb
SbzH1sjbOSvMbhIaFSo+HBZR0OZvqlnpiOMyeZKZLiRsHOg8gk4BZUdyLMePoSWJ
fK5QskJFSEx5CoM5j59A2twiPPnTcLmtH+lb4bXz24vZINRlqQl341Nz6kPtIOqw
37aqqV3+DNML6DLwv/8IySnPHEQNuuL18TmPcQHeWPgZCnSop+dls+PONDe1ngM4
zSXRfQhV0aKnMFPqEHcGQfAW6bbx3XjKeAIOibhS1tmNqriWpcXYJWjWEwgfHtlp
zVl0AyiSTGaHSYWTLOljLlPkj2h8qXSX4nDB1hcVk07cGWEU+CcfMJ7VacqBYr79
2QJMl+LiWaDjFWLpcLECkvohMi9OcHNv1cS+u5xBDTXil+Yz7b6cyeEHLEmKBdWf
L9yB4OuHl2uNrUQ+QZS3vgtGkXdpTkhQQ+CLSHa5h7/dnlTt8Yt5ItPFowq8pHbc
ttCY/RUNdURBXT0fsmpTuKRlsaZz7Qt5Ci/H8Hy2LFjo5mExRL222HUH12p/MxnA
19qsC16gL+gTP02dF3U7LJmi49kFV4FZyJxvIQ2KHY6R0g5GES07O/r2REm8lgsT
5V21UU+NjFDU9vrGoeEAfD5rr9Fxay42WVdF8FxWaCMFOAmjShoStianlwCTISpg
RIHFcL64J3/mJu69xzKPPOJRAorvZ43YnscCPvMay/ywfik4Adl5Cu7y53YdG7sD
322vig2qW0xyJG5iH33v2biOjh1fZTx+9+e9vy3XSFM1QbaHwS+9fwJR1qNi2qEs
+s3UcCTbXGUIHIc872jv5Q==
`protect END_PROTECTED
