`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bnbdXLg/5oWB5Kx4GUjP5o8oEZbNyS632lf6nPGr3EDbhmHPYY8xare+MjI3LVux
CDreNXndzOCUFF3Rlgcg/32WjrOd6Je9UZ61bWT1Sy82SUael8CVGMxgSW8L3bEC
pFtT1gCM2s8VVAbqN7W8bbPiOicL4PLMH7UT5Yf4kfH2xks450yqBSm0UM75Z+YP
JL9j0OQ9SoXVAWeHgF8Q2sFfpLYzPZ6appY+mcuzP3KcvS3iV4UaCZzo8wwJSqb4
SfVGxQnA/v5oAT2POQe6IM+4BSCCkTrpO77lLT8nNrqtCh6JNYHff9WojOfP4EGi
kl+9FNWHJ3WOPW+Ty7VHNSUpppldT0Iihe3G1RWgTT5wTqkxMT+0c8IeQeuPYW0T
sTSHdwa2FHdeTlRbDZqhW/C/fWGdF3K01crOA4En7oqjAtZa6gItDpP4bTyHRRbt
pS/Z922QWKrDU7ZrCbXN0m/acc6U4izJmP/+Dn5eEGXzbZsITk89GT8baNXG0VFf
H6BnNc03udU6CVxGP1LVxG0t+uUcztEzKYs75OMCxJla1qjMlRzilfjj5tuEF3Qw
jC1TftPlBs00dR6tHgcJHWABCqJyJOjeMZeimwzhvjmLgGlugb5QbQFMtA5aY9Yn
Qx0v0Hwm6MV/l/DWsPlG0dK9BcfnFUJOcaAxtzaAouQyvenUVLahVgjoRTR1EBE4
FOyPZ+x7ncxmhdRFTT2xLqFXcyY6G8vL+nlbv8MOltTpxbXmiuhKtjk5gz/S7jvF
Hj/dLfZ4vm/hQe4bue3rasJ8ddP56la+HfIcN+ULyrL8rtk/ZEbkRKjPDHrOu/ne
/AKfChMh6EinK+dvlCxXId1P7QoZFHZBZx99CMSV5Cybe9prAEVsPqugfsmvDJqX
4kPqFds94SIKmrCrd7Evd8A3HRApahFTZ9b3qTZqgFSFC4Eaf7L4Y0NbD+K0mRYm
TvdOxdsue8fzKqITk4DenknhNYGdm9gXeOKlqBsPgdItXF/ZKDn+8A8hkR7ivXxE
zpSCykX47oBXTwJuhkin9n6CSecflAReMQGylaWEo3vStEiSF+GyCzqxcuCQIC9K
4TxFtNZtLwNBXfmUdBvD/T5FRxPJND3TdkhzTuWxPPbRHVwOUDjyjyqDHiK1HTGO
XYpGSwVS94RcBz2N7t5O1xLKEYLjdQhjy8qtiy/hAgiOi5O0nvOHw87DzQn3pEOd
5bCYp5aFdjirQumuzsICp+btfz0EBXk1Z6Yx4H+bk5plNhygOAxjG92k0tIApdCW
5yIuk4BijMKnZSAw+C0xFsmhjW+u76/XhRjMSsOyc3wwxZ0jlwKogtMjaTylshWF
Tm1AMMcAVfhn720WhRioH2K6r98Kyv/XEoFJ4tIgctgvNncpwUSJpzT1EyI0MPBq
YzoHBY3QQTkXFWzAGAkFqA==
`protect END_PROTECTED
