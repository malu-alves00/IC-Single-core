`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Bq7kILiDlEt6pBYjRroMH0NLfQ1saKTld7RQthXuNsscQZYNR6O10iNSCfngGMbc
6kdjDVt87pLomsaH4URoLvqtMrxa3cbqBxcBHr/KytVJEmBItbt0J9dJvL+DcNgU
zZJNuG0XbuEBO81nHmFX996yrszGrnSZwll+/63wSHYggBfI8H59/xlY5xXWYXPi
6Tz1Cgk1nRiyBhrHYvVJq1iKv6ifyy3en75OWpU/Y+kBmzTNJAGhmGa2ZNfNLqf2
VX2W4iQfSbmrrfoYpk+fMuHMzmhIx7iWy0yfulcTq8RH45Q6HelmkvFJQca9XL2H
CW0xOakEik5WraBJIIzuX2H1eujUCaAMhaM0z3YPodCgFVVMkpREZ1Outm/TezQ4
1np+47WhhwY5WOqFy0iiQ0cHZ23MZIHn34TxBHljqlTy0ez3Pbrp+LHuYKJGsKwQ
omRrYXHlR27pRRkvyVbSX6Gw6jX/+h8cYbw9cF8N/3zIRlTU2TuFgrJrePXRsSSs
M83Ng1xJV3xx0lRSYo++oHiatM2d2BBcv+Bzm3kEOgs9rcWU073QG1uafNYPW/As
b/AedmBqS6eEnSrTHZnvf8gncBkgs0gaOdv4SaP+PFN9ZSGPH+Se3nQUmtSW2Ikw
q2lEfpMDLKXziSMJXrCVncIPLygTFLS/MuUtqeDbL2JuFYTnchvPHB/yKjOlCpsD
yR5CQqp29qJx8628JCXKI61XHK5ppvr7PCx6khb9pd4HHQJqSoNC60uCvyIG3a4M
lZd80SBGgl6N8+PEOlSb+4EM2ZtrCLNI2si0R86VlMZ7gzA4fiMTx0/t64tBvH2O
VPah5kIZYQ4iC3oW/ZtDd+N3qPluaICWTHZUyZAnRaNWTLR7rrVduGI9udduNwQP
0W5PphcBoRk+xSgPKsTe2tThYTP74Um8QoN9VSN2lQGeNa/UTLNTz61rmiGGNidk
3/8ZWE8Ce/ng7mUynutxX5iwXPu1WPv7gf/QArhz+4heJxyY3xDaRtvJHLBKbTmX
KVt6ripfrUUptdvT+ef39mxjj2R6QCMjAD9jaLvU/+Zwd+RsgKLjuKH6m/dJz/0r
SsflHLohFhoPKkoxBtIxhEnnZPRNgvJjhx36qyy4Z/Zd/O+6wxhXnMZo6zctjlqa
yLcbORX7iwwzT1i3lEB3admpGaSsFaN6N74BUGiFGgbcsxfUAdk83WfN4GKVm5vi
QqVNBLEiPXarr1rQhuadJUnXcwbdleOqwVuG91IG0xujt1UAF6yLytwRN+t2McWq
yY+XkmWqFEgqTAIPAvzD8en8LOFmRjkj/AFIFyJWa/TJGR6qfQNo4nY0CtFZX+8G
jH8eTYuqZF+HlUz0MmCjFCqZMaZ8unYLzrlLXNWpa96GPaG+eLgRu5iUSaanfkt6
c/+Wx+rJruiTF+PVrvMIRHfqPoxqVrx09GjWrRpUoIGHJ1Hsr4FLjasC0AyLRXOn
04hzEZA3x7hg7JkiArVAGdii6xa99kl8K4GeY1akVzr309m7SLmeVVzlz7leHFSv
g7VXSLk7JcONMirH7Oiz7tV3fjyy/U5DBuJRMo4rqkwx8rAX7zoZQBc4L6M4h58K
0e8Ry4bEbxp/OOlHZYwCe+lyfX8z+MitH/n96kQcO/ypW7SB5HNNhns28dga39Mx
/yKo608GIneRC5sVwFZnEn308PC7ZwOjWfnVG6E9b1+TaQ+yzr26SBeXOGDHGznq
Z1i6Zl211gU6nXxORZKe76JjbaTi1Ro8NhkRNz3vBeFtu/EO2QnVKTARV96V/WNI
A9dsnvw3I/IItFEK+d1DQyAnuHmeksuQf8jOy/FnylZCKdIRfxdwfRja449QWk+w
UIOnUUYN1cs6SqRqEQ0SR4kM+tQVQ4kdnwYaynwIyzjG+4IQeqwBpzUj8fgyk5qM
QTRRX/IZj0+bAQ60jlqG5UZP/DssaNeTskmnfpyl/0bji68uJyEIVNQIMJivjJ1T
mJQX+6x///OP+7Cy/ogTZAZXb+l2NKS8Nb75Dbsat3XLTEy8c7f9diUij61XjpqD
OC70tVTOi4LxTB6CvEz/yZnjM2Ysn1zxO6WI7rH2N9GJQYmHzuyBUqrOUF+KIjMd
tviaNGQphlJ1k0Htq0N+D+f2Qo07FyayLZqVEyi2pqtefQD/yBhN5bshY9uLaM82
Aa51KjsHd5AL6pJUY3guiwmOW4MJOwESOPXccTYocKhT86YbJn79KrC1TCIkX+Ts
DsYaWKal8QAHLB7bwcR//Ga1VknIywQGQdfT6uhVJOaF5pTiQoQ7xCflvOCwUN34
I/PD4pAy6rj5x6M2klzoN2Jt3KDbrSPqkt0WeN1FM5oTb68AKbTb034+CBuhF/+J
EJ0lSH+xtKfpmmlRHfSy0KG1GyDqmfWzjDh7EuwCJzyANP5mvLLx5e00mQ/gunsu
A3DxvNTl/H1/R+5zlv/GJT9q6l2cLcPxIdB5Mc7N8xL9pPNC741LKxHkimOSHMlV
jSGBPn1zokSYpKmC2qdmi2MVpEerkM4a41Fu8HKj8bCdVdp3WFv4oxY8DNLPn7pK
0G6oNXzUixujJEgOhSgIXGAscS2cuiz6Zs750mwNu7Kff2oQ1votIZ1jm6D1e9N4
QrHTOo+Dueoh+GarnopKaEDLF0mWx3T/PhYB0zXSgq56uPNkEQTQJv7Aa1srJG9i
0ImRfZqmTvos0iEQxKyj/8FGiXOmbQ72gGbSCgeDMCwgADDEogAOltvL2JlyPJSt
0fuUdhR6sYW0CTmACdK9uJEB7k/S7T3K2X5SRjInEfM/vP5o2V/9WJN7cqzqhRze
NE3cnaq/wSmVInsX7oRl37QcGQSBQsbVWnU1QXvaYlvSOetflmVNIlx1X3ONXEdi
xTTbSeDhuGbEqVea7xKP0khUsiU/l0uVKn3b+lS7vo7b6vZaYMzY1GVJKoaj+gcf
hflxiDkIEnKrBjev9bTuOHhgemt5OgzA7g9F48jlJmVe8s/yCesk4ErZXk1MufAE
62M3s7Nba7ioyPOP5FzGYYozGoIlYTcERYp0nlwe1COx37nIGxYOI3RvI3eATybA
AKy0ibBaViR+x/ZbF9fmoLN2kI+tk8r0eNt6XSTsMuW8PWhN0oY8d1yrJ1H+13sC
NlXL5YX1MoexFh8kbV+gmdJgh0wwfTEmnC0GMSwXHgVBObC8cdEj64+hFZS/mqhn
rtev8MHEfhtk/6ZpYmJYd8IAED5ijmW6qQmtzjimJDi6LVaGXaJH5UGXQNEcjv75
uMUHsX8BIT2+zi8I5CJjucCL62jzpIFW8cCmms9lh63kM7/Y31oXNWi3562bPIT+
NEKIvOjsRsnlVAwMbnLdyC/HieMgYRByCaiASTt+594TqCpDauPYXSciuWd5eo48
b/OSH3F1NGDrQgv6VITXLYZTKOdvVlu0umPnGyThgrH8HE9VRqrOl0u475unirGC
S4Zv3FsTzK6S+4F6chPVSFAlpSHM85Eb2vEHOat947kSXpcZHZPS2Y07B8vMM9cR
vmdup2IVg5IpkeZznZVQg6tloGyPhM+hkpARsof/fpLzizUagJmIbFEta9tlA8QN
x5QB4hw14ZcDlH7NPu5BaYDxfMYG0vdoI5IiAmT0XmxLlJV6gO3UrlZnqpZGPzI0
3nSjtQCG8oyAXj+Go2gPz9UaofZ2dhgOq+PBHF9BHvTHuYYGQOa+5HuO6Po3pMza
wq+hzZWLAxMi4rtFw+3MzKTcD9obUfo5Ki/sSMiQoRyl8kLQcNpmoSham8kiSbRh
5OX1lSRr9ggs1IlquOCE0XZnErA9zzGffANfjqlb2mk1qeFOK6iCEWpYZLN2eIVB
jZybleTKZw4xmmpCLU+wFi24Jkik8sCyuy808lqADwWEArnijBL9f51bd19e46xc
Umz+ZQWbIOzb41G86qExHdLrgjsLu5Bkhkxe8tnBX67qyBvz0nqcPPSDXjoYLZeV
n3agXdUCpHCYFZNFsN3cQTQ/713j/QKN5LrYZjSx7chG3UQunhxNTONBsOgints5
GwfSvCYhPBO5HunRNMmi+jyCoxfXBDG4Fq79dTZhsBZmJro/4jKrfN69Lp7iXIfI
WYoNmvhrrPTY7pXafWVACEnpSMqom9EQR0HL2CVY/6CzRoeYitDQO+fvMPEpIw+R
oypSkhWKkVCKhbJea7xGuI/5giuXsWJOy3TYTE4d64vpsA83YNWR2eTSntdBIzlw
Fe+EO9N5FsB71bTAwmbjIH73ozBndweBI8zTLQ+d6EOmwMxQvxU/D6IlW3pSzl8R
SMCfpNuQtvMdOiZSOqQ6QZzJhsC43zY9q6chdBpIz1xqnIO36vmuRaGbSPSxznI2
O26gLrzDDF1GMfC5JZai/YwEuLyW6r7CeUFe03OjUjtJl9nj7TIHXP6Cz202sbvx
v/g5fb1ULtoSS9vicnSfSm3xTvKq9hcIystDp+jUhc3Nb7ElpL9en0cLUNZ3LFlV
1TZVQoyxtSfkxRQ6OcmMHc8u29EWdtACj58pcH95gwKQG5JG/sDANfFD6ETsD7q0
Z5XHkPIf8y+JP2KSxpJoT3cPDunnSC4opnbIm0YOiK77gw724rREIPSSDbp/aTsj
4yyFy2Du6Rzg7gTk71TP7iWaF7Hq+bg/p5XEGwAe4L7M8HdoGSGunEOR7vllD48K
cywAZmIHcbeaWd+AoI0wfzHfzh6oxAafonIQ3V4zekwyNi7DYjQ1M9aPfdXhRrbc
Fw9L2hJ6sKMxGmYqa3l5wPYt/O8THhqh606ayyiKkKNRn3/hTLMWwCQhuM0Ez3ce
3LaeKFgOs10r8NToMcmdlfs/oxCj/LfC5HJs335EDXoY182G2C6BALCX/Hmy2CYi
Q4tTOpjDi9/RKhwl5HHIh/3pC2/A5NQ+LaPIFhL5SrP3fR6vnI17fUr8y8jgcvP6
/fw5PNB1g/nDASKA3jduc77+N6axFZPiaIRxBPeEqVg/IjsGS22uSqoZrfRQAh2f
LW0bfW1cm00bQl/WoqtY3wHOKc/YtxPOMGkEbJpYb3jUWgfT2J0OmhicQicMN6cC
Rmww92OC8d7Qukdgn4oYktO6I1wX9S8cnQPR9yBEINO0p7KETKEiL6WDBQ6dH+5j
ssrufHVp+6MYxY8bHN+meJSLOBadCR3SV7fPEPdazusBrzYeGfMc7MzUHakt8OnJ
3AJndTkGHpEM1SZS0yp9YAm5SkMDKx6dvJk4xTaWvhfM3rL5khvaYrJUKePWKX6F
9w3KXfCArbfCzJtkhYWVha6hCe5YQ2d8aS0bAV1fKmpdxnscyW/5kAqOFEXj313S
m0c3zTAAlqZ9c3zQvI8nMHm8IZerpxebr2PqMJbF3EhSme7YujB/4JJ5lAqG+NVe
F/Gfn8qOqvKS5MtZ8yx32sulyaRig3ax/3ki86KpWRU1XkhMVsBBQA6DXqE7sPvs
NWeyeXMdlVd/UqZmJR6JSwiCLwTMB6PIocOzZ++FJA4jsH/Qojmt/hKZ4wU5sElV
IPkR2el3Nd6fVRC2xH5Wiscr3I46L25SePhNRO9mCLKzmZI7f3CXBGCOx91MjBn0
VU5UICU1LRWpLtsrjwXTiNoVlloKBZShrHamxEbDFhpUF2D1wd40bV3G06h5KwlY
Ri3HOTnzSW6ThI5ucaX8jEWUZAmoSN1H6xKDfGATkyLSQHxKvMZ8BWriuJR50c5X
VxtgnC1Pg7bABgSUR05C1jFP6bsYeBWW8ac7RJtNnQhWUunZlrUNixvkL+GELUMD
3cKq0EZEtSk7kbnT0va9gnGGl+9giczjsn93qj45f7gmbQJafHPLZupL3SbPhi5C
ELw0iRz1mavZJ3zk2F+8M2Itgt3BrtpAwhksdpwczTSAqRJMcw8/IwYe5+jUaNa4
xwHepr5Q7Ax4c7Plf9vDqvPZuqc/wbCJHJqYAiSBQz2+4/eHqxZQAUXmVnbVzxcF
g67igFdvc0+VrJDTBKK3efdnhrPAhXIOt2oU8uNKfZBs0o9avt2QWfRKolOv/BsK
0lNIPVFpzBRp5tpV0kEsEa5jwYR2+Q4woLXFG3Mxrb0VlltR5CAfKm9NaL/2sGJj
dC1Irnf6wJzREGsPPUJKKKNnwGAUlpNpSzu5HNMoeViG/oRgD8AM94dDsvA7UNfP
zkXod3Mz949D4+rjCie2oLzcYFUQoPQ6wkSsSS7dht4FPdf1zV+Wpf1zsMHjCdB8
dkTIRwSNlHguaLvzJJXdRV0/vojWwSiILjEvU4uatC0F4/odRInAtawIrk6Q2hSa
F0G3REqJmhhYzXr2x4Zkd9ji+NKJk40/fIsZlOH+ZY4yC1A24ULdanVcJATPSgDB
8SezMZTupUGZMJQsxIq0y3KxiAun9t1ExAyWqsMYz4/0C4pxIskm94nebpQUV/7P
U76MyJp/+xOFCn1lD7BLEUKJZMbtN3wZ5+zEDWfYUsJIMXs25Uu/n0erWVTv4I8C
ZvukJIrEZDFJwBO650savCXH7WOQrGpnyzpkztJM9/gaKNR+/Qc/4mLtcVgTksdr
BPhUyU5iC3gS/XiwH+52UHqqdgPO5p0AeK/DDEUUOc3OCTxLCkIPcjDRN2TDCb0e
O2BhrKqAV8TYoGlFPN+CmOD0OCc09eJrIUhk3rElc9pN/rcmiKzRUTBJLicUx1l5
`protect END_PROTECTED
