`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fn3d4NCeJ8/9W0P3FiBSFj4q27cZxU8aYUN2ta8X9SY7scc7bEj5E+88gLLBURcD
t7yrTJ7BAXQTNUXEFING/A2ZkZViCxTgcbf6VLfiZw9PFJQNUOA4yxbzpWPcf1bB
LJ4NROf9fS41V1itkSBr8MvqKRrEynkNS1lwN9ETRePMDBFl3Az2kpt+vUGzyyCq
yCThRUP14emYGkqDoGu+V9kaikRbsIVpXrxjw8CkO24Kd84L+4wODWGeJ7M1hxiL
IfShaV8itkDeDlTsdLK1O7adCnTy3OGesyiHciGCtaDRTWD6yrbaaaN89+JaXHcf
CD0eA9WHmFCoHeh+Hhc01/IzDKgz91gwMzV1CP7I6w2DSS0sfnv4Pc47wgJk3avb
wd1NJhCMHSZljMsk+hAkWjJfCuKygQsliDwRMAUXYjFxUssGOcI/kebmX3LWd4NF
wCfOJl+u5IwgA/Qw4gvYIV91w6peD9XvQBJ3LFKKyRbitGD5CezwvYwlWmEz8F9B
2Qs0VbVEjQJCel/8HQCCccu6uXX/+vKXhbRxDT3UnpgDwCIqKI40M0t/NtmKxhLv
wfXiuJhYV/exU4EW5wyZCfw0F0xKeIh9ZDHXy86O9Xmo0M59ThZ2TRz68x9WJO61
B/K3XlcHN2CKTiaV+vddj1ULUUEMpkBpI3Uy0GQdDzEnKepbR//NBhND1u41mVz6
7OB4V4OBj5i9SyEFpkhtH19NUV1mN2h68F98HKkrqUJq8pFg9KI6hGU4BowBhSf6
guYNK6Ly8OdNNiRm9nmnQHiYcU953qa3Px07HBlFDcOJSgnn2zD6kggtkumAs2sz
VqL8ViB8xMGFx7TCliCU2fl0c3Fc/YTOsPg6b92cMcOboF7WCdtTHjyrRgw9KYHy
5C7Zh8+CZXhfqs9ZlYElzgH6piM13pya5mKopZmJMbnHAZywNPA4lJUXMaZYO6bc
AOrpCgfpk3ZfRMf6Lxc+NqmBNCQl7QDUDyr672vRufz888zJuNcTVTVtL37UBbs1
y4uuggqOD1fY7SEBKDXjPZShoCYiY6K91ckWAn06lp0weLfOb6bpB1o7Rb0vkfYU
wgAMvYHWxxZ0h5SNv2T8HHDJ4Xs3Nlr3O71i3XpqQP+GGWcO6MjLOHS4oMAINmMG
unvcMs//mGFmu9KDY7c9nwe9tvxFTU0A9a325aowzclyANqw2mPs3ZRX+XBwi4sQ
PQopllJd4+vgPS2YxJovjupZGKpYdGtoLzYDohfVQHKMaXYOe8h9U206cNLQv7am
ei+mI0/FohrvGXDAQLl1ipA9Q4xaTc23LwEh/FYSEvn/AwFbZOljRSiBePiDiVM2
hqAHGFnsWQHbfV+6dhkuYXKqRlHiEkwniKlgt4dthW1T1BH5jEuCUaLgmUV7W6v2
TDJd4SYjCz7qvq+O450DJp87bInOzxZEHzv5gL8sHNPzzd3KAHIPP0VMG0s00om7
S4Pa00tN/Z0VlmtLKTwPz02kLb3vNADd5PKcY1Mh1Kk1EESbvwLVlq1w4Wf1YRBV
Cc03nJnDHuhFfJqrXEFUgrr7OmWZsyw2VgxCu/WBIi9qnRl5rbXuComDRPeo+wIE
gp6cVNrYgNj5nQY5jUYZKXvifnM/gnVK2pULrYLbaiXT29IVHfCcBW+9/13nUDlL
k4XGfKmi4CkozkeZ/LpE2B3YAj3NdYZEI0vNM2DVaRsLoZioIjJs4EyE9p1JPYLH
EhyRr1YH7CwHH1OcLllVMF8JAou+36r0Qv+uVZoM7gRgF513AaNbVhZHZHGxp8LT
+6RomRmP6hcaOwKhA0rLgsxPRwnVfdbrNRymDmIf7F63wZbcjhzmlOJsLJblYwxM
68mUAw6Xa1O0vxpE+cw4hH7AsennVfIUwOxXsfEBUmkdXnKsDtaBMHwxYmigdZRS
knjP7243b85434t34GJ/dU3xNXWhKsW0Dlvjz9aRTO8VohWv27lP6DQ3sGYvVYcl
QhCVfV9wpiu4BiLW4GifYui3FnDyRfsr25Dim5HkLXi749/eokmQO+bHJFXkwAt5
FIlg/l/9MIgdCoJzO7KCCeXvMe7vH9EtmiFg99+QPjp8miX37lcvUSFAvCoyAsMS
tNI52JbM8sy+1X5Amz/4TtQhbL++Gat+1zB32aYnJmxBaQ20WzHc/Oz0grzXoxvj
PBLuEhv/Y7HINMAKEzMicAdsc3PPnKq7LBzuExT66FyxiVM7QUF0szgjHNXZWQMB
HD90bF0QMvQI3SiSASSpuNaZ7mz4h5D9ve8O7SbZMUkOz61IEzkUw1VFli9BFTBW
bi1T5ilu8nXDqz5Ro/YFYFKJtqDwQWkZd4ZfbGTrRLbHcFb+pEHw+/XD5H7f7n6x
GsUB3NUhrfH+HG41Q0KoFz0aRvDqgK37ZTPZivEjoORclbmVV1RhuFzyDgqbuUMa
5HjDLe9PLi394E38+cyOdy2TQchZVUhSGlLbC6gOku1Ixju5m/lilznyfAky6MYx
66EGId1XKP/WSG6jErG8jTwDHol9lDR/Uxf2Qsgyvzl4teA6CdAi0N34rlYvXRgH
W//lQ2T0wSEV2ELVmGZ+78bmSDe7fk1RsRSoTc2N9sH3OlRVgHqU7pxw6Bo3Vuip
G6KxJFiRu/fbGGVJ9liLhNuFhe8sx5SiueXpYEweikQJZpJ5WHTG+44RtiLeDHY9
/gy4qicEV4WuxtJQ94YxRLHkQF36FBG45gEcsqdWNqh3ZH2jcPS2dyOphct0Q2DW
2xt4WdaKQNgQNcXJcZfcXcuVoY2tcWMbitCMzJn770Qg2e+xpQHiP6FvZngIFM8v
6KAvhuj1VaXBx/rcT2PhFR2YKfY8LdcKuVRKqy9RGuZpLRtULbyuG4X/ux+HA5vo
Z7RTdwrxplhqOnFeWagYpTw4flY95D1r1C0EchCLddcIuWD5IU+Wv2nmRXjKOWTq
DrzDQcOd5qNx27dFIllMCqbsf/Lo6BOKokYiHRDZoCMOZce2w1l7SKF72KEuvgst
wWa2Qmpv5uDU3zEYhyfftWURQkPPCh84Am6Vose5YpJcbvQT5uzSVTuYMJmpJjLK
RjnBmRGGNiOhRC3ydGJJgGDGdiEcS8/hiE370V6iyACgJ654NkrPqQRMmOLgYg9v
xh4siVFKQNycf2BNyFoeswVtuLhcKIei78cWOG4gKT7XHmj7LxqpAQhxgjtAl7mw
Hkcw0RxITLxCFX3KNgl8FivRlqvO7/bzWghqaZ80VjZ2xfGeq8rKdiEsrWNUXWwB
Hk85Luo1JGE+j89xg91/Mt7KAQxlzgr6MjaJv4QJra/8EseDXjL0/6HwlPLEYeJA
7dkWYIxYfwShBf8QwNjzWC0AAKzqBTMSA76gy6rdhJQwYLvATiRIlbppmYCc3myE
Y3qv87Ie5Q7Jq7Pn1KyMJ175JkBcfn3Uhdly3TpxIeQWNDnJsFWXaUBWdYNBzj1D
3EE2aWj/Ka3OpvKHaLS6RgP7v5fzvkG6MZbVTqLsL0r2y4bEOKugzZVMRkZ77S3n
r+e2nPNYwFS3RrVBcJiyie0eKW9gUy3ecAvGaQ5VF1EmFqmWlvHHy4aNQndx4KOf
YHPlrRLCAXnZTE7M7f2B73bI58alsSlaFR5DGG1F+CctUc2Podzs6YE2Me8qEyGx
5gSfm586GAjG3XsUmzGZ5FYZQPSWV2D8VTL+rR0j5HV2DxUQ04u9OHrULGIFTTdW
iDQ75iwlNwiV74tCEEHhEI58nfS4NqE6P7PHjTUFfieuvzHM0rbclQIt0fPKYWB9
0P3xHyT3A25h1f7NIkozNatPXeyJxqkrKXRk0bMfqNcxmY6kbGVGsIHElseYUS+B
QykIxjyVsQwcF25EAR6zsV/XCwouNlqmA37mmYDLnvpW5WWv66ODn00n0p0wGXVK
VnmQdRCqYvhq83AD5SncUrqDfPEBdK6fgOkFsa236IbjVVuGTPN2geoWGsHXpKSw
p4eN8w11MR9ATKoraWw+Z4fdlhC9TeBVYMFTv7MFNo62RQPEpVKAn90aPEfhre/g
SnQLtn+duvcI/C6/X99wBNN0Z2oYz5YgqoP1fR9gTAr0wPFZtiZcDz1a3Ou83+vE
rYY9RfaDn4/L2Vks/amdUVypuZQWqGAkR5OupSRLEGv5MaDzNaoRRQznIzoIO9Yd
IAazUgGJgNZxKkYkp11JUiJwy/j60JosWty5MW3B4f0QduR+2jm+qkjKza5gA4Xn
Y695v5jR7Q9jBwObWpaL22jfUE3/4G3qfyGmgXi4LSFfy6XQheAAzIAIk6MheXWn
4vG5Ms+aEp+tMA85Tc7q2uSoxnh4Guvlukd8Oyv17aNKdbJvyZzXb7pE22uOEop/
qSueuOKlBVlME0UCxTy+1cep57Sc/ipgomSMPlcbz8eewfkD5l+txBkA4yNrurDe
m2PnQcAl5xEpkBUeRmtfnqNKG15aeoKC77ZqtlcqrFzkm2DPUyyuDms6hEteqR1J
lRoHNdSnEW5I8GPDxbj/Q14PYlpdpt+sbduEClwCcqv82e/oTMBUoQN6bW3VHU9p
oGcrs5dzS422YDehkjzU+w2VEdBTz2fsHRtJ4ExLMPLOJKE+reZAFerNT95ruGeu
CbGnAhKU/LQHhgUZRtrqnV2HLhgDVsEMYnSNpTIanc48EknatY+5v7afj5rVWatp
C85pN38qrIid0EoUGYCqGjvRNwFbM7WxClSg7tyNrmIw0tM8dmfxFehdtUKBdLhI
jqXHREBznWPtsSlmZYfUzemwNaA6BKkt1bLMrmzQCtPAKtXgWJW8RVeZ+m6nuk4w
VJgJ8Lf6tsvFi5SvmgBhrGBwZPNXR9RhqUUQMDfJ2RdSkd7Mf8arCYV+DZ0/TqD7
2Q1qfwzzZ9sjjdrzMVmghb4hNJlGMuEKeqhOPwcWX+h8rBsfYxAYVZc6vtt+QLyc
DVtOm+LE+G2j7toNtXGg4V4TTOjErvJ+7c2axNWguNqujcV5i+pMh83Oc9m/I5NZ
lLcxpUQ+E/b66jK+acmYo19Fv2sG5N0bdSB8Jl0Y8DUOwrV9ww9MHVgmXKW9+jKs
T8OvN36FViJySzcFcjO1OIt9I9vxIlraEHvkSdYDcNZ0SnV/5J+zHxySZjeIEbjm
MJiZjg06KWXPMvlujGliODCRlrZHvyMkqLGGS1pAj6lHbZviak1d0EsHK4wNQRRv
j6C2HNKYbiBek1MBs164Wpai4c/UDk/AcMstwPPqqrz8HSUWGvYyWnRKfuaYeFO6
RL0Di2TznbtbJ30qMvPif57WSkxGMPSRUtCz7Lq0iRchCveJUE76mGKXfmttcJyN
htc4QEIaW2pe/mc/jUfudUlYD6jjEsA2VVSHHul/SKhDzKf4pshaatps7shXYCDf
sC1QGUi61Ns1PKAIcGJuUm8hHq1uQ2P/6zGF7JPREaFTOrD6LzdH4Dwl8hOtXTrs
a+Ax3DAGIjxqzJsRvgD26spiHIGh6GM2/eQHX+eWr5L8mIXD9AZCn61TNVdTseIO
Qhy/8TQN0ypYlxMsxwXdOGph77PyyrztbuvIWRnfZGMH9TEhzamD9M4CvLRSNqOc
NpRquAir8aQRp7Hu507E7Fq+/QFnNp3k029zYPKehQEOv0u/zOSfZed/ZyH/DiBf
y9SjRfW+Bv7ujGm3Tljz8cnR9yKzMR6hAQd3QMd8TaXWCkWVqW5OOaBsJcyZMVVW
pTBcVf1ODei/HKLqeIZCQtFPoyED7NOrb4huUQWteojvSBdFkuOb9uFV89WMRF4h
dzk50NHOVw3yqbkhW7ZbqkDq/a4ScebVzKbKTc2cjR2ZxoyzUnNOV2fob1riED+I
pb/5EgLg+AGolDys0WMiGEyFcPHghr1GmYXpH0YQc0O1SWYTKyheWwY/cxUf/pzb
`protect END_PROTECTED
