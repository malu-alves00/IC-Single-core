`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nvz+0xiJVi1kDRh7JiWlwPOZ0x3NF4AX3YSFZYjUZn3T6G1AbLeiuIqXZF8As6OK
MTqJVET6Q1A6mfNxTI0RuUYDy4lxOGOVOSz0NARicUQwyxh7vUwkKmPZlkNCqdui
gak1rF0u6pZB8fhg7PUrEMKK0Dj2ymaIqPcGdpDWj9x0mhUDhibQ1goGVLgKnXno
8BmI/UcWHkdh5LmM9WF042s439rWDAsyiH2tkc+L/efglc54gX20RSMhyDcuDME7
lH5s2ViLHegylz6dD+18uoo5R+eMRCETnPmEjUpQoq63yILlvSpuoM0dJt4HVlTO
HGYkuyKK++2FIVYN4vcsihPCxofNAMdS6lc1aBU9AFizmTeUGP29xE5Y93/kL6Dg
5CCBU5pXiPA0ahn1DSFaMGxunlVEU1n5Asj8KMhR3JdTV8RWn/tDXKpDYLYd2Xrg
3NBvabgefKK2DkNpoMXHZlAOcxaqG90IfpjE1KUYpBKywiszgYKEOK90DQ8H4qUf
6tbBJQ5VfQtwvKIU3GWIGFKGfEiMxB/9PetnSFlgJMw0lTyQQygUyfC/UISUmDYi
9rA4k2nKIaK1wqt5Bt0jxVHWSikJuBZoCp8VaEGC4cEC1ZaMTMiL3psq/081p2y/
Fe0ptxt6wTRksaE2x1JMq423q0KWFJOLPAtx2QXhCBz1iPdVoCta/5Jg+k7POLu9
2Zqc+pYczhLHUft9uZfd4gNq0ILqvBiK6y6dNnyhM23ZvfEqPqZ5p9U+FrbqNggV
rVFCt/QgBQh8m2Xmjx1oQw3ISwtd6MBSYZddS9jxzGyMdHoKPSfY/6Rpo0/6xlM5
ncmK0rn1Od/w2RojgKOPB0hex0Cs140RSh0nRoThDCrVain8qNEm76UYh9YOgy5c
pMp6HKCpRfyhxRnnD42aB0FaMeHnyDlx+v40eqBdNHXC8vgY/Vm43Ak1NCmw5r1t
ldQFUspfFxSponfq1Zi1r0y0TGeHPOBO10yhE6JHFDmaIhhXObx22HzXeP5gVrzz
K8SPCe5q6fekhov0okV5Iu7+FFKctzoXVmXQx1PeYcaldQ6z8SjK8RX4fyuYs3y9
C0VpvBGsYk6f5iuxHVfLIsrEMmNaeEM+tRASlu6Y2i6jJ15WOv/sfD0P3xaW8NCZ
fZUBQQu3ekAyuETST0FM2Valg32xlmIlaQ/s0KvDp9E3kiIFinxwvPHBtzOFcVPJ
v0wZhvEcmuKnS3dFdyZ059T9G1oQzmvqx3m/Wc2eGOSICAtBDbBB4Egij9qjMjDh
Mi6MLBD1pKvpNBUI0ZSteP4raYxuG6w/kuAFivReqbY9cTFQDAs1v4QZJf4WBF0B
NAFlwGAdzyckRWIKGY1bPT+NwxoXplKkQgWMHQIzNjd4omEBUpBXSw9uJh3BdgsI
d3uPORKQzqzp8Uk9BcbsrHP6nfDB0nZLFWsn/Slxr5BS8CVgA8sZaYWaQbjHfn71
1B/f/fMyi+GazaaSydltN8oEcyfYD+L9WAlZdd1pBlrpzvl442uni26GnAPE2vhJ
BvhXIEZMPq7OrDZ95wtxVkg5YhWJGSNX0BPZ10nH2Vkbx+8MyR+FNSaMxyHWLHTW
Wlxeq4oqe7dQWUWshe0N48o+Atz9pjUOKsXG4HsoRVqLfnjCyBbk5B0TObFYAyIl
xrQ9pmjNqXWHylNYVD8j+T6CKe8O7e4FNL/TO3ibwJXCcwfAw66k70y70HXkOtXo
JGCcDneC9V4GJA7nJ9UhNN+cLEGd/71CnIrGlYw2tcJvLtYeKU8s1FQW01QoNX5I
YB0orBcLCtaPNFL+exh9aVnCfy0RDlraW2CeUd/ts5JMSkA9h6UEnLE5PiXBKiLb
xWR9fEm3N/YrmgqSS2o7cY5gPQR3hPy+74vuXlw5427hOwCvLc0KGFTRuVpjo6bR
qkpA6U3JQW4U0BF71U6Ql2BzzOA8M6RPwu6mUHaG2Vt3UvnlnosamazrIwEaAx/H
dERlQELMKvxwGBXZrIAkE77lOYEXse7lDWLLLlxkOcXHjghD8C1pWip8f0EtRDde
6o2qUPNZuyI650FY/Uo+c1fgJz/1tqFkksh9ii6z97VXkU1mMnKg9e7dhfynDVOw
2fvj0vI+5FjdxEGym3BWfqukKAC19qxUuBpATxVX80v/5vzDuJklr69KymfVroyt
gojAdN4/i7g27/rOZp+pN7DfhekjhSIIfalDFSOSzVzuKyP0qIKmYq1cn8NwU2yh
AREsfvhMNHjdlx+J5BR44tJrCYtPPshmQZpW1fn0bBpE0TjyRl4szwvvB1udP2SZ
UNumSevFXrVxYBxms6qqY0bC2M0LaduPYY4c68d2RPcbi3CkzqcjAqqRB4lFZMzz
/M00S/h8YckyDr8mxmGZtS3KVFBp/Ruzt4cDPUFmFZQweT520pGhv47+GdxnX4OM
zj+jfCOp2QeKCbDAmfZC5PhcutvQA9P8cAw1ZsoqVCXs5rav4XPjdsXgY43/XDzh
rTMe+W8c8ZHAKOuPkbtxI12q6uCZIHkYSNBeJn05iRPlsNgD+n04H0mCW+zaW1kU
XdXhpRoHe2P/LdwJijn4Path6hUJcrf1OooAvIsALpLgxPv9uSmxI2rD0tkMAnJN
XCQfQbyZKjAzbMWaFrjLIPCJ3qN/Rr/CYT1fYzo0rwCw2QlJjUZlU2Civ/71B9nz
uVDjRQLnO8PrRZMl9dasjglI49QC3egtlVWiY09MrnYZBAf84Y05hRi1KSAsKZAa
D8Bca4ulxG78UCqsXhay3jGxaHp4ev4SUnTCBjzgBqfihRQ2+477CMF4HwWf+vtM
+/NtODNBJeO1IT5CeaA1InhDbrR7BVNfttQ5bw9r6RIyC0bk+rUwqyNeP+vGcvrG
9NUe+hbc8NEh7/bCniYB+dQdqxdfNjO8FWvfxZVW+1VMLx8/tXVRHusVcMARXsvh
a74gOjeVsRbcX3Ona1lKMnhqcdgKRn3xcrCM7be6HdIMTBlqIYIGNugYjpqYRYWp
O9czfWCzCzarb02X3IkS7LaL+NI7TErGrjwshlCWWyb6nmI/54HuTNJkN7c/SwIu
+eMcZyQvTWlGqpLRdlfS1clPSxu8qHxOeWe2VK7f1tNTiFScRfjWnrlQUyyNTomw
fFI17nxrge1RZBr0WEBfTAAUNAZm2ARhp1B4YjlcUK1FwXKQf/ysA0wGxbntgKu4
UdSxprhDFi4hlS7o2dYX9QQEHbtQm7oIggDGZIVpiWq61i0zjJ/hdOxsJMWn653o
IWssAmIbbUjJBGoLg9a/OH9VMc3KgjCD0TW/o/eZiE5uZJOiFCNhwb94kUEICEvW
BWhw138ftM1zduxVA1KgZV19zbu/eGkNSYEXO+anEQhY6RmilXoTL6FmqzD0rUo2
IRtca635bevTlKnX3UEhZOWvjhJDTQ9V9EOiwV2ZMzc1TSKZj3Zd27jdvLu7PDuc
yhpVix7w804p+5NX+Bj2Q4S9cuL4UxD2FWWEU86ijhH/S164D6E/aJJWpmexrji3
25cpBTx+xeYRwH47GMp+48dnMxKvmCpgVtFCaNOKfKpFMFSsyfnIUnHwM3EWlisF
V6HY3UB8tKU5W6ig6qRoSXlflCvyYVPJkwIiQxJhrytf/qo11Q704NvIfKV/MKpT
`protect END_PROTECTED
