`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
P4mAnQ9kibQfQbo4+efzdpZcbyfmW4fMudEfgBN5enT0MywFoCb9hwrde/iYtNX6
nu9ayVhHKFww+5FoREThW/erZvZ1y4OMefi0Cdb3+N5/B9jrBIQVsVaxF+uKINDb
5tFJfmVZp31DTOcfI3nD/m2jglrPf9t5FzkJf80l4X8pOScN1j77qY9/jW0xvIIk
1kmOC82zh22mgT3tRuK0GxDjzRAc18EIoZqrTnFb9kd1SaWJa4N77ac4yFjGnJRa
rEMuBh6FvpOry6HVUH3rX5VAgdEESHkR8bndbmwXvSjHDt4WvH4zUugKiml/nmJA
0IYd/blrmHlFyl7BWnfCIkIX2E4TtOkdHAk3QQZ61ecsR1rpPU53XcE/5udCKqbM
NOHX7z3vZlrfn/RA+2Zv5zIN0esGOuiGHwPoA71dEMo/OhL8PVNB7ZzB/jywGr5V
S1cEsUUtJS/uEaGBkj2IDsS+e0t/JuC16regOhPIzWtmJW3b+hqNMsUr6jLz1iko
J8joVXapeCtk7kv+AHjpxQsfYux3aNW85ulKVbgLp9uA4/GibPHW10hTtX6dci4r
VaRzs4vkKvuK3iGsDpgQIBXjEU+HXjfCTXf8FqJ5nSeo0BOHkgQdKJQdYkI4P+hc
dyhRKhtwlTYiNE9oyx6iuz3qk2eCAx2wAIqigUwlZ5NYsdWLMwm+FjOB5kuwuevt
E73Cjy8uDOdmfuVeHey78LA6wWO7aNs3Ss87IceXuj3ihAiIZGqsVyFGdUfZVrm8
FO9XIeVs3HB3Lcsu/mCCbvby8s9gZEMr9tToHYefNy+ZZBcP2+y49ip9K+6tQz7z
vhP53cJhW/pW4rPSvGQ9wW7EOY61fmAe82zX2x65IallQUYelkTE4iOeEwbRaMB7
Iu1qYI8/R2qyU4Kcj4uOd/2emXc0MN/v2SlsZ9jVG/my+NV1Ivp5jQho1mQ3BTKr
EkK167OkYI7kTIIwX3IHXACTA1/HXYnPJIhbKnY8IQpjEybo5+2+35rlNnBxY8cV
WWXmKkR/saQtdV7YTDo63KLAmCTUL9CQJudv5+b/WI8Litvrqf+qJZg1qTKArG5e
ddTRHhsan4vMbvcQx1kfRQ42/MEGGvisKLBz09Jf7gGyHo+cSoOYoXSrUQ+3BuAA
CWl1xcvNlO83BcjHOc3e+R5uQCe2Zfw1eMzQRe5phCUXHhVOmhh/t/Ze0GzAQpC5
T5Glwb5Vts9X/E9qQP3QkirVyn3rXy8CA34s68DuHOQkrHmhCKTs9il8x3jOH9Da
ifTry42ZLOlghmLIlmX1ofc81VM9eMuGe4OKlIStww1bmJ+TwMClDXa+kOvpDzRA
+tZyP8vpaLcd/09///QYEyro1P4d91Ew6CzO/zUBIBLqHtI67Dwo7hjamm1P4Zrd
tgVCiYjuJ6P2G/igciCkSslpBK5wm+xtCfFaYbuaxrdXsJeKJfvkJ2477BSAWXhf
NHrr4CAPu+bWbTTmoUBlJP2FCjZmNRNmp6ltB6rywsCQnZ/EBqtftZhANXGUNbgj
KOXx4Lg3TQS6r8a9OQmcwhs3M+uEinxzbsRnfOeTuFjgg9JSTvXJWA2F7CNw0+WY
qc3rL2Zj+vvGOIcpHEBZCockqrD8RQWhYsnwHu6se1QEYoPwLPICqIysnyu2MWp7
o3FSEByuLi9NMkNzGTL1fbxNlUf+JO+joyfR73r6g07ISJtfKg1jrAyTsLCpRVOT
SAN4i/NMJ5Xxv3ldVYxoQorBN1ha3E60wHR+zdC1WzULjb7LBjoQtCqJpqw+55FZ
llJJaGrIWO/BBS/VGoZD6ja3wr1pMKrfmW8UCfhPR0rWgHsu7e1Gxrtw6TBtldqk
x5/TInRbLwIHJYZYJyzyhXMWdjJ0vPpCN0Dye424E1+7eHiIZL7jdBSTrksJJWEW
uabhcGtIdQfYcTCYT7pd4s/hUhJYKv3ZPTCpMbbmbUYPCaDOeR4L6bl6hCGQNhcf
e0mBCllXQKIfppajxoT1WcbBT+2SYLQ7TdtEUe3inCFiLh3BBNY5pUaT7Gfo+RVk
kpUWi7zPzKhiByp07JVB3KZsdbNmDXQpHEwd3eIfgNqvnf1FAISkn++eGqha+I5o
9CuzG5Owi+FI918bOOJffU8zSvvmPrJMIfGKIsB44f6oRmnbHzg96bc6LYHAtqSG
UCBjAmwuBHQfrTvyXfAw2J7Pe6kzDLV9HEppr72E4L3dh+YDeLooauRZpM7T+RKO
wpEudT8kiiSMBS7zIvzjkeqFPYwxrEOu7ny01tzzk2fmcf6BYcTtFq9nK4eqHJKL
Pp6G1aIXzsmV4SqSPwrDhzjny0Dm/Ro+exOeKcCVGQCoKTVYCU9HfcQV7Kg5OFLf
Dxlhn3MCqUTwBBCtsyzOJMCFQpfiM4TtSoGK5f6WuImolY8mX+42pwlhNVb2Gips
BL1orDaD4pFjyiA0V7qCHRvRP+eQYc4V3VBmzS+Qd28MfzyHF1qlRRQL/tK9EEf1
8HVl+X5MgTTKj7XWMzvWgtTBDqVHDbAE2mjNyeLhFp06M8VgqcQhX5oclauF5eBF
l1S65vck+nJAAuOaa592zltfGxRLB8iVFXFKvDRc01VzcXvaydJWq598RIL5jvo8
UfuhpF+1MqAJAjG4x4N5+tpS9bRiLl1/pia8w402badezvC/4wACMAiVs7PohTZj
zs+s0V416wmIHhGb22sMrp5QjgMjsUSIbh8NN3SFuk6oX8nZVUKoqKg2AksiPPZG
d1fsnrybms0+3/qN+DUNhwD4iCBEFKqFvw3d3594ZVKyWgL2TTZfKC+uKF+dk7js
GS7OKl3b4OKn8auGdX3qBgGgAA+SSLv8V76fo6d6U6WlyyWeFrDtzSkGvvSJFOW4
tPTYL+JmnXuZu3pUyTszZinvELCH42HIr+hEtH7BlSmZXNa7Pvk48Ljn/9bTp+vr
Fjp/A9eZJPBNc2Ax/1SeCTl/jMS3YTexRfCjcRqa9M7MsLj8oAVI9Z9BW01xyFo/
wd3+lDohgokJO/jtG3uR5dvsP4vkbMVxtDx84o66saQwoGiUVrD27LXSeP4BnXzD
g8Es49JS4W7vzEtJCnlOJch0IPgO6+/W0T1+KmqMRDm1t6t3hbEfU6MaUrWribBs
w1+wfSXGOGKaYwD6aUgY7YcCLOhlUJ7vTFPFxL27hU0xGGYz1dAr9g9paNf9MeX6
+MFZK/5Mvo75/Jl0fm4TxGXKQz8Uren29HvcJNCbqtQna1xYdFsSU1tfq2d6XxhQ
temRHaRp7vNXOaYVSAEYhQdUCfJEfR7u4aQAsKNOmR1RoiMBJYdK+3QknNbZ3qgF
krIG9XGdEpwnO/klroMdmsbms/7T8ZnhbR0MsFJ+3OAatDZbIWdxXRMgteWYYGGn
w411ExLDjb344eivm2Lf9VHEbqC8izY1pOsxlkuNx3Agk5if0/NNxUG1XLzNXs8K
i28O3MbNfVhakZCKfQLtsXWzh2G4h9oQsl6kh6cbkZw9bEbhbjJ6rMckDLlDhxQ1
JyDZzWPJFykt1LwK5wymIdF+v7EQm/WFLEsUXydhI+p6J3b4MmJLYgWOVE6Hl+mL
iiTEpF4dwEthQJraQmQB9MWLoNQyxeY+hCNDuAbf8tGzFMhJePy0/qJUCLKFRbXy
6AePvaamuVDx6u1CmVkKehjKxP87a7PZ9vNnqh1+SNlpVviOE4asOMI5IT5cU35l
I9VjELEp81trBEo8kI96Oum2rKyoG08HdyuYD2SxYG5IrkgINexZSTvoKtvxrM5w
Wj3sPC+WtXEvqhY7Z98nD1KYQAItGgUcSNXI4Fi/1XV5aNO1CKHeq6BEXO0SgVjY
x66Kov5RWekx93dcJAvweigO7ofYV/2IdIySP5ckPq8so3+NWs+OJ7LazuQmh8xa
WsBvxFYnnuIkaPS2IUIJKM3WwLc69ROslMbJ/lklv7jcoWPVjJEXHff2XQdpfFyU
LPHZd0bzoF2B+pXJAQk3Lk+HbpK/xYCcb3QEyuBAiFbU5cu71+edMLoMNMb2mAYr
moebVacU/nCNz5uwCvi9uHSJGqXEMoEzfIUQBTN+FTeAb3rZI5168hG1NVa41zdB
8QPgtH7/ihjk7k2pJ5Lg5GPNm7xpkl1O5zK31FjWbTrWh1/D+osZgGj0XD1HxCpN
zK5oNQJJLvFbFi6OkWKDV303g0Hl5sCiVZgz69/L8z30fmcPKI5uoMdj3db8MHG2
i2gRzXmgBn5/XJeX7Ou9xf+wluaQMSf9SlpZpmO24YfEM06uCqgCTos4kUQNC60Y
2SrqGxS7RdSYUckcwncpreHFWIdKEUcRhz1+/XLjEQ88Wb3aCGVnjPxT7Lw0QAVR
YTS+V2iwIZqOQemeyjJhS/Rm0leizCxz3KD87ANQfPF4bOcKXmskc4jCbYpxcWL0
m8XmLvM/w06f8v3VNX+Z3Wzb/y8Bf2VQPDO5XlXZRTG5D73jScwULK7+HQyRwkU9
DkIN6j8PTetpw1fah+fuBCohgeRmbk2s+18mVtXT8i85UTLD7WhARiAclLRIOOEH
IGejoI93h1zx6sncdIYPL6Hc3rIw+Sb6+ljr2/98XN5c/2/oejPSbDduh924hlOu
S0FPIJnwKYr0SQhuvUUuArBPhiWcHB88gu5IHpSjwiMDDQtgMrTxMvMLtmrdMmcc
E7qF0vwOKHhVaN3DGIjPwzGULfgrM7rZo/0qKZCn8tfeLu+eiSoL/FwXeRsxoBVt
yHHVSGU+T9Pfvt8OOJ+S1bkOZPEYhSY8pX5qoAeHLCMki/e/nx2qa3LXU+tT0m68
2dw0Equ2GDhx6N0rv5VpT1tyLHyV3y+Vo9nXqkX4tnHA6PqRKqJYNLmXCUfmMztq
QZy/HctcVJ2+qgh4esYWFgK76eCQwFA17GWIK02OC1v4jojmat9mosuSJv+YEjjX
j/Z5Q/oa9k+aCsWjSy9eUpZyhs6/92o0OajCkITUQ0WOqu3MzI8lfUP8jICH80zf
5wuZ6j9BvkRcWKV7XwxhNlo4LClgx2OjX4yjOsmSm7XCyr53QxpC4npraDDw4S4n
l8v1CeobgD0tVuTYPEd25DgUDJblp/9UFwBEPlsWlDIM/nCVEI5N0EVQQ4pCwtIW
HihFACOJmd0Y9UAR0YytHgv6Vq/fmJl6Xqev44Mx3b5aApJ0knrhNbsCO6ywgEIC
3N69fh22w52mb+5Qu00wbc05hT12jtvL5LyvQhtyGshtxOMnwKDOcJnl3gsvhC2z
MR6XWAIV8QAs33miGpYiSKSgwRxVGdysewKdDLok/0zKqMOeHLCUV+qSCqSIZNRA
GCrnn8lOfplitIWcsjbjnXL6KFR5tXILmTT8+6qRWisoZQCIzq4ZDsyyQ3yrWRzL
IGBqv2SvbEYmTE3T0kQv5FJjS4TbFNJBVOoZNn7L5iLCzGn5inkEB6SdfR4UboCE
+N9y6+D5Cnyydo78jyECgh0HgHMV6e2F+fVIG2nGAp87exY2eNBuYpTlY2Xgp1nn
kySwc5CCTaFswdhNvV7MdLErvTYqCQr3i4vXCe8/PiDeWZGXn6sVIcuSOQ1hYmL3
wdUh7+9b/ra/T+qSkcmcGbEiVxconf0IgeMcwglhUecLs4TfLWAqbLxGT04LKNx7
oTsxfSJFlvIqwykkPl4CIbWrnfTA6X/657X8UxvYpUgCBE+ECdCFJF7OtZAuz0Bw
oZzew54rn3+xlwzA8ciYXXPHCeucbwm/p0/rvnJdLcBESDgeAv/XrOjKqnWroqYv
kNH4X5h9rxfRYz9k0xwaKCKZWSW0UquVzicn8n5o2bXsnf/uwQVs6zjCjaVAwG8F
nwXmOXDbcnOIfwMrCT7N2WW5JiQd8HExnUmAF9guyHudmIKRVoxgwcuip/zYLnYt
5XRjQ12YS6TMkpjuiPQfJixD/iuCHC+FK/Ncr2evNN0133OWFkdlbUZzapa9bVOk
7C4p8cJSXh0ZCgzTo3w1B/hKLB/cQq8xH1pH3pihKd+vh4uzyB1SXki+wqunS4+T
6eZSsx/yapnsJTBPY/Jbtj3tTpD3kfbx92kEPf4cQI22J6gTQn6T1lVFoxKV9DbX
aC+HB1927GvY0YbrPts3L5YHdHe5an4fUdVH0SrjiZMRH/tqA0s75yn0SLv2edkI
0NVZ2QelDZxz0Ojfl4Hvit+F0NrzU7kYi3MCjS8m+9cDUxWbMCJWyoNVd0Ui1K9p
VzWfoETWKEe7HYxZtcyXAS0Re9QMaTvB83F/fGouJsqCoVoV/oHR6enXdbUK9L/1
MtjdwZ2RPktsfrIPLfnf0YT9LeV4orih6Zr1C7+TgWEMQpLNCo9EPZLS+zyz2tQz
6tXgtkN+Z/hxfOnwCP90GHgqMHXbj7YfDVc1OO3Nw1b1wA1skTnfT+QaShqdQKuj
kxbE/ivaE6i/vJ6S4UY60oXQr8RoItkPZu7oVaWAEcp90YPSaq1Ef77Qrd0Nz176
Rehz86k4CQfXzLLyIjqCdIvg22FFJiOEmePZNq++rDCowddK/mvxCVsGn3kVLLVl
mXXLAkh7259ovyO23ypLZaSzqhjzUku2pIzzI4c2M4CwvJfDlaN9b+CJ5QTs8Bx1
GdU9lP4AL7/Jq4jwzVNPJrug/+PDewyZyE+5NsmTt8VUxnnazKnioYYrWCDPMCwR
b5H/cWeFtnSs0rn61CaIOmB2NNCedCCuLbdEFqZ9xLTFFJlvwrY4yO/btmxmZ4vE
60kw7dEHo/rp80dmxxVYGYQUtoE1JUtWJQsDbpMH0TwGSPPZ/HxKMkWjK/i3Qp4a
XW6Qx1RJEGIu0/aWzIjhEUZbPDUq73XfpdsiwNE+aaKqpCIGqSFFzry+TAID0mA9
`protect END_PROTECTED
