`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RymjF9Rke8sai2nyWwwd9kGAlFoP1DcYTLm92BR19KUyfnymCjV3RZA2XiyvK466
q/bRNnTNEIoyGjMrCidY0ss4VZoHhipWhFlktb4QnEGeX+oVCFQIgWenYmY/we8c
+mKrzwcAq2BQySek3j8fckAQRFPogWl0NEMoLLazgH1zsjqZKeVDG1pXC17ss4Di
UFWsBQ+DVqEaaQpazanMuTdfZgcxO6rUvORurRgsEiU2W3eujgXFJ9s/XjWBI4kv
AMlGZdoWzwyoVgCHXgyeGdFMubB05I6/ErnKMp/PijgfnzAR4H7FbtcMUMtpxIVH
bBWd/gCCsAnEf8WEnMHgt/TYMrZdqlZMZRyanKGSvKp4M5Y/bn1B2d2vy3GfTbh7
Sn5AizSOaDzrnQ+DD/I+FXkMsIgAByjZ8HXrYQNOp5hd4yE4wecAvhtn5uo8de3T
SXPuQLJ8Ll37eVhpiuQhDeIWBF3slwWukIWkcY9JKOLL9Ja0hks8kpUW7jhrb7jG
BOTDHiY1t+C2DV/IpshAJg9c1RbQCVODqiETPl/XfoUUr4/VH7N9M8xbWjhC2uDn
b06DjrBkfZKp4Rv3RnN6EDpumFhgL1Ru2A0wzNAeNlSLgEN042+nALQ6IN4ieXLV
i5XgcAeJQQJ6/VZ/CkA9k+ZKyEsUzpVy6TdQoxXwhGdMXSSf29eOK9+828y8FyxZ
y0+9dJUnunTBU/Cw5ROnRrA6GdAEmMKdpGA6ZvSjTyQ=
`protect END_PROTECTED
