`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NI25kB2FOwNRiDq8k3DnPlTiHYw1MtuFR4hkZ+5COOXMpaUn9r0THTGXJ84W+qRY
YRoz+jr07diM5fOCFBXMdRX5zgeUHRb6H2Bu3HO0BJMWjIWMMybtFoZil6cAAiLY
z5C4ypCN43j1vRBsitVE39QkQThn43GVPqMXt/DCOK+as1Us3fGzEU7lROBoiZ2t
CHmjz1w0hvQKBy3q1omyEl4DXiKT8QqbBN+UqHhahtMnqsJDffd16xBMrPtG/rTM
4AP01XUT/5Hl0GCBxyYaBlgXYuPU6hAednAAp7+RAhiOaHqHAiNKIHT7Rq1A9f60
k12cWYl8DV3FgqzwsBq1gUdgz4Pf40u7sy6vd90HdQguYLiHAjBZFvwP8hOKI8ZF
e2NAXL/cSQFnMZp2xDnl02k68kFjDgIEoAO6+iFuZ5LHi474QdKYhFKELkegUGvA
LJ4X1SXHwVwJPK7I86ZGLSX4yqRCGP5+ni+PxtnhsmK6roAGrd+NTC/9p7/Ik1lF
dAFdJtZ+D91P0tMWrkyvwhP3fPfA9/IYI9NyJejCuBG+AiUvwq+xCroYg94y2+VV
bs/ZD4SALhuMLbkV4OBJW93SWbiZUN7eSWFkLVCfnV4g2ypfSa9nqUyI7v5WN2ev
AflFClAsvLZcWx22LELOED/1jvAc3B/thxDlBMsk4aHAiLbfNhgyPLh26uvaeAPm
aZk6FvFDZD4bsbl+mfxqCGHiKwTK1ogpN65+r5rW83QACF+Vuw7J3zWDjCUDEhPJ
rhvQ6rBfjAZw761aPwb4Va637RNAfawLmZXqe5vEYHyycBoUH+8QdwSkBkouv+Dp
2FxWIvEcyShJ0Jd+Dlgpioa2OIn8M8FzEQ8T82wPrHqyByNYZur0m8dW7XEZUypV
Ybr1AGrUlnMU9PzwjJs4l38RTFYn+P41E3LifRorui7KdhV2seqYZ0eRZkV35XRi
n/dfnevHeNuebfallXsyqb4u+u49A8Q8MgSO4gQhP+WMlqy4QtUqNcHxnuKiLD7e
6rIsR49/bEWcxbWDIRuaS2hbdWp+xZwETxK3C8hbgyAc26UPuTRQAfq0dlmSnjnn
EDLZPDUQ7LrG23F+i9G4EhdXaF28osKaFtWcVL//KO5F3qfesnBOA/2DvWQ70gWA
jwwIoDCevlrU9rpSRRansuSqDyhFpYjPZmPWGSf66tiqVQgdjh4Kx2ELiNntfYy2
xiaupXSvxfql8HhnnTdb8wc5DxCU7eHOkCp+QuJMIZPAWcmq3lJfH+tvvbM+EJk0
q1ASzLllC+Qiel/WSu38cTtP+mxODSdLS9cnJ1PzixtIz6VdjAGqdWh8SPLmlljr
oqpOGBcwHJeXRrAPy01ykilEv9rJLrmjOAwYG9U7+C3ZFtpI6uTPR6KXyn40FEw1
6+pju5Q2pBerXfJ9EdgAW4zxinoxmtz1uJ8twBM9r82lUMMVS5f31UHADiRGw/y8
o++GRcXWg6zZLJTtFB2t3hlC6u5DyGpSEXaTmn5OD4Dc2BmgPX4JEZ/4/dxDQEPm
Hz9MmieCgIyXUKt5q7kkJAmen+jVoIYbPgWrec95rwxB8NJAn7miP69rZt1hT+4z
gbhnxnZLHAOGdSqSKbjzNQyNYaoZT/Dj4XJtWAVWaCyS0+ZZlgvgZXjAHJmVs8kz
sD8g9UgGyQwJ+u+aZgBH0dVVOgs1Hpl5M7rQB34ZtWA51d1+QyObREPEEP9h6Fmg
QHMRqGMin3A06j7puGI6d/zSMkOstxpziytj8mfaNaMOu/t2cLFK990TDNEml7PV
MunppkLalWkXUy9/yIWndhvPsYcPjhoQ5MNKoXYGSCZBd0t58So0fHfPF3khibuU
kZtVSWiajkYmXVYOLFIKRheGvLRC6lEha9KQ62tIe+ssxfkPL6Igga6XGGHZ7kjs
TBBRYo+xt+65fB1r6N6YGhUU7HG9izxF4XkE4wWUJiZBMC7pzQzTiNOFRXrS+Z18
Eh9QZrfv+kDUGfetYIqLPpFcwnxdHTK7kEyzM0DbwXoiZnOtZBWt1A3gN9sjmOxi
`protect END_PROTECTED
