`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZlInbiR/5Cow3XGJWzx6V/320TYhCCQz1QKXwB+u6QFNP60iwTQtp+gTc+g0yuct
Ud7fcGeY4WteA9O0IuhKJgiaAfBevFGvxTOx5InnG1hUc2IciahIJmoNAOk9EkBa
pDmSVqnb2bIIV8fuViq2evhedCZZWUiVw48r/6PxUlaNSv8pCqBqer3+vtBStcl7
twEsoZFATzJ3oc1ThwSESCWpbm716FpUNkI4hVru8tcSPvkLbmdDVY2zNaSRCvT+
/8cvbF9EmvYvQm9GyiDuBFlmKQsIEw2TRNZ35ayI7KdjyTbZSc28iHRvABsBCdUJ
oUpeXnZZlhtoH24ZTrKt4odXwhDvA95CR//CMQoD2E19hQu35QYVffyUG271pr1Y
lyjMTseb7MvO5WN1OnSpX99JvjIx0esuoIdN1IIT2JN6U5TA48HmFmEpfJViECkW
n/SbShoAgSt7rqyqjhBHSSIN1oA79nfIKuMI2fz/vRfYIKnrYq3uxN8m5XIsyIED
o5bXckphZBTia9XW0ckH2kjB/wxXW4EFESZzyxEPKUCn98ZsM/98ggH6mRLxWs/V
h6+/jQeAdpRZb/HnGY5Azj5NLYlQYNoqSasVjWFeY7y4Pc6si78y29Wnxgu/XoSW
wIeiAMdjt0Ls1jHUGgf1Gn8ioJlUEWc3OpXiF/7FyI/3lBPiZATXXb99WeLbl0lI
xfeGZVBHbPcttdfApTH8Lh7dn/AXqk3Ex3IqXBfbdwoB2mgtq78HEP9+N4Eh+AIO
Ms6HkOK1rxIuFafx7AGJNTnN606hom0re1GCIfiKL5VZYVXwjgHHxiwoPNzfWakT
SGJ160FhMXu1kwGdDM3Z5mnzjVVk52iWJscRN5iw/SGIcZ+GBk1yIhostd1eyMfi
Kpl9aDJpxHFMOApHxzImCrqPuQgLl5BhM9dElzl7np1lAucD1Si7phhgeZmRfIQl
bBX/dNZMLYUYMmE86IEtu2bdj1IyqjrGwkK7tKa71NLgTTuHncZXxMkUeomKYT13
IKPzUsSWa9Bhrqhm5zQMOeFw14Wl/HgZbGSDi87w+/lEoIwk43YodmeBuQdnJPZ8
41wzJn5Lo/5m+FHSD7un30w+fWMtUt/okv82wJbl0lT0Oig+19LF9S7xV+5x1mTi
nEnLU2jECSpEjuRe5TUDWgHweUJrh5JoEBNAaeuaDlVoSKnhVxQPspAYsFIXx6YF
0yVr1mv1ihVMUWCoikxN9aUKuJd9Pvub4gEjivrWQJruNjnhzYMe5M/b/EZ4pN70
t4c5ER0G60a62efFe4dqJXlPUlP5p3grLTAdrIl1Rm8SM7yH92psiEkWv0iUjU4Q
kr7KEcq1htGmtuRpqwLjxeqshEdj06t1S7cQD+hJtC2yeRSjAbwyixTHPBw2o/9h
/53iivQ0v5NlJC/Wq2okyJ/LsQtlpqWYP1XuunBHaSNe9QtbHorW+o4e4G7KWuC+
V6RwQ7yT8Us54nHocUzMVy8kP3V69MReQ3vn75Nqbi6qWZ775mrgSpVwMdlVeT6C
s+kcdzvtYTE96whIQKgmHCsUrnrtSZMpxjeCeC8AHiNCPH7gfD/K9+mg/4GqtjuT
z5ecvN2ha1kJ+vXm6oMJZRNqMPyIkNxQEij6Ok1IyPUW3mqlQohEAH4vCrs/30DO
xvr9ZKyWziqA2Mnq2I6bIgD74P6G6IXyCk8mnH5Nb1S1b3p2L2Yi5AS1VqgMBp9U
8AUbMBn8NcfSMG5fn8QipRdKe1G8InLCE2Z0aa19H4dgNfdoAGKB/cFBlMVfJq1V
mL+sfA7WCmEnASJgfKRSfxsF26B0YxvM1GV5HVZsYTN1fOVWpotvcx/AkiF0/uwT
zojYDw4SqhBpCGulG0KpJ0n4Jur0nqHTY1dQKWErFyZfmAuwEqqU2Fz8WuxzlmWT
Pvi6rdma5JW/YW1yDwrqNvTIOwoJivOIBEp8rSK7RhrcT+Yw7lQcZdg5HVd3rhhc
1dt2s4qZHS8WS3W08CgRo+FHhPt9At/86jYq/s+6+oaWDUYLn0xVQWPfMZztSUXT
Pw4D+q5rCpcsquxCCjOc0VfZBUonUPzOLsh3HSP37depHa3z+rhYqQr67fkdBWe7
k65PaRBc47BvhXE7NcN0mcM8J8JAJlxvH/p5IEnm3BexpcmifwUiTy/hVuKaQTf+
fGZQ3U96mqfbgJxz22SgcXiytTNGsL6aE/FDHjHvwgn3GPHdW73Wtmnyn5AIADan
KmxXO9fGg+WM+1ZMaLcfjWq7noSbpiu6ns3oWNYLWrpfyzm3Ak96+CmwJRIQ9b90
ic7bZfOypm6+DEcHF/JUe+FqbAJ67UFbSfQLbOUDlIrATDuPiMRusy3bE2HivK1M
/1ImYSxRBzPgQROc9XHkWAESPLV+DRmjcL5zNvORpk5Pp187/M/Qu8sXqhdKop3A
/Kz9N8X4IyUHv7nG/zRyBvNG5IA+hFQyZsLWReGEmgZFTz7VaBbkAldQ3qDdJ5Uy
Qr3jcMs5D8sOml/iSxenUNJtozuS/iiqLV6USXnoPShQhtTuMK1DJKMY+FVrVnM5
RM3jxnX2GCEue1ZBDun1NaFVze03ZbW/6a42j3ptrPl6VlPEBHAJG6I/Odj1OOUQ
G5KMud3lwtqpDWTaTnYZCo8C7VLj0BWUbW2ugPelOZ1HhhSINrVAze8iEaiiJaW+
j2Y7nx0V5x6tGr8m8QXcyOw5DERfMNBgK6MHKz9mDRBKVtJQwUat54/iF/Ps0MEb
bss5NdMXOParqF1e9krAsvDzYHEGDUnGCgP4RSHD+xP6mNGTVjtINItwVvYeWLSu
ZCp3u0bkxq6QrjbX9ObOZaC7uSj20uZUAUZo+ULpDJJCWCTNhUaGs1xc5Nt8pBIg
y/vjNYyBZJe+I/EqLSX7+/inQM2SdBhOam/rjDnxpllrCG1OGHI4+tR3r4LpkqLz
d2ZwE4gTEQzGQlgquvoP33e1HqK77/cQDC+xhw9Kb0AWUMkBQNxU3/7uiU6Y2x5M
e4n6LQOrGipRBCrMJd0QS6k4rr0J5r+6+3aB36eutgD6A519mcdy0aMjva/ukPlO
wpBmPOJMlygutmEUKhJZ+9/DHC76DXonxpwJbcuWgz5NwD6zNeBYIUABxgrAkHF4
we4NzW+y+umKtBiaFFkwIZ9fMhNjRE6zqYFFhYCkuvLPZStFfMw65ssivxoILLSr
3aIfl8zdhvvSGloYOeXXKWK9sxnVFaX20F9IxIb8PqYQYTBnN7ccop2YAyjxYMVz
PF+mp6Z74O+5bcUf/RuJk6h5fkKdzqsW6Oy2WF5tEDLIJXsGMiLVJJpx9wOaz3aP
2lRYmK0UtTM99G3/4Xq9SIzmXey/Pq/XxuqXN1fHxALXbiShZswYwJ6wSdnNyaml
Sr5eJo1S8+9IrlGfsPMUbmqRGkrjk/uuCvofnS5u2+iNO/XZ/x26Vmbc2zZ+BvJe
SxdffH/lvOIjOF3DrqGA3owtQ36dIM0n2vZzSNYy9oyC2Q0oXANTqfcV3XqpUXdU
6q6cCIYG4Ijaji/yjrdttrV8ueFMLbnZo38mty6CTePQbLaawNJz1T+jsfXGBba0
o5LPeOD4YGbkBihrSRa6nkrUCamAybJdosqmhqQGjDOvr68jsWbsHNAXqVDjceuH
+giZA6PQ+iZIYa4n5hTpnk3nuVcbSfziXu83zGFWkLROyOk0AK1Coo64cbC9gK53
ZSTcdoQLH8tOnApf/Y9Q9JVkREntj/Fd32wlIlcctp/5aKIaYe3Qc8uhLE5X+f5U
1AY9bKKPqtJEqCcv5tbMGf3O2doNluerTFrwrtx3tr91tH5bXa+oEEh/aUnXqPj8
rhARVIoDK0Uw2E3GcA8bMjqtBbchosmKfoY+2W5ltutp+tJpK7ETER3NpULTBuqh
qUQWMpk7nwMoOU2jh4K0mPhkDqTreEx4l1QtFXh3poT5QFXTzesW7e7d4vyonGCs
GZLhjVz8eOLcqTQb2FyZtEEAl24ug3HXZ4KGR798uF5520yZWcIVC9oX91t8Pegi
CotLHL+IUkQyJDSYyqtyda99DYax3VhZ9PqGKfnR0ss4+1gv37GxoaYm/dQbsOFK
gEwE4UZkhwojBLtGOXxwaxs5t+HJjdJ3LKgEEM1HR3uNh4v2AORZNPh1ej+R1umG
tsCHEgHUomV701zcidC6afZjGoxHcT50yjTe6RW6zLNuu3xCDPCsbV5J9Fb9ZZS/
4KPXOwL8Cfl0LWTA+Uq9BQCqgz7mVHi0J3l6TT3UZJpoRwphS7KAHSEnm6PWP7Ct
TNO9wdZzCAE8TgLaEOgpBgsoTmyc+p5kQu1oKI670SfkVC1qC0BkL8M/DdWmrCwn
OnLp8HsRNlBq9eP2YYwukrbNTvQRdDq2Vxe4jju+TCmoC5M2r1vIkZ0/DnDKQoIL
qCR66lwShDIeJb66uSLNj3R8fXGgzDv2YTGYUevXQU7zILPGL63OyuCgxvmXfsd9
UOPhmd8XeZNG8kWvKrE3dLE8dEDaQlDtHeftPlUSlR4hu+h+yCzCsszd/FA84Ybr
GZXSmCcjYRkQICl9r9s/wuyW3Izy+HRJOy7AOnjkkHI5BMae5llEH1UiW2xxaYR5
r5l4C915Mx8fqH3eeWk6/Q==
`protect END_PROTECTED
