`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TPr2QS03iiKvOsU1O7Jow9htc48KXcYP+rLeDyjPRgYw6+EasiCYnKEE3DtoUxfT
s/eZQI4TixxR4pisHNz4lqJM156UzHYFGEsWumwcvqwZj9tjRdzJ5XKStieE0vr8
rHA/y0AdZ8Sn1kgJ19JypbBbPvTkIdVOSIy2m0KByoyferSkKXMXMFyf3b9+eCrC
lE6fBPPusqCiCk7aTdAERhHihmJxvrZFTsBzIsHJ7QGzX+wTi/OLnz/bnbhNxFDG
9znDZagUSZOUfe+eAbvVCFaQvT+ZOWKre3Kwew3z1gzsJ3gPDQsihz+DnAIVOQIc
Bdju18JDLDoX9aYI3mYXuFTT5axji2dYBOD4quk6O4buSvDE3EN+rDPB0ioCERK2
`protect END_PROTECTED
