`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VBySPPP50a4PrtpIjZ7oVN/VeRAXdcT2m1DpxOutI0Faei0JrzWS9u32P7Rt1jfK
JeqO5NfJAcmjXyjuGNdbp7L5fcZtsBu0QVUjaUrTk/28qZHZEZMs/LKrtkqx/WfZ
+uSePzwsL29+VJd2zgxM0Ry64ccqnYcrUZYle02JPw6UyxlIW7Euo7EcaxPF05mV
iSmaGkGJ9YXuHx3BWaVAdCqOKzDutwMq9xRlGEqiqb7mwCiT7r6vzMSrpMBTiP2l
cKTbrfs9uFZkJ/kFUnI9ob0Tmj5U9JjbUyVp7GNhUsseds1jZsBCNgU0ojKb2soA
WMuD0aPUoKduTDuKj0DnJ9YqoaGy3DDpW+TkC7RUzY8dfnpbzPeQKIyo3/ftmjZF
dpLMpgXApd6MYTl4wzkE6x5CTM9giBK74yYcvZHvDT8i59TJi6FYuhp39W0nJITs
3ZYi17QeUOPd35fZ7jG5zPEpmoDvi9bLkF2JKxlw25Vfpccpo5I2w41rl5Dbb7VB
42aD2OYoUZ8ahTXtjUu/+MjBeZm1R+1wbDGAaBX+Sw94VFQn4NcGt2LkMmQrlk6F
brZwh0QtD/5ldaNdeQSxspQiPOxCnk3MGTR1CJLteer5kmxvTIOOCDy5OdgMrGCU
UMeeIuAx65ZcVOpMO1w6mtpreX9atDgarFy7q9S5shTrcqTOPbyFb5HF+AQRFc9p
NhmnwTP6aQWDUXIqWmJhiRq+IT5A4MJVadD3yOm/kycYZ11ERZfpxV08wBf30B4+
piiJAbz5Z8LreZ4hInzqxtYfW8Y8sI/Qu0J++t9tYSnmxTP7zDdWm2ZPBvdmJ0aE
r+eR5nWt/nN1TftBVjNRgxZFdOHtO09Nimna4eIEdndGs0DgfaATFjX7EGBWdP8d
e1wvdylFQKNAgEfgnbgXjPrdUiiIC5k6d77E6giqJU1KfDR9/SuYGZsjU9Gahoqm
`protect END_PROTECTED
