`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QVNDRfk5AHl6ictfrJgBBHHaSJlTqYOe5HekvThrc246bdU2QPPWyVZJIUKptVgM
wMgpyBbvX9SRFtpgspPMsMRHNxNodY2sd5xDhPeRg4D+x0fdKqPL0N68waLKfa/F
MfhzLjiTKTwOvGdPBZrf173xscDxtF/njztfBI5QvZRUqKBN8wegLZ3ZwNctfsSy
ni9xqi7Zt+f7ZHz4f4B0F9IbrkIPxw2PoAehwmpESpqH9y+N+pHSo58BkFez2WxF
7CHWG/mxrHkkjGr2GEjU3E9tPRMw2yIFzgtiHE1rVCJqjHwUJNmKEZy6G+u6W4yp
0/AbGhv0Syx4TuUY7VPiKVNZY+CMLTa6YlPACwcZ++gGzhSay8aeKMAf0NuCvhV/
FyzqDhdj1sgGqK1DhKAZqDzo6Yc+G1Uu2H6xMvHnB/MvZluLyNM0fMrvnCdatjCl
Rp/ID1UaKCBZ9lOcNpRT/721hAvgIIScsmNWnOROpj5YMgNBxYfihQYTJbvFHnx0
JuHFSSU2q3Z1IaTbMirr9Ne9dfBpMo31uMWEF2qlc62DqFQ+YNloqnl78r6wryFN
dWIBLEt3gtsdfgP81FoQN9FSyji0l/xviu4ASYmdC9YDCP+bJ865or15CePT02po
sVaENl0SkYYBIhDSRGt4FYcrrjpFsVaRqehhDL35l0JWgMp60VpCkUkivwJHGDvJ
nreOFDxKnAuCp4OtvkMqKKxYzcXJgiXqhN7VPJ/2cPv9ylT7D/B40XDWM4iTJiwd
nm7Haz4Jcqy763D5c6+K7JhipfyoNK5Hs9L/gbjIe319UmvU+1aDht2ytM2QZKRw
ijyqnOgQw7BL6Ts9j75CbifZhcuizJ9tN52IaCMW5H9USKkC322lTefWc7HZ0lsB
8455SGuDK16YFPBbLSck9+wBs5HRrHeNWqhY/EYJgmMlbIsYWTYvqUAQVDIK9efu
MM9bSVcrVMwV+w51AAafqBePEd681OiSdG4CHmQSFn93etmT91jB6wYOAeUkFkDq
`protect END_PROTECTED
