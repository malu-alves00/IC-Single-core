`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VPgbRsGLG+nWA91tL58D/sBQ3DyPTLf1Oo0XXlCQdcuJsU3fWhKp8lah43/f/aB2
zklPYZsMQCObvoB8gHOVhvO5OrCEewDb4oE0KK7UGnuoJXngCNAZCkcdBvdnrgyZ
H80TfxN8R2Ha/x0eQGJ4DfS4T/vwy1dAJ2GicgwB507vQktL/25GZiAfuRwvv7Hn
dVr+n6Uz93Va2eXzXGFHXSxD6EOB6czs+duSISn100TyARHfzba+tIotHaQ8tszw
t9h0fGfmk6alowap6cIANFzUWHngxqV0KK+6j2aWmgROjyVuKD6xHhGZR6ob7WFN
pJyZ+zt2iHVwlIYSw/KNA2bVhLckhClz9LXLbuuxlbMkb+HUcdMPPYJwnPPz2q98
knRDgOMF52CfPspBkkgzzAYFSctFcUdYWVLgzhlbLOE7ExPk9nWq+MAoiU/SR9Uw
eb6jP6u9tPjR5h1w8l8oVZ2wboLal4NpK1uiyazCyyjZLsVzTWj4h3kbJkjuCyoW
EX8R4W2LACRZJ4rGzJ7583Hh7sTFaB4Mc0T7qcCIwpDwICJqjxHef4R/FaEiThhU
SBVAz0aLFeOZjRG+cSF+ToaGTj67e7fJFuLLND94vgksjCVB8Jmkp/JE0K6W3WqT
K5OA3w4N/N+RXbdJUnB+55gCL6B5oY2m+87EiOmpqaAMEJImkeaNEHnKdU9/ULFs
dVId2RKTtNEEt9LuMg9VMK9K3yqGSRITM+yuzMY+ZzQJl/spmGMy34OrRt5bnedk
m290XupI/03n/dDDmbejYNVOjDwrJNrK2qj1QMuUsvO4xii4QLuZ7yPoWjBPRGc2
s7UhRWYu6fAgDC86daidyXgpj9ZbdCOXQVetWyCfCQXkyB86V5aSHLy8W+xyGAhQ
UfX7XyNTOy+oM3Ya/HZ3UlAbpEpinxqFm7+httR/1eCc/TCGvCM4vy2GWwflAcwQ
jsYFE6zeJD/7p0n1CJdLxuoE+GJSFq9P4qusFM6SYlM6Sw2RRR9fWgvHux1Iud+N
9yZntKv00tyV6pDcypEnKqwiE+WIh1h6r+vhDbKYrZO6bkJDoyNZwEKL1cVEOqbt
oc55ZIKIGUCEbPY4Goy/Egg0ed3dqIMABl5NGD3bfW0KMfL7AE8+hQYvQ5XaY9aC
+MxX/uLp/+tWlHvmsJHKUiUC85RinwO95YWdxMbWPHQV3UFi2wZ8Ef0JXKTA7vu/
aW7XV0tHlSENw1pHLyrkMdRe4FuqaAeQ0ORwJ9mr8ALLSC+QsF/GEJxJJVaaAjKJ
ysYRm8mUraR3pwwwogt19ltP6Cc/7m8CSvvfFXekN/QkXauvyJG9nnNMfe7GFS2i
IBt5GrPqvk3Vw8O5Vs6ZExY7vutz/RXl10WWIkCmTZv7r2xFFJB2dJ0sGph/qEUe
7zG2luniGorK9eYZimvBG7tcAD1hiO+7yEXh6J6QT2OxrGmKDEgW3SZBawNpYHVw
`protect END_PROTECTED
