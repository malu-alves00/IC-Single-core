`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
chtv1NqruFF7Ut1o52sfDuhtBc4o+fDC63OnYpZaMhhaGPzPqNZxDdZhGNi2quqG
kVJNes7L5hyKqpJQ7LozTU6qQ5uMdaBBfqNNfOouOQ5cUFHdb5K5Jz4vVaXBeD+K
ZlMDS7zsKWXxPUh5v+IuuhR03amA1ROZ/zP8kBgzW4Tmc2eWmJ0q/zEAbOkbkkov
4mRmlqK3vCGibjiyTpK9mRDsl0g0Hzg2UlI88F7s8oWrIk+8GpuKPEHjjihZzK68
DnM247OdBW8O4C87uOnJ7RiR2GlX4waQXs36DwVWfv+dyZpxVj0xw1K9yWhlpdci
reiGw/8HZbfLoes8weZh48R4LrZ+BP+hCNWS9hI7AdExNbOuA81re13YQQ3lIPip
AGPqCWHuIIXhTn4VKuI4hiqdnCWxAXx8DPqhIuItRgsWMX0SahW9UaZeOg5AFGlc
cb3H4uDA5Hhi5qEL4dPjHuinSzdn+MpyZ2kkthT84i6cA3j9cFFJ9LC3wv5jjCp7
TQL66QeX9opNbweYwzkaw3bkRW8zaetzDejP49h7MUEq1+q2YBMKYTn69zM5kpad
cF+fJk3XkF+CCEy+CQdwVPdvxYyJ5uUdLS+edOzl60f0qf0NuvMitH99KjrW/aRW
nIillutywGp7iacAf8JGYLPYm+QFM0PnEeonlo6TlGSbXYnZmeQGAPC9Hx0AWJ8E
pflNy0FabWYoQn0xVmcChyxj7zsVjlGUTvg9WZAK9Bsv4n6OZay60eHrlsxR7DAz
z1/tY9ARaA3hrcThwcVdHOvJz8rcwuAZh2eJPb8LLYB5OyK5T5sS352piHp6alZ9
rCpXDBwk15V7fFkBCvH6d83fdyAAP7kgfXulxl5dUlkaOIH4nStBTtt+1UMaYliG
Md2shqD6AFQ01MpV8/6RT0mjnoQIVMgEtDK84c3QJTSD0NG5dHCZy9psKzT5u0pE
Xvc8mucN08LRkdjlTTN2hwbf0owtxHioDUyfS9PzYKzsHg4UfnpWY5Xe+X5eQfBz
Swb0qqARRJLel6o0SllqDjfijDLiKr/iYcZPjErvNdD7EbwsEyP6yAY9/i8RM/mc
w+2c2k2t/W4mfoOqR1TuCer+w5W2MZqCumx1nCvGf5C4zljcuuEsTHOw2XZgdLDO
95ntBKmYhfJtSbp2JnQTKAloMpRQImCTe19619mJ8RW2zId8ZVnrdtoBypKT5D06
OksZVGrJO5qLeFgm20L4FRApxGXXBAZdi/fzgNRM1bQebEPOFAaImDpHbEMFIp9p
d66n1TyP4zaFWg9qDNVczHuduBCvLPAX2Oxn1mDZ/vUSo7DnMGv51wbtr0Kdavyq
vMOXjGm/WLIFmYywjNouZ2hKKml4AktBGYZv3J2GZ5fQW1iZpjsGYp1l/77H6Hp8
IKyjqANVdMB0yyiXrHzkY4Q8g9DS7YM8UkklhQ013QZGXYze/jr/n964VueRxJ6f
c0X9V4aEqIz7QEvAm0QOqMfZ6eYv8tP5Madl/I7JMFrSnLgSQpWDXHr0vALb07ZU
lfqkewovypSyk+MQbpdVDjC9OO4cQpcN+cRwMujdGFZK2BZ9cRQ9yUfWI8tNkdf3
OuGVoku93/LI7qM+75jmq4dhzijPCGVf2cSiqlqozMgXUB4OCM3telZHaizJJ4mv
1FgpbVRzrmKDCT80G8nSR5fcpl8p1Rqt8B1G0vk9p9EUQv6QTDR+X8dpWYztKlkg
qncMZjuHEU9Ob8LRnjdqzp2tF3TeGGBo6kmGOJylCF4PwGb+FcyJR0gMjRc+gwTS
qL2X18NQztxHDf9oyMygNnJBzDeODqNbv+B7AQG0IICrCH4hIg5F36qq470h7ZPE
VFd0hTXVlgnO5NTWkhp06wpEAVkUGRfYAIZJGLAswkOlUomnLWexCR0i0xHaq1b7
mGZZYQKDLQnwU/FgEQrYTkfRorl1a9pxnvJXe047nXkNe9t17PehNQ8vD8rMdQFq
ImCC2T4qA34MvS0V8/Vrt/W1rnV9jGDc3C3Ynkmpk6R02Agu6qBqGya6JZpjscZV
iwDBk+p90o0hLZ1APes9HE5ax2u+Uwm1RMzy1WH1evETysqWq5T6jzrt6UVpBI/l
g2R5Blc58uqqBFp0m2ZcmxyT2O3rjvpwa4UxrKkGsryX6jez5Qf92WXxIhiMPSPv
J8q8UwkTJkJ7iwp9EictcGoypYfq6Gc/jjblclqB5I5ax3tP7LzpLiuQE2XZoJt0
7eHE9hBTiDb5tAD0NR1hjoOACHupcnZaW4+7+DbG/9k3vGQu/nX1HrEWIq0hiOHN
4Zuwz4nI5kDhDplRg/oLkK+XgbicSGPs+PWqrWJyiWvehRE0W3XwBqWJjFIS99DT
VchT+hym9W3TXKIs+rmdOcICg4ShSo7WQ+RXIWq6ujDAOvGNs/7eJ3DYTUdsUjVT
kCf+oii5suUw4asjhrhLEII2ECwNB0Ssq7xi38Dm6QeQ9zzw4KzC9oe73hv4NIX+
hJQzJ4Gpfl6Ys3gvebdW49ydZlT8EqiZgjVqSCMw9pgu5JgfSXTT8SfgOPTy9jdz
ghXlaH+JkV+tKsqh3iKVLHTvuajX4eEvhaOFrkfK08D5gmIcm4UWDWyxE34W9eM6
/fu+Ik5Ya0HBfrNnu7Bk6aN9q10evTlEP7x4t4QCxaSIuMnWzEBkrwKC6XQ6g0cW
3hujUN4iHwSDsrOOjHQYaA+XOWmW4+q1HpTHCvo+XS4P2G/W/2egJ88qme+pFsvV
0R18byVAHwVeEW9NsgfY/ulvJddbfN5XUB6xQkOlxjLhPotwYFjbvHXUKE2UjT3W
A9pvNGpOr44m4B6sm0TaaohDGXWseKyh9T+L01j5+kor8YFI7QLLoShDsol4b2b4
zfIjfZbAi09bL9YtbeAjAe3ZL0Al9V7WJXrRB3YG558XRKv4FYsyaHuV1jEmuRji
yMepfSvtxhZ3OFFqctUKubhSPLF+biQYTbS/AbFWlAnD4e3HSFGMSZCoAfpvbFUb
ct8kbWe7M9C3gF7D+25No2jcNLnaSbC1a80yoVweo1qpML+hiMOl/3OA5WILm9id
v2DH/JYWpfRO3gumRcmUOaiHqs7arBj/EO/aGRJI8AiQFLblOND7zKN3iE9Do1Fx
xZYc82PI63MMOnBKT6qhKmQ0DE59RNpDnc5BNuF2ooeMrQCRWfzbromcbuVFMDlW
MVy4rYyEAng1qZhNwbOidRWtzK14HmvV4jktqGaOzAP1zVhuDKQQl+LD5viym3sJ
cEliVx07mSw9EEpImwN6qjloNAmumx2Nysod+xB5hRMTS1wvYYRnPM5yooBqDTHt
voKDSRGthIKWno2IBxFPTfHOygRJo+HAkoTUtpZ7+PI2rNV9+DH/FBBOoo0vqqeh
SF9Xwy3CVzNX4BBtyARznKNd63dicSc+JEVL2A7wb1PXjA8gZ4PCrjsBYQyr43LI
LyCPWreVVcVR5Zjm7cSVMDRs6FKTJdJoqUVoIrZdxKtJqtsu7ERuVqSknMKWe/DX
p8rciDs3u14RjVtPb/ZmqmrIBzhEqtB7Pp1Q1M0rZ2WJYTn+QfJKs+XfitOxHO+J
ncuFioqR3l0vpUGGFqP+GBfbHgtMCjgTAp+njCGRJX3XZIQagBH0fFlQrwq6L26Z
jukzp2IK/VnLjaFctFuI+bKxkgr4IT6NhP0ILO6bWX1uEGDnHaeIQX3yjKVaM8T+
zqsSCPo/2yRkD1LSneUN5KiMVgO+99yUxdgF36VT1Dui5kNorI01ICiAOyTTtf1A
7K52TMWGhhOT4adusQZO/FTWuuGpMHZKfC5CPusvemY3sJ++WLeNn4VkzKPYvRvZ
X0jaHlaY6yD1arw+R3xF6sX6GBw6YyYL6i50+l8Jxt2I11sqMNNaoCEuc3pnhYYt
8FqnSPjo3VAVeN9Pf4GLjUWRrBk4vHQXAuTr8NgnzRdjC1Lc+2xZexirz8n00hGk
emDVmDF03DvY1a0g4F/oY5RyUmtgEgExQFw9CdTOAC29ad+jh693oKWT0CvrqT4Z
M4xEpX1LgrogvIl09jSdDe4lF/1s9jAx59D5YSrqtnJNI2adFczl4n84zhRFV3vG
QGk2CmEDxGDR94DhqjvcHFq/9CnpoLkEfZozQVgmYWOtSLe7dVnuCi0FrCa7BZvj
LuTvWY0q1YcLR5lh2SLWUvmbTLaboIHxi/fxTyIU2Htj5P+LD7xvOPQX6kJlvw0v
a/FgwC/vHoDFoUatNvrjGgjCovHm8YxkkHn3FvSE+2rcWAbNRiu1AtUkw0My/5Ko
v+iHXkMfMB5Z0DE3BUhY3yj/r0Ro89RNq8orGXsH4gtpxmTDg981jX+08dgf3wPR
x0j1mw0QVCfdmZHCDFwdK3S2J9L0rfXdb7YyCePm5K8FncixyHtraLwrWuwDLsMR
DD2wLYL9JOeQ2Ef10AXhn6FGOdHkSDPLkfImhMJokJswDr+TmPWjFIfWI7GNu7Ov
u9ZNPswi1gPWZWGmTwjVpfdtDiMRvIZA9bfrmm30olCcb9zIO0hw8CCDszfZGYbL
CsIHBujSev6S28iq9eFBSfinVCLAX5hj+TNJ+Rzd3pydnfU07bYbke6ZjoKhavHL
4uidW4y8q1tVyrKITIUNT1R6KQKbRJfFyP6tlQc6KGUVlI2r6wq4/n4xnnh4ldHX
acjkA54MJ95EAWsj0Sr0ot9wDrBb4RPz643wpmW6TLdIWEPe63SCLnGxN0BoDOuy
b3GEvHqoj6BkAi3PxRuC2wklcCNkmLo02wne+CPhOZUFVDDF6AReQFq1HrwXlrd/
kUQu+1en/JiWikIow2pe5YQtbVTNf5+vxrRa7BgYxP41AYPrAnVzI2ftr+mHbmMA
6hzt5AHHn/ZdlC/txdgRWyyFj4HPy92TeQFpt1Q0nExDSesBK/XXObFa/yU5R3t5
7WumFCw1tMZnEKOv3DQPrax/G70ua0UZ6l4UwZyPI0eTaGNC5PGYWuMnDh0mx3Nk
kR8eKmDlrxtFU9QRGFu7horNBoZMXD3lD37bA7zusA9dbceKOLPSiXYtA7EYVV+w
LdM+nwKIt4UeSGniORsJElaU0ZD/dZ+gu7srsXHmotw6lHcJ6eAH4yLP7psq4I11
ZP2QmSniRcQUwsh4akpeB7ONbz+3Agk42IbPkTWvPnEUXBYsgc9igqJ4FDM02aa/
o5u7KHTjCzGMKBRA86MXY6xo0oFhEuaYTZ9FXV/x6VKl2c6kLdTYqKvLIP5OAwIL
RIwR39HBBd3PNkgJzHneinEZCFQvS3+6rmZhLaRJJh+8Jo2BmjUY0Au27rq7IUV0
WXibRCJS3A/4IhCFZB0sWWzfmCBtyorJ0o3xj+2s5/sAAHP2XjMvoNXuqywpdln2
PqFBpO4q+hyyOZxFclu0qVLldxBiJnqsf4Sb/FG8bWckTWj5radPHJskAyqyxn0V
MA+S9GZtazUPwKkqktUEY2eqochOL/th5nIR++5ydvLFJwelxwfnubBoyxwhTwKm
icH65Iixfit4bogPdB49TfyKxzJp4iYkozQyaLBQtmitfASDYbCYthynFIr5WQG3
q1WWLmSqohrJ6kie8bExIFE/iCbh2AYqfpn97MRXEWnmS7uTRpV6Tb6gGxzBURMW
JOuQE5MP3uUffG4zGM9voFO6dybIEovUpzO8JxHFj7ovN7rg6w45GT+056tTuhLI
waTWAQTXFYbJHhoyC6e6NDfN0GIIGsSBdbV5kdrVYJUEJA7BEVlj22NxHW/9oi0Y
6xL6iHW+kj5HG0vHxAta9/0sJZ/9o+ijOmtRmky0d0HZ1V1c4DOAWs/1f7NNHc8I
ZTyk2EazME9rCJxoH0rXn+IKS9ceoo6xVXDqA1s/yth7ZlJLgaAmMWgFrzZI3Ve8
FEarED+81kzmF5bRH4M9Wu0q0ttQ34UC5RsM8gNUhyMXIB3RgzQYVAOQBtED1icX
CdUbokFCjny5JXBwhwng2RxNR4b0jawj0Rer0605bsut9NsNSfUnQfF5UNkOrrI4
KiOhZQ/c/Mhha/AWl3IzUGNvrmgSA0TtLJO/ZTbePE9OLhInVLikAotS40maHJwb
WgHpJ6CI709TmW6mLhVp2vMS7jKTi8dOKXh3ZVSEWoACx6UDR9Pi+k6prbUyvYXQ
sKI6NHGIt31wxIwKiiT2M5u59xVEMVxszjRkxzSFc83CMZfNYhRBHR1f7oDXoKxM
8NvDWeNwlLeGSelVYzpPB/wWnczC/qvUl4s1PgeuQm+6myUSSFLG2R/C1dkna0Il
UwFOrKJtg5S3Ph0HWvyn02hqds2k0c/X0+nYjv2S/68Md++++pNGfxKl55siXpyz
Cqlmzi6iW7LKjy4AFD6Pp8pxQ3DP8RvhFVRllmt0867scjBguCxEm3pD1PaxtyDP
pX+2f6GmPhejmPJIULfyfWXgAakdLAQblj1WGKHvWf6LLqWTiyWSCDXEKZadx361
8rLtenv3js68QMk2a5MQx5azSwvXr+l5kxzfOHl7/crdf+b8xQ0YVt5YM3CjT/6U
+rr/dzxUg3eeC6Ov2SsCQAPghi2RD26B5YYIaCU7USVn6d81EJ1cSAq9CnZjs/sU
LVnUHgmcz7hqKuP5SRX9wONyFiPo1DSZMSLfjL1I0qwzP81XU36kIsMqNm2+VL5o
YBcW8wAlo9uKR1UbNGYb114gcK0OCEXjkAYJTDr9YpMlLfQeB/NRr0J5FRf1geQ3
hZWbEmMuPb93splQFNJk6o8hkG+cUyBhsXJznP/S/HOGTdHBmFKlDTsslW881rgu
FfS9InbQIOTMlFrYZ5Q7V5yt0CYOJRXSwXxIbPLI0Cm2HOeaOE11R9nIYJ4l+nFd
iEHHnMpvNauXsK7e6kxXMXrKajFmOkP3oddwGTa00QU12HHq5C2i026uncFypebS
e/IlWOzlWMARyZkBtfxJ5udtYHV7ug+1A5zqVZNjbW6Xfp6TUy/j4cgscSwUZ5nf
aXF/htQoNZwfwjTAZsLlpBI9Hv06WN5ItKM+UfxJQY+B4akAWS/IrLSUX3xRIZaJ
lvjf1X235JbQPiHoD4B+10cXgbS7WZHoB+NcUXUUSL2mIbvHJY2al/8p9azZl1MW
to9Q4lFTJ+3VmOWR+OnDNzqiN8pqyN6lPZZ+Ca3Aif6vSbuIqiIbItHac0mEaxF/
YayhJZsF7EmQKpwvvYKjMJqcrjfdU80jqjiJfyo1mp0IPVBO/gjOJ9Uuf0pFEDl7
rdAIRm4LPA7YB8ApEO8Fv1nE9iv4F9j033BCMuB3nulw4krD0D8Ph+OcP3qyg4ur
0RWHQzp0r6nuUX1+pWOehLzhj2X1i00GM+spFXIfmrm6I5lvDDMf3sYYYMY0rOcI
OXRljUBhc2ZdUrfHrP9OuaH/LhtfuXXgFqJaE1hld9Uh3MURykx9zivitypOll8F
HIh8/DlDgMCxDA6z8iFQAOcFPK2SGWmQHLZ4D4+8XoVQYywVw/6txmMtkU85YszV
Ck7V7Ou3UeHny6C5lyeIirBe5eJ1x885FO1s15HDwedfHYHI0jlvIsQKArGaxvtd
oEsTrV0qbveyl4eZTCDYLGzC5q7Ku5cDe711Xqc9UhOkTsed8xHof5iDbP4otXzx
1Cr8gS353j6n4AqgxWbqcd7IPPzMtq1A2pAUX71gzvhUeIgOaYsx+TgDW+F1TRi+
QEwpGsc7SKTVL4j37HrQFrXeWq7DLmdA3YsXzZ3BCpeV4bLY1ocuBoXGDEoNeI4g
et7Pk3V+Nrwpp7UG/xG6JSeONZSi7sZCWk/aOjxQZPjOROoBEycz/+uhQHLHy/aL
FsLWleK6nysTgmnUGg4ATI2gOO0bbLTUnffseOOd5Kjikl5WXswBJi0ZUG1GAaCw
KQBdL1oUlcpTinY8fv8nGjIL/8QTU/oNtRSdFecxP/LcDOCF8ZA+L1GDtU/INfZQ
QNsOLNW1hi69AjpmonzI7+ZUz6EpBmVom5FvNLmD7N4D8DhwVYZwHJAJ0vNNSlzY
oQUwPeyH+p2ctpdHMsf1savzRfv71X6npbssYTioSV8/22THrLAMa+y9vPxvHnpy
xhlbKtoOY+vSt4oneDjb9LteXDDqBjdB4p5zhK/Ef2gsWg21LrJda3rBTXFVy5ZU
tGeXJiZnVSADiL/WC0OFtHtt2FyT9OaBC0NLlthfFW+rcgr5aPtgAZWX2X4ZZ1fl
xIJ/U5IH844ECJLytdce0A1xhjGPnEazu6M6EZ74ejhaN5vt4lAel1IDMCwr1qV2
L8EmrG9NwERWTRKWfR8m80Iy1VDxOetiUxKsrmaHyKlAky0EiI2V5U+B91MigHNm
Rma2yYR0YPmTUaHjVAuJOJCMDk4SeMMvzFbMpv+mclJLjiZObKkgj+aY3OoZDSE1
tphpnFdRm0aQi/b6PbvJ9EhxTVxaC+IDrtqHW8tUWJNRQM7wEfcLD5BY4eTUXjKL
0onEvwud/VO8uKMstzrxJsc1X9eDA6pHGKtfGpozvrMOBzDYqqa+KG6timMEOSdp
sVin1twQOMj1ezd0ZiU+tWclDzhK2yc2VWBncT0UhTocBdY4Mi5teg/kZM4EXZc6
Df6XBOczqBumwUj9eSXONZb+k7CwoneHx3Cnr23nR2Ouy5nO533lCtc2kfkowc6P
JWNeu1woAKuje1qipEQmEKPify3sbEJ1BFIMwZCqrRSvZQdrwtl+QvIcWv2jK3bj
M1Q79WvZCB+cP9ZD/PRE4BRKI4Z97zVT8CwN8tJczzwprqCTANcsb+TgHgTAvYSk
vRB3ZJrwf9e3lFDXbkS/fQkGrh8heDGkzELJ/3jvhHPwomYJjL8LftkIWEXWEqYX
b7ujRpXU134A4mEiE8E31FRZSKqTDQexh0aTYYdawAKjmgXhBzLhLSdWtcIGi8Fm
cVTvriGv/Of0s5UMfGc9bDIbiIGJI/NLA1V46lXtfuj4ey6jC1JOmyy+h1FRnyRy
BvOxEhV7R9KulodUUqxRI20GhEQRt7ipftEiKz0U73hCLu0Uo7LPxMaLtaq/PTrP
Sj9RwmiBVj6Ebbg/JNBKgVJE1lWIsHisXhH/pFsqvceKgaeIpuHUmDSmOkeN1uPO
QkUEqCImH1pNn2pDSHIEVB2Xui9ytpbaxiQUxdS4hkR5ufxqJFQvgruqbO+ZfHqZ
2m8R1oCk4wxf90lp5qOROOSQCr697QBRE/iTboyUklqxTaKo4TlD5LRAy95RUeHw
+PKx86SyurwYH5qPqB+6G0ege+yUcyV8YQ7CN4ccUf53tqTTN78GMNhxSCmhSBzU
T5iYhfI0REneVZmDVogt37VkZJtxOQMajMCqVVtINi3VcBLk4jBBwCxmZGBO8Xf9
/ytP2W3bvJahDJrsN55LxX2IChkdmN80pB4TLaMjtdmrl7FuFB65DDsoUzt/0a5J
0pZdv5PgKQdKdCw8Dm7aJkv/kI4evUT/2LMCyFkcXOR2+a+Kkuwuy+JgfSPPgwUs
DcCRyRQ9zqqpA8C1b+My3spwPF5HK48G4IqCdOWWUCR7pxId3i4Gsi1Bu/k76bsb
gjoXldOG2OgdOzfFzlhFcAGtLUOONwauE5VXSHaYkYWwyEtEpjikdj9rNrdrfDKE
ayNUDJ/iu4hbWaoc9++aovtHkqxMwL0mkrVbn2vnMY/hYhlnA5rVkZHIhGVRlpgE
vA6dNehqZnLbtIlpf7woBNFLMYSEzWRxBjBgOvHsdtG3zR32WlIAptklEb0aTfcp
z8DYy6U3WgoSAz2yNwCj0V8mCUtYQwF4XweXMLa3hK9T6Bo3OLDyBiD3tf+xuRNZ
jTas49Awp9PMQ9Fr8gkSVqDL49zPA+ZjkIwK5j9E22j1IxzwszsAXQBe6Nl12PA0
dvu/9PJ2q8CQrcpApQS6xENg/TVxCVn8/lnVdfAZaMzoO1BiGqiUBAX7wrIN95P9
1B7sxfJ1daqKYoaTWLThD1pvr3jVdD2a8r+FwBUdF3ouChhAIGm+tbFybPGXoTsQ
Ft2zWwofFIHjjMUz2WvUAGq5k3gQzT2yrmUh7dEPHYoBp4Wv/bjFwRBwE2zcp2H+
3igwkXewEpus3KKD6qAD628grz5OWgYQgcVpQ8T+mTHVvH/RfNVFfLDvFX9DCvbU
DT+uEQp5E7Ubpl60uzv1r1svnMtcBcRMpRsStQ1Y6bIUjgXLDd9TcyezZ+4IwXu4
Y5W+9V0IRpZUm50KG+ifomz6UoSnLrWo4D1kjzXrvlT5MzTGSr71dajLdGkuKRqA
mhq5OMjEp4t1gWzcJQPNGBkEJXVARQ8YOut/APCwiL3xVoOzIucQbZ3lQ7L3OR/q
YHc5XRdv5m4Lf/Ghttpl6vCRYdiqYPZx9vo5wojs3WEgUSYFDxS1RpUTZr2YW/uF
NBuiWZXfn/5p7K+9mXvv1I0i+vEcOCO1ULtUeWFVulq3WB2GOXQvtfDqedlI9GJC
P32YQu/Cc7cwnrraLAqHqse7Z8r7qWIONMCXHqYiapzvkd2TVf11resX7Up9sCdp
TSyDSPxSXETyfdIoI2Fl7EQ06OH0eeWCtpcBqD481jemp7vtijGnmTXu1wLsPo9x
qAI6+MNzAZvqDmXwfWIkqGJ4o54TfOZf1c14mc8BwDUdul5W9zAfb5r++HxzmO1j
hZ2CnhxgG3gyV/4Vcv17WdBpdaAm/Z3RUvFh4AaVWZ+CJtuoT5ZEv18l0sadiL5j
mQvOCUKb7tHdczmHZpj5T2SeybopcsNU5GWb65iVUnh+e7VtANtqT3DA4pEj+2am
tDK122LoztbXzbpmdER+keUfu1E28wPpAKhlPZ4qnKU8EfQl+ilMNlR3dghRwUh3
vfwKrtJu6MYdPSCE4OJRsxN/g6dWx6TAYNfdTtq19lhwiRQF2H74obbImHvt7Im4
oU5X0IP3ASpFnTaxl4HniZItxvjcGSDSakCDww3cRb9davybV19SdglCMfHc7yYE
8SQoUux0haHBgLc2ojq5JY2EHY7f/ZJFq4wbT+HTNI0Y/KTCFxagmyfu0iT4XPWJ
80VKyrRFc3FuvRCphr/2VttBfMA6dmUMsLLRzVSH9AQPjXwd3+itAk4auF/C5vMU
rsLUzdxzVFGWgFAgGzKuRg6nqG3t5TCakBu5DHDvFPfJC3paKy8oyt8mQOv/9nYA
6UvGjF/J+69Kq2OVAdpXGbaJNfSyHTF99lc750NMA38xppYuEOrxjJrSbs5v3lgN
EGKSX/N0NUkYiET4FedDfmeDBPaWcF1RAqOu9va26HMSkVMRKXsg+s0OO0e5hZH+
Be8HyyDKiQ/zAl253WZlGRU7Bvm1cZf7udiu81/6NThqmvky9x8YRzAU4NUIMWQ7
9Alj1Q4Uzqdjfl+l0U9+gZhe3waX53crhaSSDzmXleHUCMVanvACho32AW09Ojuu
TLhyNJW04EWMH6DO2G92m3XMIEuBULDVvejVGnuvysr4OFijTtstyxs0CsTOb3Xw
0UoYQd1h13QRZJ5g9hT25W5YDTJnhZHTFKc+j15omTvnO4Hm3k9ctW8i3jMgQTZv
uZ7yrTgsaZ0sgCMDg5K+pbtR91gWNBqW3DIvfVpPlPoiMQXZcd71GQKTqDZr55YG
n85O0w9KXEFbfOLlkP73GZkLsY76p8bxPQZITuCWUU5T6fezVMVJyz5vcTWGIW0w
hqe9QsphQE9LZIKiNjBfiovpu+m1t+picLcodipHE6nc46l5zTVIHiWddtM9aebK
H9fPWyb1dA+7xkd71N8Cc5jy7NFKShNIKIYO6aGs6PG7lyQws4OLpKEyKfBwKRzV
ReJp9hKQnNZd7oOnr1gl119NxTkUTch25W0qxlJuRItYIRfE/AnZHAFbvbg//HUA
RoiJBNhEBQIYi0yEFabhKyOLIm6/TZ8VI/7HFUd8NRDsQQHaFPod8zeWebQeke+t
xP95jSDap+OZQZoW+vOy+VuS3NHNTB6bkgPbdMyeFR7a4QotOKqlbBjw0aoIfvnp
KwwAnp7KkeS+Em5GtcUzFMIgZn3HvPwTuyD4De+WldzjIzArv+dfk4ve/eZdBFQg
u1/ioziM4Pqmiu+Z3pGpcNY4BZv8jlcp/CLuSls8XbquuUEfRtgTGevW4dS27cnp
CEPyGlL8dAYsMs0iuHugLiQLpIWFHS3dEuxFz33ngPf9h6uUEKHu/NxrDkLwNxQz
NM96o3sWsCEV6xUWh3cjalkLCtF74pvKGedyMmbpFfne4aQh38FzvPcJRQvtZaTV
8KKgRD6SDWhevNRjlKcyh+Ntskl0zlgVtOGMQc4/7WC9TjYYhn0I/yMMtB+YJUrG
lldDzAUt8LzM54NAE7bs35HD3RMohJEPk3+PB+ER8XAyUd5hKUzQU8aKAdISnRAG
OsHwfKKgSJuezrdrLYW6MmNdVCWoRhv6rKxSPodIZuhvYSN5VEv017W+Cx0DrVmP
hoxTgmMhpX3WRNhx7edszBQQSR3X8N4RHpLlaMsHKkhrTM0EWXEpHei9gNCOpSRw
WuWujXZxAg9nd0uqbeiuBz8z1irPfTLZYgNfAiNLmca6J91PjQOpcBVmLH/LPgkm
GHaOiTQrwMxKXNsZLV2HLWhJ/ei0UhzUHdrucviveKr430gF2Euvqc19o1uAMFyg
zmtM/MVaS/7/Zwrk1CLTrcOjvgwqrDXoU2GVKOv843mwA8Io/NxaMbNUk12iLLC/
WqFOTP1+cqA9H9gU99wQFeHrtGvuw402+Qd5l3Tv1H6peECPy/cz+BS5pgD/P22h
Nkdy74USrwyfiNBHgr3lLGFrA4jQ/SfPDCOoXjddvXnNHkeGj3Cgypq5sqR2s4vP
Vj1OaAGB8i+DieQaHstAyITfBwbbJWKspt1HuO5T1RTJFVN4D3K52QkW9NBqDrKV
boQH3YDG9cwD1SBvGy1UO+RMZMYlfVzkQufvhUKze/W29c/GkRHL9S6t+V6wh17E
0oCKwIu6xpzGlWOo5HHcv3Ha0hi3UsPqoRfttkcqy7+Z0C4NDDcqb6QE5HZXIaHu
fa6egD9xONFlkbmdE6ITBo2IpSayQ5+IIN5u9zQNWNNTGf0yj86B0QPa/da/wzWF
wRlPY6MCzXImF+EWzUg0uIZQD/s7NaGmqZtky/5wwrYp911kuO0/dVz6dlbjTIeg
yU8h2UfcbTymIm6WNziO29HHUFZW6FMgmwMK1xtvSobu08z5Kf5JM25DyukOXV0E
0q70xFkmGvPVabLFEySnGvoMakFgUw4ISacFIPXl5GiksPZnIyjlhaJUf3erZC0I
8R09mgS0LXPnNnv8LzidHjJ5MRH9yuElKZp3lSrjRwKAfQtIJltwtNlCBUUyulSJ
mMpcOpDR1hmQvDls2452GLJEw+4oATiyCeooJ3SYr2k0rg8EY0AWHhh3CGkyRJCL
1VswYkSpZ3GuXunUGqnctSF0EnXHO8+YZMPbJ/8KPohdknW8tJ2LEicHyo+Wm40e
teoODMflX9DEqn07uRNyWYZf8Mqbhi+g1HoRjWk9C0cVbhARYkRYChwZl3RHHEyX
CxVNazqVzBrLxd8gxrO0jhI8vNe7qFzwiJujUzATOShX4RTG226LWo2D50mf/Bkr
6YfZVX8HnU1ZiI0YYbMnkLwms7i9KT0jZWyucbkHUW3QS0Oij0rqQkK9NJLbGMbN
8YgHFpkRzJ5XjegrOKRCShjyf4kS3paGvt6hTZi4RW+lB85LeMIJM+l3SoilcF/U
/jWbZffQM35dQw/MlO0iO5CE5CM8bx/88Dfz3unG7CYwzMU12b0wUDd6gnE8s/zA
hFU9VS4QRCDROyy4TEm2MDnLKuNVE3Np60Q3sS3Za5GMVPfTWlyFz4G6RIDyeEDL
OBQv0M2nlLJUzLExYmRI63y3sNnlTt5pZhOauPjBdN2+zWnfxrvmfZkDSEbMi//P
Rh8Qj/w5WbUT3T0y48GToOww9oKkIvgO5DzvRtBZ3jBoPPV6FbHMdKz3D6pqx0ef
NIblKCBVkjk6M+89fXO3xfHGSl+Du+uCbABBTj/UMU71c5iDsKxGHa4F07b+c1CL
kobxaT8NpcSijoKWwJeIs+sI+WXz9JozIqOo5/Bmq7SyvIqs1ssR8A8yG6Cj/JeV
O40/gW2D/ic119gG7sGQg5IoQTCEmV/YXGyColdXSfl/85iXXapqzAA4rbK/GJY0
jY/KoVTj53TbPc+mO9JN7XENqH6XL8H1IP8oVW4rryXUGcyrHP1Pi423RtH7oTRD
GX8QSKmv0t7QD0v4oo7+JGxueBVxO0L84iQMmRF398uyz1ZanOu7IMXAbfL1PDZt
Cxha/9KH5um9WH/ZCgn3EG7uRNxkOG1BsiHMkylHneriBquhGpBO0Td4dwnIawe3
7jB62eewwB1dyBD0K5pW5TDtz2OTZKFH9SnP9JC283Uy6nuXOwTH22Vt2LUrKt+R
Q2+5Iq/99LkBCIvAnoUq+WDnU/PeoHY8Vrs0C5kj/ZCZYqYPzDgp6lB+BNYZN7gC
TD/vq2C6zvxvJS4Fqu+htZ0AnYtLig+5h+XhZ7lMlsFab3PjyNade69yNoNHD4Yo
lkxc1qGcqk1BZTZdBcfX4SBfvSNO2MYwcSEPC0/l9ZE2rg784LdLU1Pyjv9an30z
B12FJIx3RqDUcHSCbLmd9jhC+7Wsy0A5DjUlPtBMxPOykTI7kvQc93Q+NsBbKiBO
oNNDwRdAaM1Ea9qcdrDxWJdl8Ta7XlafQKxYhHxq4oEYK0Lsm6K0i5qWG6vm9AQ7
7OapzonQfFnBFtzTxZzWCo4jOqjlBfvdhcbBK4Zo2WbyUg0M23Wo971isXRNqyLg
S5CnIjCo8xlfWpZ6l/iYIlgSM4qSX37ZRR3rSIeC6gAbhRqWrMM4Ep3iSiYiv7xV
ZwpNSb45FYOi+wctkg1J2nPsjf6MD9+99VByOggCgBgCbx6QtbvH8zzONVhykuKZ
EB59Yqa2fWW63/ZKeKx/8M7SaOI0vtl+/v6Pf3QsA0lNNxo6b880yOH+lfJwzzDh
5luLbp5Fs4niDo8HLUEG0jMv3ojPIXLJsqT18a1l809hv20zcAV3R7HIHkkLJnNn
uTytMk0bK01UtJ3x26bHrkf5296EDU7wJioQ3bMj1HOfJDdE57qNlEmNN0C9kmSX
MoiVGeMgxWwm/u7JOvDZSjDukI9AY01pgopHAQvXu35k3I2PE8NbCgzItcq1wneI
Ij/54YRVjz7Ru8FYytpfZQBT1W9vDgETet6GI7HN9J4vRI/ej9cQKVklzSnHp3zP
0naebsH3T+BBMbPvuAZFksO7M6sDAPhfBd3Zu0sDmWQfV7JUdqgXTL2uuMh6uo+h
prJlNcBMuhM0U50HIQP1P9BlXkI4MikJG0dYkYE5/OeqInSJHUBhtsS9dDUSqV0W
EBRtxUIfKhMzoqSa13pMdkq1yoZpsFSisNgLnftmRhksvmQdalfCU19j1wAtMTTo
Jukn8PbFqkdqnxYgenphlvQ2vACCSfyBS0x+YT4Lkp08smBuJ+hdoJOzo1f8hmUJ
XBNM5PvwCL6lGSQC+VCqbQ+qXbDb6wkLzjAY/RZPkAScPcLSLsoErSJ0WNK5WURZ
eCHeD+pBOVAsQENo8X6ELJOgDjGXO8dQOnqi23vZ/jL0zJ3Hfgeh7YWdtlL7LzGT
Y28jKUgCQ9vA+3qO+kp1zRlrXCd7gOTAkFEoCXdwrjy+g2NYa9Clw6SFytoXmM8x
HAVoiBwYiBJuOJGK+CqWO0VJLq34g2wOzn8aOyFhkQRmFwA6S01zTZGnWQn9UhhP
WjOo4Vd3SKColkGWy6Zienn+WQJz7Fcpu145qf0K/Vzpb2zZdjg9cWCj7debuG+S
L5aGaJeC1iUjWnnAgYszanldQGPnQ9mlTu4dHfXQ/LGjwQrmIrGQ0eN0M3STTE+Z
MTqvSnrvU34I8KACsBwaIHWrqMShk0Knckz2+zqpANsqsF/bVVyczUSEyyJoWoC0
prEJusMxqCfNK94iQV6YBonhrHb/7zkfzemv0b9xAxAnzfI7VsJGGrEH4/H3wqkb
cuu4pPgY0CrJiuHLzZwq2SuVisr02UMJHPF9+lzY1AZnmkZ5bfQTiZJ/V8lP1FpT
7kBffAl8CbTorJ7kmzuMqwe5ixCmtldzzr2DKu2ZaT93+S+zwacjJvCg25fVCfF/
Qxu6CVrfv+qM+zmL0huvEsD8zuoN4LOAqg3AsSajZmisXZE4PP9TnqNHSNS7FvsQ
hON55nKG8T1rko1pY7Ph7+LW+Ecb7MQAU65AcDokQVGK3cnZX3cIXNPn3y/MyfWL
vMgn79RFAwtNFSZ1GrSuIF4BMXx7Qelfc9uhuuTAlRRrjWEKDf78euYfnOo3m2Aj
sh7f9+bPy6bERUcVNJYbqUrW+HXMR9P8Bc/n86GhCskW1LZ9w5l86hKNaVTSHAMa
uHWxQPAywBp/s7ivcsnytv7WXfCT7RLSb6Z9lOyIQD5EAaRWVTzmtq0SRMLBfS/K
DvQ/ujcoQEa/yVq89fZbz0FGBQA+ZS92+Gt8nZDCbpaqI6IghumLAdNyo7X5I1m0
Tl3KbdapmDjeKuw4/WBzqYd4ixaszeVyROM7M1Argju54a/WwKOlfGBXZaF6fCzG
8mYmUi4MJwtW/GNGXkuk9O2cUlrBVcjbKWeXUSWmfJenlO78afoNpTQw78qCF04p
XHa/vmKF9twptH8ngkx3a37XTo7TywACgf6PgZ3aEu7T/LBVYmElBqS0PItXu1Ia
2DL/MqWFRZJmyvnj2ji2oVtl2YFTZlUCDUIvYYVdBZ254UM6FuljA3Ar4he0B9/9
ufnQAsL2Ewo6kjEHFIkpHdVfnvCDZNyogie/mxGNKHQbBm/mpqb9ArflzHdLaY+/
IK5E3KMMsF1pqZvGSyVzvSPUNxs8+LIyGwKn8M1wj++RWJp4pOfbujB/8z1QQDYf
IjXQWQJhgX/ChpuCNmIpFRWjQTXzGGJYUs6//vIqE+L0xOiQlhA5gZrJwDG/FlFs
2NOW4tDe7RGT4WT9/8dOkxYoiSGgN6VlQ6i3m0Gsp0yczp7JK/b+1oZGC4TaJmz0
9kmyClB70e6tx/tDbpzrfbLOC5bf2tPLSl4e3zaveNkrE/bcnYPvabVSZd3zeF4Z
2Zpc04IPT9m0/i7nhRKYMI8L2afqdcPpIN77NHVyuiR52COAH5UmTh3KnT/5Nii3
9sVfznYnVg2P9Nlk7oZQAPJPHeSqNAfkDO7rQGTAafN2kZg/65Oh/+A49p9kyVNx
iV0X+wjKOxWYqvBBkSps3fRKMlbkYZu+pqWKRBMoyxnSr60TzdqkBPnFpLa3HzRD
cDXfMes1mpsHWwTbatiwyrvLvi6bSCXjS22/tpDspxX3F3tpazfmkgRCZXNRjPLQ
slq9v9fwvs2r4bcfOaTDgoIduT/C0+zVP/Rb2JO8zHvdZQxXYoNcMPBpcnLXvtig
ECymWi+WjjSRqSyimQ1YKxuoQjCladnI13DT39/7weegygR5gapfzmpvAijVJrJu
0YYQpJPGD6S/JLSWX4COQOkt0iKlqmnHYmtT7l8uydsfP6p4nhGDzrXhlgLD8zJV
D4+CyzFYYm5T4TXpEuvXTyZ5nf/I7RQxzlISa5FzQAsCQtBssFXF5aDO6LhzXVTJ
cOfudesSFMXFpoFbTXS57qSJmjeznyr9CE1enjBKW2//NVHWqjXaZPZ9LF9YTML+
CL2I5LZ/Invl2VBZQBy1XcLQ50BNaLgHVcNKC7OOD/YyWL/xI/nEBpP9+5tYpxVG
10Z0FHoM9fSJTjmbyjOAs+Xl+DGJ6TbgfGfKAeOdiMMwtFbPcos5owf41ZK175T9
zQvjJjjimd6U2X6HWW7U8cWvpRsaj90b8qKc10DzX503t2iuSqq1xrx3cAi7cVza
zk1mfRfmM4BgIU15Na9CzxweYHt0fCBhGa69rMbeEzcoHTQdogQtfB7wmAV/ATg4
hwpaQuD3CvhodWXgiW61jJJbaz/P7y35hX5EGMJpJun/ryT1hJqmitxncLJQtnIF
8IX3YyleuarlTsOmEHetYULYnvXBgfSIVk6jWqkMDQ/RjclnhjleLs9OdyHzrVmq
cbiRyg+ebpLgeCWuM4kpvJUW5Iwy9x7FHy8OYNXzcyIg9iLWGYnxMq2pGWaZK9fo
jr95cBSe2egXViCPJW6nbBuquvKBSFF7wBW8AzWIAV7yKXiqB9Ho/0IAhn2xQgV8
ZbY8msTrFj2TqDaCib0b4YfbMMo7Bh0IdKiN4/QMEzqXBZorxXlOnWI3prIZ3Gr3
Olq1xvGFks4q3QMyF+Eczp3F4Wwd5TigutiUoYAdk9n2UZdM7wVco+XBTlp71CTB
XSATiQAtyrvcMH636MwWlxmQyXGcPXPlRaE33s4dndemh+B2hHUcubhhwXBkxmI1
CM83YJhWOG7nivhCWQnLjy/8K1CUioszHA/w1CteEWw5MSERNbLj4PUypZL/QVuw
mnj/ZuGN+mQVKaahQUgQs2MtD8sOo58+/C6X/nAMhhZlEqY2jRduHCSqjV9dKAmW
pulKUfuyJhJh08qXSr0qudZ51uWcM1vsSYlg2YdHTRZnM7hh6zUQcjso7nBNgYy7
tmEcAD/+IUJx2sQuCTkY0Xzp+6sCicumtJlqSLLxcV2GNRnuSx+D9tw83nZeOQ95
t4TQ3oMh1mxJFXl8iPzYMXe0dXWOjz+B7mnjxl7DltCNjce7qJhOYOZv+sljhE07
o1KyrOnSiTbSdEyL4nlnTu7MrQ34NxCubtYtmPt1wzySjp2DNK/CwfI9VJB+pjv1
CBpa9RrHMeCCCtdfFLNNvofD9/vFwWPIzQgn6cb2tAtiwYi4VAx6Q+3jE3Q921Eu
VpAXEqpgU2sAC1olVJUR1FN1MbOIY96L4W6Z3sga5DNHEKp1UaQ8XKGRXZGK2MSZ
xR/Jmx406uAom2o3Y1CjyZXpmuw/inPGsUktXof0C50TPm9eDDrUAdICXZ9ua2/8
IFdyGVmgbgiawgTloLAzGXYv1H+BE8SoTkq2TDUubDDdexKhJDA7unlGKGMK4Sq/
4nHuqbVHuUSDzZDURnAsAouE5Q4YcJVXbSsdwL+BKG43q7tIADx4QRR2xKVIc3BW
QSFZ07an/ZdBX5aS5S35ThD7TBBmYO1h1m6ydCj8EhBs4J8EtYiMkXE2KdFyiIN+
QEO0661dzBO1/izZYJYoheR6TyJz31bJE4hwJmYKn6lS8D+PoBApyik0ICV7drPH
c5jqH8Q5e9y4KCsWERsse+hFAofTMRJwq2TPQpmLJO3JvF1uukvpSECQeDoWoJCx
oZVy8cFsFy5dprVG/tWnwgrQQJiPYmemNSRjEHrqtgPyOUo4afDltiUd3mSgc2r3
PjWnCXE6uYZkwZpgbkpMx7X1A7NUadgesePA+22bwVsqEkC2mO1G4/ihYzw+nUtW
oF7XrdBwwD8ngzwMI6u4K41ResGhxmJAOV8CUyDOZGLEDzACs4RXSKfShfWeDrGv
snItP/9rS0ytY3N/SmlruOgSlDKukvwKEg4kxFKouM6N5kppyWqa6ezImXsYL5Ws
zbkxls9EeawGKNbXC+hoXPWb8W4o2MkEsyTMmQATFN1H2tCd42kIY99rKHP182zg
UYUvNJZWmj9CUouIfXT45mMoPZa1Re6dExoLbH9CZl0JqTJVgQvpGUVkznVI9VxK
e8Bezg0HFP1bBQLmaIRrKkvNt8djof98rJ93xxVGU1oImHLr9jTo9f4NjJZK1rT+
DBWSoWPpkYoFrZIEvFt+GxCK4nJjVLPoruYUUMhBko/qeqI5458a9dG1OFFYJsKN
6+TSccCRbwB3RIqgrDanDlPBpXvoNJNfngSBrLPErVQgUPPoL0GnDpCGoOlBmmky
j73jio5dhbFybq1sYaBfHXMBB0x+f9mx9HlbYZeYECJR6jBzmHDjyXD/Y7okTJU8
tNW7Q46oe2hp3ur8oCawqhTm282fYjFa9omEcXQeiAuHvk60qAAIwtWHL5umhYka
yMhqJCstnPnyoFuA/jfVsBKlJ9i5pxiKvYZ/yryXvy9C3z1CLEhwwnveUZis83ev
X31ELw+RkpNc2Eprf/6Ayyfa2rSHdAkczh7b51Zh6Zy9HrfO1lA3C4sOlG45JKZF
Fl4TLfGeKWPwEj6ZLgHyCPNofXKTaWNvQo3p96n7d5Ak0O+gg7atLS/NXrefuIfm
e+9DJSnFfEPdyGALRz1rJr2PSAsMgvotdzQ7sI+Hm86iERG3p0Y2aiuURMWQC374
b1tpi7ColunrPgduXBOnpCG9nkB+OdtVcsYfglsx4YgsGZMl7uKGbPzMdm+SX51q
JA5JN3wOz0lF5QNQ2A4OzwFON+eD2me2qgqsFS5zMidoUG5FBmjbxUnXXtKprr9h
AgEqTCxPqsodKWdc0j/3LX2eCOr62+xGUJ1jwxZvJOIRDRWkdnbI+6F6MhKE1BPw
J3i5SQHOi5BlOq4UP4yQggutNC4xF4xYJFBPZnMS/BBgI3YPhtk1j8Kx3kAUd/lo
V1p0zULkOri+i+riYOyw56mACt46ucCU9dBo4JXtpFC+2VRsU1HTjw+b5K31fdSa
nmF/t+l879XzPcGchQWv9x4ZMsvriVBkwByMenOjebuL8MtM3tCJXWwwL8uKlaxe
zbAw9shyg0R/u3SoaH3MpgluZvf1VQTgDrNd+TDZZJy9Aji/pG5z1nzjoOFLUEcw
9GAWbPTGx0/bAvZdPusOhc/jEEBDUtHSqmJNIvncMrAIEIbumGl+YOMUTFLIkFRT
sb3CVPZZ3z8fx1e4BBioltwZ+KVJqM+lakqjfZkFaUbWmXSVqKVh/NCn7hZcT+rY
0HyYgfRCwg1eZf7L4OQiqAmTnPf+0Hf+lyKOLjrOmUD6kdKuEkpaIvuvS+7wUMc1
FNXreMDf5P8O088ftFYMU8+n2BJt2ZpuB4C4Fnqw4gke0x/Z3+BwyZhMbaNUxL3Z
8NeVHNEx1uEtmoSs0sIZ7a7R2dn72QA5bG/jB6WChYWOS6vQOG/uuyU3rbMeaX11
dnC47P5dP6NqjCLxHXe77CXde15ymVhnJvXk6Iluu8R578G734BhceYnzK/79yQD
WC+Sf8PHyI4auww2IcHb3V75A7K/CIISpUuUAyYIPC5/u9FC8qA7WcaPZKKBJFbu
rlr0RlKGiIeCdkxKav3bAfIXrQqIKCuVQrrvgnryZ3dD5kV+Xf8f64oxi7yeouWk
8jx2/wluV+HIfVJ4j/RR6RX2vjEZJ+OBaITrVjq742k++uOyyU11dQ+PMPS3pYKC
q+rnYuzV53IFErdvFX6uWr3OC7W/cI3UBMi8XfjLwpAbxZJF/ekPWDGxhLh9LU3+
9MNU1wtvtxwlc0jDQqifxtTOCfMp9UmZ3mhyjXFPehq38sEXUKHS0JDXM9ICnqc/
ubYvQ+/Z6DNMcgiYeJ9dRym10VPV76ZsZ/r0W8KKwWj0EWXBGpTQHUwoZqtKZbVk
YZd2S0V7osB1wXd4PKP0m16cTz+fjqTiq3s/yvJTtIKu2ZMTB7c8CfhonrLtM138
olerSTTKlhg51cbM+r2vYxeOPlsaMiqmeSQyRUz0S6u6zNqgxDI/z2EhiHYN8VpS
FR7t2xwyKHFlf54IC+Q1l0hTabVC9d4zoPwZGmefEEsJobEq+zMbbuytzDg7z/5b
xMBIJ1VvQQgzdCk6tD+QCz18PDNyczC7jvmYLp6vKW49rG/YgHkfw5s+1Ka5dgPb
/xsJ6lWbAqZdBG/3lnO4knScsE7A1WWEP/q6NyVGpBcjqCtwQxCqNcI9IxStIyvK
jRe7mk6LHSaGTLsC+oAf3tnhwUyCoVUIKKq6OWUmpaTfrXiR0SXQPoZVOl/kSiEu
OlFfvrcfYq8Rt9qc+AR6FtATSf+XgVnInMgpKmmq09k7MPi04CHi81dcPdbylLui
MGC9Wq7WwoshrL8nDQafA96mRxDkd7dkTYHLTbSADgFboidwA24U3Egvz0yTj4C9
+Be/xmqBiJr2vR48C8zKjnpRwIGfACSwuuV6HO0qngqPZNBaS+u2h8Llaf2Er94+
Jp/3EBnLvZJcXhPEd0QeJuTFg8B60kMdoEBuIsbEU7BNGMuzxt4LPPfI/JXv5rfO
+uw9crF3HtU68gDLMhxcsttXwedcuBZhPl9+56hF2XD7l3BF6eKDwMgLTiJZVPrM
uw0gIfrRk7YtKe7qww7kKoZbMu0iXLv5jvD0lPirBf4jfAT/a8suwj+ITXhBQJRT
T7OO9C6qv/drTJHhHmDyPPoLVFDhk79zPArAoHwiv8uCQEjIzYIXl05QLGuYE0Sr
lXV9y0TSC6fHmzzln+MrskoNsXGkvsVkmTdngF6RMpswmDY+LD0wseAJcZYcOjWT
4JvFw8q6kIRxNAmstAYaVlthZt+hUDoDT17SsbRYywv/1aGVHCEEKNXNTR8DPGJF
DQsbofF7x84lARXKI90ncpJzJEovb6Bz3hVJIRopcHA5qsVfG6GtUQXgVhg4cM+v
s9dbXterwvcxBt9OvRBwEnVPTHKmhk2M/qZw+7N8I0RL/EpC90WRJ+u5r8O9J8KL
/b1F3WUQRgHSI8X7muuAxjroQGreJMq3HIVpZxPfyNcjxIkTDTK/u89aNtx35Xb6
9wnCFpw+5E3xW1VYDBS0Bik596tExrLyakg/2LCfHJtmgnkYIcyff7KbTL6xBs6F
S+gNIfKoWbKy2KbyzcT42MlPAp0TckKMJfr2kQwF7xgwub8DX+45wQnyWPccc4lz
AtoT4vAT46MpJ1boXv1chIIfAEm9dkI3rfv7vWTeZXEzhNdMkqbwD5wsE6E28T/3
UmcekpFFm86G8urPktS5VdWiPqQsuLgedvc97dORhd345+KAKQR7kMjDc/LUnZYm
crufZmZ54I+0LS5rDsrbhCsFlo3AKvBLVvqXP2aCp6EZxCi08lfd5JEm9Yz/Tldx
qDYR2q6D8wjEs2DG9Nj5dRWSAQ+45tr5hOAbnRWagzVZrLPvd5W/b3R0pYhyrAAa
MukqM7UVG0s2koEJo3FO3nVWYePpu8dHmo37IrW71F2Fm5EmjkkJkq8ZNeAtj9vz
yBXK/USPhfCkiqFCxjugnrcBEZuerLMiitU2bq3Fe/h1/pBbS6PWOv9gBgWReR+z
pp4oxccVpvB5xmIHerZto0NgbaLRCFBH30WKuuHfr7Z0jhUsBLrfGHRB40X0gHyj
g3ekgxVJ/0QgE8IprxJsDp8j4p4zNytduf92Kk2QxEasrr/7+NDeahumsy3X04hi
NeuQnw2VRGPoyPa+82SkndLSI5vNgpcnarKY8bL2xvAVqbGv4qb0X0Dd+1w1c0Yj
631PFwU1dLE3AA9KYv9823jK/FdaAez20Nyf4b/ilgLZ+rMlIDxjsynIan4X8LPk
rDTgogrGAkKlJR1o6fij6BqBKdz/RZ1ACbfixWyG2540eosnFdbankeQJ/BFNtza
Xo2WhhGkZHzzeVtcF72e7uwCI9qJNt8Sbh5emi+lfZH0OJjlWSD7GU+3UzdgHxvl
dFpLHPxCCho/9wITil36VgGTvqIBiL2qVv8AcQNxcb/0yTeR0uny32ZVdhDTfprA
ASMLC/mx43LZo0zlKFmL/yaJnCCTxXte0IpB0qjOph/B/kIsiomBHe2PBG1xoNvD
pOjZYOy+Qetzoc10j/6cOBE2GhpZK5MYRS1BuK9ysdSDxc6eEz8Rb2/YcSTO2VoA
03giUJyJ4m92SSptHU49vLfm5x1xXhqskM8ydMbIH3Oabuyf9HK2yrArvaWV8hBy
TkycMC4ZvJt3b660VOlD0NQGm6mDMU6Q5+QsdwoXguEdP5HKNJeBFt4ZdO1eWmYO
DbPpJwKG3Rbol9BD1E+AISh048soVHQMQupEJmRRxDmCK3EjoQyoM6dxcZwmzJip
fAA2zCW/D3CSqWR82S0TJoqbnES+f6Hqsy4HimvuYG/HNuBrzx/2pY+R42NVatTc
vqy3+RY2JPgUGyaS5PzWlCK5Vq7DQOsu47SCyJeg6+AaMjRFI/vPYRuqydffVprx
EFXku7uRMXZLBF/vdPKP4jF9iNID2G0KRYqZ89dScTOExqygN150nmiz6muJs9SZ
wv1i8bi1Rt88pHVUY8Dbm4cWX+p/AoHy+lqx99dBM1MBmUWQO+yDq3V/BBkq6mDY
R8xMMZKdXRapAGzqc/11tJymD4N6z6TD6jMkdI4GQRdFw73zOIecbmdHTXzfnY+e
c8VavxEE5atYcH88+bO6V8xEtdCkHzjKksdKF3lk1hw5TAnKOjDjpWBwHx8bcshM
Bsapnl08OGLLN7Sk3/O8Kfv08yJ9ErgQaVFLcQQBpFeIh7bnAvEOozayJhMa05Cw
ErPDmxk+az54kvgc4/UF43eLpYoCsJi2uCCHGm8rQsYIYZvct/cn2TZPA6WtcAsD
EHxxZ/tQfr3yl6G0Z3Ev3eWGtVXe+AMFdbi0z8kFqQmM5JlaaP8ZKNiingFvHH7z
KaBKo4LraLpS8UyZdRME0mwdqPVngv1liSVTjYzTpLeQXMixhPp24sc+AHvZoJ5h
rZp02GIDyT7kc93KM2QbvPdfqq24ObD70zQk10veBraLsngk3TRuysE8tpPdNAZK
aNtf3DVQolzjcQnwhfEdZml6RK6+eaMfWNv/FNUveWx49m10P3VSHgxH9mBgfa/7
rPgp3mi7ApLdjcl1agvxXckRnq7ftYWMBfdSdrEoDUb7vkw1G234xekzxwn8BSv0
q9jkTMe+QzOD9oJj57ANbWw5IBfmglwkVwto1xbtklJ1ui5I3BJtH4f+54QMGckc
GiIfCjapyq9wjrfYj2jwo6+3dsaeZ7ezpK4TwwgKMkk0UzcGNYnRQAP+mdolFg+a
aGIMmqkOea/tXBQoYPH4+X1XizQ+9z3lNyVMDHdW1xxq4PyEhPWCNjZ4fzMJzII1
mcGSyi9+MAfK7FyqIJfwhi0936Pe0rtPBqGvVCmbnB+1efbwj2P2d5TRrHKKXs+z
0JwVsACOKr6qnv7aOZ+BG+XngLK4nuZROHfKrDrbs5LW+4izyIbyBEvWPF2xeNdV
kK5JM8IPglzAm7NERvIIpRMdcqKeBFfEOJ/qJl23oLmfDlt6FnuvoTh4Z1Gdds7h
6CfFE3SkFxIRreoTRh1xZ4xuvN0vwZ50a5uxFQq0sSYeW0+jDJCGVhmco/8I5HYF
dfVEL9pThjDYayKoxKRyzgpL1Dp+ujF1zcXXj+8pATJ6/3mkjGMy1m+jkTkiGwgg
D7HJqah2XfYzn89tCmY8Y2+WcCOgpu68Vx29sknnBYpEWo7JFCIyEpaOzKYZH/8L
FBad0f0ov7/cFWumHM7Kxfha30cg6QjmkJPkTr+rd75Ul/Xn5wzOl//VfgKPfkJK
RTKpepfwTFNMLw8dWT73sh87Fh6NnHjHsdogsnotpsfzvudgKkqtTX1jXZAmXGmV
olDbeOBalYQk+Np/aQNTHBMYSFnpzWDghL6EnrsWNHChkpNbYcpUC42Fg1/szVH4
eOj70k0Eoq+kX7Y4OSMSOfzOAVO3IeVWd4a8pv22MkXOQ6YeSe9jUwiiD2D9w9P1
mA1jmOVuIDgumIuc4b6OqfvQtDtNBPkylF0EEzaHgYMLVcS3jwe1DLDsUHotgkCb
FU6QN7TIESTIkd8ByooxehwDLRTHDmq6wZUCHwyULawCb7V4OimJDJJQMAD2BBEF
/zeqQqqw/wgl8iaJnDARN1zexPj4fe0T7lxqRAizJoxNvaJB2AX6hC2j3M/Mw8AS
H7UfpH1SXwKasTywkaHCdJJi+T4RqttdHGN3zAXsFjY9vavN6ZNaIfzXy2ed3PM+
FIEz1yAN23lIKmiySnJ0ezj5MbAxRHNjt5x647XRgaxtekMCIc9up1KNi4T0+YiY
tyFGq6HHsA2a+Lyidq/1qN+jn8Upx/uV3MkkBo9s3gEiTfBSxDgVwvl+WanYWZv5
CiAbwFUWkZ0yAvHU0Q23iGFqf9T8eLOTNwdT1Lfw936eI3OYXvZtkoPzB9uYHobV
1sdcqOdpQjqtXDJzJzlG/TkkJpC/0jU/Y3LScIXm2WbNq/SgAxMLdxBt2PnNy2F/
QpL/yIRMOpelSASGJ4ujesA1GT1TGWl6I1fCxJyXtsM5AQOHuVmN3aDOnAwiwAjR
jMbA++6Q4iwMgE4ay74ce5UimwVwtDFCHvb5tH7f9Z7fcykpWbXUu9E3hj7irA/x
L0jZYfMkY/jjxJkCwR2Vw3c/HWEvQ/nKucfEKzcix5f48/INZ6N1t6uyu1Xj6TKQ
iKuXDhM1B3vSwNryt5pWgzESk103EibXWszlFRZfw4QM2xiOVq32BJ+gc1tdlgMZ
YytKktZvsMg0x2IOsQoVSalhett+T+dtRelfwE7F4Utv2L1qco66R+VM8h3GdTg6
XmIL8zg8JrNZTP2bJA5AARwhtratkxUtfZ8jMx4VFEPTIiPI1NYJM7HevEw04MgR
94BNzzpKksgP8BBK/iP7nKNAOP5WC3o+Rgkd/FTK3uHMkWhYVeP3YC1k5xKX0EJt
INSnI/yhyuLpLNlec9H1J+ziOGwQxt/UmI9R0YIRDthlTZmcEKsORynIq3w42f+1
WeWf8VStzy2zzqjZfrLF7Pk4DE6JptS2G3mc9A0VFdANMuENcfJ52Kfdt/wUHEZb
3KV3/f3FPn7ahG4He+lTlnKyruEGH8ooErWVynczU6R6Xz3tzVnFKjJP4920gCDP
NOSXqtSIBox3o0q87UTzLaPKTffsbNFMe1wUDguPikYRT7IvJuzi48TP3JItgMfr
QW6sj2hAuSS+CxT8LHYQbeyjp3RDruOX+MX2GZ2SWLoHhBZVrOkchQaiGEuPe5Qm
fmm/NMH3TtzNdlVaGy5XIjiGVuWlK+HfB1Ex97TMIFq1b/obIZX+4Uls+WY0UDol
JErQgbzngB4D3lmx++BF9oQWIbFgF4/2ymmKyZcQoODIDE/Rv6DzHQQg8t1KPG/s
3Jtb6eUus1Fh2LB/9n9aJjZajI3hCyBDaIFInP2abj8ipdrb5TyfZy2NItKAh8ff
s7bNyrJ/ismfyMgy68aLBJDM2tA1YOeJE9xYlcqeAb9dwANi46Bvw8N15Lte89Lc
pY/0ZXL8R++MA/+jxqE4FI+e3BuQ26H2NN3FpTcxzwcqGtG872X1X4UxVcyf1DhE
xQy1hJf+t2O0I/LnyUG7SMRgj+Y9ylO7zzCBSsS2wqv3RSTcoNNX6MH41d1MZ21h
RVLOg/AJobnl4cvVw+e9lZ99KiPMjy8ZqN3rB9wG1z9kgXwTD35m+PPw+HlxQURP
gSEngz6Bs8OMX1d4DfCszfVV4tzdDqYRUVsX5dfJPRxKkiEoh8vv0Z52bM2CGCTi
37Cs+ViRVqg5pIWoUzh5sY23Eu7L1mOig94B+a4Ryeqd4eCw6JghZIkc+evnXRfE
KByDTybqpSzYiEY1pTJU0EcjcQQz9s8/zhRASPWSrJSht+yEkcx5eTbfR0dueHe0
33LMLLOnfowIBzuRU5FyP5Gan/ekPJqNHwCZHcn7Cic61rb8x0LacV4gO9n7NMFK
fxp0nSRnonSSK3vUotzGd1hQCbal7Wg8Foch9bArfiw+IkDkohh24jNhviRk8NG+
rdc0o7U+rO0E+6EzOQmllGoyycyNAf/y1mZc1yHSX0DvqXQ9yX+5BEPCrnFrnonz
wRFgXmdbXW+9hhv7tFKch7cRfkNuHZItBEGDzrUOu2F1QtgqfdhxuOcz/57Eaybc
uF2GhyvBq3uPUYfxW+9rt3NQ31uK6l935TcihBywPI2/AxNbGA7pl07HCS3ywqJm
yJFrZYFeGNpdgIR0Uwig4RDFbSDRmL/rMjR6LZ0plWGQq6qjAk95L1NcWi0Hq0v+
csdeG1htpP1T2SL7SvSs2PJSK64HlVpW+pCTLYIfxy9AxIMnWSMKh8C5lue1pUku
p8k4EzMAjo20fxdChecnlImKTH4AS/BsZnbLGXT2aNLBTKWLb4eFAtxA2EviKTwj
ZQNUYV+L7Xd+yyTAV8MvZhqs9EcUyJxQy1v5fERY9z5w5J4/zEirff20pCyA9Lpk
Sg+TXUf/CSkvFrxo84DZyl5dG9HKTqG/qXvXOUbIcqVGX04IkziKqL15F3Xak166
aNtUp+CZZookv82JbYot0lAqsOXS1sHXXVgNHQ5c26FL7CYdghTgxSeoE67kzu/I
p0aSt53+60/i2gOBdsjGwNzV4ASHR82pbUph/YygwQhVL/EScC1EI2iSw2kfdsVY
gDepTA/cEDFVMTeOZISITuN59kayPGFr7NdUqcn+450XeuwssPNtFj+G71ESN/L2
3gG0EwkUaJPcLkkt9You/jhGDcEOtNhbmBcrUxNXAShJGpwOAYEnnwPeY4kyjRJX
3F87ygjo0ySSKaYp1Vlz8qyehGu0PC3UUSEDk6ADaokdzyZu8mPMNnO8OG0N0kIZ
+BvV8RgE2hYonQnyKgbYrE0rlhiBZ3QtwrMODaq5pCJkSXIVCmDeWlZgDKnncnQz
oAWfU/7rmMnDxNuCKVpopsS2OHqWILo4sPhUGLjOwY/S+25wK8ji26KcPw8oOcLT
wPhDdJHeoyfqEIwDpqDhw6LkD3/mO4JrU+LVbHxlFqrMdb4a0M3yukS5c/zSdGfZ
pmuswYDgQyCATQarTWpbkSG9uOPK2jqsmMrVUq7reA3nu2rHbR5NkRymfS60bFUu
0S7YNVA3ymYBm2mwB8FEGpcT/82q8MamqvONsTu6yc3WdKtiw8DoyvcVQci0rkP0
ilMIZh2hqNRC1MeCQdgiektwWS8iRN+hdiQCNatrSFBBzWJsBFZL+fswGBtrZS5a
eMC04WvsXNYXMT2vt4cuH8JvP59vnK6YgRxOoazDP7D9muF2eVnLWx/OybdZv6hM
RdgIMlg4qicxJGeeMYogRlqCvZCAcqLXGNez516+wC9WE4t0u6rEFdki2SIaXUFX
2KITwvd91OGielIm7GudgIJN4Ezxinxw/qEIbO/M3GPE156N5xWnJfxayAHFome8
ymGQKMshKNxS6aySY0ayLvRLfnofzCIC/jYEf6Xexsj8ZYtNoNuNZhwu5kx+m6mj
8CwpBhc9xv+6WxvQWZRQYWnqFigyxyemyuxuQEmVMYqaVVlFaiH6SX8A854z5m29
PJ3Bw8E4pyaZlQ0oRLdy2wx/8XnlLjxavfxjYQyh+wHqwbHBkWBdmXbZlFGxby1Q
+pDNYp8QbRCyZXGCVbkYdMZJjwHwEYZa8VqyNCyLXJCwNLWttLqvGFnkD7kAoNK9
zQwMXZHfZ/AUs5b4aCyBh20e7eI92ZV0Zz2SgQm8fZSd603MRwXQQOOH79inHBQP
0UzsqUrXTQdg8N18SEAtNXhq3ePvaBs6/p5LAsysyttiLrm+H7M4Mh+/a9H5EIU5
52kW6/fGKT8zbbOEns01Qx4txv8L+k3JaufU3AY8H9G1zQYgTIFEy9+HZ+orajmG
yaZgShzK4DCTksNtLS542CB4cXsOIJLCfK5V5mrTpkF0sekROJeGQrXw9RFxgNSI
yhh2asrwg5pd4Qk/xffCMdjBz6iiRC9TRoKE5/6buOFS2xs/A8GHdPjL12KpDx1M
ZeKgU+OcC1jgPiPsECa2TWN9xWc68bn2YJ3jp1NuyeRel2SnH5d147dygfM0yqUK
9vNPK0S6Lwk/ud5mfUrEjtwAG7/e6jYMSibZMEPxwBpkTvmog/e2PWWYeNTyz2Iu
EjlsC/8OiQ4WXoCf3u7nV5W+t30l1WG0Kfz9fp1mpxLIsDs34j+YQtPz5KJXPhAJ
CsCEUgfpMjCgPoZ6X3d18W0NGhRPhdeg4vYTUBAg4mlGavaDB96gedZ2cSSCYPz2
g1DMY+gkRDzyv7omOy0bN4Cay0mlBvzcbmDPanbj9rOYyQqoVE8B6JQkSBG05YAM
yPExi2+GarGHJ0eFQLZXNvcqIFFho6BhZi0F7jz2KlFANEnqECnXvchRDBe2sZnU
Oy72kL/DPkes1K268hLLhh09NYZ+sP7/VdUZD6+idVrDfMKFSHN9xHtO1AFSDsEk
4pn/kURikrkil07Tb9SXOCkf5TRlNOdcnBqIXKnjP7N/+662jK1Jx3HIGihnKS6b
lOHKKOyI3Zr2wzEQeGfxFYVcTeUrIHreoxl6cFRtFMnB9SVFSKMezojRfAb2r5kC
MGoA7VPVYNTuyEE5SA+Yo/GeaoRz7/lzTKpwYO56KVL4Ztr7nFGN7XHprmkzYjQi
zUR1NFypYO8T+l7FEHbNJcXQz896YHgbh3B+TKG2XD1N6riefNOvsvZfUrAniZ3Q
Y+EqU8dunOdO5B6VsY4IHvSQSwMFjIra4UUxA2FUCp8gwkbxAD8xrSpR0R1pPTYR
X4zBsMGoPERwDo7/ZoaZoG6fVLltvFm+SpWSJLDTrh5SUdpAA7f3iwEc6WnjWnDI
RvdUWOYiboN00pR2vU9zbZibuJWz1yabuMLnabi0nz1Q7A7CU5lkwmoKDlEKk/yR
7ryh9KpPQBGVxNVZIt4Um3pubHeF/W+lrrAytdxPEdxwpvkdhdtMksST4oBJy7LR
IUu2Riy/dnJPIimOhH/MlBzahAhoiu7/2FZ/qj/FnaHBCoXgKyExtEatuL87evDV
0Y46H+q97N2ejv9gnNDlRYqkE55lKr1wvYpclP3S0C3niZjDMNJJKslax0z3bt9g
lEz3MBHo78I+3ugsJZrDPdKwg6hN3ZuEpIs+AjllC3bzVE2uXu8yau0IBCM75hrt
Qh4Ryt7EVGsvVFKx8J8yArWwfq57cgwyfCb+wJ3L4gYzmqkwhoZgrsGgC7hIEhhz
0mtvVV99ZzwYvaZ6hEcBiFHPsfOPkn/kgPu/h7Oqu0CrFerCdJg+lGKklW3twOcs
Xjnjk1MNTZc+FaPMi9pBBFlAW98UKv0ghxlPxHmNEHzJ1tC/WCScxH1oElZ84W0a
HnktUJWL9H/rfYYfqr6zdJeuTf3dD/3Da9/DqrHfs+GCtm7im+gSF1itxFoOyb0z
xs3Aw3SyEZkIg0IbXUa4DwmzBxIqvAfVRtFAn3LG7J9AFd/+Dx0IC7rHmA5MP1Sw
+o/QXUPR9/2H/fnDRrIkTzsrr9z46e4+VHAeUtY0PWETSDDcIAizgRriv9icDnJ/
kqeGVc0pUyK6edsovknUSCoFuzTtZe4NsAc2iAuvsXnr1Xw31MOC+58Q4ZP+Mbrw
q3Iv1FDfr7hkOwCMSGakvJBCsURxn+E8/C9jA5DNM9qALbUkLo1osDwtIpys7kPf
9KYbjiw7tFLM/S7Sz7BVwIMC9yUTP34KbWVOrfsL5fxQ9FYzYLKWD6Dy5dSTzJeb
3REPuZSZ4aS1WluUUFJhV3fF5DC+1polRFyRKOpH/ufPFv1OpS4s/NiButkwTqQ7
CktYjw1Jfpps8XlUl7nMHWV6D3njvF69+JV7/1kkMN8DNpElyG6NS60pvJkZ21B+
cIvPJn+UGIoX7KaELzf+ew5Wstd76waR5g+yHFPFEj1wsy2+M8sXbAJzeKY4jkRm
bWA2rF/YQEisK6wNFcwIBdjUsQDjcj1jev2pJRTEsx4xIZ+R2jK/sn/CSsUZEU+w
z33kK32zs6WBrLjNgPdpl0kOCDXD3ZKkTIlMdENLglTGS13FwObz6WkaobSr18tR
UTcoXgoteMfxIhdd1I+y79ffZTdG9jXVSzmQN2FG+8h6g4zDTud2VGMXDbHn2WDz
R7e3lGfLPODQL5b3+Nlahj6CHOR+xfzi4ZxVYX4bkP/BFEfe1/SuvbmqC1d610hC
GSO6Hivlp5bhbzEHJhcpvPWql54oMNPiAaafyaNLxhsaJXBnJ4NuTIU24smIUDQv
MTFvR9ZIKm6bYQW9YA9OuP/rHOas0fyIi5WuwDvWV8n0jjQXyZ6tNdn7Vew+ucSL
tPPS2At2tFESuT/xDPtX5GyDKg9W4ueWw0vUU2NwEjTLvfUKEXYxSZV3tBPX1O1Y
/poXEjqvnuT8Q2X1/49rCAN+ZdO7WaW+0Lc4yicVCKVikEG5qYbe/KXOG6t923Jh
uKcUEtjm6WnaqXsxW7Kuih5MjWQiQ3CecctI+e1GHBRH34VwC57GMp/tDOGa4d3J
lpj/2QfVr8LNIxBkhd/npTRaNDtpHBG4a6DsWK3wghjijZo6bFg23EgcaEUIOeNt
04qzLPDhulH25xwVJbn1FD/EOPMWjZXbYz3NMxRhWXblmccdfg6vEz1Qv96aqVHD
yfJCf+A5j8OH6ObktDF+VehqdW2i+yfCNYMoyfdkhkxJeRAXZyCauVMfFBh4jvns
jtTU3d3e3poBZbc11TKH769QuvjVdr/nbTlHTth6VentUCgppIqSoFcZytt6Ioly
dbJW7e518vbL42axyUUbTipfLfPHPJJtes44vI2xQ9+nhaA86gzs0AUwaUgvcHar
zWwgTi4cKlI3r7BF7kVmviLDEe4QaNWA93xORKr1imOjmnzGVjtXGJuzv2LnEbuS
sheo3yhGmBC4kYmFFo4JoJTMK/Pq7PSW6CC9O6HoyHNybjD9tqjhoLNFSFSUdQrc
nkTorg7xHztvWYsuw/9BLz7X3aTzwBkUUKvDnNFBOWiPUP/0bmvZWl0+EGbSCjV+
bNoDI0SOCdtPwX61ZthgViSw3jVfr4s7zU9718XZxwUFQjh+NIFX0gugdQaS9cIb
bLIfLqPZpalehbYt5fJ0OycXlAB9YRN7xcdqJyPFzI275dZAGnbuHCUXVP0vWyoa
6lMyPMVhJlZi0bIT0CPcASiqj3RpoMERX7o9bBxG5tuVCFWk6lWXl1O3X2yMf3sD
DWyfVMr2uguxSoaQqpdD3PI5uY+BlvXkYwAql4sgSa04UdocNwT5cJz68/SGx0Zc
OqcwAHg3JmMtmLnvNg8SK3nmrGglQ3ejRiYzhFEn94iw61NYvK6OC3/sjtDtg/bg
xpFuU3FbzjMdYs/A8Ux4X61M1JiP/beFUA9qeF7b9IPDr/oW4N2uraWubu1H1CxU
TLNpMIDhpsnchDV/rVhfX1i+qzZdkSVw84fYA82sW0KhxwULh2hDhWlQ17XI8Se3
sSO01LBi1B7BGLfA7joNKgDPIbP3RrbqqSJCkT6Wfz5p2IezflylnOIAvi/i6Nzl
wh+ncTpXSR5ASDABg4ysiNZyGa6aVzs6zgSsHiQPiRmnwjNSW3L/YROPclVmaRFw
ark7aIWgP8vTTGbu/+FAEyyfMu0WrzPOjeYlTpGOc7XSCDCCMM3tjGwExRnfRFeT
1gWNhFtsLyPYsmGzu3fJDSKyqdPDeEN6ZMAMCgL1pqatq0b+ZGFJGPCwlqtcu9lo
SN6Z9v1tPeXZvuCE4vl4olRrXhDFu5hV6RtxoKjLSG4iGhCZO4p4r5o2I/o8B6UT
cZJrChBXTILH5NBq2NzlM/qA516uqNP0zzJmQXhRIPyh5N3a6JsWQx5reVkp9eGq
TU4aZREvetzrPSIvsK89C040e3sSLmsNpipZ8JNGRTiwqfHpm0wlNM64N1dtNdvg
k3MsgH3gt5Q/qhKcumkKRFU+rnisw11Us/I7YfiYFWLi/Z4fjrurZAjaxpWbwUXI
xfBSxN7Wi/gae8ZvpcYzWuYlHW6dk/d02IBvwSlj0Rk+YCeLKz4w1MMRU/bfNazC
a00QiXZ1qi9i28iRwHRheYXRp0BetrZ+Dq7qpBEJGuWzNjOKPOaOjkgKYp5Yp/Hl
36HIFq9JEu7JHIPhv9mHH7q4wPIbgYz28LCpj4pjw1+DnSH+7BN9mIwfPqdzkhaA
Ay9C99HS/KLkGGFG5FD5oxxcCRRhjhNYtlF0Jw+qAmkHx0TS5BvShse7QL9paw17
iWRhyrj7I22/1yEJiZX0J3Fr95KdEOdS3BzkaFr497OGQfpvQxkgATonh5bxTcXU
3UtHmuTeY7Y6pnKiHS+OBU0QyZ3zdRB2Bc+nxIIr7A8l7fRbFtLohkN1jHLrYfgj
Ychh/Xvk52Tc46oAJEyMeq6cFTpipyumi3lQeDZBXueYZeYhnd4JZZ7HHUiUOfra
zfYHKtcEjjni0B4grqKiFSqX8XNMHE1+9FwN3HWLUSCdX6CubM57C9TrEUAX8GY1
zH+5tq8NYgEvZjdRE42aq6ItNA6nHLRd+l5Isu2ns7g+W08AYq2yKXsfMxcMhlMd
eORfNar5DktEKLiIQ6Vpl0u4SJIh74vPkY2HzDRWWeZkRAZdLBxIn85csjXN4HyS
R/1FkmD7tjFyvpKaKIdS4qi//0ag4+nojTwlLN6WKIHnXjEbui6luUAdGgBG7JCY
waPgez4sSe1X9jSrD83adhQSATQvgzxNcCeoviwOay9SlBThAO8RXcu+Yhy7HdSt
H2x1ddRNEzHnvR1qRbxUpk09mTrwWG+d+xanvxfiWrrbZ6QDSVaiVmazQu8HEsg+
y54fBcWD8JWkVAPgY95b++KKIT7Xfv3zB41t0q4pfuMzKJutkXFyDa1nLfX5gVN8
BpUx9xoOQDvQWCV3rwe08coNvMFdHMzkibpWYlF2QFZY9ZOPmFYg4vsNr4Y5BfbY
DbtCqpxQTQXeOHnmBF5OXx1JAvj/SBiCaCYO09AaTWLRbP1EIAfRkWNawmVpdXSK
EiCBC4b3vYE6dbcC02tWVWJl/aRzBd9URqr+TGYo7tnDdHiL06AxSnAS43Vl1DD9
l689XBbtfFMA1bzeWXDoAWZvzz2IpBHqCBVlZtrFfLx9A7OM/niD4hYSCYJDvoLf
4hysc2wvy6ZciTHa6c2ob33H8CRh2SlI6CVxN8PhQaWbeV+KlJfHZPBBkyIVmDH9
df3qjO5ea0kawjWm0nX4MG9pDQwV1GDaH44WdkXMMqKxImiq2b52mp9soL7LHS1w
qGd8y7BOlZTfP5mMgcPOTDh5YDPfcYouCimFNmx0HrOTe4xPFrBRAvnNeKSUakri
KknZH2DWLIE9esPWyY0qWRTar0mZmwZPCxlwamrcu+JVbxTCXkurD7WojGATHWoR
whKg9dFqDfkVXL/2LQgNUueemwLeT2oZWwFjuYR8PJn0fIkaGAW/neO+ZtLHXd+3
uU7/hUjdwRJDO1lwqxTCdhN+cE0XbXbM345gS3ikjIUe7df/MOti8FPJohkMh13n
7yIEaHx/khVGhsB7IZbMM2LtqFDZTGYZ5I6sMZ/3MGoAOF/jWTZpeoAVpQO3q3Zw
eKH7mymhCdXa3lO8KeqE7NN58Jpc4wKb/JKPL+3ZzET4bR9BwUbNld+xAaU378xW
v2vt2qtgAHTDEg8+NggZMGDwZiLpWamwhHFIfHMclt10VJp00kfnnmAoiWk6SX1h
H+lHvgKDuUGMYi6IZE2WQ4CeOwri3k1ToCjJ5Qsuw2un4AB9tFK97N7djVFSI79y
4OqdbJyztAZVLGnWFGePwkDkpeaUltzpOCRYN5W+aV1+lomb0BLvReor+GMcMWgi
9pbSxIZDlIHAZKAthsLXdnVlQV8zhPHmt8dgLIB0/2kCkm61ZvU5v2rxhiCswM8x
nz2m/nSXXxjMAxuhlnfU22QdHNubyV+618ogonmncEBzFVV9+Muf1/T9sJ6KMtns
diDnvrgcdRohT9Q94gYZAq2nmW13uXXuc7COStZI5AH2APuE+sbXQMhAnUJF5GrC
ZnsDd4C/hnsPpgNS+adKv7Ns0Uqlgd6LyTzmapgjj42GHw95v2hYmiFlw+duu7nM
omw9gM1UDuf8g0mjcFAqyWfseqJxwLyyPl5lG1YA5dCRhCUOv1Wv/jBGB2LxxvUH
WPj/9qQo0oFSoJcz68xwdNyzw94mD2TY2sIOJPe5Bv0gJzT8WeAYjpnkDOshoK4X
FidAka8fqVyeV3jiUmyVOLcOe2VfOc90MvEimP1OG4x8gAQSC/Px9RLprUOYHkt4
XI8gORmJ9Qq0XZ3vN+xKW7JHpQYtUtnp6R+KDipY8SXSFizcacA2BsEhGY60nIug
s6Xhao3PbV9Tw+tYW3GF0EzjzY6hnswg8lEdQaaGwxEL+pSaRxuWWp411yVGrWej
eJ/eWC5FKHm49pajfEBwtHlHGwp5lnk80P0Sc4aOAzy0q7Tn89SyZWogsviaHxwX
G+0dddb+69iJdJm9+8IvQKgJcSm0yiXkWAiAhoAorXe4ajXLAAQlLgcSs8holL4E
0sieeV5fRjeQSldARa19rldTUwJyoYJbQNRPMlbLWlNiWRbjtySmK3t70P8ndasK
3js8ioD3SgwfqlKkCkgUkDdaQIc+bc2sW31iL5DLk60c6lSX5XeXw3pWMtZrZfrR
MOHExS4oHoz0Qh5TvE0+rOhCGIgx+xAsmmniGhikCqWaUyOhXd4UMYmj3TCG7OC4
vEugC28lI3LzS1Qi1HKjF7x62TxMA3ZoJMEXR7vOWRo9tWbWJm51YjvEHjx/fOUz
wnii3EYrbTpveOTU2A9ymq+iL4T/KK4uH+hPZutNPNvRZ2Cvfhzl3abNWX2sq0Ev
AOuALhqaGinTinZsu0LIgKqhkRxfdOd9i+Xf05t9swXdj/6YYY44sDFdUthfkjwx
9INFknPGxo1N151rUc0FiKiCrAirCZ0LKWDEJxwmKp6G3MeAI48aFteZHR44aa0d
By2TOryxCkfem2bY2jbeI0Iz+rsLX97iFPM51QCDuQYVxJpYA6vKVja6FsUE8maX
X5DAjlfJrZ6zaFbXucQyr4XVwj58g+Mxm8Jo9tR8EZVwcOubmh3SXJpAacGnOuV4
Wmz3BywTpIuQsRqZAeYHJeGqx+ovv4qKTKNbWSVAkeHqcBM6Ojlih/D95BgMBCHH
fQWOHquppt9VQsWwKYumCpDULm5N4exYIvSqgC9hMsVbTB2PcwOSae2fM0NO1YBe
Wn+O0JeV0kZSQQK0hOVdF4ELUyJxUjYcFpmxckeNyeFv5BE8zRcDioPgaSJ/XCWw
fUNfEJ3Y2kAnKbb2VuY+OynMA479wGlmRBa11dtMLv/tEYQXXn8LFL95hbNJrGhp
wCDUv/Ir7s7ZxYM5Y6Sqc6KxCsvib9Ya4Sm+Yfi20tEWl118wD8coUmXWj8GesIf
VHp4TGlkKxq0heE4TRd0y4eNXQ+WbKj646jQpRUAFuuuQ1ko2i4u/C3DG7TWsXdf
kxa58VaKbq82ivTXQ2N0euwVVl3X7Z5o0BgZiCEapxb6xHVulONKMvEdCoezC/+X
ZxhA/0a1k3m0CFAUkaTamE2mYle4vzGJJKXMdVH9JACH1D9FpYCDI+VFC+kgPPU1
y3/Kq5puuyn7nZoD7tzVJ0I/Y05E4qNAtDtAuKqW/lTQaXowALFRRmUBZdMJOQnq
SXzOhgEfXdR9Q869qHA0VY0Uwwg3pZ92+gJSDTpQmBfBH/lbPthOGsAw27iFqWof
0WsnKs+sb+zmZdcyQuTXbxMrhFIjxUHo5QQh7ptYCKM3WLwikO7c5FstjxQE4RhX
HA6b/cbj9ZpAlIAMufgLJGxzW11RDfVS6gLEFMbWBhin/wE7YkRj7uDGGgVagY+I
7wwIGB+/UFu5W0PDdB6WtAfcddZEnvmubaiA2V3tOHfJK4TPfmiwPJt0QfhNtJiO
no9QzkosAHaEURCnoSnM0YULbMsxDS9je0CBXsNXfLnR6zuMCIiGrgSyTIkan+om
oiqxny0r23Kl0As8ejh+ekOqRKjkqyd1H2OxWs1vbxZ186Ufg678+RSGW9Oj0fhb
rpaog2TjOG3FNV/czgax7DpfCmFQRSRi8WYIPJ072tqNUx9EsZPSmSxG7IJ/SUnM
ybaWTGsvziIjS3Ktg5YInIJqCiM9hYABQJkaZkNIZmh5SZk6otT1OBJfKsCVihD0
ILlqwwn2ZvBySyi1Q22HaZ4sH+9L7Hdm4wJQBU2V20tLNnUx/niiYaXFhJKE9UOd
gBFoK58a4Ibv1Udj0h0Sm4JLzA4lRqDqLYSo8pAx5x2HF7Pe9Go8oh41KIHmsDU7
8dvaKta3Mf5LVpitP88Cf1Z0K5XkJub7RkwK+F4t9ozCmFQ0cUWVTZPVKBFbSRN+
lyhPNtvYsRQNZ/cnWsdQWj0mhkj6hTErIp4MWgjIolMjB6JFyIghl5avA1lL/xLs
R0mnX+rz+8X8Un1hlvJ/2YPhSvufA+QIBMMcvMaNIJMUpYVPH8FbfVIwBboAxD7q
MCyuIX0eKb09cED1JaioA03QAPRXUv1mMjXoWYAKHXWkLu42IF4kdYFTux5NqOp8
sGJdZWrPQNcKblJh3cxIi7StgySXJG+YhDn1qZRsvBwV26IaZNjbrt11HU5G6OF6
eE/yb5YGLnBoR+1YO2L+CkymJYilvXlHk8QMOBmIjHYAJj+TIvqsdYNIoxi/zG3I
jvZcpd7dpQTldvPT4wXdaYCm1MmSnCrXtHE9bIgmY4Z13g/8zcJJBhpypjFAnVmi
+o3dVQOG5IqRCYto6Fjlfk/jfu9Vp8iDhlimJ0jLfgeC+gxgjmaqbmGf7rS3Gnjg
jr+Jv3nn5vSSLSE+NEVFe1IEt+hF1ElfXcrvoObOl9TCBDskDztPaTtNVQnpKASA
myYE6HF9gz00RI0hUNyFvBkFqGl70jMVHA2I5utuZjzYyTygMN/U/SdedpOSSjnG
eCl7LHcVGj8kyxx2WI2yDWM4EZNkFMWTz3nDZByq+P1GMwmTEmQHtitxlebVw6c0
FC+/fOSzLyKzC/Ozz+HkkrjEXwjE1DCmSu+vhIA52T6YodhtEOTWqAJkvsU6Rwcc
Jyq4FjoJRu2TTMW5Jpbp8Tcbs4G4DSknDfTo5LkEpmQbRgC6GjKj4+2fPFMbEDRc
ujgw8ZzA28o/ZpC/18FZnfQXt/ZvrP3PzkO1fZB6dA1gBQK7AbsIrAaYP1bT4qvs
UI+dc3CD55s+igByrNzoD+hdp1E4SZP+PGYeeUDUKYwfoKOf4lkaQhVVRVmB+ZKy
NlEeGjVm9K5SsKPXDBVTEjXI2Uxk9qFUUGpvU/Ke68F9tWjE922BqtMev98QXZfu
bmE+XJbqBt7ch9XlN9K72I8KtkfaCq27h+dS9TfW6Tb9tuu/iDcSuHdgMLkmubg0
S7SknGont+QeFWJQ38MIAjnU12aXnjd7OuuklkktV8ENmBQJG3w+X5O22xisBXk1
foPgb8H0w/BglsCjGDOjowwW4/n/UIUjFQ+1DMoRwMymDseVOzIt3Feu+TWgv10Q
Ma2UYiUxbZEA+cdkLMOXwOedzf+fTRynNuvsTDHosUlr+lHtsJjS4dKUoke34J/u
I2zm8C8YlCO7hs/wkvWdrMJODWpWuMrvJ+5LnpUENXDRWKJPBoYZgzVX8BH5EDor
Yo8XG4Uq5D79Hsemdu6vIa35T31/GA1sBZ9iEY33EK3646iTzWqLw6Xkgcqs/za3
MX0qBxKtLqAUkoWjE/LrinWDP3Myzcaj6ftpxrem1L9KVRnfPx8ku8YEl8Qx3U00
xib/p3R14GlZC7Jfbpz5bzp3+J6dlBRPNPnAP3hvyPgN2ORFQLFo3bvvJAFZ3bTU
ywOXuMxRjJLtHRzxyDlqbvavzt3VMwcPRWuNFqSP5dufe4gcb5m8GB/IBvkvvpuU
zpgccuXxh2+C/0xb53NUS2FaUyzoIfuFiHH7M8jIGIfdsFtVZKPMsEnCi6Ac1VV7
c0843hBwV/9iWRT9JE4MaNNXQUd1FNzZsoAMH+R/pltAO7ht8exxJXwxZm2loZnj
33CnExJQIsUeFk3kVv8CyLjwxDNXmMKwpo7oCOxCBDjhAmx+f3AD7bzwWDhuhhFi
D8B2GuMkaGdaUIwN36/9TmFFugs/FmOgY3N2o0fzZg6aqPhLSaDrl9ZcaEMaiiLL
yx7JUoCoB2K2WlankbiJlz804yDjAfstmY1P4Cf+LlwsbZRP27It/uxMAO3Jse0e
De180wYczZGQnqnRMIjaL9pxvWMTPVhM0UoPNpw+NqCQ9eyBf7XyKfoi1tTSxfyA
gv64hKQXhVUCLOl5dwOww0MP2l8l+AgP4vC7KeAOJj4KBpgLX0p+5B+7FuinCvcR
Bg+iG2wt1Og8xCHFIzRwRHflIeeJsldl0Sin0bRshzvpgOtSpYHYgBOVw7SC+mF3
LhgrOphEbND22b2c+odaogCXy8sow+LhVODZOYMwgXtPcf5u0tkRWXbkpx9UUuax
8Epx2mMa6Y7vIcHKU4VCfD2CKFy3vJnq8rX0tuxvLtdL2/r6lwKSt4gakFm3ptJY
Q7AfhU5bmgU3huQwcUFxiIo6HHK8KPgYKEoFOHSoSNzdmjgFSyh0JsELiS2PahpV
BmsDhMTPOTBd+BCWl+AE1e0/+RW+KBJA+VcT24c3zfmXMsHWOewhv+sYl9EBxxsg
03xY636j598NDqPoOMuRmj+mPaArJC8A+8/aK5nsobr26Bqioh1nPmGfLHQFQon9
EhqojIAwTfcOQ6QNjBVtH+19Z8RFWN8X7yT6FtuthJJHBM3qmwzyI2JBlUOXMnYs
+tsyWD69YMaz22lHjxv5iiIrNbKrchYbVAdAWVjF1H96dVx2rbGILrT54bUJ1N22
bJViZu2JnL6M0fP9W7ONPhbwU8AxwqZwoTk35zRz6yxBKkxEp4efP9MyN+1eDRzu
npEAxEnzeZn/3lNhntYoAku9fuZkEMlNDtixr5OYwZj8t1vIWx9xC27lmQKfq6zd
ONoNbI4lR7ft6Gr17xvGShFh4RxIHbhLwJ6sNKQlCt7Gp6VNef9va3OHhzUs8qfc
x9GELkdWhD40aipQn1nq0E+R/sJEeftrzBF4e7WJZ6Dev2y9n8Uvl1ImYb0LRyrG
3QecWIO7AI34kx4zXyhA7rZlNFDvtFRsGwdI/sviIygyN1TUhJw6kJPk1CKdWw67
Oe4tR9bo2JyGxVvAdUadVWMuD6R8qxgOIZQBCP7WxdVrOZYFsIrYvrgjBJxjh0qB
Geh2TxwXunN3LHtIdyj5xhH+I4NiVpIZPr/HVwp2616YdJr4JfRt6KMEhJqCJXyo
N7KDxUi4QmqF9Np3AbC5HLlsfsu93TqLhkusztZF5Q3ge0m5FN0SDpyRDlt1jQQX
rqLGaBZJXk4l1vsK/pWHq7TKQX2xtxQtpxfbZvlN9xv3jTKIqy1dbPls3U2g9va0
Txsn/375axSdU3GJkIxIna6W8FvJCZBpyNh4FxD716arg8nALMZ29F3K5kEwvOBk
bURsOji42fqDkdeMQAyodk1jMWi8usgufjoJ2nWe9jMCql2MHAxw9rhAUYk/xmtL
vkWsyW/BERCcqAfs1PvXQEMBXU1bzYunV0QCwaWCw4K4N4nFr4K5EzxIAAD/Jfr7
vDzoILqJbeQyexQ8ae1EkTilnFG/XT4ix28XaBlK25KjvvsHMzJ+39IQHM9jvXY+
7/2pHI2j2ttr6uyy41EJ9HsPvZ1PNGCFxCAbD/Nu64dEYVdjOeuwVZSYC7BdmeI/
speX6N/9/7ZN/RClOzhgpRCa1kBZOlmr300oWHgjWMQZX2eRejvoFwXB1KskQo3U
udQ48xnm9XzKhVQuBUrXTQ09MCUwr1lMxXsvR0Zx6WOht5Q4MKb8VIJOPHOqaSd9
PpF6DfhjjjoRsf0ZzfqTms2C7jh2L9IRQccQ3PkTQcu5WBDC5WcA0RXVM362xDgg
6MC7sR/ju/L5keTKWX/FXF7M7QxDqa5ELthP9B1TuhRk7QQQ7HdrFzNHL/PN1c9y
QxbySMSUtDG2Wukox55EWh2PuBDZheuTAPL4DWUDHSKHXlP6gBL1S6NTkj1OeP/O
r1hbrTqPQ4NSUBk+2Y8lO5Y90wq7nXlb7hGsVaGihzzzAAAzotfVk1YDHB+PqV38
CluANeeb++LGTTxesDbTUs4rJlAGs52Vqx94+62bGe959xJAR/E+xdrQ0DyKD2PK
AZkWhe2ht/VlzKxMwTsGaiwqUBgvw7iOjRfDM+Vy8/qOtN9cTzgBYe38h9mZLb2v
cNKUfeYZwwNSzb/VyayEU8t5MSDaK9hp5gyUW1VQQ1gzMY+Nvir4J41U/viUX6hd
6E43qw0Be8p327p+PaLwI9LNchpXRtWt+ncDkbzxEFFXXzhU8iTXrBbPxWqxqtYr
DXZkF72Ac93PYwzPDRv8Do4zpWyl5mNh0A7y+QxjQZOS4/y+h4tYmJfs19otFIDq
J7U8JHMPoBFDhOMMb37teU6yQ/s4FJa4gqbUkPJmgKenTCl3fN8xqvoFYYWtm+E4
sVN7XFuRde8Eh620i9a9xS3Y5dk//l+M5yq9KbuP0QIg5CIylD6oyQWCmWieXlt7
osSedecZ6c398ChcjJnWdrJvrkqtz3yZdfjod459QS1Mmc6C3AuMUNneCYOiSjQR
QPwmPviS32Ds3foKsxT7n44ugtNONnqDbPq/nvy+bcPNbqboNQCleOS0MdrFFQbN
RYygaKx5soxCnloP/flWvqHZoR5i44oxc/uxqKzDHtF8PJqHR54ABknC2GzeW/CU
OhVYAZtD/nbffAed57H6MLTcVpcyC6898RqiC2XEifpLW/uhSqnulCWXHst6mSRy
yPX9HiajSP3/5nQJahZYM/W++zq39R7hDJUmavLeHG11/TL2OXyMCMKqJvB0hCIp
EXFPZ5SrxrfeI4ywXNwA9YudaSLekK6L/H+GrVLdRR6MPUzDAys17dJq52YDnvVX
piBSZKz6ZTzh7xgfRuK54TTlOC8yUFr0Ec3//AZ7NW35mqp2AjzjQr8XqttPrtU1
HNK8Wup/luFrLua0SpZlfwrvZCIxdbRwIgGQK4q0nQpDDJTR8Al12CuAXRrHRo/r
7uy7m9lNOZZIZOnGoqiDbBtiJ9ye08pkx7Gu263T32EhjXenCGWv0FZURSqY6Enc
2aph1M0m+FWxeUIlHtOXYbEn984GkhO6gjSRYITHOW0X57/Mik1FWudHHEGWelQ+
O0F7fKppEsfFaAkKjEcFPQRG6h+TDH14tPO/Z0NH+sHnR82KdBrBBf47ckGk60pK
aE0c3T0c3oUgqDG3XjoTlRvXZRlsbE+YmLSWaT1B2qx8MqlwvnCRZZ9hTeevZdtb
UEWk42K2KYeQrP6IK44vkbknmJ05YVbxobYQftErp2DuggX8PQMp3rd1d+Y4aXzh
UAN424S6jZaY98vtsyTgdLu68R0EpRsN2QPOHKM3fRmODx0D1x20kZs2rHqH2MXe
T14pFg+sgV8ZNIcAnrXUuR5UyeN4iR3ARGGE7YsV+x5lrBb9g//EhJu8E7Jf09lw
WIB4Q5/aixi/iuK+yMlFp9O4j+PngddcYlxZyJYhYon1dEMV+r8IgWNXeOU1UHUc
9sYCxNn3bTHaSEziJgQ+SPMDHn4RevNJ/XSqwmT/lE9OYr/0r+PfHOQ0HlYjdqVJ
l2ppyQRB4Qw88W/Zewu1eX+tHYRcsSDEaCqqU/5A4jmda4JaNUdI+Jn+Ogm82gOU
jreSqerBtEnLx0fXApSj+jcYclz9xsiYzUjbogsQRIilOBEDrltYJPELyub1Vf4Q
ues5/CXQGrTXSO7Nicacq+pkN8ICZqsrmjRLS1U7J2RAILsNMLSSiC0rh4Ni3TDz
+DvmJEyYmf11xFq2LmbyMdN2UMzWCAUFrR+5OuXmV4/XfNABT3HOi3C3LfQRFfCk
tXTSkaoG5Y3Nhe7X1EBoAxiYRL5mm6wLrGnir4eGZpnhXh51WO9xfjVhiFWL3Lt+
7q3FDdR3dbi8A1VJCig6r7wIOcz1b+KzGP6QVsXcU948ISKs4hYN2sr6hQQhq8nT
tjq8/1RsllQGZPx3CrnoAPPW3C836fFBmcwNCeq56StVkQic/7xggefdkZW8zo5s
/SWrl2h4cHDAC46wkR/tnNEs3uplDj/OGWFtTRU02Sanw5JYU+8ZyZ/MYWkuRxlj
Q7m1vVDf/wKUcECwrE7far5NlWS4S/HzT6yprRLRG2e5ogrVZniBpT+/fTfOGVhW
EleIHpQ/FMFx5iNP5e07ftlBx842wZ/GCyKpv0dD28w8RzfKruZRD2FYEheZKD6Q
RIGW8djWw4q+3wh0BiBVX74b2TKx48lXsMnNxSzz2Blkxk7o1G21leKntZWcZrkK
Hxy7+j5EnkXSyJDv5Exq9rJYaUv75wSPbJYYTCMbB8zodz8ob8fpVISsKNK5ZGFu
okPskwV2070FYzNLfamErUICqevpkXatqX4Geo3ZEFsmHoWvTdiDnonTvl/us97B
kLvJzDJDFCKaYZ5YcWJQ0JnWdvQkWTa16fJ5k4myoqp0GmR8MFhngOK47Nm3N1aW
QXPb+ooww9kPQa9sFzlcBPYzVxej7iZ7M7adkcdUPnJz+8XwgkqwKWgY51Nwrbc/
+uXta4NMUkibcYoBdHUlUfoIL0nQ8dmZlB+SHxwesLbKwjRU2DudbQRLGD/aGuGi
8hu7DFlTGY65wzz/xFKFOMn5oSaR1hCyrYrl6a+7daAybuwEtP17j0T4NGa/yp86
rHe0xvUy8vZ1PdXdPnITzBfbwezcQfmN0Rbd7HnRnnJFfU6imU7BJWtVKgSWK2/X
+ujjX+DmcLfCS6buEsdJsjT5UvCc9dLuhlCVRFne3qSWXfQ2ZVLVZKgMyjclucxG
UDfWankAIxCRbCsilGm2cGnXar8nTIJnpCsNe4u5NzxLQteUya8w+Olgv+fYaDdF
/olC4TAB3Fg5zFB09njeFc4j6kdMp7HOCAesNDaQ6C8nhgWOJ5gM+JoJ6rw9ZoAo
tZJ+uDIKBLOJ4vpoCM9fl5E4t4l3snV1pkGJbgSH8vUYEYBvhhTV7IBnMmo47FXC
TquD/3rA6Qu0C8COBK6h90KAQfp1Owbhchhf32zwJQXiSbxKAwIPp6ZdNjPMqm4z
Jpt8SyGGvs5EilNxRGoqJyKzJ4J4dLwzABF9cVEzQWItTh0e636hNquVx+wNgCff
ObzfZN+BFZTdFYKsOjY75QyP1E8HAJfhF/AY8Y9wN4y9EkmPRdjyFPsI/IvstwGM
NQhdfbgVEmnTVLJJhAPTpk95MqWHf/5S8fTkGkNWXd6WddHnKqWG3ewr/zFG4j3v
jeBSJShqQuWX8XZAKixOtzB9XcwZwUC4OHt987IwDHmeIeTFr+TKvWYqfxiKI+Nq
w2thrAjRT/lvug1nrm23Ydyz+CEaK/X2TlVpHlXbC1YYEG2rh23ks7xjF973xakG
3FfoJNkFcLwKaB6YflUKcMM6oHQ4RRwPUr0LDlVeyY+mFL0EB7eJh56suiw0DCb5
Cnf+dr+wyIZdxO9DFR9eLZeFjCRF46ysvyHB9B6k2nkTqYlQZofpUZIyXTWDMx9n
DB+uN5jqTZjcKzXvHpPq9DjJQ2WPVZdG16lHnuOF8ueM4fkl9G6bcZ3pYZHIs7Fc
VTuw9iN7DTld80n+K8jdvuQ2m8YfJuWhAmZk+/QJfSS4lvHvRGwSSsdtr4d0mQYm
oBZJE4WVu/iJP7EEsGnmPISpuRdlp48Q6ER2bujcRNMBY5JfcxAFrty1o92/u+oh
/cp5rHkKtj2ft0u0Lml3Hctir4Oi20iC0qjyKs2vUWchIWVMIU3+CkCaG07C11dF
wUHh4+zv/jc8v0NQndXOCYNkHnw5nyG7gZnUC3V2c66ESQ6I6/Q55aplU8CFt7pd
BRvjtHIWVVRj7GthaH9HB3Oxzw9VDmlRI39/uXMjGSZskyTpbTaS1lSwQscngYrv
30hcpS3VP7LUO5xJ7P9ElH0UmgVmL+okAIX0SVjJZz27byyG0+2byX2RLB8wwKQS
GUVhWa/QnQyVIOow5EgHqqk4DyB/9r2fCf/RppKWEGxCJ0IsWXOe3A4vElceQ5lA
LGcEWf4lDIhS0mP+5ayxPG0jrj9aaBvo0yFuFaZ777UJcPZKjv2xOVz+rQ37sZNF
NZUFyzLtxmdqZjqmSVJMnL+BifguChgnybfuEfiIqw1YiiBDFyAT+nqpmifhjrTE
DOB1aJ0peizNI2kfM/2rcRwxMXsbq2zkYJCryqfpgw6GRe6lswjCkrIshCpIhwaz
+SjPtZr9wHnLZaMqXVdZz3VWH4WSUQ5IUD4QWXxPLSzDY+4Wiy9BjUYjXk0UeEMN
nCBUeVE541dbTBobfTK+J3Nc7ggeXIgwzd1rDEJPAeGbvT9m/Mv0h2MRxBg2EAn2
xlPCmWkTaX9Dd2M8uiKUmhZy6jCIEpzKpBPNyBu1EE6m1WIJjuTxGpjtvl80I+mA
ppC5FOkvZM0mJo1bT7hY8bB2WG1PytojPu3ykR/m2qM2UCSiV7r1+1ZRZJixPD2j
CVoipxPSpd/x1jVy4TIMDYKE9ZJZdFXGzi44BsnjbruKsjw/Bb9zA4gxVQ+T8+bd
Nl5uAD0MaR1XSeQl2IsZzeFfMDZBW98zViQYsos5vGSn3BV1uNEAtFcvYY67238p
OzxmDnNR4YEqqLMIQ/Kq9+Hohc8GN2KesxtuuZKWx53ZeRiPRwFf43NMq3Bw8Q4S
QZ70GiFnJQDh+cxO9btznmbu4/XZLnF3HhKJqKHJPnWrlkpHu5fziSShNvxHb5/o
LdojpbHX6DaRscIS6K4Be3pufSu/kzTVdaRVMhCiV6pPfz/Zy6p29H49V4rFD0tJ
S3aLnNUZ+C34SEYHtKY3fxmUs+aYkPPSCVla1sTEINiqZmH4HWwoWBfIAGG/58zH
bbvCjO5OxjapRvSRpWybD37eY1D1qPKIF9YN0haaaThsM40EvhwHDbI9PW2U9IOA
2ru6Cw40HR4T1Z3qRZtg0rIwODmythqFQw/8GP6r/d059EWBwT/cnX6hswwO4R47
/iHz35wBgqMqj8eNn3kTSQcWS2hOzlhjjQ5zHv1Blk/LlKKMJ3bbKBxkH2l7f4Gm
B4jlODz/IS+Ozh8aHY0nBPGkzVc9jHV7BS3QoshDiQeIfCHtG+HAz6v48IhPZdb7
zrGo7LTN5DPrHq1RYkV7MCRic3sngJPp925tItoIr9NjVpgV3ZPPF323gKcG+v6M
2EdeXbTZ/+68L3O9+g7L4Q/UfCYliAr/t2YYNGCmXkwIWxBace74CdNrO89wscdR
lAF5UQtNYC1V5tXeZA2RZnbldX5AR0GQ/11PW7K9t0EZO2/LPVq3JbVtHNxMWu20
NAMW6/129aNH6Ns4mBfD46AzM4EoCrGI866kUXhljEFJDOk7dRUcUKJmY0kuW4o7
uFIx3CAy8ZYosXtz3bvv6cwLbYbQ5d+KhZTmKF9s6bobz6Xy/N2mpxab5nrynpco
21kIFSlCU/D35RtPQMNuh+gg3ejp86mj1z1FKXE0VvjiKUsAE+6kLqjz0fjbis7G
XclSK6+yNuvSzWVgr5h21KToDhpLYhCvUZU+nWsuutEBdQsZAR8fUtxSomWeP0eY
9IKkZB+fcOg3gOZjGppHxbmTrZ37Q3L3556/dcbV+YPd/Cl2ER2XYmxzRQkgS+/M
bcNwZV9kxljGFK2wO5wPrU3iMqYhEimADcbm5RUFA5CVsScVwWeMibsyrBX8OFpP
GCZiTsQMWfVjxOKcM9umiEIuW0AqomeVFLPLLnVlF2H4l6ahpiOpJ2qLwIfcMKlD
dFJmvINXHEND/lqE0pdFR6BZR00W/RSsHHWxmWuzcnSKY7cAtH+r49cAwuXoD+7X
aeomsEHYqUwvyBZ0CaB9iTZjjpMYXYFm2aD9B+A7/+UN+Y+Ht3yom4hDLbI0mHTM
IxvUJ+f20E1uwwAyza++wq8jz7bbGCG84XvOWCjOCmjovHxOKbGGXogoIKliDPbc
oKYwfB2F+9iV0EOvVr9IkI5hdudWdqTxsdivHK/b2rt9lmA+ZlnmOOeA3CMo2NNH
Y/FsUSnIJzL98hN1nwH1UGEdOABZNoHqPaBc+1fdzrsXZR00v75kDO1iUK8RO25G
4gYOGHA4Sdu1ZQvE6noFiAMYgR6jPWzRXLoYjY5S0IL/Rvt4Fqb41TqvzUuwsUwC
yJJPTTUpHjjojzqr04hiP9F19vODQEmbSqZOPUaGUqnffFVybauT4KczCdzHUt5w
u0pi9aLy04aRz9MHsdSQHY7R3Ofjiotzrh9gqAW4A30fwc+uUiAKnH9oF3PQyR79
Dl1262Ip+Gord6HswWtBIIRQ/Amy79nwDho5m+9Tm85SP5eam4ZjvbeDVkLJp6uj
Rxpidn1jQPWz5x53eiJlmJULBIMGaN4Gu62vNG24l8H4xFPJGmBZGASYWS0N7D9+
sZMLa6euKP5wvm1IGRWBlCHfCkOPkMivHAD2K87Nh1Z/Qi0SZYeTuC2F6gJfklwU
GQ8nN+6fXgmCq352kpDooNl3V/OxkgkMJpeE+fWnM5Efl/uDil4alWnF/U4EJAht
sN8BFv1HcBLM20cRn1vjLNtw741NsgxT6iwbIzW4TNSSotfZr5QqYquLYycyuWOh
F84AzdTwbAu2Py8d+BBC9WDfBRWRgA+jiJIECBE/OMQD9r3v34NLCJIyfVi63Tkp
J+uhAyQL4AtBB/clzXDIALw8+itLURtPGmwBwEICeDOzybECVv5zGY+YGwcW99rS
q5+9XcI6b4nSxAtaMZLH5fRt8iTCiJE7Ui38Mq/3VMpV0gN6gYH255cdJa+Nei/2
M9K0mFabWEDP8otY5vA0AJ/jJWBxaL/wSK5v6kv7nmAJzpJ8+Q4fzD6/h/T2W6aC
pjwKJjjsVWjbvUInfTMYBfHyJKCF1DHJW2GROmbLfax731yatg4TQQK9fivoGkQr
n+iRmmCyqcGnnPoAOau2NXSPFbxzde5FSqH+kx9oF/HsqdFaD6s8r+8SIXzl9iQY
xI4gWSaRPRKzMIxGjF3FZ38qIyatK2DXCUWWcLM530J1y/E8qhPpcRZUkE3TCf8A
EJbC1O7s1x/4NJTwuQCkuNN1rNq+d4pY9PPIZSoav1ANnvRFV65p58h2LmxzUV2r
Ut7hmUSoMhyqJIpcDEGS3wXgRST/IGLxnLZyt46oXcreEQrk1WbErdwFUkr0PPKI
aiUUxJZrhMrmcANL13HEteBZA0wh1no/Ow3OkIrS9U06sCU+nZROYzuJcqjRluF6
90yFXp8oflRIYAm8z7FMkRTTdKNkUl6q5w1rvRaQvLbDSPOpjSh8afSprvlSTql3
UTWeL/HYxB7QcamXjJG66uC9nOj60NYXoJlBg18RVe17FoaMeA77ApZR6KP1cHoV
G06ZnyHRYw3Q5Mh8sbjnCW4q8XnSbSGzjhEaaHonmPqVoq/jYQV7BHdhssNYb4fu
QFfMjqfVlFXBzj6NFtBPrUj91FMVuVSMu3wc4wLXYYWdKEI3VIwyV9ZTtN3ng81T
a7FrHW8bqO5xjOUSCZXyQ/2nLZJsVuagk1M/+1z8iklK4bOTgErJq65eun5vM6ct
ZhHkOsxzacHe7puigHxxEbmWW/lqUbCMs94tMEwktQOkRsOnM451b0OtycUhO+3s
MbN9fCx8lc0TSDlLTJPpNiMYacSk+d1EFpaAnP3iV90acRCapGydAyjK9UKjrNpF
G3h/e0uBbbAUoNGjlE3LYd3W4QCcvSolbP5bF+r7aWesiNf0gGvGbIIZY0kxZCIg
Og9LXYOtikzpqAA0T+ikvORTaLp86Mg4yoBJD5tCHibzNXh8VdBgvC8QXZzgiYi5
4iqCAmTL8ntylMMUlPIpv5sbzOu1QAEDZhbAjHRTPDWgwCOYvxnADxIp8TwHIKnt
WlWFmNLoNxyhPnjlelgqrFzEgwJL3rA+tWIkgsumD56x1HybsQuQZKrwqM2eLa80
1BSGZNcLwMyLGrLkvD4VbATLvgBkjCC0tGidD1n7Ljlhm8iyli4fZDdJ04veaIYG
fntmmzEDK2/ZL0msyIk/qooam+E2HoiUhgArHWspz0HUeKvQRBVEma/PwZb6vIOC
ldPHv6GweRuYF4UFzdi1FUhvKFu+ypZ7u95vrFwK4O1yB2BMAuEucC19J2tD5lW2
I5Z0NMd1HU3rxZ5B7Kr3X+vUqbSQqzTMfI/MTmxi/x3a2o+e4W4DSYPwRBklTptu
eo47hKbVX23XovXsqvWvwmBmnNJt9kwRQl9/OiO3DD0hdZRK/r2DKGT8JaZCHJ/O
x+NUzUYpVWggDBKbq2zWJKZxGQEt8zdElOASNS6Ezx++kWzvokuKYmJGRWFoxrj0
keGRi294GYUVfxksmGFcuBZLNcULjdzDmUshfRr2gwpVFBIDRoI6L/XqESmdlk0D
X/8qA3wo8k/BNthG5SURIf096+I5IxtdfKnOFu2vWO0SpDkwzL/zdwnOHVSIqsQq
BxTsRNeU4Ci2hq1AcaPXmBm3oxBXP/4DO04Se3Wl8KzLtf5xfksd3StEtQW8x68/
6tQ7mKFBUmw8eUOIkNQxKAsvQt1TqOSrvJdk/jKxyUEnJWBrh5Rt2uAcqZaLGsxA
SdIb7VzYWNYKMM5iLI51lwCac/xHzl/pV1Q8DFHeMmon9wKyk8v6Adrx6kfpFF2P
+atiVZJ466idzs1QKiscrha8rTUuHloZzcgp3u18JeQXn/DGc5WJQ5ssZfmaj2jG
Gf1KJY07dRaGDESX5xvGe++jhgm5VcGtcpptiGCo9Hv5ByQ6C1CQdqMYhVMGykIh
q9B6q1J1phw6CCzzXnmXE/As3j+aKVaSn6sRdpUIAqlTSsHSi3PunfZII++hb3yz
hfGOEltIb7e/eY6fG3o81KE9iTI3uLotlMorCD+m7J1/gD+irHhFDaKmIKpqwsI3
Z0kOH8ubXa3uZ6GaaQE5RqGBOJ7jV79FrL1kQ4yBxsN7UKOxTowE82VrCsCh3qL2
6FLXkFejGDIonVyhv+OLdHzZQZw9qFRuwWn1uu9p6P5ra0U8fmWn7HI4KVqgSufY
593pjYKBfAzTfh3EmI7u+Yl6op4evf2U9f3Apkl4PmmKLOn5qrJ1Iz6g/ZKna8bZ
pA7DnxoxLDmDSTOZvW3VUM+dZl16MVC+GS5ojhSnvGjCU5yrWglWUvekLzWVmpaJ
Um/H7BmKCPLwgSfRRPaM48hDtJAkeY/Ezxv/R+IxV9XmTgMS8b/19bGGf0qmo8ZK
i4R2XrbXhafscniLPQhdXWBFSjRhhYmYXjIaLjWZqwHE6Nml+GoQ4UYxKc7UpTG+
0SJno4kUK8EIqdIWTLXDzoBo4fOlbcT8/YB0VrkrHc7VziEwXhlxtDMbaWFnCz2R
9MSwFypVf0IPMLUI/U/42zWt2bXC6oz94r844YttK3VzYGn8BSVVihQgrCcDW/AS
jOuJOmaD7x17Y1EUO23uuB8gDppTq45P0M7HfAZVq7OvnJno8OzsGnJ+cscaH+dr
W6BVrnfNEhpruUdYaiB1OQ2bwSPmJgC4jaDFVFT1PtXIvkZzHXBc0s8YTQoXwlgi
F0TVHi3RB4TXozPl86b/tiSvhMKKpQ6bhzaI9S5jAgWHg+cyoP9PWDJveYmRKDWF
A5zk+ykHwfBgkMX1u00ZOZYuAe4MG9dA8SGhz5YWX3CBTTkcfZ9BIjsMJetvV7i3
PkazPiRJUPCqq+hLf0hIV7K8JaDlTZiWpM3ZhNSxbCtlWYihqikDdWvFGsnbocyu
GKvbYdTIHhFii0FIZvVp07HEwePE66WB02klvsO22V53ohayzHBuQ+XecDzyGu5D
kXiIH0aJDW3D9QNm2rW3EZj6sL/8xDg7ifHK2oTyM4Siuhsyr4LvLuYVPrRTBHsT
IocMHLag3mKYfNIzPz/cWoPERUe8OAJz0Z1p/irFXKSOg3hCrHUTpIIDezmY+5BV
4UGIcAakDgfv8jF/tLYml9a5OU0XrzLPKEJLo3TdFXe3f9t1wKk3jIb7/KfnJklK
No6UX8YzBSww6kY2tcUAf61Ps9AwfDDdHzwy29g+7hvZtgVOpCEnqAE59kllyfPr
20PRRCiA08Jt81DCYNni279umYwrb1hEs8CxlQFzNmtke97qZMMtizjSg/clC7PX
1yY8BzeKgIME1GUIc1XGYKUTKNUk7b2f+TnE0Gvzs9IL3wh0fr6ZvGVtDLtUExZS
Q4H3ItQCuTGrRh7pmO/hVUtQ58ofET7lnw1oihIXaa+rNuvFGbK2fhC4/idCTrSJ
uNTuoe0e8yVxEvJeON528QFlMG/5v9xmRhTpgd8G96tOtX9X54JZHOFpUP419gzD
alSHb2hkEFjm+AXuiVNtVECcbNzlQJ4aE208LyBMzcCrdkR/uNUbcAH9wMZVo7ui
kOMVgCR7pbhvrWPcJ44CVkA0xZdcdV16A8XxhYKCbfksmQM2hOORbQyoki791H+/
2t+uFzS1+WjVnvjycGFSi2+8WOyriGOAGmSid8/744EtvGYNIF64fWYtulLZoTT6
RZgmEeekM/5/pdCzO6U3n2YGqhIueTISFzMuh2LmFbERp0oy8d8ClPCfw69TAoYG
6J1jfHt9tEI0ZSmidqIhJknZOgi7Q8aYQbGHDlCXo8nPzo6fxgsdJO0swJFqTBUJ
GVREI+t9wmynDlddcNhjPTPkkTmzfkqVBBv7GVhAFdlKW1RtHyjqQAN/J44PiTVg
DxvkxciEFYIxTfWOuRO/B1L4w+NiBcp9C7DAOM9Vb486mvTN4jp/FNGG9MqjO8qn
ltiVHCtKbEDdHB57OyIbf3S+TgKNqqfqWaakwudOJuGO+swDOpO1a/dUL2Us81FJ
0EsE38WZ0L1YsU8ow0HbTdQ/Qvc8JYi9twn+dAJVOjzRL9lf/xv9qGRNZJEFNQPK
V9S49YR1bCYy8RnKOTptCncKdKecKJqwv5VvLoieTuZIy0VMro7+phM35Wo2PtzO
7zbxHdbV5Pv7XzCE+leTADUMcMHSEHFaSLoKnhy8iFfwNynTso1lhm6DKtJwNK9P
TVy71erhjfGWFx5Eydx4dKQAjmdzjseODphXDMYSh3bmev5IP1rr7kLP/nzVOpOA
x4O/ec4QnbIFRR6fgoY4ohDg4OlCuL9RWA/H6YU8Xr5SiHtvRxrl6Nxet1mjSoX+
PxCnZNXfKjKbkFgQTQ/esbB52FsTO1/qhU0Hip49iT4TCLKsiV6j1D5x6UwvX9rI
PmA8p5BPJmGHkgnlqC0idd8qGGsZBqTRH/KolTo13c09LKKgbAXSJWpfQx4/83q9
ngGYtctcTxVMTmKuxqJLbrcWclaZpAOXL8jUDrZKfST3LXNhPiAYC0Id0QnJBY2e
rqfwU6zTBKUEQ2i/2xJNyW02hjxaZAZXMBGbRk+HmOj5/bWdfX+jWOXebJKzQRCO
wRkuObVUk9HOsChp8hSlAlXZYGTCu8FSzXXBRbd5lnXqmnl4rRG6TTXGis4lrR1d
ZdGa5fVcOVV5AmaC7ZGuDF+d9nBvmAhjns6xmYrOIxT3I6hMJTadsZwNeMeIzV1l
kUzc6mDqvvPe1wK0T5wXgJkT/2ECEzwW6FExUf35/MV10WC1VC1zB09E+KHE83y2
vncYx3QwEKCPLjarAouCvuSJar4bwtQsod5VqSmKF9qMZUmsW/7+YH5VBlfEFVLv
HoympZhBqsyVDWXWiTYl/rTrgXFlC6ZLsfxqc9lzW0qnkTw7onW64is1AyLSPj4w
P0MrXxUdmcWdtkjBsc40GbYk/UlJEthG2K4kj+nxjQn5FelVKNIkK921NMYuZ4ry
MeH7GHoP1Ax1eoYHSZPT8owgUMwVeKHVR83SwqghXerrRok6YjBJfVW51QsHV019
fytZ6eEhCTZIKaLhnP9i4n7qVjDtCrdytHgiqaOy7Rg6/Eqx9Es6XsEeS28QCgCt
j50KprVSQ7dkqDxJ9zo+uXq0SeaxfhtjyJ9qfk5P8TibdObWF9n/ZUBD8JgCMg5V
pA34u9nfu2i+0y4q041H2fLpuHwBD58OVog6COPnHA24CVGZtB3VuV7G55wFU0+r
dTP34EXHjEw4/AhvtwRyG3OBXVKh7voAHCkMftzKLZAcxGg8FYkUnX+Df64wePTZ
4OpBl0Zxma5p6vDxejSdIsoVsWdg5ayCGhkhkdAUYl9SjMFUntOWMRC3LWqUWJ3p
vVy0Tc2LNnk3VA/yUPulNkklMrTzl4KCDvTkyCyty0PfkySM6XE4jQDENvxdkZbX
l53Hla1+dcrJOj1cMWGQ7eg0HvwoQQcnF137REcZ2uPCgduBMOu1gpQhMPmUf0HP
IUuz+O9/mU7jJP0SZIjGe2pyqhXJbxVapBqcj2lrlbXkt8UULrROkDg4mGa9HrVe
pVKq3kakQuf3QaZafjgnUb4upKb4SIM4v7gYfAhPd2VTkdCrqKldjcufrigl7al5
cYccqG3X+8Hn+69kETkSMqc04LZBqV+UsAjBw0YLRX5NkCM4K7ELrAnJMg8SJ8vN
o9NZXO/FBjA8G69+hj4Am+EkCNQ4ZDjquUXqjLnHbpEVFQwUOUncypyox0rPMvqv
IK9NPB/1AhU8EqGGl6fTCfaOSvGcL4qaioWnUXP/ZBHXJ93yUiQIOKcI+RnniMWZ
snbMk9cSyKWoG4GIu96XKiTUmInn5IGejc1vdNBFTfXHzLcgeRNjVoUwWKgKZvNt
zcpitvgQHfJR8DdYrocqsu0uVBjqqFdyxfu6igczefuK6XrbmcmFRlBHsaWF0gZG
UQKjHiUEe4rF2lxY4+xFFav+wlFhHlk9kv+5PhDxgT6PNkh0C1XxRube2SHTGBgI
79i9nej34ehTBA+TgBuuVBMEDaqYq17srz03wwgZ0n/f8zXJh52a2eYIdbJlBMN0
QslK33uYy/gC4vgigfbpF+YdePmLWvM8JfQz5K5bl/PA5o/Njw0SWJZZ2padAvqM
lGmG0TNiwAmkM/QJZUEotw9d2BOPojltjIF+FvX28jHR0zC/XyYr9x032lUJDjNb
7SloIHrOaQlAeDrBNH5UDWvXJr+72WfjRSSOaXmFfMd8oQ8MFSxnyy92OSyTAfZM
EYGOLmrU2fSGXpkZSy5jLXtm9CiIFhwl14Jp8vcnwHnY+Bh9bnXawnZZLWPhKvnV
MtxTc7Ue/gSBZzTAPx8HfkLVgr542eGlSVr9aSyHq3oWVFqnd1zBn7ZcPv203TeR
xUvIOY7C/5Uhg905FzhDqUvdWsdom7WytKgMTjhPRBiBFveCjFVDlkJMnSTgqq3B
wW164TTRycNamHvkd1q9VJCnWtgFndKWnzJcHkopqnsyOkJcnEI75+y9kI57h16h
7cAPHgg4GynwGMlxzfcbwqNZGFQoqUZKQh2GP1uguXBj7ZWQexXXXoRDkobzFM6O
MNYPO0h+XzeehLOv+8bVVW6LQpIvlJSlAySx9DdQm9DKOCLEgAC5lG+Eu3Mz8eXl
NuOATEcORGPtMe2S0qGhBRIqWclWoS3IHPKKmvOMI8HFAFHW8ebX9my3fE2D36lC
fmQVTvNTZzzb2S+Zy86m4quMzbgpx4ir0jACrIU8zs3XV2D3UljhIXPRRrjYNxx4
VgMW+tJgvtkq0UGJOorB+6u5hAdSR7TDNXgy+VQJzlMzg3F1HD8V0jBh+Dv08qDh
HDdrshPC4wy+nhzGgWAV+aN+Zy5rA1LrpQ0AnhP1cLd9DG1BYZWEPgYpJHxu6dUT
Tecr0MjCHEF6D0MKeF16gKVjDj5qHFZDBBucpjvHUr967CbkzpeALX0svXPzq5dq
YjVi5hAR+CYDQtxVr1bPBD5gJZVOx6NGE3jMxfE4VLah7WlRN2Bpl49T8SBUpCkg
RaTY0do98BUMcGW2jO4CFPuPjWa/zNPGW26cwtKpyR0Gf4jNn453V+2/nOPa4vgc
EbCE/bSiQQ7Ee2A6LIJed0kHkRm7GtCnU0UmRljgy+FWPQ8hTVYPVkvGLWJWVKXv
NbFQfUfxSAwWSUEz+hWLvBpPh7fHitZI6F/grecA5FKe6X0I+bEOsMbmOTCu+nhx
DUA3Ke8WLJVSRoqE2Ju3GjlLP05U6LiLK5sp7PCK28IjrkXtxwDM8x2DkdPiB1cu
VHRskpU5nrPt0UR4Dr7guj73HhODu5bS1s3HirWsbD/Mnbok9tDAjr3LfoIubfEm
UV+jVgJi94RsSH1WPt2Fr53E1Var5b86DkK5lCutFcMibE0EM0DQVVCNIvSJHk0R
wlGu09EDXE37Z+0B2Zw9v8+aD3HSY2h9VzZC+ZXWBonyv82clkA9PuHIk5wE5ush
8mycBXAHuyNNXZ3evmhuCh7syi/6/XnKNadoq1Lr2i0759RspbyOf+ivd5FcORky
ywkFdxrZbPTuHc03CtF2ZrqdzWjTjPZk9cYb0v2MO8N3k+POqxvZvuLrABim9qos
3BQuNRdoRP4sUf0JsjTXB5izCyGVmcu9nqc6AAZyFIr4o7qREuD68rMmKMBUczOQ
nZ0QdUUvdbUssF0x1/IKiINPCLYNEHXo5dQAQj3TXrncfHVeHVBBYRiVX3BZdKCc
VoN/6adTl5/Mnnl9g4ODnq7rOEPYSyMvm1nJ8P8dgJmJp/netxVkvFKYJvp6v/X9
kBg3PBpUvXCDRUYzEBKM1J12iHAYSN5ga9KJelladEDcyox+p93fU0iwsWpuVNC6
XBcvjQUxzx2IfWnBRMbjhnguEn6D/LQHVkzD7djfBoez+vW+nHH6MIloQ6fMka+D
SRQ/aZ1DQ7XSWwnNXDpJ2kOnNeKmvsIAe/IO2EhVWxkzhz3tsbC3RssW7oRuB+x4
Qmgc8UXYVxD46muknvJ6gnKoEx6XRtLr3HEPWewlkEu6DdPtKcmR/J6/If52tIDm
buWHHlmaTPhiKYdqNhaXWf2+EyX1Apxx4u3pSFZB9C/VDOcfw6hITN3vJjccRBTP
oVoS8CIiNW0bWmcRwfgSlk8TAAdmovysymS6q4h8Szd28jD/Y+k2L36g3qlxM/wH
afWWLHaQrDwJCEf2L6qayn3HDUqSmUgdEdac55pwNpdvLO1bve9Fnxqd+sBGXZ2w
B/qCaIRLQSP73K8hTBA3kbW6dasHkRIsazSClemRgA5RvyAixnocyWMcnjPAhgp3
JIVE6nXhFgGAlWrVO3nhUFtaCdsO5VbswdVbBDqk1LjIjCWzWPlLSUKubVUVVy+6
cZEnujO9t5wbNTH7Jf56ClVLVU4J8Mxh8WDqyYfIMu5MA4QbkoLd5s5XJVzjg+y/
k9Zw2+Wr/k/mvxGa/4aYRma2CmRfQRWRoYIFcQQcgjiZmF/HgL968Y+ejf1iSU2W
iHuQHI6GnKY8u8p7g1VfwDZikG4gofSqEDRM+XYCLjZmQgwYDC8aj+L1NURJPJfZ
P36RrotzXcMwa9E3QiFUEJb6uGbvj8LnIF5rfuSqwW+JtqaNSi4JW3+Kxz2/jWPg
RWdURZELixcIoeCC+Q6PxxBTgx35CHL14AocOLnnYHR0ZoYaQQQwK8Yri5z4G23E
MOls+t8zmrRB6lP/Ngy/OMV/oP2MLvf2UVWJbsRxQhcbb8Jqu1y8kmJEkSZjxZRG
AOb4PT9KABMdzALUB0GbFc842BXGvF7tcYwU9JQqgYgOmeLHgcNaCTG0mVLW7fTa
AF0tTzoe4Y+TX1/i2i6XkxiomAn/3DoGQf2ZeiXeTkkRPJHwuN6S1rxSHw1btSc+
PUOobFQwufkbTvwwMEY/rDGlX3e/TN7jGLT6EF95zStVZFczC8Hif1m+JZnxuOLA
LDuff6i7IiKqCzfgA8GdEa/h4hOdPwgU9CgU7h6jOH1PBOcCBgKku75t2w0r4T1N
liHduoUcdjrfFPxhBzRtkHWof8qKMpP+PzHIvBDGi1tfDR+oNr8FtPPfL/iKiJKT
XGhLl+A+r6d0tN24O9skI7X243TaqCLLfKdzlTYVPCAxH3o2VfUlEFB5J2W8hkAQ
Ny9iSVBbCIkXgoqkfr6YqFeky5CVNCEu67Ti9G5zik6d+a0qi5k4lpJzhySpP2wl
WaTqk7ZXj7IT1mZT8rf6SlkJdjX1g01r8KXiX0NFF+Mal7DsOCehKtBAKHBaqohv
4INWAYDztgVGz7/+vyMH2xVGvL8tPChbYzVNj+2pPdClsgOedMvsC55tBbQHRfi4
UyIl9kAHp5QU04B5detjPXOfTo6DeE/LOakkm2O4ESq5Ur1gxOXFwS6GSpSDVY3q
PzPOol2IG2u9vIWDyERiuJAMXTgCsGZnDBezbVfk8CC3u4kbU00jgRNagBc31hLP
0p0FguSE8AeUo2X98RhNhVEWTbrqXi7oncOHsiYdVlmq6Tjn2jEF5TpN1IDiBtF4
JnmZU7+q6qJR1uc7k7ZW10c/63Pl/v2TULjfOUNP4OfjN6kV4tA5n528gGDXyXoX
tUq7Y5ploqa1T+nLnw0OLASk1EMZi0HPwmQTLq4VEtqtsvKYGPaY5T9OJD1lKi+c
6FyHZaszbPIbE7CZLSnCM+0CGBGVmrWq6EuN6PPRT3c7SHWfwX4ESF1OPzZ00omo
2krhzAY//vUPtvglN4rfjTIsCZq+PRo0qvnZ6X0C+HKWQySjGj/B+JVYQTa06e2p
tBdl1Apphnr0dN8pTxUUKHd6Au5AG3xNqWnqjasGShfCb9cY2OH8dO3W9jT8Tfyk
MOeI9hGIkFWUTaXIa7OWWUOQmYoYgf9LR0O3tXLDBpT5iQqh++C3Zg6wyd6znWP5
e88wW8tyVkgwhma37AtqEgqyyjlHwXGnzrzyC3dHnL4UgcM8L9cAAT6DKIOVhydR
K9Glbo1ZPGQyClXQD4g7fgMG9+MZCacblwPLsLr+9SQwN/vJH++vSIYqAftuCBf3
9wWar3W8BvV3qGQcQLj6c+Av24o8Y6iSygwkgPfn4n9v/ONS6oT1avEkOwaW+ubG
QRrmtvJgTxlfTVkPIla/PrgpjCaN1JWuqvbPxnzjm/9CpG0/W+TnQFLZ4BlTUr2Y
W4yZ/FS5P48DPGLnM7CrY7Ge2ixA83sOa+aHux7as9Ha81GKwg4OdB5ZltyMg2SZ
m6kDKYGzCKUQnx1inH5/daV96JfNbwbFQVvZV8Lol2E7dZ4X3uP6Ar0dDYNAs1SE
e9HMfBDvd/0xqUNHIzqkbavvdfhAVi95b+XUN0QefwFfLzDqXK8hw5uW5wkQqXQ1
9B2sGBJdyFFybQyHgBtKne4Y+ECxdU7DOlJEQTrSvSzR84vKQ0VJgsoInRGjpyiE
uWPr5163ytJHvHc8fPfKsKyvurIeuxOegbWwVkpHkPCe5HyyeMqoShJJlvzypXAH
CEPVaXTfusXDEtiT4I+CMqUhWMp5mOT7ZD/ggVVljq39wa9xjQkM2tFTBzH9Zv4p
F9qqRKb8HcmnQbYbSybT8LS5lQBELOwdEhQHMntD9Bno7GC7+2KU/FAltvpypQoD
cy+m3u8pVijK/bYRTQec5EkGEukMF2RZRtWvW79ODGuJZ1reO852drpnbANxtiZn
HfpB/HuExKavoASdeznSDZjiM1fL2B58enrWXa+aeUk7FVc7B8lSDk1lyJ5W1qOu
aLQOku2ERLPHrSzAuz5Txz/tVpSXT1x39vzE7oV8MKD4Gu5p5HB2HaTRF84DNYmT
bBdQrCHefk06iEk5Q3ezFGfDKTgVpiL90zGEiXsbaKp3iZfhDGilmyFIOaEuI09X
gWeZxodrahcG+f/5tW67vaLJFQSATZVigYnmYFpyyj330QeeC6Dc7YuMsDBRArUj
AtItkUNKmINnVYEu1CSxJwrlLVOlrEa4Xe26hciKAcMOrZ/I98PkAl0BXdZCus3H
/Ktx95TQeZAeK1+N21WZ3pDWTtj3kb2mUdSzMLezTKa1o55fU4J+Gwgpz3YfJUPQ
uXTRwsMkg95yslRvkjlogzxB8m54jDDHty5AmK40A0EVeSO41+29VEPXNgXHs+Kn
mKnlnLGSzPs2N2MwL1HlX8crHOhlm7onbaRtlyJT6lspjETXTvgwwVC9goKXvkqx
cXkmFHJmzI1OxfUDAehdXp94SMobkOsvJidgRJ5GrLV8Hl/55bkJ5ESYe5I+piWE
2lwe97bFFW4KyBS8x5i2kfiFlMAP5zHH0Lml+HaYxUIYlekOxgO4WiSNvwPPNGtY
ErNTzhzYpcu5Qu7WnbmMInEw+OoVaj6eEmXL12maO2npqbmVSjnFxuQ4xuhZH3BZ
sza5lvO1TGXn9kJ//qiRd1MfFe/PIGd9ij/Z/5hgLohxKMHwQgW8CErkWNemLvYR
IpIIpPjwVACqppsEKPsTHiwHa9IoFEIjd8BX8Nlnnb8MYvDiba3odlgdsvExZO79
PF1qyUpb3L0Rdght+0Qy+QD9zp3q15+T/wPrWtThjLtOS/BaN3XFkJa6n0sfmWVJ
BMeYvA23+Edppy216b8zvy3gaXMcqUz8yqhaVYnP8B4sidyPUhgBnYpTjf0fz1xG
4u+1O25dNyfUkGShnCNwojzvdMTcHZL1xKszGhRnGih/XxL6YWab5P0CguOjdLjO
o1Yn5KUroAF9blmT+dLsEhG/qdG5ai6uyV/RHFhLX7NyWtRtbERRqMbpuSo6tI2C
O9P7Y5KwHMMIeXhfPLxPYRwRrt7v2yEuO4+QAoJr+fapPByWgWjRjtLZ3nXVVI/+
8cKNZUS871ky1xhKEVSbT/wr2M63kV5pCTx7UU/o79CDIE7qkgyJOkpsahn7x7Iq
p0m8Y1N+2QHPzE1etUD7dkjzneaiorN5A3T1VXgeuG1NJDfu5vZuMz8xaPmIqdWI
GcuFVxwtJUK+RT8yfwiwR3dJg/sHNZhq5GZWfeR1CfDf/d7/bRzRiDIiP5mrNiow
ENjrpNBgiLpe3TpuXvoxMZhdN4gscm+q+j49omCxhE90i8CGhviA8IrFlPIdmrNE
48O+2F3FmNCEvBINOwCI4G7q3rL8BcHlsLKxYHpDVnPPZNfB6KFsQYt6cGG4YGOA
LO8OSc0rqaJrotcU5XEkaMlbbhCzeqXPymWJS5dFZAPUio0DcDO+2oSj+gJKaPTZ
cK4WM820WpjEyz9IW2aX2JdSWPQQBizw7f5MLjnSfcmrZl8e94aANo8H6FcOpdUD
VJOwGbbXxJTeCWNMkQDfRD5qkXhMm4eTJHi1bIWXLXDNfPYLnCHSccb+CnUPGG4y
pFbiSsruFyR8Vg2/Kwb6Y/YSlD7Q/9qGTb87N4N1Ilyfj+/arSPjqzLZNdltky+S
aG6VTTtjoaZ2+GENJRkMMrycoH6F2eTLWoxnjqmqWQWcJH9QHR5Qz+noEzXM1lkG
jIUvL+vwZdkL0nR8SCjr1oC0IvDQ/LO8bmEJGeBeqjdJhOg+Zpoo47lfugKHePx+
AbCrukewUbSBMM4N3O/e7BHGNZpx0glG59NYXztbJ5y1NoJ+NcNjszR2TVtMs8Td
cev+4VnUmctlCt97BhL1ZAYxXHSpOlNzkqbKQjOm5+fgJoc3c5w5O9/bVwQ9Lbpi
b0421WM2NdT5GzqbQQUOn0JXAqX8H1x1aPOcJRG1GvmR3OVhzJEiMb1rUFD6FNRC
UQVbXr0sVLTV3n4hqD7JODzTb95Voob6x5vrknd70r5bzxyZJ3HZ6RHmCvRv7bJK
GPiEfeNP023XK5+fX47phJxEI62tubqn+OLLSkHcxppDXG2G0uuCKf1ugLjA6xVB
Oz4Dg00hvz2zcjgRs+59XVSLxTAKSvjDgoYjeu1nwaXj3uEFqMIRqjO0Mn9WuDcq
t5+Bcy1ROkqo5XTjH0t4PEoDhPh+NSLOZz+UgE6jBN9hOcNZ7b5ZENFE+67oWwMI
eRnPw2zB8NMig1jY+WQrW/YW2ptuNUgOzzc4zJJBfi2yOyKU1iN1C8y4IdwYm9Xp
JUPB7VLrVIivDzg7DsJK+25D/+FrmnQgnbaMRf9+h6qbHOz+7hCbwnZTon/4pC8m
FCQ1qYR10EKHx64MWqWQgNy/JBKSRDAwxZU0UcRzln2fuMGWsfAi9hxTtN018kQL
r3JjObgT0XyqRJe1gYx74kw6D6KgoRemeQHHeg8Zdp2t5BbCTdM5vfu6KTT4WxGc
ac3gk8/8r01BOb3ZFmKGLaPixGYDnnkSzzw7cZqlNd0uKx/wWo9BeW+crVY2F1PS
8+tsIMB2QHitQoNTlkqwFa3C8Xo6SdO+fI0COpK0NUgA3ZedpC176S82j+/9N3KW
tuZWuFaaQkkUXO9MO2excYwbAHTGk2z4eNxPkUma/oNF6nwSHDBlZG6bpzX87CjF
AJa8/0E2rR6N7bsDAStmJTLy0sXE0jJrkOBrUS1uMuH25hyRxVNlrUnUK5607Rjm
jmcZmobbQQeXDTNzLtBPCxmiBfQDyJ+Ec4PA5GPCJahLfzmynIEti43cJjOJDfFS
PojL07UfXv3rBLZHG+dal7hMiu8hX/CBiJqR5BpUB155I/ZD5cOW9DuJE7ujqAWs
0jQuMsO6n9Xm3dx45fycFYh/sCjKNaJ+USbKGbP89ZayndErnt/VsaRtnaBlUAsw
Lxbm0e2MsF73OTfm8SFqym3+GFh1Qs15rwfRL+0kk4ohQCacnKDbKrLjE5737wm4
EiyCiNEd7cu5gccVDRC8y6Lj6XI2HHUbrJfPOZ7gcuOAUit7GY4YwIvuCRU0iij1
XxUCPqquurzh8yOMOzcnGJYbA2HU+QZQGa1l6L5Sy1b1qDHVpAGmuU0nin06lqbs
IS1AHSxsX7QNMIPUkncDMP5seGEki9OWKkBZfeucpITKWZTa6UL4Miaalx0Q8/Xx
rbzXFPn5kHGzF4rWdQDRCJH09sWLO+MVo9B+uSPxhTdseJxAVIxmc+qNQj3mH2Bo
QsECVYMoU+bc1WFswMV9bvrqDXyZGTpJHP3fO9XGnpBLMdvoYx8yIxuqP+BLWVfn
3t2Q2e9Cx7GrtQr+ttNJcUxGWsY9haP4fR/b+1P89tiDekDBTBr1+xfSLa90lKu0
tX2X/5aIxcBfkh5/EZ94c7+qDljALmR3r0eENP4GYmO8V1u5jN4zz0z+xt6B2xJw
nGkBQ9l4JrFUf/+zZHCxaut/cLZAgum3P/jjhFW4lZ8xsSDmhHYG55pKk34NrqCK
sYPZFx9BmPDd+d+4Nb0B64yeL9nWjHTP6omeb+RD+FkqXrbmXB4WGI1RGZogMBjL
TLTHSebYv5Zkq1RWYw5KWHBANT9FuKEVTsLY4fgtqvj1r4dahj7BU8Y2KLZNx/GM
8nmZWA3igsorW6cXytoTn5FTG0TMWunyJlEwSBcxYnZ2H5xKiNeRX1arbgZzZ//L
6BKKTlLDKfigpsCSuTB3jiWws+SQXk/QyMO4VfcB+cMMtBiAsnXkGTESk6MCo6s/
ymIhV6D3/zwIW7fzju3VMgVCWTymxNSK1F3RUireSvWegRsi/y8knxS/ETXsaTrk
6k/bLsnKqYbqY5RCTEeJ1PVTjtZC/t0mo3au3FXjkQLUYsACDR2z/pec9ciyfFkS
LkrQQERtVB/WKu/95Eq+IMbjnagzCsYvaPAX2yt508aiMpGsPZcNg2qOlVlRtXhy
h4EXJzs9l33L0r/Q2dK1+MREp4XenZt+l+rulWDDKbmDH1PFIsgQl+LAzYSTCzHO
XdmhOC1+kFX6t0bGUd6+uwCXfcqXEexJD5N4reHB4Fcs+vSmpx4gDp1xLvZdCfSJ
C/o5o72Y4fSpQvW5zDpGXCalUaLcEZHjPZA5RZ7U6bD/QvkmyNSv7vscZK2W25QH
pBf6bgMpuLMA3zcXxeumKmaJOWO5dh1gXRUiXiGwqxgrANTKyurVgXjOuYpA3/b7
JuTGor37CMive+J6D3NHpPC+HTDri9WxKt48MIytT4VhjrqxJw8IVu88vVG5y6U5
6fMnzrCbosKaIzHnSPMTvMyxeTGTIeNL0sIBgw4VOT1FKC1KYOOtWqWYopk+ol5B
2UHbJ1ZlPkF1lYYfPRk3E+m+16rd9Ek6J8SUO8dB5Ys7wuukewihlIbb4ATb7twP
E3eHf8c+nqWTWEVPTyF6W9QjCnXvDxaU/z8eNAg2uUc0RXZKCVIaQm0jATSeRhYi
8YXExGReR42pDhBCktyJAmFSmALeio3DuzJGrIprek6KvBbLv0NRnQZ2HFIm726h
oOKU9zUCSlO9/yG+q+p39AZ+ZIzN0XoNl5XAnBJY8qHNGkiRx84yVWE86NhxoFR4
vwm5Fnk1UBdUOz0MSzqk3wETgV02/xN04ACW+wsRjJaQRiDYBliVPwWpJ2T8/ynb
WtU831anCLvLjyr6x91e8xfUtdsADaUIOrygVqlw8dMlYWf096lM5fee6oKw6dDC
01wv8zFMeUgIOF/1suJZXpNuzlvmDR9pqo01FVXXDmg6/6EDJ8RwYxlTheN6JEOc
GtcmL3ewTplpa1C3elZl2vihRS/LlGNRSTs+PzptDmtmUOuAABDLmqqC0iSVTMt4
8goA/GTGVMn5CjBATVyda65dNL4fo6FagW2AMYGpJ+rsbowiNPDD5A+DMo9I7Rwk
eLhFTyTwqQk+J0QGJzJaNmqbbmnnBRjNQITa4EfyCMA3gzY4gVNh1D+P+GcCZaJh
f3hdTk4k+yUEpxC832GlwJsyJjxqyqo5LjE4CMUDxZyxbvqznSK+rBCNa+AsMzUL
62Oqmeu7IRhzSqV5qpIDbbZofZj7/U5FKRuBNVfUlXyVkINiz8k80gZVAL4G/ha/
R6xonGmQ2GLQCZH5/sPXt7GGH4XBrhQQEEhQ0ksmq/O1fv4VypPzbsG3QTMTrFDa
2QVUMvE8jt6nYyCnG3W0NZMCB8bJMgr0q87l0ydPZRS1MTTVVDuo9qnJ0JcdfHUu
HBf1PZ56KKQkdaoQQF1tEqVN9+pN/3phfBykgBlFK112NNHR6tJIFHl+UQszyq/L
UjeDeJOAcDQA97DHK8jF8vqWuc4YGQnBa/LbgG4PzLbgVO3W60x8p4CJrVMbgBr6
G2QhZC6oIEPKRzlbu57cd2A8VhNFRK+Lr1PZ139W2wd7B/TOaVd4w3EhSN/tdlYj
LM7PRAlamvxwlsaikZ2ccKrfyYY1PsDMEJMXxaHDnZ76dBSsMr861VOQWQa7WGVg
Pzs1z4wh9h8RzFiknqiceyVzOLcDmw9tL6cGIXybLNdhTWWaE5No+JmrgA45RR4U
z9XWN9LjWEC7SpOVX4ztYZktpd6ZjcJTzS+3YtsebA4BGfGRtFr/lvETsDeA9uLp
2m3r2nmi8NnInqpdYAJPdwTX/UKG7J95VSZK86hBx1BIfy67gqk0LdbWQXtR9kkw
8TC9YEcRVLD/TyJqTkTa/O39yBVpl/j+0qiDzEyKF401N6FZwG26+NeJdUhWs/7V
Qec7TRikLkcxPPYq94W8ExPwUOu4PaXIo2AYqWsjLlm0r9ecWeMVc1jdTOrM59JU
KRrIMUGtsC8nYXE7N7O9Ei9Bk5okefu8kwdJrFij273kIrrwnldr0xN9WvYq3Phd
IzWMeg1mpPnEVpt8NlAnkMk03iY/uvaNBoaXMNlhVhEdHdNodo5STjcCgmlGQpBk
EIcr8TYHdYGXTfpheVYx0okoSbKPBPrl9QDQRIwuQLApR8A1V5u/yPLrxX3AGQ8K
uToMZWPzoAftkH2357atqOHMyNV7ey4m695aH9VB3YEOu10UQkyBG2AkBiADn52v
15f9IFcgBuICXBq4aLCLRD8WqgMwNOsaBFIDmg/JqIdJga2/l/2Bkk/tlsvuN9gq
laLVinsqnyOYA+mrD3MhsB+cj+//EdZJnins/VG+4Zs1gpWxXS1+tAyAm6HaiVkj
3ZLpKcSC1W+s+XnQ7pXOpWW0+Q1KjZodZHRSGbpE2kHaUZqmBjCXhS7BsV6F/EGX
ueduWU0xKAXp0KvfRg44TZfm1V4MfZVm7ke6ZLRA5XC7HqIxaVP4QLYn8GREMHCX
b5nUnAr8e3dzsbo+e0J05NbUfNLpD28v6GNukeM3L+75Tp88Xs9EeJ/WKbR2mCvk
hFiI+/67AFFC+pFwOrouyJCyYq0kU1CETFrWxOyMZmPJ2SK+E3pFvlTPuAKwQgRe
U0qQ5CHpvv5qOOn372RNW56sUoRsHOJ/xyygzZyfXbES2TTveAl0ADvJsjO8zt3+
QwP5xlaDi74GsW4dD2p18BOeyZP4D2heUZO99IopNb4hmU+V2uMpyxalvWx4F1xS
NcxxxwqLgzieb0oQINN28fHefO5xnM9KaTKEyp1GOQPo7I0dnS4AuBHT907zYM3w
iWj9ifuA08m6av0b7es8h/0aCo1o5/q109uLjckpYrFe6Ljt8Q93sitwW6pBOz04
JseMA2dUvevdJWZG9qWUHzWQ9kaWscrOVTTWCvYnwoLLupe9xRlxCwZsGuQu509/
JBpVDjQxXAgz4JHap2HV8dxVALdx1pV2VPiPnQKV95T1UXo0e0WKz5rketwPj2sm
wsJOC5ISw0kMAKavR1t0PS/Kn9K48WBQiObnGshPrBDADvmnAQmD0NVnaRFTGC9N
5QxnwHoWoX0EgktSBRANrexVnqyAcjIb9fAGzv/zcO7V/f5SxEIp1Aa7IBoyyJ1F
0wn0Nbr/8NE30rEwk6jPhEsrZLz7Y+FIe3Y3UYZHbN2+SP3iWTyvroq3ugon9/i3
d758O7KMFPlDV8YfW1kbuNT8iIsJIjtcI6hhJOVAakzqgMAwb6KxC0AR5FchyMEY
0m4sVDog3BaTnqeKvWQYkpv6o4prJvsDnkkNZ2L81aE7L9ltvmUN6WerF1HefgKE
LPtX4eDlXGvEpjvKvEcHFhfOeARpFa4ijShiIVM9WOwASYHndcPH8g4ubRmZIUTH
PY714a2exQJxNkTY+SCpy313yshTY/PZ/eIRJFI1pgJwBuXf7ILIGwpWOnK9b3pv
yupES0RaGbuAGwky+zuUWCdObw5X8PlSfE2Sjhb1HJ7AywL3Ph72FxadvrSOU0ID
DSN4wTsz68TDaecVqrmG8/7pN+0idemZBFw1+qu6laGqWw+QVv5q/vgzxcoKI/d1
NlBjV+aw8l9HfF/kizSXKqMRP4mL8FD+iXdHnfg4e2Z8NPPRrVOMF705p+/RGV/V
380+zsqk3eSEGM7tKSRU7w9cSzJRwqIKVbeFw/vAT5fSi5NI9K1qioHh38I90seK
T2+7a2syI83urZpzZbuzXCJQHlWEzqRNsf20qoAX3fXyjOCHIdTl7hUUkAOs7KzK
QG1fN53/14JKkv0DFTFHDYyeXIXAzCPC0IFVRDMdAAFglE9+2PMHHzsgQxb/Ecsz
zoBlCbK/aTkKX12xfPDs+HYPeN80jUJVGfdtvbzqjagb9aVB8Y7IXs/cyIcDrd7a
EtWsuszFZvmbwOQmrVx1a5F76SDB0BmNRQtjqT1X4wz6WiX62Szh3Rv393Riag1K
rV1mPddwHefgrhY2+4wJtuTb/BjdCTELUwVG9+r+HPlDPDdq0I+6qVx3GAt6r7es
X/HEAzYH+3hJB6PvgiDgZEynZ5mLMiX083A3eniDagVTHKQ9z4s0g7qhyC9cJjDf
GIz8SUhzhFjaCDLnShvNPlZ5ob/WRhxd7ck9QrUelgqQYD//s/oJRoS/hIe0ZKEf
cgqb+TLVnf12PggGFfaz0PyKcYlW9FyNCMxP5pm7vtt39NgCJlxdNV5CyR6ANvk0
6hclW0cs7c9x3hkeM9aFjJulUsLvQMv4U9gvDwE4BJNO9xvFza1XcOaOBS6inD/C
AnOW+EEEua9dCIWN/FSe1i/PtIl8Ae8KAA4adKMeqeoN1Ia5S5qEI8i3g6Q+wvHp
uoUy1XV++3MhEVlaLPJ8PlYrGWP8LASQkUSrat7h2EOV7GoNu+r2f0Moh/0CdNzq
G627s7Ux3xBqrJJD+hFO2dNiZdFF3UKWONBBLkLc+ddvaZqiqP7ysvXOZAnTS+FV
7C3NZLI4Ds+NLGhJdnLi2IGQJjRsRPncLzInuew4fp/v9Oz+iucG2jpndcLrwP8y
D3vQ6791vikEcTgWYFvQUCNBkuu4Ngd33Wo70ZJAbR1627oL0T1gTgws0X4J46jN
gpdpIjvaMjc4iFxClFVwRjrDXzRyb5XRwCtaSaw1bBiV6a0sowrcnOu1QeYEnpF2
ZxxVCrFP4ji5FafHPVcADSp5E3o8KMClpVKquvab84d69D4IPw3Cmc+YsBEE8vJ8
r+KMaVVJj3mV0zeMetwNf5CxOkmoCcY8BIavKpOzS85iEppht9IcBZfxQjyDXuGV
1JIuAsCsutuXyUSrMm9+79wjtXSsO8MYzgg3EPFQxqlftTtL2VXj7L+mOrQQ3Vnf
KPYzo/wsr3SY5QB5FUc+aNgOqYGsNJjNym6P5V2qyGLJ0TMAnr/k1My1uBva3vc5
QnY0IYQLkCGGPBVpYB7vK+CcLZZtBG5FF9EKB84fAOC3mW67qggHAat2UngY+U1P
CB4EN5tK7rZ8pXHUzJWEhFHomZtoB09uBhDyPOff2tlw/mg9FTDQszlVcFnCNGcK
MoQUqdeFvHUZkRNFL2HaoZZf6ldyUywDRS4/GXdySu+uPYsKqIJEkPuNWYTepYH3
BIQ/02cBVszFyMM0VpSjwLwJCR9BpwyyDN/n4oZqNEZRzCCGSXAml/cCEuqGXGUJ
ybBLN7XFj4yIfy8wwisa9SL8RF59yhC9n8JbPux7pCOD331c2HR9/DfhLGH3Q7QV
+MG10h0NixJPXRUTLK6QtAt0zWDCYehCjnaDGCAyhaIrb4Rd3FT6L3aCRyRiL43U
O5v2eKARA7/ozkG6fTfNPNUz3B2r6buAh+q3pGm1kUEFW6pe2TzVgRCWWrcp5giS
y4ov5mmztK0Ti5UMwr5hUOtgx2tQsXFvkxdCXyO1owTO5qLv5wb62jZBGApYQdtM
+9Y2PjjIC1YI2kmodJ/ooPMGFrGdud7eGJVMpjXcI/eaTJ3rfkuccJaNxDHNypER
lvVVnAagAkEWPUENjPEMFTqcvaI/Wiqs29hzslyQ/rDTczmUaqn7TkrAFjZvYqL2
H6XR/UAS89yccJfRj8IrTvn8maIT88KoVyZlBIEFvg0+Si7/pkDGuCwJAZL2q6Dl
rODnA2Td9xG13qZqgGHv27edZ+lR3Cd0juq9jA/8aEtfvOx0UE3ECb4vUwE4FQzo
DE7TqX4FprhbdonRx3RmiCVWmhFzIXhlGY7a9zkTNMD9jk20mnEuLAnveEGVEj5+
BaK+gunUZqY7IuWpJzplYoggpdWgV/cW/0+/SbjoIznh+SGi32WNz5a9rpDFJXl7
NTmZzR86VCuwxUOMfvaT8cMlnspvq5qc6kTEUGpVcgsFaRUJG1xBvswPJeg7L+qE
FzNIyMxzIcPNmPBTjs52oxcAJyJ183viNIKSkXOiVlnnBIu56WsNp2oOq8kQJBut
QF6vP8pKGXMIAT94kkN4L9s5rpUtjw8F0u0ekUZHL7Gy7WARICKQIZBnVxg7iqPU
8rIahYkWO4k2YpwlVMkFQeO6QMLRDRfUiwi+fLnNAvNhsIJaxB2IIaxvZyMpaHIY
baLlywerHu9bGckE3PMv1QP5G3gpx+GZoPdST1LZcuV/CxI3cDlkBGkkcVssDqcP
zJ1tbPzOh8S05k8fWMJHpBhA59qnqvJetluFYiY4mlPiYidcm5HbCo4V67rZljET
Rk12Z1IgRHO3KYO/WOeye7t1+Ju0Eee3UDIFwCt6HGyF7aViB1il9SVew844x/sF
sLDKVu9VD50NCsoFDpjswKbyAyMDrJ4RHt658Fzdt4q++aXk+YHfSjXh93YpzkSW
kwwherNBF0EdB58vowgG9MvMRFsbVFrj8fG9a4Hw6Tqanvrkz1dWWKdS/WKUbdSP
AbauV2ENVqXKNjYUCGNyW0JVftM1ViHxrtiOFHZYsuP2hOl5NjhZC8Lqi9aTfXQ/
21+kBHI5o/wiphxF4pQLxOq0mLFzH8rTpzMcwsSmaPmIAZfNql9NgjXUh0JcDVKm
quCdw5K2EsdMDVTO+YzNatIO0qKLFm19AWEbPA9uiCnh/P8oRrwy8+wv5YtSSnKc
rvyhNTm/5+u9S0TT1Clw/ofEnjHyMyVRHpGAtHL3zWusBKUHNpstT0J5kKgUC84T
M21T1s3hugyc+VkhneQzp/u4pr0elvij0392MaFID1KZbqkhBT2ury6w3B9mzSJ9
AFImSFCvMX0nmPYL7B8InqC2mx59NrFTPlpFvH8HhmGQ8PNL3mCd78cPeyFVHT0F
UcKARH+n36iLt/1jR08d7TE/xHAgE4gZOcZcqzVwDkqlka/qP6qg+nMcgS5o1rqH
jc8VmJDlpTYtp6/H29sJOycZGYjppPBUK3F8TiNVVIfDwsC2epoxGoeGVyL2pbW8
Ju9UrKtGh47NQ3EiJG/IfhWo99vABfzpfQDKCMmnCkYqwYDQRxg3tXPol0WB8fyT
9i5VqeK0trXbatTCfrTmXmCGl3S38i/0Uen4NqJ0kVBeZoO4rzOevv2v3/w+BLkx
2SJ3AwQjbThGPUPOD+DRnz0MVVNQd0JIoyxRthb6+xozEi3LfiPmdgGaiaqB8j/c
K56fnkbYDdbQoOCl6phLsLx3QZDYS3Xx/SMaEUPP1iNexegG1WAAMMheHqZhheQk
fidyHqXg4HCB9VbyxW3cHgDRPB8RoL3Tg9VaXtkaMFnnttEvBPsCxW+KYlDn1Jif
JfBLgJ41QjOP3EKB25zEGbgKQyIX3W8NShm7Cbe4g4I9CZBvLJxTm+LSzZj+4tOw
DR1eDCuSn/dgF3WvcIuU08h5hCuV0u/+uT10xFhxNwf9Lo7rkRT69Hf7vN0CW9Fo
zYbHx6jH1M4EqrkQOcPN7iPHzrV1Rx5oMTFnc4qdMALZqo1GVxcCwePCF2UByJKJ
RZ8u1KthCLIW2Up5QLPzXvb7uE6jVh8VjIY1N5NCWOp6BwbTWls/BwW8OJNPfbsq
OEyU3Dn29FBUTO+TtWg8l3muH3/FuixIgK6KFT/Kkg+uW+v3kkppc5Ce2byEdWnT
tfGkktU2IksdCNlaxZW4jEYZ2rcxjZsYUyYb+faAW21nmj6ClTT9LX3+kQdNz6hu
/8nzWy4bf7ZOrr8nrWnT241TAWeed/KpkLhFpW0jPrrsj2m5TiUOB52c6pHF3Kr+
beadXXq+6i566j2B96sneSwFoktad0MkD6w2hYZU2uJbbsrVK9niQM9udoycPSpE
KyJJD3LfjODT81NFjyD4F3H8wL2SZyea6NsO/9Gh4r2LOTWMnXA9P8Y+ofdbLSw1
+Ts6ORNI017cRqXzVC/fkBxAgGYgWZPNRzZhRcYuc+ez54AxLAKO4j7WqR8MmnFm
DxPDJfjkXaLX0KRpz74V8o1qKqtokSjJvHQPRi416PEKHphdrGoGSC7D2tBPS9/v
Dmm//XEu7K9JQkRkDE3HxyAhdTujtW38C1xlZEcDbw0BBMUAVpQHRXnTh3BRQjY3
jNPq3CVbx84QqcXI9iVuOG2eUxxwKEXKoaKfCbcdMYaElBDUaIBZeI3iydZZqKhs
FzVPz9FuT4XlIMZrURrH4bE+oljCicDTVrpMn5jJPKxBK62k1szPbo4XcbK1v7w4
gFGVSrivU0v+v/gfIBYJdRMoxuOzAlQuwsrFCUmySvXd1hBRnKckJw1hOYWlUZc/
8GYC2T8ZscYqdR1SYiMttgpdMA8M2Shp//XDtEEF5koYfuvO7W7DqNCkWgKrOY4W
4fmMXt7R9/MdyelY6UNuYvISIaY0Ccz/2L+9c/oK0TjzcU8fRl7jjx72T+MGU8Gp
6uj5xWRNBVy1e1vMXFw0a6IkM7IXOmJvR0yI1VcGLjCroPp19OpN3FiYoR5kpLJG
JON2Utd8EEWPr+cKMwlrCiBved/xNQou+smMbtXkMvLHH0xA9Xn+PCJBMBk43H0+
acYVm5DNhtVWzsez8oT3vVFID/BK2mWzMe8p/Kcls/JZxnoiyKHDj3gO8ucrRwCG
lYKGUePJdrqvTk8qSUDbodfr/Knftl+ghVMfE2uIF/i6uRdQZwSZNqp4wFvvk057
keE3L4jEPPZu2vusPhFkYQ20nTE++0ipSZtL6P7ia1kT/abAxcu58VOpevZsV/Jn
26/rJVp54pIM3bHoQgM/rXaODSEzyzYp+4fy3iAqbSmmxNa9PuRLuAyAPoVt6Z3I
BOYAbmcfWmDLQqmbXRZBuXY1tLWKnQgyWTrcDDfneUqIcRrSLCUs6hWqqPnXmQBl
L4DY3Lnvc/d8U3+EyESvAVIwNwS/t+oBK9pFRb6F5H+DXljS3XyfGUpuGGEJ7gSl
IxrGTNvRz8XGjigMmg0FV1/1UUnw7FxutInl9pNHhpq60YCAEB1QO4crnT0JqXXw
PdErk+2E0aYJSb7t+xJaHkug6SXIFNIykr8Q2/EUfy5MX57dFOf7b9zY5Dkn5Rrt
VMgI7Ud1HYhqcZxwC1vX1QjAg9tIHXOFQWCngXT4TUTlddaujf/EdY8jGvx8KNAo
+qkfjhjh5LJELZ09DHFqBsWMOp3zUQlamhdZm2ucV2O2xhq1Xg7hYMkpy5EnLixE
TQtroFIH4+5+Hg+qehIvY4S6+GuMh8p3+h/ECFzsQAYbgBoUw5p6SofbIlGdrZqL
hUph6X7/hqt2uKAnF9FfUlZ4JM8IS+CUDmGd1zkHdapKgwhe4w96iljTMkzWB744
kiOjdGbEpHJTG6PTnjMsfGjs2O2FEfQhp51ZOuqrxdSONxU9ROAvfIVh4mzLIe2Y
nsq8bKSTvZAQnOxXaakSf89W6wc9jfFveUfBZSdditwgeg8e1gRvFGDq8JVJDGsn
EF7JwW+H1OUKJsWD6p0Ja/C07sFKZtI+AmhuqaDwJ/NwUGFTHyQBltUmSVrS5rqW
ow0zAcjjij8hnBfl9A4Xt2vFX0lmLdMlSVjN4aUFYpXlVtxTFUu7jWMWpL2bvip1
ZA5fyw7jK2fEnkLegRUTfWqnkFwcJvEsWzldnmdL6JXqzdyCNzT7Re3IUq5XWxo6
pPMLJE+UyHxQBwpyRmGDbJt9DVWkDmF/dP9M5XO50nhi++tvQO8ApXdSfXWint0M
kKLY5rzTLUoKmLte7PWpz9C25ORarofc4/W8c5x9pQIf4+gjIsoM8bUF/52WOOL2
t2U8pj2Bsd9fDCIHIA+1osu4Lo8a25rSWIsWxTK/35HTe0WKD4aDffpyqwWfV7s8
oKzrmgbXwrVkJI/Ir9SrM3WtsxKJt/GmdWRGAAzaaq/8F8VsHxBvjj6kmI4Ei47c
6IDQCn8uPsKkoZ9ifQWTFLG/DBqF01175Ko/6Hw5J38baCiRNk2ZUJLE9hBOZI1U
BT5jLf5aJtAtrj9C/nQ5RFGnf2LVuda18wpP/hYFpx5NzkQR8mMj5ztiGQikdlJ/
o4YB3C9J+7MesP7wD+IciyOW7sv1u/4cWCPb57k1MuLiN3bVStZUawxSAYshDDqa
CzQ+Twl05D1nPAA8iqsQRps+AkQIBjLvKGLsZaGWvzhV4Uroaj51yOAuJzsj4X33
Z3w0o/qs00OltnGobA9anGaQsNWd6+h/zmlm2+O9NfRMdwQv17M22+EHoqYnvOXg
Gjh48iqXHW/PDWVH0GYFbx1Y/OkMUY3vq4BfR73SkD0zeuGrAwdqUbWan/2KuEs2
+pZapLbHI8JxBaBK6QRJ6QXRDWI9074xMAL1r5iqEXSdOPKuMstIAMmaaaCnuM+w
kLv2dPtW7qE+/zFo4eYdAQ+8PmxUogG7SmM3F5O3Z0nJpgFwiw45sAOZS+W9c1mB
eSG+HDG29R4MGs84aT/bepNU80XVQIs0KBONnraXcCvtBN9l/Ed7j42GR0nWPz8p
hTJD762/aeeIVLuTPRzW9qsnTpruxKwQ+wnD+cXqPr6dSZp+L5V3CyUHgt5SaRR/
HYVPhZkwBLqi2Td3vxKea5rbyCITBWxLh+fxAJVdAciCKePiIFRHYGwU54LbbOe1
CHVLUhyZBOisnktm0WRcL7G4+6Pn5iQ/tW+W/HSVXDM9vpQQHASX5nppui690J68
r+uTyzHrbgRtPar/8bjVvOyeMbjy5ZS3fGm85dg+g4RFXzisIkgqo+Wf5TUFQwm6
6+VKZHNYe00+j2shMN6k5ue+6dDF1yrxaBjz0XsjKBVzAOwHLM0qVnu6LdfeZPIF
GfJmdfX3wtcjUcIaIc9+3wvdzoT7bIgwiNANBYJ13jGhAEBE3EuORs2TtfJjez/e
byNQn6FkxJ6clEqPR9FXV6tVWcggD5OHg/s1Zi1VX0I1LHAbod65SaF1kJ3ppcRx
dq911OP5rbuecU7nIF+v7nYMqTAou7yA+7FxY4I0ZRfzuH0eJkD/iqMnu7nnPBF3
v+TJkwH2s0fYUPlixigYmvdS3PQdQdc7Swf1xeo3iehmZ8in419JyVzoREOS1oq5
H3VEFteDS4sZwEZey5zmxCPzI3IF3X++ihrCJc+J1KwtSQXyY4YeBTF/yRWwBXOC
kVLeS76Dch0mwoT/VbpGo25fBAL8Fpo2q4zICwmdY8uZ4dmn7zsYx+R74Q/YvlqP
MmsBWuG0/Fbel7WLPFM/LoNbkRo6UyYlyJsC+RQ2pjexMScGHAqSeK5/tRv1YxC4
IDkKst7j26fzGdHDF39EZoJvW8y4NApXhkAkU9RHVEbnTPmwwTN8Dd2/GNjvMbVk
/saBi8dxLZM3CwWU0HzVRF0zM5wMN54zptKmI0+TXIZ7t07buCj0WdTgeSyS7yF4
BOSGSEIW4Th4PcNKmIZgnfp7ifo0BVkFE/tccnbZvJO8Fk1ygEjCt08o6rqa/Hp6
P+dbxoznP/qjqnw+Zaho/SQGs1QjDogWL3xHVZCL+Wbme3NdTqLJA4xw3SX6f/Db
eZN1kuoYLry2oeakbwhwVB+6qh3JeZlXSLHbnsNcQE0WYlSgD/LSNAHIxzpK0Tkn
yhyFWBDwsaYH/h2ZQcJLVhuhLLw17N6CjmNuw6mH5SiwocIU1YjedXE1sOgh/VlQ
48XNA7I+GkAvUqYuUTZMDtr9mfURmgxe4tVjApjqwOggKm3ydg5q7h3L1gU0yVp8
udZld0qsvZoilmAbo7EKnPlYIbhrTWVYAo8tUAo62Yeq+TXn5a84HWsiPtk7rzoy
+0lMem931E5Tr8yWhmme7ugN2xJXQFIuI6NgM1ysP+f9GYYb5UUW2JCBRMvx6XMo
ehBDFn1YE4Xk52ABV5rws8TS2KsRfvSs8yU4u1LgODAtjCGqExlmX4wBYM+lElYc
QWdcJji4mbc1/veVdlMBXdg4vgbkknXqs10S5XGmxJVnZeLfLBCq8CLksHisiuU/
V674P63bzFRnEUPO0EBW77zFvONBRuAWQy8nKx1asAHQ1X+97J5aFSYqyM77IzhQ
5jc0EA0eqdaYARvukntDrYsjmeI4YIF8GKsoChFiyrgZnCMi9tix0By7TOhlFKMj
VHbf4gyWtC6v6/f02qEStPPYjoIaZy+uPA0gM62FzXN3nDuZp8oTWzvN/B7ed0kc
2AkttQ7r6j/TN6BGV+S+qmrCfPiC9/vWzMKW6DgrkfcK3avGJMihIh6NfzkBKiiL
t6bSC1wPIiebE7KbZ2155E1kQHI9cs+78GOz57CpZOh4tcpDYIytofrNFnMBzsJA
noUR0FpU3rJGYfqP0jrIFjk2Dizy65DOXJhShGMatctv/0aKn+HIIl/tZYTRgrOd
Y4/Q3BbKVjZG5akDL2rwgkoOVXPgNwPYWxkTnXqRe4qmxyKFv4Xg7S/b/ZYSycnG
mcRK8R1BcX0nTmtuSLDjXKvjW+/pYxYPj5UXfIYZFa45is4rrxr6eUkj6Fn3wz8U
XSj8c33lT3WHwMo+zxk1PgA6LSWvjJb2Xs/C1kntSAZQhF3d/Kguuf9Tt22OyE+q
K53qc396r4evNEsvWHNv5d2sDFvbOELmHQTTze0jeewLAThA/4A62NnLZueR2gif
26o8iQb7ToWT35668ZcVzNEj1TPsVPqQEhcgd5W6ZTad7TeEptABbZyIbRyMKIPG
4bBJiy91YZ0bsOaqcoYykzKrVjexPM9+RQUe2Nxmv4beYmzsGWPaMKoIVHo73zy6
6TX1juzMbuyzOevvbg0Ak2nqLVoDsPc2sk9ss0S4qEay9pLPSHBLzNMN9sUd5/JE
mt2nwwdmH59ptVslwOnwMCkIl/kyoKef1TTYdBTuBdUh18v5c/b+VJfL4eWM6Db4
s1VGHq/iaix+BUBEv+FwKnRsImtJ28/xlAAuF4mZEAeA3PxADWAxzb4VMTFYXeDM
zcadccwCf3CGJddVDJpxgT9hHU9AnXj7rvcNyfxebv3gtV+ibQAOqaRR1jEO878Y
t3ZBvE49lGmemfjQjdrwTHrViRUVtVE1xeZgqUuoXniwrsV66G3mZ9DYUb6+ZX9n
H958XOmGdA2cVuprV/A5gtkBSc/7uz0/veOysQhkqi5lHM06VHl3aIyacZX4KnC9
vZvcwIlZ2byXnuBDE9cnmOcg7f9/b22aw5sb2x9VIYWxz3U3TvPgrL6iE1MfouUR
t7TxDje93F7A6WVKwbhRTPoxv5/yQ6TckGxZCMDf/1XJz/2r+IBMYjkdqb6SmItH
NNL/xFslnYvMxg15RrrW0QF9ihjj8dEFRI7CKEkuDpnKqa9Gvufc2u16FtbZz9Ca
sfOBKaHDUINUjdcXC0yyRLdOjEcVfOqNr+XEd0oolmUziuYn/TNWZYHiUXTxmHk3
dwok4lrE0Q79c5+9dfPrCIa+t7s5J0vyZ6CsyhIfpL5uZ0UaKwTKB6h4cL47LlmK
7gomEWhM70UGwN3BTlYApy/5coLhVz5jrZI9FdNswIMd0yXPajDi8JOirH+Il0vd
UO8b0rX3WgbBWyvx3xrrKlWuN/bE9oimFt60vPrgYJpu3Hh37SF5IYDi8ESUu1xl
w7fFEj/cROi5VCSq5tQo0ElylvM5naIURLFfG68IBlk8WIsEriPvlrlUxWRF4Jmm
e+kRmpY7/yqT5VIfHDk591So00s9GXe4m563RSZVUH1r2sFuHIa62nyp8cXTmL9T
x2npfkOCG5kLN9ZetHKDw8Oq5IVayI+TrofkRpFUSgga+jIEBhpg/7R1AYuCUHm8
uWA8ru76DanqF5n0Dv3+8VsXSv4FROemGrGuAHlNf/JhrJU7EiYPT1o1EsXOu7ek
H471wMfBdZOvIreQbthvXWN+mZLCor4GubobZOWRl9sQGclQMGI7Eq0vcj4mSyHh
/jev8aCmCjCc8R+gqYgSGFA+5/c4KKOzXDV85T9dkCbbL6AsEw1Kp09TnDaS867W
kxM+mj48vfralLPcVXMs6sPd5B1nU/BRjY06souJuYR68gIUvd2sp10Uhz4GCXAx
0/xIALgDpvf8vUSuomwLp1RyptGAcav5SPPqKk55wm2RbRh1FhtBBFqG6wXD9A+r
GUiwcOlyZcv0vknNs3yDV4i0zN9LNY7zFJn2um8nhfXknr2pr+jfBy92bKMAEcHw
fvlhNy2v1zuoXIVnzV923456+N2cBdlpG892AkU5kh3XvX9zpiHqaABJUORBI538
6LG8x1r8UJn6fwKjbhzndwrNgjkOSlJBNHhwKGgWDizGsfOO5FKTWBryGCfhlF1M
w7EO8fGp+8QzTpr8/wHpeveem2ook29schOrxgPD2EN78d/sF92PEygFoUyW5a7/
sv6au2CP6ytUmn/yHFEuiWuIT8GomFJd5HflSX3Hh0JTxLQFAaUqnnALlfODMwKx
AwYhxvsVb+qkOeU81I+9cYqFkCmtobiAnhTs70SnIN9mhG6vIev2CjzLrXDULxaq
JhaUWzt2gvnflB/xwVMNEgPHHh9x9W1LIykGntyC5qHvHq7Xh+jXYE8zCHown9Bi
lhhm5uBMaEsyQpu5+UsDAiYmLGPurJwwN9rzlYzcZqj3xmbOzhGSzeyhpKlcCdwr
ObR+OScwtUWwtVTO6ZF2P4foP5OXpGbEk/I+bQv9PLqrpg6HiCBOvfMckjuR03vV
y/xaPsVYEF+Wi25gMcxSVdvTjyiMwFKXeEJYw3RcaL5RQor33pzAr956doYS1dqo
aoWrfjTsUwIru9O4J0QtjRqQVU6MrD7I5HRKcvz7Yi48R/SQzGMxwEbjh2Sqd5xh
Mj+mkOwFiHeJthf/Ux6MuSHiXXGWWs+ifu4iT98is4MO0/9JVItpok8F1ySK9xlr
jFgTBK0T22VXgbICUn5jS2UFLfTkVDEOWDbQo5DcRtCGdjgJAgaR9ZWNdWJyzT5b
a4vXowWTFNvoiPNNEaAizmsJ+tIE+kucHsOKfMVsI+vQRxZ9JoBm2g3gDmtJCbjH
p7DbVY/3CxeVs2ZBA2ot1rkjrcyw++BDhYO24Zt8svlNQXT/xYSYttKZBFsvB231
6kg2W4/arraQ4u3R4O5LeTiLTKjZbQ+Qy2LHPj50heJd/oWEWa+vQRazgwm3YaEC
ZmtJg5iNg2GVi5LUp2Z53Z7ksKcubk+uN+nj24ZuMV8/cEaSO1uLPrMnlt85FmNg
KKQvAiz6DIvGauAUTZelB6mPE4Ir1kkGv0KwNsRp4SECP1eZGkNKss75oGFTFalZ
JYfXXz0Efu0/LZ2t5QJmu/MSFFxddM5ZImWklWo43x1QgG4eqK68Uptkm71pAOWZ
nnPGmfaMlFVGcTwGIwvt+tkwe6nlv7nirVfRegBvtfpvhCWSHKy0M+smvyjVcfIR
BuFTswG74JYrbkoMjk7MMKra9O137btZ7hLBJy9WWXr5rkMZzo1dofCOdULapw+I
YIPinqyTJ/OH86fzNy2dIfUD3KkSj5BtKShC7B7ez4NvsXUVU1aeG4hSixIJTTYi
gCqdkW2erijB2uUFrwPj/tqXq7AoabDCp0acv6RHWd0tymmcg4SpdDsn+4gPtlU4
u9gMOxc8WWaVS0sJs+xYRA8JJ5tF4ObeM4uadwPcpJHGqs9vSuL4eCtokr93aXdy
RSxIq9J6oF+UHU3meE+3G8JhAOPRmmzCtj60FMRo2NrtLCWWEbT4VMSnL3++867u
rci89NQWoL21XXjJVIImjqbbAPvWSAuuOnx+DSnrOcdbYmMef1DanOzjGGkefV35
Ka3sb5HbWLp/whQEGSJDN6GteV34cv2ZZudtwAUJ4exoZd75twrt3XFpGW/PUxoy
BkdoAtjqx0w3JUN9rPgEiqi4yUhQTj/ZsMnTQtq4F0a2V3Nk+WZRHmDHGYjJraU7
VGMV226o7tghsys0hYv5DmDHeDuPh8CKAvV4QCYMmqM1I7pfJVYNT4RuQnunuY17
m94btQ+CLZlYITpic6KSP823WqQh+EyacuvoIfZoQj4yEMj5Fc8f5R2ZZ1+eLQkS
iZP4kypIyhrIAmHep9CwTcaqrmtYbBcYuG2b+HUFXGtDYJfjV+hIjsQtDriP6pTR
1eDocQYcSTCbtOct5piSjq+SF/Q9KcLa32Xw22myuoa2cjbn7PIewfaccBARi7EO
f1C2iRHRHHJG2dwD7SBk5zA9ist9bizBVzqKdhTUfe7SeNFL9u7f/ZlgIEv8j1JD
J/4+B+hbhhVFdcwjOD9ANzqYVruOGY99va6g1mcspjq8ZEia184Es0ExpzG244/x
ng6WpHO9oqBp8onDYdq+Aqg3KiopxpRNaOVYuzMaIRkLF7lcbk0aVzzUDCCTLlaq
6Pk4ySKVHNIENv1o7dk9WJWQ+kWCTs0TUKn0Y9DdKOP40LGrnlNZYe1J0VrXhrhx
ji8uJ6Vfc5WEhqRYG9o7j+G/rCyK0ZW0VBNZc6ETq2EpPJWl9a23tg3KF8BI1Bz+
g+alYouR8ROHnSYkqc4ElPJdsTSlk+QF7kouNE1ZG3lTD0lrqwkcCnFqSlLigJZT
4mPbHW3Q1I++dSyTv54vbFdURkf+5Pydh8eGDT+oyF5W40nf0YmACgnA7TfrmFw+
VyIIIMFlkLDXfPFoLDMI/J6ZKrbQ9/NXfQxuLce3Y4DAxAS7HcTb0+bjVNuHLvNG
r4cD2Ottp+4bL9KcmqG679UtWHBP53+AYn03JpbDq/+fBA33EOduPbjaU19K1c+g
WPqv2nMOkkk0batwEeoJWXPn5ZEHjowgEK0Q4skf3n2x2cS+DMSjFbM2rSvovm83
rVBgdJ/GVjCuk/zmglXVZZJcWH4hPstXWCjabC5QVkYAE5WZUEWlRGVGDejO4FXM
VHZeaVafr2nLRkihWq9hrfqyJwYZ9+xzq/pYD+ZaAwrsll+Pi+MBGIuY9beFIEzF
Nt7Asom3VHmbyjslsWEYXqWMTUxUUJwxGw/eEafMykY3DxXi/i019YexboGV9s44
2nfW+KKQj0334h3IfkYrYBKmoCsgFUN6Enk85vPab8Zo/FF3Z/04gjFOwaegpMGd
r+WIT9qhp3AQ9+5kcysq3vFNZt4vtVLLc+hmgOy9ekjO6eOxqVAMU2yI6SjIv499
2lfX6oj0b2QoY/TqL5YI9CjFLCgQAsgl94TVZmSeX4/xaQcqS/AgYT8H4e0L61l7
yf6JSXRWy3f9rn5XeESC4w9bINAu20kmZISqszXVrMI31gF3hYecTckjw7dxvy6m
boSKJRz4evh3zvdRs0iE/AzYKkY11RQU1MdNpvDVr89AUnZsW8s7Q46AiCxWf4wI
KKaD1c3Mo+K4ekyMdUKPCQcXRwGCZIkSjSHmHRstGv6JmZqvZh1I+2QObn5L7DPf
xYA206IvYMhIwts00bqQ9pgkrCL71L0wIfoet5iVVjLjG2BCogRjwf8sdoQ2VmSJ
Wvq4NcWU0w6M06tM70ZiC0jSakMPtVusXxAxwXzS1VRNhXAL2QIGAUnGj+s2gtwK
efwY3utF6rGlznvQtGQiOy+UnwlEt6Aw6wApI1KFAweRsJKUgEdaRqgiHc3iGXKd
bq3RnAcSjKfCqaUK+VkGNhOWn1/S/IHjw/YMAaRlaD4Ir+LLGsrRQG93LX1kxJ0s
E0yrn81EDKJ5XI1+CnHyO9AC71a3BfukBz+FSbBPvbCxzzldySBifY9et9cPYkZH
HEviTyK9TvhqYem0T6x5rr4UJrd2cNIEXADU6h35wfmESNcl9S7aS2CCuSj5ANe2
tVlCqlSqmWxTMC3io1nzSjDQVx/Ac0W4zcPnR360sUuxR9/ZV3BvtGUffWxxet8k
gaACOBSrz3Sck/mLX5ZQrrRn8uIQ89RTRlUvlFmrZOeha/wzUlPKKkX368KqeDwX
teqNq5nrnqMFOvDte732AA2a89yJ3jnJIa91EUKWiXv+8OF38uRBqRQKUP3gclgZ
EWsDTtIE9ibBr7a/5FdJBp2gcIpg/8C2aRDKSIPw4CN8NbT8kgUCv55CI2KA5++L
C1TTJzm7PLOzn4ojFmg0avrqyo53DZBxEyWRCpcsKCBkci5Jyz2IsNn7njVZrUrf
7XL9sjRtysXfX1kOAsR9S/gXGqZanXbITtFMRckbpC+Dp2AsZZW5P9B/xI2Gjpej
VvPcMGbQG2nWc+8JO1yAbf1Wz1EdExb5Vy3XTM7LiEaDGT8l4V95q7NFKg3hzCY4
GC7Dcw+v4tQDW5KJ6axgRaV1btDG0kViBizMjiAz/CFQ/oLfVcHGThxXj0xl3e03
higXp3EsGw9pD3XoRDy9dwxRPCHX6CBs4Ze/ue0+w0fKpwfyqecnQtnwruILzRRr
1yspZwfmJ07J1A6sciGFL2tEimqNV5QEAAA58Pd8CrqDhu+DU5qf2Z6Gva25//nX
OXb09p4FM8ApHFGXG+pGxbtnEVi2o3yKZX9QcRm1wC3kesvBQ6B4wa1d6YkqnaxO
0CnbJlTE721y874sVbmGW6kMdzwvZxxMzJQvl36b6idgedDJqHLsnRitssTZMKCz
K7ElqoDKuv7DI0ddWaC0bJhBJ2mrLF13ijg42oo1IAF44tE3Tpda0n0OQJDZcMUu
BLAt/G53r73aHz/1nnBpeOuJhvx7ZTnMKCcXA9wB7V7XonYQkjdDdO3RA25QWgDT
XfMSAjx3uOfmFpgTOgWTtF1SuiHawFeyFrx9J96n3GrSv4zTLumgOdHPId8qftV2
d3r9Dqb/BM47zgciAdD1d90h/tVwqiMUz6xZ1FtQR8PNTsmxMJjLG22yS3tWhI/g
zqAkLC4fL800uzxXZazblNLDL3IWzgQyDrc/OWlfftPmW6vLZlU9EqkirahDy50Y
j1Pk2vgXuAGGNyn2mwbX4yPX1pWQN/JN8+UcL5fg6fcTt2kQDnsjrT7DdFp/vZ/B
Dg1DxJyIlqEEAkCMWT+Zxc3Y+19AJ/94tDHio0xpOya1IWfuYRzilXssGKoM7/os
2KWDC7t1dChb44LTtJ0mxqlH3lCPv9WVHjw2FAB1h3s7dDAVeFePgqq+J1A4MD7s
b1oiAcmvTVPwJojXslbmaxGlbKO1nUsH5odhP3+bwnKTxvXr5tcUNcLVcsyk+9Dg
qkWErUUWU5IDqD06GVHjvk9hXNz95eqmzIfdMBjA8iiyromwkIuVxAQHkCT8UYPZ
Ic6f3A/Uxji1PpsgWBEMsO/z+Lzx8kvEnmSrn4oSkAR1KuefADlhca/3VcsnGsdG
aSCG1c11QSA26XS2LxAbjHnN5r7KcUnAKOBIdrYLN2kADuOGjwoxXBRNMR61P3Aj
ORrkIY0oCl8zv0zG4i791jyRUYRyBee2o763FRZFdh3QD41M0hM0zMavjCF5g2Ss
ikBgoG1zt7+NrXyAd30VRHpeuCtVebZrmteGQWnhmjVRdyTZUR6//NmqPfv3s7A2
3lcCgXURcQGCggLXgwaXlSWyhYkqxPd4RQEly4Y9nA0JGmKHLq0JHIDzz77Jmtil
yrnRP/ZFabpnvjT7wC236P2AvrVXk5CbFKn2QrXO3rFViq9MFBqDn37g3FIvfDpL
Yxs5IVYscAvKaus4+lUUzol/OMEgorS0SB6ySklBnsiYqt4B042Z4xenVD5lGq+r
YvyrrX3wcAO91KiM1xyHioUvuaY+BbhPjTYn+th7RmcJXKscboTkZKfkS91ltRXT
y7uD8mYWjNkuKbxsfJH0a77qGJAy/iqtLPuy3IMeqczDdQAvMCRyA62jH6qiIneQ
gUOTNdFZo3rGrAM1whRa3GFB6pwyQf6PsBadPMQ6FD/0gcfH6JqRDhfq4iTEeaxG
P4yTUne8eYdgyyF+gc7ZjtZMDtYUs/hxRjm8FBYKDCfWdNv4bbyHjMGmyYsp5PjG
oJMxNwksVpL1VfpHrFjU3P3OPiS3/t+FsL4iXBTOwD9wMvlx+dTfNwz0+arqYhAn
lcxoB6L9I8OtMTgo2VdUReZ8aonssW0qR5GRWNEqBGFQYVfqr6X/lGNjGzVsSu5+
/KobfyKn9hCWxfuy6a+gNJ2SVDuf9m4xYJyjrVi6WIZ+kpcOgCzXMlGU8ET5awP+
hc5WAMGeLRpNtdoqI944i1zZOlantr6aYC7I02pPRgDuHMv1aK70eZxNZhaQ/80y
J/AGRERJ4epjLCvG9VxeIZaobKdg05/wdxmDjA1TXL3EarW15j9Im+6a0RZTI0jw
+eHN/7pncEP+jQscCtHfIm0iZsF2GxAAkwmZ/bqGLJ9xvR3z190CKCdgI1ZXMDtG
v46CHmv53ZNzVQF3xNOLWS+1ad+EIKk4e3jchS+7D4/PHoTYhfbc9v091GitIBHf
Pmuv1EiXAtBJgy5pI5QMHAOKPx92keO+rgniptOvp/nut7qxgufTZ4LP8l5Cg/O3
VIoYodpCHdnCHELlksLUijjcll+snKq0fbLVJKce0aJJxi4HgWQqFdaU6uj8zHES
x3wHsXBUOpcZrn4MpN5Y8s9W0sQDZW9ZjQoT+/sjRKjNWtoEAS3IzyYRCUv9jhFm
MxeWZ/LFiccE4gjt78voUpYSOXJsZ0cm/4TXluTpJH6u8kRXBliKv85zUlQMFFyj
XnQv3a8zF8woHe45aSQ/cbs1yEUsp9dEV4foXeBaN9DMNdoIKRSiaYKJhTzQbMrr
R6d4XatrhkDeloAF0fRSQ2C340wqfzRuvGa5ShZMV7Y9BVfHmxRFcQD4hlDXvcFG
SBQ1d6bF7cfoYjDv9S+bTkt9ybPyTHBgviTAfgj4hJibH/w5DPLUwsFKHjy2okzu
3oA5mrAZdsP80ViY5qQ9IkUsxdrdSJWsondHgJTWQ3pEuostX5KDsJOp6Cqe66o7
tfeyeMeWjZwKTf7b2Qf1860IFnokPoDBrJ4IXdflTOqaTu3hPw5i3STcLWUJnMK9
VKDsE3S+4m+sjnzVI1dLGsjLASxZNqRzM+suMx3hv8JrUFmzIHdx+eVd17Ga2xIB
eECDROa+rON/Xu71LZLcqADR3bROoxFqkyorzYWPL39XuUgiRD/6BvAWp8RMHmZZ
RKNKJp+0hITQMLMx6WMkxclFKkDFd06yDwJV3oevsgu3V++LU9HDB+ssDl4KtcuW
fsPaK9LdTLTqHEy4hGU46YoquN0l4dINVLDrvADMkDS98TtEqs0bNesF7c4bayQa
F/NAjOMr58OPqFtRUexI5HGUjUW8uAu4MPI5ulS7/jPF3CzkE2zQaVI7Q5oPJMYZ
N/g8LsTRtlpnKE+a2EMzxeASQ5iNhQa03ixn8mFbd+w3myclW6Bl9xWS5wpuetTG
iz+9rw/eWpwnWyUBenEPztzZvXtCYc8ttf6CFGQBxoS6QJRcEFkDK6Zcgbn7GF2h
+TTPUxDgbP1XsmkwrBSK/D1W0BY7J8OLgWpPKCsLS4cN/JfFO+W1QLMkeyA/Lm6Z
yl6KQT5IiWW4+cJHn6uEvBRuT8Von2EBV/aXyh2WVwcv/PmsQkq1oFKCpghzusjT
kL1zmolK7ujEScn9SKAh0fyG5uLO3rKaCEwf+6VQ9zAQAedRgqdW142Gg4L14RGu
I1QvKX6todvjicN7tR79aK+F9O6FbgDK6Xk/ULjja0CpMwNNcToHl+5x6Ya/kWh2
3NLMItf1bRxCqmFi8QGXQnTgyZVkFlu5ByCHJ6Wn3vvkUvWDyblO5A6moWrWLfvF
vXP7zzA14FHK6RM0T2lDHZP8uaMs0BRyEc69RPCNX/YSyir00JkUAAPyiUOmjfMH
TPykmus1j7P8NqVbwKirg5OYRvZ5hV/p+kve2EZ3Ju5NuNSL5s6VgUo4AC+TeV9V
dkEGGJux0CQ97pq9QJ4cqnFKg2MvNxk+A/7zSJ68bwuVJXG3PZqR4m2pRROvcQh/
Zo1orOK2ho3avuGK78pb8rRnLHq9fJlE5b79pqgmRSIVEGQxKCwV7gtSMbXsUeJx
FQ606D0G0p+HPZUZmbRPUNGdYCmn0A/Ei7Y6VDhxd4BOHBX1VNZoHg4N6N9D20Gp
ljA4Xfd2qioat+rqgDUc8JEK6FId3T9o5BvZYP9WGLK6Nhsd+83htudJgHpKJtel
cVcfsloJtInxiXfo2MfWR+p+VhEADaJJRIMuQ7UKYKMfHLaOlE5nmQJ5jrntY2To
ho9h5CMRdwizMQlHZ8pf2gDeSAXSMouUnZp8ww8F2t9+FEWLdARRCQxCRQQPrwh0
UD79+9T1bHKuyXwZS01CwUYdYpYwDHGdW6xFytEalol06JAzfPqNNnSQSDNvpsyC
mfUz2cGS0PJ79piuk/ZnR5Z+c0Z+eO0gsYAFlOPaGQhNsSKWV4RPBp7FM7HEJUGL
Na0dU0hwmP34BzFDKaMJ+LCOvxEDVUHtvAkLT4UK0Y9bt4S/dA8hMHwQBrcnc9kz
Js3MGftV2zv+enO2e6CbmPGPHF7wp2mf++JXk8imQicrY/IAKwFVl15w7UXLcdo4
2uBpE/d6ORFcw2BQpU2JvNexcCP1vxMEyuHgLi9FDk6s/tx85mtKT6aZYG9O0nx1
d72zPN6iFefNB/hHUf1VisxAaN1R4K52dpRfd/68sGESP43Yqe9FjpCtOjXJmfbH
h63w/eOgVYK94iX8s+z8RAZlJOF6a9gBkgtOY+m3ANFiJycWivDgnR/seU0ulQzt
fyv0PTf2t6KsuIg8XovBJPi+xQCQWwz3SjQ4xREHg3izTdb5kPCqWtp+JrJMXAM0
yQhLICXkFagM0I509hmzLBRpHEMpSAqSO56aWc90FtcBjMIkK0Zbh46bb+CdTJAo
E7ww7u8NVYWSe54crzBr4taLeABw0B1ycNJRzulv4YoG6eafjnWtBQk8ZC1iHMps
/hEGeBtso5IvIsr6UuLBvn4+rpQaofAuxL+7w+ZJ0u9UQWRO77Vn0/cotI4FZF/C
ouf5AXowZBi0Go5MU9HSii99QUwhjUF8UlAejEA/WVVAWCQEnVSQfD7DG10dEz+C
sNNCPwbqLGXHbeAFvlDmDQVbkh+FEFFJOgQY+Ix9EVckQGT8z5wkpIxWNp7ex+aI
j4yZn1BYC595gmtg6ACJDpVUi0WAf4RxKLwfBm3tC7vb79vF9DRdGft/mpySE9sz
hfDlUPeq1UkLEjS9YEhXCLU4iYFtBX8Dr0ULgWCkMI5z26MRG5wVifxmRLc48ed9
Wve9UX5vnjqLy8tfOC/Vt6P/D2RXJ7spAaI8fe8GzArbpnjUuJEx4p+J0KVtVdSS
VBZLggWaMzWHz9VRktWUd3XeJFd8f5vmgaLcTa7A1nBRPWh2rU1++7MeHU4MiuR+
lC1QuHl5ZSWmfyr0wuj+49qNT9Cx1nIXh759ivAdHU3g1UbsqNo2i9n1JJ7sQ6gf
c3deyT5TUb+zVfgUWAbA6FBBx/2qdIZWzh91ksXxBtZ+Fmgi6FnCZDt9Y1JvGZAK
MoA7aSkd7e766Knw838Cj8YOPkonutRCIMw3M8vwXbmf9piXlyZlOoXm4yp8zzoj
FJXNdOX22oEvH5jISDzKnZDIN0EALbCJR5kUoAYyxBTHQaxqW/SUC7gE3bUz/Zbv
GXGBm4QXD/FHD52xagA5sUfls6gd/MonKtFGb8WuA7g00aHxd81urTL9dOwSpzC6
H0z3JKiu34jkGKsPwgTxVRl6tmJlK2l7O5bi8in3+eGI5Y7ywkkpnJrXGxA2qmen
hrAaUQ6k6MTTY++tpj0Qg1ea8r0yY7xnKdYHGAbbrX2atGBgaXljXammb5qkuuLp
4G7xW1nDjP8kaBxVIs0DQftx+a1iAyVkXBGvTIYqyRU1X6z0X/94+SRwmKc4Lz9L
0L+J5dK2Hvhg3OXXljNx8cT/LPrYtJOp6nX/Bh5cnV3uqnE54Ub2048PSpDiCv7o
+Z3i1l9pt8Q3WSI6Kv604rrDKP0rV9pKsTxBfGd6lDmFDRULZKMpjdWJB1u6OU2r
hbTzCGZPgklTOdoUZN14AkWFQfs5PRcbaediU7UzG1pyE/J7Gaal9P+EckCkbbmQ
vpmosXxIHX7Mfygt/qLAB90mH9oCl4fvj5OtM/9rKNX96zQLjWvksX5RYiU/RuJf
pExrzonPJHj4SCPxGoeQSN3Ths4m+xU5PVddjA5F4UHpT9WMzvkldRiWwiriV1kC
8Nwy/8lejzSG1xQA9cPm/Bc3PsfL1tQIFVEWGu4kiGttAjM/9bZC3sPK9FGm6k54
8nZhcHbCD/jaNUvRly6qe/8Q225TTlsAuSddacs4A9bO9m+KbKCXQxAAVdIvjQTS
GP2kjVB09L98ldSkPWivg2DhirjltIvOrqIwVslj6G2Kz3wN6TlzkyZiHyoEE03g
EitUJE3cxTQ9TBK6S95T5NeYsflL5/FvamzMaaS0Jdpm3WwdrjG1DOgoxIV4t5iU
LoxJ0ytd8pyN2ThIEswP+UEVNp3zE6iPI+UGwii8EitOLFxksNAO4/jKRtFggwp2
BNFJ7RC6PY+h+gwuFZbeN74sU7UUALfBrUvOlIR8MA1207B9VQfTknHfbM/mTnBp
AoXN4cfrBni8ULiIEKgAevSnHMe9aDTbyPrm36phZLiqkeKfaK3PiZ+N1ZVCB3GC
JkA+J12clKNHEwEQGaEsMd74mE5BZtQCaK1aPQHdi/TcBfwt5+G0y1I7bqQNM7+0
5dV8qYXAJZCNsmpO3t1lCZIoa607XbsiBjJo1HBXykeCAlcQLYMxRwxnxFOF9DnW
CeU1EV0m1eGkWCWWXp1rk+PWSDLYIlJTvz7NdvN2IvJRPqIkoElBVNcRTlrcdpoN
w1f4OEczBYINJyF3GhClWM39T/msJjTk5UaIy0xBDclniEYYhWocTRBUqTSp84I0
1NOi6o+spAmtCG2H62nD2fLw03omV8bMDXBiP2KHz/hkqjnrvn3YJstKRPLq3o6D
PdnHVGTu0BzhXEzJ+BE0zKAx9P61rlCCrZXLeL1nNv6Iobi4NyBVsa3c5fLE1XRt
kRF25ZzawrEfUj5BrtD3TT0rGuoC9iAOqWoOhRR0so+U1fej0jx+NhygG+r9tgq/
DU3j0r2U0/IVS4lWXZrG4lwyIJQY5+psCeNL/rdAVy96A1RzamEzqoY2s0DBv1WZ
tA1lT4RjeeUnLgW8Dt3iwchpEqzLWfMqiKAj+xMqRysRyfukutMGRW1TBIEfFO6U
bO8VKgmE+oNVx6iwv5kVvqcaI3LpOSmyMZ/PBlOk8uk2Ns/0HM6PM98G4BlHnfwx
antHtfH3nkozWFoGjZRpONuPqHEmFqGwmvhlkaf/xnDezNjuW8GVWd65FsnnSh8D
Bn6LYAnqtN1cntxxPpefp5IXANu2XKC43xpm8t9piU4mLEt0tzrMlMhvLkLgC1IU
vgDAxJRx219OCXeC08tTYWCEaOQziPI1WyhZp2eS/l1gPKYRO6WrbE3pk7Owqo3A
+KNEXejg5DnUHyZXiw4KWxrTbAkHFRexWdXXkSu76/xSSRC5mjS08BgFgZZpj+tG
7TfCvCKpEBc1Gx6eTMcE6vUS8kIJMZX+kb6fzFdhCmv2VFmlzpvivF56SRHhU6yT
e3TmPQy7tCtim/sZOVOoXrBN7yXUkTFGYkvWSTyPpXpMaqmwsmFRAWkEygrrl5zI
OJWxt3w3iA4io0diE3EpSVWdYjbXTu4B2xWM00rIIFqb9D9aFDM7Ihsly1NKgMql
PctCy/qXn5w3l1dfNBiUv96wX868rR2acAj39wrxE1/NDXmlywOW8BWcxC54bAwx
qFarZIol46KRU/1AvWzhysu8ArAC91MnE25oU1ZmseyscdyhWRe5wFQX8HtfFWZb
kZWPqbzRLnP4lAXAUq6BRac+6KVMLBKpIL6uItso73jPwjBKgMobL+Y8UqDEbC0U
UvbyR3zoK0yqWYANDNS+7P7JYXT//KsvaiDFFbdoe5EAiUOuxi9XUFXm6i4TTwqH
o289udCOWwSTt7u26mbYYqanikVtr+/liNQgvVM11xWqTZA6RewDqSaA4SDAAia6
E2wjtCXaaLIP/ev4MZ5h6kzY1l8d3PNfmFEwVS15ywXx+QGYOoN5bIIKoMj9HZfd
ViTiEcsAR2Rn1EeYDbbmYeRvKh4WhAU42t3V+BrL466NpFzfyk6pKVy85L0CR2Ny
emIFsjr+YybEy7TveSnUszsia6rwfJJuzLKfZ1GKawgJw04PPm1G/jlXOjJKrgwJ
FM+sT7oowOlHAvv038gPUGvP312ABYD+dTCU13dGx9q1FSKTZuG8/QcJYyvvM03/
3j7M9WD8Q/Vudi9QVT3lOXVsAotPRjxl3iwZq29Azc1bUXMmfqzHOMkxAA3ImVac
LDd4HlcYhAmKYIJ1ompp7IwUMQ5LSz5koBnqOcKf8AXRhq7Fx2gcUIfatzqsz6OJ
VKuj+/NaWoxThfDjG9lmqnRSnnw6A/0uMWz4SQ7JoHdXziKSaurcltPIdLaRybgz
Is4ZlJDSIcvfslGpM2wx4ZIQMoauxoJJtLaw/K+KgeMKwpB+7+hUKQrumrVwlSYk
duYE7nPcWpgbZ/rmVFTHuW+CXM2fkIPARFuGN7bQQee+GENZJrUd83Uhpv08Y/Ia
OMIszsGvkl3Z3N/dyLal8KZ5ySwUtP9r16DKcwkCm9wQfTmnjCmt3fWYPb8/IqJF
eNNji2j2+uDLVLZL2rD5bhaTrDRgOGLeJIMAim0uxMxSAfoL4xeJefk1dR98hQOi
jUhaudoOcxa2MTVtXXWKx+n1ua2zWKo9Fr1CriwOxqhblv0AFkqVvV/MXERnIshE
cAlNZhSOW83L97FTKy8h/OwUKrRi9ShSZd5VLYFjAyZdZsv/KLBA1CaevCECjpBr
4Ki6T4OnE1oOz3GRP8C3nV/Z5pJg93NLKR1A6jsDhr66L/8NWrgETTyor4vfmMrH
bkxLzlIG+n7inkK8kP2J8L5iz7pqaGOjt8JDuF70GHO6O6/CTaWfWZBGjqT5rAiF
JUwDtd7ww3/D2fp2TPm3a+cv0zWiUjD/8XtRFaMRjHSMIK9DsB67DkxvNbqNozr3
aQ7SV9aCO4nGjZpe8ZuBBp6pCBIsnpOhP54F/TWAntnn/Ada0Llv1wTgz5BBZmdh
7jzTtJ5Kxv+sIX7j8Kt+GXWqxZ4d3TtaFWWyTc7hEMy4P4EvFDvzkcYvD4YowlQ3
4cc1EvkOOABbg1ktn6nZhYM/aIDc+mzbJQlk9IM8CJYUFtieOLUUTwI/xUVVeMk5
GJ/ZVY+I/QqBmdPLCvc5FBc9r5tw/wrXc4a4qyfcQ+9J2P+jyiNcFC2jcC1IE8Tc
wkkuKV/Qq6xUv2m+Ako4C5lLyWqWhZPqOVxWG9xlsq69839OD8JDo/zPGETE5rz1
EM8pjOSyMqhSI2UrB3eLDFYV86KipKgauHUMcv9rSOfGmA4Xdry6Ot3gPQtDHXbB
hfyKX1SsIPEmCV/c083ggal7IwUxH+cgkULFVnclwuPnZlih1XGIFLyl90/a3JWA
+4wN5nIx03QSGHuulQjT4pUADzSafTtQvtVyXiFO3nRij/JvBwkH4mrsgcknCf8D
AA/gpaHZw8UxEENXp3EWIKjPN5eI7W2lleRVp2T+VdPrv3NP0uMyIxCIBBWzSBwD
9NCvEP//I7DcI31YDOoUfw03QezpA50wBDePcEa6bH7HaMjU9iioi/UL/EfiK+oB
NR7/reQSF+PUdw8cqa9jcEwuXYx/wTdPQaJ912mHKClYHK4I6P8xGr4wASnIlcw9
BFv8E2eCzEeenH9xI3GtBFSEcntDaw8OZkj66Lsee13XcErkM+Uy9ER4Rbe4kJ6S
EMByP9iN3FLcEBv5lzM+xDG7yk0KM88C1odSCHxo9HE3+/4siYK8y2EztkTwyGak
EWnu+E5xswyYXv18bAMhIDfvqpBSmM40FYs1jQdbpoljLZWcPPdk9LyeT3Gc7nqY
+EqXeXDiCmqkFOIBfAA29ak+JP/V+SJtdPXKh+RmtC+pvQITC2wr5zHn8Bs5cgL1
UvTa2g2nv2LmVHt1e6jgIuhAQ4FNXKXbSm5eGiaJI56sbobfJ3ZsZBikOskuZkPy
ViwBHYOhDf71gyLvojcR9/oUO3rXUsRLo5/gMzwJQ4z/kmhPL+UKzA3DNjElngNt
MlqWK69wIuua9yPKJi4m5QuDNoDhx+EGNaTzDJpHNNWjyuHlz4qHJAr9eAiMICQU
ijN+yCTKoDX1P5uxU7FhdPscWlrVM1VzulP22+PwMLYn3JC7XrA4KQUyJV5pN4AS
VwUCTJFShoOP8gILMXjW3JM/z0yPCsBAvJCtxk163msV5o7hMlcAbhe0IJupWXRo
jtJ7ELzqxirGDHAsEPdHPUeRsHvvKDTUHr1Rzd3+I3CnR6ZRkxnHhEZ8wSBAnpK+
iI74NZgnfkRR1ZJ95lnlwkoAk/SLXeaNU3sUwfEYmGAFwOZTnOP3aoQCZdi3epoJ
Ug49pVNYgEG4+AfDy2PaAievPiln1Rx8J01Fbye6GsVKTHUi3cVtJ4edvmVGdYRr
lVl44mIMDS708mmHzYDFoOqGFXAeIzOgKkEVlhzX1/Y6AReuUHoCqzjaHC7N4xyS
qMtDAbsKmaqS8yEhFR04CS4jNjjlNOMXtpPHsOdSszT9qCoCcPyoFPRGdO/ZtDLS
TsT5xUepM/NQMC4SNjR6sVX/uErpb8hecycpRNCrWhV76jXw+MsefTS1xjwJ5Yq/
y6LdPSvensEdxnEJpShbOlPiKbr9tG9vGAvjLSz0GV3f4Yvcr8YgDmjCqqjLL0Tq
9JlEYyZmLOaQJnyhxuspFQfSKy7MDM21MNiZCFTGHm+kBk7/Pg7K/Y0hAkXjguO3
4GWvFXpP+3u241gBzFes1NcMAxqBo8NbM6B9yO6crCTxTStPZH8KgIhRGJotWY1m
89buEypIVZgIXhkLYXNuCUREkYDDvLpdfJUiswGXqB5/4SbZrPKY0apXzTF7aRW9
nxLq8H9Xq3Z34UnfnF6ZpI/ePbtB6QeCvuE7CPNtXI3XrfcvVo907Iuc1sqz0PFa
fpQFRiBS5tRH7G8aUqcdUZb0Xkvl23PhlWeJ68u92NzplT8enjqLbhaKrjQkStNU
+uNfVf0VwVyzP0V5Fujz9es4IXXDGhjZippUtTMfoDBfRFz/Ic+vDRwek2mSs6Jw
sgJxmcpCLqQdbD2da3PJhxTbIKhYF4AjYvHTxpuYWrBo0RFSU2gl6Z7uY4++Utk/
0/eYA4joT/+eFr4feLWD6XSUCvZhTqTfrWlmuyR8bQEDtXg40NdmoJ/rwvZTgzJR
2NeV+wsjWp1UheIZzJAaCIYIFSw1c7NCRETl9eFKuD6qzLD7eHDYb2g4adlBH5oy
Xl5SlOA+/5Ac6DR/jPzsOrYsekDVL2vQZ1F3dIN573u6CfcfPLErUGVUi9Xga9XQ
17tsCfx0dwg6jLrWyVXTyEUDhBJfLAVchgtY56286E0949Y01e04txOp8+b9h+MK
6LXFsQHaAsPf8BLb9nQksG5bOiu9USHXazuZij4QbAbVO/0uZ/m9Fp6ymZE2D3jh
Dps+cKijylrQXI5Gc8RrFAveIgDJ4eJfxs92ko46KTUwFTQ4L5oPFHxMseZWG5Zw
+cCHCR35n+qudZiUq6JU8SxsYIS3bRo2cMouzeRn5ZjFcgNDDFdw2CNcV1GtwuH4
HJUfQPTE7P6E5m5sQXG8rVY7Wyg3VP+qcX5YzPIrCCz995TIZ+UIdLP2Qy2j+f98
QmaIw2A1+zh8PL0QX4d4nJDlaeJMLGC5U+2FIP9YWE7ffGkPGQTj6ZLmqrJBxrJ1
wwXizMswciodblx/wp2oJiIHTWFlodEv3S+A5eBJazUDZiDcZiqMQK25OoP9O11D
LVqSWZA21rDs/V819P1ris3DN1yuCUBSVsBUPYw/zt77UnDaP+P1u2uQHNn/VzuR
/CNWodYZgX5rXCYGUa1YAZoQ2y29lZKo33eq2rM9PIOA5sKwAPnkIiXwkjBIaSE5
jLfkj/2T2d4Gwd1UP+f03D3TWrAyEQ6BfI0cnoFcYzOvKf3fok3owpCAaA2RouRp
3Vl/5613VBpNCTSXaXH3OCi9L74f7gL5BbRtj0TSqSeNS3W+muA1xffhQh011nNz
5hnUC6FLISS66NdZlcrMUdCCp2XGykZkJrEgOc7u0kmPaowbLkhJUqZE36gCVNLh
b/UFhNW18qJ5SuaZn4rtwtWMIoRK97WwLtgnGxLUHzTfQb2lFu5W3bNeBet6QZhC
Umh/iiM6APdHbE+jTEbLtzTqKkKYPV2PA2t6dgUizxiUCcCytSKVw5PM54yrrFjA
lxK90ulG4rgVvxsHDsqN700qVOo2/mJGTYAdS0Ze+EMNP0s9WwDB8xWtu1l0FLtT
5ZmuYPYcPsbU+XFpMwv9DsyZRHOq66P4LQUbTWqx6675NFPd5qQcifMM7dYNZYNk
RZFI8roi9Ng6K2c3sPoPKlH6z2/ENI4N/M5xYMkyWUAIabvMP4Kikn3t1cklRLB7
Bkby8ooHN4WcqiVYcuqzGc3JVI2R5+EFMXSW66XE+lPoSFTzQB7z1Qy5nmvHyzHQ
J8cADMUBahXPqflB/xDFhh8dzXG9NvmkdUMBPAg9DyO8i+gBqryqIRzU3+hVJfan
4sTvdJ544GIKW3RrqRABvjAR6jkWf+nYSKLW6adeMm79nZwVsDC5er8PXwaUCrsK
3DE8GITlbgKPDAdGgkgDBEhjt264rzI1sCRKRh3JAWKAN1Q3m9YlbcZcWb2Y8D/9
N1U99jX6r3xyeLv57OCuwGfZD4WdIrb7Fvk1gAxFF7P9B6/VTeA+/28fdHik1Ou0
E3YadNp4taoDfd550Kz7p4T/Ge82pF6Y9x6D7uJWAoPN0pOXpbQ4BROqsg9uwyM8
IcQkL+ZAwF/bYg0O9g9NKSydIV9C0erS+GCyt+yI6qRaLdl0PIfDy3HC+GWrUrTn
V+8lVGuRV+dlc1UdSigfaqPSrZm3XYX5YViDNKKv/KRNFLTZMZ9ccwbJMtwJ/IaE
kY7wtEKn44g7vChcyBT/Yw+df1gYZCulvMk0xOuRGwXQO9m1JMynD7QNUqQrtAU+
oXHqyPFPHs54D5b0OpQEydUrIjihDGWah9D+B2XCjEzfHVURRoUxlGO9dDJ4ifiQ
Q9vFjiVGCpcL/mnuctdzKzYiH8IxCR0YjSCO2QDSomcwL7P1FwTBGJ3njzz4UpVw
jZD6qRA/JUWWdRi+6cWU6v8aRHJQnFeI7oyhz6c6E8AoIoBvpNIHXYc1r/KPgWbk
+CrWILo/3lU1N1bwJrGu9qZpWAI4A3NeaI+USQbGD/0CJIKUzITKAc98RpKnFrjg
sQeEXjBQoArHxH3uUQKF7AK2zUrcAWEQjkP9lC7k/egTK8cjf7O/EMzJZSjBDiHw
XjqjZ3asMdDK3UH60UOj5yrMqO/ZmucEr6h3DulvNKwt8cM1sIt/bpbOxCInHTpA
k8K1rYeuPAk4+B0OYpFW+jFT7TMvfcBzYtz6vFIYrazWgS6HU62pCBsnrv7pKf8G
o487cNWs9Qt5+Pjv1uOmPUpeLU3hEoGpH2YPuVDw+Xs1Xvpcl1UD9dd+N8vqBm76
/oYaI5zO2uPmi+6ir9W058FdSgPU4YXhV2Tfm5VlxP48wVHJcIP84WC9/vleaaB5
4ePS5lAro2yhL/gmc4mrOwNrKW1Kf+hFoLTkntnN+EZnJHyv5iUI1IbcWlgMstfI
2x/zXpokrsCoKyIMDak7NcjTLf59O9OEzIDQ/g7JODxmfVoYIACHBfxIVnnhUn4Q
pFxY/d3uZ6kFY8BZ/MHotBjRDvuh+1Iuq3yuHxQPWiCWg8PxHvnv/BFToGjvSnCr
6LOZpIurfQkAHR9UQfHXcnrQDde9yXFG9+d7AraTetlsxOTuxzp8fSyTuueczENm
cBSiY018+REpw1eX0dA82IJ27A6TSv59ZcUzJgXTZydfKePfYNom5S62xbQvo9pY
ayJrobDd3JBw9tEa8YdjU7DIHZwudspQV4AwpssKDzzFhaPCplZiVPJCSsz0tzPh
ocCdPppS66Z5JNAncXxyV3zemRi8U5SY3l+0hiZgnBNOxvtR+Frp/wPTCyR9gSHO
JIOIYlcEPSlKyoY4k4NvE5gzHTbg1pOVQMyqhmktsp312ilcBAuncckVRfCRqJTW
Wy0aILEESuATbHj+Ic+4Bs0XXNXqI7Lp9PmTPTuK9s8VsfEC+bg87bBDELs/qBj+
oyba8QVRZbPA2NnmmCugX5j6auYmx4pggASlNPYb2LH9p8H6zvEPls7hD5Pf/I5p
w3tQL6qCuVgYdWQYX3gsgTGjdyg5V1HrqYKQXwe587q3GOq5tZuoSacCOlr0d+d4
b1x6SclE9Ht17gbrCravgmhUG5Qi+AZUME/TGq6mXnNy3vhTqY5i7dbeqLAa8JUT
4D4D6/FL6SJmf3ptos7Vb0rgfpGxMDl3HFRYEioE9nn/cqrwRAZpV8vARVPankK1
6+BiQXTCIFMU61l3+K44HK54IJwZE1TNI3G1apkXjekCrIcoY0qxXKubbY/VyWxY
608Mo4kAwVPkOzDmdn6odNTqBMYnZhznMS8hPj6fJV/Sb5OdlFq1FLNxkXEzeHWR
PkFmhXYATeqhAt3ApUmNzpAMmOK5B3zmYDWA7vGsMSSwmT4sozfn7trbu/wfgu9y
BMvN9S9tlX8IJsQChplLGCgVgMToReYbxFvWoCsp94X3JqoIOvHZXf+KURRywWFL
cyRXbro7nyElejocyznF8oNVyJJqyp+VfWC3IJrrElSdBqC9nL4Zd9frKOtyH5vT
dRsSiHs64fI2/Dy4oErD0h6OPbUixXwazqsGjZ1eoBN5uVDrssgyKh4ITgsk0aKS
EcwEBcDDUBT2qGzInkgZCnY/cH8hX6cvksfrxes8IxpPnS5GEYRVDBK8pUMOCNX/
JKkCeiFrzldbVOuBdAgvNgKZlJGtKU7csjcGE02Z+e4/UWHEJsYxt9DjFL4LVPs8
ygSsLhcn7nnK+Vf1rkuvNYL6Ghr7qksoFvK18h0ZhBBGZcCzpOoaD40FvFNb3/3O
mtUi86H0LBmy9gZ69TcH2CBRCkfFI/uKrgoxGlGtZZi4lQgFIYW3Uv/C6d2hOnRM
pLE/POoG5n16PalMmkz2P6vF/4DdXzFQPs6hsEw1XZ54ojBGezcuFdaDc+KHTATF
2UNN8IGvYXQ+givWxBMcPklH3XxLW4lqiFv5I8iF6USFoongcvz5L2Wmf/OpADS0
iUWHXjLhFkU0PmWrgOhOUDvFDcBe6hoa7q2/18QqnVc48G0VibE/hmGPueeoDUTQ
MURLGheSnDw49+UFZ3doyFfutj1RpXbKAs2HbQ/AhlClzJz++sGkdx9XUbThnkm2
YB1DmEP2S4oXju2AoxunvVsb4GKFkQL4GVpL05EUYpK5Vresrxsg5uKOUh1ucg/b
CAKLq9CwJ2lhQKX2mxeiRSUyL5xI51PqOqdpG1lqK5fPt9eAxupVGILp80KUQr8x
o6q84ncQAXRUlGVdhYaZMPVO0odfYsVIVq2mmm/B4yf1rhCOjglETWPHhcXk5CgA
eQ9oU0irII7wKpoXq92e32VgdbBN+LR7bYU5vU4quKP77NxQOExftmXwxZssG8p+
jPuIv0CyI1XK3bLaFfytL641us6NAZ6WpW9L79vFetK+QtMAOjNYRzjYIGicTSTr
pac4TFaxuecM/OZjGTNaupmhJavz6NLGW5FS3lqF9MUAvBhRQXMOtCu5dCt1xVlL
2Ry0s3KM3KUQ/FBw7XmPdhFV66kfHtrP0WKNZ/aIgDeXZ2Rvo70DVlGyg8Oorjp+
h6xfWRCbK8nfekxu1NsIcfDFbEpHRwR3Uz/t6DYGtKVdulvUypjsxRirnFKUTdjs
fG9T+EoBY4Y26moWY4tzTFjOfDb1EfKGc/E89PjLWCdExi9jmf1BdT6yK/Vo4582
kJtN7hLAwCILtiF43YX8sPJFLk8LPkNO14Mc32kufAtc/d6WBx+PCZm8EnjWTnem
Yuf4sUnUedRzFwYwVzCNP0t4SXN/da139O/bcBPGE010MkJUKPdTRLwPpygxAdXI
71/dKDJ3R722BnSBqooiMR3+DpvgnvmgakrLeu6fAqAJa1KigLILElAq13cSQHFB
QUOCjlox42SnyACUsMyBhaPGgIWLQQjXgU+6+UPOYH0TJqW/v3e9gyZSnspQHFy7
xVNvgjQByF+zY6K7OoLVCVfz+69/sVv4WBVX2GE1i6g8bLxKdZzY59F/HPw+drgo
wPaMdlJaDtNyGPcoiCVzIkwk+TDlCPCSQOOd3zdz81XCsotbPZsrBRlAE+zeOb1Q
O4Dii0mkBRJaycQbgUyTqFt9TlON+A0FIWMoDcpgk3b1K+4A2GbtTFMGkIkyAGLP
KCRw3HNI1P8PXNgVz5okjjeywRjgKTp5pZsEwP6Fubxc6rBkqtL7DwhZJD7DevaZ
hEwoUy/VgA+dGkTjX4MEyAiCWrcUYDUVnQyUCMlZz9WtlvH8FXQw1YfuJAO8EUK4
efYom2Eq3Ix2dXYffgNni4KmEV09OKxrVZ8YNuExLm0GmmzOTSnpZNvWgiuFGW38
sbWuu0mdcf/RtjhTVVtAmVWX8KKhLzMGpfCbXRMc/Xq9Rv5/XLOZHfNK85y3hwev
j6SPkip2/0HJZgq143C5A3B8FgaCVXNDqchfflJ+TC0+hwzLJaicvhY4zDf/YqfF
NTpMWx6idVhs0yMOFDkFRqxlInMeXDR4LUFYvLM9oZpVkXx2e62yklS4aW2Ikh03
XA7uAg+PGwMVkPzI7SQr51ZEQXFdgqBZA4IoetBUMEzpse4e9DDIfcAEBleMK3SQ
L42geLs8kIihs3XPJ5t48yWdVM8PF8xS9VUgXtXyHRyIvOVzibua/ng6lKq5ifgf
dmYucSf9eSVFNEC11NydY8plOjrrV5Y/pgcRi/5ndwr+x0sNxZD/das/KFKRiUOz
gloNAZnXJk3wbFROPdaFTbPGjcEMDpCqDFCwTkBPD1XTD4VMOOimyYE0TNOcg4LD
+S20lBQJmjrSZM2Gsn6PppjBKMm8GAEmJtk38JMDYOZjkI4zIYGgbwLrLVd8JNxA
5nSC0yh3QaUWB+oxfrATyIavyrWihw+B87mWc4AHYB7gwCR9PgqfV2GE8Kz36gr0
UCLrOIvf7khS7ierPko3sAOIIP7ygon28NUIG5+zWz7cxQAV4HSAUWeMPw25q6ll
G8lMATs5eX3+qNOAauOS414+N8aaqQr8fSaxmTpBtiJTEadr+0DR/ErloHzhOz6z
EQBw0jvDUflJLy1gbcFfaqA4QCWJMcgYoWdRVOSdZOgQdLyPD6AcF6DZ1Eb8AjXn
fEVB/cyANHHAKKAeoOTzxUB5KER/ML5/S6w/3trHduibJ8Y0X9jnEq10E1NWqgNq
kKB6D9MPmjL7nBLIbsE2JKyGPPFavZfAwtNL8sakAv/9RNeDjxrpdx56hhFEo5u/
s6i601tyWE2w5dnVLKs8nwGoXpirggNKHtOFQTY3AjWVecuk7ZXFaKKhkiTz1qE8
uS7oxpgpUoXqCQ/3YOA8GMJq3k6R+KGz9TF9ZUVOPqnn0VwZ9nYCyJqwWz/QEZ2r
PyNfvlYwK87hJpknsyvyP2fSp4sgHiVg/q7R5891r1IynePViK8OLgHzJ7jjIAAk
reAetRVzPxxqEBXPFE5zZJWlDvANtADZ1i0sfVUwtvLSJZLhB46eF2gxdj+PUG7u
zYguiB5cP99dqF3sPjambMII9X6JmBAVC2HFLStDonrSL1syfWcX0NTNrrkKtUVT
uxOZ8vWl+bqgdAyFDXzm5xTaPQD4Ec+Cbhi7+XgOK0zi9PXsdURKRKWVNG3WVNJO
mNerAKLgniuV3WhvDrTfNyv46w5/cy6bHDJzx5f+0HNqla2ayGqXGyAGI7l4xfAv
lLccNc5kh0oL/Z1PQENgkU6ThpxE95XJ5h/IDioOkK+kX7NkM+pT1rV0ccFNpz5l
Pq6bUqOG1hyq/V4NC8i8OXFnIwlBhzxnaWRgL4weVXVDRHWx5qVJZ47tLYxTe50D
0nfxUV1xuNbImG09y5dK3ByCsVA0Z0QI5nmjxXGwdyUXS9JaVRzM6y0ywVSEwnCQ
41/tLU7D6M14K3NLMCYSaHUALv7E6dmIbFh0JO5UmYsgZ5pcAknax+F/tjySuTGE
6cEJvTcs0iaGZl/R9CDwatPqXmqhn62qJgSN7zocGl+visbZQru3g6piPkLkN5rw
N1t8/VRRBffV5iOgDRJzFx8OgBDZNZ1xvxYrOZNB+npkogHQ2UXjTDakKBFTTVWQ
NOu4iUn/yYxmERqhx3K0I1dpNsxjpyJtB89d+wEM8Rr+Hkateqfvlwtx7h+yypZJ
F9pfbMdDV0PtcUm8IY3XeEnurzT9wqSIDRBoGrVcBz8XNMr5VhU7IFgRsj5L686e
d5YykHTywPhmhv67HJegdnCwulCa1ndpf9z73wSI1mvoMP3JHuKcKMUC7R6F7F9/
+OxEDbD4qYqAjUkyz0s1HMOQJJQZdsO2/+5ElecnRbGlPFQ4qGsYssosa+s1+5Nl
R3RX5A8VurV9SK8F9BmJ+nhK8wLVZQ/7CSmdfRl+rL+1fls7ScO+4lR4kp0We3mr
UuigFfc1eDm7lIMSevaiX8jL2/RTi1IUog/bFJXELELZwkoxh74hhYXzeDkTUq/u
Yhgb+q4AfyYBZ4u+uagtqHiW5aWK/QjBoZgdWCIG0rgmoHZniQLntgy7p1ctqBMA
xqiOf6UFuc7tUlFFQmsx7eMAKeztX60mt3ZPU7/K7AniPEDcZARFsgCMF5OauZTG
wHIvjwdZrzPDCo3C8/GMcHCnjP6quBMxea3UtIbeU1YUIB3EptqumwZFiRXg6K6l
AKeSAt5drCl2Um4/oTqupD8d+KKQltsq5VppF1YKiqm+ZgRqet/cJEAH/sjnn2Wp
KWoT2IBXJBBlfWhH76/GnjF15pH3VEvDt161uSynmxKkOcBPWNX0RheBVGuAj99m
LMTXxku0n/DAhPfxSrlNHQssO7tVF7VxD3xP6i6wwcgWgCthywLROdTxOs6t3eN6
zFmwctZBKRxbyqe6rAWKZnazcJxA5MSIE2N6tqCK40/t+O2aSwXp8GK4WZnhgwZ2
jxqnCor+CWWthe6i7qm6rxHwXmtoLTtnH4c+epTBOYLQZMECea8YgYG31kvJMH/2
7KIJgXH5Hnme2d0wD7z5ePwBrlnGvG9OFfQ47WdD0vhI1eLgczYp1PP4U1q2UqI+
+Acza+GObI3OGus3k2DvbDkNDygnoOXFAW+H0FTrS1kQPVysQGHPSyGcPr+mQDYE
BLAyFyXYXGVrbkQ3TUkR+3kz8kNGQ7iXhvS4nnXRBvms4fiuCQLNW2gS/ow+OD/P
SpQGYxryxsIHFRsDuTATnYxEY4Oc7EEfDFFi8m1as6tB8nfp7i1ik3Of4apBBcg7
gwNTsO1RpPmA+16gyuNLqos2ZykV1gdtWWpzcBpypaqlXR0BeBKs6/s1pvCmAF0N
HM2YnyUSfioIiNDMv4o1/2laX64rvysyf4PVBSlcI0qrXKO7+Zc2t1+7km5BPcAP
WxZoyUUirZ8QOhXFhr6x6GUkZzMYxSZyh/+RfUk/9Et9MZ7/QENXk+j/Qy9ZrqHB
gcuYpm1+66Pbyi6PnjH+Fl4d9VG5DUuwkq8069kuHyfBs/S7uSpSExLYf45XCGRV
aqfhkRZJYNJS6+X5ZHEdmCK02QkNy5ndiyWDOtF2bsECAogdH1aEczXPmADEzM+3
eBTtUfB/V4hGinOxkwpeu2HM19/3hR18Lq2O7EmIAuv08eNZrBWU+UZlfCYXRChu
TTCkNEcnAlWH95Pn2yrfqqska1HTUIzXuXoRHZBwZTt+te0elE564+85VKXkEs/Q
5MEGMVCX/s/25YKFcp+B2KYD2m9ts969D9Aoh938vQEpJqginLfkflIYQnrzS+6X
EKQ+mhriT2OZHL5fvAOpn7HUUa7bh+0N9tSFf0wtkC2Fjs3wUsp9cg2Knih2XySq
GxBKpmXVBRyVvUlVQzOtIP2U9GtwDHkV/D6PwO36s+NucaXPoaO96jq6m/6Ud/Iw
GX8yQqDyMqvGEiDGJxVrf7hraIpQKbx03rhjFdzio2LYWFphTq3+5sTWg6hiWg0i
k7rXv8787sDxzZABd6Yu66PyLHZNPcHJu3+wc1K2kNJVdAHsZlDw+0Qc15CWRhlC
459B3704ptDjRkkKrufs62WYBR9OxXS+Z8gnFEnCen+XX+zvreEEVp37oYud8RfQ
omI8jyZNJMclGYCM2iL+t3n1wfBLe50kUOmDfsdHvBXZG0tNxNCg0s3cb5Jxb0di
EQXjZzpvKkC6Pf/n5LvFxtaBsXNSZwR9o9KYyeAsDUaQutR5x2N4xBkYRIsgLowb
rBjcDJs9lLpUVNcG4KvWtVywspadj9fS+y4JCYL9MY+5KP4Y0fywIJzQCL2WrcQF
8WgJ8bBaKUB/q5x3VNl6eWJ3dyaFH5jIIDZnxcK/IlDvR48lSYJvoMaZt5v8tqNf
4J+Pk99KDDWU5Bfn0BIkBumMMX6E32S3H/kIrmiDOyDj9ISlyRiXi3eh83yhc1Lx
G7h/vrrtWKCyLwpSx5Z/Qb4mZbUoqW3nhlkI3vvjTvcKUgfXQ9oL+xM+C72aZB72
7364Jek/VrRJEL8p2P5jQMucVTmuIsvKUurKWb0NWm763MERK8UP1WDvoF5TMZ0I
85h5gU5NG7yqv6bYR3XEEryQVT6OR9JRSsz56BIcKHOFLFPZmzBgYra18e6/brjk
HXqtme/QzDWqhgVF7bzxCcMoSHdsHjFg2bsn2dPdNHV72dO7dGJmpBAVnajULWe9
2rQqDI4XBuZjqxdOphZJoqQ/KR7np1wPK7xWyaKjeC5tG3+EI9wLyHcfgrL+iCv8
DrocnJyzvbmbH7RMW/qtPtuQD8wlDQv8CtDqx0GUqGwk16z6tyFe7XpMuVfjiDCX
OBEY8UDrPOnVb5wH1eNVBK5Gw0gBbXmaCU+zk4O+Ao7Ag9DSpt6WWi3m12wt4Ehi
6+iFF3AGRZa8zHYYqfjmrrxrZPwo3cfyAfHs7q21iVgDmtNZlDIv2xmPbkZF2LYT
rIY11aDcBoOu6CC5uLJsUXOFYmTzlqD+ZLLBKxOChQFrmIut8rp6a1ksqh8w24gQ
25LLXpy1rmCyHXMmtQG7GiUwEZTHh5pxr2dOA3vCA3fhsskLFHyjFQodHVyRBTPf
F3T/+EanFbSh2o9OUDWjURipt3S21j5p7C/+6g0x6sFS4i8Et403blTtrt4tKcmn
1wI8nzOjYFdE2o1MpMhRhfpKAPZN2mBi/V/MTewVHD9tQqXZ2+OEvkYBx35O5blJ
oshQ8ETzM71OufY5BwnNyWe0NWdO2Sl6RMA7TegFOy2Dgqe3vGLLMVNOpTX81ST/
ADyuVnsK8MyWlfOlXV/6dp74dt9OJXctdAkBRGPrKR0t+lupm9reJdR+jyJTCi2K
Jl1mAPHVB44Y3LiLALLwGaTnvbecH8tPkEy8pM2kreAtXu6QMryasNDJsRctcrhm
RCsxmoBC992ul4kKlqy6/ZJCKGcwp5Fvl4RI8huChsaPetszPocoRRkWFaaDDmYm
pK/Y/EQrZ78iTda3FIi0FCurQIB1b8ymHYXKQZ8D1PEF2n0SZt1X0nDWt6sjB4IA
+1kNPZMLK/9V9u7oO4j/mZEjfe24ZhZwAb7LoZQReshm1QqbPsyTXIDnGPgAsQ7Y
+Bau+0kzV9fRrNey505vt4i3lHK1bpmzKJ3yzDAyv4ZFjHWibc/eRbQO8cV71rHX
0h1wJ3bXcctsH+mpJMp5iGwkSrhgPxteGiX1b0wzuyCrpZzVR6k0noE5Z71FQ6TO
XzO9dvxobvPQ5Ux9Rp1beDJsL9wOYORbzj/yf0Fa4hFw9OzWZ2wHclaNuiFD3Ln1
8u3B/4Pzos2seXACbx+wxLjsZgh4t2jt9VCULIurdBgITugjjMp/8QNOiJskokV2
fM6L0kXZhMVlmgqzS//gaeExVkyqFKLSNuLmI/lKaMkS9PvybPNlhwBN97I166fv
QxY3X/QEfsaqaoUMxv3MWXOpHb9msJlvY+BJxrlub3GlPpHOXZ0CCQzNbMEwMVOm
JDO4LuAr/hIaY7CUz1PkEy7HrbC+TjLyEQwCxp5XDKn0zBEMaeN7N1TrlZmhSL3f
Bz4vIJBeCHDvuLDGPA8UpqAYkM9v7iMkJUSndJ1ePM6GCOU1i/P+hE5hI2vjj69g
qr88dFjbj43ZkcsXzpbf5r0Lu7i7ULJB8JzezIX6hb4R0oX6IIFi+gd8oIQ5xEKB
+SP9BaqEqFrYLteclAgHI5YIPBjl+LHBAV9FeD/iXKFKtJh6LKMMOKVPETgxgXni
0FF0gFetrgwthlLakDyslDNEZp84PGdBLhf+0neHEjh9CbvYtaveSmHrAIBv+dPh
Q+eVeW3AWUiwbADFrAv8Mzo8yEobOLhJOLKCyjQxd5+XnoOEivjYtmlVtkFTrU8t
nZb8BzsyuIb1rrqqO9Ch/QRRs9zY4ZObIqfNVF1q1Il5VTn0mdAI9aToVQ33RDXw
Gon1SVGW4fcSeaCIlzny50S9VSZg870/yjmXJDxTm+PQganX6wTCEcoCxPcXIncN
DNbgJ4r6sC3AshN6vyRqHOVPd/SEzhebi9ycWWDxjCozc/qzMwt3Icu+LsqVjt3u
O6/mouXshJgkgNk9Nt7koWSkrukHp0yOATwROZIgGS+Ae0CWb58JDCSHTXAcZ7iN
XxYAf9VoZqU5Fv8rYkuuhydhsTsEIQ6HATunxyuZpATCZUzgBVZNVdpqRFGhqgH9
2so3gsU/v57KOkgd8W8KYx1/3ZIMfAeflSVNHB7pS9agThPaR+J8pgM1p3QezT50
OGFfDZXmp+b0SwPpuJuoAixhjRVk6M4Wsu0kKHnEAKj7/wuGpPuVSIrm4KYlIzNP
RRMBC7veiuh/rifiVGFj9hg9p31zOQKZOmvJLzB+zVOuZCKiJ6f61Sgo7ZN8KwLi
hcuFu6zhoH9WQa0STDdfpTT2NcztsI4zAw2NBoKc8z42LsVweZemvVGNJ2yWn286
CVNmuac14/iGBBgSIZaMAXHR8QeVsaJYWDAJawVadNEb5JDdlv9ko5HVblDND6zl
/GM3lVA9G5t1NJ3zdUtCzPpw5UskJ1Fhcpugg5j5L/LbXZoJ3X7WS8LQsGdVxmIv
saCudmqjQlFnQwC7kx4PVbWPOyqaHz6yQqP3muetR7cWf5wKLqA47d2V3vau4YFl
Ft+KaywhpB0OyecU6f+36hIIRVn5G1wHzywFz3DTcE7Li1oNRDUgCbdN7Y+uHUbt
JATL7OzLsgO5lODJsBnfQvKqL6990EFl8KRC3tlM3eL2ZO6ksI8+zr1YiolIZg/W
/irGQRlEpaq6pOb40vw/W/iCXamY+/kcte0Rmpip1Dryvoy2yxP/b/Qpi/FiyPxR
lr+ylpRJgbtqsPBeW9mkK0DbXdW596UtxZb/K+kxDZuMgTAuueK0H+ftJJEIWbTu
Wa9i4RqqB+9ZiCtmVtYwMyP9s8exWvbMPV5Y1HAlxVMovzdTnhF3/FXNyAvB1NA2
hKBFFChaimtEvhlOFRj8WNdl1CtwUHxB89eEBxwKm5A6e483I6AE8a0YZIiWDWp/
6UZnX3E0cQk+pIs+BuQ9mwS0vAuGCWbY8dAmClHHnSX/6GFhN/rcTFhRCUnPr38P
dJGgt0+0FvvJzPO2T2pOvzrkKfde2oHhfott3keblL3bLRxqvTJMV0pyaZ8E9jD+
vnc5jXYSQyCdSWoDNc/J0NyblUwi1c3R5L8eZU6BPnoFhTLqZt2nRBE3bpkiIx0h
796nj5kR/2W864En3a4ex69MHT2twYtNMYUY1Qsx8xv5kv0aLl7lXJV8GCfTAp6c
VYn8J7lob1cd/zv9O+GY8evfSmggVd1y9edF4ptudzk6GKihc7Hc39/aT+2k4Z0N
5uwHsR+ll6+W3M2UnJTyfGwassuXJ2DSgn5eeDooqd9s6SAWq1I9bocOM/hQhYx8
WcT8urlGLbazQ1fBfkMz6ZQjzX6G9SWEg5W+nKsharnHvMwUtIfaFUyUx7zPEA7L
JtdHhrWz1yJaBFNEpS1eR8X+B3t7qKoNVIA6E2X5Mnco83vx+f42pGpG0N1j4xq4
LCE2Sb+U4ORjY99/xC76cP2ge0tt0vjMTPBG21A5OjXMlramI7wP3CLP0eHaDqQ0
8Kj16Syr3B/HwAatboNw1FAUvc5FRzLrG1enUj+Pz1FWo170WlEifnYCGZCOMTg2
BUYnwF/XI9DpNvjVerQgRsmJqhe1vAhstVFak42ysxPj/cpO2KGsQoqWBnxZg382
DIJDKLfiTBp/3ddX4wkLfYmsDuBwGDTs1b35ZuvQ/xEfIpWqnUwjSvIFT8gwNjjz
/1SG21xGu2os2hlLAfOHZ/gkRxIHVA1P37zN4iHNNy+ZBIgQqwyf5ph3ZASfDLkI
4ayH9e3bwjf7A3Xkozlu4SKWwCvt7wYeZRBkjV74oqI7cT8Dek58POWQ7S3o9+sp
fyghjRH2WWGzj2AMd90liZqjF1K4HDiUYoc6zHxzmWF6z91qan8kakeb0V31yg1U
pbiCL4dUg19lFtPG0zXuuCcNIfI9w2ztMdqohEJreBkfeRkD3tEyn9LS0BCW5GlE
wjsmo6pMsZugNvx724RN2prTtU5YW0RAZSJEeDSt7TlRZXqNsDIywqupVMGUcEJ0
mTP7CGGPzCwGcS5ScPE+OxI3nwDuSfFdpf/YZJwEHGdX5KfTL9kNWATavLuROuxi
2cD9nocijMwAM3yJLYh6WVLyT37MHgVcooFfXMOBb3CoooOyKFe08oWNrHuquw2c
hSZTmjP3eWFgkv6FjEMXlEu4uX1Gwgx8/dobOD+zbkcL5btxVEVNTVivSL75V54T
8W36738OI7kOHqQoxO/6Y9EcNWRTqrN0I4VYZmJCJSGi5/F/YdevcHD2QC8ggB3v
MfF4qN38eoy8/Bs+8mwUjWs1dGb9zvTErCMUUG7tjGr8S58Lmg2+Q/Q7S3VXbgKg
94VygX1CAh00L2mfX5d6vBjip9NcwS7/e/5WXbtIZ1nIJfPv6cSuSrP9PUPWpot5
MG9RZtUVLxT1TfZ4ugwtagStisx9GbI2+R0FigkfysZLHkGJbCI8exWtKbQZw4mC
IpIIYW/dGYexBZXQhoxgiYgLnXkJ3gIb0L+G54RMwedUM6ZmCHMjzgyhBLPJs+TU
q7iO2wAD9HGgdF1/FC+4XMEElkQm8dLLI9ZvBbvj8ZuatFTl5G3U+5EBQSUWK/ir
47aZ4dFN6wlnXmiW64w+EShlHdf/0YzgJMqbd05qTZrD9J1wTbpDkqkit6OFA4eo
KfWeWhpMaao//A41HfbEZ2vAAI/E7f4/8lFxxv9M+vOx1dh8jrVN2Sm0tuPT+cN+
6qRUsyp56o/FJPVedv6obVDGYnOCjJjTjGLJOEc3fO4XvMfagnVuL436vh67G/aR
hXPRLSvHfkU4NmaPfYswJ3KtDBQVIXlSPBVnlHbHx6BQqdyDAV3eAJnIAEYDWoay
8qqdTY8acka36WOX3Ayo8BNr8aoM4IvTNtuH2BCjhwBes4UTbGVzWh4FGW3sqWQR
7Ly5mnJzJhvBH1Frtnc2tI0trvT3W3LP2HvQrRaH4RfQmwNRyDYZXI7RYV486Qig
IJ/sLxhshxebjwXzYNWaKVB8E6S0E6JmSQLMlzoW6HSSJMXVpbQJARAEZ61lOOi2
K+JhomiR9uDZlDy3crN5//72Vo+FLU7D+cJ0vIyTpwlPSoKXV1DVPzqzGLV9G+0k
0iEKdRYj4Ohf3MEUoP4zb6dGpp2+OJtRl4fc3DrqfuQOq+BVWyqjFZbPfJ0ii6e4
sDJF8SoQLDCruFSDJKCAw62azYBJNjZoA57KC6eBhJJRy8cw9XGvmN1hfW8pBnfN
NJssKUh6BlNI9sB/PfeKDuz26Bc2OL4tvjhOrcCjFUAdR2/DAFX+bceAhyVGTFED
uRdgQsi3sZstArYcK6DHuCtZUwISEzCl6a72DmKL6gHYbfE5+UiYQ+vhCqqRl8+k
n8NXk5zRsg7o+jcSamAe2VwKdWcQ/qFnQGTAMheuBiXZ9rj0Zu942/G0v8z0ogd3
2y2awU0NiUvM/+eR+MLLuYqblkCjiqlwstzuuU79vynmPKgm+Zx4fFKYXbrUMlzH
aKp/42FQde1iyyuVrm3TUjMj1EFpjw7oxIkZ+lqOk81cA9Tbkei2NX3Ij76br1ua
QEztqDDALMJOiUFgt0GiNzJZN5AXv4DfmhLuETiTRF8LSIG5JouXURVZsebzDo6V
mEyROS798dvyB3Iik0snV80qewxB43BbvXPd+kWw7aWtdLnB1GYssWT8TIm/wKWq
x0rB58QpFR25DJ/90h0mLw6KQNI52EFm7YsEAVxdbA+Ew+yPbVZCBSk20Fy8COYj
TRTxTL8OdQR5IKSSUMw3RBBUIATn2U3iDIcx3f8DxXahTuzYv+FAtatPTyt5IYdU
dUEXvrv8ItW7vb6rhQBExGjQlfU2AHkKUFcLQ1tX7YEui75yiEtX6JpRcKM6EheO
7KMTGGb+npe6NXwazM8dCZjqFgW66YoKet08oLFOt+hf1a52gJbkCRlYaRQMqj6q
6eJHx+KsrdNl9KBUbl8GGPhAzJatS2XbzgyzHBqIk/e5WkRg5DC8sZpOBMtILViv
4KVhwCojhIgYumyyKCChJueUXEFEGz1DyxAEeRYkPRCXMpLVqn287yxwbENhDRgO
KbSIUaNrTjc+VM+2/EvJJkufyFWXRw42iDpgaKvJdyAjG/KX+h+jNKYk1N1+lK4n
BQEVcstNBnl9cGmXgG5iFjc9za8Ncri/sLB/l674RVHsn2/cMv+95x3SCIN4ifU4
/q4eSK3LK+3feLgJdZ+2ur5SkevjlztLv2FvslB4CGCwfYX8JvCO3nMmU1MpIZdI
DNG1qI/XPX4toQZsGWr03jB5TIY1oR1DNS2lb5Rmp2AubejnGSNiBpDxocrVxEye
vUtB8cDbN8cs3PpDdVTnAgnFrdSEVBxbM3InPRXHNu0a8pis6qDoOK2gvXyOWRvd
IdpO2h9xku/zUGIwL0e97M+tFiJzo80c94vGYKGqgtCOTlqw0XL8J59VEh/H/IrW
hjS4R00j93GWy9J6zR5GgC0MyvmeTPoBIzYCAqkgRFdRlKXNGZ1ZE67rJtm6i8lW
hP+PR3j9D5cEW/UOudCALXB9wSuF2s8T7BSx0GjqxT8IqteY4IEF+29WcFPWnjCv
5IjPua250GQSgDGZv4OeX0UtH8C9droxQ0+0A6vzOnp1iWsioui6HSoAUu44p0WQ
oqKofP65RUPXHcGZKq7zcFvfJTXLaUKCKeUvZEhyy1RyPSBek1A2hRrciAjLLLfi
kKTNK4wH7WCGwwedjTRQ4dEu05KECYfKqHONc4rSFw08rIIc8l5eKirctPkphjUk
3oKhba+NJeVlxcCcjZyQBJlmJJ/3ww7LkFSu5mnrdGX2CO5jln5834MwrY4f4OrS
upkbuAvncDCGHr0iimOisEoSb12jA5qt0bJfQvSDiC7cakiqmrYRmjTcfw4OE26k
lb8TaPLHPa+j/TspVvF2/Vgo/JFjdNsbY1tOtQpAzJL3od1cajX9FEyJYnI/Sj/b
EKxHRSqW8rINZEhvy6+7KkqWgRlSLY3PCOFuyfj2fT4rmQlsv+DaxA7ze9gvq6dG
8eZ8xXz3malPgew6KuSiy93uf7q+pZ0Yt8hyHXvc1tI2tChC8o4JGzhVF6mGkKDW
Wr6X4ZeFVufZu4YTPFltyIJNmyHwcb1yOE3k6/r5tcnr/FgTXF6kCy19Z6XCmJ6f
xVRgoaLBoFpjgEBPEebYKaJD+8o/0dDTrAyJzwB1EOE1ShgwqH9s9AYw8gOsdwG+
1Uta2AyrIyJPtNU93URAUfL+nzO0mpoDT0B1cEklA3yxGy4e5ROOeJ3+HzHcOQQy
3KmJDn37hMQ5OO9qUxB72pWvv75smT5TlWF92WR7bvN1F7HEoGDBCGNrzyU/E4S/
jLrXevvji/argS0oq1xVzW65M6QrRnJX8ezybDH7L2ifbeOVKdtWE/9RTaurY/uN
zN7l1eynTss56qqIdySIqFosbDn5H8P9b4zkkQfaUznHbppHce6iP+Z3L6psyhrh
yx0Hw1KtIplcfv51iwnkL4NVF3A9QtaPI53Yuopt7KTqCn/ZhhbKhQXJTPEF/N/L
Cmkay/JPPgEpFLq1SzcdJEi+Zx7LhGLzkAd85/MMt74qjx6TTAJPHXqLaxTomHUo
rdEwTdnQ38BmEza/gKV8DT4m5gfupCWlxZrIp+Mx14RvLIJdsK77s1W2uOl8VMZj
4CZ6ssm1MRw2ufPyW4EC4LyxrKzNbNfHIzrPazKhE+Rmnr0h1p2o4Su5UWx7BWBb
pRaA+kCCbR9ZwUoKj713N/h4hE0QnBXRmFpw92eUuL6sGPYoZxH4U0yMc/LJdxde
aWwcmZayRWCaUnxFUYUdbui+W2jgFZYhl59wU2RLkcPbZVnxrZadvWMcmuh5wE4G
f9LHRY15EV6ieTbStB4sAwpSP28es5eDWaT3Lmxs+c1WssS4Qqqcz+Mi/CkcFIaZ
kbBRbtjPs6gvhbYWJRlgynJ5b0RSLJsx5uqrmbZP6GiS2dGSXAkFo82Qty9RWcM7
I1VAyg8A1oTfHxPTYcl6LZCesCy/EDsfI7M5DXETZcA0Jt7w1ZMHRqxoiK88s9rB
QmNj/xaTDqLvW9EDPS/sUdzdcqmC9z5YYnLtgdxv/L8jULPvh8N0mgolN+fc5v+7
z1wgsQOTlY5TkJTUKLGb4irttIQH/7nhnDAkIBoxp+7nNI4QFuWbuOAnSN+kkrTi
UGDA2jv/ykHGyoiuXj1WbJPUXEe+Ja+1naQNArve7xxRC+ZbtFsknLrgBYLbknwK
AIUTawdUikDxA/Y9n+s8XRM0wk4Bo9t/VCPi9nBHuAcgixAyd2I2yAx2VKBpXKJO
HuQJMnbLcaziYZzxIT3pA5M4H8LQZCaRY2eD9ND/rCa3jSuVHfwrmHQQjvMRZHYT
mNYJT0KC+1uTimS2vGKeGdEdyakWFzH1icC/4qKsmzyyr8PNbYEM9nD/D46VJS2s
XvZ3Mg5KvXUbuQ0ZttEnDtshbhj4akWIk+d+ZD3eXtd0qv/5xCW5uBlT+Hsmwsqs
B5m3t7etP+YYD9nyqEQ1AqhMYAwqjxB6yrOT5n3NJUYeYDLvSJ2/0jlwifiPl92N
LVNLQBrh66tUSP3qFwhuOC+nYYcgt4SKOAsybUanTorJzMCh9xB/URCci2db1hOz
XNjtJbau+6YJzEfU5KKQCyg5rpG8Bm4Qb7Dl/gsGgiQ+4MZAQzYi8YQA7VvQHkB+
2Mj2dCWEcgMugwSQJHhbgO5I21DLMnnwyJ1yZMLH26vU/RM0OZNsiC/Wv1lW4qFd
87U+d+Tg30B0aLgOqXG6dvnlO53vt5LtsyRr0+WD4OSkEVQACzupOls4XNp9u9Ml
fLtDJlFPvzIyt/aC+qkMj3asqkSrNQUCAfOHf9e6yuYxLDz86LWZ7BwtdJPXJzhj
iyCUbssFSy7Kc8Psy18kIS66wGr8U8/E8kyKZI9mgZkKAfehtGAIiYULLCmPKpyh
NevZ0z9hT8jHGGS3pbFJYoMSsbKLFze6xvMLlo88NpTkCAH35FTqZqY4XmoykwA5
1/RQCoqasYIig6M8/qb9avMGjLf4uCxqtkthc1NGwYRz7ljTxzR79cS98NtiJ51X
6E3piYxytxRlvovJJFRNBpVP8XWyenq2W0WE3biSgj8g3SiUqENtBj1/0Kw6ZiLg
EvOWsE/CZG9XKlT5TCBDHVlAngXEZepo9ClTtLBwItCDNhgAk0ObJ1HNxVMLpP6U
57z+mRqcNSGuOZwfqBfXoNdHONgNoggN6T7iK2dk92gwGHqjdRMSDjVy84BaDQc9
ecHarE0wYVuuxy8knNG78qXWMZvx+xe08LyZ7hWF9txr8neAadoGg9WTuOfNwRrS
k6NikzNAw63KnUuDnZuVNzgEzLFpgd1dbdvva/S9AdVVYhphRHzHcZl1+zMzIpdZ
vMxNwrBQ8FKYDbAuz2JKo97zuVFs26Otji1VcAdZWavcu8/0hdtVWjzPU7sq2GL9
Z3AhXVk2ECHAiaboEQVxGvpEsVjesM3Z61Q84MSoQSUkDq7z7Ed9FtjZ9E8jwcGh
NlaiepaGi3UwtnUvZGbhLV7K9D+3x6QJapkBgeXNugezowGYFAgFgSTzoQCrlKed
hUnali4dEBhTqGKFFnI6bWKhoQ90IHZZW8fsBEps/SGQF6gINEdIEVpB18JyqF65
kCdRYzpWve0TtQ+OsXRk182M0bPjWQmCMTNcjA6rKbiBtTADpmrMkHn+ErcKEGa7
OwXmmh6aV4SiXeIvSEWKLoqXQSFKCcdmim+e0kZo4RR/lHTJqmawZcAWihrP5P6S
4jmD84hM4FdAx+y+fRZ282KE0O1qvcl5IRqmDFGWcvSDaUeX5Ogo4EYX6+Q9G3CB
IQ0YFSd3CNigLU47r+u8XiGKpRidbLYe3o+EBspxY2DGx5UOwhVSOfrMt+qWj2mf
vkdJku2iF3AtZaeW7YG6cA1YpXsRPJUS7r4dlbVxa8MBBdbHAcdg/B3G8tgS19uT
tUKpjhMkDaflomd/CpD7HtIGM3nBJ6IUJeuqL7Fchv9dTOetNDGKHVVw0YN/Xlc0
/DVW4PvtCSkDawfIt8v7uJwkfW1XilsCZ4TECH11XxYJYhZCR1YvIhnlq3XnIApK
OhrJ8br4wVc8mcltVo7VZgTqgVGO9t39BgAoSQJ1hpgKnfVL+nUsuadUAfP98K8D
z1jOt2atJBtiiobjgFpfvVQASaozJ5T5feIuaMHoVvKl3HTHHaJf6pgHLjgsqKi3
4ZDuM/LzYP0YpC7OiT/ZC5rJ6vohLKcCiAUwJDJCmUlI4lTlhtMG1KxshcHg2NPV
s3wq1JNXKddDtIIFRqxLEtIs+mNGzFU/R94dOWplHvudCrgDEzdNzrOJOBMZtz01
LuTBknybJMEE1ZOQVN+geCs84QcpPDhWhIago6iDnSDx0G427xZNK+3A5Y9+dg66
g6BTA3DBaud70udEse7fjGmckB7CkuPJpwXQerdbT4BAla/6Y27V3zEOfQUgc9Ti
f6RSa0KuCqAzrI3J9VMabRXjt89KFs1aRdj4yi1cqh1cAat3CON2+iL1k6xwVJTZ
m6sGhzpl0gk682adbkJn9vq27g+NdXDXDAW0hHA2lhhaDRHCuH5wzqxtzdebnnEB
RunajhQTOL2D+EmJeHXJ/ExMhX3s3rBXSyxxMHNP54OXyJoclSv3sZcePcuRPkiq
JqDqb+hLQh8evsh7n/RGb4kr49GoqkhqcfhZYQuNE9MyN2ZIYHcxXuF6TWVRXj8I
4abL8U1Rkd3zdNzuuGe4MbWbmSHKSt1oRmvCuV1SVNQEEi/KLlClZ9VTWUiTjd/J
o4ltgAur0g8qVqg6wvB7mZxyLfHBRsaIuoH39YRXPATojCb2jMNtJ8yEaZoHe5YR
DTI0e/WMAWb8BE5PfuT2JcfDwVUdrCwJCBXpU+V7gpVVTVeXBqYS+QLa/ZuxvzMf
4tHsKtTX6Ct4jHdWTErCu/im1Eb09parZuUxRAt1Bc8LQw715kki8EZrfYJ8sOIh
AFVrEBvwR+0+ex8KRbgzJmyywbeHkw/BsGEGQGZZB93OkxIBnkoBMPmo4Wycn3bd
9ID6t3hKjCXugUj51nEAFBAJFwI8N1jDkXJZS0RXSa5lyS+lr6Q40xIAR+hPSEMs
LAL8pjTLv8J0CRlSx4+5AflYlJUe/TjgkoV2BjAmLS1rXrKKk0VZE+emiUupyPE7
2u7mTyHH+tAqdqV4+5umyYmqk0XSReuRNdArFGDHIQ3cAel0vwnFO78JDpFpXZ5o
qwL9vDjGxyGCDUseVNsA6yrjActXru8arlpIvl5HgFCe9z8OgRV5N2gLLlEU1MLC
frFOhwjgUBYVm4HURs2TGcTwYEG2RvXKH4fwr51R/4q+YwwaAmPaBmnk6nhwjxMD
8W5UPSuObVTFzK3xvjO0CP12JQAXNhRo1XIeoxyPXGWhjHVcNTpJ3rxSVajf6l6T
oeeyFctMny7FiET26EdYNqem8UZ2z43LGDJrc3PoKj6x4mROX8hRDXb9AOp7i2Up
BqB7G0gW8ugvDFGlXCdEErq/yA7JGN3HDcCn8YQtJmjsFY/ZB1lJbCSTGSO0JbJ1
yHMvOlu/gRxPyDYZ/bNU1/m3p5K4kUXc9Jyx0HBQktsOml2V3Wnk1ViSJGgVrqw1
o7s7gwOtoxwpfVv0ZNkLidyUhMLYZ6qpdP4pNxe9V2USazwWEYo1pwILmYVIiert
MkZlsln+WTbmTHx2yG6+2M1EvSFNvdlK9QKblVQ5ZT0JX3KinUmi8xhlC5mR0eoF
tUzjLWqNKx6I/LNARF1aAIJC1n1l5JhV+m30s2LfAX5KtbOP5INBVO/DOjcP8ORb
ak5BSFANeFDRvjlueuyPoE3MI9F79Mbsjq8xbBUIo5SrKHTRVud/EpB7lmcSh2c6
wEagNjLvuo7KsPsKTSXl1krhWCpkuFJ052iGpz/xo2wYLF7X3RGtrDseR9T+kTVF
cBUGrXdcvO2Wg6lF+rkkcLWM2FohJcOo6iDt7a3J2WllJiheHlcXvQGaQVIO/cLr
DXwS48XuLfYD9yzKvW91lUAbw68vGTWr043t3v13M8LrjlZy25N8Qsp1VmAsl7lG
HdYWZgfMJ1Oif76HRDYNQl/8x0Wud60FAbw6bK/UxIprC7W2HgjDuinwdWMPQmP9
tCXJhv6GW+GEUPfV66LVfTNPMuzrHYxog8WXTKgCo5XSjbVug835IdZcrXHozMdS
jY9qkjCFspCf2GJMSz2essADozyE+gOqDb32qLI+YsFh+9igYh0sbTX/BnjWWi9z
puYFNHaArwdULmsdrj1jKcvyBBaGFxpJkHghdOu+QU392in5S0Eci7gb8N+pWNdP
ButyvF3M8jk4V84MqU2wH5aXgfDvnDDRr9DeVVBY4CKWCB/nVBzp3DiqV8AO4tB9
gkPe05AKwFO6tUzVxPY6u0GxVzCdEiweAn5AcEB54qyHi7xwmreiyVgLDtCHjELi
/XS7V56/svqHnq3rHoO9geIdnEzwkJWj71qqA6S07iMPeqtoHSTkMxi6OHJYlLVj
PwYvxFtgCr8WheIlFl6CjxtRRvLsCe0EfGC9obHcFod8laRcLqpZL30KBLYJIMt0
LLXcWtzmDK4dYGx62nNGu5mPj/3zrOSeCne/uu7v+bgl40IHxaBFmADYBG+Y4iiY
yLHzQF1VwElg16A7hZktK6jTZnDL3lXYmiyPHElxfoqPSHZ8W7kVZgK0T8jKyp6d
BfpW3cd0Ont/00Waju9MCXuAW4wNIDlAPWb4qTqIvjwGHX/znWF0tpjz97F7SuZD
vvHFfRFlu0EqzJEEIyCOBDaCtFhKXSyp++921Mttoxwc6SPBG89zKuFNzQK7ePUg
356Ja5SNoFzGa+Tfe3YVxW92njU/9afVEyxK8hJOYQjeQ37dl0DOcHhjpMlA4koe
LwubMDL3KZsX8+68HliCksgMCXtWrNbupWVKsD4ELZ+StmQuP+UxIekvscJ6I86z
clBQJsf+WzW+Cnpdo1XRSG+uR3umIegdvRjqAEq0ISkc+94ZcYQXdF6siEA35Xtl
KCVj0c57mLMYJhrlwtyC84bMF+vIay1nWK8lOTCejezIY1SyC1sNSjcbj8laMrNQ
ZgFLyv+iHykhykwQnPeDBkRixIV/KvSLTsigi6SlA0zD3l+KejhHEvGP8H76CqoK
yZfXVCav8FRRJFlpWKWtvXGGtc6y+WqB+kBnN+BjdFTn2YHivhx6sBCsiLV2tyQD
e3luDMgkMhK5oW8AIEeNpunMTD+pwqz/i/773R3qsZHugVzExAvQ5Yhp5DQpchJB
9ZVFobW6Qo64AfoFMpwoUv/WKIXSlWFwNdr7cY0IO3g/sZjaG1fihyn+llaSLYCW
UfZ+6sBIt0mJofKV/DI/p/tMyaMld+nwzUXzaXIkqw7hD9rhQiQSW3AkIQjBtjOF
yMXB0JSe1WC4lR8BkvgnnfJ9hCSZOvVRfexOXbw5EyvZyCpKziJKtOykaesf7rKA
zrPsZqR96hIfIoMefc5ApxGWatppYSjFIzFrrEIiVStkJVNjT0nwfWIQXfgwDMEH
80qKQb9xJKVnx1KWN9nOW9fEX8PyxDJ2XvCy/+96sKJX8lfMsY2oRZfYuQMU8PZD
n0ccnFZ+zDbM8Aiv0Xau1TiZ5AhkxwMVYEt3Qcnn7G9iM1HFY8PkVEz7k4p2LDpB
TIFUTWNI6SwiswhAw0lq2knA37WqaBISZ09dH3/4MJh+zBI08MLqgefNhJ9GeK/v
Co43stRrPYHEM2Wcp2YnwxjF2kp++glp4fDLySrcYv1nFqymCYDcdO1wzbSGiIQV
Y6mV4fe7b6bCKgLHyAAK8JS7QcCCVQbOgcnv4HySVx7OVI9PwMHQwUIncYt18KgW
4l7scfRBq4CS7OvYKb9zb6I31w7cloCdPTXhhKEtwRIiG++VAWy0INfDsOTf8Mru
uMY3okK/+R6635futwkhpS3qGlbYjZpWIb8PSIGcXOW25ciwdd5a5tuOOxwgrfPH
HB8TKTFVpXEtMnVyOufLqJGR+dwvX0NHH/T+BL07VPTFOg7udCYwX2xHGMk90FJ3
NG2avevBWpx/Rzw/DP3qLC3VAcXwMetM+3g6L3GTJG2++fwCBuGX4CtD/62ymvWw
jFSHvMSup4jv77IWYvaEaZjh9NDjQSzsGSQ79Gp5jf5tQc8bzLim4zXfCHZMhXd9
3Ui4j415o15QLoFloRklh4kvgB1UZBv3UdDq8yuTNmdkSm+PVPW0bHOhrqTurbZG
V2WNJr/QV9jtF9mhQDW6fz82gKva82/YjuPqFLZwn6fz39tZEC4zIYI7MEIk0K5c
o4VZI0dgRWw52zs7MPySDtPq+SfFx4tAZPMOxBMwRVvMelgg5gbLMX/6EyB2ypag
C38h6JA8iQxQHfo33iZ+iKgoZrG3N4wAb0FQqizvjxEvB0HR1T0Lqj1DwEDZeJZ1
PbIydvKa2kQIiIlXwv1zkZJGZXSFVF02YezuYJakY+oFy+7ZW4hGs9kyzBf/5/Zs
yXX3rBDIiw71n+q5wBQJmZkUp/yP720bJ1LCLXtFc6mvs119ybRB96NJs0Jc3BWh
VbEM2eVyAARxswaF4mP4YW1FXck90g1fVAzeePlRec1l8DCD+L1DbATYezvDkzR6
zb9LVb7zCZMgx7EGyiEHmtrviWBi6EqtNP9jA8/SzGuTA2541+PX2ij+nxXEd76M
pbQ+bT9hl+eZ5/ETPdlm7ihmrTrHCgQVipALqFnoR+ggPSV8i81/RcFYKHAmak5m
/GPNzxaS5r1qgWKAZGDwMbTSastxkdhqMYCXxu1MghdVferClGVLRGt18KgSiFcQ
qAeGZ7pwBu1qTVkNmgsDNeC3WhS+AgDhn9Uyijm5gLylcAq22SQYUDMXnDR99OmR
rLJNMjOsACDwO8VRD/udVZDTjFSl9C81/V69IVjTie8wl4abOqaTzVQBTUiL09SR
BEowiGGJC97bZoht4B3IsTvXXC67DQBK+5M2DqD4Lox+y/bEYXf1UZw9duHd0qKK
7yJIL0mECcjjX3cISUgAAgw7555+1eRQHuqFYjiH7MoL5xTFh+Vcg1zBm+K/k0Qq
YsYAE/YComeakB2sfGSdwe+iBRhL3ePsYbcpan6GKNX2miMnisqt7w/SYLxBrtly
eI7F6Av3GbNHbGMGd/fVkS/lnuhp+hznRcmgPn+gTfGzy9+JUS2sokDw8QXwMkEO
30Ph6tLlVxlPSWb3R4Nz0jrglxUn+L84ZEqutOL83t7ON/Wea2NteSGs4MynaBQj
iSIO61uw0ylbK7uQyPfyJgJ2OGyVhdbVn/Cl7x//QY1NWBqEgMZXjnxokaPbBe8C
W29jNi3I+4E4bAn9lzST+AOPDueYN3yXE3ry+k3sCt+ExKiWDlMCd8pJvFulm4R3
8Gh6Pk5uhrea6qD75QcQIwWiSxtDrQU9NWnoc6J8g/OK+ME8OUk/jPvYoaVeVveN
W4ztxL/qgzN/uvLcJOP3TLyeEQqcjhJexaBmJ5c7MSBgn778Elcw06HEW02on54t
m4Fzeh9c0GxUsyxy9UeqMNd/mjzZ5z7kUmJn2lBZQwME6A5PRbPct9NBmkYFKizW
6wxiSSG6FAuFn3uuJtvKaVmRMOrtQb7D8MtzWUG+rkgGs4GbLqRk1iCzz6KbH4yX
w/SkH162E695AHpwO1zGthHFyMadzAGHaJq+d5Wnpxz6igWVculjTcEkIyc40gde
BxNfqHu3XDHswdcdDbIARt2nGQ4l924t8p9gs4xWhw4Yx4p1qav6AP4xvtV7xyEQ
2/0WiQVsVBNj4csh99a0zrRcVi+8Gqw4Vdu3X3G6YGyUqB5Yu/DXvqsB9z6ujj7h
T0iFDhKr+RgL9pDLnL4xp5moIdC+0s2btjJMaCc2nCaIM9cIMsDjrifaJfcxGkii
KdvUi8vp4fsdnu3k9e5K0X0ArS2AsEIzpJhWFYORI/eKVCQcq434vm6KxMUrPdfV
gjReuOevENZbZTZMM39V7bSrw380DJUVsxhYYTxPKpSQcSN6FuxUgfLgKYCmoAB9
zakevVjf3mIib7jzrpZgb0a2V6/2ILX+vvO4IyCHEVBkOVuaZV7x3EzoaPjrJcQm
SqgBcoSoqLYdMLRGfDKkmJ8OsIII6ynTyJCQ/wuVd4qzwm4ZP8NSUpubfWX2Jh/A
Hy8QcTZeskBCD43i7nnsKgQBg//BKq0oWoZzoxsaCi4XH1MpAx7UwJaMM0X5W3pr
WShfbc3LkKKbhdCJg7PxZ8X3o8OAwRnzPLdPjrDKEGBgoOoSzK7NxMc+iA6Vl36W
3btFx4v1NwrU/LGiu6Eel/aaLGe3WHuoZrMF7BIhdpoKSY7QBtbc5mQMXQ0T4AhI
IP+oP1Xe36ym6PM0gkooMjl/RTMpR5i7PFNRIOS4emYhnnh+NRoz1pNlM5hqy62W
CnIUjaf5z9QGloytfgd4mWSMPjorkV6VlGWFpx/I8+8V7arucSc38CO0jXdG3Wtj
a2HeH2Fsn7yM5UQF9S/SbsZFc9/y9I7MvOspWYygoVWLTSrtzn3Ax84MS80y+U5f
uuRcCGegQI1unAAYdK2BxRAQeoMePs7UUiHxmI4gqxe6CFcBx21N+siE3+TOL/PD
ZNsYv9Ezq5OaY5FdW9JFMYQbp03Uy2kBVe5b/hemq3hpOF1JlD8PLE/VBhn7pxvt
hQyBfPM2RTkt2QiJwBqRzgBk6+TORe5QQAU+BQccJD/Wgo+C+IVLy4xfQnCUUCNA
XQCLAZlC5oyLsyEkAu73LbTXIMvi4P6Z7N5MzYJabPPsxqsGleO1LHIt1CK4desY
fpOaBy9o7nFJq5tqeaXU/bQ3NSEZLPr8VCcizwPxSKAcfPiN/YXZZqSIh9vDOIxh
DDiH4voX8j6HugkqmTLHoPxHmFbpfKIuZgEaRpKDUr4ylKm8qR+Csu7WgIUJNr13
NhHZaxSlDigm2cuthnCESxDm3xED1jFmAAYn96OOYzhpzP8k0ViWdmh0iEXg9UlC
6zapihO3VGMI9lDt/t5hNYIDcNekZZKvHJg3ruzOL7AlC4Zq0GouMi4P391hK2s9
3AV4tME3C4LyuGc8BKSi7x9CwGG53hL8OSUlLYbBTLIgxVmm8tCnX5zRCgeNDXja
83H7VUIZlx6C3vpfrGmwjUV/w1zg30y33muVgcgQcLlEFDMG2Cunyl9lyXDKyNtJ
A2L3ZFbXyzs/suyQwedaBi8A2qxM6tF6iLEXv33hTmDMHhJqcjuM+wau4+m1p4QJ
3enrH74rnIFcD51p+2PAKMzHdfFhui6pBMVNK3nXLbP/TlHV9I1NeclEtqMC5GdU
1KGs4GZc2S2DoRGdqxVLjWcGZYv4LyA9l+tpBeQI47ANpjOk26WSgT2KpekviQUE
xZnun0Yav4pKS8wRnceZCwXkZqxTU6TFXDVlY1of4Kns4ZEsMggWLHbS1AwjFi/K
6isgtHb+mYnkhikJrfW0UGfNpr2idW2IbS8VRyW/pKTTXnUkU4dXG77fFH8L5p4Q
4W3Z7Xjq5hsE3+4JYYJO1H00rLaVM4kyulb+IoP4spxZJeWSwAmOtXuWxrJaGzcF
/hff1bPGJ5VJ/VN+G0+i3547/afY7XojuzFfq08FtLc1SJr5gQ5a+N6Umth4bMLy
fyJCTpdSvNObepNdcctyODLLFASmjCvA+3c6lgHmn+eIK/0DtT3B8AN/PvMv9Yx8
hol3Mc0cDVboruAJvuuU6oS26qgfKmkqfDgpYYqKVKZBy56eAAzX/923o7nxZtbX
TdBv7gvomv7sdBhUUxuustrWjnpY4FBUFZBv9VWc2DDV0QQEh1tfZ0Banplfe26O
4rzf99RFjaxJuGFlOQIHmPToPKzBK8vZvYilWtiLti7Of17wKNCcPfgbnbsBLFXL
2xC8hV33mndFziyM5Xw2TZOsemOFIk53h7UWZjBw7KJw7+LyqLC3FGFO8O61Wv6M
FbiGhTPyV5s5XWtBCOLFq1bxmqdsOOWWR/NRXzDoNhy+ZqAw1Pe8tezbvMiR3/MO
7w0lbnat34ZIIPPjAQJSYnxO0FF8gzIT4mWiBueyW5l+NRAipumdmNi3H6Rf2p+Q
ot5Ymccf0px7JznCM6ysEBVon/fdWevumPuSXfd5qSLfisWY6Tk6fjna08oUmrTk
xyUaV0jlFqMxvTcOXLBYiLd6EZzNvgQzdxZGGImqIR9gSW/FEC4wqua59TT4E2rZ
Wz0UWgTSrmDoVOcUKahCcVBlFBEf7DPcws5AyVOhm3D58Z4fK9HiNCZybI+iGNtD
wHVYdmXgxxKOUShgrMZSzFC0Pf3OCwPPFjVRGUQ8PSfi1jyFME8/jmj0nBj8CdwM
rNH1LGw3+TvWh5UhxLAUpD3u1BHjlbKceXfvCoEBNkra/N/qcOgGG4oIOzIQlqeK
EbTOHa1SCPMJOrC7bv1D69sWKM33lLc9nLLw4cqiJifyhnyQ6cHXAZS9ssdhZKJG
1G91euKmcTNDDvtmZakzaNJygMPEDjTBNATUdxB8HDAFXvVhrv5WUSdRDReEhSBi
wSr6e9AA9QbGmHoa06j7zzcVykKNS2VHAatHH3y+m8qrPPqLGe3G7ECNQ7PSvQ9l
jNcpP32seyp2Nfl/7AsdHLMJDuTVrTxxgXANfxXb94A4Eb9bydTKsvAxNSffDIjx
FZt81vnrkMdPrPTACfZukvIY7CGb2Xi2SOrGWjTU/ognY18SICEMVIqeC6fYPvyU
XQ9rHjcpIWUGh9hw3SCT+NcxtaHzQ5FomiG4E/iMfVGOUHm7y0ENzbY/WiOy6u/X
jUBGe/xCGwnkwDTRK+Q9jsT5UUKWIaVOUhHQISCDGvDZcZFdQHPFOEdP6adFkt7n
rfLMUTcNmm+seF4++50BmGGEBWo7b2X0+PUQqpOb3q8bkXbU/zYYSUuU2N3kF5zM
ld6+Cj8NnO/24V7cIjfjlLV/O74TinYTsJBtSJpGzdzKUd2BIBVWO+V0oEnR/Feh
0a+O1ZaRCC6peavPfmUzrkMIf2JQB4n6aK0pHhRnGSjMIXYKT2Znyvk6s4XPvmvj
hM0K2vONKaY5O9TZphtvNTLmL9gdIpZNhtgCnpDGvYtPyFb3QS7LK44DPSMSIrRh
VtsSIBS+OMKJFyqfku7M6WUnSuHfV/46XIMQpFevJr5XCLfyx7IqQYZdkBH+Ijt5
vkUNE2/RFZoww4TSJjxrdElkrc89tX4QvIXhnrl8/nQlVY4iF9cNtV7gaI/dg2I8
XSoOfty3Pwk1Q6a5SjWZUD0ieK2ChTu+O4z+ED93ttW/MDuP8gkuZLlqVHCDtq0X
SUNznOw3CYdn7A5V95X3zT5mD1uUJh9mfjUO5eh5MTRlVbYL1ij7K5zpA6OAa9FB
1Xe9vPKFh7T1rs2On1v6jBjrcWcSGhhqcI4GwNjl60Jg6xOENX8iRZ8C9fPQw9+w
rInU+M9sC0SCRPO+A9FO1V+pvzJLmzkaQHinwXEgT+WpsMBgrbQr9d2YU1cc+wRQ
HaaeYCThu0nNG+rEZvps9i0LIfKiNyIncAxXjMtTOawqk5LJn7DR/bEl6dqlWfzl
ClLvyPczZG+ZaYrVZ/D2Sxlz6x2BgYIJpH6TtLoOa2g+YsfkZCv4xxXBUSH2x4cE
LcycXJNBJBuQq8NAiRXsGRHI3k8e7UQ8CxBV5MJ38EUF0Q5MlO+qXdsSPBgn6PZA
LBN3EW4rDLFV2SQS0EaWd9nFdEPbc9cIqvhmvcE4D6wl47n4tUjxlHpp+LeN+F3X
HG2/71GVK6SQyeL6OO8UU+t72Hhi2fnCHOZDmw+8rL0d1ffwDllHJF1E4S3ksW81
HPfpFWcukYA2YBwSIdXrLF9VJKMHVsXzmtYQH8CWBekY1qWHkQu5vRh2Ne6c1XDD
9T/HG+id+KAEWRA0QhU6mp8d5gGxSaq2ZviwRjakmZ4M2NSg6msx63iRrudxgtFx
6XGeJFWxbJb83W0KyrXrxyvf+htrVJE191Aadtp2dcjRKaNEo8z6CyLXxaBHXVlD
wUDgyEteIb9zC3oK9axGRmzebfnw55XpyAdfon+JpmsK+869qsxqvCEcstQI589n
kg7pXExskMbVRGpgPjBK/IABg6jdXhPCB70siK1Lu9ppi3HiQy+7ENfpjZrHWxRx
OIGQ2KBzjLrKlji2GvQp0wIMTLuoDOXDBOCljM7ZneB8Ee4pd+0cRC/KNDykFrcG
3xxDhVouiJRU8bP//SSCa52aPXiv9TSUGl/Wrjm0giL5asQ2Ld15/zF6DEG91p34
IeKQqIu2/d99pP6WP6G/ZB/aWUnnDruh15CfflmBkf6PRvU5xxZeZABt8At18hSv
TPfr5YIkH53skgbU09hSr91jV0aTrkQCkTlHpIwOak9HYmzRtvwI7xVGP9gF3PaL
/fOZsvoVSctw+OIKvzk+mZD0Q5znBolAGsQtzpqaWN+rUpfWXE7e5JVy6X4VVsMH
MeA1nDFzp6s2w+YCbTfvwCZotbAmro9Zl4G79BcqewE8CwtGAqS//6pVQj0zflYx
CMHUENEgZ2hwvSCMlEv1/1xOWD95wkCdD8u/MGcwQFDZrU2nxOn8R2C+gPWzsxAn
+yLMjovhs4iyVkvBSvdO3hXGzlxJcdpt/UkH4tDw6DpIGcEgsRHBOqc5W+q2s8Y5
GGrd0nTvK2ocGOF4mzHiZhnmnD2TWyaU8Hb5E3nWJgpO0O7OckOZXCG5bxrQ2giB
e1BUAtmFRYIu3ohbo+QH0MT8yIUugQr0qj0DctTSLv6Ngv6fW+gbv9SDGjPzxzva
F1Dwb6SCExNBreicrAKBxipmQwDEs2sWq4JrDXzCq4EI+yCPBaBcwm0Yfz9UQqhS
xDZcUyXxGC7SIeSk5Sgf9iK+bzA2lpne4c6O8xrkwHZVWq65btGG2IO15YIVIv80
xizIMFCPVuIah8R9X0ypeGY9KKDBfgTRBYjP6yyMgReR3NtMHAs83ErA4gJdPsXj
ZijVwnYI8/i08UWQZHAG1llsSQEN5somoMTDGJ/qXe9S7CoCBF8r4F/ifVDzE+q1
eZekHiWtHdMnXtJrmcv6NwSTpaAaqM8vyBnJ+Y3EtgluwsFxSli46OmFNdKIjNaU
TcL682fuvYIslsha0u+tRx8OiAbhqwHn3SBfvecCPyEDcaxD/x1momEgQqGJOud+
VCsZudaTT9ugzE3pxcHGRxH3jwarjN4CeafED4hGp6kjyKwFuipdTujFbiBY4pDq
70mB8YCX20K0UHrE5wTBaXIH9GFGILrhiEcsqXDovWfEOsEKB0ZtJDn5/LLqeC4s
cqcu0WV4FDMhRW65jKNbDvj8L2FKpBeFWA10+EgDfr7pNrLYrqznc4l9oylzm2oO
xfxkEmV7MvUgjvFd1/xd4oZ1VHA4L9zHo0ud6lQVusI88vOS1UeWOaC+lumMxCum
htaLPPghsXrsepWQTIHqMmaNHpwU7birMn1Jw6Z1QaqA9FNxNMfGU4/6LJiQrPRy
MBlWdIAqmCkrqqjM27zGGggRgm8aQh2IYeSiXekhfrAJf0NchYz0POhJnQEojUuq
8qN8maDKAWi8WaEX+ee8ir2pJY7SbARrgTnsNbVLjjXLIWW9JG9/eU5HS1ldxGKG
ERPttGdxYppYrWPWwMQbwROUJWjdYHqWnWhEumIQoTURoig6UYHijkBelVviz+AK
gvDEqjSBJC0KoCRkwTaXDGDBC6wn32pDwv26kJ2+dF1TWB+DLUFCBOjJ/DUin+9Q
6TzZvC7CXwakdqjerYjyaUX200ag6KVrLYPAcz0Xgwt9YXB/vAlnLGWc2RuQ0Ukx
YS/p8Q0n0XGyixOd+CSm7xlCUqIj4YkYHvlLTCkuf3JOR8DU/QBspO2dxUtYioLZ
jWu5SzW6XBqxVjXiXepIJBRhnHueHiXmTfkLevnBFGeMxS9BAtESWK+LpykZKQ9I
/CvJo8r4GMJOIjfH6Q80LWT3/0XVZmDgDDFqpd20WxjxNOkTWUAXBSZNn3RPBkJp
tvbKYltbW7s+xAjI1e3H2NOMcs2zpkdO7lhRXZoDLz6ZnPvOd7yzqG0IdLUtnAgp
Cb9qiY/TH7obFj3rdM/Wi3bCAmkrk1pgm2Nbud3bYf+LRMapvUfbp+j3sctEsuAG
agh1pvZaXXOTBmhaTO4HZPiv3ae5ZQBcfo1DlhD+IGPXhUBTgHFTXxoKakvnUtJ1
ShW+mL4+OjaZwkeJPl5Uk5yeEMs8v9rN9QFoVk11ojQwpuoJ8WqJMUuPf1CvkoOC
7Ov4h5ppqV/QpJV9IIhitb6Usvvu3pa/6iq9bqYBoJ/X8aQYG2uVwr2Df6ONWUUy
jQdPyAA/01stQWlvQOmTEOkh7BrXt9eC20ERbD9zs7E1i3aUwW+5YCjs0NUY5I3h
b0GA3758R+8EcqQuWx9SFRweEtC21BBLUWVIRPNW7J8awrCDZNLAgqKxGx8Y2QYf
kiOWWa0rdXAgs6+0l0ED6AEMyQeIB6gmIIiydM4FCHyLuj0YPZddZhmEz3LzDVxz
RbbbYudK76pDI23VYK6ffMlRGW8s/QsJND7c2r7qFXzS2TdXIbXiIkss/EjQLHCY
sagz4SYYc2cYiVfb9YLlv60auPBSzUMW2InzACy/Qa4jyr5cZUuGVSFLvL35vanX
iWZqdZxWF5Fv1Gc8gglpYes2E27DdHLhMpA7CXAfsBWJYZLXcNwrhgTygr+L4GnA
vIcgfuOrIUug0OdkhWariBJlGHE/MdTBqUku+ZSwvvKYRe02RTftqs2ERRd7i94m
h3zuDi+zXZMsR1gruzfNJwiYp/ZKNr02HTotTKiU48AuV0Vlzf9iN2iyok7VAzE2
YaGc10iTSeWM/KFc6PqyDLeuAu0g/bnQOaCdr1a6bfeagVdxX/2gDYysYDDFXyjx
ExmYi6XgWg11KgzkviaSyLMnvLl5esSoOUeAl0lzP1c0h4w7NQRpxgPT6l7bSMfQ
1JLpuBqZqcmo6DDjKsPqw7qIXPcnuRwa3JfBm6HbXv92pBwFjcvUw04+ilN4AbID
5IyICOA59aqli70ryDFn8q5vy71CBtVJDxY8jSaOEXoCk4gJLaJor4DzEC64i2yD
k/JCtFHbx3F9D5mzOxfBUSYEwiN1YBtOVKAlf1fjt1d1lJLPgnHutda/0TFADcEp
rJNtKAsB+kcbtS1y5hKnlhooeScmeDZBVZfwJXeMm8cxJuVU8B0xoxVjPGlvDC3Q
rstssWfHFZcwrzWkHbZ1jraglV/304G/Hxjwjpt9DPdLMr+PrIrLcOaj3BN6jyXe
fa0ULtIynWf4p+KXla+WFF2fPltCW0JEOCH7wYfs2ldxy2nhf5ah8ecC6EM5KAXC
N6bqLwD8TkakO4BthRkUWII2aQzHectnJ/e+Q3c01SxZ4ZS/0QgWD6uauAvPV0vm
2ys9R/DkFtSPeb4esThCgrXOkRQ3xc0VLKyhqd0vOK8vJS19OFklZEGjU8UKPYjf
j0hBdSmFR/0Vj6MuoyOwbyQaQ19URWepfX+RLEbyNdTm0QgFO9VBexWuDMHDponH
/bWP9UATvKbnwkr3xPEjHTDqVWvsG/rp4dM2W8PfBTUAYoHZizFE+TqqjQr5HMWA
t03Am9i6VE5IwhwGDlEFbXRq51aVIsBzI1HW29IwaIrDCQFnxzUXacZ75nfQ8gRM
UA9dpsI3peQKeHJpdBn44rg3TXN765RIe0R5qnre6a8mhKiMdN/cBy5w77zbh5s0
0jcVHp8Cjh4MZEWU+CW1SY+cqMknVegB0VDOC9ddyROWNwHRGunqHLo36p5ShYsD
VlJ976jxFRi+odquO7DYGW11ilfhu9CsUMlCbU6gtziYdGEqihy1nqblW9YvYpXJ
6ZKrELjkJlT8d5saI9MYIKetKm0H2tMvnUfXdEwYA3or6U4VOJ51Gfci2xzNIVTk
5qeH2MucOkZIKu+Hmn1tD37goaIdxjDmfWbyvthTBXdCX7LACDSPVmkPP8OlKDIH
LFu/HYgpOBOm07VYrjOvWJQJoPIiyCnKix5y3/Wpq8wj/lZSBXiDfUpl9jDWwT1Z
WkPZeLq88DcoJBFzek/9EK4b/3+2bZpIMqgSkSMY7cK60PNzDAJRKWUT9njUqN65
S0i+W/BFFT+QNJetdpn5cdOEZXxqBbErhnJEzAFWCNAA1FVSYkiJM+idXEOaPxJK
U8W0dDm5eFpVk5k1gSLWsVy5tD0ydcgOuq/j019R5CNm36fF9TDzSUtNchlHrGNN
o0xx9ZS/iTtgybOumn1r0nnX3Li0L2b4zHq/9xCWLCsWE01sUqkmVrkusXKRcuBn
sbY6RUGgWeHhnKOrnUdQs66g+762/qiYch6Lta8jOfcG1a6BYvgtXFaMyHcTrs2T
ojeHLo/rikxZFVLaFLDzQoS2sPTgbXhcn15Tst/C24rPP4uK9j9sCFSZHlERwimS
fxuLel+AQFjDHzjid2XeQ85d2W6LXZwgcgBNCim99sftDh7EqqulikenNIyaonHH
1RPkUE/wdjP+OxoyzogyasDuWIz4OZjJXxo37F7zOeKdma/+BZBkdj+C8pe2sygx
SPVUJ3CWpJBmFKTiiGljpKu1kAY/hL4vj6o/IfnAe0XhEEXuKOkptRc4rS4WslW1
g2em6egbZZrYXFuW+ZSavp/6PnOyBIfLyvMQfae4CXhX/Nqdzzs0mWXrxQ3LukVv
dWkAmgrXHHRSeE0nm0Hc2LELXnPPjH/AsxtrWq3KBHeYCe/raz4OPCL2+lDZlALR
yivNFa2w83U3vVnlVpvXI36dXfJbftANMrSwd3Ri0BlPyHjUwcLjdjIbhIE53/kq
M7IMKy2+jNOb/pXZTNhSCsF5vbvDg48DA/mj7vxJnk8Na2w2lFNUPh2nRxXKEZt0
aMhzLrPUQlBz82wocAnxQA6wfEOtiHzupXhiXBq46CgT1Ex0uzNr8YIglyBd8FbB
qFtwlixe+XAKbEWe1DIuKiZzOqDdYGbLN83lLGqwf0DuPfm18vE+udJkHUG456X3
ziTgUIOf0wlWQ0W5UavM4Q3ddzOy/EFcxkoGt1t/XkaenAlnvvCINQ6Kl+7Ks+pD
3Yc+jIUQyDxWPGZCQhJGXVnIMvHRr7hKQ8QvVpQE/C7VBioujgYfMwAuhpUS2p33
W3z0hnfW4BXn+9V0kC/bPFXEnv4xCDAZmjyRJsCIQgaJUt9H0cF9/wJg8XeiJ48r
MkDQyxAP8S9ZR4ccTE5Jvcgt1XgAcQbul7Q7WQXjeqNTEuBIFll8Dd41h3ixk51q
7e7OzHPZPThmbtWwOXpFYn9+u2Xv8aZ5xIvdtdHT9GlPJ89ysk2PToX9p/77YnIj
0KFk76OAgcGoqec544Jen1PQJN7aAqR8W9NRkO4QyU6DVZfepnC62fDg0Ure3Thx
N/VzrmdjfH6kt2UhjHLgSzngSQpgMGalhSzA9+RpRTdbO5nMJBOS5UUdPMOuIcPQ
FC0NX9NOPxRKoAU995X+377ZfcTZctTCbfPjpQx9eYxaDyVXsY65IJzW0QozFsSQ
Rm0kCofQIs3goDA7sV+90iC0zQWrKPFl8K+VI0CcHKhQpQWlLdjqpWJzkXQH+VWT
MoGqOGTeuu104mMxqIXUjUtr0516Z++p3zOK+akHoC6zGM1TH+DLQ8OU/N4u6BLY
H38msai9zh2fjv6BRBw//VPahxqtbnKLQL+O9UcewsB1Uj+kHLRt/JwqQEQOPqZW
0eRCuzi120m+aGydIGnofn1pl5iYAXNXEY/Q/UJf+jcq0m4B7uV2dzx0SiMkiBJ5
qg9zge7ABCpZDrigbh0EPdMOAQoiyPGYw9R6DuO48ZEW8N/MrCanTPKlAOLxBRPm
FwaGk5GMLen57AsqeSo27VvNrcdXumRjCOtOhzCRFUh8lUm446uF4RQNkzHrePN9
bhP59wdAXc1wAsnkV075RgRaRUp2eTlkX2atcfE3ZmpwP0AMrOWiWem5arJ1sv4G
dpHPzcEZe/0dUmwJP2fS61+y7dws4uZYC91kUFc0pbmZnxcy25BvgHNslj8ozfph
P9gCfsZ8QHucBy9+Tubhd8vnNVyjHNFS9kNs6XggkT4s9JNYP3KPGne0RFBwzh+W
R/hdzmEebVldkavbHC6w05OktLr/KLlHrYIXP31EBilhfB6kImiwOk0mj3orsSwn
c3pacIyoSXYf3Hrn1dtTwzLXJEzCxG/0YMLllku5LyeEaFUKR71yp9+H4c/oE4XX
iB9NhYC7nCBFpbD1CI3nAukf9F1ldnT+yODegcO/pgLmFApZa8ZqmBXcGTYaw5WY
+vMeYbBj3yJaUWAZD/zuHiou4kZgRGiHIbbDACSjpQTM9onL+BClvNUab5GHbIKG
3LOh+Qw+/Gh5O4z7shAXh0tRJ0Uy01uf57YmOE/2Uosj1uw0zB3Ov05eqc3YyyGX
MjCUN0/4sf/214hDFsIqcVDnvFQTeGyh8Ey8In88nLrD0WyJTnW+lzksUyEWrCzj
qsjquMBeAr9jdFRU1bsNP3D4ieNom0Cvrl2c6MueMn57+BHhiehzeAd9qyB0K0V8
x0tCjNe2+Z1phhQdtgp1PYdTdJC5SkSc0SjU1EbURba5N8VugI1V9SV4jbykLEbG
lWNDPivb32enDiJDl/kErNurC/3H5DBCABV3uzVeqOaM0WNpNwllzTHgpeg584qa
SZffqnwTwWu2eWv7LlZmRaOOH19bOYcxypbhp90H/P2eJ+S9bg4VN4oQ7AbwseYA
DOVe8MbKRXjqNL+oAT0ZAAwJAte9vUd7go+WE6BsTKt+0KY/czkMGrhIy0QA0sql
gL2jE2ipE2uJIPCMn8Y8OeVPntzOjIHHxfG3d57faqBID51Ej9DYSgCthd2WG4UN
9/8waCWXRM6zEItV+bibZBvXhkgIqkDxjuw0VFk0Lxjpvqpwrpa2jAgJB6Qm39Eu
IMFWniihjlAp4ghwVGdOSfsJjB7zMYOZ/itwjsqfjDvs8i14Cg8WFDSGDn5sw5mY
gA99emWnhEnSmtPpcpQoErNYt7aYK14xla72PnXeQaH6Wl5cJ7ltB2bHQdCCdxb4
fRFRJKPrQk+5z7zhFAfb9VXc6TMZ6K9vo/OGS/MDVTyiIE+X7lERGJFfCal9kGKe
S7YSLUFfgJMI03rLvgd6cUAp1pS/JMGxKQXyl7rrUz/sCFU6legLNjf+Yfc9aPzW
ywZO0cDbDGGXSw6Q8JxZVtuY4UfPrTymglJ13jviXkY3+7oOjIV29jyrBc4fsxLN
Gr3aNp4HVtrJrA8ndxy8/rQecoAM7nhc1uoVe9LOF0sHLZtljJx36Uw05of4LXuV
6/T6GWVM7ouJSnBkmatdldFCI0Xy9mglhUAOMh99fI901T2qm63n1jYhvwrXVdre
Ey1uYdrdKYUDJlkc0W4ylmBOjyw6Hy23RYh08QEEwXx/ljTdf9YQLp2PIdNc/dLs
AltVOz0Csh9OcPTT7vctYpU3dF0NTgmeaJ8puNAwwu90fre3ro6UqFptz0UTjONP
UA4zlMimM9TRjMDmMwleHM9RhKhM3/mQzEPT73O2w+mDKdYJhUMWgiYfavY5+rNL
F77xmAnIStDrJ8TObwoaGO+FYZs97OngcGOHXTiooOua3xUUNivE2CYwxvKMbwbQ
tIM5BRoELnX7piXuS/B42h0xKscfmUCShnOZ7AHLNltVsdbCtqLOxaU42sHpKCek
2C/VA/hgAZnseSZN6m8tRmBbOvjkjSZRiLiXDDhJbDoh2eoGezvhLS9HcS33+j6R
ppIjZwYwkHaPILrzaqYQPsi0Oj09r6SDVVkw5EnbbLNO+J3yZnuNu8j5wt8AV+w2
Js0IkHg2t0ReWenrU5NIsNPVIzIYqX4xXvQz2oRyvBZ8DmehykIladN6NcFMIuVX
VOzbWiYO+WGouHzyzRzUqFBKP4B+uzKNaQ1wLDaS3xy8VFmBOVAUA3Rh/wn6yJc6
v6CLFTYaPPkg3oqcjtW6PUj9ydjqHqloXHbNn9z1aiEuS7BLsvkQ/69SXv2su3JU
pgYCHPx0bvbrhqXdbciSOWBqN+OKGOMRLPWezgadynqkME4LBDqPQ6h1KUy8/FIR
T3WyxMS0UIRSeSn1GIlpAg5gqSBLVTOW4I8IQN/VIcTJFukDCq3+xE1E8ZD8Ae/I
bKxwefuv8zJLXzH4PpO3gKQ4lzPBWlrpItM5GpCyMWWyikllx+j2K4B3yy7p/d/2
KgR3/ngllGEdRZ0qZw838ZkniFac9Gw42cSTxAn7PTDHW9Zku8I4/LGQulfocwT2
OjyWn6BAAyt38rLI7NXPhZ0ZDAR9Fhn4klsghOK9/Y+d23768qrAEztJLNlrzcQw
pXR2KA1t+AVb/Gw1qSd3h3JmnC2oxCKAsetHsu6/DKQqX7oIcdGtEoWPDa98pGBj
LHSAY9+gupDNiAfp53qQ/IUWOVd85aFaX6dRPnklxjlSyQKkzX7UTeu19V//29Ma
jA3rFztblrnqMNZBLlfWuGhSnpJfG0bDmDfhtiVp0eAjUQj9xJpp4uhRC3/xMhCd
9rYvAImkvwks/nh0nlo7PEb8/EgvjmbeMLHjjjwAEh58Q2qCD3eBcHLUOc9EuEJR
71tm3lhl/GXDS4l+cyyXIiOFNRud/KXiXxp5bJ/AAfDA3YWrE/A5JShQjKNXcJ+n
aWZ/haKW9TwZjnJt3DjOe8PsuzFASFJGE5o0zMfYPJpux1fV6CJFnYcX9asSjK9r
uqas3jrLdwIN/8MlTVP7bJi+4R9b3tvamZGe94Q/YLnfNNtpd6dL7SEHRVhNKen3
pUK41zhNSPtbuAVQRbgJdcisAtk9BUhwm5wU2m6PyCq2FoJ0T+ltQacNXgPUl5Bq
YrCjGad+PJZrqzA2ggbCiBjU2n0pfe5P8bAG4G3X1MfOQdyKwzC198kfJ18Az/7s
W3DFYjndOgR4KkebUy9kXX1naSS1LI77za5BNml4o/60rQvbkxTGfDBB5PZORpuW
h7Ht7MnZOWAD57NXJzdoKVz6WPN2RWIe5DABdksha9spirn2iqZDqnDfW+vanBn7
4y3dI2FnFYgSIcoIXOpsPLlKxL1mrXAoNe4J04Ha42CADK0QBFupIKBTWWnas0S2
GljaCkx1Y1vcSrNTuIXAdPEB+ZrY8eZDVDFSYyP+AJjrMopYWYzauHDM9U2jjwwq
VYyBp12U4IQqqqwqh/jcE2CrQVXxpyi2rrRZUxsxVbZFXZoNVPZUCWJPLEcBgloF
59EIFCjiif0DWw+N0NEqXcaxfZGZvLJlCZzZYcSnTb1O5Duwq02GOqp9iTb/ltbV
QapEPtx0rvXXy5p3QWs0U3FHoaKctDP+C0DBK83+Oy9OBPGBjamTjshWXB+GmqFb
bjohCaADLWe/emzc8/gdK0jrEwYAmplzeDr0r7hv4WxWvx5Nntf8d3Ie+2EMRIjt
xsqJBvlef9Gf4t8OGgFrpcxAW/j8WHco0cTVwrYKN/kD8v2WtHSaxYf583+ejXNl
jaQyw/bIy1vMIutlQdUXy6v8hXztkYaoS3ibZ8NhJ/lnzU3fHofT5JTmR86F0GOd
KoNxTPZF8QXdAANqE/2Cf/Y3vDN8DwYIMk0QZSPz8vtjRRhCl+3RFfA5PddfOCfz
9tu0jqWeTWBS4JEdISB/4mGCOI0YSBfMDN3RU64nqWY2QEttpa5igR+B2f/DqJLu
RAvQfsDjvsNlhqr9Oxjj11tFOKGvNsme5lQJOB9kVmQdqJmM/amDLFuPOTQNqA08
H6KZqweVvl51eAYcfGISJ7Qhn4NPRMXHBSfihX+cM1hxDoEQ/jje5TiKb6G18YQM
t4OVYTDQHiX32FC4dQX1a2tecd1AFWr0HwMR7nR4EJn1ExdPpG+v/NGvCRIPPdbs
JaUijLkchFi9XFeAjKrm6BmcjTArwIIF8GiBF2MGUPOufHwA0eocGZhQjQiao/Xw
zS1b1UC9Xo8Z+z11Emz6CHwHCRie657AHHiftbMSCAdUjmxQSawvsmFdUTBaKXhV
HR+Q/EIJ/xN0q+lKe9BiOnawBtyfopTmkVcuZ058bTXq+ZQYmSo22MmOkyBghcZ2
t74YkvhJR7H00rVdFmkchzAiZUcmXW6heaYOUjhF1kb0SxLm+5U/eEdw7rm49j0Q
Dh+lPn+IHBKu3bSP+yiyhG9+gE0iOweE3ddzxAiSh8+dKC3J2dcH+b0xC42hhF5K
aCaQF4dPOA0DYdbpdUOKXfJlDXtC0UFpTXZLbPHaKAoJtsfd1X16+zHKuEK3ShQ1
OMo73nO/UvFrOOInpigsi55Cnqzsx00Kyu3X2cP+GtON/DhiCvFqoerP+3wEM5+E
stowJHqdASueG0vmJs8QFDDJyfJromWRJBUGr7Y7geuLkGYWoFyIPa2vbE2KToTV
grgaDpGeGxdBVTD9OaQ8OuZAa+Ao6SKkHA3zWOw/qq5pzckLe3UnJIQORaOJ3AR5
YmyXLOEUDvHwMsnByQ0XgkB2sx4COGepfXE3m/Xtww/d8Vh9Hc61gqnzVOjjJJZj
2V3FDGUQgmUIZnAOTk8RQRcFJsspOcjuyJf02bnkJykAs7T3QT+pFft++Y1ffMTF
+At5s3TOFH6DQjaSeNt/ZoN814/vcEl5Si9/Q2RAIK+pg3y4uDJWXk0yvKn3PyJt
JI6LqLLEds9GUGuDFufnxMUKIL8asjJE5Oc6JnxIqc0aIU5ljPx+jGI20QbvAfG3
btXx/u1lH+G2vqco3ay9S+YlLCGPUnERcLQXva2UvqHeZkQYY70Mmj+rsyBKvfsE
1h17NxUA1o81BKtqadwRCfxO1HuG5K5glKHP48OaxxtcqLVkAlTLyo5TP32p/Zj0
Vc7EC9c05KPEGmNJB0nyxIzUburUBTGRYoRg1bK/MolM8HGOdyv1Qf8puBDhyzfm
3ax5UBPLbNKcXVGFbRAokd+aMFG63LgwP+A34d8uvZ8inb0GRCknBRQnavPjBcm7
x6yWPoqLePuJILzyR3ZQdHB49oyIl81EVCJ6cgvJQnrNp87gGNVAI/Z+RYesY/d0
rWuRnu8lWEXzhDDiJhUL+YajdVcgC4vk/mxy9HAqWEOgJCMP9i0VrUGXXJSg6+YR
vVEz3Ni4PZqrfW11W2lRSx2trxbkLJN/lAS/h+pijeYwzN1UAm3FqBlcXdTEAB9I
OIScP7kVBvnaJgUEvSWRSMGZomg5UY/GCVIQXp6wZ41xZ4sIs2EsZdceiHJz3BWc
d8DwNvTW7ljjbzvrB/xoKIFi7BfPg0rcDjKwy5uJV85VkrLSDiIBcU23Bji5nOGC
QAV9BMKqMJcLkf1Fac43ohoM+rbA+woFoHkjhzTSobqqaitjlUpzjpXsQt764/JF
3r91SLipdKH8X5xfvYgAferDYabQ2NfvQFkvmcODSxcnUDMJ4CGh9wvcJFyqSNqJ
Dw3pXPOyk3ZqbQ23WQdLee02t75SYiu27iiiPonJv8sSxpSA73BhPXfLqbl7xjbs
o+zCoL9LzvR0DKRzySpHSnV0jgfmogDqrQ62AX+v4Yp+y4y/8J5DG0JWxrOY6m5R
+7Y1GdM/uO0GTHgxjBpeWzZVpNbaPWRWcVACkFryh9+eGI0vnO/i54rt9jf8gAmi
9nySFzHvIie//Ej3oZ8gp7xRZh8Yf6equ2/wS/CYqClG3Ry0h2ikKew3MLBtYweL
5xRgTrlp3tARTh572MiEzK4Jd6vJ0cs9uWMkghGdwtaCnfMzHu4TLl1sm/W+QgKQ
4JM6+Z3QYxGhUKTgK7datVmllUgCbO6G3BBSVdOuigRtscElrS25hZ766qdbjcti
rpxJbEj/LyuhS6A1hQIaSS50NUJA27c1ppW4ALDLMVdXH6hx/bsJuK2RqMOyvRYT
1RTcOAXwxt43IoonsXIy7tJaXKc7r84M4DUFdIesxc2SnDI9rf6laRn6T6S+W+dv
KE6MBzz4nS3msHBE0Kpsbhe990JC5M2mKijVjSmr2EtbLCjpsn37ythaHBXq3xyE
IEUP7SbboAeDbt4oj9G8EcStICPMJJBHl7Cy0Ih1Eju5sq2KSCbuBddI/nAq4GgB
v7HzO+519UJsNvtsRJDuyhuXBcNKOaqkao+NIwp3oC3DOd/i16jt+rodgllWs2od
gRG7sEdjrPnBP7Dp2DJToXyDNEVPg5HGEJq8mVLKP6kSwIyXWWsytz1T/P4vaBBA
YawLpeyItaFpKOsoQhYhc8SwTYzYbSzx86naztvmFn3WUE7Y6EgVJOFJvX+8wcj9
7gYjzG1EUQohwG6JvkzWQZychXbiIMgjN2y3cICRr3Pdt/+jBqoh52sLKvSZaEwb
AN5ioQU/IE5ozB6gu99fbkF/B+9X+ldiKaUXgJA+JGTwx8Bb8aNt+LrYxtjrYhXB
L0cD8Z16O9mjvz15PK/VNYKBLYmH+ZYRJL9PO5pHZoNBtPQMn6XBmJPvJSSiU8IZ
8b0fvVS+ESyW0yXKieVI3GCcPZ1GXHWiZdQcZ9Uxht4/nmwtI/4fFhTQdL+qEJqG
qAS0oJCNsklEZa9JyJX7vPle8igpk8rVZv33KP3q2RbYLfmpuNm2wv66/x9BzOIM
X4daj2ZOhnehiwP5CHPuNQsUm2Yn1kPnbhnsR6RkPaa0lzEgVJBbqiHmhn9ZjP3R
wCDeMyKC3uL0PrSEyE67eNSTTavALbhXI8RhntFWmjdiQzGVT8m16jwlNJZ7SqqG
NuCXc5lsr8X6mOCHrKlFAwmiO2jrh4DWMjnlxl7S6f4yQWmk42vHDER9OtySikQu
kFvm31D0pKz0rcng43qynGsR4Pr3u84zyCNznv/iwCGR47eREwhDkaG4/BZj3bAp
lcHNoL1XeDLW6YwXZsV974GQ8YQ/nMq4D+JSL5XzqR7/695lNT5JB3q/nB7bBDoj
bdSNS439D1/aaywgNzKuAz64MgNfSUuRfMjgfN67QorTaA80PeLsgzklIzHvBWug
hZq1WPCikyyqkqOk9OvBP0SIn5hcc7jdv2oAbJCQPGrx4Yww8P02FqjTl35RGTH5
xJ6gTBrPRAlvHuvcRjaRJJ5Ni2G4Sj6TYvLFo9hFNcmMQR0VRD0BEhA2tBfkhCZQ
RRO6hNV51BE1e7YHv5Mj6eQuDL8TAjM/NjGf4KfRB/j4q3Z2Rb48xY0xkOzO6IFq
iDqKcChUCm5MZrI0VkX2eWVzrUFUlVqKDwT5sy2RRDdrH7UifGon9WAitj4zENji
p3ArXelfy3XIugmqLtkPdn4apQ8vD7xC+yZGgj2o5wt75lTurYvys/fywPuB/E/W
7RQ/EY7JUKFpbBuzLQI8W8uIxZVXtpJu/aG/s/uu+OD6y6WQr85GojuzMaeCMBBc
89GwEhfRkk8dbvAyrK6juOc3gv5/uReS7ZJusstlq7h9GLUuYJSTU5a235qmyEK7
lYw0hdj3nDTJ9clO25rB4CVRlvWhabeL5SxK8qhKjzwYRTzfbU6CTs7pFCHOsZ3v
AD38lGP6Cj7nyGfePrfp65JT9fmpG1hI1KREmrzF8IGPtOesADlkoUsIkyr5cMoj
bQftXKkhO7K0AxVoXXKKJhAQiqqvtOgIF+9bgUbbuPR0FB31uvFJucHjAMYnRJI/
/pyQkONmcGU/cLiv/exlDGEmpuPHxpCgvGfykJWlvHa4E1LY2yuThaOh7X98cIsp
0Pxk3v+t4yEUSfg/vObGVYbhNAHpTHTdaJQ4g06mXZT0e36IUz7+gviyOs93xp5y
AAk+pf2RpWxS0yGMx9+SV1gZK8bSNHFQuo0jp1UzvtDwVZBcdMJD6KEU9ib8BAtt
CQBVODhVh4X9tuygoTGH+NICLmjFThUWuGttXDI42llaqO8IgcbEPeitckBd7tox
8SDYEJdY8tRcbDcOWGW/2yLN7tucC0nGFqUfwCM5i8ogifuI8ccsB1jhXa1w/LaO
TmOWyPHSdae0mGWza+gnqLbWB/ZgZipHYz9GqLxZB+Rvf97c+3uCBIlYj9wjgi4r
MWPDgvEn60mVfK8Cjg7l2Nga7GglYiICTj2hWPq21yCqXt2zRMkva3gLXHR5TZzN
ymeS+CLp72wSXY8lGWRzYbHBBKF0bTj4XHl34tz1dAakehj9weqPUVyJRqapFcmh
yuKDSyZeVmp9SlZ086tOY5QHW6UdSOuhvVI2IAV5DBt7kHbTIh3LGQDLpAPVIdRK
AUk0C9hkTx+hndhi/VEVF4t2bQT0l3H5O4F1pBlHZvjG/NBSEG83hKAxo6Wx/MqU
nPoQJWjG3graWZw2QBkQ48vo6JtVWvvy3soKv9QUWgH91eD14NaicFxximxES4am
EYmoNknQUq1H5BrApwiH0iyvQK3tMOTLZGWIJehLHk6FZ2W5vTcPyitrclYltex/
ufFneF0UzHoCMgEsltwAXR5y+8Xnqzy6oB5mWHZms+FrS84WPGAHqZQ6sz8GSa3D
WgG3uLW5XgJX7ed+aZUKOjhRFqu3e44QBBRf/4gOZHRkGuKJ0Ssir29PRc3og7Vv
pz1CnKzwtlYmRthgQdNaIGLOKcFwNveJYVkVY2TfFZp0XNQpQCALVGGf/5VxdDZa
PzXsq+Dv91qzAaeTVVNXXxVpszTOrsAsKRIPxzIXfCwJoV00EVhPESbLCygyDNyx
XsQNaBlOL0ls2WC7X9hu6Wn5ti12tNb5ffqbR6OR1YA3PNWSNyvfcF7Asw64LMfk
34DKqrFHFaoq4qh8uA5se74HizNMLRs3ZkoJWncGSnFoETIOt4K+cSE2K5vb1MHo
nrMtct3z5jytgHTkRfd0FFUHru0dEojq0TMCDO2yuj7x6yeFgnGMP6UJeJ+LyfQG
ZUIei6x75jMrpb3TS7n7fv5MSqE2+AwiEN+AhBW8L4otTDMUp9wAqKyge/jny121
fdo/hg5vao+ExWIiKdSWHREcQ0Ip0nhyMxybRF4nGUxcUFrnYpOJaMInhC2PjgxR
4zafF3t7F3kdf5oMlUVqhQUwBnasjtviklvf79Ds1DQ0lY9z2gjV4b+Uunx9x4Ft
ywLotjquI7RsgfDpGK9WL1zCbjtW2xOaAllgbmBaUkvyAkz/XYO/9DaltR/4fmFd
mzcwjA0PGsffEcR+wILq4Yo2RDXx1tAz3RDRZttA9qSKCW27JBV79g8GFJmNDPZI
e26IS8Cqf9LwZCtsFRzV3lboKZv1hNz0jsNx1Z66BoAB7TW71fsNFoty5DqAtnO4
fh//G6blRxrtK3MIIbM3ocGf9EjKfPpJw7nlaZEzx76NYA+q0FjzahN/atoHOoS5
srq/7IlFxedAUTATdRzuMmTyppQCqZi6+dKVLED4uagFKgRAbOKiYcHwlJ0J+R3C
Fy8Up+TaByBMo4Iw2aX0ixVLbYKZykb/8aneCRspoUbd/GfuAb1VJ8mCYAk4+/xz
HnSnyla5P4j6xrt3fuEwcCXhxZ1LhBAWZX2XdgqC59nWBdxHB7dBEQaCcYqauvnV
kU0gYo1kxWIyMjzuSvOlDvhrL4ghuSGeYg4fABYLQSHGJDzg4Q27Pg4OmlTeKnH9
qGCn+zRxB2mqNgW2KHTiJOc4SI2kV6ZSTO3gyPSjfZKwvljQwekT7rydltn+dF1j
cpYHJKAqkhMvSkw8F6oacVtvvxguIg0MqLW/U3p7zr3i5YWcyP+6pxKLyNr+Y0cL
xA/nFSIyxZYb7pVXTpudLJRLLm6Q+EnTjL0S3220q+zVwdnPrO2iRlrxyOMf9g26
JSVQjLnkUBxduollmGixs5twKyODe47+a6r8YcMOJbqU1D/pwF4vc/B+BkDIRIRQ
z92mQzkwSjhHRnPPLLsRClkDIGvt8xirFtKULtOM41lRibThUECEof31z0WrhhBZ
5D5buOc9s7zZ+kWoU7rl0W3+qcovEg8lEq20xB/LCwPLEDcBjyILTatRE8k7Pq1k
Xaa39QzwmZXVfd8maKmttQBS7mgd9uCn28MsS0Hxyfv2MA8psTaaP07rhT5Y3dmX
05d0md5HFx26M7hcYuGVGLrrvKiqEkaacfEP3t9Lg5Pa/5EQrIydcG94UzFzGokG
m5YpyLbuO0eJvXgx6XNaLVkl8oB74FqiXt9BF+raR82t5uRZBr7uDsDZnoxGTJGp
SF/WYeYa0QNO2u/OfuZHuwHu29UwRLc1seA16IlplbpBcIqbQ88muOS0ToP4y4ga
taIH/wZwLLeJPhcCSAbgozk68/VpM4b2i9OTvxQVKVSmcSwZkJKfNYuIfva76bx5
rwlDDaeEVk18MQPZNEx/6E5SoSqMaeRKt81lLnvz6UFX+LFlUKMl/f0nbXlIzafU
R3XRXRX/TM3feoybM0KIriO0ZoJ9z3co4fdGvkYc9/gZg3MXePmqfsv6Reu0spoZ
Miwbgyt4aw3YwQ0e+OJ7JMLBs3paJsHnOFk93gp0uUlYj19hJIJdTUYktzmYwbVG
LiwVk5HyMYSj3StJpuxkbkstuyW8Pjs4/bqDsRa8Yuv8K4xd9DUJCFWnwYtNRqhb
tMHaeTYSzRHA2uB3ftXv9DYH9NeGvZOD5deso5vPeM8+ocqeac6/1VBaavHGoz6I
zjKofS6NyTkFfXE+khxZoaFnoTSVrONaOGXV1KmIwPnr/T3OXt+r/5JnbDrbTvJS
uU6UTrE401o7zxH96y1G/5ACR7FiIoeImaqg6ycxhe6ne7w5WkpWa9aognPvkyMI
ZE7fd9fGQqHLJjKkNOHT0VToY4R19XpUue/4oqJJ6pB2IZbc9sMlOXca1z4YzI4X
6as0HLwmMGb8sb+gZpDcJCF+PJKdQWKfMNOXpAoSyATs0QQpOfesbRr9QbV9Ofb/
BrMQkYhYGckJ/KTOg9L73/NR5CqM7XRAN1sPSg6RLffa1M8olBb6UrLbC6wX03vN
ahU4jQu4uROQ3SZQTtrADg12wbawqG0V+Zxxaq0GVRbyqOtePuY44eq3XDZuyIL/
nYxUqIfBuUCFKpAqIwn6glZhaiBogH2yAdK/WXBt+9E4GsOtlmHcmOuIRxmDtUzx
ECftBvCQsgYtwCkJmX18dUdUXbiqe0JkTz6dWSyr1jG6jWKsd+Sv4P7ZNEc84wwd
K6io8Sp3horrIOsKs2nOn2ACks1QbNg5fi5/Js6Ba1Ztp8tXz12QJPmyXqtvmS0/
Uj26Zav+CDOmCPv9y4+8VBcwGC2OhlO4y8fmg9XdB+YML4CJCs12C3yEj96UdJMF
5o5uuVk2v0bmxS8PvrZBhx4fV22V4T2n824r87IfJXHFaJANQC5nlKqcReMSxYLi
BCgaGoPIruQOVyKKB/SwqKvr7n1aZ+h61cIQR1J8iT8M/nNb075frJD0a9irtwQt
3HvoJ9GmQ/ZBvUNFAm0CxTXo2WlUFJQufs8BuCxjTMsZqFn1ok71DrooMuCFZ4ak
WtVo8Kga9uc95SiQP4y7NopFtg37LpuVsSmepjtVvsPLUv6hUQtxWFmKkQ++2SxX
vVbKqjXsJw5TScCSmC+SABvmZZ98LPVdzgOCzOto70Jzc6fLeLSknVxw/qjdZrAH
tz9QO+O86vohAlSw1fv3xsYkEx/+SiwBwr+aWR1IK1FUpbhGfOQ6OMHvrywniH9L
VroV+NLVeCoaGfZQNWv7xhTQJfAmdtGrZ+ft27TWq774ZyZ0WDrdW4soYvUUFsLO
oiG0rXY+Pga1OIZOO8Qg7pdX1o7KgKp/qSJhFlt20otVDvm6fe/Q6TzeJ17eqo6H
dgb27/Peb9Lx/YGIVaBjAA1rZGRGLXOVRWApimL4ZsK3/8/VnNtINbcJhPe39+g6
V9ExbYI/rBgNG69FD24rZ10NtS4naSM7LIfITdlYpxmnCsAdk4UF1vj2kDxT17Lu
0Ts9lMqcDyyBv0x2V4qRl7fs5L0cIIDNPZDwUFVnfvsIDXX1AsaMSQ+vhSE/3XSH
LZ9KoelKU8n2IR6I5+WYMB729DYaw3dqXAvZqx3qrt2zGeMPUQXFX/cwMXikA0X9
es2RIkhDyXVpQKdgbLSu38cY6JPsc45g6O0E2y4wX8qJZWuaMSptAkouof69CVid
oqTwDaMzbJNgEISFGSa9ZbWwYAckDWUsMtPdz6cFAGKcSLYzY61PvOADoKHiuuzn
P64uqWV2wBPallrU5M84GQkEOwkTq06Zhr2SdbnHccD418E4v0Q7aQ2KR/UyEv0t
CJaI1yVMekgAYlOAyDdxSIRiv9Jl4+6TJSK4HfzzaF2gd3iv4ihQSUyu2DI+lZ5d
uUjpEykpt2HNGaNtUsZWSIxcbPdWctd7Emo8kcva8RjPDYlpeFkuXT4pRNtgtvu+
v5W7UCKxVT8M8+gOMbDCfD6Jh/+UaOaX+CGFJZ+vl1HE+1RoTU40/mPYyxKirjUR
L7mAqADeKfOc+3DRtlc0qZXcYwxoPAWy9FMQb6309xrxW4NffpV5ez3mhyVrd89F
MYTfMgpG34LnBuXi6Oi4qAc9IrDuebtTsF7BT71yz21ZuThLpNVZM84jgbegB2if
upgSvyq9ZmtNj1A802ubCnPPH8C91mifJru3HIhVZLF8mJePt/NRF3gEw+rtSLlg
APjUIwlkmmZQaccYx8NS4k6h+G3RzJ9h/BjG5K0xrtNFaSLgPIPqexB7DUjnAYGm
RQMTDbDdMaLwUX/xx8NhJBRiDlxoPYRgNiDzRkqSaG5h38Ui4buZIsV/wuGi1JSR
cX9MwgM/LevBrW4txhAbVkzdJ+kNFZpAWdAQScoJ7wixztuzVbMBa/o+AHtWmphW
tT4mNSuPr/ivSYzpGcGF1S2DxHIhYf3EDYbzkScAaOPz+RupGkrT3lFkMORuS01c
UwsqSRTiW0HF7ZJH1LHJKNThJBVlh5bYWZfUr+Lr36EW6veQCqXpENqEf96kjSis
44Brb+SwqvMwLtjymdcStJoR4x+WsDHm43WWMB8c6+kjpIeYxEOM/I4vbF2PqJjO
geJuLByZ3t+UJOu63XWg/UPYoLqsWx+lF62TDRH0Sidv6l8GpXygZ8UFZx5ZuHFd
B8fkObyO+WnJjpEAi5z3DBugpzMSARsKNxHAOIYjW4u6jyL7fX9W8Hl6/x6ZEEVs
79NzFTSOHqFnWu1TVQ0RwVw7suKEG7sxySo7RkMZpiVXeYE7ShBcK45C1lWeV37s
35/5zg9AhQrrFwoRAAD6r34R8bXnQnioT0QiM8OnZJC5tKU8up+T92Hei+pMUqXe
avop3hKkSNmzktw8xKsF3+zgT3DnaJjnaTxrOL4CRBrRrbCvyGktm05OT+dSerTi
b/O3yEV4IaT01UJBS9Ap8bXHct0SkFxI3yIaQ3gZu4NqcbVLvFa3v94bS7aSizoQ
RJx4CN+pzUhLX0flrQSVY62ZHI7B0en67NWtbluSmWkabJZ7W9U600IR1/6PGkFe
EgGFl0Ne0s7GZOVtFPqSs0T2AWkFNnlBrxY9bn4kLGqZ/DbkYhD34vcHCYQisJrA
dXdx3nrWVdroUvuUeqoaiUxeGcmokLqIOJyncjlTMtSxTDHIn+Lm8ddzKr8bGt4a
/5VV1YD2d/7+4GSv2O/ablctuqK4hKHgA8cm1XZ3N90L0mnIlGaxQqb6/7ZyUR+y
NXEzgzyW8cab4hH07I0U/36gUCVx+N1cL7VidciO/Zkneykz8al02KL3d0mESjil
8NchJKkWB6ShaAmimnCzaq2Wzei6GZRGeboyVsRpPFqm367L3iAHqBy1XTCblo/+
ul6+6m10WedRAS5ZqCnVQazEN4yyF/80toMoBTNAYi3kzbQQmhaTXYmFKJzR0aZx
ARa+5IfgG9MyUTaSugd8K7RafdefNPSpA1txmKhPsEqM+i4ah03HGS9LA5nmdS6R
duJGD+cCF13WPHy1CwddBI4p1sJ0scG70Avkkzyt6aU9bpmGm03Kkm0KhYUUSPM0
TXmuRwDlQjB+WO03nzp7BRhGSIEgg9u69h07vCkg0yjR43biTeRn4P8roRKGQW/N
KRYUZXlthCfscAAUg3IctyHtlXhOiwzCo9gWbR1b/dVGRmAdvsPqeVqb78OeiTzS
r0yXZ6GnZBK4Ejb/+uf+OgppOY8ShVaWaepFQe8UBHvf+aBtE91PLMo7hNNKQBmG
Tf8nm8TaXzm9L0z885L5Pf64RTp07jFKwZ/X0iQYL/l+H2tRVsZCt2S9k8ammWXl
5LJMwIvZTCmCHa5Q3c4SRU+rbcN7o37bClbrnO/BFtxmQnK0cYRvKLaeFuhMvUjT
1AXGDOIgz0CWWsDsWLswsnebW8UWWvb8zw3/QE+LJ1vEKooZYfGgHSYbJRZDsbU0
+dAXEaumoyB5fpGOTi6AKpS0LYIuLrkXe1gf0a3uGaHtaxEP8BsBJY6fBgXonnxa
QkPjszBUik9LI+4fD4EoVDhJHVVT+/ZsVGW0xdJDYHgIUlb7xAYrn8yhZta4mL4q
ZqvIKxDG1Tq62UecsWT+EbIx75Uo/DQTsgetrObhNYJ2c4GIuiaDEo24p9ejRR55
NNdYHKQq2/kQdFg4U8TVdahvZwIHyq7vjfdP/FuxaUw/O6bJDXauInXL8mNjXzqp
iqC4MnZvj5ZQfDx8MzhQTiv5UHKmOwG2tMK08jFGpQ2yVFeW9av1qPncgQrETlmf
zxjZJfIeAfC6dSeQCWsh0bkKWQCrFTHP1eCfbN/eTHXfXExkZuuhJ+zYflOKYICv
637/clj94Hu4LaWdfr87ETi0fjCtuuq+zDX45smdq/gCzc9Q18v0BGdkgQW4BqcQ
d1aQNbTQHZqhqxbF0V7RoCoZ/CKUX86xXcGNYjjsbIO2FsZOeA0XjR1q1z2AiOyO
RPwze2/quuHtVfW8QnUCmsCv7MQvC80zG8kdJ+ULjqBUHAoM5rVNzI8icb6VOyjR
ByRspWwiau0lXF7hOHVshbSmgvohgdk1FwoXb0e5vNOnRSLW/ksLX8TWPRL9HxLQ
HF5VzAutOJt4/BwLvKk4O1pNJ+ZDr1+AlAMYjE7Wnoc+vkuemJg+q5t/p+YIB4I6
3Ql/dCFzDyudgjKVPR6QrTlBJ29uRFodlGsMrlMLm3wympJGQp4aSjzeFEA8WRyM
4dZy409/4/qkGfaBbva6cq47+G9OqxU9yZWPy9tM7ORlUlEslh5ctuCk5/Yvpkqb
TY2oZ59V2NtOOtkH6ebUE/PiLzdcp0wv2/xChjeW+8WAdgCj3GfLA7i7TTG0ZK9S
SaqqlV7SJVpQ361wGUz0oSU23EPapetDZ+OY2Do9jmFDbwKYNQIgoJoUSdGJlUnB
iUFsrHF+6EloCIjfutb+0ES6/bYpdtJchexUWvAf7cg4fJQW31vBnwB1BIlp+q5w
X2Qk0vqjeZE5Ly5DYsc/r8jD5Y2BJlr0kFgOt99ljfdJNrOyyZA4XO+H9KraMpi2
Gz+MQE1WH72gq6dAHapYP72xnK7tuqP9vqZHfQ8hz7eT8DxXjGpBeudY1b0Zly3H
UhuViSIM1VHM97trhX9m+ARYtDFQ4n9II+HvFnxbdVxHZdMXPbfqp1GNkRIXfOzA
jvjohujC9P1tQF1aYD5kvLQDSCjOi7tP6iWu1Ac7Kqa0T1w9c5U8GtX1/jxhuI1w
LpP4X5xth5DCCDgl6iLmFXwJGkt0Q2LSk7JNSu+cRKvZw54K5y5ET6PvP28x9J7i
D3UrZ61WRfkux7L1jYI3V6k/bBQDT3qwY60NeJUJBQ2y78Xb0Clbb3mFAg6yGnmH
5AKxRrsQChJ32jzRGhxZAmfMWcJN4krblcathsrxW4N5yhWOB1cnNLAoMZvZ/jG7
7ZU8+oNy96oL7/CWJ+qUZ5P9VLLw3EtHhjF/UqocrVMIluU2i55E0vZd1a7BrqSC
wLhXe/SU0lZSJaJ3lIEyAp49L1dgdpG36qhqaJUb+zLcp2q8at+18k3FeaTo8XSP
7vQvWa8UoqSy6QJD1RvfwNU97K2lLkpesT2EyFw6xbaRHLNtkbUaBdC5ovMNRjYb
PxGzm8inoXBhmUAQmq2gJdHHwQEgKkcDc4cMuceqJbCpoWKb4N0/Gj6XJptJ6cFE
NaVr9vj7O3fRZR6kKVMAUqSj2XRV2oJq+hMmJOQI+jC75xqNvKSGHylPHdYjDkkc
Z/UwMYzmzfVV2LsWEfut22HZb8DAG7N+fR1ZGqrNNAR8Eypd9mxkFHl7QGD+iC9T
LAmneXJsybXFBS0MtCub6NAq3xV1YboW2fpa5tO3sglt9D2dbHIWUyVGplpkkPgW
p3409xh35UOiIJipPY4PqF2pcm0FmONbsW7LkZwNNCsGcgekihCvqnZTJOVod5DU
7e/dKM8q03o9jM7RkCOUSxvQuZ4+lYOGTq3ta06C9owlUpkjjfmMfECpnKo7gfP+
pV/4lao1qy0fDHNVQ0BsRqGCBZHz1MYKfD0Ilt9YenKNDyfaacj0+jV0DJGLm9ox
ZPbSQMOt9jM4no47B76Tf7lGlsv9MuyhQwo0ry4CdamU5OTSxIerxNZX1Y4JWIZx
Sf6DLkBwEHV8CBEIdCIBcpbiVNb1d3FYBBlbRT54wiu8eYTUR0ZBeBKa9luOwuUO
z7TrGrb0+hayo9Z8iYNCfcoha5k5M25xwsuvCbxNxrEviPmmxEZcG474fyfvlGUd
mh43VrsX/1/rOb0WIq7f5Ti/xEff/I02FuF2tbVON75MO3Z2DJRN8lADhOKyOxum
y5AeVI3fALZj+uVjsjrMooBM+cPEJpEHR7iSs8bJ347gjNBEw3MxVkowqqXpyhCJ
JX2b7jYvAp+7ldVskdw90j9HWv9utNukDNx/PNzCQ6f4vhipZHH+cs2r+AUuOYi3
qgTzGyyM/lstKG9+HfIL62vA9XVbLFoYlHMEV+F9yJcPRErM01OXfkr5ZMWSt0Pj
U4NbQ+y3WKjQ1UBj4MILfhL9TZqW9S3JNqdbNz3aeuGiFmXfL/JQlIPokBZmiSU3
bSHiY2ZYjdadvfCXNTSozyTAiDjLJwopeInj377XYOOgbgWfASJraxfHEEPg8XuS
gm0QBjinPmE5ysJV7F8X3D1GQPjbpjxs9EHlU7ykYk+FnqAqBx4145zB3dZED/vI
AWmGJEDxm2E6JOexKHf4CIV7o/UqZfXwTMlYi/yR4Tn6Ej26+ZLh9Cjzob9910Rf
beFCPa/l/54MKsNmunoNMzh89+Q0w6wOGQGAOfQyS8xefJHa8jo0cFcuobohCtXe
P+C9U0JRoh+Gy07kVBmBA5H9TCoSLAnmpGy6XSRBp2g1E1Lr9nuNi5IW5kuSGCzV
5CCMUFEkTcgkNXKcixKkVTQHAAvVKpz3RxaV9MZyjtwGGd2frQGEv47QYZoXggYN
AbFaWJ2jRXpW13Zp2WO8HLPxXmHYHt9Im7DU3K6ydF+Dwk1O1r9bzKCpjrXKgPIe
jhMLdQ9nXMV4iqd0FK45X6W6IXhTog3F3U4oXFloKUWTl+YeaIN0pf8ZUR130Gta
Jz5WeO/bZya5eS62vAqC8KBz9WmCwf3A0dlroBllY4XVyiatzpeHPc87W43uJiO1
oECOShFvinvGmDz5JiLqU/fqrBZk3/9/xw6yevoXpn2ukq898NtNJTj0p70YzQVG
jjY2cMxi/oXDiM2t6SxDO01OIKSwSV3ni6yslODdIAj0NkQSJX0NvoGWz4PrK2iE
JGuH1BQgX/4/dIu3kzxfBGnxJiqy/IoL6ddC9xTXV5P4SQZzkA0cwcmme7Qg6FIj
7QLb+fRFhHxMMp4lWdBMvN1LHudI1KS2CKjDuQhRaHxMswmRXHSZoB3ZKJ0QSam/
aQ66bY5Lci+7aQc1DoNmzChRF8Dp+e6cs/dTzvEdsbMT442fLp72AiplyC1XqRz4
KXDpbZScIIqGDMVkrdVmCjs4Z4SK6doTCIB1npDH8+r7I5MgVp1UAtAB5G2tLAhq
v6GIAk5j4ptTNgYM0l0MTZdm116vW75ZgMlc2U2w4dlVn5MmzFDe2YI2wqXpJlaN
MpPI7LN48MLKwlX3wTpb7P+8Fe4q9C8WKPNms5GPe9I0L+eAoMOrniArMe1yxXfk
zg5Ajj0ZhpoNRIyWArVo07anCrhKE24MBmxHeJrRvLalWwOo1nlU89ILxCtMT3uN
V6+AjPq+lGYxiLJynoxi3K6wCC1oOzXbs5/JekCD4ylU7eKlUC13QdV8lPqbjsaR
8bk7jNQvzVPNGbIrLAW4czHZ8x7xba/y25+10SQRAToI7Qv8dP0ms3iSXSt9KPIt
sd7FdqCguyG+yKMeFoU51q3TdzoAA6dS61sRhCBY73fzIuCL/e+WOUme+C54jv8n
sT1xiriA6CwsJTRFvNlE1yEaYzSOvXgFeryltoAXIAZpQ8tAakhD25cCynwYDTL7
WEqx56zPQiJbxWkzdvWNfj7CDtVF5+j6jMSHn7fepoF8lbYaOqrURsTa3TdT+PLC
bqfECqjPOQOCnFf7ihFKKkGJbYds7EzKaGAvrIHzyIhRqXmrNfgX4sghdwD12DMv
WZNTPANsWYODZS4ZGo5OBxbFayxmYBkvfSTr5p5fdTZQuphQmILAn9uOReHi6BUt
7SCFXsJLJAZC777qkXNv6ZW/nIou/PH4MAs7CK9PxM7hPWNYZVDUnPcBjgd9q7Yj
aCHIiRTMPqpPaF7ccKje0Pnnzsv3u5c+l4+9lMWBKmEailrf6TPBs3wl8u0LBk7E
HUKS8nQA00ilaLrP89D+jmMeABVWkKhbTX+AEhBLgPWsmc1EUOAirzrUNvBQX25d
2h2s70TIFjHsPZIS4Vg9p3V6drNjMEyI2GYdjJyGutMpl2qfk2MYEZ3il3Ha2BGH
c0Aa6Rx/cWrahnlBWHb4v0CEMiyVXLwF+ikZEJaeU7D13dV8+FDTz1FDeBNaG2qD
AYOUYBoFvOezbAsIDoTTNBV3pGKKsj1dMIAEXmWJcYPpGcYh1H0AukWK8m8b5c7T
W33hf5hxSdoT4UnXmUgsz2e7gycfVAcw20dBQf4HGQ7yjxVfrJF3Hg89F/p2CjGb
OoZG++FRWW4RzHygmCSYsbZN76ul5W6h7AsBbdDxeIxAENquZMJQPacKudgOA567
PmUZYMk7oePLkRsHUfm4IgMaS6W9VLWuXDTIkEi36KSK3vnFyN0lYWxNUAhI7u6F
7ptJVHxZUxiPgbPj005xvLPQvkklqs9L97I9Uv+9a5gij3G8MC4Cp7eW2a2vAkn3
PrRHOiXJ5G4JxByikk02ycxNgI2V/CabZP71sQy2iWa1W3bG2h8LTKDdypc2ilpf
Ldl4JdNffGx2g1r23LcjMBu4Di9gs1lLYZe3O0vvG6+QsDeX7qgPTk+KG2Gbk9Af
wTSzyxPuPjFeY42XBcPBrQXrb4bsc9YRwxuLVlKLA16v8Iq0CzoqIGLvKLjUw+Mp
Don4Ol4DRP3nWeP7G6YQZ8HDUKt++MswxEYPv9sg981YSegZz2y/5MYPFxqkjjDI
QHOqh7HxWt2VxGVSHToR3sCjBVpujb8bjocq6DyP5/fnRc58L2nWTgRRrLbLN/GO
Ekvffl3n3vsCYsBdmDpny885FNrdNWGVn/2ggV48jOr+nePNnnopDoo6HxvvRTmO
LipAddq5koS8x5HtPry1hitWeJWhDeyhsuygDfvgbdJs7cgc1GTZQ8FWioknMquq
Zf+DPffH0pGkLceJU2UH/vb1KR5TSsQfNPqpOBleU2jk8j/N95zdr7e67i+eGInk
l7axVQ2e/RN0sVHc+4v4PKp6g5YzragdHVApHNCVKwblfo0b4RgKfZ4V9rCEKVC2
+i4y8v9wpLmgHF+C/s62HJEL6PoyO35uHLIwx/4rAo/qZMSSLWmp+3zgcAmJwjqS
ynbrBSEeMV8fmHWlNukgcQ6Iug5HAIn1/FjokJ1Zg/U0MvL5YqyvLhELSLFp2y5q
xmrBXtMnSEfC6Hmc0dVnXbZK5Bo48eiUAyfe+8x7pYzOrg4xA0vc640o8g8t3DFl
4cgmv6IpamhMn8i12dAC3J2Tr2KcKMQ+tAwyEHzJkA20LRaSpQxMixVVHRmd8CN3
Al1HC5tpIsNahXDQvl5jZF2ZA6MhnKO5xk/6ZXwwf7JjToY/819a+hwz6/bGfEyE
WNZQ1oth+c9DuyJmJ27YOoPiP8oYwYCZ9iOXAmSQI2efmyZHOgSrqsCeBwW1Xa1X
YEkUMreyjr8/PGEUCQqtceVfkN9+d0XZDUeGH0aU8PMmUMLe95ktu9Tb8p99LjRe
wkBDB0XbD1IB7MfXvhZs7OkqxGxx3258F7+paIhMBtVWc4dmnhPa8oAaTk2DyqkJ
dv095I3PmycY/kZsvI5yNuUfZgi3UbHVfe52zyR1u1Ifl1i04B9Bck6t6mxthsJl
khF3i2LaUVKepQG/f66SY3haVuHZiYeUFJMKww7qCtgdP6XR7FIiLZcBnDxd5GZv
mXn9mgThzmlUwhx2YhI+sIv9Mi6i2LrqJIEyXD8prZv4vzM/EQ6sow2eLRiYrSBu
f1TFmmPEhDgpb0pgPcxOlqIDKY37I1DvPZgX0ZhGeVkgxuxkn17o/TP1dfk2njTC
Vd1oeSuO3eMVJ8VMcYJ4YayIObJXjaSHH+KYQbxFXQKx4uJXzH9F+dfoKietBucE
2COTw6dfrLq2Ep8E7Hb+JBWdcBS5q3wXPJrp8hongtWis/X0AHW3B28CWHuWN9C8
1wXnApvCFxzdFsdLvGoodYAl/yrKTGekShUxFTa8huI4VzVP5oOGbaGTsOv2PiR1
697Fv0A/0rQ2wScXFlw3q1vZpqo7V3lkc8Rykx4QqDZ7pvCEs3vXATduedbCzC1P
rfWDrpby5qFfL7o2srLBNSbQuQXbG9TOb7PPXdtsfdf46M947Ik/x5JOY6z1EStJ
JbIQWwwAnAGqGqOeShWo4S/Um0I99hM6UzZzDY8NorTN3ovMmycdLExy0RxKqEZu
rMuy4vnm3S3cuDX1cBLl2ipVksVXiqKs5w0+nmFvqjYVAJ6roJ7ua+on6/EgE6rd
w/QLFtI7BVYv+uJufqiZguU0/s52DhONFMGZq/uQA+r5HzpQLjVVIa+Sn08X2Oxg
L14tCpImTBh9QPXBJjxX9ZXze4u0Gy56fwQvv5IUEheMjiFdxkyCW0XfnN2O/fkI
gyUJr/WOsOJ6aOATTagpiG1cIKCUJ6STubpBYO15QLrj1ggZlOM8z0KhNrtmkOJ8
HhvLrf5tB/Sq3xy3vocrCfprq506Hfgd97kA+vpYZo2nYb6NaOqWVFjj+UglK/b0
ZReiqbFMcfvW7U4Vk895Qrgr5DszmJzKP9E+6KJyerSRRnPhl0PX9nUyJNpB2+wc
yfO+lw9HwzXeoZzDDPjVC28FSqyPKAoWDwUg2up4oV3pLhdUzpIvg5kEHJ9iLfdL
xgWhGCX6C+1nN7EjFRDJvwKAa0d0NgVVo1vxkFVDKjGkQmC35dqU/ujrwAlv8/iB
7+Z7hnjwcZ+g/xGhv0l528C2yboZ09fxnd7PJDuNLEUkt4mfy8Z0vomzRnhkcZrq
VSL/poTwLQjORzmtrKdxdiggN6nvo7BhVNtda+orXSRtnUSGnwkUJHc/1tdixzZv
prSFC8q4dquJvYeD7C87z+aadaYjVCFlJbZi57Ly1fA/iSDdjgaCyJbnnFed4eDV
0N0tL6Pi1B1hNnLOUyMa90y+6SPjNn8YAGSUTE46GaNZEo+49CJVAK5uosZOG3Ys
b0qrRg2BVwd2/iKe48FS7hhHx9YlGvsLr0n7+WfRxQK2XEXez/peBYJ9PLI2/bq2
kYwMs7tFNmU28l5WXlmoAegT/FnfSCTohnLXPTVxYqVd6v8MTmN3cjpzuDC7yy8B
mNS58/SuWV0rIn6pMWIs2V5RG4EIGjmY/s+Pq7JcEZcXV6qx5Baw9jZZ7f+pl6Jx
rKzi6bROGWcVLmc6lcIuhTUQtgDZCAX9lLQsbf7xl+5UdOM4pPBioY7kPNObZsP4
QL5Rxm98rXEhY8mtgEenb+7sctjbOSW8bVYfDIH3VXRvxXjZT7AZHLOw/NaDYOLJ
J2qrGNZ/ZTpJio4F6dbKfieeUnM6bSVoEy0et2+SvkFeRcZ81DZuwQ81zxewrzlK
fqe9uU/ykQyIUavKNZEdBvEeZV5FYqoIXY5IgEXit5ITib04hGzUxjmBma4emYdv
uakwNDf8CvB5nVV/o+fB5j41SF47HTVrcQ0l/+L42Myi1oVTFuS9NOkX7qgns1sT
1BkOJC1f1aNUWOK7llEoAVEsvdAwx5wfc/N0puaTRALojT2sVi3hwzgQ0cxLYkIz
+qhMNwFc4Yfsft/PhjNCYMDWpCP4tndyBfK319dmzCWtUCuelrZojlK/6wKFegXx
i9T13IPWb6BGBoIlaBQENcMDLv6DoNS9ABCBcxWmwiwGqVQ1PlE0bHnzz3SSWfGm
zehgvv1SLbVzHA46j32BSm1AbAhmR/QtFVH6DaUeizlCxhFTWTXPl+LyTLDIubAP
6pPUgD4jenfoKOu6IALKCPi3Z4BEixOKxKIGUQzcBOeDuwcZyeW8/i0qcsKtwmTx
/4sVgI0rrY+bmf2rQcjMHP8IpVH8s5LKNa4yH1lmSCUjwgpt7PYXtqWQUYwDfyqi
hAp0YxzzufrDy1gr9uo64MIVHk8+IBtm+Za0sBMrfbaIo6taQcjSabaaMt9w/0+X
q6nXKlsp7huCHNImbjuJ+LJIfYXjuhIQIs6lYjIv19rclKPTZE4/pL1nCbb22m+/
xp7WwGatI3ApyUq6W9KllCv5vVQ8RbVtLfXuuNVY7Y1AiZm90Xg0QDXi77HBY+FI
SvM/vFtBk29hVb0MdMJBtCPWFMIChfGE+amGnDgxmi2gUuVu9hFnM7ecpQ5ctoGD
Wgu7G90jYxxcj0TSNnzVTKWWmo/pkCsvdMmIiiJg2nJc2e3VhdLkaJmpxXhhTg7l
IgDVei6aJaKjhaAGr4BSjGRE1JPnysefrmY7zGsdxSK+Q5Gd4OkMMCKEC0yXlMx2
wX5JI2NnX148Bns0pt84kHsZbrpO9nUsiIZHUwwYrM6DJTBRN5s0l4JJrv5Z1qrh
uw69UMgJYW45a1uz9BXR0lZ4TdMyC9EAsVPZJime9y2eyzB8W1dmTHfCCGg3gUhq
oHJ5ZTEmYUZge5mOMYbeOpe6U64sKbV5n59qRDq7waN/tV5YVBG45ACyX2R3Xgky
u5GvYnmHNst/2ZbulIOYzwKGh/JfMYiM8akwpLwaH7nMJByyEkKND9Bc5qME/IE9
EUeJHDZkpmJlJ/b+nAzCMe7NX7u57YmacdYHa6o1zEpHMPUVcWOJqS3B4LVmAwCj
EPqHFE/401yYjafYr+fY1DQSWFtJQXCZ0Cauj1/UwUWrlBQzI8FGmB6TPNxDA5bx
9ggz8+ARZW9BTdYyZoMPo9b4c7WGfjMjbyvq3PBTA1lktNM47jS5lfsZ2URAJ3Oi
JusULlaVC0Td5iKTAl7YqIAfCLw8dN6iJurYuT4GZZfhNgMVnVE4hlqPF4Xo1fuq
nFjjIi9BvkxlIezXk12ZMV0czXu3Yjga2oIK8bdNTzmIYSeXirKf9f17w4zdi04x
hrwSZIpjPVbiwFXuiino7Bk1HCNPIFeFlbikSzTZTgOtiQLSChxrqp/nTDDfmHYt
l1FKJPDp5V2tJ8rHud+e5YodcHykCcy7Yasi933MRk6tUaTAT7Knjg9ojpzkFAGw
GR+a1tkSklDnEoFNF8AJwlaquu8SADsR8S6XFa/bVFKRXUFURRsezuXZzz6bkV6g
vSrkckRA/S9bDmyoulEgVchVu4xfk91YOa3nGPZAPk9izIGz0r3hnNPV8mvzdz7k
mhXmeoLO2NZwFa4Ic57dgGtysozc9ykO8heMm+nhSYdJ00Q71gHm/tiQ/7FHwvn3
6ruVKRk/MSlSHWJptWkAXnkSzXe+FOf6I/lpFOu8W51wxv1Kc5YMzBVml/u0zayL
FHIwUi5zNdryLygPJiX1qzXt/N04A1BlLnvDUq20Wr8d57wXf8m8MBTkdKP3VQiz
K569RzqmiHREKY07opfwde+KiChOxf8sSHKkXTcTcZ7SEIvcBk7kSE8XviIQHUTe
fTozSt6GaRDwbD1KIyy7DEOjTeWe3gq4HdsxtYaTY5fPnOE/0Wze5uCfMXJppTRY
H9iZavc+3QY7sv9laejt8/HN6AgOrqlQRYkCn2/EN04WehhlBiihxXqgzbp6kc3U
U8PTr7oqXH0Eh/7QgHGI/Rs2wV5Nfn9OwGDoauV3cgPMwml5samDRMCLIk5Jn3Wi
a1wrBvRtzfD1kNPx59+6OSwm2XEhweAbf8J6hWrRfOjAXGy/UzgmSN5uoG7Cg2C8
uP/AcCMHJlBPmNXaUOyTaoVdAcH4MHn08hlE44Uxs6B2clJ5rzWtsPVoSFfh9CJD
3JUYzRZziYcuxgM6o9rIxNHjWZsBRNwmcBMzgoGJw9p3YBXJ2pO+0ND2XcEcbEja
e9ViCBT7sOcaqcVeocvOTLXDwQ2US4cv6IVsCPZ5uNdnTjqirk2EIpZH4Rt+ECMe
EslKWgngWaig2VdULk8M80mNk7okprxsj4rCp+OCvq+lL3Wq8fnGdvIPqxovARMm
5BcuYonpe21hCr04e3jGvLY7mBJ+zeKrPcnECJmq1OEJP5DMl7pUz4zhLxNyxb75
HuvI+IqMsTARTnYhLDD/uoReXLdjC6zszpsJpZwkd5+4Bw8bDqVUkvr1g3JB9pGN
s570jwJdj1rHMzCWjxYJ3ccqg1+5Dsp6mDeV43b+eqPhAsEKbtdjd0RFJ6wmhN2s
rmAQkJRhxd9Z0PMn1srFis/bWcTpgrW0cUvs9WtA3LmM/kiZOG3K/xSYv7bTx8u9
H+YLqv7blKftiDmJhM1Fv1GBnLfjGQi+u3WWe78/jO1srUtzh27JGnP9zxWUmRd4
NWHxkk3Zb18bfX/FtAWfbPn4CSBXI7rlw7FWViRWGMUEdPnh39bpn/hAlJBvpoy1
3QRsQP8DM4l6R3uRxo4K2dBho3QgrSkppaOFvykV8Q31Y31rFDFdk9xC2iM2k1vr
rjTUovwAlhrK4tXogeyp1B35vksPw57Pewt7G5PkIgWsdKXgxYASjqKsavknAZ0t
zq3fK7DDV2g5Q4SQ/BccsMTzfR/h58FP6KRYnqa6Zn/GB4Qjr73e0EcFJ1UuQZos
q/DggUAHMCAxaw2h5AegJEoFNU/n6236XI/nzMM1LGbSLzQOA2eo5zV4jSTrLAAV
Xs1doDGJMUubJursi1KykdMkf2Y5a+Hruuif2bCX0swo8+EcwfAfa5HYQe2wSS75
JgCJ7X8t92xF5Wi5b554cKnhYgYizxDaDt8oKlVBMyiiVzl4QNRN5UVZQiXh8P9o
UL0gKqgrhq/oBnLpaj4nrH+/2kZW2+CWuzI3rDToFnPCExdWXttNH6o3fsB77FEQ
LdFfXrizenLT/QNzYOLDPQLcyoyia3jeUKLGS6FdIxDRWkVxMaqMOfXimMIGFlAl
PyT1C/ezJ4jwIlTgbMQvpq216rI08oGh6GcF2RAqhHfQQi+LSAQnC4r4nXrBEyHa
paCiQM1J6yU2KYafXmMH341BhcRoRVNX371KiJJfzQW83FRm13FS3vanRgysC0Vz
zqw+7A+Yd0iuH2DC1HwBUIn9+6wcCFuX1jXs+N2WJ18d8NSv0tM8w0zQAi0tT0lY
KL8LYaP9IMtCyzlheVXWU8mrGm/AtwrhU7GFJaX5gNRPq7zbAeNrf3eMS3IFbOnE
QsJQ7/cNpv2FuZAJmCbR7ZRBMFMoxSQXLq/1tz+6HMrFByijL5x3IYEHP2bArkLS
ZxHnPUVAPiIDPZRye/ZWq+SF6jU2edw2tDU5YUgt4TGmUq0Kc6LU9It1w2GAlHSe
QAJ/ugxVWxrgVSs3AOkxV1Bfwnv13idi/DeNsJm2/HP3uh0QPGtcMb8pT3yIi/75
7SO5clw3mVlrP0H34pCiSLeFSkKuDDI8bCm+6i8bhX7WjptVcbuia095BgibvJmK
agrwseZ4rGRJsjhOT4DdWcTc8Q4jvNbidxgJnzjrDIrR99LTgwRXFA3UpOfulkCT
FLI1/aVPBXTNhflO7TPWfrqw0Oo3yqrQKGWL9wfbroQdrd9j1nb25EEsj3rpexux
WT8juflrrtVXScvzr2rnhic0BM5FPYlNeZo/kUohoReGB53TFzLp1FtS7B2hvxJq
UWlnysdUc4psksZk06Q+u5uEf36nrjj+0TGbwu16u8Nxm5en2njvZQYmLxYJIKW1
4YfVDTHtGe9znH4GcsqMR2eYEmIqWc1HjrzxktvxVazZOL57q/ubDTpKU+ONQgVA
cY984iP3jFqeQc9WFWF/3cpFE2YMTPJ8PxTjY66HAz5csyIdgM6Y1TJ42Uksn10M
lS8UbaVtC0cQj7MEAZPxxiKoJ372DFCl2O9b4FMN92iXwRPKvt04QtqGcZcCsr/M
n1HfXjmIpLTKesyIJx219/+1uHY9xvJnYOCHimIp6FVMQ5Xexhu1annl/ZmEKs3C
BcSyGq6c3nWDUwgLtm3A1bUpmMEnvMQGsuwaGe9CyBCDWjTOSGnaBkDtZJCbca8M
SSyZrTwfw3c1yH/zeyKKK9EodHYff35Ff/zwQtRrfrSCUrypJz5IZMg0VEN5WcMa
/lYIPDya/rK3S/RxgCbENI7SL63CQ+lfC6kO1HSEDu8X1dw8wSl/9uAMIrVqHkf9
vfzXcwggFkI6ejawHw/cOAURYw1GgqwvfyYIioC115UUSBPeN748Y3tGXl1LhDWa
VSqsL8W0x4vLtMtNiGjpomMdrLzkALHeIJAL1wG5E4D3yXcYmtv5OwoIL7yScpIL
vCRx2rLVAdjthC0qZws+a9NogOjFcQvWLNTQHQaFOdeAd4bwd8hqpMuSxVtkRJ/e
SRj+0NnBRhn3f2L+zShcaQcGjljSXxshvnWBUezB7qbjsw0dyfpzxn/4YSsW22GB
ym4M6QlMbkAjsKwWrGCYKMaEPpSf5OnXw8XlqThIl2fAXzRRnrxGKwVgLrhq9Sxe
e2FuRMlnqQZhbSQuufplbt6F5Ck+b8yaSRoxegWGtfG7OtZjUlQy84lEsGKiKxdG
lsoRwOKFPAqt4vwCYOTRK96U0Gxile+awaizeOotZ9Tu5yaapp7d/eXhwqKODL2Q
TLnIBfHrxTYaQoWKJzRnuBwO5rmUCqYYW2AesjzC1MBkcm74vLWquGXemfO6+l8p
yxlU/APj0SGvZKsSk9TuHDWuwl6rGjZCYUmuCBPsTIrow0ZKZupNOiNDY615kjLY
EaF1wW6Jol0tkstj4jAIPQ55pYMJuMVOAICedf2x22oCoYiboBMZpf6MRIGnOpE8
D3U2YheLYz+OPsGcuYXm2ztRUwY+LUXxMWnvhBl27j8aCbAc9ZJ0nRfl+IDrPYj8
fcNupIMuJGN+YzrShtrupU4jUYb873ug4V0oH/jMh4ZPNl90BzBoHp3oolSGxkVg
BnEYxmu4G7aHFM4SVe8j55zSBdluzgcFZa59wYMdF/7iEFMGZiMOUap0slLrOqjq
HrJohzbaYMd1dQSCoRhGvgxB0diGiv4j+zkGfTdd9vEZz8qZtCJAROv9i/hqPnwn
l9DBzlhO13bpm/wesk0q29+hb31SOryyABUAQMbgs6ls8uV/5c1+WDV4E7ZNvJj9
0yktlBbLiZD7TKGCXP39gPsD9E4QmaUOIETkBnQcer95Gm7jAG90XbaX3POuTads
oGkR5Unq51OIYeMQ0Ve6OJiLCuTQxIMM4V2PzVCQG5Xpdw4ChhTTY3Y8HzXq+uum
FXqQ+Ywg2A1R6sMNnDW5Ohdbw8ZCOBz4q1mU5r8W4YO0T6+MeJpQQimuBp+Aa8KZ
MEWI6bOr0OOtpX/M5qfNctfJD4da/IfqIhHKxgVI4+kFiHX2FH4ZkaswmgfaJ+mW
DzV+q92blijsdSw/QEiAcuoSnq2AM7bfjDnrwBgGb4M7vzuKAh5KYWulN2EN71LL
+T7cMJ3YNPOPqUv9Aazv/jBWkvVrGBU4lN5/aN58ltssTuuAcK0//S8p6E1ocZUh
iDDdsCJWSHynMBt6/+r3/QbWXsxONEkODuL1M0ZL1dTsPQAmiBu4D5dWG53+HDD9
2zQR4+XgZdZI0kjVOy25RDmz2lr6om7n2UkSf+WQYxFtvNyGRVXZRTnJcIzw+uOB
8IeI1sZ6rOknLZJZh7euSSzaYPX6Cgu042mL3xuFUxmLxLVHlGruKNEtLzxAwiZ7
cxEtPe9SPHUyrwhwZl/UlLfsuU5b7Z3zRs8myoKEFW0BXrNj/PL++Y4a3gCd1WR/
yT2lkNZa559BcN5tE8Xxis9qRhfB+qR3vjaCyDQ5eKNH0lAu3W3x2IcKTRAf67Y3
zBrZImCYb7JQOAoFIDLMnXotSr38wvW5efpsySgUzC99R39xp5Gr6aUmXH7KgVXl
vtahcaUIX0Q4WsIWz4OrZlpEBRQlCBpEN1D80lTq6qu1QD5KjQ7Lzw9XHGvSO2Bc
Ts7MYcJBsXky7dJK3XHZ/pqS0O4lWbW39LtNHeo1eMSYvUgW+D6IL0mhbERcrahT
odYAJIyx5+BwM4sIE6JULd4vlRNonApcqYdl/toXQusWiS2+Bs5/SKjirvv6aicQ
6peW2UMhg4xyirPkQ8l+kCaP1PyFQfHLe9dWmVSzgsw7286MCTj1xXEX1uqNAR3X
qMvWazAfXnfS1VoNkCdxIdgG4hZSgceGtZmPN2xepymiTSSWEfRmjTfurbn0VQLd
t3stRVf4vlB7YHUKYSp/PnoASOV6tzp8Xf1GI8WRgejDsxZKmwMabgiKcOMO3UsQ
i3TezS1LntSI0waoXC5qcP2rXeZC8aDCK9t/Juap5JrEVwWXjev4ADCooz81hrEc
GCwr3Zs11d+EAxNHawh5G/WuMKvQqIGxcP4+RI6G/rQcqBFCDbmMnc8kjYIwepSn
kfdrRnie1aSyyLSfXiEQjBMYNXn1/qkpq8YxzS0sCZBHelocL8Z/jRj1kouV/MTn
9QqiPzVNZejK17a5g6/EJAFWGkaag6gZa1pP405ORi+iQk+MgaAsInBktwNff8w1
25j4j3fb1ZWDpMYqrKPpyZVzfo8El5QsWxbo3Adtty98ZQkUzAYN1IfNxqjLjNeO
/rddmx2y/bYZ9tF3i5eRAtJwk5+X9Pm45rlp/wTnBZYYmrR+u2SCzG4udVHvfxyL
9YGz4pMgHDQLciCMRT9fMzMD23S2Mee0zGsWVaJraSrDx8P26gOaH2KqnVfY8VJ5
6Zh0pOQNxe8xtinLLETO66DIVASyxb2Z96+9h/JrfK+G2xZR11wo2QaBDg50EhUR
vMXuTJJeCE4D2frV/yWjCiBQHsPM4qzD4sr9dy4VIDrfxIOVonLOgo6v10Nv6lyw
/L13Yw34ZH0ErpyWEVQHbgG7ksvLvoMTVHhIxMFuNErY/U8sfeBBwrwZG5xvY1ej
dbyDq1k6HSEEs0GMN9PBYlUiDmVISx6DXbeGhxw6Y2MXD7tgGOK087pDUoioWoPg
EDdrzELwwh01FKvl+HV3Qmrtk/5LZU2yvwas38VQZDnJxxI/BKjTtm1Jsbg56Cjq
wYClEd2Zl2frDTVjCXLtNROWEnWbnT0d+QLBybgvZNMs7CarknqhwwbijNNkeBm6
KkOkXETFXHpUvOV5RoyVBm+qwNn95mU3JcQdc/mUMJ2XMzaFrwP3EyeNoK44DikZ
x1EgvIf69ZwhK1Tr/dml4hD3BBuuNc5ZlsA2iM+J5JM/1kyWZQo9tnIfZo0ZONSA
Uuv0o4QvTuLm1x6klUrTO7z5tvJ6dFogaRtf3Q5mVWXa3shM99hX6KFBqEe6wb2O
W+M4VH9VGO74RO76yLidM8q5Pfw3IG1+WpmBIlZHtub2Qb7A3V5VmPq8n2umIb7P
sT6Pig0f0RORezzaSM/ND2+pAC+rUH7+AB6vO1EhjA3Z180CsJRmZAp8ufYNhrUW
ia2l86wX/0I7bLDBvgcqa8cCERL0YgsDbSrDZ46QYOtD6Eg1164ksQmzUM/3svlU
mQobFAh6M+R+zont2Qlp27LUbDYk1QO/uIghWnA3xxtH4kK+Y6kVRl5bzZqYdiPK
poZKac1rKtpNt6/uLA0s7XBCWNtWLFZ64gIsGRiKMMU7rvApaEjow23BhJsErV5p
qO6Wg2PbSxAGaDqxwp1xw7s/RVTj89anWVXV6M1hRdCl2PHmEUOIfFGgktFRon7c
u0qEFgo+0p7tKULZh4IolFO3u9xDs57iNkbmZg1hrmCG6BfreN7pWZOGC0S/sb9x
q0p0xX5hxW32fdO+SpFoexOjJ6luXpSwjq0LpOUyOFWUCyvR4jLx9dlAsKsT1Ij3
FPhga3V7zubl5chdshPs4f+QZstJNu3rlir9AZmY8K1FqWzsvosXgG2/KFlZOcYp
dcS1oM7spjXqVW1hoVy6GbmI+Q8GhgUfZi4woGeWWQ2I+RlygzJ3dgbyTGvQ0dbF
CEjCWFhDCeJIGjfHGZnhLC3OOkIkD7/4jgxGwNumfCibCg410RBEC8efzCqLRRJA
IBYmco3dqDn9PTzE+c9/lTyrQBYLTBmul9XNxaHILP1tRhBr9h4NEghngjHWjKRm
pG8n3QJHk9utwczW5WXRvCK/Eh5bda34AsXH9GwrQHCsDaf1voCNO7TtFUwZqVFM
ZhBe9+Y6JAMZZBgn2UhfMyrkSuXuF3ygSiX1ctBBn0yXvUgKIF/k1bPdKfQp1x3y
CrRpAr7rhwGYrQewGYh4igPRsQB9nMG4kAP+sVCvRWv1AVNd5TuYV150B51F1U79
nlJxIARl6R/euAmLIgF6DoG2lz9WgWWC0BznP2Tlga+yUpeYRLt6XuWyZ3fJA/Gv
NbkQ8YVDq3zqdKsDVxEkvTYMcQ0hA6yvkm/dpqszALP5ZSsTVFxhBq0VFoUm/NyK
5jDxR1SbYTvuSYafCky/OK4W4YrOU7HvakYvugHnjDLmD/t/1ZWzLbJpHETGRD/z
vAHSGOAzsYTlXQtlZQeb5+Auiw6E9RcxmUFDHaZGcHk7JatXt8PaFOi0t1xKzuos
OD/Y0+QWlMkSGQ5z+dpEPuCHh1VDug6TD/1CkGwwa0S01fg0hOeSt6+4GRa4joLR
IiDdSZrQONpLDeAAdLVpI4u7XZlLuyJ47PXSlfg3DNlbjEUTY0KMFgIntEaBbvwf
bEwUS8RYtVbP7hFGHABfAayb39U/ri6FwtiO/9t7rHU1wumb5DWBGdODeHa5eQht
1bKNYHp+nZXLuRpnl2+ioqkg1h6qXo0Q2HE00vklyRrxpLkveKhERIm2n88BKD5s
xvNfBPXKManfOWOIY1FDMoXTsPlobmIWRP+g5uXuqpF9FvrYWa+dH2WjLWLHHPtr
53ZMdYRmQA/iG7B5ITB2071zNl8GOQKaa5IkMTFGxyrQNLdn+hkX4DVT36XeIcZQ
Xf01T0H06VvmkeAf4sJxzb0J1PUO/X9E5/+vz57Z80t7BkLUtwXFsxb0vrHd7dGn
4TMs1iGQe9a9Hgd2jLvc6exFRXIgVzryTNTIrsLz99ZD79lu1L6PRuVDNhh1j5Z6
xweVamN9Icmr/2QUIVbzJnbjdz0BlFlMOM0z0QxMbsclHWnSDRbgG1P6ED1D9ioJ
67ID3ji7ukuNnwPYiYpuKgsfEwHFiijF5G3dY/wn8b/pDe5Zrp8qmX9f+ZE6qG3Z
68rCytiCUL/7pFK4fbFxetT1SrOY2YP4xifwrVOSRmpF9ISk4yK2oXlONnW/tO3j
TgbkMSVHQiJFjiOTJbE5j1ZjoOqR+dYnHVcT0cpCaxWUrBoUIKWN4wIshWHDY0zW
bpfiiPXTgbnytuYaJN8elnft7DTTFNI2fubPmFzeSZMknpfmPNM9lr/GIk3JrfWQ
WaPPBhcwl7TlaSfvPQQXgQrjYT2HGsJkijsvZYvT/S7I9SYQOkj6KQSkQ2Xjppbu
sEJ0fr5iRLvX9wGPFmt1sJu/Sbr/Bk4ac+hm3kPy8PaalIEpXhYXsh3hnzGIbNB4
NQS/sYoE/2fEzMRKfd8AjzrQi4FrhtKU5Ne5i+yg3Z1MpDzJArFa6XyP0o3KibzN
qXcvCNDz3ScS76zHa5DqyI0y251vArM+irA3mnHni3fnHEnp1sDyligIM6sWsCHl
Br7RiZUEK4vOxfUnLieN57aZB+3BB8WH53TVmf0XrhDnzSD3QX1LFBOCCJh1oNwK
AEPlQDGN29qhtLO/ptbjQ4I1BLn/HlAZjj04WjTc46KAwYjCu15r9nk0v4NLeMlK
j6mx9iQjt9+6BDIRFuZUW5Trdp/J/nwVsUQknenPmdAIRiz96xGJ+9eNvZay9crr
NAy98GLThzwl5GaevLitaKWoD5x8ZIjZtyvgainmiO3bO5/o454yox/gFu6hBEvw
KySKSv2AiwbxjD8Zu9wkOakCwHVVXwKDSWxTjmeMcXuvFLHYCrrnP8sGk1z6cDpc
CVL7Hir9MpO2UQ7s9tT2Y2Y4sLrcn9QzS+yhip4GGGWOQb8HluKJdHgwBsqgd7iC
P+BqZvuC1FrnJnH/yMOYfuMhbVSJw+MXdAhy2zEP5dJw4Zqv3bOz7V+MUEQH80Dw
taYYDu7dyuoStuqGu85eF/fJmkhN0QR/Po5AmPRZ09kwUSLbjlRRXX6gsMIAEe5c
i2Sfcjw9NhZB7nvOnmrf6vrdbTQfmdWwFLmiMV/rpZDFqYrfr/AzYxEpw0AP2EfD
77QAPvakna5tWI/FlBkQBIfgYRtmwqyTPFmD1RhyKstCEf2G9SFeMjtmD68JNahn
EVzD0he+YALijecCfrjixhqgLlL6qB42v767mVnUWKxWuA6aw3JfsDfrcwohVSbp
USCGGDlBWYepjkTrVaob7Akz8jdIScL1jv/MJDEqEQawL0mBkIDoqSEF2M6JrT26
V6vsWo0jVxXjJVo+ObAYs7jxAoUWE1eqJ3WpZZ2a5fIDaUUWYtoJt307hFQsNguG
UQioT1PDX91Y9ZX/1IS0L11r2Ptw1+jNGbV4tbYMQpSYMI4rfnhyZhTYdLzqjlVU
HAbkGRMoD4ZPHaT3msfznxwwecJmHMCHnucoNRtJTHUIMHTsNVDwlA9AGxXnnzWS
SrpruysHgYk5SjK3BEqLbtb49dNA9gxw14Mq9CvxvFS6GQzsP+R2316gDQvCBEXS
fgD+aTRJfUVOCDm6P6TetDhD/UeOGmgOz6LEr4lLhlMz834PTR0hDGKMxNTnu4Qe
AyDIYnQuL4PfgwJvfEtCSB/mazTFjgYaza+FN5GFGTzAAxqmq2HFWCrjVyHyY1QE
QOGKC3QpDXELKwD2acL6XQF/rwWjgxYaDJOTsZUWkkyZIYTJi/hVsP/1lNqEzV31
MLeX/11U7USmAYHmQeVZSIMBSBTU5Epo2Wz8x08WgD8DRtYpvuDux0uV7kdER6jH
QpIrvYE56Ya0RPUX7BuCbpNrE/gPxoKbPuHSGwKmNRWra90TlOS+bHfbdPqsTYBc
Vi3uBztXwu3OhJY/cKRyX7+H4k/Nf2drBEsyRPC2WZNzrEV9+uCllLKcxjRsklWY
hldtEFJY1OghU+YcmXfb9rLvAeW3xUGBW6YJPeVagFWnXoPdG1Ej2yLwcgmqi2cz
1XRf8ZNt75V8MZpb4Ut+yyqx0Vsd/JNqvxW9AaoXoOlTAQwVXA7uzpYPYZR3NKSW
TEs2niM3E/Fq02jONk/4FvsOrMAzIHD8gPUZ7isthnJY+DFBed+bo4bjbJlST83s
+OkA+4ua1eXdVHaRowTx1Ko4jwBrMkpkGH2MiuZuPLtBuJy4u6ZdrX6lyVYshlW6
i7oHuzSNxzgAu4ahiy7tSd0sh1VY2xgSRiN0l+Tkq+vAQTYKyv841gJReq7SUbSr
pgZ3uhQ7tp7Ugbk5UrchrVdWUIIKZoPQgVhge5vPceyYPSNMlM707L4r6K/iK/UB
Mfwu910QDn5heBLoiz/ogWaxgCxvqOCD/bk8cUq84hBPfL4KmUnkwpGAhsYVtZYp
wD/n+/GrBOcJhDYGRxDPVdtNeFtqWoaPqLOBhweyH6nSf/QbgK9luNSwGOEFVjsj
6uffoyXpFLcuTGs+Zbm4e9uLkAkMQ0T9GZPb6zw8g0x5unGHaOfRORxStc+/wqVL
wqa9kcIBAacm2+04Gtis99VKAsppTOazGjiXqhPQq9bqJBo5+ZQsHLVWmsn88lUV
ChMfa+yef81qY2cbW0Bvm+XEE23Euw9iUDrpK+j/sL1+rO/xSecBMFgadwEojBYB
GfDKg5Pum3/7BDqvsjbld6SJ0baMC/Eq0T26wT62g3UqW2xFPiR0Vyd/YTGv/cYA
ROxWD94lwMCqNpKMnH1K2R9W4s5iuOthQH7OutfMrCOIoOGNYEQS1XhuVAFjBuFK
BDeiUqStF75b7ZM6Hy+oxZ5a8l6Fj4pFNfN8qF0kkCXqQePq2KyFQotTPvUhPpgx
XHsdp2sulKnpFbKxM7L46gjGk0rLB+V45t7BL5X+lXCEtXbxV6kppDTrlQ1JNY30
E86HOxCtImyS49JH1hs6DaTlPB+InGgLGnzcvsNoWNPbwVXh52gkH8i5fmchEYSn
V8vw1u1fcPGFJdLGN8JnhhgPPxZC8bmttokUvMVfXvtAmznfTURfRUKcj6+3128o
AbFfx35GvC2nFVIBOB4e542fX+i24f8cwrbHKmGhBC7IAaVunHBqCyYCxa7zS7/6
ElVSboT/MzPs1SFmnsAG1W5u12odcXvelzHYB+8QAJgo78pqANabe5GAwn0uiPrY
AHqKd3hR5K+KRAzbY4D4+eeVHckjw05Fwz16K9Kt2v5EqqE2P34jYo+b7qxDXL4o
iQcIa5co9+RaujQlRNfu2TRhlmXQjN8TNJ9p2JR08onRwFr10diOhC41kAtpOqWc
oXcxNyoaPIQgTlTc9xFTzVpUQMYR++U/kZtzRZw9wC2m6ZeWmUzWHZ6n3JTEr5Rm
1vjfmpyGohs7ubWmYzDcH3B5vYEnu7QdewD438qJsasQ0viuf5IzC7mz0HWnenXB
J/zwxXTXUQbDPZqUxpz6NNsMaN/cPd3ac/VpLdbZOzOjJB1RjcRGniDaDxevOyA7
KVetA5EDa/4xYlVouAWj1O6zGahgovP4aRLiVdiwxZmHD6lMis978OdBH8BFHQwA
oory72MM+ir2k7H7i7QPnCLU4BiMyBaqi/qQPNoQpMYVNROBEShu5F9mZUXlsDuF
7pr5ksJtW1aGM1wvcVMGochezPIHx9Eir8YgkVwgkdPP09gOtKMC8CiRnZ2xU/1c
8Fp3AA0SeANz9ixOx3ZKpqASeImReuA/r+MXPDjDZk0A7sCI53JV+QcD4NeQiQz4
Nyu9EKrKTrS3PmDwWe6dFyAqjRkY+svq/IRLJjTZMX2pKYFKjuIEEz1ILCZIwTvO
InA6Bb+V+patZeMdLeNhVcxdRZNCiVJvJMZTSrqIcmvqavmlHbq+/LloB+oVKX3n
D+8xQyh6FmdC1w0pFbSs+LOmhL5ElGvJrcpgRHk2X8IHzpQoB0ZtCL1v+tN29uYk
nwv2LiUHGuPM5tP/taVrB6+bHlnga6ZrQh86WnVYA7OdYi1NXcezQdg+ENLk+4XI
dUvRIsQPG5jeTh2ATkf15OZSsphr+fq4TIDgsg53U0tLjMP2QgiZ9oeZlTlfBOJa
ygMAit81oOgr/I4FsNJRLylr86XB6LStkkFKthAcTLsObjqCUCKZOEplNsSndcxK
/TA7PRni0j0RXVotXgbyV/634wv6RM8Rb1/b1+xkUq2CfbHfbHSOcCUYgAuJgVbF
beP3/HmuQz1Bx4se+9lq01RP6yRIaOWNsMI9uVMpTwSI7hRM+S31yDsGNJ9JEYgW
mYcJt96PC2+4YINk7mPs//VzQqsgjTTB1D/B0PZk0ietHsc4g0akXO3TtvFwunES
IT0sgbAqH2SLsU86drAWAKWXFYMpybS31ucxeSuUn39kTbQ+nZ8ZZGwjd+qC+G2X
nSIhzKzmdnqo9Ch3UBQCTTF7jbr6Uca/t69eur5tlPc9yLCC9dVDiIhRqZR7RoBO
5/L0MwvwgXaiTpqLGudNs6VwTYWvs47JTahvHPqtM/d4pCfaBMK3swxYjL202wq9
x/ZNIt/6GClzxSqaZladqDbfkYExABXBhvsOUgt0IgRTILTObTs9V5wrNcYdW/R0
CyUEmKgqXt/JWLIg7QXF60zq3ux6uHclOiADy4+kE5mtXlkAeZMx/phl9u8TlnH7
XhJ5obXQ1QYGFp/2k5bgWqsHnVxcEmv/x+6pfhRXHrCVA1fnWeDHwdbBhaBlkUrP
7tsZ+qIsL8jmtMp6n6NiQOmhjp45Yld2Q24ODPT38CQLrR6wVc5jLb1nhOfbFL8H
0edyi2zlWShQhDNtwwLbfKS6XZ+U0ate5b7dA24f2NStCEeT82VovWyy/KgnFfh1
VHzlqQTZqmR19X8ORuzzvjnbOIj6kBTLtFhFIoJJC5sWu4hpmZDPCWRma3DWZfOx
7pmPi1gqZ8Nv1m2CjG74FfkvdeaYRGCIJ4Jb/0Qyo9/Kz7EXSRG0w7ci2JKeTBzo
QRnbxyk5flC7ZaG8icB3V+B7VS0vyRPc7tLHEEG2l6wPlfZ/K3s/tED2EB1FcyYW
/aB3zUQB50+SS9Z6780Mhy+qn+imlp5b4okd8hcAfqhi6J0SYXmKV1AzB0gREDDA
uizaGqNE6FZ+fYEkogbnspGIZ+5pTbU9ji3cWuOBMeVh1a4hzHBzwyp/7m3JYWd+
7i+xSeSr4bVysF9GFiXubreUj8l1+BLeS0DpHcAhxlkv7pMDE2vGX7Ve0hJbduaN
O0rtuiIzzH5okHFEnBwpIKzxTGlNkOmchT8pcK4lufpvj03xjNjJRQsYshvxWc4r
ffH+bPtu7gUjv0HdZa/q/7lK7tsUqwnLfGm0GDSMEVCJSvml12ReL7RDZWrUIqyQ
2vrWppa/Xg1H3yBPXW2+1GiWb441h+EmbVAuFEDQEHq7F6n0xc/BdHWphFWum8Qc
ekml36ffhfZ9dIJ4yu1YTAHoDX4gYIQUhVPJQrEXH14f+BF7pXpj2lSo8kr6SU0a
vnOJSiCdQwWZveQymXtGypJNS1ibJXdjoktpKsyrwblnlTZ9KNJDJZhxQ6Qb6oId
zfdKoe+Xsap3Vufzt/R3DgOjtKVCSbhKl6OXHi7P+j6sGDmv9AVMQfRO4RXn4A7c
TKhlc07P8IY6yRHUjETwAUzhz/YhbgCw3js5Mx79mC1M9x2gOGhxJIl02lKeySqu
w1bMO0VvjZfeMhWZJxh6naW8p8DX2/Zh6zECHjW372hvIpAao8iZJLM437TKVEgI
cLm4UyZFbyacd7/dJVKEpNf99ohmj0EifS4VNiapYUdwwrlhWiTVjxjO7OO48G2E
QFJ4ma/pD4q5pwur3MLM1NkGxULD6eYR7Xhl8LN6AjSKqwya3ajXNkf4GtftQcCd
8gXj96CrXY1KWjlcy58Y9YhspILyyZlPtV+8kItnbpBs3NLNBKelBY78DtK6rMlZ
494ykV3UtkLcqoUnHZ+YDTZo9UmjTKvxLWrCcpcHWOcqOUFk1EQIW/cBB06KrATe
4GNChAk9EWHRZcjTSKSjJwzq5XaBTURvlM02aVsEI+88Lk8pixvxwyq3if+XngVB
yuLdUNSqr/lMgVEqYg/30J9mQGemjtyUSoScV6IJ+Z+8TJWFrR0uMiJCtB2Unl7i
oAeOyDQNim5h5W5tk6K+H6FJXfHwnqAv5NvLCCRUKp5lkHWKl2Uwliphbf7HB0dX
CZDlavjo4ilStpjJVzVgGE3fR+Uz8L6sg6I3SLbFT+l67yHmkY3aEe6BVxp6Jy+E
rCn2bYSPDdPPCB+io2LKxM7OJtbqdf8NMKTjeYDS2Rs2n7JpKlEQLOKfC5lArVu8
uWXtSQHN4MO6dM+fuie2QPB4WooeulseKWH5dlK2R8batO4MgzHrEqdDJVjNE3qe
ir5I/Fmql2Oeeg9mv3gijrncRoHuNJC454CWKKl2S/8+uGPyp44NEQlhrA8Y/pIy
DmbLnQyQRI43viUB0HQJWficIVD+Y+4VOz/Soa3pHh9d0SGS3x/9noohjqkcSnyl
YjhVlpigw3rkHIkSB7wSLYgb7Y7gzlnxO3rZn6cir/9V09V9r+PoueI98344m9ir
UTci9aHdIVGSSut9jXTReUH6fh9uO9353uxg1WTz81mX7vnlvAbkqP5n2GjNdpMo
yi+3ECRGhBICnhfeJ0ZqK49F6xh/PSt9+9w4PUS+qbimPAsveI01RKy+DaBCy65j
hd6jJYEKE3ByqXXrvQmz1g6ce5gF+Q/2kpziENfidqzxdByyG8HvEQA/GS4Mj1OV
nV+5Cvh+nhvjD/f19MqIsSRCMdKL8ZXa9anKtWK3AEMCxEwPKZ6DjLLLMS/t9m1K
XRJQ9AC8Ro2QPgruIDayogmu9eo0t0EgLQgejFJ1aTlAs+QSMPLkBMGYbQhnVNwk
x7auFAI7doqsJjssc0cTwaj6gpjSEEYVTctMPQU0UWTOjVZCoP6pzXQsujseKY1v
dhh+ZFt+WArtgSKIi/PUsAo/beru/ebHwaX2LnnfLxGUwuIzqyE8gesjeMCejy6/
2BahLq6nMbR7zO35Jw2M1j1QHeBreyuaJDwGHj/OXswAH3dun8ju904uj1nPRs7T
KEBTZJQeVU0q6Aq0gKE35zmBXLaRdD19d9XPGAliH/4pU/sJzTOM/vD1VCude6Pk
LLchSB9pel6lWju5Kyj/SLVHHoc/s5So7YbZpVuWSp4mkulLh7lK1tOvcIaXYKFe
KtTMK7qWtEUoHoPrwiFme/wnba955Rg+oNN6Z8X/SoBhBeG8jk1/XAOtES3BtxgJ
IT/JmgP1+LZu7JMofHO6L1xThiyXDTgun4RdIq7dy3LAtJ5cdvdaxvSEur+XV6Mi
m7tycATSh+IqYr0aEC7B5BC8jVMkvdA+jIuu1SHGDWshuRskhYKI9XylPGH7O0U/
cjzF98H5FQBdl9g6wPaInMBdZmlDsovqHniSUgWUoVvymHkfr2IVH6A1z+T7h+Sp
l8r0sUcxKsL4vtGwxRq/l3bW656j9L4eDhx4ojtgFuKwaN3qpgw4iKr166KuzOYm
IrbYWBRW6oq3yNb9gFMaIH/rrU3Et0q1nPqJhxaNpNp/bSxkLMURTlb+UDsdLnF+
6KswAL/G+lGEBiW7ZT1C4Uj0V/DlRpFH84qDE8LZI4Vyn2lh4x0XN1xeBRt8jPT8
ZaUlLoqDDQcmFpLY91THNMT4Q6TgRloIbEaF02U0sT0P8jetdZ8WEB/ZXIqB4qFe
O1gIFqQUicl8UbPIlAYhVw/ILbE7F61Uq5qhMZpc6/Gp1EuyP1slXvlW2zJdnJe4
EjkG9o7LmLZz/H9871wOgRwG+O+xssTPh5r2MiKz/yNLc5LZZ9tW5UDU9Gf/uYwC
7rEmezOhINaOrFvwf4a9ggl89T+RxDwTUOb+YOQvpzt0ABvlPaBeW8QegvBCsCa7
4+Jmx7RKSfkUvgMtzlRqeT1B6dVbUW2seoP8a6zTPDC3cKDHqmZmFGwY+DMQxi5o
anXsrwSsaTKq3bBDdLoklgpz+LpeB2qQ4pJH/LKcrAHbutMV+WpoljIWV9/DhQ2P
FiBY90WY0ftMrJ9tVgZpk9DHQrYR+Bf5fbtLkeDHVSfYi/5AyfLf5FqOQ9DgtA+4
Uxau+9Y5pEQ9xFMDjCah2nDXWwU1M01Pws9bdzaPcUW+awciPB0HG0+4pULVJ4af
/BY1gzQMrwEkyFsla5/kfgmhbKWu/pyBHE2x6kDrYsSNjNo6ZuEM6xH1eWCJOqv2
oNHKRc7wns3OzjzeWoaCRIeLmgEjGOSfgkPT1T3sLkl0mqTX6eXV6AuGuDlrz9eO
RC/BCi1Hre+H57tJbLCsGl9lzFe8+KoQdetyzQeRikGddofLInYqE3/4e11g2ktM
hNJ/ciSr3C/OKPgEVZRkJyk6rjj2IsYpoq74UUWTStI4ioX0ncvjBDpVeEbJUyLH
du3+RjOd/nL8GNbr//uRTgrNfeAB6LcBiU310pfEfydVY49FjWeqfNxXaj/ojU3y
QXdQ20v7YiLcPr//A7UUxPMHWA1EB4H0qVfLMGD1+loBBwooQ6dc6ZME/fTBbZ48
38tcT5CFYrElmibt9Iw1n7hGS6x71h/ZFZdLXfUpRZbhLyu05HsUTskSF4C/4SF5
UQzyaisM3di2Wk+iKhN765xvwUFfsK+SGLPm/gypjYOJ7m4Y7D4WGNG/izRw3b93
Td6RCUuA0NbeyxeP/GGTQxjWJ/gFJM9Os9PwFDOI3hKBR8F1/RBXR3scL+vyrEKD
Eek3uG/xwC5+gNkOpNrEq/X7ZX6D9NLzRk3X/Q7yo6Xdp0B5sRTPKmd2YVMO8c6x
WSFAnwAvlSIWFhsUq6UqmVc+rQhmWiTCN/kXDAzhrbI6RMioJUleUjbZT9VoCr3J
G052eb5A9WMkDn1Hz3w380UmAL6pJZ8TJb0kWJNZBWEtUqrXPIh28ik9rqkdCNP/
C6oa4G7EdPzVncR50DUcZElvmcAgoJWm48K4gcjqaqy46IXirNBUE5PGlJD6FRq/
K0vBS9eZ/ihhB8FfyL/IE1byN3gKW+Thtb4vzuiOowyCSpwuoyzpOhU/y81cWdiG
b3sAp1/+cdet5tCWJZ6X6zVuVVfAj69XJhGR2Za5NFYT2TjGGSde18Z9QIJEZGLQ
JMtMK0WK5+cUeQYHFJ+VuIgjQmQ/dGebb1jHln+qYN4GFa/ZfjF6P6b71SobERJV
SE1YJToh/HLQqDnNfFPNWIwxN4AjNyhCGauLVHrseu/LT4TEJn3KQlhK8RdsaQpQ
TOAcAo48B3bsSioxwR6inKYbLcRI6DZkTmF06KTaFx78IwC5zYBA4LuC/feVXIUP
sAqLrH6Um62s1PVaXv4zKVBBecFL4tXG2LykeqhhEiA8apIw9IB+hv+Gp9gLOfDR
0K0TcGeevjZousNorsqiq7OGgCYrtQoHpz7uh13jCMQP/DZ/WrvJgdmzcofae876
S3tWDtY0Q1quomrhIMI1SVnVeu7p8nAXW9l5dWqYx4tjPbIDeRgObNRfpq15c9Oq
elQ6jlQs8NUBioGk+xpm9+F+Fb06mXupEWy52IY8flUkuNiiexgCodmrjW1jtRXk
axRPIjvQaVoXPqehUU1kzRuea3J/uBTzSFsjzVNtX00zl6KaW+8uqrjVgha5vw/r
nCg27QSdmy2NF7D7SOxGX2Na+8Rg67MaX+qpCkkZ4KxwoU8etbvBOL0Hqj3SXvnH
ufnfEpDfnN9HP+04yViwshYxeIuBV7m07/Skw+aHIh7UbIDdcPfYt0r+b78ujw/a
fMphT7osLdFbY+0Jdg/HcJ0++aJ2ciRPf4oP50q21QFcEJ5iHeWP3fy1XvXsGei9
XISo0iVBO3q6WUjyqPBDoiaV82Y9DmB0p3YHZz5CeCQ02UCYFMlOjyA2hvmIm2xq
rjLtVF6dPyg1p4uUx5tsvHAATjP5EodwSEWEHEA/SfqO/ZHb21hulHGWAOPhcdK2
bLKWQ9n78WIetf+KFccuAFRdxJbenoLIUY5GxFVVuQJ6s8fZB1LHL3LEssD355zE
7njaydYmVrzyWUTSzMr5M+dUH1DkDIw0y2RsLmTb7M1kPqGK7UaBIkveRY/I3+M8
jGbe8siEkO19LKL6pFEcJIoQlJkOqMlLlPzb0XKlsq0lmE1WYyJkm3dhFHE/GiF9
G6qJ25qxnRmhjlOA54ULQcjanDeNtpEOKaFsFcP+SAgw4h827mnyIWLz+zQHYf13
G7slryWHuP32Esl+Uj4ccrlQWPjK0yzTpbEDC9BcKy77b2khcLVIL8ze5TOnZtpV
w9MTbbMlzwPlefqnbejdLMG3jQ5NTEGaLg4Dk0/UGX3UTINcwMi71KP8g0iEU3Bk
dJz7ZjQnMTDZsuBAGEmVPKgAd+B2aSE2mWUitwIFHXWsh3NZuh9JJjCksBg/sW7f
DBcbXJKI/e74rYAvcPmjuEZ9sUV6MzQNrjFEJhKcSHNVWzmDU2zBlNL/kZ/JlCid
i6UK4NJJKxRYj1qUktccv6p1vJ4CbNmQZzEHUp/CATTxy0nAbxr0zEYpf2ATvDA8
tF93DquThQAkUI8sVXIsi+nmJCLcJS+863BWu84wevwYTYdVWKHkhNKzLEBouWkE
A3T3F1Sratdv1LnFJzd4ehtc6bqtkuEEVxhVflMca8RuYAGAo/07/NBX60O1TeWx
wIx5r1WaN2YWMSrnF8LHYIX5+NswWLUa60oqTFOSaXkOW2P4xPk7T45F2cidOydF
s7A0nUbAB/dP6rpwLAI7Bc73tfcXb/QO31e9Rrhx6Li/4T5bv0hTkv8ewENtDOhL
D676FvKAnR6NbIEV+lKeXlXyjzjFVmudc63+5jlkwI5YAguah+XgZAKZV5AJ/uu4
SEcTOUIY4xZd6oAywgiahIYA2X8vUuTwKx2pv6VhAz05z7UxFhglljTvq9Reubmu
tepFBTCoJyiGXLdj55mQ9cKukStfLtTC5Cgwg8iplKpjmBx701onP7ljfSI6l1fA
zRiedY6gmzwG+CDoV5PoNtpDwaNIjpCA9V9Hblnyhx0+GtKFLQ4hUTQPK48bGHpB
/EueLJWWoijKcOpKer+lN/EnVxFYKRQLNSq+Y5wG34g9ETKV65nDJuEXt9S7SmS3
9h3YJdYnZGxDOCfaX8b9bX4T0KDJ8GZ26E5rJR2aVmdpwhCDIkYP1DHdhDaAVx8B
70mpRYdsVjGDOURGBbfdCytVoCzuWKWuEJlIjr5WpbLy6s5bdzoi2/0FFVmzOg1d
1c+i9be4V8p3n/MTZVGLzK/VMXLWdN2SBBUtbunrGvuGaPodaZHhmelvRzZbGwBU
08yEumEP30EGg/vUCizX/vsCKRAv+56kD8xRTcsA6heAcaCfM3hlXF2fh22Xj16R
gW6onDzIaamWQGtqTw2JmnsdSGVyqqn9U3fM9uAxEYzdLBX70PQfn1n2/+HENBUC
oYqdocgc4GtmhsGuAkkKEQzUU9OGUE/fXGXSADNcP6XRvUEJIA7licV2sJEBNc66
D+2I+fMXsPqoVhc/mselaRipv2ERhK8fAO9DgH9BveBgPr4dp9Au2pXRy8g+Y+XP
3ZHcsDtkGIzXXSVwTLQZ6b2evJQIJtUJjM+JTrOZLoBHPW/F6Si7VHFuHrOX9ss7
ISgzWNHIX1eUszeMTZfe9MAXLlbRYVtrzq6AivDFKOO63/1PV7jZTNT3YO4hG0VQ
y5YRK02jw2iUqYdWblu3ncRj6I9rOxQlEycW8iWx4j1QEzN7I7cHUVzgXYmj6Zih
J0IEh2O0i6KfVtyJgRLGMyxrzipkfEQIVI45a6umISF+YuT9AR4zyx6atF2ph2zf
39e/Miy8W+RlHcnsCFy4kqA4jylxS/D/KISdziMSrJ+m80Ol7th3Kk+YM9uQy6HH
tn9SHVo6wEiJOmV/5fITKw4rMGAwt5QdPaAL6IpV3MXzj7t8LChScNUafCnx+x1y
SpUu7wjbCsaGd67ESCl+J3yEprl+4RQm1I/QqPucSdvwDJTxBTKxp1UjC2EbjmKr
22OOzMVM3EEKiiCM1z8fa1QR/PGbCBqP2lnA+6abeyIfa51kBryXEpEQ8ovyfaR+
H8OV0QZKJuz7jMi3uLpwPK8J/lPI3BosLwJSU6g3QZBqyMhwqynbKsm5e9qvhIxI
Z9AbA3a105rDuYFz/dXwR9+YYWNNIi7T5mcPieCiBEn1+nMc/RrG7vFAvkpJ+K1L
6tL8n9U5rjJUQ1ABUyD1fF9nhciBgE/ZYwwddSnyo6J3qnFaaPxETOQApTYFEJ8U
lMdUd63xaOmaL5HYtJE3txYTgw13RiURQrtlXckN50He15gXJq10EjSaTWMbZY3f
H9GN6lowqnr8zcWpjAfUcGZkck49tx5XxLccY/7ysOGEbJ/fVeymvwnZ8FjhiaIE
f61wlYtUbV8vZPlQ+GSz4vYKGJxj4Vle3HU4y/zVEgM6+yeqAhTAg8Z4aPtwdvLH
vmCAqKwFUgVBPlrfb2TKxi+2qY4mVQ9g9s2Uhzw/TMDYgPQ4w1LLatu/5guZbljB
Rc5hEarwi+HBtSjbJlduBBD4ZREFT/oCQtyf7+N8UvtEhZVwgKlAEwq4p+U/BYNI
TB6rEzM2vBiIqnDRLnSREtZWZRoVClcFupsakp41efkuqQ+Es8plH2tgr7zFVz4s
/cgZPhBS2G/zKdfNzDwEI6RbFvi+3dwYYo4h6Tu9yYxB0eAxzMQ9dFcwsxA1A+w+
2MSI9VBraWpzeoZHWbxoaw8qsLV7p92anY1kCE5AisTqhbE/QOix47uyo0SrXKIm
J5N091oj4hUTjpUNwTC3FN7EDvWM3ngzNMuY8+mLpY0bvJa/rZ683XLu82i0HyrF
i/eJp7Kz1jVriO/NOSsxX8Glp/mM9+rmkkjGzZUbAASgVe1ALfSdZV+f21W+iAkB
i1zejcMXQFiPRsl1ZAFDWMUJA5PCXMQcqdyV1IBrkCA1T0I97tK78y0y00yEDTn8
LH6xZ513/3FmgA9Rpox2W1TVAWH5WUExVnCSdqvcRP6X2JxmS6Av6IxMwmrKantg
h9MewyntpSGtCHoyC0+JANCqjk10BHvJcbI2vEq0i1iI/UgMTAYTpm9+FBJy8yld
7J0uPcQS8eK1aAj2KGMw18a8wZB/BYOoUZNn5DqAGcIJphD9C+rYQO/6zILVe7jq
oj33FFDqZun2kJwoHbWqz/cYXY2r7+cEkk1Yt+qucJFOQgHG+x5VuwVPLQP8uTVA
ov70P7c5Enu3KcjJDsaknaXlxiWYWgDdOTTK94WVX+eIEfuO/yyoe03yVtwlFCD3
Po5qF+xBvpNtqwpTlP5/FatMvMBGQCcoRME8J7mNTdIw/QDZVh2HmtgOF8liJGCs
ISaBFnSnebaFZnQ8gNwQR4jiIonJL9YU/dPkM+G/Zc8higKD7L6St6VtBgyphvT7
72xAZXYl1WRlymJvN+qtH1hvQZnPpqkzCUmOwtK3HT1nyVb/a4b3y9cW/KmD5dbN
K7eNsz5QXjff5cWS8IQZ/+mtN7bSj9Uwas1i4K+sDeF+Zli3FkTQb3R0nb5TD2XN
DkMOMEkVZNW7lCKqo7V2XRqtRax8zZspZ1rbVTCXRhDLR+K6y0z/C8mUZ0IB111x
G7OG5yCIRbtL2EFtrUs0l6l2I7BegpUTi1HlrMI+DrXUFmqVMWl6bR6YU0szhyJa
Ggg96SAapSzTJvjRRZkWhEaCqCySMsI4+axuZBJLlbY7vClTHkqkCvDDTlDbTzCg
HlyhRZHVnDurPhv6Z5pcT7fkwFnASi6ntKlQ4VYoK5itTCzwRmer5xtH7i92V4gS
K93EywPBZ1rYS0mDBgZ9WrgDNSLMNsuXNxe2dBF+cU/DbrK/A9/7u3OATUWAqeoz
OJojX+doNhHOPAJuS5VR1cW4bqrRD6M+TlfiWGoj/vG/oXfj/MIdf0JaqVT5X44z
LcnbvHtzaAtqRLvZjlFFeRrFyqC8GxW5bzjVfwBzpC3TMlEmAyiDEmRXrsx9dl6Y
IwpUlO1X1QtmyAy6Cmr7IL1meLL9N7xSYWCBMBbI9cJHICRgCXfIhPBKBDhI0dIG
kcNvtm+CNM5EDEeFXbglG58/8Pt6wtawpJvdzwhBz/l+E9U8sg5Mhy1jJvwJ2Ptu
ArqJinfP2KOqdEkFbFIZcpdo31SzozctVUreYgciUZFw8VaMgLa9/qgRqdqeiH7/
GlrMM2cGpJDGbkpUdho7sCzTJtapYcrxjNIBncAffSB+f8TjYs1jmxG8qOaLpWfa
6gkjiGHOqdrZQxlaS7ANubNcH90kbw/k6I9DcWod/DzZ8A59lIw2vAry1sBViinY
XB+haChidTS0OTd0XouRo8rYeONGKrxOPOfMnejclcHSj++q5oSSTLcD6hPUpysi
BIjWkdkTC+psHPxbcdXdNXw53GQ++ihlc1vZinso0NH7b132g05xCM3ggzVtLN6n
ES4fS4vn8iaszAvym4+LEYITkD9zEGWdDRy/E1RDHEd2pNsabDHRbUzvDM2LpD9h
niuYFKm/VswdHX0lbGcVmjASAdW3bvh2VDuzfwC8Y/KofrAdY0sUSNQP+6ueaJhk
R+XDxvnLjY+NCPJ8B6PbspGGgGf571fEAAFwu7j0Gv4eCvHNeSMkNqcD8jKwVIKz
r3Y/yUIh300wcyh0BBTr0ojNl8YArWCdILRkKJfGTbHvb9TrnVX0wHoYohskLAk8
9+tfWLBA/CD99GUOJ2Mf6r+tqIyafrkS22g7uOXExWywnE6y3CtgKrK3x26Lyfzc
CluTwD08SpCkdvlng2v51R4nXOmoz5ecrBzSUUW5YQ5utlgI+t2BgFrdkjA9ZkNw
qFFpErx+/BKu5TI0TKoyAY4UD4slJhUY5eGHf0e6TLHMcUqF5dWa3wtKdaklIUgt
QpCX0WIC6sXVFxva2H9rJG57VK5yvgzkd+NtBVwzWh6q5x54XQMtxo1NH64poqmp
NKsMjPjYH6kfvB1rNXy+q2tEmapJ1gXZrERq8Ah2AldRgQrQISiUGZ8B4YuqkpV+
S8OKkgH7wXXb3IXR4K9q9HNirD9vfovMsgBdxpdnqQcP9vt+VSugXTV/50ZkINqv
JjVBimpsguqYVo8h7COUBR2HZq5YnBmbTxr1lIyNYSArY2bV9F7pkn9zp6qLz96M
Kn65jiwBOHh2F0evx+E2oNLHJ/wHg35PkU6P/6SGVKJDxqfKSOU++cgoXulAVxwk
mV8NddQrB5igTeudHnWN5v7F0yD7cZpmCKUVXqDhTMBhDfod/NxZ7qbYpxO7ezYK
DihUMEjzTxWMGJv1g4N+6cZEq0GSy4qbvweLV6lwjHtUlEEbKGoRahOGEGsk1qtz
jrW6X7LEoqmRaNsUvlgxrSEvZPeZY/AmuY9pWAeH1dzEj2LXTf1FvC3y9+Xgtcy7
Mzku6NP09pD//hJleM4FkChXeQWrgv/aSsycUTbAi3RbCwdXvuKrbSG4pw+MXhJ6
I0BYDLg3enmm2/Ciqd0Vuhj5cNvQipOW9CkQiaduyzyQF3/cMcGyYom14nNnutiI
JcYIMBIpq6CeXFByLu6T7nXEzwFOIRhgM3oonggVtQzW6T2/o0N1kQu7PY8qYm7l
swR064lYrCrqr0hp4IBWYjpCh+vdPh03VQEG4BQknZtuJdWVs06ONtb4ZzjisQNl
KIIy7/fU1mOjrVGNNPonXuSe3Zj16a497JmGWWuwT4QnqpcSBG6hpelvawFngLF/
aQVhkYfOIdcnfd14UKEIAEnzEzkZqmFHDM4r1Tsex5qenblnhEJ3py/AxK4HDQWB
V8nramzSyn8YaruM/3T96tnKWV2IHO3ygfTzcBeRWGoi5J3l6Mor0GoCRt07t8FN
UIonBt6N7xYy68o3weAP1KfG4E4M8yJx1a8tfS6SOHOC838u0H7MtiUGkYsgEsHX
bBrQ/NvxtSkvBLjucJ/8Prpr6SUBtdHvnT2QptI749xgtodEk5PXbrt/RVcwumHe
QAJQaHZivYqtLwBHMxP7gnJHY3iXghqW3ge98kJuuw67ipGNxRVWfnmSQmkb+ICI
iIIM3AEKOlTOlLIFlkEWWHiq+42sKqma2CWXpw3J2SODOz6N4L/j3ZCrIknLHTao
oAt33BV4ZO5dkhsin3i7t8Wy2u6gfurznMebZNDeUQwj3zIpSulITek/FX/9Qlws
CnMNLRXFiCkDULHZnatL/iMIHJPu9Q7t3KaPQ5/5elvBT2nC429idkgzSnVk+Qru
dhK1EPOw551s33/wV4Y0ZwiSbXfodzz4z/jAVw8KAuK+5RoQUpJkkrHoG9NBKQ/A
6cZIl3q4xE9Ifwo1vMCdjT07iUU/88oBjPeJkys5rFimoHCez+GmWb+W3wlXdA1b
PAk8lKoz3ZX/X8+ONHVhtm1NeD8ep9rPZglnMvOJ4yrqPYsw3Ffh/Xe9IwnxBrFp
MKeMeJtkr2rEqxReQGXg7qI1LftOSftEjsKHV6TXcagC/o00mBHBatN3A9gU4zzB
7NGe7iiQVcyDuZP9o+jJRR2auFl4HWk1LLswyINXdWgGBkq1ZBfG2491Qf7GmKzj
ogFbEMlxuakMKpbAx8p64EXnAucSeEjkgto/KWTGMUESPQ4ccqq2Ee6cH/bxOzGG
SFNRqy2ynNFsHdDPqoiY6l1D3QHekYEexaTeahgIAd2IrP6OpCqxUz/PHWXSqRVN
KSO3irUzFDhtiYzHP9c/W3tud2J9Jep2gOBSGeYA2bt6Dt9wEbwPyXvpQhSEv4Qz
v/WLdcUi2lPA0vEYd8e9lc4CXgKympznXUEZQVOx2ghbZPdUkduwF1MFZKhPQwOS
kN7uFKns5pjd/QNm/eDDFQf1WZdM/QpBeVX3iLWugs20hzPOIcFsmd6awIcTDZ8/
Qy7m+7/RHrrD+Crhrl1qiK+KcXzoUtV0JoyBJS4kKkUu28JPqe58EpulPMKsgs3T
Pcc3k3cOhURUVaU/JHeANo07sfegdmBTFvhscn7GZrBNOMqEyufx4x5OEBwT3dn+
ojfKOomv2kmBig3QVcmsB9ws2egRChBRzfxbDfGrrKaJm/F/KrU37pB49p4q/pg0
eW79LahwO8tITj/LyJyQzQ1diaJEWZ/rxw/SZ2a4brexFksmzip2zQYk2xBqurTh
NvB+tFmc03S+aYdbmpJneSXBTxDgHUrxnyv4vnPzy6Iyyw6bh8lRiLexSje2ID7c
2gWLk5+Oa2tf64HYWJDrX3caCdMLk/UWxgiXuAAIzjy2OROfRq+qhEYR7U8RsSsx
888kV5vtk5cSo97Qp5oc2yMEIFtx/8EFlas3AP4jwiKPenFMr5nVt6CySaSTiIKf
rSJ8tL2zZ9szwtvLyfl2/UZaCiRH+kO58amSi/SaO/UIqEaTXWwrR5D7Dt+AIdst
1vv4YOXfliUHOU/U4xTDNmYDgovVvHkWyxLuXIVPVnDrleaC6cVz/pPm0bwuF5zA
TSQeeqkMmOc1PZvSZdndn/nI/PQ8p/xmHRgS92Qpd3VDPU6lunYTZz22+Akzz1fm
tdwgRavtaxv2p2UQNPsLW+8vFzmvZuxDlMhmgiMkOmsWNra2L+QOc0+RbKbnG2zx
1a3gLVWYBbTI/2uPEvE51TsHjUM+7uqBCQaZ373iwqslRRO3hyQICyU7jbnolYPN
o2IaTE4MlSCHrrEDpQcqSVRx0Lzjl3R+qVOrBRvRcHz/SL4jip2LCLHsQfR6HXqL
6pp5EQfMLVvDJ+9iYlWfCq2QRGg6+dnwOy3zUEfWeBtz+3YNgCY6ILf8f3IWtbIO
X/5P6Gv/ilfeL4I9sWX/T500o+ShhIow0QV9Q6GsIM2ZuiYeOIu/DE5mBqlKxfvF
dlLXw4s+xMIQqfbi4FKjBp4F6tpdQwpGwjvWLjmolKvjfeVJUl6EndbTWpB+lsiU
Cxs9T1csqqSw5p314J3VNT32a56FXokretNrvHHJ8Y7P2e/CHVI+DPryWuTrowjg
MfASuw7zbwmtxk7q0EFYpx+3k6n5PoQSaa3Jm8cGW3sh4n3K3J72k9airEdPUoj/
Rj2IFvXdpe9XA90JRXeWXGKaB0JvDxNWI+SZih1b9CeBIhw552WQBv1JI3eRBBVx
dKm6aG5sQ6OQ/aI75c2K8KnAKE28Hf2clZ/0srbp+arnG/rFaOCFlyordyjGB+0W
9BsvOk4v3N6I2T+yUdoKPoaWff/fl9CiIx63KcVU7tIGPu5ILMq/9msDN/Toahpn
WtwLa4dBsRmFktxAyEt6NneZuV2NCw0SQSw4xbBDAQxQVongbubEx/QFhASPeuLp
iMN+qUyOsRtZva4cg+3HMufoJB/1I27ukCcOjotEMteL3LTCKC5gK0q+gH+MYWX6
W27e15CJFUBMG9snDf0BQd1Zzx+whovqtcawpZ0d5kogMceRaJcT1FAGOyCq+9+3
H9WClBg82Rq/K0xxHhAqIk66xxkgkmWKIMeK+412y2MCq/LNMLqsrbw8Tixb1uqU
1E3SifHoixhPazkVlv3/QmGuhs/5vWggKxAL4PCZK34V+OgpHu4W7pXLbsovlg7j
fLM4qZf2KKTx3jHKMwy2qwEvZYm0Z2lCfgEZ9jpTE76dkHJtd05niMVc+/AmTUwn
LopEVOEFJ9twJhAYq78VDALzaKhN9FjmXUbnc8+ORja1pF/xI8TGc3Wa7r6W4+V5
u7eSrTO6v8IGrBr5ko8+uDebKzTLxoXgrYfj0eb5peMiVN4oey4L70SLS4IjXEVl
xgjkYcEkcIYTZYHuitzcpqGS7hREqdy751WNu0nJbDaERsuXWzPJd2C1sWi5e8nu
cuyfNt+pF2GM/zD79oq/vLtMTQWHPHkggjngpnSpnJFV1nCY64WBB0TtjSE13lyz
7p5tEsWTI2bcF5Y4uLnYQ0J+azuBULlhPHo+XqE6oNVvew2LkJmtkEnh5jEk9sWe
5uwydCEvoKRytjYueIQy6buDgJozxflfl2eNU53CgU3aVCofX4KTweSZ2dzQ23t3
KqnWModczb7+P7nSsMZHKMewhYC5B3tzODiSgiAH9QY5AsaeqAlmtW2825Muhors
cVA3+BXFiXLxcIrL0ii8OAA86Lip9qS9InSE6ViWFIqAtV1BvHeS/nzDoEqcjoky
6RO/cI0OpfpcIdkZ3WDTMDPhfLURMYU4GnEKAieBywNjmPv2782H+s7UZsJ96Jk5
zG+iyxQygR47QMhEunMI2wi0gcntDVcltwK1Jy3wFiXB2Zih/pXlPDMBKWqmIna7
0AnNOEvRcFNjDYKmHWD7MummurNxW/m1oohfPUw2cP1trmHXzZ+A9PWG8UyMqzms
T8cYJPLLhgcUbzQJx//WDF/grRnoXd3KB/5vhxMqEYw7+2lsCov7MXxYcdSaG9k6
IIsyy6ImboJLxeJ5cwI1yxkAXkp97GRDxagZk59dmga2SEKlpSeHoZWVTS6zbVFr
wB5OjJyunn16+gLk1sC8s++ed+k1pzg6WgLOM6hjTr3LJ6jEqJRn5FwehXb45xyE
VFwZYB78KZPn++Zmp8Mk7LK2pJZtb49P6XrAyO+j+femwjKCRUGqE4KSMlO5/xBe
D9gkY6x8jjFBWMeeHZ/ZMzC8NG6GD/a6KMT09L4C3AfXsshEbA+fMSfDrEYfuqFy
fUk0ogcc6lceKENEHUeK1aC/Po4ZCnBDmGktTCyGdABo+4cf6g+wPcBoLwKKX1na
YNq9xGcB9Nw6ZqeRIl1gzwAXtmlUNJuP03AdyRCrePExYfuUbyjWm4SBdxYdt6Ld
bQs9z2nsuq/aaaHVOfoB4McSepDjtI+1X0Qrlxelgsg+WB50cYXDW2jJZ6HbgFsx
U2Veom9eEZ7HTGqDIdZemk9M/gYgJbaawvv0YJzacbqVdlQmlpSLFj0r+WzZoUYM
IJP/rf5aky6EhWD5YpAb4pGqg192qyme/q60dzjdqQoILUrH5NdBvxR0m41gSFFs
NaPsHCG7WWb0h65on7Rls5iYZImbMNOYKiCuZarZe+pe/gbyeOEs1CR/2n98eGXI
e094h7st3Yob+J2IK6UY4rqzQyu06geFTAip/BWo01sNtIsONYvSdGLrAmmi4EyW
/fhvyC+oEoNW4T10eQjgjU6KHIZ/08xOX/hec1Rjph2t3YQIHDxwi3XvoFrkMlYQ
P6CrNaTeV+x0CSBxEBHi+so/4yLyFHDl9qXBCVRakZYLRQklYSCtSwJlsF9JScUW
9A30igyjCkiJLMf1IZp2wDdO+zxwtRzGvS4Qk/QzEK3551s18TFuX4rNbFPl4Ao9
rux5OtrdXbPT5SA/f5tyI107PBN+7U48cn5LpQxf7qZlMTbqn95JKMFBFn1+SRV9
PwXzgh6glRYaauF7WtQTvqSCHgpJzx4QgjL17oiGjp/H2AjFzQ2FrYTdSOZys5p3
UJeE35EfDOjv+dgbJBzawzaC089guPkReMpOGH43wWJyomVVx/GuucrxvOO6sONR
vTMOlmJ4HBWxvOTXuI9TaUYJyE6S5vDpOgw5cuA7M3GBxadl30u6BgxDmz1quOt7
h5v4x1HvZOOglrCxbONVgxMQH3qvGdbufHxaGj4CqVP9BmSpZMpgTFb/jAXRnz9W
3bvj9Xoi4+ZtAmDuzFq7fkVXo8+/YAzoIpB/NeR610L+//HbHk34FvW1pbgpp573
CURMKlRB9mSTAqPO6kq0n8zYr6HJEcgKBXv9cTQ9d+CN4smtAOaE6f05H3rIdeRE
CenOrtQUEPqskCkbTwWEKrVbKC36lWNIaN0YZJsN7Q+/N6ESHfGlh9VFlwaVBuQ0
1gfHRYl4yVyUJtQOylW/cIeZxP6dZqcWKJgoKLAaZgK4FxSplCRpUP8LRL4x3rlN
6PdQbvWibD1MyL4UXAhLCMDVGnTdtA//NDR7eyI0R1a1+qc02csNueEAogVlc7dW
UXKzC8FENu0AS5WNvtYo4+SutWH6bWZKKZ/6OfIfTXh5mU5Iuj7jgIIfgqevJvei
u+gdworkIUxMFpRzzPt8IwDtadTzniF7GQUFySD4zHPdmfl+IhveesNjblB6xclq
eTCr9kKAMfeOFTK93tktVc5s0PIJiaSxLtNV5CRuFbNOo9+hE/CN9bGTRqpJtbPh
xk9OJxysEexahiV0nfdYluuStwlMjrYI1NBxvd3G4+OrIl/b3vFY5F4G/eUzdJ5V
Nishf6Fswcvd9mpU3qbPZBTi7FCBHaZw3V/A4hbi6cvSSA5QTw3wfywdTbQFkUsm
026crc2lse5r4Jjr+btae44hv9ny7Q3wwE7saJIeCT9k3VKbmaQ6LY6VS4twM5GE
ZJ0+v9Nx67WAn4lPEgFwCO6S7050MkzCsnq5YwVZGdRwOUoJdpJtKXQxUUqNHzvG
Rlz2NeUKWgv2E9AXCGoUz3NyGPZW1VstBLiz6tOvpysXkRvgNa3UkunIsLPBiiqx
poaKZU769Q4xHp6IJiaOrmX0M4CK7+WGCUrZOQ2Z/y4xv/WPpUjvCMKNUqD7nmli
m17TSgMG3jNyVmmosyZMtKCeSPnAnj9s4mXCglzUoXqJ7XuOJXFlS2b+chmuQIXp
2To4sj7UZhyDa8er367V1H/P27GdsIE+MNZKqe6tF8rjUTmx2Rh7R2g/e0zTX7ZA
AUqF9sHL4WNrY4XdOwtkc1oxakzcVbEPu+GGKmsRdVIVQJYCX2QGwKxT3huyOgQT
HwKzv8lG/w0+wAkcEYdm3WRe2fA/WC7hUbV/ZXxAMro32MBYl6JewlgiLDS6cQ2F
705tqQTuTu4xT5VQWrU0WOnmU67jpagL5QWDRbP9P/O6mVG1Wwy34Tv1/OIs0s7h
ChIA7UhytCIzxdt/MqG6nFqSDJuU5n7f3AIDWB732YpccBVcMe1IUIMpoTI7nxol
8NOhgqeOl/Zjulkb7y5rWRuM/rydVzX5VatKCmKUqea+0WFa3rq/bC2WmtlC2Pkd
pA7s4abTriRKxtjaXLkqMszaU9xYDVO8Df8RQ5iJLBGvRZ414ukIFDjIfiJ/f3Nd
ANHrCftt8u95UxRmc+IC9IGZIIw43nDqhIhRVW/KeVC1LXpeBChVicGB09H0gWMc
xsLGam49XjS5iiXBWMOcItZKO5BMMN+ktzAacVHRtoB4DF4yGQdn38pYtqg3nqTZ
8Ctro3wMeB345CWOl9aCr3VZTynM8tc7F5oS989kEAuJZDOkjng6ZrPt2dSAEU89
wNraSHdotY6wYmJZxUonhSVkqWndyaNzdd6WNjjVdJOdijrRs6PoJpZY7f/zDeM6
YDkbYrHDxAiZ6Xhpaq4l4wqH+0vLXgXCMrrgQBCZzHbLcJSthsMwinsdF6sLXg1t
bD/I9seoqNYy4mUDieTNPYmReu/Q4yTPl8YU+8Jekzo0Bl4LXpipJjVTK+2BYdiO
D0ogBiHhSAmWbeG5Hy6RSfmfkF9R4gsxGw4Q7G8987vJukx3Fd9wPF7XG8V89EVb
UrZryYzeCBQMuHG8+P9w+SUoE5iop2Sl98Feti+qoMWyiuENJHzu7/afCggsBfq1
/f2c7zG7A3MI0phnp56rrpy7xS8gWCPs0MKnVsHJ9eWsxImDFuiXa+/IsLyIUZSv
eVkIvqGDilVK/Oxx2aiXJzKQldm/akXs0vxgosmsFdSGdNu54gmp27utpeC46Ckk
a/+41Ud9A64ZiUnDx2Zcl6xC5BSnlBtiskpyxCZwyvB2MH+jmT45buh2cioopUUu
KZJu1DL1+HlA57E2aNNiA0QfL0ZDJvomEfl1Vkf7r0ZD8rViff9ZxX1TrNPqi92n
uLCx1rq9NVMfokBFy3xwUMFS4212+jWcfVA8RT79L6FL4JLXmka+gf4zPf7Ik+vd
mHupMvQaFWJNDtk2Mo9oa51estfpYrxCTp1298nl3+oAjkaC7kFAgqzbS6rthYHf
EGtReR7ahHBLhmjsHjnVI0/Bm++Oi6PxihY3ZFZ8v+5oqDXqqysOkeTmv3FU5oVK
3Msuswi/nFcZcgtLX4BfdvpS176vIkh4sMSZpYYKuVq5w0kkN1N3sbGod+UE48dq
FWzxp9h7Fs5+XP9xI8xJFUuUCFr+IIrWPepBbWJwiYKw4ZimgrE/ottdt9HZXCrz
pnHz5KGzQ+4XY8k9kPW0jihVGpvYXSavFTxl4W2/i+sjzrvPO2PINrE3ZMLlivSJ
eeKyH0qVgT19v3+ctSMDFGZ9/s3zgLpDEvchLp2LTpUckTm+cqtMAHUDAC2kV7Tb
2nhAW71g2p7RYgwoDRQyxNXPcv4ATt2z1nXr8fHB8lv50Ie6SzFO6E0k0eRIJqaY
7x7iU+f85FeJwnguOEhAzIypurTBF8qknTHboMt7+OBpHOwHJHxcnahsKt9JjhwP
niJcd73juH3n5r4k8qYyqRZdAvfPj9eorMJZRMdJrn4lxUIqKNWRA+5s95dNUAbp
WGS4n2Th/g9Mx7uI1xQNSwUMfiiP4lhTSd3OjHhy6tlREoj1btrqNW88KFJkT+p6
Q49p2XHUY/YblykRSq2K7UEmdWEOrDK/meNI+HVoiM0ijOLzj46kInCu28lv6TcS
vJsb+kNNH2hASREPmcq2coAzHFEpmcojKwVQ5zKhXZ6PdD/kWYsJLOIJTaUvaYAc
sS7n/ONkEbB4rj3G6x4JWJca8qB0PITaZH18LxTkjc9HwqibpcjCPnR0dgsLZxKl
Os7kdyuK4WJ/2h3amfxE2kP0ZAy3aZVV/djw4C23nJMIa1oCAhF1bvuCN811NDGG
UTkNVMPOTEzdCKPeZ59+Ap1UnQv83m+dOu3Dvq1X328JCyd7ajcRYeFB4n3248jx
ZIhyBEs3jPbf5Fl0N9/kBLR8qwS60pOVDaJy7FEjf6jIn0AiKMYNuZtN75ECxdJK
AdNl/lSge6FtTzKtxWrxeAYmwTyPM8QtrYO+operBfRTwHiSidD0mm+WUoJEeblI
vF5XgyPMMKbCh/BtPgEA7JsZY8WROJPf5QdryHJRabkvIcyQsbZbFq0fbyYf0H+Q
f23Y0InkQoWOaG0XfhIfe4osT2Gzmc1XK+cs9syDqXSucw5FVizVxQyY57cAyepy
LFN0KkSTJh9LiYu49nmXPBLKnfKPBhYfRsPvEV1n0W8/Fg/VE+DTBxUs0S6waz9g
u7BXk+AvVMMzAmF4kH8QLhjq/wdnv7i6ipgewhrNgepawsN9fAgFFVW68D6BYfh9
qGWcNfIgdPpUrXOu9/9g6uGM0z0WXdmx5X36c7xZS4fUs4L2NI2B+Fc4l/UAQBqe
W1zq2bDrjpmVCxuxZcL/H1XeXD1dZg2AuYeyu/7RssBck1W3DwsJ2/eXkFkv8xuC
v98ublgw0EdekrQ6n5qpvlBxcJcnGGy4NePuTGyw7AyNLTZv/uchB9G6AiuKAzBr
uLeSxa5DT9rj7nCE5vVwGn8QedrIIkdqac5Gmw28/QHEp/AL5bm8/XucA9uFTQ+c
W8banozfr7Y41RbStBN8LXiJ2SriOmq2KqN5IHUegzF3up7xH2jXzkUHryZRi4T9
kB+X8PGrB/Ul3rga3gKejMfXDssnTQ5/gNgPGCwdrNFMG1U+iMfcI3KrTYQQPqSs
VX3XycMRuAizvUzR8bSAtJqqK1/wgIbFqeVgsjBIuFNy0/pdHKuFmGeKoOG9ZajP
Vu2XuLVoodwXPuQhfPo8d2/0SJoGWZoN12Es6D8mFIeoeE4RfOc3D3caaHwugCvh
CDtcWVQvMN2Z6BEvrrnslkMa+saRNp+E4gF+PBRag1tklVgeSMrzIXH1ZbaGJDL1
T4sU0xfmCNAyvd8lUX/JDNeqfMlqzw93kMLrtRCzcHhlbR66Fxsz6nIPv+iYWnOP
h0vS7GNEal5lil7KJKyQNA7RmQIzW3pIvPKFR2qBmhcYrzEw69RO3blJ5YENAZwd
8gnYinm7F9QFEBgIYlSYcGgjWDJk14KfQjacR3ZE9XWxdnnbef1vac9BrhrBnWNh
UgEVZ/I+qSWmzAc7ngYqjnqA1b6veLBMRoxcM0f1Ov6sSUxdIzN3y3LK1257XMpY
Sk4xqblpPieZ1OsBTD6LN9TnjkAt+9hYHyrQEkgj7pupEq2AUoViN/YsqZga3/wB
3vhsHxPI7920Uuht/bhtgrXki9xUOQqubMqNgKKuWjY8RIp0KdMI6wAj8xNy/duJ
nPe3tUcLgOFT5/fLXd+O2FA9OD8ne415mFVGnfS8bPMZgnu1L1fMHk7ZKo7RMrow
gk7io8KEASAxNeOjjLgHsKvdIwH7U0c7PZzcwgCr1Y+LvshMsOdG6Xt9v8kyZogu
knKwx4cVavTseAnwk0NfpIwa2ip7glIDjurhOIgaUIrk2LzI+PKMRfknK7xGw3wr
8vzqpPRYlTIdk9CxyzEuGYBMn8GsIBzJne8kiB9ssicNJ8LxfEVCWnDN/Ei+cvFm
7L8bXkkmcg5/A6yhbCxfLBCJ7nQjHZgiGrOuFANFvhfPfZtsp5YnJDI3Z6ehjO5Z
OnMd62JOD1LBD2rT5HjV7fnTjY0fPUtNtXwHH/CaG0N23xSmzkn6EN+w8AaJhFIb
LOEzPfgesdaRymepUAMN8PaRZQ7AOBmbTPUfRaBnHlGAkAEkRUOQx8SS/NPbClAd
5tWxTOWrvOKuOtMug3N7ikX/2yeUWIpIneHynxLsuD5IUSyVuh5XZgfQUPm9zaWN
uxsEXQc+IL4Kge5/tFcHz/uTuIE5N84o4bzEi0R3tXLj9eGLKo7xISfLYE8XhUwP
G5emw1jeJv2o/14SH+1hmYTSVAtxKNUWJezdR2ClQkUGhWFtfwvW29v2b8Ju1kkb
k/GIenyPDhG9Yiwury31FGsZzkqgvB0k9nfQwXSmmQJNhnTPQ65sfBu5uni3K/jb
v6PERwBqEJQvQGdQe78dECc90IG4lQnmD+UbjZfHfL6lewbgRD2/dtEKPEjNd8Q4
JjaQlElT5GcYNEAtG/LPl/HIKBTBnnDI/Gofu1LR5y8jEj0+m560oI2qTlKbwFO7
x6vp2clWZsela9ByGj8BF9YYCEPZNACBRthsyA7Q9glpeGNiQJdhsIAk5Rg4NJJj
zItvJ39thoRGT+k+10VZv+2xAYAMfx5SgNgDxwzqA8tmFle4hgnjcycR/ibZSYCl
rpaJT+gSLMSzk1rEBJg/FM7U1wnonWdCRQt2eIMh2S8r5Zgf2fyk6FGETQlTC1VV
DUxzgh7kQG0lwKWQZ3SuVbC7pQ/Vw1sb52H0rgGJhaJuocXlUqWTiOVzaZ8tktw9
6OMvTfsGdfCNwyhWpcArwXJZBwL76r+5mwyzESvw+n1v99yQq4MGi0AGib3Xkmlw
egfRSbcMJ5D3Yksud+Dq/NlqkJMe/HHL93FgWvKck6gEThFI1ILQAMwjk4anhbM+
q96/e+MGb5jWFGFc5Ed1Ii9XB6kQ1GRDGp3K+U7Lscvm2OAz6Ek1T7sqykJuPNYE
cbnDU9xUwnSbt8Az4mLj0rwrStWAfP770BWL1FJbnD4cQoo73gfQfgNeJpx1Yi/H
6mKUpDygXgTRQLsGmV6fXf002vHM6tB9GKJk1T9fjeTZeqpXcl6/aNQDDCrHOW0t
BPBTMgXjyWH8V1L4MjXjFBumzQaUvKRIC24tLATcavCqwcQ2g1pyE9lEQTLKUigf
kIkWr3koDPnEaP+wgCyfrV4E2qVMpGZ0UhOTmInHp00pr9nlo8Q7CsXZ4EmtXDWQ
fAqgUnZubz/OLxPZZGAQuO9Uu35/eqgR6IYpnzRpM5kkY77b9eX1lvUzNqGu0mzG
BDANtwUKTJqpRuimpnuVfXelGvgGqsoPqHEju0I0qn+DQx8E7LBLNFZIMa+ZmvmR
Wu3TDa9BsGblXlJsoP/GYQQ5kohnM7U3kBnlRi8TinlfgShQ1o9gYKhdH1oyh2Rl
CCcD1jumwirQ0fa7MUgYZzooMbgB1EqIS6K3OBetX2KzbydYNBx5E1vvGEegY6Uf
IFF5R5bm+vzC4Cpm+wo97a9wpoQhRf+leUNsppRsYbnymoPku85pyBBURolDzb3c
lMeczP89127ZENoZCMNLSxiyN6BDdU0MX2nfqPBCdVfZ9lTFSfNoT4Hnn7icI+kU
QNwWgO79SBhK+GF3RZ2RIUF7Yd/t0xGKe8y6uKJMSHeEtlwplYjtbidzoI5/RZyK
08DE/NshXeZg+92RmkRt63GkECCVEeVALouDcrG5qaDoZR4ttOBAVY8pAAyD2XBb
v0zmJkT+ygQ5fTGsck0iR5SjitUQjB8kzStMbg5GoL2e+j3XFmRnyV26No2K45/I
mHdqecJJrpzEPuFRAiIkbkp+Njl/Aha/0t+Bi45W+wqN4BSPLQjofiV4zXf73JZa
hLM1107Jd8+F4cM2VV2zRnQpxHM+AyruOrgU18Q+MqkuSEDeHCdw5paDnzFqTC9X
d7253VNhnqCkLe3BRjFclVom/qtEi3nQroCb0KSSpnQ4QmATNYMQpPi7FqCEu51v
BvJ1O92CTnCrc4ihbW4qE9BgcV1uyxF9c55AGxCzYP6tUuD9TxbYyxvRIB9x+Kkb
vwEEfoGTcFvkUL3uHLADm5md1uvPnmqgmpYTcYz47rlAg4wR7w3NI9+V38q8/DoT
z3HOnBIw7PbjR0gooFJ8l1X+297C3PBb9bopT11TNAKZUf4AJwy4avKzTbA5D7JJ
F2g/rAXp7uUoLeDct+u3KZ6MFaa4LHXaBer+AreKL9KEaYUcXqYqnilhUo/Fmlzi
59a1ds441SHpCRfky3jMwOwCDpcnnGawxDGQ0qPKS2eOqyI8LQ4/3iLKAZPPMbro
sOnfH2+o22hVDgf0O5n/+XRgm9lDnQsQH8arSnLrsmjwZ/Jajo66X8JijraEnyYX
Bd6UH+RS/8NHQHJq448d+SiwsIvVeea3ROemDYZVvrwT1p8fTi+NRhb7UL3lhm8O
AIimUjDt1srLlZLdKGkaIlw0efH8i1MPBxdovLuccvAUilSs11WXqJD2Vz+qqW0o
Whtpok1OIjeYBZKFr3Ek7T2ev79dtVmCXGiyUaghRlmb7rOu+dB3MtfjO+5twg8t
PrC0UqGot0XE6yvND3yc/ks9wmIsWrm1XBllO/dMJLkhpKXE93tD3Ifw2i5bYCdA
HCAGajwpA1cE+LrTJr4Y+qNjGIWy6KqmqtwC9AMCnt22/iLT8kvAAPen8tA6K4Ud
AzUAnXNNRsyVvJeYWk936Z2nTDtosHSRvFerFKD8CgDT8ZrE5j35B7v8PPAQgp/T
OALqr4RWNLTb/8TvMhBt6ZzTIiTML8vXsz+HqiQ9k9Zq9NgmkWijUPhni2hY3RFl
5eD5smqG1t3iZgyhwE50zGcYTVIMf/JVZ7dDN3JsYqIsSBLiC9Mt3jy8Yd18Bd8v
mhbUR/DrEW48XnN4rXZF4Ywx7i99Tj++d7uxYFqqEOzy/qAC+ZdFe+DGxZxK8Egx
d6OTdTbTSnF4gLc7LKIgOY14Is6y3lkq5R+8lyAgrlLcidwT0kEbwPTLJsHuA0jr
G7l7YgJei5EvzUWLDfH/Fno5tbyq34HkDDQmPLyopY0/uA9lNZIW4+QlWt3Xd5jy
xZnWlcIqL5Zh+T199fzMerblNhlEGQ7A0olyxhmWWI0qoAbnCaW72RfdsyyAl3ZY
KZhi/UiSWRBSDgJaaKF6UTPYW9UxZuhR1cLm39EDXusx1U1TDMdPshb0eq8S5NQV
ydiqwJR/XNKtU2tCEnMm4kFRJiFbeSGmSf/4JOUhUj65INur4o89ESso4NZvbpCO
ByecUZiKGYfUXs6AA3lHA/vHFNY1o7BvnufA1BokchF/3gA/H3vVZSuRdT6/vnI9
eTJRg4howgKTXRXTPprUxnQFh3Pdp3Cuutd4OUeA+zJ+TJd+q1laZbPzaaMnmi63
ASpv7+woSkQkTkjpIky8FPZ4spLB3y9Rp+/z07Hf7/73sA0I3QicRGDLRPkeUyn7
Rxerhl9fZY+STHUMjSzl4jx51sDRUMbz9XaGYDL8RiM/ZjdUgxK+/idgkhGlm7l/
7Zgxdly3H0IE0XY+CxXnI+78iRHPWCY9pZpLIDpA1LyDR4rouIXodaWWotV4IPZe
gPa8a6fPwL5C8pOXJIFgNmqDr149aA+l2SGvrLRzzylqnEJcmU/EhMfvTw8D3HUo
9WVnditwZLrmkxBnbucj9WXri2vmEjT4mfL6qAvfXRsk0B4lGKcQDR0SDVLPMW7o
ze1fTixD4dJiw3HmaiycuiXNedHKZgg7QzyPmx/Rgc/1aRxUGbsssmEVWE8VIEJB
+vTBdrBwmdWf09QAAcm/sMWFv01fp5oThVkf7wPiSJ0p5qFVYAucGvUkqh3q9PMp
0Vijq5p0r/DfFpY0OU3NAjU9vApEMjHP48ACZflIqu9vvr42FASxBD5vo8nR97/h
NI5aQltSXhmnJpBRiHW8XKqROfBm6SJwIhm6z/JBqzYiWLcgqgoHydhdJavzVXF2
BwbDDGIRCsHqj6RnN6K+cWAZLFD/SMH0KCP13yX9V7ynVcCeMB8QWSVmQChI5JHF
OzVCoGvxbdjgthOoB2NYfV6IagYJHgFPPMmRgxk2fX41c+d/jILSMwfSWjm7OtEY
igexYipk+VgFgC8y2/dNAk9UJ6ppQIR6J6yT2JZfohC8iGnkihu2sYPzjJwvM4Dv
PxNXp88mKEjcjHGOys6/mpnnQXp9eSNaROv5DMEkdMOdhvW2QD4I/fLQeUfyahsK
+0jXpFbxj2sTFp1I2vz6NIFWaLPK7p2shE/hd/4DrdjaRANK7J7YM0DSzxHLwW2I
38zhgL8mU8KXkYGbq6RfHjbPs1Zaj37LoerKGA13A9zHfvlSCDQwVx7I1gDdkh74
tU1WZHKiaN52dUmoiSvA3kN7MaGI7Fciqb4sRSxg8yOX6oI1qb9nevAeojHIY0hG
KAQoyYxJB5919yfr79ID7cXo32G/J8ds6lPeubgFVMb1N4thZjHdetnwjaVcVzN9
S1hfMQOpHb3yzhnKIdMGkrn1hZJ0z5QgXRfxnF1x778d92Z8InSdiOLci8P1bU0y
2W0BkDbc++ltER5xHLV/fuSC6BVtG3wMjSPf1ms9CI/gCG7adu49EUMjFojRaWj7
GMQe0j1e7c9klsNaKHrSccvX6Bt90Nea2OvVWpcMVp/pE0YSfFaehX4W+tVxW/lU
jmjwtWxuFyvLvUTQZ7SJzP0/2QYUnkENuR8l7IRPjuSsanBy9WIU894TBQxEIrGj
LxiA3VpyYxKeAjIzGGDENINcY8eafj7GfACEnkQsZwxZbK3u3OrKqlueUdZ8EQMy
8uPvvCmDrMCr0EYN3Z/PeH5sXMZJtje60uhQU3gGsDQiJUOK34oXkDTC5yXmxGqR
6XHHkNTafHZU6IfM7A7V10jOEJZCtlNp+cYHXtYcMoI/x9EDtIFis5VO+MGq9jWI
1YxzrIM0EKMpK9VRMJsAM8rEayuzDRyIMASk8sf1jVbH1ToilsgF116hLxqTksnt
emnNEr2XN8eUCjPUddj5l3KaFEb8jKCUXQyrtR9aSGIK97nvY2C311128+fBv2NQ
Xg0K2cuJ5WUgeBFfDoXx/v+mXYXX6vJdYtmIjw1kNRrtJthclMaZJZ2cZiXeT1da
mt7vqAnSd9sL/4942G2WKa6dhRwhVLbkuZD62RyfstaZ0IJFurs3A6ubx+cheCFS
2EuOHZiUrCCQairFWcYYx0f4T1xtnrJYSGoFBHt+Cmpj1QScfLhMyUEUrSNowLYj
m8QFi0e3IEAfsb0FSdnXvTATEdBn0DwE9yPaDLLeNM4iWSgvgvJ3n/1SdMox56re
1VaQDBTq5oKZyLDaNi5G+cBkkxZFJPH2sYwqfWwjm50GDqqZELHL6DZfd5aVKKP8
nxb3SEXoKJUPYBpm9wi5JXIXSLTANYmDGgh0V8lwH6CtBBMgi0KdveicI7TIRVP8
PYV4tehhk6aiOhJePMDyITjhCsAEFqOrRoDKSu6hQOhMaukijDn/gjdF0/Y89ZcT
4REopaSaQdn4sDyiceAogjp5SY5g5n86X6jtRxn+v8qN1APAUAtBqFVmB7ABEBiM
h4TY1bBH1cEqJRk1KTQBxfb7ZnUn/xo0HGgRsKSrVhJwN5V9l4VX+snTaPyHMbmJ
zo1uX0QL81TUq1fzdaRoBFxnYSP0omuiond/rq24gApF0DcaDcG6XV8+ASBspGqM
EZghwKvGKjoaV/sOfUckQNsIsCQyA26+g5pliwNMVYvAfnze5hi4l2qAY/jAJbuQ
Fb4QgwxoYwA0GwiqOrkJX5MNW4Jsq1qw1szqKoRJV+mjdfzM1yTdn7s4QbVduZ3n
upTKjSUPs0bmmbOkQfCm9rwlPOr2VdJzoWr0plIMsNMY7r8fDHaJBZrJ8ttmSCCh
ro62JFVuacLowFC1dx5srImywBUMAOpG+M5zyw0xpVAOXu2Nr2jeTp8yQ7DWxudl
2xxfIFqzlOiIpYrIJ8XiV25nRVqKKtbscbcc4Oh05FuVZ5ljQB1aZp5dmY08Q2HY
csqWElX9V8dEtX8QeHaMCnsBERyIASoI5B03rRE3EqbGlq8oSNc95K/hCoKD6Jk5
wU5ruq22PVqsGEYrno2iCy+aPNTVq9LQ9rPFmZqP3xFOkJhG1PE4Sa5XiWqQK6E0
bm7kl+533UgRfuHcCSPWTYwRvR3rDCgIcxQyR3VuI+DHVqsaFQYkdRzWKtxP4UwY
qUyB0WzgDj9YGE55uagxf8a6C57wLgAfgxgyhXi6m6IvEmLT4DP/sJL0lD5kZk63
MmqowoQ/6Ukq16ZaRnc9kZupx5RU9KFbaKETLTtJHjUJLCjkdB6gemDmelPhINgV
jTNn5Tn6QE48WXATl4tRwneyI+dO84/8pSplfmGLCUduSEDc39CArybiaTSOp1MK
ef39IWyNtidwFq9spf2e/bFV05TjAB3y+7tcSVRynuFb7CkdFSUeJc0CFz11aAEr
rzOhnVY1fALowOnD0EhMLWLJtuvd6tWTcAK6F5Cew5QOJuI9AkYcIFB9aBI4QBLk
s0ymQGvzZz2fznRoJs4Fgtw5rvX6wQkIZR/G30pKoSLuHcW32f6cnW2qg3AGQylL
+eC+/ZQUWuIRbfmSCCizoPRJUiQ3DniOC5IUY7Lbvw6VdC+N9Wol0Y5bNeH4BP16
FfO+2cnY9q4+1mG6fCAy+Y/nZ3/VxKLr9rkFGKRWn5Jn3Ee7CGlmFzoMbbFR9FKX
YMRtJLiKPqHjCN4Eod8jxXLEgVKvpWl/nF3w3DL9+4fCuBPLO1X5xLPPL/qomRcp
YrfBoWnFIRVc3M2PabaQBt6qDmqLuNhD1u7JY8EWRZ4k+OzZXMirhJm1B42KyZAH
pNe+GVXr9geNwA5qpY2CH9VuA6EapebZKJS3XsmHdo8RYzeo85fTfbKZ+3dLkjqI
mZlAzFxvO4H7OTDHfk9KyzHOps7I5jpRR+3i03hQ7ixFbDmFqGMCON0LgjHmSYIX
gTIobameB/mn1N9aoYEITdYGFZrY236kJuz6BIkMpft1QhWTdfN4mDPJb/YYQlT4
TDhC91pTS4l3kJlJgeWHFRw+qE91+L5DGAQhjBwMrBk3YoRzq1tzYJRTmBBL+rfs
YF17PQW/EqNEOIA67H5phMPqdAwYWf049NGtnMdALOy8OP3oBLNusMwSWu21H7fG
DQ1+fkebshfKhE5NELT+mFZnGCSUYm8V/cWT9GCpRWMmMb7Dg+MZcq0iTdS8hA5X
gTwmwA14sYdNXqaQKrV0zhz1TcFOIYmUIZOe43sSx8B1NmLIVQHV7H5V5jtVE8QJ
9zOu4+xxS4/cJ9eHpymkxOaK/c+dL11vdue0vzE/dXMPv0EjdqUxyvFQh/t2luI6
/jOyHEz8LLOJHLXcAqXyIErf5PgOnJnOds+Fl5Aj2Oo3erevi2rkrB9euSsu0ZkY
91sdNprBjAyZ40xtHLceeWzTjQBWmc7tmf4RJCogA3CfGGbO8AJiu40k5eJRktzX
l0IqkcMTS0oIEr/jWTpg5+KuwMnK8sUMa4O/5iGFsXf8zgmKI6wX1jUdAyoj64i8
2MQ3EJ/doFd/9zjMDYtHfv5XsL/cmyWEGsc2xSw+LJzoX+gMDwyUuTzwEVY69qlV
PcKlrDXqDpuDW1ECy+pkhMUkshVwkcF3yaE333b+J50vzjJPiQ0RHqd0qd8h8eh9
T0YP9UZ3k50l0WDl1EO+NR1UU2abCu0yvueKxxUSfqm8NdVOMqv6w8pRh63GeLGK
FMMkKmOb65wWYTJ7WkVQ56PDHpM24c6ElhJsEUb3HZMRhUelwK63dIqT1Jdmx1XX
gwfcFfzZ0WrVeKMT/DCUG3+0Bll3NFBA3409hsdc5rTZq7rBGETT8e4O+XRTpWXM
YcmrsCRN8ETFxU2lf+F3g1jDaXjvqRGfy+/b+x9pYVlsZMuzZ/6TBRiQlpLGeHYv
NcDlqa4Rr0LEuJYan/CS0uCepVSwidIGrxnf+q6eaUMrvn7TcZlNTdUnMvTR27lS
FCeVv/jmOLUipBjBRSDpnNStX2LjpDf9jscFNGit7TpIAeXCgG5E6qFcExGHuf8J
BU3A2y9497/eJVUCakhc1O6jAUgnWTMGA1fmXI5m7G8KEqsq4yyoCbVt189+52qH
/+rsHlZbiXBd4Kqnu71IpqWp8wdIO1jLNKW/jiogDnV4EHoyngHVCaWsCqrEg85w
a7m4kd868avBiuBZvnYUjoKPTvRfdgDwq8UixHtso51x2AbQkulsJ69+nbaCyvJE
HKU1yvuoBvbaunTnXtVLlsn0Q4XZJwK9rINu0oezITeIUnlUzo7OixCG3UZizrK2
TyClxJfN8Z5/pkukqD9Flei5Mo/noMWtJg9MM9AA7S2CWLJYb/b/WpDLwxETVqZ7
yCMlRy7pnA2IOwQDSYvjz5U/ZE7rdBrjuJcJD1e6xvyansD4PE92X6FU0Lbnarfg
DUQdPrw6w2JFBYdrQOV/IO5m17XSTIqZE7KoxTgTtjG89w1gJ3+2u+/lhNbr4kSv
sVyFyRkJAcyCl/zg0GX1FJks1hjn/0+ruF9nMtfV8DrHw2teB4V4aSKilbiZzU5n
TDVvf7lkYUUC4yHN8MRue+14UU7k7UFb4m7VKHSGtQm94e3BoGBGNoHehMLGlUnb
ChJzW6F/wB2DAIDP7o0GmVWi4woC+y5sZQFFotwaMQgA5dJ/nuGR754yRAt0GNdB
okYPYUpwEFjx/i3PVX4FAuKdhftRrkDf9zYKaL98DVXvfo2upLT83o8cYegM3wqG
lP9UlzS+ad3O3CB8hw49RmWzfkqQ78FK0SpC4Pktj1CZjS9eDdtcCw1j8yAxCMrG
8VOm9CiIDE5ImgXXXFMjw+mh7jUbTJQDKoHyOOWWTDbqsWCUWOlUK+Edb8BWwMPS
rCPwaf0Wv1n/Y5IefaUS6VKttCfT62niZznWuPujJskiJ5D/5WsMNHvg1bV+wj3W
8XNFK4zm01+K/Ol/p1frEcWM1uZ5c13qeoJZ3p4eBXrMfz2cLwp29i+nsOejNjph
mfNxCuFFjfXy3jkDUDJzOKbFBaQNFra8JABWDFlhzjtD9vj8NrrAULB0cKwxNCYv
DxrLALBbe9Zd7IhTFJTdAUIdkR0YNd9mH3XQKaGR7Lf2wLQaMCQaS+KRPH1kV8IT
FJGUGjYX0vVYZCuAxA1qU9t5kxxMfnPVtIhgeXi5y0qvjuNTKKCBU7MxSD3SjUQf
Qk5so8lZlz3zp5shSRd766mY31Ulf1nzPh403gMGnCROH7WyR4fjuLLwNEloL/3a
eZWXFdHgW2x/zlIfrrsuH/pHLr48dgAnkYpd9phA8SPhAOlZQ9xR6zyOzg44Pcjc
+Bjc1z3OCJSPWzlpfsBL5ZXiFvegsZGzd8Q9zZGkUZPVxfSXE0MPjASkkvyoScFt
3KXPpUG1W9eY6qKLLxPJ3wqPwY5KjquCnMXptIEua2Yjr6ZUaH6e8Aa1Koxn61nj
hhnoBV+HiLrmBb7aR6nCffgCP48dwzml7cjCUu01N3zp6uqcZ2nwfHURZqYWH5xI
MCRlivDUNLigkzF5c73YTMr2xhOHct9DS6zn3UcUGzgDSnpjEYxd9RClJF60uBET
j9c7/B52r3+yiQ0WVh910qTd94XbniMk4R6C2KBuqMvGqLwIpMwmVoFBD8CeXCWQ
e9OnvGMZ9CCYFQOWbpUa1VMT8yxiWqee+RVDwj6xwl7lckakSBs/7pUTI5bdlx0Z
QY4kuGcW0t0aqyqp+fn2chXTZ+uO+6Q99x8UkEd7P4UwJ9EAFBBHyHIePj0b3GMW
qX3viFgaqr4F+wHhxbg5e9c5P+fjkoOjme/oanK5OUSEprjbfwIn13yKX+izFXeC
H/5iOvjOls+nOnwFWQF4AamF0SAdr9p9hghvjA3UilEFGFOfl2HNLO5F8QYTkbTg
aO9dtKsPFrukrb+ufPCo4ozwXwt1j7tMClVozITNHb4GuxkZEtAM/BpVAeSCPqI3
FhKuLazTN8pB6C9YPhFXL7VfZELrjZaGZ7HDD9TYukWCdIlcGb0JO0Q7eClIhu0R
5+gv07WRDE01sEKNvo0+1hulgyGKJ+UTkVKyoLcJD62yvf4qHAUZLQGSAT/7wIXt
TRDYdyfY5NGDPwFnzvvLvxgHV3nANpenXYWQC65o+WR/cQCxeqIQCzafyqWgAEWW
eHv1VolWadK8c3oi3V9umIzo8boauLpuIhsmKx53XDGWsUyhjRayJYt/YfMFW3ne
Qk+umGhVtf6oFkUkeU/oIdKkmwkZTIuqP4ZOhtOkRVLXd2Kw1z5KhexgRCdLbHgg
QsWr1N57PqesHmAxthl4UmOTxEGGPsbQQN9dTR0yApIaorNxVckCulj9mTVUT/2k
cR13PcLhyvd0Tv9Lyd+rqij0N6NJDL51gTdpERNzsklfCl59uy6dPBVD1llAGLMs
MWARSWwdff8JpQdi7pHvWbDfVVBG5S+LjWvDYLuzSZ6R8qPTylgSw/prakHRZbP8
dPghAWw2ABqfSTys1x3SpiDM+Nqje25Ngk+9Y5HCb3X2PR1fJEdgrqNcOta5loJ0
AcDuVio44G+dprzbHyZxg6qPc4Wa8El/IaIyg76pVeYH5d0aSpncmbuhrcz020W7
rghWjzAXkDsJjSqhJuMHdytyo4Y/anN8mANZ4zP+Tnl0ZvntzypEJUJYQP6plbrb
BfBOVYDHvSQizaEbFQy9fq3EplZt0yH2+LNEmDG5z3bp5PWFQ+IxmAEVLhQd7GA6
LBvQ0b6TPdexkFDy0s9e+2P0GwbXv8yRu+MCe1wWkPWixXH4u3lTpVnzmErlYP7y
2UseVMKHDyw6UzMesquMQ8nzZ+EGc8u/pBtonMIhULUGYwZdfDPPrhMmpV9k987O
MSIwrKUj17ZofAc3cotYbN7YZLG2TNyrfG7SjJdxPXY3DvWr4rlMWo4FuS8btSpg
0r0sUUdMykMSO7RYApHG3YPocgrObuu2sSwY/jodGy8n3wyNmYVLlGsBF/tNlbqE
NOFuQ3Nwf6a6+X4DTwPK1Ka9Cj2lo/gJaaJ5N+NVDW4Y+TvUo3LU0cIPFHFLfLGY
vfkp5HDBBfIl/axO5YZRiCgaDQ/+itIv3jeqY9Tgdhut9V4nWMWhTrLD2pVT65Fv
RuDU4LxlyVqgAy5hAbsSpr1CtZtNM8AK4q2YvJUmKOh1r1x03j2ot9k4zhrTU6Ur
BrUrGlCPuZi226uzPjsfeXL2tv0uTTL4D4IGNMhKVpBX3nYwMbtJWjbF4wirTGFX
2pkZJ6Hd7/oiRvGqbo6mSoClt1PTtcXe2Tyq/HzaHBzBZ+7I97q52RknMN/2ju2j
klxnj1cW1lC4V7FwVOA0HuuR/LFyt99eFP1U+k1x+7VLA6b3Mh98yKFLBFNVohcM
ti1xk78syRZacEORcC4763APwYHiA6pdKG3eaLmrLLF+C9+zkxQp6P+Qdt87JE0+
r7goSaA+4ZfK8ig4vDl/M+7ugX7OBi5BSpgJzksOhcferP+F+vvcL7eMGosvSUAX
Mmh3lt/gp5BN5/YGvk6B4TTstHt5WIUaoh/kLgIOOf34aRZFJvoDgaA9wZXCJmNB
U/PtK6vHqzPK1pk2XEjSMHQlgCTR1jFPeEjA4JcovmAv0HbIbe5DEaocaYj5iFoZ
ClUKGOl11f9OEAjQlf8PI/K24JSvqc4dd54y59V7gPoqqdxe05nHkeSA7s5OIi3G
Di0xqeGFASJTh+u9tazzOvRUNIB6vvbNcGYkZ4RbSSd+V8D0r8Ngl8xjLlfeujfg
b+ahSqwxnrx6MImyOhigFWUe+kYnjMy28Nm39Xq3+X//Mevv5YH40T9xeE84W9ef
grRBcybDAFLjE3R/GH5wcu90f/yERhWGNNh2DnoNQwG6rh/l6quJwr16CaBoSujd
+SE2nbgy5JLWijlGKqCbGX5BLty3AIvLEOaQUKmoPkb6wTb4NGfkVIlpX8z3P6jB
OrL+YvQYDrQrNAVS/ZrAlNm9MSfMogDfUU27Hec3Ilj+E05lt8IG8nWwVCJl+25u
cf9Om6BZXvfeIWn/0JvSJF3PxFd8ZPKlcyJMK2cegwABkMoemz936rShg5hH+ryv
OaFu1DCp06BKANZCBlAdzrPSpdMZbwGie/KILWVYxr3DaCw5tGxE9hIhcpq2lW9R
8kO+vlvGWEP8+L3SXVGEP8ZaKqsDoCL2+zViKRJ0c8gPOyrIGsz+QSRAwfGsIRZ1
E9ICy7PSS6jM4UrKZzsp7oBXLCLrKoLjTxlgchkSDeV3rXAZWX5dFce3B94+hmvI
v38lK+AZrmDgXjV7C1uLaE7ofIK+mABwr2v07lA9evXoA6Ks+XulI64WPvAUzBwl
8gzsbRQ72Jdk+Es4E09YvRE7uQqdebCgltdmiHF/U9SSFD1KRw703pjzqMrUIQnZ
pcs4EfAGWGCq63QzkYRpN7QsPOogA04aA3Bu1+k4nwquzTR4t0KqU0LEXwQNENzv
aqfni/Ai57wiLYsSA/nUQg+nob7JKPrCwDfntSyI4usR8uTlckWZjfc1/xUJKQJ+
Q3os+dSJQMLrS71qU7TqIGxG9n8IH/rIhpBJDM6OAGLUOoTbcnkOcIe5DllHFE65
/g9GFrp/+rQ2NrVo3TXaPuRFIR76qWIkdY5EtUhnfdC1utQT5A7bEnnuOD+9Qgdm
iQhQ/Axrh2V/5pq9xVlpPEkX9Mw3HsKsOLYtZ4GlLVj+4fX4hsVvOLrWS57CJh3+
hmuBnmgyoIQ/7aElw0SLI5/6lWeVSi9UIqS3byIewsCnNHQLQzLfVFj7xoKg2ltK
kIQAUlY3QjwOFqe6UQzrCGOG/H2h17m8IAM1OA1inV798jW266hfD4pxbZViXh39
OKRQVPW1dr3AZZdWWPCBqdL2dvZJIRx8xlMI29bhrWVlUx/pSxT79FKTKz/eScHN
+t2DIPLDKrml/ThUTvI2bfujPivib/T3kT4N845Dpy+VK9ytHG/CdKdxdRErXq4H
ZH0f/QFJ7TpSf89Srow+jYTwPiyWFWca9jMAxOp3I3VHEoYXke0tAjJUjHBGRk7K
TmrKO4VJ8aOa6U7gUUmDxHWoRzDLmf5Nysgf7RJfD2X/V6zxJ+FiiUgYYTqQAtvc
8u0vNn6KcSStij51QCaDs+puw/gWScgRwVICJAudQhJD7dqgKQDCtbck0ylheOqb
aezpCUS25FCEdhAxDxFFFNEnWXg4leJaRGooiug95A+ZteQuj1ewovT6iidef56W
0YRy7jEmqlTtwBgvXVK5eMvxae+Obbh3TRnOIEzTmQY/4LLeYwXGyoqJX7YuEuq3
IeWArCXAjWjzDSbl3LaSMlEU+v6vOrg4gHvO2FsbY5FyfkGIWV7wirJNx3rH/Z6E
UeF2s+3r+HQKsKodEqlCWzY0iguk3+YS7kDq9eb/3Fpwvcme7Kn5Z1x8iPQo1vTO
VxrNlTqDLNOYMG7ebggTSz3DrO4hTh7ha/JD2xPJ295NRp8vdleAYl68C7+Yj+iq
l8/6uU1baO/INPt2n8iYE3Wa/Xe4d477x8CYzOWQ00KPu1lLYmy+HY6lhUNoAzgA
IhUMbqUXvab+j7zYEitQNE607mIdUI3m5dN4JHnaxnrkgouw/4pc9Zd8fiGZFRMC
vTSmXfZ4E7XdSAyOMsZsQ3iYK1INqlouqrxtAes2F2qC5by/samnz0TJFsiJpS9f
l2WCTzcoWDWlolq1B3DOVn0qwoFaRVS+7qM9FPw2TaRblJRKaT9yLraC36hIgXWG
jSir7ISQihVYcy8VJXbbRDz5QV1N9hif+jtlsKnCLMw+7DJJifYb3idJQS8fa7BU
G3ps/2A3OHtD53+Ja5X4YT2PD5+OmACt85hHVYQddMJNckyAJ0U72moNev/keR3b
OTNfT+vMjx4tLEo4egb0vs0VOqCJxksViPyUN9WJ//GCaiNPIV0l9uafMKdSH/aA
0XaXirmqnc8F08ZE0UW77dQlcBdFNnzjsivPkBp1pq9KpQ+1DYVU4p2tbgJZeV2c
Gnksro9A9lyZQ2y3o3pk5wRsKxvxAV4N9UtvSym6UaTD0jXrXa/BDIgnrsxB7yiC
DX/kfl0R0O2NIGvnnevXELE5HiSmheqjL3la2LrURh1oTb92viSq80Ky3kytfQLP
sUuzJRiyfYPkczYPJi4ixiNnAFlwbyBtjLSdaHLpC8yAhPqSedd7kX9IlbkrNO6o
5Hv3RZeCx1/cSweGfqieZCDm7vUCdUMY7MxzTavSOz0rKu9tqaDdnAhv+M2lwZyi
4QoAd2yZbIobU6RrrAdb3bCr2RBQrj0DN0/llVmHorCJ/8tJPi59ZW8WGc+c72Xc
eUsY4IvOOb3dl4FeGSH4mZ3C1qoGdpDFrodE1jwRVOgXbaUvdwN6NS6yQMUER7/5
HxUBY/nxfoPKHUfl9RurURYGlHB5GxjAj9FAi804OKzCqcpcmuPN+xL8vnXnd+Ls
39vhRmZ11ogU8/7EW3Iwc6zv6PpD2m1zXboipOjwVbosd1u1ZnMuyGIt6OiQv6Yi
8SKtxll2xfjN/llN358jaeBpAH3by+6V3BtB62Y9QO6xrP1g+j29T7FitTg+8zQR
NyjGohcCnFUrt/kEg44F0Q8XLY+DFQ+1bR4mLa7Yk/JqwAIdPmDHMCzTXPvsasFI
ZYQu5pRaNiXQPVadPn6ndKlCJSCueOWcl+XVnTN42rhJ8OoHrF/k5mBCIu1UQYT7
R45BeRELX+UrExKyCyC6c41AoeBIrQVJ8Q90cLI+4/t/hW89qc8Ih6+lJ6WXp5Nw
kNlMJXXhfhDzHOzNltLcKMnwMorC4OaGEaYpOGk6qLCoWS1cKZ9t6cq0l+QKFliz
vgnmJdvPJra61QUGNQtwR/pYoyR5Cp17XXbY0T6Jh0HDxL4DALEvjNHyLa+Zhk5O
cbJsL7sIyWN332M1I7eM7yeL6iVuLWWbqvMTef+5bHQgRBh9xLNNdA1dt+EFDl+O
fudKEOwX0lg6Q0zhwoHG2FYVBigJkg6WpsTv3/l2Zq/V/5BMZPfTDGAOJHE6QrhQ
cIihiy6x6yNzSgoXGvJ+9/8GcZltVF3v6AnrxP8VjWv9aoEQbOh/rbPave4avQmO
Aknmg4GTkFgBjMgM7Bqdo/y2PBBvFRuD0b2kZRq1HYQZMVgsRnMskYGOOREqj7aP
AQGWUxvVdgqEDZOiMdqWARlDIbr19WDc/XX0S1QCEO8mGvluzqZ7xpYDGl7Jc+MS
4KA0Tx7ZoZzbfn4j2TrKf5y7pglQZtejML+5U230VsatJk3ROGqRWcs9GFiMRZqI
OnWZwwtakwQiQK1nvPughIAxZIzw1UnXefoT7zo2I+ZNcprhrUU3hmb6sbdliTKR
ZCjXTEmiz8YRAllIqme7jo2ewCdEKvBFi4qZK04XIQ5ZPo+wX9aeV6TbNg0WPinp
/2c6FqMDptgnNFfpIl+ppd5UG+sHWCvuvUUF0qPauz96qrLZaMeILfodY1Qg83SO
Tx2gQ9HhesDMveDZVZwIsQeTxWXJrPVmQDeRX4ZJa+LYKLc1E9m+9KYlXknS5uPR
/nvX1EAEN61G6fk2OBLIS25Vkaeu3OMVhWyEbogJXeWeRQP676XzXBAAL1K8P7jX
eybKuda6Kf3eeQGVmF0tPYmC7SR6b9e+caVH1mfcqGFb7J8GXxsCHDETWx2lJVyr
vrGggg5kpd6UBghdAAzeye7Y212D1pfUspypzV0U/EBCqlOzkOL7tSXO1/3mm9wq
fJ4sl8FA2Fb5HIWrfiKShnjzQapnFjHvMoTx2vX1GYFC6rIsF7baygqMN3z4VByQ
n+a5eSbNlPKvoZrZmC5Xpy5qkrVreheYaprYU91FqwyvVtD4EoFuFWdt2WIwzs+H
lxFjEj+2N8+4yp7iNshQLKr5C4s2pkyLaXrde3Y6swj51V6rucl1YtT0A97d+2Pa
uCU2bAn76YxLglGSTeZRhyL3MQom/1Q/k6yFsO61Rdnl3gvqgjwJi0AuZHvXdN7d
1ZrSCW9Ujq4m9BxX/aeH4xCMOGMqDCZJbD1S+ASnm2CxVcX09cZZL5GpcuQuspua
0O6NBihs2e54LeJp0FMl5ZjDcAIxrYUD8QPbpBbi411w3RGv4C882QJD4ZGU/J74
C7O+3JiJb4l9imiagdAJ/QbHOFa6rbjAmMQoAd4E4pgGRQ9aGgKBz3gxI+nEdoK8
GL0f2LthFS2j/exOQXzv8qbRVMjgehE4HGXRJk3YnylxZCC46m2ZQMdeWgMKgD4E
tw+5+NAM8YYkyv/Y5BbRVQUfP6s9LzztE9ESVQt6Uq0HO7s+aYCg4v0ho3df1Yc1
S3gaoxHz3ymyOP+3z67johBRD5FjsdC3sEJN9NUTWLk71MVmhTz6AhrLG+a4frTQ
bkfpwm6KDQG877bmfsAFmy1ncEIWWiffzeid66mGWLrAehSk3O1AqGpL05KxIoRG
7wXuoI0R1ZlvQHG/d5078ftjiCNY5d2CM4h5yFkbV+LRgFiK1tblxyUzwLO4eXEU
AbF+JmZ0+7k57M4f5cFpXwrnRQm3COGbDNpHgyeg1d9cqvTfBvx7QjfgXJXzJGvu
Pp5OVkyggA9SLDX+N06PQV1GPrDY9QQgmFc10f02jw8NU8hWJRNFEtsoGByYfroL
fEuTdpTHHO2vdugy/OEW2wlgsH90dBnJnRzD5MZ4eo0o7EZ5ndk/wAkYnqvPelFV
TBNinTpM+NFso/41wtJl3LwhOQP2pWYNUXZKoPatpqejJpRGkXceeP7UKhsNhdWm
qFAPRr6f0wHnk0h0+Mr5gULGDwjCBcJE6OI66AkzwYg0K9XxVV8NpzxwaE/qkN9T
Vjm5jHOc8z1vbAMb6DeEM6HisP52JqjXggGK6EHk1ZyzUCqvBJAgcVF7/eoJTzcp
zwaaZKhrSoS1UmtdQfwejFHMbMgbpUI+17RfDo8jtd8WhEi3wBPCRJSeXYhspR2U
9u/2jjom+vjPmnsWmHl85dXrs75+ZYOczKsLt+RfsIBo4uOfX2IujL39VmIHiha3
XeskV+CPfDMImgJ/bfQHLgLIDoTZDSl7O48IwWy+je3NttrhqBYe8GHBcpvE07tk
biVAtBKFJ82NYR0q2/Sj5hPnaZPg6ubjBpLyMzagYTkCumiq7/MJhT2FGd7pSKvo
raJp0mAsSWNld6bOCuRzggtl/NC1dCSqJ3vkDLnK+n6oC8qrZ0xac24gPaoyTkcd
1f87ILYu+fntDWJh9uCv2bpy6LyYldS22JPvph/DnB2SqVWlYQ/8iZ5+BqBV6n0O
LdpQ18SheT1VzZ1aiKJCz4jl1H6s92mcSz2cXs86BLgX57JtLT8nk4pUCJMtuBE2
aOuASYTk3iCmhsby1TInNDax/BEl/XN1jfgLM+hJUpJBEMNBtHl24twgDgdhth8e
0Jx8a2axggsbihy8KofbO3APEhkCIYIx7g4rQfSsPcLGQo+P0FvlP7tTcV6YJGSk
Y7hDoAjTNUK3u5R0lioXIcOmUT4Bz9bN5MOmPofxfchtt2wImXSL6Cyj0XYQG/MJ
ZyTyJoSSPfEZ22h6sgXa6FOwgR279xaES7g9/170/KRVApy1eybeeG8ZGPTXAQvx
HMUi3N94aD6hZzGCO1UgxUDooLoiavmtsMCRkOJ4VweuveJifL3XhONS355feY4g
hwKJPDnMwPi0xOcGNVZsitAXF7OsAGtxT+4NnRaw+ydoOYDkceGlOSw+/8fP771E
fQyeK2LzPlHwkvNmK7O2/j1J1LIeIH4gT/rUsnimePihlsSoWoLEQb+gOPhYZRf3
iB3d0h4nDbbre4gyGOtDR8LVBEoPaGYsFGMjLPiNsW2DOA6aSdddA2Ox+2aMeTTP
/LpW4NOgutFUgbORMviLouNjtwNIKFlt6TDyCFc7kgt9k2G2/VFgiutSvf7kNXMP
jEWD6850xEh7bIvhPOa9rWtuZDfMlJ29TPytm0iXsPK5jSWJ1cSlwwft5h8po9Cy
MdsNUFTpLVYsWpwBwetNeUBHG5GpYg70u7ikA6j784Nz1jIq2o5WDDlWkt5blNKL
iv0kFrP78aZxP+pVPu9CBMHl7fsQ3XGh8pzPrEINfrOgsD/gcKmJ5W+jcLjoPl9V
blG3njR8jBUNZrKDKa7S2qUsqhW6e9msb3oxSTHabyUZrHW4eCBpmCDlAYNqXph4
ZpCC6PSXEza2PD+RALLJh3ZQ6kACkyWllq8MllBT7kOLqmOPfBqIyEdV5UxW9lke
qvkdEcu6R3sIAmUKH9GKlmiOvBs7AdBh4x7vayDcNgZgAYLuATNHGZTyqyR4cG7P
a7Ex+6zG+/2uPU1S00n9j+KRM9jV9fRB1US9yjHncMF/6ZKAmcdbisacbtiua+62
vL4dd9Qix7Yl1MYX//fg3pPdrjgg/5LYIragedANsVKoG9eAxJkqR2Hdw6tYRSSa
iVZA+RP590TlA4d4PfDlXtja5b9U71RlCCwT44Kamne8dVeiDfvHD6Y6h/Qnzbpz
h5PWNgCD3kccoFGra0yRKv3XQbUS/5dqHGv1UxyI4hBWSqJFUfx6IBZv0zL+DX0K
Cd3pdwJsTzqp4/BLaZerP8OSmueYg9r+bo4Daeia7lB2JykxoT/ybDF7JG8kfR+Y
Rx5mnoxfSWP0R6NNLhBSKe7poZSkAUpVr9/Joj4CHfxFaZBeu2hN3Hplf++mZeB1
sH4JQ+B+7WMSMgguEKwV3OGNJrTRm+XdWWie4UacVhm5zWpKpWsSs9JKegs/cRWC
7pyjpZwZxMhbO8q2X84A6OtzG3ZJkrbCWwADyOVO33sqI7NwSwF7XlgUdvcviGNn
vs96P9oUUnlCspw0lHzvHZ9uRKf4ZgyIoX3JHBq5jUtPh14pYf1YM+Yk3Bk4PhHh
C593uvqDCm//td76gCAFVnI6ABDd5w2oqPsa6Fb/21XTYAd+dsbyEnIC5oi6pgoH
UBje7X89YH31hjzOet0bNAmpXyNYFGCReuwxiu5+rx5TBUh540JIN17r2cyiLp5f
umCaz0EDewwUt2eVqYvskGEDdli/VH/oKUQXxdv8NJorkjPc0I0ioh/RQZ17s4Bd
cjQsGxr+jQ4Yd2kVKK87ixYk1oV/0n0jQlSmkQ8ezr4bP318bx30W6FkAupA5Sff
p4ipEhRBhEMc6w6rqiFDmlRP5e5DAF4RSt972LplO2zhKD4B5g+JYTmoUFnDbLCG
0IDtHH1R1zOKxF/LM01MCPcJhg64biUQq4FAKvVILsVDvwjeqvnN6pgMGczsQwuZ
Gmn9U5/HDUrrvTEGj53Fi2r31T77YRynu/OKTtAD3mkW2fSFz5o1qqVK46t4g8ic
5cNt9sp7DB4DpY5JcTkXP00L142n6ssFkjprZsXmzchJ0mwFEHqQI5Hv0SPoK9fP
1ygVlXuhRrpQ74lmRXjn6N7pzbiFYx4GKqpKCIJpzJJlx1IzhbtYvLvszjH1wti0
FdagPL24g07edTn3QVqw+CQ5Nc5pS2OTtsULBc2y2ri8Hc5xZHaMwTRpFBknRvYY
kLRwmPX5KmPZjEAtMCSgWlFZAML81s1/I2gl9SFR/lNGJmiQGT/D817U74aTO9ov
14I7xJZHo7LZ6eWGYq0YBdtjUoDvVHf2EPKPZtAFzK4Nq1dBLuE2vCyOCjkhyn+N
dwYsNjGZhnJ6f9xBy6UJvbUxTGamWjc+I8b0TKrQ+vhs8BzrlORg0z+bq/OvjhKm
Omz9nIOo38I307t8tLUwllnroGGJRWpX+M0sf5L8yTndG4l1ogeEOn2e8yYuf96g
EwGEn6ByP+LrEMMKZh31NIsl1TUO4qz3nNu5emFSwsVG19m9h5djUrYpEmveVu+A
kPSSHmRMb48BNPEkkEGV7+R2lu+p8mremGJ3Pv1HI31LJs00ZOb9ntiXMEvJ8AdW
4R5P3BE8pfuaXLOIQdWg71IL4oX2Et/s9Fenm9MDWdrUjspQdl/EX5Ryga19W2ut
9okTczlvY6Ej/uBDhGcfy/KwJiMEiby6LAWefkt6nuMtx1+sQRRnfQnRQI+t5bOm
6N/+3FFc/jiDNe+3KJNNvZwsGMJGbXGrgBF7/Ij2Lxz+GytiWfRh/q1vEhL9R8EF
KJnlKDZSyFGgB2iOSLbQhSAyhzWLam6UFowc1lP0T2fcHdbvpXpluX76KZLU60Bs
IaB2lm1Fu6HvByPljnONAL09zXFFsx+sMQW+avysEFjesi309HugB0iK6+Gkxn7W
1aBl/dqAVkl14FtgwquzYAMf/SiKSctif9KW3or2FTuvIybXod+bCoqCluIwqBxs
Cz4SQfLPRJc1774QVcG0g5IhyvJxhg7e18Y/scjn0UUOYq4gc4M0QZpNZkwqBH56
q42H3la/YVTnTBtI/f5xbWmA3d5Js/lmnIJRUG8G1o+vRefCsdNsqHqJRBt+jBuH
vLyky6PO7P417k/NsL1LreJYaxrhlzG1DxTVVJrvQE5fAOTL2CA3wMSpZfNj9axe
FN+Ol9/td0nV8QdoE0talPInbpXmDHC37OloVqngGU1dOofGGreOUvUP/IyxNegg
sgjt8mRJWoxwtCAEjsKxwEkGU6IkddM8DzF7d65eBsMDv0kVwb1Ra0e/0vj7iinI
vyRxDlL+mDjJkExRoSjYSfqOePgr8Ss1QBkJaFTNqenBtL0IqUI3LDwoeo6DzwA3
16Xy2hGC+7juTyEaUg4fjM8TMCtRR3vxG27OuvQ9ZiTc2/UzI+v+3ttw5ZkFUYtO
fPa0I2PBufavCXkGUlscu2M8r4bz70HPjWMn5lSVGBkp84llFux7sP1ngyyAb4Fb
l+A3bZHsMRBMHTdX2AEax1JwPn8poTGYtdoIy1HD4LWBdvdqmIvUb2q4vmI9TgX7
glWE8oV7iYvY26VzS0cs/a1zNs2WiwVnrAnRl/ZcA74i0UZEHudkQE2HXGjmojrR
URWSvax8lTrjYS+QpEx1E2CMSmEmBLgGb8K7PCmYS+0MO9dna458u8eQVSt3lQFL
vQEVQ0/LS7oWop6+9BW40CaczeVYvjVao8EyS2TOfzAOTyY9bNsxa+Z121afdhth
NB9a2zYn0rRk1XQQ95FS4tdZ0mk75i8H240VjFx7igqA/F9wrfyZzNYwm1z83hqe
m4aMGL8n/QMK6tv7W/ZoHL8JawtKNM8dby6a0ObQXSVv1/YNK4+jk+rexJIBARA6
TT2/xSSRzQGhxTfTHo/gxjvqOi8I6ssj6VLoAs/p5GnZc7y+8TouhTlIBg3hIWiY
1BIxpDJLeKLX4+geNe9J6NCcf4Asug+xD6+jSm62vJdoHcIt3BOHfVYqRclFgd3H
0M7uaUeg3CSEdVbLVRAIABpyjTevY5ZGlrqq8WPDtjBZq28Iu1w4tcxtofTo1xFi
Q8/3rWzzrySHXtvtrZe3Rk4AC/cat7zi58Qca38XnHx34iIonU9CanmzVGUBeI2O
IPOEw5InrFbK+W5LIFfmV3RE1En+UE4iaje3XawhpDLB5abAlP5MTVohug4iyrwB
XAmF3lSZr4tSP0QezsABubtv3vJdMGiObuFl190RFXnAFGg0n6bfE3A4MIeZ7I5M
tBHQkXn16ZdNyKJe9iEfhAcPMGzFkFCA7gVrbsldTGL96Ovts5SGo8eDO2Qp5HI7
oSfBiPgCV1neDg1FcaUbpM4rmbkMDzRtSOpUhH6q46O2sTQ7452fHyvuSWu8RBQ5
fwWjOuSvqkr0n2R0upQIE4WpaP9Jb9o5VhjkHlbQzjgEauBZGHA+mZSsLUBrxtOy
uvCvw5BJsTNAdyka9cOpNkxIdAwVMEpE4vV2Y6s0TJYjCDXHSsnPNsQDFJDmJzdM
v38KwhZLrkBru9TAnebBngyXuadoX3QIPkFeazHWrgBAlgzi1+1rzYBHv8f8cM1k
8AIB41zZ/X7Pfzru/rOTvNgA8YnQrp5fsWlCzrDn2pgXugtF6bE5qMSn5le0PjYq
dgnZBcsOY31/4gwCNBIxw9mOV91vrwydbOsKs/eIr2CqwnUtqZ7gnVNyPmxy9y+x
8+tuNi6WPp5AVlFtpjLG+22ExWXMka9Sm7sbThNI6meyovdnZP//4Pks+i3yzEiO
+5wuLTsDCbdwykxblLteSFqeN3ZppN0K4H8MPeePmJ38YkkmLwU3ytzZbfosUWK+
RGSPWc4NLDmuDdayl3zXtjxkaWt+16Rc0QTS6Dtjz513Pn9EHnj1an5eY6zMwunP
B3X32v76mcb0pLolH4tHlwl7j69kEHkkfXa0gepUnjT2cRdJ2Pg+4nn65PvI3dO1
30STwpFk4HLe6fIsOI3izxz75nKU4qfcNfplaciuj+GAW4CF3YuOaPUwYoQnRMEE
AD1//PIJckvXTUI5+0WEqzN/ezcR9zasXMle57wsDsBYZrjVT6VJpawpLb+bsn0L
T6aE63ChWx2TVofvo1IEtySH/acCiWUdRJBx3YS5jFZ3aYO6b8AnOyZYfUHHeknj
puJbC8sNRuVsxr0REmiYhtoYSzcBtvYFG6014NwxMi6q1pRBFLLXlgNsnxNjCzw2
6GtAOiIlx38MC9utW9FaLhg+N/uH8k2sQHnXe60Ffk0oketc1YSTkib/MxqaKxH0
EE7QiV4QqXhA6Y3To4Qo9i12dTutJ79hIjrG9tWGfIXRM98aDjwGmXEmaa9G2r0h
yf5LH2P+JDK+p2jfrPopfVqJYnMTxjipn1husYLln/Lc9BaPz9fLHkl1OLS/fTS8
3iFOl03yM9sd/FNgSVzIIUyU/P25tJvctOEEgX2kysAwfSNpADgcX1OjqmnOnUEF
a85wS0J8RErxIczRCkBX1W/nEYkUfHkHj2sXGEBodroiANT/H+eu9AR/D/lkeVyI
6rNBv3B0YpSv56tf/CCAfTfnOGS5Q1oT1/JW2IzF+r/sZUXNvF7ay5pNWHr51Fgy
wXxCVucFHV6u5jerCK7OdAlsTpurtUiU2pScxk7+4OKzUMJC6mgVwQXsljAwW7af
zh8FUvJgNiVNkE4qYxDHRuBnU6P5DTM2E0wkdbycXI2TPTXxErwawn/n3n95H7wL
dE/5AUJtTY+6Ta1miGEBXxuysREoOynGGN7QJMBOmhFO/6agsfpE2xz9VAt/6THv
9zSVYgFI2UnN0Ig7OvqbWQN+ygiHl9j1YmU51Fx5hV0nteOWb2HzE2503XOmTf6P
TcysOWJyje1dQYbJ2326PDisLGwEMZfAaiuyQsDNHGmnNWFuF0vS6Z6Cc9IIuQcw
uXx5Mm4MGdrIMYJ2xGDasNkUumCS0SeG9stKwtFeByoAu6dQNKE69wGRLXtOzK6g
0DJpp8EtTdZ/oRYzSjqoc1XIwpzFVYJjcaaXxIrb6o7JIuhXOktWVBhwf5tX7uaH
zLl4WP86n8YAhG+7FCMfF+OF2Caj3JJTKdsynJzOCGHiJFPTsqsDhhZxA30ujAh1
rVwXCij5+KUaDPuLt7cCkdZ8sNoILbdOmOwxB9c0zYtc0FpP3q4aKHb5WDUkFeFY
WwhPmzoLCKg9YN502rW33FOxz8rBnIVtupQEMC79moLDP3L2atbiJiiFu0cFoP3X
mqXdabYvB3gLgnDJE97ruc5pVPOCu95fVeL5NC5C/1NVn9f9Ps1BFwGf/ir+2xAW
+hdN2ajz0K7l8Hry1tiLXhb2lDlEIIrkofQEhk59m3M0W/mm6jFEGs1Qsdu9QXPv
9oKJsnYNrt3hvEaB5iDiMGL/sMV0SdUrOUXLEMVTfNwShj/BJlCFhmEWCfUvljez
u45xKAYa91YA68fVhnfZggn+1kLRB1Bnkl0Jo1TR4MRe/qO+HHGpuzAbrOdVOdOW
jnsl2GRSmYr3QtwpqMLVMtG+zBqrK/Tjm+cJjJ3/JUbTRABIxtjKjWallqIF+4sf
km+LpWTe/I6FkRkVslNAw3UBzvzRv0oLVvVcZd/ui7NqDV89p0imaLr0HXwSLro+
/FxKVL6A5egHAghProzqfYvkM3M3tmAY58lgGeknZFfhkpZgP3qHjSljOZa3NQB+
t+sxesAzvRUW0kRqVfigJ7HbYqIynLor3DXPV9afeThJpgPNjKpA5TJ+lZvO66fS
V+2M5vUUU7m2Hsd5p79IHyubd9k5gxJMD5vd+Da9MehMcWid4BCA83ikar1xvhvW
YA9iXPn2DQe8P78BJtL5AOsIKo0D+KgS1ZWVmWKm/bo3xee6jmN16aIs+ZyebQ9y
y9ULY9qyx7nuJ97hNj9mlAEt9IOVV7HjEMInf25kLCkXXM0sX03dnYKUjDty29fZ
dg3ZNy0rk/BzRXWiMjPb1pYFPL4crw1RIwo2JEWabr6x2Kk/hR8ibRtB35c61BBi
TRtLWNW1xLsgnJ/lQ59cmNrPdXYBrUHzUwOgwIJ0iPv9seE4/m2MGLiySZDshxaq
1yB5s25cDrebm3c01hzH6bmsLYMzfKQF7xmG6NGK3BpECoqSEqXNLMylLoI4PGx0
axDLwdWiZg6NvDmYaParY6s60I4vqxy9AvfJSYBotP5V6Vii4g4mrARDq/VY3yQX
sulLEbjdA8yRcpY7DYhuyRoIgJA/RIhUDvasxffVQvX/W5/ZtKomD2EmaDfT6eol
hzMS8QbLrIbrTyOK1PkViatyFHSSNoC3ayUrcO0n1AoKH+dos/laao8VKZ+gi29N
CmhyNiNnRn9tm59lyUIHCoT2mXonyiUSGnPdJvV1ThJpPZUrNPCkoPK95S1PW7dv
MTjZdssI25/acueB82CmdQvB6p0Pj0eA5kKzU5R6iPMBA8WeNWG0a2QCNFSsZApv
CKmnLQhuco7+kT05tEnWlhQfQ0WkiDCbzIby5DBaN5MXifiICILmHnAS+jpy1A3K
bENYqj7Ve8VNHuyNL42LThRtssTsjAUdZtmEURmuCNa1xJM2xKNJfctKmPs78lBb
MrK1QxCNzj08C5O6CMbnJCzHAR77j96HRnFmjAxtIYjPfWH4RNee5eazmJKCY8p4
QGXTvAIvhmUizsGefY0WXrIdllswdZgqe7DWmBfTCGMThrgB1+AE9kQ4gIhPA9ji
Emoebc86DNyk6Pg8w1DAVnCnBW8By+Qj2YtgCZgn0cXOaJaSprooqM/6NvQgMwZz
hnbKdhaIXv0ug0EdglmtNJYNIm5liFQgjE4I0KkutWCvFBHZbSfEeypWfA176xpl
odF/MRTKAYvffFUrherokZqk1lqqb7YUqitvazkcOxR0iowceQzy1veDUTXKVPd7
Itk7OW7GuHfDNdeAWmd8vLUyL6wZFiyJoIaa9LEi+2fUiL5MJoTcqdx7AVnJ7Bge
MXuTF974FYznY6dX31x0p5SXtCaglIVOBFIJv+WP5Va5ARSY9mnFiTZ67nr4U6xw
tvqS8UBCQgswWnlocLlvqfaCBEMeop+ChYZvw/h6Kf5mjqOWNQIy7V5fp+knVpBA
tOWCsUdQLQVDByYn2an46yJ/DvfzQex/AZUSkYjUjHEGrpC6KdKgiIgpNNUVZngH
QxyA10U6Z8XFKo2q//U5PjH2exDsQmcPBtbrGoDbwF3guN8d4YF8tmYDBFPhtoR8
hLrwXRLcxFaeAiCivwgBl7zpcygCIcTGaGAPOkdtXK5d1QvL3EbnNoMOk7h3OaY+
YjHVXL4HiBuIMX1ZUa2T9Sy+OsLe9YnYhwbfl6zLXiBMHx95k9GiptrMOD6SPPsT
TcywI1e81UeGSQpe1GUejdphz2K6hzInNbqv95pe2KwE/cCuzUv4xzGsjStIwuYc
bZLGrzLggpx5HRKHQeXmqEaWlpl1LM5T/QuXfK69tczEH0Jv1MIIu1WRs/3lkOg9
gcU5hw2Y/xkRQ5lo3LiZXPEpKGdyKsrDqQOGBObPcui/Q36dN7hKrKJxMx5R6GtL
WRXUMGHoEFqE/WJzxyVi+UkHZlsGDVxYJepEcyBupKYkYjmrzS3VeXcjJUiqpKLF
QOAU4Sl3+AHYk1+Q6q2Wrf6KLV4TUbWfprh59U2fFY2XN+A0zHSj+qxW1beYIW0X
tIdaSBEdoYFgRLeHfaODEDYSOVhU4Nlmy5aks/a8CBHrALF3tc6VYUU3bO8Yxd2h
oVxIEXybpW2i/yOMY9A7aDZrK+K2C0aDbSYKvxdLHsDo7Dhu8nF5qe6TIJhdrg8l
qSjOBTwikJHJLmbXb/onW9QoGXwjWVXuccUgzu7YjIlhOP+He5mnjYyKQibBfpQa
TdfaL481FFtMg52h0VkshshlZulKWhzGei6/gUWNNE/npx75cDVu9mktpv24CaYB
Iefz/46ldxLen9wwLyfExoK2Irsmz4ytfvUCj2sFJKXM1wpLKoY1m2dsyQh67OIU
oUQi9NZumoCrG6rZ92easx41xX5eJt613mFPE25OUan4K/zXsh2wq62C7LY8+xKT
mdlOHTWDhm5Zn+ihT0qj//xY9nnbhmKL45rbn4ohIXDNEDzJeYf84tiEwDi6FFX9
RtHCbMqoSWbMcpMZT40BT83Iq9DDO7kZoCwCADIFuhal6td7+TCVwkCGkfWojkKG
rDowFGyPHcO/4B6KqcREs4iBDC+UAQcVYPOjSBHb7tH/s0MNHeonRKCZGPF1dIFj
bqnuzzMrDMZVKobqMzhL5bS7lPvOirfV3ip4fcrRQlrj/Z8QDJ84iZ3vqG3FxmYe
7pqiERkjYItWeZzA+7GMmSTuBg7G7jx44dhdvRIFpDFoWAhVAM6B8hdJwtkLNCYJ
pCth711iz+dvnOW9N6OnCKN/PPGMmYbsER4SxYhC3NZ91tJ78jHYKiEcDMtAs0rU
xUhZVsUReSL23SVqH/bOZMqOz/0cK4JRkWQelomraIFJjaU1h6E/VCQPrrzcJG7R
KSq3gFKIYHRy4uXy6uvwTjeJrMHDN6Azj5Z1eTLK88QJf14uJyhzPpaSw0G5SabM
elWBuDHi+PfxWt9MHMq75WZoTWDVt6VZLcLIB7WkchPQASKoNAFl+rKqo0zUNWSK
Vseab2UymKEEcr/SrcX1+4UD2tnoV5ac40ues+Y6pgsKdl/77eJFpq2gBWB4DBvn
zo2eA0FlsNxlTXcN50Zy12c2LjeWjhlwSGWKQyys1xLOFavxQdzc4LID78ZUbz5c
dZCwwL8dNC8kZtfRbTBvZy30b/2UKMG1R6NLtxbHSC8FY1ekBsrMaCMMXtJW61YR
QxQMro4YWm7EnMvLdoR98097Vuhhr8+Oghz3tVWSt60/iQ+FdZCapi0js67tBbHh
Ezx7AgPMlVKALsDJy24wwgTD//LGfdJt5IsgNLJ8jl0b7rjIW6TCbARZP4AyLLjZ
WNorC/gNYe59U8CybfuatOmPOD57oDzE5sfzBiS4eiDzm08Ucruv6lS8f8lJXfR7
qv1SVpIUzFFTehWpwhCqiTuiv7eEm7E1i9iMkByonBlstxFp4/KPhWNCWPygQBb3
g7kaLvKvjCIyRk7qJ9m3xkuNlKsb5/jMOBwDJVvXvPwHziJ8QeeBEnbL9J16mV0b
Mco3RM8gXz0oF/D19mhriGX55wjXkd8wJ9oQQLLhOBfc0A/6uC7crnddv5P1ChP1
0iVNZAfwlYecE6bFHzBrwF6C+Nr8CniwBXAVPZ6/53r3g9ht8pllRYXNQp/o5UjR
tWl5GbpGPk9HU2i6jg7jwJ6fi0qj6b55hQjG6ecUXOJ5Ap2+b957bdQ9jeKFO8aG
LRQsfdvaNQUQZ3YvzAK7r8sdr8M8ogpLxhqca/q2k57rO+dBvfWlK6Pj3sx1UfBL
r6Cipnl9DHYlxRVynyZUhHazOPRF6c1dyUvTmVnEWupKm9Isg+mAhcn7Eng/WaUf
CUh3/c0ov32UmKvvzBETI5hnOH5uGLsenTUnVS5on2owZJ0PN/Rt4ZXWWjV6qeQr
nTBVZh7rj115auY8hklyStgFLvTxJ4F1w85e08SmTnULzLkwrP4h/n2u1lAnUuFX
5r2KiAE0nbTQb0hERz036eC3+8flDmOaAH/qK+HOWpS5jYNZKdu6SWufhOcITmTo
R4eqvXhyr3fEtok1ZmrQhXDgIhvlFMIl2171/b8o7Jkh5LzGPXtD1sA1FkHntLS1
Ag8DKITWpDBhFBPCm0FE+qu/Dc3CsQ0WRgJynnZuqrHtCXdL34ZtrXUK6Yf9hUS9
u0RKF2XbGVAgVfXDbegM0oY+pyfMMfuw/LfC7dwBg8USbpf7psfO2T65w7Vhofju
QQKVfcPzQOLp+TCkh99oc/3OPXOqLr7j5VP3WXNRO3CR8JzXMT44ABn91YIyjfA4
wGYB/dwZv1RJ+LGVaPe+IsRDOMolPcADn/XlLuh/L66dyS1B8XJSwx5sdm0ATe76
/7DmcMeqZ+G3OZSqM8s5ZewOgChD0xrCMZh305N+ygVY6u+cXStNdldYNevZvwQ6
zCtdB2EJf/+agxx9GEeDFRkwAmgZXEYao46dLp7V4TIsikEd+1bBc5Ad5tyT0Stj
M+DYcqtHdr1dOCt/hG5wox4KMF98g2crez87ROObVuzk9zUn4/j78Ic37wW41wS/
xwyNbUU2jO+CesO2LrTMwvipJSe36S711zQsNg7ZHPT67IXirR6vT/ggTNU0+FiX
7N3j1hTFhg/FA0l+eqJVvp9iqf2nASI9UXaHZ/V2rQdWuTrUSUhhQnzUDxJnOKQY
JJ9iSqNzZNfoWb26OsmRz5gpSS6dsk0qNciiRTzGXRaGOloinfaq/uiQN3epK61d
ccqAROt/9smml8hTWY2J24HGUyvEHpDoD4Wruwdq/uraa9e5WSnAbfHvyoCtLMlT
6Wp3vwb8bSuxrbycMB0r3Xk6WlnLhvbNsQmWNEFwGouk2nuCfEkBk3FdFo0s5NKu
mQCTfXiYHjz2C3IfCutqTm0gDcQqWNSKNBPzu130zo5H+mgPQRHojynTfzidNnOx
6yl4wCJcQ18eJ01glhNquv1Hj0OhWnJ9PPZwIpldiGE1Sv9JsmOs802eG7LXOAB2
tdIshJS4qjlEZXSF+7TRb2BnpXuYu4CgMyiGqiP43PkRfOscSltHL4mp9zrujVIs
x9pMBjOal9TdgA5l3RqJfLG701jbDV3DzH8ZT05o24hFyavBeLcK8DeblpPFzsMG
zGQDAZcg0i/0rmiM/ewKBt9bctFo4ohAmJiN7sRZgvfEiEhORPk3rpXKO5UAWu1B
rueXS2Sb0HNaOvR6dPKqbWA6cIVU0WG+fc5Uy0HMdHxv2akC8F2d0csxKiJUTPNd
a/cYZL/3Vk/JtwGDoFfNc0x12OwCY0BvQuEV0L3rN5uaDyD1cS36jQkE263LD4J4
oFK1QPLIXNMsKquQWsrFwE31JQ2kEoLLskm0iqic0h1nNCiZIkeBkOOUEqN8l/Cx
wqjkBWtunSfVIgeZAqUMlmYGEJ0304+r19r4HtDfxjoaiHpomMuGRZLOqltP/2GA
vUPzcxuk6ohDpMtvlmfQcdxu1logE9OQhDI+tCchC9wUYJKJVTLcd37bGYl+Qhzn
UnfccYbCqqLvHIYbCK5zcgqWmh4ePpxQGjit8P/KOSwPgTW939uxa1TDJxiFjTMu
WtDECqU/EDa+E3R605PobFaT8vh8GyH4z30pjGOlUAhyHLD74bEFotkOGW92BzVA
vl42s8x4KxqB6np0F722CwaNuVDdsauoJGD2SEfj4aGQuLbxi/ZJMrAsx8AdaaAK
+C+korlJV+f0QoF8Ci+Ko2nua6O5zwPMD9XZLnA6IQd6HJ6cJoxM7Xp3v99NRHwU
iuxTvNtGPieCOqJZD8gUZF8CUt8tN43okrxH7BdeJlIO3Gr0W+uaGu0FFb1XXhti
ZYhXuaL5AFq+h6Vj5mic5DQxgMbHWFJLiHYCLtqGWgA/948gJe5tDPbB5IghJzK+
KKm2kip3PT5iRZ424eAa/HzRgwUcIWGyDjHxa8QOfWjmiW0BM+0J5uhzRu0e4hls
3apMRJhHWqpLk3pl+Z1IHydMjS8xZIdDjqo5CeNvGmzFuLBLwQU3E/2uCcWVrdf0
3E1AdYj5ea+AxJopyd/LX6nwT+Q9PRZvNPi8jUS887W+THT36lTaLksfwyfiFnqa
MxahDDAZ5EnW8k0gqXLHJaUwHRyTQvM4Onwm/fPdHXdaAyG9Z67/N66GVedH4cvD
8KaKmBDEpJzFBuVIfEej2133mZ9/FAUScg4ReT1pSMOeCW0Tqo0T6AyAFgY+FcuZ
Bxefln+UMCyNvQIMv8l4b+hdhozB3vKyZ/gMly8fvf0GYgelu5x/r4cbSyjgBP7n
D/BWYjWszl/ItEDZ0W8uib4OZUX+9r+gosmOfpc0w72uzcOVGk38HIwQNHGsFqss
yEGHsCGAuj/GiH61YtxshYO7d8i2Rp2ngeTiqh+k2gg+RMntnyzyaHIVbpudztY2
sBAk9BF5TSqqdmHxu7a1ha1vkyr+sp/olp3o47R3IUwYx+RAG0+MuRxDgVt//0dM
ee53MQJ3EsaPKbr+FDw9HFubYQOdjGPSXMxBmWrB6ywqXfL4UkIzI2sJg8AfOT7t
8CNi9zz0Gy/7BuYOxJOT73m2SQi6WTH2xka7fWa+OwWnEy1E/Cr8PAps/C2mpd0k
dsrg4GyzDOy/d5IIv+Q4a4xf8jsSre2hYFavl7tP7aIWf9236EIg/V8JgDcVbJj2
3ED97whMSgK/djj6fW2WZR3f7raHiUX3dpGMV+SkcfdRUCatMeD6DRlGegqUjyS9
MlizHVDLkX86++kNF4MM1pk9yBJ+S6VIeDK79bmD7I9WPhZmU96itLiuNQ8Nx+Py
8CKsakyH+gEtc1WhljLYtHsY3vAE+Hy6QFl530zSGl3anlvM3wKYerkdzkizF+97
SLXOTBzTMeeN+zLoVd5KYDCJsYK9D2bzFLr0k6SmxFQ4heMP63SaZncCF72lZS+z
arjx9sI97ITrwEsE7tXlQdLg42XLgLY1TgDUeXwXiyV6hbMTeH45GIbIZQJFsC4j
1CTz6s4ECcSviYmVPFueT6/tmp0HosMxOZrRnMPMKLRECMs3R8qsoJVa3w329kl5
I9UxYqEoNMSqKDBt6ADkmxZ8ZAPshT7ruYraEQs/WVa6KQwSrKoXEg7YwwShL8dE
zmnUP/b+yBeJnrP9GlktgL/ibPunjybEsW2S7H03q9K8IFBW3UoryGxxHMsDq0gf
dCK/UHB+FhjBgAKbXGBthAY26Is5O1d+B/CK24SlcFaysKQqkT3fKpXb3+FVwJ7U
DWtFyekrjdPiuKZ7Foe0UiBcdRAgqvPGdmkIqHABBETjo3r3GuDVuWXmueKl8XD0
MTFfiliNWy5oQMFXfBkeiUqqw1nIoHr3NvHwSSRbAsxW4cwJyGdkXQjsPRCK6AMk
0KSxNVWb4MhsxjYB/ewJGMl+hHTH0AguJKEHATer5FFNF/VtNNMzNNMOmCnSncDy
fun9TM+LLeWV9qM1zFIpYuzgDHsiamo4kPwXbgyU9oQWErUCtsXY7FP3vv0rDW2L
pLoeLkLD6pEOkJPHMSimTi1y4PVmNjTFIYQ4r8sJTl+tKqbbgwApyR0g+QUi0Mjr
SNlXMzVz5svd4/3rIbuiC17gLVqdurOhDWy9cwGB3azevtqmA8YujDhPxmuvywGY
XVLAAHJkXQK2QNQAuWTpxdDDif6HVAdEZBXQVtNtmDtUOlpxn7xvj+hrbYxvGz2O
tMWeq9V3jnTqTceEnvpdmFqqgZ+reb/d7RODxcm3p2jjUHkWI0tyzwUna4lvgNkf
T18ilnnIUOiXfjbp/8Moob7JomM2ECMi4c6HHeWX+Ac4CyN8KOiYTpEGUmteOzL6
59RrtqGrEAVVLUVqew9hR/94d4IdeD/PFm1OBmn+ruDyeIGdb9Bqo8yCQMFsbbwd
NyDJDyxJmeAb4sn77aEJKJN2PxMy4KiT8Y4yNpb3g6NRnQxYL9AyCLOXRJTF0Vvu
kJYHCld/rAYPij1FBpnl9lD1OBeaL0JQaaMfu+qJNvjFYzPx8HprERdWCZnwXUfU
l7MC3SODbK4uelxo/sn2g7bdbFZjj6Twvard01HeF87zitoeWpIgL94nAQlbM4PJ
WMnig0hBGB6OwIxWKs+5vt+3Az+Ywna6APxwP5hWF8U8DZkWV/G2z5SQr3mewXP3
pIfstPHvE5bakXuXQYIzS6h+LTi9UPxl0dp7616/3n5n6sY1lTbC1dbQm0aeNwGk
nGjTnB3o0rudMuG7yA0BKWRy65tEzk7IOR7BV5WGmSivSNYXX2UDjZSvIbrY8Atl
Jw5XSV9in5R5g3+GZKYvbwyRjW3UHdhjmO5C25ssq2AOrZ9iF6M05k/MUP1eCzZi
FOlmqX8CoViCLXuzGh/88lDrQddSh79UFEyfmx0wvZTfWNxc22sbaqZKUi7iRgeV
VKizwORWCGxbfDr3Mnm4YkA9Z/i8WYjPB6S0fGaNRVhXtDG0cGMvNhFekYBDwnk3
j/usWMjVEY/AbxX9aISRYfJEOE1DyC1uV+LlZmWtYPn0YarjecfbJ4gZURlrxTa5
711++o8gE0fnwNfWAGj5eZmZyAkosbL43oyqaiyc6LTgigdEC9f3ZBi9wHHWO4RO
MwqwcPhZWj7ea9yIxsVvtuDg4YMbAOPLDSrv9/529JN0gGih2IELH+5+tqatrlgz
fQ9ExSeqKEj692nQYtGGFoZpj0ot3Bal9SGxUA15pMFmVM6mvpJU7isn7vK+r4Gk
663pzBEi1ZXRSp2RNU8qUUVVxB54t9Krs7fnpjrzL7TzfCuDyiiwxk8ZHZyVSFLF
cO7YxjR90M7/xrsG0gI5oShpMEMqFZ12gsgUU0NuWmRuSUt7irK/fE7OktM1Qxns
1h+Vfx7K+Fd2l2wyLwEX/inaln1MfYR+MFQbtb8mSeQyBKgww/1ZTOHsxjrCS5QA
Hvtc2hyPQoVhqgLo8+HnQfLNPCXb4NushCYfDe/1YeHxAPvE5UnXuJkKmnS0+QuD
7d0MEmLjPJXNrEYtFSHUql+sNu0vri1VaPSmAA5Y/CyFCygDdlE93c9KnKgTwS9Q
CFLuc3jO0mWOmK1+k6/S97R0WhihKNX58dUTV8HtfIpmEYPTeSPqtD/Q5TkMvcRC
6FbShEpJb4D0yoT1uzyr2z8+adxg+3+rie8CEj50nzWnZcK+dtM/4+90GqjOys+v
jU+Zd1O3/ETC74KdmMvnCPeSSFFm1qrMosezyxG7X8ieftGQHzVawtppkHdCN3UT
PttldqDcoBHhm+0+Cg3qE5z+nPioyjVSIYiyzkswfVI308Op7WyR5gTTC1DGKXFs
Olmi3KLmXh0/NDdRpWyF5jfWtrAfZKQhgiKsFVtjUFtA+yQOv/pp9oTMBz4fv5ww
EmSBbpsSZ6lKwoBF9NmZNwBl6rwnybGcpFx7oKT4xCN9hRbR+bH2BzxL2UiiNn7/
zrSlPEQyg5SOzGtXMY2euOPvmz58A1Sew7SwnGMn4gquCY76sNPZouhyjPMRh5ks
BoXHStsWKj/WHsNNPGKdNxkvOO7nFVRes+MctgWizRuWxMBOPrpKjPuBnylYDhWQ
nw+3VfUIDCo6XT/2unUVjpdqycqk+IWFEwloOjYgjkRUvCbkg4BrFpyQ+kY0jP3h
LzaSFLIb3QqW0pzIwcMovv1vhnsGDGO4aiyDYF32KMfbhndbQDgl6IC8Go3gDAcw
gEKS6Tt6ga/wNhx4jCJBIR5RX4IRhCDxJOP3HdrT7ox8lyjj/NEtldNdhaBuDnZx
akKRyJcacvZJZaQWoYVAtOGNusOvzYIjhIzVNM8SgH5HrGvGuzCV4cu3AK3CmCqw
5RCObKkmnlOcuKMPQ0yPVOchVfm1cuCqoVAseyIK77Yu3IHqSdwwLwKNr0Ao6Lq5
3+LIGU9ecIfjlKBPZI7eKPDCGF5VxCZCtNz3Cw//kB8v6heBF2YCah+3ROK1L02g
JyCEyqYYZIX6n5kHjwFpFirP8Hk+JcJoFpAyJ4UOS9awAwDSb/EiUMurenTXBoCL
njHlpwiWkAIOkWkPsEHfVX6xQo9+reo+gvH1D3y3VLVHfWEpCIcppM8X9Gk7uJIc
204xinHbAE2MIKl/5z/TWnHANtqBbFsR9sNNLaE74EHcoBeyP4lCBpoJDbRsT4X1
KQQVsVRH0vuqtfWm4jmzNEojgue7MsJwQBXXuDAyVB3ffjspLXPnyDGjyI4Pi+DN
tYTYB/W/jgQ+fUMR+EtKwoj/FH1FMBSC5bw+3KKrTaEHWEOy6gobtKYGODmyeMHW
yRfEOzkHDSOWMUmn+Mbm+gLp2rynlhdZ9z1lEcFsCXKYqHyEc5FRsLyfBGBrJibV
kv3MpZ1sHhQILrFjuosWYipasCCFFhw+/Pp3nPF0iSnHH1j5FvseDs4lXcOteSo5
Y337HhL3KIgvyyC9Y86p8hQ4LsIL5F0TwXy3rwxG/PRsedH5Y0s2IuqFFRkzSIQz
mNofcZ6aAbtqnJzJIJOZmWT8IqFDtGxUd2ZBSeAv1gXdqauGPNwqrmbQ7V5UUcJa
p1HalnsR8r2f4zOJFhbcu9PFH0r6LgtYxsXCF3h4BH3LcmQEDJJTF+eQqyxwQ8Je
+MnNEZXfzhpAN7AI3WIYRWAaGZNSU6Bm6orRkakdaXgCWKMkpMm/xSw2U4x8d+ZZ
xQp/zTDtJqV00xaLA3u8PasYmRCHF2YXhELA7xY/CYtuzmrtWsbXKatjyO1N6QYp
Gfo1vbHocbcGYgjnLT1VAz2yF53R9Gj9ZXpWf4Ofthq4iiT/PB7eoiV3K86j74D/
yXOmbpV8C/nlIaIWcuZMy+bQkCSSkU0GSI9QTXCMO9u06Od9baI9RMOup3xJ5vRg
O60Wx80T5K5S93haWi9pdf5vfNk4rFVgJiUJGdNA/qTSxjMveSa3aH9xL24YNkpy
N+Wiuiabut32jKaaPEmdXaMCzdfqbE2NoCQkvEeoOdkeYr//g+VajsZ0SJe7K/UD
yBK/tWjWCDREwZJNmAKJlrca9tfQFOQeUwqQqlS9MnsDwwq89C00ZkiywFfkrTlN
YG7lP1b/qtiHbHEAy0u/6syI161sPvbb5M9TC7lafU3TLj6Wi2OBanV9XZnyVLzC
KtqRf1qUTE4Hy96zYjV8qyFeKYecFgq+5GwqL/dn1it2JPbFzwzzpbPlehNZq7yY
mWNZGGM2OSS8E+6INf1B++Wby/jqgooVD0OppGIHlVR85SvtHcjZWFtbKRgSngVv
zLS0dn67t8HiZZGH0dW2sogqUozBSAouaydAprTQJhTI+BT/gEODcZoEUEbjbgTz
fxKSHHFnEEwGlREch0CFfqh/YqlZJUyhwPfJoGiAuqXWZ9ztPVoNdOVWx+ZEgrjg
dA1mEeIVl7AOPSTUoOO4GCmoFv644ykj4fKfRDl6Wdm1onBrrUdAlOc3fKVzGfv5
bcf8e0GqxvXB73YqpGwS+HDk/NtQgFoN83moQoLHU7XGfpVgenb3gEcCYYW9sybc
F1icVQ7yD2oU9IW1cWGAxdgkKIyVr54WaZeapT0ZbE80o+56y9cWj6WbKguG1McM
9bTuoWQpNZQve41SLqDobun24FHeAFSEEgTHvrO/yyM373OrNxo56jFysJFoO25v
CLOLmwmJCGyvwzCCoT2oaKu6qXeq+owA1ypSDMpK4pCy9uxZHJU+bzRpy1Kz4AB7
+ZCp6jlDE/2EPHTBhDFnmGzH8uOIdIDw9eDd4/qiJmZwEXClvPVU/oBk6RAD4zOj
TmX7NemvSvNwBUKgdAKJg0RbDkdV37tj3UVSH2rBBNk5osrVwdXglGXpXxhfRcsa
8DjEBneqHtxuGiksiUOK7oacDWI0v64xKDHIfZLCA7tsnEPG73VSnjBXHGf+3dVy
T0wkslpz+Knx4hrWy0driyI2tco/sySRXjqgfXMM3Qz3F46A3V1IljSm7nxCZ9m6
DyNiPUdtX4tMN9AKi/f5rQc80y7x4xVdSgjfEqVK9Lt7HEXKOhCtbD9MjIlseBLT
p7M0wlCr33+yhvTvvQOJtsMh6J4SDd665X4P6yzEaPVNpz7vF5V/tVQY+8HyNhBC
XsntK+hUgkEWL9rMljcc/k3Pp17DUOmgr13cRbOrMW7UIXUxJGrvnNrEBY5GK1Ks
jXuA/0D47aRpMYGjf8tLjL8VXb3qXu9aPQuCwxDTGAx6mmQu2Kl+g8d7zvYvNOaW
ehCGHWcC6ia2gfLYF59n3Bk2sDLX7W0P9efIs3D67mauhlAMeGntbCeqNZKLxCsx
xtEgo3V5HFDmPKcwG1hm8Bb6SVOGYcYkKgDe7vugN45caBakbV/vLloHQr31xJEl
2go4K7GhuMiIAa8Qa+cl2OITj4ojUQg+CVj/RrtmXDrlR2DqWsR2ssputipu1fdp
23Ier8u9H6l7oWI285qAWWi8++jrTzA2m53zxqwVKJM1ItYh7igHVi/rig4hv+rR
5O9m8WVkP8J9mn8zlUWhIPLk17Bs8vPsPMNwZA6hQfJzVAUFkjnXE4Enp3I1+IyC
eB1zAINdyHD2/G3jPji3t7wL6gKn9eNJxhfYcjkhXFnMZgJjnSJxucve+G7ccEpZ
yONLKFwgBghtRTqqkBUGj30rTipo6nD17hn31fC6iQFh0RNxUAFg/PpeJoDodL6M
WxeZklFqqyxF0tdLSS9nPQXbYwOBX4X+/uXgmKsUa2c/cFCgbMQguDmvEZy+BnEP
dOX8eiuJ8mPPHXqT/Bxmv/FzZOPAOq7Ms9ltsp2Ui0MOeJGWcHzukARekjId1lrZ
RPS3MmOCH85DE2Q3lKoVVkkwAGTmAAz97MvRzdTjot20vYbLXscp6l2EDFU+OMCP
CLlsvXcdFb7DHbB6ze+6Uf6F98cuUO4SyVjME+R7I1gwzy8JSCpVZ6PuGSRljPAb
gFgEhKe08hEwa63B2dT91qgyO3xxRfLfYYQ0rPyn2r4PvgSpKYnPi1QxIfZqIbfm
2EyHqwYgq2UsCm39cnISJNii6btXPzN+VTkOoKqk9rRcX9y1SJj0sGXwnuIt7rIP
h+bg1eBoSOS3C+7qGtnvnkCul7qaIg8dfbr9RQm5BGtmkxIJUHrEEXF+ociSyDhD
3jo857S3Mb1Pm20ua0/ZKwqAd6Kca0sbYW+TP16G0SRsv7QcrqwihAqOYusqH0m+
e9toopBa5NMGomK4mLX2tfcuIAdYgUtNywanbCy3YS/sJ4SsAy0bjRKFlj327ICD
px8Y/8321HaHPGG47tlQ1TjIrxBLulLImq+fYqTaxgJY2o7YhB+naXFqTYZ3DmY8
yDKOwLgcx1w4PUCC/GO08OIcWwmSq2l50iPiaSXcMd3zt5+TMOZXT28hR1FE+hmT
cePy+lzpTAH9ZNDBtr4p3eg3cFlKwCtlFdbgpBmW0V2cgRcAt4FBikyi7ZNlj9ar
vyKegrBtLPWjduszHYr53KisDQ50w9350ajYw4mtBGMSGGmOiLcHl5hXijJLV5Pa
VzEsRRx78QZ9JXTqeHF8VCaUh96ccVI7189Y7LlUqAPdL2qRsgEXdZSn847aIAU/
xu0XqYhUyO8uBc8n2GlSh4ncVijuH+IHITJ70c3tEuz9lHSE4d+FuiepT7S2Sqkf
PBwYWctrO0FsGrK3CyJ3vzNKLDgK7B0klUQZyDit/Ailo2ikQ/j/45AC2QpFUN3B
7VOM94wVVqO83Wdp9iW4WJYiyh0WYJReUJNfwB1qpyRBEUoJBMMensjWGx8oxJV1
j22MUYwbpNz/Eyq9dvTA4nvqkNJIgQraL84Wpyo10KbCZxrrLiVCfAUeI/0eLcRm
1KahQ1ReVzVlQJFMVOyuX0GnN/k7y0CMGeljnxQaIkDH6mtzu25ZENYkXEHEZC7Y
9/r+9M41uRvV4xO7IUc3uD6h9yLXWZRK5N81h1vR9eGqrXMktrVVnDyF723fgOrz
evkBP08heSpr+Y81bLDTGMANbnX2QV631cZMPXm8qcag48xOch7DSo+bT4R9vav/
8hJn1Fkb0zmrUfjZ2esQA2laDgahhdlm7h+x/jtHZNXc89nicDvOr6ntxtsk00Ns
d+jpN3j3exO7bH3uaDgaFmHCscJluvHOyCdnjmYCH0walHFYBRVCJGnwWpsaAW4R
1gTBdiIH4o/mEbmUoG0ECKmn68m4WvXlc4Ab5xCHMkGsjMSDYaM7dDilTnws0agO
S+LKaVPeS7DCCQqO7KhsBk/7yAMWKmg40WC7GwiC1hy33UoKLfnEKa9nZibvbCqn
m3t1TwCodxJGN90FaVIS4LZWVpassmQews9Nzctpr5c8TK4yC9Nsc0RVQMeU9IAC
vfDuNIDB2IZfjW+2iLJAT7b1kTqaIeprK/4YGU+ElZ8M73DkxG/mXiw5unqGmLBI
XNvVZg0SvpU+IHz/ovPtbxBujUYIlJEBg4XCnQ68/k7KPQGuoh/Z1SMkh//5pA56
i7GeZMZn2vl9W5gHpJzytmBNXOQL1Znt/ojmyayIjVM+L36P8KNu0unoc5Z83D06
K3gtXpRf6aB8XEwFHxLRIJyug0u/swyaMtJnqAgwvyPj8CMRir9d/M/8HLk+M8yA
Kf7laqUg5pGZMDiLdY0AvV2bXx30KrNgVk/qsOiFgMWg7XdR2xtnwGNjwcbarZEL
0H58D8AF/isANOPer8ezDwJRa/FGVkxIB07N+Mmr1jsKVioWGOD5+mMOeAUZ4ZvH
fJlokvt7zrg4gKFqD292lEojAKtpatCi+S9IInYP1vehs3aRfi1PSZYL2w5HkLtc
bGGtyZLoOJfk7mr5BVR6wFVp01IX6UGeZRxLHgK8Tc9Oq5PBZKueknztbuZGKTOD
zACGupKRBTIeFKE8zLgWDssV9/1XV5Viyt18qu/za2cbOYvdfuoobpdIxqx/CEmU
lAIfSPa/hzKBEkIFVbkgTMiBRghi1r9xCVf/H2juXPKueand7bgD3B95PAVUyhGz
nSH54TZygi/+P8ea5/hXER0XyAoeSxt/j7ibPdcdfZdM8pgJ537wRSEKUNBghCxm
h4WvckIJbi8t4gwXCGCVQgi6zprDUtReaG6lFgF9HMhIbAsJiEdvFk4P210j2fT6
eKrdgwf1KGsO1SYMcwwenVw8njhae+o7oAmmoF4Ib2WUjliiG/UQ17TM0zlJi3au
voXiVU9DtBiusTJJH71K4UcZevm1kBLbNT7wT3UlIgDKIzauBJvRdhYTQIqMNwLB
9lEJ77ohz0UUSvy6VbONspNlc1jt9JAxRkIJetF551lvxdN4fz/RsWmTfJFMBVc3
qzvU7zRyGrIOUNGDBRh7a6ikrqdGOh0NiH04zYunpcWRaHaYbMn7eDDQwRP1i89X
KnxGa5gPM86Slpkl+Ee9wecRV0ZDunhdvwKse5bIMoDYLbxy5SNAwq3RyKg94WNX
iqPUQGJZ5QsH1sTLWJSCiybC8C+57nrjsmIpR4dUqv/FOKzdWT9HIvDBrx/+7Bsz
qlnUBitzfj96H34i0r7y4BGJWfaZavzJNGCJWwULL1c2U0fLijNjI4vaMjrK7oI2
kE3qKDR/rjhcPBmCo6KyMsurtXQIikxL8hQbfXj7doUmdHvnAgB/x9Qf/4CGvAC/
z+uEJxXoecwnmawIA90slNg448cStsIdsbk9AANcHIans/75YYCoVjeYs71NQthZ
LfZGLVs6d7XsA6qimRY4nohG7q7DlQeSinmWILvSLT38VeVA7CtWSx0PXHAnRA+R
ZeKuO2tAKZ08wLneIy4uUMpA8nMJ95i3N0TEfIbY0NbiImvufRQ0XKFBooGMyBJg
aJOiQtkF6B+wevZTbjvTyLwZXzRo88UPPWEKuUVEhYja0LlHglBxBZve0gBIFe+Q
MKLKhqi0uM3KhzaX58EPvJJW//5o/sBgJYI/4bL5IXMOffxVyIeznY6a+MNj93RR
rpd3mDWL9sBxeXEdAWjIj1fpRLw4X4QcxAK5AO+UI1gEISOO75mFFzL5AO3RVRd7
6wssKauBq9tmpTXLrFAAT4w0BVrYLOHLyilZ5EAOulXdj+qwPa63p4WVoo/x17ng
CWYGxdlGwgJ12iOlaGwPsGexvK6thK5+iUPYUe2w6QjIqG+VbBsYsI3sUPi4s3dh
kjyhQLNmQU5tu+U1kS8nUGvukXptP+gz7P48Sk5L1haE06GkckCrYAO2xHus+sus
0Ao8dCMm3dkxAOUeX3if4MLENl6lJGM3hBa/JjAWxNZqI27ealZhb4pQ2SvOrRxd
oMLfbYNg2XDlE+P7jNDzn0nAsOENGP6psC4JPUbjzDgYB1AAgmWHncchHz7aEnvO
1dQkL/ZI5oYAa6Jvxsl4uI+BVn+Ofg9AyOM1GRK7lKLNZy/j7GiPXlrkawSP6kL8
LwXSEZuBX/VLpgeoBH/ce1FefR6JO99kY6Gbym7BBP3dTK+vI5JGv2uSinWCp74S
zZh+TejhvFw9L03KNfs5eWtP1I7miB5eXUHFvQ0XDw3sEIiaGUfVvqPbMbHqoCKw
wvfDDWVet/DLfkIjp/HwvkZu+WEXkL6lqywR+eDfvjEdavcPuhuN6DoFgfTMQqJo
yir6gojWCBuiBKMKnBVL1XMPqE7Fuj3cpbzsyQV6j3ezTeTiwT4tN9Bj+vfGllGR
e043ibuiuz9D8zBHHGTgsevRxSPIMHD8ZWkIld74C1f6adO1m0KOjSmoIbofv8v3
mM7yLniCcWJwx8brF/Bd4HmH6aqKKN/Caka+AvxUdrZlF3Y7ELGxZmoimvrifnFt
LGXVQPFMc+lSTEa/mZloI92B9Pek3C7ZAgbznQVFiXwt5Px/BtzmZLz9RXTSNYbI
ObPF+VaWD0Lgbv5fLw273b9RbrHHXl1kfmuWiLiyd6GbXuoFehZ1Fkq1CK4OBaB5
lXgAwag3ywSQcTz41pSVTLFugtJz0ENGh8pSWSoWVXoN1u5VGtWmWd+vubmKYGdH
J199uNYRtVtpxytcMG7+P4vAoviBHWVPfdiGafFe10b+VQbr7khWAH1OeJiGzSYZ
g3WmhRlT4h3rHdrLr8vIPZPn2FMnFLYvJWRZK7+i+58qAlmCzG52x7R3lMQWkIO9
V8wq46BD8XPBSD56bn1kHcoZnvJhcLkDMi3aSOerncK2rGmRj7/rtdHnJcqGWeEK
ZUh6fwf1og+7LuEFXFd1xCkuBBKI1wxMkHyfjZ58vNLUvqXvQq8f+IW72v8+2MIT
He9N7bJJAKLBmM8lYmcLCHG3GBXXaUa/GZQPD7oYpBlepyu4iRaSajZB/WNrmapV
j2omwob+KvVyX08BYt7Th5ziqZelKVHs0cyim+ragpeLAj23s3BUDC7Fr88m7StG
z7f7uGXEAteG4yfUeK+Kgj++6Qm4CQoGfNvVcMhcXQInVg9B6dCWqgDhrAM6oomI
znNj1Jz422O8Y6OrNDVE6ZGHlHMM3y2QZ8RgZuGtYJX+X71/GUCE6JG8r0ImAtXd
0b6RKOMHcyUl07F+F/Lrtf5MMksjhLqeAXPbt7QShDj6W+YtR+kAUurVzyrp/Okq
PqeZ/VG/NZhkGPx3i7yZz3NEf/glWOSOfvamp3BPOAgEtfAnUeTrsbTnnq3PUlff
xPyABfe44ZOLf2cuEuVmOafZSB3cV2peDfEWBFEdikiAPhZW7U97aiNhOqRxGhF2
nnYTbgcS5QyJPc+YzoHYKtyEbKVeD3oGw7TKLTc5/SBGReW32nG99meB3zXk17KR
qMZKiCvb6STj7rEoPUZ26Ju0j8sneTHKIcv3hiEh6p7S+SLIEM031F6gstlMRqnR
6HSAF8Sn+V+nX/C8r4iJRxSI4eCIEphw483rsHmKvsZBW52X0I5/VnN2O7IgICJ3
+KGjcSc+lMoRhJ+cEgGeNfJfz1sGEqWMV4w4AbNiRrThDcB72INGay/LXoTL7L9+
XcBl9LqyxRfx1+sItbher4U2iPe4zGXKfkHbgY6ximotYWhkAH9GzxOCr+LUkpbB
m8a5/UH6pdm+ndkcrVLGMPSt4vcU4tKtzDeBwRZYdQzx3jFZPS4GN+m1gkg0YnnF
nrMZVLE7FkhtaJw6Z4bC7dTw6GYDxtN7DFLQUKQQQH39+axPpHl7jT1q+bV050xr
FiO5RNwiiV640+/b6P/vmdMLWx7FBTvGSXS1bL9xJmQcmGdQFcgwcckGhMltmpem
59295N8Eq3H6QPQ1il5wQ5xgQCN4I+3/CXIp9wmoaOZR854B4VEdvgMLPkYBgGaw
ka68EMzScDWvH1c7rXaext8pKA+PIoaQxeJni+zjppA7faaH1zX8SNdetzLuIdIk
5HW311Q9PxKnohRweEnz2PqNJJq5YRmfn5AFsn0C29aPl1eSp+f1VVkMv8COsm1D
2YGlikLJI3+G4LTsenNB/blxLilH/fCdLylAmJ3/l93fjV6JWaf48SD4Bh9KdC5J
LceFnj9FKkzciYpMdAyahs8hapSuxV04PIymguLMz+VSQJ00AOb7jMu7HB1NMg+j
TTrKiCNh1WTeTzZW+c73fKhtDb6HbNZ2uNQjTvmavZYoPhACyfQsVfAOsP+dSUF2
E9qFblKPgdGisRIi4ZR6fJPVzDD8FsLy+0U5MtSErDYWIRW2ad5oVYMLGZB0Yp+C
Hr18jCTT3fmNi7Z7sEbvHK3mIeNs/tH+5bRoEhzwSadUoPX3FQmihaGWTvpkqf4h
vlp2189cjLL56avc93iS6rM4iPT3ngFNnGqM3CV4tsp6UogxEfMf7vRUDVm10Uqt
/Okgz1DijPnCz2xxch0y1odqWROOD4eEULYi2fTVBL7p4PqJZLCywOqOIBkGcyIj
CsOiMuYjiZOAIsxrV/FJAJtpnhWFJ/cIfay9d6ie641amz9mxkC++u6qas3TY5Hz
AjTuuVjFTbeXN8dpWSKMXFKCSDguNlqsKSHA6LMGmbLNxMWJkWAohiIGoWFZh3/l
UFwQ/cQNuKEW7q0GQXCBlOBQHXQwxAUiwBpUgyscShYWRHUFFA2dLM8FOjTxWZuu
28VPwGqIxIYuKqCt+UfTIM+U6szCpYOaWmCtMXASEHHblogegKL2zJDCCjdHSLww
QsXnzwVR06+rTXEVL0zyQ8Vr6jo/pWL1bkCcojKThAVE4HBpthiGJQ2v9BjjQwoY
hFJ60za/SLm1v9L4nDca57Hr6gyfhrS00uCzNxkZPyhkZkWvYxKcfYzAKx99qkF0
tgj+rjHysBeptAQUS/UeuafPOYv6BJ4MZz1/plKYF3L4gOyW4H4SPVYHgOijMuqr
rWf2ZDJYdVCKvWp7i2HHuCmNUAlmy4hIgg5Zp+YXISM/AsbNkg9/3w1S3r/Mtksu
LHOI75qAYmAQzL8wZT2p/FnSmMff7UilQk3sPc4NBR6rrU2IyoU/9YghffSK7TwD
m0Rd9S13jEB6dNIA5WkEqQ9+am3xXJfa4RgZ9MWLTBGhnGfhI1D676Rwnk/ZKt5q
w0D5nOnCryoCizHeVznA5n5is6r4EuW9rilc+ToJkNWbh1w/B+Sv6Tq789An+Ewr
ghJACchSIIHlz44E/Rjl/ZXJa/JRAcwUIBCki43sLtsgfweb21iz4ca6vaWDFeqI
y7BX+i39D7jDmsmPdGfONC45p+XC2Lyx1lyk5Byr0Ylwc/b3AaVhELkKMuHuUMa5
a+WdYgAE8bSrzo4tl+NMDRABqUKGMw/XZHp61pN2EnoT4kkcYUpSIedvYsiI+9od
KIYezV/g5zKjNQM6eu/8FbsuCHXvIlPA/SRlJIXTBngWp2tI9w7GQ+LdqiiCoLgB
ZtAdY2t/FbAcyF2em7y7m8lz2KKepfivAvDH4Jz5E1crEs0OUrgqWpzfmcLJM+Or
1AY0EKSaCfYuHYiZykOf2vCijyWKyrH6ERuA6ai+MYdnn9z+6G+ercX7cwyBYN0e
3Z99y85w2L/bK6iw2taeEOliWy+Jy39aHC1pu6kqDYV2Jk4fs8Hm6x3ZAMTiLijn
HwbmjrV/WknmVaFl0BOW11Xtcb7IMPrOpB6Y5fQl1lPA0c4BPuNQGbOZ4CfBC39x
ah6OYXxk/7rmgrq6ujXtsg5E1N8OJ5ffpYSIZwhipk9nSjp+Z5tjzbFp/C5EZJpE
QLBi7jrgBmmm68PuCLfo4WVBU8TWaA1ii5l+0qIom5IgBa4kwQdf+vXEneLVvIyK
/yYgbQCNaf/Rr+2SCWjMQzw5wUHWh0+N0SHA0fn/t6l9A4vUp9hJr27xDk5aDTQ3
xv5dRY8iY4IKhEk+zWTmo3y9KuF/F0KG6xnZAaZLBOeTUPV2hUY2N6vJpZa/OrR8
ZydCURGze7U6l6tOEElFmIrkf8zwfIWpB4uCJ0l0OdB9RA7941y6Lw8tlb4Jpwom
aETRJ1LTBX7qr0/oh8E635beGmKGmBnUJcf9oWL3bAPiph4gWdod14kUAm6uYfc0
3fC8hNYJZCWwfEICbaNUC2L7SCDcHndd0R7yl80I6eXmpuXkA/C9hf2Mr1/2HGdk
n2QHXiIko/rADN3gX3mK2BHQNPjI9Kt9V+ATykpph6lokMKtaRuILKDfn+0KzY4V
0+XgG4n5uOuJYhAkB16E7BswJEzgbOY1Xuny4RY2NPFFNlH6GFgdpyKQk5sHGW/s
lcoA57AwV9xDj6vD3P2rExq/ZzVh8jc4QIeEnLl4mEYH87DO56grBdSxurQ8JfQs
RlkWvGSL2ntQZ08zZuREEOG+GCqy9pdjSy8oOXTQ0k+EL6BITtB5GI+tCsVnqEJQ
zeR5zxeMNb7lLkXWhnQ1XNMbQYdUToVs5S8W76nfS5aarJGdVE7pnb6+C2CIStFi
/YzeNI9ewFrO7ucbEIXyevDhkhkEYl1K079Al0XKuCVV5mC55NvK+qAnZND9cmmH
zl42YpRSp2aEf/fCBgraoUA8zy3rhCmryVEegbs4ko59TuYNonJMkuyDCZF19gr4
lMYPfhHlwEO6xvGlNAp3Afo0NvAGPsM1vDpKcBr8Eb/Eh7JytIoVJNZpKeCBmLfr
67H7leQMDbCLRcMUmEAY1ZTj5ZMyfIkezO1wIk0AhCTx6j9a0mKfr6TKsz7l88H7
2FLKwpPKkyadeiifpwQlSLdLxGaPnNzkH4kCPulhYbgNSe9AsHAy4jpCCJ7l0sZv
ACUr5eUQq4c0MJr49rmGMTb0fXAb2gPYwUrL0NFaAbr5hiIj5hFF16Ps4TR/2pX3
dxnMhx6Ynb4S1rNeOjdb/BraBaymZnl4sSEB22ov/MdnzjIJPqM4Cjb2eTIVOsh+
OamSgp+3sdzB+vYf2eGUR5+GyseY4fOS277/kwn6p0RAvMl+V13d2hBWrhrfhzx1
dQa1AocmuR8vXDNC2VV6RvmpeFKqPO1d7IiDTLNHP1OFIKGBQ9SjwJrFG6jG8F+/
0cOV6nVS/ux7aSxeQY8wkcRPFNuNOoV+L7lHXldg+x53gVbEsVj1L5SzGqn2zP+x
r6fI4Bu5rGjowKVC3F6X9yXJtyYOT1RPyu93sX5o6LMKenRzR+seFWANOZShQcGl
ZEh0+2c6DFAl85Q/soWgxJ/eXv8f0APBVDZgMhql0d+w0E5ZciOncyyWNqvLCL0p
EeelaSb41xCixY6U3abT3A2389hvArbrup87T+lDW1HzasWG6mVhMyU//NtFq0wZ
7G4DGL1zLAArzf3zZPhugZCE6HznCJir6LqVZjgvOhUsvGKCdpuFUmeaTB/tfjkA
XZ/8xUIx3jH6zqFgEDmel/U86YiU4XMzT0Sgg91Ir4YZiEukf40mIE7Ch6kpnA6H
LWVFQlojjJHNVAhwRZVPE0l+Aq0NfkaWgA+B9dY1fWvQgWVXygI4Ji0okLi+DcL/
q6qZLkQFPJRpNnu7GqQcio5wTPZaSFS7Was+B78wEJGcF6gzlCbTVqk1rb7eOfjU
ufCxOVPgttZpzDOn0Eu/4g/OFR7VWV3OtIHvqRG1lRY3ZGxSjLoDZ51mXGenxR4M
bht4SfT4jSD9wba40LhP13DR4Xhu3QlQLd+bf6nZQF8W2FiGwktyaiZj9eGqDKz9
fpLefFCGV5l9jQF6KiE7np9Z/QJfhUaMbILxOPgk4yb3HA9QDWx/CetKYGtIxnfd
h6OborAnT4aV7CCPatLUdTpA/ciq4Q/vC3fcaI9eY7UxUVYESvWenczRSSV7Mzjo
5XP3/vTRZaLZjohCX7ewqCJV2by90Wj3wRz5PeMg4WbQ5ckuKI6cw+mYhhgWBlm+
mHJ+swCewy3WPE83Cgj+64hOpTtZooY8GIyixOv0QXfL9MFU3fa2RWklswXDMNui
ZgmDqA20bgTWeu8LRr856PsyqiORZMFvr42OdGrgnq/BibBkjB9Ay6LkzHsCm9Bw
Zj+hndM3elSJZZIiyG6OzAML6Tw+rYNyN/9V+eE3i8itKHRK6NLnXk3Ytpyl1Zke
kdFATuqn6S5vvlc0pKFC4r+asvtZO+5ghv7sb70ik3AJs08mC5NbS0qku96Nid2F
5fNHEPbK1KeESevVM/KnPSNuHBa2qUEUVgjeAgrk4f0GCyRdivjeymERujD5iEWF
kLcH8gVLlqqqa8wfpyYvYOgGjZHIOkQCb2XqK7iDPodRg/e0ODI11iTuzchoN0pI
JbJRipEom08NWuIGkKTT/SyK3t0S34bNFbbqQrchDje4CEoiaYW9W1SoKb8c2bAl
3MEyx8URBfDF0vLnb/ng3FwEtpWjLlLxRoAXjsPkybjlfrZ41Xr2zvoQ4dw+Ntgo
P+dC9+cB22+Rn6A7HCVvh/GTIloF3hZPZNrThlrbUmZNh5VzuYT/U8CDw1GrqvR1
Xe6m9ktxqerJNhp8RE5fD+cWGK5v+6BjHR6B/+KkRv81goe4kLmcl6s8gdp68Mud
Th36HSQhrwYn26cvhVDrQ8y2EHiHIu2727jocW+yXdZ2G21TSTvgBq52XlvsKTDV
grlcVWwH+ENhXahjCR8mY+m9lsu/k8njrIxBhOhGRd14Z3fmJleI11udZe8m1l5t
+7ukmE7coMX22a63aJGOgoE1B2eBIs2why64znE9ijw7qz7QsXlquw7pFAgB7WjG
4oWMxzmibYz1bWpuNgRow8wNIuQCjM16wQyu/nIgHwPapdcYIS8qSjW43LplnJ0d
FlZSypmdYtn5k7+e1gEvPztMb8TeqH9r/ycf/Rbk+KyJypI2+wifd4x71P27ASKE
eAVIW8KgIWY4AcGSB6U05R5AtiP5dQpabDvVhyMGV3uNXgqzqa2K8oDNHzQp7XAC
8knOFfd9Lc+SdX+5CDuO02YP+Hu4w9Oh5G26tbN5IwuZHvABAc6vlsqrUKuaJaY2
nk6nODb843KniI+QN/qO4es0ZVStlkCjNjyFAGl0A8YxpOEb4fLYcx8Hjd/6RgKN
tmDqGvWxbsECUrC5bzJViLkT2bAe5BPYZjDgrjHgFAj2+Om3IIVUd7eQytUEak3W
7IDWyJGJpuE/hObE48LhixI0lPSZWsELN3pwTK4c0quBHguuvMFbuFBdWV9bljtQ
0i1CCWL9RlB1vW85MKWHffrt14BAAV6MS5+746XKm93qNNWD1q5kbe0HwlUOXH2C
92K4gOhipZEWmozJGnqT8I7sPj17RxmVrav83mvi3NuUHTdJsouXVt8H8G9doI9P
5jqQyOpTZs61fHpr1tc+rhDqmYjpZVRK1cdxvI+8IxmpiXqwiuY9sV/SSIlY1RXe
RzufCpxPK4F9TZWeVUdl9Jp89/UnF+ODQo6vtekhMO9qzOD82LN/Nv/9vg0EY62g
5YOzxfB6ZPEa+6EbXXf1WefFWnn5DTRxw8bYy9SFcw2xRsqhyVGgN8kERO1faAmY
AsiDdqbQwOyH4aZyqFuClyl1UqPU2sXanTVjBlbW57g0d+z2UV+UjT/tGmb/WFte
7y9JXsY6lb+EnvR7B+0wWUBYxWHq2lOrcBv0laPetqlgWv2A1HxToy0ffYDwKXaW
gwAOTSL+nBOMxhTk1Tl3zHcT5oUndsnjI7AT+7gHOnZBLgHeOEg76+hQfG2q0R2W
mi7+XE4SD+kYUk0mADkoTAMln6yKg3joRZS7ckiBBZTEzteo4DvVuYb7Lbsvae/R
2ceiMBCTDj2c+8Qy72sHujAri1EW398U1fygKaypRzLAwnGMPUitI87IAEibZJdi
wScl5z+XWy6GX66/XK0uVGhkrrSXZ6lQ23VwB6O2FqU7azn1DOa1Qnd9eVUTx5GP
MHIM3qHqC8IzpxMAI8TnmOU8QhISf8J5g7mkXgopmnnjlNTdELqLGSGpAXrcl6iE
WlpMLRRH+orGx4TfaTLCZ+SMC08Pvm+T49OmHBQNwPxH7XRFIJ9NVUllRt1JZnxx
zHq6S/FtkWxwNYWxvj7RHHKlRNUaZekkuLl1axZaIbYX+70nzO1MKN8/tA5u8fnw
yXX9grqgSS2cSM0fi6+0DdpXX7Pl7iYMMyfeZ4f1zAl5KFPBSciwKSGNW9pfRkYc
GR3vl4OG5mMPRZNPxGSMWPMbIzP7TyEDfB4R66xpVrKXA4XHPM9qWoW8KEGkEFfB
ZlfKFo7nPA+3TRPFVnZLKGDu9rfZzQBLC9tNdH8u6jdiorGinBOS7GRSBMRV+aGL
xs32VPJzradS+AIhyle2cjmwUmwJUyqKutod25/1/amoKb/d54cuTY/vACEC57M3
HiqsRikevEn0+6AqhDRysIABaXifITxrO3QVZ9cXqptBzoGbUJHj7Hs1UCz5okoh
SXrfg4q+jVvvFTX96oQ/oJH+LNQIHpyrZDWM94Q+FUHTh8lxQ3xdfKkOXigo1Tkv
MTku17+GadzppLZcrHO1mEaEKzHvhQu0N/Q2KQprWVBi2vzBAHHNC3AhKMbV1PgS
p7picM8nLfWN4dLOGqLLHxIKVbshgJsdjN/SfHYl17YeUugW6izIJtfKenQK2QTv
NGWZfTE8osykkhE83Z4KD8uJ7ai7qHu9wPQ/oigm7UpfPs+5faoGibK3mF5yb3OR
Fkk4LwJTEZxFh8LG4DGIn4e9BM8H0FxZaZp2ZEikiUGddu/TSEkg78NTCHfXbNu4
rmgfAgsXILTodhhPhzC3Qp6fD6wQQswG/cdniYvOevMJC/wa+2OS3AEHNTjxXucg
Yegzn6EJLY22w3OYxIfGbojLwVZm0Tc9u1PVeAaSZ9niglvcOTNDa6y8rMAwhbvt
WGJGPEplwc2Hk++tSDyeSotSUgZPJPvAjOQW6qXl7U+0FfBgY+rvXgNoJhGsanb1
OlZpIzyG9vW9UEiKWx3INpgdDS0tCu651ETSpAaRppm4Nogh9VlOC2sgyXL5CF0L
Iv93Lr2jWAEm+IEV66z5ODLNtXOrT8NR3xssn3S4Kb9Fn5hp79UbwOzDSqp8x0HR
He8VJkQof2248MpLLC0u+5NEYsjmLJ/cWR0T6jDlr6KVmOLcxj2cm6oO6dq9DcTm
ill5cS3TcNmwl5kPz9qiANpCU1w3IIUBsid/C0ox2m4Qp95EkwN8lR/5NYVRBIpV
SJl+6kRKFHO+h6gI89rcgxvWVTsAXSHKw2GYeWOVqAwqj18Lt5VH9onDkotvzXos
vE3hUOzotAsaXPzZck6qJH051IQodANopZdZL1FYteDa8SUvtwjayYMDEsh33PSy
R3TXpblw7QFE5SPS9tNbMwIVMFeRtZxQA37yN8+NSvauZXzag9RFF/i9noA/ZfwV
k/g+r5VDrsZ6uq31r2D6z+h3NzSUaFfDzOUxfOpqG/dzV2uFk52yNt7PUdf6xj3z
uQ37DZoexM9CZgF2x8ziPt7gKXTrOgvxWTYoMnMhwTCdPdR5XsJ103vEY5+62BOq
SIh+I4xrR1N+ta4m/Y98TqGw5thot2rAdDCbIfrYBsY1OWgujeXUMfywqSFr732I
qwuZ8Vi9z1ggi3dqALx1EHoAAt/8WRwfLYVAiphZ1uRLS17bVz0qGRonyfzJraN1
lwo9wUzbNOy63+Ik7eroeHURX2e6b2bDzGLsgbPng6YAJLlL4/hf4REycJqbLE83
vqGs085MKqigwPvnMTL4CzjrNpv5J7kHQXND9C5PE+4UriRGE2djhOfStSQrhEQt
pddurQLfrMas01AYVAakddxKFUFYMgxZkpCVg3ecw1dOrSN8P8GJYMHFp4yRPUEO
rZKpnn4JTXwL5DNLjw6Bk13tmh/5bTxpdTtykCvouC7Y+YwkhVHLSsmsMZIDNF8w
LgfEnqnt+5URm6yNwiZHjjKt8O2aW8kIbXGR4SZesy/lVILV9ifLjeLlbUvg+rq5
4Y0+GcYRm+bVyKODW5AHdOKJ6sY13W2UVuuu7Epm+XuY4n912yZH3TRad/7pXO3Y
jvC/kcG2x2J6cgzPn5jZDNxDUAt+oWGhE4cIqrpoM3pBVWoP264I8aajSePir+PH
vDrIMcEkG8r79Zr44tdN4MPgEvZkrX4EdGzCzVPuNHdYrMUjvbhCNQWevZrhACBJ
hKTsiq9qbYkb0RB3vxB6eWT37excq+JzFQKWBTdZNbjj0ENfVVNWLGB4rA3caXDt
XaO1SlRLihiJlvNV0h0zaZqMExrvdWTH/mbHAPRxjqhOG5bc8953kYIMfVsNdAzq
yiOLH+isj+EOEj4vZqIGMzAKc0cFSXpeYB4bBSspzkZTu5ktYZa+Dw3dlDCEn/0c
4nvrnop13kAUxWoy/iopfRq2QWInej+1U/wo2CqEpIjGAn71oh/fOyFtNuh4sLzU
hMU1MuKqOIYLxfRmBs/XHWumrgsRWUVTs4k+0sRWFJ2/8fY3R+GA2jqeBCimOtLq
laSnGbycBIgwxbOZ6GXkJxOlVi7gYFZ/22FfC+wRBPTamb63U2aWWd2TKsnGlZZD
MLlg0NSXveaOssRs92c57f0Vtk1KfHr0ewyuHtgvubZcUrECQrWPVGLD31/xW7FX
+5ac1Ntin8aZSRUFQID1Oul2vbz/ihIY2fT8YxBbwqdtifJqRaBxGnvBUkuNgM/s
qCywFky6kQBp32rswt9TNbJWEaX/skQwIh9hcoq45L2/WTJXvAIVZ55n0OgE69HK
wg3WCkuvdalGBIHS8B0CYNk4oZSPb6v0Ijqvmb82ASHxc4ksuztieJyvFofpO6PE
qYJ383DXb5cRH4gNVHz13pDJ+4Pdw7BYciu78BZp7+9WoBpcBvVdvzbglUHcAZy8
pb1Pf1H/+9crPUsvBXPO09z3VRk0gIK69szBJawRpS+XE6bZ6d+WRWVf7ms5I4Pd
BnFznIr/8rxLaiHDZuoe5B3uJGmrozZGhWrUmhnVRTj4Hpir4xJduzLIukGEzFJ2
l7obL1Z9yQQiwIMWaoZtAO6Uao4y9ViI27ZlzGGXDsHvK03tO4zQvGpU/mtWSzDI
BrqEYxtAchXDxLWu8Lh+hGHGr8R6X//ZIWt8HNxuTFYQH57TR7q8zLW34GZU2/PB
S9d/yzbR/vckuxsM6UGjD5GUCotwZ8+jO9FUluodmWElyJa13KcZJcGxf+aehJAB
ke+LgahAIq4fbyyxsNeAwbsx+RoGtuzeU2l1nPsDLVhuT2HMMmeEg+U1huutIqTD
cWl9q50xvzgaX+3WbpA/XKH1YJD/TAexrsZ0whejGyqLxFtSLIvTMW4MIPmxMhTy
lyHAbMaDKMHwteYceQ+coOGutOoSpUjss66j1R0Ua5H0O+nE0QAVjpeHMwE96W74
AZ0wvKyVLySNgc1Cn8Rmw19lFRYoUAEJ6iVvJHL+kYHb2SldTLIrhGw9MFfNpErs
WhLUmisJjNO6iaBysYVTCndLw1LD/gl1anh9uW5eJy0IXw//haZTPQkAu4HyDwZ3
slSUziNxdK67+/xAywflPYVnjMNX0KtbikA5VKh4zZPnrE6SHQFwRm3WUfchTJ1I
OQ3TZcjUDd0ZSVjSS8fdrts63PBSULcMpHBmxonRZhilw9RLaOpBZ74yv9eOZRcF
Lu1reEoS8bejV7Kvd+AZbA0dqyoHg6Vo4am09Is2lUEX/mvQgNnVnQdD30oJ58Sz
0H8UfrEYvhvnqMV/OfJh7e21TMMlPRcNFpAGwfVbNbETl8rMlJGMdSKJ3pJnV0+d
DI1eWKbcFAMRVUHXrHVVuhR8ncEJ8JSQ+u+5cHs8FS5jo8H2k7IE3gBpygoP3hFC
u7kT8kWJaf95wZlvKrFuWu/Ot9ZabQJV4einj2duBl6JKHpgJXCzWd+ZVq/19WC3
3p8v05Ly/PXeDIh1NINFSomIeeGwqpeN3NmRdJGotgjrgKV9rlW1UT2ClN5FNRdh
Ck8ipW5MNZUCtXyqPvoM6wiaRUQTx9gMNjdiuivQSpuncY9qfWLmv7ij7mjBSb+W
Gfs2vc6xKb3fWi2R4IlC742Mab+0LzqqLBEjS7e4tCmvywVZ6sjXSkc82Gr26usu
H4WuMQj69HYIHY+DN7I1bdvYX5pdRRKz17ADjArLUnCLnm1rgv+1O1GQqjUbrzn2
4k4YEchEvVsbS8IlnOYoAzXyQcTuGbarzEzK50wNsAkSmD//cWrbuwW9dVDwkTaY
ChacxrxjBCkaPSXi1DSU+0UazDtsHFIexobUdwDO052kAOtbxwr5qwzxAeMm8ZIU
LCqzaqwmw9wJHKODSe62WkYHm7XwtBTz0FENKO4UyU1SAL0ta1gBjUZcczJ+TAIh
oJxRSjEssfNy7ky1Svt5CIW7NN1kx2SZY2h+N/Rhhk/kwAy6Duw6jVi8bJkh2f/A
2mZQyXa9TNPd3CrFm/QYjU4moj9e/sL1cJBAXAET5Rm+GUilSGW6VxwXnCxa1xTy
q9nePQzC29Ktwyz6xxjOShDD/JMyPc2qtxikNtPSiP5InnDK4EFOrlYLKr0W4TNk
w2yUuOIn7TkR2Ll4acBNy5SgUhSyM52DH4+VsjxO/Vn3tsqOy9fl9Lp3JRbl0D6X
94r3pZn0JbbMM0kAjchiyBSr2IYGlUXBKApHvv8y39tyxRs8cmjI9Q2r97KTxNZ0
YGSDG7DbqFYWkfH4TGiAJ9dW4JNr+oLOGDNuSLg/9TPMdStHWEXuMN05sXHjq36k
H/Nyqw0eHDEJMvsf6w/LiAko4Ef5gfHcR6N01iktyqi6ezQ6DileNYX7jt8ZArot
wErbp+lt9c2uqEZxWCfs1c5/A2U2gtP2AbDIZueFXlB1mIy2gwUATMsbmmQH2f7N
tycX5Jh80TkFJu8/KgGeQcFwTWlDqyFKNimUsqU6EW5Jg0nUJakqtSW0lZ36TaIk
mcEwTWhIc+kq9l6ThVQn4hQlwD5bvm/LPsxnP/CQjsEEOT0GIPIRDJ9XZOv/izHH
9PZ95eCpY2s0ztYTz+0Vu6/Y9odWXxk85EJv8tN3UUSBGL2+hsJAWoZRl+T6eono
6gOOMlycrQf5rxW5tKjUCGAWhB6m1cTvpfRSQpX4FCWJuW9xovHQ7eDJyCBe6bms
k8sWO/X8gmOdxZFd7shHLfu4r7XvO5qi1A6ixVDFB7oIBheLfHTPw3qEx/VaZjZI
mdtI9CmiX8h+vAS1yzYqVq+2QUnBse66zyToMxzUMkcmuOuUwUFtLNiJSXVv+l05
YhFmiYPgH2LRJ5PB4LSHL4is4TVvR+ZGi4fkpLyadeVm/2tHv7DU9hUJCzpTW12l
hNVd/C7aWQ9zyu4k17lLryYiNQXgieMbHBfveQpbkJJ2lyyBi0Zcy5d1zLGA+bX6
O8R+3oXBKv+2x5Ip54f/OXHQ5z4rb1YzRYCwdC07TYPxalSoa5JcITprkDqSm9+2
JFP0VgBpflcMN3jLI7bDpMnpapqJWzxk79gI0+j8ndg8mv1iqd57Drt/srF6jlWT
WCgh83rZ+5ceaMv4OtXGqExAOsNG7z/TaU0xw80tEaXocuhTu0U+Ya2TL37adJtc
EwC7X5uxSPhsxG7J5Up+rc7BghdnxoBVE9dYLf6t3MFLs/fTaEDMsOW3FhhjOsFo
ydjRt1nnDFKRnoWYKhZRFU/GUwfIXJvgko0qOFb3xaQIEujommWdRt/Vn8Mj2Zyl
kXrYG9kmHAdum8IRZlObyYfg8rNj0QhQ0Hb3xh0hyx4faRsstlF3bI2aXZz2ZZFm
QYsk0wKBR5KB5g4S0mVRMBo76M3C8idIePOnpqnz3eA8E2KEaZV0YhrWNUUwmPmF
gMZcekwq4a9mnasQzTIOkHsKWBe5kqfnXEwzWhesn399Fy66acEo2FGDrmw2jddc
DThB42RSJM03AvlMZkUvMWoZ8RWlwxGdRa59RYtpdRwvMiTVQ5WsFsXb+oEjw54O
x8ainUEPfxVoTi3h7Wf+HXJ8TTsxnlhNs2WEfG9s9Sghk3vnz+mQywUPuIdfydwV
yojscbANd87mr6puh/gEipJokCyVzus+q5fMfKAaHX4JSz8PJjtMklGsBL7exAZY
7CagO4wkZfADIScWqowIg7mzYpbQtjeRB7L2uyFf+xoseJUezAUfO/jChpUNIHIs
MYMf76yznQFgLtI3WXOydDrHWGDoMBPnkhbXUGmk8ZT2SFehabC/mCFAYkZc2xJf
i3euEs4r/nrl+mkdIoZLbVcxG35+NnGI/wR12ZP14BrelSJ0SCiJtlejzI0YDlIK
4r7bzH/BYkX9fhaWgY5h+zAmDiDUv2v3claRrP/1f1CQPkHV3HigPx1oLXPpppqY
35WP9XMUap5rK2fsPKPfqCluiPJp5lmB8nDAl01vWjJA/jf3z/A92X1uamIcRyT5
Ae+CnmTawRFCPTcG3DeWJg7ZYO//D2fHQKQpSJrA4B+BlO9CLMs9RWsgm1Cq2IJH
d/KX+R0dM2MRFayQ8jTWOi6Xzfye1hPZ4NgWgI0zTXKJ6fmApkQzUU/zfQnfOxrc
NmVMaXfIvIXTC72SNpqg1EQ1SI/Ledk0Eb5rlMxNkf5Ngs/CPYSUpgDrttCuosT1
9InMFiTYfYSDS5cZTq6EQRyCcqf1AxCzdKsGqnOxhoVRoWoA6C5rktXiN21crIFc
7SYOXqE9zUM7c6l0qWRZyl4hmfwnDi5DNbi6+/VVNQpmw357xPdc9CWhY+VsOp/Y
S/Yg//UMlIj78/n1xfcNG8pwHxdbiOE9fSsbuSSsdi4wtsGl+NkXeDNcVAeJQBrW
rcSe7PsIv2y2K+ki14ZVPSgmADzSPEgB7i57HfmIQoMaRYyq8XA1re4cZJ58lMTa
aBttQ7TEBlXhZ7awZCFpghC5t3F+PCtxVqEkdxTeqdwJ/VShhWlaimadPlFBOrhI
IQsOSINU0r2eC2+IAS+AeJBAwtAk2xXZiMFRGjsje3GCS9/J3ycss0KUWU9TqYW2
hfoIAApLmmmi9GOISZhmcbPjtGg5kPUFzHt/XJMNkA1dSpw8RYPvMJS6qrbaKCnC
coJd0cbR+GOYmpXuFW/paz1TOxPqUvOTJ3UadELVHmXxNWOLf6rg6ldhQaCiD32w
bsbEvVTYnhL6qwJMjRjw6WqE91cDDUgaZL0aAR9VtlO8Dt7bJpfnMhSRbfRBxF8H
5D2MQfGEbxfRLZMVMuAZ06DqHk6GE6xDuhexD++JfDswY0f+/HTaQBKFZwzBWC7W
g1Gke/gA6hhdGKQ4WGG1rHD+NcY5SRSXILhPU2lN12r6q/eEPngatW1yOLSiI+WQ
1CWzVLXnaJoY67CvS5q6Wz8zRH6cpe/0kl246kVdkMccO4oLbigserm+0MkJllFE
QVyv8HJayBdHzX6fx+YUmixKSqQvjucHJpd06LOml8QQzZhVQvBFGbChpc21Rz0t
cC1VEsGAAMI5qq3A1j7bUDA5ybydJ7TkcaVpnNm6p21xr/eCbFlG1068Vatvpteg
cILENscizMPavStLvbQvsxh7xpeg61MSu+mDGcHmowW/6vmjj0X80QQXYjLADnrO
4mmQ6BZkpqw0tLobhyCcT4IFZbaD5obrFeoriQywCvApzhPNGyoZ2G1mhvtR6ZSE
FpKp2uPj3+Qkf6xwspM0/vNN/QAWcBhLLwPD9047zhY/BuLgwwdE+KJYBULHLqcf
5XFtPWkhxcu9feDD4A5Y4cD6Xf2CZtC5r/jLLLjLf1rqnHTDhfnFtDKJmGMNog2X
okYHfefcE1bH3B1q/yWFNwSsvBmfnvjOq4wYo1j5WsRRQqe7kVSDrBKbI4n21+cE
XvWtMQN9TPh5vzJkRlPbmh8lcIUl4mFt2XFbTTkhp06U//fA1PfUfvZaYJFVXqIZ
FUxlMIXak5jaGvhH2FB1ExgPApHndPS5usl3w/t5erB0kENe/azhdg4uxI7UnP11
8Ez1Dfc2laRZeT7d7kMzZsvZMUU6z8UrObfL4l/rSho8EetI7zTfJEuuKAUJmedU
9A21Z94jQmVdVyVyrq+BF9M3+Oe9r1bRke/Zf4BqbNAvRiQ0lKnhll+7/013YlBo
rfe0BereChwz0anA4CtM/dOq7eUOJWcMGPTP+qJM1hXofq5DF2jMEixgJ2a8x39R
KxKPH82Mmus12e86XM/6tWW987a7/vLYYreNRQAeIghYER+pc3SanvGNie321wPm
9ilvikcyP8ReAOLiVvV7flVp6LYJQIx8zOk221tGtpd4Pynl/V1vJoQJHGa16pxG
XqblLeJjs7x/9uDbKxrygYSIXKwPXP4+e5npr8aUobtTXpGoWDcHaTYXGoNddVib
XToRgsvWrx107UszzT/G+041er4vE6Von1jHPoeGDOaL8BC6qZc4eUdKUB/iL4Yr
MzTLVCrxmSCGgZaI2oIagiRIzlyvD2l6rSGUAEQMolCXJMFkMWtoisQk2ZH4sIeG
V+mpwAUqDUC7AP7VH8xWwxcIMENK/tHX43dKh69eRvImc5LaP3hSPBn44W2N7jrE
5uac0WYUxsnCMcTiE6KUhE1v3tqmYj70veZNdzJvKNDXAo7OsEsCIbEw463dykYE
t7Hf5HYJqAT00dtJX2+KkSVSUTI52bOrAyUA7Mi1OmHmHCdx2xaixIAhjlPVR+eA
Vospq6XoDPx32KEsY7PBaJNUjbzIIMdjVx7OFdJNwjQVoERBA6WQfwxlC7w3ktX+
HD9mZ2R7/cQWCo4B9Q+aTa/g9POSDwsSNssOHGhBqXQlDMG9ehUl8fcWHQPtbEHy
vlHw7eCuS1g0MnehwhZAjD9LQ2n6Pq3/hezGcGwALKdHTTfmdKKW4VrcqRHGJ32m
Rb3h8pf20oSKbrDDTWpSrAxsuLr71zaL9lVT3d+5Dh0NbfQLE8q/Zcv3tnKIuLYg
zKbjjsi+SY1SGlvAK4TI8DrGW0QYpnFO8985rxho7NWDqaPur6ZwzexE0aVO7m9N
rfufCRpGjFbywNWavcoUtMoXUDFaSbHWbhy98mvWNBeQpsNjG0+EyDKnSVd12BRf
R+JASr0dxfqa22RiOJw9QuIU32yM2d+O+0hXO6hDWWjVnmbEfgmqxtdkRU1wU3qt
6JdXDuWh8Oat+b7ZMHRMWwkG1oz/i+1FoWwiA32/yMUo8znLT+Tc+S/30YENt/h1
NWEJQORwLKTxGT2kvBZRoz/9yRfH4P46hQejNiGFhwQAuHXBVFSGd6BczwbeLRSt
EzjKhov/3MQVaReyouyavLHaIUdQMyt//vzT47S2uQsbD3Zij4q4oCrfJ3XDW2wk
h0Rqe4KgrB4tHEGw4FLxPNd1u9unNtVn5U9qVnixJnoLhcv1FGK7751nE+IwDSGN
wn0WnE6yU68yYeGKK9YAGbYQqX2C0PqYD+j+9Me9GDe/lh4HJmVh+vD354PAZ+jw
PWSdR1nYRZTYw0aaPMbJJmiRVC4ziEalTCh8mvhHks/IkNeFRF5axRTj24e6hbp2
rN4QaLG7M4QbKxeABlZ7Ap8M+0/3t+gHXdIIySdBes2x0j9jxVdiu+pofoY0KhET
DWUtWXxp3GMvygrrCYetPosdni6XMe+bAvZm0N8CI5ebQkP3RxZDbuieaufuIozS
YKTGBwZPako/O/OIu88l7AMPeVPfwwbCqIpCfcevslWF6uPPzAYX+ZPfD1wlMB1Y
YFbIUrUdA5zZA2zWioevYHyNpoYMik9Jc4AUvmZfow0bEstM4PHtKOrfkomayqAx
KWDZ7Nj1XPNLK3R4yr39dVk1eA6Ot8MZVlPgKhPwKvRTdJeEAAwSO4WzQzsMdtl5
eHrbE/E+5mqW9G6OjpJv/F4k/5IkQ1n8+miGVtWasU1cfjk9C97iRqIlIZ93dZ4g
Lan5GtQy/+4YFoXM59myP5PRPov1cqbrTrFT668kqowHlpgJxieocKKnB8vdfafu
dAb5AyFPFQCycxKUn+cvI2NNpxGlhk/P2rFzrDECAPIYr4Nm2HOILHs6plG+Ksyc
vvOYilMwmEtLJIsgqBqokm0ZdVqoTQi9D3wAomjEO3CAqhXW4jfbTe+VKWYr0GoG
t4E7L8CRCD4EBIUtxGcY/RinriVaPNDuqWGwd7+90JQxme/RKwtDF1VQQSdwHwtR
TRMGV5pcXraz1s9shgzwh7uBcrMzZGbMd1nVsWVA5dgDvaxywOLkm5W9OlImmBK0
F3gEYuN3hHEu07L1L39yZat7W2QGPQBJ4vrfD0nKwrU3NwU33pCkttLDbdI5y3f4
DDo3reZkbfgpJwjElRQ5sXQsqf9O3i5Tx0egBW05F6C6MyN+1l1e1dZ8YYeWcm91
p4JHdxMeRrPsaMla1DXM7pitfMSP2owf/AH4MgNoniOx4hwKxBA9usZS9TO2ouhk
kH7WcTByqQhOoUPelZkWWXV3rcR8X7yMyiRlz4Lc2UWMswmwStT6PRjlT+KT0wVf
fWKW2stNMensNSCm/FRO56KBBARgifgicgn19hOiTm6n0P2qvYAd0dBqFlFEY+fa
12PagCpVw4MHOKH1cSeRYCIQxPoerQCPGW9Bv4hY0dvhGvLFWsD1YriBffmdtSbX
w1Pkt23/y6nvbwoE7BzhIs9ByDAH5roFV26YmrIYxlUrxdErQpNe94OrJ+SxoeDX
hkPJMv5NAS3xSzUIjw6M67jzwzxt0NjGbmnL8CuC5fTHl5Qdg39K0Zv6PtOnXzT7
I6kXPsrqo/d6Z48PXtu5SaqfIX+/hCqGAJlkIDM7g+iA9ty66Pe6oC/k1YMgRaHo
Cv65S4rxBdhjzesy1Exeiz8rCbgLpa6uaSFpvDT6WHFsyBp5N/74LKruQZJLHaeA
0iYpW5mtNxmWl0HAepwkdidD2ckifkJe+qANOlfzAm9LIEPdu0mC4rlUefF7v/QP
2MjjIwAgUHOCWqGkxe0UBSB+pw2+3tKlnhDfNVarBu9zMpFXBfRPFuaX+z6CtXQV
It06ccrzf0fTFbfsjlqfD0ZPqPR4lUu0HX444E0cbkP54jRc7XPY9TNjpPPV29ok
CB6zJt8uL7EUKdntxp+ckfyhhYgmi4ebO3BooC8d24rj0BJtA3oW/8536+AUUpAb
qeb+hP6mqV1iOosvMjRNYldFvLaW44lCVCdHpfxU6Njhxb0LVF4IB/41sc05Wy9q
wCZPcpURsSuf1SsM4gGpe1VJ+r5K6oLJcvs2XJnP23s74CSl1RimDYVYhA7JL/qb
5LR9DVPutN7ZwRodgs9bi14WwJDDG5KpJyqfRCD0A81zMfvYppy1SNL1HuxXEtIr
42tlHfO1GIWklA1ifE0rv439PWnvd/t3dVyNh2rtuav+hyUKG+/+t/68+QYa6CSc
dAx1UoF2e7Uuo3uQNN4T0sGEEGVJ3ylWwu2rxexNrlk26v3b7C2Frv+kgEo2t1SZ
4i4TLA3moRasqNd6LF3DfWAfwUiM6mn+d9PqcI/ycuVq5WG7Vlw400fvw019U+VW
g5Xy/cgiwdirzvtP7wloflfVybjuDIU2YIWcIsjLQb8Mr/6I/Upxe3X104jRz9hs
avp1pTyfUmvyTM2AWH9Q3KPvlHnTicmnp0z+nFVXcJz8br/fVCWAfljUnivI8Jrx
QkGzegrb2yxuSjBeugunwlL240iy/JyaLZfYgwb4Wpw6cZBROoy5xQ9Z0OgTPGug
95t9dc9VWP/vjqH2yRogbXlPb5cLISUx5aYgnI7tMPntJtMp0MZWCEdQjEv4YTcn
2CrCvlxgqMm99cPQYFTQf/1JrEYtHqxZqyVnpbeobmy7GcuFLwvaanLf0RKy2xbd
eZWFxmRGSym07d7pj+Tz9yMDDsP0dte/+wGaf3Z+kyrt4SNUYBLDO5LyF3GnChvM
CIi1oQun09979vFdKVHCT41HnvT+Z8nFaZJ0wpnbR0w/ZKIztu8DFvw+m8m/m4FU
Gwxh/Kl4nDTndXtJetYNCgzzSrVTygwAFUw468ZMK2TISWROAntceCfi3C3gM2F+
SKCtEF8fxNOvqg91MGd2JQZ5AQgKF+TYJxeDB2aRLyDajUvuh4vtITBS88qglqKI
wUm2WIXxDNc9FOZgrnEkiKYudjmx/NadXJCZopGzK5VnIsCgvNYnM/85elB7LgbV
WzbX3iU8UxqOm9FhN/UMLup1mXwtEDkFVlx+J+NHXgaTyCo4PVRr/fgzvd/LQALm
DXN1vZtYI8htUfYjNpeDX6iRMH7oHGJAPl0OrS5fGNyVyQWy84KNDG+7gcGcCTXV
C/DEolzdFqFxgFWJFsS0rW3b5yJL+9dP73HHrHB9yd0hh9Mf3d7l3b+NzhSgpJy8
xhVhR+yYhHDMxvPbhgtjbpD8VDzXcLGNX0U6jj2spQqyWxsxEiNaDJ00VxH2KCDw
5jCx9PEeR3oOg29iAoZxhfpFMAwTRgAvYEip5O143A85R1GKQsZohd5s/4eZaZj0
K6zxxcUxuIhv7zGWph1dW/hc5AsoXRFTot007qHpwqnoQ8VSCB87P/Yi0jh7jaWQ
6nXbYYs8lww0u4G+dmtz01ICjdDiNy8s5iqeNc5OJ01CB+BNNlwMSAumf1Q0wdra
kEpCxvfnWajE8fdskNICuRvjNbawJbIp2dsODREXeeXMGqgY45c8ezepPRN0YQrN
pvh+m1OfrfcEmgkcRKHgPVtsXvHgctxLEZfEGGHo6RMKojt6zAD94KVXOykBMwqY
Y/kKpD2iJYq7BMpmSUj2Ln6c9qYywbVeB3rce6IVUJ8zmfHAIgLlNyfs0h/Rt05+
Uhkqo5HSxfSzJ9h1LXmCZNxliFDHfbekNcdNJibvbg7XRu3jSA+dpS/DrlJ4ivMw
Hio5yXsQzKfIgksrKX/Y8q+xRM5loSPBisNhAuzHx0xj6th9s98MOUI2cJxLtcmz
jGaT2zAY3ZNEMWAMrRU7QPYUiKOXKsnhry+wLYFIYQMqaw54MMqQbmiHhQ+w7GY7
xl+SmrMknWE315zfR85H0HUHTUYzD9s0QKCULEJu5CuPofW7XUaZxWYu5t5yD2zw
+hddVX0/ltTJPI+veX29/lUXT9OWRC2nAJZ7TbDqD2lqiw+fn+kiTB9SbkfnXYOs
QiNobBhFH5GOcYIPh0mOqWSqR3fDQnbIJjgX6n62VjwWUIDatdYk4lPKvcvv0IEl
sdib775m4D1H/wtMBL3yfMf9mzq0BK4ofF11BXr5Yj9t+8RMHjZMkK/5wx1MslzO
3wNESKIwqSiZbhBnEscGz19b0H35HK2DARt4wNu34HdyAoBCV1qb70hrTvi5UtIC
DIUwYlUJacq45KciUg0Q41tfMBp2LLFxcumsZ3vQUIxVYb31ZP5sWHizVt/P8xEd
gKc8yS51sPmR7fiyW3aV2iksYlb8l2CyyIC1WyuqutxAXSc/z3KHlxCvbbPDD8lh
qim7ng7HB4OasodK8NriuPLSNonthhgx4oeCGBUO+6adOi1aluXy5TLJ5oUY8xmv
6hQv3ac+M3+mwW5BT1zfkdsG7jUlj/r2Fw/2OIba0qcIK1JgUgUvE0cA0lD6xg6/
PLHzNuXQsYrsMtIbfGOL5NJQmrwPUiFFWg9jrIdkuQSTVgyhkMVLJBpuawk2Tpyp
PNdrGsvsLR/go4MJZ+wceTDHsNQtnkTxn+qEWlh9sk48q8ngOYJsC/Aax+TkcowX
v4IPMadTwGEUYLFOc2uGYCJHmO2Om7iBjtrlUSLy3Hrl2OkMI7HdJuYeOlGdUO59
Ey40bFMpZX3S3A3YMvhZ2e4ReSs2w5bkPwf6S0RoIAr/7emucdLElDvMn5Omp2id
NQiTXed+gU5asTagpAssfxx1BKY6qE9loOBX/mtOeYD6HhC8KgOYF/Q+AoyyTu3s
SO9knRz6z5w2IUTF02XKRCMK5KZTXKBv0qBnMJqTj/e5jFOizlM9Su0FooZDw419
eH2JEQgxeg5A4u6Ycu39X9s8UBBxp5eHTRKXYz8A0MalWRxDKm5UsTTe4ix8zGWy
vm8zRQmlDgLjnZMdJvmgV3pL0k8MppK2nj8i6HfANe0tFaueJ7fGxpWSrtr0jYtz
KxvXTPO8CZJDb8ldVqe/SOBqgkZV8JLHFUvLjvb4Kb4lT0pXI2lAFm6nzTb0yFRl
1mz5XUUpJgCbXFSocztejZ9ww0WeYA74aIFl22zylxCd0jp/4iehvVR+NrLR5xEr
tfOAT9KoJzbs1hA8hePdHqyr2RTz4f0Z9DfWNlNHIseOSQ18UuF0rv3tvDuUydwg
gz1h3FfHY1O2d2FKMTXedWj7YeFNe5a6rced9/Q91TwhpjGt+UMAgjoPnRzdPTZ9
J9ysODAx5Kl/BzzQHxGfFo4Z3Lo69kdNunZaqT9Ep99Y3aAiPmgFd+S4lnKJNJEN
HyJHIC/VNw2Ov0B1eytlatytisohNf/KxM1D5Te6iJJocrrwuy/RTYXKpTfxOeep
QZD4WTZ+ioyEf7QkG7owIfMOKBIG9mP6G+4UrQoabFT+9pgEJAO+pMGbl80eY72B
wnzQNaAD4bdEoBzKiG3AhHOcH1Vw01SyeTcZdiuH4cZEqneXPg3CQftpou+kNvA8
J6R3yEZyxSnKEGVx0Mw196s/14dsAt1jNag6nePNvy7L4xZ/g+ncBOKsSq/PLVJP
4q0Z81fIsHmaaS9qKYo2fzKRIpXAfvwYDBD0V+sN10Fe0CmDxSfovZ69YDTGXdy4
fItxs0pgo6tR+XAuBNorbfObA1Ra0HA0dJOrkuzDV9mOLjxSu5E/uM4NrjpyYViW
JubwM3ujqkGBqVNCbPtrJnEtICxS2hgNrViekq19hpFooZsiQSXx564MYBAyfeVy
lw3UAJEDxpeyYDUAZ+4n9UYK/A5bJ8qTl4R560ZfmoiQmojcmeDBmaOyZB4HoXU3
2JsBvS2GGK/mQAAD5ks8r9HNOJmAQZcOTe8nNKEe3MRPAqhmkMNjshXvLaq38Tms
bkUFLDi+1L3V2Wi3ILAN49LA17Z2WUL83Zhe5gaGLPVa/ybaD1/pV1aVbbjP4cZb
6fV/cE4c19wU7DJfId+v11ZbkIU/9N1IwYmwm5vJ4NuapveDJbMCn75IQRWLyP9H
KkaG/Fy1GEqfPyfz2pwshhQUMjjGvycpl7wxFjrFl7dMSH272Kc0gHogj0wvdIXj
wAgCi2lp0uXLkK+7++xmSa4UdBI5s5fM4PxYxVGLuFxnth3B0Gj+j3XCicS9lU4j
/7tmVExVq7jO8vedWt/zs/p8zGUFuvgz3tpoQMzh0a7faIef5hSP2VL7MawadDsy
/49ueKdSa/lZ0bwhfO/5xje6bzaYwqMmC8wX65jxQ0Bl1gGOF0gcP15XPVI8tn4P
iFT0QO9UzcpxKbR+CA28u0wYyKijXkzgHnZfeJvKkgLqWg2Wz84MpAKAzrGjbwep
w1OrNSry5MM3KL3UnZf+wfIrsr/o3jiPl6DPG+4Ji+6ppLFknxuEwPkjgaLkOTyB
wu4iE9Vxwj2YSyVAz0aAlifWvKv1yFnAUygARpeBY8w9w+lUknq0amthwRGL+6gk
gL0/W3ZQVXEZ3dcIx6i2GYhzWiAqfZGk6Xvf+vVdPKWVQUn1RnuLix57WrSFg4qk
9qswzQKKWkE+NhWzrn0klzbvIwRS5K6euP4DyUtWLj3UDZPBH7B+XtTcHWO2QgsI
gNMohHzuc3z5coehnbBSgmEGz5EDz7xZgW7bSdMvn0boMoxK9HzhkFNFt3tWSQ8R
gNIdgno9Y79xeNKdAFtDDuhR1fmXlMbRf2DYDjfPPG3BU24hXHppqLM0tRs1U48h
vWlrhJJPKHqWyNsn5MjRy2bvwtHiydQLCTIK4wuWDayYzEIUIAtIIxbk/SCpGOX9
L+C37al5n97XuclruptuuNVsd1FqlphzUytncxkmNT82C/y7y1l6/99gkkdm22FX
qfnI/Ue2Lj6j6UXL0ccU2Y/ZbPPkc40tCpjP8Ionou0V5TQzFRVmjNpcur4OP26P
7lL2eNsmR4qfVKLlEnhvqRocHvI78KvjisF78d5XbPz+kzF+GoBjxBsdwaDeYOYQ
sXokpyXrbO4TSitLpelLAAl/Q+R/m0WSKLOZ1ylxB1ArpqkItHWK32VSW6FCNyK7
MW2Zz9pZQvvZ2nZ6Bq/N2fLAi9Z5iT4AHIfGu++qtqZFA0ffaBToIbzCQv8pVk5q
z/kPEps7QdiL6c+2S+l+SYhiUIQuOakepiFqE77b2Nr74eIUvXIDx7MpAh548FIH
a2/CHx1cNBHh+T2Y7a3SEDVpjIYAVj6TNqpZ2C38F83OpxW8vBVQe5zJUAVQzELI
3gUZ0SOz4285SPACzMFalNvseFbKWWWEE54VxRpxRHsKt3csvW/nzHXXIaHhnWai
w544N66o14Djd8Qb0wjpaaEeXCyoY+zeev10nsqmGVQntOOtqJkguXywtuDAZaPg
7RYKK7Rld3DzXgXxzhNIR+BVwDa3Yvpk/QdN6fIR88OEcMAS7HKjeRMTSVlsSA9A
HuUQPyYxo5UO2wsC+tiqc813wfDRc3U49tuXKfwIicjFo0S07Jns3Qcs5XnocAMM
aPv+HD19GJ9WWl6tNtzKUbQc7OvCkVauqoqqaI6paKQAeXGwuRDSl7x1RKGHFjY/
KDm3zvQLeDKbNAjrD3d1z6BEFAWZngsqA/nW40c9mj8eIOHTUqueaQ6sb7OeKyWz
N25Mm5+UxmF8RV9vNXbv6scnUFD+/VFYiDWY6U/IhT9pUjweDtjSyGxyitAGIQuN
3veTi6DQbSKp32L4g11nSFlOvPFr8lCs0bLZxNzmQONhNPSC3mKqYbExn69CXTNb
ABzCHZQ9Gn3aBD74/q0AXrPXecMui26gbBNyl7Rq2NFBDGCRKPkUJRrTDK8O2Lci
UPY9MKxVDvKB498WBgpXGBMRY6EKRKtilDLVzJX2KAXAs0IwI/LSLUdqQAPAScFn
r5a7uzWzJcjsciHexQjW6UiKFUihQMgf/NjbYgRdZ/5mjXBOzc/Ec9lKoGSNiAeo
q5IUSt9xgJPuxkb7IQC9K4qXX46vzvqGysPtwIxvqrqJg43I7vnCWOPDiDz/xxJ0
z2aS/Q3twR45KKNN111Taisva/AMXm/FR5bZlBsGlH/2Ob3zGmgzExpNyJvTZ8Bk
dJDS+nXaXoffQOiubudLxExXZzoWIG23bW1nHpigjQruY5YrLaA38LiiurVjjg9Z
PWLuHZOn4KhZS1+ifL+clpC/osg8i7Asg2aT9Pu9ChU5ytrPW7UXwTdSbTzfqMZt
CS+UY5IVLlS23FURNw+PNdbRAHsSAyc/ecVy7kL7ukBkpNrA6V9T59Qa26XWHL7r
g6F1K1ZBtTAnZEPm6ExWlQ+wma0+5haA2+HYrvBNn6oed/vdSP1pI0SFx18Ka6VX
kspF9DSwcdgiw+xG3/cUOhigptaefunpB7krRTKoVGSq3R/FIt/no3WGOv9BZP5M
cqbO1fPVP3P1piGgDK6Cule3jhjloo0W/VjmiYXPYqNByud84Vji+fK5TgL4Ym8I
DhQ8zKmurT5584a/WAbtsKcT4/qFL7dwtBXTwqKX6wotS41wh55hONDRThdio0yi
V4NbcWaIJinNiu6JdMGpdMkpQ/Krpy2Tt0Qj6rPtVnK/wP5/nAJcFNaZzYA4Y7y7
GTsRR9KA56MEzJlO2OczuTNQ1FhCCj6lkXYOu8P86L69swYxAogZEbVZzLaHlzd8
lJ6JxPSZG8d4BNOFkQ8JqNQugZ4q206snNlzw5LqmAfMPA6xhWKd3eT3M7yrFlyZ
acAHaH8aJzsFFZ2QYbeaXEyZgrN1WtyZZvsIBWrEz5dPAqQefsOk45S75Pjrkh5f
XRW2WNPg+TTfKCgOcUS7HJsYk65rturXqWvG2PJUwfUi+yqwTNrF/CuU3b93gJXT
OOdA1Qs5a7q2TysLzcFzS9Ko1SKACeyvAe37ghg4pYG5e6TRsJJXiInmn1Ydt+bX
Wg+X6/iaqTAbkTgmUYNOiaHgPO6HI58Jf611rRZmmKvNKz5K6TnNOnvaeFzewVq5
2jvqXlkQdi316PtIBpVhwR8X6NEEgqj3x68VwPD6K6OHLxgJB3Zce482b1XyEZmX
j5jF/m78Dm3t731OED6ap/p+l/Qp9GWDecAF/2aC3FZ0bsNmpf23HSh1W5nhpjEw
vAk8mETZyWMqxvB8pMxxGkKhupwLEE8NPifey4fFSA0rc/wy5e2SW6922zF//BXN
39/AQTpH4Lbef614yS2zHzqFpeliyaRA9+Ld3ZQTeztGaIKAur8uiX1+FhMYO7Nz
OQX1rmAbf6sa8hsDCl0f/dXsL9qbNKa43n/YHoZEREW/Om0Ggv8kyuPcehmyKWHG
+jPj8cv65mYFJGmQe06FzRCMB5ZRpdX3stiGC6GvWOTfZiPSFyK2ssGETyfQL3LR
xlOwJtoVdJ6UVhN3EzgbEQlddheE8RW7K1fYj5m/SALJdSmhWmWuv9xckYY3JZLO
vrSEZmspP1uLYkpOIj0O7DkyLJJseduuRJcOF8EMk9Qwd8ajDTFCv6OEFjcH1kX4
wVRypU9geDTyCGLuwx7bNBy74SKXkcRtgw49/OUttdmhjkXHqqTCZtQHItJwVKln
415yQkMo65PEa/39VmAplau1Vx6En4yYSygX5mjQ6u3nLdACGhZNvrMHHvSwyt7l
bX2XAY/8/IcYnbYD48JgS/nHkRhTOPToBnyFL7Zsd8yq9vyV8utl7PI2Fvv0Ty1J
zk5idmusEwsV/AjMXYXiqtahzcz0pAPcENCUiN+cDuZQvprMMlQaif2sK7T5HNjs
uRAzqV7wML5wDMjIICIAtV0G3qf5E2NZRN8T8UMvu+nj95S8xshjjcgFaKvogUHJ
dekQg2018LjtzfzOwiuanzlKNukV2Yy/8oyCmClCm+7Lf5+LdWLIUJp5vl+lJMKI
i/C0giIepOzjE7o/i6aYdJBXlFPZCihxbK75O+Wmcpu6jaP0y5OBZAnaSwBU4yZR
Y+JkZvJQMotbeISkNzmeQrnCFVGOVkEAgVqhYPgZwpNcQaqBMS+lA77Q3VImeyBW
y29GtrCEgvPx0rvdG3nAfziLWyDJjv2x/0IjSi6dPg6IRuYoNqChjAQlU05VGflc
/mg3shdVXuOaOOrBJEu+NF1DZxzBIpCOrXkp4qIrrRhy1iiyCRQ6BM37EgCuiCrd
8UOkdsRvRLNgiDIbKCJPG7xtSERpDSwubZEmOokcUCDd3jzLeATetFUEYR0wolIm
iaWswqQ1U6T0lywpdYWHB9abIgb7yFWxe6aPbBPOTjMNQYny/85ypeTxItNJOzc+
c3r0Vccu74Z0Kz5q5ygM0pKahy28+XZhZ7YO0IWzdqxoZdyG6/WdqRRlI+WxI6YV
o6utEGgpWLcd9FdUJi5SGiVnGULSm9zujzp1TP2yLJsQB/rRvZTYRl2UNDF4YcQE
bm7X60Vxv+q8g/Sw4qZncJDBOeTxN8GjyVGkIAfrGP/Lo6yUT+GxWpfR2AxFfOtq
Wh0f8x2Uk/pxdE0EEMO4mguewUdIpwlrM5J4grEuS8cmsO+aVTgRm7BOqkxnutiN
0rHysA/s+TfLKgWWq4flgCUp4XJyBs1X1vIrwiY4PDE5Eb+2mZEgXzW2c3ts204A
dH4JqlA+LUUIB7OWou48yWwHXSY+QijiafF3ji+78v2kRk1IbwG5dvqLe4htJD9g
pV+Utm1gJT1J/ZhLQG6wT+kh/pl5ty8ANknKPXKeFN5pzrQYOK+EBvr/QkidKkd4
lPvD/ATNoIaIwlbNVU7kp9cu3RfWpEFb0buirTleCiJi7utEyXwkG2cfw+wc8hde
3mLOFZoVSdXi4z8VPASzmBRffrODZERFLzFG5wSXdUXZXCzaQ2dyFal5GAp3cLrw
su8IvPQ6zI9yDU3Vr6zzlGSWd/wYQB7HIbHeWUjoRM90RaMgfGOtI28YGnVLS41z
0ZCEZ+b0m6vxgUWJrSThMr47X8EF2uTO0WsnfkQ9Ebx6o3lsLeS3uHJtmKILoESR
/Ci8SAFycddrIwUJfRZzIpTi7o+v8abjA1l8P2zTsk4Q/aR1WRMdsMlflrXz0SPw
V5+3DUvTI0HI6gYIc7Wz9MYL6SZlvbNyj3inK9ke4ceqAqvquaen+mez20oQacZx
SNiKhzkNDPAj0LLhPzB4dCbb0wy0jvOQLqle1sZ4usBzbRNmkzK5mR/IxfmDxa8S
0dVTEi6IKfTcqCZ7sE3MWd2aeXuaXBdsz504ZPGvXyhVi6/lzEHOo68cnz89oT10
1r8oW/d31aHDIYwi2rkwBI4n04gXN/qoLoLzdqsrvOnsG/mUQn34ba/J9c59LniB
T2SdR+CROTbxZCX4vzdC2FOOxfeZ2lj+roPWE7hWVO06lRXqB6q5AWOPJQ0ArKdV
orfR2YI6xgJPfk7AQhNn+PZeSLiNZ3Zibc04oPkVf0rFE30G6NWdEQJHNNn7vObv
lfLOe5siCSxlmTTBsHeUVMWwFuqI92BDJq+Ddtso21HM2ozIBSEzwxJSNwwftwDx
Sc0L1UrDLMy9J/8uKebWoUSnlC1aPggK7CmgAE7f3ji4Si5Ct9M90VAkOOreI0aU
xVUFQRpBTAa6b1QetuuV1teJfwvxLgbBXNkpO5Z9emb1Li+eX/PpmBJ20PiqfSc4
skIG14InCM7e+4/xu1jzYU100Zq98+8GBAcGE7LWEfWXSZmNJxqWjjNXEr9zCXSi
MBTuXPeVsE+LfSmXztrUnBIyMFRHxiBzFQRbAgprmGoqMQ5Tmt5YRkbYoGTlM0kN
pgXJEGmvg3/DcfRuZEDKvOWx3IZFPjtIqQgTj8EzLy9CKzAT/hCDri+sjZSGqhbb
SGE9vXwwKWuTLPN1EIKZ507FUnzGsB7GH1048vWqC5qEFE1xLc1pz3qJAUuI+rPj
2ppa/+xkgjQoag/hp32T5A+oTmx3kC7aNQh75N9z0phpf3vxJQ6Sc19KnUPjcVXN
TGPTT33zfJrDIikkqOq60VzVu/FUsoYLpjMmsHVdnhBIIXLU8IE/dv6wllHN1OP8
obgUUcD8SmsUuM2JcJrvIdtku5kPMuSi0TVLKMLU7+xKkgqwJfgdX5Xa2TxwDvlE
bMTpRf+URosVMaFXHZFQjAbILLR51djSbk3g3Ueh2zVDtMM76fWboKyxALGeDNDR
/6vnmZkG+nrNWH0V5oGv/1AbI+IOF8BdUb5N4z4032uYkwc867//VTYFxZGzbCVT
LgmrJQWT/68KRZd4LDvrLnCJ6TTNZJFOeDLNrB+dAUT2p8HTaEVB48I6f6QEKzVk
lMhfQFh+bcSLQaIrsdQBnJRrR1DqiB254oiIbfN7JuupVyutKDXRwchR6uczeqfA
j+v4bES9j1OdAv+9qPCzfshwfSEQiXj940lYwYVQ0VCrm/k66Mx/Fz7PPv4/5HD9
BZnzd3XCz7vJthtarlQ0XSFTV6vgh2zP8Pt1ZhBsCpAwscNeTJ30fdfSad7Xanvp
RTGbRIFd3Hl/x8N9kgOkRc0IqKKTdH/N9e0WDcPoiBeqLwTxBgmrFMsaNcsZDvl8
Rz1Lbbyyf8bOnC3TNAIxyqDttEHUw0amAcd5F2+IwIkqzHcBCjyuk0qp+GXK4JWj
uVjl77xTDcVwzOxHr1O6kvfSNYpsZmOTaXOixYpo1TVtJwR0ohHMXH0r+h7g27EP
fMLHHWPdypu+dYQtBlJPoNGtinpFfPgfE+NANCte4HbuAl1Tl4lNMfYGuwdxUizJ
xE46uvNKUe+I9dsAtQNTpfsnCOzF8ImlcshLQKtQoCt9GR4dekhy8LTVB1KOXJNF
rNTmWiILq1uwJ79uzkSAStY9QpEWgOe6UKUDbxRX/msxtGGojEz4Ccyw0O3duwtv
7QXXUnn22/CY/25HhYXoj6YKVQHmF5lwoV6Z5up56CmEnh5ITP7JBmyndBL0fjsk
3YUPMBQKQC8Ect/Aydn2YqjM6L6e46do5VU85Km+qiaCXtnE6hZoc53Vb+jf5fwY
JhpQ/K8JsmpPQAywffJBshbJGbzV2or7SAwe/BhLm+4RdUHiNqCJt92tULTdwd6N
cIYuKH1/vTI7O9v4it+dUi53ky4574X1Ncot5u3+pvkVXL+7edOTIET43CRhAWFf
JpZ8EA1oR9RburacD6kGEIGCVL59yRflMDHJNrPTSgJgynjkJ30Q8EkV616soVZ9
uaHYaTa91/3uB70i3YERL7nCldv7wlLcNsHLuT84Uhsg1i863HZjmod0ftMf69c8
iyOIPW8WqnwGlUm2U31taD9/nABbkYrdtPiFuS0c4VDzJbeokQSG7YL0+VmYIgAG
E3hFh+5+8WkU6FnUSOG4tCSFuEHnVjO+9tjyXnde7ONCp0C/FTPhusqmca5CIUG2
2JryefC4IxJoKTbd2Uzn4W/7u6N8t8U3QK6cgjqiRKdP5b7DhSnQmcoWtTB+BXiX
Ntae8eOfu7OfQRZaq0zIqWxLD3Uu4q2BA7nNHlhQEpAaTRAPZdHEQguxdZrxPyJW
/7Znx3dL4HcIpi91kU8H0IOBu1heDMsGVZ/Uptyw7FVq+f9at5ReK7rfN+Cy56Uo
3M1jxUCit0xeAq5G/QdcaH7CiJm09NEBk4JfLceZo49GSGQ5g9Ok4K+A05Rv0xpK
1MuZVpBdnCc5s6ZoiMPKCvbaz4X1j3kiUr5PeWiTQhdnTMedQiXlPBgG6uVCA+uX
tePYFRUwFs0GSYaW8mZlMStB355YWVTBOGIzqNt+zs1bhe1PgGjjBFiKntBJeoAk
sQNX+0gzN5Ppwkv3MoFj8XXCjDMLohDFULUNZ6UWjBNwXzGsGcSVP3yurDsPGGI0
mg+ZPOTRfTjzcF4xZG5MHOPQFNHekuOfkA8WzFDk2hrrapIlhFmuiYt2CghdguJr
kXF9tbSSXaPlmsPIONhR6mAjpg/22ZmJ+kCr0mybzsQhWzHVsK6L3dBTwW+ysqxi
XUJNYDc6iN5NDEhcOJ8pf+83bMKu+rtXjFNVfHTRaHbKXX+nvGpadDZpQSG2roHf
9U/du1+Fx1QCyBIFOqta9icT9oGenU9TYdHri5gF0AWUlf11JhDN/NixFrteGttO
FfrpANRxZStJ1qRcvnwI9e47jB4RxM8wWcR7mi2ujFRZQYUJipd89UuZfHHTrhmc
jCsmmXvTw4fgUeBeeY9bw1ZKWLqHVP0SM050wYpPimSXpJzXJK1qfgYNfeQGPvQf
Ctzb2siHWYZa+Fro0HEoL0FI+JmKTqmoMu6vZ0XOJGk6JGbEGOYZmpbb5OAyW9o6
anjXnB69MGFYJowxsVOlF0A9IeFpHV6sVQDGLVAqeUF9b1ezQ5ytcQqfVzn0y2lh
ZjaNlrwg+E0yruupdjkONrLsvCCd401/KKlnvRXU25EuuqucS4kRYDDGsg4jGVxO
UxyzDo9HTJv+ip6R4TmPbkQ69sVrspEKCsJbV+2/SkFrpDcyRO2rac2oWdEzZ4H0
XEAmWB3QQX0N5Bmr/5tSW45VoCl+yZXJDOfJIaS3F0lye9jyuCMkkI58WY6kq+Zw
afdP3RNeD7WjCdCNScNrC+GmGDmrCghkGWUZhl1/hAg29hOI1HWpAhjqu4fI+Ub9
bsORzgRcwUcJXRjm3SBCvCcQdfaLy4NDMmZe8TWn+1DwFzLjmOBRox6fyas0nsCC
Ud57/keiuktro86nPbEAuqukupo9ojj6IjIJxkwJaOOfOnbAkyYwzyu/U3A3d7RU
ruAPGTDqwNNRCgsCvbARFfr8GDCOlyCoK6JaF5Xr3bbBtIm7GNfOOF2XsI28xNwe
+GWWnLzcztJmWlRJhZSftwb4f4F66xHvlFyvsPMFh1lEI6AwCipMkbeqXAeTfERQ
2Ni2y4sE/FFrWTfcb50cSj7jWlqV6lczkDG3DwSBiC3INnQRmQsqqiQjX82rHVT+
vQ0xiG0PmLeVmJRe+T90gPoe0lPGUk7n3bccyBQ/rQNhNncj107+eIC9rZd75xkZ
13xaFQynu8cjuBGjAXF5c9vAMujUf3O6kaKZ9Pwx7h4Q/rZlkRa3SLkdz9uqj51p
X/8jB+WtLjelmA+7QdD/dSNUDgM5zcE887lY05DOCciD7m2bbdx1eK+Q9+rFt83B
OXGVlx/4A8Y74aBauw+QId90HrXQ1WkNKbGUIhn6u/ggKTn0VZoKoJnvENiMgXd9
apheUFpzRIhiZCZLGlYnDFhUtnvMUO3Yhw7iKqopBWtXdR9IDeVnZS/070fy0I8c
L6BStIPi/fGzGatuPiQSXZVNMmw9/tQYZ77eGC92PFzwkeekxe8LUa0Jtx5iViUx
SOqVC+VTiPurKmpTQsPtLNJTaKZIG3P0qjtrU0O+hCMXGoURRi0Y1vovfiD3UIsm
Q5Vh2ovQF7NxGKAq51QQGZ2ME/woZmQnVL6sJW8zNjQCQMk+sfjUbeHCOWqNpSY5
kD5jFRG6qx7EY1gCMgGPO4cYnYpcFKYG/oW5OlTcmFOFJzzRkziIUBG0EPHrn4UI
ORFO29zHERsFktbnL1G+QK/jKBxHSnwXcDpz0AGo+2JDm8AGZl4Lb0Cm4+BG1gaE
2ZHbZISWYxMjVGHjht7NA4ejpY2oON+vIPzII+6C3h/SqV2KgKNRZMprE2+8fSqD
zAio0P1PdrcZvc6zbdikZaE53vi5VUX68SFHHxhHkx0cRIhY9SAS1iPlhUEsd7zF
5BjZrGndAJZ/OX0GNZD42OB6SlM2X6ZRKPTlCqAPoF11gnUEeW8CUV/UkUGvyaDl
X6gB+mwzGOwI8JbxlzeKh26PNrxhBkIEfteaWINSrnxngOTVKCgyrlUsyL4AJ2mP
HIADkeuL6hLDhdbeO8c32fLBAIsfZGdrzsQ7ZfaaVTl7Fsnp00PgsDy36LOcuX0l
3HatjpXTBvKBjEjCgQW07qlwUTeZgMZGVNAFxZL1etUEN+CSmJyKaeIRS0vGYjcV
yMcET4pueuRZ7d5rQW1ZhS6E1/SOdTXhL4/J4xxIERVnPjT3qbXmqUvOLoZGkv3I
BZQj2yMzYshVYEDCBqL7JguQfPsVRFkA33hGDH3Z8K+5a4Vr9zdsRuEibA5wLfTp
/q1v8kthENsOjwVMBLFdwUkUJepoatMucwApNlL/KOPxLazNhxBp2NICpHk6S88i
FY4nuRJI2dTLoOvGv/8wiHJT+Yfi8B8HhljDIbO2UFJ+W3YQjV/k+r+GuWURR2rX
qZsv7z/2GMjUicO2b0FpWBsBQdtd32rFvSjoCkAe1qK3U7QJWquC42MV9aO7y55w
HLe7FhGos/jymAbP+bxsYziiYLlFjuA3G+pFunKj2Q96CZXGuwKVQWK9R8XfHXP1
HJ3bSpkOhtDkmGkHsUAYfbLtyl0dUbdRkOKmXEQ0NysQqExdkRiqu8YU02YbGIHO
60uu5pyNe8UL68eHiQMfu/QVr5YTsFxk7JyoNfInMmwEF0ZcahyTGdFFVMUGXpVu
8ePn7ymfUMuiP+ElBt+tXGyyHmlUM2RgAwhSvNvqmmMNuUPtxQosptS51qx09mUd
FZH9qy4XJiHZmRjLyAjZQ7QkkKMghuYJF/jvQpSem6R9i9/k8f86ix4B43RGihN0
w6cGGYaaSQGnzfuXoGEEAYTvjX/LNlbKLEJ/nJcBO7KwcDgBmAaCIwlYIkRQgW5F
GCDukgd0s+2FNJeZqV5WwlSjKjp7K4Z/NAHyRyBQmL1ePvEOSXxvNC+zbyQvb6MR
zRGOmLMP/H/LEHl2oywHijBw/2Ljc4HiauLeMmQwVT0hENpqzC1tMzTh0OPLMZaL
RjCbwhHpRChY5doVonGDBsJXIn18W2Dcn+WtiIoTySoseEs4FDuUPtp0l2dU8iPs
6uI7IrIHC42pcNPJmxp1Jp+wNABbzSNtcOz73//cTSsjH5Kafa3NXWfigWXSzzKz
aOs/hCX0NbBwMaNrj1TAYWu9jYiCOy0ceajY2LQ/V5ufQA7V4gurGQdyvkTCSrX5
hdRA9vsrJFGiwZuz1q8rSdXGsh7inGxVsEPOabbAE6In9KCVdlg2c//ry2IdSonW
yWFmKpq6xHNNAnMQu8ggj27BKBOJ3JeM/TEPTBRNf+m/Wr1Pncadg6+o/vfyredC
VhpFcsQ8oR7kLs415isCIBNNaKHtVDAIZ8PKQmWrRMeegiOdEkrExHqqDADzZpQB
ZmiFAVopsuyFwEHAKU5mXCbFNbDAi1mZHefcFOQf9wCVjGvHN6vASx810tildl5s
lODRU6xKez5STM/MstUj2rseVLiFZYz1VnywAWEFPgqir9hs/gDQQBDU0+ph1I70
Ef4Dig7AYoF9ys5axuX9CwSbxk0HYgZRIpidbOQvPUssGOqSJBHvLTgDikD4XDIR
s03SUBl4jKl+idfHP6zQjwWiSjPcuOWHubwXBX1AiSp8H6R31M8m3l2aT70Qr53s
izs27c+4IE3PJ8ZYZoaTq6NT6ed4NkXYtj3/56tBfIJs1eyqmoLlLKTQd2bk5b1u
iMAjj+wlLRs4SbjV+9DwQ67LMquuPHXkSyEX5fexDQawj9TwJj7bfzqQI7lfSwtS
0pe9QoouR5Q0No2Uaa88o/NzzAwOIXryri4mctWbs1Ja7wz97uo2AxuuE7L2mse+
lLaQ64n7bptHho41lSaVTK/gKl6o7R/jU6hEOt7dcZ0kXzCa+qTMmo/DmAhDbNjU
ofvKw1SOdIuAHbzSJdUYYbis6II7WW02R1Yt4l0xzox5xtAXXq+K7CAy0gXvsdXT
DHrTzI3PMm3MLGl4RqVWP3WMMPTPePPkmyr/IzdJgIGMbZ+zwBCQqmkIGb00RwMr
Jhn116uOIIn7uY8X2iqvi9a/eNSKv4rclX78L34PPxRDNDew+ZGJGTEZ3qsobnTv
jbZYbZOmeXSG0WJiOimqy+Qh4FQ4jarleXbg59Vcw4+Egm5Tc7wze0woiLpvzA4R
Bmk5MMpubyIYU5AWNMdR5KsX1H8fzzkh81ScstjU7J+0+3Spc3/GxFBzD+xLv0lO
JnsfdP3/2ULBHjUSMAxSYmbJExNrognc/ShBwVVbL8C8KHBZeLfyQplm1FK4YUPD
0Z5nkpP1Ok57Bl++VS4eGQaXJkt1Uh/WS4r3SFgSxiOWcX8mP29V1Vg9obgP2qFw
3fTdr+Bhg6Y8ELM2swDA1/S1sfXijBOKE1dkYSrQijTRO7i16mWXH0hS7Ae1qwl6
64d+lnEdJR0j1z2/BpWvEcYk2WZkSJYEbFKrxm1gp1PIud/YKY18yB389wtkc/hd
g5guvQ7S+mXNfVGLzFvJ/UBmbj5MnGQ7Hv789kLNTK5fOX8lZFUfQTkmLZAj6Mj5
WuoZyRRJovsndQUTKMeQn1SntFVZydz0PI52nQ1tayWFyvNRpWT+BylLM00UbmTK
fQgnkqR3r/LU4FWATK2F3GTf7UTcM6gRu3LG0+x5x1zT6K4sdwZaOeRyIcOp6THP
hajN3tEuByoAi8qY+ibj7CvdxT64k6KUMNMu5PuHMKo6ltEYkYoUBYtS9xKXpVj/
uV1J2NEjReRl1y656oumEEIpLCUWB59S293MIC+J1qGFNGLOmNQZUSh/JtV+jHnw
D1KgiyTTpStJJkHFvAfgj8l4DGCK7dbXGlMR2XiuOgnlO1a2JiPT9eKcVmCSEcjm
azJDXzxfPrnKM9YbXzZTvSL1yHYmHaThq77zw+FtK9BvWWYUXCXQTAQZyUl2NAan
rleV19ftl34FIbM9F9FHhztggV2l6X27Zde+o8rf2d7Hx5omvS0vvkhaAX8OL8cE
R44zmyNQ02RvQHsOMGC46NJevW+rg88ef2mKSGna3nNTL5LVaQ3Vi2m5yjcmDqku
mnnj2guQadkm9IbxcxjjEcMGVlZTL83B6eOTRI5AZW/XCKsJa5CwmwCWil2FENUi
kUsTV7HRCi9PzEpjinze/2vRBjizgVT0vJXXLdvk+oekrTNHiVgxRcxqQ3Ai7NWx
llVPwGy3Wk9llwOXXJnHdI4nM6lCTcxEFsVJA/WTpE231dUJFEZ3V+3HPIWP60v5
d+SmgQ2aflwTMU8sWiLKXs7Oaf3uioaHJMVBYMRCcHFTJFTKse+wc8Wy9Hn1pI4S
UE/8g2CxDnrNsPlzvqcyqHeamYp6JmeSMzDAxxvEdtGsgDjVRyL9yIc8TFMwT0fJ
3ozcZfzvTqaq4SFG/fGWlzDvM4odmNvcUbJhO3Z7+Q7yZvCNEdoS+5inBvoGdKZn
AIt8P7OXE/8KUOy9n51ehEAFW0b7gTBUs/M5Oa327KyaoO8J6Nel6/B/3a3xu/g/
frw9l4d+Orb3RJfuNzyWoNUlyPJAd+kqT0jB51UhMRtG5QDaf+atXic08Dx5xH0x
58AU1i3v8NYa03SbmYTYAXKbh+/9n8IwarTLKpN1/vvdq+VYeDd602ORWsLxi9QX
TbdJbg5GZ73VEzcEeoB56scieXVbDXixTkiozvyxPR1VEZ7QiDGE01Cs2ZHnBPBz
H8Kp4uUxHOJFYcQ8Tr0e6le6gUmpt5JeYrvdxPb0jYB3yeiLXQnfPsXZPifwVYzF
gHxR7HKKkQ1NYZyCOtbh1zhzhheOajYrV2vokZTZEqZmNtCosXEsimoE347Pomv1
l9GfJL+fsCTqjStyNzmjjCYXFbmyIckdpaOeAvGIzVHbvwh8J2ivNheYLZl4bWlM
ch8M6OZrwF9RFpGht0XTy6pT+bq/7gQpDnotS3+RW0Elcevmwo9jG8QlfJK5D2/D
mtGvlEJFPc8XjOAiBo7uE/ZVrraErWDFSuvvV1IkdBJhbw5l7ixwstX1Mqib0t/O
g55Q4dijE6sh/hEeJ7O5k2UnIPG3d/y7hYGD+UG8R61VGCf0/pue9oVa6X383V/j
kBXyW1LxMuu5qgh8nAsoB0QesaNGWYBHIlfrRIkaK0Yw0E+qhVNEJsg40x2+YRVG
WbJjqIKIbI3ruOwwYIk7kOGD7JidM4c4/uJQp83u0UeW8JSu52ws61RX704C9zNB
oRnu3eW/UgGIr744Q+WilSrBMEE+Njt6d6l34bsA0RhOS9BRm80/RVA4iFNnhmFm
z5e1EgQKKm5YydyFCGtBaV7iQ8ndbzpPjyUxxXaEUsOUZftKnxlcyN+DKWd22JIm
kTqYe3zM+SkoprEHAL5FgReBhxKzv0xu9SGXRTVKhI20qjyXO9TI//dejSh03bc+
XhiE8NM+BdlJurE6FpD+vNXz/0YT5HTSeTt4xYhIacY2irwdZJONMfNqMf/Oaf3C
pBCFOHButklTuvyqbs0d9uEs8hP+gzRdWNfRBSy2zmGWSURX32yNYCWbh99Tk+vS
mRD9YtGGrGESbcXzxif33yznDQGC7WVIGY09jIt09VdWsDLEoMUucZiGcVR2tSyh
x+9UksYGGPvgFQIWjHSfcSFx4dbhnY+SbBo+k0cNMvNyTnqCufsw5Je7nvBxrTfg
nf+va80TOI5gQAuwLI1bB9Vu22Zbcnj6/JoHtkXanlLzLPGE9FwUOQ0+dc5NVFGi
1RZrV0jfA1h1EGsVNpC/iKukz586+o7ZCM29oHnfqQOKaZPAb7b7MXuYZy/MOG8+
L/qWGwbiBjeXJwZYkTdiahxpuW458OouqfFUO/ZinbZ68KsBzkPlnYUNZzUP/A7Y
GZQiD9N4iJsjIa0TveEIepa28twTGtEGyR6spz1+6P4EuNzw9bh4mbaTOAEvz0Zz
D8n+wktkZPEHmBLR7uf9Jomy0GU8N4Jco8LVC8HZnSR2R/eR+/tdgo4711j40eUo
PXT2o7gNdhFjwFaSTrG0Qc1GtbN9gzB/i5MoAalyXGRLEXhltMQPgAqkWQqMnLIg
KZUjVf7UVrarBxej1rUOpb2Vo1fr6B7Hgy56OH2om3AJZBMb9Tba1SUo4ZfskzWq
Gf1u8krBWHT22PM+eO1c3wEVBbO4ThHzb+t/mrcc2ERa3CubTsWH36KU2Quw+3j2
kQGGeunHzuxj3dFXSfTUeRdPq/PbeERsQ4pLzmRdOLsLJjJ/jCQ+6LlhIJ0BKyE5
lv2bvV7Z2+uraOCx92k1dCFO06P+061eZ8zbO5x3OBf342UbJqd9QOCR7FVn35BA
wePOW75/n+hyW/xhzqd7C/nLWYI6sBFb7fhQyjOQbJdYFTmlfE0eIDPEOOSj3Dg7
XTtHsvcNlNnXlx+RZgQzZYDIJmnSWZu8UVyn39SFHTQokn89z43mYo7c88lFSnc1
9PGlPa3lwpzrhnSJkMXuF4K4DId4dyiAH4xcAyFmU9Jxf2Vqj4oEovnLnOhtPlVl
wsHphoA8FNV/iy6M0B+u2+YIhpbwPz7P38ieVLM/QFw/9pbT6al12NdNxLsIB16q
vy3BYasDT3jiCizPRGb5fKDZDh3oHN1dBgoe3b2hVfQXnxKCp9aneOQVH6Bm7Y6I
1Z1iwSbsjclPBJNlYnnEQ/b1QM/wkiHPIPqe0uPqcsXFsW6FDJzJNHtWnpiYf7Cz
2+3WAuZPlep06CGIw1W8AKOZtzDdRphhwuLXBQQUhgSx+FtZMOnt+VENssellC8C
D5serk0Yhcoa9oK7Co1+87CNDspgovtrDaitIOZ1/DMzXhFcFL6sqNgb/oUAzl3O
7sDhGhg+W4dn5UYhHfcQY8NvSBXalB39RuRyOf/ALDRgeenYBgBPRLMfy/HzMP7F
HmoEg2X/GvNQL91tjPxjBhhMW6RsCWZfam8/LO1IKfYluh1UTp4t2+P0QmGE38zH
MCWGlRNeOftoj2iQOkkyqZeJnkJ+uIu4n3Uj6vJIBIgy4ex9RSB492lnF9lRmWY4
6zD7I0pO8QUckvTLf3zl171SlsN7vAnWCZWCdq3LNhi1IQ7KSR9E7cPmAr0Y1KEq
rz0IK1IoMfQeUNva6fMKQ+ZnSJa2e5sKlYFgwHjXuvtK+tn1xCzTEA6mgtPK6fYM
qXzJjSgDW1ar469BGdKYLUdQQG5kDZd/VRBOiq2oO+aV7RbNCL/zPGEEHwNt0oam
a/eBUdXULsK6JOo3JnQQVnMeOk5THXvLk7ME79HmsGGoebVyaJDSsnK9GZfCwTgy
3hDdFITuAOfYAnlpi+TcfktezQhAT1cIZ8Bt4BQFgmUoW03Hc26CbLTO89LSu2wv
a69aciPs9zEZ0todA8lsrtDn0xoNJswJUZKljdOPcVx3A5kvQIhTvxS7Zl3v3CsL
pfs6nHT0vEs70zK2RVnYLVux2VUmyIYuNWsMj3NwXKrbp2uhyKTIB8FzZcy0ayIT
QNGfDfyPyCn29ruTGBvl+eItzwLOfY+dAXTEJ+6S15lKMji0ezQHEgl8CGoUKO/y
imCzYIVlbZluP05AtWq4j/R2LvhVES7KNesNJUKZWN1pzWrhS4SbKnzcDgJrWUyO
HIYQ/sKzBiN6zl2J3NNr/H0bI/lHya2tLSO46oghhTI3FVW6UyhlKdJlFInNm1el
BpV+oK+QQ48z/chNcNhffKxNIe+GfLdOOmQyJtVkwsnU/AplfgeOenva0YVIyE4o
+JAjFYkwfLrX98o/Y62WGbOQun97oDf3qcoc64PVrRRZg7xGQLgeZHwSBvzkX03C
ehfi901YXDqyQ3L9PyH+0BnJZV+44wNyxbyagNJlTg7fdQc1cSmH7r2F6JFu4Apx
jiWvcvAzjbm/WdQfIyPUxNzKfKAExdUFDL9Ph00HkMIEov7HhWwFhws904fyMjzX
ghUbvLBUFAJT3mJQcHosHRg4SKRdQXO1IbzahksndnH9pc0qXtfM5fRNr+LG5oOp
C24p8NOKRW1CUx+tqOaOTeRasOIy22JrnnM7eSnS9IcV+pq8YaucdYio/RASNw6m
2PN3MR06aRaRQ0T501P+KQMar+SKmKS9uMn1g3J16XWODpZpcJ8S+lLQGP+L2e/I
4kJrIGtKcGXttrmUhLz7FjsVNkDqNkuw+RsN/2Q1CfAkMThYLnxrw+32cLOmbVJ9
S95rXF2dnNjNmBaIbBwJ5KWvsx6T77r6Ujtr5Aek7tq0kfSCCTJlN2Z7CwbXCUdH
rEMwG8AX+fRDDT1NFc1wEWg9wRGMSfkM+CQ8YJ2tz4NKYNFpQ90xAKvPrSWvLf41
aDOe7wd8doosRnW0UhkxKS0y8xlacDgXw0XfEl+ZJHnOjoAfe53hh/JE+vi+raQD
6sHx2EY0m7u5AgwJ05ODZdCEjnc582SbPIsz03Shu3Tt5S3xPni7dih+pyZ0wBHA
joCJrlF0/2f0J40j/3NTNg1jEuJ/zzoVkh8x/i2li5PE9EH82Xc2U1bI3ioULYvW
u1GZnnOn9k3MYstaiOweUC5fpL6jg2GhJsnNlj6Vay3xBC265bobzX5Ib+E4apDg
MXVbHdWeUIiiay2tRka9LvHLImWNh9niuChzBb/dLHFORm6B0ppSqSbiRtMwRqK/
lnsi/iSrzbNyY/Uuya18g0W/IIMg16+w38OZKITwH2WY0alf8LPZTo++N/V+3qN2
7yJN4m68sFdwZENgxXrV+XqSMAO9czmDojGCb7AEY4tiw4MJ9Q/3krIGqpPgddDF
wM3Mhph+fWgsQ+nnchjxTspmnrGgPcCs6H88748sj8H1YuM+trPImzt+r0dkkNgy
YDnNhQNdtCd3VmH6DiXbTxZ2GWj2jITE9Q9HZL8aZXSF/9zfkxCrBHWUgK1GBeKm
g7Se69pDF6YZ9qEEkSB6vT7ZPcqV6xTEKE3vG6M8mz3LtviRmuiLC+3jRQhdXwu2
pPX4keNdW6M2so9AbKLfvJ5oomhPBkuq02//LvWjo0omDIyPSfGsX8ftIsoK9eO0
uhfY/h6SoEEE5P7UPnVh+XhyoutS871CB2c3jgH34iSbAqGIDGhGArVZT6apT7M0
6702+41ilq9YFe4fM+jb8SANmX+aP0YibZk54Ix0DvfcwYkfwi1Mm2GMNCXwdNYV
Up5PHWFDv1S7wB1biS9dxKewyvDfXwSRYkLQEivlgeFBwjTpqger5l2mHXRTMfT2
2D2sw8bRPMBvIwvFGyz+OWHWmF89Ry/YTdxY2aVLREfKnyanWKnN0DhSJImHrpGn
i4Vnz4EOrHxIsJQJAQEwPlHu+d211+pRVqv6KIjILirQHjsVyV+X2+bWKVLnqXVp
zU2xFhlqTiyFCiC8H7vqA6Niq/xVxxPJ/TWIZrcxVh3uwywcw2NCQP35rH48ZIwC
6WYPA9I3KDk2ZZe4YsrvDnd17Pc04dvlorfMQ9UpXUuqMtdTBHzeisnKfgrP/j9C
8/AMN+U9VVINc+SPvPfUq3Uvhfgss7HWgw9BJXOvt6wuJW0/fCvVPEPkUZdQ8qmo
sQwwSYXpnkDBs997R0FGvnSf48Z11QBui6HwbJA97mvHLpPvEAoo7ite1lXphIUc
VDQob5rX3PHrN+OlsbTp90SXfOx1YumYFMA8NEUBC4O+QcTAA5W5R8u2HCKfz4tv
+J2PP7CBzHFhmxQaIDX7gxFVI5Y5cnBMFqXsCgwle7+7WAv5DIDXzNk6JwqEsxwA
UxnTe15NOodA8NZMXlPRdNIcTwJAXTG4co1DmAcGxhvYGPniw3svpV/v7eB2E7yJ
t5BX1+tsaJkArPN2+ixKwg2sr7T7y9dMez3YyAmS/aRwgatQTEoEaVUgk5wAPt8H
lUHY2VGEBSslH1S/2Jl16930RH1554nEKQiOh9pTsdbNwwmRs6J0nQjJeD+2TRA8
BoDNa2HPvNJzRfXN+VlMqbS7PvinVabt8PugSNGKRCTKDfBvCm78oakE3cg2mwBu
+/ThVCMjVYvojcfyr3WtNN+UsyDTGSCD0ACOjtIYifxLWQU57W26zQFeQr11fvPM
hbWbr1IIQ82zxkDOMoS8tayOfyDEabSEy09KehocLdhTcnZuTY2PQIiorHzJn/eN
obsuD7BvyTzvZlYa6BeKfW3z5RkZHVtf6vTSBOyMD9wa873FXyJUWd1pr2B48p88
tQBvlXqWXHUJ88emXqAi+bPbixUmMKlAGDMnsMGgPGc7OK0SH4uqwM6wPtGKGUkg
QlSfr57ctjHe3CyhiVfFhQpqVzeaNNbpqmBpfPxNmWBzq1XtZBdOwy7yHTJVMQ2O
ToEPc9ErWimAEA11Edm9NpAaCNtmPFKhwXqigWpvJJjwS8JIgfS/Ksk1tk0veSEn
/BWWnTZbwFrHXNzD0zMV1nedHClqgpQ9ZYD8+1z6dhH99PiGCfGMqkFJGseHJuE9
+SG9A7oDH7zKLvVoWe2AhEYKNm6G3xjWeN6PAbFjH9H4MU82doOpjNFBDUY63bsp
xvKWiqUh9awUEOw46CknJf0K7bSA0yeru1JeS9ixNrLb3y6K+2HYsteCwqWv10nK
gXhRQHyHpWGOwFqJtlMMhvFxRJu6MBzKutPrLoLMDk18t39Zgf5oic4L4RqUe2Hh
+IDGf9nHA/SIlnsAds8KydiRtql2AaXSxYhsM0Xc5dufbFVIex9X54hyjtzSfCU0
/fMeNkxPA2O/pZajglv16/LeWOhEyPV4CotMreyQWnqLFvy1gnQq3ZEqmFnu9pnc
FA5IpcPwPuRXadn/GjPjXfB2qpUGrEGP5B+X3iGkJWs8P2xz+/emxKwW0xAfKaFr
RCsSzkG2BWd0euB72U1IVxLZJL87doW2mJ73/ccYsQL5Vy3Mcy8orhZ+p2J7KLwZ
qbtP8HbeCygtF7EhmyiVFeRl9r7B7dAcsNHAtGHaO5jNioxHlmIFzLRodwjwZEdd
o9CiSZ293mAc/2dVUK8X3kukL9oEjBaB+nRuR4NwEZwrHV+p/rg9AYXzcSUXPeIx
LLcPyAovkFELwE3PiY8NK0+CHlu8TCGpE3OQjasPOR3kjwFJ+HXFfvz8z7XU+vD2
EM9xGbRI52hzTngn7Fs9fb7UNeBQxI8zptCjIxXNU5FM8eAXwDn4p6n6k3vpu+GC
nfnZB42RDw4QzpL4Ge40Ti0U3v/brBgPd3gSpd93t3xz3cvu0dG719guf0NsNDGt
nro/piyKf+NAwwGJIPSdjrYtYVskXHTId16ST73dnpWtbWArH1/u0pqMBu961ncB
R2Hm7hFf7kn3LuWMJBQBHXCnWbrPoSyM3DOQaOljeTvjbnjpbmBagHWADb+w5hdT
tJ8maFJrCTQsLUAdL3AoVqF57jX7/EEat8q93Sg5fqBO8kAqv9JycZpFhw65220X
K773eFEfLfclPWQixeM3K/9vta73bNPxOmvBerhrWTIxy3BdMcDNuwi5WLPMHv4r
+IQ4nSEFAFSEq29AJWmVrSsDSVf41ZnzN+/agjGCV/BPd+X6RwOAz9UnaGb8ml6M
gn6Npnqp2Cjy1T+Esc1GREHVCYZ2O0oGvA3YeYYMs5dXKyrGdj/ZGqyv1naGFYBq
eso7wTUkBTOqyfBJe5NF4C5J766EoU2K889CCCRCBu/qWE1Vd4n5bXOnYwDTw/Bb
ruo5jIQQThY8K6LXvHDR2PMT87GVqBgURs/Kg0nixW8WwV5kLNJLOPAh1TV7mgk9
ATY9mw1z8swOolW8dmW7KygpwhXEQsjZZMpeLbZ9Ej6Q4Imhi+sD6waeH3D9PAo3
oAI7ZqAYDBmfEgUhgtnLUxS7ImgDMxQj12dWhS0jD03XQpxA1d9WSqVD+PsS38Kn
BfI65JYlwRBDM6FD/vhUG23UA20nfiVyQ02IqvZdOjdRw3RWTSkMia4qgzHbQUaO
yBYemrsBUx8E7so7iM2gYuCuIQM4QS5Of0ssHjh1DKimzTxn/9c9dH4hay4v7IVO
Vz8fnW4f7Zf+9TJB5HPMf3JwQuBcBSn2V/2cgyxu/kNra3Tb6hUrk1We1CnP3qkV
+KVhsaJGtgqVjcmEADvHQGdrT7ZOablZx3UeHoYHRUJ1FzYe0XluYXUdzjVGyafx
f5iInTIpVQyOTejaZsZxch/p38OfE5yNaSHuA09pMi3Az0yW4wyiCkyV0zhlyZ/c
5SUtMzvxleYHGRr34FanU+xUPiut8X8aiEhDBW80ti4OFlIWlIO7+bHPMnBbQPZQ
SGCT5zSwX0RKxH338fIjUQAAp1sBskRqwRA5yT/JLSzuxZfm1qBNF6dniH5t/xZw
VTk6jgOEVP+G+61NjfE8f0CqdLHtFcv5j1vk8k06byRKXESqA+mwUuYxps2yghhM
lYjkkPbHS9N7VS5PfbzrvBjZXjEovJ4nGicwFQ3Ps/lyN18zYPrd20JQQEhCmK8C
sWKMSWHxwweERAaudNkOurElOo1L7lh1Y1AdwvgfQLFtCKALZE33hwkJSOCcEJw4
8Ptjq/dWyk7kbiWBbqb6wxoUy237d2IPrF48zilWfUdpcPs056OXtyfzoruZzkgG
mcf/EMgq9LhkuqUKtMb9lBSxIWboK/rlnSJ3ZLEAYJzGlwan/GEvTu0Eqrb8nki1
2X/t7VBLsdKkW+v8h9ksn5kT/53rwXRcS++hs/PlEDI4bDGLz4p/or0TSKGjeUfu
GnWPTAedjho1sV8y3D22p9VyiODJqabbAyB5E99hnr+RjYsyqAJnYL/2cNeGnUtp
KRGZZGRu/uQLfRS3JcZZs8jFS+vm1/j9J1npUYtNn+F8Ps7MAtC7ceuvNBCDq6MO
a8bKXd3ZKVBeAJ+czwT8fzR/QpAz3+IvgLAQKvhXXPD9LIUm1El0Z7e+QCJh8bcU
T9KBrMHbWS3PS5j8JooqtpBgu6P31K3M8LKhsrGRvruLLXM9beE1rk+7zJxOG20r
2SW/OzM9EHik30UaSoHvrLknwBS3XCVjRgxVs9VthvupKle+f4lUMJ5Arr0pj/nf
UrrxPMaLjxWjC9iZxR6s7e5H7/lSyhNis5tyyn7yp5nzCQAkA7dQjB9V0sHgq88c
Fy4EtcSdly38Wg7Rgt6Va4bDVeF7y/wM0f/tBEjfYkVMF+UajVCFKoWIprXNBetr
2IfV/eoPIR+bfMB64dpA7LWhckSJLv7Cb8Xw7mijjZ/5/ML1wKVJPLwxg+cAomuf
8aloWOn8s3CpX1US2X3L1MpJY70mtrAYj2R6apSABpjzweZ9Mg0QnOzFLcLwGPtJ
GJ94sztxg21xoojLjWUw6faoyEOS2+riAjOWF18ol6pYJP1eSI0VtFqm1dbZ+CRo
S53E0TxeiqRMHIkT5PhPoOP6AJuYErFMYuEdOV0DjZV2Y50vM6oaRptNAl3XDrjK
n6BA+SC2Qdxb1gabxDyCNoGCfkp5IkwE3QAK7luuE7Ye+XpLGuXe0Lmz3iitspxn
rntcjXNB1Q73jXxLcNvIns4V6VXzafCyYz11Vxf84WVLQxh8R++J98xMkUVa6JVZ
isdCEUm+Zf1c6IcspV6SryviNgWDeO71wXYIeraCeJvAx92Rg4CfMnD4bFKxg9FE
h4C4gA4fHgUrfKc2dhc2UyfQoSvWBaBoGUcVjvlK9haQwb1eXMUmJ9NC6WSe7X7l
S8H02JDEy0dq/+OBFNuGHfinRnZI7uZf+7UF+/yhrnszQH6H/s+LOH/Vf73XrfbG
q3SUi9YbZxeov7keF2090wD8fSkRDGERxYhvsDGe1wzpQGBQb2LeYGw9DE6LfMtu
QUJO5PBczI8pCXHktkn69PO7VXqWUdj+ZWfpME5iXx03AARQ3j12n9XXcdSnrYAs
eVZudQJ5goD/GETWukDD2WB4EOwyFSUDpGki/7Ji15diMtnUibR80YHfJGYJuL/8
dk+9d47TCZm75PK3zFaPBVHCRWbLWAKfpwLdYHJCaGBhoz21jQ37fK+WEqGYuX+P
LF1g+IWt3G4W1qHO4yCc+j1UG2hZouqB9WwScvhIYg/iX7fprXcr0BMsbIJtf9Si
ZIFiXv8ZpNdiqN91gvmftuu9rVMObAK+AeIFRYioyloGJJ2aHb1H+rR3gbPx6Nxz
E/N87J/MXTxKkrWp1pNUwNgt76IgHMax9pbX/NKw2qmaJn5Gy+SXkh7dJG3xJXM7
EOcZhJhswLoFfZaUZPVHekacxkx1Vsjui+8M31491BK8Llre/x56RjpTnlY2ALMI
trdcD7eoba+EdfUKjWf8SrDY5CtoVeyo55HtemmhY44JgZmQym3lB0dmyCaknZ0j
90V5AQvfWK8Y/yp5c8yftgGQB5Q2j+FwsRTzHfVdEeUgq15jGF/gwx7Y8mByYOtr
JgSNJlovwyg7ByDHX2YEWYvr51U0DpHz7Ed8ptqj5j8LEnb49GEazBZgX6oUq5mD
03lVaVj2QjnrcBFGR2dUX1th9JMDaDs2B3CWpqxwZgR0/Kh6cRBrF44Xh2/8fVrx
wECSZuZ0eEJ4zSl5ldjrC9KK9aG8iqtCwfI+ihrY6eNh/AMbAWCNsJOLIVeXC9jn
JMlTnX1uK+fVQt3l5mSTGgcvS/JlySvEOf2tnwT0pa/eIPWHO8lGjKYqRqDkggvP
hB2Jcn38a+8AoG1tlMQwXx2CtS1GmqiOs5ZwD7ZgUkW8OGauHozkBktEUasV96mf
cXtf+aAZAQkpQ6nhUJPpgHrF9RjcoD7hPqUmPZSVgRuxxjHnLEojmwQRU4ViJ1I9
cGeEEa98+mCTKwtni9KfQWCrtDh5oyIb1fJldNIbIo4XC0S+UjteeZrksIbaiV/+
92IHB84xM6d9w9BwM8GCubItZqrWzg/Mjxo5SFoqBNBC68/Wv0tHCW1kvVFpHhJN
H/iUdognHIFHYqQrHXO+LGeoARVHpZlKTz6FCFGclHcbrzDc9QLkzmpd8b6zTTa8
HqJem4/jg/YmC6gyahSHZIJgjSsB2qnl5YPCzbG8ApiFW+lEaOBKrg029Nsik6/k
ULn7Ek7m0MEAKkn/QuJVNqnM5SYoJomrL15XMfRiExJ0euPy26gaQfKG0VxaL+8M
h5CDVvkNRS3nhzWBLa91XUXzvnBAHcOXnG00ZWf30oDUAqPxFRKDLKf6NESxI0T0
s2QuZ0yzQwIarCc2zHKUK8HYtZ6Esh5nJvZVXBLIGlNmwRgHRm0ktVnUVVAL6skh
voCH6e9GyigBvosH0MDpVBIPl2zcdM+BeHccN6DBGZQ+5Ij6svqzsK2A7mYpb0g/
cyuAyv6joJ23Eihlqb1N6ZPdSJBXTwq3Ifq2ST5vQz8UF6junjTsImOild1T1Ccw
+ZM8ousNjwCp9+DIysqmMhQdACWrhielddAO1XcaZeSOshhx/9/Efl1DAVyOG75g
Kqx2B5f/A2C9+2rbDm30sD1mPsjzPncoxUZATAwOuFQ2vPUSp1Hj/FtOmKDupKRD
FeMhgFjtADrKRZ9WXI1o0JUIMVVm/R8VyIq4mebcpkK2jRBZet6hZg8Ta7aSvej4
rnl6VXWvGolaqBD4ZNVL2VLVU6z2YaDoWEp1mIEtvTzUabLJseDtWC+6dcOZQuU8
dTnbSuFhMOfkfvh2FD1TztFQgIUvm7SVs0SGWf8gEhM2lJqwZ6ngHKdk2WL6PrNV
YTKR9Zy3Bo/RFn8HqbHhUkBrOsI+sMOlIu43+Ouwu2TaJy3qi92pgBH/kllayrs2
ktH2QQktcEB/KzI1ajcVv2Mi5BmAxWlw9Fm3bQGhRjnGQ2CoBC7U5Q8Y54HjSA17
Nq36OCigUnIYyZMe2g4p1wXEc6xWZy/aEJDy/FnWNDoAvjXt7Jvt23K5jo4jCKOc
1dgHMV0sFQGHKolfBFrVaekA5N5BHmODo/GLKp0izjXzM32BMG1xAvYmPmiyNweY
VnUtXdXT9PRJd//dgFHIqo7wDUrUO+o8OegOrtrBLmT0/DZcLPkrKPz0DO1jDiSb
qFAulJ3m6zadlZu1jkOL76P3VZ6VFWXDjdfH9H3rW2S2EcSwdJv1kAp6WQISWyie
7BAnfzoDaqZLgbq8S6aLr9o6ADf9nYa+EWvfjvp1oQTUOU37DsvHgd0sZ+olvYvX
z8l62cNl1/j8NCrd9AFEkQytXyuW10dYQ3YYMW2K3q3DEEFv37XbkY8kAT3Xv/vH
yXeuNj5aJM9LfBBxwRXpJnSo4kdSJkNnNaTwrCA/FHE/ty11YQjqVKIfafZDGWjF
HXwgYRmvaUT9Ycj1tjo/+ZJ+1VBzoh9V9ykHe5Pdv9OnCUHMZDqEu7yPNj6B3sFy
ZD4gnNbg+W0fjGwvrbeG26Se/ypllwyfBiQswruKS5tDpIDglnJIIgnKGNejF4mW
tonQRGXhVGQDnjwOENjUWfd3WAOBdFG4Rq9j8plPMBkjXWI1eR8WZT15SNTfQN32
ZCi7KEl6QT1ky82ms331UHkM3A/w2iq8PjbMC1RmyXvZAFapi3Sslhcrjbr7Rkfk
jvYpawmFtqDg97P/TNBpLM5pFmzGe4h9EJ5cB6mZqLiqqylXgqUwjVsVQfdT2ddE
YYthn6TTd5s494W6Gfv7flXCkWpFiHNVKB5ksctCLQsf/nVA7nRSgYp+1tH8cGIG
jHOgVMQ8xqt1oUaGBmFGMJfzHeZRnJgjp6fAh9IFR7bnna6FD+joAx0NYbcBk7A9
OF5mWvf01FfEi0P46/WOCM90CGKLGq4CB3Ko217bKiit2rgZzS4yYy4EXBiVHwpK
aOfgfVhA3SrLAsNvQrLa1L0Bma6tQq2hkscU3qYjQlKvwoyQYu/Qt8WWDcr3q02v
xYHPHrQiG/TOkvWMAYdVzOaHngYYAzUgnKFW4a2EYLJ2FydTkoYW0UhVGGglL/Ii
jSXpZpbkP9SCOGwpFSV5sBhprQHy92lm0gg2vJkQbwJxdT+Y6nUZVlU0GvZVuAHo
LL00lTvQOB8prjMnRI3NfmpZW6cU8V1Afy9RmHaNuB6wJPoXFemE83Cj0i6Vo+ZH
p5ND9T3lRmlpzphX1E1yTIqMpI1EY6HGLK33DpQ86xmt2AFxuIE5GvA7vWLRAFid
3k/IRo1vYGGN6fdgkyymeUCmmFUBM8Z0nliq93eaeKSwoZCS7AegJYYoHRuhNmvm
+8LkY7GAcK+HQWSpgQxNKU4zfxc//JlzADbvjONTbxl1f3Xrcx5pZ8bj6kkEh3Fi
+4MiU/omaMk85/2aeqq3s2amp5aA6wZOrz4R+SaIT296W9IggTcHcfRDaR+yavD+
FuQPyiPleb6nZG5+2qjr9c0Y+pcTh6omGnMRxxTxgdFTG8gSDx59iTXlv3h+ynE6
EvQdVLrnONoq5H6FONpGSlP+n5cqgv7yIS/+K5P5OW6dF5H2ue0LJ9V/LigttTBk
UlW8zO58n/X9a7UJT5tszZMylVU/YSXw5lJYba63zzreGPBMd7UYZbA5IocHJa0k
w7RS6hIDiYnhnYqN68+hB4cYtaC65dLtswOD4hciG/EqgIOueWazJTLSOJK6BIeG
Oiq5LMiatYo/qQGnME+v3SJ+ZIhf3mVR0g2DV4CWLxBKEe+GRTBRmvBbDIE/oL0W
mwQh7e0D0Q/+FJQh+5tpUJKdDU6bILKWWL8yZT8mSw3PZuCKOhd099BPQMaCukld
IIb6D/7Bg5dmrBAimUiZ9znfJ0LK168538N0uiXeC741RnNqeSkkKQ0ZgewAZdKU
DBJaqcBQqDT7bNAx+FPU19odP/NiMbutuBXxOwew9wQN8mNZSVtyR8tSJBlG1S8x
Vgm1Lk4rrevrM+hxNG/5Ohet4bKVvCp6GaPUJIv3RInKKKVp9brPJzPrNyK/M+jK
meIXx5m1deqNu8ca2w8ENApmUH8+Pqf07rFaX8zTURpqQaEmDECDBUK/3xJvWgHM
vITfteyuXQ/dOnk9PjjYiCP5HIDzL6ddtIthEwoLCZlyTbx+il4UwRK4ZOnSjndE
IadUtoFdn2I1M8p36Y5jdb1xF7r/TKSNBzXShG2SC9zVSdBYN1CLv2c/aTjgb25+
6UU/xj11akTaeDn/CT0XFiTRIFRNG5TkcNNp5tcs1/Wtzl6BenMvFqbBa9NXsftI
yWCuRyG+S3b2Rhvbr9vtt1GAxSj/6fZ8LMBzVGAUMTgW4DKC0tK7lo5BfA6Xsnf9
9mjpxRH4IH/UaFOudri0JTAzFa4yMjCKJkiNjEFzXOj3l4VPPlvZCFssAl6Idn7i
6QcIhPaPbQupKrXDfET2YjkQqVoFAFMtMsl5EQUbZhB7bTFsM27Of4y23Obu4rjF
i9CYSd7Ll70aAlqJlMYhAYdLxWeWpiQBIJ2C01CEyafCGY6TjtTrD0fdqmrHNiM6
waXUzJf0E8z85s/AZroORzS1IhEKHkGussZm15zQLweQHKwWVgzuWIhanHwn+MKP
SfJ6PAtDga1Kjv7oRNKiJ/8BRaoC6PZFu0cu/Cl1GUYDkEYfrSFwPnmOd558rdj9
1NoIjLuj5a1EqPZEMtUu28jadAGM7dXgMAOY2GjpOgx5x1/o7eMvO8V8PerQTDAx
VI1ydVTT+nW+zva+4hrTI3KuaYwUVGmmUOIEIpOrg8zbS76HbhIbD+xYggUmcajU
RBT2XvwduYUOyAaPZTAmTuayRefXxMGoiSRwj8HTC11+l4MJ5qnn36yUjTWc6Lz+
AnTOMBPOYVXtS0xC6XRYJnA38wc42vK7F3E9tx4hgFrDB2KQa/DR3jkJylYxyvxP
gX3ogByitQRSngSBvCqBc4jVOyjvm0NXxifAWJR5+YLn0kwvdmcXfbiExwc3oz+f
3g2YC3uijiqpqm7hmLFhi3ixrsDCS46T50fCCPc1uuCjbTEKGImWArN3JRl8kwnu
+wUu7ZnHnIS/aV/HjB0snzoMUd4vQHFwUP9c+z/Y8ChDVxeZ7MqKzUwCMSRvL6Ux
YIvwPjFN81iIoPGkLpyB9ClR+hVwZYDoz2+rZDt1yN+gR0CVpGpaeFzyQRCfDRNA
GBLSyBOd/R21D4zhoSmGQAUI7x9tRU5aU7LNoXVEGVXGCcrIL6DXTbl/9gP3hawd
8c5Kd4pdkakixVGe+e2SeuDsZlKx4o0Vnp7iEgOFRE4GrSTxavwEUTeu+klOLqcs
GkGZlEjF6wnHArXDA72FEb8OuuiG5bjjtZQArazq21XFct+ccAqVJFpOrGSJ7XEa
oUCtWRbP7h3IECaY30Hx5Hy4YiehJb7n8WTFPfgCtM3Qqq5oenjcuvjj8CoLP6Fr
VwiilNSvhOCfkSMH8V79ez52dICu65stWX+qOsb5S7kaOvvkzOmwID6I+hE/iZbD
kw1lNr2H7/zSvfKWfW2WIFLz2lXNJLknF2SfB4tjum8UWR8UxA4fF1M5YJzxOJQv
8/ywL0B+LvaFMiAcSmsnC6BVcmSZzJu2YJf6Zx5YU4cw4ac6KCJtqoVfpSbqscdF
YQqgwbTkGf/i0bou5O5gLeabvF8eHDJ+L96D7t5B/k98ZhKLZ9XN5pNAte6gWEmu
LH6E5j87+QQQxyEs1g+jYGnh+gKWB9G8mjZbaSRWcw4UqAxAI4KqdBE3ejPCUo3C
WtJ/4xA4azS6W2CSXfoMTlgUnRMa6OVl9F+EqherhUcS2xLdjf6mc1ZRc6oT37fs
dq+9WxnbB2o4spfBg9rqSAIqgNn2crupPcTChetpHfqGM5bCF1hrxaIaG6emFiZO
eLIDd7GMB3gv1ehgLCRbT7a+fFH/fc5aQPbo8mChge7YKdLAd5IhzmtJ9OKnc/Qd
cKTcTTJ/nxQKkxqRkjhDQvUXHJclOdA7C12hYSGEG7ounc9SzucgJhcAR8F7Z4k5
vNI6aYlFY8l3ak1G9KuE9oG77ATy1QPPcqDyBtSqV72XsgjWYNqSZr+mJZ3uCGWn
zD5b74RQpBuZYcr9Sf1tni3kX1mm/OTLi6+m3BmBoxbI5u+Lu27Xn8oQho2Nwo0x
yIAI+b6nO5BMg7BBQov33oZWDa5krunqbC90NdzYV77SczkkHzyHmbcyLt3dSmaF
lPDQhKh3rjJn0sBabW9iC/92rFvOdd336Kn2VNVdwxXVzZHNZuVJ3LLLTkefHL6E
GtSv0wM0pn3Mx2IkzuYeDlMASml53l1+oa/E4eMsyAPEttRkYAWB2A90H4ICscPR
u0LEcFDAfJNbtuazAXRrPOPHTP6jFMWoo0glcq0ANq0UsJcvpv9BPgMQBFqEnEhA
c2GPWQOSSkBF3mVjeTK9k326KcO+qFK1ZQkyWsYbwXX0ofUlKg4cY5GzfzKsbxC0
cFFxRe+f31vdNGhHRa7DiGa51e4SD0BbOxwISadpb5B81/UdybK5msnbhsz8lVJP
dySE2ldBlx24qUsC3ixljUv1iuxHWGfFWrTqgPoJT3DQPFk/CnaescyMw3ec9vJs
cR0eaZ+b7Twrb9R81WTBltvMtO106xtQY7SiI9DXi1mIOttm9zyUZWM4hAshVjra
rSstKRiK7tGAXBr4f+19SeTGnL7mEpymudI8ylOl7hCx3iQfvVyNBNcRpK28aYhn
vRUnuhtZjY1MHfyu0Sya9JKknNqYAilaWWs9tUtM0kgnrG/ZEDmlNy3wyPdqWoad
/EnvU6bBYPKPy2pL8n2rR4/KexPNreXSK+xzQx/zk9Qwpe2pozWT+1XJyYciKKrp
OBDgrdHm6gF5qS2qNKT0Qnrjr3LCAx0PGw6CXouwABkT1S1TWNrsTIve14EOmA3G
xXlkzfUoTgI1IB5mAGq/ARBKcLLBF4YZvm1voUZu+gX8lEgTBN7I9BhFB4yIs7jM
RYGOopklPptf+4RMn8dSFWjATAmgnE9dBBmlS8Z+60RrBueFA4s/zGvDjSbShfAU
ukAt5vIYgp31ikBN2XYK3YJjQDhz4jmSqxDmauYvzsGk/dH4U443MVQ4vPvWpYlj
Yu/FE8G6xBNlb0XNNfTgA5f9ZEDUyvEWHQiKe2qxgSzTAnLLH8g3C+hHYIqo0t05
JLS2PYASkXi2rOvgP+HT6kA1O09ovcEEBbdbpLnb4jVm9F6yCnFhZD8vtxoaOhYa
zJqTqtkP5pJbFUGY2eDzeb9kD15HxGjPwW/AgTLvqE1hboRRptSXmNnTPi2EKo8i
0bDyvPbdJ0nFEtgQVZnWX883OjRljQrFqAiKnXoPxMFoAm8gwb0a+X3KNxZEA6dG
pBRkmGNow/RWf7suh1fjwrSyEm6RwdwVugh1MqYSudxWowQiNSe1eRhultcxXMaa
sit9A6qGnorsaZRIf6x0v98/GtNT7fpwubpcIXAGG8/7926zQzG0ZJn669U+JadW
5Y8u32brnfEsFuOwAUbQarZTYoTG7SVYU3ykg6YnXWPL4AZKv23GVAwZ8MuQ9+WV
PaQUE/D4X9PHjPGu6xodB1hoO7tQCR1rWIpVrIMe/iAjRLigHIoZMzDUmTH1Wl1F
EL21LR48KKlLmSL2pMHHo1SQXM0JJStj/3vSe6ErSl45+Ksug/lIpMqCr6yiav+Z
ZijmyAGAngljS1V+EYhfeDVt0ursd6jJHq0CQRoPDiEA9jB8Sl4oTopcR76qp0Cr
BC1S4UkIQsWNs+9AzouP0RF/0eG4kPaM5vRUEL+DvTeA9eOX0mInFn/dTIlHYFwU
hlctzDNOh59BB8R7xhfPgTR455SEX+nN8vf8pt45zVyq6BTEJr00NIEoMlN4ShLt
C/ymd05cX5D/kZ91+0OHfr0dv1muMyciEvF+bXsAkeD9r2VUlEzF5D0CHgphthRW
+7BUc8MJ7/9YCBJmaa0GEg2x5MEXIwVv6fnToHoiLeaF7rJ6kKqu4x5bJ+XL1Sga
TQ3jYQVTeknbYd8M07SKnV3q86/pHgV+Q9/UYlwCmsKTq2mQk0KLNlKgHIpLBbKQ
X0nZkaM4Bcl7DyLQMxi0/4Jg5r0bMCgj8R7Mx11BQVUZKokwn8f57Rvy+uuvYlXu
wl8DAwxI7M0F2s/JAg+aPv9yEHtbbt6wFN2Gc2P60AWxRhqnvAaks/6HH+WigRbi
UJCR1EdetGRN7dxTqb5GEiqen5LwlbOe0DV26DqNvuZa/JcPEEir8/Lw1cBL31QE
CMmqru7d5BeVmthRYq2g+GznTju3orqWu0Ow3tYOAuOS1CVrxq4t/MSNqVKc3GnO
nxnz0wrwzJIfwVoGLDWiOLTqgspCe30auWN4mhNiVheNlni7g3ycFgLUFcGE5tK9
kizo4sz8PWy3cPNQ6zNB573ESqv4z0aePupr6JoZX7K/azQDfMgzvdHTLoT8QWcm
IZ3G4zSrC4lalFA0oUDPj6eWWG2XbuZg1GVSdXC15cBGXyXRfgegNulhkRm6ZrjF
aoQnVq4vWV+66OG8Jn0maQ6jQWnWSqcUePfRPYCfxfyOzqZHQawv+wGMopcs4I8y
mwlPKq92qrApv5nZ2+ioYQFYRJ+yVftJcgepNwoUi4DNsmm6CnxlMi3UXIArf3kt
q5IT9xIwsGNKMBRKaM9D95U2X3CTb5gY+9bjSVqfAW49mfgd2hxMVc2UHtqwE+lc
jILofrT/FKG0avOOnH4Q+3V6IPvij0Xtm5TnwJVUl/nGFTEmOELUMCIcmiVvVQ4w
7AHSQrZ4nCxpQr1WKhv1cw8vfhm4KQy6Sh5mPorMpa6gQKbJVL6VeP2XhRgjbpTs
NcdZt37EHLNHRPY8z16Wf2GOq2Grj801jR4khJsDRciWGywauH8AzTkUsBYq11Fw
9lxo8+UO0u1cm+lh5o9kywfFpKiQTKbDXsR0l7C+Iertv8DwGtvZusgJ/N++X0CZ
tC5UjF3G+437bjl9WcPyrYD+7p+aWi7+3e++VzDEozlHe2h2hgQI/VPalz/DYtWB
aXj5vwASoEZF7UiMrJndhEVlKeMIHarF7/9TWc8e/mEP2RmbqL4DGohnb4cnWwCY
EaZC0BgygjuKtm781Xozraprjya55H9KTbvqstRvLqjci6rujHFbkU7PNX3YtNnD
5TrmIPrgP/1IeaKPNeFMs+7Kriryah1K1/wL3uFzqephyLt5tTcKUIn1jTSCPNSu
yufDn05dd0I9VrPz64wILaIxEs3Tk08N+bkAqMNi0s9E7E0k3dEriR1hEGzRahvD
2LW18OnbukXaSh0J9M1BkYJf1CrynloDO3YaicRMfVzOzOrHq90PGi3rvbcFTZd2
4YGVFRzoKAaCYlL3l/hrN2J8sVvBVCCAjp8zHebIWY8ZF/Af8QQKJAY8qwjrATI0
1MPMNkjJDXcYcyKUjTpQ+9K6Lzm67wVWOA3wmK3fwb0YVhWy7lgvl5VQgB+9ExIe
2K6fmeycFIiqqWCnVS4kB8yW/UXpI19tv46xLBu9giKPI/Dt5ykBBkvzfmBz1928
RLoxEwQ+N2qkQF/NnghdlwsnTMG7/fXJmsCBXac/gEvGdUKPmZ7huRCsp4/gXiHA
PTnyI24N6BhcjvWTL8hwGyX4Q0VpudMpOHxlrOwRiuwd3bJUC4X3EQ1BQEnLOMZb
8bCz6e9LvkgUGAKwXIVXK2EHajGCyc+mbM6eZDNDRKUHNfLpuWkXVnSUJsICsLwj
occ29LDhLpjwqOFIckrUxjV+HMsy1Q/F+167C/ab+B3ulDCUJOv4N3MD8szph3Q+
nKFky9anDCCy3/3k0ukgLc8pvABnitRJw4vMA/a3Zqdm3S7N6dHByGO9B1uTFZO8
r1TKlMQ7IULhsBiJdw1fRkHMcxi7kUIO9E7Um2Gsb7vpU6G3un/uAu2bJXvqGo/r
ofMb5E2s2+qhOCPXK1Wv3WWXm86apIOLc29CjQCwsCMHmbruJ3PMYrxg6WQLCnFi
CAersaMIIWDNt5JwkxmTmlLMG0D9hXqazZfCU9mW5zeNVG/kHvZyOz6xzVUA3vjX
VhcQfmRrl0e7r1FLh0RTM1oK1thp9SWHmKN5jrTPkttH9nG2zz3g/6Q069nJRdOD
c39scyrL7mvNoOKHArWnz/3lgSw5h7GW7cMX4bRg3jwgIMq6EABkYkNGVWTsoaf5
c9e+RYhIlK4sf0J295iKvXTIKTKH9M+LxKULDAKIuyX0JhkKlYIioUd5Ywau+MUc
SNGyKXFeKrwWTxo/8BdXTAb17SosQuwR+iHnnWW3aCMgnodc4V9BeLT0Hk//vOeW
wWgjc+DAddAE4MizgwdEuRjUnU1p5xa4WLXj1IW0GouqJGglNvTvVK9KrtQ5hEMh
29/QFd5s1heQZ8c5iwzWGbg8jQIHtCeuWMTTLztawX+2Z7sf+BvRp8PifSQtgHWe
UH5ZaCTGPrtpmYMv9x1H1vRbtwuDFu9xR3oIywHvjuDKuQqxe33hfWivpUYy8VRZ
gDeWzZLLUr3Qx1lGMy5gz2ovdaQKVcVaJbmUfBvO2Vg13ms3oi7gDj5sY1ANBOzQ
EQd1saTYwE2qoAjJBLIWbeut0sMPDXBV/SxUMcT76szUYUywh1wzFFN5ubO0/P9e
Y3m6t1CFKmZSLOBvi17fWgxgqsYPkwFoUq0NRES14YqHGlBnHL+ez9E8NDumZMfq
FaUCNbxuYvTi4Y7xTrkPD5pCg9Su5NfCuoAv+wC2N8gE3TB5EZshhXk4oScxQgVQ
pTUbbTPeYeEkc4iEaljTwWj0Y3lyEYUOdHOI3/YWNyA2fVhWyeb92U1qvfXqyEaE
B8xvZ1/WkOXW1+NwJgIVzj0Qxir4zKxqvYBVKL5UyPhg608PUGzjwz3QsYL0Mnin
ZoB2H77d0N56UabB9emTu6fn7bwzUT/8VSK9DBZu3hanZzTejZMYpuKbYCrQe55W
wQGYizac7zBCkMV8Mt8bEMeTu+isJ0WI7/Us92rWh95Yu91fl/8PGOADiGAy5GKx
CHwa1tNTVVF6bXxNemvW1NhaKLeYSo/3ruBhO9H55Uqgo1gLMQA7Z2V4XbpDtton
nAfj07e1k00SkUanoDFEQOvw3dhZFaJ/sQLFP7QUczKlMG7w5OH0VHseKzNTyJPD
+ZYUaZ2U1E5z5cgRpKAxFAlDJypn1OuEU/UcDoC6kIx0TuPPGHf+GyqttiYLkyDd
4bNS4X3Hy2oSFNWdK8zwsp4wW6wbn5md/ZAKr5pltoUnlLM1PzIhns7/FBzVZTXD
4EPNEs4NMCuJRCNMbcnr+ZHQ+XxmyX6MRKoS5avTANoDTaJWtJn/YNmbDZJairrX
5oPpIjzmBinBC2D7Pkm7VVhiCGnM7PqqKUbII3i/EC0AQEzw2uo1v/Hu/LhMzNe7
K+7Z68Mwm8h86zp7/kH+FM5Tq3cuQcVb4f3C0Kx8zQOQRG3MVKNDV6A9PUzGeqQf
ql7po4C7F2eW23AFI8yIkg67k87/uaGK4d6ApZlF07WBGPZYy3E2SBT9FS1AUX7C
Llw95m9efEh+nJ3GCzmGmiAaBcBekOhcecIuVt4IKYAr32xtbetYmulPFQjxIH6O
q8P0/ATXehxRIqMxog2yvKovx4LDFcOR+0qwz4ijtpwGgD8YEW1iaPDnQNqVZWmp
Ljqbt6mgmqFDh8wZuvn4ngHLFQo1T5RLR9xhPRtQJ2r6YS2y4kl96uk7zJmaNhCZ
JtfxSjPJI+XQZ7J96DRLDO1sbt7x470ggtSgevuz7ss+UIjycEbBBbDc3uYDq7Xg
uv34bjLsEN5bEM2ynibHjGzT2zrgo2geOAwrCxD8eLiYytcIgmpJp5pCmv3NGRr2
xOexVNsGbOLfGEPrd2iINmsOug0+AVvknx+suteVmx0IHYm1lFDX2Lj0V8EUw4EI
1cJuw6uMwGPQ0/hghehtFrlHnedD7M4gTOUu3wIpthqqiNk7rJWnbCCmlabvI5OD
LVT4+v1dCz+FcPJ+c4ddyizLH0OUcEn3AB6UA7qnExcBzBlOC9xHtH2famw1U1pI
pMuwwnDbR34PNwf3mE0CyWUKrD0w/1ycunjiooKrJKGZMnc/MaM3DBPOWW4jdkG+
h8GUhvhVVGmS49jzmfLnbRMK2oB+DvUq1MkJ9elmKgV3e5OI8cPPWv2R7LSse3FM
CmgK0Zo6zBULtV1zdxrrbA4W70w5ajhiLh8ifdGPEq+NuUolW60xQgX2Xdo+lYdz
QygSlKDeJ7y0RuRfGFSFSrtRQR2OKmeQpZ4qPtI7lf/xbk4MHW7ZosaOkKoojdOP
0r9BeAs+GmnWUD3QxIgmqbZeFvRrgTehe+ZbaPpuY8flFzpB76n2jvNV53I2xQLc
NtDIQYb0gmNhfgJsR+vDlgsDweKuwGKo3oOHw9zGETkGzwgRpHWU/wJxB5oxOfUv
x6/NwmR8gLuJry8KO73sM2XHyjKMaMo4/c3495WORapJ6xu4+j/Q3H4MX2eBxNjB
DCpWMMFrDJmLamxvsoAyQDcOpioy+GcfuNRDlswB3BCICXfbdeuH5gtWX3gKKs9k
CGb4d9oQWabpzWxZxqNizkhs6QYfVEWLTM1dZ+yIBTZUSIZm6SYO/RshIgjBp2bM
oremuAui/Qwk+tekED+58yG+MoypSfhQ6nPMAghqz14uiEy7gXyLaIIckU7qq34Z
duCGXHhBk3LlNHPLg3Af+XD94jbiKweO65nx9ws++OzashV2Wlp7orH1JY+l3LIE
6lJr8mkQCXE+E+272H0pKGmJkb2HSQ3QXI9a0xLiAYgcn5bzx8ghIvExmrZlCE9p
oft5Vk9QQA6HsvTUqgrzDqLqZM77fLRpplMNC2bxl+w6PtOuYyPV9YDcAo2U2GKW
gXcF89A0WzLdb3rgE0UlEMESUDTalBxxh2o751J2rZvs3JQQEHB+gDGXyL/lJlKW
RNI6u/zlVopFqWjhdewTfKxyi/zvbWJoN+zJBRoXK3uS4aR4mOx7l4+D1FQJaK9D
JfQ2guSJhNZO2vp446ssdLn7PL2mOFFgHDiXzwdsxfs2FqaAKycZpbqdVS9N1XdN
aISGfdfwAXEN8JJNHsOPU7KkUPbJmW8onRcnT2liwOvbaEXEGikY7C31heMBdTWx
b+fK9vfMosR9I+g/3FP/7dy5EBEQiGWOyZVCEIRrwYITg152EBnoJ2QcYBMk64Jx
BOs/73K8fbYDNwwqXSb1ecaMz0hAsPiv/ckeYxJUa1bSMgdWg2F3mEu+scFMKLIC
Hkp4bNLCmBHwA5Z6h6DdGBbT6JVNCSZGPjQfmMFEA4WQDgcbMFsrIdtn36YIbF81
yvsM378cusO/pnRtJKIP+NJbL0RTx/wOAr3yNBd1p0r/dv8BJepBuegbCVi9Y8v0
xLhc1aSblmMSysGaG5Wbt4SUeUBfo8mTCrxxktHDiS1VkdKnsDbM7MDk/Zh1cSXm
91iQm5c0tom6ugIHl90j9GJoXxEuSy7aUYcb66cGryJawXLGAA2xDjIsxqHWtwub
ea4snOhuMzNDv1W9vHsuTG4uZ/rZifKsl7ncp9XO0zTCRuiap72D95XImORz7rI7
l7DxXamez2snc5bTxU3DAkcsxqjAmcn6ZB6ep4a5/LdvIYzR2OkWFE3Qi6Ay5/Uf
UlKDej8N62LfRFpkXDZEJyeU90tjLbX31vqFzzlid3dEv55A+1hSlTKIhLYmxMwO
T8cYWguK+V27ee7O6YcNzEmxWgHscEbWaMkLk8SqQJhdtsWuEeOI6+um0/zcMv1c
AMAiNYRkOOyvgc3q/AYgH2Er6PnaLTwWVjrspNZjltogNrLwu2oW90IItnK/x664
+Qs61CoHI9SR5dDCM9JrwkFRa58W6Bgo8lHqoSSZ1rdOyJrK50D0EKowmgzJrz0W
sRYl5idThV8tHZGojFHEbuAu4v4Loq8qR8mMVzGNUTKDpC8u4qZFy6GXknvluSp1
ajKmtUA3SEJdWp13/K2+UOb9CI9ya4L0ggQDehkQAEppKDGh2+XKLNMS+JT26MP+
fmzsd6h0l3BrvjZswHp9/ekVvO6AjtQP5XUZVthvujlyJ9h6jPfd8jwO+cWLkFqm
2xekt/6TGo1ZGbwIYkiKVjET1BckYqGPvEAwt17nRJ1/d7zoFrfVfjqTagnrdDEq
QIqOdVNeaxhywEUR2x9eA+TYzV7HTmEhs4Jv+FOrXqaKP5J2Z7Mel4GcRBcbtrfk
x3IjZE/N0WeEaclHZEszdBqDNjz1GKIcWirJDA5fgaE28xvMMnWM4uSrSA6N9VSA
+OnhdUqxEhB2nhViiK7kmsX07WlIjqHmYxyatrFJ45N4/EY90sFebwcfjYX1ep7w
urwC8STrdwyB/6SghR0TB0PwP15tnuvpGIglpLwwXQqO8Tgl3hbVwBLDAx6ZBa2M
WQ3T01K8OWsVk66+0Wk6Gm/8dWKVfSbs/pfX12v4a23fHpi6qd/AGj+UqoVRsvsd
34CpxH+UWTixQtIuu5BGmV9GeK2yB5QrA3mpE1LPgD8Jl8bROGKPn8J5qERIt6xk
iAJT4FnUvuGummIhLNcuNHPpTH3UqAYgLM1+Nn1RqoCVD29dXRCBtGJD09LuxoHu
+BpFu9YqGitQRlLruVVcproi286c6wr8rZkXpM02pJMKQ9iXTf8cyx41cX00kG6l
6g3d6h2rCQyUCQrSOVCuXQUZdytx5uhriJSIvwvDvHmlNmKbtCF21JMH4QwcLpWU
lF8mRGSoJMPqX5MhkAGykM5wPhXMvPeYRtl+M5msBKbJ06E3QdHINLJIFSVEP/Sb
dy0OFl5qedha2CauurIQ1TSkp3sIPS1yPIh47Y9Wh8K0Yp1+FthKacCkOgDRP/MR
1IaQGU2NcxKV6F/ukkizYBZp0lZCjNrSq2ZIrqt+dKGDj/+xD21fd3srkJ+qQDpO
xWWip/zeSJeppkvn9TsZNrLAkQvct1SBvbf1pGjmx8xvokWEOoKrOQeIQylXvCXC
lpaihM6cbClh9idTeDpncBeJUAEHHQWDdtvWJANFsusSIDs5eFyax1zGOxrnRstn
nLZaIyM7RWkme1mYM8hFGhhFBqFOkLRzrXNfIYuL5MUSCjEDrhhIN3s7d0K8PYd/
g3sbTJZ+4Gdy88sfq7thQGhyXOjds3GTwlIA/aMcJ2IEB8Vo9cFzo3PVEMWF6Ruc
/GuAl9cj4QjM++LscAvx5E2cAo/zYwPiBLdySUMC0F6Ispa5IWKk5KxOrSww/FHe
rlzv3YswW42v1mcVnhHSwOlivQIcZaVE3jSmd3BWnUV/ZZDubAA7etvZbi89LfRJ
jCmvYYEDQg54cdX6JrO9fQ6sEQpDgrUEIvLP2C9fnc0syrUSJyktXtf2cpXe7nZE
TXKn2SvkFxzFACCgn94JtA7nQMV5JVhA7ZQW0jW7kGvgWkhKtjjZUFmIWqaHtOlc
MqqToMm6nVog3k5mIJKa1sgGeawL9tsrrKR9CdT8RhX0XRVKGwVQ0H56hPA1k7X0
nUmTN3Jm4j7CIG9p6CCqcBR7/Ci0AY4YKXycj/5K6fiGcX34X0c6zjRQ3a+8T9kQ
iY3FHF/vwgLUoqhU6uFBu4XC+cbJvOZREcyUNG/o3d+oc1jOBj+Vd/xIE1m9BJyU
ydwyPqIqhJI1WmXZMkd3PAtO+K0OIZGSLCKe1kvTVUhXCgppEIx4fdsbF7iVQdpe
Eo56meUrT1nb/8pyzJZLiVj0R3rahMZYLeA0ZOBZ5DCibU+F+wR0iRRIdvdc6hL+
574o/We0YqogOkrBZTSRig==
`protect END_PROTECTED
