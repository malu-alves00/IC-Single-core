`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jjctx1J8YAqc8jRBEnhZPIgpEOdbDVjWes1rrn67x73daQso75QOBkwvtW9HyIMv
pE5cK1QzXf54UXpd7G8oiFFq3BOHn7KFnDEu9MIbuu8B13hVmo2dpS1PNWVA2/CW
Nw9nW8SVlZ+pZvg5V3I/Vtg3N21tJNrmXneUNwH7abybpowhIm0IjbEUVJZRQQSP
HdVg2O61TJDGwO0VibxvOLkDVnzwqi/hYLCRQKuWSpfTyva7ix+vG3iaMKPk02K/
3TlZ65lhkshraNoWek9WT4ECDetQrvLZ2b5qitsUAIuNWE75vBrPxTOIij4y+Uoq
gV2oLEAtqbk6yQQ6PF7quMcYCDB8EC7twAWdd6pa8urVZGTGw/2OxUqKN8I8wL5g
L9lMv0S/Z5asEXtUzAHyQWvLJ9cm33i7Ggdx9PEiJegu9hoHJjtsMMJ/PZqCA36G
JjJw22GnL+Sni34oxQc8XKdJS212BsOixFmSXLfJ/pNk3Pgx4mibAua4O4nWz3dQ
ZzS5TaeFz2k+UJGcbJ/xCgOvBe7xvsNwd/WR4VYqLD2tws3KFI23LsPQBcFpjZ2p
NNt4x+IyYXo+AiC5qi6DRATN97Z4wx/UgzShZBTywmCZYII5+99/v0bJ2mrCWux1
DSw2iOrbwwRuc3zFdBAkvqSBP4WYR04gsRJ+U0qJEDedPfnqzdLJ56UTNB+t3d95
xeYKRortm9Z/R1V5xqsKhyqubpI5FJPtr/vpFeKkdoQYjiAC1uYaMbwHvncmlO1M
ap3thpWRZ248h4RFBW1/ZRg32t0vcwISzN8eVA64uRZoumPpFMzhhyR9yDQnOxr0
WsFNOoLTV45ogAXJ61WT3FINCdwAprWrkRI5Xp+qInbFSulUdcATHb424qd2l8nP
642j28b54l/eh+5rqfDRAQEMoXQskMZa32mr+Kw45cdDxPJT6h12wDLQVaaeZyCQ
dd/5SFzlVoKm5JRqzfMXJYpSN8dhMq25E+Dc/q+RgVQaNejpQ0kAWYnKeMfs3OsB
kFfLjjIiPACuWT3oYr/YaodsBaKO29XBa6ZT36OoYCM=
`protect END_PROTECTED
