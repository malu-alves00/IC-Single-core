`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HgylzQ3+SgxXNxBiS5SauW0mKuqzMK9uogKIA57TUKFF5ui7Zb3ObnveQG/Edyn7
RN21RhKgNRAD5RunOeMpxd75NXcyqQ5mn37MyOCnMDhBeiaDigB0sY+h8oq74Tq7
H10F7Wo1vR+O5JAFE+BYPMdAkwpCQJcoq/llSjNgAuLvouXeMhbXKdvprvJxAIg2
Y6RVJCWae2PfEDvCTHFJ9H+dQ7tzovuPvosDP/JgAjG0P035zVrxYh1VjIxFeyzT
DCAS2JTgc+DY2/rYxTAZoynkWAq/f7HcPq6IkhuZZ4HSuI+4xLmobb7nKGoqMGzn
wzqrpMFrjh3AOCpkf7dNqpUYQI7i88ej1AKiJBdRKInGjzmhegvZ0Mhf45fxNrnJ
waOUfT5E1G5VhTPwNmH3GHc+tFuJEG0TpED6n/EZY1GJc0+ELbfoRReqqzmy+LP0
2IH1Ctzu7CKYwfzT5eNo5GZRxBDrK07yn3qG2hkfFOyhh4OCENfJPGWikwJmm/qG
m92L3FIn0zYGnqx3n2Fzg7DJtFsJPmmC2rWkfIkOUzUtWhoCcQQ6CEyj9M55rm/K
p763YB21zIO66yS0qeAce7RUlcdzOjLqS2i4NLW5o7UdCV1von3+eGgbmCFEFuRX
hcav7WoN9WpTNE7qIW5xpmmWbnbfsvE4EmcQoUMgmuLaGe4ApPmr/0ulBx9Eonbl
vVxqEl+fQoNHUqFvD9S3e5QqhzfVW4NV0w8+BPF2hs4e9kLX7a/xmP/T533HD5sq
huP9V3BQswVMqGXFzhvsdXbO1plDxNs4lOpGcz5mjF6R9Hw8DM5eIfyCWTXvkAkx
dVIpabWRwo7ozdECdY6vi8zNquXfYYWv80ruQR8WvMjl7zarHUD0z+lWexy2r0wN
31JF+UrmrJEVZDzOONtpRHBqEy+KgiqFqQKTqebr1Tg=
`protect END_PROTECTED
