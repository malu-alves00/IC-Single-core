`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Lg+PLiYycWD3QZzkru302q045UC/u/EiWwO1hDJucAh0115vshWIZSF/73F3YSHc
psP0yKeqtMTvL6mxpsILbWtPzZ3xBhX3KM+eNmYOwK8KeMTrbfOA+Iq1DQY9o+vN
y2ZliEtSw/pzsCYn/KKfirjNhpTgoEG6Zw9G+jdOX2oiranYN6LW0K3B+dJ2YZdS
NiJCKnbwhhzQeOXmUsxhnmsySTlUEE4W48WGQDRITuxEjcBXcs4eYSsFH/3vGKEx
mBFzDNEg17Lc311awnISowcHFn4i7TTQPPUYZGGNS0gDEvSuAIwBrElkKGm1aubB
QhhqM4sWwyvmTdqzzcV7yLVlz/sFJxayr6fYyzXNoGwBHx5rmCk4zqK0KFmPu1xU
Q+ZXBfcpTBcEpX87qlSjpPCw86U66mlyQDFaBsIdRUkl4OfFdD1j3/YccuHIxTmr
lRvMWN3wqiPH962RHBRc0P6Vxnf+UQxWkPbBn/tH5FRXAjSm2GF8hcBbbKH/OpC6
`protect END_PROTECTED
