`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WnFIrkiPubju0QgJ7xmF7emO7IsJbDlsWHs8PQZ7aa4vElJCUJ5HrFZtr2zKZtEn
Vvk8ti2i0T9hiX+Ud2uamBEMUFiQxGYHu1i8J79lN13tu0wAIrVYWiJV6gy9HDCt
gfHrA0+9xy1KEKA9AR1nsn6l+tQsKDBsD1Mg0xj3NMWm86+8MmoWaBI6ZdQ9gt6k
UrTnIgn7l1RmMglWRJDK+xR4rSocpXA80D+t0W9hHVmF+zIKZXEZx4v0C+lgKPsk
CotzRtGMutyvfM+kEir95aiWtEurQf7shcCFWF+fa692KKShyuN52orEMf3qE+mV
uuQFaxEBB4CXqPyk9YQ7r47Rn/VZmvwB/2yyOH+EN4WpvZ9dDSqOsCap3G4KbEAe
GIueiESZeF6bjG8diOluYA==
`protect END_PROTECTED
