`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kikBcdCpm2SjfCE8ibUfihTPBJKzyyAIuwk0cxaRrWdb3h6WacZ4uSnRsFfy2XVX
c+srfDX26tntUQKM0fbxqOgda2oZ1dLAQQL9+x7S6jw9WkkBncWzVzilik1fuY7V
rofTHXf6COIZ74BiyPb2r/A6e35jnLiBvRxrFdOMcj34yuPQOK1PC6AVpp24z9kb
IZfvzAQrmSqn6zeYuipfOaOc49ff8Ky/vTvF2QSZaj3ygFrAlsjhNInM6HW7TtyB
FX3DV/2+LuuOfn6SkBkVnEJfleLwLa16CiWg+sYq3sGrU3LHpnh/VviK1odVkEPM
hzlmEYQh/wjQI3PkY+cXW6+GnG6NKWOn3TBWe4AjhGP0aEqtfDp+0sdKSBzRpc4u
avEeMru6zU8ZwX+4MSsQaDxXsYLI2r5IAWMR8YayphaoXX+NXE8Tln2ATxqYNUC6
UDXS0FiSasOA/UqVtFrC+ygQkFhOnLJUJCBoNhJ6B6zMuPYJj4ajF2rYhxmcOL37
7Eq3jS7TX5ZluubGfHA7EihbksjVHHtpsMPmrK/dcRrxwZyKGRpsP87nHThVQYDz
J57SmlZkI8BVfeVzcOeGdLoug5QfCtk0Le4my5AHJi0c0Qs9zEPhYYLjY2F3qqXD
U+BLx9/s+FDwe8/yXaNfVrkG5XTU1FtDVpS0PENAOsWpyCa3BY+IPZDX1FsFW4gY
yFExruk/KbxqP2OQCKNPCkGu5Qk/eighL+8jzypZhC8RMNxqQU7Dwhk8w1/GL26/
gkU/p20VSHFTLI8nvge4EUg9lvHQRcMwBxVl341zvDzZgTiBsmkuL3C0IMEcFaQ/
oVEuZdS6cc6ABMt843dfFwY/u/gl1I/Qb3/upK04j17cvsDz4TprwkW56Hu9wSHP
VePXVf7QiDtn7bElkTRhMWoJxa1eCrp3xArz7UCCzMK7nRTJZf/ud7dujc7QSTrJ
LjCIvf0xFH+r5+zge6sDAaKc7Gu7EpxTuaWPXYr3VSB/IMrDoUpCgAw8KBhgK3wC
fg5QeHmyejFPn6/+u2a0KXprrL3RGVab6V0dl51GQGFFQy9AXjXkx3qkv15YcqaB
HC45paS12pmyyPD7pEd3d7kps0uIGiXUodLSQVKecmge8wWcbTkmNN6QaPA+tlR8
vyIlOeJFDVFxun6oRiZanywU0yL/lpDILfQyBz9boutTPSvgv0gXMbfjW60C4NmP
AZea70CWHC2yfcFegiLSX13hKZ9CbKnlESmBMfz41VbItx1B77Q8k/RfhaaT6aHC
OS8lioVXd5Y3D1iuMQux/i+Sn7jNpI4XHaGVjWifOD8PKFfX5MDoj98uNkTwOI4O
dt5jRGoWnKYqzJUYsi8cAPJDlpe7qfg2Nm8UDd8Frx52WFpsHh9ye6MHZhUdOcQg
3ztngyVdVuVOYXmxwXddc7cV5jVwXvT4q8c+T5PvTqVCt9eT+exSg/AaLkGkGe9M
zHI9YGZ4bCtZ6Ku6nJA/TY8+/atvbt/KLSME0OnGEDwB7HMIKa8cYi+h+NspP0ry
yGs6hlzoWY9059caCynaKnhySw9tREqLVHUoHSKctyTDLTJzXZ94GH/ntBl6CAV1
hSj7Fk4Hmj7VSb7L7ul9wW4nN6w7gqVykJFsXZMXYq0a1QQFb7eq2BKGvbfZ80dO
`protect END_PROTECTED
