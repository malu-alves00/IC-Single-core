`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OBxMd2sqjvlj+oiUOl7U9xzF5AisQ4AHqH5gVp9JXVsP1bDgND9jP44AemWtW/lC
qtXLRLVs+Ri5e2T+MftO/PzKQBiJFDMv0iZNtmEANUXZmZdy2nwhvMlAfIwyySgQ
vFfaMP/RTrh+Zwv+us+yT/HGCm9WEnla9hY3XIGMY/TJnSWNP4GWpRvvDMHq7fMC
yOt43EreP6X6ldHocDUFhsjC73H8HOf0Ql90/iNJgXRD1LVSzaM/Fr9TIZByshMa
85p7W1INjnY4V7Zgm6ErCnMlVs0EhYlTrcR4tZogAXSEfVuX3dS+fdrdyeLIo0U7
dpR8J1fbxMz99iMTpEIPPgpSA933v9GJWdXNFI81bohFM815bNAViwRTLCGn8Nlk
KGcJwo9hfwBtsoDuuD/0TSBoOD+PxgtL3ucT+Jr4qd1yfSAjQl7icno/Q8RS0JNk
HOn8N6sQi5+v/HHwue/a78aHltCRpyvcc48FW9fw+oc=
`protect END_PROTECTED
