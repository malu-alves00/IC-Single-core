`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
P998aqwTx8IRZzUHCTy1rJIp+ZMb7siqPmpklgvvl8m7wQhg8XokzbLvofG7eeod
y9gYe97IKpGRYWSpLQB/3GsGXcvM2CXtTr0iDf/BXyF2ScxVvFsU2oiJ3BVx1rVt
HbMGxa30ljQBH2A2uxMMPPFMlWRMWC+q/v+VSBLxMZM2DUM5G7rILkPnuHJVKlI6
/GHSmnVqUQT8CJuFrSlyLHgPDulClz/DGUZNFIgNaDO9HbumiTP189OmVcZYH+JD
GSlv8Ze05rSq15LDaTfrmF0Z3OTmq+ch5go13u93FLoHTy71GIfEH61UzIURUA0e
TazQSBEFV8bXyN7R3EDBwdYkbKceuXWeQ1TS6txTdxLb7HBq19eUWvwLtaZLbSVM
hhf9oBLwvh7bF+Ts6EllG4Uw+V3dSKjbZaqeVWLIfxrUUcolNie3Xblp5XXJmoOg
T0N3DvJX60euOuF9LbQAsJy2zbPdzt9M4gxMUzl3UEzrBr6gAGcxF0iax/0W4FqD
7VXbMKFN/z5A+VP4cbbL61PS2KUyuZ49Trv3yRmYQfb90GQvtvTknjkHQ88CePx3
hJe7W+Rfww1WqVdktiekuZFTszaaewjzF9hIrCsnOKF/nGo6x0QjeJJJFIs8d8KQ
pWsNxLj6XPeJLwoiGvD6y63tcSUbiOjmIDRYNZK1/g1X20S35NsXOtke4JfOrrjy
IXVyUW7MTvm9VNWjhoNcAcLRij4G5/C94FkzXE3JtTPm7YhTF2kTRIRS52Vy/I9b
mr8C2O6dbF6Qzgozxb0Z6JPUDHLE95k6bKxVDNh0Kc0P22J06s6EC3PD+agUnCuL
/XLIZDYdeGabnacljjzpevjxdG2grc9uc5m931pzCmc/3qoBlLlayDLR3cNPK+P8
1qnhxSamoJVsaRlLJ3U4QS4qfYUtXSv11tMzKkrMPXHMa1EsVXslRz1ll8lsRiPA
TvPBwDR69pDfd3yijJwzYgG8qnw08xAV5mDLtBisXCqpmFJtHD1nIoP4eRq6wrHa
WokfLM1g8FVAO07chvRJarMho59SLzs00MIUsIAl9+eEUJajg81iHLDOYx3rtmQ9
71F/I5XJoB/SzXQyx7qLbrfS9T6UNXCodz+oNKiHzH0Cv208yDuHWYBL7TxgB3fQ
uP/NIIzTxJ6N+FCNAFCZxmIMpUuO2VNq0xqewOA/r5s31m4AwxoexqKDwJBGRe9n
IAfcu9JIycUIK6Z6cVibffwUGzl32eWv1j6Y5ceY5LhNcp2TE9cw0qkN+vBPQOln
9vpelU3opU2uJ1k96RuFks2lrHtt/k5XagBTuchI6BSySW9doAmpPvWs/JFfWAu+
5g/HFMTR7MF5azqyeAgTOOgtJIC6gCFTI0IcZ8uU5EjglYKtZLsa/tMHplbkGPgZ
q6TIdR7x4epRTBkz91JPCGKlw8rz3VFHNYepIkaGEJbw0jDJrEddRyYETX79pfDl
W/F3cksomN60eV4yYEcmZFw0zAi3ab4UEd+K9TNYm8NIPCCgNsuowsUQaGJXJfL6
uVG8hlFGQr9qTAIc3Y1c8olOKYoCjRu/ZMpYSQeKs+7BFyxXABE1hIScu+7umC51
8PwxnuzRC8+Sbp0cyjRz7qUbBYl+bK7XJjR+N2mvpARDht1v9EFl9juMKs2W3a5c
cOo4c7P2bc+IbjcXSZ5S+wYGlG1p72atFKQtu2inoqwEK8JgRj2hIUaZKEMiCVTE
U4e3MSv57nW0YCbXjK65PNwsEdH6OHSSEdEaAP53vuKVQQ8rRr6FYARcdgo8WHWB
CQF+sh/lJp7uPcMpaqU9/Nvep9FlIIuMoq2gHgOeu2xnvyikuQ55vmVPcF/WCQ/2
nUsaWSxM1D1euCcLBpKIki5XsN+6cJCWI6ip4TT5uinaMnzfXczP1M511N5LrUf+
oA4ZDwfnYnfddcwfvn1oJdZNDAAK9II7WIJYhpWu8WE7EA43Hf+7KqD6rJ1t0Qb3
gLeH7JLA8zTkjULjPaVnVDqw9RNug1UzBZ7IZTSnXKvNjxIqnHEAEyaLh/E7McF5
zkM0sVmEaSP9BQAAE+pKg6CblExV5LOA8L37eDBghqcWz2TUxaQumKxw5TXtx5nR
kKzTeVkKrLnLH8aI64R3bOLcjkZ80/4uhqwxYj3ORHXtos79n9C0ZEB8xYODqWSa
rNxvwo5OwmN/ewo+JQv/t5rpDoZIfUD1YPcFSn034Kv3MUg0gcHXPr7ptqLubzjJ
T+LsEalou86xFY/F/U55zOPvJzJgAaP4V5bszQQ4AzalYJpsPHtM6hCUQXlrF4pe
svNPQFcPXn0AHzN62/UvUFPijhPis/o2i9mTpJrcWL/0qjfjaNlefgF5InGyxYRN
Xi8hML+vKFO6hj9bdBLS4EDPCSAqhX7WXHpR1AlR/U24lyPlpxQy1i4GZJpFtXrE
2/POo9KkJYJVqnQHchW8vkaNP6UsQHJ8uQ+mCW7E84g=
`protect END_PROTECTED
