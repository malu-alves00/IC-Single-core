`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UB8Hh8HpZtqP/pu8z+LDWkExhD6xJ6mklh4yldkxAZgutOhvu73XHeyktW5Wm0jP
xJxDBQ0zRlZmbWm+jP9iKD0Ygb6lPd4L6pN/i4tcv1RXz81KKVJTkVvYdLPxvdm0
5iIv0rlVgEsF0SCGhwM45sJb5ZRRb6KOoI+Lo+mStqthjYMbDL9obF0AuQibTUgA
Mh/KR74hcT4Vt2kFGgr2fu1/RLm5qievqy+u/ICI7i/ORhx3Naj9kmq/Usx4lkaa
bqYs7kDQkb1UJ+zDgqQbD+JTc28dwA548p0NxqWHNl+0heLRKbCMbnyBkvR/fkZc
cccUc/R8E9vdGqCjVN2hY3fktGUsi84x9Z4JURuj3VK4lF1XuwBA5ac4uGOfvYFH
ILT2ad5Q5JdmDD7nVMf1mDwe44QlfvqE/sVOEVRTxXcPtONc0eEz+Shf8H0riAJI
9RwcaVu95at/OOY2CBGFJS5tHAZhBjnnBtXMh9qlxb4CiwaphpQCA+cPByDG86Hp
qFILuLqAhUAY6k5tcwEk+SmoaLvEf6Gcmnwz14F4xeGSe8ocY4qwHISb2rqj1hoU
fopW49s9TglU9LjvmmVsfDY+7pwwjGmJaq1OdzgqbDUJsS5W6xrijszrZg9v9EGm
ci26OVFPOhx/SOpGOAHt0VzhnqrySBnU79qHHqow0B8X0lA2mstpxM7KbJCniyTA
5X3YBZ5wohBimJuU9xsKgq6Jly9m4j+MWcVHBGjUbtCvroMe/eL82eeMI20ImR5O
EUhMHFHXljvllPu9/VWcyYWUmp08EytKg70K9waLp7N1NU6sCDylzAAxcMtV802T
`protect END_PROTECTED
