`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NTsKzcdcqrIBYM0AJ59xVBzEzd/N6t83LVzpiT0KAP6ici6XZsEAYmT7ttdAzFfK
JSILGzk9HpcN8V9zqHjOqm5HaS9NhzE3kcCAolbT7BK6SRdT336lvk+aSZabsoZY
0pPrExp2fzNiCymppcQRh9jUgbtvDMsSHVCmCF4CpaNY2zfO1Tx3MWl3SStf68H8
vP46DkmUS4JR9f8eaQhbM7he3x9JLS2/99KPA/UULG8xxMOoa+og/nG2Lo+fhlnB
hCysJP1XvCs1ffmDewihECH3Djkop08knnVgs3RJEZmlrICyc/1CHbZsHa1rqgdh
ia8zvD7KIbKXZRSB5kiWD542BDJoph4BmS5A6qzZ8N3qR0MfgYwyP/4rAPvaqh3j
1xXCt+rPGZX5X8qBzgGTfA+SlT7yTOS7EEEIimfkdjcHdmG0B95pmAY1zbIgNySG
1Q+Au2AdWDeagWqIuCkpa+3w37zHoJhaCDNON0yaoMC7oA0kmDHts9phglZ6yT1S
8G/keId6bdBlYSHrkoclT+/P9/r1Tdl/e6EoffqQQHHrBbwHntlL97f1uJS9CiMh
ikd7piUpVdJF99wL7MLypu/ip2AY5J9irKBSWJh/J9p7VqaQQCMOTpudqQ0QJ7rW
uFQDJSqnwakfk2fOdnt/vY/JZY/92t+0I5w2IYKYe9PEBCW3mcUtJ9tnieiT+3t0
8J+yW3yGrIoNaAC6DvvTnYZGLrtVbIP37MjAvDlM4tFAzyeaXEG+c1/PL8LW5+WN
dD4n/fH0thPjgjzMOSkj6U7V/EI6IwFP4tya28J2pp1LeX8Hvl+AIyjd68N5+z7M
NY6Dhx4uW9HD0PiLs6tU5V/CLAsiy3+65+mwZof6bfgCz5+Rl/1yNyYp4pfwC7Ou
8F+xmfolQYekMJem+gCWQqmQHHiXVNrOR48xboM33maynFbPvogVZLxnbTbUhIK8
kSYP/fnkhpP4V7kZkuPjqT77THHB7rMZuwbs0vSzNDviFCAsN0uNe/VKDaXzE/Hh
XK7XG3W7xWuGK6ginFORhLpZw9DVcSLTnSpGagZZ38kPE/VupAH2c8ExE5fPlfZj
YD5+BYY8pJ8ej1Gmj+LLi6+cNUTOvMhGSht8wwo7PUzo90jIIN/Tauj8EisNn1py
N2XtPorZ6xSmP1uzdzNARTLHWKQK6v5I9ew88AEn1WVMnq0hCnrZUQO93tYIrb8b
P2N3rcBrgev4bPgQ451ix7hhPDCON0mDSsSByyNa9Rxq/y502DIWcNMGqWtPDboS
eiR2S7KEli5+Rn7IQ/7XHLB1gXqsNJgPxXImIahV+eGmx2CnRVtrULw7MSoQVMze
ubg2ZtDVF6RMAgiLn75Oy4uflm8KJm/Zb7+LDR/KZDV8NMogfm2ZMhJBXMUbsyyL
JRctmD6EDUFEJJ4/MZWYr7fLazW8eIdrzkaXOHRBDx4MRQxGUQCjrW+7l7U5zeZo
tu9sXKfSa8GTozMFHugZK/2XaVzlirddb+usnRGl4+Upcu9xtAchHVja4wkfl6tp
0gZhrZOnIXxPDz6u9NjR7zgLbjQMUYEwWxGShJfWibNr8FlUUEtoyNRuLU9aaYXi
59Hgz7qJq6Vz5OAr7NNOBMP9wpdAU+qKpJf7iRuZn5MKzvHWU6nRoJfaCyrBQcCp
ij9BJdLTOM/bAZyKxYz+7l6PlG13taQtoTdn341V51i8vqm1GLF16s0v7RUa3uSa
sq8YUr7INTmGmiYc8xgBs8/Zxg/f+/stySM8Y35FGrGmTjCsc7Jw4DfXr+R20eVH
milbIq4XUbzjsebHJQLPgVF4dcWMzlX0HIAXm+YAG+ARCK9qPXtMYJEzz059gg8z
2BhZgtGk9sG4BN1OL/HH32JbsoMEQI4jvR53AHdRyqeJ4nnKN5bAss7gh3G7tjYJ
kaUisavp9g7m2tfc5uv+71VSqYppcGvi2rjxB/xcBSUj97HbB/EQw9DzE8tTY+Ig
bDZBUaLiQErNSrWNHa82Jh681i+YVqGzY2+EX3aC6TFmilzqkoc4doH70boXQjBZ
0JDtpSfGrGDxrNc7p6WEtCgZe6j/tiuQWzuXDeNRvOwvxmUiSJwHmcQOJ0QtcpO7
rx/3eBVvJ9kPWx6unlzYmxsw1XjxSljP8reTV+XFhuOwHy9fcAwbueS9vDkumIKl
mOSSdikHicj+i5K8cAZX8cqjZ23JP6xvAh/OdHPxgaUVD/2zFGKx5w6jZvV7F/Hx
fzDCzFoD1DVrpJDoKaeIvzg/aearmDg13acGJucicVFbE6qoaz6XA+bMiZUbl6SQ
ln9lHH5VpDi3HK1lA9P3me1wEAGNcBrhUk/cgSGRxyyp/feNliimML0uPs5Nr/t3
tn6bt0qxrg2BaBj0Z6byjbby3YPLOGXNVRFlWEFoUNDoP7wmgFNMWxETaIkhFgCp
4kOar8Us/2bFdQ5T+0e5/RrN9ffIXxqAia08P7n7PUjdrGPnm5wnsxSupS3N7qs+
Bqmb00IpTPDoCLz/tR9N+eLyRKm9GYwqgPkcrQQJY2G8JdfFHzb1rzPONGoEzRj0
mMiHDV7qXWr7GYS9oDZYymut2aJvauVGvEnV+dts18N/zkGjUbyIQbiv8x/mYJIw
4s3aUhIzX9Brys7rh9w3fe7ojYbf9Lqo9A/Loi2jCr2cEhw5mUlvvG3TBRsyL1xn
tXRszGKbo1vtxBUDwJme/eC41LPEk1XoQKWSrf5i+bKmgaplbFdFhgQpDSyPwY0G
WakY7uJnYBqv8e9z0AajHdABLqG4P7ixODA6jLT2iZSZp2VLEtqoUZ6n1rDts28I
fUFJa+lpXV8jxHcj9R3wL4spYbHOJ2AeTIeRqiQZVAgCoBi7u+MnPkHVjmLT7b4j
UnMnCGVdKzxqUpqtX6Yi30fV2kKOpMbBbEzWeP6pHMjzEY3HP2GZkski0lnI6O5F
q6W9AsteuE5hvWYrxK01lE7o3+znftdpKkOqLdAYpwgIgy/JnKeFMcWqB82w3ZWV
XItn5joOope7a6JycqFhJHTFEIfsutovuhDIf8Od5AFQK+HET3yU4dqj5SZCHTPh
QZQXmNgIIUP8hf37cfjB4c9TqJDjTBRT7gwtYzb9ShmGRu4ANgPsKRJ2AIe5bAjd
QFCeJEyO4Jpn8nwslVOV5E3xmENjZmBKxl0e/pbta6bZu6jvtFvP0aUe2ChEAKsq
bmS0qD4Zd3HQpx9TNeR6Zw4jOGMY6LoYirmEd7rNPtahZo1YbvUkmgwJ489vI3nJ
wyJ1/02iUIVZuBUeC6IOxZVX/YPu4I3NsSmu4tw3D4eocwsMzYwpj6sUDw+5Swey
7K2KbbrxwapLGxvZhj/yEw==
`protect END_PROTECTED
