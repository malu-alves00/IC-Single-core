`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MwtHuyR3TPhB9/AUgCoRAO6tRxUMX6SF5cc6aHFx5gMM3NAa6st33Ck6XGaOoqfp
dgXODKQeZNPDZzFPNMzpF3jIbJUbYaVF1F7bKL19ltMuhz8kLyHB2X4oYict6L1B
vcfHhQ99DclkXJfQj7xodto6petbQXHUiWV5tK0SUf0Ig23RzhPVcPB2p2ndSVEF
qEUA5Ge2g3J2OB3/4AwLOnu/5bxuvnKZy68hHjmoEU2RiMg69BPQdk5HRWfhjiqA
9+ldpY4L/ub+SC33in7p21uvGKmy6KUFexRU52gnUvMw25hJi5X6aOrRrpa5RK1s
giqByF+p9Ps8D3IlUoHIlgfXVZYbzpEHT9ukB9WECvcV7F7IFJizuCB7d0Zfw5g3
JsDDfONs7toxDkvC9hY1PAbKFRxVVBGCmJsJhnTLndrvUgj8AOnprtuqVjKzdxj8
uoPXYudhH65ml98O6YaFCKtT0c79rDAyrq1LMafagg4/Y3jtM48udSws2bWIaYbZ
qLe2kfIawTjPAJwZh61AqQi2iCr6BQB4qAwUZ1Z6hiO2lBmVvXpRk9vU8GdnCWcS
wNs9CtfPLINymi3vTAZ3ng5ihCh3q8A4TCPkdpQ67ZQHe8VAT0F/am5Wd5AwtLOf
K/Srpcc8FVDHyCNRsQ5qiRpSMpmwvT5CbAWgEppCodKoZct+zYee22w0TtJQho9v
o6ld+q6HoQ8h6WMwdR9NLWGkw5V7Wk8nrsW2lqw6RhdDlaM0kMlg7XhA3UPBmNMy
c0K4n/JZ3s7VmIBMUXb2J8eYabwPf9f1yxa6CGb0VgOANhcwHXixhzv82pDMbGxu
6+mRFdl3rRG7hifrncc3IJnSFQBpkXpSU26crKtt/92fFmKcYEYgBTAGOeVfVpcV
Srr49iCXd3LEaf//3abatbSZRgOVbG8mLf7kCmnU6D1rhutN6Bf4ngsNltVoKkw6
hlSe6oswgIVkUIBycoo+HhQTfVQPFDrYtPjgh4U5Bk5FKjTJgAfPH3oRuVE229Tw
zp9LwtnHgdmDZiSxeNGS6vW6Dw4V+IecE+n+YHOus3SWRPxxPB1hiFg1nrR61Prj
FpaKuI0ET22fX435fUU5OPQziJy3RzdWu9y2EBE9cqMVmV+3l6I6J1m2WukiwglO
tsW3jp5zIr2yCKhAPF5GTfN2eoVyq8gw5+rgDJSHLiI+rxNdtA7DyLrHk0/1WRIU
NpHWwK4u2IsQUTOyHJvVP4YOEF+NiviSRYY+wjuOIviMEpkXo0T270hWwbOa0XWc
n/oLI+FB99yF49m5IG579XM31Xyue5TrGa1vVE0NH8b6k/fn4mMpZe9hUFj6EThx
YZOcP9bOi5+a4+VjOmpNwW1oaLfVEPTCPufpVMtyrVxSWfeuVJCZcRcA+Vt6WtDl
iL0T/RANHSchMUdJFltZBMbrkCVbjTb2p9EKjnK0sTflodsspGALoZRqr37oe8d7
b5Q4ScQijtPcQrvyPbz5xEEifpG7QLkKnTloGgPCNZZWPjUS20o2YkX6+x7U7k8y
WbUErGiTl87q8TIFBcobo/tthSaDWkmlhsZHERmgebxrYWoeQ53ESSx3ylBdSWdc
bc1mzeYjwRvB1mN03IpFXXSUkyZ0L+tiu9fn/C+dBEKUBCquLEpbSNXY4MjwpXZI
FfbnKWi2XpuLY83RVqevc/rE6WZwBosRAVvq1s76BUiCjLcI4GaarQXK7+g9qMm4
KeeTMRVDVuuKXkF1qTreKtA+25+Y8y0T4TiVYHzbDMnkyZGiYg1dLLVUlj6FCReY
D1cS9KwWwY/wmDg3+VJIDTpWFCVFSZcooNg6+DTcTPtUExCQcbJGMN/kVfNE9vo+
I8hZ44GAURUgQHIrWG7eF4B0etSbkNdwsIBka7I7sV7snK6wRC1PyVuXbSrLN/aS
NzPyc9VZg+lg96gmmrAPdoS2HZ+d5ZPjs3rciKaaqvIIAGWXlOussWtT4Azo7Hm0
dGvhbZAVKRBOj5fgfgRGlFpC1yVjMaRXzzmdV0c5UdiZqRgo2Pf0YFzb0jaLZscr
cec6akE9kvxZyMjpnGV0zPJl2LsybJx/s6fDLr7B/Kpdyr7KXrqGMiLlCLiAPMP9
ZS7rMRvVm94NLnzSPzjBk+qd5gia9e+k5ngDtwiDUK2oaiBGUYGnA022YQf9lbz/
JqzdQ4o4Jjmd/fw7AkWdZkYYxpglSt8l9kAJ0b5/URqQdmOuvkftUKPcvxQQ/uQx
dPUV5VdGzK0y8EdvOROvBdfztCLZ9/7sHDv5YEBUyqssZePF7FnSQk0QavJvCqUU
+1CnedcxggLsgeywV/yabuxdb6VLYhhlKtNeRGrq4aOrL+1ZEaMwftbqffIDuYAh
+yoa8tQwOQKdSGQASddQN5uMxt4QFt+9EOyHR7e82r2NtVfaq2zPvTrKQ1SC6QPp
VCeOu4Z/EeOCmbCK6zy+xOjDSaBvMXCE5u0dPvODy6JDVmS6d5yPdk6m8dYdXIIl
ESjZwqhBGpXACH0wTNSpQ2G0tCxMyNeVLRsMr4foS9rJLMqLtGcbbsGonxr8oG4B
i9msN4/QNCjf0pC2SZdWDWvpsOzvDHhvf+msCZXKJv2DXxNaDjmzvl1Y+Q1xWFE7
lunOdugCQscTvb0uLgYNviMUcTU5k9mi1LysFsHpih/eAcU9bWDGoTPZJ/OLFWQl
K67OU3hef4BJ/A56K3PrKdRbxC+PmA2kNof4kZfaT7nuiNpSTVRQATD2gsy8r7f1
X9si4ETPtKLIicYXbzOA7JHdDpQgcElNHTmmXYKsboj3uuwtGwjX1gi3dVA+gQDD
H0QfArpcNNmOEY08S8FaNB3GBRasuBwOWwTE9GaC9bqWkJleER06RgH3g5FvqYxe
spV8rXfBiALZORK61RMboj3DOcO0/ChHFUnIf2xvV+5lT7+rM8FxZZliPDpA37wL
CnGkpMTPvgyNAFMgbjNdOr955STWki4V0D+zIGbj+YEo/QldWLrB9WGGPLR5LuOX
mE0Mh6VmrHtgBbyHDhXJMLLz1d7WuEYICmyTlCgT9/NqmKPImGfvFF1vBU1Iif7l
OvlFrk7331D5zQuvS5YC/eWS2TftmmWpauJ7MawtUMWK+2Nv/x0Jg8eeNnaSJ2lC
4lFvj4q5KTUCURhRy2inYTdR5D7ovHtperLMiaz2duIuBQR333Nxs/ArWujcZKfQ
b655f8nwphmz2SKyobAwelVAfFAT1RsVl1dWHWzHWC3j8RffYnmvud7GXNTe/6lF
xZ/j1KZdudIZz5whnuTIrjVQnx3A9X4SIhoo90slA90QrtYTaU5Ifgr0naM/l/s7
1Yp3igkfQu/wJPRUNHmfAY3YF4lGxCcMfjtdVbObxZs4DK4UIfm8sXbzwFnosidY
/iSjtJCqiJc31hCzpN3S9HeASk7Fwkph+JDZZjc91VPZOgTFKmj+WpQwc679Ev12
aJY4Wdo8zYpY5WdybE/eAmJljK2StJU1qBS1Bq3/M3O9O/DUhSZltbEAuWovDTwM
qpgDlkh0b8+/pyInyAFEa3uW7i9o9Rb0fVbBABMUaOMCSXI+++6BVzjV98Nna+BO
D9rHPuAMH1u8q8MDqLngROkbgR8/lOm/VyJKB/yIfUFw+KfPBr0if8/UFc5D1Yan
qBLknmu2FNQlwlJg3+qig2ZVLP/0etCOIuIIYeq4+D8qfaYE0Meeer95eN/VMFif
jfSZ7NACBhxOhpyES31d4NcWbd2BpKYYUZE58JhlPMjTI9KzjebY2DMIIfkZCD4b
hv681YVZhcC820Oldmu8I9s/PjEKpmIzVQxAX3YMmJ9h0a1MLNthu4d3GaXFmZOc
3O2ldi8Zo/I9Y02xdN2m5FPuv3G313jtlMgzjw8XbyTv77zyxBPB3DUg03aUWD0V
TmJ8TcVeDcFZzUHtxX4okxGjEfR1RNQShxIRGv7qyrVmAP2D9IkPvRuFoQzrA1ZC
xC2UoJeEy2Le2je4Qubj041VRCsDJLWfbMyFKB9oA+zIxsHbSGPh5hGNbO+AyIA+
Hzr7k6iK7k3+7h9iAvJczItnvF3FeICaTUi9zyPT2qQm/nFR7moRZXoUvvePFvYB
FkN+k8wgsProcfYiHR7YTP60n68h3/BS1v/X0esFloLW4abpLAtJlVd/v71rUY+E
DDxgWmAcR2B5CPjlc4oC5RYv5dqtdS0wsfbRGfyechA4Vi/pVCbq20Z1xCS3jspV
koK6JlvTq9Scnz55kuoz+EKKoeAkg4j+wcr/fxjE9VKCXNxqXJRZ+QKvHNYFgfPm
EsuevW06cBVn4GWPAnRoMtGGgAgnZdrxBWAeX0x11rBZQ6ZHvwlU7uElZAKga1Dk
fBIyp5XjrP0+wuwkDKWICmLU7quMzPOULhDJoV74ywwl+gtTeKQcjxhcvpoVw/25
DbCOJZYeFAdO0O3kBed0NmDwB9DmjEXf8jPyMiUt5PctmTKG8z5P/p3cJaNmryyg
bxu9hbzlPlrURA85IHswAguN8Z3IGjD16TXlHz13HBdMlGbfSIrg0ALJpA1nI91X
CouJmUImZ/qI9R2O6Q+IxJzLw0rtF+OBUVYcTAGB7FmPK/H2ewS6SK/UprXDc7Ap
g+8wdCmj4r6bAEcALTrvf9azAJQKwsjiwJWmxBilAn+3nFOROnZ2yhtTbYZ3P676
hjFEHWATWRb4bekJs9n/0ll/GxwPyOzA4YotcqzwjJkUZ0ECy8kqqI4FmzRAzoXm
kdPw29G6ms/0q1Tzyb8RLrrARevXAyRlC+UzLIfHwqmoidT+xd9PGIhcI4GdgS+0
vDdHlNQBcvcaxJfZ4eb6g5OfOseUp/WD08B/uiAfo6Uo+ZiR2yXdpGN06qE3jxsg
C48t8pNi6US/PcsDBfQPaW0PFcqE6V28ZVLmGg0VX0osRNauEUkvrF5bEhYpJPUt
KmeAeh6jlk7fBFTqsQ4EcOatXFCkWU+Aa4wS8zLgQ4nxSkpldOpItZldHzFz9J6v
+BZSti5o+nhSWdF8nlTJy3/KCE5am2oBbr6sTZdQzokTm3g5nO1cUa3a6QKI1m9j
AS4rczvQ+eZkIYvLiUeUUg2SFMDXvZnvjjpOW3iSIoA9AH1DMQZBnIk8XkHx/A2K
F7wdKd/PzFwkxiFRqtFFEpRlZpIEqJdp/s8JzM7No4m68janHxT0ptEKZPOGRos2
2zBl7HnBHuP7E2kX257QuhmhUD1rR0wsrljDjgMJikGvDL8ZPk12unAcfYWcZ5Dh
+iI2Owc889S5k5T5m53G5n8+gRQMUqR1+RVIPJQlToWwOD5zdFvgxi2LdOYJudiu
xa4Ik6t8rP/OVnjME9D9eSqTIy+9oAxtKEHwIkMZYzrrqHX0aEG4Gw3iqqPBCaMK
n6dyxoV23spV1J+Ak4aZvFBbuwrtUVwG9HhEYA2Gf92ygnSEukZiE6cN5tfCJcla
4uqgyH4IRcm3FtbD2LLMsA5izM20XVARV3Q6IDeNUnDzIpL0/GeacXZMOvfph+Rp
uuQo5xJ+WmKli3CPDNIr0E98lPmAYH+Ub/JwrLjEAw6Hm718GRR+wKcycjZhVU/5
UrzCEmDIW6S2qxIex/q6bYoiW0vNAkK+CVMgZVderLmKUAKXfKSA5+8mZzjaHPgS
FHzA6zvzOsLvWINUeEvcHMT4lkvbmeHIK2/kqegtCIIlXNOKRg4lSDquw0OQMP65
7+cyjQk/p4Gk0TagTvMnigUDkkrIZmDubGb7wvHOHRD9cS/YGLNxlVCvNFlV2PVf
5inC5tIiroMVdS3YDhYURXDa/mZH5l626V/3Mr3hqZgG5vF9N8ANL821dNsZU3Vh
1+1Tsyj8Iwv60cnW9q54mXoQh5cEXSWT8nXTV/4PpvPGHt1dR3rxO/sEo4ni/uDV
tBduKBWrS8EjWJGd7t0VY5c3o7/N55EcIMcutkWMlNbKU1+NHpVCEU9qAIYhpRZ3
sNjpikkPO5vCsH9S1XyrMfcwU2ZwCTgq3fCzps1MSUx3W6Qf/16d5BkZaS0YFawX
FwS+OVrieCsyhMbN9ugol2UHcoYl4+BWR6A+qAJFDQDurEPxUsNxUXlAL+TNnC0Y
f1gcNW+6NI+dSemaQ6/oBSG3O4WLY0bSMj4BYekulV3R3LVxEyoLf/ENzbM/YsHk
noWtdaDQyoOtCfcpXb0U6T1u/EJTrjkt6rziyzQngappPX0UPoMU1NoJACC2aQ+U
HIXJ8R5Lxdpn08sABuzXTPCoJHqjf3R7s8szffebSbYYOY3XxYREPfQiqpK22Lwq
hw4rkIV4UxmRWLQBMjaImUAFwPnFtRzb/+A5ylWDd2ehixybI2kE6MUMFAj3mQVM
Olc2Wim98u5jhnEhOj5Qt4McwtviAxnlG+4QRvLTU+SIDrt86R/aQo3zj1r+H+xU
+BTNno5CbbnKTZS9rGn2K3oM3TgtF9a+fPhFhGD6c5/10nZLVCxZb7Rk46YRWYOz
bLfLE3iCwnHegiZivO0St8AL722iGJrXUe6cTOxCSXJD9i9VO5aDqKatZq7ih2L9
E4Ofxu1Wcifl5Htc8kv3mcJVYPnCI9AK5uE+UeRQwvRlJ1Xr4rWJajKOzwQGlyUH
ru04J/xyBDDtIMBjt7cQiXGOGwP9IooADpzTzLtk/rcVJorsYlaLwJ0H/S7b7ACE
nMCCfgrICOIrSswwV1ol0T3Qx/FFRHjaWoIA3axRWYvr242M9ZSf/19XXfesSIR7
IZUWDV4kMZX6JiNw1a1zcptt8lhGkRjs7oluP9D0EPadPDyL4CkdLo40+EuFI2mh
7POHLaWTiWIUnAOhVRJ7//um01Y92qPZrqwbTIOYpuLsxcpLDWtw8GzLDkfWWFCj
+G8DE4O4NZjFVK0azTd83De9Rdz+1LO0ueasVYQEgQAWJzEbYP9jJYbLFt+Cdunz
QCejbFNsNUg5oCubfflGD6wNNQQtXTtHECAeI5hrIMD8Anw53kJDsdceH7sIV1Tn
uUIvd00i0izqAn5Mb3ZKG099HPXqWfI89SioKghzfFolmJfRAzsNh+cLSJ9WAxhs
f7HEnYf1W9H4g1ufr/zr1bhn4km8zHfwApyEbH5hDgKdDrhp1wppR4H9cv2qLoMd
4pu8YyHLeJgEEN5d0hyVToLU4nQ0ezod54dXEx1xEDZXrT7AQUCLsbYtMRft4z1/
z9fqT/0Cj3cOGkm+c1SvAsoF1pIIockC8j2F+ONW44Dz2KNjglO4bDqHZj1BbOAG
F/kBxkrWu474JrgE2Pu2zR/spe4pi6AeyNOAe9PInQ68d7b7lQ2+EMi66IXXz/tx
nhnfSO8vIFIU0Vcw+hY0496dBMRlvGlLOOPWkAavp3hQVjWiNu9qVEJ8MjNh//y2
zKjBqzN/+Se1UHC0RQswCR9BMFNbG9Nu+pp6yV/V74mQm6XwwPcoE/UMqvVAo2/h
xCHuJB9xmZV8J9jlBMfi2jTRq9U6Ue2INgWF91IDy/ktS8s16Jf1BQLpUuE5/RWp
cnw79j0WtWAba9PBNq/jLzw8zrPv/AV2ndAxyuZ8C+CAatG4uArERk/3zsrOnuvz
9YZg9wKCNJITarHEQEu9fPchzaQkIBZTt9DNmLOS9o0LPGiVGIJz4i/BJWPwGICR
cdD9zUh0i2J3iTijjvjgp18jI/TiCa9G4NtZwQ6INBPMPfbnmgzLAkiAMy0ADu0U
Kpw2oSumu/NqXeEDVu4h5HuquSBsfO6P/mpKww3pLP8/BVzSy0K9bD6WnFkohGMw
dr/rRw/7ZJr2AYEJOeVS1ncVvNcZr7TdIxU8l4NV1NrvOTjfweAR/il5ObD3sPL0
C8GjE2WpfKgZ310r3cQ7buONJmxCZBHTHtI+doDiYMh+k54u5Tt5fH4MGmIb6x2A
+B70r/My78arS5syncxpQnBPgLo8xH5YYu36Qo5X3OjTmuBjAIdxba+yqEvKnlDG
DGeeOhmrAI62pLPyRCQ3ZSQxwiz4iDkmj903bXbR6AId/TyZcBsiNWqIyKSHkuDN
Ey3+aM1ofj5NImBW3uCshhDuNWxxZCZCqRApsXXTxD26d9m0IBPEPypnhMToDq+h
f2n38nL5DdWZxckevmGM8ifqzicXXuObAefi7fwAhLEvVba1SDfqAdE0mOijyy08
gaiSuRvPRX/AN1ZLxWO1hsEyouM2ckTsOclXpp7dBW8KXnBaD+tLFuTbSyI5DAak
uT2Es8Y5SeRNZKdLNMfGgqKS9txjm/tpWYPmaIyDsMIAAvPssoPBM8BgOaWUyDW/
748wk8eRAKg5B26H5hzTP/bikpbynANlUvVnTKJf3IY2GY+jTDwccHs1U6XRcX8K
tZ7xI2MQPwC31oYZ24d10/ZwguHxMApZyRy/LDrOtxNwzMs2FgoIGov7B0AKvCG3
JOasKjWjRV6mqSwLWEJlK4f6eQhMA1CAGVzjr8qb0TsfIZb6YVSr9kmZgAtHOdzm
IfBARMwbCq6qnRxhRQaDOD9rv1MttP2+e+EqIDF0Q68d3vXYKDMuJXzpn1yjp+Ly
8izPoiGtg2AowNPAIx3IZXw5kN4HvP+KZDnlzkw9AjM2gSZCTq+IgBWwrVRN6WGG
L3ZeyghvY0ozdbbS2E/+JMZKUJ83iXfakQ2FxLFXoc18uQPIaCuR8u4IpOmLyLEo
e+q6qHOe82ZvoVBjKoqCcRxdpLI3jL/m6kAqasYv7NK8zc0iBPmwGb9+OPMyGoay
Rlb906PgMGVEcDexWtNxwvRheLfWu7v6viHcI+EmCDut5TsjaZJYGarSQmVpHFxz
tdQbTzcwbxRTj0oL4Tw5nrhQLuGIJhJ1FU+o/yafNpSsGYHtwbJDhfeZD9BJ42HH
PIz0k1Q8DMMuyikWW31oIWTaGD7DvIVeH4+yWLFNVGtW9VcxVlQfuokhiUz5+Jxk
//sYA6wx/bK34/UMM6UvNsHlFfpIH/faLYDChSC6kd5vGNbYNZAfBTl4EPDR1jZn
l5JEVijV1o7rZrNWwr9Uglj2zOeRg9lPdwf0Glw3QKs/YgmwyR5dPJI88izyvAdP
bN3+g+d1a1xLiXm9yWFNAoWr/5r+QucVzMefGj4zjSlveCnfJJFMdJ4GBGvUx4CE
5jF/cdwRoz1IJOoX8875R2tAz8HtUpaOR7YCkNpaJd3nEJb0ZYhWTezchHLFkdY/
TJgDPWaYXNQAKeDonfL6mqygKRhiATUTtKedje8gvcMxeIvO6rWfyhffzWeiNxTC
T4RmXIf6o2sYwGTgCH99zV7JNf7eanMIt/gqm+Ol3xDY/sCpetJWrtHFlE9V9RaY
jyBGzZrOPPzOW4zF3NkpXQ1QuWmqD8PPbUIal5mgUnO2lmj5dCI9LInj4Qtgjjkc
wCQSrankJOCYdyRaSgkMy/9nuezZhHcYAu2QTMDk/lqGEpf0eeHPDpQOAjJgFzpz
lZm8uMD9jjo7Y4fN6xj0lEGS1P0utgQfsTlqg2Tr9Op7ql6bxZIvXsKQL1+iX6Pm
ai5mOcAVRQRkIT4MtbglWnnjesfWTtZD4Jkvl/1W+Ob3aHu+A/Hb4gdK8/yjU62l
pMMLfiOqwRfcWFnIMbpnhUuyXlQ1AF2sm1lEJe8oFmRM6lacxKpbonYovJIUX2fI
WvKRm8NJJ5GCI2rv1wDTGyhGz9drtMxd3a4ph79xFA7T3h0UQevNAaGfUwds7TlI
MAjfK+WrMpQ6R/1dW8lgyEdASJ+DyUCFICGU0dcFzSOjBEqJopWFVUWQfgYmwYJH
RMMFoWY9KI60MDIeUM5fP5zOBHn8pLYsctoTbneI1EOCPXHvsarbyF7ymjNTl1jM
0pNAiOfKGX5gbN47E3cUfDNKQ638FqbjMP6/Uwkoz/UOD5/Xz313uuRJxatxlS7D
7scZ94J4/AxYOoeGs0fTD3X3XUP2HioZrM6m8RgaE+Ljtf6ip6beU+EL8KuxdhME
a8lMDuvlmHT5uccYu/DrojqoZNXuPwjf3xRlbduRTRrjKfcdDomf1mAkMYXGmFpP
pcWTCK33MhPV+p7vxAACQyNb9PWUmBl05Xd471SplVA0IbtelFDAtcL2mbUF1KW7
dAO5Z9GiVjgQw19fnf5OVv+Iqk2iySKPXpK3YXyjzBR0IynskYwjgpVZKpjfm6C/
r7xdCv4M9kjLT2oec1HytvDu95SyA07HRdWxQ9hpL7czVzgezcSWCc20+VqG/mSt
miycWy5fmfKy+ifuOvBdZ3CjHSQDQIAHBFvlOXusTTvuWcgX+gkXvaXxLvNsCUeJ
5W8nKDW7KfkeuqwMeDHjYS3aUSLr5y93TSQhuG4Jre6dYIVIuhHg3COw3qO4SHVM
9HoMkCW4uEqyWWAJgulkSVfvTmoiEf5Un4s6A8ADcjW5L4yX0q/C5r2AHVOBmBTD
Q/ZXXKGSvpXnlqfvRzEPb1uGm0bVZ77yfmhXWpR1dBznY4DybTQZu2IEtGBE9JZO
hcEQDlGa7LSaIblNeO2icJFJzSFF5vfQC9U+O6o1OxDZg3HbYDQC1LdIfaHkxR/5
Cis8Uv6wRqieNmkrm7fRIW1wvtkxvZHp5dTzEuxS9HUJUTQLf0JeqEgFHQROq8Wk
zhm8PfSNqXQNytKlEwdP/z66I1uT3plh2ksgDk1QwQOkKqG6gvgsozq9BnJNicwY
EJfAxPFAhOy8ifZZ7I1OLIAlc+3IMQpUp/6ZSM9mOk06CAVe93YoV1Vc6N8OLsKZ
sFA+dUXlDQiatm7Sd/hL5273I3G4pIX31aUABEK1RK9IzPXj/dgYH8ExLIqcHE+r
qF3Ry302E9eDer/ga9yRuAZE9kgqJwePAhQyrNy9PdJqYPZ65z/Qw3OmpBAgw2tF
FwpNBKBRPZHO8DxPuRkXW7SiD2jpmRPCQuGPdR6aDWxPze5MASzFwuxVszH+5P/Z
HZ4j2+ymjQM0I9gLG73lrcIQ0WAs5GHhFzsLWwEEmE5EqtNsuNIx0C5jgPQLiOyw
P0QTtzVBke9vYLkr1YHZjhSU/A51ZJp48eW6JUS/06AV7A0xfRhBFm/YvdGE9ZSL
BgS+y5cOBNd1jgdCOkSVQXgAKvm/p7gZFIbBRhjw9EMA6rFILacJPo4ksNIFJcV7
bUsTUlcDq8gC6Pz1dSNQu3d0UBMtyFDUQu17aN/LMpwOcCfsLUtSgfQbSzuBGyHH
hPjjImNvrz794GxSt7Um9TsP74mYZVwqXIF1UdkI/j8oI28kTuWkSW1DWqMSFWhf
0qzwnZU8Fgcc/CRbbDz0RlykvgU0ETZvd+MTy94g/PCCLBsmGAio1OU5BUFmzbhn
jMdW+cY3CzuQP2/kvx4lGojJzWjuV4gPC1DnqzUBIn8A3cMI+EzF7KXcoxmKBSuv
klSX2dOeDlKBX0rqXnr90pt1WW2Rq25pwHfjHGVjdLxrV+cK7lPH/veHhkbkwCcp
ACLimEHzv78mavkdES1XkNYjC/guzYZbEYiIOvRBs1eJk1UB28A8Nlipphf14oMl
n+L4ap7fRKgU4bEyyZ97PTNAmsDsLQWLlNnVAIAvK22o/y8eEac3/+mkosICsGTw
bpjXTHRGkv0ruo2iK2AahA9dvmEXO6r/YJFs2qMaFF/THvoSVg+dZVrMi4LsSzlJ
tWpuSdgnoNK/O5aZ416W8P7BG9sOGII5rnj02q1QKCZOnPlH9HiBAvt4Xzzj4i5M
NWWrrHZPgHYbGQmmrNr3WIPHtfIKu1T0KORXAzUZ+5MPcNMhb66oDNdLLPRfjOUv
NyFlJr3YdyZr/aL+5GJJU3ztIG0egS6woQDLiZkXQFRIW8PMLKYB3WhKTkY1cW3w
1Qi25xZVoRlgVpAPucy2seCPkx+qJsRgyxj/pwGGLvIdkQ2ckepfy/R/+STvz+vR
xky5gJPDQmKgQgwNp6oYVXOfHZJW9RC/cKqTK8lTVuPT43O1WymZYKa7JjsCisKD
yI969aUMUwzetbNa1nH5upL0/3/waZFpC6zW59Kn5YBlkqmISD99++y6R32/rZ8V
D+DJs65dneRY9UpzcfqAsM6Ja8dLEzZp7HxJdB7s3WPCeP5pquybKI5fKOBDKa2G
QAxAvX5h+TUO0U/6ZtSfZy5droD7Suih8wFCcgF3W2Cf1MRT729r3xAdsWb1TUEZ
7uQ/f2HyjQGP9ymzRClNmXIMAH6Z2dXVatKhVN7POI7Lbw2PqYbyBGZE/JLdvr4v
R8mQF2fz0yLLuhlFMN+ySzQRaG3ECNjv1JzRseBg+GNPtTi8C9el/Y0FxshZgy2J
Y9pSerc4uOoG+m4m0aQiKKJkDa6+aWYxjGp+/QrANvvNedRNC5w3ObB/rqaXCWK8
iwv2vffvUmgqrdlMdkufr8oKZtVydeYhAk8bqA0A2y33s+SYLKsa8mMKPt+Zoayh
EWrNNpkNMNVo9/UGTV1oq1CsNlTxaDJkm0cqeAZYjEgob5g94MXtZ8v8V+gUHWyw
dzd5Pr7iyZdLSUqJ1Ibuf836zqHbie/GwinIYKHHKgH/uQJYOgSxe+suCJ7mTJOp
56kYLbPaiFnPSRkxG77E/rsjNcxNOiqGaFNswgcP4KbgXspCfJu9zDr+7qOh2BCC
i/F+yAWeQg/eoUdaBBuRJNwSnLKgCez0qf9xoRMPd5bRBH8wJOgJgHWGfBzDk+Pj
J+OIeF533qiUerGpVzV1loKCyueLCoMM++4Sz/22O3U56H7hkvwkC7RJD6avi+nQ
SLmthJZVvTdRzqFAT+Cz5+Mii7dSwHTIvv7hNWtkIyR/mKsleixfi6Fw4dkof5BV
V/VgIDUrneP8aJ2SyOvfAOhiMLt4Smcd5UIebuLX17TVcGX6oRQ9uW7XbkDnL6pz
j3/lloZSt1Qj7A6hRBvvvNuEQY4I2KHidosoQjsm2lHFSxHkyxp5QQ14KABZQokN
sNFV0dzHrFenEtl6mBXfU749rwQr/qO1nBF6yaO983X1mE7DB4tDJSP8zHpkflpO
Tqo+j/BTv6Xhnoemek/9TFvkNyl+sCTgOuEFCRrPOe8x0blk9nO0OizQstKFAl5Y
9kBqp7GtxHvzGNnp7u3n74Wmwi9pbPUiFK8kaaFgpvTG+jC9aYqrDE/mosPKD7eG
i1sZwF6bZ7P9A37K7YNPTcYc4ZjVlHy5Y90jMkajAmuF7RAWLVYb6JSieiefx3xD
qNww+2oMdj7poxCnKctCmZ2u+zw5QTm/QHDJuSy2U+KGWl25d3/OVWtRLoa0yfy2
M1Fg1dk3pITXZZ2NcXXM/0QRaJEsAg/az1pDKZDZGV+oIaJTIs4OLqxgGY/pkIRB
G29zlX7fSAowWv/qhZh6fNh2WMOj9FWlOKtilTsiixOWr40kf/JTLfN3lzVrDiyc
XO6SNEP0ZPIROaYb8AK9d7gGsvytHS/3rWKcIOvODibvSgrjFdihSg+KPav7+qLx
NJuk66woHEp26w1L19opAdSrOEcfA2kb99MZdWeJR52atS4KZtykw8A1oBQ7/LHM
jUh4EvX81TrBwoH/MxHJ5C1O8b5XkHE0bCamA8Ouknuvt7Z9dw0E+S8pZRP4xT4r
nK47KSLZiPJlPvUv6IWGOnZp2gA9SeUT3MqmYYIMxPEjuHE/e0EF5H5oD1xxb9S9
fqMjn+aHzlCzj5c+Ilh0m+TZrbPtd5zGHhLhkYEUwgOC8KYZYgwaQfGZx5IssyCL
JapTkOcmqL9BphS33nCJ6a/+YudVjyY90dNdA+Z5W9M5YD5X/e2aonEDd0CP25ks
Ynbg1TtMe4AkaPZdeZAYsZUkTb59ec68l4JtMInIohHNawyibntdpXncpF3lCF4b
3FCLUe9B8M/wpjXk5GvtQNdnnNAM/b/KCg5ZrtmlzCsSzwPcUpHTRI7Ez0XjQdFB
zozbwVBKLoEzEnX/wYqGwkhH4kFg5qJpQWYsW1c5YYodDbpIykG1VipJ61RE5mRT
rkCb3Htx547H5IBFDrG5Zpwp7PlpOvm9t50O9h0+C0uAHpLK9+qv68OIuaNNrmQj
fFB5oTIoo5pM754qGIV/ojzsEheZ36o5wICSE11Kq2tboWvdZlWiZn7ZwjOxafLF
70tAQfBj50tsEtS78Ck2jYm7Q++DVKbaiSzYj8ufpeS3rJgracumiRnCtTPDgk9Z
hZWmfpaWHlH4s02Lji8Bni+8k4wJuhc5t8HHEqjyJoOb/XcV5IEGSZdp5evdE/sx
qH7iciz9fJ5RqRw2I11tTPfZ4FHs0FOR+zjCfjKyBOqnNXpCDgbv7jaMT2CW8Uqu
vfK39kCvY/7Daz3uYNWv8fTVguw5ngzchEwAuCkV1MHpxOU9M+WzJnR3UsJEygI5
ZTNn4CyK/rg8XTz1awvbjZOQ1mQFTiZgYQ0LYy31lQPoYSX8vXaREE4HcCMK1qc+
pODFZ36tPtvNUIak2GtfkDZRGhH3+g7/jAlctL+iHcC/Zp2DDOQSkyLDHshKXfuB
7omYht6vMIhlBjXhhAAe4X/IyWZCCUk+iESikTYEqFmLUNSoYpzsqdwHuTq97h1I
52+9ptbq/NAWlYTS7A3AqPte6pX+ADqJ1BuAY3bxj9GO0Vf8wsTosBWuES2YUmGq
e2nhLduamvMX9/FKlj+W271uOGmBpcL2jDhc+l7rZMKaYGApGDIcGBDhe6FuIC9C
Fnw9YhNSgnadVx2IaLgV9e0TLDY71gd0po6dLZYc0CYehxgPjx9VOHIFNCSY+xJC
6HrHHG47Tz7aBomR29llcXm75Qvl8srqFOyA0KlxQ0qpbvgADX9vwetHUFnTHrDG
dUHz7hDbVGNzCsH46AftXESyogPopRogi9wOm5qlXmgwcSj7Eb/08ASYIciTJFIb
3XGaHBlpIqX70N6Tk+g7owq4ADEtO+C99V3Ra8hUlZX68m8qrdc7udoPEUBRPzEN
HxMpG7EWtKHib4iF7XdA4KWELTWdIN0Kb2Zktubp7dPnrX1Ipin630GoBlPhnIv/
dCX4MaiqITOAe6NyInjFJZQ39x4FVfIJiS7ZhU7Dl1EpHmRUuODWsYt21b9QCRBl
EL82QOrnz2gcNoxUqyz0PMVfg6lVDr+W5u9Dyzd1YPusu/lhY5FMw0CI6ZupJASJ
qUzoc+xi1LxW9udmUoODFISljoFMFKxFewmUDEqa83OQLbQMgGu/aba/FMv4zNOf
SzSXK7gOoCC+R18dyuAGPUoeY+vSOcM5exV0P5knJRzUQgiSad2cxUQZS8xUr30f
HXdR/RMhtA/iUYL5FLN5tgb/TdfMR7i/Y1nzQJLUMlAiuuyLG9OgIT/R2oAZTXPY
sFHsgx9spoGryIq0waFh/tZt4Twmo+pWfdE5NqQSnTgVAHyc1/aqEFCbBcB4kO3D
tbVJKGDYqlub2l0qY1Lnr7BO6I9DPMtwYM0X6SozOwIVsxW6LLvmbgLX+iIF/mk1
BqM3iTMcW2a9nj5EV1qSOvvGrBoHnYeg8k1gfxuSb25JeYJ0MjArOjjGkFgoESgo
IjzTmerlUBJxc9pabcCmYRQtnC0+SHSwEcRrjy5KiS4WOziid5pWpf2IneqCvuuW
jdc8b2+7EOZoousT6egL49tSYkFo/NnHTChpOt2DHiM6vDg95+trApaCJPMrhm+l
LJ8KppiTYIVPVVJ2CX3vRofmW1S21D1Zd3s+DWiEAJH/UsJsZgqB3Rd/pZmAoMYG
cLDPjJd75rUAff7R7c804Zo6QqdSQD7EtuKoy2l75IKjeugXC+DlLqEvy3o30wHx
YKkcK4D+8ehzKoiVyNHJRHAT0Or8ew67MVjXcazXqw097lVjh1lmQUwD8V71vOly
1NSZyT4mjL9vRkyfvxKM+I+pwqixUdACAHIhj/QQjJde7SWeaaErHk7/kAOymbbr
w9tREfgys1/IhAqiWF2IquJuoOsU3QP6tQlIjzHSP7AwqHLfPpzxi7mnNhQ5ksSI
wemTS5SCqWq+YWpzo/uqUhjRoZwGXdkz4cwQsUtU7cXuXRB4OHHuxg8weVarsgm7
6QLy+lAKYbqXdKFuaHLVwLtnnKlRcLyOquknmMOihwBnbN2WQC/c0S8AmcDpkFkI
8/77wUeRsXIHKyEDYUUh4epoez5ksCpFqfdk072Crjcbw1Cop5sOUlsdHazTihnJ
KbVEFBKIe+UYI34EMA/fnJFb9McSnFeQp925szU8dU8pLRR3unq5IkHG1SQ0nXqu
TnXFSul7qF0/1vQs0shZV/6TyJUTa0aheEz9vrXb+pdF8xhV1ayEkHJBenAwKyeX
4SWdnZYMSPlZm4Z/vb3QRq8rZNYKfS99GPHzK06Pk/ZB6Jtn/SlHNWTyU6gbRaHA
kPBwGxltNEPHwqZzrHjPY+e63mlF5g6pEJU6J2UwZjKSQw68qqf4vLH9080mwYGv
zKwOGlQFffizqxFN+6NZVyh6T59TlIkbJCyhd6qswBHHQTwB5+jPxtd/8DtkUYrw
THOcXraE/lxlAZq4P0zUMhakZhtTQRFGUY5q3AXNW/ZTtBRuWMk+qhOPSy2hXhrY
hLN1a448Avx5DrJ5Uf+EoNV8ERa504I+NNUbghelg0nBorsg+xXUF2g5tGJYHc5D
gzlISbn6dlNXQMRCBZLzw2i2GJafE1kv7Au6kzFYuBLE4jTuQ3DvY1w4AfquWFwa
Sm7c9GaTC5Cdhbd/a2IMk79vUPF6sIDgbM3uhU19JinA8eUFfsb4uYEmCFrdsmvf
X/ItF2s2BARxVoKc7IB1EfgNoA6tq8Ee8wxrLFDjwLRMd9JeSEWdgkkjx2NAJnOM
oQRS+qMSOWegGHOHkcqZAWlOumr9KAJ5rp2ts5Eq+ZP/h92JNBn7E0pgK94i1aU/
p5jU1YqaCW5M3PocAXK+GbpjiaPnowJJ4hSMf9hM9DsmPCdY2gl/YJjXs+EY5R+L
0ILFRUqFNEJ4hHpstNyOCEyNR8/yqS4/Gmk8GxCU4MUSa1SDiadmwIC/ontNpFke
SmclgfH8pibpdsUaDtm0JqpPPJQ6oUdrSmNMxCn6Zi8nxOT0ZmoxoBjDPJGZhVbB
un1jp964iQOcnw+1zkC3aRKDNwEIKgwAVlRexDjex+t9C/A7KOfHeXyzaUan4MpN
6+iMdCmobB20pC7z4VQ9wmsd16q3HWTQAVNPykbj3fLmlO5jrQSCAdJBriEvXl4/
Rndr5ej6Nlb7HlUvmz/exPSnCv6GJQclw/sbxY4p8oiBDdCN8F8A9AR/7LkLXWop
8Ac7nWRGncZZ9UgyyKOg2KlmL7E/SwfemvSl+nK/MiW5QAP+yFeP8BH95Al0tdtd
K227OY4yHbBHHQ9+8hIxzXAyfscb9Gg7sHVx7Xy6LIIrDPqSYOOq56xgtNln9cgZ
fnYMOg1Wcu88sJTXZww/xKMwAM++zdVA6qA1e9cEdx2/1hnG35FHdpkKGWALAp5X
M9EQZtilHllnjtQ2VtzH7qOrjF9SOFmWghnSmaNR6/w1vsUyRn2gPhciakPoTNT+
qNMFeVa6mxtQ5YSF0eP/ChTcLj76OHGLnFfOwWN3NLa/ooS7pwycqGI0+oEv9tAT
WFRl/xMmEIOtIfvXHTZKn5m0QosKj7mzsc94pRxkzMFqPKyjTeYaLOcWEr6Ywfez
9/VulX/FcqEyFQW2SwsU408dDzucNDYf39qe4KKe0te7OhmowRmLi4jhPyosCLbI
JJXOYUGySLqwIVXVGVdJs60CVbam3dR4mcnGxKpbh3Aq4OCA4aBLRiT4V/3EzIjl
sZ6NwFIl2HmBqUHEIgL+eEsW0AinSDmJM3ztyexJuxWW5T/AyqWb6VUI5YE0qqCC
63F9oLuIX43ON0g3e39XNulA3b1f5YD/gGXDhAXOUCAh9aJxkh9tTozqAWqjXfVs
bMXewF9Orvekw1lItvQ14HzGmKb3wpBKYvoa40tUuwbwyTcvk/cGWxGvIVsmxDAE
LpHHMuzCmaCzmrwFMOCpNFsEcahQAAcS1qjZFFo+rzH2EJXVK4A4jb9/BRUVYK7Z
zkzMQ3IPPEbQiJ8jriCIglMczhqbI+dUeSWTmrlNfuZ5l+xOZnMwN1TnV922gq+2
tz1V3Dhty1RaoEQekGDfFeoFUkkvPCEBgv3nTkyCGWp4T0GUYbl542YIMUdGzmoA
+wIE2vu9GJKfTwe4DO8dJjfiMZ8dkmUzw/22F79gjjx6cIo5pU1fAJx+ra1T9AsV
kcP6fqtTVBqI352BJEFVpJeAV8p3ZDOqKTwX4a32YOOSohlHYBkwqdipU69KKfcu
gYP7lmVBDj7zsZ9v76rOVrWWODv0nsWoIqfgNg8xQbQp/x1DtSJ9quvk4yH/o3Ko
dlZpyugxUOfbzgOdgHNJwqeSiS4g0Db/oEbp6/BPE96zwibw6n1aiNFMZe6bkpVP
f2l7JWbD+icmC8xd0ryYE1lRrGAXYaV5hZKql8Zc0vfgREm2RP00yPhmGycN+gK6
DddxwdwlrPVGKyGUUQWIuX6SaNPNHHtxFu97eJrgw/glkynQ9+HhHZs1uukzWZDb
uqxNeyFd6qVL7VUOjMahIz+RklPllWiNrB6AJxcS2ZV5m84InHstnQf7HjwbZT+E
9CkYRr3LscJR1t+5zbnw/gFxRYIfLeMniEq/ZF1kl+tG523MQAAoVRzK+AEnU1xY
n5sZQAbz6Jm2hXUFJubgs7xic0fUIGsFabsM44aVaJKDjE1DrP83q/bL2UnF2/to
xgAgTQWBZkBEBHX76fKaPvfzQcJSi0hxmdaocGYhrdGoVgVMbVjY3xLuwmqOmnsD
uzCXGW1SNPfWFs8OA/NazLmliwvsIlWrtK5bjwjKDTpt8/ISXTfi/Wcc+RK2XO/f
QOdxrjQ2S1Aeghw6BscnPaHgaKaEs/4SR2eV2KSQCft2EMZGygROIe8T76cNKRLG
3rJfY3gChPCtmtltK842aiTJvgYS1blfGvCfcgkcMNqCoSgSyfSnnTIr/WV9eUE8
YVM1quWEGAcuw24FZ9YPgdJten5QRIiEBQYV27PbAXfE0n+vs3yLAj+S47yJLzZD
9mFYu5myS19J0uX/Ohcde4gCxToMJlsHRlVhgnA3KpAk+KlKb6+dqrboREHrpFtl
xID0+iX+Fz9qWELcorYc4LJkvygkBeu67AR/fTG/KnSPrjwudoNidRiLoltrHObA
z19asqGvT04OViId3+cnKd5oDcIlTz3/GEu7RFPnbuam3r/gy8dHrPWf2ZM3xGwM
UCh4TiD/fCXBdxIVWnBfMsT3C+JqzOdsNWsNw1KI2YDskuCNKUmGnWF6mtONIkd+
2kEWfSvPtECI6r2SISU6zYGNBpquZ+pMkywMpIDYm/jis5zD53+hcRDqEz9I9TzG
qWm78GusS9M8/t7FtRsKe9JkD4XdSwaCIoAzFajsAPq6Hh70PXiuXGdp0tyKLKLL
iqsE6bes6wiHY30SJVmNn2yfZyRC0cIEm27RJrImMpkBcP2hH8otkcOCuDYSsZas
1xCS+vsAacjsfP+HyHYyddqqSOot3KuMCGQImvbr2/2g/wsEv1fnOJkiaNiatHdO
fQvlvj9rFHrxhU9aDTPgTXVCEzS/pF16UzWDy1/YEdRnyRWsq3XuLRXCu6ML1BkL
zvsaLI7ssMuylDIABHCYuvc2GnPqqZ7V0Tw4VPcovHOQulSmEK8dw8tDseimszCX
ts8/6XovfQUg8qU/RCOy6OD2BU98J3cnaUN5wYixjmOZ1b4BRFIDevDFpx4Zt6/E
cuIrw2JkHJbEb6uCBv32TodNimsJAvGB4tq0QCgH1nta77kLeL7wHkQQ3B9kon3X
KRaxyA4Cx1+3Vqt8DJndgsL5ImAChGCAsq4y72o1oy8qUg6Bu4gYAaiuq+vyjRee
nFjkSU9Xb2OOZturJ7T9jVGYoPk6zZKMyWR/rIu4DeN/ql0/RSSkXnRluBzV0hcl
PeFtmP/ACjJesd/DqJ9DeHM5p+ykLS4+FPs1nT64INOgZjDEnaryEgYy5zvBrKH3
8VU6ogYOEloqEzjMGThLGiN37gDZ8JE4J5t+9iEmsd8EN2z4FvK/d6rPDgigD9Ix
SX5K8rqE0YZ8s47oe3Fan/BegTBPvr3NwktvMhHgV5Dy8kmAxksfrHIsW5BEYlsR
FeVy7VsOCJlPyUKT6j8IFHkTGRUT7yeevXkgrQYrTHqFpZwzNG11M/YDwHae8+UT
or+rmhMjDEi049MDoHVlj+CW9nVN8QCSpJ3UMLGUKXHSt0YwTCKlycu5VIFl0jV8
VD5/hbMh7mK0XORrFmcbozLKTckuNyD6sUnQD1lS/7kCqs77ScnQSurl3H3grpQG
tc22jkrLSnzlvjtP/cXllZ4OlN87o8f5uaPRm99OkmfEHONfEzF0rriKef4u0Ezh
28Yk4doPKfHEGNwWuAVGR5UPbkydpgCNPhZ7jDc1YStnk3YD2g3AJnMGoZjQD08W
LSLWQPnxz6PX+CKhDvGiu2iVhTNS9u833I43S8qe/gxa0bn2Moqytmh4h9n4k/SB
xzYGiDQotFbKyWX24IbUTjPXboaf24sS9ugnabL2jREJMpsQRj60r5CyF2SYLbuT
KIAo8X9/430Tt2o5/sNWWzL1SuBklpvLx8T4oJbc/rYL0u+t/KeTHX1qhdZ+zvGf
ssJJ9Yv8GGIMht9WvrJhycEEbp6OKnLZy3oDcLq2OpZrhLU23q4Fz/s5KHcgqs5i
pB53jAy3KBFq1XyNJ0iU3LPMq4VSZ7YWxai9PwhUDstrEz9xdl17q4m7TjmZhhl6
blArzNj8bB/2ijI+WFMAhbYaIrHBWw/9XZ2EG7VrA7LC0yC59Ixg5ZG6gZlnkHk/
PcNF/R2lLIqV1li+TXcz3ZKqnd/byq3Vn48DZEZ2K+6RxiTOX1BZqNGd0LIGbmBl
sn7qiPyqE3G2bDriTJufUvqYx6MFttCURe50Y5Dt/I6v3PkUjZnLLHX3TNL+gSwV
9tpymsRqoU7pF0+L0ODvCBIXbatQ1rFqaI1nMTrLT/vYKCy3hJn8KMOQofptcvA1
eE813ImonKfM6IsHGTiOCMTAwHO16CcULEu/GxICsDuLj5xNRrb+6cp5O27qP4cZ
yvEpDWQk2dL5QoayVubvLJDlsZ30XDzzRM39bmkHdAhouH0u8q9ZeQ20Tpw89vXx
Xv2J7R2lEU/9fBPDSz+96wNBWgPs6t/AdWit5xTPB5f3cv/mAfiDCb0Bsz4kxiAm
RhQ563rifrdII5dcBzMKAha2FQD+aj0vAWPtliV1woI06PymB1RmsdtZrwttYEbH
g6Qk+9yyVXyh0Nnl0FkB8ZVeq5neWXvHbeXR/9+PagvVpG0Ozh5vQIF6qF7FS204
V5ZqqpAJhtFBEw+iv8tcPpwiRjlu4CAW6EfgzXJKdroGrleGolNy03znsRtvEpGK
nDcE9MsLG4G/FICp1QW6ivrUWuPjlJFY6oajMO1YlOI4ePXdijHuMjM+UsBIgnPT
uEMVfVERV1+aijMc28DeDC+W86qb8LKzhjp0Omj+oz9QJMgQH1BmhgSjM6+C69C4
3xA1QTXbxVlVC69HbWtsXVzMSE0lqajV/2lC9Kkp5bDqNk0+AukpcVAlWySBbzc9
0N02IDwPfXeejm87cGuQDJNMYdKqBp/1AI684h1OMfyy5vU3OPBqQAFK7gez22Kr
iWdllndAwhc7mHxbe4jpfEigGw5XO4/mUmFe4LNnlDgjBK7RVYspBESw0SBg5HdK
PHK+jIXPMdj/CHXRyTeeZIrM5dgycOE+P7ISLDGvoWzq09Uy0zqv7H6+6QsKntsd
TMES+Pm9CNIklAD49XpqdfENRf+rwyrNs6fMf8oPLOjQisbqHFre1AC43+MNVWmm
nqiGlaXuFIsNSsNumMWg3wR1TymxgU2bzuDZZkMhvk0Y3Rw+VcxTvxAmgrsoZXhd
O0pKbrg1LHVoNPT22xZTYkcZHEfIskggcHXluEUhmqx5NwwDxuDdwRdBHBYyvdOO
4TfRoGzAc8Vt0F7fS4eYn6ruUG6ABBlCo5nC9WoKKmDvSFCvb4cwjPXrSbb9iG1z
3N5keas8+QAhuW3SL786QQ9yK3eTeO6zOYr/D7uc3btTDFIWm228PxMMDUH2KCmP
8BbqideRg7AmBfwuQ1cOrjW+Iw9V6bQgZHlHUXzIDROe1edgC+9hR2ys7ackF7iA
pWi8J+2jJhw0uWX1FHshrLAAXPd3xYKc/1dHnLin97dn12Y6H3brRN+Ad2R/Bmzj
1gRyf5NGVUSCb8YnJ6wuwpKyIUA3BqKunVbyNSb+rGrsG4zdN/FurrJ4LjarirA1
sIyMrIpCX+h4oUSsNU6N1MX2Tda3HIJh+r6vO5eUU/vwC9TSrlAZ9Q1Bp87sjnDV
j/irCk9MXMyvXpyydaHyykk7N6LblBApdNYuuGbe2XtfXwQ3myIwV3XkkEobgD6y
YSLraQglDNiy541LCxOE21H4EFUKQ4gu5IW6vPBwxMDFTUWFq6+IjTZDGsDwBzgN
91kJAJAOQlfVLqxr/jH01+BSr8k7+l3+H9chCXE5VO3Gcl7SnNDbvBSNO1Y0SrNd
QmI0mCbpc5XgbdI+n/nCKrJoaJo+qk0xW5nmmnR8RLcaC/M/CNCpJ5IJxj6m1CBd
fwPjMO1teIZkI74aTpTkGFmcPyT6VDt9Da/hysRH3s56gReMnQooZW5KfEboA6qp
5XiFqL+i6EzJJGLVKkNZtX1O57P/7UEq7lpElu3qDaOE5EOdASZzkMpyHgn4YwM+
N7IrR7B2KSXYsqlpzex5KVa6VI5XH/Ds+G1shUJmWQsYWkmgkjWGRKkmwI/MCl4L
vwMvBEkJl6A+j/CaSZyNoTR/NvGZh9IKZWY86Q/vFNb5kXpyIRFkuhP48OAzTABD
aPVbFJz5Ykaz22YIqKdIpi5In+Gj6tJvwcXfy/KDOM1tMdvXZdqxS9Mqrjpd7WO6
O/C5cT50rdowDPw3wa9TI6YuxqwFH9lT5wKGNiDA+ziOMVb4bG0AgbYjRSHrp6ZK
hekIADefUnsXBVDDydeUiQgvtbOqnVf+7+8zjNpweNW7LCDOGKB0WmFh3W0kq3nj
BmNSvUu2Q0JRjxIG0V50iftKtR8t5Xw7Y4MqRNknOloKxeCbZa0O1a5vncNCW7/4
+yo+kuBntPstw03TigtTeIVsCZXzCKqcbubYelkkKYxIwoWNPWNgXTc05dHsYrow
c1SUt5WTlud6MHHgZ+jnk/61d95LML/PFSivLGhAOUtdIIds7P60HarGsJXgKZJT
hlhYjV547WBLn7oNWyeb5OsjR/wVso99Nj3Hs05FaCwd4aDGQzJ88prZ94BFwjZb
snboDbCSI5SJmas8RuEmVe6uHUGY+R8FBSc2Fbo5fg0bXt8DG79v6GQb0n5bSWJy
le7QVsiRgqcWmasu00eCvE6TVKxTNUijJr1Qc86u3XRHQ5reThPyfA1Gw6+xTR9x
6g7NaJ100nCFyzBCuxVAWzhMvuKuMQTBWbqdDMYe8YrOQqV6v8sTjVv55yH4Z1hF
iKscEEuPEdIpdKV1f7+qwQblwIS9Q5GJeIzBmyUxyyhiSl5lqn8evR6fML33XMF/
E26dIVni5DQiRMtgRBUUimpUWTHMR6jnwV/RWfzx5dnxjGfAaC2PiJzcNUurXjqT
bBnAj3JtF/pVWDGyOWLXyEAWZvq6pPL7iVXDrRHQ5DBoSeQbPVo87dmPsx+mhznq
t50cY9Q3r4VTWcTFdRZf6aEbloFY/QXprVrek7PHzwB2tMRFxs8CyL0dPbanQdRO
GybTE4HGKhN4PmONxDfyxOXE8SPsk3v0+fJiKkdV52QQFS1n/2ztxilHoedBQxbx
+mYx2DPqxTP/NboHd8tu7W5NdUwR/qBu5WevNzopZJqKnEPW+5GzyTzKyvDrOo5T
jNQKfUhXY8PNGxgb6kjssLKeuaMt1XXh8jfYduEnrsnVFnAULwu7GQjg3btA6PCF
xHHNQavRMpFMOQDW7+cIwGX+2fSKcuzuhqU5Dd0etQWmxnou0LCU8LzTfqxyuUX3
P0j8Bhjpbe5AVxDkM0KlX98c4W0QPBOy4irF0K6BXS815Y2BED3Qmbje94OuO19+
Aq+2DmRXboikH36QxHORh5clqar/XsTnaCU2HlgRPJ/tGKjuIsHP4M7vZhc961p9
AzSwR6R1Hm/uDlCZHil8ukc22C8hcugOCyItjKCUUVEPhgyuSmq9cbsE023OQJL9
uUTdHBOMOw3xRjYUtxKJx0o9OY2JSBNINx2WvNlpRhS+uPfffUptLhzafN/kB8Ec
gU32bzYEYW60fvhA+5tQZmiicKfL3m1MG4YcIGTwWAxobwMduqvEKnHkzifwZvHD
vLBCAXkeV5gsd4lIcxt1Xm1DIIunYLmVBmWm2qstMSmmZW5kt+q65HVNU475YR2u
xxs6hUlU5SBWhowQIw8fEblZUIR+ewWSLsjWcB2yknQVG7RD1j1cYSn4//BUqGj1
6MP/+MVPWfVJjIfrviIoScauS/X1HrS4cOiCzMYOfU+WB+0Qgv+Vkftot9ScDNt6
AcnNZPPthSeU+SlaDz1lKEuJALLdVMLPQrdeUjbrl2+OI+7Y3AxxHiWISrLSScLq
Xt13POaLRJXgLknrgM7+7aS+h5XtPVboPVogAkDHAcYCWibo3m0MBEXo8VH+HGCF
p7BIsYkZABdot2M1YTUDYQofPnGSlwI2j3We5b53iH69otDNE8TXKCD2eiDxXPdy
359MEpzTzjsprg2kjIvAtcG6IZ+XBDrM9BJ1AK0SbQjj4x3O1aHA/YGXfMarepw6
ij3sZQGGinyy9Wpqk7yO7OXvBUx9hp4MLUry4lNeYNjW6o5Faw3vzwGhUiQf9mme
qL1NIUHukMVJpfzwxZ8VKFcBBT24vXBfIwcpnaU7NRfX6e0iCuvgL/Y2QbI+1x1x
mIckgMLd9OuubQzWOiInSVT9QCGkcvrrVuNX48gHwarPSOjSDIxuAzi4KlykPI7D
9ZSBXHZCo3gFTQM8OEK+NMLOZzcuaeyGThDsLwb9ixhodlVjTxklUHf98oLTgTkh
RKei0V11Zz7OzfI3MCxIndW/87Fpqj6fijAq88k2XXsD8Tl59neL0DmjetS+37M3
ZpZsUV5rFl2GcQomcXKwQGxmG7wyFJBIvgOZ8ZK/oUXb9kgweM/OPfcNcT5a6nQM
nkoGN0GKoldzJ+jNjMosjG4huVrMEO2GxtgWlJ/5bpjCpSWXkDXOoJxL/q0+YBpz
iUsUT/3Wr2Tl9zgxykcTbXU2URBOoGfsPeE61Ns9qTp1Wj6eq25hJ7L5oGTAAGKg
bH+1s+e7xLzHXtSg6bkn041BQ1florRB2YCQKTUemOG7mrl8JDYlkC98mjHOlTpl
/UieK7qwIn9TN1HliqtI9lbPik+mTH5jAywbeQO7DuOKWpSGgW06wxyALQYpJ0tj
yEkiTHCKVNC40u/4Ym6N79OBtAT+nA6+7q7wyNEubdKGEtR6AVB6T3NKxCrCBaql
HkdP8FqXYPrWqbZF7alZX4JcfzRf/Y/IshPafWcumnpvFEiv2swRvbLrdKEfJrPo
vx7PHg3Y4/rkEQVtUk3DWQ3RqBOq5RMjUq2BA7nyqhW0dV88pE9T7OQTRzQBJAO9
aRnaEU+wSFinBkTb8D8vEiBH7E8nZ5WIEGDftkLS3V01PeElkFovebZXSPyGmE1D
fxZd4rkAZAgsbIF8CYdH7W8icKVFOxLD4SK/X1eXOWfuAssYc485eSodVnRqnx6Z
zafFXo3OrkqWelXyje7F08lwmW5LPd2yO2F7hDsOzwCeORhXcOiL99jYGZDcMrhK
FqmYpsMLTmX68Xmd9OKg5/by1p8QyTa349/bhUojs0jQr28pzABx9EBlAIhfW1eS
iThf3aZtEZGeULCG47Zqu9Q2N3JkgsbOkR5mJ3UYAsaPURwKOQGbxf+nLxYfBcZY
A582Za2m9Gt6wzwk5Q2kygTAfvrM+8ZwToE4ebkYKbz1RN5x4Cko4O/Nf25XLnEJ
pJ/RLmhU+rjT4zfU7QMtE0wcL4pFn0fWWVZK58Ojj/u5tPbiJ527Phf5THndpbhX
J2pJRc7EW2YMCCp3nfWaaFkHjv02NnMxaqwfTmFXeSirQaYWgQtL1s+Qwl4jV0Ge
IbCMl+3zLgtIktChF3NiEylV0Js9XRrU7tdfQ8DObnUBO0r7Ju4Lhl7MdbtR9DDt
i7XX7ZXZAWYqf9WN/x8C4KU6Cf79C5s6acq5CcWJcsyV2Mxcg42ubhBfXdbKzgLw
3IOhVY/JOYXmBM3ta2TirvBqYlM2kveCtLhq7kcRn9uDNEelST1d2By6tmmfOvjj
RDCUtmnQstXJWr6JvjaYPTczxbfg3Y3t5Wnj+XIkihCFVKqOs2p/cJNuy4wD6wq8
FIl8KAvu7p7d3QNdkfXtQSbbmDNmQGVWXswrHGcjDdO5J4UmSvrFmsO0rp2tYiQM
xxqN1XBuiplw/7zklYDgnmK1jjC6u6zwgf4FWSfXXPZIh6PlbLSVPquDW/2YbmCt
yJy1UwiMdhIdySY9xahlKlT1rflAeWGf9LWqy0OheVn5Nm7TYNRyMXXDJwlEIIJl
nGkS2PmN2WmKelvIajM8X5q5QpD1xVU8NknaXSgP7OIa7Ztg9hBFxOmvmkePQQAa
kmLGYAsD4zOnJ51CBV//i3/AYGWMWQDbI+OSMgLhZIn0ZZc3JebffLOYWDVQePfg
VY3lhv069QGEAOBFR8ZCubJs2TyMiynYiJVw0CRDW3pnOWNyhu1A8EutzleIlJaN
kRCPREKuuXLhwCXpIXC3Veuhh/l/FqIE5EC+E4bX75y/9EMnczyVFc7BiUK6ntqo
uEnvReMwrhje5TLID5raOMZzPDdRAFpLncOcAQqVcVpTSm1s1XJa7E6a0Kvcp33z
NY8nFI/dWtTDlg2Z/8w4Ob7+IRJQtDI0AFwn/jrjkrJBEllFwdIXqQ1xXMrL3rjq
gz71EnEnGW0djWYvsSB/rE79jYWDjxHM2CfnwKX48vbhrZmCqVgGfGFvz8Y3nAzq
lMbSICxyzGK92XIANl6szCvSNQuBkY6Z7IfbvoSP0SFsiPI6gpOZLBkvlPfSnfe9
UCiFrizqMaTKqZRaJomDVyfq86Xpi63hk9BKLOyWP6E4jntG4wLpke7LL7oiOxng
cfz6RNMolHFUzaS2vfU9YaWZjd15/JYGBwkaB8xz+VlKYYKTGgG+v+pWXKL+ItaE
Z+sMLzI0TPkWkU2X7G0TILD34yPyTuwOYSCGyE4HONCISnxmr4gVxQcFL3xgPEXR
RaA1/Nsg5dD6ic/8fx0eVM/zs37cm/sF1XgObNKvRUjXN2DVM8IBjbPDuk7jXSvn
sFO12KytWtHjLfBiv6gB3AYVqI+5VEgmitV1bn9u6bAY7eggVbtCLhkyZUz0u858
hF9jC5cB+41sbYP1KiHzEp2Qu8Qbl4tF93NoPfd2peKrtf9f0ObXpS4c1OaVUm+h
2/I7xYkSVvL4JATB5AxgfGRCg2LWb0mwwno1MnTS3U2chAMP/RwRMC+Tp6Iq4cRS
AhwihhRDtOzd/30YUv2eTD7Mdg9jCd8Ces9r/jnhuT8q1RB4VFdhOCRSU4wIHqj5
JAYJ1/m08/oLjcH5evNwZQyvK8US/zDQUye3rhSE7ZtAKzFwIc8bzFvAKBUZ1src
TyWnsBNkyWHia46CTWDfx2esd7EuBjwxcdGxMsSDwFS6mSDy8Q0TDsGun824tfx5
dRzg0dd+VJie350qDNbWcdyfqhTUL3kcmIV5EC5rzQDggb+pFQNEhJmdNSaEjSXf
VnSvJJGIayIq3MbNQw741AMB9cbTHd6obSVzKzN+rlpdwLpcLy9qeY/WyslEZXHn
qBT3+8z5ojft2YmpDb8JFoA5hjqDPHxjQnAQMprHPpPHvpKWScdO3OMbJXVjd74l
1H8s4TFRsNLRMFLsB/O/64gEOIXgE7cI1fA+1Xjb/BBZ5WsP/MbKaKs8xulsXo2M
ZiH52MowPVZZUbDytf4gH/qSr14A2K8YADLQEr0QtDszq5Af132MuhNXAaBKF5JH
YZmpkoYrcF5pxSHoUK9vpefnGDNu05UaAMwnQhEHgMi4ZJ3lV7xNWoXAgLkaE+Gz
xhlsLSdeoNP3jMu+ntKT7J630LRoPi08VO8Q6NXbZ7JNysuDvrsqC3fYmqxjtj34
tZXU9DsbtucfMEc0Qv6jPEjT2YVrPteFf1KDqzMPM0Q5thpQ5vwKGe2Nfu2HIbC9
WnR0mQ1JhBq9lSA4HPOKOha2d7EIz7zJlfchjeZYLfYKJE99qunBgNHXs/ZSryw9
uMQYgnbXWEsjz1NO8hZ8giGxadTBrM/ikceQioq/XLhLsb5FM4FFe+HCzabvmdA5
C8SWnpqdQoo6sOQSGnzUHfI/KhCzCM8M9qsZ58WmG4EjruHD10JFMzOxOa/if+55
rF8DjZQxYgK7TTguixD4Qw4sS9lhHUfjy2CmUzgewMDM7xQKS3Qz0e69DMqqKZd2
TM/Pg2R/AS8fAY7gGXQkfbFY1v9WF8FDrCSnTjmU5rXQkXRxM7szgOh8cOSiEcPd
MkZHQ6kK4PJO61u6IcNrNpEdmRCalHMA13XuVjH4Ult0B3LiRyrUlcQx84Yha+Kl
inm0BJQyclynWvZWAmpjJgLy/tEZ4BZKO2haVjiOS47jYZc42bAe2DQdpKM7Kng2
d/12tudaKAEEtl4V2DOMRbvc2JbGAANhLeLy/RKPF8lC7qw/nyzoypDf5ul+hoKI
fNq1LFfyddEGOkRWF+1RbKucX18WtEjV1c8oH6IjvsXuMpvCYAS50ErX7t0c0q1d
WHbfl4NaDlBBWw0wqu2HD4AYWTqIcYxmNUHqrkcFPJjL/bpvwxwq7LZpswmj9o2D
3i6iJqniFxgcbSzM7xbHfQtAPdLTDP29MgIKyeQ6ACWeg8UDqWmw0HGIvdNIKuJO
OkAK8gCCxFUKIJqF1RssLJ2FLaihzNj6EQCGRjSnZuJ6dZfH4Y+aaoEfs70ifiJA
HukGl+QpJOiHVZgBCMqaq1yV3jfyjL41YZO0b1E5uXh8YyIgOeUxvZKZtWxME1bU
gSeErHGSvx1vlxKMuHvouq8hUMKrEj5BLbm0rxkiODrox2t3JTGPEoEbtlpnaQDE
VKufJm0PJuc+3URSOXwl2174ePOSqiUYuTTesgPgTCKotxTZ/VFJjp/Jj5tBa4yT
Hji80L5szEB90VZwVZjvmP3LoC17LxYsHL06Cx9dTi0xfZzZ1Qzja/bG9773Xu9d
TH4uNjw4SHt+PFa7B9ZjZlyRom7jor97K9GcGIO40M9pID6iHjWEdEDA7uqT2xiT
G58iEYRmdGI1FiKUlSCWeu60WqST2EhuG2/cpbComaISjgrIfyAkJmXmu49PPHXe
JbeDe8e50i/vMhDEfRuV4aud/JNFJ4fCZn+/iBLPSpVUDsZ8sXfNJ3CQuk5Ovvl2
f5AffeckX5fOvaUCCK8hvzTY9ExD2vqMTUXLcEdiPY1AFA4vwl2ympBWoFuscOH+
JYSZrTT63NtB/oPBEa5ZS9rbJfs70AmaXETENfoivnyEPWzbqKnRh36z15/r/mNM
xNBnKZrOUBc9o0FwV49Kc8wNhlUe4B3ftwzkgBxnTEtdBZ6l6zfjJZA6FB9ctMdc
NRch8kX2OAworaiooNlyNP4MVDsZ3fYRSoeBlBa8IVJiUEkBWOQ10WJ+X7ToEhHI
ghxAWoPBiBIB96XqJQyu7UfR0xW612WPflFqxkRDHNd4ZeGvpzzUxSkYiGkCzOwy
WTAPOgObDIdfNCZ7Abl7oUwpo+zZCkcy5HJ6xJvd0XAW/igFDxFh/0rxiJJw51Fm
LCkJUs7bIPEij5hlsNdXbS9wV+W0weZkZdlK5B3gK8Eab2j2W+n4GVzJbsuWYyPP
ZlFZaClZ9bN7HavwzTnx2kBAy9JI3qTCllh0c4p9m0r2ob2K+aeUfNEablfnun2a
7Si0KRWMVPTSw04JJ66qztArNkH7PwYfpU3fPN6zONlb3mGnJunGcwv646gECTFn
0Uno/qtUDjnBDSG3tDwACFTKX1Zctiim2FL9r8m7OMHCtqnWlyD64Ejv2bDyR/Gp
CqZhZQjqEizUR6GIWF+MJzV2YC/A7ydmKvIU5jT7IGrC9oB+cb7RSyq5tjdiLyiM
QjoROSolxGVM+V0mrGNh09HRipkaM+JJOBy2l4TH8Z51Bh5Ybs5ZCcj6w26u9/vu
7Mw/5ikzYEGtr98m/IXCV1cHW7c/fUW/hgZtLs+xGtkdZlHGKyhRlKNQ1v7ygQTo
Hok8xL75T643NDAGNkdaIdhFTZu2fQK22dkG4r71CWSIkKCh8c+8wdbgiiKN4aK5
lDP3PU84PHUxxC3bpHbkD/KXzQxZOCt+94PiOU5KqftT8zqg+8Os5twMXd87VEMX
e1SWYPgl6iElUFno8q9y8jDoStU3O23yHyJ+0gsAACR42q81HQnA8+fJqtnzVZfI
ux7uUkwWXGVpgCsu5odoFC4eFKBFmgV6WMZA2vm3y7e7t24wNCUjHj7+2AucYyzM
EU/MVCSnZX9ZdkLYAOGT3qxqEaxPTtwBnJWPEUZNvPAIjiY0Rbhmfi6V9Q5PhdZC
6POYHlnat7EEd6huoSQKFGCHDsCPBlYO9+tzG95zW7ZRWChzOAZhOf46+luf3Saq
VRaKjUKOj2ByAa0t1cF2JKkDDIh8o0nLAyl9cdo+69QkexPeeY/Ro7ukBIams85V
c8WERd05qNu4CnvllUAGKNHqi1RvxOTwLr/3yDYT2M7QdPvnIVCs63YCGkC9RP0/
hB7JfoR7pCdOYowyBLD0wNccZX027Y/jwVQRt5ohyYDS4tG+iEUD9wIEyK2jGwDS
/etMkUDpUNBvzuxkFFQ/7z4o/mqs7egQ0xfVds1yntJAgpqK9Y/074zDR85koeKn
8+DDc+pDZpgImM+xgwKjlB9/0ki0Q9hO0Zhk+U5gL/QCZeIg8W0iKWxO0zrP0X1j
yoO9GruZUcn4oCHCyIWBz4G6dDwYKk5NRMrkzfP3dfCITI9CWS1BTo4VBKiMFPuh
YL7sxMefVmS0EzOusD56ibx9UBV9QnaAeWiv1SmqtDZOkZkYSoCPjevZgtBeNG31
Y2lIrecnu2vMcoJtTsqiAmIR/Tyf2b6/qYRIQhtXu7pOtm03j/MHY6JTutfBjqdh
VfZXJFlh84w/qmnqEkY90fjQHvymy4rcv6LOBn0UddeW6Tf8oTsVlw+UP9qzMgxo
7BJObbm645g9vB3bEm2hrEVmL8Bm0yNndhecBHdD4om9SnESwmxxVd0nyTg79uGT
LuZgR+b9ryfq2IG6j3HLu4vjeQT3CyjHzrkZj6DQ6MSYXmgCpyj16yETvjaUwd3/
qHbktPzGddhBXPHvrAjmAx5wNgupDAQK7b8TDJi+iB9ashOwAr7/Qr79O5xtKnLR
LmgU66aWOyUT7ms2XU9CrMiz/vDsfLGnyjYV5+5fnX0mhmyMNpak3oRjTRy+cZXZ
4tCgGDXxj9umT80MRJpTslxIu4ph3KstlZ+fQE28z8AAaRF8BBiUiDQt8+ktuaMB
3axaO/zHloWLjhvgJY21qEmRRQaKHGDZz2Ek/FoFgCTDTtJcI8V3DBihBYjwCu2G
yHFWEsU9xOsksJ/U9TapXrs+36r1dej8F1txGWXuORcdwlznbh/ax2Y78+bV//fa
KcQTQW6PpDv9rPI1WgKug7XRbgdteLxPYqCAA3FKr+FqxagD8eQxCcIkfNJHPTaw
mBMZ4eUIz7N8qm+7ln6lZWgwqkUgHOwbynV8S742QtY+IT4Gggp5u0tvSEa87GPS
hNweGj5wF06zbHIwVfvpK7BsWxuy2vMNUJMzYnKAZ7/A02EY6hcdoHYmtO0N2dHP
szfywpgB6IYuXYk8gD4tiFJIw2KbLyOPtpRuH00SwrOCSFZPfSuZ/11RKIgdais9
7E0aowwiT1qzKnVmspydTezD0T4/M4N4ezWfr3c1GnmiOPoLimJjE7rl5+yg7DJy
pn4GRsFiDaDV6vgl2oC1P0TjEareu1GzKXv3NOK+qMB1Z6M9e2I2SeBQsW0I6hDg
GQNBkcbd5nqRNOxPZk28VoUnm3p1l0SdY2qnQCTrcu0Nr6TuYYLi4mvpqIYQWmbp
dl0bb6SaSI1y/Ik+OJBmKyIlLrkeytnqt92wdxjsKaAq4syNwm58ENr9DzNVYY4q
4UckGZCy2WLrT/vt9RdQ/S2loNfddapUvd8EMimbVkSaepaOZx2hT9X5UHKecZ9m
EtXi/xdc77bVNqYxhj4YLT8iTUbHT0o8CwXeddsw3sgv1/7YAZHFB7c5BbWziKCr
WE7TQX6ygpGYlUYaddhjH4C7AMl3Ipu5RcuOFeyBM6XlX9NnQ5CFAX7W8UAjtiw2
YyWOn/UoubWvoIIgVi+2fXqHYk9heImK+0/y2W9d+I3JVS5vvk2LMGKNyQuL07Lf
Oc7W+LQcR3jVmQNfMh9RYdReGy1nuw3Xnwkn/0FXW7PgNDHopP2yzcZK5VL55Hw8
oqp8MnAJAr0BOLkgLmVZBI4E+MjCS9fcN6INwJaEHGBZhSgmvCfXSBOUhJ0FqGrS
cGMrhhPzoTmTce7IUMPkHM/+87fXFt+EDHpDkko+YbWL0KH3l6pIPt+nIv+uyjgU
ImBe7Z4xn/vxdDxH5mzLs/0bHA838E4J/htCOwNlmRwK4epAc/89ppAc+tEfWfWg
/I9XzNNvL/erfK3lOT/spuawQYrUdI/85gjoO6yTbRbuVqtqOWI1BMdUGoeISvAu
ukm3ejUOOo9eZgL+RsxyE1rrovJ9EQdJWU+brhkN3Y8iHDD76yFUW2LXnQRYM1t2
PQnHPWe/4oBQDj+YlBTqcTCRSohaGO/wuqIMYcAa0VVCbo2eNvjtGTuKRbyfKnuL
3q+bbqp/dt4xwd6pIAof5UOIi3ogtTDDzZkwEy4o1YsAz8UnarLPan1KwJeuE3bP
4tvNtbcKsHkLdnPLB+9NdHZJerZ2oOWSoEnqT7KiCLMZTf3ZD4W5wFRIzKFO+jG3
YW1UFVHo7zWPifM8rrt2bTNFzEQYppmSNZYI3sFW6qoPY+PS/OJH/E/Bc2CpX1Is
5m1znzVg23HLuIJeeWytC6WggacHIfonGFcx9kpPMLhznwR09lkB+6gOk/kaSq5x
Iwu060Q2NwoRn0X2pDxKIM72ef2/sOjZyJ6ujf6ySi+cIO/bzb4IrkKk6Tsr6d+8
LMy30h2ttNoYR0tOEZR18oS+gDeTm88lXE0Ge7QA8KXc6pCUuqAKoT9oJ89MLl5a
G7vnMU8ycXRBplth0tg0llvPMnPSKWz8hIOK56pwUfyPrh+RBRGQj1f7ldpVf8A8
9o8c/eYnJzouZgnrJM3VUeyU9rmD0i7aRXHsawSUDlyyv9LPJk5U/6pugBiA2bub
SeoyBnzZJKveLvJBSnOtLvdl3TRDfp5ka21N7WpWnf/SV30XN3Dl++R+kXA49zgX
t7QuI4JWR2AsboIVzOb/vqJfUhNOn9nhzQyTtTWNQq/4TGiFUTZAmqa0iorA7x2V
ID563jWwvGW+Px583DFp8O7KiDZlIvakm7YAwMwgt29A9c/nWZaFiVrW6xR+sET7
+ZhnEIMTGSmIPyXGuHvzxVLjh1bFjf5xKliZhDqdPPVGRPjZCPeDVYX1CBrzEfOo
VO5gQFgz2JehNh0m0Urt12skTNKpgJf8ERtH0cEyiVTF6r/k8z53AFDfGIylx7Oy
Edu9nhzPI5wqk67c4QsNglBS59rnMh/SIZ4I2xOocb1msMZbe9ePlqLX0pQdi20B
pCGNrMTUpheuK3nUUz9LUQ32tp6WFUIpNR+UFXG0Y+DJrBunbcHZ5VAHZyEVyGvn
44VadU/JQ+h3vZD24pD8lt1dH3+I1eX3EqbiIgQam7nexi7S5WkFR4sunXsrIxQ6
MrWtBdxQDr1WaLBvrjs6JlrKhCjQlKA0BTEnyUysvBE1X17KibQarZAI7gLboTNF
ouvrdvT93gMEUNZ8V9Cj1xB/F+BMNa05fwvLqTXwPAItXRFFrgALYLgV2hpkvpsZ
oo9oJxRVpbClYmyEhCUvSA3drrxqBYOw3uOxfRxlyZKj47GcejHJgWWVEwHafyV8
2gH7eLRP1ySxh70Iw4xsuIG1QnjZdmrb7e2YCH+xcsdz2Wx0+vsqBEW1Rwu3YB8v
GmShIvLtm1GKJlueeKC6vVb6cLp63x/Mkzkw728D6pdUka+fnLxFv3S6RTsu0M5N
nKo1CowQjiZ1iTcObpyN2OqZFB1IYWzxPKzQG3JYaztnm6i2mB8OHk7Xw4INWvSi
j6iwINQHiD14MbqzUAoIKLd0regEGjuH71cZ7HAE/k0QRBi63Xwn7LM5/2w8+Ww1
S1zb5H1HmGj9U7pSS5QxXT4m5fpQcYgmTvuhw5osSxTcuKGe48VrTYhOO5+PygtQ
6KfmWRalm5uUez9pG4LO0rNwtabbMGvxTL79Mj3EFBueYTAUBX2TtRsIGtp2Ayco
2zsjei2PzfJAfjGpVBvrTu+T20EEsDhx+lwvfJAQuufpHuMx9aOYlyMlKIaz86hw
EqaiYkmNzCsG3Avhzqixtt59TGQhMUfDWcRNFe0o+JQ6sSuOckUiI6DexEawEHAQ
hg9/ftDfEgQKSSVLp/VtrRlcqmriRug/pQZ30tdEqQJBtJTD1F6JFEwhjgnAJvlN
7L52XQsaB0ovArluqVY+yKRBFMKmk4a64AbgzWhATDpBCBEBNqtzmV55nSnafD0I
CagNLuDh7I1bGjasDoexz3jKL+UHnOI41386l7O3X7jX/J8WdidF7PI8VY+2ae42
MrF4yrU/oAx2RZuV4Y1iYwvNbHSaqDMWddXzAEBeGgZAM6wQgre9GZ5hpIA8GjwT
k07t+GMb834foRibrgoUJFnK0M+rLICZHv8oqGyQaGf+lc1/aezeE3pFKc753gdN
9o9WieZgIoYVV8Z/Bg6aiSxxrcHl2dcFV9G/A0gBKfivXlGQypOuTjdDfhckNmBC
C9FBv2tnZK2z5fLJNHaE74cpUvf45dt7qae2kNl8xhLfJzk8/7yARwFzQlIDlgB+
aWa1QWwaHqzqSWTrawnBJZfhcysMdYazbTzjQa7SxNGrkXfKf1WKz/S1/osnYbee
n+nsDhgH4kf9i0tPv7g+/f0QTiFyhoaAu9p3GR0giHDK8ZNefrBWSExpvUN6g9+3
+oDJ4eNDZqGl1ivwm5lAIF46c2EF18Foommu7wB+ow4W2FfDZfR2pEVnSw5CE3xd
K8ouqMDWYchwRWUbP37V5BF7EZ9K254MPgoIt+2Pi6Q+AJ92sUl/bbNQPcOH/4Rl
VdhunhoZY/f5G+xThzH1zwNO+yC5tVGS2l8XIli/TzorEZmWtD5ZP4rFl5peP4WQ
qjWPsyZzzRBIrBOdzuCq9B7ABqPfL+MpTWFCW7o17Firb1O95eMjvTwPowUR19iD
mRmKZ8eSxr9TaDiJkbxWI1ClDOvuGZLg4JdLdWqn7SAPXWqLbkdpJ1jW6OOTX4xh
nbGHIt5Ux1lJUKOieVXufZNkB9f1o5yWfu9l0dwf5kHOJ/fd8KHReoE0Jlc27d8L
aNky4xnP8rhFGnmyBeSsZ2VCzIZy4LY2U8IBVHp8YUzkw5XWHmdwuLC6PobjrzGo
Zjd/bc53xRBeE+xEzmSPyYPqjorg3/6qXTyrEzFTuTHL6Xq1RwqV70e1J8PIutZS
zgqIahF5hyx+6V1Z0BwGhmj6ljD9vAclT/391ZO7m+3Jf1XaWS23hMBrh/taATQE
1eXvoEtzTWsLmcLlSiIZX9oJuPmDJnMaLM18PgO31KuDDGXWVuD4+P3PCzsHvYyR
jl1ZQtwxyXsx1eUNC+8pnfB598QhTN5e/FAhDObe7Ue4jYEw1QKzgqNthRCBnkJ1
9KRg8B4Z0GH/hO8Nuo6CV6tfq7yt8EmavecGrwd4yKlbPFyfzksPsYEpNjc4xDC3
lYP/P/0kI/5701It0FRhIoTYRXxc0oZbjpNMjsnAUAwkhNgHH8dXwhGIMv8kCR7W
IijuutAXrmoo+kT5VwrT5+fgKNXcc9DWPEKCmM6DwFHR9ySVWS/wO4HLYaco93gp
EEYeaUmogxlRsDo0PL4UH9RDK7SCNJ6Nk6E49ZNiqfqs3itrbTty1Wp/DUl0lrLW
xy9IpEwftDsHNGxR3GyvQTOnJnsGjnL+0lKoW2Tn/6SmpDfR3cy1ykWSLAUZg4X8
+Yf/FFgkeXUBr8aEtWdkIZ1liTe4if0cnpcjm0uKDR0MfxI2wlGStzy9/fcwMmqV
Ieo4Y0OfHphVwkI1CDtLNEwYxy7Xh+Ii9qDeGrS+HMoiwE7gJO8KGHTu43ak3tkL
VemCjQvV29OnPKfCNdUpxcC5B2LaR+LoG+9D/sIgi8e1NDbyvFf0n5bauwifZt0L
fzqmDv8Yzkmx+Y0BdYLq1zZfmYqohRskui318U3DXlfHyC6OHUOhIVKspuVQVfRv
kGT8RJVOqdAKcHrtZIIEs9aHxj3RX5Cq0XZGOuDOmCV9S68bYt47tThIm7QDLCE0
wmGaGg3LPyV/rphmOGMDkumO5jgST3mqYQmABeWXUkDQqIhUsG14gN7PyVEx7SJJ
H+nwrwxRH6DLY/CQAKqVl6Dhfa6Ka65bla5q+GIRiV9OTihJhvjjJgQnAvz8k206
VXMqMrlCzkcE2n2pv1ZpNsAaDkbC+DyMn1jOM4PZuea4GHnTRIZtG1yBcEtnD+xt
XHPrXv4eGJeEpqfDwgiWuhKtLNZ/6vP0FzaTsliQPRijBsSqT0dgOe891GaQMI2K
mRQm7bZliT5vX/phfZLUeKbhjRfDDIw8Csjnx1ySk+nj2jfdh/vX1KC0g5O4p/KZ
sZD7F2YldWpybtZx/lWacj59tJUrsFMFL5tYXlYHr8s=
`protect END_PROTECTED
