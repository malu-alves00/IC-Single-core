`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GgZypw0CjdoQGtTpLBspuUCX0uBOQxRbBS51QFjNwVTTipFGK2s0//b8AVpMoOSt
QlNtYUU9+jfaG6cP9xJ1JsWQZWUA8ckC8MC+jPkxUVSGwwNNqmASUvTUoO06FNtB
36QFAR4h126yw8Qi9yLGiSahRWFo0dUFlq7O4lTJ4qqpYkfQH+yXXG5miwc3WPRQ
OPns0g7uqFsOe7hbmLAU2tkItyOlj4wu1Q09GMaZ/3CszbXgwMFTibxD/QjWmIzc
+wBCjm9nhUZ8Y8S4bX6zJyTSo9mjFPHNKJVQCdw966pizWSiXeWghih1qpngBVTI
29cmt35OhYY0lDEMbiJ297iI1KL61KhrNBgeebhmOSWb1mvs5nITYFtZHxQ0M8Jt
7f1bPFm2ujf3kf0CYQoL7BrB6Bm/YETpcNyvxccANZHPrMSRhCFfU62Ssxr5qjsc
MVqSCd9o1dgbvCgPeJ9KhratONufaBvtv5kkXTf0Arlv2QHgThyTiubeKmvQ7gKO
i8hpxqgXve1Hgfy1wAMYwmTUDF5HjKp/UA5HZntrmj76yJ32jJKXRSL2Aq2HNpCQ
mvLF8wG/kJ9q+/vT+k4u3sYMIA2ErAT6h5pOZDVmRMoq8oW1bG6EWxRSxeWrJr2U
GV5oDtkn6/T16k7pqzxypWhnXAuIrgjTx9tDqjyE1nT9ndx7MtRjLcJgSClMKncR
z1BpGSvJy4KAYiWR4rIGADx+z/PNibAhFtvmXzzE33vI1hezLDuiVAfoAM2+tKKX
D/6AGvvaYSSjVh+hLuTTb0OuqFJP9MuEXdZfJE6dQfjZPonTWo83gbek5D0nSL6X
YHwLS4G5FOXHmJ3lhNsGR9fb8mVFywf05ibVvCxbLvZBZI8rpPI0QV1SwkKtJKji
Y8KQcdrGDRw9XzZ77Lm+GJL1M4kLkm3BSa/ULTdr3QYWrA3evydY/gLcs7aIpjbY
ehKtLmZB5jiH5V9/erwGe9z6AnzrVh0yZ/UTTgXkVRBY+qzJnJ4h1vdpEUHZLeWQ
k+MdhfGN/nB45I8EE9Z1SUnMClhWaijTwWB+yYvnX+OLR6Wrn91Af1AqvfF3GbiI
EmOHReWM7E6ur3Dn1hbcncbqRRtna8NA6t5yDLzr6eG5e9QExLrbr1nZ0qVGG/ow
qreJT8DCWRAOBcULvgkvZ2GKHM5CnO5oNR0w1Wsj+eTmrB4OWZY9NXyYNXfYQlIz
lXJKnCGVRiPnI6Va9EYgGeAz4yxB67H20I15Nv6BGyly69RH5W2J8H9YkwTPsWcc
nuNpKYZoWeAsdmU0hwA/KX3jwWlMgYGSHOy7+3ky0zRakCZAEuM9z1w3It4+muFb
RhRtsw28/V+HCBlnbOHD/Hcq0v62xve5uWd+6ziWCR2nzQ4eJuMxyPHwmOx1fMnq
M7P/MWdhdbHkuOo2jajAmlI9Biutdr//WFiPIsPHLPUGt4csdf85aadD3qXSbzXC
ePwYBzHXrpvhN/KFLXh3NtaUSM+htUNyyK6DmhgDE2nFxh0s66FcEKbbvmt1Fe6w
aa2mhEZ6eC8Xs4DTXkwiHo7Hf+ipYfww3s7dxVi1hVgn22v7EYsUu3pUqRLZ1Add
oLFu5Jaa3ILRxdXSD9kPtpDLjhr8eil7wqtHlnv2PmDfFfNq/R+Ji29F/qlPO7Ao
pOoLGtlZckPSc3WFA0JraZ1ujglZQB02frswTDEs766OcXeb4SDVAlIrZsoiSEKw
gyezqCxWO6NJGnl+b/aiI1TW5g4jzcubbX4dKu8/IogleZONrpKJLYR6ZYyyN29J
uAc6UQ2gw5Md/ECBgHcMCqMtrTmIsF/uNYRugwbfpddqPSn18AWUonEHw8zdwkkA
Vg8gGD8ypC5nWedby0uNWysPnU5BAy41QpK1HcBjt4h+hY+9zwMxfBwxUx2PAmH1
h+8WkFZh3KIxw80+wji9V26vKyOTH1GZhOVBs8iciWg=
`protect END_PROTECTED
