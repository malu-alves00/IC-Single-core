`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sNyBU9HJXT3AZDY0uD4eU/I6l5sdHeTBSsIk3uo9Fb67zJqDu/TVi1ZQ4D+sicBb
sHqH67k8/BykdfeqqfTklPYdw1RLo/ONXiK9Sl8U2guIGb6lcckMflvt8wuuJHii
Ant/dkXjRZLos85ffIuQ8D+0UXJmp874vYu2THPGxgAmALYmRnN0tONZqPr2R50L
4NbSKcx5vUQduW0glvq6E93KWBzznXXtZTgRdkt6g4907i9sSSmWyg2jHM4Ob6W/
fIltKYrxrDZ/Z0mkqMsSXj/mSR8vLQcxgndZD32pf3L3QLdravdlD85QRSpGTJx8
LEUttBFZsZhpnS0DaswZ82Pm5LNv6s7dnlrHbsv+aWo6jdUofQjMVKPWbVomzTzh
bF/lm550taSH7als9fmV1AmdEq9D0QTrAWVFACAj7FRTzFdAjTZcXmxF9hsmlGqk
2rgW0RabplVrzynKVb/jNSMigRAsDXSLzr0IJBawEmP7hfgFrK9xZDXbf1Zw92zt
jvKYQVgAOjzCUZQ7HDBmgUJzcOVz7vhP5efMfowl5pTWq1xqcuaRkYzjjhQlHM6i
ujPK4ZXh2iECmlT3iiaclMC3PWpd+xcS8crgCmrMWt30RHLQNreEI4ieaRQrgb4Y
SD17i8BNqPRCfEyUTFKLkcClmB/YQwCk6ui4UYeMbIcmlMBNVhctbJ+O4JFcuJ25
LChI5BXVgtOKrSDymcMtm231U6Se3QjNT9rfXvxe4QNJnj1aZH8yHyFlqrabMZVA
Y2oCuBLP72PgaKvb/dUCA1ohtlJ93QpmCWkjARpVuHdC3ZXCCF8CayAGdb6QNynQ
x/BgMqKaNsMDD0XhXZySYq+q7Zskr4bmN4P9y0TqkDMHufQVuxq128yOxTtl4JTS
Xy42cVEeR56/XwHvThFIN3mphi3aKQJYPQqIeuwulLE1XYG2tvo6+MAdauUXABE2
kcUegVvyTRDi/Poa5c5QPWiS93Ai0eYrWIQ7pRkgTkd0JUpLnNLVTpoC9o4M22vn
oQHP3HHvQB1uqIiKdcH/5O53qyPHjatIV7Pr5yECGioVU1TS6LQMeQkNChctTFof
tEaBqdxg3ztFhV1NALG3z05BmaQk+Qk4B6U23DRYu7Th5HuK7IYGgJbUOGfNILls
nJQBNAnlYFEAmnuxi1GuN65tO999oWoQXJ08JofFnr8PRdEQs1ZGX+0VXxh+PsE0
5jlW1HIFZmoaKSS2fPdC9QUJmA/PYenx5s3xSElXNIGQHVaf94Rc+soCa6Yy9atF
rY5hMOTX6ZFtU8b+b33sTGyW69RXKb3Lj4+2aqn17RgQSDLLVVsHA2Sd/4zdzIl3
dtINFCe81q1Q7kFW7jbHSasVqhdmoSKePAJBxUxaAncfpD+8UjK/ZOGaCkVAJ3wb
IaQT5eu057GmsDbW4SI4XSQ/cnDFAy854A6IDQlaazjrELG/2IgvHINJTlW5BuAw
wBLnu26hoW69PloafXTrLLT51yOxFQ7qtfT1b5wOnwMSThE8aah3lYtL2sOWozbz
Mb7evDcL5aLsKnZlDN3LoBdLz/O5+3y9HGMxsvBGuJleoHeuxIBWga5HPU8ttMB7
sYUceeEz3P5mWt1CHdsuOqZHeUwwtHSKsk1ppCG7nusrt2eZdDSKpaLGBxXXuKOV
0/H15PBZaiac7UuLXICYgAxrpavxVi65mIXn2nP+NrBF83Weanap5oYx1Z4uXnT2
Hi0U6liRE5jpQ5Fc0nvllG2a6h2NxKmsQR/t2lK9SkD0fi0SJGPeA7lqdlb8flZA
c43W+CiuulRYXjd2F7+Io2huVtZMC3xrJMyweGIaeHZWizZiWUt2DwDWPL6jv6gc
BbvIi6461ek/7R2tT+8mltQQrmikz86acRBNN8FO0buTNNNW1mI7rsPIg3iZWchB
5G4Nh7UJK966Ee177o1Mb/wfkEMitveeasODGE3lOkiLlSWb6tcvzcRjnjXx9kYs
C1fQj11/myxgzAxt7JUfSiPVigMzkhQ8Rqw8Q51UZ6V7YoIHA+Z6zK5VYf5TTSlA
2d2T9vTv06d9g15+SHfa9X0mi8E2BfSD913caAupEVwsbV+z44QhnBv55WL+3UXS
uX+8+HUmP8lg5ixZ1RfJr4Gw6feqinERHrYhh3iiYEDSkguK4w/JJgpEPgcbMLlc
eLXGeT9VBovQPV1hJ8oL3IYNS2oh2/JQVl56jKYn2e5LSe4mUaDf8IElR4NPUVxh
B4kE515Dcylpi7s4S85MN/L98w+EU8S0DIlqbUUMQhEtCroxocBCEqtjiDuGxWqA
6mi+RFIEwJb3hBSTez2We9PbbmnV1fs1m9FaLwX+xbff1GP82HDIpZV230kGQo+X
IdvBd12MIRVeus7+NCx1XgTnbn8g2nzflD/b8nAOKjmtuIJjZ6gfj7GfNRCitTY2
fEo6NFirxIc+lH7xaglgIAanthUwO9JYqB8/O/Vn9TZwbAC2fdBjvJgNFMu6t5gR
ZqaqhMm1VAlCLWXoS91JYDMzCl6aTtsOT2FfzblN5eI3evbaKVRtsMBG7JLAJICb
j4pv4YpdP4o7yPYIDvWiGQaURIWHwn+OenRXD0EZzRTeH4spJgLEYShXMVkKOSPt
LNRS8P1HOOBqHbxbauPLua9ad4IIJZMg75zaj3mPJIka5yRgqLoaTT7fveJf28eq
gGGud3aGovw8aVStT8RG6bb33/0Apqk78K+IrGB3/fwp46LtB3litOajY9TGvsB8
dd4lcx+gT3CsA9ggZJHbsK8fMHkNKnZ2Mbyb9rHAvXb/ZLZaE/c45V83cQX8VbsD
nkph7986ZTISKzI7rO10nU2D+7Bk13hVulithxJ/pkvTvjJrQsMRqIW2cJmWcNEj
LMhGKgYD/bKlfdyoNSJLIrg2APctLnYyYxJUtG24ghLd36C7nHNeSAh07gXaoz4j
h1B1YOex+Rz9rGyeWxFFjRzzdAYQbWfS6awS9LunpR3ybdS1jAVGs6SPsYaI3iVA
28klObECZgN6sIGAhbuyJal57ypRK7BuIz9x9w/gDY5AY4EzSN3iufOai7v7NkXP
8E7FWbne5Bfmpzvjr6qjU98hiYbTn321GheCHCvn62dwnVEYk3BohK/EP3R29Ibw
2mgkIl2h3MSFDr5CWbH6RbIpZBjQ0SiawpKFNRqL22UZZLets18uIRWEuz0eZZCk
EQ2FHR+6VluYsUYOQktwdofxYkEzpw6CjPJfpu9Oo1lj9OksyG+IwAQdQ4+89hJX
L17ZIV9Ueevv3ZGlNyfsteyf1eDX0V4fPzF7+ud/HlCZLocvJbEpNBtvPVBtafej
u6ODNGI1ZY75nj9/G1JzJ1hCELHa9ISDA+G+NVetyOVKd5E8liDahGRVrbZt2bN8
/qsddja3Tu+aZn87fcpNMdcRnQiax7nXTrSWaCJxxzlokiJqQq5mkFCHkh7pmO0J
SX06u1/PXnejOMc7Unchuwq86/v0fY1nUQMB2dMc7PiGJIFA8IKkSHHOgw593IN+
K9Ymdw9P/mxGJaVZwfyDZCNR39w/A958fezUS+Dt7KuywlXSsUqXdZrL9vvYIk8u
L+9zUKWhkO3r7WBq/iin/ZkEXc9VP/9oQE06GOoxxtu8PVGhdp81ornBKkyyNMNp
lTL9pe8wEOa58IBKhhM05u+cGEUqISvZ3QQdNDY5JBu9yvi1gx2eCVxUP3oEDQMM
nS2tMWAejv1iQ+eacoxp12EP2yjndeiKsE5tuZKmybp1Br4B4H6ozMIOciRbMAzv
1pk9xSAlaqNLN19O45OLhexTC8k0xT5854EVJzwtET4WJnB2gB6FQnqOIIvPZWaB
zK360zK/bERs2qy2EecDb73CZzsu2ywb8Xxe/ny2ZwwyASFHwqqTkk7XAjRFHnO2
P0U2fcwLc7X0dC2+3Pt9Ljmu+odLLfLUDOSRwwtNojjksbPNegzZdC9NHbMNVgOA
6DRsI7+oYlhhfMv04i+RQcXYshMLMOHNgDd2gsA0iaECXajvypHfjhcQj3xT+LYy
LHFcuNyZKPV7EoClXS0Ud10CLCOoxeIiKaQqGa/bYKjThonO7bN8iK2DYuXCpW1C
t/bOlnJdR7jIOPvhqeRDl8oF6s86RNOTUlx/KcC8h/dK7tcNNvOkDOlMUb3PjWCc
c79tdZXkPIK4Fm/Y1/54obn0Onb7Husd5DiB7s+NHCk2LMOKBsDJyRFkh9b/ub++
ljDMbG+uHd0DBfphvZjC6NrLVfkETCSPM/Vs1zP0Yu7Bs3yVca/xDPBiw1KH4cF1
/tZZCoKd8YpKghJpcuMyWaVCGfHpZPCKgXmcEiDg8YsyP9tOXZ+ibC2tYjQZ/GL4
O+pcoUiTk5nZ61IooY8Kxt740uCkm5TQ7TWYEs8wVNqP14e5lXvG8nJavEAyf5f0
1DtlwVH/Chd8bltvGgmsxIxpfFdNHwAz3rWrS39Wt7okA+uwA1X2ZNSlo8CzkLiY
DrooA05Lc7yNeuhx/3Bbk4llQxntKj/Ft7W9s8oBz5A3cjUhV7hcFw8UvAKmyhnO
pEWUrI4o1nfyLhjlUQm/X1MUvDUylbrZNO82vpCC3x8UkLo4o82auqdRJqUqRJ4T
GHQFBZLU91tBPIDReYY5C2jQQ8K+hd3Q9dE+p/sDVv0oWNZMxPjG49pb09UKd+X4
FqmwaLDe18621ZLPhYptkbkzuMYyOekq7aic9JNyGYIGvSYWFSjc7+itew89eD95
IdA8lyn0WEuUco57Q1fOfUN70m1oJmzr3/KlZ0Fsy4wK3CzWJwxQPdORYCx7woPV
68kPkbq8GSuiDP3SHHaOIT+Uznk3FC66SjJLj5Yf0ePI65fE5y+o0YBldPXGcwem
HNLkVjkrVgelF1Wm5sEUXM9VkuZz7RNcAt3J5z0Jn9sduNtUbSoAW7btvq1U0NWR
BLz+FwACAcV0br0bemfZT4vBcgLnJQ/bKbDNlXXQRECMClYVCe6tWjm3riY+VqoC
yot+MVbQJ5D8PWY/+tyNow5n7O/lMrrJRLSVZVvEwKw4mZLZhncD1V9XaqG19pwi
+Hq+Wf7GRVVVXQSd5apWKMM3Pe27Y7cHpkvzN89zk34t6zaVLffyAQxgoVL8Pl3P
tdjxxRMjX6ra0ra75BUMpMoafthDV2qOGCNdBEFSQaPqQkMC+UCLUm8ExXGI8C5n
RVmjnTR2/Hi75S5we+8L09OwYnfWpwiqXoJGW6l6JNvoJBmE2EuMSqXQMGlUpXkK
F2llX4l5HVzsyFXbuKpRpq9cTHPcKZdpBJUEATOh98i9NDD1ke7Yd4pJ++HcR9K/
oz3z27oTY2Ucih6Nmn9i4jk+Gq+qtB3Sy0gthf22oUtZA0+3ytC4aDfV30hx8Q4t
2Kpjs8X7rCtF/nB+B9HWi9LYohEisdFUW2kdl/zaIhroES8jYJBHBRjR4mtBunTf
siMQcrCOqS52ta/ib4UrYMeFnQ9aThwLqSEtJNaCgDN41H/DVyFPgXXoNwHYzoJ8
IYLahCtCVfwXki14LA47XYZzdcLWAwlnFy9uW8gOxgyiUQvnRnyiHV0yjUKrdZrq
Tw2rvAWWOGWXz/cd9M2BjWpg7SAHL6lCJSriG8jUai/IbAwi8MxrOPQ+CPaZpgcq
6kegDkapv9p4fMZ8D/ZZIcwQhj4r5M/LQ5vq79tLGyzZQ+Lxh9IoWAYEF3asWI/d
rC4SoFOYSpppHk4RHaFto6TAbW34tyjLrUK0mf2SRZnnu2NW00bVE2+1VOmm9ZZK
7y8pOumo5Yfqa982QpqPc1xeSNa1TrsCzUEgovJVfaQAq/tjzWrG2727tZsc/Zvz
fD9SExLa3v64RPoeCxKKndxdQi9WabC5x28mA6ddgpVHrpVVDy5JcOo2Nbr87joS
MeJAxo1k5VeS5bxbr5ZdnKJITn4sCGi9I5IZtQJYYszZaMzrdTU8vnOqF7jACIgK
Pi7FPr9rcW5NxwfqNm8Tk0GWVMUOT19BHZg2iCY8fSIqpV88quFiERVePX8CGTEA
xBIWAJ/PfnxbV7+tuKERyRGEF9NxpEFzXBHbRo/VXMDk/5b71Fiu52LK7x9VK9on
8BomV0xkpU/VQ5UQWU1jpMPWXAwqCuHI3fYviQwgpX57Hq0Kl8sOkhd3MdyhCMKm
IHR0ySe4pqJYaa+pSlt6dbaWRg31hRApBJ6YRlIIGOVMGdEdpWow3ey0XyXBVeWj
ccZ99LCiDLUW2EJIG2BsCN9S86liVjw8ndoB7s0PnACfPwyy7vtX/nKHKcgzY4UK
rQcVOUkkiQvcFn7IsYwaSW+j8SMuKwjPBAk6dNrP+UBh4hCi56FV8chIN91hcu6W
pOIdjvwoaoU9mQY8KdUGAtA0+HoCBDY/iTpoTaqvzMkn7//f03jsKhTmwzKY2bHi
UY9k0z0DYZO8iYG75Rd8i/kst+zgBBDsTVElsXibf8wBOtInOjDrP8JcTD6v8rk7
SUc2XIFO8Jtm32Hn6TVwQYp8KwuXpD8hR/g0SZrjWY3qmdBfIYS8Yjcm910sSg9L
TnGYlLxMLVeEJd30FUT+PzH/6IsWZ/TU5Ex10nkz/4SCuRTQ4Cuyj70hB9BDNEkX
ZHABLXUVwd0JSraq1JwqvCRRnSbdxdUYl+hReyBWZ//+nu1E/Frdc897e1r86nlD
T6/uNubuJJ4NzsbJYV9MrpnjGjVxWU/GTBUFdgxwsAxXCmgjtf++b/Nze0Z+gGXu
EFVZk66Md5We7SAj1eSEkBkJfuarPxfyqKdImznUrraeoAxNwwQshkLKy09OlX0I
o8uYNOAdH0xjNQuBUNVeCt22huVBfgh9ivV5OZSQgrco2HUNPY4M1r7YJWKWoKt5
uDSPqWpMNjo7wmZtzg76P3E/HlBwx08T80CRgI4mVeuP0117kh4RedFDE/PLd12F
ENhIMxswr3OcTVuhn3LzsR7YruavPDJlk6ZourQy9NcFafwKGwPIkWcNGeBLgd1K
fupiHyjSGPgrYJJG+Ov96v9CmEePpAm3XDUbo9LROdWi1nv5OcYVYgShQDDaG11Z
bl2lHjEDAGQSQq6Y2ZnfPhSc4wbbII/8jUKQdjZ7oMi2pvOVnRlQSx02I9RjVA/V
u4ui2L34kELNVancqmgXF5qUMc3ae5x0Ukl52c7PcX2Z7vmbgq9eL9yjK3Gof+VI
VrnrwIVkVJNF7vJnk9xjlrT5i47JwWPyXDZqyUmLTQ4I1ngLPZ1r1yzNloeGryHj
E2p4/kdXtW+O4xvQtM3WVQKFhXDckZe8mYCMf9Y0bztVG7sS40BcWf1qmPnb7xTC
Qmtt62vKP8jKGI3I7CuD2o1gTN7pn2toq6C+t/YRrrFbGDpgHsptBIUCOgxQq62l
pNax+RRl8RZnkSCm7D2oRuFNvaGSlg2+TEUQlTL0CQ6iwR/sfAy33CwyIuNYzQNy
IHihpmLdvgR6yqwGzZJWnxUAUWfh8k7faXdzPq/ha2ALGbNoDdK6hjNKnvS0U57z
Ajh6dbPj1chR3gmULVv3v/FoRn3eidI30c/kTtVBCajKS72ji2nOLgSTvKkjzbsc
SkNbot4wQHPMZ5VSilC73eDvLyL3ppexpC2RTD4vjegNZ0/kjbAlnp3IXrNOlOM0
D0+AA+9LE18OHwfdEBcl7ScPJZtQAsU6HhsLhvm3BcPz9AP241OHA1EQJOTz0nJ5
xGTCzTcR1VFMg7HXhIvSC+zcKr6mdj8Pm5nbQOBH4uF95wRsTHOXwFr1F7M8eWtV
z2t+sa27gw/BD8E1+kTo72uY20lQSeRIjQ9CAXWer0QqSEg1gkN9Q/EQRGnAOjU5
aOIZvn4oC3kCmUCfVkF7X0u0ulW5jxXf0SRs0KHIkodEixomj3YFDOjCboAgM10h
8iGLrD3T4LKuF35cIeC6zudz1SnVC7dXNHBk9iR3LMJyHgBCHxTFzz1LNOX338km
fx0EDx4isws2A7whEPjL7jtJ+KjO1mFNYGzCFtG5vDkqTEVxe5qQQolp85VtYQn9
/v6HttORuzfldyJsdxBoMXB3L/v+KeByq6hmfXzXzAS0ubdnQWcU05fLRN23AZbe
ippLLPgeUEfrEMgRfG/q9pv45ip7IttY+0QGQEq7Y5BHwSTgMhXRuW9PBJHCkRu+
/bxdnf4xALMj9nvOSPsChaGExhydL0WpYKCS5ORBftjy4K6xFtTnFaFj0O80QUG3
4HwmodZB++2B0JS9yQkoET3sPy9SudP3sLe2zpNjITG9TUpe8DU9hlUHYmzQxTpq
ShQFHUoP6MMJiVLt+JHgrrCz4GfAy15Hu0QSgzJuKoqC4q8mkOAIwaiup2yUg9S5
gdVU4QGnxBXzKpq8zKACPYZe1Yi3iVySLm2byj39GGynRgpoPGxKdOPIEMcJ93o4
aXr17QZEuXJ+ojn/I5cJ8QSCAWGzam8fjbrlVS6AMjhp1B+w1UIFW8qcGDvVvRP6
OhuYZHUxbGdDLVbHDq8wczf7j6qryPqoyKKJWw/rQI5wCJrgsf8uEzOLNvU2D9kS
mYAhmX1EInuXjEy6BeH1Qrdubl266zI/a/r67w+hpW3PCFl8gAisO4mFhZVEtzWm
lzU290PZkCEo/r/TxOYXrWAvuKhysBZmKryKs9JTYk8bt12yFMl/851w0e/In7lX
DE6hPNUebABw5q7MJmt6mRMz23KJsV9m32NEz6ARaHLXLyAb8hBuwQBqpEHRnSOj
mivNrsLG1eYY4rZRU9gcfKMKY8XN/+8F0sR7S0l2/c1kh4/ZZHv5tajdHeRLDdP1
JP9Q3idusmxhAieqeUsxA+98XNbiRXeTfywVfCIiw1lACPODg8isB9gGwFKtOy9N
fTOTLbcZjxkYwy9P6f1j+jFPS+CesN/5LdwwGEgdmLtYZ+VXeRgmclPLQfKFTsai
lKIXcG+9xgsi2E8sMVQWqcK0DxNGFYxbTYudKo3F5lrXMrR2pz7Mpo0S6c6WklTj
+Y5FJ5OfGWrMsn9FiatdjdjP2qSz0PFay7j7hLQ/V/vOqQGX7Ur2b1fu1k+Bk7vb
p15KIVltPqQB7eszCYS2kQXEPGb5CWRxeHdckJyB3iYq+a3Is8U65suhGhRRWZyA
NnByjieZRLxL98+snYVgEBHTnh4LurKGRIW81ytZEAmtC8ovN4zGTuVdz8dtwBTu
43IjGBvLNZy9BEaB9aO/c+2QzY+K0hWdylxkH27s3pgTOS/rAB4i/WSDo2mirYHE
uLgNwl+5syczV1Ss/2HWExwUFM57n4b9+Dja/ZWJWexhmKlvQlEkgX7PK8jaZcwQ
jb1ioraFL1qc00V2aRVxnBZfWhRe3w5fldsuOPVu/g2jLZ6Q7ro8BCd8VFp7vNkU
VnXR0ED5Q2T0CW81vImz922JdLLlyLtbDplUHpymbKZ8jjAQ573DHnjIRCVHb2XH
RN3M3YP//udCZUgI+0KicAWg41TZNdYmvL9bz00c9KuPC7VREqjjtzr7jHBGZsbS
tYIkO03zHsjRg2/nW9CIULnHLmpikxO6E0wLmeMakT4lHxQg5dMRG/tOmfYv1INI
ZzfBZuiXSZFzLUTJws1SdzJHhc1QcvFrMZkF+kAaJw3BAicno0twNLCctCsA+viP
m3LLt9R6SIulbvLdU2W4HPHilcnkjVNj7dQ5jn3Mgc21aZrgTr8g0jTh2Ix7Ar1x
xwfauWVRDHGz2Jd7yG+Pgxtdkoq4OhJBpokKTwUcGvUAJJOHt9iX3PHMayNmR4y5
+ayZCP6lv+vLvjMtOa8fc8tGTQDHTqCxzbR4Lv94LjMNLs1QIK+LJ+meRTT8Cn2/
JrvyYd2a67PGJ9IrLdxXzmMgknGVxOg+2mO0DqrQao6sMbV44HJwIx94jFaOZ6gi
VSfBr56UoT9oW/Sl7Zuu8yZoXr2mDALQU40P1vJkV9LeVTe1iyHhYzifD0txFOT7
9I01Z9t0qo4fMqG5cCxQSjvARhN6eEPPDMf0+Oj7yoLXrGRQaWnR6MRHiSfcWm+e
UlJw9Dh8vItMnWwEYsVv3jVs3cVosk1I/wV4WwkPz35qmqPaisrpZ8Dt2Mrs6Vnq
2n3p8ohAduvvJx9xno3dFjyC6ghMeVJh/toPaDFKlm3pjvTlImI/rfJZCIiClaNe
PWcNckP16HovxzTWLPQQYpwVRVZXlkfAtpFul9MvbrSLTsj4CRFV+FByQybv9hNl
f31r/xZ+rkADPYEKyZSLTGnOTEGAAfiB3CeS2UZrHs3bB4dSvhLnCwXTJYPBfty+
oIpy2IVgvqI+lN0phopXWapAlsKx27J1+moOljui6wzrqcRMv8D5azetrfq4zRbS
8JNF8nyZWWdtLbj5vES9Roi7eyptpdNT1nNEBXK8vLyA4HePQ8RjGmvCSwiZmFth
5mIjqVPg0ynPPsPM2c6TRanWuD2u6VZPgiwk8N36GM3UMMnmO4+LSi+cBsaGbXLO
T9BLNw19pD0j/Fj/M9Sl2Q0nxU7F6ORiuESiFMMmMkVMb5Ou6Xw6Wo/6zuEpfb8y
p82CDtA4N6bG0nyuC/FH2d4Uq2BrGXuXyt2XnT2oJnmQ8KpVRwIl8rOYlozLpet1
blVtijN3/oSSYYAXKZq6Fv0SxBR+3ZjDm5i6txrmds2HcmKwyLHxfOqAPSQq7YwV
XtbwNM2sOgQIWxOOnyi3SnAToTzug464m4HP9KtMo/HCtNtPFpbViT8D00lJGZ2E
AJ8SQ46Coou6BuqHvgmR1qQBnXLZaWGsWHKVmNQwT9zDAyr9OUHW/T5e3Pdw3u0D
swTVIJR6fVJjCZwoJhVecxV28IXKo23X5HXXxoq/0z0Ha3B71gQCwY11ySHT3n05
zDKCPYsK1eJEsdltSSncMC98Xcazki1xnfaR7rZAIxZni0/rJW2K71ZTIPPPG38W
XHWfiPFuQCfdPDOPxP6exXHthsLPzJd93Tu1QvNBTv1nBGkRZZwgznkQwFvX0yhr
CzGqB1Xb+NtEAdU4j2AJSkBK++kYR2xCAA1oR/U/h8By0T3LpcBPeqbK+0svS4Nv
9G0l9ZLP3syzO221s6enI1nvL/t88nZkFgElbTjmxuerFYz4jFfwkR9WAgqrkjKF
tHkbqEm2HF+PdVvMzPSSudFThk1DhEsdV9j1Ak2Q+ihk7hEsIII+ZHzqkEdrW+H2
OElgOgGTgXiIZlfPifVi2VRDe/kiPWCtUwJdJ3IXhOBe21JPfaCoBQPj9ns3OzsT
Iyi4nTpsjpWH624iVEwi+VMxGV844f/SxMbeI/9htnV6Z6RFjbT6Cc2RNuFivMR8
w4+oriV/Wa2Im2cjV4Y6yR3CmMdPtAH7ivGtEyRDI2rjn6RPV5FTFJPafh69J7KF
lciP+Yd9xm3WIiIcStlYg/qtJfeEmntbXUzxTY+gz/fuACMnUwV7p6WefAJgDnbM
gUNd1RSBi4M+64HHcn9JyZP00IJGJ8EH3ETze7qIN7XZ3Asym6kQe2gNPaDEn/1E
QtNEb6TWs4i3b1J8olu0RaWHajHBwZQekUFZQm40NTqdDGvxBOvTb7IW+8GdLgmU
RBHT7+VBuBDT4DEJybbhnXrUkCwMJj72sXTlRexx7BdCBrxLhYvTy53enGmqjrb3
eYyJHahQqpIc27KfwjXLZHRpuDTOLZKlucypAM/J/gEAVVKWm6WNvvIDJWw9Dmgf
ZGGmScznDKNCrew47+ancL96+mstRe1qeTzd344vIhUs7B2vRjnm6iNb1mTlHQxP
1XMZ5/leqPGaLETBDaJb9A+wWV/v4B+QqeOMhb/6ysu6CYJDVA1kBpZBUkwjyCsw
nHU3lk/f0kLZPSaRM9ePEvQ5F5WhZVU2tQcHJ7geYvJRJTe25nYmior2Xo1Zk7zj
imUGqN4P3DRtBvCvxbn0FOzg0qXeNrdczJsvmU73CEIh25GH0OryRWCmwUtsYr5M
LoVvaoGtyZjsOi8iHksgSShVPmICOVtnDlWLVT02idDgecgDXmkR4r6pbBaHLIOJ
MyUeqTHKJy1hbgtq9eiQGEKXkb8bxMFGToYSCcfjZr4jc/uQo4vFuKfiB93xSUy0
B3o0oYYE3qAS/9q3yd0J1K2ddqeupyk4oawqlME6Hrv/ipzdI7+luyTuI6De8cUh
w5JPYCV2/mFvY+GAIWCan9s+wtOFadG4eWb+6H+Tj9Ahe4/SyHxLTmyd3FxVYLXL
sV/gFvqN4OXP8bxYz+UuCeBsqTACo4wzQrj6MY8+/fesT8xLW4TCIBHexPEWvB94
egei9xxP+ir5NSOcdlJK9JEmR9Qb8WxlSzvEY8L1Y5yZGvtnKK2/ORRNK2Ya3aDd
ZTlZwAR1RIzMmnGbF+HyBO/W2xyMe+ck9qv3PSQmCr6irwIypN16+H0oJlu5S0oc
+HYwgXJWpwN28utPx2+77O4YDkt6KavMzw2+j0gHMBdFmnneQbgEWB86025JjCQ5
n6QmxLLSBNeshwCY7m4vxvNFqy9WROm7gC6/NaoJZ8ESCD+AD2slhAAewiBNeBhe
do5UpPa/FQhHo4+74o8d64iESwW/CIBB4+FcZCcNS4p3w2nG7S2dVi1x6ADFML30
sgWd+qG/UZuIwPfIiFTnibAtSJ0Uf1fAQATn2dLOyhmPo0tEJjUiLqovF6qfa5sp
J5QBA/OffwHihMpST05DSgKWRTBoDSwg+7P9AItRG48R0JOCOcMRVPQqXwt2Shcu
VigXtzBp0xdSE7nokmIg3r/zNnRm7mn3r8sGXrOfIHfUM/1CrbxH/9k/1Ml/IsH6
gV2Uxe5OqeA8wThba4DAnPoIc/Ti4WLCEO06ONU1DmFFjEz+8UWC3SOIBwa1cEzY
93kCLtFSSkVhy2liO6Zl/HNxhTOs7T1tQAgU2O0mWNp2OAf3uLRf7SXREJzxf1OM
sLLNhBtMBfFvOHwzsrpOprmZE1FbrUe9RWl/P9kd+iyYlAkAu0IvwEBhVQPA5Gec
w82gBKRncdtI/JKVB2LtVziOs7tjlf8wFWlhJhJcxcBjpblkWrKNcCaVihKjDElu
NlGzpWYzx6K7YUgoz4uuz7yEU2X0C2VES6TqimQONoF5iqlVTnrR6C2FJuJ23h0f
i9FaTfgaUzVdgFD9pTH/1pf64QIVGRBcCHXrIW2+mk4po4J+7jBfAkxXpTMmlDuh
B8CDEoDpLu1V9aJaKvTVBiOyGm0Ej4EFKupQM018J+2UI+PE/bzilePQD1TsALXb
mAU2+Pc4hmnpQ0JhIQ16kVrhQUXcxx8jXtF0RsQIl5XZKzzty1W2LJAgXjgrj3U5
pcGyIAcLrXwDfdxhJJbg7l+NaEx3XeQ1YhdABYaAYIQaVLyKA/3YDzPwenIAnRdE
yFCA5HgsMkIjwFfvgUn299x//X/wAVXEcZ0Ct24V609XvDflYIKOiJJjMffVdr43
7XXNYBh05lbbW1GHWnRiTQh/BLpKutN5F0XkW8nYxuvVTLMs6U26ylbwzbqf6uur
TQkgrDIWKnxIyXBG1TAj/AdtW+r9mVXwj7sw7qj6ZKKEhF7kNqpeZ/e5LDAR1N+R
fHpqb0yIv2aZGzAZada1BBtCjUlFXyHoHwSANDbWBtbTUhgPUn3umAkkMrPvwzbC
JpylEw3XF7K0IWB8wmZJE+R34jBJrSWfEjMmzemQXhanqHKMHl1Ry5DLhLJ/pcdJ
o4oaGdXqiZ6zZstbM3UuLsnfpqgVZkxK3zQTpzC9z7AuIufWQKsLahBFJnPuVCla
zR7RerUtzBsa3T0eQqsKQegI4pNnSvyOtLR/C2yyBqW5CNoXzJLvXmmxl+NSnq4u
xhHDbEbUpLJw8Oqrrs+g/XtVvncVFmazGUmoZlePs2c+Vm+hF43vF1qu4z90y5rO
spN6Uf9T+sSY5RkKT0iIWtilSLtzMtv50awGoXyI0Twt6xlLGqSi7RoBUODKyhJw
iJByJtXMXDBWCjF8D84iT/vTOf6wvE/Y3Ipl575hahA9J9otQmZRoG+RCuSR+4LJ
U7F9r2WXjFUU8bVje5VtA3GFtSiWM+U6/51jX4kkiGr19a2q0RM2z9RiU5RKSxmE
pfajjV8SyObMmQcxMNcgQvWU6zGMUDRue1iKe10qZmi+yu4rx2w/4Uk+UzrpJKo/
5qR5thJiGJEoq00t+tu03HJMQ3DEXPH+56bbvLTSw5T9Rw7n2n0nPt8L43cjx/XT
FcA0IdIwLT0ZUajZcH5cbwl9qxDOpYGvgaGjHO/nhWXu3haukBkPiCpw+I1k0we2
7UJ3mOQLgv7xLRb2AL3ENnqQ1iCbx1AUUmtoJw4XffGp24aCuVWCnFtTL1WG7LOZ
oovS6GT0mCnAEAJJqMKN2ntYdhsQrFzTYSyXAHiXRwFowzqKWyyShNhVuOO59TpF
WU4X7Xr/1n8O8UK2YllyKGDNYTz8gN6gIPi1XgG21NiciNOl6GLY6sNvVicGs3PU
jRfVGshHp+RxiEAct1nYjVV7FzxHXnOKQHCNI6ebbEcFobZWO4X+iCr4IckQnrMt
WTOo7cD9D9oskTlsM/g43f02pklKGaVeL4anSg20GV9CT+z9dmZoD5vsYBMsvoT6
HgvfqemTJGhw6FTyc6u+EtGRYhIWVxmQuJXeHCi5iP1mmp1naQcVVNJonppG7wal
caBZQNUqQAse2LaeFf0BtrZSI5vdMJ4BAsUtd4AbXcS52M95bu8+rpL0mDeVX2Vi
irix6v6cgqzbUPr1D17hz+E+g5rGx8lFtXI4iZiMmPoctWEj6h04YC6W+rpM29Fm
a8IMPKRYjchWmHdYhEPiWU+DAFd1QptK6PK0azFKgL42ypXBTlhlhMZ7d3rmO4Od
gwL9Y4NQFy/Sw35mMCLxKRE8SCCc54DrZ7Lw4uSkolPF4PEktgmK/jA2e5eJStl/
V7l9DfYO9zyR7vun9TvJYNT04dB1vKTUaI9lo47X+rt/C0qed2kED/y97zvTG/AY
3KRAsIlw74qfYMpx+7+Qt6TJaZ/oVJNxdwTX/PmOxUokBdjYbwEd9fTCbXazi7X2
Ix3ts5LFJHU/ruAF+Gu55eb5QlnJLIIRD5p9MspGli4CSJjdgb5GH+ROkuQQNLKz
og4o4KiL55Z2QeE9Zs3mqRoWwdfQ4JkaqAumy+/zr+ahf6tFwjRYzZlbGrmOGJzi
QOPJ8QDS+/W2+FJc1g2w902QpaLRmh0J3TXGajWQw0T3UMQvB0I0jbnkO0O8tR13
ci7X8oSLLPWKrYlJ9wk04BdZw4nKogDxJ8STtXi/Xu7YN1EMKDVC+1d3KfpMW7fH
JGotE41KrxQMrfyNcdm9X5h6JLmS3RQxWE9RRRo3jEiDwSO0UBp4YTnlyYKF+fPa
qPMCLiR2wHvHoW4qZahAJ67NkuK2bLnbgwHxoVgwKYJ1MkjUMvTSh79X7YgH+UpA
AlrBDjV/V0jJV7IYXFAlPQk6/1Hcpya5VRDrbURQuzpDDEc1d1giuK1WgA2WnvkF
3O6GLtTka9sRl4sq/VYnyuqfjIscVJohvVhUJurj0d/8McIgPo58/UCTCZ5svkit
u724pLSjF5sosUgE5cZnygYQyohvdoiWaFGQ5iWOz+bKoMyp86/pxhHsT1bPS75e
RhYGqnrG5QbsnW1W9A4k811f/w7LXOY2eR/VHamopX3KaEQjRByQkFdHsip3cMc6
I1vUJo+qeWkDoU8wdwTOsudmGQ7gFUFmZjkxvjlGJ7ymUi+OIVn1CtsXgPYnxP65
uRHMyiJShbKrwBcUAeFKovtv7LBTUtM8OFIuKez5oCWtcDpb8Kb1JDQUK2Bvabie
dxUy+oDBMJFbHk24YPTbYOwDo5wQVqeBkNYC2Enac7AOO4qBXnOQrS8J5TdRx4xT
AOCX5GA3hytvZIZFck4yP9bS1iAxz7YEMubkSjCax4udL6P3joQQoSEoIvehXIgu
eyP4cY7SM4S6Pbc4R76YLmli4wLp131YmN1myh3Y3KtUO5rtNcDFLAtK/zDym9RX
qpWnYJig4UDQ9ZKDdF40iUdlO8d65FifbB2f6xTccjyo7VGSDwPhdnvJj/YeH4Iz
zQrlY8SmwdVdLzDk5t3buTgnEDwIV0a56qJqo1PJYpPZNbCKQHqiDLlPdcZ2GjSU
E4nmuj3DLH4zaaAtc7JtSvSXuCfcaHTHYF7GVAODX8fB1rA4pgy4p5AOd69jnLA9
Z3Bju0aZAOFGO6Zap96Snwj6hTOBK8lY3UIrcewWkpW9nfKDUeclxxR1Q10cWWPp
vlgTUl6LP1oUKNSugbQYxRrEft5sFQRGb1hMrR3DJoj3YCwxAEIHBh5Y27Hc0x7/
Fke7ep/vIffr7qJc9kZ6H1sFDRwTeaaQzpcbAp29XronkZ3HLJsyZIJZvO9RC6yp
ZaeBPUEAg7R0rteFAMESV8fhrqmWKVICNfoou810XvfJtbUoD7uQI9YtWpbU3+Mu
ynJqJOa+8bMQwMNGRZPNQLN0oHjgmHz0MmWjP6JSSBNR5YbwkwqiElt4m+NKuOr+
pM9v9NbcA4X19wAOsfsJ+dhSJIEKZs0bdfcJ55dSSTIaQHTTlFNYDsJWRdF/8/cg
fu4KOp/rxk1fZGymj3/LoUKvQk2WDFqZ6qsLZ9OCTKKWVnrpqvWu8HEkATmi/x1N
g2JfWdEt/lsGEtcw/3tmqEG+8PqrNWO+spGl3pyh09o8aeshEdCyjFnxhfAyeQNV
aqJptw5cAOVLjA6bp7srr3GljSVr4Qh1zO2Zjz5/7foF8BN18nJBvLEs1h2x+rI1
cFtii5LxD+HoFm5eUBEb74x9iZJeT4DuETb8nNoSp4An3P5NDC+DAiFk0gMs3Wzj
07mq43sPvITq3wXiTJz3lMPozLfH/QYTJaBCMCucWjTVy4pqJ+m8QC577xlSSafU
BYVJvEU66HxLSGzee6RXHZ3PC+ngFfOh9DHEuFLUyv8kxphcHsvdsx8EQmWcXJdY
SzY8awSBPV5Ua1CBYG2flefOgu2cPq7bW7/0tobNxNwDkSOZAQa3Ok9yEbeZhNSi
RHQJUPrZ8f69Su0bUCeE0/WjN6ar5/hbb4fYrEDcMCdsJDaXbIj7OZE4SvWkDap9
zQ8pcGKxnKOA1FNsxgZDvA25HSZU/Lxv37yjtea4ThtX6aBibq7s/O8rHQTTuz/o
mai/MiUSaUbMdU6opSL69Fa+o4LCD2mJrzsJdSkex6H7BYE158sy0EzBlRiDlyKd
P9SM24F1qIcCtC4Z1E+2uAG454x1kmQ0Nz4BC8PeRpkK1jQuF+wYxb2T738W/4iN
Z3oasBgiRzpuGegnhmUZfEuEfuj5MCYfPRAPWS81Z0zqfmYYf/8z1lVDhx/f7sEO
tEHcHXvV5zeDByeJciYmiR9S9EWLJZcunbeGfwp5hfs21s2gtQmcLGIMwl3amH4/
NlsxX9JZ5v4oF6VJwIBSp0dnbQLpRP5w9SEW86snf6wxGVNNz3UQ8dh1hO4/d85G
dA4GJaOk8iQA5R2YAbTO9hT/dTJB9Md9QcEsIuAmEF5F6h9UUM3xoWoK9XdaV6Vv
HXQGuKv4OIguOeYKFuAAkByCJ5Oltp2jo4ZcWbWg+vROzVAZ6QHvJV/Om/R1H+aA
Asbxmr4elv7k2Ph9GkSyvxJutvtPUSAxzayAGh14CUc87+dTFoCydCaBaOP7JLq4
aC3fOm98qexxXK0UdCYfGPBZ0ssKDI/EMzM1rs4JcUBqAVxHdok0swxLF7lWygP+
LlT4Jeo4zCBTwhG5FOKw64U3YcCUYNZ9yUE5qGhdIFGln4Vwjoers4Y/TLD3hMs1
Pt/+KHFmBeqhB7rbbAUySG5llvRgs5VPPRnxluZXomzKJXhkzAaHlq+K1sCRvU/5
vBXQToyg0t/Jq6JzelFFwzPkufebytVaLInSwb8OZBGtVRX5yHNdymkBjknhF2fH
M9H5mWgwOQps4t1NSNicxoQ4cX6mN70Rb1ElS7e3aNfm9OEDlnXCU2P5tBM72Ssp
bRcCPN4kE7ASU6YtjmfMK+dFbTKF3HR8SAgQIE9EPCsLdSV2sxQw7E98L4/uKsYf
CbFNozfSC3kiS25OC1WfbtIWjUDbLf591+OWhfAq4U4qaOea7BO6URfBr1f9/Fx/
vHwSI675WfAuai/hRtGRF62L9RuazkbqpiDsUNYEObq+NiCihS0rmGhW2pc+sqgT
ahDswLjunLpsMgJra5K2KWMPIVbs4/dJNauopgELmFOXGLcETne+zh+Veus/tpqa
56NbLTjoah2UfUA7g3OS963SGElzzaQ1asadAi4byB3Ehtytmv+d0+vjI/Nngby7
DfcprvgcsysyOOvpGq8i5dNr5hrrV/yhHjvEfCasrCxYtCEQcModwY0nWRJOICV2
Yeo+Ar4XCnYfZrnEamci3Wb8TokxfnlWvKBYhLSUIdT0JjyFLH4PjDdkGqnIM84Z
kWl/EA/4MN2f6yFBQmsPAKrLNcS3YMpYPTN1jnGLtd8sD8b5I+b/Jl26Y16/8H6V
cs6IfXWE/JNyXPG1+Q+UW9FTwtRkWQTvmw5d8+TunldgD3YQadAJN8wygvobo86T
JwQZlcp4A7zo/ANgNGZVX0I+mkjxNwYHDTKFSszo8hyTRwiZ/GRvwD5FmGjm86wI
cEMu33thXJPU7ySWHKbRx12tvx8fwiScu/Fg0602fa5Gt8D7Aq68IWeOnzLjwGSJ
ueCMPPXAw3uZ4YVgYrt9zHsmcni7J4jYXmc6BjH/rulWpQJVLKaKKQvqA39543MR
ZucZ3O9+gYjNKrkVyfmpb9VZPI2QYHu69p66KCU4Vms0iebOHSU905KOil6fs9mi
Xhep+4BGyx4wb54/NkPeWA+iNTci0xfvoaKeQl38YY354z3Xzkk4IGBactMbO30t
i27KeXSJBUcjZ/DagmtVY4Sxdpj+7eVM2cbnVh+3GTLeynCfZx9ukwF6YMf1+Boo
B7dYlxi6os2PuepC7OzwM8YCrbjteAnyKmc9C4xNMD5A4leuC/WdptWOutNbNNLx
hT7xHx33cqoBnxP8oRz8lrlSeThC1mp8SbDiR1aYHajR+5jltRgueGs9zuOul0ZT
t2aHS1gmSN3XlHWKuX/Og0r1gIJfsdxk1m/qbCNe10E0M1xwWyRrjHBznHZCE9x+
+2KHTknef7aB7Fvep6Lk48xKfjx0DQE+FxZEJgKJG4Q2a2afqTBtV44n+pSVzf3i
lVzW6qprjDZ/YSNu/92i+CvmN9P4c0BwwsRHPmgsw7oxm/q8/D+GR4gTRfYRPuiw
OnItUSA+Nihi0vx6FiUHRWW+RsZ4M4WSqaVSMeUISFjIB4tuN+aJSSCfNnqQA4kN
FM7G8EZPZBoPDM20ISXhSW/u6w20jlih7LxeXVxNq+e58RYcrG0hPffp1+lQsGgO
dbzuZB6xuGQqbNZRPYZKxpahrq13Z4Yd/oC0JqZ/hhTw5vB0lNC31TuGcuA5y5DM
iXopsjNuUYLVBMjn77xmqvAZtbC8QidvgYACDlilVrXiD1ZugtmfwguQrp5YJ9Ya
jCixffGZPot9ghy93QgLwViuVbmHVmexKFfL5/qFN7nO/t1h3W+RhCFibiNxVY9W
3yOGSj6/q8uTDvFLFW575nSC48Kzl7m3oXJdGs20S4uOH9fo+PhoKhb1fgeM4G/c
124TtXjdIBMRKJU2hnTADXbZBhZV7xYGi+sg38ObeUleBp2NEhNN9ye1OyGdI26R
mP5dCV1fcltQPTWYMW3uSCBgVnqX1XK3V4EjW/X+TGrYXPeT83iy8foSGWMMDNLP
Fx7IamPtZt+QBeF41EF/vBEU4kDUEDH0rdRcl6Ha+qeJVLp4NCtWYet0QkaNIETs
4aQO4BX5QBWIEmzlsh1eoNE8LuBs218vHwfzQpaMgrAw3O+wdJ+SaF6EbBMq+7pv
IfEqrkFzAZWUdOJ7mKDFl3Li707tzj6eoMvloyBjS67vHByzSYdZabtkVfcrqBpb
n90JzSCL1zyHnH3Fb3RTQvU/8ZKIGhCKuJEpHwXiK9Ao86wc7/IT1+K2CscgTXMA
CRsCLTib0ztFJTBEvVK5wGj7j586rVhsvotKHxZDTvg6xnKaDs8OW2UQfv+Cm9ud
7u2dbQtuzhIGONE78eOauZ+7nEup/F55yNoSLNrDbtHrIYGQx/VNbYHbCQRfbF7I
PqZijvyBGtdO2fRecQ0t14M0ldukoXdL+ck8+sIzcrCs6BJKR8PDdr5TnPDKsFnY
B+lJb/W14sro009WVXv9nX5HyCAol4sWSYXTc1NNRQ+VI2plczdDzdIoY3VQLuu+
z9JmaMVebuOzCBYzb40s79uj6scwUlXffHQCgniXq+XNwE77vj1NjHcQPEjDlRep
jjozmdWtpLJbQr3sQJ9cYSCkIr3uZDx/38UflQEHEvBACWz7vFHb/GXtbj/MAGx9
HQKwIAiTNblfO7JR3zKOipWKEXbqGYxaoiplmrAHGtH5f2F4BujpZkCuicWO5upd
eK0wstWUaTF6c0nbBQCAptMOKbPcPuT719e0TN3fy/6b+/hQU9LFP9os/8BzENnJ
B5xlY5TY5C8iQTD5LwGJSnKx7n9eHn3HGMd7B3sB8fYCCdAJGiwptvsr+VJochhe
MvTihSOc14m4U+dMTYYy+Lu86iC5gZvYjeMF2HfzGqYQfFwM3Tv7iqUrWS7z5FiM
bVoeFgliChaiRZqzOa9LiwtZAk5cujJYIEmonT8iXdCOH3/2pW8AVs6VVDTZ0FYX
gCfhZnYSK7mj/x6BxwNdxlHAN3IoA41quSivtXcBP/DJEbkeWriVf4WftVM9wcRE
TrcZ3TAtQmBIX3fvKnsn7MY84GU0GSzgX4UoKGv7TsBxIGAOR8BhaALRXYmCa+4J
owxGSv9prY6+/s49+CWJ+lVy7m1jTlHXVIbnEM5nbTMgQl6szMqkY3QGmwP3KRja
JV4mymi4rnbj9S/2vZBDugXOL7/Px75C24CBEu/FmSZeH5vnn3CnkPFZrEsqGgfz
cghybnJZtLXWm4VXEvXBmjQKWYjNG780HOmYgfJ8RllD5IHSWKBJIgGWcT9xl2IX
wOmN4nF6NOZImU2fThz4CY87Lzjs0UmusdyerP3SlnW1OhoFQNJvlibegKHZ6W9U
oBq5bORt3pD2yRtItjeq0N6CKYSKXy/MDa5U5JIqelpcii6T4gXetEWrcWX5BmkV
zzoRCEjLR0WgkGLV84K8bYU+ek/+iEzbN/CVbLvrmy8fCg1OyadzGo49Kb5QOng1
nRFpnWU1jdB/nyymRGziGTKtCSHfZyhc4p3YTFMD5KkI0vKS3KeNGT3twwqlbnF8
XDj0axKUtRkQy3EPhi33Gde+AC2lkLmaAyMH0Bl6J6SwOPVYkUXZVNhLTvBDVpo4
olWFzec8ulyWhbWm+jaqJ2XrWnK4rKwp2Jn0BLM8pK08TwQkuR54ED9LNxn0tImg
aW/pXlbZDJn42kZNggvgk8L1KTOZelim/ooMzkP4mKQ/OBtHRP8ZHAv3k0JCmIKZ
Z4eQSFvBW0zc4LZffR0tcgEd8NsXG44MvsdXc5rpTHeLMZNX/i00YYzhgpql9Ibb
II4qo5tI0KEdgk0DsWqO0WYyQhKc1TA0sdKt0sE/RWuyzYlMUtBXdqbsH/ArjAlo
aBqI33TJtoZLQa2/uiPwTY0Bm6f1K4NaIWyOx4H90PiKDrQgsZZWVt9tAuS7iJ9v
qTAePLLie+h56uUL1XoxzA1zNl8mnoDP8BejL+HCb7mmrkSoSFPu9tyNOJHhDuKY
mJ0ACcJuErjlloBuwPmRXMnmptWDxrxfPOvS/wk4yF/JpY28tFxah4eBCL39cxYi
L6BKsa1lgm4OBQHgsk9BQy9xiEofLXL8UPqPSRd7hJ7vZTkN9itWIZyMQP5EodOO
b+oKoTrtOmssYjvej3PF/eWp6VnIfDdQVst7ZiYq4e81PkcXy25e530pnSfMsfoC
K9OzWIJ9Fa/A3taGVbt8jWao73h4lE3KxtlLqjDPUb1lDWdlneQr0agtUjhqzFfR
Rcf7GH21ztOXihBXOUeCHvnnVDULPXhoINCRKI/EnZXJmwm9AB5PgJba2iP9R6q0
9QbbFVyetoWdyDgPe3IHEHCmPV+SIueuw/R8RyVnWSrH+a8+exbzzE/wTq4eYgmq
Jr9FDSHFw35DOCiITvYg0tDfYq8zs817TPVjfmp3NO7vpETNTaD85uVqUwfhvtnc
2zAxREONclaP9XzGD8hgN9+jTukSUKNuXFV7on8kco7XhtEg5k+ZOPIcWbSqQmC7
aAvWCdcL11Q21FeYwDLXSisX/kJCDvpNePwIJxo85BUgPqoj/0ypiE7r7jpaO7Lz
9u30lwQ3F64+JV7PCI1Zwlx7vZ/JjxKFIYDd8AwAJeZ42IvGRI8kcFh2ccH4iqok
NQLHLtzl4yaVAMmcDvZJQUl1aPIbs23CJTR64IWaqk5QZkbWtQvZ/ud0Y7h3x5BA
Zg1QXVq300yBIMlAk6EY3+7dD9zPGUB0l45q9Y3aNh0QmcRa6co5q9wDByKnx8DC
EqDMFOldsyV7+uYWss/g90buo5ZQwwnbqwbmYqN3Vl8bewLTiYRU61jd8D2C+OGR
fzVBv9HTnmo0SXqYXKiweiRTA3VYCGCjBRMoAOqoHTRNAXZFpAeahMOYzePGFvSP
WhEmXXR9KCF5xtdyEQs+JjSb8ORuy4Z0LoWeESUgMaVIMykxJ1GZ656SZmfk9eLH
oYyp4w2o6RNsQ6Vdq5CSOAuAQ8udkk787HM9eqHF35NYZehTWQbYrFO/WRNDP7aS
23AmhSQOh+3/gWshKQFK59prEKWD1bhzE6Q6uzLcaGvOltgq4hWrl1hnlJX7HeOJ
tIa/B1mwEFskqDrSoKgcl6SZ5SqTuHQCHVVyRLWZ/S2m2ryncro6dYQUWwOgHXQA
yrscKCQ2Tb2r0TsxiOV7PBzYj9IAoMh+Iauk9Ux4Hkex2n6z4eN20AAiH9rW7v/D
BCEDescLMWaTy77ZfOcWx3Sl5F248hKlK2X5qSDEEycDpdCH/Odfr4OpIHOmVm4R
LBS204LjAAGIou9dHf2YBY3PRPKq0FQdW0Sfol01pCofFsPBU7LQ6hs686knx6/e
0q1oQrydp6qU4ZnUpik9MOdU7pPAh2jVgHwT/MWFAStxBuTsmWvIOGw+XgjwmLu9
TPYa5SJioDG8CT4T+Cf/NuV9zaECiaqX7kB+qApSZf32fJ2qDF7X9eWp7f90P1Tj
InxTc8CNxLURTwO/d/rBv+01Em6I0q3lVUfrhL2iMe9g0RQ+7wJooQ5SwLqba9hm
HzR+Pgbn2AzCDM9JlYbEaNc+C27MF+3gGrSBnJ/vB5WA8oiA8VhOYAkBwObu/yhN
ASxZPREv3EsInfeKN2bAvQR2j7kT3dOmkUcvnBEnmYjZFm1o+P1/X+Mz4pjftGv0
gqdg9aQcmPyJSXVRzpfhRxxEYfGXgu96UKkkxjWVh7dIuFGsA8d5UQRiygkzZBjr
SLIRjhz0pswv3N9B4WAJH1qPB9JHcC+MSIayEkgK9fsAk6k0ZxFxkGMeb8bnmvEP
1YcExzXqBegp0n7KcNE8hPfP9sclV9EjlNCmZG8i7sY3hILACPGjLcISjRdiWMdm
kLkGZXf361r0eQHqhAtedJiJUg61GfU8T//sU3C7zMq8H9LZvHJ3o7gVSN2zhlQA
XR1WfUo2ZCiYFkZNnPNi4O6zpRyLTYREZX/pvmY5M0b1HDaztBjdLmxn8Rbf3MqA
U+Cj3l1Rs4OIX83tv70tmZPpmUnWsjJTx75/oZ4N2f7Q55h14XBir+QqZIPbqG9E
zjLueNpOqAnCkdoDqhkkPC6H29ohTqsJIeX3P/Srze4LpiwASRHA79nWWQ5dDogI
p7NDgorCnCKWSk6OOCRNS3wJGqzSoTwXg6cg3VCPZKVOjDRsVeRsi7wYIFLA7wh6
zsUkhH8+F1RkagiYvVGFu2Ac69vsT15T1tjr8kDR4CKwcaa+piQdgccyBdzqCcaX
ds7nsGjU818i+ZDoBwaZWsQWOKxKGdpNazQ3kFrebeEwCvvw6N/N3/DZAmFYY/Do
ev/7AT/wHoUbZ1dt2j9SY1zGP4bPTT2FtiO76e/v5/UPzDTLfLGxPxK919dC5TQO
7736bLlGLndYGVi3faPOTcCJGfHKQzFwGBwm4PfXe3/rVEXAu1tExKau2morT0aE
QSFlW3YXJOBwVId4/xYGR5Dq+/XZx0v2lWgLX6acD6lP0/ZPUrkI/qGrP8ccJQtI
koBAPU7Sgnb1mSmM4XzZiaFQCqaVffvS2okcMySO5MylXpm4PBoiE5acb70vcXVE
f2g9pubLYlnrWDTn+Or6EPAYT8uiBywGHqsx9jtWbN7kx/SUhm+hy+j0F5z+07Nh
lb7Z7sZaFoDxgbXfjETcHdIdiLRsWY+fBXqnAlQ6a7fZGuVyxIfQf5hHVwOXi8+i
obFSfzG8lplfWZpm4g1rcK0odxsNQvqtQ2VfjWLUy3UsbYViclfINbJLBzm0J1EZ
dLlWM1uIjs34waBHzyVvfar7AQaKknl4PtBsRjTNGOUxWIpcNDfiSDhWAGJ2uf6W
n0OCINFz5yk54HF2iS03CrK8Fevo1QQ5rLQ0nt9GhuqUKXc87mx6O/VYLNbHZv9X
61wRt3ukG4JJyCxSSGaZosLoaDw9yIybHKeD1kfiAbEWWQAwogTSMhZ1DzlBv4yR
G8lfsApZwPRFHWsRo1LeEMB49F//jHnlYItyM+KewQc9wOzhN1CkjJiaTI9PktO1
XE1BRSJTDOJoJ+s0NJAibwYe7MlONFsL79ob4jTzWcPEv6FKtxJLFzMtjpUsv22v
QUKSokY5k8QjSjkjYyWfgYx/HxsjXYWJrzhaPJefq7ACyYxs+5j1Basig4k2JSOV
oIjV622OpaIUqA17BFiPGMNp4fUUoTvbIBna+UjHkAHZL3iG05HcMM4asinYOaRj
PeuQh0coTyPS0X4GV9YPZBQSiTRN6aHGJYSjTIUOGWJKTJrYBvUSSRjC8AujCzmw
04Kg5XeW9Sfl99eo3lVpeQFxy5deNBX+nELIZ/WBsgUvOu/hlVpR5j2++GnMl6cn
hz7xPnEwGcAorPP9EtplPD0jh71ODHkgLxone39DdzfniYzogwgT/LWaVyU0Ja5c
84vCjI6EgwlCzafhg9cHcchmdMHEa2eWOJw5zQaySqCgG8euLSnU9Y+ENkiGCNWG
hBP5rpBitic+8cgowTfGWiPfQVXhz70ATGRg1Rb94xGrb22XemHsS2ZZGQ3c6wdn
VWmGTsMSKR+7yv3Y9KAW/Z8pBtOjeJl6VXv7iwrphETmB8GoPISZs7xMGxwBsslp
i360ag3sd/42niOsnhPQGkgpD/PnXLatrWYvq8gFoaUvzvRdICTDzRPBTqr7iJDE
QvEwKxe343n8i3FZ1X9IimVAfo2cLR75BfgRnQYFB5F66iWrlQVRaMGnUSzrqVTb
ke4E6XEUAIJCPYC7TNf1yDUfpCb/eeNVZu8vfzk3Pgr9QHWSgOVSPlYKtQ7CCdZB
qtZK/JEXnGI+WhZbR8qFQWhGYOEYurahCfjI3ujyd4MRXHr7PnpWhimllvSodIjp
kKO5Rwvx7a2or8P76OUICWdPVpRpAavGZC9OOyVBAq9CnrSIBGthbXqyV4K6EGyH
nQmUZu7NOskczDWhyxtgZADRhC0oUaHBV4hlM7Av62rS2vjUKZ+TDWHrzIisbXFJ
mv2IGWeQW/UkcJlUGogha+5bTLWE0UjYgpTrNTCT4RCdj73wsHp+TItO3ytf+EOv
6FmXZWsPSZi7zKbyH+kp0G28lEeE60o0kiXWK1LewMw1m1x6MMJlIi2YhrTNaEdu
3ExtuYPp6mnSDjQouOUa0ZaJLT8zUQk+CJR+mjduFkhOAP6MlrOV8GG5NPEH/svD
UD5xiNU7IiOO0jP0X+PpLNj0IuYVtiVxvt/V0q0lO/0+l+3djXba/GHFKZ1WoVHW
puNqLB7w+xYbUjJZIOiRsNQ8xXFCpweYdASxzqNPUFwXCri8uOD5e3rnoZCb5LKz
YlSMXnxN3RwV590L6dbmJs0E7Sy/Hak+lpIhMwYBSyUwuGYl1EH8aRW2oP7kplzu
VSlE8JCuG/8WQ049BfgUG7h4tVYtd3lVIWAu5Mc8PDNBVay1GJuLBhWmprAK+D7f
VfXhk4emu4lAlpTM/ASbTB0a4/x4ZBXs6AR2DbxnQrAH1XogMef0LxYwvvIXHQYR
h4nwFq+1Z2oJ8VoaLxcxQHD7p3Wh8GhmcYt3f+Aeyn/MUe03jQGUQp92y6xb7wER
qNf1qjuxHNHj70gGX3PH534FWgUGGIiH+hh8glfsmeML/mrw5iTYyylTewsMXuei
tcIPu4bevuEtAdV3B++Ncl2TNVAJPRBDUpsAYzbhH0HsU5npEKYfxeqSVKuoKZko
Eh+Y7qsuye24HM97L4b1C6k4G99cBvmRDcufL36eiNEN6rOlW+m1xrRMCXAsBAHK
vRZ6UlUp09xWC/B41gIRh6QVw4e+PdZlIVUoOGz5YT9a0DJ+zAnqUbpzdFOC+J73
6sApcx+l5bfjS5CRfV77oxqZBohe1YEdZv7EYZTjghKT/3mq+CuwTdhEZSLWtlRy
oA4cFij3rQMKBsalDMvRQOXfp3CStVt3lZlehFuxEieuI0HTeNWT5iCmY8H4cakz
nwM16JAT/rwvp2TlADn+qJHrVHKSAI1m5sjsV9HR3CxkTL2g9P6Nx+h/iMubJD7z
Ji8RRQwIz6M+hpIAtoRc6L2utHlFMyuDOB8Ofd/Tv4QNQwlCOtz2nmCi8Oglaiti
aG92osqDCKgw/1KeTWuDA1BEUepOd/6O0Ogo4SOx5i4JEVE+mFcmgyPG6vh/IG6l
QTVx4SdM/+2GwLpcPImc04RL80OfUu4WvO63F1LDoa0oJ2MN0ALdqeYUdgSZ9m2A
WDumZuvO5hSMgBWjv4cVaqQ2cT7jRoN7AJg45PFpGJDSFfKmBVCYye+Ff0WxPNR7
68ePG3uGEpAbYW7jErTX3Sqf3kasSD9BuyesU/OCG8gt3MCFNrHgHROOTd+ldTXO
NyyELdpwnf7A72jrUNiwy8EUEoO+xOIFBntY5ToQ6IC1bZh9mn8Ot7i3lk1XWcVl
KoIdUhQP/je6zWFxhpSn0NQrqe3Y8DPPSegbSlkGZPRKqzbS6K9qoU0FjMRHrgOp
wukYki5uTKvRB5v8XgE/RJz9+f6PE6pCXO2DIpzvL10GrN71krmbH/vm/BhWvmEg
J1tjG4xqVwLH2AN26Cnm+gi6ghK6T7JTS6uC7ivfchPKrP1oKGabIqlBIZm8Y8ys
rq5rUDHauTXlyA+azdBxWFkkwJeGXp5rcvI4riQM/EBM9w354J/D+wdoZQBlWqMo
PzzehPPn6qm4AeJ7zhYqScMW26qXBDFOfBGtuyJV7XSR9II7w81ryeLjKxVC+QZ3
YGkA0ptgbMGNdhV/akmrJjkq95Wajf13SsHHt9gYJyj/F770gAp6ocNJa9KElaJP
vZdnVxV4SBNYYAf9KaGhrkAKNHpVNZ6ek99lTdXrfKVcjQck4cIGts60f0UrfqP5
gqauhcS3LSkM9k233fhPryvUTQ5xzSPK7LsZmh371x2WHT6NDjEFt+ZBZUezzLTz
rkFMxQ08ZsI5jHRKgSVofPE3C0C64p4imNJlUFzgYmzYrAQCRWRKh3PCj9DSjPoV
BsvMlS/e06xurhYzAT24XcpFU1xp3iw1aGtZey5DkGz7efla+OV9yz2JDDIOdCeT
qXNXLPmQGpDt2XDEm/CPsbFfQ8A00k0A4m91ReFYeKG7uMHvGVqg21MFuJLMOKwm
kxKQGsaUR3sRGD7rDOKxhymbEF6R4cc+vYqV6eQwfRPjZbIarO1HbfONbyZYKxfk
8eNl7/IDsRJ49taa0HEIdTWSolonYUvdf8bYE+6fVr0AV+3sZ7CBgK189cojEgm+
/+o1RSv471lBprXdGFfNxuKrH44rwZrVs/yNDILRWRMm9w+n3KptenmoIAXwbXdW
RXYydO0Djct/W6hM90GfMBHeLBiWaCgbDWIBeNMmLAnknqukV+B65kTmRxQQn7v/
M+z4Wo0HP9c7ojkAODcY8YHmVZMSLs00kGAXbxahjeHnwrXziCluOg6ckQBV02bU
hDvz3svcbxm/rPLUVUyGsTEzOH2Zk3Wn0jS5oLUywLK8aTI+DyDlIcZMQj1QRFPw
yoIW6K+HGWPEBjeqNEv+ZGsPxUlNMXt7pXsBE8JKh/vRvGf9O5JiUiiR/9uzoGQ2
XMhlnLXr7SHAlTn4+iAt2bNTSuaT52R2X8hqOlADdQmIIJPAuRCAIJWpywZJz54U
m+X8toeSWbkKIOeC3iRiKONR+FaadTY9/LFaXa+uBcvwESPeLC7nuHh9CnV8NcBw
1ygsfFBA4RuMVwQGAgLikKmJJDVkr4uPstr12bynoleXCgE7HxEsYKC5ftkPDzuB
MX+b2MbLoZSjxYvhtRBc7GvVKoPfMu2mwVUxOY5jcGAK0ElxLcDdRlihCPLFQpEJ
u4xTgVeeSlw4YpwF5FfwQOX9o1VDxqf3FLJCiOLE8g1B4eLfzSzQqCcs1lNDSFxJ
k/4z+v3ai1tyl6uNqgh0poAstHTwQPpNXdTRVmuDzQFJXDnzg2LrgF06YwHX3cV8
Nq6gdckYE2cYj8bMgs49W4Qni8FzyoTmyjnlox3W7EuXSaSqWNUZh9nXqhv/fRpS
7fBwP42+BbmuqBfM3GXqk0dcPMTg/WjCLSgkN7P7egi6R7G59ZbPSFc+tsw8esb8
vLlLimO74LnqqLICy3WnBb9G7vB5i4lGU+p1vifA9/LOYhrs2+V6c/JMMpYjDcDp
HHX5wP5xSJ00bAGUnSbKbK+miPTS/09FVvTnvR4XtboD068lG1/BSbV4sDvhcEFx
vnUMLEyaJdyy1vN4cdFDSPXo0cHI2nGHqkxd/jrR9OjW3P22Q96PmP9ffkVogvWb
myGnLT/Cj/XN0Lr8wjOPWAEESrSdKGkF3801d10q5KfqKXUlup3NlTvqC3V/atz8
CZPrrMS2pVA1acUaB+madJYDtKUi2qyAzkLd2iECUtIuFhLw1fEbfxCWAB6Hqv3r
kRZvLUP6Gy4CyvBz3HuugwN2iimGQJAzalB33WkY1LSTYXnQ1403pNZM0TiRHG5j
hDiR9oYTynPXyVzHAJIgDubHbHeaV0s3kSspQyYjyqg/00Yz89CuDAIkyt9U2+n0
rgWgybgKXuoMVxQ31Bmset2oXxWpoSqu4/1qgv6KPQo6X7BaDDexPkrtq/B3AmKN
Ui/RfpE+Ez7WSrMQcuhp8xRKNmO0sImq7XPJm0/98xWMW9NmrR1JJ36AbAzRzLxE
lrNWLI/Pq8kan8XIqodJKiplbfn8DC9+zTlfsxFhAY1BDpT4A/mLMicqWL+iJZoI
ex5tX0P2m2lm3+/ID+nz0pnm819zdoasrjJzl8N5PfumxSWSwyTbG5MZwjhs3dHx
qOyDq7nYTjFqStYfuw3ArxdhMzb0DJw2B9pu2PcFob7P8hBm70ewMDW8PPlwWrcN
I4LXPhuTffyw3W5hIvvGq50s6uHbZMhP9IpaapXp+QOsheyHtIRrglcZqAKq4iFZ
acuozXkcIsOBuAjQZ8v9onGwgYhlGftM4n523ZMEFxlNVEFmBwzmVxEHhOtQYr8/
9T38c/OpI9JOgYjQnofzvMUGhxIG172/zevUG3oT08wVvyLY0nHSsOGO+MYOIav+
g63nMsL31kEIndFhCw58GcDypr51xYICG8iOP9qTOHWXsarqpWeCBT9+0dXDwL1W
F9AqiSfKqaZekuVv0BroTXuQqk9DHYxeiGv9bMfQ6KnGIhnVmcU07V7jHNGkXjGl
M1+IUM7DEE0JqQRjFiLyP/yO9bcGTtmw5wikLOL3sFbYcgMZR7WD6TC6jX11iepm
11EyJm9qQOaq3aqDxvJddpqtL2yFY4VCx6n/Bvo3VmUii1gTmtJOy/drUlV5tuRB
8eQ54+omTsWXN4VWU8GdJ43qQrdFMaCv8x1kREuzyzwlV8eyFsMnIPwDWIar6Yvq
uMT8Tej+cNMVyhneXVbmlLyac8Bmm7y7tK/R5/onU3ImwnJb7n8sFN1hwztv7kIu
xpZMGYnr9OtGajT2WwQkKEf4bG+DL2/a/PK40Rt5/A4o5n6agP1plaNg7+G/QC76
ShTJDIAfsgdGehNXD6GBg7iaj1HTBL5GCeBZoCA+OFFEmzrVsv9k8kLkLAjS2VhX
yFQE4Agxa3n4rJYYohJp6WNrjRkJ0C4odzCaDiQgIN/1ATphCNc8FAdhBEfoCfVn
oe0fjbmGirdKsJHsilI4nibRuGUZx3TKyw/VP2NKzoxcf/BnRzCMlnmeHu0faOrQ
T29E7zDKsE2Jqw7RFmAZ0ljWKxQZEyvOc9LrO9x2qrnkNqymo79aHiUVMGEBpaSh
+nk6KObaxzBWmI1REXX6sf8QfIuPs6zvCBdEVO9ljRP0QGXYZfqsP9ICBlMsXJWv
2mATvD16vjzcew9pC6Xpbn7Y+8lNIjCXMNKa7TxSCz1fULp4w1VniFgruRJ5QS6w
SZwoISR/Tog0sofV1DHo8PmAfpMttFUi2/sUUzByOt5hnAd3LH5koWNdJo74ZCd5
tr2D9p0fhn4XM4uoNUYpG+ErYVnL2wWKdImNRzKCtKLi4Bh9hFUbaMQgzdLqA9x+
cIGe6dqDzk/DkEuLgqe++Q436TQmh/GFq2TxqiR4srVfbl2zlPQqsNra7TaDZIr5
QUkQ2+tAdcUD5Qx/AGRyy4LWqxRJJnOW+yOUkUxQqqrSNgBEndGIO8PLrqhWs96J
Eay5OhZPPZMVyG8ezatkyMjj3/XTPJxp/Tvau7bQHlE=
`protect END_PROTECTED
