`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FgFp8lI7a/Lyopt5jkXT3ePnwkF3FGANDt+DS5+EUiGXqxbck0VMYj9xKsRSR+lY
si2NkkPmyiFZMREWgcYDCkfXqpXc715Ce+8A9SBwYewdqfMcAkUXMdaWdMie44rz
tZlCpT+wewBfH30D8sJtoN/x2eSsL/AxbkWK5QUPeyF1/S323+vbM2B/IopHHYCt
3SlAEkKWeXfk5rALUQ30+3dl5Hi7UcTpAnUo9nYCfPBhrwu1Q1nNiic1HrTaQkTX
w//FowGT0bbhG6zEfGa1Y+029LbNRMlDYx78hi5pgoAke1axLkTZT1LRzZBXBiHJ
k20wap00qrnQCD2NNbJWbb3ratLxbkhVT2mPfpbaZ+psreg5vONpoyNHUtb1NYsU
YeJrbQJtFxq78BtFuOgw0/vQ8hJWtW24dok+0l9hotlIHiKc5NrSks5YeEiWcf6P
+/3881/zBwEM7YXq3SOwXAqhsl3HMIJPytou+CpOsiLuc2+Gs/9FUi+bsCFKGTRb
iugelqjOOudMUu0Qz2idEPUk2m76LUKK8AOJtn+tfZAY90m6EvtOOLb1ywxyQAW1
LneeQqbARUlWA2p68fADLo4pc+8y+DiMVzUnGX+9Lihvv7GGwpo6CVAZ8Ut7lrdr
IDF9Afv6EupvX/WJDLP5NqukyYtQGR5kflZ70kuC98w2saQnGLvzo33eP5gRkDaI
CfXHPierW/GwcwhPArpRAv/ZoNzd80XZiY7LCNLSMky7QH5efdIUwbJ08296JjlA
zHBhHSACz/nyUd5vVFf9R0JpH0ucN7u6xrDUg5y4npBKnXkRxqAtXWwpPTaYg0fZ
bBaZF3AtUXJVytVLiAoWNNmvumdbAHXrSbjE+Vfu9mzXuzp3HLZlx2p23Xueg73I
MbaL46xdimjc6rvicAjBJy6fsuECeZxJKT8c/MQQBbl4jVKRqNYfnJ231b/pc+Uu
Il6hPEDAY+P7cpitPn9uEke6+IfDG1JErY2w8IYG5o8ZdHWxp3sAN3uTcC7zg9P2
iS+7ud31uMn2HajIL1eIMcnGT7KKAhKJpSNXjk7BY0k98TOJIEklu2dOH87yMAqu
8pPEuAJJMAdT4p6Xj0yywUotxDuXSkhL7zSr/lxqvxYjdfkqmh3S5xRfHiW123aZ
BEGStTedz1rw1Ikshc6AWoqjbYbq4n2CSp++jbInIRw/sknHqCzE21IbIZW5JODm
twcWKYaM+ctxn+5wLHD+RVXmdxG36zO83xDyKuqaeOEFDSoMtntGU0NiUdUpNqNw
VejfuIzmtYg5bBvsfxwQBnwrBHqPU1DHXUY40MenBMOa4LRJFAIMc/aswfUr3S0S
6XePG5kIuZqTso9ARW9FnyPMlFbk0ubkZV6Zn/ymKi8XFJ/hJVzWSgHbt2hsgjpi
X10eceVZ7EsfMnG5SMU6LYCD6lOECWSZC2aT72nHYzZOiRBoFGfgOx60vhMnMbdE
o1dUhqE4FXZc9wHId2xWDiTLEWGnRRJRFMgLMC4Kxrazk3AwewjTqLJwHh5DqemF
pfd5sIgKrO4xOyi6yhZBG65i7hImB8lKjSBFItqCABl13TbcJBoLSfwZrgibVLvv
PbB3wJVC+s1etGUWnKZis7eH6MFYJpacjFo0Ky8B/yYmfeQuj9fERIRxbXCSZxZh
BxfKif+QQWZIJnEq7OjE6KwWeZD/Ke870ga13i5csoEcLJc/gJ5fsiKbSiCbaMS3
QnZ8Uc7V9owF9aKB1xAxc/kOEhDBP0773Z1fpy1orUD00+nysbRxKNE2gHAjnVOy
ep3i5Sm53AbIWTUzoCv5+KK5OXpIMmwUAp4o8StKwVxqi8b5XZzXvCVFdfsioFRb
imiAnHmYcy4AC1Rhx1pfHJmro0YCj62W65NsSlYsvZplxC07jkLtNmpiuqqgZob1
WtPJxVFCSDJ0nI7VEV+7FMxABCoIw6A8Fmefr19o++p38E84vs95wG7+xAxDPI9n
2BkrhZ2s6jT6MHY0Lid52GzKEiyy6yvvh2DyYYIuXKSzOMaZt7AXyAu3cYAfgOBY
jWetwAS4xLroklcbvRTVUk9Er6owT6cF0ZqTvGLWGfIGUM52Q/m/0myDv4EuccaH
kyJqwKq6MDsFjuYcP7lcv3fuhhN5F0cc/eYkqrHOPOj4RenDz7vOgKP4kdtVK4A8
JmZfYUda9U8ifF/uhrrMHOuYr/l4TQaY+RMq08nyYi0ZltVnf0PjdNc9FAr4PxG0
stcKtkc6UbETVzhZwX/MQbzF98NMy7ri+/lvv1lUCGaU3RX3ljqradQo4e3rAlwi
mL4Ew91f5olSUkM1XDV3uxMqclbAn8JG/67mejrtO3km6+Y6SKz17f07TeBUg/dk
zaxQBOViAATkXfmnPdfi2dTZZ8FT/CC/h+csDI218Iczl9ED6fzbaGBsY6SPAsp5
S9Yqomn4f2dDFV0j8ii8bbJihJPuKdy6OSOzKVi1ooGSApWkqASvCdNgBQ1YI32b
00GLf0569JrLKUam6Ns8QeH37zVkhta8QN5wId5BwSzSjnLYgLs61CNEHwD+wQmM
i01oJiF6fp5kjsUKNVtQPx3M2C5hWUpXaCHJwnmSECt+Wb8ZDWZbLKIKmwVM3FGW
/o0QpfH71dZDciNuqz31XG/Y60MpMZZDC/ZYm/S2L34XG54349DyqWecwh4iQOt/
uK15udCERtZDQV/dq+OOGl1oaq0UivbWj7TpKRGgHwe9YiYkOTb/ja+dl+jD+cuP
bgZIf5dcxJxOX97t2b4NxFqUb0n0K5c5XhYQt4MsN6v0ECx2aH3ogN9VE8NbiTFn
O9eQEi58UDM8DLXEI9c6uO/wTmlE0UWbbPDas519a9thDZXjvz7sU54kDBwJnRwD
rHbo91qY//sLdr/6p4Ya01vq/OJnsOMU03l6LvfN3hgv9JKhUaof9q69AIxBXU+I
bOcmtXOQzCq97L7jZRrqpgITqu2GUcaT977VbKkyqds43f8frVCHBL+d/BpRV9VS
8MCnXnZsEgZfSyoiIzNA0MpYYC2DZTCVKZ7wZhKtL637i386xMb7htUmGBEGO7bw
AGsow2FbyBj9YVcfJwFjr44Zz0r7Oh2QY6zBEp5GFdKwgpgOT8XehIe4us0omE52
pjuvcmw2m6PS5DaVc8ZKKJW2o22v2+0N6rwNE2rLwH2Rv3PGnYIKs4d2s3RISCT9
hXg2cztStHrojfQDRalFDI7lfi0c/OWyOHLNqgKIlKpR2JY3IQBvf1ihwBifNE+s
evbq7GPZLy2pCMDWw0wvvknLdfOSLbA4zqAVkFVHTast2KjqNFLbL7/DoVHmod+b
xqtpWzNXUs0eN10PAEwzL1Ouivxh8J1jCRmlkYL4rLAgOeKpl3sMfXfeijgKPMOy
fWRyU/6G3DooWUKX6SRr8n7JEYTgH/OHP3M6QzkX8cA=
`protect END_PROTECTED
