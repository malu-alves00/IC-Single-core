`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EQvReWPZA6tTh/lhCOggNPAfFT62FIfdoBOHhNMjOE9bGXzgoKJ+EQsXjh8q9oPS
STdACyVqNU5dECYH3fRlVgNbssHOKPrmF0Y28L3R4KP+x4qPbOdAye+txw/7Wjxp
uVfRw3ei3RP7p+dKhlCZnTPmWQbaYIxHYCBRvGmjgpkK9o4tOoTnmclIQe14bOG2
MLRjv46CxktFmBGmZvP/LH1w7HErfFX3TwlM5SkRY/ZkQskNUQD3gsh96A1fU6zU
H47T/8HTolcYP4KVX7yg/LzHS3yYW5xOKxBJ0UauOUzHmJz9hU8TfZEOqKpS7uAt
VM5tT090LdX8Xzy9yyYwTqEHZcD7dKDe21ET5TPMYcBz2Ir6p1TS2Sp2/Z7nnvxB
XHWE0Btusu86qvPFNaXPR37zR90nIvNi1nV3vVKANNw1TK3x8VnebTdkn37jxU+M
Dc+ebrgM6+PwykBjOZfKOJfnmId2s8DU8A8xqZmkLnA5Yf9rkwt9A4zxLjQYDQCE
0wUCuT+XZqBxcW+MWLiQIvUcJmgA1U3J4CzTsDqj4BzNqn+yDhRzki0qPGj6UR9L
F2+WLsX4JfstDr5tn8R5HTM57osQRMkMHPaSFy0ZNGm9yt9IcOpYhHB3qVC8eabO
Zr+p/YELLdxu317N86roieSc6eYBlCPcGukPsvjGh+HjMnMvPD2rF4s/L+BIt9lQ
W8BXOQ3vr16OZ6IuLubM98+smNQHa5yiERPC/YdcDXT273FlBPu60E4nIoGMUwaM
UDvpVIEQqTxHNfVKAk4IOJqhgRjVui+yQ2935r1PpBl+E/FFmMRKamk7EgfzxiGK
olMtiAh5dSipnDa0gYCEsOLe864csBxSaHcOmJWcLqk=
`protect END_PROTECTED
