`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pBmfAqqkfqLO7TqL5tAy0zaYYomBLW55rLLPM9eLTxK9pzt6RUpN6nMhPrc+U4gN
jISacHYxg2/rCXvllzle3kxrmNNmyGeMbtqM+WnQBuY4KcfyM+kvQRxTVzKyweqT
tkjX+GRwIFqW1FtQb/yhRT4CbqO5xoCae4z/pi29tMO29LD5HN4ieBQMD0JYX9I1
lW2E8/0SFfU77AvjxuEVPPW9O+/kEa3XfzwLX+VDn3GWYKplTaiaM5xAvYwItr3i
HNaVpAn3nk+JBNl0a6qIyp3wyeK1icFZpUE+ZSPQPE8kV/Ejq+oYAhHUPS+40k3P
P2BoYN1CcQWXQahIWBv5ooUkBKNzgJE+NWjoATVffruwTFb0Yq4F7Fs90wh695AO
W7UCCF2Ahs/8o2vIRBfjV7kJpuySS26zEvA8f6tTfg2HLcFdtLtSg13Jxb9dUNyj
gwvsSYW9et5DXoo0/LnXPAm30lVbL62l2YEMfvLA5AKht5cLjkLyNrhM3sSYRA1y
tDNCPpPIl8OwZ4rHRZ4SIT4+VInmXBB4Skewa354Yu6QmGLmsUBEmAVHfpWUOeRL
MfdLdTWgJ0Q7a1eC6LZwod1o3Hj9BS+E53IhIyRqi4kLU0p+8LJF/lLEQieTF6zB
x+nTIgdr2jq9BtyX2mgLh7YDJhN4wpXEAZs44H1uR1vBRyBkQG0fGXN90AqmoFeu
iwqbw8/zdOaNIBhPeHIpkEW5QxardD1LIOWezyKw3iEBalQ29lgQF6LHv+QJn1hb
La0xqQc6aMHRoVOuC9ZZ5oLGYVGuTwCnqS14fmByBokmIG3OMrd8DGuxK34lIaxH
WbYXjzbV/VUcFUOo3Q/ocCxoC39jEu0OiYmhcQbBDqrj5QIRK1vY8oBmFMs1SDaI
EmBZqMlz6J5qVfTT9QsJ9SKgfwR7T2OT9WJYAhBuSd9SMJN20Ok/2VeHTvW1bKXQ
zxBvf40xhYcpnEA0+dC3Nk8P4p0P01+yJJVJc/GB1tCFBRQC7Pc3kMxXyBO4Fmjp
Nb2z88Uf6u6detI6cYomCChrimhMNtwpdDA2/TlaLaSOlde/5oAuoB8yOcic5f7c
CfjrqkaVROmL+mRZHTp1tIWit8+kc2+Bl/N8BGTFFYr+oNEiOSbeyDLDA+xAn6hd
aSk6s66jdg474axcSWOE4Zzfkk8oax/ApoPbrlD9v4csVV9JZlKBC6TJw6grtv8C
WkPoqT+KC+R2m06AcslPEgYUVu0cBVXhhQ4xrw/mfEm3V8Qy9e6IOJ7JGB8PS2xX
cXiA2JmVDn/w906xIPYdvwGBcPnm4NQZ8tkzCDNOLTCm0DzmwC7ItBIuinJAGLj9
+n3KCUQ0DqCgJyg6opFh1aj9wCkjxJfPy2/RtgWIAGIkOmxR7QKee4nESjavxlFy
QZeE6my8VZFTUnBsm+6oECQLz/31kM88tcsbweTCPRWF3hr8Kt3nDDhsH5wZJfPQ
nm+C4hKZFKzxOlUzU1f8URSO7y47zHjoyu9880pOXSzG5wrzUqXR/JO1JejwI+bf
Xr795XnhyZrWjndW71zhaf2fwoMt6XKLRieUkJsJAPapx+lYLY0/whYunTxwqoxn
zPwZitFe8gNI3GxtxFUN48i/biapNPQbPdwG41aVdsFONWIhrBm4aQ362QXI3Z63
PHhPhR+Ly2bFno6RhdUJ5yDtuo5WGKcPw0QYFq5b5nJEdytKGpBUYT04B0ry2Kvo
y/tLC/Yrk5yqthfWurzYfK0YDdlvVe2mw/Jlri5yjgRBZMHrbDO8IbEmaBaIwpB/
363gt8beotmgXebv2+6YTngRzda4tq0bJlC3h6FqGgnCCWQDvTCbx4Nz/rKugbWU
vwICfaXyTmZsk7mi4+rE/brxVXdAxniFnv7k2+q7Vy+QSDcgON/c4FF4UGTr4yya
ZwUKfZ9w3GXkWubMfIGeQokCtUwM6li35O1gWpYVaUL9LBM/ngPiSuEzpi/m96/W
OagAPvLQIWsxuybS24QWuDMwKO84d2mbyL7Xpf4g/mUJFZ01ERciQR5pHm0CY2Ut
IXxV2hifZO5vo2eiIyum0a0HVsHgaWfXxSum82Z/lxGV58IDRORys8N74cAyGxLV
zmdMbbow7BE3cUzKneATJgS1TbCbLkfJqvO1dfGPrV3qWYQWRTTdQ+B6RrgBOmlV
WbhMs3JfL7Bb/VBQ72DGKHuIaksPNrJWSxX+O9xK9njR4Ua09JQoWlK8f9JhAuWM
VjUKY3AO78lF/QfRiWidTewOyMWsFPyoSW4kG5tXTnMRb0wuNyYm0XKU2SpyoYXo
dJJ5EG8eM3BGZZ6isK0AmlJ+sX+pOjhUcPSqgqgxPDNlSREpN1eXi2BLMVeVWzlZ
iG6KuKW2fo6l3mmC+Drr1A/ujRcmxlvlkzlBxGkmjFWwt/u1YJW384WupZRWNOj3
YoRcnW8gGgZLFAG3YpXLXUCVoweC62+yB90GLNZcymxjmreHjI26tAAPj4G1xFpO
jJxL+ZAKcngzk7kWd6rsCFcD+yK76E4TNdLjjGWSJ8xJKJQBQa8AfNmbRg1WDKa9
/3FMtKbDYlhQth1Z3afJrRilnsbvYFwO9IvMlySiR/lVxF53ppu3+xSn52qmTtdi
8etqOMpCn5nt8n89ob2j1rs+AcI8ia0v1r+BHW+NgacCEGNcMqd/5M1kMVDcFP/R
kGJ5j2E3WJ8ZA9SlrgZNnD0vYGdAg+A7f2OGKUklH9mQAshM+x5bFTuHwiVW9uUe
`protect END_PROTECTED
