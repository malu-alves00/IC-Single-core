`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3qoMti9MyHh7pZKhwXQLaMP9vs/arO6nEWO8Qh848SE5NXTaFp4EmYtGgUweF8St
m2BGX0vLxw9nzYmaJngb5S47f2wRN77+UVdi1T5xXjUyMcGM61AizCKc+wEtwA1r
1PsyZEEntF7b0dnkTNFYxS67nMmV+aTsq3C2Tn9Z2kanENntjHjfYf+laFirbZ4H
qqs9TjM2Jvj3Yo9jdU0VraHBSbpF2pr9GdTQoDTYkDegPZdCmluY5rgA1IAcPE0Q
vRRJ28fdoIzgvfaKa5HEGBsaiTGViY2ZSJ1hSaIYwCj4dfU2pWpfkFIjhDetseQk
7XNRwL98rvHm4qKB/TrHVBqEqDeXNSO6q6WYDBQ1c5gFIlJ+deFGbhkgkfBNg86v
bHzNhBncAnfDQWjXHWG9sCniwjgV8acoenrO3/N6kLS2wmG8mBaqfntiVkanCDJc
5B7sth10CMp/T0DQMrBJWlKTVRRcY0C8zccVDHXYa+rg2q+Xm5qh3ECCefk7c/pj
OvqA6SREsHfoY3KOvrMal4Pu3mtp0ajN9j8sLiPv8J+YIn1S5UJ/Qfj0avDcap8e
+lBVJW++zcAfEl9bxNAUBg==
`protect END_PROTECTED
