`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lI6TkwABQrXpt4gAmpmsopSt3d1VKOpyAp/O1ikt1mlZCph0VKiA5ipFHlq2y7KU
Zm7fsR7YlM3r0CURUkE9ntxiUCs7ldoK6LvcWN6JfGLeTpram4q5iLS68+s1Z8Ct
I7Nyy6xZFNJDDZEWJqz58Qk/Aav1tlfmVCldq1GJknEevZyf5JgEgzj6yPuq1zXS
4Na2uaCkzEqDlmvrghDnbyYOihbJB/78sH7dUZjyonvSIhTBspRGnXze4hsqPQmK
Z8G+ZUgFIKbk4gcRdQsTZq6pTuFW/rtRi8CYSkqwrs7xivVgr82PvfZ16eU7vCqh
sP3jS29faYg9/2uwAvicfNjlW0UnEGcZkqnHY3r4WOdsi8/EwzrW7JSFdsHmDxlL
P4v03sTEOAr4vjaY1jfwGaDV74CoMOefyXcKi1Qs+YmRAINRT+alkTkZLePluaa/
R3dFoh62u94Oyb/sAJgQppogGgLjXLxxMt/fau/RDQdWD2UR2BSaDga9Vlu+dq1F
34joOLQT14ehKFlQt4cZ/AaGyGHiM6QPIZTjj0gkBr96Pd+jdv+XzRh4BkD1o0+R
0fw+PYRgu47tA5XEmQQ4/MS57QJ3VSeDHYiRJjuWOZZbBYHC4eZ4RVw6+ZkeWeSt
vxM73kvk1CYNgKZ8Yzne1t5VJgXjBcoinly5zt23V7XFhuGiA9l9M8+9UbK/i0kr
J9giEoUINDF4mH0Mbok+avOTTFM78j1wYTs73JxnVtnIz+MmVK3lVsReV/3SdBQJ
KPLo/i2opZ+AFp8bv33fKLJdSyjDmweheeWuwO6a696AXwDeYmVdjy80qKx4TsHv
m05uA1A8vQb9BYpYbByXerA72aX/5Su5j6/YUAkfcrQ7SBZcA85gOoWxRZBLhdxG
GB/GNofCwMZsgyZH5VoUJvXx2jva4baUBOsia8rur4GWjSd5piI9BY+pGqo9cU86
ckzBvC+tf1Wyx1VUY0I1atiocrulWnC3pLn6nAXJKrbUH/qlMVnJbDUBP0WkjlLS
0Ybe2lZqc8u1OPI5/xIW59AuBc0HBcT3SHYGZ+arALBb3ouOLexJ/S3+V2kpECOT
VokeOPdiESdhidwuduj7N58qESChQ3pDjY+Ztc4d0RrsnlVr62RgJMWFU35inGmv
Mna6jiO/ivkKUJz7/+5Q0EeK/Yxc7x4azNKi+a5Bw/uzdk1AS/GPNigMP8KxsvmO
q+/2Z5jdL8blcIzzMKYnYESUo7SGGAZxn9TR/FZbmAGLVVNcv5wNJq9AAm5oPdlC
`protect END_PROTECTED
