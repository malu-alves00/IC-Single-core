`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1f4Y1V1QSlyNpIFV4erPa4av3hUSh/4od5nnGuvBYdVIbCdPhJcly18QS4mYnwJt
vNE3vtl78Lomhq7t/ERY/KAvLqKREclqREZzxmblXMdXTFleuS6bX6gAZNWm2oh2
r5P+2W6uBMHIwFJlbvNyc8JKcQju2vnKcgIj1fuMCjzD3Vw5IZdxzxHFihlwH+Ff
w+fA+SD3rGXVrmBTaSLEWk6k6UXujAzcj9CeP8CV2NBnsWVKiCZ6s4AgEFb6HxUT
vfh/1mZHnQxRMwvE1yaSUlZxGZs2w43IdBxmatMRmKBQUYzhQzCgcPj7iKImSI02
Nm7UXr0tBY9ya1tnxyctE71YJl5AJhjvh1nFTD5L+iICO4Pxlp+p6XKosSehrTeS
B1ab2aiWel2v+/5T2FS5OpaOc4m1dODbPZQz4Eyvm9YFBXwg2ASkPh2Y+AlX66C9
xiZpSv//5r9Sz6KVYClX6voDwBbQYpaX7c4lEUcZJBCu/JCJjO4+R885tViNHRfS
buGC1/f4l21Ibc3aEyWdrO/fBVxsS0q3ALmdKD1dtXEzxe1k1yKJOApqIisiDHln
caJaetVTidnaMai+qNdPO4x5ff7GhiGTJWhnu/Y2iJ5h77YJH8UcSASrjqIztWgX
DkFaJauI5n0JIkUZdhOLHuvwvpRZWqAYQrQTBLlue/peNY2qiLr0VZPHop9zbqcI
SVgsqtQP0bTnuLY10w/xyrUzZR1pv1wkk1/4cGXzzMlzK6aUC3lczX0MvzXAITnH
NwK9fT11uDXGugq1tnJaPMZlsP5hiaY7fxRqluRwKEGdSXoB32NnhX0EnO2MjtOJ
/xEbwLpA973M7pS2uPOqvZfrYRPdfVT+QcACyAm7l2F9KNrqY402wKIVGstvAuf3
30ZdqBsbMnIOJWaXA/NMC/3VIO/dx70JkU0FyKRP2UO6sKjLWqeoKMu+Z/fH/JUK
rlGBAWcOymZIoA3heTQ5+Jur6KkOmI6yejtadOzgF0i3dhSX0NVkPowNDZ+02Him
NGSco1/fe7aJf68P38CcG5qBU0i2lqYPRM0JF/+IFknH7LQ9qr8dTP0jOVnouWRX
GX4EH5gE2zbqrNbv/VFMaUEsl06ryW6yD23UPZ4axfZfg8TNYL9UpxyXr8Fy9UuO
JkTtwlb4EE9hLLxYB/Ftv08j/aSeSuQni5lQcZmzmrX5sdl8dwUkz5UopWjaFvC/
tK/zzkAwqghreBEa/Yvbxl006dO09Gpd4MneHd1y4Rv+Edccko9nRjSl42kX2cU9
zu8JaDU+j9BsndbTZ/UHTDSg1UbgPWTa5ij6iZByCcML2s31mYff8t/RUUI2gxhr
UK5yt/th4XJ20jeqSHZchQPu4jX+2SX55eSaGqaG75kY17ICbFJB7xUwW+l+Nq5x
VCMyZ8BILzTXEkoK21Ivl+KVqP5yGPimHNfqMFO/iHVuGoX9CBDXnVxUKwuI78cu
ebJSfYGjlbI3kLeGbId22+JLqsPbevzq3N+65oNvyMqwZDeS/Obn9/m3ogSgoctQ
`protect END_PROTECTED
