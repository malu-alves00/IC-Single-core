`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EV9Jo7xoW/h+HKHQpOzse/fp6ayZzmabQvfS3wuTvdVOsSKgFKoR7LOLueS8CzLQ
FnUwxu/MrdzS9/VguUeHUnAUZV3z4AFcv1LFdE5O94lH1DWzKj1VdLcfFr9Ms9f6
iod3ncQ8E2RcOKoMRcuSNWNLd7EirlOFThFc9AYXuPCsgCo9KbVASTOPuKJyYMoG
nn54K1Hd8lns0iNEEAmzpmIshasf/53ysb1WAiCL3z31aUaJys6+mrEhAW2DeLai
43Z3ZRu9DcLPS7WAp3Y3rZVRXRVbUC4J0ky/Gm9+40Ax+TjUnA82scThNZmmVCPm
np91Z7tSjRxRrGnm2mOCZgc+yl5hTSIkaQ0/NeMZGEki5mAs2OB6r6nuHrB0Zudy
/TzKM/rfXyNu9x9l3ADCskH06NOVMN73psoBcutF8os3PTN4UZMH9+LlaxcP+rpr
TjBwgJENWW+fmVvv2f7s3NBlSp67eIvXMFaQPKFVt7gK9LIq61n0zxYBb2EyGRJ/
FLpXpfO9+q0/WR+oyG7cWoqOFhrY+iMfiniclyWUpNjI/0Y500K5xcFjzsTsGp3t
4qz8lWE+nCl4T81ELrXRfH11eO32BwSCxku+1QMceqZ4E1IGnTl/h/hREg63pHEa
id5njY0wKfJhln7BD06WoPzUFO0TbQFYX/xTxgKg7qV2RmtObBikv19610/xpG2O
NculVQTOIl/tETwMeU5fQORwNcGpSRHnUb/WqL2KMeSrwTtSsD54gAP+tz9h1C2j
TXYoK0ojcAaZCTCQY5UagvtGVxjGIcEWYblPknMoc0sLmgwnEK7KFPm3yoF/HYc6
N7BwB/2lL0eQLIo7OliD/O+nBRjWYfuCIRPDUXpnRAeWzGViya6eLcRd0LydZrf/
W7eQAXXFSZAvQsPRD37SQN2EvTUoJ0orz/9BK3WBdhPu95GmQSYjD+lphphDPUsd
IphZFk8RXYBSPN3DTFTF05zNwM2V4PJ8+nVZ4EisR04S2sKVJLhd3n++KuAQLbzv
cZsk5f6weJlQ8raFbnWk4SUzWEUdHff5Vtw1KF4W8ZjhrioWUxvg/yl0ImJiRJqu
zkA+40JdxQnqZgmuF8MHzrOZVL2HwidCm669c9YcAbE7rVB5zoYZKme6tAy/PvAE
krf4gQoS/pWXfUBWhhYXgQjoBK0U40t/I379lYOG1p4o8y2IMiZK5pSbre4GKaHL
ZvCDY6yegM6rBYqOcOeOcWfrRYd5uddebR+2NZtzwE0PH0bjxoUYFNJY3g+MFCEH
esqn2hVSipxPS5MF8OT0c4TvZJvBHhQrZHE61wwjd8nMud0p/RLe44HOwvUZrGVY
bCEm3mcgiJnlz6QUo5esG+wxlUP8SgJHAbrC+U9HPcV9qAbCQZz93By4Hq0595cN
9housvJzUJL92jJkbBMg2wJcNLEoFzzysnrH9ZcLTJWBJMk0/cxUrs+JkTjCbe4f
Ibfnqv6d35S+lfJz2L13WzHTb2k/aTtByPxHFrpAnG0EgC1ghIaJ36rfEI3nvDl/
nJaoAQFM1r4Tp3GEsLV5+CsvPLcescECSMKlfk3nKC8yFvGiDGiD2xowbKa4ZfU/
CtZADIceoneo3EX6qrjRuZIB9B6iDFs2UpbzKLrI/eqjq8GT5gbFKw9dOzfna17L
83cJL5qlL/xfIB+BXFpGHvNFvbOwjoMBS+8M5O8ihoQ0q/yK66n9GWqlTSjmOy0U
/4ZV1k5XqGtU4TD90ar1zEKHGg+OSNEJMOA6Uzx2OdC0Yum9L1wFj5YUC4cKdxak
iTGChpTB936C2eEQzmy2nHMNXUtLy6EyCTg6/eRUWmm9eLqgOH2rIaefEEb/CRFQ
lmZ85JGsLg/J3r1X2sGfMiFjrJQFH3bovttxWt9jrlFkA3fnofUHYOIi/Co2XqzZ
MCP6cr9t2gK7hIAm5uZtjJnvJc3HrK6yF5dxmOigAyePYz04FXQNmWCY/V0e7wDj
L66yNIcPtcPW7rYIGpyzqxtg68knLE5yoGMtlNpz/1fAnh2FpbGlYvmVI4zaO9Dw
I2T9EMr7Qus2SvF/0lPGA5jWuxH7fTu6arlpEjJ4ylhlMMzVqKSvIziPm8oFVl9I
0nzEV2D9opSziO4GNqTOWtpidgFL2a88OjAu7GjOBK6XjUwST0Eb/mEr6ihlV7Jh
EyMKsM0Zhbquz9ZabwR1/uH5rtFQfRQDgEOdV8v/YaXsYl+ZXTX5HR1exUOKzdMN
jvLz6eUN5HBimG5pL7P7QK0yic0/BkykMShBXUOzVz6uUXci2hB/w6B/cg6+u+WH
gNhkogD8Kcn7vzhYxqJgGBNXKjOrl2/JpBQorlojt/nhfcKf3kHhWjszE6IB9B3U
IGDf/HONYDKNr0Vcp/u4CsFAoV/0hfocDFX3T166SvVCvtQruIqDgE3VS5fVH1L5
fh0iYUh7rylfq1InktW0zipRtTknXtu2KOyU6QV7u4A55C7gZHHfE7I1oyVeL6rl
xJejZIawYx3Y7mLhWVG2YzTIN5o/Vsa++UgBhKwsK3Yl7sUau1us5laenUj0fxlZ
9D8hHXHV6wxNeziBIr7353EtFAkIqDxYSpyUaBpFbzuybFcmehbscn2S9VrxvI3i
WH+XAFr8rQVpdzVGqhbQcx9h2KNApUFLRMDFwRZqE7UI93NA5ZvwgUSBqKq2e6UX
ffs7k9KoNUkE/kn4ZGB237kF0PvAoPQTmQ0zzpsadl7JbpyXzlnbGXa/fKPKVl95
fvvLIyNz8Qz/ZnieWpTB6oOqlimP83d/kM+O3u+uPW6fA0tHOFrfWVpvowLgz1ln
qTdzJFCboQ3QuBA9mKInLsmEQE08ErqYFh6QwPX+478CWZv2Caxs9mIsu2Aiy1z6
3zuDqk9wc6Cdjs2RoK+LcNwZ3/emsawDyc0ooEvZyGvozqjliOsDTJgc5mqgolzJ
+IONisexnJju1m9klhyT1TU08wiGribAGyLqwfm7jAZxDEUyTu3AE+hSEgLGAK7N
tapEZWI7UmmgkfAGHofKYXOZ31TLcwq2aEMX1FHgaylj8dnHFgwNyI22fxblX3Ev
08ACGhImHYO7vKC4kiEAjUcb8tlFG57DSu1VYz3IYE2poSImr3d2zKzUTGvZqCsj
RFdjSVVwiNrki0+SBMRcvRA0vDAcEWhHNuqIr4Qekd8ysMSH76jULEgfoL601S0J
MBj4izAvlHX7WMZzNmKuA6x+cf19MfgTBNfq0NTxo2uz3daQVXhkbbvsHBJFjW1m
xOUjkmBYQQCT1gmtLpOdZVGMcy88pHXRmgZXiEtsOyq/GGIpjsZfpNROyRZgzl8/
N7NCmcpXqSppC0NuSgyk/lz8DZE+VMYio5yWomo8ek92sgsB0SEAj1UW1Sj5bl1U
VXzGQ7Hyf1OMHnMCoNo02o4wjx5QbgolH588G+bUcC2+GL1mRMUFpTIPlCQCndRn
pqcPw1wHjkAe1h9xXFIvvWZ+VZBbSk4dig3/wOYTGMzfo3bxZQ7jRiXNxGd343zV
CJ6eU0pfhrx+JwbznM1EZTcWm7OrsqO9N99hXgdzwHn3fvVs3AMvc4v6IaaSMRiu
3HXrRiWk8L7H0AxE2KOIbIpdjW7gc8hht8wfpcmV6ghrqhotem9B+jUeoH3mgUn4
eFYseg/ZHiHSI4Oapw8I4rcan+IetJXrMFH6RgOkdWzlfKJ0pVd5yImJ1WTNKHoO
Ajx1b9XUHhKP/LyeYJfinU1co4PEHQ6oMFn/FSkZCuZDvjC23BIde7pXndWQFOpV
b8+/Hlw6zK1vU9e32rukqFIqfefqbSJAGJ8cUpJ0Qg2SY91LZGk53xncUmsMz7Ut
jL/P9s22y4fiXYQkvlH1IPPWpkkO/YjrpJHnTRboBSJAb3H6JLGti3Lo5mJVaBsy
z5jPg1znim+kmdtIlAALciunAAArpaK57tg9zob1owzMQD8JRGdK9BFg9CzLD1l/
BQe0KKv8Tp+GlUTaWyw0EtfEIVLM8op/FBUdXiu3U4nWc9ZFUJ3DxpvvOnQ2IHuC
E8KDULeOwVfDhubRitC+09OR2zvFNVqRnCQj8prdAf8crti30rJpQWr19WsV6jZ3
e5rjUZNNrJjtBGhnkO+OivspPuMFlLVq0xZZ3EACWDqwEDRl9YnSR4wNWbLk6ymL
2TuA1jiRvCexKSWQZGoiqrEpUFArT3Q/MW6uq9EUiTzyxUpmmQgrpH7icCwrEL6a
/QYHO7NdIcFaFDey0Mh4IlAxWHiFR/TpxlEvSRt95a06h0HzKG1URavT1Dv3Hz58
FZuqYM8GQxtoIJogvu7Bar4yIg+fizWYtrzlwF3By9SfUjOGjmLQbgI7Fez8uUS/
CLu2qFTwMjJsPywyQqiGEjyK/tB0DpJRwaQpL1HYiDUfGmfqxPIXlc8DE6R0y/6F
tJ9pNSMMjSys/7hff6UjjpewurZ/9O6Gkn1jCr2wQFf8GxzojkNVDL31NLuG2FnM
41AtYcehUq/IqVVPAuIPPcM42L+D6GG0bOTDEA8cImtzd/7NrQfP+JZmFKQHFxIt
omWJmB/83M9dCuiF9h99oMkPLAjAq9mpvsN74qYLZPkqnCxyr7G3QWYK/1AigtC+
fNnw1jYqIqJuHctOLuVKERF5V22Wg9eArBXHkTjLq2gSi70DpwQCP2zUxk7uLPhW
pgZ3pdfXIK9slYWKPSUKOIdst9RlwIxEmFu7yCF+Vl1D/2sB7bvJkJEE7q1LKBND
M7xm0ugnCeirdjl2ckJk0ppppoENWM0Koz1rAaQ9TqKmXoD5yaNPnonHL8kneCRL
hwUE3Q1bYUCFIziwwPoXx37vPJmoSvN4upqYauNIYNzZK77JR58Lqxtb8I6+EfMF
QYdQFsfJgI90BI7dUFvVB0Kw51M4E4xtsc53fhIDH5tkmD10KS7HO68NHIbr+Sgw
G4h1piyQtof2emhnv6oPBGh/CADiwEEMptVSpZXZ4ru31Ii31JQbQZaW5hc5IXAP
9i7XI3JlQrAS2Lk2bQ0PmTU6BqZl2qA0pMpMrH4bJCyL8VjBiBlHco8H24N47Viy
hnGSUgp8qTZTJkLBISUok3REI00YkKSOBkCntAd8ZBeRCHbDCTEt3F94WB2n3HWv
N9If4Z97AtxyuyvjYPRL5t0Xnf9e6u4/0CnbkaBqsLlUBdIlFJcdp2PjoU03xD4r
NJjazyiYnx7TBjymKbZJ1xHWzrFWe8FxyLTODHEOwdpX0WBpaRiSqLr+BIxomGnj
qBqFlN3+HPgfjUH40jO/igLwYodSB3iKz4KRRqJ3HSdjWDJjebYm1ChL2seEQGT9
xchHnyxpfhj2i/44bHapdCafy04GHtKsDOQjgWIlesHMvOsZaTO8J495W2GewFp0
rOrXKieiMIZPJWNoXgsXuu1jLp8Mgaz6LJn9aGP3VHAyEg4vFRhGqe26t1mLCo4N
qEDSrb+bCrL47tS3g3tOblhjR12jXhUsZG9Xe+Wohpofj/Zi7gqymSN+A64Vhs+R
w7LNqxoFp7Xap5DczIqR3XyCXijUtKJRI6ilntfN6t/T3akgi9VkUELedWuiKyCz
mymFaya+dcp/PjQlXk3ge6PwcDrtArzlPB4StGSHxg2PY3RHLPy80IDOz/AYo8Kg
CVRL2hY7jRoVe/q7+8SkejSY+0nm2mRG+6ri46k8xBjC7Cqeqa8rXiatuWJ1L2Pq
PQcMTJ15JIrcNXM3ABqFNTr9RWpoS+4XnaQm0DMC/JbXgfoXjW6dTfeuJ++IZnv3
hC8jeA3PdSffqgQl7Joha1jR55k8AKkO1w2OtxWWQ8QNWQjWfwz/L3LdOM8cWxZD
/Qa0Xj3h4vKBvrQ9+TEneB8CbEBBMchjU6s+3nMUbcFuY2KndLr68qg1++zGXJe8
Wzx/B/gGPB34XxYZgv4oFIefHb586twrCG0GC1h5A6n+Lm9CKyxQgg//jHyfFq/4
KmiWrCrbKkrO/q41HiyDdutDTblHbCv+f8hC6ZXCEn2Erl0K/luV70KWqcr62CLO
EUlYtQAFxDKvEy/fuPEDY0+7FgY376RBmLTas1C3+fGy63covvEkJPayAiwJu/aA
89SrAmtSbI5jXwTorr8b4q2mbjHeolEq1UTafWRtJ22DG1DYr1krvM7TA5OBeBhw
qffQHg5j4UZAjlBIeOalSkoFj91BQYTx86VY9DD7PrCslfVmksCkscr/A40PCJDF
AiSkK1j11qEj1SqfRIAI+Huo9NfmmHHHM0yTJs4YQXt1dMw9JJVM+wRIvgpgJdCK
X0QCE0VAwTPKYru6yTHh7zXovMvhQIV/9SkSZUuBRcleS0bl+W2zD23vsftCh6Gj
9+C3ImR+X5IGvJ1btKE+cEuOfxcI4twaHWF/N50Id5ouobhuDOQTNK//inB9aR33
IugitQJp2ShE0w0hO6YZKHHGugwfO1sneQ6ZHg5+XyTGjONXPSCv300z3hbYz/X8
Xa54yjDPQ3jtuNXr+0VUQq8NlfC56nRazDCLdWZfFHxV8RG6yW0AlXYgCvTja6UB
/WfzhfDnTlNRhqBIUVtMssL0vw+yJNFHtJhc+3djGSL1xChLKfvOoSt0GV+hVJGy
1Kr1bxL0lfidUVFEsgqbEKo34v13rEbdzKrLlL2K997yE7r48RLtCXQSY5JXdGU5
52OM84uA949x66wvRtemOtChweB+CRt4REv+1a8w+dHSMidxvEGOO4mr0ntxpuwc
ELXc01Bi/WOvwsuGYh3023c6nqK23yHGrR+8juM8YaFCI3m+XyICeEw9pFxJPpSE
Qh216mKET8DZvQhDpUAt7xcD2YuOL1cBQiMSKuip3Z4r7PCgY5qgy6Q2oBwNVu5X
poZOKPBA0wnJyCubHUB9ZJaop/AiS+5O3IDy/6EBW4zQ4bQwXvwrDE/aGLRwQ5V8
KQVCdsGP6AwAVpL/TU6Ap8RoYmfNLCho4jAg+5r35wQP30TutxVtKNG065mvTG1T
8+lQaMabUDQyx8Z1tar6t9G0yhi0L4kqQAs37CTNVfK0SeVNumlr5N1zfqBt0hT5
61yLrWzOfRjHePlm/HTPfhOeQxySEZe9y1bb8f5eOFFdUHz2E3S0pe55RiEvOJ+z
C+rfPoTVJUuanKuNs2+Eqlkui1Lx8/Zk+3X566jtVCIAVY2K5qKfuteIRXOED7rS
iSkscJDVHeLS1DPVYI7//cZJosr+uwGrOszAfQGBMeQk1UUrQH+r4lZ9/ye5RpTk
2gsAFPFvRWy2nI0BqybeKEiX7rRediqc9TlTFuLcgJlrEhsOZ1y+7vd+muitt7Uz
euIR0L4CTn9EVPGKIR6RPxhVZsBSFVs0XY6ykqpzyvGDvrx37E7EfGqV2GYenPOM
+E3gpwMdVNAZWun985EmdV6Fx3uFRLQW+j2yinSn+PgEZ27Hfskp8qXdMRtw3tMw
eYuzRpTtvcDh8P9b+qW68QyhuuYNmogrSThdmL1Liu9dDFJUed6JTmG6HyQF4Y99
IzoGAxnxvshW8UDuH42SIwjTt6V+dxJys2BOvqzCTFWFo6o3IhnuZuHmRv8cRAgV
Z5BfwzN54pTsNMa0/PAyb+amCqGy6pqYdcRuifIMu/H33O7xwcyMN+VmUwueDBc/
7rGqSOBiuiN6E/B7WvGZECkfoii5+cL1Uv8PsuMAP1fX7Q7l6IAnQ1i3BPojjx2C
sf9oyQjSEfnvvi+FS7liSsSGDq4hg4CcFjoDqo+gcsjXbfM5XPe11LJpOqn2pgYw
9lLcvpV/k5SOSgodSeiwoVqZfvl+N8jTBs0O+qbAaIham6bWWjmj//I551Y/9zfV
TFFdlcPAGxBk9gx7hQP2EIWzmThld6UmhNVZTh64n+kD9wsRRYZf+n1O/JpcSJ8R
6Cg+vrjPs32utHhEAZ5mfWhwFrTNu6Q8xe2DOLtVZ/5ny8Wz/g36zowchkKS/AX1
0O7RQ0dyh33ywLFcc/Jdd5bKqwExpjPMVGQUdQc0MZtu+8VRPrC/md1FEHsqBswM
zmuaEUQ5rYriGUA61VjHMiqdtgITF6o5BAT+6uoWqvcNPzAFAAZAR/+3OX4YQt/z
ITnsXcdjbDxPD8d+kb1zWsULAGpnEK0APOhlhLZ+AqKZvYBAmLI0w7IBwsAWDRkL
YBsIxg6kJ9jpvzOnrWEH1wTrEAfs9gnkAiLN90zW8n0chrqCkP1Gnf0lQR5wl+bW
T2SArRTwkxb1KjEXBmwhyESY6PswM6HLfwB2ZNoQUP1O9/1339vxk1bD9JhzHsKm
ebqdUsDTQaRYRvZT+/061yzna3+/8LLrY57hq9THMTjxblE+wU/MNBq4DhuTNv2B
oYEMKEJdhHanyz9W2FOfYdRLopQQug0yVRQC4ezsv77DZHSLGX6Bb6enDgw4iz5o
9vyLKXxAqYfBozIYMmlPx4xkdQAAn4voRa9qGI8nlFk3lHtVdqH4QItqX8rkDUEG
fjJn6Dh0lCG1nW0hD69BskwAlmLrtsXEIa3LyCtuEqpmC+KSVlANLHfdu72CXBl/
FskL2NcZy4OfhwPCNEkpasXWuEQsgiJBrMzbV0dvDi3ProDg+6KXUmKmhn+/Nkx+
JAFrfkE9K65DqINkTjP4Haq4+Fmiwz0y34QVTni9ZYQ9llaLofWYGQbPeaCnwV+U
CpUX8cQ6j1NZzuyZO3qieC7UeLOwKjQoVJM/g3cid7UB592VsUh0X7CPAM3fXCkC
FeVZjfhKpTbEiNgjfsGC0b4uaU85Z73CRvntx9A4X/j2NRKuGMiQU2S+eMbVqjCi
nNUSbrVWFHSGmKsRFjqebmUegi8FaMkieE3Sd2q1vGZTY1FWbj6rocLdRkihMqLD
1WFYYSdGn7YktV+S1gpmM/iMK9Epqp8jfzGSTCwAmuu0TwjIyo5gFhEZapA8BLkt
N5B5OQ290jbkVzbmo9/ldHDmyRnG7RJ3Ut+qeOWLzEVWImabUitWmlg5y+FHhCe6
aWXCgr0bvX4js20+SqFtTomA0TVEVqLw/H6EEkJG6EY7cRfrXzpVFIwKWQoWyqiC
3kCM5IjBle+GKAM0vBMTZqDJlzAq8PH/dgsLU+ve68+CCnpmcVECt3eX5XIKDQfb
YDxaCNWTIxX6st9LjYIKvHTBiGI9CGuqYXHvK15y6XElW0TrpLxy162K06yyGLkT
ZcrfRp8JVbrJVD2TQv0uT7lWE8WE6ljtJqspudJeNmHMucW5o63WlrxYxgD1+ZZR
z0M1H72dYCmzVlMbo2sMM4pZg/ennSOcGhgTmGpRoA9PJA5T/MR+JbRPJxRg1ZOT
Uw8mb1vBfLuVHCsEGunDRktiRC9hCGzvVC9MRTS8l9z0w1VEkBbhKpU+Vsf3EUUX
W/puexwfMeIeMrnHLZzzoqfPLopYMQa6Y28FWKd3kd2W+8MRCPPFX8vNh9pD0vZs
qguB2kQYMjcsj/lU+BHUJT8K+vu5so2SNhpKWmSnb0eQZF/Gd+RV65Qlvv+USUha
F3AQxi9IipX67UgnHAI7PJBCrkIs1vSzHDIH5eiddPixu9T7gyxo/CHpGfyav1q2
r0YTe78rXPnKO6seA1PeriSi4FV93zR+5YlOqCEasjdwSk6gdO2KPqz45AfBR64m
RH1ds7j7IA4Gu6WyYvQwZnv2iQCSjSjvRuEa3H0C3RTYgofLbBAl8bIiaLKvb3EF
JWK16SUc/+8LW4T3M1HDAM6S5mzaSFjij34Gh5BCIsSGqUwxMfY5UIbZ1nX0DGLW
mAZUbnuQncnEF5qUqPs8b0+Tb+CrnvExDhQ5UNABVMg/ngrWnLqB+91C7ezpeMIP
C683BCF6GTg+TX14NvdVSh2EL34GMoInPmrfiNNVMStJI8orWuLDjQyXAtjthoWk
/JMMppiWkw3lStuaJMVY0ypdcY/DSAybb2sqwCtGUEMfmKM5GnKOwkGP0B0iV47u
o4jLUzmOU/pl3KKZASoBDG0Vz4dVvIGuYAw3Q0z20RJ/z9e6SQhDqTC5pWh4jirN
hJ0Imlh3gAsR6yYb7VWr7TG8OoKRiScJJY4N7NrMQ+80TFD7g6bataMAP6651i2M
uUBKZTJFuUh1YSQ6s3mJYRcFbGB8XTMiRiA/8TSuQNRzgqHNB0r01nknJHW+0HDb
EOhDmsJGvadCLajSrdFiLIogia6eqcedQdUshGtaWyqa6d5PjsUk17rGBUWQsD4B
VDwiYFNtL0J6WDsFDIrjqDpFctUjWPSw6qYvJILVfXCdULCAnK45Bp/6CfSQPXiX
EwTBIRYrcaiH41UEnOdu/MPIhejRA8YcKbbcFPRlVqAqd/CCi7LflK+/drghZjMb
LcM6LpaQ98V4U7IATigGt5i93GFsrNFhFirE7wRCwh5qlVzPDLiRIoy/DKPAHCF3
C9FI+N3v2zb/IqyWUMDCgPVfTQNmttUvRfIipUvjh7Mh+G7zGLxz4g4FeKqkJ6sX
IW380D+ZkDN2DbPr2HPLSIqm3BkzwXic6SM809Nlx8LDVC11PAJy3MuT31d/wDG8
p+Zlcx99pWBfx5L8rD0JM/vM65dyowRlUMGa44sB94gu6UM6yNLnnwrj/9q3yISv
jTUWw9OAhZq74t94TIZ/4AGQezZgQABzHQVQUIcVU6N1OGaGTc6ZgF2nF/WLaGiv
0K8TEvlJ7rTXWOXmbBuOgdCeiY8c6qzgarT6s8FdZJrPq1QHnBQqQzzt9d2EJxWQ
4ulBJfjG3t86mjFZNKVqPSkKL1UWrbU3cgOn0kiZGkUpAjvECchI0q7wWclXof4j
0wFpw6HdcwIIfIkSCcXduv960kJ5VVKKSlv5LEXWUrootrOPn0ko8h6OGz+GHBx6
KRb2Sl4hU//dOvPfPgRCaw0OngDbCeIUjel+LtMoXQI47cHBphh3oUPf1IkYmLpw
g/8pWHVW5ZvtoAagQTABqqQrFKf+ZEEfS4qfO74GBhE8DqYXBx5yQstuQEbVvKz2
OOcsnTTkzlyxV8rz3ybj825i65TKPaF9WfL7coe72EInnTCEzNahIIxAK+mb3Q5P
Bx1sDtmQk7gKD1YO3lsq6kUCGjrpJ6YV+8OxWbN6tR00keyrRnbWjpT9uN3Up9W9
4mksqiNN0RqlhrZSnJLSACqgcTbJjxQ4+TypornPQJeuov7MVWQCrTcxSkVhV/mg
xwRZQY4IDPq1CnG3zTjyKVnqEoWGO4FsNkbcqUo5WtukXBMqEuBWQlCr/CsPxPFA
SodcaU+7Rw4dyNHZmkxmr3Mrb1TSU32844cQQpOi+0b9P6sy6Q9Ufn/AbP43ZSms
T0fjahwtVEHJqcGLvH/NjlCo7fIxW/W33PziuNfUu7mpVpLDejV+6Z0JHfGuKeNS
HJZhacB6lpmfh8By+Ap7OjcelIqBS0u671p+5DoT/8JyYQ7Kx8dsUi6koW2h3blz
RiYRh+UkuqLDynV06xYuLe6HQ0isy50wQCfc6pwHE6Zf4XQat8XO9D9ieDvKYRgn
yK//bIZ4BbfBk0VoNtMc3yqpvdG/dTCRmR8WfIkNIDIDUCQGUJEIZmhp0zIjihgr
kiFha1KY3sWPVUe5qUIqkn4Am+T3qtjeWJfDp8bl48Hnm/1y5ZEv/7obagXK8RX1
nuoulJ+Sz399Tu3xU2A9zdepqa4mf/4fvCdIBFJTedhb8hXI+LjuGo6e1jjoKAgn
Xepya31mHM5Fnvi2cXPz0Fmumq2cqtNERqHBBG18TzyWJbbso9RRxBhTmiAD1fkk
Fn+sNsF4arfG4xk2XxjadwgUQ0WfTJNW4mx1LaYGbvuSkKJrJOnGr18aRjRfHqAx
N44uXY7U5wNf5+Vfsjdt3zPvDLrqiL2WnKHfEhXM/EUsacguUg0W+hfvLlcIUhPf
2m/N87KY12590zNNYLtIWnte9zhf/HiONZLwWtXXKmFekevXcItrGvDXMzZ1Yv9/
aX0af+9LHOqwLU2UCTASIhponS+cTsCRp9WF0fwhVT1+WYKWQGrxnJFm+1CNn4RW
ceM/E4oh2O8Gn9JcHi9UW4IlU51wh09rzcdXRzaJPzW+AoO+kmpUGZvTdy/LMSTu
uSc6StIEeoC6cvYrGIgvpWZck3uzoyywVY/ssArhW4g/UUKsh7WZ9BK176+yFofY
L7n89Kv7hJ0HnUqv5/12YPdBAY2/U0X+MP1paBlnsxd1VeAjKH4Skad4v63G2BZ6
6c7K0T3eUQRto8jN8e9r3uN1MatJddgVBPNeHks0X4ZqebghbfY2YiqIYZzIeb9j
Oe4gSQCUtEDJe5tFQbzBCZGs6NbMGulyR+cZVHN0y9gdK3jjIVUYQl1K7CdKbLfn
w6m3/8j7fLF2ScMigqVkGum+8Owsr4jl0jQeRDZa1uN+tkm1wdsZlHJJV12iQnnZ
x2wzRVBDyeBQfRzo154VFHiH4qA9Fq1oWs7BGO376qB/2b3xodFe2kW4c6Kp0zD6
5NcUjwq7Ji616Ivc08fWyrnqz5x16c8gztNOPdSdhhzd65nZh3EiR/6ZNO8JKMd2
wxwgjLL0cF5kwUgvACCTx+7th2JMRQ94ksfMAtR2P8Rw+vSbH7ewa5C6dwHrrfGs
Ro2Vi+ZyHEkTg5B3Xzk7aum7YcEKblP6CNcIYzX9FBXqH4h9waBpzzYwTsTeAedC
38AWB0Q6nV/duK9xQNvo6VTTk1bI2V6pJSRVEnwcYikOW4gzCIIXYjyEPw2paqSw
bgUhLx6vAxz1hBgP54HOIGmD1iECAS0IKPboZrlqP6Cfk5A/2B9yrhjmjuKlS2pK
/FBUBn6Wx7rkw3RD8lD/jme45i6K/K8d2aGqWtoViG5jNpbWinpMaTTyi9+qeFRS
irIwJncP1EZH/gXiXGGWCGgQZ4xRH4yyGq86xCAA23zCAXfp0pkdgEkP9sDY53du
fwtE1biDSlCWml8Irvlon4HOhn0oxDsB7xcsamLPTDcCHXsk5PhAqxAkvucm4Eme
QIPKH9m20vTfGce4GDCnYkeZODYjyqAhBrT86mNVrjFsPp3FAI3Dceky08k0EV/G
v1D82i7lKbemj87xniUN7sjdnrcF8KxLexf/9fSL01ltjeQZCBcnVUsIg5Ya1A4t
bl1SMF1UI++vP66PlG509RtwXYZPILSTVU0xw0vY+ib0eujWjk6fOuscMQknzFIh
+rTiEy4382qAjuaTs1fY6LE6vi511UmjKAjIR9/31U0KyWSMYr8UcIHvoNjj/J6E
GMP+VUkfEzK2CK6h4HbwsHwhyTR8kU7sOPvsdYWnFpzNP0NlZZdKY8n6K8qlKfRV
kFkqYiEDvRm8q/hBXuBTG4JVbGpbI9v2PrpcNm44mgiSutkexfYvF03Zb+l22bQy
cqRq2AtYlugdGFChUQ6VeJowZNQihn+0zxmq0epEhlwDoOZijn97dYZUZll2aVJA
lgvSBAkyu+GTHwHzdAUjPMah9k4nHuXHBILgz9wKh7g/sZYnP/U1C+g7Arr8FHFh
r1f/vkRP7BMrDEMDtveLby40Ftoc7hNZdoasPtsja+mSFs9NXuaSDK+TCH/bhrOk
49aM3LqUC56vKUCh9CtICeC5LiTAe5uR6gBcPiVmyr0jPXgzpd2JqWxbz617rCvv
Ox3++Lp6T4bl7IWxI2g6pjRPmNh7qUByIOnT0rqYeCeG+7IYFCo64V5HgUMVY1/D
kUoVTWu1Vb88KC3eykASIujFtjoG9z0exxVTCq3IY7Yu2tvtOdORUd/Ol+3dw+Y+
Cu0BBxdmoWxEZYq+X/zFyIrRYc5SW4aevWl8Af3vOcUIiTEYtzjibxA7QR7pi2br
EECIxUXanp4mw4O4S35xqn8c4K4BXzVUWbDjWneCVyUsTpH4tRk4tB4tzRx7Bu+t
MfoEH6zUwo45Pd6jj6MwTQnqLtN2DEIUKxAF8Ja1YxeLotMag2nCrgXl61XsAU+0
z4errVywJyownxuxig9SIvQi+f3IZHdfSyUDvKBOjJBZhXxsSE6x4J4rSMDvCtjS
dJZdBvuYpjFKFQmdtkam+fELbaXndlPxp9TKmFkqxRySSglB/CWWNLEnX+YbAPiW
iDKcQVt2uR2QvjTCP6E4PDegarYjiOikStF5bXOf/JVpJT429chfKn1kcWOyRdh5
qFCAoV0Z3S8LuIFFGPKAsd33eroojGbbebR4XC/y0NvaNGBxfluPSb59e/i1FWmw
FwMuxqsZlDJxsNRC4ARcOLysnu0rIEIgPtbLtZEatet9wPMAgcsXLZeCO27JIwGS
txv/GedZwLXbmMrLFA74//nu2yoF+WWgo56v1awfzel0D/uM4lAcBrDzQ5Evkse7
VPndTPkLD5APK0B1lVdes9VbIWZvN4bXtyS6vO+CaDb6T8/CCwUOAvXcU13i0ll9
Y7u6cfJDeWGT7xnBF0Fr66Ob98oTsfCc5wjOlrlhoKYRiMZ8HGTfkV4fw2izC2Uh
cQ0911a/mMjnRpmV5mDbvzOCueR3jMZDig7pA3Mgw3PuLl2LraPQ7C1YCwmlrhiw
i72aTdPRVWo5zpqO5dI2bw1+aJzN1UrYcx90v/7STA84ePXR1qjdsq1M/uFLn0k/
nC6S75+sht1h3hlsYkWaiWsUSJ+YSiKtNPhvw1/47r3RVeLQvqVUvGnNSjYb1MJr
SGzQjsJN/CG05ImytMSxymk3UKsTJe80avPuf1EZcm3cbEZakbiHKB/UA3dgIUY7
YxwitQsSTHhL3CD1Cr+MKKGGX70zjwcpHsvti//HZ3hPFyeNJBZ03UJDeAmh+Ct8
qClGPFSXkTicNobPS7+6v+dd603iTWSfACKykkYrOAxuiioRWSBH+1GVmuUj7wy4
m+2HiMY3iTo3jSOn5lIndu7t7Pa3yILN5NJEOENf0+KIqaDutJYKxfebFczNlVp+
f+EedJ1VThwYA32wRldKzRb1pDkZNw/xJ0D7itnwl5ZWLhhQIlRtgqwP8lktALla
HzF2sZ1FoMqcPSYtiIZTI/mylY2qsgG7q66HQM/9HySss++7j+Q+cHIt9b0ZPUQz
yvrh6+OVRg9mtKHBrqZQusQunFFTzGq1B2ByK6M+rkxWhEpMSgEsVr35xCC4ZiK0
IfBk6tkLonAQW42aUYPSz/J1deI6YE6qEEwvAEUwMO4wT9OKZHZiKxuf6AWzHcwG
70fVcGCP0RK2iBBxuXOx8LOvntp7xmFtsIt7Y/mfQDhQMlyeK23KkO4UVnIioWJj
wAOG/Qhao8voI8voAqrTU1GK2LbDEkfFpk5GbDcfmNVG+ANSd9LZ601BPgfodyaM
ZXy+Gvint2FI0UDUXfmntPbQzuIAZ5oGIKXNeJ74JmY1xxtvMufHDMXMtvkzBLmq
ZKfGOCdvpnjZXjg9q9LTZ4qVn/BPpfRdWFm0jl8jJB4EvDoOUSYsgoQOHdCYo2Wx
/x0vTwFisAf2VUi1e2O8v23T8PVBEa77oHgbhscgQ1i40iX34ylS+5ktto/mwUSH
lAYzXJAiNmPwpKL8KKlh1GvKAY8boFlsRsn/+mUBOeaA4w1L7fllAfdJyl1dlkaM
ICNfq5/KJEFrgXwZASBwjuqZrxwWsawOyK2mTnZRvs0mkbamnzvRUeIulMJS5pW2
f4ZAWVibIFbSTF5G3HiWQiue204LiakaxSRRPZZGTV+csGq9h2O2leUynWVDpDJC
mFweOwGUPNtZHLHjoOjQrjWz7FTFAekJC/TvI89VVaPfUbiOs9Y7t7/qUQcZvBIr
dTu+TQB2D8sFQPDiiuddPgbkvolUTEaOcxnYAbz8JByfA6BUaYV+/D4IOlpvHUr5
KK5JN7HcBVSkuw1BPXXY8T1YK9pLJc+YiTqZ13U+xXDGXuIQnMI9jl/zjUkqe1dU
W3nyX9+thqBVsz27xSzHUuGWztQHS/r8Tj/BWA/JFjVyUd3kmFOX4IZtCJDA5AnU
oVLYk8zRjVddJIJmcy3dJLgvA0dUue4G7HCJXbO379fSVMp0o0dK89sW7wtoGA+N
+I+ix1jHKib0SE1aS3PzQrQrlBzAK+mCj+CMyUsJGYZROCpp8Vzc0GweoWcj5ipN
3kooSXEPd3I9RdJDKayFNgd5+Kgf8OoBmJ9Q2qusWYnf9y9V1hV/a1LWKLzGmOY3
BSOSnwtGk/5BJFJzfdMvECnBK0b0Z4J4h1w88aVNuHjPsAzPHC5PD18PWjki8S7P
nlwftYuPocYcGNSiCUaQ+FQjqIjyttlVDtBbWorNtimqNC9EV71HcfpEvJbQwmbW
3QIdI3YbAhr/BjZlX4ZC7b/zm2l3StG3WdVD6kadwLJ+jWM4yeS9otA9ePgqSdEI
bFBwEx6fDnR0JQmf1BSeOyvIOZNUEZkWEMUhSttzsIyngNyR+BMwHAsBHcXuINVT
meEOG98ZJUsEgRT6a0SdoIz19E5qGrGRm9IUrJCuW84qeAClyNSIUjOHPEi94oRL
9ghD3apuKbJUbeKp6BbHA95wbVJcxJN7CY03YpjtyG4AZd77H75FqZKeJcYhl8NF
X4iOBHKgSacT47lqfcQwS0sQxFINBues9MQBe6kswWGVyNYcOOEpQ3tOGeMM2aa6
kNHIn380P5YIs7p+/hCUW+4i4+tcbsBDI6OCWIXW9stvZ3JY3509zDqqb4CPJFv3
HVWWn0GL9T4WNb/Lv5ix5YEXEip1GQBiTirrN8Wa4+5y93hL3Xbtq4LPghNKeZ+F
S0HfEZ6UXJKO90t0O/23Dy+p4h6ypp14vpizCBu0KTDLw8u7ubdyYzX6yD1MS4Iq
PHThhsQHsI15XZBwaYdfNdT23tTKJZlsLicCZsJikMxycq/3SAlsfknIYfeHGlpQ
EkKe9cEGPyHz08s0oUvtQ0Vt9Arh65xNndOFINozp01kApCMzfm8x+C2t+euT7nu
Nbbfqce2PyQHQX7B3E6iLmcW+m9paIv+lEIrz2YBMkPiMtxDlMGqKoQMx294r5T2
JlXuaPd/sCtl73F38gdZi9FXrd1X9IS+h3D9+ziZ6XV5dfoemJ8INkD2ZvQnCwUL
118XC65TtdWZJ2vbjhfMWuT4F7jjXDBT4TXoQh5xxBdrN+cyVorlqjeZ4gy7nCQM
Y/su4jSQ/SsVHpt4QHxbMIRTxZutUxW3W7628gZCFOe2hq/3PWCketCg5v7jaFg+
jE6n3cgPwyznPhah6I1edQW2eqxu+rV0SbVx/FDBZhQWZFKn6zEI3WAe1R18rLk5
QJR/CHp0z/9eVC04JGCQRDbeWSg69ySurZK4JpSTGJbsnjJsdx7Fmk61JXtxwCaw
BTESaY3+MNOTsf79pC4fit/I8aHr+MOk6jFV70MktQxXPNvl6Ox5JVSBj0P6ZUK1
OKW6py9md/dl60vHU5IZN1bhQIEsq5WkZB38s5DsLy/4jOMAhJa7QT7u3wIEw0e+
D8tCe2US+4T9CxZ7KyGnIslA9bysHfTpZ/nFsYpy2B5VZyYuBeEWnqBxHqx2ULoa
LuBSsmbqolVXAwDmUlig2QniXXmHEHBoaBjDN7JaF7XAef/BRXnNjLdGwh2m+Yd6
iP4nSEWgItiNB6uUEHzy1rGAvpc4Npu/jCemNk6XYgbDcpIphB0Yz6t9e89ALV3V
Srvq+CInF1S0eqcM+4RbGus0tJ1why1v1CpIfrBr65REIXlIRQITIj+JCIZBr6b5
/nLno05gmQcy4/ofZAQxbJPkAQyu+geieoASVQyLUd9tracLOS0+5CWF8Yb5TTnQ
s29wU9dQcLMFC+hDuszXwBzouCNjJq1QeiCiQQi+ntBqfQmcZht9JNnuaeUzwFe+
jd85/pei/e+h14JOAvC5fsG1ix5z+hOjowZnqZBvVZZRcAt9A4B2bJszli7TebNV
nIAe1+AOKDj22HmAqkJ6yuGW8CLgLDV8hwo6p6VNawQfpgg798OKaRW6JWjz1a/K
f7E/jC3Jm+6tlrfPAOxAQfwmfsh80ga11q/7k7E5LxG9wuxy+0NLhCl8URMMLCGh
Y+7+o4+dTum/d9P5j0MX/QwrPiYab+SeGlLslSdJs+yehYLtPqJGMeIXKH1EY81s
y96pwKM4vjMCWPki+YbPIzKSIGj1tDfldlJfEAJ2DgMbPN+zG5WCeutsfiX/39dE
G4xCPa37eEgGsM14axW5LDRKBIHIR+lz0dDiCskUNXPko78B+hYJm2ZM5GOjvCZt
NlJ1bKB7gIOr8YLxtidMRzdPdrnVx0ogG7diM2FtAAe/w7qCjzrpMDEpRXllL6Q1
tJQIlElQjT/39TOG6my7vPve/orF9RyfBKHO+3+DqeJSNDILhem0KXrhmZOvjyKc
LsLwAgUjdO0HebLhWCodlIfb1B80/pJI+fYPg1QlIMB78ZerjDs19IK4LeDW5px8
2HQpGKcNja7RTzjb1k00lOrk8JFifeJXK4Z/mSufFJjvEwjI74OYOrqSlcJijN7a
FsZtuvRfjMwPuzhxfJUvQPQyGR1qBp9s4FYfgVGViEJABP7TdMOxKz0Io5FHYLzS
HQKYXDvonW564U0k8qBH7gGwxGazQhutBup+6WHrsI0ZdrBMkrA3pVllK5Q0XvgK
/Ip2eBZfajDaKP9Of0yPF8PQqg3p5wzOIYHsBy46QgoBYboRs1VDRqKnbH9nK+h3
vTcOe9w1GPY0ch/qkMRVMcLwcgWspi6u/0M5S+pI58viAxesWnRciwBZSqGF2E6Y
0IllN2lDk2gS2pzbtgG7e+buw/+gGsarrVAuk/pAZ8Nv2qAvMfodlMYlK0defx53
MIBauwCk3GiRvvVSyz9FqZK0QPK7FxAhkfjsw05ZdUE0xDh+ZJ9LyRbGfXRRECQz
XUcxDlFst7x55SCbFxQkp4W4qOfD8GHX/3Q1Cc62+9VOnwKasQCCqQ03+44SXEEA
UMcJhfEWH4jiPnDsoyiwqAVC2dpaMEQCP+lBm9KeytXqjyVKTl5YdWkJ+9pcMbg/
yFAlXyL0lQ/q8pNjI2LysOe+rPuxDLIU2Gvs7VbiObuujWoExDgP/C0NilQq03ZL
iO6GRRnkmaAfQvVzIDqY1J4zmc3XkzTEKGo1Mfl2yShSDZRaje4i1c3p35nag3gt
t0L7C9xxj4c+aHi6ApZYsjuYMOsuIEGj4FHeSvgArIFGIgeXgc5tJSWQta4nrvtR
HqT2sAcXy3hsy/uOK85PzwkQTkySZSf2YPe0o7PvmOl38DgqcD7cxLS9nYtL/bEs
SUbz2o2ZcUUbHSZrETEl+4xaS7CDDgOBmC4OQN8fZpf+OcpLA10U9BNSEECbjyDU
G8fnvm4aXAwuS1kY2gVFY4TYRwsrhmG1FWh8+oomp35Yl+nBKoGJqIZwbhdR/3GD
3WGNHMT/sfSjzCiK/qbWpDPtN0pJA2yJ+3pb1JtyRIzotLuw1Djj136HbgCqqyh3
1We0x/rzZuXJUZGBKh8DBz6CYmaDBr+fI4+Bz3uGsBANkkNn+B9FimEOcAGfRMld
ASQ9K5Jj4aA0Hrpo3A03eaVMmVsEQP/oyd+O1eStGvdg2jJ4LCCLGBjX2hDnUdrX
lrv8JwJLgw1i+AITw4SMnyr8kzlj1Q2BeIRGkFnHW3dTf9LzjI1XJDs/W+yVfq7M
od6emJJbSfkSH1L7TWgkRRE2GlU1wDef5dp/uRoaAUFkq7FsDtz7nO4jRD80Xoe8
URnO/azG461UsKb0H7cUzy9TZ/H+bO4k81/e0e9aWrds7v0tMda8fdomn3BfhpRu
Z8LPCSkFvLOc8lw4uqHdMfc0FRqy7dsaufI2oRmIn1CXWcv+xJVytS3FMg0hLDnZ
STJuM+RD8tUPSYq04fXjy/lQv7MZvdketg0YnUGQDqb8Ml21KCcKornqyt1Qnzpw
zaoJXetB3WTfFLwDbdAJgEpPu5WIbF3Yimhj48bpxfxnUE9AGO+EIEFcm3iyXpK4
9Z+iwiMpiDcVlnuqq7wYuTMmovyS+4un/c1V15XIwZyBWBGyqvI73cOGiAxVc0J0
aW/QkGkUn9orrsQHWk/KzIY4EPaKEYs+DNQBCwCUFphv54udwfzxlV7/koy/T49q
yF13hZd/SQlKfscMMR2zXubs3/vVSvdS+U8XBcQX6jvVAX8FTMCWjoR3I04NRGFw
6lq9VWg2oXsf7GCdqW9VHkiCx0QUC+oERo1iNR6Bus6tMUL41gFQ3V5usXynQy/H
pUSyVdoNlBvKZkibEmIlAGXaEbSb6udKioHWV+HO6T4d3xfa2JYnR04+Enz9XE7K
mlS5WkAOEHatu5tprdamhpifL5ADMaJaCTsZKElouV58/GFm2/muub2+Kz60RRfW
ScBGEnhvI3wLvZILvmKpPZ7mB61Gh1QBE887XwbBeisaTrwOJGAmJLQjHOpnCt6T
35DeZFUv2eVxyHNLmUuguMpsGJyho90gI3bWDDFl8rusgm96vkmizqzsQyia86S8
+jCmXUr0C95deOzAR16mMmfQa7KdfC5u0efWoEzV4juKIA4aJ3eCMy6gF/sZNwzx
cLotLcoxPNdv+M4mTcvT0A2QTff32Ecjp9FcE1DefB0niB943GkEdZhbzrj1lkl4
qqJIpchUvuJ3oBbKPP4ZEgNy2+T6RFhT+XYQQuoKQOOqrZU2IXiXQqWf9D5GG/IH
fO2adWnDuAZgi1MxEeSkPWswYkwczulcLHlA3rLx12ng2MHA1dOT/HC1zqtGFQ3y
FsqSq9EXAZWPsdjg4ip3jUEIeVJwYml2JG5xB0lLbkVDXPSGTQgyurKIpiUrLeDY
eFtIvz3a4F1QI/6iCqQyO43Zdxr6EVRTEqKTLWbIk5HZMSCM94pfLYWMGGpup0TS
pIScrTKdnnoGkYaIY7q/xpHn25a0VGYN9mRlNsfiMcuTUxn5ND2qjEpM5C6ie4OE
DRT2KxkxebiIsZA6Za1UjKGehDNypWdoUI0r3HQ6piEQ59h9Hc2S4Xsp4GjbhtRW
Oye6RSwWxHSczSGmo5zx+3kwJr4N1HkrMTqnTB20bdadePUwVovHUCVysGY5g904
iBznESlW6J047iThwKGtpE2KMFLrv67OOushrhIaOqQW7fWn762Rh8pvxzjla1az
wGcKzWph8JmS0zWs2ao3ugBvIYOYx+lWQnz5fbfhajvtHkBvJhD619P8VOZ2MNoM
GwO1L7ACGmapxRnQP6fZx1EHVC8gSsTFAf2OZXf34KN7D4SECAcct8lh3oBBEhCw
VEkmaOpYPF6SegGk8EdKkBglcQ/rHo0sktGj48SKiPeotBtt++3IHCoA5/oBNC1M
/aXxmyOI/iw5Wo0YoRBgwtgO0C8kKx3jHrWjhXMfJ/0SjBvxVogGS7dNKbJfZbSY
NF57T460dZBAFjZHm3cCsj6LTSFYWHILJ+JKa1yiGMK6msoTRS5P+oiVjpmWKEC3
QFL/q8GHCYcECPZryKKVXZRh7meFBbjlaGzNFhsG+ADGYVKnZN/vJEA3V5R8HDMl
ICx00LuMnHfQpHzGngAq42Gu6iTZQDUfUmLsyyaQHNB5a4lwb1IUF7ycl8D2sx8/
+eAEpDBhoPlYvM1kLLoJePb6mJnQkg2kyTqeMQKeQ5WGEc9F0B21t47+jAAKdk1Q
EKhflV099qxQxuDHL5g9Zj34XT6PscE09zalqE7lMIyeRiHohOi995KLZnYLQwxm
VGn0codJ26A+inIotIQNMyCanj3TxvTFcP0A0HxFPw1JKKZGs7ic5S21w2m3nZkq
or9/eaYUzKR5XUtbFPHLwXDctPsVnPgv5lTKPmHJSdIWBs02+DOirU5XnQmMbz8h
uDUWobV/TOJ+Pt1XOfTHJkgYawl8bA37xCguDEkSKZhVnaIuVd03AtXB2alGiIx/
tB1YOhQZxZg7Ku6xZVLwjqb0fguMeoPnSRMpEvl13s8cXG76aZq0lUAOivdKY+YY
NL+7JhxrmpGHrJt34F0FT7ETGqxLIWXxGToEO91pnuwn3GVmdhMjqa2smTSN7Gt5
PEgQhM0KMJDVb6uCuzJqkKVMmcxfA2zE9YI5ypPQXKVOn5gz3TlmYAZBy/G/6Bxt
K8TRJVN7I3AuUAeYhzGWwzFApQVOMqmh8RXfM8CDHGjQ7328idCwukMM/mCO9BOJ
hhQ51D2z9nfA41B/KDuv6EU1R46OKsesZBKXETFoviajg/EJd+PV7IBgrFCLTkks
4uOOZX1vo2xIjclkxDd+HIBiX2Ukoi3X0WjI5tUj4kIp09ZLP9fSlD0DdgYLpfF8
8nxXZAocvVlk/6scC4zfhViyqt9uhe+IAfvHTUOSHoUmKzC2Mm3kVw4vTPM8Yfep
EN3Ok9gMH/axbvLBVP6h2TiQhploTeFMDrg+3TAshRv19njqzFVxIJh8+TDHuNGV
K8KIYt2Zsash10T2ccXqYUNorIpoY+iwOalcxpea/kgwyBCLr313UORsjLU9TVsl
DKFHYtsyuhvp2ErR1d2gF1Mn5iudmAAQP/8E1zWva7xg3vXGBw+Sg1Qmhd/up+K/
EPNht5HTBuco0nsRK+EfBuIhBz4Y8HgJQD/HmHawRVdgUF5AEQLQxhnPKPAR7QIo
T9Xd+JX6NXOsfmqN9L0Ev0+hwkbd0eobfrW/qDDwCtBIo39efEsF1HkjZCL05Z6S
URVN5l16qDGORMqxWfUaY3cPG/EPmYhgea2qidryAI02y2+sbIgKAuwuHBEYh+QP
qC9awa/oldmY6Avkk4/KsIQY4ag8xpsJGwjtRgncG6wK8+sTFr2WUyjc3RB2WUDU
ZvbCjUfZ6VkOBrealsyc//qiIWNMsivikv3pZ65euSfz+gW+SskhLT6SLJBQAhWH
3M3zHJPFOxaOfHLQwQDc4E8pRKG9rA1EOYvAiSlAKGyXe6ZJy3Eai8LWXh4WoP+3
uYxuGYGluqYH0dKJX2dbK/Nh1hIYCe6sU4QxO57rPZNtHmzLRmDq4lf24d4Z/6tu
9gA5FxBsxB+F08FLiNtLZEZYfDXrqPK8L7TfH0qxCZvT/RrBnGlv85lI572k6sNx
PcuFKFVeIP47FuWaJJT0rRyEtpk/6SxeI94e4Zh5EW4oHyQcrK65+1bcyeYddpD0
a1dGJ04837SByhoRvXryl+NMkywfqRr3VNxtIOAM55JuBfMv/HyjAGK9Fdn8ujus
/2es/GCE/Rwcrb4qTTS+16jJSAlblDIL2RN8nS6f/YVulLrBz1LrbnlqENrbZssE
IS8psa1H1rHHzs+j9O+KUNDIQtKWiRL/OX5BspgzO3Roh2nnRf9uCHldHvCgz2sE
WCIs59cqx/MPPxIyB/Gxp/3wNKnC+Ilz1dcWSt/kS5EcliQnbmxc48ylvX2GNIOs
136Hq0N3yKASYZql1RxFWNtUcnq24gB7roR4AIP/mAtDK3Dkv8f9sFR+XNUynS73
Tm9pCHnr0R0685/0wEDbFFxVJ6ckIGngkbvOsGtG0F1NeXaUgIxdA4cxq4fEQ3QK
TgPTPa+wFkeGuttOrOKFra1/sJYtgAPGREX2D4mqg6EavJMAv/LDU9Mycq5b/bxs
bAmYRVjruqUVyv4StxtXKz1cV9iUd4swT6UaAokSZI9pVUYoeDR9cEe1rFujzxjc
0QvbQdWSCRi3xe+e7ao15v47BPc0atMo/9XPHACdht0uQVuBP9ZtjPTXdrUcNmUe
Mh/hk/jdvdU38xq3xmP8YJ3ShupDgGGxRKMVBeVUbMgBdRlvfUG/G0Zb9gwAO5xz
78aMN4AObbFxqNbIJusHKw+hVPmLqjqwH1XMg5BAb8NGhbsUEK5HmXD0ts8/W9ka
lz7dcp3NRwpvZ6lAUX97cp8H3TnDdusilq0xFb93O6gV7xsTWuqkfr5rqaFfWwGS
d76AH6/FV2izeavbZUNlMfmNio/1pDfB94536ZaDmbNRIcmQ8ME3a5l1sbBysozL
4XL6S64v/U3oh8u1NPu/NLwvd5iMI2j48UyrXo5HlO5pPFFytyPqcEY5A4NCl/OW
WB6rXU1oJQ5t/ly99aPxVv4G1v1EnB9fHtKxzsxz/auBSlslvvVEVzLzql7iau8k
Z3ivOvzjMPa4t9UguKuDk4DnsnjvEkH1/2HXjZMmWMu28i38jI60nqt+oxVO1y73
C+5O+Mb7R8oO3Z8nAeVnAk1IDHI3TLfjSj0W6jAfm87lwSsSViuM/HprZdS0sHAy
eFSUytn2xrN7MIEaMD/epk5/Ii/RQSXRnNbjsqEWN2joWDY/xgCuaantFzqcR9dE
debpZ5S/BbZOqgn1VXTYM+X8xOnw9HaLd4Q+2RwksqJWbl2Cc9uNHdSYc/cPdMdt
/vLR31QjQr6AAGS3xtjbxOS60pik6prREr36Rxg4pW13NAN7k6O4Xk2aCy0XD3f1
OexmeHKcfL2rHILmi6B1GzozDADxfkYJZ5sLOK1aAumetwMd8EKhxI7qYG5SMMbU
AA2fh3SW68YO8S6J51XRjaVA+tJb/LDb9AHXjbYheadmIU+VLwtnvNoP7Z7gicRo
YploA58B2PgJC646P+1shTS3acIJe60pwaS3QZFcM9VQAnI5ipO0CWhNCzmOQ32L
crJ3VRfskhBZFcV6h4HRTJqD+Oq9aCK6cosBym4Ik2c+zV174cn9B/2twzYWmaXA
S9Elnk/wEHw1vDL1KzisBCmARUW4+U6T5rytILNp7JvnpH8IPkaYVShIlCXCsvmU
eI28h3CT8wDVlZTSgHHAVD/AXHuD2lE/zXTk5Q1NgegRperQJrawJnAI3qZtUuGl
3ZUvQPTEMNt/JYzw6yW/6LItLhEC0Xa7NxlQ8QPUUy5DamPGSSkjljXd4etoEf3I
7RR3i9zlUyCIoM2m08CtWA65PiHX4EikM6dBjsqRoS6kwJBTfNw4Gre2aSemk5UF
kC/jmkYaaXGf/IhQqPzvAA4Lh9Q3oSGO2s35jRG7FVZ5/20gSqPg0JXXP6uVd5tV
zsVQiSNfWgYaufSqi4PNNyixSJDnEMdmw+odqBE2v7EJjjbFU8o8/AV/luvPdWk5
1J6zccZKCTBAFFEs9IyDoczjF/jvBWlnl0Y2l9bhbq2zM6U5Kbl01oyP9jdlu+EF
ysasmnjNiaOCHbzWW6RyFf2G8pZyrdqlptB8+PMkj6y7tKCMV61zJH0GYKYtUK9o
YU6VvTtJRlMSyBixnCKHQOlqWaYTsnCWd6vqUZUV2u+HKAmk1toeSBCke6GKjCLU
L/G4LC7aHttscSWBVXl4FzEWh+rmJmn+uscOOZ7BP//KRQUXoBKTyLyzC1YK+c6Z
VG9Taj2u9QXuIbNlHaO41Z5zFVO1zRDwHNSP9+uBtuBli0jQNnl82mq/QcQCXVGG
5aIw04+J2U/+b0aatUS2zTIeRGprQKSvOgEDf4vMfepG05042RUq5v0jikFTUMpP
Rs9r+FFQlG2HxMW/Slt8zleTaO8mJScu0eF46+8sVYE4RcdozW4Fo9PHy7ZVA85R
X+hPwp80Pbabi5uVYFDjZpN9zPHIP0+Tp8fYWf909CayGKYar/RfNrAXW6i+vpq3
OYcDLe6fEsTu2lPmOfV+VrJb8cnSPP606WPndV63JVMRcye0514LHtW0DOVk9NSU
f9A5e7+Nl7GHEb96/o4lle9PGrOPgL6cp3tZtn/RKKN76eWPV6qkOHrgN9kHZDuh
qHuTpMS/hjLS10TxKYZboA2Z2ew7gZfxCCHfgahmbm3HhOj8vbNJ1bcLjPV/mwvl
PyTh6o8OTTnFPt2NX0rte3zNXwe3jGmGqFCFajxsMLRs5gnwIPROUmodSgp0Kx0v
jnhUFF8EoF7c/tfD42eJ644UaZoUqBImJiB81aPc5v9wVl1gtfp4vBaiyAasP06l
YoYPT5Xrfmxgi6evplkUVcjGi3RTQ/zCpMhgQukIlT7Nx4NiJxEKFK2QhMXMmSgH
95hqc/RAm9t6YuwLoDlyXOnjijjmnIwcKXID4XNRzNJ/jdvbkN7N7q5r8pNTCFoC
A3IWXQ2DZM1QITpAjSPcjY7kca9fbwTMfwWeahyQOpuK9YcC6t39h4KjpKTbk9eE
IOV9xw9/M12cXiU7FIIdOiFMoOKLXCQJodYRqWPNC2lSNiW7HeGsndhPX/FqbG+D
USVuzXcLmGyUAFuH0+aWejcQEQIu5ZwdXSQ/n9CSB3SRpr8js1YERLeLW0klA94f
63Xi2x7V9NY7smgShKw99bUW7H12ktEAC3iR17su0ArXYdNxEWAL5x72CRWaqRaz
6pwxd+PUey8Bt63ksjuOTjcUIS2lcvdFMqACwxmoCjEogSpEGgV8BmkxrcBEVSti
RH1EYUGYRg+AX5T9g7FjrWxEZ9luFuT5HvGVKvF9QfLdsDiHpC0e1el/kMUktIsl
SG6aDX4adlPEAsw8ufJe+YwleDb13EhupqcjxJHl6liVzM6Pof4i7AbwwIm95Snq
0njFy9iiwQ9/H//PZP6rcgEVJgMQnViCZ3aR6jqW4Q6troOmN30l0mtdgBT4GOco
vogZk1PuICj6v6b7TQctChTDXnbiezMRGV5zStn+3QrrbUA7+LvQv1s/Y8Dv8m8A
9UwEqj4YYA0WT0wzzLJFzTJD7Ba1no9ll5oF1sdL+ef1w7ato75dEHHjEqU/c/Uk
tKK31G/ULLsnem4zQPewW3wZVkpsZTehoaM0aYy/OSjvJ6e8iNZLBOojcekJSfIR
yCi6e02rCWjc0xHP25T4XI7qo335N/7K1cnkT8xaTbGwNIiHv/XaOwuZC4tHIu5h
kGvgElt/Wf9CRmrDQH5MFH9HrFdNPowhuilyJPZ+NwM6WLBxX8kIUA6ZzfKf4TE4
oa8+jqUCchkvNNXOdh8Rvc4lcTKYK+rrOZUfz2XUikhGfuyKwsjj/JEhqxU6sVZH
Ej3aS95MffgE7srVssV68uDRxMSWyfQXfgA12dX12U+nsQ1jMRYSxE12CTDmX7e+
oaYSnsGI3+Fpw1vgxXmPUmakeWcGCwE1K3gDohlHQwPgeAvS5ruAo2vMeRtNmQ04
A5bk2KAlU/aJqtM/IE2+4feeAIa5CnfHr+rRYAJB3S4Uoydc9bY055/TDTX+w90s
jyPc6niv+d5kd7Gm/uZlZwy9KnuzaDQx2llftjvsZrr51KVW2H2EDvnz0JQpcc6U
RX+HN+hcDuT5YhlhcMu9B20lxtvaHfB4mbIfWSj+53tu+I+koGFLosGy1UgdKhHq
f/1jkRPxnLEWPiD8btLbzDZpqrKaR4YdYJ4qxDi00HNmsiLOCk7RtPSHzlkSYqBX
CF7Kd/OR/gRErcrs6q36Gply8IBEnIPc1WpUK5hH/hfT+i7JjYd1IXGf2rV8/t8z
BjLYK/rbCC7UTSHYetrI9b00bz2TySPhYC+G5P9/kshusqHtgZXr9RjFvrKwElYS
e9P8DipwIi3sX4W40EyZTHqrifYrAXd2bS6pfA1fbeDtRVCcFhM1UP3s4nw0nexf
AWbYkPmdyWUIRmmZ8KuYVYOYPoNmHNkEvWlUAXL6lt9S83tr2g6+yq6g6lQbBc8a
kA8alEMHx0LnbKBDcs720qYugZjwx6snlYRVRetctmfmoTlbf1+IPNvXB87Q+iDI
/eIQu6qcU5p3IqDk7f9vhfTgW3BpMrdP/cwPXsc8IGVA6b34XFKGm6RmMhc4LRPs
nHnZTqCGTDjzw0ZRvGqa7bgYWH3mxhPl50JWM7lkQBZlLlqeyGvtdMQ0XTWZJNhJ
KFVr086At1Z59LhB0g60/uXErbBa666rqRy2F7e8MBqj6EVng6IFD+jw7nmvZ1IX
dDCToIa05SXqGSmnJbKxdYiRTy7lETlu5ayZtuFTqnMeWQYr2Jl20IkZ8a39YLfv
2eqpjQoanvLGfm3D0QpARipaS+PXfxPDHlBWOYHGL1F4pDKmZOc3+aiPKwhpambp
e61XQK7FJ9pju8BB8FuBUG+dGEvIAXnYPzhngIJal6LnpabqvJrHPSBkBkLOHC+m
7I8aDioXHPvvy0RaVrblpyg/2U5p0nGfvo+uBnyyrCqjFzm8be3so9x4kJLjC8R5
tBZLiO2mL0+ariyWhceLMbFmN7Qy+bX4j5kzJ4wxYsmtyoYicC1Zlh+yg2Wq8bbn
OExriv52U7/1m1ALrW+/GEenUQT8ND93Di1Y7e7/Jr3dHP9ejbJ264APZGgmONuP
pfPKUSzQgrlDWkUg9h9of5bGS+FRZjIsmXNrbhURQw6KpFZIwQ+XxLNrhbnIEWsu
snMIrQybNUkKSp//iXFAsfwsYc3VteWFzxiLhDzGZ7T5V0o7Skpgi5TSzkxHKz8r
BLgmqSt1oDrGYybLTaARDWa1W5ArJOXOwUMSNSLCZ4Hn/99S8NM19/sYAvKjIqIv
IDvQ1hJ7ymZ5G/A1PUBRMfAiOyilzWUHfEcKJAqgOzfWvX3gXPGNJZppXac1ewKo
b7s7yLMLMmaOt1UyAb9o9fOTwQKEft21zhSNKcFdBa5M6HYQnJVpMJi1ggdosu51
8X6farhtmRxdy9hiJSpLTnKyT3lfxpWOxg9UDSlrP65YoPrwIJTXYLe8+nasodtg
UO6V3QyRvfIoFEz+bE6h2eZS1vWId9vavCEm0BERkxRGiDuxG9rckJ+QqggULtlx
3NEDf7g0kLJrO6TBv+XfCHG+Gq7Xp0B9QoNqR4lVEO40VL+2fs7JzgY4LKq2FTgr
qMlzIf26JT2roMXWuLgIPS8nMCUxse5UtlrHXlJxKdQPKica9o9bX+HWsTbsmk6e
8pmsOJzd8v9GoYdId7tt08CDICYSfYDwSwnhv8Fetn7AJB4/A434m6GvsJYXQph+
hIMID1ScL7Q7beiAGWsOOfzkDXW2KTSpTMJ1U6805D7+6xGZqgyJquTfpMm1k+vp
bmGW7gsBCdKtoDbnXeuD6pbSKUpSMCErGXwKLeIDlgCXwy23S3rC9RdBQXiVq7xS
fEKPbiNP9ourLpdJ4f5S0JYAA0GmIKNzmN5+jK7+g1QWSqCk1bEN6jH2k9sOHIWn
IyqCveF5fR+dZJa6L5rL/bFPtHCYQT68d0IemHKHLNSo2/rAj7V2WlI5TVKlHREF
dzvy7PfsyCtzQC5MPGqBcS9eSXXv/mr3jEir5IVWIyhVV2MbQlF5bKLut+SJmGPx
lYn56Mx/7uJEyIFfplYP8DKhwDl2Oeqw4BbDYc5Yxhg74KV+y5f0vyQyfc2+6YVG
/kB/4Qx/KHzQfX5vANm2p411eP6F91F0a7LN+xUAh/ZL1pOjM3Idosu038YQMQFH
++X9VMfhHq2l+EueQMEaaftk5WSiv9aBmlQYr+tZAzG3Cb6ibRTjJvHI62LGHPvI
SFWWwvYXq2TkpZm99KcsxvP9IDtqNnZWBf/kjoHAkLtom+AiqNv9Dl3PHyO61vAh
60d9t8Qm39hy2DBGDxPm7uUHCM3dyw5Jer6iczk754r5vYcSxbgGCY2xr0SmU3kD
dgJF6EvazZju820RVAEvLOdRc0BGnZQBTbGTy3do0OIutzc2UZGINlJy+jy9O9yM
PMc1HPi3Rp1DrTmYAB50eegOhF/iwGpmWAmXIETgJfZhVlWL+6IMxzR5VZaIswO2
NLWilAQfwyTjHgvXfI8n+MNd5cdPS8ba92aZ9SAgHnLiTlMb6/3KUW9dADcC3BGp
1Ug9Q/vZhLjHSYOn5hfBWXEaMbY9nhKRWRqO50V5Sc591IqWWT3DaeSGaYSApq5t
LdLHUlvZC25i45ZnHN5r4DElTze2s6UdaSsxqi98XxsAU28YuYrF4BaoFjUE8tWA
q8yyZl7HO469YpEQWqqwwwTD03PDM5mdcu2V+cxps4JNPHBCPwfEe2GHC0DR+b5j
3dwJgeJVZ3S0HOtPeqVgUq140zr8voSta5hUu4wQ0uAdFsy+pC4cPU4eTMOa+Beh
Ib+7K7Ic91NEuNh3WFzsp9KggfM7clMWE+XIQpuZD35Mv8BA0Ki+DVbfSewWhDgu
dAXkpNHZG8/rOaEf3k4URbJEMeUecxGYiH46WME8/qerocJ7zctzNz9kAQTGAM1C
ZwLIXziNF36EqS61OAPVSHnDp1pGK6ylDEH8b3wOpKcxwj/t/3ubsyZRzXT/eTyA
PGDKpDwouMUwQiCySZo+BDs7fUW45VbJ12cAnd6B+AIRDTTB4lOsdI9OXv+DqHT2
qka/8QQ9ZgMOM+e36gcw/qUwH5OZud0nAGLtmw0jhOgdudKG6G4kO1cLqq956lCw
dVYxGIUGs/SOT8wMRVgCnOaaWtVKTMoj45vkxEHFujx3jn49C3dqiO96quNNAYUu
g7zhgB3RkzpmAP0jP1y+zSEi8SLzIBZ0Eqzj7arsFC3QufVsC+UpTl/ecmUH3Bg8
1EJsgxb/YEDn3ndXwgkXMU7gjTSX52ANcaYWjpWSp7aqFOV5vpC0fo6c5Wpisbff
SsIF/sjd1lkKcOYpCnzJh+E4qSzjN9OyaVNjhTe9vCQ4Dc01gx2PUZGLHZNxx0Vy
OGjTHEnr6efJyZ46AI61Khh72pgkdZ6JE+KqFFu1+aeUqJHNPIl7XrFaA5z2Z9w9
qI8C6/Zc+MgwIX4E3hYOiy9f+cVtbW3ZAEhAqpikCwC9KR56epPYXc/H/6mZtZfF
piLsAax1c9JEYif1AfrhFlCOFzSnul45HFiiqpUFEWmP9Dc4PYz7DCeeKOFSlPP7
FqShsq+mFnFwRU0/HJujwwF0SEIAR8rHCfxJ+YBebfboY/C+sX6YM0jr25RaWGgK
UI31hPh3Mn1VUsRRvqYcvPMcBLzSLVpWK+hrEJWdwA3P/zdZ0zKQAN59E2EWywwt
U9yRluz38bRi4QwsPVwhEGdNF+0AxPQABAdbdZB6vw2SNzvB0FbVrMeNqFOcP4zw
k7svb1wLUjAcnq3lM/7TNQQ15YXXtZWvX3KlRvBddeTnZSUkvtPIB5LYDPDpswva
koTmOXd/YQMAgUwT79FA0olVzeYvC44V6T97hb7AdiYoNoCQvRRYy8mzRJxTrRz5
TibpEl2fk4Cs3G7KzB5lyPytLEE+aiwFSvhdVfL7bzpg+9ipG1QpvbvqXywN1OF/
9VN2C/u7oFqFKjgbYErbteLnjxJff5Kp+PO0HnMBTwmi11GkMf+n0tUuJ+qBGF54
RP4dghZh47o3LE+PPUOprVa15KZQxpbWhM6Tvqd7R/krStUVFYAoaNe2cJrYelLP
YpB49gDZWAWFxyjSnMIHwINzc9T7cGQSQhqDWV0dZnCsBLGJIZ/NSw4GQFZTMDh4
Vgt83fy0BxNS/RFXspwRuWwitbsTEoQU2eFqBSoqAhBUgrTkEgAsHBF/EsadUiUb
C4tuYgIIX2+kuejvqVD3pcYEHbDW+VzD9cgHizygtZbgU6Z7iXeMvIyDA7sQT0gL
HB8bgbFAeIuPNKWOln3Ll85tLGVj+6grdZk0mfosPr+ynaKJH7GHaXmgyQeS1fZU
/erK4NDMbShPaT8AyAleOby/CaOLCnzPSU5hQ4gm99m4MOrnGdJ6ZqvJup2D0ZvC
y06CGqwekF5TFee81LYgG3FMUr7A2dtit7IrIyBEtIeSIKsgsfKpVXlxQzzAf5mQ
ZkLRdb+DlVuJXarlLv2/ca3jCQ8H2wPAI9dE5F28rq5CdnutLVASHetntzXIkxy0
9697cfECdY3me98E0Ja47w7FvmGQ/XWrBWcSHQnvHQ2mMn8vAZjogrhv/1MRpC6J
gNYcWBWAGUK16z7AyqBNiWPQcq0CJ5de7TIf5IjmYa0RzDd9C9JsJxLjUyXe02Oe
dKKeuTg54fOIiwaby4ShUEcmCtIxXkeqOwlTFk3Jn/e/GDKK5xsloDS3Rph8yd76
ie3810CfqPieuuHUOCBDEfB1xoW4RVvYoabaW8faoFkuvhS8sAr5wcGgHUVm5jM5
Qq11HpebB2OvMTUYEXDS3oKsigGP9XzrCiwDtUKuCgR4N3ysKfHIdj6F8KCK1UFb
npban9KIa9SlUSQwl7V/pqIte5yBD5gs3Xdql+oTVWDrPTiUrtVmUAffziKNXJkI
TIrTIm5Zy8aOGsqvbCo+n4CWfSSLHi81yvGshOYCp4pAZBRcIcwpaV0OdwzT/N57
/IyrwJGhbmEcntCbfa+7uZO1Oq22YY1RXyYoEu8F102gdtYU72N1wv4gUNuuzzex
+1iWK8+JozftW4BKDRyd+f2Ih63QElPHWGgj+yrnKkQlVmpBJjtrrR81IDB1/phK
FBtl1MKUCtvpH20xfYgC/JrD5o8yzItG30ZcpRWwxGz3wqrLrvR0m+Hvxu3EOsWL
DpEjqR9Pq9S3xR7RTBJui/S4Ig+6fFFZeknOl9Oub7X8jDjTET8VC3KHFL9Z8QgF
mf2ea+JUcqQ9pIaAm1QwMNToUP+NgJ290mjZVXncX/EgTosZHm0JivBxcnJP1NKp
PNHh3g+dVl39uQCiYZtNT3YaDCJWzZiVYUnmyj4Yg3kW9940gvjUlpcM7C1sm/9n
A/o90aW74UZGqTQPt6C6uGzeW1ik016cjLhEQMy974ZLvqDXku49BpZpYk451Ygj
IHRNsYvCGtNNe1qvwZ3G/nbQHzNrJMi7FUT2LjrYq2fC6qvDdkcxaUc8FzX5HKy4
3m6uGlbBoDNkCrKbItgnuuYBVF++Fzorl1mbVjJSqgZbyRDpOYg7GVIRibHmM7hO
HnMHHIcutP0zy2LgXcOk38o2MtTTmLma+U2HEv2Df/wK5Oh1/6VN5o6kb36SZQmW
rcknesqNjmxJvld4KvNLcU7Uoj5hkbLwXs3m1c6VoFGb56ktgCS5wgbkva3tF3/k
ZFoPbWNEa8ZxP81dZOYdmDtsEb/bxlcNSWRHJny0pJf6iebkXhvUyg9Qm6KORLHE
3NHOQa2nGp2BuUNe79x5Iswocrh/+XEFgR18kB4fmQAwCf96YNpasEJ6tuH2DzFo
kib6Pb2GEFnDIEiU9leabtw5ClflsDWHytdkP1IKHYcbLy1CWGiuJQeMfw6Tfnf+
WnrD8tH5GWrAxf7Mflthu6a0B+FE9bKIJ2s3tKD94wvjOnU7k/O7mMpkBslt088F
PiqygTj2aoTqeXZlaxplBX2z3GmAM0rrm6KlecODXtrNEhdvtXSuNiHIUkFziHPq
Uc3xyjHD8qOHhDkhUuES7+LbL2g5jvI4XLVTs3mqOKuM/Y9SO7pkiGytIEW7l4pU
nnikqnqKgu1ysmiuBTOKzRbzdMkMg1YBlAC43u+2s6OUmbwwhxWf1G5XiA9DQtBA
5gnxwh2VmLcOGcyOaDfaHq8+LsV6EmMNlLnJH0dDe7r5bz/RQXyNHzwuAlZqqeVb
PB7Zf281rzFRQKpxMWukj0sVKf04owznAUkWODFIbG1a8l6YdG45gcchu7MVjjj8
vv6IcCNfcm8ZEuhxP0VJLaQI6CqsJbGUXwxhfkuc9GHN0swdz3D91wTx+AtKieI7
7YwcY8OnXMIATSNpOONF/eJY/cVvk0zvdkIxgXoM0hTctEHxRRjagRPTuTT8GlAY
mtdXQ7m/mc+8p3ZZOrElc1yAW1EhD5yDCQXSjeVRxyFIvkTifzWdCkD3qFtnMxWo
jEhUp1i5epwRxKAAINvs5P2WjgU+gyLGwdloSmWytn1WaF8XYXOC1xJGpWXc0ubk
LxPLEtpO3Wg6poXsFxmUT98McE0IdVa+PGsltTZygUHcE9NWni2SviGYPJfBKXcL
nymMjGa/xu3nvCrl5r7Sp1pmgleu40RJFfb4Gvc9kjnrX3RdClELTkfJf+UwsCq6
Srwvy7O6Vj1EqAvyh32OQ5TD7z0yUheYMlx0nRT3qRBV6X8MYcuJVAIajPetakXp
pp6qGm11QfPKNq7fXrF5P3+Pt20OWbABKxZwkWv23KPU+kh9QJk5JHo+GQlT7GbX
rvHjYvIiOfxe8IOZ8c6lr5d6FfZqZGBEWTSPbH7OEGXym0Pn6aCCKsKt2BTVlvxg
0FCxRGFES5bPiQlvgrHSaVBPrOiYAdADQJ6boN9ywXJ9LfQvhcTrAMZrptBa/Idi
oGIE+nKxPhfoEoSFLTvl4ja9NrWsiw+vYCxztlMz8xrwuX0feVWSWr2F4KiCn5xM
ZoE5AW1kabNV5K6rCVJjN2Lp5U4ZHUrK0JpgtuS+srgBDX2w8c4usFiCqtfmA+P6
riSxrI/iTXoLTzwhbyd+/cQrI+J5fLqAs1szYA9/A3ADLvObfirnTUYlKG4n7fhr
spMoHxAfTPgycK4M+PRaiVc5b2YSRimRvpgbUtvfUS+RgZovuhfJT4TIHtCzNluH
o9N6R2eNIPVfDeLcpGkM+GmjDiOZkjvpfw82gFlxpi0HWyvMVRGGbaGz9+daB9KJ
bPmAY917ORMsjIc2ng6to3XqTm2g/Ret3yedKyUIbcFDNDIIbnEUp/ZBdv5lRPdr
mzv05YzpOvIFxjzi8GveefxdMqZ28AuedTg5Wp9A9Z8woCVteOr4E27jLNKD0HB9
d9W10Xs+/5pSivGauIk64UVOE4G8sDjUz0/FBcrAskmcH5CPv4/sJW2bC5RA3wQ+
/GyR/5gLGZpWGBtiXC0g1V8l7zIdwhFIpSydH5Yh/UwSglcWAEPCq3ZfInKD1Eyd
CDvbQ7UKtVrJju1jUB+58yOodEmsB2mLTg5W9jpmBYMdcMoVRWINJd5J/5MdO9Kb
LEPCl9tyExelcJpMjkx54PCvK2ErzdK1tkzeapLJdBH+AK8/YEOJfIFRCGHhbVy9
9gWaWWMVgtmKQeHApTjbZOlcp1T8ef7839vxz+sksxWatLDK1cgmrwhJoPsr4/lS
+lCGWHJT2PipiqwGdghYxDuYIdjMVAuMr5sTLx2mPhXFs79I9TPXzXM5mj+wtrMe
jY9q9l1WsoUK2LaV8jq8ZD5fGcgiW/QtvY0D/JqI+/5mWCZpAHAHBpnKGJYP0M6B
xz+a+AEGorv0R5xG2KUWBWT0wex/hfdsoGm4PhLCDrKYUR+CprGQ41p4JOKWyewb
bfMW9xi+C0pTGDiaBz3Vna+sUktuzYfPoFMm0rwcxc/uWYvlIRf0Nc09eAfyg1Tp
jBzAas81TMobHkOdF8KCKeIObwn1QLV02w97/QkwFToHUktKLJdr4Q/Wmd3Byk/0
dycKxWpdsS5/ikdLzd/YjHWuCgxjiROgSuC3Y+Vx2xX8eMA0x6ydF98nRx1c7mML
JeSkddN4Z9k8uKy8oSwPtk2CWgpc+MXKOU22jMz1IIxOsTRg/gZb222m/3PhpG9Z
JTvVknIBxjDnQpYvm3ncFhafYgCk2lMn0xh64dS1eGHlV3bfleck78KH4qPc23q/
sSuUKkoRO5lIZG385sSsD5aNR+g/qZwYCbnK6CCpbPpCpNn1G7jyi9siA7F1Ve0D
0BxLT0H+zXdgp/tTsHfxNzS51wbMzMkqyUDXNhdNfuhaMFOMvfRDa4NTEHiwAnr8
EmdCyDIMNTv79ni45KiHNnVjV2Iyyh8gWZlv4XfoZhDfif4+RPRfsAIMWanCPCNY
jl5Mle6RDQ2WG/iSfSAEOVuMfw4N2OMSi90nFaESF7YCgBnquJVnIJ2mc+a9wtZx
qBTWquW029EZGGO7/onQfAycEmcCCbxLfX2ZqlKtIUW40XESWMUbBhrpn249NNA5
w0BC5iA7MNHgOshLJ+Bppjfaq11JqhbM4fp2ziwNV6Kan2Ub9rfju7Gpy1gYmfmp
3xrh+MVd1baiJetlbIdEnjwsejWH/0bRF8m9p5ly2Db0hF+8mauGRJI4h52+sV2k
jDk4Jry71jniPYiYB10tek6sRrEE2jaBlOwpNiiHn/FfBhVuF7pvmJ2yTGV2gdTF
bofkHhykcBbyQ56IseOEIOKlWibvs5oKTgmoSeFBiRRtreTxBba6E716foylze2q
oa8rtU69lvq8I0/lNtPbQWV6zv5htIVskxbVKgsrQhnY8nkg0yEfYnHwYgAVdErf
29Fxv+Q6yLqNpwXxhu7QXQBXRlxJyROW++ncmHtqbcHyZvnI9zzxYor65cik8F+z
PO1rQ9r7pnRRpQc6WXavgjtof9hrPWHaXxiMoPK+2Z8hOQ1/6rQKUx0B6oOTtAtc
h+1LCkiPlk9FMLB62k/e5ArJaCKJ0Ltkb0QWAFgeZ+11JMScS8umFrCT0umIljb6
fXMRLw1Fr8KmlbMKQqRx9QJmfJoo+FiElZnComEnhdKQxh/vXJmM+ERljyW8qYJa
bWpU6KYt6FkAt6yCAFgjgYzhNdHOVuM3MzVXKU0Cje5nMsZHmVlH8dt93iy1hEnq
AJxh1ENngJPNGRTKEsovYVp1FeyP6hDv+sC5/444gnhyGOPVefJhSct8Gf+1BAWn
LQIO7hVDvAJAs4zeD87+xfVQ5LYpNrDpSQZCoBtUUlN8AnCGH4vwQbqvqADBTBDj
bdxSdyoMlKv1qD0vfYenYBBHUNo6pY3QO18InivpI74qzlQrlg0mhZjDwz+xgeFT
ZATIRLePAE1/TIaFstovc5bwZCniFtmrCvQV04JJqhOm3tVF4ndoFb23bzSxjBxj
OtDjFkjzW3t6KWph/G60cUqpl8IKUs+s4CZHOzDXwakSFen+NK1uxGVP5e7225Yu
SM/zJBOqOPL+0iTYm3LvuBT6IoSnFBEsuDupS0/BiOhnW4rPhpikFdaFm/jHD2Iv
x4/en6jqvWKDoBVNOE68EkBiGbiEnJ5uD+X/K2KTEONBBwLA+i2/RLGqQhesjah8
1u79vc/gY3A2wIw9XtXujsWdZ06IIXT+oVOHyPWDGzW2VEfcuRSRpnNJZuY5fsG2
Uj5fUTd5F0qcn4TNbn6G9CMowLRMJAYymKQoTfsqcShoK2XOZojFO5xmluCLlzMC
ZN0MgDo6AG19NRmWcPbqROR9lQWXmCsXXgzf7Gut48vYMuTQQHHmwkesLkRbKepM
iH65C5CyjJUSwOtIHNjkgAAp1JekDPxRtyAKFlgd8rNlF6xINHYsG+FH/FuAYqKM
/x+aUsd4nApT8zG3KNkaLy+kQLwlr60tVxene92OjZbmB917xpB78JFhVX6tuHO4
Av72vCVV95VWCkQN+94HBeKW8tQKPnHWTXVChWF7Vedfiw7qzyFpAZ2vN4217Dlw
3tV5P50QupPcaYa3AHSWA3l3PonqkqCs5UKGhL9TYapNPgf0xH/nkM0TNAnX7EJn
PJLMrA5h7Y/r4KZ+b9mJzJ+bLvSAOBzckVitpPPSfxJe8cj/vfi8pKLK3pvbbykF
3et+yqK/STjMnGRk22rj3wbFtq5r3m6Z9W3I+rv5QeFI4QInxZ8XdCIgO4BFjvN+
ww8mN7Eo1/DQpHBqIP7h8NFpM3zfrEtaehzTzS2hMzlKOGnAlymrSTDoyIz6kj8V
loKM4TzNAGxLPabLNi0+bC7Fel8MEqAbB6qAQHE/8ULYVPMc7tcI1/54QikBkM+G
ljCcqZn3wQSx3OqQx/jV2N8FWNF1L0CJqQpwG1M1Gj3BqBAtbB5fZMD7CODjpeP0
7H/xO/74p/gyxEYs2FtkEZhcRk/wgGpTybMOCpH2J5eJvdvQpyBxDVlMrpKExysK
faU+jRgWIBq5cG6dK/NwfveFakCKW9IfT6pVsUrZh7GjtHKuWL6stlF9tTM2x8VT
SzfxnpX8TkwW0xy3hysEB4gPfGz1oHJN+iZWcL0C0BBj2U7x5Fz03PsfBYVVI1C+
fiHtaux5daP/eWv7Ohfly68bAyaimqe+x86JQ/nKuPEJb0NWzTyVE1xhTYVbX0WI
pJacb64FTZGKf7lWCC/0ZVM5L5gUVoB+dBXbxtrJwlmQUvFXslJuJLAU1wB57AQl
LGUXoVad2D70kCQ6I0YkoLLkhs3QbdW+SZcsirERbhtxIngWrhR7vVktMlP7MmJ5
Y9vlM+TJbpOza+yXuw/fi7XWiUsV+AYtXnD/wN2oUOu9DFBVnAN6mbyk3kbiYU5F
isVm6xWiVNZ0eAZw9BgqYkTichiTA5mfTNAkQ+Dj4+GDmYoRtOVufyewOR7D+gRj
F6+2g/vha591A4gWu0rdQCL5mF3zJeypfIh1Ug0yFH0kQsGJt/m2iWTggygfhbQB
A5cBExOVNII+UYfYLCDbrWVjV9ugldLhWhcx7s11zfIQGOR8Hip4obC81Ux5acKs
fziukoAJzPamMAJfZM/p4GfdEgPJnlC1Nx8bSfJ33MXTAN8IFWjd7TJPqWmVqbd5
41d2hEU+GiMZzxmxScUP0qX25g09QIfDfhhRC4cI89TJ6XqBBA7v1+PMLD/l8obv
LIEQx+ZzG82qz3fycrfNorRgShhvP1sEjQaR8KE2QL93xPKJbbWyL8IRkplDqtuM
W1ABLRAhumvASDK2E0UXlom+rb9M4+hfHfH8i0u2mZ5DL3VJ3nL6qJVCaxTBNAay
yhDH14cs+jqtGXmBN/XIzLEPH5f2ZFMAVxnHsBXEcvbNvyAi1I0ixoGEPbolpz/I
o2J7/TpVCxpiP2eNmsOMPSaGcz1rZm+AoxTJN8A1Oe6tJ0A3S1QxujUMka1Pu+HO
JJaK/xNAiLABRsd8Q1mvOKJgz8Hsfkk+JEiKVBcVMLw9kanLcR08B7VHL1P6HuHK
LFiwDZxt0VNox61jXB9EXLg3M7/4PcfXXTATNYpU8/JmcBMLNjsvZGF1GrW/GbgR
H+KlU5evF/P0TLpucYFa5DRM/048bzXrkZJnaBVE3qI8ZYoyikhxyEjlWfQVatF4
J1SRNO1l8Aua3xvj1IKLJgmmOZyyOvMDS+UYsHToIP9dh6irtMuySEtR9h2T8Nip
R3mA1kFa7TVcEyQz+75K/UqdTwaIidW+cVKXXyYUVwTaHuviNRFffMytHf2USAV6
cM9A8G8XblTBw5VGccxXaojQDrqY8fCSMu1kWqvI1eqfdGMa5zC8W59mow/xoeBN
7R/6SPlqr2HNcwo+RXICVQPTbBhwUam32KmBKH5N0aYAOgeZ0xQpXP48gVLWcb29
NFHvLcpF3arrjL3O3stGJQeUhHLJu+fOGn9zO4PV94UOf2dR22ov70ZTm29T1cv3
9M69oydRoZwe0Oh8knfF3/Pa7RKWJkE/GAfgd1AZGEiu9y3Sfpzh1LsKmsfq2Ura
HH0scFjRV8zfcXpDAtHrA95a0NZruR68PYe5YCrJabbDPeo4rTEzQYGl7q7lYfnD
eISEK1cwHi3GAF53s3BaY6+qyPb100N4ke/yek25313IeFHTuZ40YG5mCg/D5mjD
pHnOxYWKkOQSFF8Va602Z7LhlrkVuHuqkf3wp4javwPuk19uzmS4WbBCkhL1QoeS
yXLizDd3t10OH2MhjTFczZFaTPQcPz+eo0LbHvCRGZYUUWUc3ojPK9pyDL0vCqnK
0negvL7joJIQgEYa+T/veVpvOtKtoQohjug2dgVFB6fpZDHYz5jcdSuclXLiwNDJ
r+dIqK7fI3V/rpoL/W8A2rhRMIP42vJqm7XqjFzhehPsu6oeWWdiRXUmZtyPQ+lr
d0psBup7NvTIJ/VE/qLpwgvy72Adm/SUht/XIMKGrjhgNvytzgXCojlk/DJeFi4x
HLc+pKFWRBWbK4HoyHKwAAdzIXgPgaDexdXDP2ejtVSqwCT9oXi7hU7IlHYLOk/R
wsGjJP5SDzKSfb8ljq6SGJgvG0tftDzh+LxzPZq1pYHt5E7L00funQvl2gteKIcu
75Qbsg7273uscOI6InjREjpk0Sm82rhO7qX/ciWTWl2zW8qxyu6SksgA58CIyepV
gKSyF5U7IBPg4xn4pB2tnhgU4GWU+r6EcEWBfkifZp58a9sQt7ZJHJdahnkBLn/F
D2H3tzD2TbazMoewlrxMMGMbVNqL9pz7bI5k1XLHdZ4IkLoin1vFCcC5T6JjccYe
jxdXzLesaThkW/VGlbPmVvMm0GUGi41xcgdsrJ8OUs3OpB37sfg1y/htdJgwdrQK
mI06ptmNl9Fa1BXHJyy1wXtl/CunUKX60OmGtNKrnIn2lnv597JdlKdJ991RFzx6
R7XNFoCfHW+kqsPIYIU3rIXFyHBS8FypwiA9oandnDeS7GXmYyLbmJH4GvIPwgne
QCIlM2Ng4VlIkORNYH9nahLIf2vj4QTyCwaH34T0OhWIfatQ+ci/XuN6pd+IPZEi
ECwZ+PqJA8dMEJfxq0i88MCXbp9gBSScrARHc8Qv+8dIXcD6eTxt+AzOysZZPlei
gJ49YT8f0p3YFdVGjunf3NJPW11SxN3qBQw9u/h/kKO6ymYskI/ecAcwSNCYqdJ/
oSBovL6xIr0YE5WjKBAMuXJmRSblQTdpuTaBp99Grdq/j4FglBWlDCbxIyRkiAaD
a1IKrc2JTUx73q2PDmANaUglnLbkw3pnskU1WivyKrEJr5+qApWgEgQu90nQDn7t
gd1DjmX7ydX7qQWmcz5neqafDMDZo2DRjwqQniv2/P2Q6dT4r0fCdWIO5Hyjn9p9
i8H13zm4a1RJ3yMUZzyL+zrVqJMjsSB7dxyMCFXEqxkiKRD2d+K0XMw1VzESMW20
4RkXgwfNDZzfFdQr0C9H89QbiQFNCArYDqQNpRDtK7uWKdVn9PeL/6RacvujrhAJ
gxf1++4WwfFTH3dQbSovzXvW/Q5zCqFxi6WSdbdi76in/o7CI5pu/pMdp4y7xHXH
/sMN7aOMvDfZKZqOrc0DOaKb7bFlovzmeIdJdanyNaxnqz+zw8fPVoRN2DE7NFE6
kGG1HnQljFWSCp5yhwvmLNUlYJQBAORdLKff+ft4K7ceeTyAsTvJHbytHkx6Ggo2
25RRRiqh0ydndrKO+jQc7rphu5tRPPdF0RFX1q/2cclNMXPodjykIo7kOq/yyMGo
5P8HtTEMH2Xhi6K9MYZK+8UpWfoRnTMcePd5HsZRhK9cMrhotC3PSKDQrmUQKP2L
NIGrudNtCZIf0SRN9eEkyx5vC1G9s+KD7exnPYvZnrkqVFYm8BcR7WSzSzg1Keog
0jAu3TDT5RYmTBaoSTNq9Ns2hg5CEtIQAtD5yCct1MN92mxDtTld4OgWW66w4aY4
AKh2FQuxLmxd1Col/Zy/dObqjoKxNBMSxvrOc0uUj85HbkHOk3CktGBpMe5B2rBy
f9XvJbVrbT7BDyxxj0TL4ZXBVhYqGEindFF07jqR2JM5HdeUWm3npf5AvvSTHV6M
zBqNFkQ2G+zt9q31odAvKhWun2zSTZBYgyIkJFKV+7jkI2VZwCb2iZU6zxUgsXs/
ypAyJ4PJ//KC3TW7ADwCutETYZiOB+vi4QsKkT6nEtJCAiylY7TOqdcRdPLnD1B0
WU3LLJ/8kuEU2FXYuf06IJ2jdcvHaHLH02VNIpAUPoNCAjThrLDxygnZUhpfWqG8
BATen26Srx0RBCIxj77OvhlDvxJnvIUF82cDRUXtOHpQcfCUI6/TdKMgDx6WVPqB
Vgj7U4Hi/EC5yT32dZjVorLJFfmz8/QaMZQo53eSdw8/Wb5emSmMYhEsdmN21X5w
KB8cCjTJs2haoEm6fiQoI0P5Jh8SYKrGZjKzyAR+IZHA4H5gSBYvmkmU/hM+5faV
WMiuGy4rdqR2swnZaVI/9RnOpZFouIAPK3TnxAc2rpWmJmAFHLCddIwZg+P2/SrG
DpYYEvZeN7zmOkknxj8WiQ==
`protect END_PROTECTED
