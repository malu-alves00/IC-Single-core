`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Hmn8UqjCm1AhU0m4PBG1/UuIikfkUFdGR9MfFXWUbn3WG/sOpSzGbDr6yGEXUuXB
0N5NpogApN0/n+qYxIzq3zZdTN8dgr3nfxSM36QW7MSWMmT3sTDb2VIOSBUpv486
CkTAUMn5UxMXB7KG4yS0eBnogmRQmCO60d/XOoKeaQhiyVgn4I5aSLW4qV9PcnZh
QHWZtFJx0y/oXG81uzEeLupgPwP39JdC4eBXczXtHEjS9zhFFeYYdvf8MqZwCmYK
bhgr1QEAwSarHgnHPDV42qptBEgg1LRPc6n411BTc5ss3R4zbD55evzGBMSSPX0w
oy884Qw2uBgm05+5ORykagK+gFCRVOu0W5/KV5oYfqn6Grm6PbNSoUbzf5L4kpNl
Q+FQFBNqMeaVY6bche8uDRVYOPm78SIJhCepXW3py9R5MwIve84HxJcBpHrE3CZg
KVXxYtMSmYSbqRjZ7My4Vs/+WQg+JviLym0EUpj8aFML51KVVOvTUuiqmhTX/4f3
iT+hpBt7+4ZbPgOimvMDqy6mW/hVK5rQ7kMGZvTjIjGkTA+ZCMYKiW2mak3bNFlJ
dEyCJ1587woW4+n/5aPTZnkSiwzbuf/apaZLviB6hYc3ZuQoE3YJnDsVkoFBD+rS
VBbuPj/wnwjjI1//Le4lNQlPBu3U+M5WqITzPLmG54CkeDd1hZG64fOutrxRwKYM
eRUicFE9ELovfIpsvdlxKcmoAbSix3yuRzSJMrWnA3Zu5/TlnBArrVRkzT3pXbu0
XyHyeOb08G35tMVfFhwzKlpSdqaq92fRZPsakP0oZP0LiCZjx4Fz4e9TtzVv5nBP
hG3skEmQuSj0cflEpcASUfAa56NnF/GM6nP1pyDC/eaDqvvsqBfiN7IzGRLJ6NZK
51IvHvXHrwGl/n+U2A7ZPVgKPmq50akSTcbOzMlKLhtbBiKdDocNRlpN3gJ4fHeS
tLCOXNcI2wpWCoCdwWWLIZ42vdLqNLzFZL8IQul6KbsGu3OlectfjzOBXd9wbpLs
26wDwgIn0OFf41tVCnEtdenZqe+GpxmgT3tSj8QjkfPatTCGF+MWONecB0WVV64+
9/UUgugmbSk88Hbvmwl+cNMlp9LUeM9a8JHoJVX47If7MabjMmj0B110VOwJy0v5
Iy0zhdm0ZC4AKsQf0I6Xfp29aGuk4OmWnFyIKQzrvlAcgN905+zFWWKETWc9Q9Sl
M/hmg6vlMXzQAIXX1TO4NYZ72WbzloApRK7swyVNejcQujbJoV0WGBC46ldP8KIa
mpW3EaBQRbBURi7+dfyMLhy3oI5djaGI0jrx4MQitSTQO7hKCxmNB42Nx51g01oN
rNaH7v4+pz251BuJYBF2nF5w5W7gUrjRxsBwPlRqeIY1NYmUA+iqrFi4fJo35hmS
8BE2oBwCsRfUdcCWzkSvOBpNBtS1w+GWM05wT3oIxjzIDdXZ9e63ViWRIpVbY4fT
TkiD17uPObnfBsjalZ+ltX/JHFTvMxBfAag8DpCoyAdw4ImLNw2V8Est+OZiCRX7
dwosIcTGb3DtEj8w0qmMnSQt2zc+qgNBviFXTLUndJc772PTBaJuot5fHsb2M+XF
Q6yC5Epg7vMss7f80UKQ3s+WGdgvYOWa5w9EY7jLXk3PiQPxetujcoaTiO7vQP2D
RYm34Ly7Rv5gyCsgym8IT9/OY7nwjr/0+bAFjxyUIWWOGUnQ5xAVKBzTRP0be4vI
e52bVL6QsKqRNi3ZLe/PBc2gP8XSu34x64jKyaQlfxiRPHQ4UYo6BzCAEANKHMEq
oL+NTbnlUR0eERURJ7VH2v4b26V5n8iKubFUxJlAiRvMDp4aI+KFyoEH16B1SLDg
BkcE31NPstXvqYm1EWrm+YYi67YRrHvJmMr0/KJyw4GK/4yHTA8sir263Ste6lsZ
liPlzy/3cWzC+guZRexVNJOeRzwotPmbikEerrOFMonQbfFEVH9Ii9ydFEIxfzTR
zSrMrDXjqTGO8HJeplGzJ/uQ9MaqxfDNS3F2Bv87jcnVOxBQ8ljoZacUOwo5uyV8
Q6aLugGKNbTwKMfAq+4AjE+9QbPN1TUwZ0xqDcMLWGeSrKj+ilLpWBeMM8S+Q7a8
yQZUaMvmCtZDmV6nTJi6CWoelz8IXOYO1/IuEhM6BgZDVX/XZJhM3ohvphOCsINy
7qr3EIztNrRoUOpB0enNdJzaLCX4/xRjvmtRm8CvADV6NM4Ykg7aksTSAGDy/Itd
v28g9C68Tc5/vAEASfNOP/BQwLZQwelnp+ndsJMYU6s0gW1G/VVtvI8YXrbfovRQ
by7GJ2Utpkjt7rqvxXTqO4JbQFQOhMuXM4lQrSWYJPs95geh3/HZicvdwC+J2xqM
oZ9pWWigFBWPAFJIo5fn+HhPwG2USbjwfs9dsnZ9ilGxv0xB8Iy9LGxKb76y6GnS
AgwPHH6+zw+Qx6YDuyuDccqj9O3hWkKsFySglo8PFCjv5cuTkN4nlL9hFHE6D53l
u6IPd5UWh9WRGCdAlcUlrI0qRY0u6+GQkh/wVp14zf7vijeyyyv3mCqKpowf7wkt
zkd+oqFwec6Mb42WGqSRpUso9CKqFhU9vVQmThCGr3hs5Go2nXGy/AZChXPnuPKR
qTEfFdH24D/9WXBwfTlHb7JP598iTIxV5bGytt3+D/OaEna6zzi+q1BKvdgQsXCm
x4lX5x/RDwcXfubmocOsEsPOHYQMXYyYArpubxMv0091HteAgxLasRmD2MTsFhji
/P3lHTRMyrzLtV9ltRp2ucDW7CeYUkiLFX1CHfFlKe1loOgJcEheQQP62yusSlJU
HyofYRGIbicnajR1JcV1X+8GYNRzWmADB9vpQNZQBj32kdQPrld/UnvBbF0zZJmj
1o+BRwNDu+UmFnnNvcKnvHSUWs2nQmKabWvnzK2eNp/6kuEzz37vJSrXhTG3S2j8
S0TbdJKnjc2aRJF8Wm/9XJBY6SOEnlrdqejizjxzLcbpA4cZ94xX8pUlr1owfblL
yC4jAohq/2x2sZslObmpM789k+LALYnclAJ4pcuyc5Jsbo83Mv1CimYPzUE4PEU/
YG2LVj1gOhfgKvHZ4DxxbKNM9yJx0vjc3Mv3hgsu+lX08PE6JIN1QaJjzt8JuSPj
u9M27HRzWBKMIlT0pLGdZRSXIb7cyQ5otTCpDN9DkeBQFn8cjfuAvfjZ9CPMH0Ek
s/qSg7ohTJ1ammjwGymsOJM9z5vOfRyQH8yuhaeC/PHy8P62K4LWeSMKfxYzxNWs
rj8IfdL1KN7GIcykJbV2p9bvf+4eTdzAjUUkwvamyuMsL57NQtbgYUNu76nAUGdg
CGtyry5dhiwpnGhMqTQu7rfYv2OG04MZ3bJBGsa3MOs9p6bFY097Az2KnNMdMZN/
YUjmDfUlQ76GyZTHRf8xnTUy/2VZnaorlpouU6lZaEjdQSzzlQxxL4cJwAOjpwpJ
uuxaO6vJQeqEZDTp9UxC+cI+mo9dQprHG6AudT4gUgN1ANkYs1DtoKdgbjhMZwFm
Tj3scaVswRY4aMlNqNaBUbYOnOG9/HJ5aNojV5AuUj85OghFrJCDiiSTNqdgoe1+
b13agOb3pasFZyblUK406kFoz861TC1dcDL9B7oixCsSzlh3NPfKEQ0axk0Iu7yU
tfLPZiYqEDmBF6mPuhbfth2yP6rCL6SF4aTO83hd7HdNKPtxvm3E6KtLwh5I4GEx
6dCPeaDzoSB1ev6etT+26dU/IPXjPJ1fcyeJ4h0l8fVg3CAImkp4S9xYeme1+9Lb
HsBAwuX5IgwIdhzIbo8jn78Pqryi6oiIlPEySbj2BU8F767g6aUQ9MwYREBJyfDI
w03QmJeCkWRF35SBukvyyOIGNsvBs9ZxDVJK305YDszgs1RbIaDr8KAVre21gMRa
+pG9vT1jqXF2n8FuSX1FMF+M6E+31hWOg3By4MCByNXDe5Sz1UQVNLhmVA3Bkepr
rPfd69rKFrtQLUzVseFWbTO7D0vsnKj6AwT2kq2dRAjNFtezfKg4q8SptPZvyQHo
AfC2kRAcMtTgcJ/qIl93z9mT4v6lFh3fDojC92PH73vrWzZt+gnnrCuuEarS1Pkf
pD77qKiPYh2Br4gKF0pDjIQSgoS2GKg9oR3bUl/aOa2qRbM9xnH2gi3xsVsZz1BV
tAg8C4pdyoyvRpt7Ct2YYhjp/XqThRfdX6fWan2QrxwGOfECW4ttDH7hIKo7U+BS
elJKYtKlbtKqmNrtU8N5sSqQ4uVdk+jkigsMbfabt5IanzGf1Bzy9xErghA87PgR
DKlK2RG0HJZAaRsXlaCBKuiPKUiIbh8DlNthjSPYu5IiYL2KuoHwp7gvYIAtSCcR
7PXsL8LJhFDCLmoTW0r9umSYpH+b+aJTSziCvFS062cxLV/fdVg247vBvgbuvvP3
uNffB84Q2/p88dlIjWzQKRLmthWSWOD75XZ2gHpQb1r2cNxgo4wllX5J6T4u7M9J
BAKgTikkfNKHdb9FgpcaN7BxUM6G8Ormx2YpVrvb0liRAJHkkOVlUb4yIfzwP00P
9WY6BuCShCzK8SEQQi/2CgVUZZQuicZ7xkcyjVbkF998iQNVCLVB08J0l0j4/sWH
jOwV7Vgc2tzZOIf7CKlO0p+g8T1jxTeDKOoUuEpqNGlug98SV2s7KYGHwKtNifnv
01ErxY574sotQua6NiL65rHYVtZ/t2NKHZWNZP/VzzMNGD975CL0w//5LKcAeU6S
SradPxTlCp1uvvnzJfbtPPojHZr00Rqi8oMGo25dv27hYgG1ya4FoItaHpRbV+9v
mHp9LfRospRsPLzW/xUMrTT2hot/slFHNDWLUULQ7QTdCHUjYGMDQdKOG9fKoNQD
MDH4NyV/J2TKZEd+ahB5tZqXfyKqHSwnEdC1Hgnd/XZQbzHeZIH/OLLyzv4yM6Eb
Z/VIhn8cJeInc26f0gpzbKdohoIn2JxqWFw2JU/L4ah1TbTuLo3SETV92UTQYtlS
m/AdK69VMa668E4HCWl+YDMdtCZN3syeiJlrOSnFBc4Fw1Afpw2VLiQZpgiZ0m+0
TXXziHkl9O5OIF30ARCKZkp7X5KamhhULYmSeD4T97Ug4qjuyolwy2yacPWWwDXP
uoidydHOLgHtZzLT9IaSxYFu0vV9hbm8lHUtbOC1m8rdTXUN8KpgthvSdvjJB/EU
tr6cOm/ReYmJt5ZLP4K3acDOjDQx8BnKIdUR1FTRDIAVcsRHob7IQWzJxru2rKDF
MSLCqAeVBG/IkVqJWdpsHQ3GOAt6rYhbyocPp6evGSiKbmFuMYnU42I9zJl/YjWr
f1ntEC/Kv6Jmah78IAL5qMQ1or0SjCcOV6EuMBlhDq02u+p3rZFKCdRC/IDRk16H
5heo+sjvwQEGKtkTJTB87gZtRcwPffSTbrj0gMYWB3C/wU0nBtenN3Mv0AaufeLZ
NGIwb3uQPdqJLdZWrOru1bP+eojviUiqvNrtU8KDcmvMUtZci4ddY3lTfPQw2UZE
hWmxiGlpjo2/IsoBG7F392oO5xzjN0PdfpI7fHmJtteBomm9uqUPSSIE1JQ5ywhy
Q01n0XT/SeqUrRLIJQC1959CFG3IvU5c5+nMTFBCj4072jX/iQgXCBUIfpopTMEy
u/p7wG6BwNjCqLXkPAj64WxGAdxXEjITs81MoNnBUjdncRo0buS3/ofBlGcjvAG0
K9CUpHqUWMWgddtBk4vH/mcC1BCzmzSU4EQxvmaZpPq8mLhV9jnWyPEYXlE8QO2V
RUpypwCq9OOJfmOT4Ox4JpUZANrjcS09Q9GGFpuMf+Git81b/+sVAaOOt4CxweaF
BsE4FMZpasZ/TFl15Qo4zo25NeGe0cKE9586u3iJWuEsfwcVj7us/SOe+wra/j9X
cEBWe/8sOTVdILKCDZ5xRpekaRtYUxU4Tls4ow4rOiPmx01nQJZK6FTrXmxeBeY6
XTqYcDrTkxxAdjiqj63Rd7cwafYuemJY6p0YEm0dgY/7nSTY27BrlNMjEIf/jaoV
PR09Ab87AEL2pj58fZ7FIZ+1ljsTfTQuUsPoKZozUmL2NEwUGiTlPYZLafLAW+oO
4qJbhcy57ddlRuzpQrO3P4UUzjIVkO8nM2thQl+k9Hmyh/rOYPHX738CFR7xWhkT
+AI69kpZ9w7JWNUOh8AkdfLi2P22v5/2yJHq762iePCvhUTcTzhbD1doFsZ1/s+I
KjO6DL9egoQklpF7K96eoKLx5g5qCVTIC0ecq76+rUnYDYEDlEPQjFXiC+/LYSAr
GJJioYZ6JY9Wu2B+fucZp0ZaFZp2ySEtsdWXMqOAXnb6gLhFqPNJ5kBUBYykYTTj
8X4w69qZOdT6+wddlp01fBUOg3M9gr2xP7wb4P9icwPogyTH1Twzi7W13vnWhZ3b
X0TplXquj2FYAfg8CawZkdHmmx5c3AcAKXJ7zXuCh6vDTFrk+XTfAcCTJ2xxePU6
0Yrr98201qzWloTDAep9q3D1BIp3Mug0VPqOXYPzmGHR5HIf+c7trJHY1EfGjUdi
LvV4AF0wdJkmcFC5rwYxyvBD76xXzNBZY2O9dgJfBLzyEtd/iAxmszdxaTX8+MAE
piDEZsO7J69NF6R3iNhTomLzY2vjjJVGXSjC/z1cNXrt1dfgy3lRUflFiworccVA
KFA3TQ+x2UNR/0V93vuqVeUJyzdlhffN7HyKlESsYFRmxS+P/n+ZqIDa8OvCOFcD
ZIWBFhVGOXC3YbG9OPJMimMg+stoFvUJvGa36FZGLXzlvFLvysJjvNA+GQgfGDN7
BA6BJ/UJaBno/5Yx6JF3pD+PK8F1N6nZ25ZmM/VaJqEBSaPQwmLZF9Gc0V3FGdpH
S/oqp60TxPPZpFcuy4fAEsG68uJXhhmOKnQyojFlN62BHONcohQVE6wgdrXNYxrw
C1Z0psWrMXQfwdvj3T0z3eTubkjglocCAowfHytd6o+Q2N7tJ511bshBD3mMnsPi
aoBroP/n5z115NHE0GyavUQTxNhPbLJYOFztn25b9piA1UrD8OHX6oTBbWbJ9sk6
BAWtsEpGmLDQcY90g9ULTNdBcqEXCw+XjiRCJHXc9UdKRgnNYfxVg2cryuqQwljh
kWatVuw8j8FNkTzevCj25zrIO+sbuRa7gdTS1TxJCvoqFkp0+aTYJT08Ws46yQTh
5h0+CiLDFjfavN6Nav3+FYatU8lwc6hKgpATvCBL9vDqVUapv4b9A0syX4BLSIa7
pdzz1Yb2dNEOZ+lWDB7qSqB3dn3vi+dugxOisFbovwpc568DWWrqOxx3khl4no2W
OkUXAIqBZxcH/lLZTFln0xI5EIr6OAYB1YvRM78hXsT8VeRGDa9USGNP7pwqJl7K
/qnUxjigWranPweB1NxB/RVq/jLirLOY5uwCcjwdtOk+1xqLQSABzHRhXIB0w/41
JhEP9SHv3X8VkFquvdY0gVcN3C+NGMq4VAH6CysEPMRnFVf0q/70qImoPR5ie/5v
Q3L40EHE+mS1YiAwILDc538Qeq96/0aNq5vsOudAWIiqzhUB4Gl2RRgOksLV1TtR
kpDQyw6sOAptNidXaD9+o4ITmQlK2J6nuZEY3Zazx5MnOjHb1QCPiKsuBYuENTVD
J3MlJJL1yovrHgEwk1pb6+Wliuc6quYodSnZdXV58Mo+8d+RcszuI4SiQaWnYbc5
nbT97SB/2cP/5LWY2cWqkBopYGo1P5P1oxSj7/WvGhZNxfPu+tnJdqKsRdVI4fpu
c77HmsMPoblMiMqHDvPBYZcVHeb113mMmtextcA5R5a5CSyXCDOXXD8CkVjR1IgC
cNHy458auJyOqB+zEOERsNkEmU0B1te4PNSmIAgTH0ubDqPjNg7n8Cr9Pienhawn
vlP23vgrdmVDdV6gZVrSxq+X45WbwnQSz1zdWWuEC83tg+/Fh9T7LokA0JGeghZq
3lM4y5+faM776Iz3CTQn+xd7Ytk1dMf2XHWm64W871Kd5llIFw9UO4a7BN7hWw+1
uYL1DBfErFq0CbEI81x5lBIqg3F7JviVjUPJRyEgy659dGzp4Tip/xGAXvJMBWbZ
gPuLWncmGzyeR7BU61a+SdimnXrfFFnGMjFHL3/qCbPJvZdCXvvaGoZHIFAp3/J4
pYmN6h52c+4v74xejy2Tnm9vV6fV+Kts2Gfc+GAMxaj2uSWF4kF3//QUExpe1SiZ
aJ0nB335Zkec1D21Stq/kLppXT4Qk00WJ3Gkty1xwjsuHFRfohUgFhlR3DAzLIqm
mKTa7+VmBYexBvC3qB+L4q8cwemMv+fSKEgoFyAEuszqXJ6RNQuSfz9vZ7EIHD4A
5HgZz/yXxH0ygw5R5mP+qMtjUtDJ7OLpbvrAdE+jJUraxUNJt/710NdqOP6XjmgY
ltwMq9hCDo46pQLjZqOH+au7wbi5LRazgVcXe6yIGnRBfV5vJaiQRuwnl6fP1+dR
xNkp0xf4HEBLGM7ZY1H53xUBgzoDd03rkPANDXAjuZasDhfiy1V5FYnPi8EdUnSv
0oUT4oRir7D69bhpyfqyvc+TcWl+6s+4LwcCeslwPasCfiLYl9sb9Bld8PL+G2De
Vl1wc/GR2X8CypBiSM0zQA1N8CVB5dtM6usV1poh3gPBpqz49AZSSQaplZ1JKemi
oq9taOkYyPSr2bac26J4Z7/eatFv0pod6PaIKDPrRTUHv18luach0vhZbqj/H6Vs
3Ghl+eIyVQsRLGPvkCmOW1OTnE0iafHS9acO/QLDD33xOYweNZs3FsqyrQ9W2vXh
M6MklnYFqv2MkNr/E14JiGBas7JT+z9NXDG8UvFcqB+D0HmEiTcADgR4bush6wj1
0nQql+LyX8sIwYb+XYocfOnCHkmBt8x1CMact2cymBnsWKgslqt6TNMCsgd8YIlY
omG4kpD26HP3JY30iORgZBqOk4LbTqSIVVyM6aLXr4NFKhPB0DTuV8osCh3QUclV
j3geFm4geV1TH0F2DVF1Y7FyrrwY1jn3mKVXMWKVyQWSzXIV1XUQMFcF/Hq+Pj+X
rL3yqPpwzcuTJrMasC3n1YbibCb9iSHEIeWIOtGvlie4pTwT/C0+gVubxDezj6YY
XCQViHgEaOO95m49w/AdIQeapQi6DkIeFoMH6jYYYu/Hsv0fjc7+cXf9gnx79KV1
aO+TacUipGL/ruyGlpbX88d3+BtiFshSbV5xTgn9KkQNjwbkcEQ342B18FqyiKfj
8F4cxYy/fXU+XnyZNZworym6Nje0DD0SBHmgarLZP4JDrR5JeaFDFmDEHWxb4mwk
C3OsqqEsy+INGQSudXlrFNAxagT9HnIGkRUzcxLXCVqQahGMVd06qoAzKN9PHMKn
Kf/ilDa8yOQz/c9YNUdVYmptscpxcp46p6dP3c7P+dUkb/DFF5Ab2OlbufRuJi2Q
FJofVFVI/ffueFN9pFWHck+7Ka93o6cQC+hPBeBrbDHrL3q3CMqd27BbJXrBe0Jh
z/IY0SBP8spIsf1GWLKijfay5BwPGZWMWESX7XAnuLcu/7N6/IFn+UMKcBB4vK4+
v0GUH9w7/sipnaKypkvfLwvFfDHONGp+oUXflJ0bzID1yxe8ZYCM4w4ytYXwEkOK
D9EW+SmeSPNI4aQKC5OsIY8fMjqyrA0iImdGxprS2Oia7vz5Jbsw1khZDEpmQOLU
Yyz5t/9tCN8A87vmN17ryH+IX6l5xt7mFwF2xyxhJqB//zJ4H/XLzMlDURZVdWOe
2fYb7I8IgrjoJHsyPKrIqpczedSIMw/OuQywDSW0+Oq3DfX87VCs6wrSLvkvEsvJ
TiGAHoc7qzCKbZ5C2US8T/qtPwi+CuVWqX3aCBlSoTtTTsAu911xuUJLvM9ZZd70
m8dL2P1mV1D0y6owFmSHGPCXgtGZr6NONkjxXxHe6TmZcm0e2kMHN7Q3vEok+lH4
4OvqrQ1VKi1Q4ZEwCUSUK7ygpLBR5C6XfVLFHJnKXlDgsuspvIL275eoRUHrdvPQ
vFS9lXlzOmGbdNQtd95QdfAiUyT5giFESszcjHlkjkpDjwHOkmwWbvIH1fyBWBPY
GGgMP3isiVOFuYm7ppEsfcdggsC6vz2gAiKiCUsmsB/jZHTlYZtaQarzOvUGWLKm
34LPBoyImKIOgNnjxQyY54bJGC0Z2bYat9Qk4BKqaA5vBuXV2AiytoQ6cUBgpjyd
JJfsbhDWfTobKJae+DYc4cXy6gSY95y3Ir0ng8/4xiMSKZ7YPZFPOMgVxzvXo/vJ
Fujgu/Ru1duCtlETEGY92wEK6OTJOdNC5rhtk1l1CeZOvbAe8sib4yhkLmbTFDK8
MG0h9lgpvHHKkTR4KX+TO076S6nohHdkkUBBf/+vTpL5FDQIqGhzWfvRuRF0E095
sPSrmenYXr9tl5j2K6SJ/3zFmZsiIBEChQVNHN07Be9lJUwLjq6OAGa0IZptJlmz
yiwfmaZcY1o5xlDcncLIvgYqqreGvRu6aMNMPBSYqogoPUfpUHfyWn/eDm8zJQlS
q8QINPHZ+7TU2rK/FsGKlf5J29aTw95nwJyoMamktxEaiph8oppsfkJAiMk2IpD5
Md30tWj2oKoecIhgJzVHHhgsPRwGtjSnYhax51iBH3PzGq0yD/RO6ngbbLZt8k3x
ghgqKIR9DDFdCzZ1QVED+iOg+q3y+9VO8aWP7eO2Myh8y5TdtiXXzKlWnWktAtD4
w4gjz6f7Nt5brnduJdD0/T1vpTzsi3qF2GvSyJZELa13dBNiqksMYnendFJsLhMe
+LsbrRoDLb/X6NSLYxYTBwSjBF54+E3yQCKX2DMrlK7DMbv+jcK7NrA4zJk/cKrr
mYpLwnTFx0EWz7y2bwSLFxz+H9rprnUe7opUvy8+SRMfSzxbP0K/cj17G0GeG81I
P+ER6cDn+bTGRDDj3BLx1SPEkgHNIRY+UpD/ExSW/M+0QuA5/L6ut50uZDXYcr/D
+AJbkPg1SNMjKpjIiJLF6Bis6oQzjQeKLBrLrin6nHwN0r2HKmzR6oczelbHfWTW
k5de79t+FdaeCrQHvjQRKjd3BthTrQrj1keA7PLvAJtfrA5LxgV9yKQ5u5VNCtRb
yA/ORlF/5s3s9ilWek/d9U/7e+9lLP9rKH2bagVDBq6Yq6NteOAvPDaBgOEbUa6I
bUojw8EMwT2cvVY1Ez0DO/T17+4rRup5wGGBFBZwsQfpdZ5HyjvVkBU26CEeUa58
qPAjWX13MHrkXPQLuD9nYzNIdAA+G/4PYDDhgLj1TWZa//Pol2Hz1i/gzwfI1K+Y
EU2pmcFHpIqfyIulq7X/SZ9+VQKjdlYNiiESqrK9i+x0dxnunHlk4q6LSZZGKAmh
QLRzN1YutdkFfiw+7XhsnIzOPn6KHJ7IxIbWFQvKDSerPqbkpyyNf7bxcYjFTk5P
L5s5/9aDRjQRDKIuBvf4kVOt+mqM/Oq7V1pwaYAZ+lStrfKjW7Sks9QFWL/IjeSH
W4wlmioo3k/vZxOOH6AkzK7YuMDldc8dp81Lp5EGL3kgPmCJ4x1Rj6mQdokblAiT
9vjydIaPkZPxs0XDLeVJpibgykyUmzbUqmwb2sZ9FGF1wiDUoyi6DMCttx10BJlh
m+BW2tXa/ivnoUcVs6lRfuNyy53aj5nNwhQv7epvX1nNp/3uLblSKtNfkz56vrn1
jEZbZ1l81Uj4EiqiwkiqH3D4Yb2wXdnK6nt5+AZS5q5bEVzSSGzPTWyytDvR6DPO
4YPx/v8z6qYGYiOr3+IBhBa+WzctQZM3fVO4+oQqxnTUuSxstfffUQteCM+bGK6b
sO5276o2c1PmFRq4UvaGenkkyNkK3JL+OTa3B7GCP3Wrmhp6XuoGHfBku3MJTgOU
sBXXuMtXMs4xgRCk7OhBtDE3fDIU5wVFIYyeCvYaWJNV49JKbELA945z5kOss+Bj
GnBc1Lirge546B2eXaKQ6wYhonJDlD1s54rCMHSMNNpDtNmik+0d6MC7LUGa4yCv
r4LDul/h1lsVdY9CzRqjXLkvZO9MvYvx1P6mEzdCTYtcO9dI91bw2NLggT3VoUu8
kWAOE8btOwFEksZGJRwfnFY/uv67QhVQnxeMr4F/r8GudCfZK+q1cFciwTLINMu8
HSaug3kYnJoqOH12BXbZ3h5uEz8fhT9GozktlEsAfxy/w6RgbrkgagSnl5leQD5L
of+cIDaDFtlvFAWva8dgl2ugDQki/CKdPyNi31geQLQDmD0PrH181JStAB2pDpyv
Az85BZojl8XQL/Dnyqq6XEIHhFPnkFH0olxW9jbs0y4hkdrqpNNXnOOvODF2tKHJ
8GhPEQopLj+PF0peYpQEBXOocQS5Dvrynan1Wwv2TIegDMyTnyU8Svt/KCLF1QFf
aEtkduzDk6SN1cpZg3lD8zFC2Wf/1al+0VUVyaKwzthIIcj8DzjvbABpjjBreGxz
j5Aww9mLNLDwG8yADnjxBYcntjyuCF9YOio+R5vIO3tiAcX88bjefKPq6/8fWYvS
NYeogt9uwORu1cZawz3NJNvS15BVcyt4EwE1v2d0OW3w6aGmXzmS+itYOP4GEF9B
AgqW5nu4iUgVvN8mclzJYK77FKWDmwHRbgeYH7Avxe2VLPdmR5NV0hfeDVOTInrr
YzrjdwJTeoPO+D5mjDwKaROAj/MUPX442r+WaRiiEEaRY3RJ3oxwkqnlNla2m/To
Gp9UTpHB9f774QvFRfJblShthH7JUA5apI3G5F36UZizyvbCidLJDPib1MJFpAuV
OOi2CSlmV4ehGwf1o5+pspsMbqgkYVy/u4vqOrX3itb82D69zQPi04HO+AW9/e1q
FawqskBeH+tSHr6PjTRAr7cVz2KJZM34DEJ8oBoyiA+u+/+wuh8XHZwdN9yNs3vB
znN5GvhLxNmDdhskc+7wzwWuPi4EqkxV/HupWuwD1nPX39CnHcz7hfuBG1GRW4EF
FaFJUXJAe4VQH1AXQ5PyKqewupQezMnzlk/CGrfrM9qbbvBeZdP/FE1C9advCu9v
9sAx212Db7B+fLNF/gQVm7zzfqmBSoFcZkhzaSGCxcVbyuV/5G/VLHDhtsxESBmd
mS/YySrYlgEIwANAaAjUjQidsuRxQ4yos8tjs1Hq8/8RQmxdTtOUPKO5W65aB7Wk
JduCCsAVG//O0VkLpGDHXbR8dViAOBxSg0FHpvpDYgDi7vhHX2EsOBqt8qtx27Jb
4RITXTraKtyiFJIivN+61ZrFHzpcAx43s0WjM1zcX8PUtDRmeeiw/n9fLM6YDp/u
rzAwXdo0FXEbNXw0o61RpXk7/divUWH/nbBqLFpgdGARiZEFtgy5Dlv6EzObokOS
mjChpIBtmjmloWSf1cgGZ8+2cdnTtjuQRGwBBRq5XbIjunuSw1a4reb/5mybYdso
UmGwH6lnbXdmKKNzcY2uqCzkxMtyv5GOkDHb7Bvgoie4oj+Kd/nTnpoxzPxfLzzw
4OkoQVp5/oXdXyMtxsZBz7rOQBXSDMHI5pW2VLBEOtGM9zKfZ90KRxZ6ZbairJKi
qbwJKCtH6vhQqu/LKP33eK4C8CWOH+CF6Vp8Lk39bsLokKZPp6PTediVIYb8MUVD
BXfjXcih4cq/XuX7cZPecbM4j/iksS6G+ZrNoXpyUBDlB7tiXk68P/+xdlw/kEIY
V760a2edtGNEAptZ3VMpw2nz5cpKV3aw9HL9TU1+NQ8j4VcKNmUDEVixrYrCDpLC
2ay25bEdXX0ufvw4Kvh7eEt+hKOlkFPnWYkZ9grWQ4rVtPt7pQ8fz5qbjICTYZew
5wkZuUbgToS3tloB+kMkv2FABc0/BBAbo2sabmUC1pL+PEMO5XYNfEvXOjNIPlIB
FACua5iqxEoVYE+Rmu3WjDwLCrumdMjdFGA/ZiQ5HK+++LK4GmvqP/bXmm2Nqs1M
Q7pLbnhA0TUW9lzUyta+eF0gkR9u+ZloVtdMzEZPB5k48qQwMgsjdeYIKhknLWXu
feg0WSAsAzvNEffcDtRmcPgZkgxCw0Fcx1rMMhlFr+rO2QpUIwabDyVLBKacDX3v
c6m1oEsF56yeJyjCmC44LHSyJTqKnEH9tBIPs+wbUeNvsuTDsIMXRB90eB594hYH
OsKjyfdtKi6uWjII7cfDjVUWJEI9arNnpkBAKfj1HDBRA4zO2/D+15Dj5ym4nd3J
gicsNKv8wjDP12RAfwBRVh9bo1L1aCnIsQW9zIR0Rv8Od6zK+LwdsuqIhYnyBC6a
7EfBdvlw/77VOwxCxje+YFAgrf0YEx8NDjtuas4vVbmTRO86FyxojYg0H7aREiEl
C4/DxCkkdinWSvoFgA99IY2pIyrLmlxYnx8OQOrzQAmf0KiWNdNXkO4k0k5Qt+xR
SJGj5fekRx6mLY0SvPkPv4a4bsb71gO8UGoQ6rAcbZSeWkF9omATM4IbmREkadGC
E4pefwdgjDYQasePGP/kratClQthoWethSomQFDFLr/hsn1VqIPSTRmGEaJJKJbI
OVAQ/ZYeVQC6qWCQPz5lmAaKDBseF+Wzc6IxUH0w4tGIBEXSckVYQDN+M/2at1DU
xRYB/m+YZiDY8ce/MzGNQo1OnuRIJtyT/5os0uaakDfQz2+7QuMklGdXqf5R9Vuf
U1Wd3uDD8cqncV5JA33qB4k8zdA1nYmaWAUSV4X8P/hsjNm8Bxjs41Xq5r9Io9oh
wl8tC3ssdl/LeDY5RU+Jh6lYewMr/+GgV8G+Om0RPI17kVPYCeTntKX3Ejzf/Qy/
3mcqdPNK8UA7pzsEkzojLlZQ6/GEQ35+CjNKas6tB+q8GzKdwZrGeZkJJjWmbjkA
Mwx6vDq8YOCGoQNBoOuivVCcOP1Db6znKSl2306G5K6tCx0YQnvNzZwGCty73+XR
NCKyqs0MnVVLAL2YcDNx49QIzy5AIBfOR3CTTCA1VCloKy7kms4qXM/6hZ6c85GW
0gwPTwI0X6ShOQ2Sv3ZODqKLfp26go56XYlwzSfTcvlisM2LbOc61Xc+WgiNR0fB
Dlc1p7FFpmHxHp3mGlBI50s6pIuAdURh79PFv4Jw/h9vDefjqYiZUkBoN/84L3M0
QEOseR2jr2vkNmSW02WJUkLKkeuKnLN8Y28Nq+QYIOlLDjqtBqkvAXKJhHRBXdM2
c1wSWFRylO7XitjFP3O1Pzxy/0KqNDQ82POAPPq49qz5MveWMYeCEwCgWSzGMQRz
q/MVxwDxrN37QHljdrImyijUu9XZJTGDYi0//bgOAa3SRCFfYji3XgSxZB+/jNev
2MSRhOeFOPocr4ne4Il1gVDDh42lj0ocWzuWOam7H2gmAJgQ8O3wauyqqeocQukN
a4MMxc00Z6+9DADWTwyPUhCaiYYnEg8yIz3SJRf4ITqNiO0+9CcrYHdtocG+A1Nq
hrdZCMm4t1scl9QaHW/3jEEd54Hy1g0aOjQF3u9FB2iB26firoSen+s7ksq1Zv8H
RjQyE4Bq7F9Jm12SgydEXC2cw8G0gYUk6mTjBDsYzbHNVAPzNs7vGPxUPxvGrAxG
azhaa5BNyF2OdQRgSSLlj+dEk0W/Kd6ez84pFp3Tgcv9YhwtvRy6mxYKoyn19Tft
SATmq/XRZl6q6NQw8vKB5lgPrU/brmIE62UunwSjpy0yBOsEzqxvaTXzEmWiQgJQ
HHfVpasgrnY4J68UsR5XIlgCXwnRKXyfjCOCda853YoiR7c6YtTN1OXS6sf8RFWd
wwzO5pcD11MrreFEdl4fiAywHmgVYMX8AaVn4boqE5QzqG70xfVTxs+nShdPETbj
e89+Ko+VAGadAasXI/M34dhuGmFeI50bbUtObNFtG6afleyWKaTF4AbaVdHKH6Dg
VRE8H9TSloRFOVRFv5eyJcQ+NYwmsiXODC5vluaDZDfL39eXDRY7OS3p5/ZK8Yhi
oTaRDB6lewDuxa2TxqAjFcAkTQtZ2rJrZtvQjQcPJ25sQs7vkvpOh7rCky2DY5oG
Ib1oAe0aq0nBXVK7LWTem0MDBPldGGyQon2ccbqVJnbNmc7j8gCPAr+o7aYIpQE8
2/87+mzZVLwUWMNb3A9yUViRhVge2CS3zegJZ3T8aJ5F3WIZSGaZbV3FpQzrXBO2
w5Hde+zD7us1IxiE4CA3pb8t6tSmIOB7uu7a31TSHVwg4H12dzl3YYRlmD9Bon6l
BbQRVNHlfoBaJ0yjEpSpRhH0gRDFx2ptf8wIYsybzUDCmt0n96PMogRrmLVoTt6n
Qhw2Apx/48Pj0zNm5r3yR+5KqoZQBLOg5PWotqgZIxioA0mVzjUW4yOy74razrL6
KFHW19tOC5imzn+vR60iJl3USXYoUjS1/DgzZY7REAz1dGS2ygjY83qCBwcEqnFN
xIqOW5Acn3/Zmv6IKKVoCDUDI0wDgrmkv/RBFJIemwm8zGuBx6CK5xcGh+I1tSC2
KNMUkRxsDZP409kgC31srEeKI5OYujPxDnM21i7z/ez+EBl2WUv+OUdHkuhOogDS
82lzemhWaMKBWLasQjf/n1sNTV1sykDTiD2O57nCAzSurnlGia6Ne4fFvlGBNymw
aY2NUUhYzt3kolInTytdrrB72lMe2rYPxrrq4JM5QM2ZyyVw+yiHaDPAtK9aGNF3
s/wvLaD40jlxC+XEatiqI8YDVlgn7SdCaXgKKAZ0uA2U7O0Crl43xLeMgnsv51Ew
aXYcGD48IUqFwOvZf7kQLlsgdgG2tLowqcxWmORNUe7jj93ge7iMjFBAuwWwqhYL
F1IuPaWw2Y0z5YcY+cv3vU7Jiqmn/pc22XOhnOegNbMOu9dVHzTUgqft+542b0Qv
WyKB2hkKWBd1m6dRF/o6x1K6JzF193p/ucE3JvA7EiCbpRCKNGTejCr+HEjgAlWw
v50jhsBTTmhydPqnacjf69Xs1gYVa3vNSGMJxayJJoGsjwg2P/P4j4sfDRrW89eB
moFXRD0SQ3e4frjDufnsUKJAGT9xX6nQLiAFnYHiSiby8i9xZ5iiZAo1bpB2MkzS
OZX4xoqh10FEWMyiAHuQUIN+OCG71/MU+JmpuVoIuOJ6R9T6abrULJabKZ8KubdC
V+rzSIlE6WVkictcY2nmnlHD+KlwoqGNErrbpL4JJDJRb0mxAF1BLgxkCKpfIUeH
9VtS5VNtR4+PFBog7HetjTTv5cPxQEwT4bWBVU4nf+0szXehY73GPSyw0dAcSU+R
5u7FaiLwDz3fmK1G6Duar3s0phH90tlL8qkUOE41jKEKh0qIkynNtyNHzoAI7GXU
1p0Ul1lVebSBuXnkO3M12rAvtTWnsikvM2J20xa6pDByx/lhNqCL9K03lHV8awYp
1lHiYmLb44x2D1ax5WWe1qdai9+PHQWvTMjk3FmAl3nJn5L1bQoLItYYdd2BqK+g
7OhHYQ16a9LbUxo6xlf3DKY11zzMzBrAbo7FjkVTiuPJWVwlTOSYUOqsroU86W2q
rxuwCE/1/xB25pk8VrGDCyfvxlSQ3g8pUAHiWOIZePzfOrZDSSIYuKqNnY8qHtEi
HmAiifoSVqRePCBVyb5NN9IMJsNDIgP7/brQCjeLerpNwQKovc8xuSv2tHy+1I0S
lisYcnJ1G5HSCYj2ecDu9/z/ZLfy7lwPrQuzVEMWyovgofYpS++f6NjkXAIMqaxq
3ZMyt9eIRXsBh3sKc/Ri4Q52TGOdbfrqd33srYZdRNxrzIk/BQbuwvVtxvIENJBg
tisk/4xkhR1RT9LzAw7SzE8+nf7fkwY4Urn8N4yxmm5lqzzAtz3SAZ/q0f+yw8eh
g1H6KVSuyBo3CD4KD4lGDVhKN+oksrC9YaMjaTrHFJu4674fUFLv7Xy1Ljo8oBTZ
6agTNDx46C6D4Xrkk3F74fM5lxMpnlxbxHRypkXiBnPGcyJcRl+TB1cbYeyE5mHL
p4BvOMczRml91jN4aHqSzn7yzS2/XIPs9bWNTUJ1AhK5r2JTprr5LmIhT3Yh0qr+
jJa2Y9N7WwTHEtRlinyRNzZv9JXO7BIKZUjS2k5AE1dcIH5+TEaEAUe3gVKvqRs+
WfVJ0xs4VymM+ourS0CiKTUyQLrsOBQ6tTdWV7cqDazC8n/lLUt0KYj72zd4YrSM
4mgzwz+n3mPxFMV+U07pcGx4fg2PkUG0qYFao3YwMJxOQdmOhS8SfKZoNwjX0IPI
cH1RXhWYr6wnvaHLXnMVt6zfQ5JfPTVV6kpHnA2lz5zQwQzx2DFV5w4AmYKom6VL
bJBxroZ+Ix0jemeNo/3lsaK1uHPaFwy4P7NRNXC52SW7tje050AFVcKlyy3tY9ah
nmYhLKxyO/HI9PlaXs1X6+/cPN5aSeosWICdcVXDPsab/LbJ0lK+4cZrj4JoWomh
mxHkrEyUtZh4K3YGSLjzQAuOBXfJU5srnZAyJveFowwwF1HTAROY83Xej6/ThWbO
Z5/TxA63l83VPJoVeVkui6v+isin8sxArMPE/aLYotq8R7TBYke0PkTLLWQjZ09B
VQqyCPK75FE7WmhP0EpQPuX0j2wPo83L/OalzMyHKuvHVi3VIOHyTJR8enN+IGjQ
METeDXrhtE6cLliU5i7b86hj/1Bb3H5I9kVbcv73W8Vd+kDSUZ/DW+C4VfEbzTVh
1jRVI37FG7d/qcWxE6n69JN4pU7wT7l80QsOjyMzYPtiZZrNVtJ3yoSx0D97UzEo
z3DTXWiq9HQFXRnno2PCFHQ1y4LPcmrPg9Rv5PrjvkDA+TMdbN+8qhX0YZA2qrKP
xr5rYPNSQH6uD7x8hV3GyEcFJbK6BXuN139uXy6QzGGThDBRovZYWO8/b3aXxwbO
WSEOMwMzbIVn+Z3r/IgjX3LXmjFpyGW2lGG284ca3I0/crekNTcryvVb6uBhhRYY
+C1/ySiW6zlsCVKlALAenPPcF6ek/phZCoWde9i5QEWB7dd4k03LMjUV+pAGqStw
nJifnz0yBQX8eFdl/+lGreu52OODDhEze3m6z6aqrahP3pp3sL692IGWo1M4MUs+
as/FfvsNJ53zxvOTIYiwT98emjnFAOipxxeDXF/8fkd5yuOu/aROrKIRU6+tZnLK
+UtQ4XjpZbV4oj73fKmztxqNc3NioXiRL5PcclQZG8xTJjF2Ld6RwG6zudQedI+P
9njjuSGtAPyq47pkbCUcY9TId45rNSf/6vXqCN1GSbAStsyfifw7m0EsWup3iJih
oKqSVQK6ZKank0ZPa2d0yMJ74V8YJOk+5zKbSwtlHExCK9e9DzfdyLnT8I2YMC9R
B9RXkUGdBtjsIQv9M8zzfVyyt1JX3QqAlsNT9AzdBBRtwizfBcaFRnbNt8LblB/P
HLuf16rB+J8+PE9B8ryJDyjQLE/KSyGLrA6gAVX1Qt6Ln1tuo0sYvFMQvGn6OLuC
VF6psnfUKQK4UZo4ZYM9YOOzPiu+O9AgQEjj9ILu9r+UcWzs6GX3blXK8+oZIzNt
4RmG9ZsjLw3cx0mw2jkcr0zJ9l9c2yaJgUYIlcIMaeh6PdPEqZZu671JQaZAqU5s
b/JF6o4eziXHQOx9X0s/29GDnpKsPoQVbGOPNoWJ7WCEXkVdLJcxLukIDiwdSipF
5rd/1gdYNrNOTJRPtDt6yKxDwvUlEDWbYcHrMaUU9Fzvq6duf2xvVBuACUL9fegV
N5ndDhcFI0pYmNGWj81R/9zGTnPotkDJ88v/LUW/19URWlo9mgBWo/iHg9Kv0TGT
b3DUO4/LaKjcnG9/hmyqttwYGC6HMfVhMdW51r0HBoPbYuNXn/9BSssRfoEaUHdH
OJrSMOGSGJ63IDv3++dhBcob6Fhr/2O1lKZAdePtkPxEXNUPEXbzj7ppl8OTgVrv
qVk0F4p63gu82Q+Md2nGYCzr+ndbfSiwg9IcJKml13l/qmNVJOg9EWtd+C8um/Lo
3Zg+Z53G8rNsfDG4jSl3eAIkPrLzKlaXNBqWQIkG3LqlbwZS5QWeb5FqMm3iiMsm
PH9TvxsmMem6QHz7iX7KzH3KsKvO8c0phkvDD3ZaOr0XV5CLQd8L/aI2M2TNK3Dx
DhST5j/iTNUTW79uH95BZZ2JPqlP3JRv3VGyz6oHk3GHfkPsqgNv8SGxsBpUSFjc
aGdUfKVllrJpu+TmoctaK0gDE89I/PVio05hxOp91beDDCYzBYBHD9+Vclx0NJcb
TO5SzljMb8tAEYsa8OBjo47o5vKW5t5Jy+OX852Elmg0PpfPr3nCs7ltyTqzz5lo
bWwqPDePuUZMn0/z4P/s49EZCPJz7jDOBsED/UIuOhamrXSwGK48bql3D6ytSmOp
Csk6mP98P81onLF8HEkdWDFk6UHx9Tbv5S7QNOlEQuw5mbPM4GgAa2r8ELfiC8l9
vdz62IrAW5kWKqlABCa3mTmWAYns6MvhIgsXirqrdxjjnoPb1UD8rwPKCzICoQw0
QbFtQJQvkWJrA2NBqvXHvzB31D0v19IEN6c78XDxI5wZ3JDDYSU2koI/9yt7rRLJ
zEOYTuB/7CyxYZQJfHokuwpjtLqnzglrQZ+TAKzwQ8IJXNhc3oXpXC9raT24iL7e
u8kHQYh/yC8EdH8q/9azQ1OAeHm5sjo4eiXLPd7SSxISe4fLQla8ul0E/bccsF6M
jkL0WrZrmvv4aqdwoYWraWLHQhYH9nxE0rPL8a7AtW5htQrEGCM08ELw/SgeJWb1
2M9W7YZkR1GczCaYZB2mkcKYMWRI0NHl/0Db/6Or9zinqOgD+eo3pGPgH0aC0coQ
CdvXV09z1vk+xTLfexc3N5LI6Tq3/uaSoNHlELT0AcP2mEMae86q9W2Pkmwqcn6U
Z3kKMPI/yAEK+ZIdliGkzZjDjd91cS24mRbKeN3aqa9pv60XiF5vARCYGcz3oloT
Y7lvqupBwVW4Q3BoUhaqH7Ven7BQMnYXjKifFErioTz9G203YjoX1jiR9CcvlqNG
fdh8lA/3OcseB/2++vT05wyEVVcS4NYq7pzMa+PHvhy1htE5vumqk3/gpSPJyI6K
tS1MJi6TXusFlGy1+KYkE7Ivrk5O1LfIA0JPwPk0dzaMYGeLIfthuPwaPrvA8xvR
Zf8Mm7KVIZD8aboIW04BIdp02RV2HsxXWkWaaB66Np8Dn7Hw/za//NaOqv/mtuLT
O1GWgGf5h7Gk9eHnWv3lfjooNNst3ukvT72SpGY+HyASPLoDXh8yXh9SP3wUHa5z
JAbEOgIDwb/e40TzvFc09F5P5uAOGKWzGJ/M+MFzVNI2VTX4RjGXAEYlAgOcvObg
WZlTffcGNDRa83Zx5ESICGWYAnG+Hdh0qWY3r0PPpD6qHaZ948YDljZKnX+699uc
mx/5okfeFkHfMcH+s1U3dluMETFUTdcpQTzlcSrzp9YQMJjBLSY8EP4gVLSiR/to
acam0T0I36jP4SvVClMa8oYCWOwLg5yryI6PVhYwv3IcWlGgxp9gCOulJW/Gc0Ns
p0T/uocSNzMFQdZr1sHWU9NzYECd0oJrVyBkvenZ+9CcJXlSvoq6iIYhwF73GESi
KcS4qLKrp+joAFWZyplsQrg+MwunL2c2VYyO6QfzvA6hKAfvJHbZHIuXjJRwSAdr
t6KbU/hchWfTS4d13i7WLVivgKbNVfB/sJUYA1tAC82ffq9DDCtIM5bPKC5tWq8o
PjJsksnXzEalfKqhI3FmeBdObenLddqgqZdF0XJ39AhV8YMt+WIHqpJpTnxk+dEl
GvnxtsEydAWeIMECaBUwxxvNruFr5m5pAlcBAZLalHg7B8GfLCbowpUmL+0QQAE+
5B04rVhiY3cIIZqXexUiF3D/boUeBnfUPxV+25Lattw9SvDLmNlbl1JOyp+r8Rbm
khE/z6jEQcEEjwvbSu41WGodtUr7PbOXh6HYc4PuQzkPUlT6AIdX7ZlABp2MXYbj
obqpIswTn8yDj4RIR1Pq/ZvArmRx/gD48o4ewLNm/3ITRdDkeK39GWGj+aq3vm2W
+MgzLdr61vBxT9f/YVIeaEav2LbDStO/rRgX89cKU0tKltp5GtYrjtZyjoZzb7l3
Ttoq2Iw6altjoKDcAZWN9lABwfTmXVCCs8ThsG7fsgp8gtHpt+EGV++iHRJH+uVb
TymKUydFIJnpwCM9QZEjSy8EYT1R+tuyzctayXfE4Mp9285xaJZx+uBf4yO4OIj2
30arlYBEu1KjP30TsMCFjzlbNW44XBgZye+rW9HiCF6/sVTYf3VWSU3rJL/8+Bfn
QrzdRUpopsPrM4HfvjXW2RyzbhcInV1mEHNP5CfROwGYle6iXI+vleMbwJHlMrrT
2Azy0nwG9cw5Q6RkZBfCZGLVEuoWFD7vxEKvb6Zm6eY9yNWAf12wyWp6L5i11Wat
YbyfL/RtERi0vyn5lqID6pNSfoaWBM72fFqJhJlnwwzZC0qcJ4iZuLcuoyiSNK1W
5p4WvC9AFnOlb6vCPXbBAaHXPxZF0NtTbHs87f2fu9N5leQGUBjYWQMWyZBc86I9
Vol7iE27SBb3ni27uI2SjSUDEzLF0+kEy9p44xXKzREX4Cx6UNQl3d3NSLLM9+UW
D8kBBjSMk/ZqCIN1KTLgpROoPQd8YWmNoSalMOJ0h3JIP/zwJNiJbUEG+YbHPvWe
x5wuOjU4qJkKNFpcZqv/egKbK8jYyo2DyokAcoO9pVGJPYpZcvTzZlZxO/zj0oSx
XhOLe5WBXo5nbsXARN319mejUHYcpvZbINmS30GEtaSjWJ5WFAd8B66H/3Qzd2IM
KYWh+jLxmDSwxltF4m/HF+dI8+GUR75QvQDfWi3QyRDD9FY1FllqqLkMA//hFntM
AIVgHJzEhum7rYDT3q3cCRzDDDbFPpj319r/9PREfnEXvugh/V1l1MGzLLfAuFRP
wXPwhrsV9zJBgV5MZGnwy0P54B3OyIHYh4sxugBPbyzoq2boIglLzSHcTCzZcYfi
CfoNX5X+p/IRM6hvPe+CsakmxP0svDdbp7MxECoMZoj/Y3dKTG9euHfLf43Yo9su
QK4S31JZdHqQz6/9DW4W8GiWmSBqm/5fuIeBgPjdBOjAgQhOt51Spj9svXS4JCBZ
SHWyHLzi6Isv1uN+GGCipKhLC3+SeyuRI9Wf3t3gakbLuDLUvNQTIl8wjB32vRzo
+FkcqFtn89Vm6CWr7B/h/RFZu44S4QGfgX7nxXYtN7ii4exfnO0IrYTEUBFBe0Ku
GvB6cQjsADHTxBjz95D5OV4B3I+iURH/f4rDTJjrqllx6JgnKCxWWy8pJNOY+ybT
/CTEnVWBI+wTOpIA7eZmJ8OVwgr5Ab9fYyTbUQWOgzAJt1UVWZI4IMs23910BAiZ
YvMxbnbEHXgdsLsXqM9sTEV6ih1NlnmZmpWL3iMo0OD07Acump5q3VQyhIt02fIp
c4H9inxfszNjl7t4+qnjYU3a2d6DnPgHQ3KI5e3oz3DKeNr6K4Ld35SrrMGPwXZr
gnAzIh9DC9xifXpNv4oNWH73O/Q/varIzuug8Jl461IsS/VxsfTyhkSIRGW2gbBh
IcLh5ytc1pD7Og2xiAnAmqVbGCZByoAXZuv9goVyoRdpRGKxsId5nnd8X3xrOiNl
bXEUis9OnOA6TcNzCoPRKzmJ5E7jj7R4heqVzR7rJRpBoZGB/KagP6WXx1RjZM2n
EPGUDgMxqYLl82PsKilcU/8NFaEecCoZkrcwyOBd5Qkc8KUiTMQOWjCHVbw2nP1n
Wam93C69dDuRGbKAl7hwaE2v8hJPz39Ek1dn3cx08Efdw0+PyUwNMimPk1mdpjrm
7iU1CJy/tTGbt1C0F7CBDFZt2jHYoEpfRg4kGVx2xK3sKXYYy+LpB/hRh3QV9BfI
MYSYeSFdsHEabEcfXgjeWkCTUrTsZ6xV5LU6P5TBLeMtMw7DWaNbQXshK6QQqMZ3
ZBW0oDCgVIhMjN+iOkjW/Nc/lQ/PSq56vE0S4Xd3TkxtTbpykOz/3Ik9L4BzYP7R
FLY4aQUGZxRxqVJv0UiLemYNvwKEFuOzgiVsZv7WcUWD+UliH2Cmhv/jhY5XMuM6
M2xjukFGtBYblMzhyEg2/TMBlx4fC7jqRYnA1vBRE2MWg2a8JoxnEonDmVWXfJAL
EF2ztZN1bJ2fhHvflK+ef7EXIq0fzEMSctzSA8uwxY4EiP0cSd1rRTX7UrJOU/Ig
YXRveH1Ct2JHArfDpyrPXrxzqfmE1vIX99Pu2OXNR/JIZZ1hgvCkAizPz43PackU
cDIaG8cGacLxUI4a4MsY3O9Oz5bYurlgrqD72t4y5RLLtedP2pmHLmxbvsLiQOAi
giWqL50O9rcGgi6eRSE5IYVhumpraFWcaYgp8cVxpi7bI3O7Suz9NDT8jo47SlFm
clvOgZUV7ZWtM8WISoRIK1wGbzNinV4j8ujqrxU7ZoJKEeaqlnCvK8ggw7oEDirs
nBxv12JjstuCeupPRXgbNxzCzIMJuxAZHhZiYlXnXf9CdhShqF+0dXtP8T4faJds
l/wSZOB66K0h5PTuWgpnxuo0pjKyuBxLGgX5hV5FMSka4fP84G6ZJlYG2OidT45S
+ENuaDpKjnSoPNzryBOyeh6LX8Z7kVFpwbyXlPBOdfXRKr/z5LiMoo21vO5UdU3J
oCVml7cp3MEEA0hxB23N87U2MNCt7JSz5kIz+bzwRY8g6MiaJT+eVdgdsueIb6IC
KR3SHxymp6pT8DQawCEJgGMgrjSDzaOtoine0QnjCPAcvK9GpQXZO0ZsA9Tgdh/w
0q7aVoFQcFmOx61DWxOzE2yRNMUlCWEfLpf8jpQXJYrXpY4HTeb3X4z/woggB33W
k6eGfslhl+GfXYjQWo0bAtCFvj4uUb3LsFs0Vkzkte4imKvZySalUVm1YBfjsmR2
OI6/VXOXsSdXQvjdJay/iHLyreTGHEKs9WD1o4N+ST984scR0vlowkxhU8bF1Mo8
f46VpXBqXrWoUnP47TATvHxQ3WxU8JsuJdM21ar+NCVIBbXZG+Den51vN2jqJ3mD
16bsmTnCwNFnb2YghC6HOWWXMhpPTfRibd8zXG43tIM/0GGuZTsrziJX/bHvesuZ
XR4ToJOfVnmWcU9PhHQG6C3dU2j8hld2JrLfmoa+RuiAqNmBe4WwFjK2OLxGKtd7
3mqnthXr55dWjPVrra+Y2Ydqt5FPwjDlWY8l49u7lQp9Ib4YdPm4JK2U4sVBtPCl
GylAYHdk7QXoVTwumlkjI87Xlr8lKr7aQb6OcCuB8aamMHukyJOwo9okLys3903A
3tXJYU6RXepcTtj9CvPdxzW6gg2arWuOIQsjwG7Jn0eg/GxgLQ4n630hFbsVE+89
Od98nZVjxrThMDPfUcCXl4dtJEOC1boQFRMuJW/HuSa9o3VgjegPRGNRrijGWDt0
UPMZLMU7qQ4x+M++RNRjLOR7XruzhBZlpVVQveEsHGcUDaicT3xDzBTAr4C+leFp
ZNW4B+zICAwvSOWBfMGq01Fvm2qpClTV5ojbEfFRw3BY2OzFUpf+c4X4QEcywmWB
fgKIEJIYndfBpjKG0WgwKiqlJz5bvyYaQHopU49nAoanzEyVCwA+XQTjluCtpE+V
9HK36Ix1+ziH/obePO6Ulua92lqoTAeLCebNj5XYgBro+hGuEi9Hpv17EfRvkD9q
XyuYCalNSmfY45bcBVk63xjQ9EDME5Cdm+UQ1GZzPxXMg82zdS0PyQ6QJ8lOfUf3
8pEdneI1Yu+PpD1o1vojMmVvbUpyS8OON86it2A3JHoLaD++CUazu0I+Ru4NAJIF
9FCHa/RDbvHQ408dKs2zQtg6JZ9+a3AVzcYQdjWvsMhhgaBweZtnf3tG1DtG0e7r
+wxh2C9fU++rNcKJHIZ2KOWH5kBMiOw5T7XNIqZH9XTId1dDyDobtAu28V9lHcRw
nj+lBWb7Hx1kLJN8k0SX/W2y6qgTzzOcOtHnR4Q1/4ojKOPur2CCt0T63wHjRi7D
5Rx54cIzgM3I2QF2fSaKJgU7jSeee+6M/rwBG+81Qbb08RO/0fj3LeCb2+H4fWLx
7uSlLPaA74MVSr0/NiVt9D0UIsKrbZfK2jOLw8d8RSJbvXjgqAw5pAqZXb6w0iPv
hcgUwwTDcJOdaSywm9si9v/mli9AhKbZRT3vcNPawfhMonKkPeBvTOrlGeU/lfdr
3+hkZpi4LAerESEy/OuqpEbhk56AfRVbVR+UcolSFMRkDiL9rab9Xpl/R4ppuqLp
xA3MhH/ZyddnD75c+Lq8EkxTa2r/sMJ2Bw8V+xiRtdC4nL5W7Pm4/BchAgJyK6yD
0WPwvEnciQRCo2/qwtABuDwa3snsTsBI+xtKolYW+a/A/tU3Srujw3xTUbnHzTmb
QCJJXhBx3a47Y5azJkSwWkTk4NQLDnwnn+I9bqepQf+zKu/kr631z2V5gaxefWLa
z6IaAAP4kOZ4DfLne6nXazfn4yT4LiwrHfnkvhCocEuogZUoH0AiMsDrvvsYkw08
+8WwH/uX8v9vMEfSMY2NgAaCmtD4uBRkUfN5DIdEuGrZHGGE22VvPv85zYfHU1YU
tCcdJ97GzgwVNyYF9KszcrrgdzskWXaNGNmDw0ieLa3veCzFRPbfw7dUKdOZGhlm
WW2HSZ5RNuZRN9iNXXC+FeoQS7ZOUOJmXKgmyc75/uY2eql9jKEcPgPDoP2hiL2b
AQ+h67YcXOYPeD2xOMjGfgi8rR1P5FFFnT84tJRFH0aiqYdko6sf5N679s4TZ6wz
H3E0hUXlY2iR2m0k/7WorSGyT/kXFopVMojJhNt3e5vOPKSeTAdgOaU15EFYGJ9x
dcjAt9mbqjgBx+Vg1axMrrSkMnZr3Ezt5NyzXzjlet3PNi7ZrIEgCXzWtdkkyt2+
+szDdkZnugi6cjWi4RtknM8sd2j6tXBr1UKvXduF+ogCqQVY8nx4EiM3D2+rHObI
ZuwvpUA+Z1AOs1Tzh4eCvdq/L4N009r6DF6qQftymsh46ZxP6F+O7G5T59Q2F3Yj
gwzfCOxW9yHoT+9F4PKiVSod3f+kIn2ZjUOviowT7+hTXjABcYo6qtUEciCrSY9t
c49megtH0ElmsT9kgT8NdTHJHnEstRRrbKlYUPu1q7XPY42jrNlH3+F/NckBscAm
dfo9bClPJcFYG4a3qx4fQFBCu6jKrYyFnBcqZ+aGK3co1ZmDX/oBovynTrnSvfOM
9CsqgKHcrcd/RFpJv/tie5w4GpfLyOMgqlXDqYvjm3yTtJxZnEyZdmAwp5lZE7Q1
PWaVERJvJYouIWyVYhw0tpsR/9iUgRuu8VmPsXIRkKt5S1rlRZNgTXSh/EtfFXdW
j0HeQexjoc1xo8rNE7vX1Kpp5WWcOEaUuN/lAZR77hqHRX2j9F8C5WJ+QXwLYiL8
rhS6bfJSm1aqnHWG3gM97JU4+k6Ecv6Cj/tdg2Ni5xjWa9kwJqIEr06vWH/eBtlJ
zximSZctCce8mCVcnBZTgkjqa4sm0rLwYOOr+TqUMdw/SdDqgaEODgH9R7zoZd7U
hFjBGsWP4mB6gf389ost6eJrPji9krZSQVg0yopvbFiZ1bNhskENG0JAL/KBQ0aN
iZiArNU4Na/FXEQKF8dcaLyyY8akXZ9WaVxxqIXzfSNPzgDO/sXJ8qdBljomfx6O
bki4ETBEnKTQj7q7NM8T9xoTKLZmnuwd4e/QulKnQ4J/wRbmQVVEduu00DeNvj2M
tM2Xs1PvzGzTJml4jxvJ6N+97SuT+z53xqM9bWvtiHP+9pFNkc6BIXjSllm6OFlH
DStuWWKPhyxN+O+PD5RbUFTyU+jp0Oj/BhHk4wsEvDesNyUjZlFPJP2u88Z5UlC/
dqlxtPi+VPDCEKqQTqjIF3z543OS7EduuBTodeRNvc6YKeeZ9Tqo1+gTpb2ficA3
OSgT+YBXH6RFoUj7xA28SzSZzzgIUrT1H/InS/jkwXYnan9cS+/NNNmvkCGug8X5
ujTWGjuQHeR9eb2u0V44Z1dZ82+fF3O0CF3azHivYPx89b/PYENHOSrCOmsTlQ12
nYT5rc55jUPVYwKz7ME5mxKVOvDmUoNM7DKo6UWoZOVRAS0alt/91zGrc/59NNfL
OsEpTW2xK+BM/nyeoUlGP2dFS/9qvHaX9im3TmvNNNgrcE6CQfY6xvT5aABmJaVD
2IivedqeydLcqYF2O946+6Aomina2YaiXYtJtr1XzrllbvENIz3AzMQp6Eu81mrV
uMBIeh7gcEmAYtokU1VxoXwKkhX1N2SiOfjCPmb37Hq76D1HxTNZ8IOMX49+1GzY
7z6f+NHlds4BMBj2ytjHVShQ44SblfJj/XsZKPW6VTiSQ7oMQVBERJLyEAECuOXz
4s0MUmaAHH8Z9CTo9hCjziG8caUgcQA87zuXKsZP+eUMFv+mpEfy2Oy0GXESyFWx
ltH7+sySRBITtUnkodwwfVmYTxtWHW5Z3puz9HKVn0Kn58rzkJnokQgYbo/ElKPN
erOUJmj0B1KPYz3qzbstilsBqwiFY6+aDCgxi4rGRen+/aHCP2tDvAz7t5tEfkQk
Ibyec/bm6Rbcv5QXy28xru2HRrADRIExaxGf+TsQ4tg8KbGd6hG4GZ3eRLF+qPyf
ON8rnks4F7NKldisGXAz4kf4RwjGU68NF6vN95ecpm9CALl0YXnK/kBrcfHAzf3+
2+691cZqoG3g/jCk3i32Rrpg3ixV0PlhYY6Muiu7t62lMVg/o9nTh4u5Mm2sxtKv
jfeErAw8RVGZUWflkdvRRmo/hjTEOxq3Y1yrBEnaSbx0Mi0St4CTJ+OwQJxe9Wg2
fL3B6N1rfaKpU2tg0vZZBuudp5QHkuPn9QkD2obt+QgsYLh7UzmHGnG66eVk+sQW
5AqRKEe8xz7d5do8R8M/+JBrFwD+Tz9L6FXLGs1mhvmUrxENal6qVsAM0mWm3RlL
GypvCrpZugUxRTmgp7JNVVrWufKhEYbIe2TTsOrT2z2WhSE0ilkH0wV6Q+hw87hJ
rMd/5Sx2sVfFX17G5UtRIZ+++RgE8+F14x2DqN9+Xx6+pEHXludDWagHnJSdK5dx
LeN4UHV6clvl6+zBD+3+DzkEJ52wAGRdT/rcy2x0zWZPtZJOrdu5TSX4K3FBTqfg
t3+pw5fGTicaX3vLB0Dvdy2QLP46izOk0v1sA4WFpx+YYzKrh6Z1aoC3/8yt/lUb
tMhHhE9cyFAfoAEiVqOJAQmAKEiDUr/TyKo74zjHCsZSzfutC+pOL34q97aCdzyf
uePXUdbUNUU0a7UZ6IxD54Hd1KZyZD9A1jyIGB1w2Q2C0chstiLBnK677Og6+V0x
MlIiiCTALF1S2BnZ4cc+14p+nEhDeWS8hgnpbDZW42ytJ/uT1vezdvwB33E3swcV
1V/6Fbji9j0zGnWbrCFZ3AWFmIPrEoIafnjDMfxczbPuVso0q7Kv/9N+Qx/Mf98u
fDNNaW1NPL1g0e/W2i9yTgMzcJG+C+IhxgEi0TNX/d/t9E/k/PbGeObF9aAUnZoS
L+f918slh8ui1JNTd//88np52MoFgxFoyBfcq98OROvs8/F03+CMG5CtWM/fhgiU
KVEeBwnbl3hLM67tjPzi75sfTu5zashnOs8WZsJTK2du3jAGIMxPpqZPr0yGrwqF
xW5b13jZXCrYDrpqo399Nev8KYWF9U99zdBGI3Z/JrhqcuSoh0dbjOSo8jfq4tL0
0yZOLqLwUvBfg6t6p4Ztu5k244e4RTZrzCU4HZxc45GcAeu1vTJXFtAwa6u+NY5p
wH6uGMjRsAzYeNIMUwiS+bz/SIu2eRYhmIrog/+nTRzvj3J69KufX4cGq4x6kFZN
ymp7WzWlDkVvIgHxSGd1oSRBDoIj2NPIvfMEAnNTAlNEkyEgE/SRxR3R/HTci+C3
dikvHtiL0B54/Scp9Ju5y+OxKSCGXo26ppTBx/B/C7g9aGn6fqwYAE8qrWtXMtPD
SRESeKj/dMs9g3cFFFcyiT9FluuQyXb9WrUZbEDFaP3OmMHv7X1ypRseUwhEubf3
TQxel2lV4bVk9AuqN7G28O/i4yba9u/WL6EkoI1o0J5+ZcH8d8E1oiTWZRCY8n3y
1JKJZpcs1wHBX9PkEFxDgRfXlkXPxDsh6q/9ldfgS/6EVI5+iS5Tfy57BPYAX8ZP
fOUxRJaUsbmiSqyd+sV6H6QIWWu0MHOWdFAqgNuwA4zRmTHtYOaGZ1VefLFpOlFV
yYQOULL9s8JpKF9isL5SXF2DzqfhynbgDfZ2i0I7SmsxX9ynKv+mSimxzwwJ9Vp4
tM5NJBJ2iRYC6fJTAliaZu/tHWfDeW3lLe8gh1YQfKIYRPi2nuMRNyKHDk/jG8mF
qdCAL5R4mETaCLiJ4zGVLcCkAf6LPGNqCuCUM4c4a0OkrWRmdIKK2CtW1MgXI+v9
AC2lpv+4+SHpKD/H5iPSLM9kq2+iNedIoR+vEa5YTP6IXGSZNrA3LFSOmaQ6EwqZ
w3Wnmyjm4xwWJJhpG3BVCyETJpphpwoizw38T5vWv8TSctfIdW3Mq+ygMyA9YqoT
TivxsyhCUd+mR3Nui4veiKNwIqBmlnwNwjAZT22vJDGQYvNH9xtCtQKBipRBYmXN
b35rPuXQpTBlj3c9y/LlAr7czNk/uDGkfbGoYfgTSoD3siWVFtMZLrsWbSeXOk91
EjE+NoU8N4hMp4EZyu198kn6/I8HOPOMjeBmToyzlyNfsZj0iFwrzwoteqhDGJy9
1jSc/9zQmfO36Cip6479op4QImki4Edp9otHTaFhfW/ft8OljBtwalWKIHOXoiCx
K2aLvM/nnLsVVFMjboLLOP/fNOk6ovcucoHa1ohJuGB3UtAuGgTYfgCafcL4LEl/
W9GA/aUe9mx2duOnQy1PNWAiCdwDhLc6DkLb2Vi5yNv2W2BoLajtsAgnpGMJpnJQ
JNIqURS6W66YWSvtEL+KbMSKHCAkLDr2ZfoUtOQtGSG5CKOnicavzc0soKz3upD3
mW+KfRrDufYaQnmTw13gWycta7QxnSDvDoehm1ytzrk03271b20+6wxe5sqPvkPs
PyrCn8pf/XntqraQe/Fj+r6IRU8pcSUltgx/0Z8ZUQjxOocGZXnr9rjJY03vQfxV
/4koP8eBWhEIItCOGTiMjOq49nQccidnSo0VbUKjfAB6tFjw86vnReztNxo+m0Br
xlsAuQjkKYNXDGAp4YqVN2d4hHHtE6NBYeEH+45/kIgcf5yhjMx6jJLZ9XdleF5x
FPjaUPAiUyXPuPYpJf6/F1ycrp5pUENDwDvMkZzxIhmODk689mtX6tNzLBGg174T
hFzVLrzKe7RBwgISf6S1wYkEfE4Wexvwf7MkQojQ4aLTxZ2WnCAH7qlm3H7vjoFE
Q/29IGdJLR90U1pZzsGoYkpZiBCIBbVF6LvslDJWeiEb8XcUeoRbi+I7qK5CPrfd
CVRI7cZTLYSJ/6dBofVau3iV/ej27g3ds8f8P6KAjQ4STyD0B/A4J7UKaFVTRSUb
JcCwknQZltP7w4lnjOeRL8yIoco49M5jYiHvEDCI8pWy43Hg1oJIs7fjVYSC3L2s
pMaWRty9tRnv7d1CPs8D6lbM+zdzQyLC2nmeDCLfaY5yICM3FpmXQDuGt9+wLpi0
nZvo4Cz02iwZzS/57GhUaXz1gv9OcAz4y2JK2x+y7ipnSMACi3mnShU8c9RttKUR
bMcM5UW8auyLpUJaNS8H0L6BeG0hW1RTY6Te0UA/D7dj8+fLvJtqEU6X/rS40W/8
lSfd3WQNQ2mHErvwLgilWXrd/vk0GrkproNO9hQWXjCJKjCY0NLZi0/PsoGCIt61
tIcJaTsJaOZo53X+ikMLYRiRp2hykefCwZGWjUNEmFF7ivplxatNCfqHwlwe2Xn0
zLirHG0+N91CkmEPC4eIH1+1QYakG9gsk/+PWba1i8GLbeAbyKissWVt7uDjPDfA
0zWqj76j/3nzwEq/9MjA/i6S5c+rXKxrV5QPQlcFZ0YeQgIMIwx8VgoVE6BsYYWW
AeZyAQtg3PLifSzpADaSkZClrsbW/cWihnO0J6m/o/NiQsBafinK9cM37y04Ukx3
oVQ2Y8rQB7gVFCnxoTFcioNK+U/wPw5NRAaO9Fu3BgXhKz9gyLA1qgCnkI0zL1tI
ADuNhkoD0hho8LvQHOeghmUb09kic1WTV7YH6iZbz3FzU2+jpYmZhKXZ57eSNsQy
stR03BYnM6jrRBQS6tabjeFVJ80kGhIa/k/QoCF85z/3Fx5gs+z3G2u8Kt0Hdpyj
kuxYC/hK4vZ/e+8UXeoIH/decpwtkiUzSbi96bwUMI56/2kffmXImyzC+TPI9Pcs
sAq/hP1wGOLfK2NqUezq/F59P8eqnC35w0MQeya24Tpn8qcy7VcK0Byx7GbgL+NJ
qCvZQjCg6ZWowH3lYdhOT6kWSr2Pn+f7VR3Sd18q9c9Ib2RVmCW+tNs+Vy3yNDyj
I1BZ5U3HBr9mUMedlAvi1cc1Xn/0LB8bN5iR0UTljNJ4+jZoBno/FkMxAPS1c0r1
YPSHgWuaq+1h5O4FIycHY6jABA6nmgr9pZ54vyIYZlVBFNZr+2jgF34+L76k8Iaa
FisSdavbdl24zPH7kPYUhAOMoaGDgNStOXe80EBI5VmagGLdYgBa//xmm/nl6wm0
hsrR7NBNt3j8V0MdxSPhMos/v/BEVjgEyObZcpM7gECL9slaUA0hJLcLVPMnUk6k
R2FSJ6iysWcUuQUFmywdcSP7xOGN7nQ4G8UTRM2JZaB1Iegm2UgobLXqFNFJqBP0
7Ia61WIz8gIWb/X75DHYRP8An9qJzED9tIzkTSZrga7Jx/JZqbkwCaL8etpP4N8D
3K5f0Q2KqDywrFVTo2tm7UGjqV+a4cBKN/5G5ZyOuKzeRgqVOOYjZbLiZF2r26DT
/10xrgC+Gi8o2RUP6BUS/TGHnIEB76oZ6E7yimOWC8co0w1jU63oTVo29dQzai2d
BJwdcfFYXzYmGZY/YqWRRjCM0Xh7BIGsPNdA2KnkHC8JCxykl6zGGI83ijEkUWEy
NqkZCfJOKo25knTL43vBUFFQoYTiHvPkAPbfj017d1FWo6tDrHadOZsDFDiJHMcF
OUoL+zez//FjRrQUVPXECcjrzmx26eyr3R6QVuM427Y/WCIHQA572Ho61G29Q+LA
4IrPEZzOYnY9J4xWu7WRhJ2UMlP7q9BHEWYMnR2x8Woi89LlnDXkUH6lNZTCRHPU
QmRzm+jnl5BVLXBLXYDTNPr3B/Q6Rz/+tsuEORiwjXreZdd7VYM04VaJjB9y5hRL
C22+6evysR6wDeO8Q9+hcPBkEil72+pjIEht//+mPH8UJ8vM4u1o57EqzPOKLkgu
PI7Ytr/xxCmXM9NIEjhpxweVSyDpk4GCXB0NQAJobZmbxa0BpfS3y6px15O77JrN
CZxHoqXFRf+LBlMsBpidDEm4DV/epHd50iRVn8zmwkwSxrDyiZwhBir7jGDhFB09
LisSjwW0gdcWzKbeOvJhemfTgFZ8wlTi0pfelip+OCyMrXBHF2LE2rGuUks6w5lh
Wxg4EIUGD6kck2EuJTn6Z9Nyvmdj5/U2qI1I6hgTgwlJnJ7LVNxPy1/sI4mwZPXd
GtkzP1ZpkmXEV5Dd7SYY+mUAUcsqAFkQxqPwbmmUepC9o6QJjgd1UOvvHo0ZIGW8
7t+o49BUQpkPInFIspALPX5AYUeGahs4ZG8PMJhcUhLRTm/VtMXDTEyFqork/mUv
IjJxYkFI1De3qG+jNHO3WuJP2Zb6gLEaKqqYPes0LrAXlov/xKQNqSxcXXifkxIp
onek1YQDxTPjJBPhBUjb6V0VmJrXi+DX2jcDfvss7Seln06q8bQ3PcCSrh3kM5r6
Ch1JvE48GwozXfWf4vAi7nOKrPdqy2nGvhiCIAMANj8KXyX4nZCTCs0jKFsTKhdm
B/vE1HGPPKEN0V2iqyW2byIdLLxUEX6SbVpITiZhIRNciA5VDZk31nt1kniT3rQ8
8a39GkyUkwk9lic0Mo4W+eQcJp+I46mZ4+Vsnj76heeAQDmJH8JKR66cJ18/rGIh
VaxprmiMUkoXwGJ9q82GhQz1v9E81bN4DS4EYVsCxIT3TWvHdjPA//8JrfKEeqHD
S4Xk22wP0wpDgkgXNFHQs2yty1nY4DAIECG2ZCrYAaQXHWw8sTuS48AxZ9uao+ju
iXr/wnEFP8t5gwbW41Wkp60XpHgQzxAGSdjdLypgRxUGn1owP3zxN0uVn4lmuyUp
Cr/NL5Q7y+If22G2kfVwAF6cRBLdx8sXF53+0ko8Di5z13hh8q81qt/A7W0zljJJ
yHBuAxVd1+bSuqa8rwO0kO0ftSASY4J9iQA/bG4rgYAuPgnU9bOwjNvqaSw3GPVU
0xzEzxUumKXaL3IJ6LypIhhC4u6rfNiyDZDBxslOedZSy7vZRz6Scti7xK1n2l31
65vR7nMCPtmDhmfgcKabukWxdirjpoEHF8DygwTkGSIVFYPpWcrX26bz1yAO6Pl2
vJ7FTpFLYyvZ1gt7QibzSUy8zE1C2S4AueQ+cwFRLeOEXvXnr1OkNUMpWarRUSaq
LQpmb+VRa0Ng00NmNCSwL1IEKuaLX0cE0duwnQ/GiXVNvMQTQ7UczFdpzE79RsV3
4FBBqTt8ClV+1FdmbyWPy6gLDHPP2BFdSIlevJAke5qd5qplalmfYtyYZj7h16pk
2WuCCa+kgqCl2ck5QLlrSPSePYQaSKhwJbf4hLA+UXH40tmgD5nPc/pN4RCBFWP8
D0VRADWdZiePpXPw07OXFUb7bUSCUWwlrgJaaP5n4Dfi4AoeiOrXercgeNkt+S8W
8IN9Lmjv+3MHyCh/JrGJvG4395y6oIP6sgzK5DDcQAWN6aHYku2sH6DBvd2dtFem
iiu1L53wDIK2IHIePZ++jOZaH4+Z+F4igzhO02HzzCLiMOT9v61ozC7/mkwKLLPo
edlxP1ul+W+SdFI05Ib1JNQUL51JuqiiCwB5QdZUdYYuQr4HSVHtVnQ1ZzhDxscX
RETCoJzAx66mGnU0KXJL977S/EqjOKk3ZPcPFjIJRbIY5Nc7X7oULXtKRxMHgAan
NTpqMpU0Siexmh1CZ2PQbn+/iiIngWE08oBh5VNds+gSkRO0D37QIciPXXMozvul
2Yn4Q/NplNyDL2YJSfDt3/0wBVYEmtSFgS4kfyEbwmlVoUcGtN2626q9s/Isevfv
GOYwhB8H7AOdlhpoGKAykQxARwt3BEvSnyV1L2N7VIbioNiR5XtGJw6Nvb4EXF1F
qM4xTOBN4F7RCaK/hKuCFt/wuwQugFNmX82KQwiwZJhda7xAamQEWea1UsgF9I7a
BcGTFZifB6RXyr3aemA1DjVaH+4orRp/h5zvBT3EWLcnNRkYlglIbm2Ezicdz9P+
OR4jeRKcU8r7n+o0bwQAh28y23Gq4ub9tkOXQ8y5aqgjloUjo77T9zDVy+UCpX+R
T4RSi9nWiLTYHPPdmr3Mus7YHYZ2huIHJH5c2ABxIwnB38NWwqpUDeiqTomMoqZy
dXPyq4Afqp6uYhBB47QxVby/qDrJFUtJkxlHKJhWtUmIsf1lYuekFGy0S1tBHdYb
N/c2R+e3ImwhhqdSo02dN3LJ29pBkK7mSIp/IIOCvQ8TUmyBmuRNX2aaagMZFCRV
2638DEFI3yIxh5Cyo/XYgbEh5RsXgIqxJg3xpLcW7Q+v4zCX99dxQWwkSd41Bowi
X/Dh9qXPKAVQreBQJsXqHnfOO/S82LAO1Mkr6sWnCEB8nJ2qg+uWgQug2/9/YmgX
Zpw3HRrkQmeea7AiiW3OVhLOp5/DmIkwfFs4Vw86alLt0UVROKxDY93AbCbjevCv
y7icJLAJrcRm1Lv8xGbOlGr0EPgrXFTJfSyWie2UHPoLH0ANOu1Gm712RdkDPGMA
xWcAkOzPn44w6oSxGa5km0Lui8Xmjrtfg6gRdXs23Eg327knaQKQeyMj157Mt+c5
xevoDIrET8utjDcCaFEl55M3OtEyqWEXS5APW7csqGretKxz5G3+YlWnLtmXJ9+P
ePahxSscXpVS94UdgLk/LK1LI0r7W+KVWxQtdpssziuX4jVpTYjmVZM2Pk1RjXBr
seuFfBW4vJUxludyHv+RucvEwcpfffdu0z7tzncBIo1c+iO07uzBZu77ekwDIhJR
yE0c4uuCntN+H/t2lM4GCcSLMRLBoILJT9mmUgrltVLnSWrgY0dsx9cIuByQd5C6
JwmtkhAUyOfe6hYtmbfnIGRwt0GNisKxxP4GickyV2axYHKt/0g7jeum7bCBzlw3
yscaOgqHh23LPGOBK59Q4H9VsYzwqqC6wXSNY7g+rpW95+7f3T02bUYddVI/VY6Y
gzYT0l0dXH0nS3sNADvfnYC7aQfsg8RYq81/ULtYv9gmZN+XAyMiYpp6BuT5uOiA
XiKwVAEIclFkFzlsW5K37ndOZZQBAPNLIjO2Upyo89FnZjH2KLWHruKmqFLPjHMR
lhyxE6m9z4oP6xwNKh4UP0yiEgksIJGAVduXgZuzp2XHHKfqqpLSfTE+ovJY45z8
YUKOQYgJ0SlBwd/Vn3X3ENMeUKYepWDi+wX3xawoV1J1+hD5t6SICcTH2qVBfo/v
iGyF8RvZrjYL2wBAB8NE8Vm9jcU/Q22Xx0SYbuh+dADPe43vCUbxEM4mi5p3k9tj
s5xBhAWwMALuZlRokylV5ne9lwh06Lsu3rVp6x8+B3OHCaOFF5yF7P1T/HHtj49L
kHR79KtCKuQCiC25Lyl9HwKLkxFyYKSw2GcIZcPvs/7U8aW9htv/dxiKfRFyH07l
Bj6NOiP6aE1f6QcKRWZppuRY0XRPB0quHakSgJcuZmAi8MwUZyOlG/2PJ+mk4nMX
SYFD8pkKYaABWH55alvbdddtLCaJKMJ2emdMGojWGMeMPvOH6FtCHujQ2nVHIsCF
BXm5WYwmsQBm+kXv43Ru8Usxr9WtFMgbSTPjcCoQd0mdFDwCcRPV61sE1C/gDWkB
IOXUYCmJoLONaESEqQAYvg0RSCYq4/vo+ll6JbnVmP8NCn+VeziE/OF829aqZU9m
ELMlhGqBBCDkIUkbnlYoa6hr/e1vmtPJMSpEgTz7rURbJ5NkvzwT434XhETZg2Fx
TMiYUe8z85/oMYlxSXhDvH6iYBioheQmoeDY6qPTuBXYsXTMnhnw2C0qLsuZN9vX
VGpUd4RsrKdDhC6ycpv5zLhw6DkWs0c6fR7tfSVSb0TQoAj3dOiZBT28TCSVPrDN
0Yi9f0NPBevGCfr/yc7kIHwe7vPLffGx/L7Gvo4gRnYwGagmxIijSSyoQhqmrMZP
fjHMUvhmblbbg7E+ZO+e9ofVORMEreAWJcsLzyR6Va6jtbHO9C9hJO4m6UO+3001
Ekl0QpzUqPedo5nsF1gzdAPVI0qsg7ecPj+IbucE00l1W/KZnb19XCUN+LPPJGim
qU9OS+DmxY+bxwHVyiy8Ry+zyt0SV5gDH1tRfZRSJhSinZPtCv7G+62z5oioQlWa
TMUUAL1vlH+OQQv7fjXLFlwJUVTo9b7TYkT6kVW0di74TkIBAJJWs4K9yNGmpeT4
hcPCCBRQHV7y8W00XDYQ9yDv8aS5BB42l0TA1gUbnMgW4hgIdn1WrPhr8YUKLwF4
Bxl2p8HWTi5cR2ZVQgw4CCmoC1qzh0pYi6nZt99KHsa/JYZhGOQyWHKS+aZ1lVBy
8AX0fOB08jPeXdHMrpWXdtnjj7/fm7FzvpGzPrshSeQwyzlDUh7r+PpnDIU+PrrL
pRqywGzD3GGG7m3nB7G3cfAz1+9THBCtbBgFdar530Yk0D2suW0K1/Rf/92rFnAt
qy1FGiQ/OESpL0DoJIreNdUgf1tCasGrCm0u9Wrajkm5V8CkeTrFx7HubvxcquRi
kcE4sKKU8LNmlU5INCfCgJ2GyZEojl7h7IBZ/0RCzxChw5guMvVB2ajGYF8WceiG
HQcD5PnGyzkrrH/q/XgwKiElNrmzu++4On/k7Yt3e7rSdfx6AP+Pw3ANihsSMSjI
yaWhQbyNkzpiO+FkqRRfE13Y1s5kZBDH3xcVCF2jgt/eHfHHjwyvV38sGBKuRmoE
+fOdgEjPyIoj3EGnKI7k+yqsR6WiE/QnS7RXIMLxD/KGlNPzx+nZaU2mJ1WP0S9k
xqoxGDuaHxkiftBB9HDlBBnh4uTsjf7dqBeSXShLXileNel/MYMQPforoZXam65A
sMx8+6Fj+B65hfhtIc5NyE8MUqt+t3aaxFNpEcQkEboL3fmbqyhtYDQFIFNPnuZ2
ZET/SBb687/18V9VsPoYDYbCzhbUtHCn5ZfYbmxGPPd74vuCH9ro7VxHqi9OKPfu
w3CR4Yrh+532HMp3sYemf6igcmpUWDGesbcD6Uz/01M/Mfu+/gUx/6d3A07SgfKM
hRYqva0myQBiU9OnZyjdXJ2s5ZKzS/vTsWpaRbmg75EPv3RHP6JQE8IWXRqsJVPE
1hA0eguKAtWC1wt4wdyz8RHOf77ljkObTU1jd/dbDw/BWlEX716dxe0t0qP4jO+3
jkRfmf8a68/Nmid3ED/T5I7bmcuACbDFtodVAGVCtilgIDk/jezgSOEpaIsWXg2f
cOPSDZWZbfbJNoNYIfbNdLZMYs4F8SlTuj6k0lVkeyfPOzC+nX/bj2DOITNG0HWl
oZIMnGDko1ZwQSIkheSR7fKioHDMLECdMtk1vN3upbxANemj0cgt7vLHtxuO5dRy
WaqUMmeNMAl/RksEAwOKHaox+j8vdoP1h1EealoMGnTOhdPbdL8bK99C0EnNKSF+
+UKV4kCMeey53Bnb4MblAMGm16svEyo7NrFPt4EBC+5/YlsprNA+FkYPXRi6k1HH
J/r20ZsYn0AKYo+E8VxAsyGWfz0OgAo+usnPcuwiKcHD5LRoAOCCpZ+r5zbsjgzN
N3oK/x8wHdrYtn2+OrkEYbE+fOo3C/NJhv1ughmlX9YI26vyuIjeWu42LRqLj/Cf
aRBCoYpvmEaI4MMShSuhYblMmRm+iiUl+mTubTlJTpRVXTKHy0s1C/gmjGm8BRc/
tZtjl+C9me9KXMAiiY95ZuHLhWbyFp1H4nzxXJsUoTKwNF4I0HGd5yhaoLd6cQ8d
GhOpBmVEbM1SDZheAfkUAIPsoAW3PfXVsFa1j/5jSSuuVAtiZ5YhdEgS0l4FNR96
CVBOnYzNMhVkmQIixqMebP49x1R/K2cXLhn6cx6lVDmb4ZLfW/U5jpE0dbcudHYt
98NyXi3QRC2Vd0vPpsbphJ7dtpuzJJXm5sC/rgYWu6PR1BwouOrOwU1Abiq/5fgK
OgTTUeQgVcimT68GzRFgksvSXc+xRfYpoesZPjP9d2CYviGLtnaaJfyitHCDsWI+
DSFtaO+fpvt6OynTmZNngOrnOXxpUj4ELcs/OatGd31cuxFZYj/gQI/K1EDxC114
JXAbiupIqpTUx/r1Qei53Q6qi4HE6LNzNfCgfQjbpuQKNQexPMRGbma7gxzT3rnA
mEjxjDTfGzNvgMzeFDNayTjwKsZx201X3SspJ8NJqZ0bJ+BMCKMom4QHAKbdPiaw
DiiRwLh/akzs2FyO5UkD8JZ1ajiC0+tfAdN6b+G6MTOIgGFTpobT4dwrzinOA4aU
+G/JggDz14DydWAxcDT4j6usWkbDCOnr9uS5PX/KoFOVS4DH4b3l62om0G3ZCsoO
W4d0Me8F0lBOokpOZMwMxewuY6FXsg1tFKjxCVfss+r7C+q1dKcauiNZCjbjuzt+
pNbCZz2BnJHkS4hJUp58lZH+8eVbBeEQRTQiv/LFzIHpYEr8vfFR5o8963DH5VxB
mIvZMjIRkuygBOxcFxx0o1xb8L8xg+tT5UqOE7L0OIpRP8BX4ZCufIu9h9cPvdqT
sIVfWGNkZupvjYo13DtGxM7DhzerL/UEO/xhsUcQRkbnxYMwIaw7NM3qAoUlXJEJ
IEf2Tdeg4NYJGB6jN/+/cu22asRVK7yGRn7CL4haEdoMOI9RCLBN7K1kk27gDX9s
GEnzpSZMzWDSTWwSWCXRi9e1VtxRauSK9P0k34vR44PUHqmEUBeZFBJG8ENg0Y1y
P9OwA1Vi5yUjQooWrfnzfxxHaL6/N5xBxR6mMVmt3iPMANaaqWi3+APW7019GSrz
6ZEScSYtb2ltd7BpWIwehHw8bHpivmhJQpW39Pbop7VhfG9MIM0e0rsDKpPuEY+i
+452+sQv7AvNZuKsm05crG7Sq0bFEclPY6p+q29RpOYhUl3iyp/DmvxcnMtULlKt
z3QRRIXF7u6kFwacqZS8JG76QlBhucbQFTbdm3fi3YSrLD294/CWa4C1btqjTXD0
pw2MLzqmpINXUJECDHcaOzgni377dWk/5Qj5kjADb9YohQssiLIv4BNzp+szTi0x
ve8omYJI29V5lGH1cpbdPDPF/papUURbMEF2u3xVF92DsZjXkCcN+UeIxrc66eDv
RNwe19mdtBoVnixxByGpvTKhUx0y/R+aI6YE40sl3zzFJCwsq/XFi7p1LH61I4JM
o87CChPREt5ZAQYfCXEKv/eBAUhYJoEloVP2cw5iWC9Ie3qk3WmFASAYj3IgoGGz
ZmSN292w4beLYZXb0pMpMgAPYx3YQWfE2RkqpBrRJHZM1SL8cNjQNJXWlBhO/08w
6RdxOoG5G4EH0LbcGpcbnr2M1dvt8Ej9OU7Om2fVy2z719Zw7Mh1XeJ5EoIysjVV
SKUWesa7a0w0l8g71+DIDLxC/bQC8KCDQ5qz3KgOMDz6T9QXqhUVwWRjxiSQuBwe
xvbPhlSWkhgcXtMh2ka0hGpn7D5T+/varIwoOCB/YlgjBWoFXIpxYMAa2JOYiEP2
1t+vHnBemMiX3+UIur3ZP5jbLsQVjYDTkfA2bAVxOIea5iqumspKMA1lx8QnDiQa
C6E9hvusOmnr0H59CRucXe77fiFe0pfbb8MNQ/3ajdH2UVFxBr3RDH736cFVYHN0
s04fP/dkJsKy/bpea6i2bq56op1U3igL0/YyiZVOjOhcxD645SptGDtkiDWTcX+t
7Z1ZwEQa9ncCyZTIeYO5BseLtHlckQe3I9FT7rBQog0FFisraeklm0dqpzr/lmUu
7I4L9c0TBsEtlWPIsx2mEb3Nt6KK1a1NAijUFapxFoFpAERFNNUpTuRpEyn9JfLo
JC12uyL0B7kLTNW3nySSBJ3X55AHwPl7pQKhG0Ne/rmeQkbPRD1fFBoRWR76ALFx
/xjHNtaeBcfXosl4up4IjhBnCzbrh73/Y/dvYDiH5L2j+t5RfrZL2H0NWYjmrNa+
JIw5MslUMCwZK6fV7wktBCRqGtyH4bPPglXNDrf0n3jLzVk6HFcei6CJSu2otTHP
a+eTmReU2tMzpgmlzcuKsKNqKrEryjXpiYqTuUkWzXphH5uvORR2MZBSSo4iVLw7
t0bBOjCtt6Dj/NjQGSgwemiIkDQ+0AmmGS9WJsSq8xVPl9JddUjG9oQdELQk4E/F
wK9pkVBocbWYJtF46A6PauhvgGHuds0XtMbxvcwxkguV0o9XWcFIucrO7HJxQMyG
mzzTBaaane9aXpygCi1WNQ==
`protect END_PROTECTED
