`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
P5TRRXkom/v54nAXI9nwWZO4n4Y2wReZvQQ0ODl9Fyqt8ReoL6WW5cVmZgaXmY4b
HN4RKKQCvehRQQJElgkVJL+bsXll0VwMrI0SsnC+mkm6MgWqqomyMFOjDWTaOBwH
GN9vBKVgY7lIt2d/1G4Ow5FDt8FjlgQ+zYnxKo6V+iuTvMvO84zfZx7SoxDI7Raf
HFNkCU82thfhKC4T5LY28OpGNMd14+B+E6BqYBNlWH/E2N/1s2T0J/Cp2F1KJCY5
QullBX+1dO7MZ2umZXl9sDnNrd/bx+nc/Lp7IRjAx7Q0DSwNDfSNoq3GXZJRvyrv
Fo8aR2d+kDmH9nIgKQyETazn0BW7aHBg/Kih6ETzxxPP4ze1y2js/46byYiy/E73
rDrTMNedj2q3tuNsI1M392KBbtYhokX4fps0z48UkF6V5BgDqAbGiWOjSn0Ciu7m
iMAiOuQNDo9PdywnyCFgalrG/fvv1U09ci4LMSGpgSGZzwgH1JUEyx/oOhZK2XK3
4/Pooz9a4PobvYANLyBKizg673nX0x0lLLPoK7wQUhqQO/Cze1pM7onaN1g9bviv
tKUo4FKT/3/k9Qtjj93IQP6W18AC+1Atk2cON8Ig0uBzYVcQ8vRU6LTx0QGtzS7/
WA+srW7F4N1gI32N7/UpjxRz1jH09P8CZgBpAqYLI51yQXLAPw5ybcfrLFzj9euJ
RHl+Kaca/2/tZqoG+jwmKlJWMKn6Zh5k1c9imXhLb6TFtXmgbJcgM5C6xifNi0kH
67DPemdO6Tzfbiyb0EVLuujux6w3j0Wh+uQSg0eSf50NPk/8F6gjc5HVD7W7v5M9
1tsf3Dh5IOEmw4UTj9hlNfUgsQ7RF11cxwDnYCkvl+MACOYb8O8LLYkr7jPopi9x
aFFag8hl0bAMtO87w8pLy6g1OFJoXEixTb1SpUakY6eksw2V8Q1x8A2mZOvjs62Y
rxXDeIh7q8gTMmECJ4F/LYT9e9SDcNKQxVOKq/0x06wk553V7RRVNM1WOlO0IceW
Ys/7cLB8p4PNKM6AQ6tbL8nM1UGTl6PQjOWSEtP/NqHnp6N9Cg4XkH/nCqmHSG5R
9iaTBUPf/JAtpCp7BaTx0ndbyJZWqWYIBlawiYr87giMD6IZoD0PQktgGgG7Xr1S
fiOOOe8lzKvX/quJxvjdHtNTD/u1ktu49hjc0NpBqIf40NFfnf0dPKZR/0bWfdKQ
w9JdWqjfvE/Dp+2jabiQpAPQhwIBbMuDmGgKYFQSpWDgFV/+qAmC2jb7e/6kdNvw
BNhNlkYWMEcKiqXzSPr4zH4ehAkNON7dbR6CNNNF4sUNPc0Ly2WOdvVo7SqhvS4s
ubxe4amyAqUMLHXLASRVfGIVYfF34AYL32LV+Tb4KjniMYSy911KDtUP7CcwjnVc
+XjL9S7LzvdyC0SfOywXpRGWmW3YyqpS/MaXCggvvOmzmImvaUaWtoylPz5iFZjj
uu+wm4k52WQ1cBwcLgyz890HoGwWVlYlTvtrt/NxoqQOvvXmLR+FIQMuLbCG0kOt
vvjUSfu8TIEnUm04AoWWP3hVkXHkE+zl0FY2iRgsoLAke475EEPU30cdES7a/qXx
WmxeOV98dUOsGWtZXDBf5MrpXauc8Y+U6QB6et+skBa/XaDHFmzWsgLIvNgBt87g
g0OnxY9rNn7XrawrfOs4PYVxfA90vYcw39kDdkM8lpUOhyg3YWeph8REaRVjPy5j
wy2RP1UOdOdeSiAdCNcZFzc9LyM4FMx5a2+0GU22EDYR1FcGXJpH09UNsduy/Ac6
6JTLYHOPj+++dRnPyCuLEDfjKdUxg3mxagKsNeVSpdEiANSXDKZyy52dU9Rz3GBh
LrODYwpSd4ziaHYfFdXjhaj6ZbEIOa0K7pkkjJd2vgOr/9vFa5myKjgNPTJ0XynR
eJAa1HMdB8sYiz37n+R19qpS77lwpuv+Bw2Fs0wWQ5CmvLH+owUFpBVlcazsSfG9
L0FJsLFnCWAZ6STGwbXFc9ZaYDcWuqooSx8bvAHgKQux86fUrU1RGM5zRw0pOyaL
Wourj7shgpah6pHyNib0SvKw9W0EtPec9ZzVZcV07G53o1iESHrAu72tc6F1sIpg
AJv2Dny83OglBD0py0FvNPZwOzRGtttKqsrGKYGWouCrmPeOEr8OvtTtC0smQ5bR
xYYCyxWwSgXP0YVPT/DsgjJL/zAX0byOlkEkZp0Zkp3GnZjTqbcCb7L2Zb2djXEu
flmDC3eIRNEQ3pWAqqfKrC4kB2dVYFt4I+vfE9dxpEJ+p4M6Yj0vvXchFgWTwQwJ
wdBOYuRPYArAxVxSpVXb3Jy9zDJfCG+laBgj2gD6eiVlBem3PsqZvynp0uARDCcS
aABTFmmRGsleODc7jyDsx+UaAKXbm7Xwf28zaqQzdELBTqqnG5JSGC3/4ECj2GTi
7OOdoMseIOAJQHFbejlWXwTMKB4wQQ7H0FAYQ4/o7KrkP9Picc+7KKF43R9iU0yl
1KP9wEUlFkpkZdOvP2WkKGH7LHapMv5WUz+bsIzjqqY=
`protect END_PROTECTED
