`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FVwQMs/9c2FPnIWTLV1hvSqs2oBO+QW+4eaPMtBTMMyUH63GqGP/gcH6jwJY/2P4
2vv/ASYw5DtwnLtt5OzpIbHwo6Sm0EwoSd1Q9EmjR4Cu6C9WtGn+/RHiu2qiiJu/
tKbnNfbO81pFiJhbQo7AyDXfAeW4L5980AUNc6MbbLRMRnCCZ7l7g0N3Iqf6EDrZ
ta9POzlHCN/C23A9X/AwWjuI9qm1KHXkAjkMOe6eDszgTBdOV9Jx/dH9QVoPSSVV
z96fkkgIbrWwmgMI7uYBk9GiWbvdxAyuaOC/yrXDTsIZqsAOReB8L0jvSE3YII0L
eVFA/8jcICPikWk6tD5NIiRCntgu7Ly8J6BFee7wvvUxBiR4YOg2yfkt4irHLU1m
N0ekDHJXn2Dl1d4mAhSo+w1qRBno1+5x8yzILSk3jJ+oUSG5PCIrJVzYIZ1hrsv9
zfsY4zTFJ2fBrIwkq0rsokJzpZLDhDkCRuDetkceUMj5nkBVCHocidYVO/UcnUW1
k3Lmb4f1U13TIdnb4C3veE2vu/b7If6sR6jgAVtPkVZzYRZqZEafB8VJgResTi9E
FgbveTw+kMPFu04ISGSur/QKiU/IL/f5ZdsjREz4M8tHngKZ9zMKHv0Sj5uuRcJU
+QJO5oYAshUsC0mjVCl29mJoAuZtuLlNzuM2oAqD7YaU/7CTtn8JEmbAlixi19yr
4Ahp5CzEPdAkREjLvDaD1BRWmBjIvUfuFleTixADEEQoMWqdHJzlSHOOS8tksnX6
XcWZqHMV+T0ZR9m7Jf/kGNKDgEuanWxDAknsAAMqj/DFzzl0y2J39vj5n4aPtTBw
QlNACaKhAfVGcSwXJ+zLYEwewqWGVEsQMmFkTypr8Rx/VxtYjqxG9AKBCTGPUHYR
lDEV618uXsHOVrDuIVVINsHQCKzwgPS9vbzE2BGGARiq1RIon/z2oWbmOQ5rwlw8
jPkJ8yZtsBvGo7HooPx6xf+65HVhISx4yZ89k9xCYTZ1R2laIW4dzlQN1GKR1DMT
vEmeYuKiEPf9JzfhCCMnFnA9/VgHZeoRs+eC+mWR2uqKGbS44zcw6uptUGeDx0Vj
vso7mQYZUTG+3IgNutNArcNcmM9Ia4NlGpK/FwrIEjPLBXOKTKTRbelghe5wSQIO
KspC+ZpqL4iVXbPuzeI6vIZKwyLSVjKL8oc2Be1Hd9rLnCLuHt0CZePnPdciJTNY
5HzieH3v3iiV92pDWWv0jB55H7VQWSYLWknvyVfmW/5kGvWWDO63SrkV0A80IAKu
saYgIKb39uevWCMLNG4Laz5kCTo1Fxv5ffDfVUAz+IU/J3HBPyZ/FJ3h8cxXuphO
OTHeR/NNwN5JXox2Zh75ZCr6IMSpFlP/SCS2DNIH5HWAtEqW+A5Gfu1hPpRcoaNw
62DpchEmtCkegUWpabFhLDfapN9ElI7YY+AKwqu9Qdo0JsRwLJ8XUgK2q/SxzuB1
re355kp1vJZKeYI9PMTUARBc+F51c6WFDFYjk9zL1bikeBh5j2Iy6B1yyiAmwlzF
ltPRprjZsPgx9/JJS3oCQUucF1sm0borkDlfeaZLIeKhtpq57+Zy0BqdvLLZuBvJ
aGifQ82qzBgeIC6gEdgDKA==
`protect END_PROTECTED
