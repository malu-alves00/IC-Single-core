`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bOFuWU6rlDh1BiRh+KKopllyvdLat25JOQ4WRjHBYTVLl63+8+fBSOjpZQ6VehKT
iOXZN17W09CS+E/r4kMHuvQ45lL3aIPplRqbus0z5+YPFEOO5orAs0WjanFOrhmz
uCqcYgWppDchuaJxhO345EXa0eAYZbuFHXBPOfiupt+QqN6uBhemIKkYOxLo6GOL
3l0zugNcn9Dz3gwKMwgkr27sEjpZlzi2RK48K+vP29VMA6XeySMDtZLz98uPIOxC
DCpZVa3hc2idlLNz+ba3bhDd1PePDiID8xzXXsSkkCgkFBJ5/kXbv3TeJiLofaAW
3THwxGvlmt8XeymJoKu8dpRovLFBEXza9wA0ugHQV3T+Depk+Jg4yn7OQ4NuYyzA
D/gmDS1f1HHLtfsPHwuJBZrYfenskqN7/1hXVA1XURDbLJyhcB11b2tfqDyZSGkU
uUHiOVViIQfO5dGO3nqOGRRadjJSyNzgBaBYn6jF5aw=
`protect END_PROTECTED
