`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jizRnI0Wai4ixWMr3bfEpAw29YhDqUYVS1X0Jr73SATa+sUwvXhFO8CpipCXsyEC
g+At9q4aw7TQ3+/wq4kRern6fOU9rnAN8gUk6qiwJHe2gqfCUVqfuNt63N6elO11
BrkVHjQ1s5JmEUsacPjltpJsgaEWhnhFGdXmag8qhPIgFnKKUaXRxw6rgJ6UXZGV
Wlw471XTE332/4qUa64KkyzgSsy4onlZBmHH62WsHPwfBVnfCT/iZMVXMpoHtFOu
j1l5Y4QnIPYAyn7FJmrs5aIOLjbzREs077Ge4FsEjpUOZhz1ea/MRyPYIYyDGdeg
gB3fgIln3YlfETv1iJf/FxxH80thrs2I4oC37EaSNS92YFsp9mw+c5td1J38sonx
kl8D/fxErx+PDJnLcLchhN284AyT+E9kMAzXfJiZLT0E73utM8tcP34LUdsJ73AM
hdMbBcumz9tm+6+xdjFnnBappf9oXsPjrkWRDjn9h3sdCzfCJh1T8bhpDXTX0UuX
Q07x1OhtOuafDq1eX0ZH2VgVleaE0ecbTfq5QgIeyh0XABP/T70NrzrmwIoepR+V
NnxsU7RK6XXvugU9SloqiMGqdXtMKd2hh5qR2HrgKW+krJL5yilN5eebZANU4GhB
dRwhg7PKfIGR9GkB6+cLhQ==
`protect END_PROTECTED
