`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RftSQUED+QTuhfYBROFXPMm1p3CznlnLVWZZqP3xTt6Vi5D3TG9p4TOr0nia4jqS
lj5fRzKsgr7HiFQMNBiDx9tBQN/5WAzaLIdow4rwSQUhYBwGFModaSiKTv1QPbJS
pMHACqRWlhjq2n1pKbqwYY+9jeHqhrOQSn3TKwHU6HmHcKQA5ZgeGKVgoL1gDTyz
C6pxxRvIR0km5Kl3ZsgAy3BsmEx/RAULsGyvNyAm4WCnOzwjBPyu/n6SCuUCiK0B
MbfhaMjHSccC8Zl7amCapHgdzrUdWWNFa9GaDJiByfGUX8EYhyKRiw96srU2dcHR
kAnQstK1C2aOR0GpHBlPDQ==
`protect END_PROTECTED
