`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jOPtcPolOJrDpeuCL0t3WhTtoWdXhLm/CUH05EP+ta7x+c9NDDBWWsysJlHlQ11S
4szT+x0CCfTS1LZB2+IjaXqzYQuqZlO1KbOYbb1LuAg12MNcjyD8Iv/szq7/9UXO
8DHmQIeJRbfhTcgt0HL0MwF52TOfxJgROxjrV11IZiaokoywlHdg//378r8RY1En
2Hulh4xoU/OqAVd/IwTE5VMh384cuk1nD09aWhc/M/aIyQ0FxqzKRP0zV5LaZWdC
R1U4B4fMbwtAUthhIcR7ghfGyOxKGleO7+LvKq+VdqilC/pKMmYadsto56CmBN5+
WOEujWgtfomFCO4Q5WxoKeVTF+jYJGgh00Ey1lZA2VJxc75NzFDbQR7v2tSc8HkC
xh15gl3ucQTFBpsBPHlo2L3FR1RKrnP/EFKOsuqc7A0IT1s/5GzGS1vWhXy0k35T
yfX+v2z8gbuUR7lPCnc5zNOYqTLnlE6dYAOHUvLxOcIwIyY9BBnjo+966E9Pd9sT
SUz9lI6dYpwaN1lEhbIMHzOpyUO23SqGdb5zat5+daPMZ7ndLI9ZDf5vZORbqWhU
lDf7Aq0NkTXAE7w2Z9hnS5PrMwF97TogzINu+bI7dgT1Jk5OuBJZNWQywHX1giTC
ollEiDxTtjI9WPwsm94WgRSoO7dXIewT3nVvqce4PU/hOaGJDfWUThizpZe08Dfm
Z2CM2We7CUhACih2GEkhLy7e5V3/Cs/Cxy8IFP7s9oIXjONcJQeX1wpfKcgWJmp8
uhLFhg/GekXd4bBVN8BwPCqoJjIfYYzbYUrCvxqbaPoYYPygxaGnJWumr1oV8jJu
y2hE8x/EUwncaAcGhwZIFeX5Ijt1m5z2LM9z/4YwPv+ykU4eQTOFhQfu9yGzjox7
eYLqYiOXcvMTeqYRsJ9hjIWVwTcRkvv2jIUUDQSBsS65kcY70M1pu9H65wzOrwTs
1Du1z/u5qKT4qUtxyZYcTLWPpujIo3QUXiv9pQAAmS5MG2U+A9tik4A/Bop05Yvi
Y/GAQz0mAO/+h3eWNE5gFKrpf6cjQdprfDMhscyhiaREq3QFTIpt5dAAiMl+kcaC
cEnjOzjSPz/l1Tz5Wzj5Ie7uzWcgFp0L7Di2Ay9vU7ixSFWbqRJxYeV0hEjSDigG
JUZZIR+8fAmA8vVagjF54AaWaDxiNQPn4bg67U2JKw8I5Z6mutHMnM9UAgFtz9+y
WF+ccnFtQ5O2pnagWdrAQkjYBjztf23b7jsFkXkDdA/0c+/QVpxQyN5+jwS586MZ
oWymn1sfsG0BQBkAOs+B/4p9NjW0U7f4yx5eiQ9InGs2Xvf1y4rAPZjAYsrXamLv
`protect END_PROTECTED
