library verilog;
use verilog.vl_types.all;
entity cyclonev_hssi_common_pld_pcs_interface is
    generic(
        enable_debug_info: string  := "false";
        hip_enable      : string  := "hip_disable";
        hrdrstctrl_en_cfgusr: string  := "hrst_dis_cfgusr";
        pld_side_reserved_source10: string  := "pld_res10";
        pld_side_data_source: string  := "pld";
        pld_side_reserved_source0: string  := "pld_res0";
        pld_side_reserved_source1: string  := "pld_res1";
        pld_side_reserved_source2: string  := "pld_res2";
        pld_side_reserved_source3: string  := "pld_res3";
        pld_side_reserved_source4: string  := "pld_res4";
        pld_side_reserved_source5: string  := "pld_res5";
        pld_side_reserved_source6: string  := "pld_res6";
        pld_side_reserved_source7: string  := "pld_res7";
        pld_side_reserved_source8: string  := "pld_res8";
        pld_side_reserved_source9: string  := "pld_res9";
        hrdrstctrl_en_cfg: string  := "hrst_dis_cfg";
        testbus_sel     : string  := "eight_g_pcs";
        usrmode_sel4rst : string  := "usermode";
        pld_side_reserved_source11: string  := "pld_res11";
        avmm_group_channel_index: integer := 0;
        use_default_base_address: string  := "true";
        user_base_address: integer := 0
    );
    port(
        emsipcomin      : in     vl_logic_vector(37 downto 0);
        pcs8gchnltestbusout: in     vl_logic_vector(19 downto 0);
        pcs8gphystatus  : in     vl_logic_vector(0 downto 0);
        pcs8gpldextraout: in     vl_logic_vector(2 downto 0);
        pcs8grxelecidle : in     vl_logic_vector(0 downto 0);
        pcs8grxstatus   : in     vl_logic_vector(2 downto 0);
        pcs8grxvalid    : in     vl_logic_vector(0 downto 0);
        pcs8gtestso     : in     vl_logic_vector(5 downto 0);
        pcsaggtestso    : in     vl_logic_vector(0 downto 0);
        pcspmaiftestso  : in     vl_logic_vector(0 downto 0);
        pcspmaiftestbusout: in     vl_logic_vector(9 downto 0);
        pld8gpowerdown  : in     vl_logic_vector(1 downto 0);
        pld8gprbsciden  : in     vl_logic_vector(0 downto 0);
        pld8grefclkdig  : in     vl_logic_vector(0 downto 0);
        pld8grefclkdig2 : in     vl_logic_vector(0 downto 0);
        pld8grxpolarity : in     vl_logic_vector(0 downto 0);
        pld8gtxdeemph   : in     vl_logic_vector(0 downto 0);
        pld8gtxdetectrxloopback: in     vl_logic_vector(0 downto 0);
        pld8gtxelecidle : in     vl_logic_vector(0 downto 0);
        pld8gtxmargin   : in     vl_logic_vector(2 downto 0);
        pld8gtxswing    : in     vl_logic_vector(0 downto 0);
        pldaggrefclkdig : in     vl_logic_vector(0 downto 0);
        pldeidleinfersel: in     vl_logic_vector(2 downto 0);
        pldhclkin       : in     vl_logic_vector(0 downto 0);
        pldltr          : in     vl_logic_vector(0 downto 0);
        pldpartialreconfigin: in     vl_logic_vector(0 downto 0);
        pldpcspmaifrefclkdig: in     vl_logic_vector(0 downto 0);
        pldrate         : in     vl_logic_vector(0 downto 0);
        pldreservedin   : in     vl_logic_vector(11 downto 0);
        pldscanmoden    : in     vl_logic_vector(0 downto 0);
        pldscanshiftn   : in     vl_logic_vector(0 downto 0);
        pmaclklow       : in     vl_logic_vector(0 downto 0);
        pmafref         : in     vl_logic_vector(0 downto 0);
        emsipcomclkout  : out    vl_logic_vector(2 downto 0);
        emsipcomout     : out    vl_logic_vector(26 downto 0);
        emsipenablediocsrrdydly: out    vl_logic_vector(0 downto 0);
        pcs8geidleinfersel: out    vl_logic_vector(2 downto 0);
        pcs8ghardreset  : out    vl_logic_vector(0 downto 0);
        pcs8gltr        : out    vl_logic_vector(0 downto 0);
        pcs8gpldextrain : out    vl_logic_vector(3 downto 0);
        pcs8gpowerdown  : out    vl_logic_vector(1 downto 0);
        pcs8gprbsciden  : out    vl_logic_vector(0 downto 0);
        pcs8grate       : out    vl_logic_vector(0 downto 0);
        pcs8grefclkdig  : out    vl_logic_vector(0 downto 0);
        pcs8grefclkdig2 : out    vl_logic_vector(0 downto 0);
        pcs8grxpolarity : out    vl_logic_vector(0 downto 0);
        pcs8gscanmoden  : out    vl_logic_vector(0 downto 0);
        pcs8gscanshift  : out    vl_logic_vector(0 downto 0);
        pcs8gtestsi     : out    vl_logic_vector(5 downto 0);
        pcs8gtxdeemph   : out    vl_logic_vector(0 downto 0);
        pcs8gtxdetectrxloopback: out    vl_logic_vector(0 downto 0);
        pcs8gtxelecidle : out    vl_logic_vector(0 downto 0);
        pcs8gtxmargin   : out    vl_logic_vector(2 downto 0);
        pcs8gtxswing    : out    vl_logic_vector(0 downto 0);
        pcsaggrefclkdig : out    vl_logic_vector(0 downto 0);
        pcsaggscanmoden : out    vl_logic_vector(0 downto 0);
        pcsaggscanshift : out    vl_logic_vector(0 downto 0);
        pcsaggtestsi    : out    vl_logic_vector(0 downto 0);
        pcspcspmaifrefclkdig: out    vl_logic_vector(0 downto 0);
        pcspcspmaifscanmoden: out    vl_logic_vector(0 downto 0);
        pcspcspmaifscanshiftn: out    vl_logic_vector(0 downto 0);
        pcspmaifhardreset: out    vl_logic_vector(0 downto 0);
        pcspmaiftestsi  : out    vl_logic_vector(0 downto 0);
        pld8gphystatus  : out    vl_logic_vector(0 downto 0);
        pld8grxelecidle : out    vl_logic_vector(0 downto 0);
        pld8grxstatus   : out    vl_logic_vector(2 downto 0);
        pld8grxvalid    : out    vl_logic_vector(0 downto 0);
        pldclklow       : out    vl_logic_vector(0 downto 0);
        pldfref         : out    vl_logic_vector(0 downto 0);
        pldnfrzdrv      : out    vl_logic_vector(0 downto 0);
        pldpartialreconfigout: out    vl_logic_vector(0 downto 0);
        pldreservedout  : out    vl_logic_vector(10 downto 0);
        pldtestdata     : out    vl_logic_vector(19 downto 0);
        rstsel          : out    vl_logic_vector(0 downto 0);
        usrrstsel       : out    vl_logic_vector(0 downto 0);
        asynchdatain    : out    vl_logic_vector(0 downto 0);
        avmmaddress     : in     vl_logic_vector(10 downto 0);
        avmmbyteen      : in     vl_logic_vector(1 downto 0);
        avmmrstn        : in     vl_logic_vector(0 downto 0);
        avmmclk         : in     vl_logic_vector(0 downto 0);
        avmmread        : in     vl_logic_vector(0 downto 0);
        avmmwrite       : in     vl_logic_vector(0 downto 0);
        avmmwritedata   : in     vl_logic_vector(15 downto 0);
        avmmreaddata    : out    vl_logic_vector(15 downto 0);
        blockselect     : out    vl_logic_vector(0 downto 0)
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of enable_debug_info : constant is 1;
    attribute mti_svvh_generic_type of hip_enable : constant is 1;
    attribute mti_svvh_generic_type of hrdrstctrl_en_cfgusr : constant is 1;
    attribute mti_svvh_generic_type of pld_side_reserved_source10 : constant is 1;
    attribute mti_svvh_generic_type of pld_side_data_source : constant is 1;
    attribute mti_svvh_generic_type of pld_side_reserved_source0 : constant is 1;
    attribute mti_svvh_generic_type of pld_side_reserved_source1 : constant is 1;
    attribute mti_svvh_generic_type of pld_side_reserved_source2 : constant is 1;
    attribute mti_svvh_generic_type of pld_side_reserved_source3 : constant is 1;
    attribute mti_svvh_generic_type of pld_side_reserved_source4 : constant is 1;
    attribute mti_svvh_generic_type of pld_side_reserved_source5 : constant is 1;
    attribute mti_svvh_generic_type of pld_side_reserved_source6 : constant is 1;
    attribute mti_svvh_generic_type of pld_side_reserved_source7 : constant is 1;
    attribute mti_svvh_generic_type of pld_side_reserved_source8 : constant is 1;
    attribute mti_svvh_generic_type of pld_side_reserved_source9 : constant is 1;
    attribute mti_svvh_generic_type of hrdrstctrl_en_cfg : constant is 1;
    attribute mti_svvh_generic_type of testbus_sel : constant is 1;
    attribute mti_svvh_generic_type of usrmode_sel4rst : constant is 1;
    attribute mti_svvh_generic_type of pld_side_reserved_source11 : constant is 1;
    attribute mti_svvh_generic_type of avmm_group_channel_index : constant is 1;
    attribute mti_svvh_generic_type of use_default_base_address : constant is 1;
    attribute mti_svvh_generic_type of user_base_address : constant is 1;
end cyclonev_hssi_common_pld_pcs_interface;
