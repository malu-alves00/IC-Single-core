`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ONTUHz3GZ2eHen124ivUjUqiN1fy37fNYPi9qV0puZs41RMkKBvfJXxfN7ZWgSWy
YSiQJmOSJZuTqUs0dSiEsSZ7xHn6xCHqXvjGCeHmXVipSa3cSeLJB7K6dpzjhlQd
NsL0IOVm4XEtJ/vkSU9tox0nJgTP8V6srunNX35bPxDxMX2PC36I5BWH0hxPcmaH
TPloi6E8l2jTOsEj6sVGsSYK8UZ+8VW9N/0gZL9Y2xnE4/0abIbGkg8b47zabWNq
HDreHaEBI/GIKttb+zb0zLa9zcUbqK8bpH1bXF/raZeNZIEXpx6diKiOFu76pa9O
WLxsD/KhxYvL5kcdnfB2a5D8HCx6NS/qtqKINvlUS45pFoVMhpO0o8XBadCqQr2r
2nqBCOhrANphU9Yf2coOTYd8TfHqs9Zvfl/AAY1rE+078N6RIgZKpsbVsJIkIm4w
XoWv7l3800WUgLWnxzManGg5qxNEWwPZfzD28FTLL1BImkPuddZM6/PUwwQLk5gx
FmDZ8BCJ2YO+Leod9F1wfhzViduUm5G7bE67/BCej4vMjoIdTdjaAGU8WQVuz2Dj
m7utnDy0GmKHLyTNnXtXdkq2BP6S1NeDPDCJUy1QeaPgvQwSvs+Ishm/07Jj/AaX
ZYXSJC6EvXMG8irn4RvlNIpf/+fUiSYaATIj2mJFet+Pj7eaQnD521PifwNXy8Cd
MXpjjfCRynq2EVzcrIy09xT4ONVWZ6txXApKU93JHIdIKyZG/w5EUfv6KGIaWtOP
3qZtcxdaulrG4UjlZpsDKys5Yn1CF44TCWmysw0DKhu5jHVXYdxmf4WRXMpMba5C
5v0oAjzsDHXHxZNJv3YANIKvHEe9uazyOTUbbooiD2A8OG1XZ30LOBjUBiWYf7qb
m0TtCdzO/9Oy47AJYvwIzpxdiY0gWwlUo2iiwGk/bYsF2hwB4gIChZHeEOXjAEyz
X2vDsTXYXJF4zzRX8aL9aUEG3vGM7PpvfhrcPomaGYs9GCCFBTFqzM+LeaqYXc4l
P0ZuyYUPrfKBVbvKsVgz3MNFVG7S5n9uJPOGnkG+drNrJv5ngdO0uM1Rtrm7QK6Q
CkPA8sPQ/iLubszX+axl4N3esxC/aWezWdFigrR8uwZrhVnVWaCNaTHRLfWtay2E
baoQ0ogFuoo5eZ9eBtCMk3HrcJeu49JOXORpeoiadpUfktvI3mYvL89fPjuo04B5
0gxAUWooVVU1hq3H454www==
`protect END_PROTECTED
