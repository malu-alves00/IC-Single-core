`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6e8cFWoPFK/AFDDkAjMC0R+eyDPErO1eRYarJ5MS2zUPb+LGMWgHw7H5qCWeCSB2
FdTdmWpK2jb+rjarJYgkxxnRM8oGBIhiMMYh1nCFMLMsoMP/rBmOBOLCH+abuhWP
HLmKkKMX9xU2k5ejNTsf/xs6E7FvvsdtMm8uIAufbCH7JEBBlbVVf8qyAZ3k++1i
Zm16THc37FNiVy5JlLmFh5u/SzequNiljaa9rkKcC4PqhvvA7TFnZwjPZSGr2O/q
L3sHyHZ9nXFAjO02NshMxZYQOeP2/8v8WE/oD2VC9jmDgvnb+tqMRRT/bylZFS1y
UMZauKWXrxqsw3+psv5sqK5baHxzk2EKs+3xISikhrnHUbQW5dR0yorYPLKRdrum
7cNeOZEyLwk3LCveHr8yVG3sTYodzB/JeNWxUHkwLD2d9rW+W38oamC6HeIDoVVO
RVtcaU966PhX1UIr4JU8HvkJdMjPulqYj+1tES8OcM9VatPRIhyiPWsGzwYjFgfN
tn8+ecHQiZapXUykhlcOjIf0OTGWgf+ZdzCT1JwwzRC3AnWNgkY/1x0JIdKKUJa+
Xz1EENu8yG8g8tEIrMYzTUCwj5qL4bLGFB/ZEr5rswwGtIbUm5bngTHwvv/ZApWw
Vi0vTUFKezHBPOVyFu7h2GYJdAEp2tPKkF8UDpdl+AJ0M7D4eotWJSE4d0P8p/ra
hk9PS7MDMb2zqc1GqVxJZGe6pwCiZ8oCOyfWlRBgGt7z6PlhD1uMX/PxtKke+XsM
nSj0rCvCWwhwhgm109a27NW6SdGCcd07DicbS78Ac7IsMHCe344DOAztW6WtzWDx
tLwJTExpkODNWbbvm5HUm/rPxQnIgp6GIPVy8zx3gFxNzQvUywnD9zlFNxLymSit
tpuCObEcrfR29LQkeAWc6seK53RP871iEqvNxoV7Z8X8t+KIOc8T7auRY8BgJZtk
EhZeJQ5YvcAG2JjgC2Xqu5SY0fei6q99P2wN84Ht/bTb1vllqp9xGIEHY82OFJZ5
ugtreuQH8yp3DiRGycf4xPHR3gXhUSH/INlAGhXdHFAo1E5tYw1rZzHLlUvtrt1d
+12qABIrFZKdZyqzr6UJjVOEcdB2KaloB2LJuYzhBbelA0r0mi71k26NOIGzv+3k
jhQTTdUtOkEw/mZa059JxZMtM0r8FxccrJttlS4z5BzyLAM//spH9SQwFWQRpiP6
ID35rKJchQ39mSkDR6Z+HTXqCqRkHgQfpqrfoP/FB1sDNfnLhHq77wvIrrBND+4h
J+iDfL9mGqPWBcyFmhC6NtfcPWW/A+Q5umBli65dt2kW8pZKarRhpr6urJ+RdYbV
xYFbpYYSygN0bBv1r15yGzgsAHCOINUSlynCHZGnW/zdvaLz/e2pKZGBpyre16Mz
b+g8vHKX1AIFS867rn2z7OCI1MI8IcSkh0ydYH1pE+zQOUw7Q7FhRrReKnSrjq1G
/8/5r+HdDzauxmWb5ejjJ85x4SZPCvIm1DfBXVMfEpkhaS7QAeCUjTP7+GOZVeKV
2vSbhfA+KOGTGx8E7M6V2TIVDlr/wMVjam81/adJ7rHCdxisHAYZWxGC4OTAjnsm
mDxSzswhH+cv9kC111eJrENWe3STvbi3D/4+vz8jw3dMOnrEKRi26UMF/U8lB4Xt
7Knsow5DRdWfK4kZlkEQFIe79UMeC5xKZB6X3te6VYWeCoOH3bXy109AcVcRSePw
j4R6mwSDv+yK14ngCQiJV9W2w7M4eSdVPZXYgqb9F9euKUqs5qZvaBPjMMICagtT
wOwY1xmCIt2UW1Gky0lV5BtMpWNcVzd1EICb+WO/D7ibrK+GVKntBKnqr9IGc/mm
qCGkkojnvSruSrBdc6rJvoUrgn1kR5oi5OXmiwZ6Uaw9ZVAIvEb7lYMPRFzIXIxA
/k5yTaEEmZbO1UxDrRzzO6Fas0p15n8Wrng0Yamk7kiNqOLUGPUyq4OFTARbkshG
u0xF+qhRvC/MM00IaRvOBkSspEWzgUEce3ccMlaaS3z5AMdkHjrNIUaM3K5VajI3
wu1Fkr7EDFExG9nQ42EQ7oHzd2JwBpYmrMgXwo68mBwdTfRWZA5A7bUclyTyU7m3
1554ODPneHuq+PT82TPYML2GnnNqxWVHJAIgx7Xauo7oibfnS5z9iQ7qH9Fw/83z
3IRWoNB87AEMWmvUP2jlIwQVYdWSDIQogd/gMyeBREB3NpZi5h1BRi9Tz8XN5RiC
0iBGSR4dbieGJ21tcC9357QsIyRWqpz5bPeqqxaY0LRi2RyRHICo+DVrZcgoTeNb
GaFunDXFnUttLvMCmDICylowAF1UGG46X4/cbC2XP144sS0o6zCX/loXgv4P3JMQ
8iTtDSzmrOssrBGWEupL/QvN1w7eYyPnKhrkuBrFfuHqCHDKxsgel1SmvK7EsUIu
HU8xe8BgdG86Kyem1l3PiI8W7SlKjng6yzGc2iJznh8e5o+naG0eIKJq2CSequl9
OipP+EtdyxxqDi2gk2Htew==
`protect END_PROTECTED
