`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6Za1O+VOS9HvHcCdo172uCn2t2yN9Z2IcBCUEe6AC6wAeO0CWKwKA8Gae9sBLS9s
yaPqa/C0wDES051qarp8XC/UJ5pd9fF3CXDRrYGq1n2Z9FtzVo2DBA5bHHHFet48
oza5rkJSahDmRjgbn5Y2tZVoAkj7F9oBVRZdhPkJVGT6EXVHwB4/E1t6M8c1qOSp
5HPjYwF3bDHm9ctoMLa+ayzauzafESSmfVcW6QXU3TWhYtXuCqufTo54gEkTChaJ
VnYS0dNkMUDvXPTEh0rJBM9pxuuVal7d3n8l1tDToUWX4g5lW65uiCkddtouz8lj
nOGuAOMklbPmuEtBziQDqA==
`protect END_PROTECTED
