`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xEf1mWyG4Pag6VShGjx5j+HOgQbUrytaCTZ2DcrZJeYz991X+psZ/kBqs+GtRG07
zzlOQTdVCqRTdjah/UJdNw160LKmj4VJUSP23yUKuwEYKRESp4W2ap2R9bnZjil9
+WqR9s9T7rf1qR98k4cFnLmkGzNlSfnpnFqmrSyPjoZzYIZf2cy0dbhLToScA1r1
XqT2dgYjYZyjD3HxFo9yPHlydyvDZlLI+LMGXhSQiN2ps4PPL15l8YuzJudlwkIw
4UIfqIJaXBeQy2z12Uwnvu137MX+rXjBZQaI7XVAvbOHiRxvck8Mdvw/Og6kDVtS
JFjdXyh403EqCCemtRrmvQZMCAEq9pI2cEcuR6+eFn415kP7dGOE4CMqBVs91O35
7kQV/17HMdZUJ1UQAOK4A+ReehsuQJt92rASO3VcXQjdpzf0MVtnyaOdX/wFxs3y
UFFcDyqpc/78/LuFtnDjLzkIs6sU21zWcnAn6vRgKvKpqtMGfcovjV0Vy5l7Bp10
oNYKYeECYf3JrdSZv5jwJGcERVL51voUleiZ0xF5sdXDi7w2cNSd6C+Wphxo1B0f
MjKg3Nzxm0idpiUiDiF3269XIcWO5hQJ0Sj1r+wxrwaWmNT0jVo6/HJX8JzpnBts
XzuxUzp4JKikLC/VfVeZpfuuRmmiBS92jBPVqYdVWMRxmNYy7ni/eldDT9ncWLFi
snBKG1PLRDvSkqAtmCTmDPwCXiutWpXoZ/oF+QXQmV0HSpbRH3AQqcJC39RqPM2v
wcD9sC5zmM1MgyrU9c0GbsvFEKyIDzujK7GjK8M81kSoxyJ9RGvl5mA2A6/aem3y
8nFHGHWQk/JjQwvoG4j3iEfqwPb691c17h1JmIfUwxxj2RSp2UQPrgzT7TbuPuYO
ghRK9MU4nCFfTWjMu33v9VjSqXkrJDPKdOFyJ9o1zqY8I4k3nYr3bn5CmMD5CL2a
3JHRLK1J1CIByvky8Ci9ubrx31SJ/7bj/58EMgl+GV6xNtXunGtmJ5JZYQnV6tRH
BZ9eCTJLlICyw97GYtR8VpsiBFbCk9JmqQGC+8SkR1oA/QI1P93Z8osKC5sQL3LS
UNPyWSzBDJ12qE9o/rPRonLzjzQ0iEKugiQG9l9D/sBDQAUZU+nf5+asvkYoQaxT
MHl0JPtvyd/tVFA/r0lgNiVaic9EbiARLXeXJT88S8VHk7beAtNM2GWhtizoblH6
8/jCTCu30c3skqj4KL+fDywPYl1uytneHFbBYqmm9Z+XIrdR9PSJM3/3cx1oDnhT
bz4RcUT3BU2A6kGnN9ptNGQasuEUXocZxDLqAHI1kD7g9hReICS+2YVOlxR80Ktv
2fFnjMG/3vUB3fDjIp24doUEufh1q9sgrEMBP2D24Inm/xNZRTmFo30qvioiwxbp
ITYjEcn8NCoHgRgNzIrabw/dF4eFdprkKL27q4Q+fvH9ia2QrZ2otZ0vMsyDIzZc
+PLhWTWDc4F3qvAQIQtNJHCX1NL4NLPp/DXVk6xNUy76FRhdP6rIH+1lU7SvBdnQ
yCviZKBQciaEeXA2e5kj497sxbqoSUoOfuRaWAXNLNw+MR33nBkZ2ypD+cR8fhFM
EBgKnCxRA+q240/fVQ1S408cnRaq+N5ptbetRcJpgMl/r7GbDIEUDD+m8dx6MxF6
R4qGhPUINzpZCNSudBipj07F9rfkTCIxklIejCXcMgZfK/gosabbtGpuxtubTZqf
0hkAIBEAbAVbFa7SHnHIGxpmzkv3i6ZtNKBhxNYO+t8Neg2o6Iv+GapnsmgmwQgs
K8B3v81oj+XNhCn9n1cZpNe2FREZNVqtLJNleT7pf8F+hmOWMHW/rSYNhl2gRi4d
y1eMEVfC0BuZtRjvTzKpvYvFGVVWmtCFsCGK8Qv/NhEYZG6u+FoEeD+PlivwhNuA
OBf4TRnJ9aEOOsotJWNGkJz52n3+EYYl3JTHwbNS3Ia3F5EbBvfc3duchX4hewBt
Cs/O2NTPy/Bp/RU2cqKn8t7vP9wlP/LQaanzOtOtws7aSXrjW0ED9YM8Xh+Ae7T1
g3adbBE7hxTyJ9AyB85KnJHjhyHPdTFeP7xSDu4oKkMwdIaXGVgagv1jYfM1M3bu
bAwe5/ewiJBcthJxHVyNSkl/8ogWd3eIGvhBk+YOVOFK3Xj5JO/+UL7/6tpfTbt6
inmLoqoo2OzrQw0nU872kmtyJ9pYdRUQNNgLnROCLdKfQqy6rrVO9sW08U/wIyL1
Kqy2VxcMMOmJINjRpoF7s4Mn0k8JLvU2+Da1E+Z+EKXg6Su7EhpD/FTSbht6X9Bl
A7QgNXVry3BWKsJ3IW+xNfQCfq+hujPmQmTS1oQ8tZRXpHTH+E4RczzgzX+3hrBd
NNvMeTkP5Df7YLqmN4PSaAXZ5WEIWqkPWmRYP5tFqE17ag8i69+CfIaTMCZDTu8h
as+/CNJLJZHcfD9YPqmXQm9+jpkNjvygBD7iXe/SWGfGFFPTu9KkKmaTm/OS1xv4
360ISL3kQV6Tj/TaQYZYQ3I1PSVPTqWiSbESeei/l0+B0lbShAd45JZLtm0c6JSP
EFc45HLU1cI6Xo4fSlq/AjwGUAqBoS87lNYc8rgrn5JZ9LNBN/6EaZoiLVSNTypG
D1jKhFkfZ2IfuEhteKKy6Ny7oZkJrpbMZ+zAu8vIIMWvGYe36XqFv7o8w7uwlnHt
0obE//cUj8yZsErOi1Via61IBNl/3oszXRYXQYt59RbnLqkE9e+DtTXAG9KsBu7a
6uIUNaWUYBsqhv4NOIGR6Wt8TPhCW6t4DISXBB8fOCl3x7GqkuXGs/OBEyc0Hydm
A6o3YqpgJx442jGznGeGartJMngHafmKn4ACy7p3DYHi9Hx9rSJeUh17maIDavMV
cE3N5yK7WoVtZ+8Fx9fyhGVmax+SSmD6Uq0F3QKJamxWw8ENZP3SGI4OIERADCo3
euWZXdZtJhJuET3N7r030Pa6lctvhvTxuFKexShvexInPSMZN2Qc6PHBfTakIZ5b
YX+lVYp5Df5DkqARLk5IFk9gFYvFUqYEY8qINqRzYlAGIuOp83ixpCtgJkv1roI7
WY930GyMgXc8ChVc4SmBxcmyGBhajcyifNxY9MXkC/YIqWuwzfwinrfIYT67giPi
ddCH7WveR8JAcdMVKGWg3EA1F+smzFf5SPI1x0rL0APvYvxlAEm7FA6Em2EvjNbg
2aXGuRn35qYc/VxJvkpyFQ/Jb8FWr4eUS2WyI99QsQrse1xZzl2QD7BF1cp9fpr+
twCYG5pE9TxZP27uq5yw3m0LELcBQJKEtds4WKnp4+80t3HItihijD02zV99cZVZ
dFfLQwi3yRHnNninCY5sheZzuKva5mWk56Ff1EE44WbV94CBDdKuFu9MGSgBJVf4
eayMXR0nKLUPguHs7MdFXMlRUD2e7HSUqHJvXk/q5SlaZYYj2Tn1SChARMc18lgz
WynyiRkKyHLw4w47pEMq7vGjKXi5jFrWbobsKPr6/BsIRQefwm8ZJMlBqhpdEq2k
D8UpiVDFhnV7tg9+7s004WaZwf7nZ9yh25wOcdyNOm1RQRdjyakUAue4/OSPixH5
sSroIbeKibfeCXHtOHt5JRPZdayklWpbaDQwt4jMReJk9udGm2NU+cXg/QyaXhD3
vmDVPN/yeUO7Kh4QQv+m+O30YlJQHD3BSW6SRno4tJXVbAFyZxb/C795Bc2QG6YY
LcEy/nSVmaKpL6CNwHgwebMiW4K/bUJ5JNQ9Kio1XvOJgHLte45Eyo26er/EaoO+
LGWkv3g/WEfxUZm10DN9EoZ4Zg1DfigOO0tFXu+Q4lp/peu7EMjgE1i44zm+sYo5
Mo+I/DUdjYAnDLGuRV/3PjO+IjvrMgqCKSBzScJIRFxE3lCXjJjMSK7hMG3gy7LO
ePJkJI+OEfyh/X8FC1gGXRbiXzDl74y+swv6o8nMKrcALozEb/3DQ8hEfuObmjcw
IlwMvZeVjiqDQNo2P/WxnSEawz4YxSGd0yfZTlCCOr7ACAUKyK+0EL6HY/EZD9dO
JqVdqSsdcuG75tfzdjObC56IPvlEoFudfPQpwjOFrNFTGU7H+LCev3NTqZ0Dn+SU
cELJFe7MNYmaMigKuEKVvEJEMCF4EkVsJNJJUCd8JxdJS4Q3uAHaR/0ayL+TVnvP
vefupXPUFwcDF1NRKGS/bx5wWTLzqUY8NfBwSySUsXlOeL9nqw1ETE2o+bowLskq
4SJWMgz/Sucuq7dvv2jZ5kam/8d+OuYZQ+YZs1hVfGpO712RnvQ3NZ6gzSTIzNHb
0pUxA/+ZAoPLsshY75gwli19la/sI9f0+BZxVnkLdV5n3NjKvY1Q5O3WbXX0+sTq
jYQU7gB5c1cCEE55iw1kqbu1nQy0z9fSijao+7+Y51FBu2K8jkwlxNSz+Hfm1+Zg
LTCZM4LOL+SrShapLQVZOZ3lY4V+9Nlvo4/0+aw9MAnkP8wGE856wO41VsFkUlrc
yqLfb3Tm2WKarYq0U17WFKQpbnc6xDMTqOGdRTJ1qtlXA6uqsicfANauad4lq3f5
Es1p7713UBaV4eSjos/EEWzxuiDFRra4imKKYfCtQaaMQOF80yO8kFOi0GLnzkr4
M/JR042Zrk0h4RHxTlOMqtMoPWfYpsRh5hoPNnzmA6ta+b5G8Fi2tS0Ur6SaflJ+
QuJG70snXZNxbpFpLbLW9Kqz2QDI7/i0VV8BNOOu65uCJSb/ETLWzk07QP1OX8L7
wjtwP73vZOJK1X+LpBRiJjofHfxHjWZpbVUCBvq/oCNbej4nEyB6FgYDECsH/Wf8
TTL+Z18T8Vt+B0kMaS8Cu+GblBPuESDTvmzka7CY/sAR7yX4hi0A9QIqijMD68qo
PmIMm59K7xilQFklNfvYNzzv1CZw6CHJzX158odv1lljKowil2n57HUN5Pa6mX5+
RBWtksO+R0FpnIcUmRH9e5rYBpcrzECg3UpqOhDPrs6yqLGjuD6+E9lY+khXYQQ4
bodA3amSe+uYtt78cec1rfjYoUoxe/nyawdTnyBJhdV//rKY2AZwb0M6bYYh2tbV
KhQAo4LD9yobtnX8A2xyn/YGbQalCHM3su1mDfXJqE45c2mVUR72/6jCdc/f7oVY
i3Eix1bv0sc6a/MUeFn3rcMk3KjtCITO+3F8yEjBan+BeN8PYLJ6+KMdUvy31g77
CvftIE0sYZSW3BG376B9m3fj27yMqH0bdpzw8YdXFpMLpVl/Zt1RqOWWmohPbjQb
NRETRSHvSUX22Gf6X/IpmYeBilKFpPby4nGyUZJQt7CA5tIaDcnhefYdsW508wT6
hLg8oGGhvgY3du3CKUnb7I1OlF2yA5fWR7RXjzCr1HzsmAIjv2ziJnH5Czz+IlKW
26F2FcQggAfqjdJZSxNc95ZFLbJvUiiYJqefgrucYGaqdnkjHkls6EsRCdmOJMLT
8eVnKt//EWVTaQ4Bq5Y/uNy9a9vc05vJVVJdyY7vwkirkbbHLF/DkfY0Qydg9xvJ
9nP/xSx5YzOF34kjPAb/gTd+O653siXITdMYPmHVOxOJcqULzxE6FT+M7ih9TgOn
lxnsW84llKc8xSIEDdpD+O3UkONGb7K30VhfYY7sXwF8MK+gAkoLqkww7p5POJbd
ZeZlXni9GG7ERGWREGY7IwGtroZuCSk51duFmi0aUcuiAK/VkVUee5D5W2FRAiwB
s/yE9yECc2TK+N1WOZQfD3q9BmgR3a1w9IZEVt9xXyyPcbPCfH1a83GI2kYzIkra
i3ZU/UrlXm9xlRyfo3hSX+rrcxx4bxCyhfgjVOeSQ6sp76+fVuMgKQBfOTvOUS25
F/7MzUbP3mKhzRJZaxyARXH47e3O/FOzNuXKrUu7sgRlI83ZjLr3bat/NIJbhqAr
0E78sivJh0RkEZtwwEj0caI5/y9H9NOpnlwvFZ8AgtgOXFvpgc98tUwnFidgFHIW
M36u+kTBcFoJvf7WywzjUECPjiLE7ALDw7y4eGnRLnwzEVFtmKbo1FIOSAhr29TY
RPlL+hd1+xeU29UByP9oOroOHE8A2A6JGvoHAINaPbq1Ab9nr5TRRZ142ztblSmF
3aIvh/29vWAV+tyoz9m27MgIpX1nWAItghmAYQm+iPun76JT12Ob1w+qengDKxrr
1jAoHHZg02x44pH2bPUQWNycMHMju9VE0/efP1RFD8JCUITclf0SlISEGu2knL6c
85oiVOhwr0p7UfKSis9X54Dlz4OJroRTvyZ0axpmMO7tnco5M/gjlHcNLj2Zj5n2
6mjQWR2Q7oeBO4NCNrueC5J3Wd45/K+khLQysXxZHZaiSnbzJzJtmRTwdn97uDBa
utXYNA+VrY89s433PZLZMkbabVDxzJ+hTe3CkfB54ftPrJRCkw8QyXD7CJl9FK05
+dmtV4K+Lpq32zFz3dT3IOc1ARLEmmGT/rMDZxjGh4dLyEDIR8dzhO4GlPj23yvY
ZRXB0m0ICGmkD+yDbqU15wUME0IVBAwsO79/KvqWLshovix43OoXW8TUKwADL5nZ
Pjjc9t9SL8Gd9SkoLHQt8nhCPn0b7ZUjD/WuOX60uWat7FywsPLI8U0hAOP1XEcd
QBV48z2x+L/FFTu8LV6ypQ14mNGUo54/gSNhHbccGJ9YYujMOv8ufUtpGImchwM6
L6G4WYm9oLH2ijloOs601FUMp8YEixqvgly5vJj70fJvdTPnm4WPizcuXiuc3x1Q
yMVvUGmZctkzgGZpaAHcTVe4g5MyonRkN9nEHp8WZ0e7JQS1VjuWrJWoBEt1tjyk
TOaFbnXnZVcuikj45w0/K2vwzfHdLC/AZwp5Pf6Nx5GW6f4EN6FsCw50N8dQiu0y
mg6HjoT4oyd1xj3aKWrmr3E8YyW60OBtKakbIbUh2oc=
`protect END_PROTECTED
