`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
u99A1h5ESeBTmg6OYoNrhsRiLkswUj9fYrDB5I2yMOTmovYiJWf7hJgNdFO6Jm21
Fut+vNdEzQw66D0HrPxF5D0JtviaOwGO0WVEbE2a458ZBTA7zhl1HFerl+X7wzZ2
gIc6xykozLLjevfBoLFxKwfl2ZTEAk36eDObQgrYa8gunAsrZl0mF3NszOj4wEty
ary+/LLdq7BC1XeDx0V2KaVX29vTH8zUYWXr+DIlaDbyn6NF2mTGZ5801Gk5ZSkH
Hyhc9+M+mmS00AjLfQuT9Eq/mCpDWEIPA27BvQBJpJzgx78B5pflIa5LzBZIRgqL
dCBcS6oJFZvHlpbPVP2b/QcCJrpHspN4J5aMDF7zNgMYeTpBeqfpKTLwOdq55MKl
FUJf38dqHg8aj5VavVlH+8xsDcDz9/L21cyHhgybGI6LZtb7ZBMzIkL7WrhoRTNl
VWBuPMihYLsT92McSIgQsZulT97fjFDg+nxcjp8DvQgIbuVPgK7xLmOnLCwMq/OI
BFKGMqlweLMknqhwWRL8pih9eNDQMaz1BQHITAy1kNWw3hIFbpwpvpGPlXsqiSWo
4MLgo8S2IH2rGujcj5bvPgsB7bzywxpc9AqG70eNRzQ+7uQHTH2wg6GgCF+HKvSd
Y19Gpb6Mt730VlLW9XTVL54G10UmYhIi0t/jtLH9DQmNFi2enADtllfUtozYrZ1c
e2nx6PjSzimRMa1yhnFqdmCnUmD6RSovWsJUGhksPIBQItJg7UtUWZITK80lcVFN
IbIpFI8ZkaLjupP6d9iKuiwchPETCDA2ge5eiFj+t8I=
`protect END_PROTECTED
