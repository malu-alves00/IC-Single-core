`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
azNgkx8L8fyuLvg5SOx1V3MtUFaVJr1FQnHR2f5WH5cBNgc5vVeDTsJePw/U9BA3
Ai9uL21LpEBOKWT8txEmR2/81MzO8eAIdk46U41Po/2vGFebZwiAs14Y5n117F5c
aYTc6h6sArpcYt7BzZzF5c77WOI9pzSgTioUpTeii2af2YbVPD7TuUkCK755sF81
W4W5Qw0fdwOycsdXVE5PgamAVTuNoiJXaeHz2miMLbfIs12E6yG/eDMKwF6vNgUW
C/sCV44F5MhBljs5n++LooVvQ1FSQbATQUG+lp2cRTenDeK2R2So1Y8qrdE3MufV
z0Rpg4mGhsLEDu9PtSJewX/ijtlIFHSng/hElNaTInbf4YKxkupzKDL5IBykb0v2
gQGpzQ+3KUvg7g1V66PMONtux+1JtXQQYFTLx2S7utjuKBian0jZvBoVKbVKlqEI
cKSWJ1aI3sqSW2Bh7rlL41bMcBnqcuZXg6p2hlnopyaqbWPQCkGA8BI+lvS7xmyW
NaaSnK2GwtjpvYLJ0eyJ0e/T/LSn0oDVgSWa6yFnoqHFeQh7sdyyq+kAhVpSVxz+
ljEKJvQG3KC3/E23wLyGUKi9BKJPfmvsNjiCdc7SYvmkZ7ophRuEW+Z+5cc8z3g8
/v+q1jkPs0NDQ5a+8KVqe/bvX7xOhwQemhwQxPFp+dsRGz2aRKFmEHvjp5Gw3thh
e8h1+R4kYNDSeumLH2+EVYnTZTCjJRLxI58x8TEiHOiho0hFs5DHBulD5DfZlQZy
+eN0Pme0FSCRqQmtYDGn054hRvSuadsLca6yDfAgMKHQFfp8TjBPskt0cSK55W5Y
gJ/rv1CiyHf2ioyT6Q11Q7Z+AWriGyi/A2e7BolZLL3ew9b5CCR7KKHbTPiGTQtZ
9CbqlKraTx3/a67QV8Gs2xrpYqWuOsFRB54FQRYsTyE=
`protect END_PROTECTED
