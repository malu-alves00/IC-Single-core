`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MXOVR7WosjSDftgj2kJs4puKA7Y2O6l/BpIzXmoqkDZ1N1oSS0h30/+Xf+edxjfl
TDwoRvVH2p1NZuJCeFioL/DrNlBa+6DcE+1mrYzaXCcsvAPo7RLcDGB3GmDeQi1H
UFEjVv1BYNpVhxh83YezDtBzLQmjb815Vhk818jQcOStLgs+I/9rmNzqZwthIZv2
zrai5rSSlJvKgzi5LQq85HHNNMWiSd2le/BHngiAAj0gJOB6aPsnbNIJUmodMYQ6
Xv9HXFQM9wW6jZxNCtLGNwo3iyY9eZvTpoSTyOzHGLXGTKlInRgqnDZLP15Q26lO
ah/trsQEr9I9/IbPTk0j6fpD8BCkb5ABrZQ4xaMtKFeS3xFmmAmuKJvYIUJxOPoN
LSnmu7G1ky/2iU9UsavUhLo6VFkJVOoTwEPRtG2tSKkVqw+z0utxYJKI/F2TDYCV
Tvh9+HKope7Dyp72Im1qo97zVQOzoQm2/UE2DWYmeTOPwZ1/M+3uxES42ZAPQGJ4
veffa8o3xGJ0KFmcEmfIlvmHTT1GR1URFDzqU6yQcxyJV6wb8AJPhI+qp4YEMgqg
F8OS7j6caDx5M5+KdndzWaLmM0dFYVHsERIpTFAUdIF4E3a1IgtmFd7e7rRFmJgY
Q/JQOO6yxmzihE9irA4xWP8JHQJ3RjeByFoPYOI+Bf1SH3lXMpoUJSbk4GFAFUqY
vDuoWI5kV80FPt67i9sVPO63mZPCIMycAdhxmcBySVmfvckbF6Ee/58k0Xg/Emxu
o8D7skmRKonigd/NMfuyi11qJ+Vq2MBY/FmdohLDD2JzQ3JAWNBsTqN9puFSvdak
wkFN5r1K9hV5Xc3+NX5q4QpIPx30tj5UyZk4L6b23AdR1AjF7QYQdmcNGH7bp+Qu
87h/5STZ2cL+SB1vOrXMpxXMmkQzezc9TBVqpArfpuNTJ3w0C4I+bW/wD+sKNZxi
uETtkEL8pD/b6+coSmNvlkQRq4TetiTIRCY4taOk7RxHpJUC0Ux4lVwoG+8KUte2
ppKlnTKn0jPAfqOx1mtbu6el/CQ6jO/abPMwNzZy749K7nQ1b5nk4kpGKi37VNeK
dqAH/VRgKA6uF9hqFlRGwQ3kMQRhLajStEu17TXQUQqjisM1xyuyD/O/vJNe+12h
goBmmiZThG+16mtKG4jWf2dsZAo0JKmhCnNHKhbPGD/+rg+nFqGCz9X5WK890d2C
p/k4ceeXJjs/HlnfsjIfyrsf3uis5E04hcq0sxnGhWcOzGz0soneUJTpa3M7OFBn
XF1mZRfGejiIw0p5WywsANhZK/8jh6Vl8nIEU214yRn/kfA8v44i72mlsncrS4jX
GvzyB8EI/mh4Q04P3ByD6JES9i1dRCfXFhTUbXGbjt7OjTJCvTqHjFRtlFaHwoST
pZy89zXsG8CeRBsji0F64osUxLTEOwnbwKeaa5ZFPWKDCihPOOEK1G144JMymmhF
JEfPXAyG1uUbE8+XyoNGjJB1gpIjE7fX+oE/s61E998ywggMxwXtiJ3sqwleIXX+
ITKmVGepWBKw99ch0sn35FpY0olhA/wEt/RJ07AFu2wiFVqiFmYjyh2gM7QSsfOi
eoSV7ya7ozS7qmkIykUB2l0th/r504z76cUJWZ2BXFUFpwvm3QACDGwDfbl0FSFk
r+VcEPtIZIbZf/vxZi2tD0X7AVBuS0Nky3Ng1UoZzzrG/ht6Sg+muMoeu/9hm9nd
JrI7bdPxAJcxRhhGYgfe5EMf04YdJFQoqlpjRmZHGnqHsM+KB6wp6gE/xO0yCmd3
LE8g62uZKeUAiGPyCbYsflHiOwb5GskklY/0J43Dw0xrzEnkTRL90kMtQCsWD6xB
A5wIj9Icfc9ZrZ7XmDElp/fyfX6LmKANWB9LND9q5HZIgU3ytkbfcBU5FLfSzuea
uKtOY0nxpQN/5GiLdCFJcv2mRY2nSl7OapbNJs60qf5OMESl/NwcNDdVSRHWv5Mj
HFanddtxreRRliKoR08mwZsvGHz5mIfSjJ/6iJ8a1pJD0nqlo8P6GS5ktaR4erJC
pAyvDwnf2Bt6POevYcQbhX1Yd2bbkJ2gOCADsPQrVIsCshdt8JURzvIsGaa6SUhs
2maceSPhCrV51yAd1urAy9O8gKe8iZSE1kRz/KKn7XR+n+YVvjwOuC3ckIowYRsK
RZe1JGbB6TcUJWen2p+3jAQWTH9/9DBPaQ0b1SPMAUCXzPGqX5IMCZJ2CWfw1bdI
TZOKpIEsruk6npnLu5RPDOlPfHHodyC9gN2yen7G9u/IstUJewGrjESHFAZDDVV9
548csoeI8NqyX3XGO4ZLxOR2ZvTK/fbKbh6zLatJex10TcdaN/mYmtjRoNz1jUcC
c2HHaVXAREhRUNn5eco3LOSvHPU06aDxeAWQz9AI/XbMZJ1oq51qAUJc6OxIt1pR
s3VIyprj9GshVz8eL3Seqa9M7BMyYKMVzv0oY8awimTP5XjG1oLcCt0Pf8/CO40q
IFwvFrXz9W7P4p21HN4oLTVLTruNEoqkJ/mBclql/SGBqVjg1PUCgxuRshKvmmFd
9QPiMcKbwSi0TN3RzQcXTNf/GLEMDAidnVgn01GrAPd9U1TeoaTX3FXUBAN4pmD+
NqxgTF7gIOP3SE5vtoBjh7B5laQvGQlZGKAKnL4/63awjNk+Yg9h46kSJPvLyhUR
zKMmeNbitR8Qexe96WMkYFe2MTzivLxDUzoqMtHxITMAWriY6PUdhaEoC59Fm2Vk
cUbuhu6AWrM/B3JZUoC+yOfl+Z/aT1acc/6idiwCIAhxFRt9qslH8tBFWYljMXwR
1gLuLdMREVYcCJlOKDjcg9RW/gmuqcwODVwd/4vFyzl6dbib8qax6Wn6MdBwD87d
rMqUnO5F937haGonjkowiHIAnXoNVufYlpugzl9YCJ67gSTDW91tmMdzX3uJAJQr
35RRKbPl4zu4A2g/rEtmxy+py15uP/8wEMHjRT1TdSZN5IgO7m646ZSM3lmL+ltJ
u1HVUZ16bSSZvu5cRVfR7rzagjzSvOZRwgZhe3MKDYnheaMtJe8TorfrrsAAw8XH
cuw5ebXG5cgZONK1r+VEcT12Llq3dOWrs5WoPAZvYyHSnMauQpStMOPf0/hcB73I
3NKfX66Ov1OlRW++MJXvWER6T8mtM0LzfEFVF6kBVjbYoWUB86kUzXtTBLweQdnb
wtItU7auHn987jmuRYahvQG9sc9XXFpTM0ef+RnP1/LEUi+wqf7nLyNWSY6yfJv3
dmXCWkAIWnegsiWrS258H8/TYuE6Pb/69V6/PG1MXtu7clUAjNnoatzkRn9xQein
zcvp+Gkq17Jd6QMetbYHleFiRbdP6EoqREDK0dRUXjcfQbaCOXlZL2kIwZYwNAtG
mzucT7TgIAiKaCtsTnCQnW0ESuRoyn4n4KOOyYeczPUp/MjvTp/fksryZ5VsOnfE
6/CAXRoptnQ1QKpNrI2hcaWof6XzOs9lBq1FaIahL0N/VL99zfkXe72KsFr34tq2
BRq9b5f8u5SduDkKtIXtutQDwPSEGAGQq8YzynYr6Wh4IpN+egHkvnLJg4LGsK5b
rf7exCK8yn3Gc3jYOWhGPmu/l+zEjGb0SRJ9xtzzWAmb89VnwQscS6Z7JhrNnl5t
diUzalnO259x1DCmRIh8rcaM0xCAgHC2vvX0O+teL5KHOe766gefqDLVbYuMW6g/
oR5Mb7rSPVdaUF2fbsqoUaMPQmMNggr2eAu1lFDH9MuBeNIRYc/+NUk6FeW3KdDE
PvPCa8UzwPWELCO2zKO2y61DT7CZ7gnJWBroiLYtkS4peb6olWzveJGun/zZOLcf
HOYZkWy6SpqMXVf1IXhEcNOpUmVENorIFVOeIKtb2UtGfcW5LeDeYvv+pJIJGE3U
/og44bKNdnts6Gb7opb/sOoFkzHOt5RS8kvoGgPKDSOp/Brrp0sSROxA9R4waV+F
1/HsaGyhVEHFsUY/9ndRcZEtmnOGorpQhgKVnjnyY3KPA8ry9gKeEusY5zB7Ru58
zJi9cZ6YOXuDfKELXmM2zgTZJ5eL/l427rniWPkch6fHQ4Vvb6/Oqy0xflILunEd
9yM/rBFEIxKf1ZfRlXSlCoDswCjkSHe6dAQg8+o2vvHjp1AFzaP0KEfK331nwv6/
rJ3XDoTRGCzURy7gn3Kh5L1+7P9A/z7qcPBhM3ZdfnAqVTV3oNsfbZbaP1WE/Cy+
QzOiSZmJ031t2p3NLJFznu/feq+14I1kDdDTA30opONKWqBjwVQwBPe3GIddptHw
68f4OpR/Cid0l16LPY6hDAjWF2A+mbn1mr6Ha703EGYIVz9hzOa87pXF2/IWW7nN
rlsul5bPuEra2AdaBfqZ9Q0BFVO4LMw8NeKeq17GWCywR+Dd3RU25vZp7xWzjIVj
BORfYFbZzMDrjiX2yv1Nf89khVpz1Je8vyieKBw3MvtHN+gHt26SLQGqO2qcMaGe
5Up2p7kdkFvx2BKNuTvuUn46gpnpm3LNLFK5FeBTLiArLiIgiNi7yMB2JuvKi9d9
Zxu7mZE35qNYiGfq9oHDcQ4uaNvkpcg8FqshSVn/hSevoJBBO6GOnrljLH3UsqCA
0Vta19kSN0zGUSVCJlogMq+nv/6sxLMDj8GTKdguFynkvbpL4So7KDYXoGbvkDrk
q7YEsMLA+YCSx9kT0KWBf4fpsgiIOKWMEe06XymAvC/Mp8fgFt3VPB74wxh6ia8d
EZm2wHsKf27Qo11TRKnBZSWNRseI+LfWvVT7GTWyUfxZTzco84KDE/1xHVCqrl94
XS6lIDcTE8kFDthfWqOAXqiPqeY3hNM4CWGxzKNuNmnS+AwdyGekqlt/GAOsIml/
5vGWp5d7a8MtJBOJdpdhhA8eWSZqQnQ8Py088OoVc1Htw2GK7xdY0/4u3dabF5a3
rC5wPcwK1N/g4ioPoafd9UhmucTDCpEGd20+zeYaVFmDEJWjwb+4wY93TTWpJhoB
5ZNrgfvrz12AGQ3MxcOndqS6mu2nJSpWyoL63PkaF+E65DDoPyLM2bSbLumO9Q+4
4zsuz94VKcgY2UaYOYxfXEAELPEs3FwTyGEMFwYOIf1ldXop1sVWVO3rYISExZIp
3n6Bm5SGNBjvwkGXrq2xpuO+lbL6zsTCKrWdgzZPGDtwmjdgjseEgWkeY7j/r9jd
d0l3GkrquLyUH8Bo0hE6khIGpDjPSaBauqUJlnZyQL9VDpOVH8q7i/D5JIbchibz
+mZf+H7ozsvxZywDwE1xSavSgm7BQ9GgcG+/KWvvfArtq2wm/wLNJ71VJUUozu+G
QEhjPCEC3Qg8eP41qPYiYY15EPAEKoQ8jgNpiSdocs8mZpGrOTVXt4DRn+Eml7n4
bqKIIfLN4PJM29Zloj89Cs+M57fGHfX2lBWT96FVASJ3mq4+Wb9byKCp8OmEdGLC
HJZBy5PYnRljb+/BC0YazBDcHw1shmYkpY8t76VSYrjoSjJDHKIRZ8zWSbGF8w24
hgXQXfsbBzP41lj7vrbFShFLkoC+KvgqovLdItKVKkiJlUXGN3toqOawo0OMiI1m
nDyZDCmo+qM/BTYKhWfaFAxiD476d9R4CaVYLTY7xHcuHfgSJsJUTrBhc+GtZ0q5
I3IhUP/CCWWKBqC7ZVWYbObMZ8BDw7z5OH6cEKZFpJBYi6FOSzWTnZheXgUIx8Ec
Ezsi5XJqq/oU/s/kQKWtQ8Tti7/qnF2bFzTTLvJcJydU5ZVegBTLdkb+HqM8TKeY
qiImlSrziP495xy39tCiHocwiagSem++eMzv41zFTtVzbcwr+pAV627EFop8l4V6
r0/tEa2d7oS7TQKwD0yUSYoSCCVrLCR1EUfAgeEwVOg9FebKSt++s590gqjiU7YM
sCzDvjzAiDiTXZ74EQoXSCzj1ktv6An5OkvXbbxyrEeV9EVBhOkoJQTXICcycenU
d/lFK//QvHoz47veUsVCwCxQtv+kKIDEk0r8QtObO+yVuKvRhR6QIakB9liwXSh2
38w+fE+Rpm+EKRclXPwq+pm3IlFEnFaWC8VIYqzzXNnfQJ2UTN0sUVL7pRBufGrL
Y9TzVP35NgftDE1myqBT6OOq/2tXCUIoUIsz8ZnCLOw6Onj8ZS3RHEaz5wvbj0IY
Q5W8+8wvc3Yoh4JXD/sy8SH5y3ejwn/c5/g4YbE3nH9cpd6nsoAQzVT6dLAWcksO
H3EOvP3ezfqfsveocDaqBjayjo3qgrtroRe4AHP/ibyy4uiT7+CyWs3QdFnTxwaD
Po5GnHVxRmr27DFKvftAw9aUgHDfFdMiWtucdFXFSZCMXtrrB+9unMOMBtX1CMMh
7tDSXD6SdoNJT+/+Ji3itSHgosB81ltyv+EKGn4puCttvmNvw6lCftlPGCnFGR1Q
bJNTo5Wpj+SdS7TdeVhJzkMquFUYzgfzZElOr13Txz6JY4BcWzWpkAXQm8R1uvoj
miItS/iMeTfotfA4NZeXZuVpiqQrhjaqtGgg1ASVb2xFjeuJJUURc8vaFAP84StY
LMZEeeERNW/j7cRLuFkciSHAJ89/EEH9JSSYZ9GWAlqYJbU8LzMaH8wu+f65hd5+
pmoLQuQ5fukMvgyNpe55XdXwrEf2yDpgMXB2gL3BHDRPgl4p3Aabil7rgkMeT2/B
aMRhm/CD7ldG0HwonVUthsMfzS6asUfrhhc5OEXGfML1MJZbvqW33GSDIGJ/03jC
1OR6YuI/lmTsEjwpionikNIgYgSjSLgCr37uxMZ2fotZ6OrpFrwGvETOdzaBVtGq
m6S9sr1eL35Qu6w/T2Fvt0wJhSx44c/X6IPDuEcs6J2e9evF6dBtvqnqd4dxn+t8
N1Ye8qBi09YpLXpe8r38WhrfKyuFyRqjVQLv/8QHyuUjcuqchPOiT7yvHipoLYAG
WlkNCQLK6NaS8IDbkNZ1/xg1fGbHYa0AUcuX1QRl+dEsYoXZ/ge5vY1nTOHl50HB
TR8qH9CQizmt4n6E+MuNZJPIRNaVSpQaQpkf+ITmyAIjJjgFJUSuvt/5n/ZTXELg
am2HjYdnrq0Xriqed8yAtaO7BIEb9EkC5YuWMN+KL+EnGLt/KW+8shP5wb3+coft
iJQ+xUXOJwpvhgtyN4ImBZ9GQCDCTnAbWbu3XohEHxvNpVQbXrNIyTZ5OE0l83g5
nBgjuGatBhwqNzYCZaWuGcdXkQzLdPRYiSQTQo/YMA13ds8OIpUe6pA0Agin1CYg
ds79rAGTBkzWcEXX2s0TatjJRvmprah6XAP7XZvm2weZShoj8oL7YdOCL/wMCbIV
+oxjvnB3kbycoEWQ8rwoEzzwM7oV4lSDL3+un+kHibhaRvzwOzI+jzIDdRxaigyq
Dzj6eySgd0mLkhVkFyVCUECFsQmc8EQJqMB7Td1BD+R0U4kYxjF9NkXn7x7xfSkI
Md8Wpu289ef8CRQBi4H5xkggTRJPH9b3eu3HcfTaAr/g0GzILkHfKTep7a+RUO27
e8OVPcN/MnVuj50fnYy+cZUzQ2je07qdbrBr7JzX2rJ4/F0gTMWPz5HD7A1XMxBz
j8a/xl95rYrY4dGGQnZ7yeK/O4ZnTX87umWhrP92qEuH7UOEjJV2LHpotIZhLOZV
3HetE4IKIFZabCQqh+bcVmNqQlAmRlZwWUGvol0yFO/D/uTRGl6U/6xue2C/LrIp
3y7CKmeOyC/Lsq7ADfrnxOoKpf82zWDCuRpX4HUFDmT8F1I1NZEduhA6KmhAosX0
GGaVGyoNM/8CXYjg9WudaVT/+Dy2OxSApYD+7Wgr04Y3Rx4fXVQraPcZWhsFYW4h
VExK6NETmigYBh+UnbeZs3jCyt+ml8ve3PpoMh6flLJQP1tEiinP5QSmfKBVNBlZ
WFitOO3crSxVALuHgTM+IVe/eJl7OCos6ET4WMtpGgUG72Lm+AWKV/CW4IuvOlpL
nnBAlQESTtoWiL7eTYy36g==
`protect END_PROTECTED
