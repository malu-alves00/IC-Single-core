`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dBuo0gKqx7cZRxG+T406RwYcdVDKQk76/g/M2CFbxXJWa5IMLL86x6Q3KWGSFK1E
TlRzFUXyTtefyzWRH9i/HOpVvhTvH9TcYHoC3vYhUNwTQ04NpUiEPukmvBNsI7JT
RdCTYNLbCvBNOwiU7EgV4n8mMnzuxX3BufHz+KBLzqHNwG6YVYSMINSB069lBl2Q
RIF7x05KDEgwVKuekb4ooXXIreKcZqFv3tqmMmF7RjW3YYM3gQmf7fy7OcimosSg
sjaoheOUGjuxlJhvw8Kpued5ACej/Dewz6qXyXEL2Oq9YWC/neSao9nUas17evDk
CNLrjacXDGbgic9zQg3y5bK2NkA+ADcGm2ZuZE+4TT8q+9VxX/I/5pcJAnBJbDby
hHorN7euJ+s7wqudC7we23QaL2NxbpkyfAcf8vrxmIhCWqVZTf8D15+I3cdlzw12
xLv6InYr4zEhaVn2esl5nQL4Fk7xjYS5c9rtMxcIv+RX47U1KuPAo/QC+zaDZyj0
lMUUQHaEjS+zBpnxEx2cXLX4uPhnw3J0NObxd7wwDFdOWc3eA5aIqcck4N/eomie
sXesBrAB6606LI2jwoBOYIc043GOGGxH7gKjTZFVJXDOcyNyiCEq1ZQPQhXAp0ot
SordLvLfiUUw7Lf3lPPtbtQJ0mieCwh0zDdyy6yl2ne2Ce9H/I3A+NnZgfh/crWt
5okQE6g46yZb6heuuEnxsMXGSg05AudzEET/AtxrvdqR45wp4MfUXFOCrEQ/cxgG
d6L4bGkerDxtfB8ZMNeGBwQXSnc+FOlbHWxeDfLHY5MmG1UN1x1iVfbxgwoXVND9
chbZCmbwMcK7fU2kZbfUD/r9b7Phxt8RXbusEhHhRPvmMIkxqp5WZqDCBuC+qbmG
VwHdaf8VbJUJdM87owQQBo6v2A3n54QT0QQxoSGyALK+rNvTaFOOAYUL4odvx11H
WxLMahpr9HlNC7qkcCtr5s3n2LESoT8kXvlBoXbepq/GRpEKFtmJYc/pknSYeofP
Mc84/LTpucTAb4UUoyHx9wB3cGEH+mmV8Qt9l1ZtsSemIKUpScHkk2DptuhF7+F4
iAU9ACLFrNv7cM4Lgywv0rfgIdgpcnVdv8vy3La3J60aR56klpYcFQWlRC5EgdNn
+YjMnwa1yiG+va/PkQnc5bpKzmegfXYD9BveNP/tUNtovdgamnmKZ7VWSoGFBg7B
xSgxcxBV3Pc90tvTjnK9UNgwoTziUahbf32pISV/vfNMUBXX9aWptBtQcicMyXaR
Rn16436ifQNqAwNWAOwViTC6or6pBKprpqo2AVlrwNeRouH1xXEVdEkf09ptvtF1
ce609MRZCjGEs2aXvd3p6VbqCRHZo7wdWAl+UtY4KeFqD66nMz7y1VsKAC+562++
faKpzkxJb2madtFPl+qoJhKNtAOR45VajD4Qbj9sv4Ia/2UrxjgiOlO9nl7n3duo
n8CRDrCFVu6UM/oAEjb6K5vlZUk/wenETWF3XTbFZAXa62pTjSmBXf5F7pQPEaYR
+4WKifTR9BXtil6bGsAuHiJSUDTBLhqOv03kVUS908kOOOPkFe4nV6/VRy+MEmAb
1O11ppHuhDJUiFyoysmaUNET1qiepiFs/I9f8W0amnkWYtpKBmZ182P65VVxYUOt
3swd+DmdT3hntKXjgA0cmVU0nIfIUx2CXs4j0H5p4FRJIfJQbctl5v6TM2LHk1zg
oAwpYTLFzvvvyO6T/8nsurtDaQQog15TrpId203MEPvG84xYVhZMI+wxw17wii3m
rJ4spKFH6j2Go5jdRQaQBzrv1MXnKL/e1bBpnXiU2+C0aFHgYNHa9GBhHk++sAq1
zBChKq0F10b07QLhiJZbE+tVt9bzBFTCEw5ySs6Diif8bWxg0jJ85s4qd0kWS3W5
bRVddEzla8WAMyvV5c8QhWmr26OTOdq4QgH/hILC8BPRRKujYtoHGuvk0UFvoxz8
EAmSde+5V1rAJWm/+uKLkf8qAOiC/MAUloIlzfyVPN4zWJmkkF5uaOg+ZiXtpuyk
lTRJdFeCOzDgZVVtHS7C3lsLvJFh1Kg4OoMIGgpETVlzIWDHE+hW70mBWCqDH7Qq
V+D9KSAo9zZLiNjV6yxoqavkU3T+izmFb3I9R9Q7RyGbtRptvXb9xApOF9SCheAi
6gzakf/PEVnW3TGWelueG1WjXhZJtPFwNp3pQbTft4fZtGyVf6Tpg1dFWD8hH7t+
/fdZhH6RqrIGlf467hfq9hFe4BE3Ielj3lB2BqonGPtXADZGw5Pd3VWI4YdOUa8r
GLoIpOcQPtLr0F7KZlhz6/YXr2eM0V56V9vjinGNETzS89tEhr8fuSrCNt3CxZak
P9gUrh6CeJa0yaPvIdcE+OHagZQwXdlp2kM7OBxff9klYfoBWpXVJJQI4q1Ox53P
/t/9J7NJxGap7gSWiGMsjyJ/rvlJQYBf6ZNqBxvecvBP+MWQk/X2jh4yT7DLlQ8o
D5ZGW+5z/+WtGGM4zpHsX3tkMpt5GaU9g1bXmF2ADp4iqC/FhzR2tJVwgpJAQ1co
mBq6ABNW90NDWpIzYULEGeWg0MEC67Z1HlwLs+CBrqk24xz3Vb3m8DpcIFSCgjo1
CzC5vSjB4Twfv7uFicbWgQIeAvPq+i8QtahpnvS6CWAbuzW2SiNt77hI49EIXjLS
gl+7Cch1hV5AmxJg0Iuh5IM86nrQeWyOTWrwBx65HuV+vf3hGhClrDKLaMMtBkoV
3adCFrH6O9A3LdmHt9dRe7kjfSYIC2mfYMktm8AGl91EzqmgGiHcdthsXyHAdz0V
FXhQMIUCvDCMbQdmO+40s4HK7mssnQiOYvCftJyhwUnCqZfJzum+pcJQ4pjNSV+O
/TVqWzjeet+1lst1mB2xLv/Sx79SPWbErBGNaZOB5bJvbIr+T6z70+08x/mp+mdB
tdPWR1zbARHmsuyZ5nDjq3Jd9VqD4HuTMM9rWSV+2uQBm+pmpWn9NzVcoxYS0rba
tO3ncjq4LYQ+Eg0d07cPqEqEmwWj2BZ1ABvwPekQwcsASEVaGqoyHcQlzxlu0UXM
Rc7gvL1dLA9ggE2XF9slQWN72wnFxTEARthAQoZfimST5YZCTKFHHMh7MKcqZHzl
13urNrqV5IpSGfmkBNgiwgp/5gUqHMe9qPOlZNnbtes85auJh2sX1az8XADlQUU7
MkfOdtfknVu7l0gwITCcNXRf6FD6QH3wktEgJCcYw31rffWtvdup6p4S2S5FI+Q5
grf1mceIB7Xs5X/fGzehOpRLFRoiVuxaR+gyrpwgrqR/uxRp3NoToQh6f0JNOsi1
RDQK8pBTDvlCOP/uftxIQj92D5l7YuhwcemsVkVgwzfJ8N1yrm5ZQeWfM4b9bqt6
MpPODCzE8o8lICktIGsVSNLxTHBtsKmtWjSpnn01z9n9YJ++svS81aeJH80tougW
ZnNP3gN3yUyy4AAXe/wTfJ/U55eVnzXRZOpNIJqukgKXa9sHSQD6wz8jxHE2m8iE
DEBfFOrabV2+1G6qqj4sJiAMlxLDqWStreS4KU4Cz9w61gGwflDIKmzbu8m7fnBV
vOnxo2+zxqYLUokujpee0tTPUz9yEfHbBsEg+F4xwgJIG7sma2bHnN9a46ZGIERv
VQor7UXEfTC/Zt6HP30pzQwA8Ime6CyS93tCOf9VWGQkgTbgbiSvBSRodbVq2kaT
WnU9v30jISEN1yIM45NH1/ZrxnRxf6fpzz6G3R6ovgIfy7CsqJgDEGa9fQdlOH5X
cwC9K1RlgNXgVgLNU7d1fF2vi6QKVDheWJvQbUzg3IiC8VwyNYWcHKIDesU5d4aK
VCI0XFqnQWH0UgbESIyvUwhHR6kEmwdzD3GJqGN8qcSnGct2PvX9RThnsHUkMow7
spwS474+B+UZ5YIGUTO2yGK3aB+qV0rXbiW6XmB2zXekgBu/eoN6bUV+dun2LXXL
XivH1RMTF9ebVnGqpPPorGMawodxhHfah9ZoJDW1Ga0Ri+ZAI46iWps9KwIIIogR
HfpAaheEReqacKphivSlnxFp4YRJDkCYSfYjQ8RgrEIs6/iSaIldeT5yH5dk3CWJ
LruO+9rP/bIiMOc588KF/PFmg2zuVIzjasTXCqhYrckiak6OQe9wj+iUbtkdNrpI
AxhkV8LSjjat+4MeTdCJqMQ+HXKqgahAdYXaxZwuKwPq0C5eclqrtFHh83wzPImp
bFeKP762RQ9BXOmE0/6Y8aqxFk83/ilfRaeaAK1QI83vwZHKj2bpW7rvkzA1Q+5/
bGbe0TsNE2sg23wOjiLYTmM0CRM/4DFELysTDYMd/UJk4iEvEfLXwgrZ4nC4XbzJ
2iEAjCqVuc0bhhn3RZnYXVJtSUHbawgsRi7mFPt4Vn3RqdJ+gw2eVdji5BT5t0Ao
90cIn/wEUF0noPeJfsVeFJQ1bcouQKi/3alPjLn3eGw=
`protect END_PROTECTED
