`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5XPNJLVTYiUo//D7ucIGugFApenj7/FxAHCxboqVyQzvirdwd8kb0nSIiGXuUOYJ
yuHHd7e50tIn3wJTXtSAoRXXPuxBePfEpk24RoHqgl6cf5P4Mpj3Ka+LePtGYb6+
N9/vlJ0fW0ohjmezwajLIBbdqkAhwN7UvRw6kyeee+1LKtc47/HShnf5mzwnYHjQ
dRmniBghmGs1A+ATbmKix+dKTi3nYCNL5vZQN+dybv3qAq5Km6DkJzq+Ypa/Afoz
5Y7bfOdHEWdVO3sj2cJN1hpB8TzwgH9iD3fLbZ787TSqv0sJvJpnl1u5uNTeeviS
XPzhIUhoD8yYzGg1LIlWr/fjbVCu8D14VMzWKQQib1u2Jevbs5j+HGfDWpEvfB6Z
P06QWYrl25D5ojOUmfr3PlBCtjiYzpAnGfpGKeLXIlM14fIquQ7U9YKnE7wAoPHg
sDHa//CWP4xMwmB35MKxvakSEJyU/04MbxBPrRTXM/mrhgtpQL6IJXThKVu8nLJI
wS0xA1OL0cvLJp6n7X0VCI8Vg0rftGCzCo++FLZ5Ak4H2iourSk00VNXZALIjQlh
O3icgC/BuQO1VOWP8fYgQgfxDLveJqWobk4Qfyu7R7itawGDwd1eSsQBCFga2cVW
F61ebDiCmxGvhMbZDO07UBfQhPjZdCvZwf1z9Zq6bJOXdbqcJyjxSQm84fpIVGn6
FSGLw4D7yM/BZlOxW/U30V+1Ov0hj9NOq5/XPze/8aMnMK9hxx59fLmmtC9SEgN7
WctdSvquVeD2KYu76YVgOEqcJmNZ0j2QsmXWUtiuu6/j6qMlM79+nGj4tzkLL6K0
kMCcZnLVv5zmDNVeTuXgqhmCp1e9DnEYT4P/AW8IPO7AkQDGpKLF+Og+Z5xXqJ0U
OmkJGn1+2aYiDVMAf+AnXlZNuD7kKQpCawel6q1b2yvrhbBQwAK/DcmGpVCWIgo3
AI50QbmL58SAFhpKyX92r3xbGEUG9yHtAuEl0ClmYALrfVxm2dfYNibvnetl/HZo
e9W0d3wPzmbVMfNgjjFcy2zLq8vu1CVa+fJceMsFuo8E+gRG+gwuqaYfNcD04CSk
jscb7FCYjScaeYpUoNMRJVlcRMR8w/W3kideSRZwzSg=
`protect END_PROTECTED
