`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8D5GwOPlsZpbXZXtNAHZGfrXzue2C/h4xMh0t40s1q7qTenuvB6rermP5/ZC8SNo
vSBGJqrycabSEYWLoPJODU+Tnda3duAWOULjfABcsKMLZnKWUu0u5PHvdHypBQC7
23T3EgJIhEj1X8ws2j1pASvHlK9dTp2RjL8CsScxyOGX7sl/pOSTl/rQguTUL85E
BcLRfZXfnDdpwwrfYwDSE+5Hgw9p3QNzk0UsHPTK2nfOGZc6D2O8VSYYESoAei6/
0dUvDReyarwAxFpZ5tJbAR1gakoAQBS0aUdVGaHS4LLvQ1t8bodzSG2tLQMfxZkC
sV7Ix+ayIeXKNGnjchLKeXmCnyEwGOCGq7Of3ISGKPK82/psCxELpAiS9NFpKz/J
76NIcR8E4TwoVHfPmz6MJ+QNoXyLoTbAe+6v3QbNiGr69Xhl/yFePk38G+3cOMiH
CWN8mxlMuON6xi7DPZw1ogFt9dNnqKClx4j53w3c5kz1Qy9FU3wKmSudI4IzEvgu
vIo6g6Pn/WnW8mKD0SrMPiFdzN5DQ/8fbiNam6wEECqOdinmUPA/nYU9pNzCtO5+
WJANTPdxwgB9xRj4kw3WH+zQddrqFrT9JPN6kjBolAQcm1QZWzjaLEclbMPTkxeU
H/bQSqL7pHs2OalmdS3AJQnalM4ncCKzzooAbmvG6hacnvgsMTdD6Y76o6K1BA1S
URS1LeyJDFxLi4a8jamtiYci/11NB+ody/LH9v8JGkatt8Q+7DDUSaAvrs7llwuz
f6ut7HM/XqfLq/5iFtP+Nx03XqPuUnL9HM+/CNNKBNG+O2xIG9MP1Hq+2i4VqteE
M3rWzCg4hUl/GkIeNF48Y+L9qNcWWTrmDZKPw0KG2SjtmimFLs93vwhx9AZcdGZi
+Uyr5IkV/b+0g1rJBihXvwcVba5LO+9W3zOBShGKSSSir8DODoynHad2I61vYQtG
v0LTe9XDaY6pQkzKqYxnRHfH8lvugpQKR5QCjBwrlHrVla3nrZZrJmvYknBhWOtN
GFJViGmgB8Mtj6nCMmreh8bDxRkv6O74TuZ1ZMO9yM25oPUwigwbMoDEO/nzvKcu
/01Ja+mHXPUOUp2urA5uxPHUTRdMhQSsgVvQg+ZjA7VgFOBntdYHxD+v+XuIOnWH
KUERQzohWkIzY3YwpWIlIFuE12lxKjbqxHddN9PsSBnweteNKZTipdnr+OBVEae7
1hCTQFkx0RN0gVWkMg9TCgkXsWuOz1haSnD4irQp8ZLEOg/Mr/FyQy36Ptzc3K0+
8zfjR1raUww0kTwh9nOVxZnVMUeJq0sZNXkGsy38hzoxMU+dbmmc+/0/mpx8rEom
c2iF3Ef6iHfJYLdGULa7T6EBMQaEt5HBiSNjbnaqRnMOFVpzpZwQ6151eu0cf7Nx
ddHQakqZ/2lcRbFT9kDpJrZqBb8bGjpEvYNjP4WLzPia5LrTpE36wsFgNKVRPO4o
oMBQhoaBmaQbmwKz5JQiF7aMMt520MuFFHYWk/LkbgR0uF+q5ulIapg5zVohpQm4
EQo+0sK7H65BHEscdUYDI3CbcbA3QSPwKBrSmJQfWNqMxPGhUWZDIub9aX23tJu9
z9lxbxWi2U/vm5RriS3M6yzRXlbDOUXlo1KNHMYWKNwq7Sbmv8nj1+xcsh5wr0bn
XKwsxj3LOFBBW3gxUDbgQdDGAYmfJcNCgBpr7EPrJx9klZ2k+/QcRwBmQ5HvCykG
TMW31f8H/KBSVmFTewl6cEf09UtoRTmFxX1MWL7GBdly6QdlKhhOKUcqeZYCxL7q
XaemHlXI1vVpkXjj5vEbQgnuZ3eQHDwJc7j8gjcS1W+F709EKT+mjqY44ZP1SLrf
mafdMCHQxXDOkR7FOLfplBqcPDk/iO8l7ugq6J2OAh9h7wt744Ep/UwT5ssZf82V
qHVenu3VoFgJmvEv583nAHaZlHaurA1+benmypaIvQlyN2c/X8iMzhxNU8ka3nkg
dDd8ViKaZ4iac8K7l0wOTC1fEfcGUFOntRlJgiWhb/QtYeOygNi1QpOvBX6EYweJ
vOK09Sl8vOsBomnpL6Wb+MIB40Fq6cX9Wk89/0SZXgDZDADMOD6JcQfhDnHUanK0
JScHb4uY6gNNq1VTaD4mQq6zZ7LMenx0SFX4p9hYO8FnhwuK3sapxLLV4yhkSrMw
3dKkGNHnjwSAuZACRS2Z227CJU+L8rHx2o000WCCh5bme9oSwIKnX6m06kgjdbs4
IL52HcghNRJpCvrY1tKqlMaCHPmmiZDO+eH7wmNmutnF8XIXBXrsd5CiqTkAnRWb
EeMdsNUtET9oHQXWbKF6ChR5H4aUYzNz99CQRVgMlN0v6ttAGdvf83vGDKfRggbj
pjtFnXOH5GBFTqYs3SulMKWYo5RxKNvsrWoc5QxbVFanaHMFKeW5+alfdN83VEK/
AFrNMzdepAacIakp6w4HUmHav4Nv1zHDOhozfZ+CAtuATNhDAbVkuxzrjRT63EiW
WOnZy8xI961/PImBBL2OIkUFI91iAyKyFPg4GaiqCy3W/+fYQ0+8sSo13xtanVV0
ofmOKrJDMxN85FPBYwTUiurcI4wudGWGR6Drm2mtJ9+yxBHu+Y+iTNeE1zi+gyns
7yo9RaUt7RDFek0njw0b1wE7RurpNBi8hC9lmjW7s/3hr+Pe9fQejj18HHVtV2YM
I41VsLSeTXCeopXSXBOak2plHzCPEzBttOubW/emvktqztU5MrfM7wqP2bb3l8Oo
nF2QpdJv+9ZzJCf40ZqLBSfZsJwZeZa8xEgYK2GR1Ot9p8xJSaLU7UyRIHNPg9LN
39d38Rj6CeBhWY69vYjgWvgCWmOQS9/4pz6G68p0qiE0M+krmJnYifzTPMewYZwN
sTOh6ZT2a5r6wPqOhnmgkeH1YtMPhE5JQMEwy+iTSpJOtHqhNAr7yJ7wPmZ16uxp
j9IFb1MV87xvkOkeGpgTvRv8smoSy1WB6a4d4jg0UweZ7KNIOd4r2qqpwtpGDxsx
Lk/hey/TIotrdQj2sGbe1hdEOAPDWC30qtSgWIhX9++FHB1xLg1m/XZHtV+vOrq2
S/ypdiltib8IZwiziBjZp73uQ8BztdONZzMgkVpc7mBR2vcIu8LFxovHmYPdRyho
/LqEE8iMo0DQiTWLpXhoD+Sec3R1tnVXmrY3mqY73MC3G7apsiQz/fXugBG7UJDo
fOK0joXkCWDhnqD7F3V85njRx0jk7qYVpLbP/sLnxYQAzIFtdLOpqdWuFcbA9FQF
XQs3D8EN14wJ7lmfezFRYClkREIOP1Z4XFhNniIf3+CXp2BRl9KGONuQB2elwtQB
RC48rDIeGw3kzyPofSNMWHxWhQLH01u3V32HT3X05uioCD+z4+rR0LDJmjiPOVnZ
nL6bcbpc7QSiqMX58oUHbaxhh6MWgp55qGYerBv8KKqo30Lcux4i7X0VurUJGCrV
Kw/U8HLLN/Zc2p8rTAv+rKylIgdS83uJcsN9AFxAWYDUPgg015lcw8Cwgr6iwPII
IG1bZ+uum6MgQIU9KyAtyBK+x01sdzbFcyJhivC1/HeDFuiAeTcyQAVMiBa+K7HW
Xv+VsgX9MyTuS/vTrTBjZU1aiTqxjPAI4aHpN9ThNAUHuEzCMlgwcl3dIktuTxog
VCO0RSHExbj3bvh+2/7N0QAmooNfyOQfIw1/AIANii/tUo53zp1F6kAjwbY/2rvJ
JEuf/v+xswoR4ywSvmgVG2BlAgA37LsgUdmLKLuHvI4haTdXEanL2SDGX8NlQvVw
6g/cX9nTRM2p9itTLtXRHZv7TsDbnajkDr7jhEl6E5kCDEHY/j/+jXUMwHkdsvb9
aa8Gw7nFX3kM7Kdon2ygrLhRPqOmKFm6aF/frnhV4rXvIM4XCp+UbxaefFXz4LKR
+wuz3MhX5iIaqo0GGLYzYtMDDJKMTcGmeEBZqsloHJyQiHVe6bqAdN7C4oSaDb7e
FrhcMmDWfdy9UlHvMnvP5lFHc8wsA4VB0Tg+W4kO6wo=
`protect END_PROTECTED
