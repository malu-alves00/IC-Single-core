`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6bGyFgXWdj+8lMrcbUH9MlpzRFmq/NYbOkVNZQfM8KF3h9Xl/XksqWYlJl7wh5wL
A1Muz5QxlZu+ZC2RiLQMFgie7Fa7B/ECYpsb34qMhA82opUPGfEAq9gufYaxkRPb
QoCfxQqB0cM26cLtWbub3IUbAnJPtAFcyNgLx5FwnReQktv+fAoVdxHZR1TAds3n
lLvnVjcPncEt9MGicYrIkg==
`protect END_PROTECTED
