`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hq+63d7y2vX5ymOjj45kVoW6po4rwhDTRCY5cWkSRL+YKWks0ndtdvydx7D38tHJ
z9PuTq87rwQPCbmrcx835QQ5q+DwCOUHPz+QLpimjCW2arejrJ1pykt1aDoD45ZY
OUs07MmjtkSp3upgU+mO/yRzLEhtOIhLcmSELw9Grr/jY9nURmOfCZ4ecXEr6MLi
aN8aJ52nMq7vMmBdnf1O+YvcNuJcWarorX61csp8yNYb9dEDGutC7RidWgCZRmvg
iFxLdDp7P4sv4mHH3OQkjtZ3A7ricuVedQiSJ1zAafVvlvcILOS6NVl8XFfSK3Dr
jfSMWvMh51n5+4PM8m8gXDL7b2Q2UyNrKPpUDgeeEXu7ugyIKTmcTOfyLA45wFAJ
pigN3AtMox3/tGCxcYa641xcv3bQSnUpLP7UK0xiYsZdTfNk/fTpsfd2CgZMR+fe
x0z9I230BKU4AvA1V5i+rpWYoMv5OhR8QkmCzWQcw2P/TaJObW2tHrsmWI6YUr5D
56fYrs3s6Edx9j+Uxc5840FkpaudHULVFr/iYieuocFho8bePz1GtT44cOYn1sHM
V0LnABWP6SDkFDxvJlNl2eABie4GBwqWdMwhMhOhFWGS818Nd2fbB4OIHW2Jx1g5
U/DLhvhrA6zd6jfDw2TYaWkuvBOI+2StRdvrLfTeI3OVHUtLqXZI1eLh8sKDMHAd
HzJy1kuB9pv1mzXz3V8cq8tNDhvzb24g4IEenUilX7EVIPWn15KadiFT6t+mlcgL
pN2HOU2feXLwdQEpMCkmtTye4vdsyVNIxD7B7YjacWeViTNGP61UIA4kmroe/eiy
mmviRSzO85v23m0TL0VNFg==
`protect END_PROTECTED
