`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nqLktNVJhYY0xLMIe8IWwxMCgbX90i8Q7HMvpBnA13KUFrar3T8GbV6mL3LQ36rX
NsRdOBn8cVNmVWnGSTYZHpahVgH1kGkYVTylfCoIwn0QLZUaJSFz6RFXdTHyvYuy
kgFaqGhZSBsn29+Tl+zSkWldZJL2BXynTL4opC4CmeyZBGWBmvLL9o7/mYzM3ss2
TtusIBIVxFat2vCLZk4zC1LnJPpfg2x9iXIWfjQiPdg/wxAZbVSJip5WoBIK7lql
h/XhCYk8qRMNJ3tEVOwSiuYJ22GjXscWPxexLCpqGzQ+6Hz360ZrzzSmAtsC8OFX
KzzPcwdogPc+sQDYd+F0uQ66v2xA00FisP8+VmzFjrHmyir5pIOKrIrvI6uZ9YGv
liVhb+LE3HEuecDhnur4VnTrs+vo+7PAcJTG3stSARQsYBDhAmp+MAHQPx1n2HKn
ksbPv6cvfsiLLdaY/yIr7dbFtA7IWE1bpFvqxK7UGuE9ewK8HV/rCd+9XWBeANKY
349GxOSeWwIPHDPk2aTXJ00NgPAh7aaZzGMPD5IgSV9qbeJZWjjMNipO2E3PIqJO
2AXysTADZIL0jq6OFCSkchEm+7Fyhd/qn+unmer558KiWFQYBTht9oFSs4DstJd7
cbHvUaX+TmvIYZ/OmupjtWz1bi3odpbAxAVWeuaHJPdbqCAXqRKEGg+CM+u/meKj
XUYDsDP3+bWJ6x8ZUcRtiH+iwRGf8l+Fsf9aaItTl1bA+nD7KHQ4zlvgC0pLWbQ9
wk2nWjVvQ5AJKi8GYQMMfD67hR0VHurlzoA9l0w16nN2Oy056SKK5OQdcgOUnOPI
Xg3JtWbY/tzTktlZLalH6drmbgkYe7YCknMBhpeHMyssaiWWZMDRyldsIW1Rw9Ak
VAC/0CXq162/Om35qcPiN+ONNV8S0/LJA3avTCvyA5vmZlpZqz0Ejo9xcnxEN0Wt
4SLS7uppe0ibdEvB9ynVrhE0fSK1a4kuyFwN0PP967zXFhkf7SuGd/UK3frZy2fT
p8FZekTE5CDu6NGuuNZ+YAsXihPv19wymzEYt5EVVdXcg02ZQ2pexB7xuYeWg8uc
yfko6U1swNRim9kRVVBII4B5EQf4o83X5xe50iXRL0dzrLmIGbACR3gDfFBXV73A
FSQhaRRo6LYoc043Ev5VI+248Hp6qzwkrZ7cxkovDYo2Q9xNf3dd8+GkcU7hl8XO
cTW66gMIe5U30VCLQK03SjcZeboVwEL5lHV0j+ERL1ciMjs4Zr4Z64lNano9ArjV
lhWnmbk8XLs89W+uG0hWhKgnz7t+UXbRElx/W3oQc/04hjziOAsed3wG0TYGbL+c
U+6q76/Khy3gFR6PgPbHGyNikO9LSqN0PYM7LWwtNm6EKEODUZ8xGTwfG/f8vRlL
i9yymB/yd94gUdp20sEEJ7hAGDtHWsYmqrjmtNPhPeBC5t2zmeGcbJKjApzluH9t
JLNzWLG47T/1Wekfamq0KuyZQ594gliYEEpdtbhw7biQHK7NEBAQwFA+SaO3POCE
3zFYuvHg41c63U9R81kJ/jSgVsG1rw4QAVMXn53cv2id8qIuEwcr0IOvGTE96gff
Odc4Mh+FXeKl9ZnNVXmZzXRHukyrS5av6wUqclC86C97YPy1YG+tuhm0FKHe1v2X
g0B3F4QME+zdk9EkbsxwsDXwNW79SrysRnWWzC35TRQKWeJQRv4T+YxYS7g+XgHK
uHilbN9Z7WJ6skxUxofEIuFm8Wu0XdFUkSElNYXJ6dXH8cpiuiwHdDdKSel394OD
NhjJk2STKg1I/8VXoFUwhBlxR2CpyL2XJ3pPAHeuCVS6QgO4Ud4JbBJn2Ftz/Rbt
PT6Kw6rnefval5lZ8RiC3N2HuWY8IGa1qGFj9f65bhGR0G+tHMfk3tLczX5LZpqD
FSFPKDKNV0t1KQVssMIw1vBSyR/UJIK8d3w+VC3bafyDHHckqRQw2KdHy8PoxTux
Osui0hx+D9WKDJDZuH1NCPc1Km97IKoRF7d++/0HwwL61/Kiem+geiNo/H3p9yqV
HqAZ0pB1I6a9gDZTtB7CiCc5SQayfoTey2lgYf91QIwMXH9ck6pG3AYKjBCqbKfN
B7P50VJU/fKvcIIn3CgF13Y7HNizSQyj3MbhLdBhttwjvuI5NInqfeX0HpviTTLp
yTAk3CZMFx/d3b0zflmQtcUefwz0eSLTcbC3iAPCI5TldYjBVPregYKCkqwnBWu4
Ab1i372k9o4/mm0/F78R4xAi/ft0+/S5/Dp9kHv6xUNKisVT+BHtwOCHb4kNhP5F
NEB8+x1FliY7LGtCA1MH0Dn+Vg7SVVLCzWQsyMi6g1v3aHJI7hAOC6f6HL5fgQzZ
+M+WIfxdH5gFomHr4DLejrVAMa3g4SDJN6xplpxci//5DHG4mO72xX4AHdNqowMG
nRXzHZFKPE5Ru+n0U2MkJt44XvIWBFH+/UMQpPRrLgv0mXfI/TIGFTA0v0ev1nSX
FJ0Sv28czZpad8laB0g2iqqMJqIFTgm46tN9phxGnv0pp00uZyfGlJ3xyju+tx+L
VEIQl0AgQr+o3XM9elc0oWILGED78ebAc8NDtKf7hEK4V3yHZhrrhshV448zbYTn
uE73qpzt417XzuDRbLvb8Ekj95BcNaHF9HeXWZQN8oiLQfWG4QAEmHHpeQngM8ya
AYpn8cO3vHhyX6j+pf238dGkV9PgKPxp7GPNNmuIBzNRaqECcyzgvP2lV6+NO3+m
7+u2fmU1ZhGKhHOAzx51SaIL5fau3fsWcbR4cUgL07CSwEdFv1zYUaRV3C0jZ89Q
qmyRHJm1aCPyXNZt0vbzvtoarvg0A9V0adQFHkz9ru5X91PExGEUYV3GbkCi8ieU
MDAGRg2bTdLR0gk3KOzI6n5w6X3n8K11HaY1dNRaYYiVGbbXDw4CFgGZXBFuKV8Q
EBBtGKISFcQmn/oUlPwFkhoEzS9gvBEwJOmEbKyOBCdNxvBzAGEwoY+riZVDrLM+
M4BR8schARB7TpdDrpA+ReEDnXWYVNGzJ9eGfPcznQTsrbE0nQPXAVBC1Pk5dL5N
h4d1g8Hbf0Kipz+96RnGG2verOkFx4HJZGF45SdjDHYKbBMSbsI3bFzBjgNRPnOh
SAWhVQZ6ICvYpVoCxlBpaLpM51vvahcQjOGIwkw+cvOmFokKSY4yKPbv/qCB/plW
vVrWcfsB4WlmS/yzTqEQrIlwAqNFgKz5Iz1dtntHNOFp3ctyWCp1rZkEtq42la7a
6ksz+zVQp4AACk4N9T+qJChKKrg+G75GYjzOrX8p8YkwDjdT/7lNV/vtbEZuSLFs
XtJIpCB0aShlYLdrMjhvr0qIHoS4H/Cznp4jp2AdBx+qHl7Bz3DcIcffmPULCQxo
+evIW/hWY2AO7L0/hlaCs1/aOONvFapHXa1zcgvlMvIIgIsBE/zvfeEKi1pJLFW6
GOmsp754iix0rGIcQA+2QvQzvandt64Uorht1k7Zcxzplgd5482GkS69PpnBRD2Z
vE7Whug6jA7MKoaGg1mBnKZ8Ii411wdN1Gstj5qWkvC90hJF2wrZjBNf9O2tX3W7
tTtc6srX6UvEtC+lHYfehwXEFJfBO/QUFXyFok6JmOnNfzys1PFB3IB7hgnj+2+9
d8p5Bl75IzLy1ZwGWqDHixAgPZLKObR6u6JNSDwZa2qrkXdk3ccbxlTyXBX+v9Kv
E9oOa4vRQhT5hnl05TVX+QcBFS3bK61bg35lUZOF8uu8NtHy4ZCmY+zTggNSBkT2
pIuRgmq4Dum/RHqR6wD8TgoDyEmgTAoXu9440yu59PAIwbzS1ijUEcJ1bBM2zH1B
oype2YXWXdKgCDRnJhaDvklLERIpSfIroeA7OaPJg5OaYVcoCtWz1tt5bnWtGBhU
iFYcCZZjLn/VADAzen3uQOq1sqiXO8mB/UBVKtdqSBf2uq6QaG2Ahw9Pq9vRNba8
2wUS/8jLXq+nIQ46zae/c329yvNxsVO5Wn/nxWmmDfaubwgKdhsjjPVyIptUn2D+
UqZhfS9A3QCRrytqnqNNQgBjgNw1D0ijsP92qwJAbmXWoAbPPBQk9CHaxhqElr9U
AjvboS3SW5p6ZfWKKaFP+l8vgo0Opa9gTeA4f8QuKqvgRnLec3wTL90UUju9L5Zj
/jB3Oz/ieTRV4hWW+uEvgGKU87yHhe/OwK8mi8Ay7iq2JmdXxtsKrxrVsW4e7ic4
HDrad5tkCajcfD+A0RLlv1QB7obnK4RQQ+x1cAOF7pU22cBWXXffCJyvCi6uJvS8
bZCQlf24c+AUr34E2eWExeKn0YjYpNGgrtj9eK7yadif8djOCejZzIpomBxQOX+U
dqa1c+RC+byPgqSzhWl6xYACjd9WBYEviRzxz9RvjdNDW84MpDoaxUxQdZNRO+xp
zGUIKopLZDv/+qsGmjJU6uk7rug48zHkP4xEcsSfvgZ2YV0qv4f4fZkcmEjUCPQE
jblBQGi4CYeIqMJsk/7cue5frc3BoSIjNlpQbYS2rwj9zpRzyhlhwDyKnjeiJ+9c
D/8rCd7MyD3+jxIcWlGyIVIXWqHtU+HaGtKVa6EONxpdCAymMuMrWrScSkZRyaMB
1aSNu6Hj0a4M5QNCfdEwcQ==
`protect END_PROTECTED
