`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PXkw2XZsLTIzFVpJCkZa9FSKLpvySEyBClO//K6X8MuRZEwlturAiFgXAPuIgtxt
zgsUWFfKAST32sJFU+22nzW+3SM4ZVr1+ONErhlYJmi7PjLRwIu16ydbCKchp0MD
8Eb/bLwzs410FbOcFIjIQzjgER5zLEbSRDH0q2NONfvMfTbXsrK7HikOB4ATwNGv
kH8l/jadsQg55nwmtHvsvYqobYtpiD48TURnkW2U99BYH6Qz47fTYysQGOcTeTe+
2w4iOTVvelOdY66Iy6Eyxlh4S4wXozBJudtaPMdhEc/Xc1XKtPDYFYEbfUMe9rCX
7n6oPbsCnExGItKwfU8ZgDwstMyFvoMN1E6bPFeKgIwIDmro09wp88FTK35RLhK8
23ITTaaAWXaK0zI6+yHTZwlzPHZ9vMymHZMCXHw4mWjSZXHa1setj2NLbOaGfcF1
zUuVIy+IBMLbd5JHseJLITqWfT2/YDBQI0GuOuu/QxqAi+q/UAivvub1YyrXTpVf
krzIgMrB+tjPOVRo+gt9T30rG7elXrR6oUJU/l8QGfh5/Ofw/ocO5eOqkrO5tDAY
X5lfcC8BmARQaOCITKi85ORsp0DOg+26NmHOSUEz3KrSqL3NR4SRKcOhohJj/Q5U
HpHzYtB6+iQpnvkg62G/AwHa5kRdH+SOqQveR40MOx+rY3qGUY2iyfOa6Wog/sJE
aI+znpGIQbNM9A1iUdKnX/Su8wGWYqgujeH4qbF8n1WlGrBABkB3w3BMc8AVnRSR
Vdg8IrnbXEbRb80Z/5iYGws28AkbnIpkuEznb6PR0baYw1oumam+9oEYpyzulWZQ
/mUnLg6Ljff/KLgZmKh8amdSaA24WL52N8fYrlPvQ8DPSRSiY5WCvKXiMQUhSvvy
FglbEuzrfpuCdVE7fqXwfHZKLQNZt8IULqZCr8SLXH6APi+BCj6muY1+Lt7lBOTm
sJxdScrp+WYJ/VFCqhAqotJe58Fr/mp5UWl8906rnbyzPUCQz1UaHEUPCZmwgWZO
f6WZ/z9oE9CxY/5UYnImMpPvwxApalFAE4tBKhQGtG2GWJIWSoBHs+xIuTJW0Bcm
WNG+eqbVFADgXC2/HvMJzFYvYFYlj1HhmyAikRxUbBAMOaLwmziB561RFqAGO+JV
9MQBuhwCcO5ML1q4e+nyZOoZxt41uuGQ6eIIioqn1DFatWI3VNTwunDnic+SWvxe
6LfnObR0Zpqv4JPDKheORo4mMIjj+CgvzodLQeR4jFwieBKuraot9eg0TNQYKSQr
xd6x+k3jhcze7a48+ioRH3aksCQ+6ur6zO1GosaT9ngPhNTQURptu+Js+s9UPXUZ
+wDJkA93pW+FaShC4a7z5q4RvWAOncRqNvKTy/viQnql6obyHt+MnqHlLqWnw0Kd
G0aydqNUJi1hDJ6amC75akJwu/6XBu+/zkTgbMSXfjvgl+Oz1/6xbZnQspHdm5CJ
r2h23sTw7pXD1cEgaouyaDgHnAtrdQKLVuI+rYiKBmX6T0d10HjlLcuNr5s3IAUD
+aO/WsHVj13XfLbB7TkGQA4iuP7tsxUQC+NOjOJsk9zGewMSa6C/6S0hIIgcA526
Y9ubBtjhntBTeMyoFR3jyOyGOQBVY7dQnPMMayUQJR2rkc/2gEOjmcWQFtd+t39e
TIfC+HQQaMntc7TYgzcCCcKVg3BI+6v3AUd0RCKBINpH4ydiydpBWBpjhoKMDY/3
xdUD6/WYdJIDwZLp7fwBEY6uKT80VLD/vpOuESc2lRcJXzTfm7YX6H1xWQRSX1tx
vha6LYMIpJg1tmxJLYS/g7uSkaR372BNbdGhrsrvTqraL3MMPkgM4whdnfV0QV1+
vSQVcu9hxzSTmTA0SPgI9SYYt2K0aHW/2lrU826jITiBe/RExjZvnriGZ3vdGCnV
v3sq6qQYBvQ5+Am0HxU49Kq5BfUYbVCAtCdHYD5yTfSQUoK8f4RqCEHUc0r+BqHR
IK1iYNcHJZXTavjuYm23J78CmuAoMml1L29w0urgD0uuQLnHz8GZE02sfkaqMiEV
DXv4Lr8NGseNKtVrCO6w+S8oM5KjXRGcN08ZdDouHPezJmer9IoWrP1Y+JIJpLdv
rcL/Nenw0z3eQiHrOlbe6rMxiJydN3mzedFdq3eE3lCDA8FYEJPOK+esVRHtIZl6
8hBG9F6JO1VC79bPCg7xcohNfB+dypk5G/3G7KiZX2r94DhKhBxvxibXiQPF1KzA
2i/2JIlGHf6feay/bJBgI7fo0LLvB3v3f1ZcyAeeEMha/1ZEo9EGyvnWg8W+KaJQ
FxddlMnJULKiUHtzZf8LZ9Ivj8NbwC8+bQPIuWOhMWWanyqq8EO4uWnvnQ99X5Ll
ZAqSNLtLAuWFV0OgnWBj0OhJgQ8fpaiXSz+PgQe5wiYM2gD62X4DzOaqXt87vJMq
vSwjJaXgxOYVsjLz9JVu/bPEihlmv1c5cXlkFuAFM0Avtee3S7Z312MymXod/AKX
5Qqu1+JvyP0Zs/PsdwiVDDH+u/XaBD/LZv1572+LCLNlbz0CO9EfS2QqEA/VAmoD
vRSTVPBHGm27yQNGdPkOa85GIxgJAbkvqauhoqmxzFf+xQ+SsNePST3n6O+OHFLP
J66GI+gYeOqfjl3qlsKrde9pzWGvmBKLp+oCfiQMMLy/BMbDqnu4pr2dVmXve5/s
xFkEZYxFWQ8fpRra5Cp8GBMb119h0VadtT4i5G8k2hS+Q3E6shEb0Ryl4HUels9F
nF8NAs3h5nIX5Hj0/0e5IDpyhcw3jhPz6cEGE6e0euqvDRMg2dbype75IQ3sElSx
Hw3bU9khfMTKPMkzoEWpVpSRF25o3hPilHpG0ludKjQdQvayrhIpT3hxpT0DV+q0
quLqBag+Z/qwf26Fw3UquMhTR9S5vrnD4/mRLIpq51JqQFtDRrIIbDQv5Xzu5he6
quGKylYtvj91XntVI50WTfd0ZHGM5lCqw8lHGvgRGr02vd4cOH9NkoWVQhiwsWgL
Dln72Rgensyrd5+8LsXZINGnToxz0T8Qarn6C1mg318qP42ntAA0qG8LsXBaNxjt
0JzMF9U8zCshY61FB454fXdt9/w2DUjjRQls9j+As9uNmEGXjfxqSx10CzBBb5NR
4u11cf/49RafNp9S0DRwyN4wfy6tOCKu974Iunb4zcZIZAj93MBiR8R6jGLNn7GZ
H5zdqj4kaO5vkCwuISOc9AkeA8NJtaEp1JVUSOV9WFAPBYPJ2reSpTMAKgP6g43d
gGKDPP9hOOzzoGJ3Ko6RHgzI6T5k9XU//SEHJG6ZXNqHPZfrxkL63eZUVUYOrSnp
L2km5XNk2NN5BCf+N9a/V51yKySw78BIHQcmM+BpPP8rJr0SVRPJyQMCSqQR6LOG
31SPaIRkDlyDdtq3o1yRWEzR/bsB4EpEWNI9FuCRMQdEX7BUJX4QWK5avIZgOJSN
IpzcsNX3bbE/DyclLu5xhkaZ7olWBBhR140oboduvdJYsO59BFQDohr6phHrReZt
wYw33ZEpnNxwCPu/o2zQnux8wDzmIRxhBx/6E90fgIc7ay48tQwz4uRcBBpDx14p
VsntdAlL7wDaUrT6ORceLcTuqxyK1PsZRgVvVdRof00z6qPCaF0bAo/Kuiymgld4
GPK6HnB7PlyR8hyIb89AISb/r0l5rTYOHisY0nMhaGZKTPRiyk7dB32KtlAXUDnN
CyZxwCK14ypqNdDrLz3KPEC+3YMRPmrr7saqkZPNDrRz3nuYz9yF56l3BEUUllrV
7StytIb2AulFc5kAafX1OKHwBZHHTeKPwZmM1dVa0yE+tFrdL/qjlU/pPp0Ksn6Z
AyPtUispCDxk5Tc1RebE3XGbDBeZXSOcQKYw7csYRnjDiF4wsKIhqdcb43XybTB0
cR3jbf/ly+9azGCf4Cx7JuNbWAsbV0l/2uzxkegEB3nupQ1mZZ2X+5xjJuw9nTiv
HzO2HcnUT1s+aleopF6Y2lkgITNwtqZ6t2V6z/DjCvMqlngzEKug5g6+DkPnViMW
v3TITWz5uYhtpbRcBcevrkYO/M1pYGLzbyV9IRtXu1WKScy5dqbqmHR0cvITZPCW
+BsnHeArOArfCCB4scMzymzOkGhv549J9PV0x5K2qtqF3srSyTEJ9RtuouzexwS2
MHsBEHUYaK8oztW5H2/UepUdtO+9ukLiZuhzT3727NWTKybVhYxZIU4gqUt74jmI
bFsrQVjRdQHs1lD4OCk3hQFON/mg5aSzKrilPCRh46XxHuT5iu9IXcu0xVoXjO73
1+vG28BF1u5ycCft1UvJg3wp+My9E7sQeExNj+F/aHq/uAkBPQqFKRWFLwt15FDd
q7B9uiYFxLyzOow6QcEKWxofnd4Esgfh4viJK0zWBS4CApoyKs2exVkvrmzCuUwU
iZI2luTb3rh78xXgyIjyVg7enAQbVSrlLtrCZNnQaMuXTmoPx0cUupreyoZYkADr
EeXAtE2giiBAykEkW/6tZ6UJxkrIJC8yISC2w2IEUbqz0XXfMiXWu8wb46XTuKbU
a3g4352Jye1CvFQvYnXw6G6r/57l1n+iGsdeCw3rsvv250xQVn7Mr4MrOEANQEm1
vZVSffv25gkQS0HOD9YM8+q+GlJjuwp4vrLXViz6SBp/D7YoLwoxIaAwSYyrtMGD
6EMZy7jrPgmS6585111YEufEs3z8fY4lBvYeGJjkR6g7Nl8pVPGbq5R5anm6zzuk
CDH7uRxIAOZrrHbK6q70A2ok+jfvnbgj2xAZ+fvOc9BPfyEyW/lS+gcbTDVMuQ5Y
wVBugCqaVyXX1SaCrNScwN3Xp8iUNwplXSl3re/gI7GePprvHT0UHaZjd1f+eKb1
+ufncOgIIAW6dbsI/jONPAG6kFo0I/Ez3Rry09rxDHWbtXrvl1/gZvV0us6+WjGJ
TYSfWwVA/PfSgGiCS4lsrTRwIMK63Ny3JppNyd35xX2AfA/5gyKLUkiAloZLaqnn
1YNd9wPTplzBynJP4pq996DONrAesI5eR1SQxWduTSt/gfPV/gwxWVUcFIXvMAje
C2lZ6trTo3ElxPMIAShwB/7Bd3pYoiXOS6P6jadsg8+nVFA7p9waOL2JKWnFv+8N
7WiWW2zPDzX9sKglV3NpzWvSv2LXtXYRW7KVEb72Cwk99NtYoJZzogZ3uCqGt2+1
6FD1YbcEg+6q/hnQIasqZzhSFcZBXWGedf/lmmCvgbBHsxsEl16OS4RUZ2tb1whw
X7+d6wYX5Jw0UZ1onHv55oKP1KoHeeul9J3U0/O29U0x151nYKfAb8kTvTzYCgNh
eWbZq5D+2sCgk7oaQXHyO5mxYRTjcXrZPmZe8DmOteu1bzJ+bLG/pGh6CqDWC1S0
NJBhjgqe3gJRFRzciRt30RHs+Ka9+dbVfJUEJoKu43xuckjZzKnmwvHWwEKLG5Eh
Lvrq90xZn2hgi0kjxyzrU39aG7KPk2c/AzL1a444tTfSChGCUEiEApowFWUSrkJc
pOLxnTSU9le+XR07+ZJKgWHQrdjyl8JAGD5qirSSoduAF1LpuoCWuIOBkPPn4Jpf
Q5oySi3ngyQJq19ZQ7upCRc1GcLThOK0iQzTcRn6wzhmfZD8+2Y7VoDkAGa7tZah
wy8damrF+GuLXNGPh1lbklwdFCi4zIZhfD//pj7CLClEicMM+H5t9Zo5giBQnEZb
sScMYCsnPv0BvdGTxPGk9oU555kP7300qLIz33lN1Upj72WIYnQ40fGKbNa2mS+5
+leJpNHntXOmmAT+/NVHrJf8xJKmgdwyolgR8eNaF0BlomEVC40XP1bNm58hzkn0
7tIeGRR/x/Q6MIBP0VeWkQx3QLxgTuk8s+2e6C0RxgeQ40lXhfqFy1cQap3hR6g/
Sxb4Qb46nev0oeH0NAtiPz1QYhoT91oHC6bM2Z+Y+Q4huxJGyvvCCAT4EGUPICPB
DmNkUxx7VBw7fRygI5vqah57I8pVsQ/wFB8k25Ybjnwyfoiox0XLZrb7wO3O4xJs
jqFGKgyL5o/P0RNB3N4BmPV+Yv5jzF2w2JjWJWUp08l9fHDaoL/H85XAM4UkLUMq
/Wlnmi/oQ7UDo2i1Z8zS7gNMDa2iRk+cbPcHjCZ5tQoKgdMaOzpxM/46bTCQVjBR
a/fatt67oMJozXcjxgd3g6b/+AQkluF9dlcu+49273OfvGhJEBWJpSpuH/mRj67w
MZtUV0NROsqAGGafXOgbGaJzaI699F4B/jpLziFMNmFkO2ua51pWU4MW8aaOTFau
kJwUwr9NNVYvSyq5oJPQbVzUG4ztjFCSjMsXsxTZM7yv/mRNLWqMoRv5kr7qjEdh
FtXv+4hNqemNDewswWZZjGesWzrSAnvSt30iL1DEPUNQCk1CcQ61/UkogazbQpIC
xpjOTcK9r5JkfU0nAifcjaPmkbl/gCOJM00wlumh+koxJnaRw2x+f8BOqLDnz5RQ
JJKGYb2QweR6453Tn5lqAsSnvwlSRpnzNEuS9abWm+Mwzp7VJz8KWKyckbmL2imk
Gc3aqbFpu7XoKNC2ZMBSBUZeI+OLPDokouWFAMkoZNSy0Ht7VUmImfqyAkRZWfka
RCXTupIIcWjK1I4aOExle7fkUioQPdb2aooM0J8prgnbcAOcvY4hFViWuXckjhzk
rmmGNjnOrfCZJWd3bNzG+bhVG0yng8w4vj89n1uK1Vn6UqmaU7W00uwdMbWsCqBT
JDy91OhQV9cZ5C9w+lYX8yiQ26P2pCYuYXzHjso27wS7CtL8YTdH1KX2d/EwoIAD
o5NYcdsLUuMOxJprk/sXQcYmwQx9LpRKmQVS2BVPLdcF07mvUuw+isTUp3ZoEUZe
AgqGxD9sFdIgpX2f3i225A+LSAZeqBuBuogGRsCt0h42N2y4AZeiqcCoRSF3deg2
QCy+h0FJMao6ESTKOzT6bqh/Z7ysVcRBn/9xLMrI4yizEqknNM0lFL4ZHt7eu/mI
0sxYEybkyORirlC3iBWp6YOoDbqD8l0ELvge52RJ4/CfYeqFl2IobsBhcUANG7DT
5eMGqXfSNjGgXdyFpN8E5xugVVnq8uqUeq5gMkxXgrrYBlyuxVnKytKe4fOqsQpE
9qNAHAyeaVfKqMPbT79WCcjF2MLVMcBIBDI8FLpWQ8JfkTrMW09Bd4gpQ5D/wSrt
a+kEQpc2+0Rd/LqrFVgzHWm2J9x98qwZVvU+6mvqQH2j1SkgzCPNt62xus9/GQnw
ZiDH8oQMWa1T/on/UtJQ+F8+Bow8tppdSmKtTr8xRAprkqL9ZeXKfBNzeDRBULQC
bmyDM86gzcdQsXVS+fGyUWKsm4qXfjTphDCGkJIByIEB+JrOF6jQ5PLX+t0GD2eA
L/3w6fyZRx3ZfjtC2+D27rcwG905PevdcVxdNSKAM+BdfgNQAq7ZA79B1FdVH/3k
cLW8lMqWt8ciFigdOrKFmm29+g95hGZRPiao4SY0xZodKN6WXeDLHGpLFm0vgkPo
fQBaSkV7IvcJRB+xgq2pbe4IiR/BIr9B68845yiMnV1KpvCOqLdbCYIfhziQ1yRu
hySKmHY4StfflZJHGQ4LeBW34BxqWS+4o2nUJc+t05z81aA6Q4txxC9OwZnlGPvH
x9LsiNyA9OE0r8rKX6BK2a/hK96UvBCHik3cQ+mbub5RbmvmmwfziOAeifLtl2L9
4aa+Ra+WtjsnDwuyCPSNu3SzfVzk8bfk9uludHzthrjkaY+sXDBR1vcMqTCEFxX8
+KJTQnQeYjfNrm0Pi+yN2XMYGsXVaduCVk9Y+pwdTloPtAKgNTpzHlOezIi+FpEt
IjczTYRNaJgw9pLxLLKz8bD0QG8sFS14+z4AcHV/w9fl36UNByuydJeqDn/elLlZ
xMJ+lw7XKX9/QeNuN2V4WIJBkw26VWsVR0cHg1ZbAH1jhHVGIeUw/J+4o++i4kSV
6YUtSemmVs8nzCt00OG8nanVFfJjfRQpKusrBeEdJVwOc4vbJKRrYt8PeoetCiZL
61iBPU0SMM3bPgZFJznay8L+l/C5uEY8fmqydgOH3357tByUGUYo+8PdmrnGQdZk
NfAgTL9B8e6UpiulbXNjgdrN7eyg4pQoEvYDi7kbV9xIcts/xe0ZaPidmrRHUada
cw20m5aqWReZIzcVTr7DQE+F9fSmPr322YrrSuFkVdRYsetvz/l5LDZNVw6LBJYK
HzfbqAe0/hZSZWYtMOKYG9bB/iwwCthYCac8IIQ4oIzKp1Bq0po29vOmiEMqzsvH
+V7VDD7Z3FmW3hvd2NZXdP5G4ySAM7T8NfgetO7X33Xu6HXENijcSXogWVFaRw4n
ITYSEmYTbvzonl02Aq4EiM35ysTMnlWKobn5L+DKrFHh59TVUcONIQN6veqZAmjJ
/u5sgY+bqANmIYa5UtoDSzEHTqyZNGZjgCJLNwZkSWUTTDDCW7s/CZsi6t2+nUT7
whw7JrVIrcGwl3ob6lNP15fGq+tGhHDV78u4aTz9ss9a2XK2bXq+vPdCLAE+YKH4
R51lIUsNwCg8+Pb77DrxQQ7w8/anpCbiK3oZLD/0zANffV7ApHQEHOnwKqvIVQg4
sdx0RsG3RZszdzhgrWWb6bc/0hXSb4uk0KDv+6LlceVlCecCshFTNAFRSN9E1xue
jiLLQ2rQ5yr0XBEQobJnGefV7+GdBznOnU3+6uv5+Ae51s0eE7Ebah6XJWG0UgKv
eZ0TM2bSqlh+iNMEG1Cs6ztr5kSVQ3I5fHzXRF2GCmIFEUAQf512YyJhxAAx+qKq
0cWVwdBSHszC/iPa3R1WAkBLx5H8C4gbPLWL4Mdb90asEU7828TH3/MGKwuKv+8O
VR8oGcND1df1xnX95KGQmRuYu4TR3R7R/l7oJjA08t9IedLD3oR0GB0R1SwiJr2G
u7bZe/ynylK7D/4m/YV7prfC+82ssQ8yjTzFJAfx7on3V+czbIMlXWuvWqucWiHO
VN5apxhunZ+HyUpmjauc77JLe/w8QXHhcRgMvLJHzL0029V2NorDQ+Xr0Ix3Uppy
ZzSvNLcfrXHid0oWt2D+M+9tWeiOVohr5i0jcWP0zQl8GKWTLCCqykb3FoD3KOAp
IOnj6lW2tP0feVGWNkIZGoLzSyiWgGzppqnjgN0SI0NHo2SwFHPXKEJP1oFJMHvx
E8PSHRKcaUxJIMo+3y81ILarl0ygXumCsG3nLA2khRllFI0KZ3lQScCJ+mRgV/Sq
asjmOQPO/eCd3D7Tn5N6pcI4ZS8ccr6xLNKSFSzR2BtZJ9HZV1Uorywx7NiiNowb
jENTxvoDEXPbvUJdtaxJmI4B5Tiom/dEWqnjaGsksT4hK0NN8wHOP62jJGpvq+Sb
05/ej1cu4yaSrPPBRme7o8wX39SVuQopgr/FQi1+6hE1sy0+bSj2AzbUysonjsST
SWUDuFSlk6k1phacgg2pbNBed3o94JtKUmiqMGC/uCWTAt2wLYePQ7zbTJnWdGzu
`protect END_PROTECTED
