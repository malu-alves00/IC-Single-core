`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uEgK7ihJDD5EYSx75jVAHHV8eWt9xj4BeK4sjlvbUAQFDmzbV9K7MYWOeEo3/637
zWl6KvGaPFaOhFrnXddn1DA7mT6KjEdB7qeRIbGjgd6WT9aryXIpVZmt+wgKKbMf
3dNZLn5mf7OwUkMDOyieIQ/UJAvFylRpkpYixFGCrNuib1sUmqWUmyHkuMlwEpDF
6J0RGfSEeu1tm/+FxzdxU+P4I/C+gtrjzpt/u0QugtvexJmUf9kofcHW/xhEZ4eZ
G3BxAEBqQqBAIeJB/Fet+zbeOHnWsfh59aO9C/QczDog7w8vXFO/NXCzYr4kKPEP
iwYjhsVBWJyvKAnp0ew5CsjwGDTuJcYgFskEF7PaPwN9fO1On/Fb8aoUeroqD88Q
NqOCFOSG6EbHCk2lH1AVtEvZ4r+iLB/3OKCiDELtxNUGQ2x8zWMxjpXSKNheGSSD
1eEVDIMMDqrw+JXPtTt3958ebzko3K7wwFIuf2FoIW5ZX0JR4m4/7+NKtSnh/aZl
FslnGmTT0l1SPrFT3Wes20zgofbUaFCAwD6E3y42+R0Wzm5yfsjuD8nXuLX8XZQe
bzBGk3GBgLGneQJqG0zI8nv1McqB7S3A2GBvkQXquGLgBX4FYhMmU7b7C5pc8f4c
qtMsEk0Xt0dVUnBupVsGLEpRbHg4qy0198gMhD943FJM9u9tcWL2LO82ufg+T1SG
3GdZx3856dBHohUohkX+lLTpnYlMWjXDzVVmjjS+t6qrZSRsxdxxmOpxJp2hB688
dm0YffAm12wE/jcOMIPRZo6oI9n3WjmUsh63O6w9R9Ohdeb+fb/Mjf5OkZSEPBEe
7CcgZMpHTWyJpYgeW8Vs+gG3sjj67bWLsCDLh8acLyrauc29gquc51ONbVu4fLQ1
B1SW3iyqBW79nd/6g7XHYtSKX+2Ur2FnChe8t4Tc7N1hrXkDWll4BSff3mH/Y6q+
8HIw+XHT7TzlDrKyfveXwd/6cq4l7xz2ag5Wdg7dzrV8fybXVu7kZaJx2qxKVCoy
3tDabU/7GqATgl4qYI6bza3w303PdWtuj2yo3XCM/Z7KQUS5E9364N7Jqp+SdgPj
DZALmQL7E7QCcuAgcZfLqbgCD65EcafvZ4pgtBbR5q43AIZg8leECPYU18l9vYSt
ZCuHvBNlXbhlGG2frtTbklMtVRN/EQRRebBc3E7L2R6B+Xe7nyVHMxCjRHOEK64X
GXhfvRNhFrMjwdvdzKDhPn/qQs6+PfZ3RSM18OwIm/D6TnqaIj9X3S+cQvdJSHgK
hF6J0bAlOTwSDktgbxNHDNd1Pnnp+8+MKIW42OCrlxtdr/yTTf+GmluBQGthheWo
j/p2clb86T6d2sbrt9e8G5+NRQ2VY15dOnwR+Ne2/M+YqqWr1K28ca+Yk104VhNv
pnLXxG3GWX8h5A7mp+f+6J0yzW0MXpcx5D9O7s9uAEGmN93Rs5jYcMCfa5nSz2jf
vbDlyZszzQp91vDzpdc14EnnX3I/BRGqZvbe8nAp6ENRUQNqsblTgZaNXtkE+2X+
XQQMqmnBMWv+3rIIXdGn00eldjSW73oJzfMjM0EEugQJWe2tuWqGFy+8qYxFZqbB
ED3IMjiSl8TeAZAJO0IjJqnBgkm45ycJFPXxFB3kmL5K+z2myeERtT70BJUEUERG
pob7prDqurTbwlGgFoZpQSPYpf67EZkvSoEHH8TIjbKdNc+o8xvFo2kky+6bG4vg
lGoh0wg1n66ex4GZRtgq0pdlG4hoqd0UHvnR6FpjgOo2EoYhRfNGblcCajCzT/2b
sy6peYYKUbzGa7kk8UBqLN5udgDgmWRO+6tKsU8PkQXsfvPECmVFod8F1nWfEDGt
THBR44mLfhdq2oVAYi7GRZK1yL/0WHTCx4OuMNEKfmkLRvIK8IL3TMw5kp/r403J
O/ra9h3ZiUhJ+pyvzJWYPaPW0A7tuxfJKefMWcDCwYk7F+JRPOgcE81MAo7mx9Kd
cjoVFN7Akd15/9oZ1D0v0z0FfkQ2JaFR+hTG3+bfbTOQIn0hEgyhV4Vl7ud33tfz
i6zIaLPW6h240FGeawgtXYQJbuyBkRQ7egGpBXR+W3QZyFas23/NKJVUXsL178Lk
0Ja/kVOb6qV0snYTltH7hOfE7Dn1eLDjJ3LSZIbiFJVoss9Qro0f7ALRBqyrTFc8
5EbjjHsOPNTwMbwxI5S24Es8Nb7henk0c+4qb2y4bizapvTzj0ylcIGT59OHMGhn
ZZQ172X92sXxQR/ZLlHuNW+wbqxi7ib/9xW2/vrQ6a7BwDjkpdqV9ijOyz6LlMhP
Pukzf2dW7VN2274juOXiMsxvwBva4t/V2Wbd+4Ez9l/6tzDH9iSWKZSz852LC6xp
bWfZl89Dbdf8h7DSYkR9ZquxfjcQ23B2Zf4RJWoTiw+FrAbbJlhJi5ilGEV1lsdt
GaF7eVCr5FC2rqQRe4QSObuajHR+o9xGvsU6NKuu+zJdVQOsFpHZwdU2wLyyQanU
LZ+N8+V9YA+4ZnXezoNaGYRI1BK7C6BWJImwtQJnL9xH1tYIevaRvX/BSu29ZoZo
0ceFIqqd3PcX65mlvNE6LFuLMbA738Ni0r7PJaJnQuj6z5LxAdhRdWh0rhgGWx2m
rFAPFj6cl7+G1TTGe67XQKzW1eYH+imxtCNvtdTtM6wE95J/2NMxjsDPzjLt/bBm
b2PRhnskgY4c4QPpt2Ebc+Y60465zmFovUcoP6+yHvyH3h7uR1H9SdAsPg7p+ks7
/PnnlBCZm/xJgQt7IN+uxmSg72QgayBl/2URlfZehw2Zsf2AYR6FhpzXSX6cihJN
um3hKIN/MLvkey6o6+O0vlvOHKiRNH1qbQOnE7uBh8iGWTqE5Eqdi7ud6lmUJmY5
dpr2K1wkqcTU17pJAszNVx5jIMR6UfGtrb05uAJgqkMS1aI/SZUdGeWoVcgGC+Xh
fyeK4jbWkXebP5vF/StJcNB/b1QDHpwrJkGXdTqJolA913D5GB/e+c+DRuVLjQDS
gLozfZU5T2OagdCB77ZF/plbytCPshEdlK0pwe/nbCYqmn8JG5AGvrFvIWDU385J
uFPoOVKKwyI9aiMPsCq9jOxkF9Ag2R9OUN1cDoSr0tX1DGZ9f2lWIhNpK+YVbucZ
1mHwFA/biGaMI7qXX3GDQaxuKeqR1yhKQhBhWrNOnsbNUjGBXkR9O3yj9qIrExdp
TO+JF2yEit71ZrFcIIUxNhl1dXZIIyC+OdJY3fTBTBpD4uuj90LIVCHgPSezoIKJ
syE0BEwE5JjNbWDqvd5wdLEtxjrxrYM+8XuetqLGu/pxz5Yy8UpBj9wxyPPtMiVH
72D0deTYTIpKpZkJeJgmjS04Yg4YuPEMF3nlU7ByLtJN6lkcKjNcutxebpdT9lk8
dg7tFu6P3XDPEoOqAH3yrI47ilRS/L2N8d01PQwTmQUtgUPIVJZxaWFfaTyy2chb
FSFXF0NLEfLGJlFPt7+m4YJZvNWdvu/1FrQxwRm+0ZB4KgBBraUwiiwsV3KCSaH0
u5O7NqjVZ8Ixhql5GKm6NJE/8XD5M+JNf953qUzActs25n+oL6gUBbBOWmXK//Yu
mm6byFOq29FirxHI15Vk7x+jZrTQuhb175zgwZS8qrQT68JCHEiFQJtirijdb1XX
GQPQKyZ3jhWJq5EgAiqnXajP5ohrwvfo0pe1YlK3xQFf+c+kCTALJYCwtJrTRjP0
GXQu/5CXNovL3Y/4zJsUs3W6IVfoBJAl5gMfKtgR9wQlLgMxUOKT+3m12zxd1Isl
z8kllJBx94WBSG5BeAsXNd+ltU5eygpz9Hxl1uKWQaq9+X4qYvaW3Op8SsFLtqmu
EL5gnIYl8jAEt6XWvwKfamAA3Kq1RBM0zjEx7lLUKM8Dq+IMa6bbsoigvljaBa7r
DolMPDl+AapgERbpt5Ks/OJEs/RQ12doZBul0FEjcnMV52J/TSatGYB9H6HxbIgM
LfKs41Ahl2vyaWY4QWKEGwlzGB/0Gx0sFwXfI/2vlGca4QrYum6gddZIsuH2nkf+
BOaBdMTuLHrpaH7aj4wTJk1iJBBntil1TOz4Rj6q1VvLNydw+sEM4EkbWdeS5hzN
OavAeGacB83qwCGQfZWGQBG1JkrVnPAYtJrjFDJ4ZKn8j4ajVl0vhI6A+aJ23+5S
QcHYHWMxFPvvi8gONffoIt17Ln8BtOFnAOoJmwNvK23KCx9p2VzbBkNVU9HjIWSc
g8Vpd/i1ZRHLKPXZPbtyfNH7tfjRChWTZbfGHtD8+RlP/Eu3BsBB1PvSJnEoJZe3
3ilzPFew25TRqfFn5iJTSUX6wvC7VTu1KiaiRnt9cQ4/Wyj6ORDBgOxypDlFJzSE
ERTaNEJIqbjj+TJHt40wDIHPr1GaqGj4sFozgElATft0JhztWrW0sWIfP1H4iMZS
KJ4pI14JjHA/FNv22JhMjjRVt9dQ0Lt35A4rxT8hnBguP0Qr9atNInDyCLccff5e
cLMwoTgBP2kvipcX0meBhYnbMi8Z0HSkn4Nwlq3LS0Odg1wD40D/CXXySbQc/Jdi
deKkrwtcORg74g2Bt/GPQQ99WruRW0FAOy+ebG3vFNtzO66HJVY6GJlfA46WvHGV
cCmFpUILcEHp8Zlt8eBiW2PknBZ59O6+1s/UctlMPfTdHv5PicAcYxSLeMZxamqZ
F9LwZVE8e2TFN0lLpUmUnZkxko6fY9mHlRbokXnUoleBc0vCC+jVM1FeEEWwCuDy
8XkOf5DBAkRQ60koHZ7c9krH+kymB1I2KA9nDkLQ35yWm/rIvl9ZdXDd4ZHAJESA
gzb7IHWxxc/P3WWK3w0YzCJIXDeNo4bpXMqKX26FP7LK4pjQ0PiHfWKUDZw0H8V2
ezTp4eU0kH0Msn5fCyL6L97k7Vk5tezfgySO9aTKsf8Xww83VkKdlGnU9S9MinBH
T/lG40/IrveOzfYgxP9k9UqNxzkaLu+NjQnKLVPAjmYDhfmsU/MfD0uAgX0jiMKo
HO/y2YgfDFKY16WIws3NT9ReCtD5I6ZxplDgF6dy1WmN+cO7BnO54MTvgPMqBAF5
YdlWMDCzG1aLHbBJKLumFbPONicRjuM6YboptdwM1TbpxJIdnosV9u/GQTnRuZnZ
/f6LnX8ZRuMwdpRuCPQephxtN4wmP2gC5kvDp15Dp2pE9JtXfVEUJ5DcgQzhBcbc
SD4Fv3u3HHviJOEaGwTN/Io0Ndzjw7qYa+m+08FYrDDPC12aZS2ihEd0bEInXSvU
2tEvXxdA3eKtNnPqaYd3Y4Gpa4uX/UavWAUuVX4kNXOQo+u1qcDkll3MAb/mpgnw
+7N4W1MP4e246ChyoZH053cDNxtBN91xxZDBObsWCVrhjBBXsWm0GASbwEHPzqIG
WQ/zdXH5WPEwgLrUZlSIo+x10G2TuRjcfvqVrUyWsooZqezUp2rGEEbWdcqfIpNX
DoUJVZZef58wFHV0IKpWZPvp7TavMTtQTFxnGvsct0VDlxJBU0twkV0lMKKwAsyf
D4HtWsHTfJzPXhQuO8mUij0Q5Py0UX8gPF3o1gNYbR2RRQ6D1biUOUNWdGBd1P4q
H9O8h+9dSP0KLcRanaO3XQve+79+VUCu+qstC70LOKHrUpuwRdFrGJUpkMo+5wwV
LFGU803/RTyFwFqK0U2kQHzW0p6ALjP6wca/TmFWTvJy1p3jbI62JrDBrRqvIrWb
Eoszf1XPHgHmVHwLm8mWlvBgYpvLfDSu26xqNDHo79GYqYEINMv8kjiuVnUTMPQV
M1WLX8gerIDLRbRsqYPcFItozg33D/+o8YzBdu38gOiDXyNLLFUpTqZWeBvXuF03
wlv33cHY3/dnmS3oJ2Qu29jZB5SzCR0G/1SG1mJUolnyzbWTy4EXXX115S9Q3FLI
1Rk9h88FLxldG9Y9oZG+4+CC8iWsfQEKy9a6IawgkxcH/LCWziJlSAghy4Iwo1nV
M+T8tFhUuVdqXENcgRPnF6rXqA26ByKS90x9fGQEJjlOQAlsl2ndbbb1+PUku7VU
L972Qncj+1YdaUgW/mZNlHUriYJGII1KLshekO9/OHERZoSKVCsyAal/EInOkVfU
89OcX1s8GuDH0P2btVsyy6LlmQRKGzGHP0tGT0KTuORqnhSWxJLZMnWGrVyKBu5L
plAqGdHdC2q8yOLOIFGF9BFsb5Fnh4KFgEds/1e2mVllo0Aidx/aW2KAlxyFmb7z
U9ip5fbnnf3dgkKTykXGnFpUaLFmU57TOU20O0Oe+Zv84r5ttH7nc5fgDzpgH8tW
5hK46EcC2GTdNKLKQEGN454LuIRt7q5Az8mshWdf4IDfy6sb9aYQzP1bB7TALziF
Y/8cZTnSmoxiQtrT84skcqKbjTTqUWFFYnvNcfVajespwmB1xLmUaI3ngC7fwTwo
7zcNnotk5znpmzYDfywbmuUV8L4McT7Dgxkp6u8EhAqTeBWuMAoEmHvTYmtiu/Wh
cc7Fb8uQzBZ4bnUwILm9N95I05XvkhX1pm5kAosz1eh8HQcDKiBwAkeC1lVpsEh8
T7n27nGIv6JebqutbBGjgKDGmjEtTor21w72fgXC24Z2GpjV70CDxZn5r2THFQPr
KAz8sattkaRWpowC1CKIhOXUUBdpnGf2bLbx4+VC3MKJWcSYEIKCTUeclJyVtoGa
X/fSg3Fw2v/qNuaK5nEhYGSRQykQ4gCfoWKVzH97PujhM/RkqKUTvxfk+xxRpiv4
wUBCGt5MJbd5fj94PC8L7Eobg4kq3Cd043donN9Xigv332wyOvjnaZu/P4hj3Dwm
NXwwllznbQ6xnX+YgANHUlsdspMmGNhy5mr+Dt7BauJuHJZf9dgB+ChgUiGAhxff
jtA9JupqFr+W2Tat5mq3jnxVk7e/0UybNeeADgRt/pr76eua4/Muil8Rm3sIzKNZ
Xhwed4P3J5XG4Ty0r2tos7P9yq2PYgze8uIYFZat9hRB69406LkgPGkqCcnlNpBT
5f1UZn5XKReYuA0bhzlaYgVdyohqHJBL4/lS/W450lnfPosL2FJ4JC/BpKwvLKEv
xD1OE/brW9ehJH6fwboKu7SUjRJ/cV+6z254OBA1dXIazdTp+cBmp2BYUiy5C8jh
NGIezPw2Z1GZJpzbpkA+sGY8AY6w9LeK7HHKXg9021Mf7DV6OSovQ/qRtAnGr/yV
AMHxGBlVvyR9M/ULXB64TZ1RneEfAHt9GlbqvZRKI+JsbdDOKpnIQ/SFiuGF0c4q
2CXyU2ImSDTMp74z05qV8pOSOOXadp5fCBNF3aO8av4E6RuhIhPIN0BVRb3FED+3
AwlAoyl0QujwFXDVDpCeQzM1DPyz9xxqN9m+hVx9OFRAREifr/zSYqO00tt1OKHA
hxMk0kQwYj47LH9vzfDrH2V6r8uMr8M0NxXSHCzoyXEmKH0zu0Z+k+slwRRBpqEi
3ftIa5OgokcNxdPjSc9RSGicXesGpOCmW4wDFaLD30AN3h95qsHSHAwLqBHt7Cg1
lyjLPr3SvI+abuiTwY2LHHZcYfh7l90imiTNHCzf/KHHlIM9bzsGu0XQJjj6o1pU
3MFWQfOjkHxvSYCLHcGYkwVquwAlIfHUuNVkQUDvtPeuSn6X/lTtAfQA5Ya/Oklp
+g1EctPq7LBwumj7VnCwRXEL/XeY/PAt819XSRwL7Dwd2VO0Heyt2hOSewvhWFVh
S1Xd4WBp0yzjY0YFFhYwkkt7co857DqGV/W7CV+e7n0ojBeF4pD6jbrhJm4tYUvV
FYU8pBQHBlaOga7IB7iuS089XcFrm3ehbkb3A5Al3w4AVecodtAVqtfH7WdBqADz
Y72VRkzYfN+haVcRtLK85rw8H9IchNXDMkVzURJBxeh8eq6RsfTzQKHpUmmBgT1C
A0l8Ylt+NtPMHaCAtPXWRZj1BF+fAotfsoFWxZmnRQRxdJj1tFej1av0cBkKEJC9
9ZsOV2WoNnaz8ntobavg4CibdvGEeGOfRHeXJAc2Au+CGYYtKrXe8PMRYzxEq1XJ
ZY+8vfW6BCKPB2K22Q3zzdqocJSgskuNrvzoaRoo+OQFo9wQCpQ8LfNptNuuJddN
hqsu7JTURSahwh0aIJ+lNhWk0a7d8eCEvaxDKjywi47Pj7StGHSrJIvHz8qImJZq
T9OaYchXJyiwFBLRxo3BGn52QR3CfAd6BsOe3Kc4YEY64jYued7qv9sa6H/PxDO1
rxkZXPOSHQbeJBD6feVa4YdRxSQict3TRKt9694wK/wpIzVsh8WR7urYySnmD4O1
XmgG2l/rN4u2I7zuWcQcb4Rx8CCZCQ5J7VZgTY22ydT3ngl0VFOcC5O0cBLounPi
gtqg6/V4IoHuSOxVOXAIr+8LdcfI7Pxxp6I6yyR2z1AePfnin9edUeOBf0JQnl3d
L/aXmsWCVNnGAJca+Eb9aIScOAcpuvoqXF77ITROgRozzL0Lcyx5hogYhSdJt5pN
TyE5V6vIhMzyjQkCKHP7uANTYcR+Rg/BC/UUqltvKTyp2nPzvH+XLERuJh/s5IW6
Q4Yc+YiGFBQkxnZbt471//e5S0TJh3fSiH0J1ut7Fm5Kbp8z/kOIan9bAOIi5ebG
TagZYJrKciy6rtG18DLiSkrWBLJNrEhgWCXBCJ1zC7KgmUQ0UOmYH87KXnFtGzv2
HZj+15nsduMDP8LBYJEZ/NrTr5PF4jDDhZrEPUtl6LNRmt/XR0Rm0o4srBNZhHee
+4gOjsSf4DNWZh6psi5EwkSA87jFVKxiaI5Nwc0G+8mhNLu0AUIogXnPjxvW7/OT
U/NnSOZSnwbCI6TFNooImKr87wUEV+ZWnv7x/OLiy9G9a50Eo/+xcaQX/t5jFX+o
pwALnmAriCllp1x1iMzE6X8y+VD3g1o7Ur2hR8cCnoS7Mdhgu7bN7M4EkjyYCz3W
2Q1IkBPzTSUjAZ5DtxAG+ZrJBXwvcu3GJmf580X1wBJmciRY99A4SIgje73pS47y
pGzAnYv3VjSe42k7UVKQxDalS0qv0ipDt4DRsfjt6gikTcPHdvUPbIfnd2VFjuDW
0xx1BD4e0SM6tVDh3To14LcH0Zb5FdAzZeWvgr/kBzauA8MMqiYDQTEqZbSmlsm1
MjSoR9z6+ISR2n5eEwpHUVNpVBSxixzHd6SSpaJKf3CmO4ayT2irk94O/XT+TCpX
wvIIM/1pIQectnfiEcaXpJZfUb6Qnsbfjs3TGjB5GcynFeglb5q3Ll9NYY9dd67w
PQUR8+wqwSQ8BynQ+Y20OuoqcB6cvaA9ahw87zte5X3TgYND9Yo9Y/gIwtf8FJfW
CM/Vgj28IR3HAAbosxFwf+XKW9xePH7AZoQYZKy3yKGTt53U3nZlnDV5ONPKjbVL
TEQjVyU/Hn3jjA1HGrLdlumCMd2wipJq77ooOG0X9anSuR4egyDTaxSbe3S3cxJ2
CBtsQ6WX9XPayb0z566esQeIMajOJuDzxOgXQUCtVxBY47oWj4pIvwzwAa+OGjn7
`protect END_PROTECTED
