`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VPKm8uPLeO15myfSB058qeyzWXPcHwHHploXLjN2GUuGqpOpQUOfPKIqIGUKMqxg
g14JwcYP21MaS/hYgKATh9ubO2GvUjEpRE1+JNrlbENqzMATwYGCozzPA4yRKYcQ
wlovHCKrHnUsLqWkXxwtWBxUnsltJRyYBYWVufucwP4PcgEnSR8JAvKcT6G/xVMi
Wg8p+IJU5tNlxne1XgVCY40ZaXv00zj1zzcN0nkSkuNQ+QS8AF5Ul7LAWA5PA9zQ
6g01GxLP9BRJhHlcVTbhNFx3zf562F272VwidvGnRUcWJqYry2dTmfS0K9/sc4s1
7AxmU7S7EGO+9PzTvOLHdDuAFk5IgUPWS1s4tkABEHQ=
`protect END_PROTECTED
