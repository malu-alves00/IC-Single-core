`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Tr4VEKJfqt8h4jiFCKgAV1tAsA0U9z9STfgg6oyhVrloKvQFmfVAWgl+QckAIDcp
HARoCTqsntcNRjauALxgDH5W9DQaenuVssdNkbenjI1Rv+9G2R6WuBKvJ27uHXRt
kEZSVTHCr6EbiTGA+C/7JoTQBthRgxIaTS5F27ZVuhNa59wgooTj/+BvDqY93+94
8voGjcjU2gIxARCaScVCzwIamctrabNjEnI6HHa6I2EEIlmxNWxkF/veKOf009hf
qMUjce7z/1JJpSRZ5NJMIk89WYadmR8MORjGu9N2xvFUvkYsispgnKxOQFBs1xPw
A+T87RsZhcDJY8cUOfyiJEqm8gWmpqJTcPP9WJ8CeGk5BnWGxcjNn5eZogDcoT7m
tdb0RJ+wZOfNq3hnstIF2cnw0x39/0Pry2oug9tQnwjTUAxTZd0QhrMsHXgPrNg8
prQv5AqbwYrR2QKp8BrhDzlly8dC1Y+E+/eZyp5L1x0dEMYplgwcS3+4fUA5OSvy
eA03hr5+KtcUL+RWQbh1Y9lILevjoZTNcvMLq0gXgbjT6ksFP6Yujm0ito3kuhyZ
4b6u7+q+G7QniHKLCxPhlyEePilaHZG+lTHhJwV4RyBx9VcIC5ZCKRqaqlRDoXgU
wZDKigxnNv14eND8NDO5n6BgxBaOUhcKtesjJD8taYeaWeil8asO6Ovq1Q+PEP0W
`protect END_PROTECTED
