`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CZC/O9By1YpWtDyEe5GYWi84N1YgAPBKlyXmsNqpI1oc6RxoEa4g/iE8iE1aFNRW
zOXxdWI07TybKqMyp1/qxtSPlJhnW8tdLwNBGEkEHIiOXd7dLZamZHFZpvu66hf4
rqhGRsr0nDeK9MPM7ou237QZWQ1WA6oL9uAJgoZMVQ/Ovd2BnsdA9OzguSrdr5XK
yM1VOioMsfrWPCkZrsZSkYM7pk16F/Q1K/eKWomqH4vy2kUZ0QzONxrPixLqVJOT
BzDw5d1tciA3XGhWNWSi7ZDRQHG8lqU8pn+GURJXCo3RRCdHHSRt3E27ZCnoTodL
Sd3GX5iI6wT+E5dLeoCTT5586gQ0Tbni0SQBKAOxV2L975T1fJF+QaMgAv/aU48B
mj/t8C9Rc6h3pCEPvhYU1S1p3WOANYb2fhsdKGBkKmLG/Gee0mDrzBH87vt2oqDx
S482WHWbB43yzJJu/f+01r/OSmtSO3UFgTsrI/9LFwCTe/wkRvDrALY0j6R2InwA
gX+oLVnhG1tAHCbvh5MXnOWf8W+GXGnz56r4h8HCaSc0n4oclsqqNxII9fKwsFv7
4fNP7LKDXpXi64/e4XtGBXp6iRb8ZSoLQe0BCFTIKxeaDWkfHv+c2ZnmQ+CywpzY
Cvm8g/Vr3LQPYZm2NxYD6ExSIN9Ad5b9UNsm5c0kb2gqjkbFm1n9gnTMzun4rBvP
Qb83VTqnXlzArQbGVkiZFG9IGBI5h6eiTeFZo7kqxbDljpOOyrsLtWM5nsdkbYrq
V9uDURIhL3kpY64rZsN+78WAEcsEowc0zi54kcn9JVirvYhtW9gsB4UqqzbuuPZl
p2lnaaoubcTJn7+F2xehZdeBFeU2tCQl6UMoLKQnWZZMNgZKyjlH1vAiOv7na7YM
ySZ4BwjOMKPtNfoOrHHWz2kEVJ1woOtlQ9CqxIbVPGcqfskEvULX9dYSVraB3h3r
qR1Dn2+0irel5du9CXQNKKtnGBkHKT5jPdLFRQFKW3iSWwiXOl7F7zwfhEDr4vsB
bd1rg9+jST4kQBTPnCEQBfU+M0SQF4zRWBdyMfTwfRe8H2HLgzuGEykTaFB6ba6d
I9HOIfR8e1TWZKfi8KME/cnxLQSpa7sNyQd/T5d9dBvrfz0E6vzIYzQvOAiEzFCE
0Px+xyYgWnT4z52AFOaI7rELVl6+0syQt50FKnzWBdlmxw5TOqCcMtM/ztRIl6fg
qjUvyRPlBVsYtZ9nkMWT+kRRd5lReWE/32/YjKEYJaNScfX1IfO/ZjDSR69gBjvp
LfdY0n+oqQF5rfvetTL8LA==
`protect END_PROTECTED
