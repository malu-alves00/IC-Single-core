`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vIbrE7IXJcqJ5FnyomrXr/R3ZAn28+SUZ1MGz8s0aJds4Yo4a7XhKpP7Xgqb4R3f
4GFed4/1S3eoBGhxswQdJsJ1t3qwD0UoqWgya1Qe2hDiEadZtFmPG8zmp2+b0wR3
aTMeCzs6B9drMVYXUtIahM1T4RH+CvPUwdTPhhN0pTEsI1m3l9rEx3ZtWYagZDj5
V+qoxteNmILxP33k+18Hfn1Td+zvDlp2ShGdMqca+JGh6gfeCcTyXgrqZvItsUjB
OQY9VmJahv8K1R6nFWTdU9Kp6l8naByArt5oOraBa356gvDc0xUItZhFHIuLpfxL
4Yjsn7IbusL63ZxBTFCgS2Amq7PuCTR8/FtRtPdf6crq8RrqGVC+8T7m08JuAVmj
T7RTEExWNIsCHDcqeg5JLETQN2eCJNh2ADM6OEfz9zoeVd7fh3DoFu8o0d69uOQp
9HHDpN7OHTDtS8aCmfTSLEDmp/JkPVtrgZ0sgASW8RwOpZdzZZjH39EHX8HC/Zkq
Hk0ZCEF25v0OqpB+8oEqFzXZ+wxIU5APX+kfzalg21pApiu+3+O8iK2zjtx7e8W5
kSM7zKpfuFXroxhw6bidN/mGqgLrT2LINyNxeFdjhkHWPtE6NWoNBmDbGDLCTZIo
TdeuDM/zH7q43AuPuJD2sauEK/y42cyAHw5uWNIC4bctNejTasUB095oOGv3tb3Q
wVqApdE+8bH6V3S6KI2Q6WT3NxBIpeCvKtMmYh05mAh44VYgdkA/F0W45zdQz7JO
rKFAVFM5P2PD50wcvtEc7pwsRYbb8xaYbWTJKKBwCA9ifvqo+WdvXSTC0TZxBLyZ
zncte/95F4HjsanuJV41v1X9OZc+eo0DDebG700jKLBbOteurV+OO6MFzjTdNaB2
FY4qbMN6GRUC9TfkK8fPnu/U8NfoV6twqw3OhopiwMGIVSPnXpnAPFs4gSXo/yJu
ZlAEM8QdpVTor9SqPabtjByMFMwDGxpuPrtzuiLs62QXgSnFMZrXDcEy11lLt8nV
FnPDcKRLjVOFNHjLJdjJY+oqSEWu+whxpp4lx0IBgzdHXgNCtFWPiaG8LwH8y72B
u48gsksHrTsfgduIE3wzVeGICrtvhSe0Joaj0JzocWreAqkKL50CfTsueZsIE6qx
bslWvIOdD+GNzFLoFvY99vnj5LoiJQ8xHmZMM4uKdMVxDVsERgMSziHMnXL8aAti
9oSlHuZyWC3UpGvXNM3LWVWR8oJjBqfZWMEjuwri9cph71kI2xwF6J75QGGGaHy6
6h0hDmEeoBAKCmq4DT92hH/hMJQhegJuDMuOOJrmLmOE+tYcsENoYcwAmp/6gHcd
tOqr3Z/uQCi5/Dl4zVO6e24w6Dqq8bqCyETEKQkhQ1Yw21/TJ05zhcbuAOQzRbAz
YJ/3hq65o+nAkvQA/99fWMeN1Lu/tdwHEdt044yXZN10HP7rM3FEP0ZavyUHfv89
AzKLbYEJ4Zpp+zWvMcZYuAvldtrUuUQSiW0QbngFxwFtrA7wmGO11j/DbkaFbglq
21fNTzBMTEnbPGrlu1mdBfKvcE1GJjXasSNqL/LHXT8rzv3Yqm48XY3tJPqLQ7ze
+n/LpQdhnOlliIr7oUV2tML8bUHElNS86XclRHJFwnkbYiTMRHkPT5MUkCIaKeVz
F+uxUziGOOvWhD63cOB1NLoSajckuf6w70NmILoLKRURRaE4OhsM2WBfTPxTjARX
XOXASYr3L/42kFZMOoNb75QXB+r+LvpPUz4Qk2cyTYk=
`protect END_PROTECTED
