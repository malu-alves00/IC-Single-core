`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hhfcTh+PsaLnonfH72he6XDrXvuD5kzJbKx+4n8SfIbXsRsYA1MflaWG6ca94RFK
LOKwqaxxbJfh47wBhwvv+lb9K+oWbWUtN8E80d673b37YVLU3lTdQQ/fobOZrTlU
nCPmzCZfIzQygBeo01kkXapuc2vr0/GJS/6ZyJcyIWQ/hmtW6Z+UeLSnHp/bepdT
zyI1RwctmKW/3Nz54XR3ODb/7dErkfj8btrjseSsO8fIcq+xg8aizGJ/nmfB/yGf
SnnM8jHXC1bZ05lJi1ncsOMl12eeg60G+rDhVzMCEFIK89GVqkJgpNdd33zjYRXR
EM4PETTbRb7tEh2fHHWksm3t0WQJ51Kno2LIOPJtuLIoNBK08w00pMXAZwa2pPZ1
/wuAFsJ0oRhheksYxrCAAYqynyUrIavOLXZDXfgaj36StCegYuhyLhePeOPySsgd
P6dww/e8Dbpzd4d/QDJOVr1xN4bgy6sivxfVqU8jE/jffuVtzt9lOHAN5h4LuoZ+
Jvzat2KDMeKc83fM3RqdZHFramnsprR+6za8pta6eI5gcCA1BvIyhGtAKP3GU9OE
K4lI8ETJYJqU9Vu0p+hBZDTGCBQFMYcFmDFY2fp9gZmIR4rEFiYiEAwBqJj5ACzG
sQaFmAa5oJBRy6+UwB4769UnMoT3nJCIWDMew5IVmma0vXpY7ivmkm8XlBOMaA7+
rRxNicR1Ixwv4t3OWTxBPyKwBOfWYCZM0F9VDpru5mfY0iuCzMgWJ0Rdd4MBIMra
5gDt/JhICD6S8Dr9tfs7lmOGjdAfiTJsiJWm0Rj9Ky08rdZUfIriiDX7lZ4X0J46
tOXDpHA6v7Sne3nz+8VbR4OVJvWioRNBMKZRFZkebIJAffUEnhuchdZ03Khxz8TF
4nakfmSw7QKHtlojVlyPYqyrv51il/hVhg4Z0S2pDKcr+BmOH/1sjkJC/vMskZIA
39zJWSrfyJIyFyZWVNTNRr9uPpvRKLixZ2YbItk21yuMhiRyjUOgFLtZulWjRkAG
IJG8hDpu/5qO4nx/NNPRIQUWZuSWq9n/wp+9Ettw6Eza1e+mEC9RyGKkML3aCmp9
113ej1yuH6hcuKK8AmL+0p97BEQ3UF0QXXtlSOPiCtKMn7RpxzaBWjxS4hq+23ra
`protect END_PROTECTED
