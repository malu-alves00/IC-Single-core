`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
I0RvURw9IV9K8KrD+kfscg5Qm2C5X8e+lsWTxu6TIiLp3tkBnRRCpNkqtU5arGNc
DkMzuRLieOq1iGRYQtvfJdyVLnC3RqMxBeoNpw/ziLOAiSy6JsCiUaZaA9QRWGet
zBDZPSwf9tz3nYznJPfb6gYzx7KrW/GlJra/sT3t7jv81YzSSH4wgwqMYjhBLboy
5/85WUAImwnF1q80zenETglrEXt9p8wPv3n/ZH4MMjYFkNWhlcJYn5JXk8ON7s1H
7dnjW/YqIxI/tqERp+r90wBcCRBuN4Kc1m2GSFntRfUZiSpDRLGiSGQXpjo2tNav
zplGS2iIrau0EN6oV5uPRikURO8/zwg4+kWRT55B8DUd4c4lr5dFjjwPwY33U+5t
UoR7MB3Y7JcoATULIPhoCaszlBMFgcTjRmrm7M+IYvqhDvwHk8+g69GJe37L62Vc
8LxyPWGfOIuP50Dn9HVBq0ZxXfgeb+mopO4JzGsEfKbARfRXiX73FnlUiK2x/KPE
fPGYuoHw/LXjNIPUdxMn2i9z4B24Vw4uwb47JZFQHL2B6WhNeQkUdrlK1Qwqoat5
ENT7Om7/MRJ/f9kYfGFS65ehs5lmxh4Fq0TU4XRGWHYPDElrr8445g0wvUJk1Nnx
HU+aoOKVAIIu6BTgzSYgVqS3xTW/7V8egT2UA20Rndx7xBD8VwRznc24UufZ6Um3
Tlje+4uLd/ZFZSpHUxXlSr050/o8kj6DyvtFYAyIe9vwGXqgS3EiCHobd27nQLGO
DpZmK5pK+YwwcpfLZ4gjql5W7S+sF3vjbaTkyKy8irotfoHSsOhSQmgjo3iUFGHu
eckUfK5Um9sb7UO4ga1DRclELJPywlTOtFZzanElqG3hqa8icKm+5/rjf/RPwATd
8fLOndLqextAsX/Oo+oJ5xb+H/Bxb6QzSL8+/mP0b98=
`protect END_PROTECTED
