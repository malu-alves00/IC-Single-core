`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xybO/UKCyuZGf8dJOkUJoNwwwfG9byfuUfZ2JVMXTf1zBUFFNZQwP34SYELPc+16
0jryiscDXVrZsQLdlzYO60aQpNuVntjfgifBFXia5Tq0/NSVk8JlGt+PyHcwdm/s
TptBdJV4MEBJfXYRfP5v5DzZrkBZVQEap5lERNb5rqV8WTRDL8hnMr3Gc4VF2F0B
Imd6bjOv2nIDWBE9BDD23zGy4GoGd/gg1JYHgFryWLwouWF6ierXKLu2enPPGg5D
Wccu7+CVQIF0nh1cm4CXjp7SZ5Rtzljityl/9OGIW9uJoPU2/cJKeh1GULZ8CqWi
JZ6Rg/q+c7T3OGFi7KIBJTvqG4Ce6XVBOK/7+Ue416ygE+s8U159IC5ZCzVvLoj+
hNPu7ptVC5tXoaHNmIt6kqAQQ4+GK2D1UODbvaw+HkWtlHOGj0yfOC0YHHsXyA+j
LVvC8ueiw3KBgmLwR+Av6qnQTvgvh5Bi74BfIxySq3tOA+049p5DeYF8FzfkDPq1
FhKVdZMfB/1F0cSh9d9AcB8Lbh7gVMz8XwKIBqjJCjWnVZUqwBDBQsFka64tv0rM
HoVnyQFCew1Ua4nkCwSrVtvrZ9voH2XUrylizPdsUMroIh03Y3WfscFi3SMgtHOx
9bpkV/tEul1NEE0RjV3IGdrekOaYTIIskNV8zzbl1hTWPtdnmNwwM9jGvBOIOCr7
ms15eWm3mrRAYQhBPauYjyfGJNGvJLnGK9x1jS05qH1s2EMrmK/7XtSnT0c4//Cg
PYmW+MIey+PfKC30ZgxjuYIF1yElCZdjX/xx0VEVVL5W0/izSj4e0i49WG+3QVPH
uF7O9CBoa4BTJkKx3F+pSWAy61ZxgIUXd8VQZtNP8UJllmpLuCJujHR4pI6vGlb5
at9qVktz3LSFtKZD/5Up44C9GdDFc65IyT7yB4dgtbW84Q00UEZh2LzGJeXETfLY
AWemb4tTOTttRHpklrNww9bMXNQk6XSWO2UWtUS4+hRI47WBUPXkXgbtiE93MOwQ
NmNeBO2F34lr9ij8ooAafqK/nVtoPcNBE/NUYD/WjU8O3tRMg5MhQLjA4+rOcYt2
b9EmP5d7nD9Q9BBvbanWHEugq4mLR4LN4/mA3G5nsBo7bqzSf9Isbg9T/r8nN7Nd
k33qbHU6C617YOe878iF/GXhKNR5m6QRxBvPpQh5LvewjSul/CBkb8728V7qT6qK
46H2NQOm+Etbb200hbfEqF42VJ0C3CPuHt6AJojJDUxNX34lYCNjyZRP707PML4M
PkvFcu0xaGEqIKNRYmf84Z8NW03ly/KyunOF9+QPnPxIyfwmVKmnLGIB76uj0gVN
1md3eSZFUHCjMHJLeEOZV1T5ZHO+EruuiLwmhuttGZ4XGBU43Wf/ntOKVOJCYAnr
8xzUzj6oaV8KBMlErHXcEoyep+NcCjLB+TPDaWm6TLpK+K3Q1h5lRoB/obyMcxEf
zjdDxQoLJLKr5LzlNGutNIsikQHAXhl59gujIR97eodapYSKb8jRIxC2ml8KC+zA
AnfrTk9RkeZuO2SuQrTSNgOrkv6QDjgMOHJI7yjDC+9SqSjUS/shmYE0dmDIl19u
1UTB0IndVFvRIh09bqHibsqbtjIlMRpKnqTzkX7eRIH/NqEALFOFBLL17HI0LN0O
iaRURZuqlP9qgpSxeFt90bdb+G8ZzaBjZOObhWRGEudKEO6Y7XMqBG+sQ4AnmHHw
+RWDbdYqFL0z0RkMjVEkpHlr3Awaz0FYWWgDSjwQ+nDqCCxPeEse/N4NAAFusXxK
N6QSVmkBharazd8s3Kd9Ee70zIZuntOnqfYoOxSMT8uqXyzWPJ2OXfJ3y5XK7RCk
n/ev4fdoHiVkka+XhgLAcwe0vCwkFZJDll4qlfTfb6PxWeFjW5QGhspg1FyMudWa
OpA/ErOs5NJW++m6x3asl8GlEolQEipLu6IypY2tEYr2qFR1uACfyfNNX/qLRLCJ
m/PpvlmSpjLGnXHDtLhKyLwtjrPXowf3CjpfnaYE1IqjAYWm+LFw96ui+QUo6pcM
v+O9DGYw+s6DHFCjV8LLCrDyKvVEpWGBKssxWS4VFSuoqqz2GSSJvkgoWrRajr5+
deMlH8aTwj/4Hyz8YHGshYb0TZIVbrmr1GWu9lmpVpqiHqehcEWXQQTxFqAnSgFd
vjVr0s+yWyV3mpX9MEursvbQFhJW0b8Hgad+6Lqv3KSXcMpaWANhDZSQx4vmfAJh
E/NWJMDEaMc52Of3gvRsvIXlUtqibB+j03PFuA4rJ+cOW4RFN5TFHvZyB+TJpM3A
n9m9dJBVa7KTlIE57frpC3XjLp6LiReWPiMQ4bQR8MQ=
`protect END_PROTECTED
