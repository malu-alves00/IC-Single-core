`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lNHemouegVgh+ikVquusFOTslM3o0PnGMs82Wea06LpV1kZ1YlYXLXfDyTCRmiG4
sNFS3Q7INZre0Jh5O21LkJNd8ddfpWTHokOq76BMMIWk2FkTyYPhqyJ9pqXhOJiU
qykDCg4OXThxHzbVud+rgT8HgzCXyEE2BgNWeF3HQjqAjsbw6ge9QZ+yc5J9jmn2
IKo7oBwWMgGhd03YQ+G8JpONwbOCar2swhrwM1HL9wrZWADlXv9LoV5OM+Hw95y2
RzBrfE4I/jXLkvjoiU1caRk4Fd4WOfCTvFjJYbNNB2Xehpn/6Z1nUOUt3mU+c3Mm
QegQ2G9ghn+06cnMgHZHWCfMAj3eJHKUNAjtt0ahdDOSUta8HjJpD+9F6YCo58+M
GqVIrzgRrE8DqaIY23G3HI5a6pIOdryDXPM9PobfY661rtVTfbwm0jcGZUt581s7
gUtJTFRd85atDvdTBRYZ2exODGT16y5sYKcaHmxBs1LKWe3WCKgJ6UztUbIkRyTw
JFGrfegmCg2ZvbUD5ldl+1ShLVnbEEF5d3O+2qTQKvyzNUrYa/eH+e7rYNKkMcU9
2UP8s0vgXkg54JMmHfIMY9/CwfFa/5z6GlJaFVlfmid2+enPqRpsJun57dA456fH
Cnvpz1RiqWPKnd+DmiFCAmx0CT+bKea6qtHANX058HCai578oMUVyVGqoNmzOaZM
g8ZIiTopkf6JV6WSYkjcBN7j8edw8NRcfeQViGMBHAMny3eXFuVl3253MaGE94iL
irnEXZI2ZjthqqOyx+kcFVsFRWeOYaEnzZ6XXW1PG36vsLc5kH+QyonqPbuKYWMH
LUePCgEulSc4sBuhtGfcQZ5MrCdi86iyeE84igTtBUDvMjBMU26c6/CLUHANMCiV
JV8qeUDu1kA97z0UPzc7cqJ6ek2V/JSmOCiKkofdbNa5XUqy6pOywwfnC9RszzVn
WsyUFheNdG81oQ9QNkCcAOUjf72R+QGQiEVDeSJ7yiOaK/CSW7VxPKsYFGhBPmuf
g0OacuBppVBPpqy+BAUc3R84YpsrqB9FVYxYKUCgpXihbSH35uDYqupAMZvpORoj
7eBWhx7h9S9LxNfUlgA4y0WIf0JHVpjerhJJrhp0gVJIllcYXLMLpUEjZ0ZuZ2RS
TWOWrdzlu8tht4TPtXNsDi05FhugWpRSZpt01Hr9RUHP0MX5cZfkkrrYItNatc9K
l+0crZsGlBTxMS4lFOeRZ8uv0JUFcJs2qIVfiGv+gaA83ceV8A1QebFy7vtjnhxu
jugjLUXdgvdr7odKvlJs3x2yyQdkNXYklU6kfn9mjJaR1MgcCmlKfZch5KgrQbwr
ybKpjUyLaTgGWOE3JpBEdSElitJJkRmD+vj8xTTufMigOTaNBWxmMZs4wyLTnuE9
kF0N4U1F4OJydfpQdlnhkqzyML22clCjDuht8EZF0JYQ/Q5cPGtRpySxtzGvMCFT
82tMzuIEo10Twi5AC2HtURgWy0a5q3Kob6zP1m/bSHG7dqHPmDYDzMaiUo9YwsJh
6W0NAgkdGDfjNRGe9FeS7I8+gA/Q98AJ3kbJkhEEbRVJBL7xmLnSN+8XHVNcYytb
ezrWaG65d7wZjXobBau5sbVDg3xUJ2oqwtCWwbO9mebvZ9kp9IS3fkay1PdEOUL3
YWaVeO+tLdYz6P577rgoDhCyv8bMF03KXQjlP6plUGjQx1pOqZHWgIGGqf8eyif9
GlnoAxtXCfnutqsOL+HAvL9DannT4S3yZ3zBA7WYAcd92bHb065CMBJsYffAkyLp
rfPJz/lnNAv9KW5Ai6axaQd3Zn8XeVCTmR7M4QfgaBAQoc5Ki+ULGnwcPOfk0+P0
WWaaeuC/59gDE8eSSdah3mvMXTYSNsmemF6sEB56wTwfWftlVQyPXzxWbuCUIIgi
r2Wocx2i7RmEJzN/5Oso6Q==
`protect END_PROTECTED
