`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1t8MV0TiKDnXOSmODD3wOc+d3ZEG7ZkT0hcI4DTntlQP/nL5xU2+wEc7H7RCtx+6
7oKiABgSswAejIsmjcRfGtnOXfJYjJqNQZecePFvzg/eOpnDURuvjBvqeH+gHECj
jXq6x2Fh/6FsywjeuRXKA1Lh/Ou4R8OKoz8NXhmXzUwc7qipYgBQd8w6heCog9Am
3rFAjYRhfBlqHVvOwQEDOmTNyTv3a9QqkPUdNiGENRJStE2OcHqJFX4x/orWTfvo
CiusmytsKAulUUkxqfuMDjQme2g3UIjR/JeWhxUduL03QkqsMnmRgJA56smQNLjI
Lkb3xsHNw/T2Ssmi1aP4Fh62B87IGqZA05B/YwP3xgOfcBvSubbRSPqrirtSpuFt
DdaAbBPpDHFAGZlOnHImC48jG2/vcZNI8JwVPay7LF3JZoz9TaUx6IT4Nxf7jxaR
VzpqYatbVp/BGZrP6RK1dudOEMiOFnULd1RzOJAlB92A5o2ZcDjTwaq+BSNSLw9Z
E/7e+eAB/zMHrUTTEQZgNylkbS5s9NFZOvMO9qnbXFS5fAuJrvlmnvAiP8hGBvq+
O+bfNCSKZWrnSu8luuynKtnfISm1ElywtkHcSbkMSrVWzMe0qfJX05CYipR8nPdE
D3arIhChaT86IibVvFBdEriAlpF21ZZ/In7RfbxVU5pQxGoVIOhYqZTkErduUk8c
Y++lS0XOM0s5KaoN4m8gO772KPpVjfypjWzv9M/2aMzWgpAK7uJ2oSLl1WaYXggk
NfIVkloSrI6lQfodqa4PyyU5aYwsalozCk4d1+IoyKuXCFyTE1jNQPtG97ULfCz7
Nejpv6kothcK+a6+5/7u69Ove+ypysG0wTHh+a+a3ghJt4hrIeaQLSnR5sCIsI9o
OzldOuCF5W0VPWAcPBavsGWRuPfNh8AecVzmaEKMaa0PU9LG2Dt8yaavFIWJKxn/
qvA2PS19Wdj8z4qkNrl68L0RX/c1Evc7XFiQuHk6YbZOy+ZhhnwDL+Ncc4PmEBfI
syhHnoetCn6qp+NnpIfRXB6pcSn9eqsCoBops8Q0meEazfAklHwIrsFODjRhMxSK
enNiotvoB8ag7/0Gcw9BEOuOS1ziUknpTRMZ9BYIuEBH0tKv36+j98HKEDPKz/U7
CqTfQGEzLKGzuikxiUkF7IupIGCKgvTZsbREzHCDetkHYHiGDp6xn7yz1r6UsJCG
eM+vKzVsKofzt8/MiOvgxL5hkT5GggSjAZq8kUmaFSjRCsE4D4VPJKjDEMBYzSBM
ZWndB+sKEd/fyj+clu42BZ6JI969/P50zhGDU2pXP3csq9JQuSYPVbRLq71kAdl9
9LuylnJh8yx0DEFG3+dU6drUaoITwC045D7HKEFh6PNcC1wdq66elQjj4w9ZtWs5
Lk+lBRpoovGBGeJrMb4r/beIJoppu3sI5gs1mGeAZMBVplrkqOmQNFdP7fTgaz4V
avGLbY6SA6cqWCoXWyHTyXbAiSL+Khd5/+6gJSb2xTOau00g6QldV0LmMTbnMgwp
hQRwbQj7Jj9UXqL3KmpsPfc2M0UQgmcQ2d/IV4MmNFg8oAbt2OICEgc0K3w4qMhf
`protect END_PROTECTED
