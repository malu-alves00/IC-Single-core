`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EBA1FIMbuR+0rMddLHuqCbsX0gxUTxjASGBTy9mm0S6FKIRZucQDkxAgppCgj4Vq
wYDF816sAi48szDWDXYGdOdOQ3DebQP2IuTLLJVqLJUEUL1YLop+xfch9rBauc9E
1nto1V+jZhJ0tWLQsPH3NkSMo0OuGpUWzwSU9etIXgbNR5FyGq73HwynzzxqIeB3
ZVm0Q1XCEsel6EytekHevatzOys2yi73NfqkE6Bq4FjADs5BX9CHqc8ACgg6gNcL
7iVMSFsOlgmcFr1ncNF48iwZwwl0aqjGt4hlN3zJbUcD1I0SCkjz1tbtZoPnpvMP
ER+pg6w1ukBtQD32YOaklseHMbHSy4xEuhuqcZw6qLXercRP5oywkeuDfy+YirNR
L3y/9Rsmp7ait4aF9TbreMROBfjmeVNKFnggphlhxNCoOOV0ZE+yhZSBTmmZZ/lC
F0G3pdgq8vEyPMB7QZwpBxSGLrarPBd53k6yxObk7Wh4VkTu4ZVk1PPmBP/PV41C
QvIbWEBEPY4JsyWzcEYxXV1yE7VaA/034UGvd9l3+a+aJTDONVgipddj9ARTEBbf
flcbPeIFZc2xERdb+Y8mFvjfYBU6EDWLVNE255VsKa3ArGg9gkxoAY5J8OqP5zjF
oSBYhQQ2DkmXnRfj1gCv3NVTx9crhv+C30pdTZqY9em19pNXkSzw6DkDkqFyDOUd
bD/IrljQCajNlxT9S5mmDhS7Qxkw4wrPrDhIQydFnGiFUBq31kc32hj2BONqj++5
w+atqPmsViuMawRQSf/Gx7EDRg3di9tkNnEmDH67tDm+Mw6dWPZsZ1Z/E49RHztA
wTTk+9abeghmGF5hdwaQnHcKi14TVzjUyczelxRl/K8RuhnDgHy94M8qM5r/XJmm
eKVDDKOX2X5bMu/U6R0p18xwTWMUmJA7/3LTemEXUMlVQ11sLYPyiAVlQCRuKLgv
Bs3wcf0zgJw8RPDQsIggLARlYDIc5IckZirST2b/vLJwdZ/2K5tsGbngYvwZ+uws
SD7yEMlfmF8r+70MK5mOr/Z/ExGSaZczVrfn4da8x0KSAgTZc6mZwhITgZCkRUEs
ScwlmnVpva0rFjOtNOh0Zvw+GcCf6uYRrH0KWb92PK5GQXaod1wjVA3Ima6dGVLI
svaeIPlXt+PSfnCFgZP6nFHkWqDplWZSjHNH+hYbP5zuaRTqJ6T/FFDOPzlxCBHx
q4HsPODXtpxildHaENUMXjdok92CVtePQ0JP0RijZAg7Q2SzFSlNMCe9WB63fs9h
cOV8JI4krqipw09MSgLwwAcM6/1UE4WfRHlkG/2fdFx8jahmz7qPSgDM3IHrDiHJ
TLpY5odM2oatIoNfDdMp1/GPhHlEaxjPQUjDh02wrJqpylYhsDUbkJZuzjxO5rm3
Qw/Br60h86hqlwLqeVaZ+khV7Ytf7vJSar7vgzCrJmM7O/fdRC5byfs1kxI+F91+
Gnb7KzQPHesF1p7E2Wnsrblt4pN2O8k93tr4bSAiEFhsjjijTzBPHxTYnZk7y2Vz
MAxEjnvHm6RC7/zwCuPxJBqkHEdNkaFq/9iMI2a2WbSq2DVryD/kwDaBDYYES94O
ZeLXbhRNwhxQdrYUq7RBUTHRlPdTs1esqA+8/SdCQZSYaRNro02e+kG4inYtWb28
mmm+RwlMq9LgIlCjIQeEK0As4GMiaWVMQa9uY7B5Y9WXoxUXhtlR/28RrLOG6kAi
e8POT44KXVWjGkqiIj5up7ZGNlvNmDWAUF+prFsLGYKOx8MsRIPJcB1ASE4iaoeI
lTkGDTvhJNTwo1r1VfjVNOsGm1Tn7s83jxBQMAZY2v4KtZ2DZGbYmoY6RjqqddZD
mTibDT/EtfMyg6w7u5wGcgI5lcR2+MBYrMPLFquWnVBH5JmooMJCaAnxf3bVdxxw
1uhxYZSKs5laSUng54+oOKOjd7TTUoIIUmwGT5/WfDejee501OLijYq1Sj2c7wzW
C0dzHPK9FBFYDVtyvSRtvFeOgD0cl0sBxsERx+BGed9sCEfYFj/8YR1lhlFfcFwm
pkeN+rSz+o4bkMrEyYYmm/lvZ7qrDDdzuxkSvVlSBZ7up9camWFzz6g7vepkk0c/
4f/twgemPkU18oCTFnqGhHgmNPr8EqGesXVsBNB2Cq0G/HrItVSOB4ZM+IhwEO7G
I++3w3kAWtYAYNabfNyZSf5byBkKzelyY0wUa2yN//OV/G4kBPPXo7kt3rNeuDpR
AiCsaVh/xjlE9D3HmVDPK/wOLIlzOZEcmLkNcjJ3hEuKxvNHvJrM6q9FV+NwcCil
u8TFmoKNkxMWsbqz/tZLXKaub85V15lPWkACAfkLWUjDXDBzSDhQ19isT8lW9MMZ
IaTcgBKDRZC2LyDNAYKHtqxhYzuU9DKqzXAkx4fOfMJDqI7BK33OC4d2rgtICcLN
/QWPQi15qbShFM7B6mOtx0h84dorKn1b9xuzi6TbVBHITY8DrVNzt5ACC390YP7d
TbkvbxSnAQYpRiSNTxRrl7naDVkl3rL4qhYQsFmkqJ2M5XEvxra4ioUk0p+0s369
mqHvAQ2m9oiiVlDix8bjNb/SAlq/H5cPgQX33ER1HcP1NxfZZPNIQ6X1RU4Ybjrf
gBC0VIMwhYvsen8rxYYJoZlx5YlsoGXiO9FDzrZ0vmc4Df5SHXez2w/u7OUryAIs
iSzEr1vWNaeQfIJloZPU012yXf621PQEf8U4r9ZpKOOrXmmooVVMEJimiMaiT5CJ
9YqjU7Qz1jN+BgUPlAHSapaYa4a0ob6T+A5wbewjd1JqTeNI+E0FK8gr5ChOYSdr
ihtCsx3qacFX3BFKhUoJJ3M+8TYXaV18d5N8wA9efi2lny9DWrp3kkkxs1J2N9+L
68ZkJwpCYIJsiliKhto7ARLYyRHaGWgYkzPPGskhLBviRF/vlEr0591IF8mhBlN1
eZYqLxTE6W//klE6eRCr8cTnrA2PQVnuQSOhH0ktkQ1Xgz0m4vJUAX7WdJW9jqn0
BjZlIyNZb+2KRfn+L1FurGOrr/QQ/pimQhA488PXgU+2edqj8RcYDAQYiT4fQRTS
dDzOkWxUSrH7eQN8beBs8Rld6o5wZ2qSpQkUEv+FSGqdF+EmNegcrIw4Aac5aIhG
GLJNliv+kuS8vmf3zVpuYGDUbxEIrE1YD53PLr1UlzhI8u/b3C9+ee/R224pORQz
XU6FB2i+RuFTkVQlrBZDjsXZY+VR1qQ7fDGcpFT/06xBEVJjbThssi7hPS86TMWn
O0i2O+jmCoEjrvOy6VEYDUDgSrNR5frwNAuERcThzak/MD0+JcymS9BX7by0ZUH/
LDRZG9560nPRvEz4Qd0jPEN/H+Z+rvbwZT2BWAy2a73Xy4U8yGRsYIWc/5/6DYho
3dbnDGtA4PLa+51s5/SWAFlUyCZ+8kYLBruqDmQOjF2u//grPsK08x2GudF0UH8r
1RWn61ObDM2w0RFEo9LjKx0juqIOZWlumUWUKY1fh8A9fQOxoYaFWROsdo7qJnb1
ORq8rslbkt4FZifLj0L8GqIPWhIWKFcdYuR4Krt+at6TxTPLp6MIRpIkXtsBL95j
pZqwaJ1EOUlerjslcxNsRcpZ+xSXrJyboQuFZMPKeQS1BJVHXnBTHwmWpIlH8l/6
xgIhJaF9ysi6Hfwv2SY08oNsp8iOXwWmVAaWW1ddoDuukFPo1IkrQrB8AbBNkHj1
O8qzZoVBEwPZ14OsGc4SpEz/MIviGXZqmXY9SylN2BMVnaUxgZzj8QHKfrJSWzoQ
NshQRpPSCw7o9C0Ed1yULbB0vBsJ81pFFQfsWG3WTTQdkSAlqqYMJ52asnA+qYoj
Q6yV1H7i5m40jM9dUL3kiMjRubHtI5brLZs/ndGGasCPAAAQHHzxued+5aQPQ0iX
a1vLUH3AWn9bRQe39ljwHVgVpbxRvAQrB7BmeU5foYoOECcdyN0vhrhP7XlEL01+
93cS/ZfPLKsrIMhv2EoPfankH5H4z2EhXxaC0+LKP1uenb9YpwbHXzum2B1Tvmnh
/hQG77I6kBfmo5/oaFYVBkE/aDmKDpe9XLIB2wZV5zDmRZ3ttyHU7x1M1rvDOEH3
SYPZmsCuXKPLqNQ0c95IzEf1UG5CO1TZBxJtVpPr1j9cYbIKGQ030/xp8uO3QIoP
Ae1cuBP3eFDlQt1BRVDjq55GqhaBhoplEdfxj77L3A9TXbQDAL7CrwRql+ZOVL/d
Hc+JgoHqWW0XE5AFUGTXcQQUBWkoabt0WpZ8wRTOsr26LxD3E9tgoOsluCeafXFT
TgAJqWB13GkZT613loZsZlOB9VzV0Ff7KNPfrW+mTeL9twRQiVp6ONuJ6VPY0cOE
hiC/mY9L91s85BZvmWCwmuP26tt5ACCPbJ56WafkQWDO3I6VBWYR8HWLM8M94Zlv
dkhnbJ+l0+VgeQ1HEv8utPvDfi3lWWuHKdsrsgMad+bZLaixfOKq0IfemXjjedpg
ck/mDesbg69iaawBxyDrzJHmRveBs4MFhKCdI36AYg0MSutGPBjAob8y40OWw6wE
zRh2XpAAtAHK5SzAqINdQybtt4ltTIl+JFV7b+2i/SuC+fR+OzOGrkZiNz5oStpE
Ay2GOEwMGbstg6T4tEP4jhkbVBfJgPp07wZX4vg8F3nSitXZVKnPPR5byb5XGp78
Yrb49Ur2Rs0YrOi+8wVmUpdPBYYWl0Nd7UBuSyV8DFOiQFE28s1i0qKZa/pe1Ytb
SxFMekWtHSMS928MT/oqcKRJk8yrgOzgzw10Musnl/XQUNSRsp+QINmUzx/t1HDx
QwfWhLNYp4xwiwJ+UUbNnWCeKOcXN4iZsQyAWTXv86Aoh7U4Ji0aBkiUFlWBGm8F
V9jWmlKEtsU37Nfshxq9cQc0yUZYmcjUhlXs8ENsl9m1gdIq7khnCeWTxkI74j6y
PI5QKi/boq7dvvaY3XkJPA+6vE9KeWN1R1p+kVt1ZZNuIbeEf+w1nABjfbDE7Z+D
RdSQXxW5E5GGonb5ZJUeWskqC0PtSCmQ5hYa3P96IKHC3Qqzky52FFMH1wp38vxP
gQZi6zlMkX1KAI2eI6+zbCSNji6ZPyauhkLvshNZy0fQXB7x0coXrGj6quix4h3n
YDBnHymc7kDp3JhEeqIUeAiNavrlCRTma5cgZ7rnv8lxGQ6pIYIQU1kKnHCPHxGA
cS2zHBs3Ntny0PMTjNNRnX9nqUEKjFKGoquqdp4kFItXvoql8upqHCzmrdgO3+sm
F50FHu0G/RW2cDxJ1q/vZDJzDqJrFZMPRkjrkK2cS2TQXX4rgf51pG1cE+k6qvsl
p/OC5/Ot+RuB2Ji6DaHpd5HtWnnzuhFONen9QBywlwXmoYuyhpNS7uP5n709vi0h
4vmuxBBEN5A7Ipd47EDpSFa+tc/t2Jom8YLp2fklE8SMTJ6PSFo3WaCjX1LEN4OA
yGD9bsWoWtrXa4HGsyU9RSfk1FAMGiMG5L+Yqf3Nzx/abtPGHvJfVa/ZANWqxcNG
szFV/Evw9L4DZjmmUJt3VmY+kxJS2DobFkFeYEy2FBchum24tJDqej7DoUQmbtsq
guOriLeyyXGhQYVxHY8np5hBnQg5U+CtHd0AeftBJVKie0717AKK/aO46kX+t/yR
BR81GvqP/EOcqLnPug6OAoXBNfGTtdb3EAOxQMQhNSWSdu/g5ljBUQ0uuhrcH1PI
HsIpT61mYpW2cTI7tEGw7LM7PE4d0t3BXp/7lpYrt+gZuhj+ItxmH8oYhBAju7WJ
rHJWvfRLuOi4/LF1EX9p4O3GNE8P7x/2B0eu/r56yx9VX6nKeAFc1wbmVl7Zqqdk
7plaxyhvncdCYZ0UV7QwkFPXQFdbHixC3GWff35LqCMl4hUfGpxLcart1gxTA/cK
2WMU5RcZpcAsQyhXO+QL+Pjlu3VWtt7ZQqYRb1R+tVqBkJxwrN9m/y9OhkZbHogt
ab2Ek/E2joeV2W4lugCHRAFVPnfIFpaMA1RkupySAQi1g1+nTk+hAJ25I4A7d4yO
CtonSrdPAple/w/j6ZgBzl6F1fEixm+BP/BctZUs8fOGVrII/O87vTP19+Qef3eY
kFEDNbDmIHz5oFsZwJ9jeu02VS8P0TB9nIcVo9NmT9i3I+3lQBJrSlhGd5F3cCJD
M+CF4WyDMlTU7wjo/MLU59zogs1cVsikjSAJ8SB3AFeCFLLdSDdr8CaLnDXErcga
XoUpe5NWl5LJbo/usye7KWMeemm+qpEfvNVchM32bWuqYAt09Opt1og5xdKeXXeS
3mReS5dUIQ5H4cfmxaMerLIF2rjJqLogmerZCyc0v0rshBGMbOUWDMdezRBdfjAE
GkG4LU+56HJnsNHjtsgUd3CwbzoCK/KXw56mJmGQzJxYzlsXc9GyT0gDeGlWPI/D
zQQnc1/h2U6vjNINNSLBN/UlOIFF7Andn515wxz8oC2K1ws8+WIPuUpqBTlegU0Z
MxAbIKQyqNo129U9mNE33thd5t2Snn4kCXvj8ranYzTzuXBu48kjGa8DCbkE0Qc/
tltRKzyFCS4tpB1vmm05PEgPtC4esPdZJ8Vp6JtqzDUtj5GmXWmi1CXDQhqsX6Jq
2BDDpSgmm7hzJs689MKdonHzNdJ+NwVG/iU+vYLITOLFyU5C6PvG21f4mmKbDLag
2Kwc8lYf26eD92mmPSjfrwkyfRXcB/4Z542oP4bHWV+aZxO7LeJxTpkRPnHHSQX7
klDZ9TZorUZZKWX8ixFMXjLFSTc/FMELjTQ4nR+UytT1QUijGcw8hoGe4SPJahC+
4d7p04nQQT/TsHHkgAN9K2BcCsOAigN1d40TboB9NnVXa6ArC7M7WjuQzasnLwlv
V2vjljsItMkSEmxTDWy94RGSjkxSpgxIoi6JeglaNcrGdz2zGyQEvPJN3MOmEyMo
85QoKLMmimm+/lqNEupvX2TzRvxq4kx20A6fAuRwSlT5qsVuZaCE2PG3QWLKfiYs
45YCP//I8RQfFQc19ttph7QsGiVPIeA4wSwfiKTLo6ESm8MQwxGoGSkMlYzpxI9O
pa5dlqWv2xuy2q6bjIwNG+LFOWpa/Ryoq4p1xnONr2zN9MdH2vYVQK+HSX56jSvm
/W+ZX19L9Glb6SCMbCSQH8Q4f1JfmHnFBdiHlbEJ7nbyYtCf0U1x00/qcepYg5Pd
MRiCipiHL2MtKA/4wG1KpJxisoz1hCGXvRq7P5ovsZGArBHhwQDEtf9GcdhIVjXx
4RJrAA8fAPShHdfwpx6Qc5YcSMufTvqhJNrrNjZw96vBCgjSw/vqggoebzlgP2rJ
kov5LJqD/dEebXMLxjGA2Cl9H+A6tFIZFkadB+ddqx3LLYxQIXJ1wjSSRHQ1fHYZ
bnh+aqJyXpBYVuxN5qOI4cuaoSsKRAwBXnrhccY45sj6K/xUfGOlQVgfGcp2JsF1
0m8X5+AC20k8ZkbVSKu0n0BqVjt4r+7CQUQEuQTky0TfEhsOhYHC6TFz7QtOanjc
gUTk1NNN9AaCXDlZQlcB+DME7GBZwmA8zIK1LQOTlrDtC0uFR1CJ6JPmP4PliSaf
9T7X8eFnXngYhDOKmqT0GXaiDo2FZABL/c/qVs9h+tDF27Mqx9F+Kzg1V8GkmhWh
gNZ4y8Vsfhh4Y5JmGejZ5g9MkFEh72tnlBpiomwFWHSgNVslCcQWmqn7t0MwBpfo
jHGXty55SHRv9WnSCRh2RAKV1sgc9/pV34jbLAqSNjfQ7Wd6sh64AXp4JPnLaWis
WEw4ciDmZxkpGcxC1+lFrYG1sLQFVdssylx/nTO80aOQtDOtBDUdiQOLy3O4ct+F
00lZ6WVsid2B32tbO+mUq26kVnOdTzkFJGhVpBUmfWXZz25tfO4eVle3QsygZlaF
d3duIa6hRSfbxHUdp8wI2TQK3vTodbMN/sfmOtraSh/ilJwyN3y60A0nVJFSYOS8
79p6e93xs+qsnvJEXkOaOTOhOmfr3LupT/yH1iZI15+Qa7VcWbMMJ4/Q0Y65AMwl
d0Xp0P7td6zyFCUXXc6VSIO1QnpqdvLTYwDZ8XT4VFYDKefJX4Wede7X3kk5Qwjg
nY7Ckt3BnssMtRHBIEeRag1d/2kbDn7HrbdmF2ldtI9YnGmyD+2WgU1lJIcce2nn
uwgA1058jQj6Zo6GLrha5NqJB9nADIyGkAT8KIQ4Kb+qGIOMX2HTxmeU6CjjaKMU
YPxZR4mrFfXr516d1vTrPUyBppnuIwPkjBBx2OkVFXcOVbVTHJArAe6zBwJ7jfwu
AUBDIWxc8WHtcQyiV72+HHScvRjKwStdVAQdOn4WBY5BYH+m4DJbRwO+/kA1zkg7
42tuVz4XsnBWdy1X3QQiGqwnxLYh98vWvxAAvPdH8TDxTcKRS+5JQxoL1qdvsYz1
qrK7KvIPU8U2G2qZ3ErIRvcAFJhbwcMS/nrZwLLWyU4s9FcgH4IyUhzvOMJLaVGk
uMKe0xz8CYi2BoA5qBhgfp0i8GEHOcQJXmiDfY/YNO0vcUUyWXwr5uIaplvt3ek1
0upZU84MbnKat+p7RopR9bV5GWrVBhK9CO07TGj8dRYVqO3e5Q1bS8YWv34eKzkm
bf+cnEj01BZrgaEMvV6/WURpJwsfZY7MYQNoKU5s/NCquddQGsJJGnLjOgc8lWSY
OHgvM920QKoOg69ws46O8PkBbNDK1GiDC5LutXe+jqc47e+noRyL0zVUIFmX09/r
uQbxkJAJPXVHibySzTa5RYe7lSB3n4axnoIohLgGcBCD/YWlZwltBkru+ChKa6xx
rwhugGwIUVxYiMR2I5PhBUtf10wXSrkmxd4j+AqN/lYh2te/B+Wf9yRtwNPzIlYg
PYvUGkGt3LvDERtPMN8cNDyOtH3JxP31jbXk9UbPSUAo/mf+WGZfdqaHo7DQ9MhA
OM5d7RoEuEH78D8Pd1+opPAuHDkZgjxDwJ933VmW5qPXlnJdQdhtVcbQ0KtcQe2K
qt7xW5JREMy7i+tkByqQkpss5R6L4x1JTLB5xbPFTQhctQwb6Q/mRiIhl6+8z7ba
dG3XHshmHILXuUrWzWO6MQeOf8nTbhN+s8eBcgahi4sZl+cnpnGxb+NdGoZyz7+b
pxXdZvnUc/cqg+qRU+nhfY3lTCWINIH4UYY9NDhBM7uRNZSLYp0pW91xiexr5XR/
6Ja7gqvxy2FYpKpnvcW3Y5XoWAw9JENymAGlO8m62QszzZ2BhfFXaw+gF7U9Hstk
P71ij9tzDRDJtUcUQz+vehdyVyCF07JbkKoFod3UPbJ6rjwHVnQZFY3NThSG3RON
fbqiwwj98iRObM4Eesm2jEqN8NwXDyA7uX7BDzoPVdeJqcnkuyQ7eUslL2VUZ5w8
owCuQV+tbm4dN1Qihqob0yvaqpe1ovNRTLVLBCSOjX5DNVbex39wRbFid/fzeGQN
uV3dwdulr+ODffrf97LCNzX//9EHMWl+jmcFaplnh4KeQWgfmJOlQ/oTZOhp5dD8
e4VCGiywGVlleKBXd3n2ROMtp5LAFR7hQzzjqZrsVegQahPJzOKf9wn6kw/UuP7+
tHHd7uyAPFXJPq7RiXJyQI4rxg3T5pB7YpOKdjuBjsmrYdNfaSn1bSDrNYTtYavx
3+6L/hnLDs3qwL4F5kaWRs52Hyi566+YYvLAnhgg7LjifHPIlL8NraS42IHkI0v8
xJYEbKbI5HCX8NMJsvA4w+LL8tIrLQL3haU23t0JBL3WHX3DI0oaycPYG7DdkVnW
bEifVbAQwoEimRvZt0sVDOwVKKuwhEfUAJb+NzSEMyIQTuG7Pw6NqgXC9jlHc+F5
0CR2xb6I1UxDY+tv+EqPjKffuxx9QDuzbhC3yePUyjZ/xEPogdu3F3q68HEl7Tnb
xDq32GzCZSsk/sjSczOdfo3i7Bw+/5eSXOcEODaYPZDIjnF0v0fnIz95RrU8pYp3
mEmI7WuDZG/gbIuOhR/0ZF3mDPtKKTf6v3tjqCVR5XCHdKbAYrtLHY+XZM2buw7j
yvvFnxQJr1AsTCtApnq97z/kBVkuf88WDojkOJiBSd6lfKKxn08cYiQTNBwVaIcL
KwNXNDqXAkuWqlAP/aYC4myNGAxvcYVVVxIVzZSERg2eBhJY2Nyh4doC/e0IXm/f
5++zvNheGZtQnwltFgvftWjjQU0vihC2JEeXLSV4U5qeBdJfHTBNrB16h10cNfWW
/X47LG+XShR6pP1hmv428mphj+vwBq3A2O4wUNaxZDpe5h+pIMmHmv5CUsbt8gmI
fVKceDJ21UUi4cNSTxWvhZMW1Il8MZ7Qo0WnmVZWuTKfpytVesb2z1uzGlfXdsN2
rf8+PtL+sbta5AZ5sGJurFh2ufbVsMhnml+pI6oVvsQqWt9bp6hr7qsH5tStVSF9
/+V8q3JdFQOvHfzg1p7AruOupxvbyM8GbQXlAcc8FtQtpmFOYgNE5bPSREAe/sy8
AmKmKWtqie3Toa5ALgA7/RUS6xhF0ZyRnocMAA0lGo5x6eC/jHfBQot5OjwHFMNX
IRKEkgde3XXGkgRFkKVCyw==
`protect END_PROTECTED
