`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LE0B+XKJ6BcsERAgE1DI7xQHgAHaN1MdqTWgQNPzyHT7wQtgpdeReXFQ6j5f05xU
MDyZbJNrWd2nKAjUdXWxDXXRhx9XQ16/6ekkgXDDCVKtG/sgopExZ/rZNIeD5HLZ
0bKcU05WkdRfE18jwwA/BqmCWFAaBnJC6sueYjARKNjP4II0+NhkcZjYk9nVVz9u
SOiY8+m1nRyl4QxAJfTtAs1pFJAuFGpDARRE5oYJbVxQxrvVLKPhpoil9lkSFuKu
I0DGJMa5byHWv0Mgmegm3IPgD72QUIDKs301soyGDSf+xtSmr2I52K86CxJbhnZ1
1FTo7F2flOyxP820757IlEBv3IESsznVzM/Jaz2iOJTOHRoQSY9IdZDbBhv6V/QW
uG1IBi0SCbecCPedwL72dZS/6t4NFo2Ij4TuywGrO+rkQiDeaDrNd9A91EQzVzwk
c3wtJwZ8jNnppG3tmHgabVS+FvGzvOQ+qell7vwN55GImzyZ24Gkl1dS/pEP+nCK
/cWo0vW7Il9LlhA8BWat1Z6aSKJhrz6UlkvsAo6jV5IFT1cUqpQ/HAWY6wiR/u3j
kqDmh36an0bewqrPMdwIFYNpaFU+0UDq86el5oZxHh6iBZloQUywm3vsO4JtCL0Z
lBP49lra3mT/UP4FxZEzLYhhxRSyhTNsbdQRXqxkbTe79EZK7HG7MePVavawALvm
za/fZF3Wq9YBgzI3bCujViM67I0/zbJdveSkev9SXjMt+crnTffogKcxZewEnAZq
SKvhupWffHLRsip7QEDrXZ+AqEihkVGC4inr3nzHTaP4aBByCNmXIO91ehi9lJDY
UMuNSyeb0+S9UKQQ9O9bN3vDaZSBkNCMZ0O1Ii5lbjMvEoAUhrfycDop0BM3U68O
NJks5YbWsUCtVV1LTjmcbFld7IvVh+EIBmGzSnxg27QHCRhzFjI9fjZaWjLBj+eB
zcUgBQJr9EgsVXqMX6D1gROOyZZUzmPn8Tj5kKnOd3a6ZJT35m38pHxCRUZ8oL8G
KII3giDy+Od0QvVgMy9YNA8uMeQGjUmtFn8I2/939LL/JZu+7F9VDJAFHjncrC+7
R8xiwbqiIWzR6Pc+uQ6qRxHkfd5b98NX21XpmKf7FFiD6egqCD4xLgDqO+p1pCB3
lgEhrXlfMzxKBfsQsPwg8dHdK2pQ50w3pdfZxnlV8sAt8s80zPT0eSeIyBMBjaWZ
RmfG0oggkAziYsdiHqHETEUIuEOslyjQaErpe6v8gwaipj0ZTuR9VbKqaC7T4Lzj
rRhPfclHrgELpKo50bdUdULIdkMVQaKfsACwWRDjDfUlVsSd/1Y76BlrWFwTlAhG
RwUiM8rG11qHo9cMWuNrUmpcec3QTEkG0ah22itX9O71mCt7eXkTZbdVpS3Jvfz/
aXG+WZ6KSYngMK6lo3VaBgq3Ko+ZaNfORr9nq+dHzdREKhbpEuE+PHepgUiqTvYI
+0eLFzc5X4obOVB3NuFnS5XVvFVd+jJI2qM1xxzh07jqdy16Dh4v1yKay2cVGzBQ
m8UzR+ARRzUuGK0oUGvU47uceuvvYGOUP6VALpMsz6QVW3zviRVESjWrVLN95Xnc
9/4UBItq98RyOExSPlLYydujkSGvXJdSAuaXtnrLfHguALozb39H6y3fPdcCtpVU
8ljY0Q6lQ2kZZmFlLHvX1GNqEqeoRb2TSFaiJBtOL7PWYYbvtTVfYvad+2wjXED1
85LNCauzMzAXzEr5TlBTF/AFHWPR5RA1w4xEp8PV7/E2lDIO1Zh78p751yKivioq
AgslDFhyU+rSprg4Qs0q49pzp1YBuwvkqS5bd5A05TIxtq6dgSyQkqJp8poByPyh
1sHBq5/rSI8/8FWgAzQ+AvaAM8qrhLKuIRz1m6MeN49/VDNiOr4WOheoDQSiJdPG
FvxKuiz9pI4wmFf0+te5PXvOdDiREt4iWecCyC4yhV1AUrzBRUFCYZ+Jq2i/AHa2
MT5NKEvvmHnz8GbhDfLFGK7+Da0qtXeqV4sWhRPcZAIVnxplDFWc6tztVhVxk+q8
47LzQLk4ovIE+vZ4qKlKhwrjiaSgm+ZfXCyFJla9sA+QSifXsMKAljkGv+haefRA
6BDNGIuVsKWpKYQASHNwvolBt/gDnD6qGRp2nfS/LFDEPMgzkiiBwYUt81qOsj1m
Vh/2IrHe14JI2VLfcjeKNw2qHON965IV6FwNvSPCx41KJnigPmol7826eDgtL0AL
hXDdhqOSfJKQ9jiNQkMhWlq5bNardIphrrssWwW/KY8Mmmg71pE9M46dCbETnoBC
3Z1Zd+0JDExjI7HMcn5izYbba0Boj0hQZpyRlRr+BfG19hzBztUy65FBI0xFR0xq
0zMUtzAjGURvRwVmXiQ1jZmIyObsG8gHjYfMn2kae/ZU2AdZ9Fkys+5D6fSpBII3
vAvLxCdgf0t9orrFPP0cwwvssXL2cN3E44OuA+wT9wwKv3e8ZWE2jt4kQdwXbwho
TIf3UlCDXVqQTwRF2S0CygR7p0Ma4gTHAgTGmmn+FY889QevxYaz4iSpJg6leBfC
EMIZTt0asKdsIoJiznnvBkt2DrK/3br51NqKoGq74dm9Rlaq5Ci9XuaIVhiAcie/
qOosP4UIRUzDbQAlXmpo/16j8wxxkcgw07rYW5YW5I/euoP/8eZYMgdfEbIpns6w
T7yX/Vpn7QLxNatInYMkioBnUnwtQGckZK1ZrZdWTb+vRP4dEpbVneiQKUmf5OEt
vL8yiY03gsYDIdi6xmk5nYqzXdIr/xZ50hHmUgAT9t/YGsb+HouPX8zJasthq3zE
WNDvNpiEmkJqknKoE81HqZLh6HXvYWABeay5y/qWCuhXrqMV7oLZ7pFQrTxBU2hM
avHooUdMNdNy9rHlzCSJ701Oh+3efFoyt2S+rF5J+0ghvLKUIsdzECWDplpgWpvo
jIjnmLSYPNZm9kD6PsjwfFiqocgNNh6/QwO5NFAwbu8ZU/yp8wgLbNxoLRqJtOED
Supj8j0MTvtwa5u/sgAdIIBhaQR2LtxEEmSbilRbHYSwU6c/WQiwl/M6CkO078Fd
UX7NHALYkGLOlhIT3Bv4lQ8atijLBuXB+JqIMkVaNssALDkR4drPrXLHZ1WS9psI
NlMKB6C/bldkp4hhg7E/H2Y11LlvMtcO6O8XY+DdOn9UDa+D0+ujGNIOHOuzC1yr
MYZ/ZCW6w2fq8rvnQ8WdEOfEa05EZI+YzhrLc1OAEsuIbe+cD+dmuTdp+qI7ik3X
Inw7nK7hlyjUHtCmwxA09dDXkEvQXZ63Q0P3cXTn6M7WgdHGgwnLNQm6Mwi4Tnqu
DJJzxD2ddrRJGl6eB/Kyq3JZO26wbxHjiWABC2SP8s4Pl3pbvP61ZtNLJtxxapjL
LxfNLPQoh2VtQLFcIqJRb7IWnK+MTg5+PRF4fDuDAj4+n11BEUzHbEk633u47tpL
JchLnrTgPjAVxG7jqUpt5jSvMjmbWl4GXZgimt+pAZElEi/hDTqoxkxpwonWjwdF
GBcASgRZWwoniD4z59xkfwAz7KfL3sWdbJCuO1lIz49v9/IRzpgSJnlBIrcliIF+
0T0/Bo2350Su0KcQ6fZJD7m0nSrC5LhF5t+NMYguVIeAxm8XWD+kICTVlYGMyCnq
XanQKCSh4298CFwcHbb1R52UCx2FatxV+8AJDIfSi1b/m5cveL1bsv+2SpE0cUQ5
61dLgiMjpyezmr+mX7DCTZPmWK/9qzzjfnWvii/FGyEZB5LSfTUkZRNyO8VNoMnY
fgGM0k7d5OOmXQtiM01XiM9hpG5CtnMtVSZLgyZxJuj7zd1XSvpZwdw+IiEMfAsB
r3WUXGHvpVq9DQXnzUrjY6sh2HV4P/DBF7Tua9FrtqAcs68bN+gZGiZrYYuiV6Dc
ErHNaigfXDpJOCdWhgwsVfPxKDA6L0WJsyDmMyk1c14TiYrJg/1OP8SK/VUCoON/
qd0D7i38g8dVRdZgy3lFk9zA58ZKyKY+USehGXYWoHlJjxN6lZ4g/oxRWBsNC6wU
WdgFDNIxibO4dlIObA7fyfzKr/yI4xf8RqF6MEzLQs2j3rCv9KbUMUzWD/TO430E
LIbWHWIfBdrRaGc5PPRonTm+8yObAOLGLkQB2flWtTsynJHgrUwhZ+7KUPs8wbzI
RpmwdPCagoowN44oAfzwHfSPWMPE10pyDHAxwMFm4MxbPo0OdTJheRr1w5lXIpzq
V50OEiox5jpLnQOK06is6b3jaqaM0OqbaI4i60TozWHEnDItGG00gfLbw63PP99X
tNJssPDnYFBJnYLRgCxKG78N71juH+xqSVHl7t+GinkJEl1L8qlutBzjwMk6ZIQ8
jAWuW1FRvnXhI+rtPiblLlYg2j3FHQZju5VWZJy82z2D4XDgEJxzj4OPW07taXPj
Tgv4dTwPyV/gDJ4aisiJxYcZAJTHGe6BUrnE/wfVGKiyg+Ubyyv8WQGpweKBnOLq
hlBa3jJItEq+5rrJO5PWyKexOgQFtn6W33+Cfor0MaDd2lHf3+2Mp0BE+dYWhSfG
zV5suZrGE6B0V8nOeU5DE7PPGyo+StcN88enIhlz8zHpCORCH1w5XsGlGcAk9TF3
fc0vnijQwUt8xaSejAQCxneMxSvGd0qPI0NO7z+zCz7TahoyyiVaIcRgdprZ6t+J
JOTX0LTj/bkMkLziiCmvvi4A1JVH8l+LSRaZLpzZy6pSZctY5ATkg5kqPkd3mrqX
KOOzWlAYlNME83B+GRmJeAn+yMItXgJrYbxpGoiLbj0qvDekCzDY42002bcy8p3C
VcTYYFWZa6+20snee22q6VP/0mpHrYwU7xJT/iVaybDrWAs0r7BhmrlDc+R00Eys
RN0RZvmmnFspXmAEq0ie5VvcPiG9u7d3tRnsnte+O1aG+fivTVnEnIJmmyPoEx45
TM3bEM3pCD/d9hCBdzbWoTkZlYKaXLKL5Rq7AJ6Cxe3ZLR5STPPGuqhdB/mt83HM
wHMG1JXcbhmPdgVdTYx7neWWeto3QxSTh+sXWjSCBy1a6Fsh+yiygy1ATxbbNDpC
z8m7X4TQTXkZZ+5jqmN5WtoPEuPtDVyp4sNpwyp6SCkyNcdnN8bxobkPZu1RJbuU
veA/LwEd4/0jW9jMkOvcNtvfQvd+K5XCxP8zRVzmn1xhyD1XKM94Ykcf73T5vRAC
1plQDzj/2y74WyCPBfd+0Kr+nFDMZJwMTEiJD/cF7b0sSbH+76WfpAC0i7YbXxyV
+0LwqOPVdmXk9rz1arkkSNZIrDe+bp5ZZWB4xwRQwqvxTetmfnd29FqmF7BEAIzk
WrfE2yrphnjC2kSAYCtUNviyLVyeiWscM35+ir8+87cW3fHO80/80BltQR3CXOwZ
dSp9qc7U+Dwf0v+Tzaa7Bpm7R32tY48x0McQUlHV/dDw2tukgxHZAPzYmULjRFpy
n5pK+tmLMjThBv4E0zDgWcq7tgvHziJWpqvdEXO3xURaurCp2iGNIaoVyb4EedAZ
3LSxEbVBA6k24DAdEypvt6PFebHppBEyo0U/WV/MCozbD6x0xjSRyBu6I4rc4IbF
SKxH3nhK+ecnc1kselWGaQu1JmPVeBWFQVg5BbmQTJ/1sa79zM6rE74ahbPrRRaM
AZ04b7jJfiub+dxakQFlHQrdd9eHk664AShcRvO3gF7oYRxFNnftJ/chMqhBzCTe
TtedM4eT2jWYPLx01aDD+BHdxTAehQ7sR0NWbQ4hBY6/FqywejEKAcvCmOGFyy1j
UwBrzN2NvvRxVGC2T3x935H2eOreI+Ij3JiPun7BGzTzHMNNVh6dfwWlOUCxQAQ7
z65mypVhzbfqJs9eTepU+ujAdtXAPfSEl330NECRuD7gt1VFlynnI9Wwq/zgi1yt
KnhQQlxtcHwsapwWvfFQ437fWU9K/4v3f/9a9aSoUQ1LSb8tRj2x1gW/LAyzFhsy
u0HKP22P0C8EKH6uPrhMlHuJtRcK4Mss3s1ZLU6ym4ZPg7K8XbJMZOS4y7FZPJZX
tbbY8mA/3+CNtsgFh8C5aAbGwXUMGJqISXaEq0D5D6weCJiP7N7Wj4V67PVw1RM7
379F3uMszrjgWofmepC2OcpioOqsAhO/Pdz99HHGue1Jox4nQA6KQF5CxoY4RAcZ
xD6NH5m0JsJV4bwoMqoKYuYXR40Qk7V1g83IS6g3YcOdi90WhKZkMsMCMxlT/ToP
Y+0Gel2azHfNrN3//Qt9ZY+cnkIrsjvw7qBiJWIML+g9N0B0aAp2hv88nGdU1Yyt
K44Eysf8/qSJnTqv8WJ0YCO2wT0WlhZ1KDOlH5BX0y3jWwq3LzFWfGlwEGcJNULY
RD8y13pPUC4BbAzCZ/+oqtsB81MbJ/mjDrsteH0BGoF4VIH7JVB7l4Ewcsx+RF31
WaRqLDavv6iP65+jMAMvRlqveWwI+aRID4ObGqTneoceISowfDy+hBKwtrzsRy5v
0A3ar1CCEOR/VA5Z9t8bstME+5pD6B85Jlq8pbQB4ooDgUe/v7GBjq2SWFp48loE
/Bb1oKz+Xc9THrORY1WIsKZyT3JJ9CI8NZ0tgU8Hylxt7kxsEuifAqLHOmW6ufDP
suJUalHAfUR85lVLVPxn4Khco1fLIlPrlqWl+OpGxvLDS8TxSXxGaVt16e8fuBu4
JIS98qGgfIgiKX3X2xyx+aH/fqT8G70sYlNCR44DYI0ugbHOzZGj4Ogawkfi3vp5
l9d8LTCZMIYnd7WuAv6bMw==
`protect END_PROTECTED
