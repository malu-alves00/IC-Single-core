`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+leMGtPNVN1r7PcdqY/4d4eOyTET7iphaoS5/TDqx+efLSImniXxcmptr2UmBrZ8
psNiSkwUh5XXGBDjRnqQtDveiBiQhSV/kMBjeOKpo7gKxqCw1kip1i9R7yXHW4qk
Gm5DHhRH2yN0HaC1azie3EWfiftryqA16v7Z2JmAJH0fgZc2PZ9P+BxLvnv8cAqt
CgoDSxbBylCxHABSeiRcjtxbUZ73C5j8J6Hg+jkXGUQkLZtxI/ziBQJabjoCI5fM
oAvvOi7fe404v8A08xGdteB8JUjxaiCmCehQBEzV2Ab9tlfIKNELwIbRswcHDJOY
IYs4dyMCua+c0VslXqqckLC0A8lyHMpfYoFQA+E0S7HTXwvf0pU+mAEhht+9N9rl
URnX+w6HyHYcnSTLqcTcCXC0WLpt95GuR8JFSOxASudSHxm5LfTCvcKDnqyUpO1E
6g0Ftv8RALtRII+8UJ1harfkKNzwEX/888v//5+lalhva5lCQ7nqsHxC698u84l0
3nEtW19RAgjAyuazKj1Yy9jXz6GMQW+PJVwvx8FWnZq30H8cAslHslww2JDgC6Qe
YrRAtDPg3UASfNr533JgQCbIklOvk1jbFekXCX8EtIWgfZmqT6porTPDgNpQqmqK
XvrYxB6OCo3ane5jR5Q/MjDGLorojeSlFiFuRFTKfb8nhHWObwT0MnKObtu60o7i
5AoZliH0Ub/LCKVxoGACYw3pgr50DRb546imllTUrCq2Ebcumt0qfwo6wyhYFrhK
`protect END_PROTECTED
