`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pJGOQW+A77t+jRRIi02KIC+rmnrY3eJvAMmeUY6sWhUgwEPwtx89PijI0qXCtwhe
Jqpr/DDvoWyA+Uw9wnsJhDDelumO5ceH/K1cfOjqMNlfCyWiDb5le1z0dSRzycW1
f75NMpYE9IN/Y+5+0E9jtwsKB5In9sSngMBGGufxaK3fJnXIoeaqxrOjIAyUhmkB
LnWth9ZwP3nup9yVwSKXmt5Dg8G23JV8tJzqau4qSODidgJJjnQDZ6Ls//c0iCc2
mYMZpS+JtRtrxk86KJ19lMQvr4mnIjShKL+VxYJ1UaVbHBrj2sCnmBpxIhW32pki
gaHZdyEiUUWTyWnktmhmo6tNrqtKMEnnvVMEZxqXSY1i20ZSktnLWJtDeYzp5YUU
kXRRq3pq6/ei+Qz6+VSnQmbFw4L3cJrhp87SQvrjoYT6YYRV1OyoYXC3hsKxACZH
lhEhN66d4GufMx8fkEscM9mLQ1n7moi2jpUzOW5Tohhu2q4WDpdqPAdM2L+I6vZM
LPCfK04x29u7rUUgrR13D9zxTi9Mrg8AAbNbgmY5s/eggS24H+ZJPgGT0cjYOrqu
/MLvVI+BTsyK54RkYctmzmsVf1AK/fBz+x5nwQkpuRFUdjjJK0knAu2UnY1r4o4A
O/Aha+Emap16hX/BPBQRqsqdyD6PuMhOAcmxWqyGMbBa1ppaek1K9u+zgIoX2zES
RV6Cim+zTNj99tOe+NOm9GJCi0/YXNTijO1X+no2nxyuRUzo8rIybG0QAOQ8OBah
UgTGDWkcjszVAFq/NdhW0CjkPrVYuBxkn1DGv/GrQVvWWf0GJuMTAQSm6MWYtQ6u
hrdl0/fsZEhljL6HcKE0skatKFWikLX2LR8J8nH5QbtxleDEP0hkUw/+5YB26S4z
PljU95aEvuqGsUjAKiu7MO9qno4m5BemjHGIzExykXVteQIJirdQz4DA91pYVn+U
woRNtrlQm/9IXqpeQILLhKGfHJOsJRWGG1a5+YOmEavXSp5nVOkWAiPY7VsvRTp5
+CW1ADCW2Zcz58ewnicrTTfZ5EFvezc4sY6ijfBDMbZN00icvmHqN0tKzhZlm+wG
r/A5ciw1ooaCtKSvI7tcqNFkLO68YoHD0SvkTqahsJAl441ijnHkDIwIN39wdK8d
CstvNCf7EjxxHVNvjXnQNtUVZ3LI8+608e/qPcYer4G9k9f6BzYAc36yap0ghzL0
yaPdDtMediEGABTgNnHW+hnOVeq2vQxkZH1/K8WpvKfyK4YG7Ezq3oBeyyZ9hPsA
TB2kYTuoMqRiNdFMSDojNamHA7pHm4gf3NhF/Oyj9dN3jxPhhL82NgJdX14ucek6
1DQAI4C0aeu1k9j0sG1VyH23BSyW5Po2ap+sR0KAwTMPjqtNR6i5RN0lWXQNT5eN
tn113JuTAQjk7hBLkLNVpf9Ctj/nVK4e0tFegAah3CWPlhCencavTQ5GL09RU3a2
ZyWDnPFEn0OItLF9NxeKdJGoIYKL4R35CntmtChHuNCg0cZM5lLeatrejkOLs/+K
PaqPCcOkvi3LWtcdoZsRwDG7LGO5GHFPA6z6qzdGPPagbnkzneptLa6BL7tn5uXN
zWaHJQusDx3agqvfKsUQK+8wRXPNNuQ/skMWybXb7rliOytDCkii27WigDfjE5CC
E1ZPrW0ZWUnxvnhTAfGP+NQoglMcRFJq0B9QJPyF2YPGSotN2C2060PIRR4fiHzU
ewYX9+VcBPV/Y7PCJoN/56WJLM5h4tDZ+8rIsFALMg8iRMUA9JIRLk/ptOLtcAEK
YGk9jXB86w2jAnY4ou/SlQDPaOJIdTSttEDihrq0nSj/gCUdeD7HFOhKqKy9ab3o
xSAllZ+wuRGfpsGmOR+Z/Y50bRN6n3RjVcdAINjUdFWZG6Wd5w3BmcaGwcgffmiS
dTIRXtm58Slr4UwiWK8SmZG0/QQa82rVcxU86TvtdXqHY89oXN5hqbU0BAs60R9Q
jSaDHfi57TtT6RHTPP3DfeUv43GPaeOwVJJeQRKeQt1Py/ol6yVun8XgCGoWrOpo
zNeO+DWuhSlHIXsWxGnf1LUzyIuxygH8AroQXo3Hq4JV/DtNPS9ufd7RzQwl9q0f
SuMJ0doZ9DsXLb1RMC1/UyiCr4KZOM0qE1HgyXjtOlUJrVtVphcVmHk3HSVT38eM
Yb4zakp3lTKeBXewpKxj6vFckzWkRIxwjVRLvVFhqM4ul8y4/iIb/C/THgM/86Pv
MwN4jY6qHqJqsJCub4loYZHQrgoIWqOoprcntIYyKUaHBcz5hIiGrqVhzYnMLVPY
4Z+w+vNmxGoL2tpRpO5T2HBZQWXv4mwQUSBwEoxGNft5PPuakuoxkq10VzFBnuJA
7BcL69xZPzALQpkfVPZwUO56GJpWRxswD1xiXapigjeqsGuOV0JkgwM3FBw+v/Lk
jhXH4VYC6MLGTMUhlDkKP0Y5aMFUriFYZySpOkvOyBvJDKb+A1syWdh7Ylkacnnt
TND0prIISct9LNg4av6DjoJmpCFyI+mHL8WhKtyWqssVj2RyDY/aHp08vmHtDULZ
SvR6JFkrplIvPr4CTnU7dSoVLd5K6dExlf5FehyffVInEFkGHDpuWiJhmWjOAMfV
OoG4V484L74Ej9qINxZgeL7F1aRXZ/fm6N4lM+7sVIIkadWx9oepJFks1vM4GULG
J6hy81aMCBuBnYOM7EeNP8dQT7IuD8eQgB0yKZAgYN72GA81rRqljySbCBBxgG/J
KmLY2RsLLBf0/B/1LX7KCOLofCZjV25Ac4nfitX3FBUKw4czRQ3kZcY0ywTlaqQz
KA+EXarbU2ZqyU8gZ6XN9lTiCLQF1tPHiI9oJAHv74W+//ynTzAyv2HD/VBflODp
MlswzxTZ1BEetdJtl61rlXSxNSBMiyUxVuyhhkVCXJhyAGc7OYSAw7dkV4ap9DXa
4xaKblV53/Y65ERuYNCwTGnVolubUQX7X8arHK8AQhS9Ej+JYCH4S4VQohyA7tiJ
N1bj2Qh33pFDBEd0H5+6gaxfGoGZizY/bqRj67YiThRmE8/+njpzfSvdonYJHNNZ
/VBhf5y1pPXHkVd+vNUEkBJQOiVwsWog37HPtmYD6mjptKsYxjltN2ekFqu838yZ
ionYIlhc8dNHe3f/AFnOaySIqopdaYrIeN9Z6B3zOA1MyNQBf54zb+YtAr7EzJ+G
dDXWFAzZkZAAgrOyQ+OOKYelssVgeDtDxCAlTUtICGPJOwbSyO/jVopLsv+W+4VJ
ahAkIJ4VaG5s4Ixg+HvHQsQCtMmTqbgS/wpq1UmJd0zBnQD5Thv+sxYYiCUos/t3
PDmQRcGkKdxh86fE9N7CuOMT1ke4A4dokXudOxFvyo0QTq8oNOfApKOoie084xyi
lDqkUNj9CY4NPfBjuBcpvOWD+LdSJbE2gyyU3+If70BN+9BcQ0XwsWYeRC0aN7Hc
o3aSyye7DDYELSptOue5W8xJ+JP+udFT7Nahf2/HwLCsq9rbTdo2RwKCjziJmtYQ
yrleqK3D6ZFZTiih9TvmtrSEv1RyQnkQJzTDn0QzLzoydiX++sGeKdkYlfWx+NV4
A+H+rc7zExw/pYXQnmh9Ct+9X6i2HW2QJogFgWQtgZ1V0sMInFaGhbNLAXU0kX8P
T083gi53mHxiii8+II+ME3PkWvOvKgAFSSJSl/9LqamMXSWKutBa9YPFepPOT8iL
H19tMc5jZ5K34J9lCirAjW3HJzEms4JnYOOgtR0Vio1bR/CLc1KPZwJr54681ZX9
05zn4tgz93Q6pfc/fBMPIy93S0yLOhYs/wCYDKykkHurMEFhhjpBWtc9SSnd5n4F
3txkesMEv6i0x2EeQygB57JE64AhMrTM9WqI93aKOczMZCdPKGN+TsBhacYmwrX1
g7WT6MCJnR+w0qn1Yka4fykPIkp6xwv8XisjWbnv4L+YmPZqS3zGPKcdbQFtBX9U
pC0e3xIhTiJcekLqGQmhbEhn9OV47z1me8me63woPA/Mu+D1Dlw/UPd6qqZ/ykQO
C7nNBFVFs77xKiCyMob2QUZm5PNcO5l2pUDXZMmw9a03gggWGe2IRITOjo3Yq/Pb
dANxP8dDuFnu+xokokFkmyq6Bx3nQWOiMa9EcvZB5/qF21tNr25ATb01Re+HdThN
K+RvALTkGBNC/ikgQ0NWXvX4Rvj6I9BkIZFGZka/Gn+XwGqeCX4KwsM56EOPN9xs
zNGvsBsD9iHgruCmsiC0rEWaSGWMU0SFo0DVj48wF8wq71Jexk4mP6+itFvTjvtQ
YIEKRo2BnByZFnxv5Fq8eztnLPQ4T9rPzwFy80u85N/9WLQN9qi5QAKc2++oQ1he
zPLyZJ6H1qGyS7zqag1uQActa9qM6lu7g/C4z5EfK8Ld032SxFw04Zwi+/xW1ED6
cYzrOaIPbDU8vvcbJYv0h1ll2PbZxJ/xCgtBaeYPd6cDoq4wrvYBwm1WSFQ1rXsc
hMhZBciWb0incUxBkHX1iWYo1JODM9fJh4HB5KUnRMd0Na+cbw8rUV/PSkfkHNSk
kPFzY70snY6D2ZQxfJBsV3hIEG0r2PGoG63K4SWjYBqIkQwHkeOblEZ4braiOU17
xZ0rtzpPD8/oA7rLBy8C/jmFY6a8GeRiZuYTQww6Zqwt0NtVSLmxz1txPBeERv4l
XpQGxXtcHPTL3OM+0CpSX2iIdeuvUyerh8YV12Ytz8pYLhZUMSa2QcKraApf+hDJ
E8fV6KvJNMhOgLHMH9BwQARydpiI3BLQYiy+zveylHczqFMM47EXRS+2j1VWmC16
Dv/fQueoRAzuXmzUolBkNRlUjK4SG7BnUBLvwwWmUL/zpX1kXkrF8bBB7yfqm2n2
kNACec9gkLqwjyDTRIMmxgAQPlcAQgZqdftxI4YI1fhfio1f8N63KCHkBf6p4zHn
XHkMDNPB2kNoZeIkf6iqJ6l61AbyXaa2viX50KqQE7jeb8BbH4hkG693SGspbMpS
IFmtHL2btOz/WgTr7o721c7YsAB7m57ncmPeC+xxTGKRf1MITLAZoWrg9zGpMy5M
kmmzMGuhfVl02Jwz1BfG4VwLSchxA2DOZG/8vq+yXUFbyRGx6vGviZ9xNl35bmTz
`protect END_PROTECTED
