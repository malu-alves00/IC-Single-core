`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dnZwVYj/jD8YkgvZK9c1/lnANc11tCs4PK7SaBPEJ1NZXkxU8kXgOFi56ImDSn4y
8a6K8jhq7hdDLKJ6YGFrRGzr+BqwKrrE96pR8CnsZ7YKskjL2pzxQ2rHZGxLaz+k
XUUGiOSwyKgQ2nKajUFVJb79pkC471qLKVHegcJtXreqJHUzauOZwOZA6MA7mdU4
ytNp5QEph3u3kZPWFDti2kap031J2VixfpJJ8nmde9ymkaCKrIltY9W+Zm6YqBa2
94DVsM2o5Hc//6XkzACTdlu5bqi3cLQ4wKK1l5iqEsgk1RalmPaPqjSR4Dy+1XgL
oornb+r3XjhiuXdUZRUQfvZnD0XtFdSBEm9KlBIdi4YyltR6cUqRCsM2XXH1B90k
NlEh5kOTbDy8zw4Ox0SKU8U6mUKnRy0b0TcFLy6Iu+kANPjeYdaH+cAYwYpOuKxC
9XyPKS8IWc2fB0zt6qM3GR291byZ5GDfM9Q9JdFXu7LnBFiFFURBdFnz7Sfp82oS
UJfoF6dEPZ06HfSRXxJ4+sbC1aQp4RP7dctgyHmslUo4DuYjZJ/QJS9yjhyOemyr
siVCs1w/3fKbnui/dgYn3tFDnpvZ/l1bGW0VF9GSnWUik8+fYV/YU7W/BfIGIucE
ChsOKteZIg4Jb0j6Zws1U75I6KxsS9bz4mDU5/9RhypjnBURPeiQmzjAPOOYP4SH
le1B2N06GXeoDVj4/Ipiub0w/yl5C3w+AmYwbBe8R4Q6uKplmA46dtj7cg1lUCdI
D1ooztKq/wWPlPQ2u1/2haj6xOVu9ZDnm92lBkf7Mw1BFOkly8zC+hJM0ey8uIj4
47XyDfvkkppEOE746NASNc74cg2VE25vC3CCfpNlPMPKqabsGjpc+9QCxL6Ge0bN
LXiFLDTkJtDlKtn/Nm+gsES50/9V1AkTGb3Kvj1Y8W7sGsVUWgBwOnglmmhbICPF
QUAsOsP9GVGyUepd1RWwY6DWjMVPsGNa14DdgwdQPhOO+IdRCMGXVdAjmpdUCjc7
JzeS4O8kPHjC8x+cS5m8DNzfFJb3UeDMh2QJYMNNLg6yIc0uVr/Enmasi896JOqT
/0NfIOB9Mj6zVpvpCDjqP5jIPjJFKGrs9XhI4+03vIM17qp+JOo+1g5YIp0Z4Dp2
R8BzKZjtJIEf3YIHO1RVHPtqAAluyEQ2bJ/P0ChvoGxPJ+2XUBVUcZgsfxbbqn/a
3a0f+rSC60fIdCkfNOUT2qv5P7Q+ta5C7k3T3NS58ucz0aOKW7KtPVcrdAkNEXzI
zqCCR8SjVEUyfJdt/uAsC10itDvVLBTn0D47tJLRE3kwWu2DOJqdzMf5VkCWLSqW
xv5vwLros8lX2i1XwpM7Kw7jqGmq8197tkpaqGa7bYwhkuoOyf2r8K3VmtxbjZjV
6nHFInGCeXmfHcirikMWXLwSQXpFfmbpO3wk7I/Gm7WrvmIdEmGo+9KPYnYqwXk8
IhY5PJUCe60nBZpzkCanYjTMvq5V6mwDscPJcOg3gKG/GVrlxCilCYC1JbrAM3He
A2HFCTKsgeX9TVLDX5LZ1UPBeumWvFwY21bqQdo3KXHPDrUFmqak31PvqAsvx5S9
jLRiBZrBQ2dEeAk3jemLi3LpKOop3s1/EootdkMN3E34+fT2gZfaYc1CK2fRCwaA
HQ+H+Sl3auNJ9YhQFJmRoLNdJXmp8iZGKpRt+DL5NTdUZRNti2N+HMbpb2cM6liV
euNb/tGm+71nUYZYxkDQcAgF9AGO5J9t8JYotxBCgTglYhGNXXhKUHLstWgHbCZp
fj33iNjpOwHp1Z3jiZgjhXwcgq8Y0ZHkRq3SqFHplml09Vhqd1cB0oyEVC8UqHQS
yGSbiqf3IyuI/nig77+p4+KpZca2cUOlyFzWQnE/jbo1sbHBnk6rtEcIUh6ZehFV
iMxdGvrH/PM4YwAXp6TH71Q+V+jxMd4Qw880EVCEkWl7vnl/vYCejehLl3XGtyn4
Naa9dcGu9glbCo3PueP+/1LVhYT1Kexuxz79jTCmNC0kkZAchgm0tfHL3Ug2+B+L
uQudwSeAmP1q9rmAulv/ISpWbmHd5mHthhwUu6S+xysdmYZ0KqbQXr3Jwi3aos9k
8xeVMVqNQEK45Eo4gBNrGS9p4MkaJSlOehdhXk6nU9zlxTLBEn9zNBhMvF0ym/JX
lCqC4cKbkdozqICxShm8BcSjrfWBUfklxO27NGVSBGVc6RwD7cNG/9nzdRd2sKKK
APDjzKAas6fi67TqYLeFs9F2EJJkxWkkdH/7AnYUmYggVsiYPShlfnHVwWVK2CjI
E/ZvLLmgGvtSFBE4k2vXF3UJWm0MNnwgOZS/r0PpdTu/UISdl2vFyXVN1mD66QUC
jXtXX+xuOLnXfKar7hrHDAtna5jn4Yy+wfNgDEx8lEwOuAxpMzY7NJmOTk/6VzT3
rSHYFgKvo11ys6DZXU+mcw6Fn7tCezmjDpZjIqxDBpIOU6F1rnWPHZA+V8Brs5hA
EdqacdVb+SqCB580x5xsO9UcMCYV/3ocVx9rGthol0PHO2ojHchiUV90mwwDaCxK
8fkH0ih8XeiNLRDrQBiQoZCCkdUCd3RQSYtrGEkIcXR8uhMUF/lYTjLAmpG+4XGi
8CYeQdFqeA86+Z+X8J0nBuGwfv3XyHA1BMMB+I0pw3A=
`protect END_PROTECTED
