`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0b8x/G7Rck4LGt3WpFxZ+Iozyk6mhHZZ2qSA+DphuuaIlp8yvXUSwJmX9bSZwpKx
KCwm7e4dmzAuEdCZUsiLcHQuEeqWCcqUHqACDCQkGlJ1DIQDH1WtG4QR/cAfT00K
+Wi1AWpYAt16uIxpTNNvc8mt1GYi2umtTJAWkjEzk3rfGjSF9jz1o2UyYw8P6kl/
37SHq5knt8i07yk9yc9gAbsrLU8AxBKpsO31043Qsp/9f5uuJ/4quEcMlGfRT8Dj
wQwN0ttIcwAI7XPtmeFeXquPw6Em8i18QZ2aQtgTBk2UI9RE7QrPTAHCAy/ueOk1
RxKdLWxotCno/+mxIdm/6iTQDXCKayEPi+k9k/rwxR1+ELZvntz5bRZTvOMNPkR1
olVFFEfjLOMBz4OhpMZ6ByBdLyBeNvRtxKhq+FncUWd3D4zq6z+oAegsjagUWK77
y/tcSnZTqqzeaWwScGcIlGppNqs+AjE5rurCs4nOE6iPkpVwr8FdyVQGysLLfdEA
dY/TdtZa6zcq59/FuuyR+yHAM2M/+drl7t/azh+gk88TouyKsp4PZ8j7kAbKEidJ
VmG3afTAMr3hmoK02V1lGjHRDFE3Ple0/ni+yZV+dlJhDD32BC9CTwY3dVFoi56D
+3CPR2f0RlnF5EKex7jKrLHJYcEtG2jB3t4YGkxhJkbotQ8XBv9iTeDjVICZyrnI
bgkTL3RmykNufJduEJAvxZZYq8wNZw97MX40dUaDIGdRD/2I2Pw1wKyBokAeoDx0
mUOiq8XYwcV+giB1ygn+lrrbiVo+6rjfQNidw5a7BZrNpjJCsjLAaYdek74KvoxG
GaeviUyCCr+OZRjoW9imJHizcq15hj2QkPwIEQOyILFv6V5BBRy/hbF/v77W1PWZ
2lFHYG2dZC1DF7iySzu1qerPpHT1d0zqubtZSuLhqLtKPv5WY00SJvS8ydFr/H7S
wFMvMtgH+qF8LZwdz4UZyunZDuwjHh/KsUyCMd2ITbRWwsTy+AQScnCbkxBtWh1V
EINPskKn5DTVMpOZnr4vm0yPFSskLpjH7qscVZKbSed7awFlYNSR6b8o9QT97rYJ
BYpMyztzdliPtB+6tsjQRuo9b+ttaAKvg+YWa6ys1gdcbbS2d+9cY4KmRfdbfHWz
x2A+j/2VpxYyY4I3urzZ+6v46A00Jdat67ZocT5UOw0ENShxC4Qwje7t5B1XAeku
tpbQyGD+pks0ndjiQadmpuIH+J4b9YlGbb6+tB/NdruaOSTFYkMlk8gGT9P5NXc2
kynVZgFmFKtZ0/mg6Jn3pai63YJ7hjqKC5HyhTA1oYMNPjH8A1oR9RbNiwnsMHKi
2e+wSSc3CtCtBnKmqFy1GnjM7mhg1YUEl197+DX5N5EDIKxJe1fSyQSyzfUwuy56
cFIVklS9oE/agUAclscIdMgCNc2l1w6FPczzBud5yOXC57VLAxBD6jmvfCUSv6sv
0ipRGCy7RzfpywZEH82CP5mdvdLEhNtCqQooPfHVFT+Ojzgi4vREXkjbVAEhoVHt
QTV68FUhMCAI3wbDpIzfEDd4nvm1ZNIz17cZwmBFp19GuS0h+huGC3JYCRxSyMv0
0xMJP1CdWPUdpkodoyGjeL+D1OcIwK8AxI2goJz84fbfPqmyFf8Sooyi/3ihPFwQ
VQQjmOCh5l45IjjM4mqxQ4AFPT74IVOFeSSCZWbsj0pLRD+gd0bHex+TUcDZukAj
/Pgb6BC7fWaUjdGOrkoDokp5dVt+bl7jqLl6aXQfi9KSWqqHN5E5g9jlck0PIuGt
fvayNHFWzEzjieT6YCnmQJqtpICRq3nix1SUkx/NlqYjSCN6EEDN3Pm/Apda9NP6
d2PxSoemVqiCt1TMDhrRqcnh3fjfMm56GPT+sKZCU+vKLhr2th5c1dFnTdOMradd
7jSbNKmFX+dS1OkrgQm5r69SFbt+llMz3nuemIGFc4jXlAEP6fciL5gv5jRAUZ7N
Zr5/UUF0swN2H9AsLSGqwnZd3aoP+/5LI2JwihVXBVPt777NndTosZbmCoSEqVze
t3PPucJ4/n3mIxCST+YWexiDxUGuXnoLRwIPRlpK5vbUv8YLtr02uP05re9DpaQ9
Nqqz4a2BuLAy+VJZi6odsZJSKMivpVWW/0q5wngYNVrGLIk7XieDlrzXc6uA5AWQ
gFt1XdPAHfwSZxAMCuQnMR8UgFy5Zp8aUSEX9EiruTDaHEFvAqMx3U56WxMV7ppA
XTuk6eFrPZZNc3k7XT8jJpbb5wGAqS9fRcBeUwDOFZGKaJ9pkLMiRtTsSwIzLHpg
LjsmWzZaykyDobocTwWTchl55gghIquLbepOC9tQu+8flRCBtOwrsc23odJgAiac
TJwwUcYihCOZ+0H7PrRuCWUGAtShkGO0ZPJhzTf1jwqmOrnp8i4chFLlDCgpv6kI
x7VaOgOWlNfn6hx2tx40jafjzp54cR1Ni5+VJ3ndh4+uu4S7X13cIwQqrUVcIUvF
CIDO8cu5irih5gWqnzSZjVS9+sXtvXW/mtcdKLwCE/Q11vrZjpv1RlXMZvEywjTs
RsYefXUUKWe4gHgKm8IlE9tmZqc6z4FTsADbEwe6isAQVtgTERqnIdqenP23aogc
pOY/6CNNos2TIdVyVZzUbw==
`protect END_PROTECTED
