`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YCCGKT97OXEHNodb/7Ex4IdKt9z/Bxl0xBfLvjoSXKerzgwJpm5l7EcdphLD5ZA6
bebb7xa27aqlUVS/llWZyVNvaFj3R7AYg0rlc5yoZYb+Shttf06VQjFYlW4nc3d+
YvP5jDt/80CkfV3zofSJ3mHuGzoyEiFGmm0t99+2Oxy/NBJ45/acSFFrAJhf4b09
t7pDfTB+JBp94eBNx0YApwzavI/fzjjQ3YAnOleQ0ibquHGOO5+rTQTniHAgpnPy
YuNlydwtIASOq3OcDsZRkp/WZ/6HB20y9ow/KWjOExDDYYeqMy8/pxyKP5Uu/CW6
tgGV8CrTn7NBtVeK3/q4p4w5YQuoLKJxiBTFEElcfxcDKjoMWKf+4DTIK6SseXIF
PGEdJYb7W3V1KVloc6ekKU3/r0bZV8HX6yYMqmkUu4X2IYs5LIRqNQuezuULHByF
nB+DcchWAIGZwwYiDckuwClTKT+RkNCCg1yct2YQ/zxK3JEgFSMV/eU2LXVck4q6
Vm9d9i1xsv2HVBsrCG4Zd9HdyJmqtvQATKky/5L70S53btJs4Qnt54Spg2w1hSwq
rS7Rc83hobUD9Y8j6ULnHO7ozIXPZAJtC88xis/NxsiJECFCqJJfi1J9eSuRABM6
Idf1puJ7/VUbgKpmLdYgGMfHohv9LX/bl2ir6C0P+zv3tmc4H3qjp/MXImsIfwo9
9uI30mxArgmHyFjmvsSLXsjdEV7K1kV5IPX8NxusQKWRGFwVDMvI0yuBnQUB1XOm
m41rx+VgLUHFzoW09AOML4hYasZHjcPbW2f0biiAOTM=
`protect END_PROTECTED
