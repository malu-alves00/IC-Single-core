`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4So2qFdxQV+oREsiLP4TwoQOIZQzuobdt9ck4ZUv2A+SSeiICfBe3elpHiOpv8QL
5rpemk3mD5HNgBEe+4+iCZVSnM2Z4p2hpXlOs8Fo4+Qolv8OrnEpEsVW3thYDyTm
vpz2+WYlzmTw243p/AWcVabolgpplRVYjHhCZF4bx2J1HFLVzNrvejb81AUwvV+O
ggjUECfC2AasYiHzQ+TWxadpR9utjKxIdBlDKSvFJ7p/CUONoTrTJumhOEoSj1DB
9SVf/WRBqaOUBwp4CC+Hmi2PHZTmXKU1j81p349Hc2KkdabgeE9Tn10mzl3HTjtb
TpVzF/ipw3JdnRTOT6kxxpGcfREDCvpF2EL/5xnRDLiL2rGI359RChtjImvH12S0
KNaS+u+EfT6T2wYoEEYOjfz2WKnrM0VSGCeuiFUFKT8Q685mzN2KBhGQxHTP13X+
zbNkAefym2RuYBDuoLmtiGqw6+kRBYrnNZiMoW1cST4ujc1nLxDfWCud+ct1eMyN
Kq8bX+TG38h2p0pYS6aOLIt1rWnxprEK/0Cgd9UPCAgzhLviOjgVGidJtJcRm8RY
AtoKMaDtCdOYhqFkDv3cmZB6/gt0+hpqxIEjENQajFs0IRzuCR4rXp6eiuX4bFZ1
c8z3MYAVf73BSF3nDwsoUFQwGBm+Y4kZI3x9JNjtzYGey5lr72ChOsBpoho7hzXc
8X9DukyDj+5m1dzq+S/J/yKeZBllIDnNdZfz/HFUZVlNVydTiDCM6OazUMoCHhwf
RCxjCyGtJOI8rxSKnMaxldPfQ1qLYTp5unjeENN7kBkKJVHlPkZd2vE6KUKvvIx/
p2Q8d/FRxmXtMKiKI7RK/aGnU630gQUZ74JUtwvsfV3kiB33qm3vFkxCucQ//prM
BH9rYorr5JYKHq0nBDNU84tj6IuU0cVGolPW/SrBIQ14L/xn2Mqrs2x6juL3qNtz
CQLIrWm7nPAXPGVHWOkpAB2jOi8ANRYpRTQh0xvmVxxI5cL8USByudhhdMkaZVxZ
EKBX4I319d5XINHiOYSBaDbFUSakJvq01QDtP/9EUKjUBPYO56gul7Ry1fWKi84n
lxw+F1ZFXTh6cRnipGRZ8uqZisHlbd7wr5Z9/mljQONhXX65Fqc0VX8wg0LkFNbU
fXuMUly7ed4Fa/kYP6pCpWTlv0hSitjD4lvH+e1KVdtqTvOfGGcY2pGpuilrDXGs
6Gi2o9z5MFBf2YzRiUc1JWzupboDFPIgi47HSrHrqwFVU2QN/x27PlIw2TxJt+8/
Fder6VXMjx1hhvQ4YkBn/q5gWEpcwAeads4rew6GMML6sZ/WY2Uzxbc/JDyykWPi
5eTfum1kHYJMBN98ob0dnwBFmsP0K8jYXV8G/8g3tYyIyt5ZiLOrVQ2LUwHqsBoi
jTeojV/6wWoIm6h0R9cLnmwCMlpJ+k+dLna+J2YI33wKbWidAS1ia3qNgpbSziLg
DCrTaqtMHjkARtI26+1QeJIR+v6Z1wzjUTyUEIh69v9/aiyTV9CgtM0Fv+vX7bLe
xT+SCh6RfwqxLBSx/kXds4c2Foaidd3L96sVgW2Cl445enatW8L2pUWfyWrZKu4d
pIqOjpL8st/qhHaB3dfJZuzRjdj90qmKAcmGirlEcxC5CAMHQu7XXR5pg3coDKSi
6KUPFoANuLCoUG3YXiPKvpUIhmEjqsh++ONtYT4AoXFqcTxjZ2lRNgyIkwmfkJo0
ozoX/R2Atcu+EmvC0P83/BRqVwSobNjUT5yUSo0s85ljU/J7Sbx+gO6F5x2y47dY
hfOng9LwRZd69Z3RY2VrGxkO3l4+yZvNExW8Us7mK4XLoAGxLO6se5m42ZMREoT1
2K3KvCeUWwRmYFtRvey1Sul5JeRGF8vRxhzHzD8hEaJF0TrZ50zySeNt2/x8VP2A
Ot30OtLPcDXXfl6ihgY4n4QVt4wJz9B1HuNQfNxI9HiM/hzMjfzXYJBEZyf3w3vB
JJHN2H74zE8u34x9qeTV541V1t51XCl0AiR/2yRIlO7TuyqnaSqEmyzekIki8wy0
AFNZtlZaGGv3jwr0fIaMVK25/C5cbIHdRkPicy2LOhq1MracLXILbGQ2zX+JdXtn
Oep/tRYCu0CFCZuQwqoJhkU+/EWCa1ixzcSQ+BN8hl5f6J0XbHkpDaWLYg0zVoka
+mSJRKzj30dMBWUmMqcgbmKPVMKwbqArCnVNH7rrYBxGq7f+d2t49GElpebL3OsN
pT3/mX2qSXt1TF5OvagJQHMeiylHIus+Amxf2Rz7exLuc0HUESAHTrYQACNkhEOI
gfxn2XwO88w3WgPMchZLVgp6dysqwTZNYcWifcT3wjLY59g3+Lks1IVpdiT9YLMO
0WuiZn/xUBQ9S4bLWGyhYMXd+Jt8C+4aZM1QDmeTgllrLfwrezEVJhu5qhuTp2vd
nNTSuSkKtMyTPlDyFAyybd52y9Ocj6VGZeghSKYQLVwzm0NhdhlwIb9QzIt70H+n
2hPNvZmph1IoAGHmLE9ooz0fUsGUFVuxgYC1Hv/DkyUiuCNOwYdA7Yo8XMotL9DZ
IrxECv29yV5s3XSyeR0qaC1nSYnPc084svoG9WqQMsfMeIcKy1DIBohG01hdlbPY
s4ZiUxQkzA9ymUStYmdxA0nap6hhE9ECm4XSYZ6ei9iG9IZfROc6qxoOn+4IZ2PA
kjzZXYiijlEVk2oj8zD9eAA9+QprQkCT3XzXN7C9RSAW/VrWpnrzW7hcZTAtByZD
WE45nCs/y7Wy9LpUQ1qGyF8Hen25LD4ox+2DUm4hgrFF5x5GdMpCKJgBhangKRCn
vTmfxzk1/lOHVcwCvfRwdO5GYhs9gGJLDmDmFnKz/Xk+2LLrN2HVYozKx84G2jvN
KZiAIAVDavoG7IE9fo5xqbaJIdCyni+uG9AC7/lQVES+MtCtnperMCeGEE02jZc9
Z9IfiyspOGoAkoL4kDw3MOTC2IV0KIWDqyg1q6AnyxDYiWYRCYMLW3+MmdDqfR9E
n4oLIBa1/V4n9VSTh66qr+pj6BVyYiBceeV9Vu3jEtsGWmiM92heRpxLwNe5m2ON
usjRRP6ZViyhgqIMaUsFpwJMzMH2N0IW5FXFm4t2AKSY46raaT86+NFLZgKQJzMX
tZlx4An4PlbN19FZ+glz6v71ztAYnhnsQaj9TEb5NFpz3qq3uLlTQ1S7KXC2j+2m
WsSGar9xHKPZ5wYzDeNXPxlce9m/1SKYujlR5w6839At6ic8zaCXbutTziV/V5wQ
3ZK5pQ/T/xnOyv01b6UOt9hsffFw3y8nOTOhX84F1RSYeRFdVNReAhl4rQt+EQxe
Pn08M6ZjQz25wIyW0wR09JQgyJPRP+E6LXKVw2CFMcC6uVHbEY3dDDXsI6+HJSFQ
00N63WCDvK0M35bgxl9Kk8EwydbvPbn4MzZYjC5Om1rGVCbjZR6xd0DT+Mnuy92o
byOmXBS27GZbK4CbEn47QYxtk4IjLvhnplJMZihI3hhZUZPlnhALO/OwGGxu/Iko
17psVHRw/1GEspnwbBK6Y92gPoVGX8U6Ikc3gH/HAL1C/Afs1svQ/X4EEoOY8WHz
9ymqSOIrvlzxJJuMZ+OL1LSbrIS5hTcUm4625Hi87joPAVqXBU1WsievhcLsLcBD
pUfQdQarzxXUvM5xHY9vc6u3lV6Gt6JFUm4RsRGmt9+uQ6HGgJE25/Wy7JAf3GyN
CLjRYiuGdaKZGuvM8ZLx2WZ2iLNB3iFeOPdRMzJpjzv9iFP2dPxiovRR2hh0e0A7
7hAUq+RbNAmiK0oP3r3lx4gIkobZjHbkY96XBWNxvXKoLuuVmQukrJfrIbVCUi0H
oJdkT+RcQQ8NPb9V3nL3M3gqO7V1hgGm8DErU1rGmvlo3uq7N7KaMtJjA/U9MKGN
2gpC5WYjYx6ElMPw+bWBA/D3PuYIXhcl+tkXFnyOvbiosAvi53goo0i+zUe3XFfD
0P3hmIlsRIUpQ/8RClNT1O0vPorlLGkbvMzONyY+GfGMHtXN/s25ln0yiAlnGrln
yZgMvvMJakXqIVQv2g7S0TacPw/+eoiq7WR0zUwKJswXN12D/ImPf3vDAJRw3RuR
H9e9BkmNTKfeG3w77AoOBHBYEvdkvehuOTu06p+XSIhbYBg+yGhk/9i35TG1gQTV
inXGgUqUXE0eqdQmWmUmG5lfhM36V9JmIZqUpgH1kpjZn6RXHy1iKP447tvm0Q7C
Y3nXNZjnTxe+ODWwEADD6sxwixBf5/EJp++BkYT5Lqcti3eGZKADwWKsa+EF6lr/
JtzrzLDPiy5T/DwAgsvVQyJcZ70s5f/vUd0lQp+l4NKZ2KkahXus7KZ7lwkcZLzb
98ytKEHTjX7QZkUq0nCbiFrivdGUhqDMJiRCNCg7sl/yeD8xMWqMMel11kts5GQf
L1JKYxtVCaZW8hgyWGewjMh3dx9CTdkEA/Aw/NEe5q3mlzyZS8DDErWEXRJ0mhR0
Ubx5aojBKR0tfhN63Wss6rehnCpjtAV7cJLrfFJNcgKu2Dl05xyTMTz5mLdn8IMA
GUNiYPAL8F63FLpbqZsgSNHOwMWAaZxZb4RRh3SdmWN5BnGExEypH3tVUXl2syzl
CfGi4Z4JNEjabETVrVN26Waj/6cRFYaDdaL7mFavTJJqpnFLNhAiJ8TXbRR0KtTI
iEZUDVOakIeTvzkReQETMW+11hQ0669Kz4PFzNHVASoL1nXHgPbyKbYm9Z626CbB
FQqFZTae5FlhCYdhKAf1OM2tAYXz4PEj060kkx1pbqEnR2W9ics5LAMjDrsbXzYN
C9wRan2A5k3jhkFQNFiMLZ1dy29j1pE9/snDrKqFgFXXOpgiP1KSS1JAgOctC2Ed
Vw7JHI1ao4uPcvffmzO2i+GXZPH3ibrWU49LBpBJH0/zOFiMlBTgZU8ivuwvpP/X
gH36ELrbei3StFb+6UEANEGjOJXwtJkNMRNNJJTQtx+9Uozxajlb6Uph7qdClejx
X4/sFIv5B6+/NCYKlVeSNlZqzMifxVKUoKs/3rnn3WTls+NQUdcKKpMHWVZN1p9a
dnMPmGMdODcmM1/93+wFSjW9ZR/PcjCwYFRjGn8/lAsETymOb8SrwZrNqxOW+DdN
/pYRHNgItsimQUyL8K4dP/hty7yyRGO8ffRoKgomFmORF+k1y/RfYcEQNicYixNU
DBiBKYViuNC2/A9DzN9BD/07wYApkDDhNsblg3MpaKjClpVpxf61Krzzm923g1EY
RsOOliKgP1+PfLqKPqCyM2jTmV5btn+a1XYhbxFaQ5YsDHmXDFhR2IiIR2+2S7Fs
50c7lrXQyb3creFZ8bkuPTY0IicTiNsODoXtY8DRusDLeCgFGGDCjQqDwbGgNATQ
g6u+qaGO25b1WLB7n6D/tOrnvzhRCoJlILvtWOG13anClK+YX3LA14XagLvzHSNd
oQfkfS5PvfbMbW/jag9TEj7Vzt5O7+VEFX2iQCYK+371X/UM1NqhhsQ9ObDlZ8AM
6pprFHgQOK8/r8Fj8fE3sXciLL+8TRB2zrC6eNQB4PBj9TQeQ75k+2z5rGS87CLj
Sgos7fT7WX6kMzaaPRnXKO5kjjqtm502TPFO58xR4Z0WxcS9ZeLp0aVh0vXwQYSr
NUJDEXy2ZON6/nIJsmP2uPq29dbcvT4QCK/718r1bAJ/Gi97bdp335TSF8qqiwhE
Q5geerfd/cKvCg8T8x0NbJMB6bXF5cEzX80VGyl15nje7buiETmUC3ucyYXw1y1S
LftqU5MNTDqguKOJtKS6/GP+dw/sR5lRoywdFbPrZEqO8znSwTFAiZ5HBXm+KYNa
hciaL+p+sxRrDpWG9uZYiM33XxzGJ765MDdsLEOiJkei23kZSmCPZl2ZFQmPvPdZ
lrpOdwTRROu3K1kf0VodsJO8CD00HP3Ad/jYc27Z+kAv/Z8Qlrna9PS6/r+gQ7sf
flQkzWSbMC4eh5VAzuBHsrs/2gha59WLq4zLKMr9Wuqjw3drWhOtdQUi4kUsQAoM
sIrGxwuupV9nnkHj8Xvc1wxsGF2x4TJ+sTWoqN8HeV6mfXNLWnepALiuqxdaMP5G
nIox5F9wHWiWemFiJNUqVyPtAJN8SMaRgGVH3cOICave4FWW+e+6TBuwegVyLa2v
Q+mY4WMf5uNowDnwDrx6dAlsVnwI2GFeIPj7APJUJoRuX+8Z5gldL5AtbCgcLwwa
vA4QCE574EEU3MNgzIiFJTaRCB4Bs4pFj7fO59e2d3eL8idwadPqshNVnlkhms11
c+p9PwBnDKarrhcSk2jAtf0Md+X1O5WLNK3wTbLVVNaELZ+yhY6zmLFstrhFGGpU
KDZwW9ld+h/8VxQ35QQjywkMKMJI/oX1PTwbEwrHJ19gEEAffFZ/gZNgTI6Obkry
g8QSfXGvlJcpIqd76D4aqXKdydH+jlzkgP16mP5L2Q7JF+LUwg4A14iWUSAFPJp+
oGMnB+TRov77N4L4C9gt2iew79L/TgpS9CnOgd0TfH9gLqMfu+N1UM0/WLZGnNSL
OHD6VO7dgj9wfbCjhTg77MuyaUwqks2SRPoi8yCCdhmwtn/Wg2wYxhsZzMprmW1W
cJpmIJslVpq9K0TnXQj3nMiGGba6dAt0sORcjqjfaySNfqjWmAOtMBJ5GPX02a8h
`protect END_PROTECTED
