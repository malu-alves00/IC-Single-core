`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YmJWd8SuOdTM0JE34UWe3rNXHUznnquIJe+4qwhxmtkAnfA6JwKrcvI7ExEQe4Pl
i07d3EuCc69HNLB/+L+Gt3ve2LdVm0Iq0bX20yyk3eboUz+2C0MA77ezFKdUgkyU
DNiISSjfCWnO8Z8UezC70psH4gHqQKXKerro8XMF1mtf3uBX1gONqqkRDXQW0rLD
ghITZdaqrDb2gpbiLdgQcJIzFo5knuejBjEp6eEvBjRtFuuzBC4Wmbh6Dav6rRxt
aios7DtMQT9V/Xzwhzc0CSpfi4YkcoukRLSthwSbV1Cnk9jqkWmw9d8qxuO86QCt
2Xo2wudjcpRp2gD7ZJ7hzIgiQY46aaLm8cDL7PtMWcbZnVEEUD+OXaS5/GcLchQf
r5ki0SGQpUex6e5uw3yww8Rlr2A1+Sx9T8htGU73CJ6wKTlSNtiUwMeWWyHIDbWU
bVg56lqz2Dfu4APnmcv44ZJG7u9VtZQhGvMm98AOcaej4IuPMOp7clwBrV0e463T
gN2kkSi/3Lq/nOg7wsGMRxIUXYZK6Lf4/7TJTFdRTPf6XlMd7BfMT+Kukf7yqsBH
F/4uDySVSSBgeqB1eW7AZVTA9hIJVdirAPbhCNXIU+DzPRGDBsMN/FnKMrVqQXjp
lfyB22a2lLMp8zXQbQF31BsPxUFHPg/ktCsXvpw6iXJYThX5xavSbQsdRR9I+h7E
`protect END_PROTECTED
