`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GzI6xtbBbb9NriK0L9ZMi5ZWcbvDyCag9m+jsCD9swEaG7JaedcLIEQ3XB+iA8cL
EIg15fia7DiXB0NuaDbQ7urgdBBrxMFOQrjLYS+r8X6td/iCHwCjexenBcI/O8Q1
n8dK3eNklYlURvQduTBpG5uSh7jBeWPGFzOoXEPr3glcbnH/33ligATqnsy3qnlo
kfm12FAq5zPrmWZa4Gzs/FcNCWJ6oqnNU7ym42BJDdLd9HRs4XKZhTvkv48ICy1b
GOkGy01oalVsdh4MVWknNuUn4TgSw/pY5u0B/0H9SqZzN05tPpWr6x1eYMbXtkPM
5OqOLQnLw68mYqvb1fd/XT81nI69PJF+W6OJhqOPXKckPqrNH8wvcS856ShvAFLF
YWyHLkZQOeWxkBtJz9Tohqne/iCsL9yXhqdzSuY3cd7PU8L6D32FyJNDJ1Hbw91L
SHM6dQosi8tIhd36SyJzyucVaxLIyjr6Q60NRv6nHE4Y0FTmYKgxpmHbwZYofxQx
e6X5ZGNKWMuGxzcItm6nFXzPHlzUokoF4/Q/YvQtjoTM+on8pvil+1XwH30VGyLW
SnYwEUsbNz1dY0wDhDPG7wcoAI/hvueSeRZ03qNjLVaJzFfe/m70Nx6Km8vGvvSG
RydxX/h6tU8NksFVCOHHxmxegPbCx/QV1hg/U/O3Id3AijZ9hHeN2yR9mRZK6yJK
dDjIc5vOShUzgBeB5G/4wihmR02Ln9o7UCWiJJwVRLh5Ri4M65SzqNz4nBZZAqg5
6PoONPNQWM2bXBuES1+yCAQCaMB14wYQOG9Bu54rZzHWxao7CVnHqGeUAkGrFrQ2
0f1/lNhGZ1kXdR7WetGoIqltkVOqrY+xyOWticL0cdhalboDoVitPmYF3vkRzzNW
TkMgNivHeaXg2ji+grKJh2Mou2anAffKqnebpTOWL4cHuZb2kx7H+eVWhOE4uAs/
eF/J4fQagAHe0hsCxwyWZXUlE3m7n3y9nwvqeFHH+1NkONAse1zgTHlIV1U6NO1g
rjTfMSALTMEZSuADgdzEeo60TmjyClTkf0q5qXp9LWWS9N+ivVv03/DKJcVNtzVO
9WUw6sigdUzZ1+1zLTzCb/nMvrnuFTlFuBswwB8gwEnu25Da7Pp55Cb4HkUgAVAj
AD2WwrMjzmVqHNwVxGwKzM1WHpHA0tPst3/h8zJJIybO+3cgL+w3DPS+iX+NWjI5
ahRnwkfFAYTNAvKt03aK0S1eqH/4omWqDNO45iX/9rCQ9gNaEzFzN/96nTRNllMK
t4Fc9UuRRLGwUP40MxuKKbrmECg+wwNnhnueb2HsLKc9IOqcsgmvbf1Xy7RigRhZ
jjc5TjdKWR2yRaqpYHs8WRj8NlqgdmISqQ9azpqjfb4wlJcw8Vhc9t/oNduxyZWO
JoiHF1th1aAXoZuYgX6Wnb8Hw53uKhHXVQC7lXJ3ukdui5KTT9dgpKAu3SzOZ71p
n/wMo8xZ76X+92zHQxSy/jU8vVMxPFY+DF7oIJjerSGzrvuVHXHznDNQTDelOerB
K9RvTw5KEuJFj+oMQgVijD+5RxyyI1Pwug5GDlyGoD8zpFKAmDd6hmDTVSjDdedI
Ql7018zpx8JRL1khPF/HNdZVDyN0/5PZVdBsvx9gkWzxE/Hl1BNydUjCw3ZRMoPi
0TAHqQIs6O0l409voe7NGYPJLxmIE9JpgF8ckbAG/8oztK3r605dwVf5T/JW2ITm
JE93nh5UmEBrmt31FNG5bb0kBEB8EZo0VNjAl7M+XuURnNcngUx50xUsBt+dW6Wd
z+sJnmC+iHwC+LrX7NSY0D8QtJbmyT8EKpSbevC0Gb61sFydTt4D8ZzxnGZ4VA7u
3Ud5JJcg5XzuR3EQBM2VwJzM4WhAsSxiEbnuYcdAf3x6boL3BsoEGOgL4IbbJZG1
AIGkBUCJx7cUtBhihvR6LCNbtH2+yZr7E0+kMrKJTgE815PsNfazs4mdZ+nr1t4U
a6q4J+VcjD0K4bu9dmHJNIVAoc4MXJOknO3Ri5Su2uzIUycZMTLxa25cmyGCbCQV
uoh4chApsBM+LaLht+dTFzr5eW8FkqChpN324/1FmMk5VpSBqUYXG2iCjyzRdPVH
5VlAjtzs3k2e7EqZehil/SXANKDHh9gtFI1fiyaZGQW4OtR/tMNdU3tPADGnh7C0
x/kmTsBhtr+TjY2p/YoZChO485WvkieE2M5gFOhJ1mJTTdJSVxUWJFEOCvh4sWYP
pMJ9kQhO9qNS2Rg8FHVKhl6hjyVbb8Y+9ZkqErtGfRTeswzbDqA9cWgM7iSoBFmx
oXwaOsctmOPBeDlC0oLjaxIVRQU0M0nhsJKNrk7s+7xJxOYb22SAhQtJqsvWmg//
/waX6OG11AzLa8KxhtcjBC+RSr2sZoiRjk/h70UBkQ0mCY3IjTT+moExVPKTO79F
7xg+ctoj24i34UV4uGFk4e3lnU2S8+HAzxFXbP1eHBcD3x89i4ZGtE3M/jLiZT/P
MNPd4XRo8DJ4mke5hVb3HsujbM4d0cDiCN7TGA34kC+eY+t0vjvuLqH/bei0tuN8
pK+lrODYf0Awi4q0Am4FnQrtEBx2OY5HikAKI955+GUcrYpVgIfGolsDa7q95qhW
bNvvSUrlLn2RmzkVljSa/Bv45XxwIs2iNmOlfka5/aIiVLD4PaB0XbySvw00yhnI
0gN9W08xlnfPIZfoEwrNS+LZzykAeg2S92vLwOCc8OeqhdX8zw6SV2LTkL/WhrCR
Q67XulGjkfCaEV43Hg6ySmyY9YmnyToB/dWw7kkObUaIobfbzaAZHh0PUVf/8ZKf
kM+jMBdv9ODQL7dLLRrvHswWjDH2HtamKmmY+R/QAxKsPyfGko2qVwgrtBv/5L5V
EqdLx/hradMAdjt8qT9zXW1I0Co/PrOiUD+LI1H+T/9LfA+bb/reYbF7ZPtBaVSS
BrIKDfroL4FJQyYl5CkwVCwq4/z7kAeZCSvH/oMkpJHlrcbA3YG8DfSG3FWvgGEb
3HSI6r07m5cDn9hQ8XitQrzp1N6QBXl/ZaVJ/IBqDDfOzU3WLsG4F4NcCrxm64S0
Z4FgYgiVZUNrMEg6QydRUGmKyN8/Rj2ICb7z46PyAAsGsZjgRQFrGB3YFYa2PrFh
BkCmdz5vK8gDutAnDnIpLXZAHEgONhpBjUh1dQUooeC7W2eIXSrYzyq9vQa8KK4q
V6qLyDl0dAVvsLmGrYZGcn2tR4nwldN2GgiuLYa402wTjXiYAbWzGELWe3ikDN3h
EJl8j4r52vQzKL1utf/yxoy9Jomw6LJzWEZ8ZwRLnHr0RB1sBCOyrz0MfQPI5mSX
QA/lDpw+MVzl9O6L2Tr25fm94FvEjv+QTPcq6zu1QQqwcGD/ALefyA6bZoUlZFGZ
YuCeyZavmD0W8gBHh31rjgyZbIPCY2/Irk4BXKTiIbwwuknP88nu20Gat1VLe6N8
AJpKxRgM09UNJ+eKJUN1XBurBgv1YomQiFdRtd4Z7qkt0STXMGEHTKPYA1arAChr
axsDzYhneyTsut1m5dW1dfgC7zpTbQ86fdgWw0/1iT/QQrvzVSvYqV8lP5FjpnRw
v9J3RSvtWuxkvuXCTVB9+urGfOfeQxKyGjlp0bP18u9mC6Li27z0qRlTOCB+PLJZ
PAxLEWWCNzeBAzezNXLomrRgsFiZv8Z2EqtfuUJHo1Z8oZc5ipxPGYrXXcfC21NH
CHyBJNh9IZIIRn3Fs3vgvhgynOUIhn4GIGStqQJhgrHxDzUj41kFo/LjRPaoLJ7M
oHHOYIrgvB6B4QJVDwJFYIRCJ9oS5HzPunJJLCfspaQX2mdXAe1oJx9Nuk9Vr2qU
/k19tEaQaCpum7BQQ/5uYJQKz+vLusXtfyqKDMOnd5ySnFb/yGZaP34ER8pFsFD5
q6tpknq/DDZdamUurfarn6pZ5MHOgcKWsHVA7AqwMz0NjzdqyhDw8sNiJoZ3Krgu
P8ji1Q12VKWcVqHOL4QGkDkKgBic50X4Htf6v7uP+LnYqsEWUg7mchOvgwkySBs6
uw8H21LfBCs+hVZ2G8O2OKWlDLVImNc1JTbNz6dpRi2t6WzyZlNNLSztn57IsnXM
6/wy7cA3zwR8U1chVWMjLch7g6irPLM+MCCkXk4bvvbEFUMpJYxVTkvNbYGWhGk4
cHAIBqj7ZCCr1f6SuVBJmiELJa6gk/Y7UHJSZ56VtWpjIDsZFOw279RSgif15K4e
FvQ7yu8QqGDiSA0ixs34k79juhFuy4p/2u1vZacbh/U2UXU/eNxD19LU4r/gsoNz
AQCqTVEiU8F6NRfBBTXUjqvJ+ZuLHKi1hwRPgRq7Rvoi61o/I0nmUsHfXQUqSgBF
Q5IrutlMgWmfaiSw1b8+SuwtETUYQkoPGiRueiC7MEVZPspAosm0OkrewMKUAGRV
WihWOjlRL7s7FOV2r+pBD52GC2X22s7t0mo9HaVGh73dUgildetLKHIVKjtAJG7o
dr8qEbJ4DO9yuufGrEqta3mp+bDjzmfX0GZD5nyy2TXBjER8x/f9sPgqBzeLRoZz
ls6rDZ9Zzqpoak0xOm0phw/NHIf8zeGoE3MyoCIgS2RqtNNV1EYZqVg5qOJIDXut
Ecjs8HwdZgNYJRMbZvcUrhHaprEM4t0vf2Fq7OHJZMQ9P3lxoUTLIpicr68cDdFC
xWqkg/M50pBw6YbVaeHrFNQGlimVPPfS6+jWp9pQvFaVqf0S4731EIk+tjJdagyW
vPBHHw6IlEi1NvT5jbfuYvT5MMRnmn6OEV9PS26uq+2xaGt9eUP3Ra7SN2UI2/bx
5nEVGwtzPwgFXKZG/3aK7rk0aV+7nSWC1I4MX8X87t4a5kSaywE6kpdKWAUes0Q+
h1DSDvkqEiSPmhVp7tn2+qivIJtZFkzcexrXFlBWtkyvQpJ7M8/Ha/02SiIdx/uH
1Zj+OIVK2eKqsos4xla/S5DjQXzE/ef2NwoyIOu/utrp1mVSh/gx8jgiXtOx/lWf
Qk7rI1ppL9tZ8NImTKKKxWJojpLP2vkZgea39LY05N0VJcXgEzBzmnVCGQ3RnMNv
`protect END_PROTECTED
