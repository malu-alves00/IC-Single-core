`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3ACD2EfwQjofet2YkN2GRajB3B/Jr0s3NSQcQ4Yu8I9hogWoHscDj/2NxpbSNkel
znFaKs3mpDmo0R/0qJiwfTECH7GtTbMFs2fXKKY8XIYHCMDYLZJHopkwA0t1gUOp
wnhd+cCan2oqVb6O6W96Wx21xjgbqm8mu2schhsqznWsN6E3A/w+9jI4akiZI223
`protect END_PROTECTED
