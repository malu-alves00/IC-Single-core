`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yTtAMxremmq2OM+P6NB9sRjdU5hYJKEu76nP/BMryjALyIAio87EvrROlgxkbEAP
5Q5bLvfkH1/2HOxXD+93IDnf3kL89ebQi0lFG7tTu/euUDNevylrj4Y3w6LQrCME
3+Q97QNIhf7Mx0PoJJthfkyyB8XTeISdeopQzsBsLa38AOLSDv1WePHrCdTsSyxO
C4Cp8jFUXYPLhw/7pcwMAivNfq3mEbxm5z81dnbJkDeTbAVna2K9quywpc3XGle9
9kvbPVmgdrK6FId3Fklc94kIUvChYNBJ8CCf17Plj4q4x+Luow9mq7CGixX4Ro5V
hg0Bq/Vuzk4cJPBXB4jue9nTe1KHABVdtGG9STFgxPd9aeVMd137UE+1R/BBO591
/WTmVjgeV3cP5MDS91Htz+11bUu+QajqXBDT+ic0Vb1pI/JydEPOzjQP403TKKT0
8LzXvxgM+2/KuBlTUhCeZov0N+b6Pdm8nzjKlKKK3lV8ptJTTeNV/wumDv2nCp20
1wiijAwqfjMkv/BM6RodXEtgy/7/srbuTve+N41DHTROAz+pePqkuvVIF5XU/Sjl
s2uwNlUom1nLD797SYInIAhJNC2LEvsYdSLlk3K7pncxG8eoIDt7QrGyEEYnr2OL
Dgu9/y+cSVZE8PkPowjnzKhApYeMEFmEggvyOVSbsTOcCpwIdUycpXvk728n4P3R
zpaRWBNSQvHVDnsuFk4f2/XpgcPBqB+V+MvTWz04ozIFrIWA8PRZ6UP7rzbxxa/J
c16kSi++/3bfJBSJie6qA4LE4WsxRV6kSe8S06AqLLste40qmJuVUx1JfY9269Fn
9W67odv4i+fpNLq0higJNvOONF0TrL1riBsS34QhSMham5AWNdk151VwIJjOCVlV
89UlL7lQad5H9PPpamgskO+Cmk6vIcl3ttqx6sDnAxwTA+ehRQy3eNfvmNZnU5dv
oMo+YaKCpJYKoYh7RwXoEAW65XWY+Em/+AgMZxpdQEz/rvdyw6Rrj85Zg+IQUK4A
ZmMIhuwYW8r2Q+lxDHAW2ckXKY6VRatB667ycqxoNtxLvNUWk/sAM/mA5a+c2I1u
5pOoIhzMFJWn+tDyHWYU4rBtgnfgJFpnqdC7mF2V1J51FXf+Cmmrw0WX8YtkRddq
9uGqHsp/iIZb82yIgJRSsS+R1elyIpJvGzK4ULunRQP5Dt+77vuf9PvZe3YXgvBs
bS1f86qhZl/gbjO2CKL/cDh/G9gfSpKZ7TxReZPOqpRUEGJE1WGBq+JbTPLl/M3x
l+I12og8kq7S5vO4ISyCSok8mx4AfnsZRgJ5M5ZDIdXBaXsqnWB/sXhpd+l1UjBD
EiIJ36CPIZnq2iCJPkq87zNXo8PP1vUZNMVXhJPASR8UL2lbu/D24vLou99Vxshm
uWSPoZDUttXLd4msJuLjSNF2Zc57K1fU1wfEE+N72cqLpIVplUj54PGWpIgPQZe6
Y6SaDIek5EVgdkb7ETx15ekUpeGysWYxjU8P+DOLr84+nsgNQk+P9VD9Hbqvlb1A
lY5vEVCYye77jq0oqIJyc6i1riEvEn1c0Jt6j8dewfLTFfCzhCEqH/YDz9KTUB3n
unu99rPb7YhjGhYEuyl5R+gSiGxWspXE0CQ74p3S4QK+kPH9zh5rb7h3BPT/+DKQ
9qU1TtOAqITal7qNSQywcAGMIV5L1ibfjcyAjDz5nWI8qUTmYW2O6qpcXSUX4e2p
iGBVYLyi91mb6jFn62BYKD1FcGel4qLPS8Alti30lK1K+lIyaDGImS2yaRr9OJ33
VZYf8GCSLJ4jxhqijC4h8Syp8/fwD4MiOvx9XFdD8eBUq0fq4SdB1vnrs+aQ4WUq
wqy573EpaNyN/4hiVzYQ4jDkaK/6X9xFlWlTu59/u3YlhkBXjQfsWihqwI5i1jW6
9HQ5GkBecRON5NycgmiX5q9uSn1Z0UwDMySu1eQnlCnIC2kE0NIvfJN5Bp7UWWCa
klO5TAKPy3BeXaMXAgGeNfd3R+lI5RJDy/MhLA3FjX3vG8USYM9BQz44t7hqUN3U
H0sTWFoPYX2TGcG2aynDNlse0Yj1JCE/CYmhv0dyTRT+Mj2UroeGbNH8YBsfZUM0
4QpMWPBrr/wyAQYNxC2QuB9VseYKeHIMzewhJQFhPiFfrbuA/ZnEhFAKJ0Q1tHB9
VK0oXfdJKWsbA+5MlJSJyRf6jUZhMKpX37jT02U3HJi/Z0IBGlb3/hBRbBpBPfQD
UeeCbe2+do/fe5CFFwSb7YrrdXnS72GXUt6pDUdNK2twsv6SF6/LNSN4l4AjRlzc
fkIPuIjJVjbjwyI9NFrv2TAKEBmmg06GrKBj7TA6bd489TR9EWeRwOiVbPMhs8dN
ZuNl6HQWZl+dXHpGixiKEzD+hMQsxZ0tiyaTuTSCYTthrY2bzRPrARY/MXZKD4Ju
EONEs0TTWIzb3v2PZEVYGxjpCQtRSs4db8b61AtIjvW44lJ1ISc+N/MJaYwtuwxE
MNQu13BPQMIxZLXP3T6ww8oyknI/V/QaQZh9CD+ogy3myMmpnARcmmTFOughKKgz
4temSlxYH+yqhwIxMpjMsjFRfQZGlMhZg1ISo2H16GWu+CBjA3ReHh4pAOL/7Hb2
gJ6c2HhOjXEz9jQWxxxfs+HF3HIR/hZX6allRalDIGmrbrDD+a9w9RHMyPtCz9m9
TmTf4YTvv14KQP2+Yz1bjh6GdJJJjrKCgB35Ww1ZsNuvb2vajmFA5r1Raqmz0VUX
YtnAHximvqQZlDvohAnIgD5epCB7ETPNa6u6bYtfJF8PYGz/jVAwpD2pMnEKJGwu
sT20Lz8iGzo6AUT6+AauMzUdm0bNXUQCAB2g/hlHj1CMSm/E9xpcAytsVm6R0jwp
b0rUVlR9DIIYFJqbyj99VLAStPLXh86z/Qv3N90kTvrhUcthVeBs1AYh9ODH+LyC
Jb+qkGpu/4HIj8+23jS/fqFeosNnV9whs9w9f7T/HECPjlh53kPILj2WyE1/Vu8a
VgDczv87NRzxmjP4urvNoQCgLRFBpBpDo7MPfF/lPDk2oJgYE54Pd1Z/QYv2XyO2
8vETx6WMlXuK50exrL71FCWT/VU1HisJ5/767R0Kh3Y9rsaysW2+Z9rtLYKaqYcZ
fNGYb/lfoD4va8qzeW+oTUAfDUaLNt/4fNOj6PIGcP9jxrtcfXm993+OMFxBr5yU
8NOQXfNXhNMX6E48z9CRvQjnOm5alLviMK0yMRj7p+Glt5VqWR+jjkgzfGAlJS2e
pdJAFzuxPgjUrA2JLeGNYL4ONUu8DruwDlXEuM+4tLCV4ulTtKSh1HZB2fQOxpTg
VwY6v/xtiiTMGDPNSJPkKt7e0ekBwMXC2bbyP1oaHU4UY1xSWjkyogdMlWenBKLA
tOmIeyyIjqfE3EThkhOzoNT6fOFjBROfg806oKYfGmJE2b+grv3k0rlTXzR94eI9
jWTl3BAdl3m+qSXhpu+hqGl08fv7tW4KvpOkns1e5X2elf+UiSa0PMhqxT1/vDtD
22TfCfinfg7yy+VLnXIyCnlozyDUhUjilXhj004enLtHixBg+WG8nkTsQwzot3Ww
jqer7HgpdX5o8sq7RUxLttFT/ur3d/uYcrPYERmVtrUHAQXTVTVvzOaamaZugs84
xMNqjxm6PwuUchGWicHuU93+fKUEbz+8v6ljfSiDJMl1vNTk+TvyWOt99h83dGHv
QGOAi5Wm1pGA3YZRVoU65Jup6gdMXEmEQi2gNCEFHMiTLwCbuioqpPuxj5sitDBz
YzVeRgcJWSbf84zSlSLt9ezcxn/bQmJb/w7DbATnzBGpgMPFd7KKiCz6XPa966D9
Ah/VZLIqkxSP5aEIN6QkCEtssF3POZmpcYnKbmPuMfQPHSF7CjBR+tMm+Yxg7I6Z
Gu5wBj5g1zersCUB5iKOz5uXNFC8wT3YHi+QMsNxBr7zZC12G93PuJxX39qdzpja
IsR0KLQ08MSY9r9I5iV+/8KbiGt1bXBZB124fCStwkIYexX6Q3niqxUA+5K4ef5m
L3NoyzP0b2FN5NDcLz6j6DewDh41f1p9ARAH0rlNyT74nKb52B1YpaJ4d8G51Yh0
/5nQjkd3wGFtNI425H6qfRpmD9RxO9+Dt2SwDzz9xLek4Knj+HoVRdilEqav3yV6
bEOv5hBmA3FylCrPtuAuvkw5NCajIPLKbKLoYOGYrkyhCntf75mDFHrjJSxOvsdw
dM7MVw97N5rNUFKongi57tgl1CAhVWTK/RcN0H6DOr1LyWr7jfzGwCzgo7TKm9ij
xnDSiMJyP0E13KFC+fL0SoKlZ0YTAClWJjfQPapJMuAhsuGiFhnsHgz3FiVvoXqv
XBYW62C1gVZAuCXTpD+Dk46quiSxXSHL+q85YQvyQOzAS06wCkLWKbrX9KNy0HaA
RKPObpPD7Apvo16h3oWcXU/IQkcPLgfD4ZL86EAGMgfRQhjtIhT4PjjrLW6j00IJ
wfGpqvJDR7EPvIveDrgizLrkHLKj4zupQ0N/rQg5OKMD0eAhkgbpow+PIvr10CNk
VSz2oUTAX4GUSe3x+MPY571OyHi4/ZRzDNR0/e5YbqwpdF8VWr3t+MFU6fha2+th
d8ifu+P0ywS5PeJZWAUpSkQ2NJvPtJKp5XsMGXhq6ume5uE6h/OG7l7p2U20fstq
qlX2MdCTYwG9s27rSQv4RdrXk3xcgogbapKoXPtQjlyNhcc3+CK/w/+xUWhsBXZ6
41bttLLBhB3OdWW+SeaIzAB6PLH+2CeRZFPPGgYzWB+871Cckt6SeI3UW2xmWqfg
JmFbYrjaYA3ljzHxroCXLXLNx3Wi5Y9pJlp44QppVgLBIxPP/tiVlZPhBFlxyTlV
bSMrOOZsDpsni2e+iCKVDZL3DXKMzj3V3K6ivaAhjCuAOzhq7gNrEgmbzNtVId6U
6E/oyCYPMuhcRxP8ycNeCE3HFLJvlWavdkN7JOU2QQzTUzWtIMn2nmVRfdSscsbo
9rl6vAbOg0sdw061y2JeBvch0VdmnaQOT2pmH77FT7cxgVPz5j3o2F2y99q+y4X6
KFuYVa0kKnldHGGyto7GlJBfhw1rxOPZTswDc1E9VfXGWHw6JSvyLSE4CESQO/ei
CcqKKe/TJQp+72F2cflusjDBkfT98ntJB7dOvOHLGkuxHVnW4J/TvG0UyeHmpQIN
PbcML+iLpRrJVL0Lv4j3ldx9Qvws6O8Yl+7CQ3tcEqddeU+JqxEX1yGVmP0eAjcv
gvrQn1olFLNr01ifG6s55Tve3x3UaxQhfvgdPxEH3HD+6HXKBcdV48h2pYZNozNx
Q4v4yyQCLyptzS4lWyb3xj8sy1JQSCoVb4oO70BVYsw/n1e0QfQcSHNwyifAhLl1
I9eaYjnw/5iHlkkU8BbnbQIdL5BvrLdGkDJISTcyzfRB2wFT0nRBRT/BKjZbvm7X
WsWboh0T1WoJmW4xMs8hZeBR4aixEO5QZP2aMGn4TD4Um289YdXPimjCE1JdqiHE
yzatDFb1n5b17V9XYaGNC/PkHNUnAo/G9YPA8JM8zs3qTkSYEixzIGTlN+/5CAuc
qhnRFvvazqthqnktIYNydDCNM6X0DM1WnW0OfNznTYTGN7AcRm+yJIhd9mFmviu4
m5HB/ot9riQaao8fTsz+auOZMII8ofe4a9WbZSJ70yx/EqgtsB5LqfFt9rNym1Ok
i9Sdc6+4pEcv0PEfUhlkDxeJSz2tm792GvpngowCBN0SG1wdpnzVbBCsxviZYaZM
UTrI1T85/jWb7TQgkHQTkbYTDaaoyNCRg5y06gQRSs7Zt30n97aJqS/ugAvtZsTr
1b1Ff6/H8xBVNaTjWKF3EZbS737sg7v8woeNE287qO8nInclu9fbLWHM1T3BGqlv
hdkvH1g4A3NHIXMj3wZ0uxaCLsyVYZcM0fNPtNWFw/HyjTQE/qUht7cRb17OB0Ax
QCk61XdqbQnHeDR8ZL4emHN/vqj9KYZmK+OWnnehbOl+XA1Bgn9gn4/6v97q61Sg
CWJieuWSTzwE4rYmHDG6ZjOJjwaW8a3Bx+jyTmFcui2eQFGJW9hEwggHs81CFj8r
PvkekuXjUmboY8ce/p0LOY6gBLrVKSZm1SPpN/FWWg+9MTwIOdosg7Ds1zUDr3Uq
bZ6dbVqtyY9a/9T+MdhJOPEFAqGxmVWJigXa9UE9D4tFLeVIv79xYPKuYlktIpLr
mEG78d6TFhnSRXhytgbpfyimkDKLR/c882Zl/wH4rkYk7h4uMHmwGqI2C2DkKONb
pBTfFUJ+LFtCr0lGypgVkktof9KDzdIRwcs0jbyb9dMF3Fcx444txX5Je4RmEf4D
NkCryFTjh1+WLbmiCF14uZEIrWpSqhNJirclylQC1to/WwoRLKLVfaZX4ZZO9kFU
GzsDPCzl4U9IgEQZO5I5YlPCpQdkzxTsbxZ73K+wyfvFbA1S9ekXa0Zt36g9ZQnN
UI1ufmtbp02fFDfkjL+6tIhtcxl12Z2X/FrTWVxcbRs0wai/UCXG0TOJA00GWbzV
i/XFbCrcUpgy/SNF0h4QbcztnqZQHFJkndhETTmKpHgqmpQI8MQuKVo/GT3IZsxm
TvN037guKef6gNou7xBpOiZfgea5aCPYydJLoWq+i1RKOlZzTWMHHQ0Xtqzm5ZaW
Xr+5ZsGmqtao0oR8EuUSbab2gJ5o7rbDiqxUAUwdE9GHyh8pweSCjCtd+rQdQtJW
EoGmnUjznbkGY34Kwdea/UNz5Gt9K1I72/cAWrS8lsCsmnqn1cJm7Ehn/Wo6iSZ7
o+p8eiNC3ocjyPchclM6WAIcH5xGlJumcGZzWzJbLFW8313TXGBDQ1OOR3kD4vzV
Zg4P3Qj2K1k9C2xfxcgRONJpoZapm5vD+KQSZaaHJFIrNcjQGly/gpSesTDTSwR7
OorxyQ63dTtiMTmYghF8SyieoexJyY6/bp8PDe/BA7y1KzvPYv7ld4ecVQGZyAFG
cela90C8z/p73jOseikES3Mh9sRMsqxs1EdHI2LCT89oBYqIUFqMT9l1UzZ1Tsgh
cOTB/CDuyx2hE/UNVFLuHdutcgYrm7dekhvyeJtVGzJjdymB7D4Dm2hvQJhxJbJt
p1HBHMVL26bJrhfkAx2ef1zarf/qq/ZzFpTmhxD4i0+jedMe+ZK+vUomqgxWX2++
Sl0OuiPcbsw6ZzSSchpf8ov5uma7EwhNgG1n2p4OmuhkGAJKHGmvuGMxZODUzd86
aGkFyQnMXB39Kpzzm+uT096F0fQTWqOGNyexQbpmJDEL4Kc1Fga0dfYNtm7Q57AT
rXbOhs4r3Et70c298iDkZsTeT420ymKntTEG7z/zn9OE2Tw0IlpcwmzQ1VA3ycTQ
ct+UX2lOCbBqPPEJ9KQkcln6fNpO5O3TBsPTVHoYSc8XUkwxkIhE19bmgkaLmbJi
GYNxdWxSJNf9LW0dz7Yk+hT5nojNXsfPwuRXwNRLEFfRG8yvIFaJs4kzfRaNTOST
z5gjweICes0h8dnlSHmaT7Cg3hKT683njOqBOXBc40ipv8u9QQ8pZqqg4UWgK8pb
MEShDu6PE7pXeMmY7ORb8iwVrVIyzYtsR1LK/ZOhjjFzhV4CkQqV3hQAr5YE0MbX
vJRLQbZUFaCZabky48zr/V4Vnx6mP5PEccowPyv0rXkXQF92xbEdEz3zGC1sZKdq
ytSv9k8bP6yCnBvbxWiOgclNVz4HUn0vNQ+FMWdc+cUj24nmJV0jLOj7qwEyqykm
45+MI7swNrqONCaCca6PFJqr6yBzRFb7xhNqKbtMq6vMaVM1UOC7AwtCCL53xJux
WRSGu+pmNG1h2JnHaffP4cnHwtm0j+o5DhnnaWTC9QRpv7PAHKTwzR5pEYoIA2Ed
N3z5iY4yudBY9TkS/EszANvt8F+dxMdTS3NqeuqPAyl8/ySADjEc+RXdR/qJdhwT
Rq1KME8VMUag/IK8TNRDoZCNiM+eisVmRH8mVYkDwzEiH4RYc4iDFgibPIeMa3+2
8wrk83avsPng1Ef/oaQy1P27lCIgBOYe4XIJ/6PktiiAs65/2Ncrm5Snz2AAIFqi
hDcX58ME5+k6ND91pdD2q4J7XgR/p5IrXo+eKaXuZFdrhR2lBk9fHlF2yqOuefPc
vgbpAILavWi+p+XPY7bVWIHjwOX4NYgkE21Z3qK/pxhUx512geZ0fJQO4MUKY2/J
Be9r/f1UGc3eLSFb3La5HSO7x0OnUECD1lZxJ1mLNP8V4CornmI9AVx30jLstYAh
KQTqPVc2Z+X95a3/My5NvNrX+C/61EVYVPoKpboKG7EPtTJjXNmtrLF8PwYYAZkI
S76ywWwKGkM6avdStTLocUfxtCAnw/fEkX6fZ5u9yj8P6StQreouL2rnk1us5S/t
iqaYzX5ZK/kWmKdxU7YOusZiK6EZaGft54jzdnPJNJ6GYBU7DPTZ5EDsTjDbu33B
OpMx/L7YJLz9pCm5+WO84GKNrds5XLRfxQYchjsifPjlFsmY+fo+i97PrNPHB2xv
lY4CqWzKw7/ETSwFd5UtAtb7p9V9wlUU03YzQEsF3+V1IE3+M2oUcznMuJjPjgE4
k6NyDeouZX2t0Bmr2nNjhM7cT3ZiKo3Be6D7vO4fpY6biXIFPDO5Vffr6Yoi/u6J
e4mtpb+4MGQjkvbaBD8UfNnRccTLPh8b2G0VWXoPysY7vKxNlN6xivA+xFcvoejQ
0hTO5jNeIY895EKsKCswdE7faNlcxJEdGScrXo08kEyOTv/I4O99GzM3zPOyHLCB
jj07kud3PgyvFJc80ZItDccj11/iFWAeYdodczAwH4KvoIlCXZp9Tz8U/CnNpq/p
NOff1olvc+NNN7hOe+ncfJmlD4Z9BnHO8KptDx8h+kBP0lufHzmG/1U42n5NtTZb
7LlvCpOc0gZ9awkXhkIqa2Wk5JTLUpmcsaA+c8L6yxNMTNEeTjBfiMsxRZuLDiJz
vezfk/g58doP3+LGHVosPKSTgO3qQHmX776Yd/2DHG29t3srlDCGO4wFpPaPgdkd
Tba5yVpW1753Xz4kXDmYfNqVVsJC3XuU8ISxJwVGSeKQO3PCIQIa0zjXQNNLnn0w
0EIAB0h21O/7DBVqcml1QDYY3XDsa+tyr21TGr6F0lGlYnbyoTq2AYqzk4HWgrK3
KM8EVaR6vadD006JHMshVlLn27VFHMA35K28qhdktqZKUl74XA5iKOA8vCI4lNh1
Z8kRBt5gQJg9jAG4OImLTfSYIbYhm29edRqOLrapfzMcVeFY5gPE0m+ohmkEEVTf
+Dn1DH/izMTVMiXcR5AmjUd920G9NsPj5eBqyW2VdfCyXhopf7RoZe1PfptDeylC
RHBfgAg6Ee6waqZwi/cb0qtVdNRnCbeZDnTjo+aRIt7gmz1XvZ7VO/pRp4y38us+
NPQn1F0K+uwn3xB4KDav4vYL9Q57khnBKkhkvnfVsfYmvOLDTQKa1mQOy53mXFHd
grzqabVcCFmdpMyCZTqD5WJdR3xd+/7OfheRiQ0tvsvppBqGxWtL5VsfMmn0ioTx
WR8r3NzaJkk6yyRwdMvidxbbEMAoThjkRjhyDizRv3/lce7nKl/1O/DjTX2g1f9k
5aS/V2qRlN+KXTKuvhgWvcJSeVSsDhoHogQY6Emmtip5tWwcN1SEFF4i4VWAA0IA
jrBKE0nb9SaftELGjY50JX0Li5W+XfkDmP9lser/aCkptXuDgmLZQH3cmTyqMPQX
ce5zRLOPGwY6lbQaskhG5kwoT9Je3on4f5PJVGpjbXVVrW48qinH3xw1H8W1Uoy4
G9ODK7vX73WHnpNoeiA7Kb4+x2d6xgFqWICGCBV/QbDQfitkyGUDClGC5f6F71fb
VUfyZTah6a6wtGsVTQs/yKHrFxi9B8MYMyoFvamCZ8UTqpbaf4RCXny5+f1yFr21
GVO5acwmbRk+phfqQkNAr8omyMInyrbZMWwbzY+9ivz9ib7Qx2iGdUpy/1ztnw86
za89LUf8LPvYHZ4LyylXxRDDPVAcNQuqvHKDUJ7do8WmY3OAi5LHo6j1e1LhkEGP
8cOpwm1fHjuEDVnxh59vpRDdNymA55y+S1vkWoaEuUOYIpoVi0G6mBPN9hTvcQ7b
F+h6G3EkP6QsRPfgUzcL/JSdQ9iwZymE97eIVXdMJAybUAQkCDHvPn0wF33qSSus
2M6YqWtX6z3yfaGg+JQ8DS7UoQWsTBLXSNIMqIf8EPf+AT6yNK20Xt+lwamClPSw
SMJR1HY7oql00DTUPh1Pi+Z3E2ljZiQx3Y/2l9lwws2ZDvHSMg1wVVOdi2+o0ocO
M4cM2IHv2XO7/aXLHs50D+Dw1arKGaMdxswLF3/XcgwMI7vsSnPA/vxVCo6t0wJZ
7SxSR118Ppk8wuO8BoTjKQIQZOZsXn0p+jzwdy1OioQkVC80Tf8tlNIwbQ7zWfx4
K4l7hPQou4Je0NYIMxq/82KKRRTrJGfEHn3rDGIcpgjTNj96qAdT88oul/TQqDKI
Bec0kacQqVp/8A/tE6JM7XeWI9uOuRQrhRKV4T3ZR12NviIiBJgiQj1In0Bp50Oa
cpfwLTwWUu4AGRwczl/SqCdQiMd1H/JnPHyOaX5lmRHUZC4hUe6moUqJ51n92pGH
ugpUrgHNFJxhfbGtYhFxs50TH50mAvydf0tdXZIQo1339JG5TbabX+BVUvnXpFgY
tJAMS42rIIjqCfxOP6YWSmFyPfSZ5esQ79E9zVEhu0cKBik9xry7VA/hqa7WLL8N
E06P+rsjtJBaDmpZEOQ8oa35sp1Ik7s9TdDZJUSRnfI4hYCzKWN9A0O6LUTs13rD
G6Mik4cnZEVb8HCG+NzaNiUrTA5C311BdCkqpuTzHJ2w9srGR1igGJ9e70NeCzqq
FS/NL94UWbfjiAAJ/Tku2jDOx8qqPBc47F9rdmWoHOUUzhLtg7N5DD4+6YgItNaT
57CUGdJ7CBlSrGRKxgupeZAxlB6J/rIQIZGFRrmpPDM8HJHIJPZQH7KniK9ctE/3
GvJgdjFD28N3hJxq06sEobb2MLiV88IvLsEtVCuD7NmomGeFWF4K/2jvmLKMK2R6
E8eVQViD9hENmnaHtxaYnZBqveZrCNP4dBC6FEqEG0KkVRrBSBtbBCXRVZcbuUbH
L4SjZt7hRWUUVKb4AS5+ilH5uRA14wkd3M/Z1lwx/Pjv1T3/HRKwwMomSo3gDfpL
/UrK2G7f+HZXEgMCcC7ePUk3ryq9WVBBeJ/XPP/2/cwQfbwmEKQHFLIU+jDqK9rd
5vFTDsPHlY82d/Ls6lVrpPl2pfljJzOCcQ5p6mENrOh28jYWCKYN/W1o3u8XWceV
gUqqP76HTsPSlmJfVVnsFuQ0TC2og84ZSrAnJIhbb/naosOqP4XL5DgDe+E+OXrE
vPeZrZ7Vd4eJRADM6E29DGeJ+VcXPO+QLjC6AhyV1v3P9Jec3znHJ7YJk5YzHVId
z2MnqPekmh0uLFJnjSRg+Kpbfm8q6xkT68XDjbuk2P8HImRLUhnIce6XuRZbRonS
Cfu/ABjsbMw2ZfhJDoRn742CxhRGl8jHaJF6HKveRAOUORDlFQjlx9EeahsGxtv7
r6La7pNUEIIeOIvnK7uJ7GKL7gcr1PHLjXNv+ikFjrKe+6IlfHThaLL3UYVq7jgv
/PmdP8hO8QOI4WkWD5wDcxRlXlm3fGKcmAXDn60kuh1dzycS93soxeguHyZcAFrZ
OXT8p7fOznBaZ8yHmdyiV456qRTwKwO40vnS/jgDLoT+naa61/Ka4BT8ayIfq49W
emzDdLPFEWffEejQiwhm0DmbIqjqkv1kGHiufvGifVVKF9S+9dUXRzk1AEOQ4evK
P5Q8NZqlP17GX3IpL9Li9IRzXWt8B8NryiMFWkJQp1l2MgXSOGp99uw8U2U0Pqh/
GPeaAGb17Q22CbIKu/HYYpMwD30vTdPQmFZzNifPr0bMIbY2J3ifTGBOjBcJD62u
V5JW4ImErN++vgI801zIRAiE0iq/bcl38uYumIegHR5+RM5ay3BTM2KSndcnoYHl
y2diRK64YFbZn++Gz8+lrV/5X1BcyfVQ+Frb6m3U/qXJYwhYovb0vT8znyP+siYz
emGJ8V8W5g6L/hIWjFyLmLnCtViycmgbd3osmEPKFj4kesdpfc9KHDaOeLBxRtCW
smWfs7mdEbTrtVE3zOzPONC+zQhZwDPj2cClA4FavOm4pqCBb7MvJ1Ete/UZSP8e
1cbvjzEr6aauk5phDW53aPKbXWLEwA1PKXCDhva/WsnEK5zMizooe1+efD2/gcz7
qtLzg4oCSmaDclfuw7o/LRBx+RZy+poannCY4UUzkqkYKlbknUd2Pn1NVC/WJRqy
7Q8BaBVnUjlBIRxihYoB9Sgjwj5epeBkQEmAkAxBxuOZkLG+vU2Y4VEvhB5aldPP
aMReXSh2NVzNuHHTnwlLfa0t8LG1tl9kP0BPdQxTuRFNcitJxvO4djWQf7D3ww/h
marl1vTuSeH36iyj1HPNXIJrTyQ/sA0xDfQoSoZmwZ+bNLabqx4+2jacG/IIdfio
oAoA07OUSb84s5q+AJ7vAwvAA7aIUh1i0a7fIUhkF7zFiuUVp+RxIKfqGe5aqfVB
NjbrOOWFPOla4OzUc8voBc29Y2hMYlP+U6KvlWeWrh4fTTprss/IEQty3hyZns9r
xzXQiMi8XQWP90i8MJM0D1VNI4IY8WETRFq4vZZczqZ2hZUO6PmdPD0+t8nQEPXt
RsiWkm3qCXPgvCVyDPUsfyrKTUqi5JIWgY1p0366gB+fF2fd/ebM0m54Iva34A8F
HsoDT2c0oqHezLgCwYxKfLNpxryviTcKSgcZWfzHYDxFvfuiTauadDWSwmgLc63Y
aYHpl1jnXyOBxHGCMFcbrE9LOYU6B0sP/iN6w8OSuBwpa2NM9MLj9mYSpCIhrYxp
B6LcooFbP8V5Oc2Bly63+xOH+wmhQ6abH+euIwu2GeIUvEsoZt5Ju+vMKK6hyvG7
iWKiWZaEimVm062Vt6YfP1xzHGtMjj1LRGh0pI9DMrNx/rxFfpcHII81zKNWH3WF
kCXWrGvqi59ON5w/NglThKf5DUJBQ/koQGmKAxGxOgDcPvB5Bh02kuMJmzsYdCdP
2sDIrt75b5NG/KR7UHtYCabm+NipeUgIaA+6Y9H7CDVkJJschxg2P0Fj3Q4mcANj
bA0gCJkbr6bcnmyHoF4hgUVbuk0dHb7QAXTZB2+2KORPH9mI0OI6Yyk+dTxTXFO4
3MAUwNu4p0c7vKGgIgiRUJ0Gz8pO7illJHR52LRFwZOXFLwatiWqMvs9HgrOIkZQ
ta3OwNu4Bij4HxGyjKKlK07UeXm9wAhgmuNtgHSnNp2kH9acc38CiXGzUhwY2AeL
LiEmwJdTkaa1Oxuh4mB0jI1gFk7AvsRBiNRH+K7iGGurn6aTKJRuP+W9B8cor+JT
/zjY7exvLBCWPjEHu+/t4nKLrMuOjkJKZeI8X9Y9MlYv17QxD+7K+1va8uGP6ekj
eBK3DHzdH3JmMefg9Y3thwWr3oIPo8ZzMbeW+FarqoJIe7GdBQdFVMcsAnRINBGK
j0wufkzEOiH2yfsCPiKGyujOXr4XP02wycFXGJqgSkamddTu6iF7eXidVmcFcCdI
3S+CKxZgGzNexyb7mNgbioUVgWcJhJ2jRCS+sO5IG8om3pyajcwUbgLJ/mtjMbNs
+Ie1dlSQynndayrWoCdTajNbL94QLHcugGgIxPUP03ELZVuSqOcpflH7e+vsUzhA
T3q0sKJvpUQe5Nj0uqS4OxW5lGAOotb2zKeW7Q0MvSZxaXr30VFkhZWDY5MUcPHk
es7ggGbeP0B2ElDGbWNZAvQ5uHWIATraRngwPlaqYeC/66KTeM1/sZ67UKZoGrBU
ZMQer+PBW5qTsRDPGXf/h5dbrozMShNI4QoNOECFHg1S9z1plYCDRiRArcROlYAJ
iiio5yXlRz2qRBEzCtFvIUYQsfZVZuSs4/Enw6T83CBXTfMXZqBM4ll3mqKhkIbE
r2dj8iu6D4vgb6a0uRTvK1Mp1CAZx/coU5TejnzNe2iCNounak+Ccv+eca5/TFmQ
ywiQlvsyAuCdSEZZxaJcHtD9aW+vyHj14G8fcgKTV4A4GXDjalhJhT3hDN8vdDya
786BynLt821q93nR53CB9ndeKlblgD+U+59zTpaqR8WCRmTY5xQeAEbPjNm/Gix0
Ecnz/6sf6KNGRHww9hkIwdaB7kGxnOE/mwyiq+W3+mQ7wxOOnKC7sy1rJlzBa+R4
0e2yiMUB1clo0tsKla7REcI9B+BQ5HlpsQfzTwo4Z1+v81Kq1nOZYDIHrLtepnty
g7mGH66SzJihLl8FUSWEHkOHmcJQ9oEaDNHMb8X//T6vsa0LPudyGRi6cainZNJS
U+3/Oea3nwSDxAxO+jflPBS8/ojlXhbt++mms4Qt5QXiI/DON8/yCh30TXfKlMwP
yKnW6Ef1o+pgM9DrV5957MMioH7G4AqIOrC226Dg5CVCmPXGlh++dTqRCq2lcNun
CMSrBa1IP/C/MiQyJaY9ePJBfOaA2JrgU7fCAlPhfs67uf2fmvCSJdjp23NC3MVj
7OdglTDFmnJZVTL5aALLeFxBLX662BsR7gdDSz58Yx51bu2gzdvggUpAwMImtIGi
Wnn2AupS8/xXJIeNzD3Q7ZIPvvEOuUaaAj72ic8NEjBX/KiJrwFDLMzqC297x2Ic
S7CEdYrAIQs6u87ITxbUyzd8W6q9Ud0D/oVyp7irNR6zdD2VraVmiTm76XGSpdOv
TGV568WGOv+iCTpQTPlHPPJe3FMdmz8FIgdgoXLyPM5bNWoQXcVqBt2ymvl8xq7r
W/pmWZIJ5AuQrsYjbx7olyJzF+43CV+vI0SgFVWqhVNhvyKc58lT6djOOAdeO9x3
sy8YaVQM9Rxg9CSRBOcJonQCcfBm1AM+P4To5CMJDa9y6T8+CDmfjrcDendhAW22
1Z26/w15tVqwkqlpUKEkLheJmjM3kxrXVyWcK1TsoOurmyI1KpWX10UpsfM4Cn/e
5loHnqTDsARSA6YzTGhtMw/zdXoCqDbYx4n6CAAFn6wH2HA/0b130W5Hi4N7a+O3
9y1H4iod9eJbxBy7Z+D7kDZDO+rl9D7J7XWRsbnhmdVNw0vU12OzLAzmP5Ig5DpV
dH5j+cjzDvJn+KSpaF3mzZs48lc5Yb6boBVEWZNOIKG5NNhZWpzHqUIxh4BhVCGY
43H5BsjbRmv/XWFqgjyyQ7OKkE3qh2l1ZF7qgW0AIVjkxmZeaiPxgSkcqpALiUML
uiZJE2hEMthzTp355Y3/KtsPWMVoNk7wgzsn/qXs92K/gt2t6Yh5Pm0cWGY26/6C
K8zqcPy2UE5myss1SoyiuL3nmGsA9jhOAHFuPYOoMZMnnqM4h8Ujvh6R1O2SryS2
AQ7gaWbuEfAN+5nwxb2j6Jb+7bvVBvbUCEvZR07sR/Dnzg2mUwPTWJf5m6wmKeMC
ce48qsPO3NdyqifwaEUq5PUkKz26ObUWpqhQVdXdGAaHGP5emtBJtAZl7yRV/yC+
k0c3EpGJtiKDZNk+upZACAoqzstQCyhuQ2acijdbw2rMrgzRlWMCuoVEqF3unDOi
G/YNyVITxJy+7GvaXemqX8JoHXYJ94DU99vhhEN3isA/weagSTuDg5z2zXe5X39E
hYYiMqwfoZtDXVvv+AoSf7J08x/WGZ9A+MjmWeqpXlzYYenA8ueqDIMx+tuz3aID
uyI2oE9gG0qV6QKt9vc104Z93k74qtCGQeL07OlQY7bGPblctY0qiLEoDY5/n1PR
G0faTWSoXJ8beNpZnnVEgIWwszCTVG/4IhIi41v1vVkLnxdggEmmbhELpCk9v4cC
+YeoQkLwWoMwyYEirjII2r3qIJ0+eQhP8Vr06PQ+70IYz70kXV/qRUfXCGfHQrQX
jJ23C/V0wPtKM8SN/xqePg3NWlTGXS/x2oW3t4/WS5W0E9SXJ6wy+4b5E80qAGfQ
k2lAI7QmA0H686QyMD4ahbXHdT1SPbLzDiqp+A+s4IUFkmxjJRgCSK8t9CsaPT1k
Q4I2QG+l2BBTIXQ3oqLhF0MTpnaYt+SyJpgp/EaH8PI5L7p8V8WFA8bARkAfqrGN
ErJ+6f/L5XPZbUW8ufHRz8WogpDtti5IZKesFRNRXoqoiEwYYnz1CQd9NREBeHbK
lQa75hzH7sIhxKHUQnB52vS/BNmKCASGiTFaKMqvzRpTT2dTTzaxacP+Mg06qJD1
ysj3o0RXLAw4xxG0xkVhOfRBiW0lYra69o5QBqGi42stpehN+uddt/V6INMQ0GsF
AwKR9Ic5KCHwUdpNWPKnJgE+VesoXXl6j73Sis3VfAZyxdWj86eftX9gJBJmlKEQ
A220+X37mOJkf+FFNyaqX5OX+9TSEE3M4BHE0OOkfxcIraXsNNJihFGGqC1ABNEA
BcvABYHcII1C1f18DR/8xCG/IiNyGEtQM5UJOgmRvKPKh1ZoYbSXsUB9CDeU9hgH
/NjD1YgfGLhXmTdFFLbKmAjGrye1kEDjQYwnBIBEc8e/ZNcCHc4pe+87rrK6YMB3
BkTQfLWPGh6Pa9v1LpuX6PLyQgrlzJNh1D+DSUAcsoSmRbEmaJf/7lYQ1zb5FZQs
Ehs04VtXLsLivN89TeX8A/4JAmHVTJ6qohRY3kkSgzKfdZtnvSJO2NEdxpRlVGwS
gNeC0cEJHl/qMwaN/N5cBgq0BjJEvnUwNu22+FXRhi3g9Ds5ZuSrMl/oPYIUjd7C
YrZHpsplBHxJcp9HT4kJHK15XT5JQdmSZmtPbDjhEobnAuGSVe1hvqhD4E5D8ita
RiZcJ2yTVEj9Yf2UF14M6pAyZTlk650+UD6/42k7nm2pFxhgoDf1LzSJOTjNIN4R
Z0FX+8jLaPYINoy9NzRJQKn+cj+NApuFR2ezEIHpz1qfoZ+E8mlPxvlFfj6l4seo
Rp13WHsKiWGtUN93Ksy9eFLKzUV4490LL9MzCrptqlIEjA5ltafIXXgobzMjrUt1
QCEJZtEzqGZh0zPGdplVHG3HBaCG01vzjhuAwt1p74WrQJtQ/PlP11WSQeNVa0jU
KOhA/wL0oHpx5etleNBtJzFvtNYYYg+Hy0D8guExNaZf6JZdEXm50LRAOvtPwgX8
KZFF0nDLKdrbCg+Z5fTuCu8zKDVujNiJBpp8+k54uXEuu1yDZXMdCOyzq2aCfCqa
a5IKPvvO7xSmCv0q8fSJHIJsixuUmsospOgagIQYUGdISt24DfhkF7PJ1rYIYL3e
drT9qQcT+/riUsGtGTlw1XbIw4soTtIKY8sAiBnxbeKe7m2o0LvjRiFn4lg+ttFK
OJFW5DmU50z1xtTmyv4M3g2YXYA5fRX0+HHTqxiqVKZT5b92gNwoV64NSFuYBWbz
NzB0ZHmQaezlRBT8qM01zIz29iAwfGPJ+xvh+BkWtqUvTBNDdAc56RtEs5+U6ikq
EaxMzqs15RTGSkHoJAjQvxoAgzgZkRKIZvTW15Ou1WRPuZvhe4FNCTFJI2kiMRgc
5OUl+C2ZoPHR70/+SJ9sA9MrZ3IxXqaENzWzXiJDKQ4jABjQ7RMtIUHTxbc96oZ7
+834XHPOjWJ0viTs1WWhQSPX3q5NJqY5PryedYUSRsk23nNUiLiAb7LvhPbEaCuw
g3IklnPP3arygjw4PnthLWE8PmGcbUQTEm1VN2UwU89Gd4/0ElGWfxX+qrK2cBRK
L2SIj4UMIpwBYBLU8sebUMgrQVRfoZRDpsDrCL1nXzWVL3DKO57ndPM0yOt93Hls
CGBEqJ3AX++ERlrLKqr5rPrqnC9UTvMBLI10w4/oBUyiHDp6EcsYTQSZcgB3Zlpt
xOWs/KFy1RqepdEVuZXKEdEjLZYVJlkcHVp/kCfJYodmlt9neYXI9BVflNStfMXW
dGVxcp7INkgF5cAs0eUNptslg00HxW2pw2F/jd1lkMya5gVtklfO6qwiS7klTzfp
++kcn4KUg0sWNRV8fKYIubmRX7tNsUPYK1GUHD241KND52guwgBl7FArr/8LyoN2
rOSvLVhXfypmlHMPbKBCwLdlSmQEpdHi5fzZWS+OIzwZlnCxeflJ1FYfnusn0lh+
XeuT9TzDVaWnSORElBsi9sUdp+W3ylI5kNOXfwqyBq5Ed2tPZY2ITtb/yXFz464C
nt9TEzTX76Wbcp5PGcibILYbMNQ+VCFTzRg4Ex9fUKHkuRpYz4z3Qahiqsc+XaCC
gPtYeyN7sE6OQSoPw9bxKb961sTIy8piEDgWUcSmDEL3Lo3BRIPj/OhWLMGw9L8U
tbLQ0lK3l+HrrUGJ81NGHuARIAq8OiDuQmCmrqCqvHy4wwDdAlVCiRZubgUROThb
uk8Ro3Gsx6b3anFrcIgVwV2wp7j4ChS99nSLC9aPjNwDB+25TCD/8rXu5aPrftti
e1PGjYs2bMjlo1RxGNvNcWSmg2jsrt65FJvd3xiEQq1qGmFzrUv0qNxsbYWgHDkq
M6xyv85X7bmN1ZJ0oS9QOYFnfMLnzeLJl8LsiwvBxWVSlVRY8GrJo0e78iL78r5K
+mgej2+ID9F5kiN6d8xCK0AZDCEwUmx9oac7Nmf3QV6NdwLXCBpLQSUmM32FBGt6
wvi0XzmfjZmtkj5MQH+jojD1Vk/+XJMZyqyTtjC3PTQeGbPV5b5IGaxo/MTaZezu
7nH+6otOwU50uVaEzDcHjOmA0asbtFeYeSQyURrCFSSG1QQdweeKkHHI214vk+WO
iWPhhCdI/zpZhsvO9Fak18SAIaeLzoSdmeEF6J5j+i/hm5A6yeM3DTUzdFHxy/8k
720l1PGt2DCAoyCI2NIYLTvVkyhPOjfWKYP1PWfbIWFnyLgPlBOuxBo+EPAiKd8r
AW7lp8fC8SAIGcsT3TOPsnbQzagNXxmsBVG6wKk1gYOfvbVk88aBb+VVQP7+4RNZ
5sxMYndLVYb78gysrO3ZAmjI8HKzT4tJ+mkzZzDXrSqvEfNBegbTtTz95v3cTJGU
ssAyefreIQNc0eAsp3/EbDN9+JudVMnhVAi505yOr0nXmLpD72DVaKg9LdBcP0R7
e4CwmZ6ktke9WAgaledF4bzwF93PIdDr5pqZitlYGN1tuI4laM8InE8EJyHWbASp
h4o0AXUWN+e9ex+vW1puaSpO5IPtW+CSZbcCsZJeHJyaUxwZ3uMgVwg3tzEqKu8D
0JI+lAJXBsNuHXoPpSxEOKy6OkMgAnc2UCHZ+M/vVB1567b11fErdvMPl/Rrr4AJ
yIqxnw49Nitm7IzlSE5SkbrN3a6hNh7wS0lLXrtKIc+XyRCm93BVO5BT+QAWb1uS
1uBFUIAtYEvPJsbhe4t1g0DSgKd49vfNf3i3mZQn/AjqWxtTD71vrYzIRup2Ljsj
3SijMwr4tBnnjFCu34SgB45kRtTo1gWqou08s+KtFeORv1WCNq8tHUKxzJneHIFN
SgHWRPjcqp6KukJCPzcX72C9Qfo56XWOveUXOn6fnvGzMR6Ljnkb00A0yCsKj9R7
2ZrYpMGDoYPU2gp5jpKpvRsdsDqUY1CvWCf+sbWfVBDmpQLkGVwAJLYll0ms5An2
FBYbP4LKU2vTezz/xPY3Ceq95rFZZs54ig1++xn3fY2PJpMiQZscDU5u4hAmekZf
4dgkxopXiMff5/ZNZA0kWfwOPRX761KReWCu/kqy35RxEUdxjT36tkpeLfIU5+Iq
Mtkw9m/IGpNnn4yXBKJ7Scvy03XO9nxQ22tuXEkcaMX+7TChq1R6T0Hg7XxWJDGe
3LUPW/xx78ErdGLcKCOWV8lsGZkbhg9teMPKA81p2KziSZRqiain1oEIMdT3kjhG
6LR2yQuMwWPVqggpxQd9otJDg2O8eFXDCKLSTXeY5wh3NR1ix2i+4isKqOf4/ad8
ErSM+G2KpXeiBxT3cvH9yB2vfcHaO6jsUWoJRU7bPgVStHMjpV6CYeTN6nedvTXF
Ca9QKTWvSqxEvfyE/eohb5iZE4kOzatizAoYuMLDwWrzbFIqbsvNhjLKJ+VHw4m/
AHX5k8oMoiCi4uBsVgH6HJw6x3mfu6BpitBQL9UVOA3PkQ9KgW22zPB0iUJNHkpo
qtFIcozm5fy4q7tLSyfR1MQr53Pwyp/V15tqoszqeVJN+ncAZnr2rdQMR0FH7YGe
mwUrNItTDhN0hR4M0A0smidPO7p7zdKiTGLM+gBf2qNteQmiYrFW/4DtXgJo2F6h
098LoXwcEpD8H/5LR3svaVoqbQ9U1i4w+Yg785krhTdb75FQgaX0E+mDLOJ956ke
Y2f9AIamquG0zLCNkiKxOI/00wc5R3j3AGg0HrjXQNrtek2zUYwuRP24jCojgCnE
I/Kih8nu6nOGdo672GlJvMxocRycJ/2WXwVH6uvri4DeHjMQgXSpP2k+64FtK6+3
Fw4Dp3YVw7QGwk3nxe/kL7wyDEUQj6EiX97xzNs0YQRbRsTSjAJMDvUKGzgvdrWF
0FTdz982E5rtN3rgnmlImHgntOYQ/SZcXT0nJ9I67GF0ZKae2IDBQCdFcxsWccMA
pgx0tA/CHEsqAeu9hpsfBwHwlx0EDMb5n0OasfdN4lKuNdPtf+HeVyRox+9t9QJ+
o5Hq3xMGdy4HP0VYOpkSZkk+DMqqwLFcJrLXdPZEfyoGS17EcwQNrbG0nNcsbvxA
RYzrWWptUtyeUCeG7SK10PT0EUhSRDpX46agOnRsdp0BOHf9hR5CSHrM1wgRmDyy
ONsyMcibX58jcdLvl9KcNpVMVijBe1lVKgyzLeZtx/xFSCT2n/5xxG8kW4yoJQcQ
vV+F6rMkBsxT6QSTKWafYtRoDv20ZcOV1c32vcZfbYfl1wWGzX+myyIv0V/xtHEW
gwhUZC0VTG8NX6IKAle5UZPc0lWuZuxMuBGlxFU2Vf0EH/+r8CfqqPPIC8KNQrGr
bv+4OJlquFohC4X/IAvupnFnEq393o+Z/xVyoHwWv9GeQhRqSXup++h8tzXPC205
mvrM/7QRSRN2StY+ZUMRU0OaFYaXI/r1BMDiEKlkE22NNxgS9mngYpzKb4FmT+ql
bHtbggv1IllwIfyMOzubiHd4uUygf60AQoskaWoQCVk3/nR13B93rInShTa7OTsH
g4p5TWSczzTbWCetRS4FfjJN6D09yeRFU8oMG9CpaX4=
`protect END_PROTECTED
