`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8y2MXZcrzvmcJkeeYAMLwGnaGb0Xu0l76NxKOHhGzN831MTOYWmZVn2Falxq1zxM
Ba7Mo4xuFAu1kMoyOTUIgglfYPXUShatrUAfxhsgdsMbaNHioxl6XnYhvtSW11sv
ARePHnoc5RYZgD0MMP1Nz/mlDM9O0h6v/wzWDUTF7g8eQbugzS4KTtHXOWD+k6zq
wTC08JdFT8aK562fXTs1L8BHikLNx70lGRWU4OXcm4wUIKSYFEkaPxjZI3Jiqw/p
DQQcPBO1cojj5MOLCrMONPrO1ikOk1whbIATcKtsdKH5zhUX72leWK6rz8/Bqhe2
th+dBamXdR6kDAnDCQnCGwVh4lT435CPsGkDcd3uIkKYqu+vvX1pkdeIrG73NL4a
QF9k+vACroCuXeX0h3QIU9FWJnb6ZHXGhkwJiG1Wf6OiUHhYrYMBH8PzDEQr4JFC
XPhcLxhylUjtId9wHCH01ucBhgXpLAMZrI5Hf9UFXxWpf0G/VEjLPkcHK1pYaTTS
hXxirQN4Qg4kdacNeXFMhEOrp5oxaUrcnbbU+9XBQ6IFtB0SoP5aKFomT2c5AUIo
ocCkj8aOlSwr4ruLXK1EoSMSkibaUTjuuAvuywIXDxkUtt+NOn6/h/RfKpAAcmjm
DUzIKp5RIn7oVS/5iw8RXGJS3LzManjPetPifRuKkgILFUqfIJ66PXA/BhaWUsHc
C+dTQz7+SCG+2aqZYn7bGg6LuPnOOJ1cDDhIJsyJFdIj7pJUd2IU2EkUPNTccb8r
zqm8GRiWFHD3WAvCEU9fDQNss9FLhaUg5bdeq3rTtMEAwjaM/VcmChmjosn/3mys
pPPdm34fCnjsG0LSUnXHqki88wq/epcTE05fCNpCugiuS81uTytjSafCBanfXv+o
0qA4/nvz2yLnyWQdDrGQSlbFRCMpbGIUQraaybkfUAbPEw7ZGiFd1GCq4ikDX3Iv
atDmaq5iaX1fxVhPDW0kM+62wy/3yRY54oyVM19cDRSzZ7HwFQoXse8YA3Wr4PhF
lF9kgcosH9HmZmcXdT4U9GKFUVplJKQOnktCBgNn2NBIUXMRhLPgyxOGmyeik9DK
ZE4ln0u/RtC9vQ46ZsRGBs6ogRIGB/DBDumy2DpwgJlQ0HdfHczM7SjnEvmyk0bZ
JDs1CoBR/RmNZyk31o9rLyJKPoL7vucslRyGJL66fwYAJg7enY5cwagpr5i6xA1B
953NJqAUdTYitb5/ckEIBiG86ctKq/7+2F61xQsaQBQlX8awITsVg1MyL/n9xWg1
XUQvs957AVM4xU/V8pcxxzCxNk5VWP3wI3lwsYgAQlSqZPW8Sj4wY4GVxXtV6gIL
r9KZZFCJUX0WnJpFxS9lDuY+2sRGhxW3WbXwCMB4o/X/9ypX7QT/nHXtWQWNx4Al
mM8lzpBNkt5Ol6FJ6u8byFOilmpPfFAxYbvCnOwt6v8AsQKZbQx1Bxj2y7qv6fIA
ki9aXgqEQj6cGXTsl3YqJZg4s2eoFEVAhLMdqN1qv4hgDiWTjR/U11dNNiD4w56A
gcjm0K1n5aGlCgPKCKAA80Fos4DPlUjSdYqBvwVBdAEe4EwlaRSYuB9anah2Scw7
ntynXgQ+iOQOoEzlhGC3LQrCr/jWQo2VwxJtbD04m7RGsqftytXCjFIbDZNJj0fe
aoxdGlu1ZdfHLAJIBkbxdQ==
`protect END_PROTECTED
