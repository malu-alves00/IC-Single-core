`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+BLlRejKR5LoYlgm1FrDwvesIqofJzVIb6okxOX6YiKpsdzYaxoUpgBnNGrlt6KL
FDMuiti0jveldPg6skZfeY1lJo9nCKhTV+H7qhIw6huLm2Fl4ymGQwbfY0TjhHH9
W1uq3gWQMf7mOlqR3cz/wxLqbzfEuPnwY8zEO0m78FNB8xtjDA0Q1rcU4yXXm68S
f2rFImcMrqpKl95bO0XWe+KrBGAoS8yLAV0Kih+UvayuxFfO8ptNRMRIig4zT3Im
4j/4+K/CNmMnTSATUVGBCI3zD/LXzYT8NgW5z1RzRFf81G38M6GIuMZKvtE6Q1km
wrd9i1ZDPrhUUqGMIOsTO7/zU5ZH8KZ/vE1pkbhPApKBsL1Ys+2+j4PD9jhZ5bPh
99zA68GZGml661RlCe4C8tKSx5uMnXScWMjYW3Fj4O+pyj54PWRdsFlvV1oW7vbn
dFuDqufbW6imgIA2pf8iEWq+eYsJ56r+B+SQFz2d6asiluTHZxcL9Ycmqg4E58Ho
P7q51KpckDVdKRZWl158zyuIDbsNgGxY31XmgBPrJH9uu+ZvRVLKnhq4hhqfv4UA
QvKNC7aCAArdWrDIizOAxR4jqVrtMyhvZidKxSBZP2tdmNnC0ehoKvwJb3fLeIvr
DJ5RX3cSBxwNep6kVkvoQ1+o3u0FLK4CiH3ibD2r1mzFlevw5ewEtyfkJEulu+r0
flAaDqNG3jHFUVXetVIbhPH9Dn2YYnRs/6GCSLYJgQclOEgRzZ8Dl30GmQNNHtqf
YvBHhE/T4TX2fYAB5YzLajkJRs3RxJbeqCd2FSTSLBI9PI/W9pqTKVceuuwk+lGh
vYL13Ijn80bo3hMxH3yI7rXy7oDNv2//AvLWzXXqiK/0PU/57lO/ooGBkwNj3Gd2
y+DFphK+EbnjGU71IECG3ExFmkgXnT2GAZRSUGHKdQrrpolxy3vnzuGVy0zW3ply
IwujZulWlPZJa2wBHrzN6C98Skpynhgb5hkoCTuHIHIeb43yuy5ixdxGM8Jlya2M
Na9a95LXOIJxtOpGO8mWu8k3joJYAYtQ0kmxeHDW5zQMk9QVe00nELBFJ1k4tElQ
N7EWFZ7Q5b/Vmclqcqh+OHMBhxb1Yicbq50guEQ4E6L0v0vWUFbeJWo05ICiTq6P
3GJY4hPVvtzCnL9LpwJpAbJPB6EEoynNwFhW/oRUXJkde8ugCORGlrOnMbb8oSp2
CCooQ0Ws3DpZe45ZV+QgtaL2F1sTVsHVoN6nCfFCNoI0Fpox0//Lm4vLk6txWxBU
hGqgL2XEAlguR8vB9DxDcCpSktOwcsmK/JLEs2vUIqcIByWq+GifYzCcKhcfAIEP
jeAF3P0mXMWCYOLmd0+ts23gp3m+utfGC2KwjjsjTzVCbkwVIF5xaIMAsp2Eujwq
BcJB0cvE8oZjBIhGgUlP2oRuwzX+BY6V1WPoPFQTW1UdlQ8HlY3RW6MdJQ9Cp5bF
rnK4BY1XWykYuYoB3hWRrIhHJqJOxuz/8+EG+byY82L/RO8ZVnNKmXkyCb7mzgL1
l43p3B4pYQWlIhOcF6zXXdjwZKidc8US6dJyK5gzAi+mnFQEuu3KYAN7KpSR6cLc
HyhIG7oPGmkCKPrMajSSnZ10ar0V1R+yYcTiVyiV+200pS6eLimS/7AsUgUY+LuR
QTi2r8f9N1XJhsfT8qRuuWixRODo5ol+0HKqFx72yCV5/z4Lw5VvTYApZHQqW5AL
wTvwepd9NLSSUyF59BJ7mdxDUW4+ikADEyHS82sZUO5xQ4fPIOVs1VVZXE+wJTDL
TePewC4iH/DVdxdaT1ZGGsbPxpYsjHeLWRR0xZZnl4OpSzM7G8KLSMH1smHQCd3W
B6KiopbPUpB14QWd3CZCPKXVykcay3EAyhC7iTx5J7Fxk2VOI7c9Fn4NPtSLenS5
Y9uEZFLG+EGt6FmTx0b2qZITYXjCVkYXXgfq/Fxq19yGtad9dvHWU9gd22Rwc20u
Y1xlxZU/E29wnhhIE8uq1cB3SbFwyI9RA0a5Is6v2+RPeUcB4hd+tJAwQdz5HgGN
VepKOefMVaqvxZPdUJCom6+bJgL81HxIgt2n5WCJ85qs1VxjE8bhQ78GZpV+5Ofi
910rgUq5mtDkv8McpbPZy2V8NpyWZneQsXChPRyKPHuSfHYa+j7jP6RK0I0EWj+T
8sX5kdG2j8D6P2IJQ6wp7MMvGA5ZgiC57G9SKI3qy0ugYSmHGJTbArAYq62Gm3MP
FD49/Rru1Hjy+hcS2QB7WVy5in2X2DSV7YADl2bD9fG6/vHWMrIDp2xU+u/0/WaW
ihV7UA80Xj9Hr/zSPrLeObQaZaURuto1HVamk/iF2dEDzFEZ7ykX46P+ii9hiiKs
hq3SiVyAc/CQ74IeIlW+MsB9fT3oFb61fxugMx7yIXFzzTpVkEEpbdXGKoOUrhB5
GALJJiE5zikw78IMoWqGR8dA1pmGhiHoRHPDNtr/l0/NQsAi3m1pMMRkRu30+qaa
kJOtIX4V7G8389QzTJSasDXiJhzIgpIdfrsrFfAl+XrmxNe/eFRaUpZ1OynlaF/6
NmBQ0IlLqOUXq9n+1JryPnFifBmki4diBI09TxrVaLQ/2zkyGYrAgp8qgkqrap+m
N8RBb6SUo4QvtT5YumukvAzmJI8TM3LBwqMzK7dXrYYy0J/gxuKmA3/aKffdqgLt
8fSeSUagn2a59Y1fb7clzZIPiGSLn5lIttjtTcoFA+4IvUeFgXQn1p+L6zjtVOum
GHQaQQ7PzRT7k5qCLBUczdKfbrGn71KFxffYG1nT5RZN1Hke8HgmanMXlVHQ/Ame
9uflCESFwsX2LjbBizFl23apE3H27igzJ8dAyavubo8MBmx220jtKAWx9NElNEZG
GihEVu/LE7foYBLLhWg50hvg9xR/xHayJBwsX51xALK9TxZpkgtSy+sJgyj5x8Gu
J8WGXtXcJ3Fc9Xb6GUrto8puu4d9FjNMX7/Y70bBxqVJDRHGq64FH9tijEFlX+WS
0RS+WR1//aCneXWaktNMWNtFFSGZXX3vkEItzT0KhyEzy75Mgb6nxk6vuoIBesrj
tS2wQUiDolntEKs8W3AMjUm20l4n0umacjdp8/CMMFu2lrxgGQnUqVSMOotzH31v
p5N+adNnH8wcQWbDIR3n3BF/mwRbLFzNiGh5SAEQ9SoWbkWYKHLVzgUOP9S7DDuM
S71LyARXEA8OPfFVVGJwrL7V7/w0jaUIBvfonRscdHRGVvfZqDV/QLI3lZSKC33S
B4ooc8McNMSsv+zvAB53ZURgaRcdgcPFEi9TFWnyJSauiZE3kp5uufOrCMHtksao
6WBwja55AVenZhK1RQezd2tV4pqGK8DWqhO/HVzzcUZOOedjYDfXKpiSvZsC+b5+
LZZq/54xdoN8x5IGLNYQkv0W40cS0twfX8c3aSf616jpbQiPWe/U7V66aazwB9rb
Eo8TPe1gnvjy8B3l+WsyheA2hCgznrrFfpehX2nwYur/h5V1YR/ZkPWEndZFMc0H
DkG5BsH3OxwJWH9vFTyV9pNWCLkCAlb9vHeYEauIi+EBGcgsuvI+3QXuACx2XNNQ
IGr2ZPA0Ng+MrJDF6dB6OVq0LIGaukMs7bOqtXU3vpPTgbCukHoRNB3L4R4yZsnU
WPkwNjGccYgP2pkM8kpcYKo2HHbmxxE2ApsCmh7XJvin0QThXsg3i6N6nUSnXb0W
lE2ou3oCbBNV2dEEBi8OZGRtXZ6NsqBFWtaUTLwFgYMJjUseTQfCpSE8TtyQMsbJ
pWtPGIhOuSelIw1PCvFnlzcba143wrjqyPNbwNdJULVFEjSsvfdpJAdAL+IvHACJ
KdU/WkyvFxs/ULkVuAPO3SOlxwp49sjSgxhC/8sBL5HBpHNlv4Ep8bYgFgtap0kd
tD03x6p3XykIIH6PVGC7O7dZZUjeGCOWpOA/0bHvw2OmgP82fyDwYJs7wDajzmMD
dJOKQxBdvMM6lGHY0RmNBDBI2Hncq6BWY7pqV0mXQLqWkEW/1oCwtKCNbulYUgav
ymAlu6fASDGYYVeBWObzxPs8uvEyNs/M3IDP34zxsPVriA3IQL2l97Vv8QbiA4lu
NRQNAQQ1xUx8N5rmRbF4o4HHQeq0yGjnGRTqU8urk3vKKSLGqkTXVbySnYbT+6Hb
`protect END_PROTECTED
