`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mAqpWE2Lmn+aQVSohevQNP3vQk+FOjL6V1gveNBVkkD8FoggBLIkwNJvvzwBS3LB
iQRnsT2KKHjYpbHpfKsaC7TFqmY7g1MgUZGsncfKKjjTBsFZ/syXRDPsavoD6h9K
9sliuR8iGF+p/245buT4UtYNs4DkT7YTCkOGD5MaF1IN6Dr0UMqiMepOoakrBd56
LMEoZ4w/ciNyupeq/UqFdIKcPbDF3eBt0uDZeEcOk8C2S1y25BmCgZR+1izMFCQT
0NGeQYP159Jnjq6M12o5o048gzc5FAhZ15NQ3BKtOdZNESAZS+0eApwmRyQKhihu
3t5AXw6OwbkW8+hggyj63c/CevuF/5pvtrOirUmXMzV0DUEHt9bz1ASgZyX9F8FS
woq/Ic0mHT8yTY5nw/clcBDybGv/qt4qBuY/UcYR5yDeMVSv71GwBHSyxpfaozoZ
gJFa7sewTZsGm/O53O5U5QF2D+Ra4AimwALRfGCsx/S59BvOxUbXvjPpuRByDl5K
+tnmgroO+HRR18fnc1S5qDFmMS8g2r/U7RO8wI/F3wHQZE5frcvej2c1NoGD5dZf
ZmteMmsMp98xk9gIvRVGcPAZ7UXujpp2sxy7tfTWEjbrY87rXlhpl9m9/W3vqvRi
XmHFQ4vlcmfjKlO24ao5KrCZycudVyGicfyowxa2K+3VMnkahw0u6VJPi7TjZoaW
EMTCSq/ZQqk85xUxMSrU4HoHKiGw8FRC0rmXpE0RY7Q9o2Dw7NrtCGiHiUbY9a4u
n4XmTLlEn3s9pSLMUlUwaSLkucJcq75h07gXcDjiXRyFbeTpqXRHmwoWL/WxRbdw
pcKZarrGJVTdyTWBT4DarRQVpYhpJb3r1sCIUfJWg0oP/h3CsQIypxvkBbbfN6ix
yX5Svvq74fboPBEz6+9M8acZ0Sg36G8Ks8enDxLyuKQep75qQsoWZX1e7bMNo9Iy
AKRKkmk2nsEUgx8Bnh8iJHWeYtwsYqGbiXmt0CvnqMg=
`protect END_PROTECTED
