`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IZT0eqyVmAy/uUqW8T1qWvDulb0gILbXPVorgeOFEy3uf9kaOnTqZXSVGja6gwh2
uN2pYfBeC8tY9NIj2IJy24X35B5jdQohK92BEJPV0j23TpnO1EfMxcuWEPsbvSCa
RnJrnoAqwYahPW8wzt8mUR8cjcGfFSeKF0Qrfw0EvzocdquChTTYxxouxKGlJPrj
qVldhIj/WVzm/nyVgmlF33vMUOr9apsjjYzyXZ6CXTByH4aAdVAOsZiDqEKgu+lj
sgQthsc4cKpstPc4Rp4iRTykK9yDZGl6stET6CdyhYMH+S79Y/a7gYIv4LFgEvFF
u7Kp345i8jk+G1bB+NXRm/mMiK5zTF1UKY/yXZOdkcvdd2c64a+jcPTE/grLo7TN
LPYsKS+P8MR39nVW5panb5k2IXVIzp6Mcv7erhZHJFIFdhd1ZPV77EGdFvMInnAE
7DihQlU5b4kEkYmKeVNB9dh5dxBkLK6VG4nO0Ye/FybIzRtenDyVRf5Q1iBdwH7g
tXv/SMD2L9DzQOJcV7FB/qwQphNbXxHEJ9P5Mc+NO0I3M4Z3Pw873bZhJbbqb2iI
QQfZtU32QfoNXvgRSrVcdFiG38d/5dGSxKo5Ojc/VGEllNJXV1/EjHCTytihOF++
DbIgyWXJ1xF5iqqqBIlHOrBEE891N7RhXEV3WqNF9EL4z9kv+9nPm4DSZ+Ak+Xvq
uPaZ4zNNUaBWWHp3FbS8nZNOb0zkfneOlJMyXCrKf7Am09Wk77vu8bLoS++OEJ59
jQis7HjgdpGkxlQUL00kdQ==
`protect END_PROTECTED
