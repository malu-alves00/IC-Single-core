`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UAmIiOCKCEtSZiZn15gGqNA/HRPZQABOg1++hyL5Hq7Nq2d1JKkiSwo1sgWh/ZSt
nda+pxAxZk99hP0En8dl+wXasBtWX4HBvsd0fo7dW1XRqWzyUyXkLmN2I3XQTTvF
MP73RO0gljvxEth4ramCp+6mT4U7XoCq4/DbLqcOug4DInwnnmjYaWO/TitdiafY
+IKUncw7afo+VXm2uhjY3TIn/UHrK0xUTXeyy9XxO1Nni/OtupHZwRux9pWwwFHJ
4M9sg5G1yegq/23Q6GdOB8lIxBg2OG+z+sEdQGlMWnaRyOZNoXEFtb2RgTUlhKYD
QnBareEkZn33f147ClGzegyATudMr7E0ctUWMjDTFK/G0Dm6MydyZwGRIdc3UUoC
QsckhlRc47EZqPl5kIDAiH25qHY7IB+YxcMSbgfcmQW5aSRtOexuH56e8wJi2K8z
NaRlQLEpvq8WpAx6pjG3+qQQwdPyilT1tRnTuvrBnZ4VXdN5RddbxPhU/a8DyEAk
jZDkSEBN9PosccPmSnCBGbj63p1kpks5znsm3bbT8MMaFHUn5+h9fnI09HYPERHd
N2c0NCPi30TqetaoQNJrohVf8uvV18TN+t+PIwRBSe3XjxhYZ9hT6kjVBcvQ+EOn
YJMNTKs4Tqxh8+g9gTLi5AQ/Nn+C9l4gcSYKe50V7L2ukOrASlQq29G2U6hZ2l/Q
F2gjwe0d3tZqSJ1HWaV3mK5S26LfHrLf85N/dv0U2h4e/2jl/X24gOv6ulMGrvcp
bXQLjroPbfOmBK/3KdIYA3WrsaxAXVyjiZMphrNhT0VAM0IFChAUdiRvAFz6S9x7
L8lQPklMWvXQTh3aw57Hck9YP3U2jZ5c3NrcqR1dsKnH4+iGu+V+vgBpI91SSjHG
+hKa6UyXfkCIG65MggS7OIWmdG6M06cfCiVHqkmM/JzEIxdHp1PZg9GpCTHvUnyx
TCssG16fynKz9VgmhIEbdKilXUYmSTvQlJx4bGnssp+KYOGM32hv7OtzlUBeEFRW
/sITGO0szWINLRxd5NtjLa9B6pF3CPr4AmYlfSbtukg8wSx/mg5bt/B3WY5tlfN7
5mLd70vLlMyXgvGmncmTmmrHyA7QqYIqyYOBP4Ac9r6wbNdK4No18d207C7lrPqN
42NuOjyXMFCOE4D0hdTSukFE6T+uAMX89AHAo82nMSfYs5eliuHR1WtXuX40rUqe
9WbPMi0b+rt8V+DF8fZqWKR9RJLAy7z6p6ErMDqcpeYMvAeTwpMSWSQqwsWnZzz9
nD4GGVSR8Op8GfV1c6Tw9GfAwtXnyeczBZQKhfy4LnFCHT4H+tCTqkoRQDJeKAuX
d2oRf94MejUR6YjwFuvywY/B3j/nBDyKtNn+ljeWvFx19QN6Y+n2zJGZHuwGxkOm
FVr2N9TnhseM8YgcjZwm7JqpI3itchkfEm/yzNC9jQBfncw3qzd7IVxh8XlUV6T0
czrsKa3UqxNERCiBZtbyTr9+xz5eKzAJHzkfXKsyXBFEy4W/3nBPTBrwGRMaLe0B
W5m9TwzrqpEzp6AFr3d7hS2pPDlNrRnFrWufgR0ssMboUYkQqjMofd6FG9O9I/eI
Yc44w1qnBeXy8HGz3kb37+uP657Ta0doU6C3LdskE96/2Ps5ehgV/v3SMffDsgvS
1895830KkeBI1UFkbCWf1pG9tYd5RL/rFDZfLM7zS61MgFBYKaYZmC/jdxWFQRUr
tvXGGPttkczoEtGV5uMtip4cRWgqtImI2bmTysM9fHfGFeIYqUGOWCUVPCxmx7Mc
j2b7oerq01qCZFvHhz0W9T70p13pfx6nCt6YNNJqf6kS45amtS9cpOrxr4yQ8TAB
H9Mj6DpBka05DHn6vdrK40t/nNq6EbvsxOV4APdHzCL/MHBOgELkVUga/JFrbefr
WtPqXSStyFvmsQe7MYEPYJpLSTpDwvRj+KnRD75Bkp9G6e/MtLfk44xq0WLct5X+
Fgq4C+tkuBN8BiZheqhvFBumVkiAiTRKEC/yvRLJSxPQOHv/73H8svvv+UiEne2c
9vAEBFmt8oSoDe5ks1utvklilX7l+eEoR06zMHEegTYamV81O0mSRNF5iTY+738O
NEWeF/py5hO6sViRu/X1jJ531EBXOq/sKEASemM7XulHyxPSkwTUWH/EY+zWfkp9
Kz4ZGiCY2hPvLPeUwrmY32Gaa9niMq/M2RrWX+B/HS8dZ4eD0VWns2E8wO4grUql
avBnaWcanGhckTQ36XHD17vJGA2IywDF4Rni5feGQVFgSBaasgZXnvCt8FnVPwId
62D2vXu3WWE/j2SQxlQX7c8jtAPf4bC5I2173LdWUkdnS+7FvRlhVNmLivD1hzvB
Q1ztBoaBD1yZKaHedixe3sRA5VI1FxpHvZtoewqApLv3NROh7E/dZqVviXWcEJIr
PVrwGEjKediuhnBoCLTqG1Xriu+z8/S+cbcF4FL6CTMv0cDFzAkeXTp14WaHt9S1
KUvdU3Vlq8jFnH/OUqRZRVK7j00+6AWO8dbgk+4zcNueMKY1iVHfeU1R1Cn1B1Wy
IZ/ao4D5dklO0lxx/YUZpN52zldCRvIsRMh09Wqsu5fqQrUZqddhOYRjhSeh0P4H
zgJRvgPF96NPhB9hp1fCEBhkIGQF4O4ydmnRFTAXZAvmjKaC8kuDkDmLp4lidNdC
u1w27iWk71MwknJM4B8XFAtT9FJ8Llq4y2e21DXxs4zbWUmCR7Poeer/msLF6D6T
6kYUWTmtWfrgngBgsOLPQ03mrVfqSwDlXyJiRB6Rv7Esmej/GZNDMJNBznPnIENN
DzPcp82WMNFFDKCj+TFDhKOWQgXS7QzyedbcCD+bWtQZWxdzLWc006mPn6A22m87
MxxiX0VvAqg3JRmRsnnBKBi0vVqJvEC3cu7J5y8StNX90srpOjj7QBeUikk8t8bG
WLuh/f5wAX8CNNm5hHDeD8D8ed3UUkPqYdqLxr+10qCBi6fH96wGiDTkLq6biSge
vpVcjmHhs/tXOWsZk/P7kEVMK1RPIxlvT8/0f9U1/Yk5AuZdwrtFHSQXMiivN5/9
PMRFSn3VyxBajoHt7XyU1jNk+2Kb8ns9zSI5CgmpRTW4+Iu7llIj//bfCqpVFfhW
qoygluUxl2G0WoLgBuEvGnJx2SGyXQoMQ6l/cKMC8lhXzC5gYqhJQk8jdDeuLHGP
Y8Kvbz7O5ji4BAGs1twAqInGmLm9TlB38Xac/t79vsW7PkmuH+dUIXgshAn0nbGe
cUdjEmHsR+eUm0cyXC38vWv/2pVXRlo8jXnkIi8qhhOs+LAVpqw97o0UV9BqmQrL
ieV8tIKQlRgpXO+7R01IkmUojONNGWs9EebNPBB8mz13p3AZOrA21nDU87igDWPH
q7MzX5/geCaxtohGogoF5FgROadxO6qqNiUp5I1RixJbQJp2uqawhSV71r1V/H6D
ECtq0Z6pmkTLYJkaRoxtr11W/B6PqCu5kpX2sUv8yrw=
`protect END_PROTECTED
