`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0unONXmneb3+BSvJi8hnMuY7CTkGaP3BQMQ/c2gKa1Q6mkWdspVITslbNYVDS8NT
dEVw6wVqehyBWF390iChyFhXUdhCTh2ULRhwG05uPP9E/lt4rCvoEt6EzeeLf3QP
myaTz7GgEyTDCEPsPAoUY7VgdgTnoEBU6rzXmFwUI3cZ7bqEDqAlXUheI5RrSpVH
VXG8veb35Xqh4DXgdw8iFk6m8qkxXt1ysW1qU5fNhmevARsn2XrJqVqxMChLr4dE
X0OG91AL14NEMPV69uWAeQ2FIp31mND1dT815XS80LjhPxRQFQ8rpR87egWbuA9T
loQXRs0KOkWBpqYgHgvBAUxO5Vw2PbWj3SSH+gHRDvXqN92DnpNIkS+7FXMDhKK9
NX5HEi2UmwHJ7ODrdgE0L0QLlJqry2QjeazpnN7zi+mLKwE4RRggd5cP/fiG0wri
rN+OiU1MYyPVaizXwes+3BKa+M+ALTC0hNkAQsiikSwjJ4OLvUBVSDzS5rnxTZ0i
NppoMQ0yv3+DYBRRAwTdXzSmc/gOOUQMKm/lZ8FlhGvONTQuV1kLXw8MryJh/Gyb
GloNbXilzTLr/PkbLa2bl8SP7zyOrF6hb1r+EiRxEebexuvViFa4IbdwCW2FNX2s
vYoUnvB8tRpSno7On6vzE6/dGW2Ow3w5oou3mxu4ZB0e+ntfWIrr6fdtnSNtdygg
DqWId7gJiAPTjWs+LGq4A4OoqCH5649h9gTUZwyAi0I1xhVyuzvMV2brwejJAzPy
oblnqZ/3s0McHQVrtAz2N1vmnWdyJi5RMOVaAx1mNiCBneo1/k4rKANbGZLqTLm8
DlNmZkRVX5uRYiSA/OuwurHQVC78k9HcfD+eYFlxt35z1Am+iXofp3fayb0ZlHR2
Ge1suCn7tZJPdFWCOkE7CioxojCrEMUsjtEEi1/DmGCCynQIxHOf6adstuJtqoPX
wuAS/VAToau8n8xXj1gXQXDIDzvZ2et8swGb0yC6nhnzc525CqxtEJCrL4Be7Wk8
TTe9Sq01IJi7/p2wI9vc8l/8eKlZH6XD7EEUqCbSn5O3tFhn58K8pcANWEeQ+qyH
w1OtrJZpOIM9tS2jDqVRm4NfKPDqGlT5ezaJiNB5w/KkYGhEzW5heJXthmoaj297
2ardOVXrr7e6AI/tPHam+4bd6gLilazEdi4VBtbzZY+nabHpcB/t7V74p8fD8Yfn
/3ePHwgppW715IXuAXaaoZcsl1fyEAAVq5wlP3x+OHFB47FAmOktAZE/mBZ9GjX7
sJziX3l40APBGcdyTf4uCCdJ74HAN8uQ2b+CL8o92OY+ATBbvucBaLDZMWXHteAt
1Gkv6k9ADBA0J7vJEROgOYw0By923ilmVaE9o/fg4JS2hn1TduFFxqWZUqWg+BWI
mgRpy+E4X34TFbIC4E/gM/VIEQwn/YfOCnsPdNA0zJJRojlnjN8GNL3AchtdK3xx
ni8a1O/01bZQMHSLuP9bo/lFiadXOGDEYt2ZQBjlWLORZME98wjNP8HWlEkgFHHr
r0ptnDhAdKU03RqM1isZPGQ+qNy+nbIG+R+Xjfg2o58ATtc1orWwYV8hxKLxiV27
dBCBVmpiAGtokm5Rs7mGz11D+urSwArqYaSUGYeNK3uD25Yk7alnykonCKwagozL
dk7Mzm7eOkIISHEcGx6WB02c14SonXBOWzhcwERJyY1S0eViNbYpOOQzzQowQoRR
qQYGvPo9Hnur1WcYk4I9G0WX5O18tWpfxfVlM8b/tVpe6q/IjMSphIv5MeuG1hoO
1a/Ne5rOvME7znQLS4265DrtrSCHpqwMqPj5NcJg0jdsa2JMcG0f2xtLtKJnH98S
Hyb4ElYfkI1dFDsrms6tZK/GhryDKTJbil26YiKizn4vy9qRo85cZuexy+x4ZrO+
hsMHnxVKi3Rg9+Y7YpKLNQ03+v1xJSAFB7ZVDq7G0UB8sunH+AosSNSYFTdshaJP
rn5wH9zvmfOtP2eeksFVhkl5o7EVQWzNMNLG0UMkOyMa+6KCUELiaRD9oDmeL7J2
+cxfow2pS62KzETELPojrcC9YcqkDe9OCIXbGn6Uo9aMH6wDIjPll7hB+Ypqlx+G
+RXRMiVgGJ4hhgUjfkuzKNgEvOMKBKkZLD/6whNr8TmMYJktZ4FWOBU0kzoPM2YD
rVwQEOQEL5yvj6mDvDRb2GESlPgtmefOi4DZg/uUQeqXnfoOviaTPLyUMR926R3n
3Qc1Nyt5OdySp6vRTlnniY4RVD2bw0IRFmwem8BqJSC0Ft493d5wLDQ//wCbKDRj
N2XF3eEH9u93Lizjo2pceFSyYbpCgyRS0NB/GtUYxKfVOd0Y+je8Bx43ThKx6eLW
FO/ytwUgR6ILYDsxWMG3o8rs9EgSTs2X9PV/oAtLl/5G32ZyeHLR+A5Gk5zJHMgQ
zOd/pFfB0LipR1wec3Z3MExBV7coJzSmNWjDNuDjvC2VSKWoqoHxxOF9UEemCONL
5q/gbQo8v/1M6LlZB4hS3du2nLAJ0udIlo7glQP4woLqDiV6SmPmn8yK3spnquo+
AoIZ7VTxoUOy1JQbGRKrpRL9u6bhetlIiKtp2L7/M3qB+rSOjmO0xSb25fzm+1T9
4jb8xRV10wgEZFrJ1d4sS9Z5oiKMpMa2zKj/2BHEB/xqbsRFXpGZ8qGjQ2ffAzof
oXzHH+7TKOZnazhPxLyrwT4sL12nA8RsKusl5t2NV+dOzSAS6YkC3eg7nReYGq1T
ErozqCfPe5tP3WK+m6q7FOnuay5Ql+6JGokHPVmpLkSfpxD7adUIiVgfikGLbs5c
qXFfdq7GlwMjFrmpg46/iEDp05BjJ7z3yLq2yIuI74BS8zUa3qFjpE5L+bOumaWC
juNHP/QTeiWtX8ljsrfX8jR7AXWgGjawTKYy4Mz/7fneeWAA36RZRpnrdJ8rb6OV
AOF3KLpHOUGMWf5tWm4MVUhhlsmkU4V3xaLc7e+VMMOWrIPJNiaqF0kVAsyTOUE8
CtbuB80Bp+Rh7ujPRGdMdefdhzMvSJ+6gumdYYWLSvFPdzJwufj/KD4VdjNDp3qR
QX3MEXVNS3LVrObUafX59Iy58ibakwzxbPlijXHg7coTdZSX7921XEZhho3xbE0b
btaMH0nKUHLcRAwRB7dH+bsAUUSFD5Wnj3NacJvAuzb5/0iszmupRj+P/QEEsUqc
/ukA5aVbdMQOHvsar3M2GOUboepjar24YVZEGYHldAXiYQ6Xe2PHx0DOdTmQa7TK
HIv8fehoUJS5EI9v8QxtO8zQ8KGcX6NZ7LM6gixFD+WUWsk26j1hkHsWYAFe4xhv
gso8mwtDN1DcT+XRgSprjxeVAed7mSvcLSVcnbejLtPsloCY5COKVxAAmXGZmQ7M
54Wyc/+f99XyOXIRNUPXJhoLs1dqO/KJyeTGHb10tkWwhiNoJYxr2GX56gp+ghRa
0+AWI4sq8fhWhkEYw2dDKnSzu5pJa0GAyaVU8blblrmBKSrfHDV1W+kd+6CR+EXA
UtYzf57rdQ2Q1OigI/xezELUSc4R19yfkndxAD/QnEuZ+gv/NbE58EPgHg7TiyFD
yTJFsm0L+2DVkOxQ5Pc7RhhWOXbJlPHq5FmIc/Fk263qLmaf4L1IIlrGunbobc9k
xtBXYEaYpWYUoXv4tbZ8rFLOn7ZOg6eahQcxfUlZSZ+/c08Z4ZbzOY+zvnxfd0CF
cjeCRAf1Og5x6aiOSFOxdH4IBpo+ew07nt+EZhP8i3ifeGeqpaUOBayDoLe7hJdU
Fjhoa/v3evpU2zyM6oEpq9RZqAlyWMBK1m11+oUr6wZCAGiPxSmAAlxt36RJ/Ias
euVIYyMEi81UYxdhv0tJWojv9MFKlwohcqmtjVEkYMwasPnwapLnSx3hrI3SIc0k
dtmFgUHmaWxyRJY11kdFtdPVGUnTugUnehkylAXef/1fDE8pkMPbAF97D8oxbzTg
WSVXeNfoi8AhAANG4an3U5S8+QbTiIUWlG0DEkE2EuMvegLoeSslYG/oaqbIp/3e
1dhoBzUdUckVKIk7pKkzc/lyDUzjj6rO6DSLNp7vSk0Slmueo/81X4Fus6CZTO7S
PxZRdQhBReOlNjMnOTZsIgNxWaMRb2RY0aze+JKOMk11QhhxbwGLFndboh01KDF4
/uOQSEERYOYvn+Hlr85YwuB4/ex1TB//25kDUpg5y4LWa2CmZgOqkKWQQyzwGKFZ
iNpPfIvvcvyWeg33fZdJ4UMqHY6/AfqdqLNuLfhiQHBy+FjRurZm1jJHMtNv8DGu
oHPqjtLwrRKOXrHwx9uJRXLj6CdzLpSsee+94npLbkYyUxllrf70mh+Uaig4YW3Q
kr90IYwI3ZkPY0NlQyfkrgCblzydZSewfiOot5jtqpRQ02jA5AhV/PpSZVhlSmyY
M/0zNBPcc4z/Ns+QKv+Y7ssHVI45dYbgJCUDlyNnztmT3v23stidyi5iQAqQkF0i
8Y/sC7ItXVnD+At+AsuhewcrqRKeQatzfWozjDfUvr7OvJV7cAOmH2GCOeAxEhWM
dIdm+LlSLORkLjNj/KMLN565wuPme0n3DdmAG0/lVnjzmlOIBEo2jO/QpdSFxC5t
0VLeVp3BXOfd3RYAqLGHtg61X5fWJqj8Zm4G2A6BR1akYwMX8ITTzcNiEOatOjzv
h2g5lhGeGKJwNBUhvski7jH5y/lqro8V1dOSINX0nn9mOqpMqP5gv5tuFR7pAbJv
LRZa999acJ4HYgrhhcRh8f7gGz1gt94SUgBvYv2EgW/igsbGY1SxQu3CAg6dCr4u
QJFsUHvuqAIEsRYfN5DdevY4wqeuul3tShfNzO5UbEdxmlVoky4e5x/2o7Py3rru
+0X8HIMu+pmKXy0xQw9scZtV7CpXuEBNYcksuLJetv2LY4QNcv0DBIKAr4S6jCbm
VvSs7uGKC3ncFLBPtyc/p2nFnsRcAozDqtZnwlm2SEVMyLLcaDiv8d5cASLYMsYn
iE4GXcJ0Z8Wti93m0CC9e4TqTQvBU7zt9lLxss7iO/3xNZVH7rmjNG7ZfrfWuMGX
yOdHsGg510qlHhiR94SheIHPiJ+YndyidWY/1MZnM7oAFCcbTFG5YSXfUQPBFIyx
BUizLJg3sEIulxeFyH/7dfHfgdCvOKlTq80vjTNdFZ6SHpeJBTt7MpZPdxnt0qHN
7OwFJYCw50V0/hLmiZSHgn2Qo4bbjX00ecSnxzMB8sd0uf1r2Mk6QaIigNx65RJu
Afp9D3chKMbVuy0pEz/mC+ZV/XTgroyeXbV3HD7TgS4XaMwCxM0kpmisBjmhXC5i
8fMUXexCKZtrCDnahlsTXMKbbhgw9TquPgq6tP5KCIVjOLvpSgQifBNyT9120JY/
V61lUZIBtwxYnh0ui4Y+j86x3NIyAQJWkixDruIFrsLOVw+HNm7ygN/tLPpdxqGD
c5Sjqu8NSuYTApX76f3IrydvXq8AcW3Hlg67T8yx63UDJOpsRqRCe53Uywv1s6Tf
adEr+cMu9RnfYMj8afSFCY2TvYTflHBxirejLSydKNvdn6NfSEbvKCZwYArlksKy
vtBhKf7HOHX8pNoSQQAsY1eBSlIEf1Zlsg1NMNYY/kuUSJQ8lEHRJc3P/f3Np5IC
rtmmfNAl5940yD6aB5OdBj9QYOqZ9EP+u2P0VQzkzCek1PHU+dmY6l6hgaVG1mzz
fgutbOIgNlrs1Rh1DQp6gZhg09x1U6yvVlSt/Sw0Eey5NLa1AVbJ96eYi2I1ri2L
dIQs2jo2CJb5N9mXdV0eupmR3Bo63a3ZwQOsgEfOkVTjEsx19KtmThVken5k/X34
axDKbNspb7f7UpypQMiiL1+DSGXKlGv0qKonnHKaCILdLsQelGIyDwJ6P/OEeDE7
9U9YLqmQV6+pOF6BkgZ0b6fSv1RaOJqrj1rLWY5gcDQL3vML33ZKSnziuYF4HIJ3
9ZPpTcVAktYHf6O9iJsN7pkMdIhC9hXnCMPUYuPLciXMB9yWIvmSZyYpLvS2XYeA
D82u1msuNxDPkPPFv7VzYAiiGqYGhugXkCsJoAF0dJAkxPVSdTOfgD/1dMjgG5xC
VpHL3PEo7yA1Y8XvyLQkTuNnTDdw42UaglX6aTdBj9iYOlmMi7zaPZkfIWXpUNJp
VP+rk0zm53q3OTqLDKvpnTeU2OxWZCTGdO8AW/iYZNrc5hTc/Jt/XZiIQVdtZRCO
zxgFdPCxExRXJFjsWw2HomOEXp0h1XtGplin5jRanUGMn3vcoVHE3VSuXMcTWv3m
8MveqPuRZuNnhJggcCRltHCETHAdcOd+YvjfRgqRS4dwOcKrZ3C7jWfP8FlNcJtb
c2VYM50EHym/+WuhehPV2bSbIXKTEQqVzX4jnk/MtKjhfJeutYQhkaI+gOWy8g+Z
BGfc0AaVcFKk0zzj9Vvn49vBThVsLXdgAme1Zm4aub9cFkjqlzIDRsweTAyE1pOB
c8GI9azeOIAfTBbtZkW6iq//XDpl7tezqKrZz8zs2Intht11fiDh2nkjXvL7+Ty9
74gHZyExai08ufNmZx4gQQdSI+hqb9+0DJo+IFSXoO8dcqozM/u7PlFJZip2H4R2
753w0xUrs5rUu2+9RSL7EvpC6T/O+D6jYYt6PkHRH+cLAjHNzcTRQ+ewduHOh5Ru
rn83sv+MvcTafPtJJisxtDn40Gwtmrw4flg9xHuhu85mTXcAtgDT8ETWgcLWYggz
+xaPwsz6+DgNn/5NBtyVABTR9Thy13/AwymQjwNOif2hegNtc0rf/HzxHdHSEiqA
A9PwVNOIt6z6Y3Ra9HZG+DBP3/6MZYjgTHTwqOklOJOyfIWeDAuaIEEZQZs7GSXG
xTZkKXE7iw/DoSEz9eQdUpv9u9H36Im/pMMOrhZxAHkkRwVCpah23nAYNigrKZVB
EYuOaWzOWGFpa6A3nRTsw69y8MgXvbmyCypQlXeQXQXXxUEwpC9TQrr6Vu3do4Nx
ZMAQ59zEDlbSGqJXGzPfeFLpOgNmvXC2I3czkth0Q8f1YqLqOhmEOOnLvWcX3x1k
IYUVXpBUM2DhX/EJapgbeXtT8glXUGBm7RZyLy5s6Ddh2rmwFcr4nK7jxHwUl5PQ
MoLiVvmUyvreTe0IkPHLbXZRCFO7WF6Lljtkg4mBvmnsYF3PXF4iHuflHlLDx9/p
wfzDAdfJYT2gVoCUgXgzrT3Skizkojv0Uub9b+25oyLMKto6JtwNzXCyBdMSMh8F
zqvZJEkid1P1qVom54QwGMrVzXv1Pj3fDBiC2xK0TaLosSMkE829Ne7MAN1eTvMn
88S6HHM80YjW9fidjUR4YKtoFXumbbCjYgbbm2fP0CFQ8XnTNrox05T1YIe/ft+C
sQAMELkLqxfnoGAu2/Ay5Q6SHnud/MUYhkTUDw90NHiIWtk4g5/mPONmYedijkNf
tCQHV50TWO/u8FYps4AYyE6vJ10oSgbPDY8jskD8NU8wJ6LhtIdCHxhDS+AK2vIb
SnvHioiIw05ykzVK1D9JTHnoZ9qML89Z0Pm23EgsDANpC+zP7XZpQs2shFJ7uKRC
HhIDi8jNkLFsvaGGjOijXvNHOYnbCKkCTquymwrwS44J7cSFEzl/pzQJm5KWB+u8
oPKrDtZQs4kuy1HFIQBRVFQ8ado02Ye9o64fT1VIaPTLGSg/35AW9ncYAQB04TiI
akDTeo5vQS35ypBrnaZz6u5Od/KqUqqq6DGYnocdI2Zs9c557APiphhETS+WQsoa
APQsXcvMmAIUqvL8/shCRBB1GnLZgxhAozujQSpodRM9KugQ2+4GiURuVEy6HTWW
OSQ3jk7H1B7pN1E0wzOsXOkmoNtWSY2Je1BvlUBZ8Q/PtWGlVHE7g2Jh+w4v8pVX
OpNcUDH2QAU+keHoPNK9ZHSwo68DoNIYBWsyJhV+tXh00rWL0z77iwpLCvCEU4ic
fKGYT2ikeXN0kp23liMV+hKjmLSufIGXJEqjLB9xwKEb5iN2kXvpIGMsTH7TKwUQ
6Gzzlf02kYwloTLR8Gm/E4GmVPfUm5/LN8w4FyDq7KsxsKx6rB4HipF4WaBpBqtH
IZunp+eFlfdgSBU3i6rphl+XHtL4MiM7myL2GzFntswpSuCmUWs1HN9RAEOIXRF5
4VJfA9iRoIErOcJ2krb5fN0bcH05+ZIlQljX9ZKwk+cffRBzZ1GyAP4J+LZJnqv0
7L57QoKAvYM+BuCZx2Z2p4oACM0z5YBamJel9nwWsYouqL/HHsI71DaVmShv/4bm
iCNfJAj6Xi6WXZTJGe/yoZx8aK26iN9FjTRQ2EDXADLBDMD/EQvRy6/8miGVSJ9t
yPe+Vb1cVP1gJ/+cs0fz+uBuL/UMNzc79N+RRojhuSToTtjjGYdbIj2wvA53Od4D
v89dvuCGFLmcsfGQRIDKhJsKb79Di0FCQA5wV40oZ8fDdj2LuF4PfM/nqtVdbl92
A6vtfd1p7hFjKU8yhf5kD5jTEPowJ7NKK7NPJYOJlD7TtNqlu+1NpJ30wdzdM3J9
ANzKxwNuaglqNdZHahtmBwNaxUq+XgAj+SqxnxTR0Un73ecILCWNcdTaLUh0QyFw
JpRyaXolBIxUejE9u4zaXGwxrLCeB9VU8M6LAruZLYUdOZdOfqbQ1pzIHPEkVPwa
0NnvS0d96tYPpUGWkyGi/nbG5duXiI6gBgqeU+1oQK5QQDCE5S5X38wdmyG0GLSV
dxBqzwC27IrWVlERVJxJX+vILhLHAgIAy222vrq1/Epe1jqkCFutYZTC9rCt8pM7
lghm7Z7e8trhAMvSUZrAUaqqVDTRwkwWvh5nrndQhGtHF7jAD/XpTHz8gHSbb0ZS
LVY9py84ivjKGTrlkb9vX6tbjo2jLE29cNtDHjYgbPG8FhZbXVmiGLEi3749FLLz
Zx8RUswuAnR1ALpYrvVAOJEuDqgV7bPWClD8kYndSlT/AIRTVh/cOlqN6nO2eQLx
x0pu7ijvpCFTFPm5xpXxIRd+LkiZltjG6iSsVqfU/kUuqk3+KJRGk0piTptCcKv+
lFlTDaqkxh5yNcuk+XgrxQBjyeeCBiDINoPXVglE7Qrnjjjtj6sn41ul6XUYORPa
OYWuL8C4A3mVpX3y/49FDVN72526n1udvqgdVX9ITGmvNAHgtXIYVS+jlmf4/IDR
8dinSU4RMl1RQs0noCbsZa1f3tNUgTSETZdERNchSpQQqBwoABO/0miY40DAMOzZ
QgbyD59JXwL2KRtqDKZo7z0+V3iEOoBhReW7evDYxdnBHRgdyEK+2u4K7+FT4WFL
BK8gpfymsYhdf5q3/EoUnSb4VGBAteLXQotn/BW7xQqMYKdPXUIDkOZXS/lUSna8
+qRJVKwl0/DFxKmp8eft+Ro6q42fTeDedlZVnhA6MI5tOC1I4YWiCQ0/ZEgnEyra
eVL1AwKEGoziqaNO52CdV7lsimU20c4U3R6LIaxKntmIrNB5MGV6O3dTbIJzzxGD
wquuBOBWffihBDipQJn0ghY4SNHBYVNwpuzq23aXkwhJReKPnPh6iSKIlRR6q4j8
BrSPxYNIeHgkX93VgfiAqbvzCwhWR0RMKTDHUnsxiE0PIFoJsXiGbfeaLm6Qjo47
5KzFiWsDLzU3TJDJj2pQ1Kv1wb1OaJCw9/HAa4zc/xP0AARn23gHpN+2On7cehI5
vK39PO9E0fMU0G6kPU3H0KMm1u6fL6+G3//Sr3Ygc3Y7jA+J+deq/hx+mYPCAMGe
`protect END_PROTECTED
