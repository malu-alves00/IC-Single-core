`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nEGcF/TREv8UQq3VF/n5//Qw0099+B/WjZwtMpHIGBVnC/hsvkdgCDIudvXqRhR0
UfGa6F1mepm+G/zjTKmiTmncsYT2KlpBARjnPFMnjaPs1XNNqqqVMbAOVXdG6CBy
5FyPO0jiqCCFPI2GvpAXI0GsxpicHopd40UIRLM8fMF5sqVlDwOAWixEDgqpQEGW
ClXutH/FqdxA/5TFXil+J0K+Vcy72SQF8a4LAKIVDzrGoEHNYjm3ZPxU61VAInu6
Jq0VioV8J3P8ew9ITwuSkjNgro6JS/fR3alJMKAySKmljDWDUZTan2zNibuw1iVk
cz2MahTGyXlP2Xew30ksdEIeei/db3d0vRgPMPI00azxHZan3r+GmElXVgUuGt0B
`protect END_PROTECTED
