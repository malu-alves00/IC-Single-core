`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Fgq1RzaRd28Vl2tzgFCR1ttFqOTqUQkV1twEr8h154qZHHvd+JfQ3XO1W6jlLmB5
VLIpQgNJqt4hl64/9LlEtQdcyluDhfjdpwMM6dOe5/3xQFIQ2mND8LuanAhGrXbA
3lDSXwDPlRmJXSF5WhhLCleGONuq6JmkI9x6OTQAVBEAymPwBG6jAH+JpQWmHdf9
LMuwN6a4iCP5Q6u/hCWy/NH4d4g04bk1pb1dspYRMau5Flu9lV22QoATwhg4v6t3
sDgFfF/t1AZe/3C/W9dH1VHXRDsU1pwng82wCWKR1tci9svxbyOlfjMAns1+3yue
cyPY27XMIRSaebYQcO3X9njdYywV1kdmLOGr4sWhuIeSGVWWCnyliqHuAuyg5TGy
paTUFWYpDKFZI6dBzFnWrpEGZg4TIYQcEYwreTZ3Mt00xx9E6FAfy5EP+XfsNHD0
pAm5WU2VHAMCbhn5SmNuw/b9yp/KMnFmIk1RaQIuBoaNnjewUX8QajEYsQx+C5fh
IDI8+k4uSORJ4dNEyHYGBIoWxiYqi7osg0pX98MrAKBJXo/pDxcVHvHMou+Vpgvl
KoCqAwv6ZDagy6si3kSbY9byJvdLu0c08pLQerDAp39DDVkJ4B5Abr04yg3slC0B
o3Cw+lICv+h4u5Im+a5COEk3mLWl+FWHXrUVQjivJcDrWTTMBfhkjBqYNZXNry3z
NKNR7JXkNdmLeP7FWGR9VXx/TR8zxGmOsoG8n4N1ghIPPuSr7TMq6rvTAo2u69aT
3gzAr9oUqsJNTov0Lh5gNZ8kZJhQ7bzltWSNvJ7wVyQ13rV0p2wmI921iMbbGRtN
Wh8BXJk7Ng55iC3aCrTH3f8WP0j6Eg0h6J1MvE/ZZpxTskrAH2Pm9c51HFjKbdef
fXbAvR3U05Uny6d01dhwQLImIQFWGO9XqhhPUBB1r5yaQHL6Z/HebX3TsilRDU+Q
zLSAfJE9RvSWar/T67EAPbi/VD0UejRlDJKbe7RC4C3BZ+pez5RLNWooFx9g08TD
kzxpngURCdnsCFoP1X430vRkxFJ7bZfFUjM/GoevIL+Mf6hkxx4QkA+N6UmIfeeV
/ds0lPoB2qQbGgGDUHElkZ4NSIk3J6YkSA/g7ksQPUNxqmPa11jYvoRTfpMEVh67
1WSA7Jni45LGSGBIPz2sfnpkIfsN3GPx8u0aW54F91Iy8Q7v3qdCua4HoIHGQzo3
LVQ1BJgKGY4XQ4YOV7xFNWAWdXfjDHAS8tJI+kDpmBv7pigFm+o1pNJ+7gg3V9Fb
nYyooZeAq9xX8kiFFdvTqTXKFgCTh/tCjznMnsmn33XfZTkAycqwI3FkF7kyTpkX
6/L6CU++c6HJLXertId0NH48OE+0yjhfIKuJD+At56f/E8knwVhFAXF8EdSBIgLx
unbNsTNRG2wE26xWjZjVjOpbtAcEq96ojl9AIP8yio9Mkl9VequOliRe4PLvgC2n
tLCqJvOzzV5wrm08zw/bzUb6hs2l4EX/aQnplRYsCSn8ccQtPzPytKm/nylwE7/0
gC3ZqCR8bgZ5bkq08HhsTw==
`protect END_PROTECTED
