`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jSDSOmYTeItzxWaHnLT7TRPX1PvIJCYXfqzmDemNoDubqNyVRjwDBt7swnBnyao7
esLe0citwysFwFTxama87kvNYlNNe9C7p70H4CgyezHQu6f49EjBRHD9qVoyubj4
Th1kGLFNxXxfNH4S0X82PCZaqcRi8ut+7XRc1r77l2dUnl5MgwLyByVaf+iGS+XV
NLce9yymkAs0YbdxbJ6r2TkPKbZFZkxg7oweGA3/GZ5CyoJgUUFRoMwCaXc4ptFC
vY+yBWJLP2G/0RT0Kj0t3OLCTFVzthvieG+yzQabRJ8jVz/btBSGr9Hg8/x7zQuk
gnvWcm3xWAn9DxhMmTHrxvkxQfVWnI3hUsyHOpk8AHYJk0EFSfmVxkCsom4RH6Nb
bhCN334ZRpq0Xg4ftp4FGs9g2ElBxKKoXnxjMzlFQ6OEEiROFVtu2qo06Z5b0uM8
WFJlXPE7i4NbBzr3y1//9a/FErLpFTl9oktK0Ybo8TQqH3SfEfiIq7myw+hfKIW3
iEB0+3SgdKHgF82Qxmr7oVtLjc5Vav7K1PG8X/zda26B4p55AWOfnFQXuLL3kg1T
Q44L9rec6QxJAVKqBzvOr8XKwGur5NA8N4+XYo0bhL1jKUWz8EftUc3sCu4gBM35
wqF5NTBVDhGreVC1R+Y85k6WOSCWlkg+z6XntK8IDp8cPXQpBcfm+mnXPieocZUp
luq2wRV7XqEaPZpPtpk7dXADNeEc//Uod6eoyVUGM1VHG/s65VzbCU+5ExdqRy7/
JPlnRd2pVXLbmmvwKNyoFleqbz7CDt4gKv2O1OxCAv3ZV1EuK+CUQXa3MbolEEED
G5tJgUR/ojLNeDkY2ZdTZi97ipVewQShTwAcUkoWgGGmviCspUp3m2i4mvlixQ4U
mYetjhh0aIEgMuogm/mC0j8yzEUJb+7ErQhP6Qmu55/7QRU/e63mcgTqmJoQ5OEi
ibUyY4BZD+z8No91FvOlV1lF1GMM+1c/DCz3D9IdGgvMi3zOgvSZNPmcYSjvOKn4
fyM+bgd8V0loke4nx/r0kaYF6RQ3A6Uv73ZHgUdyc1lUWKHA1x1/1xeV9C/R1SCh
nroRSmuwtnawFcrjvoKC2cuON3XHVsVByXF4V3iVRp4Y95KXi8Pd3vSzXp5CDjDk
LhVQn2UoJ/nGpPU/2nyagCQ+VbH5N6qzS6NEMUkpFyXWAtKWnxvcOHyjSPSBF2mN
CAf1GWwUM3kCjDCQlNy7EY88c+Mv4j8lyuRynzF9aZ0fDvZrtrzMW+sxshDNe4p0
+BqMyM3+SUbSrfq39mcViCEVJ8A38GqdbAu86qg4Uxmlbz449fJx7yQYW7yw3EqQ
uCtwD9EVPRzABITsbBA/fojmNTcOi9FbSPM0IcBjBwWkPcUoNVR0laju0BzibE23
95UUES3EXu2BqbBeK8QqiswviS7KSMFRNhrQP+3Uoq3+P9n78dQkWqLyJARys4bM
pBBVD7YDUVKEpOzGaPV4/gYUmpHR/ir/g4CX6YPVWmVc3G8li6akVwZ4daAHcsZk
IygHgykGlmFyf3b7eJXQoHTcnDtZUrmOzAmw2wbRvzx2PuAzI9Pzvav+EryQEDlU
gE0eQIRGE142X7wUMz9GWo27SS1KeLkU3GEx+KMmBgkTi7gowrcwHK0x1Sd1cV1e
iQVKI7nzbkOKgaSd6zU87w==
`protect END_PROTECTED
