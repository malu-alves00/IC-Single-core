`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qq9AEee6vo62Wr1jVqjyScWqI1R9cAn75p80yevxLpIQtIOq9IY+I5Z9SdLAg6df
hDCSjPdVXFqYSf6Ei2oLWiSNqY1mMjeUNdiEFXBwMdUOIjQVvpQBn1lp6ZjU7ZgN
7nfpl1OKsu+PZma6KjaD++ffIQ7MT3qVNRqoTSO4t32AY8t9H5nqDMGJ80ZsJUs/
Bm9IKCIXGWxz53rgK/GdaAqm5/NIpu/a2/PnJfydK26X17b5xkIHA1xiNueW5Ogw
H6HtMXhBjD3lhJ5HqzsuCUZYCiB1NSBnD8wG/KmqPnIzSgSdZtK6THGKCoxwp+IT
7sY1mLtvvMrwJjWLZOKM9C6pECiSf1hvP5c9Pst91T7etjlX8roSIL6TNqouA00I
rsnVSKWVmTkwJknaCqrdxpAZKw/3637eu86gphKq6IoRyB8NmHAlAsSppT/m34nl
Dl8cpf9JNeRG8WBXzuCqGKC4XvzThQeZctgIHIfHXfYJJvXHIKEp8xHRcFVaz30W
B8E78sEEx92UO+xLPdo9fWNuXjfzgmGgRfywULZn7HkqdOmGGnlVMdKvBQaMfQxv
gRaTHCShLvl4/zujC20pkhhGcPxs0HTEOWDgL+zyMCH2eC+kGHHbLLYJeIewDLGH
maZzHWMzZArpVEx5C2KQX+KFwlzxHg21xzmujqWbpR9UCjymV473kFfkP7zskfLJ
rPxcDAYp5dP3ovRfXjx18S1SCShc7e3cX7Ro7QSldWNgdLTIYi6/bv5QeHfAwal+
FHCBEQX83GLbrnI7iimHBzAJcpWXjzyIUgn3o6eeXHM2dSlQZ03rIJBxmsd6UUex
dizegSWaMpoRMse+wrYAd1b2/xURJS1M7AY0wK0hNl9mn5JVtWDaDWedzp60MN7i
UGLZ92KEKibzBx0uumvj+C9dZwbPuT3mCOcYcsNyOu2SMzBSgpsbfNzQ7F6AbDD4
tDniiwS53AXVON79fsMA3cHxCTjJLGBYlaOTHFbNaj4jVnm1cf7BjRsl6ZYW10LW
K9xavYmpeyc+Ii/L43HlNQZ0bYR484gzJMf12Wxyt1BmTCGBauKcmi8YAVnbH9Q7
58tdV1g4LfFbf3+VSZpwCMoPkT8GezYfiWe6AQvxfGT9HWcdPwh/6+1AiG8ffowh
Nw18fVod1sCayYRUskm4a3J7juFkIZHyxFGnpT58gEwWIAKkloCeM19sytsXx2RX
sbAZ+36LZqmSL4MWUk8jTTNTRtN7o51EtyauDNt6ZRa2AZjPcswunskHq3TzN8Rn
b2fYsfJqyZvjIZVDzgDouQp/Jpd3WOdRFS0iZB2yyFs=
`protect END_PROTECTED
