`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kzcDegS50LKMTH25/FBNwpiDO+/d2Q1MPqThR44/miPzcYI6MVrvuWzLRNk7Cbg5
FkAEt6EApFHhBBxOrHceFYqSWeVcZ3/LJaWBb4Ww4NYxmbEmOrI1LVpXNIVgThn5
pXYtfUwng63RaTpGhdKjd3LgoInCr995hZiecOEpg+syM7FFrbcApUtUJahWJwQu
3BE9AkUz2qvAQxfZPot6PBZhHzBywu8wj/vVB5ceLyg49UG87o4J3o0riIcT4kyp
rLkxdbSaPFrXIKGWLkJXCql9JredbUTZq86ZdepeGRfHDfU6XEOLRdcMB8is9YwA
Q/qjAKN8hG8IljzPw7+HWN5KVcM2DCqhO6CRbB6TgazpDHPu37RUVTLn8KV6mY6n
pXsQWhNKrZL2tYydJVgHUMQwfvAV4jRKhhNDPrtrfubM/QNEDfb36ke90ky7obrd
xbxhR0BfzFBS/Fl3f1F/Wb+9H45H+gMbF/7zw5GY2QLpqYbicWh5YuYdGEDwYo5f
7pwGvKOw3coy+KyHO6YHYLcHfmKCYDyJfLCd2HqdW9AiT/qd2SobFy7b0ur7hXOh
IwayyNSoWx03P5cW3ZHFWvfONmWLEziZGPOM+1Uq2exZVJ1q47AA3KvoK1AWF5g+
VYIgQ6wDhtT3Ng8kON8kcZXkDS86IA8GmKiTDiyVLG9EFhVrEWfup4elgjzRJ3Cc
sU1wVnCsS+HAZ5PbFPrhhmLml/bLlHvpsjd2/1XJpeu8lMZ0BfKyAvXeJk/Ebeor
VWWvBwgUYbKd0uVxI6sIHXkRolSF7HqM/mz1ucxxy6fd4cCjYn0W8U99S7NR1OcW
HVuuUA5tT8FlBwT4jw++gUzh1gCnIXKPoszTHvwQ2w4ZpcVZoTK7D1eTBsFqDw/8
wUN/N7aJL+AR6/2MQeiE6s8QoXB1eVxvZf919szFVp2Rd52miLnZ2XX4XKAWaW5s
FgL46Wde79Q6JIS5ClrOet9rMg7DJq0+pUlYAbR5sHD/NocikUtM9G5XFBW4IAUW
nubPQc3u6kLCvzzJoh/6f0rnqP3z8T1kWowlz24+f1/oR4CmFgIbxgZ0OOc/Nidk
bLeoVqqVFRZ4I6PlVtklx6I4VK9PuzVB0idJzQn2gr3uuIzsSZEGP9hoomeTXMZ3
Vpmg8+1ijfea6CKtV6gG8nWl7+w7CtnPLymYW4DVDWzHBhLdlCeKCX8hm7/vak09
Mjho0I0JjrFt1efCJrr7qp9vrUWYJR4/AXfCt2V3jemsLtlIkTngtF195FFnZXK8
qQh13AISFcosBRclhpBo66WiW6hStqH2f9OzIs52Udh/t/+5cZI3yKhHicPcGgyO
u47Dwiow2fVHcpO9dJALeNmDveNYkV2vG26bkpSd6tyopI1Al8dHZJuh2xWjdCkD
Daq95VFhkerzVT/zn8ZV98yPTjlQELZElWhcNkmBnJhyVfvlCPjHI1xpn/oK2OD/
fKJWiy7Ay0P0TCJ38oRjjDdEIuwfjLbhKNTP//B7A8g9ohmXlZaA3DzPJXTlhL8i
kHfPJSnJhEsNM3hCQhUyao2dyXqYZNyOB8+T858E0ttTR9Y3AJt92ZV+IPMTcJ3Y
PHJ9ZRQzBh3LnmIfjGo1JhTsiJYe1G27cAUwgCbeFs0sI+9YtfmEdXdDAX/rwJQ1
F7P647WgInyj6fDAISnw1cVaD/9dNv13zubbsGzoYpRmn8QkbPvGa+DUfVCPa0S/
+dYD2JS3Lw9RmUvWOKib3gCohi+JzvAtf6NdGKbqa1qshOMJRQZGipMDEgQTKIsz
XrNjGFLwD3aIyRRGdZR8gySZ9vIDgCTpJra0tcvhsblmP0fJ8c6ZyF0bxVkYnCr+
CKM9gNUUTMhW/RdmnuhGfOArDel1QsIlEA8vEtb3KTEPTIvlvOjcYL/Jray8dnAU
X9tgvxV42GXOmI8d39GroBn1pC59DJ2L79NeuuDWh1mGcU3E/Yjj/21FntIcxt07
lcRuIijKD4f1sREmFfVuuyQUUnc57N1UQsdgmEuAaGYwMldjU5O5X8piLKKhl6hB
zq8G7Q0dw3YhyHos+t3isHero0qlItoL/xZ7fkkHos5lIucxDZE9tgchwrs8kDGy
/NEQu8JGUEKt0iShz0//vEnBuKEG8G16GSoe1X1W5uSbBx4dp9EyWZ/dAZBLakTO
9zEfrM49qD/wiaWe6Q1a5e4p8Go8tL/vbXGvBL5TYu16+kJx7ZCDfhF0FfkFXaxM
6sdWj5keZJtVaKZ8mWqizHDpT7kNx2zO0D/X1M8EaS4IAPYlsP5RKQYaj/f2u49J
GZltRBGssWgs5wqX85gpD7XpX5mxqiL5ybV0VPNy5E5CPXEYYX3Jj7hJjr/dWfzb
tffCqkqp2mpw6M7xb2Oshc+OVAPuLknDIWgIG0vUlDa4j+ICKNI/bueJ/q1h0i5K
BSml+CABa01T1psOvdNQ+iAiWSNURVnU77BWyPRRMahRlNcSoxT35Ud7jQQSz2DQ
h4+AD57yzbaTDqh5mc8uxp/6dM7H7aRpQxQV81W67tGYtQY1BHmZUzJkpyMTSZ0E
auYNPoI83D+jyNY0tGZnDL5kkXYRj6LfnpFbNsFChwosahzXHzElYjOE2ktW1gNw
m7Z7gapv/mh9i208cFPVXbunCiIFCWCGud8ViYnb0ruHALYFjHCYfpZszZvSi/69
PWJgW+NXOX6trvsRPLGJ/w==
`protect END_PROTECTED
