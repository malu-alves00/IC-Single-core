`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
O+MVvZY9Oa32PNL1NGMXl0oEIZkVs7EjDU3t/ZHf5Bvyra/1vYfOsBROF0B8NR8S
+OOMfCeLxeCkf61hKeDYC+S1soiV4vlFUf/R9TKzEIXBLbG1Bq0tB4QeiePQD8PB
d5LOBRARFPXo1zPaNgyVrx8Xmvw3wtAiIBfyy/UrRO9PFyTsRxYaHAiFqxphGs4s
dq3x/g2IBsuma4MpPbCsyeUnhFXIZEBuP7g5jDlybRdqqvwd1upbCYAy7l4Qj3JV
yLJV/tby7c3AcSO9B+nBQJuKP8Gt94t1YTPjcMxsQO2PE6uHseYcHHePNS836v0+
4UVLpKUlWa2V8f+BNcwYaLmMGd3Dc3jqYC9w0t4E8CImo1+aLlWmBJvRT2TPb10H
teZPo6Brt+nJlnCNFq48cr2amhMWXRCl9Zfi16S42lqaHJ/JZINBVYySb3Kn0MZW
`protect END_PROTECTED
