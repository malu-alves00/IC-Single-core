`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
A0D18hHE0FADIbFXctCFg4xvyOlwnfsRiIoN5++RsPfPzY9EHgEz73W1OTXeHnjg
Y57/m0w1moSEMP9K5Sfym8JZtLRPQ5BH9gjPDZv3M0pcidSsmkHdlXVicsmCrO2K
Skx/XA+qPZ1W9sbFvRzLYhwneIXLqb23tYxj1i3b/6Vtpjo701ZvTE0Acugv3N6c
tARI7CrFo/mcXj6W5qQH/WDXn8y0V7BtiEgQMn8nQDFPir7jFU74gOW4tzasiPog
RQCiPeuotoZC1zvdIuka/vGNkxyr4TlVUEMBimc8NiJKFl5FKSQzXvxzZXgY94f0
kHxMuRc03UqzWo1EZh/yF1ugxCIvmW+Ww5fwyg42y0Y0EId8coQHGC0wvcLz724T
Z9q1IO9YBnjWkPFrWxHIFhOelA3eMHbuR12fcmcCyak3xgf6XnPjDPWkqU3ooi7B
kQguvrI7MOXEyZn8QszvFOFcPaF/fO9H0PpHPFPPRjQdQW5DLNkg8XpffuVLz9hF
OrVvpfgeojg6Ru2532yX4gzWyrH4xk2cgYREsdZJ/FGZP9vykveLiMgsyFFl85wQ
gkpkg5uDMCDjnB0SAKPDdyqgyayLEA8fW+f0cbvlA3zlRveVnFqGASgrxLFj4AA6
S4LGOjfiqCsUTH7aMXiIYQVAejEm/kMiQv5Adjz5Jfs2Fu457Qt9dvBPA12Um3gL
UAC3yWksnGseRNA0XsWbcX7uO5to9OTgibqRBZCC1x8Qv5Yjmjaztz0J6t7Z98NV
qovB/3Lp89PtQtcyZEHd/jK8NN7p1SFvcNrvqw+b0M9AA7emAhyvhWM01vTQsQO2
pjcL+5crUQurVVq0/hT2BBqSa8NBuIQxdDUTUUoRjqHQHZi+adoZEC9mcrymrf54
83AuSgyXZUVxhLCpsJGH8M08Ar2omyrgs20DBRIxw3tLQnPjxMwuIdy8W4RfjtSR
hHFWpBJ64EY/88FITSpbtJqqXlbKluFLr4hPPD+CHaG9f4U/3HfV5223jFJSpzND
mLtbQXldGXwXcvkjM5bh1Etosh1RuHfUEzpG6rxwy4043rNwJNebIWfDWe7rJKmy
sd1ROCOxu6GQ9LuUL2r2eAz0Ti0VCvRdESUq9sqIEhRRJ9X02J39NUuAYy4cp43L
/aMOpQ6mli8yfH3FRZ3EvNswaX7EULHsLv4cSccY3v8w4N5cIxanxW9/tvL5/v3y
VFPgliCgJOZdvj4UbRsxbYFMTU6g0MSEPqH3QoSdfP6Paup9C5s2TUO8elxS1cQ8
0TqQnfBAWzAjkHJyqM4jRKjWYhE3x+UEPbftJYO9EVwSEleeBEz97l1hTYmn2THB
eGOTdQRpYnPRptrpwhh4ZfCqB6MkOOMdVmhgQVGbUebg92SklUIygawYbVNoWM1Y
+kY2/45VQCvHbkC+hl4TxgBiqOBMh8agjllWvJAs8hmDeM7HdnxPRBPH3U36NiIu
rqFkC91GJETQjvKILPNZDYEEyaVJnB1NHHyvzPTTmB4+TXjX0p4gkDbNW8KsaVHf
D4pXFDePaHkxn+oL/L0JKGKa6pNpKu6M0CBqarkjxVNaFT0BnMyqlCHbfzinOWw+
wt14+L3U1YmmQKms5tj44MBEe6Zo+wXHVgMHCIYB31RIR2Z5FGFRVbstji/MqCTA
0WUutev6qtCVygbSSGGzZoRAmFwiVKdp1pjGx1gTkY9QrW1NusAJ+pUXGD71ZZE0
GL2lm542qOSqZ1IfkvoOrXpq8ZlMXI81/fEGt1xhpZwN5SYwNb0F90p7/n+sJREz
ehnsFuECMcU5Rje9mIjy9gcQe+4DGCB45xbGH/9GrnassEybCuD9b2mKrDyApb0k
0Wo8TDCccWatcFJOL9M/nqn7nTFBzZfz+I+DiqUF5yGI9XrMl1NJJABjRNTnSol9
Z9a2BlEeKpdXuC2tq/SZnblYUmddsVHYRVwph8O3fOwgLq1zaJMFWC92qnKbJA8x
SWgDPU2NCoE5FVbOyEJ2yTOX8PAQ8cLE9J74CawcKb+65Vb+0w4QQnWJ+19viUD2
mul4NdausmREHrTANwdvXbflR12kzzn1+VLGgKLk7ypSxWNbZka7Hb4LMIozQAVP
ZxEvQRn/VMQQXe5UTtOkJ/D955eqzNZdlXbgGioTKGLUGCWPknxwfe7ym86H8X2F
3do2pGvM1EgOMrYzOyRQWUeGBJhLh2TH3RTgou23duPXP7EKHcJpM6i1NM4uKsot
0STEeUL1emrBeJNzfRvvbuuV/BRZF80vXV7t1mKWXi9ywlKQ1+HMVi2vEX5GuTmk
n2rZ47D89Kh2vs93oGeyqFwySqaS/PynhA+6WPE+a4U9yANyMxJQc2f78K95BEBl
HXZNhleVys91L6KSeQy/4sqKp19qKvLGZhIUv6a3aL7Y0rlIh6UKlzjjzal4X7uz
JrtV3dIVzIGQ3tS55h4R73c9QqGf+osC0BKBG9LwUmVptSqD6XUBy6QL0nYmKhic
Z9/mmNPMxHUtjpGRu2nVZSjy0wTt5g9KbV/eyR9MdR9f2gxSpF5wyOqTKBSRHK0d
DG+ovDoRcrupCYLZp1vYSldr+jJNSbrPDEFKpHPTdVRM3u38OgEowrtoS+ElaC2X
LYT55GfQPQDyr914mX6AJDv6PNTrlHW4GcJBiPv5moWPV5Tmeh4qi7rqUBmZlAx2
P8ZlMVB9/VZj6ruEIndz4pDptg/PiY7vrNp+NQs+ye03vwH2VPsalG37HcXrLr4f
eroPb4Sc431QAktEwyrIplVHVR+zNt4O74j3Q0qM4C5+0b8Ce/1nIlK1csUPW57e
zlG/gDGltViyQfE72n2D2NpAMPHK5rOvt3ohtNg3UQzJvqG3jIaoX20rvfvaangZ
/IW3hD6tItB6ajDY3fn4QACMxDEOq/YVSQvqBF7mCckmiDr/IvNYXNOKOFlI7Mlz
sN+4wNwP7QMhgWCv1HAH50FYaPwZfZS52sJxKzx7Xe0OW4mLozsQ9iPOrav+Pkol
LszD3X6nl4Qs7KlTo4mJSQR0mjrNVJXzDmNYKK/1eMyjuCkwE+jvOMKM8GmM/Ach
GuARZv9vfrfKrMwsoRkwP4cFRqneJUgAo4qwI9gR8Q1pHgZjLYvFY7yWzDaiz/TS
eC3oofKTMXVRNtbdZJrmNdz1JiHunsYfzjXxcuiep+09GvyKMQG6pUbIXT6eP3DV
oXzje+jGwJkQK5KlX9p8NAPcBI02tB4IlBgZtgqihhxHNi+uCtmTiT3qQNxSc2j2
bDDLsc/Pf7xCQolz+K7rPMXVLChVDJov3xt1rrRJpoIhksErjyJnz8j3bTcpiIWd
skuHyA/uaA21kw6+Zo9bAzeZ6FpNXHgtrmiDh6c9DCyyVFI3Pylz57Rp9Lz/VhWR
XObE9Ipv9+ZyuREx7kwAzwCDqJCA11GfOKe/1+Jj0WRYGjxPelptRhunog76815i
LjTNp7x+fqKvwCU2LmVNWxoS91l7lvW5sHYdFk4PxBH7TO2or+nYbqNKEvFX7NzW
EkZOULAWk+pFH7uQNk31dJ0AWO1jetsXDxJI/rYVRHrbaCBC1NlUdsP4ziyMMQZi
Ri/JmVFWSwvkKZ5zznm87O9pcy/mfj5Xc9kKELLT9mDO1IpdlB2o/8wTU3EXxASW
P6v4yU9ZtnSofVI9x3RQjG1XhHMgdkKCmEQxPmoUKzgz6ZnQ9KE/RujKXWRdsTib
BvDsukwYluVw13JiL3Kpos8JUSTyJMBR/iafmvB1m+UVxQskVHhJMMo3a3x2TBBw
K+kF1k/dFxJOasfh3ZUDzU9s8ujLZZ9OYP7S5qre0DUmOc//xaqbbmJuMZOpC/ww
PjWH2+FwLvBqM7zFWIoWS4KzWwHqC4UMcMridpvoOmxyK79PTo0aNlbfn/j1pmdG
XV0bgEpDhGjUlRm8rG8cIfC5MLieZXc3t0aUlBkLLRUanMWiFJw+MvgIDZGOC15u
2F+aFAbF+o1KiZOOpH6LxOmEcq77SdwrJio6UHfkHmz6ijT5J7PZntHmwYxgrpdj
P+Z6OBrY/3oWW7W32az1b3ZpBGgvVGqv/qpNjYk6oSJDO7f0UE0cLllWSXdfsc0t
C4Xdr6Itovmps7T3BToGysjgl7GhW0HsgJCpqHdXWVPCi2X4DtadrS9RWe4XU3cp
3fw/o9g34/T33/yx3Q13rY0Y8x+m51y7J5wqie2VSOXPPglXX/wXXD3rRlrJkLve
VZqyuSZ+z76rYituGQ5pF7x+64Uj1ofPywezVPvpsaGt6yn5ZNw6p0sMekmcoTaU
0vHR4HeqzS3u0v0Clyik1rVp1Nzf9EulB6lhdypCgoabmmEtZxk/WH7J/xmmwLuz
uoLOWQJFRKukpkyGpQxKvKEvlwLf49D/eT9t15o3rooqGLxcHnTS2oK3Xq806ANR
najMNzGJxzXEh+Od6wQanz7L0dyaAflnPwt6APHDwWxiC6iqZmemRhbbzrnea2od
FIxcmbypMnoEHR3Fui1ZQlB/riNY25KG1EC2HTesXeUvGwO/1ZO9LiTghEAEy8B4
UtCMSRNqyfiPZDxwDC/Q6pRdTBCf3/9ZqDd0khda9DsxPch6vrxbXNrrurn3SWM+
yYP/nlwmhj+0coIHEYDMFvwDaxInMywvIPAkzGwO0+lGIGnZGs3h5KICOybUZtDi
sURgFAEAYzfF11G6FzYrOTN7Xcey2A4Bkv2+WN+vhSzc8tJK+uHrNfFDi1iNTh2g
mPIyYrTzEHeZjYTPprza3RXVdOi3nYzwzqxU2bEjvGIXITtHHKGeYbz7Y4Z2/9F7
PzbsCBwAkWZefPF+JZr4pm9Wi9ehGBUFpYF2frLNqsAOCqf4oxX5xr7SVHgxbS9A
x4ayIPIPwQAXfxC1yFenB7l2uW+yPWoMdxDOgFvL7f/TxjfL6GomBOyO95jHNWBQ
MnoW/vx2acqKw2Vsw7cwO+/fXVUWn8XN0z3E1N4kGrbxWq+f2sPyIIgGcS0JQzPw
9v6eyJ6n6QfLELwrOi9YROOjWWHi72szxKRYsdhzudg5P7eMRMvxdj0VqOkVL0hG
93L6lWZsuHhxMW6Ho2rTEB2T38Z7dQHcoUoTKNiNEDeiFHRKPN7GtYoDIhHgG/sI
zXR0pDuwlHS0VGZ1bKS1Po3PydcvOOcJCCvGoAKc0EQ4cKAZjiuPZDNurYk1lTqM
hDy3RFIlKXs1G9KBjZp57g/0N5pwS2cl/0e/k7Jb9raRU9QzQz/46nfsVkBkYYbB
DaDQi8PQO0kvXplLZBo96A5KFGATaONS2VxiO8NdlXRCz5XL88vCuQNWp0Ov5YSg
DiSiSO9TxjTPedZIgryUp3+xCK9kuhkFajd3LEh8O6RS/y2u67qUwkvNDfOEM6ON
+B4Dech+i79pbkbKvLsUlPvRHja6faPB90/AgKryYYiIaeemElsrYqzRmTswhcDO
xsQosMVXtsxb84VTEKUQLeshLUQbM7oo1b4dPdowBmVaiA4r1QJTvgVztIu7XUBO
xVna227v8NrU/YVi4sSNLeDIDH1t6RpJs50+aY0UShufpxsWNs98PaaGGcJmDPOW
fh7nZehSyFtcQcUx2EGatf5NcCpDDqy7C+9/leO2RvGqcyMFgsLhZuXvYpg8950f
CB92VhIy89vUKz5UCzFO9Rnr7LZ7K5nESQwPUtFgmx3b9z/3lDLT6L5dHUFhsBao
9mBiu1r1WUM9TXyGopWpiGzIPksqjbg5NSaLKxJrjPodALfJZPjkp9livREfT87w
7rVoDZhiLMeoAE/n2u7aICx+nkXfrARuKN32QfNAWL8O4tNp9wyjrrdI/rgoEKOm
02hnveC/kUBlL6zEZ3aja/jQ5IjRW9Y9UYv52m8tqfBiNO4w3PF4oJs4+RM7ijZQ
WIDyYScNQiBxkGYmuE/k2kXxCncerwNYIy51XPYO59qiRENGhJEX+Nf83gjLocsn
XOgDirBCUFOzMoJJ4UfAT5htpsUCGZIdiBaD0zUvxWWIB3WG9x91SVaJgdIG52Ya
IVWvSBKI85e4wuxokzLkSFCitSYewQDnE0eTjWJY5s674m/OpV9bWXolUa+h5bhT
n0IN7atvSd2BCKspN8a9bf9GauYahSfj3D0VWwIopA9MttZRqfu5rC2vwK63lFuy
214888/Z/Pd8NFLIvM8BEV7AlwcnCI0gn6XxUnqnKdr/aCaDitt8Fs+nARyWm5OF
WTwZOxz7yZUVNBBffxDmT6DoNuIrHdPSihZDhEwGuLS55SGHbjJSo5XGyf1yfnZ6
74XMfeK1bha/aRh3Nk/Cj9egb9uGL6fAT+p940UKEv35Uo1OklhHNlYOYFAZoSn/
UuhVjbZ5cd5J9Q/BmKJDZHbMzGY8ho1julVhjCZDljtV43bKrdBLBMfjyDTtOTI7
rDciOknB+3w6ujXYut46cE3pbwthegg1ffvhFq3sBebocM4Mcr44JIrWx07FJ3tf
tHAXXVBqgL/2ceCglCmM3IEAHfMvfF80K8Ma+INgCoYu1tnD9vDNjblsmeFemo2C
4TX6jOpGTrP7OVVrNfKSCwK0+IgVTj/CMJlmlpkFviQoIRc9jgre73JZk/8VD52a
chyfGxvuaj5BNdU4ODShtP9BZxbh5UOBitdAc2Z4MX6RDt1bLHy/YQ23utLTXCrR
sdFKurzqVaZwiqjwD+86mNkDISKBvLaEG4tesW32O7nG68Zc/fFcke+dFNyNm+cv
xbwDM/3rphmcXuUBahnrKCxOAOWW2vZrEK2X1HJhhnMz+kvEdL7CCFgbJxyKNECL
EuO+mFy/Ge0cE4OYQbeoE6Vk54/ndlg/YKQDST8G8qRFcCo+GsORUT2Ywl4t9YBL
CFrgBR5PhTceNGQ48u01nk87ETfp1jaQouQ/mCmKODnFT7a1oGEuziGvZ8CPWPCr
9MfyJbsev0esGoKbJbssg4BlmcGYoq5W2RKjygSI/ErEsQztuoAJAGxeUqYqdkpk
6XcLm/iXEfO4BmmS2wipGfq1tvRP2wuFmObqhvzqQ+p7AckMF2vNMUWSjJZTr4xk
0wwS52PGZmniPLrsL15k9H8sP7s29rUC1qeAOQ8RukcfsBcF+w9Z0LuuaF2WOqDO
kTz2iqw+WTV2zlElYaCxr0rudXbkS895wQopRugI4TSaXXq1FxuaC+wLDPLLE1Y5
M62D9ecDubfCQ1GYpRJbfI7tVolVdJEieidzEJ9g0yvCue5yIWFEH0Vc/QM1/9X/
Oi3tTCy3rLcL03vIFbWXAmoNcka/7Q5SXOaSVLI++C4rwG6beHnD0R+TIFrl9Y9X
2GHvEAyEDqeF2MJlovTQ3mVnMKkkDH6yJ7QYSPLMsqaXa4TAztp4ROhdlIlr06DV
iC7YZDma/XJzhcnyqyJGazDlGKgidpMT6qMQV1jSm+xQ+Wfp7yNtDiyadPgCyVcz
fpETp8fvBJa0SiEuhengnQ==
`protect END_PROTECTED
