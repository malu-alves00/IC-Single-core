`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NY+bCinLnh22JX1mA/0W+rc1O9/q7xqRBZQZYfRfA/MjhFyJsxb/rPlvdng5Bh/i
MikyW9ERxiBI7Bne61bdfByrbt61vCbTAICNuwxzBEyRK8qYum12/wbE1/MwcTTy
GDFo9Tv/XwtY18QlJUYhH/SL1nkkhy1T0LswpjpJoZwGOErSgW7bUZbvA+OCCP0C
OP4i3pFp2NDU872gdwm0mWmQgcbWF8cCcaBZLhbjuHJK9IMfbsZs7G5gv8xcWqcb
wbN4J6ISULXkJVa8LEnL8HjwXpvAgfIgQtdg1DRxlKXTtWbNVoh2474QlNK5lIZq
4zE5+yGomu3/JvU6jrGViWgXqOBS2ftdXCePd3cdquPStDekND1zBNdCGWCZ4PC2
gGpUTaKpImKM/5kJHx3LalIxr2gQV3+WyZ7atvGWuzOynasnpTFdQPvp+FDbO373
eP1cKoDscuuDuuf3qXaqnOnAa7Ow0wi94IsQJRkhTolKPNy/Ib2Msl3Q1v4+MDhc
qNvKI8hB4Oe4AEyU1hBRgFEq1gaiDgJdI0sJYyttYnvRQ6V0+z6NBopDdPszFlgR
8VMaakfE5yDLQtEP61EEDKj0/WDPRp8FX9w4B43vmYv+rdFZ5JJdkHqmCfKp9P9q
Ly/GOzG5jOEC3L/eFXo3RUYbmARIVpBHlhK49vLUm/oHX+cZOUtOGdK4MUHAhnB5
vAR1thTV8PO8BkInnTJiERvR749Ymyk79rhTY/9uDXMoi41YGSAgXEMHcWvWolMG
OK34d4r6qAD4ffaoVju3f0PQrb2og4JpG4iNav4kg+mSm2dymK8oVAbsfPSkCdZR
B0fMEBFgOwzK5QiS6G7CYmBWSAzT3A4pmHgEljhYvXyp874cysXdZZ8YroQ0qy1f
cg6hZhYLVhi4/oW/B0EhkzuTWLe4kxWdqog8mlX57nFr1JeNWaacjt85O1vGvI8c
YEp009hl8KpXWqXHH6YZmFR5Gv244zoUaZtlnsoXtVj8aJgicAx0RBTeQ5l2F4bR
WMrIKPOpSPlIByPX/80sQzTP2dCkrN7lX85OkdS1iu3gKt/L7HiBl4WE4++GQAkh
2Ki8zMO3clXPmxMWktFXoBesU0YdS0MEd/hTvZWlNpzC72dmfuxsjf/RvmVXqFe2
Yt72uo1VvxHG1v8EHVhngNT6k8B1C6MsQpnbxQDzaoC1GW0fMBzh8ZKZIFp2g4gx
KS9+gXNrPX8314u6DaF1tlp8OdVOkY44wrWJIENOhrw=
`protect END_PROTECTED
