`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6VWuPH7SGImHNYB8YMPS+lT6pZlDq96uvpSoEtyVYmQME/xfd3w1FcSfXiZgH8cx
ddwgkvnRknQEPm/BIu1RRsSs5PWvs+mfEfL+if9wWehsbWJtpgI8bZifnddOvq2c
yb8shitZWCOEAq6zGxc5/mRnOPbWDkFFwH7MSMsVTCGaX/3xszDQLo9t5bgiz8kH
AI/6j6h6oL4ocyg3g+JNFdMxHHzicLYea4NbMD+VNyBxOJpeHkbuPmcvIPBkROJ6
cvgP3mjgjm51w/Uk0ruG477EHn6oakFWsll+mT2vGfcAWmc20lxaRVbn0mt3Xgem
/wn3SaGNhgz9AMU2NSmLs2H+PjVNcgx752z7UFFsEoOw/AtB/p27wX+bF831CJii
wZhDVgaOR59Ar9nOOBECF9sCiJs70yShSx2I0zaUzZJsjbAF5laiOeTj8JffuVfJ
EFplCrZjyEebbRQiWwiZ1nMe10lE9jcmt3RXW6+ccJQzNtSFBJqV5d6ZPVzwfTE1
E+Sk5W8pgQT6lgtkpbb78q1hMhUs13Lj05ieLDQF2n66uah5BJjAehpg1+pw8gPo
Y52c674exqxp31LjVJDCRgtZsYxpkYCJ9qpgfFZMLq9/DV6yQScR5jHdbWPz84UO
yzG5gKI62KKKpTGQVZuHDKxnW7pxrvBBUdXCxqx2KZxjwB6FmIt214BRhUK8WXhs
32n5LJofgtijWakQG5PMC+E2PDUJilxebhBYEQp1mjxH99xHWIBTX07rlLR8jNJT
hHMI07Rug7XD+qgWEObJklhrH3Jwd48aNmdGsoPmIw2qasbQVFmH2EWI/xpdN7pm
aLGdghA2xh65FOlez8P2c8u9p+u2Y7tfW3Vv2+gGBR2nczHytjPTbCL/TFr0UmS4
+F0KOPQpY+XgdLymPqvwRsS3Ltpy07KrsSLfOuPHXWDWnh1GczuAs0FsuLH0Er4w
0oVdzE4barS72hC/7hPCKw==
`protect END_PROTECTED
