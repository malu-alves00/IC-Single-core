`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4/zJkMcKLwcNqEwD6Z2g0QDu27MUvJ3gOxw0iP0UWAn4lO+ITwNxTTNpnLGZqck2
TVmEcEmgwtMR8j03lEtGayU1IA4/VDRaV6XrqguDfbcqgj1+zMMiKcmhUMYuaAMh
/+SLNUsEuQ7P9k95fKrfpnVfjKrsJ3ydmtHpeiB9GSd4iGJQiTmhWvHSV1Zi9aL8
u6CNSNbuyLjIkTn29TngqCpf3qD3dOWVfZK6YtIosuLOYZuz9VjwFQoCB7n5CEqj
SAo7Ccx+aXFmP3vm81Tz+JnPBJHgvrn+aa4EmcAzPUfoXLoNmmSk5jdIxnrbIWgT
T/S+8UzAWKTn0+OlHU68/Fbi/lu+Uo3PYzco0pMhNQA0Qq+rsylZrgVGR8sPR5ts
jt1aqn6se8lPC1fxhNRVnL31O6+lh5LHNIfScoRxX2wyl4OAhxRaXOhyIzIoHOKT
DLPAGqAgnOoh3G+2W0IDO+Dxh77+yTqDFmX4OIYpnHgZKnbbQnd72qXgowHhAXLa
7sRfeozgObGSytnP30vN200TR8MYS/w1zyNGZfkTqZC2x5O7cl7iE12eX32fZ8rE
kQqQggJ1+DmX9AIu2yP2yIXqnHC9FvlkKm2dnUxxh1oLEsFdDOJa9dMViJMZR8U9
7s4MeW1tCpHQrw3ISll4nDeIZsn0nRo1VMwSW2YkOHB6PQ0PpalXQphzzu+/6om+
laM1UMUrmDsU5fNcO6OyDffHQjOMdc6mrB2voAid5ZvRWPMuVPOqgygcHxqbMNQe
o2JE7rHwv9bq+lSzN20lN9l8C+pwtmQN4BLhJ4Dv1V0dJAgzI7ieF+uRUjbychXb
LAyCSi5A8x4YN5KTZIAN57vWf6tzD42/js/Tkmv8KeX+FYVvpH0wIuRZQIUK4r7E
Jj5WQ8ysOQTNDTzykuiDYtei9lFOQykRYvTpXi/w3W2EW1oWfPw9lj7VfppCfggZ
L6TkUshUErCRwJE+jUCGfz6H1JUnp26qTj59bNDNL717nA7Bbjw70FDJu8RvanCD
MUYfC3fqOFRPO9lxtJg2jzVoCpz6ayJZw3s9vVPPxk7/TKUAqyYy2L4fz6S/TFyi
+O5xQebKhxMYp+CcRWMYWTAQaHCqdRLEmJvuLls8WQN9UAf0MwssPSCYbUEz4O+I
GieEbPciNZ4VZM1dkByyOMqHHXdTnlexsNNnCgBdz2VFbyjtFPM17C+EZ9Q58D0M
gi1MMSf+4pqG0Cm05dViwQSMdAYB06+S1ysfsyKvxqcMXMYcMApv9RwZ0AFFgxAW
iKN4Y1uqNOEXkEmrJXdTaXd0z9bgVhpO50acmsbbbanJWavxmhtGxGukSyn2/Hso
ugKrmgmIEPFnc6eEntGeIpAtafIzN0rN18fOHbWZQg9XVnjY5PMwoytmzjgNZ0Sj
D+FvCMB/4p1Me026LZX2J2PtM3OXdHliqDi7EfaStonKCbH9hr86QjJSPp9xDk1O
FUz/2iGXjKgr5DH04JCRGXF2/1pdylEoPMBBJLFuBvy6ztuXRY6PJSrdmoRNW36J
iy252uz+gYHKdL/zOa4jAIlxy039Qu8+dagVRQW1xV50xhHdkFmtCDI5fsnjhN/0
`protect END_PROTECTED
