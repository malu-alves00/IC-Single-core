`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aKMl8LyJkF7BcS29+KJe7Ayppg/LKp+pF07gQTPDZFao0XutVFcXOfi5eRbKSkbf
6j64AkSBnWyfaFOIcNXGrnC10lDDDXxCZtDh8UCwZ+UxWaRmfeovFA1zVptR2Mur
rX7pYoduQ0DaCBFD9SvFOzQ4IOVVUkSa4k88aMSzJZyc4jL9IFDvlPFWveDRBGoL
w1dazIfG139bS12gAR97JftErc7AakqvzcKEfwvMO/SiTKE3kNWgGOoWk1ur9H0w
CJgEX8jS//lzNvCBsTmRYo0j4m6q8CkHSfjfd/J5GH4cXSdOW6CEnYODJtiPfYCb
bzU5xDSNCpDXwV9tEGg1FaOaMVZQF+jd98hHDOxVkTKEpoS8Ve6BQ2+xJaxXQgIY
X2arfjR17kTrAY2VfihO8AK+E2C2+GZFRuG8Tm2vgN/yZlMvXx/LMTvF60LW5/w9
bOhWcOqM/0kH5tr/8Z6cDW1ad4lshoCmPVnXJfDP30qzw5oCO5uLYWugyAsIg/dB
pGqPdmiWoODBfyZV4q2W/nRD+14YpIXXwcba3QhFk+tFh1kK4Nu4P8opQ1dgk3EE
UxrWb6w+5BEPu/t4U/NRDMXqhY5EiRCf1HDcaFdYjEA40zKNI2RHO+xm6n4iBfzg
01khGtuFAJaYAt2WceTzXjZCV/PBa/DEK++hK96F+UdhG+FmopDzYSi0+HSqtsYW
V0tbbgiEnQVaYCM/4zxuxIZOggG7fJcvgEQWcppZdRK/+KZ/NrxteREwMy0BnSZQ
w432zFpiijaijZlqalgDri0V9GNhNLK/TEvtJbuvD5F1xZtignF++dsjalBoZ/ji
5te8/Dup2SWoLa5ZbecS/V8aMe9AJUOeyMxWgyJx8wGagsFerjY0L61+9FsjOQFs
8hTBZKQbC5K7F8Plm3/H+RHHmq4tr8dfuciXi07PLKKdAdfZOadKgTVaPplKSJvz
GNahdiLgNOs/MLnKzhq6UL9kyaUtwGjsyu2uue0bRngVMUANm9bCsw7IeyACKBGo
GaFvGq4ONA59uNKoSE0J51lMpuoaLVgOmR65CTGNF+se1iuWrGq2GhhVlpCygl6G
EPP85YXaXig3UTQ6mUm4H6UZjUFYVxsqtoQUsXgrKliqq+0SJQ3pJhBJ8RJkOGJk
uIbJGyL9qotzwGDPTEkLC/1h4SV1B8hDsoBdhpxM8TYrFygV/uzbmC9VUUoVbPZt
WBea9F3ZFvGrIFa+xMniVK7T3a6iP+AupEFBUeOmdbI6T7yeCDGJoS4up1NteF6X
o2WXGx5EJ/0snimYOQJBTJkAqioQNk1Ya7migO3l1baJP8E9ajeNTpCwxB+h5BOO
nlj8av08Bscw5FjhYxm2CvuBVrauiMMHLMAAN5CSxERvyKmb7UolfuJoYv4R8GBx
sztYbDHBWkbSbE+fbJjRtqXON4iivAxlvb1ievLu8NdTEeu+pasumYBMLKvhv0Xw
kbgZ27I521CYMpeMjRtjipEYHuFeAFnrgABihx4+j/pqNRTwyJSTWLCbeJQIfmD0
yExkf0cdjis1R83BFg9qhAmUYks+abxUAJGMyyie2dn058IpDoNi8304yVgI9FKh
RNwGO0/B6UDlDYTkNHsTSw8PI0b9xUkbfC7DRxl8lfe3fak1fVcZxgSvmxQm8dy0
5jM0ZIje57dcVFcFUbYqPrLyGPntoO7OWfcMCBb2QeRc0txUuUDbwG/XWg1B7mX/
VTTKDz230fID48jOQFbvQQ==
`protect END_PROTECTED
