`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1cctAy7c9ggrqK69prwpq61TP0LN02h0lEcnI4bZhdWxolTj4hubwMTdvIYU5kEr
B6L+3ACf2Z2fYDtw7KfAyqHXxBkjXuu4uulrfvflWzhPE9cPAOsev9PQvQvlhPqZ
0kyjAvEBuaRPV61N75y0qSK37nMvfh7amGlSLZe19zzTpPMcDL1/rW5KEWMqwqQ5
wIF/DEP166kennoGfFeRihzeCnGfp2ZTI9TvQUJjHAGHler0wTIEy5BFa1MyaKzI
McMQIdJcMyItQgm/3mCxf1VZbk+Ys96Pdi82HW3ny5QIyynNpELTNan9uxQpHIiz
oEi5OSAml0V6i7s59B3R1dWDmwVYU2CP1qvvUvv0wemiRJLkleaGxNVti805nabp
ZmhsYaDuT42tHTdu/dfAkx9bEzqfTBP37VHxQGL41BGp3HjupOAt8HEsuso5ycT2
0c9ax80VfsraoJOpDuzJodfoBsDz9LIgB3+99goi3Q07wPbaIq5OVj6f3UtFdwxR
bM4guO6TaxxjvYmPtmfxibXCmOe5o7JAQx31RVouDSDJNdeIzSOCkRBYAMqsPCI2
LVSNc7p5vtYB3JS/gRtUwEBT+d6sRlQ0HEyZBr3jRGTDxo7u2Cr2s5NpHkd4oqqZ
NvdFNta3QEMpf2nI82K21qeEMaydyDmrD3A5ohI4JAjoAr6qdb62Mp6TIykCmg3X
KZ9odYC0FkoDnSf10XcYaWT4tWoYT4XLzs/HGoQM2bwvS8paNlE59UQatLhAnIUy
AqonglBCDpKPThMDrqv6bg==
`protect END_PROTECTED
