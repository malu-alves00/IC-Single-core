`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Kkc9ArindD1AvggfNHhqs2cX/FHMrB52M0jqax1E3toL+DX+VZ5hQXG3jYvdXRs/
+7qrdI6tlJJ9F1qOa24xZht3WzBhgjjVMK6YJx0cTcukhbalqHnckvjA5yiRXAAL
+6ztOoqYlP2mycDfc1+GrgXsWzqMilEIdSgyPf6oc431V0oHFZelgr3QgRTS7+vQ
LSxZYp7z3Tgmv4+MvmYyymkm8jfuozabDBa7mgxZnjgLs2LMe+uchA2S30vGFbOq
EqJs4c4hDP7DoNKiqaWN+WhVSb7Zr0JyL444uHwW1aMUpMxFv5cSc+gxAKVQ9Jxo
L1cu/Vdt4ZfvwZfaSwTL1A//3raFXCI2jmWDSGbCkCm7ondRcmP3bPEAZ78+5tSv
9d2xBmIRdflAB0cwd8sGUIZnYRFar0NPbEjNM+XBYg6I+9peQBHl2Hp2fz4oDHA6
oB2EkJEHP5RZf9lbFF96OKIr+v7UQKFpSy1R6voCC3AZaQ8ViGkuX2jErWmL98Kx
YHsshzaHBL49GU9t6QpUwp7sPYT6wjzunlNkBnNpv/kCEpvLP9RhUZLUlFCIsbj7
50jrGuOxaVkYw7h+e3Rfhk2J3WyMK+EGYiifG/BMz9cT9hcPwCiicWpPSm467WAR
anvp7oHvkHMnYZwGkBJnX/UEzabU8Nyby0jm8vZFfMfZgrbtBcSpEuIGyTURDkme
J1Ezmec6OjHwqJj2DwCnXMKxq89dXlR8NIiiZYo2L7D6V9huliARNMYS4MBjJzly
uJp0JHeG5Y6mEvivY/HsuI0rgBbSOED82Z5NOhwgGVeElmlg4g1bfQTSYHtVtCNL
haJMTePp6i8KxVD2hbuveyqRjXYSTOUnaAUKzhrQQApob6YOcoJquex/ZurVcJ7a
+3NRqnyj2Lp1KFSpJVfqkvFgFmfA2cUGOX1eU6kRHndWeTupl+KV983NheU/DpIX
mtaucVD+CSMCeNBxB/ZH2ubWzoKNuw7cziDM8aDz+n1W1hFThGzzkCp9YRZpf4Mn
cwt+AgoShI8maXZ5ug7hd7xwV6H75ZEcGNnFyEFJeMEstEvH+2rYb0IIvBCK0sjW
ZvragxJuKTsx5ruLCTD8u42WP7pg/sjV2ofpEMyM3JjX450w/NDywmSeVtxYwheR
5tTkMtS+9NtLgOLLCAr2DV852OBF3KcfdIOaJDF8bDABuxqQXqywhzUcb53FG9rV
84hGlPCKl0qbwwvo0ZVrI1aFToiRsv0bw39Ho+SaxhvE64SvknaBSPSghu/6TbOh
Pu+MPjKnm08zMMkCTeN5wy/vddbi0N7ZRbTsqVcllmKMBK/vPZpUXCtTka4tKWr8
ojsYHc1eTGQYyDHX/qmiPhV2+nriv4f/sxO75OvrSmpaKJsfaaiuBDocsZeg2MY7
ioJ1hGH9ubJSRoTbihfDlkcunf9+Xvyk6y62nDyoCX8vUDVs6VhOQ1ZtiEA44RHV
`protect END_PROTECTED
