`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Y2spoDGn7ezxuzxoapZ4joD/BuvKSDIT3IyEr+Yo/xcJ+zx3IvZ/FGveaWN2KMPs
Z/DjjwQK6oaDw0GT6kGUjGIU9bONWeagEClUJ6dzJ5eSZSAgYxyIFjeC3hUPMH8y
E67clUXJEVuYgUO0rmcSIo4oI0YN/Tm7bif0pTVXIHTDiRcWGi/7b2hAhpuuxjC3
yGysHRtQqobEgDouxDGaYKqOdji2wo5dMvEp86W7k8uR9K9uSd3XZQ0otNlCDXUh
gQZYTtHyNZOTnQEVYNMMO6ZAgGtrbVqGurVZ8WRzrBopKPhovQSb0Y9ThZP/gIRD
pG1VBkv4Gp1ckAtuVQnHfV+NtnRamGt4BJU2pmGmLBf7cpjHefWmKw8XWbjynu4f
IjuncvKCTQjL3m6eoDztUi7vvExXtgADD+5BQwVPCm04fx4Z6gv+hpGpzXf5zNsr
LuT/HW7ouRVS9jIwmht31/ezlX7ILGHtOnk2eWY5JRLTTZEPIvMMeqU1NreA2QNa
Clfj88A1r/Kk+u8scYmsw1KjuLyFPSgnIXF2jR5f+reh0imSDeBC1QZ+jO+l77br
ptvgtMln0UqMQsN2+Q6QafrSpMF0yCbCzl4ASd0vBalmpu8PbIu+T5dTOKor82bl
ZlwU38CGZQk3TRcAJAwUdVl8GBKJA1gLvwTv8G3w3uVhdgaCkTI7cS8fRMnGTQpJ
dyboKAXRq8cJfG2/Gmu5GMUQNmhoCxYfRRC62ySBESM=
`protect END_PROTECTED
