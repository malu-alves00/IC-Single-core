`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fM40njLuaLndOJzSYRZvEMxdolFH+miONPm1hy9y10EWwwNvnNi+e3NK7lUzPkvK
wGEhCfw88s/Wiw+XZrRYCd9AwJ0nZJmPYcA8wEyiXjEUXCSv7MokbN6xvfUfl7Sv
QQ1XCN78DFQnJ82SPlFRjyzgf0Q8SflZU5/oM/VFwjMGRcAbIYD57WIkMN7yvwkd
tCnCjB34vyrox/EqCUynSz2KkPuOM0U1GiZGmGF0SqgV6x0nhtoAeygUHvTgAlzQ
MqG/+Q+myLblc7s4NL9+HdKjOICy+8nwgECwvHQrtadvgg3nBXxJGpE33ikR3MEv
xZmFRL8dktFK7qATsZ8D+0g9rOsHwyaFwppopCdmkxjVPg8hdVoZz5g4+0++MtjM
sHYK0lZbPEbF/02+vlhc6T5I30oMgAUVp1eDMmQEgyNsvcNqrkbwcotevTZORT3d
XAokhU+xmaSx7AG+8ETlWA/yJJx0cGmo79+9xKP/0YSxZ/PfirNWAA3OXnvs3QEG
p5qOf87269arBvyHkbMUFkGBc9Mirr8FwGCFsfj05UbgMvNsdB7lwIrk/NJoOPlv
EaoXHiMA6GDdEy1Dfcv0BH8F5LS066M7FmFhiV5RxOLyqmHZR4E/ATMCvmfTYmsZ
FJW5NB5ssHJAC5pseVZTNojDHEqgTVI/hCYfapzPhe9ywIBC179OiM+hi3yBhDsL
BF+Se3AinEB99EQ54NW1OXtrlmcdysnQEb5rF0rWIl9J88gtczry224v/3Hiy7rA
tN01DlwN/yfQbLR5a7Disho3voTQwbr8yWuf+Mve1c57QfOSNdpjP1vdjvtXwbMX
r47XYSCDBjacNKRtNXvrbYY3ENsXHNO/po/Kqj+UaS7XCYYBFQ7BDdxcMg/o3Gp+
2PjOT42vEIiGZFuSA3fOpfZ67N4GHZ2X++yoH8jzpwvBOWXrbLMR9+wBDAb0Lg6p
nUtiR0MJZ6Z9mKrVql4w4oEUOytfU+b0JKCOfolnX7vZL1YCKXoAlCshhr0doed2
fvEqSB1sinXr7g8BSK20a6KlDpRnRII3ZI47AC2/RfGGbDlrbCHRX5QsNSC4raoZ
QEY71ZqSEnxXoHwOI38CUhHi4h5Agrhd1eW8eVWtDJBYwgjYrZBn5a7/qR1JIggs
MLy8sR/wO421J+ikRyR4zPY0KAY/APqcrNz/T3L0MdJtUoyXoZe9rkjRQQouJC1s
HE+1OmAY0cHt/+YVauQQ7F3dKcUVCpUP2LEWeaSmwi5DOhupCsK9j3ZekX+jWaaR
BOa8PCe+50h6AkQHSOhENBPKk+j34I50TWYzyg04hTl3d+/Q2KVNhLZ5wW5HldsM
PRp2ZMA3/RXeUUgFzEUbQqnp/Oq2KEitP/3RyvOblt2i/R5NfosYBdumyM2SJwiU
5FhpIH6qO6E4QK1R6gvDmtPVALwvd0F1fUZPaqe63nDLpWEmtoqXUz07QJ3hxRDO
`protect END_PROTECTED
