`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PicaziBrpDIRW1TouZAGgMDOZVYwiEt7lMYa0NY+SDUDcwYNTGU0WNfEJJcxr77u
L6g8S9IeErYfOj/Cl4J8IdBptkPgYURYbidwUGTMw3anlD45nQZrlXjlVaVV5VWs
olKGjvcUmuX2xCI7qXFhyR60BIi9QlYdfO76cWhSeJ0mtCC+9UXHaXXA9XfVRXdq
PHK67OYU20VNfq6/hK/VdACOnJHh6B54+WJ/AcTTvHwohG4hxEqtEZ5SPCU7z3JF
K83t46tQ4+8V6AO1O3rX+y/9qCxW8gqvl9PhOk5+5AXhn77PuKTMgDHQVleyffas
3vZw37B3b9ZnEvyz3iqKoUkfmdQy1KAekqlF7PUCt2nqndnohaujEUljVOV8RV4W
9OBbK60PXeGysTsyUNEoe0T3x14w8tB/nWHaiygqBaA8D8KS2P6W40sw8QD8D1QG
mMDkVI+5Sca+Xx5TOTztY4Klhi3QsfaSFKDLgLRcF5Rnkk1A4szFxkLoWLTGPtxL
Opy58GaKEtY6+943tDVZnw8+pGK4jTJXsxNCGUKV3IF8sVb/vOeGHJuWQ99vbbHX
BC/qrAnzmsg4uG9HW20ki9Qnq58u+vNL6p2hcSUW5WjOendopVavT/n1CuPRbpn1
JqzJwHMMr55Pe0m3vzPQo3hzJt8l73PSNh8Z+faO3vC9gJToeGluYVgHeOypthMN
q1K6hdhot0j3wFB2oLrOzGcCwpFLABZEVUol6GrZtSZplu5Zx0Fc6i6x6tbb2vY9
Z21+PJZ+IKFs8OBPF64pOzjFvI+MOUKj7965H2COQu5Cz3eJuXpvv1v4xu9qid61
oMG0IzLOr+5gFW4rML/+GyiR65znSrYYZmOPWglB3p5dcjWldaVN5sf+PPi/s0Rg
r4KCJ5vnFwEqy2vamV63JMlJ6eAjPXzrXgRLBFdcF6twh2+ojai+QqJrBu0KK9wo
QRqPrNOkMhs6WIXfKrigJXOqvwQgYWsJuhZCEd3oIWF9djTWYuqX9XOuWa07httt
7WUjWL6uL99GfHjFOHtWY5ymcCdGQ48QhAhtSqFdsYEM/BjGHas+L0fZSOZb0EUb
B2D6QmOSGE2Vcid0wALG9mgRjHyjuq5kMv78GjnuKCMQRWmvsYrj646/9pN5tK7c
FmwieI737tMaCY5hGlMyFG1aVm4UfC2Kw2D7RlC5rLHYInhpqTXLtFIXRSjN1xFO
vfd/0qo5ehgyW0AJKuvEz8BlKpKYheN3+P3FOj00E07rcJbXCRUeMiHwTwaqpYAH
kzTdpgrNS3IRo7PTUaA2HjS1Hsfuedx6kvT2ybAJXOQHuqwZuM7vzsKEnPOSlWwB
xMaaXDPGKoc67lC/54OHnXqOSpouL5/l/WujydwzyxxCEF3P6OTUTrKrJapgYYfi
aMm4+dCs3WzK+0V0fMDuePEcdxDqQVWwdWIL9EPywoWV4kA77YGv0Mk8+2NgERxT
GPUCm8G6eh7x0esSn4ZHQH7CbfJYGn021CyUW42YBOhe3JlX48DWweDKOi2Dqvrq
coBjwsHRv88ErMODN6cnHzmkKvN5BwXKfuvMl3iY3RasiyeNrrt9l8we40KMGIfw
pKOPyu0BlrMPP11w4lVLWOLDxL1XbmcoxClC9weNMDkshmtK8PQL9oPylxeL9IWR
iXweoQYlJRwpz5VvOdgh4Va0rwyJEgS6oNrO3eUTCvw=
`protect END_PROTECTED
