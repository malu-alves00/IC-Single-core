`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qGScjVVjND6HRQTZz+qGyZgsEZPH1u33narDy/sTAjUYbbcJkGdkEj6jeDl851ZB
I4+f9fIvu4h6Rg9wXEYdc/1bFfcActhx8AZQaD0XvLhFn0JiuNW7+z9lxLmEIlxb
7UhXZ2cgCrAUOi16+uSEc6XcXCByROtf6/J8IRMPa9bKl84j+XRR0o5kch3oEl3p
SJmaWCtSofruuPIzcc2ZmQyXbwKXjDHHiqhphYCPYFCU0Dc5g/Yt7GKg/lrxuHyg
hobSjTf003CnHF6aqkCc2BlF3CIsxXwPnrkBmayT8jb+BYJWYCQSPPqWEigf1XSn
6v1YDMZUMTXnoogJeK7vEGJ9LYxZSqUQio1ZBZVeIzSPAjz5xVTpYadV7+7YWp1M
9or/NAJKhv+IbbCd7QvKTjiHDwRCMbUt6vGk+A5gqJBk7RySNkyTYo90d+HbG9is
eGiw7IqrL8RTTjuz7I1tEd+venlE1lFIuFWEYs0BzwhMstWRS2HEYhNSPoS3PJfw
HleVny/snXbQOl8iOct5SPvdKK2+lKByE3iDW9+LRrJupq7PFuiDM+lQZqV9sn5c
G+TGm331+K7F4wlDkRZBeqUPgyYFoJyVm6SaRd+lsqdFapcy3iMN6JXgU5l4qY/B
QSbsXleGK2pKYmG3TAeTH4BuOxyIaliC83+gLlnGbkFAOK1Me0Tg2/eHNpXo7K3H
XNbBcuum60F0kdvH/yie/pLRguJR0mj9yWrG+a8d2lBzsC8dL8CUhdRq0VV7rZls
6foJqFTFFInFzXVdRwlE3/YUJKn3c+8JjuMTe21psmo/1tqKw4/6QpjDxOuwyNaW
JcjWR01NbZ96wc8/Kovnm0gkxPNrPY+zOW41DdFxhmlDdlpc8SfnrvPPMFfkli3L
mX4QziLJCV6SyJtiUz/eF3zuM73pRw3MePHqWknGo7QHXuxnMwpcaZXIjOfVAg3P
/NfYjGhLFZxhiWcrNjgMfkMJF0iugSIanHQmVaHAhSZCMpBGfT/1UvFcVBt5D/iz
Gc6dL2l4q6VCn/QqM5fZrO6eGA+9SaWh3wVURLlUib+gVWl+JeaZj6hzVBVkCB2y
CBA245+ZmxuAeUeaug+CxmmJvDL1Q89k7vwOWFEPhKlUyWzI8X/gNYkd/0/kVj8l
sFaAzjS/UmgjCAiIE6AQXYdPe6fsqyUnha3GTuvu7gil9VqNEH0JuIxEefEgqPyr
LfxeOZQ7rZ49YOtD6jk93YnrN3IbgBr5XDIk+kZbTFBXQz0ywZ5xe6xnnyCA1iHK
erbvjQjO3yQl5rYIUro1kuq9lGPztAf+IcNtAzw/HpOHLQcBPbG0hAafTIn69cYp
GrbFZTTPb8XreDyfDRHi+PNuoEmXlpkW2VIn8q6C2lsbYT6jw4NtHPUOS8K7+cau
GdB4BEwm7WH4X53N3JgGnK093Kz7svOB2LnH2SuUaL7L1qclxXNizWVJZO2sIE/R
GnKcxmw3kJzePRgpvFIJcryIVFP0gCCZwUShd1MIQJt31dsEyVXPPnDYFYjWKmHS
31hi9RcwYQ4hGiUjRphXn2TWJJ2aAfQWyte4vNQGL/tPolQAZyojW/LELmwHT7J6
gbMZfQogBwQ9h64H/D/dghxLcbJeOvNbs4AKS+XkptVj1zvsceq40y2c5Sby+F3a
sIyQAPqBLtDAhv9otTzsilVmn9sUmzy6w4BfZToT/xyxlD+3Xb5SdjrxXakJQByL
`protect END_PROTECTED
