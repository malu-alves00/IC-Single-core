`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0ifKwOMOR/Wcvn4StCJCL+tv2O2ZKxaGeEIMwuLDSNagmChLzYD84VGcRUI6skGa
uV6v/lv9gk0SUGb5qktRODbXrDJ+7y2zFfGA5K8lsaj8nIFU3f0e1J2RA6YpkmG0
qP3S5QljNfyRa2y/LEq7AlZvz3D+0EmXo1gote0gReLE3N1EWHc+QZzpP3sTgB76
NUHp4UAVFR5HnWC/6ZWN2XAt+elxN1Z9F15uj0UyNx7GoJLr1foXTS8KgGdT2xRM
xXLu9NVMgI8tmYA9ujk8TxgQm3xuxcnCmJokoRZxCC+sCKy38nYOu7Hv1FGvO8/H
sbrUXRS7+xmbwRmcMgcQKzX+LveMnH+yOb6xnoErU5jI9L4iFaA0EaC9u4ecfn4N
`protect END_PROTECTED
