`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EHH49GAsSZ5x5zJj0I2JzamrxkCIMNCJxWQ8j9O+5GqrJLddc+qmGkDa1TCZ3HyS
PkPpvOogK1Za0PegCJOpPm6wltBqZWFGr1tNCRWRE4JnQRasZtqsF1zgLYCD30+1
WVw6V8jzwTlR069xIsFbrysGYuMwJz/BTckbxNp6V0C7gvDNuqkApzW0921idue4
+EP3kESttCyxYRtaRYRtta2STPe1o94FK3aQKezMgCfMvf5b2Z55B280YFqVtsZK
FcCa20LCaJfmD3iF+VTBINuAtDWle7GVh7zFpgEptX7TMi0JO94Rwyz05Vc1NK/I
6/GhqISUp538IgdozSGWHA2aapWP3pydzPErhOS09irxdgG998c0bEUMZ107H2ag
Q4TTw8xhh1rczIcTmFnY567ht7DX4FylddPHFiMzvSeJPO1dnrN9NijFfW8iJD26
bLPJIkysMl6FBTUlf+L2hA9A63DLtONZeEheDcotL/aWmr0yiZMdQmQEpwCw4q6A
`protect END_PROTECTED
