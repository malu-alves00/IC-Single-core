`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RxsNFZ93lPdekzGWyO91FNHEWJ5OqJwPh2ENUj0JxPeIUs22rufa/zqdxylNHwsx
lfTXhsnjDoHqa3kp5+4nITVnu6rkPtH0hGIKgyuDCMsdsSH+3roZxqNsP4uHtMr8
19MpLO0MVRRH5gpPDgtgwGmqSI7FqMB9L33tjUEzwFG6UwsGwtAaNGkny8Q9OJYg
yVedNN/GQCwtBCOZoHprZ2R0BAqSUyqR9DIof4vdDBNuMJmrs96xDeHV8sRH6p+e
K3FHQZ8cRUEsolkESddkh/nVM731vWt26nuxk2t4i09uI4zWyajJ6VaYYR0P03iw
0SEmMGocuuAMrzTtMrtNsO5wIw4RARCpyGxnoHauOpjR4JLAIZkc8Mb8vz2b1Brf
IbFD+p4lFx0nBpGbpRLUEOruwDoEQVjwPwArYLCZ04QZgicIKIU6Uf1c0JlvqARX
7VpaCLznki+jvSKQqBg2tHBnx8qy39xVM0Eq+T8LMjbBN2Tc3Dz3Wj/Kdd+YZHyi
eArzZ1ndNtADH12Co0haOqYK3fQJpij3dofoo87v58BLFugB80kxXj2OVx28wOuA
0Nx2uZKjSc3Ej+m46IPhX++qs74XofWdzoGZAa9LmcAMvu74CM4l+25ZMH3U1eXM
YS5QSRFdLWiDqNNAW1eQhDdcevhIhs8ezbUcO6yEK2tR9q+yLTPyOtDDs1n3TLGP
6iARyM8PSNuvQY+SA/ubvh9E59sQPuU3RXaFR6mXAX+A//n6Na+qjsG1BdM7myv9
bhf8te7HTTWMqMi0XdY0GsFKuDiMWaGbj61XSnS4+Rdh+m0Nly6gJD3NPge4yEF0
InBqM5cWxB+sEZNYwRwOUxhwswvX0/mj1XVllS+76QrT7TTOmMmHinhAmpaGeOt7
XfA/uAC7iJ+nuVoVcE3Px7bJg0ahHj+KTaCrCw8Bej1xjWPrPVyGFS5H1j2gZa5t
IcgJwXk7ob1MZSqDxkSlpKDEj9hyeb4lpbTWb4EyxMxuZ7kwI8fo9Ry14AoHvXhI
gYlJIw/MwHwtdmzDBJxH6iUywgdFDl5KCV+1TiWMwYqHAY8/iRzd39cSQYxHY2N5
43rClXMaRbTeciMoBc3aopkVL/Kup5LeX2SOTT1KS7cZlHMGtSBlnav73265JxQg
i7dEfpBZm1wYo+4L+zTeSZB/8gYT0ePc3XRPBBlGeI6p1X1XV1+Cx0RcE0wGO+am
qw6ukIzzlqnWbgQWkMM8Z3zE7jderk1TyTXbzu7YBJdxXT1h5LU22R5cXSvZx6UL
tpZW4a3sGoeJnTbQ2IftwGV7vIbdlNLkTTjEGMdUtqNFcefpBz/+9/YW9EZFNEgn
GClJs9a/Phw9PiHjT1DI3Q==
`protect END_PROTECTED
