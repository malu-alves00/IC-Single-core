`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3nHJrSHLCmFJylSKAu2COqRpKN6aevF6H98kE5o3c2x/kZvOD3t6YCpC3Fq2x/Qq
1Ogz7+pD/RAwkvdU2Ly+sbUZSTogBvcL8HjBt8ZFx30Ifk9tr2tlsXxnWiDaojwz
z7Lhgwn/Qh5vlzwk9uSl+75kwIQOc6OLJKUWeNWq66CxcFIaTt7cxpoFvSgaQYdC
QNaudMYLC6DrhBwZB+PaTvOZEJPt4s1JlY9q3reE9KT1PshK7wT76MjIBm0pacn+
M4uZxZ5kD2LlQCPBqgboGj618HP/iOsM4iLL/4DauK0kBFv+WjYkMhGKfk9aVDVO
+SJn1InKMfwxSIWQ08HVFQ6QdEUrqhoWR8X5XVNZzZAtzdRqEU0oqDMGHHMcRoJo
JSSD2CYDuXuh1rdRAVhedMcicJvZW26+tqxqD21UJDD0+P9HUdpwAe0lrBoATI09
ogxCp1+kxX6wwwutqRrkA8YEtDCDKoUiIXvQEcvM6wKvm7QtV4ZdfP0W/6vnr94F
odLHWQD6Zv8lQi9uk1kTz18lVZGWTqhiIGGJ26wNnwnEN7xGADnKtLHA4SjuvXFa
wV2fADf1S9JoacTueVX3Y6HxuDQA5Ov/63jxZGm4dN4KEv9NraNrqCl0CcCKbSH6
tiD0h9c/tztLuwzHaFMEM7I7uJAMQbsDPL+cGHNObz1cHsn90ENGRz/hu9Z9FLzL
o4LuvJ///AipZ+OCWwv0nKsCL1bXVbjLbIoeUzyW9UV386b9P8bOvntbTe4p2Vgw
9gD0uTYSoZI7oh85E5eAC+ox5LlSxkZ5is1vKfqOa6KTGcG8Q1hN1yyxV2nyPj6I
neKsMFQ24XNLWa7gc49EKLkuVqlgSJeXuSNIffa5TQ/qH7bmBvZZtQv19qDN9xoG
MjAa7Fz+H9ZJAYWSTB5v2fZOzNBsqwg1I8C4FbC+/kfFh260dnDOjffGDwedPrxG
0PyeEG4St2CvjdiRvFKcCx+qzUaxfwnbvSJdOQBKJZQ=
`protect END_PROTECTED
