`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Owj30q3vUY2AtY/zmm8l7hlR4Y6jA4m2ugVNIC1SwJW7qOK/y0wtxgQKNqXWdqB7
I5JH3WWePw1CyBH9G6pP3AEWlw0lONVl8Zg0+rscmfBa2c7p2U5uIw0QLWINL9fP
GnZR+FGqhpZU1tJWJ91tMXMOI9+GHfBgl8mT4Y7RBFJB7c3/Tc1LMktZQWVIROoH
/PODvU/EgY8yZ2YMp7x9PWS6xpUjhyrvKBP9TM5X1oBYJCfA4LbjD6qfQWaDCwQg
Mp0DYF8F1ShD/EAvKZgx6ieWS6/6t2NCWPYL+lkGcICC6PfhAb1DTk8p7ocpYi+g
WNVOz0OYVmx5WPT2c1VgRP5dr1TD2g+roPVmNhcka74Ci+A5MyV4Wn2TAjn793TU
07XH8TxjQKBLlBX9xrCqIyQVH6nbVqpu02TlM/BHvLTUL41v0t9q2X1nyiqoi1Dd
466JreOYIMPlee3+Esg6ORDudunpNGZeGRNw76/OsVRddEUXvJtrbXMrAcwhDppu
UyOK4Fmy0wz5ToHxJZy4PG6iuwIlaGhA8BRDCSB0MF+aPyDBuy5jybiXhm854ie9
0fi8s8hKyHJVrCMO5MZr/cmHd5dEXmxcP5k/cJVKw0AzoxPJ3mNLML2td/fK+wcV
oAZ5QjB+uRRUDFAZt/B46zO4Rt8bVV/Xjw6pwQTM4xRMkJE5PD5BUzcMw97v/GSz
sxr9CK8QdiJUhivQQb4a0vwIX+Uakl2cWGbEnHEPFSr5Aqa4x71ze/LrRXU47NAB
rfuQG0ofyBe7bbUiYCjP/ZJmpHRgnP8x2IcA8nKIbp5/4aHVHcQFc+cjK0hezW7l
1P7KVB8fI5d6zpK0Foc2HZaH8A9SxXmj0dUWv7uTppcT5UoooKzLauCNMcEwgIvs
mXJI/K0VeJlvWS8OLUjaGwgJAMYLZ8imiwh/yDzeDHQ88+wizMGRo2PwURANZzMm
IaMzKGHLTEJfG/Bfr+NZSw==
`protect END_PROTECTED
