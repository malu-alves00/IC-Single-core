`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KtGbIqKvrUvzvK8JMjdu9VebWk+SNVbUnvb5JffUyqnfcPVQQKuZsJu4NCJSsVh8
3y6AVZjU44vVH8+0sJXUndLHhoKhA2ktkwIouVDAN2lp23u6Dvyu83Xi9xwV2zyJ
NJjuGE41RQ6CInsJYFPENlr5Z9MeBB5WdNnRDs0KjdH4BbwT7kk2U6Lh26S/vhNW
ZWKtkTY8BsWzYSyOjq5rhob2RfnO+iIY4njvRuJeJSXHWGEVOSqPjFAbUmUkFXQr
v4L1wSrq93wDM8/9vVYMJOmnnJH105zUP1JbeBBDg8tbybaQikMjC5FMXvv9QeSx
kEDiExqrryY4XAVEGECQ7LzLpDTBidGxP7YIcy3yoBsykQq4UGMWDZPEdknX/fBp
n99oHnLR2uOraMII1xKkFXgq7KIIJGNfBDGmi5sZ86FBqF0BWoU141fAIipHBJc6
01ybZKm4VuSRcNRGus8mQXZHDCtOmsezXv14agfPxli+maQoFNv/SaOslO9uwrJa
wPYZUG5LvH3pgeS3OOYShWalUM8NHWQTKq2Cc62kklHY4iqLXv3eaB4vTR3SqG6y
250uFnpqSXGIJoKlfdgGfcu+Mp6bdVuB9/63FykiBttZ/MClXOOEfoBJlgwMc9Py
8ASLKkLIFJxIIeCEwb2piXeowbU06GZ24tEdUZ11BgUzWsoJHN3SCwDOvJRpFFqG
p5LNPGgxYx9TakGfeXg7t5a7M5ZaaXhopjezjbcJ6/6KzHSBOjwMw60Ef+8/ClJC
YtCH7OV5sMgMfWehg+lVjef6vKz64zBrlGArSC/qBppeHxuVWWPUtHLtCyvrkMH0
rtvih0bhZ8HwpsYogVf7fBVmzcsmYyRBA4VJZBDX0prfujjdkJrt68U+B0vaLNDc
+cao0APyr0fwEx6HgsgHiSh45Umqmu/x3fd5hzyTmP4l82RcY1GWVDHdZVBnqSh4
eLTchoQIgkSe7K28CvliE05N44zb9ZuTPr4VSeLtvsOHmNx7XWg0uX39MK/DCw+L
4SwyX9ke5g5YFqUhun5HmpNVfx6RaQIV8ThvVQ5l9g9Rz6d++g9ewb2E5MWUzeM6
2hK9DW0NVnyi59A5GdsnXPlERFe1nnn0O5X5m9W3+MGCSLXStozMWYgnnVJ8oyU6
Y3/yrqHGfcjrLmoQPqSNTPT7E0OiDJ3OzJrrvoAY/7qLM24k03+o1NnARFiPmT47
QxiPJYZE+QmLkfHqiV9+OyGjkvSwCwDqO8+2rFfu9iEkFW0xtyOcsLAgz4w7gvcr
BZcNI3ikrqoLK+ghS8ICflP786m3Ah3kbaqlZ7YXLGdOKu+inJ1fBvtyUVYHQ/FH
LmYHlumGoPyncRU0L1WLg4KGaC4D2XDJd59Y1kf13nDJPteZrAqcf/22J2zT+zDK
Fbd+rEjyaHxDftrGFs/akBBPSrOQX84badlDzkKdTgYWxxl/vMOfHZe9X5RXpmCD
LtkmjyxudkhnHC1bu++XH0jbvwoHfOzeUE1Q/bPgJALKgcs+F+CLoeeMESC3uxPJ
wbrcOf945DXDku9x/5QAcP64ZZ4U7NxRY7PHBzuqPV6MrMaArpI2Qm0soVq9D4Xq
AfPqk0yn5WYJs3yQ5AiXD0GpSNe6lewKSYpBcKiG3GoHjJa74+vSQ+s4lSs7tNfC
5mnlwWWpW3GiCowr543U6WGy4N9nAe2mmU8VLCOI/uaSFln72p1cv+acZHSHLHwX
7tbe+WxPQSbe8kKu4T2Kt7F9pB6yQDp4pWZGj1QbpDfmyj3PGO7Ttk02MMILYZtz
M/gfsAQJ6OBWwUqOu3SVPTx5YBCGUhePCPiafz19ELHMJc2IDZLVjzsu+Fp2ERDK
9b50LIYDq+p/WOanB2nQr2Hl+m6RxSz9YgEHIRkk4rlzPGch7x1o+mZJUIue0Ilz
qn4nz5KROPI77/sZi9DBHORsnGqTGpCUq0Ckg0s+k1wqIHg2tVXOanEcCzyBqize
yzI85UkhjnexaSTehxyxTFUrcmzTsVWzsIm5h0y41GEEME2dc7ePzwAzrHCBSZvD
PsKsSNXRvVqeB+dGSw2aw1OTeW8z07xknITiNUmDlDbkFZtbCN7VKZMHQ8FKxNhp
emYp6BAEdj7cm214e0LKChUbV1GD6XKQ0KJW2JHu1OkdW9XwxWv8yejTOKOnBC8I
uIFi7vaZHiy9kSlA3tQMCUpx1BhRZS5ZVUUaBU70CN25MUVMXL3sLeLVsTf/su5q
7K1edbsQTGpvQKkylmkzCW62DIxCRreRztQnfMJAThYjhE578mLQhVAT7CQzmXAg
EFDZ0t8MZipse6rj38K0JH3vUuJykDwMPsqOpaZPrjXjcoHXJtxFwP6/X61t0fn8
QzmqwPj5M2genQ5EF4MhcXFt6jfLuFNfJkTGhqfilMbGzq9Yw/313HIsCdoqLYrY
nCgroCdqwh3zSG+XZBNqnzA4yhUAEvQJv1jYOdft6YmKJW3Vl2NK6j/ajr7ffulo
xer7iy4/NQ/3bVSC0hkgHn/jibJh1B4qKtHWzs1Mkk1YJpvk9NvX0Qtio9RtozGH
Y3JGM1jPmfOdhS6xiO0KTOLH2yb6HM0STWYVmVfk0LkBV/HQCSnMLHAnOkk/9fE4
q6rgtEpBTgCwXsyMH3qFJK58ccNHDGIMKH5TLgsyuUY5q6nv8oHg1p/Goq6Xb0FF
443lJEUH7OyREfssZvL1Nh0TUEK9bXTfe2pHX5PGxGoQC5gaWsF7mbMR8ZOy9c+X
QRiyuEpL7zYYIA0X2lJQ6Y2VGEO6gLAJf/iVHuuSlkqinuwP6Z5Sw8vMELdF9+Dk
mq8PMJ6pdESleXLNSUfzuscVi+HzFOuFQrLNJWIa9M9L8vgYj4oxa4Om8K7smAAQ
jdnjpsCmsCpITIGGucCMYUyzFafEMfRiah8GtLmkvsIKyeckTX3O1d7BNI4RdqPJ
EESS0UvkgmRHwN5y8Un6l0BgBDjtuta+z459fx/5XxdZXfuUD4+GXeQRoNY9XkYl
BZqSiFUhMXoyKZszlesQigF4kMNSxmqrKMjp/1S95B8GNEkAg/52hj/yDgy9oBO9
ol8Oa5Qp/Y7MqjemI2W8yt57v4M63H0izhYRJubB2rHwjqdKiYpRQ0saUMIFbIMA
bpTIpXHgegllkBJxD5o3RE1PislF+393nTxPFSAu0WYVXd7+datZb7148RidAfhf
peZh5vvKb0ADWra/E0gzfW5KyrLkcwdieF/i211OF/SWqVX070aH0ew3MLQKdRfe
/7GOIJAwlseCdL5hHWbcuv3I/oJb1IPbQbG8PZNr4hM/ezZqY8AtdFhnsJV84XLs
yqIiutsZLI9NG9cQEeDEfMDkbuOynXKRZ47cT8p43+/StX/T43FlHF5En/2g7i9J
n9bDqacFyxpDrzMdQZ9D8i3Kj1lugQsGY6fdDSWsyQhYagjloigwRQbnuC9txjpl
V/temzGBHuvngU71jUEn9q+WmC7fmMFSfhRUJhrsXa50fA79vx3/4Zr4qhzBtZ9x
w/GNMwRhPzxpud3IXSFnfu1CQM0HlL4wbOgIzlzLvECR2cOowS9EAMsop2qaYM4j
GhM1+jyDa85rK8sk2rperxhGBZUTr2qFCQ52/9ekgdEgSzHSQyUU8suxTmbtKkb2
Fh9KaKbB9vOTYI80xh2A6C70v0nKxFHw1A+3A8y3KiGDqV2slWZPu1op3bnbwwog
EEbJglGdnNswyAvz5mZKyfHkbI022I1zf7Ljf6uM02xDBY4PSoxSnB2y4mfhXnnv
zwKsumhVkiLGllbOlRHwGGkZ1SoFV1TBQAR8nWfo0tfcgZ69jtxrTw1KEy3+wlle
XEb9+GAdcGNYI0XicpHVPF8Wq2ISQR4OGW1ld5EgxPGwi9i3z3PM34q+ljyGhjmF
uySqt8a691eWh/spMioVTbfbafX5C4HJNaElJe8fKtPw22eoCufFWAAdfxBBzRcM
0i2bgme2NVUVN4QHy3uP0p3QKzeUaEi/cMa9YkjC8wl64dRxceJAtbaettX3/gXM
SJhGSqtbRwSniTHe0Y7n1WHYq4F/HT9lA3Tv+mlsgdB4RO6ayMtR9FoMlgecR31G
+dmzbvEQqoExB4Hl/kE7xWFFJwXdoTOJTEdAB1XbG78jUjjuRlFv1TNgawMebiOH
E+FAcnMNK3ohmoa4sbFDpz+c2FlMDvowFVVK/w03err0TAI7WUlM4K81+maG5c0d
m9ergIdwrNn7O6J2QInd0PksYuecs+01FQcwS0X7iyVNogSujD9g0ttI3Y2zYonD
GZ/INY2R5tfBk2b5aa7lqUZohiTCiZ4oPfwyczEoCrri/RxtzBRjuCec6z0yacNL
29h2mGpWwSkSRfCA/X8XkmtNJETgv7lHjMf4EgWspkDsMnGt9WgzaGzIQaNocCLc
/FxHZMwuBhTQdWjrrD5BznToa2wSyQxRtlkIzjfDZ9VnP37FXgEgDXI7jcEx3S87
nMzTV0KcW9bk3yVxBnW1a++lEs2+hqUgnUnkDLbwicJbTBO1Wwsm71IdMDXpiHyn
VX/xCajBlcx92tqcl0KomebbnfywPDk5fBDLUsTrsT0ZAa8Owc4re49qcfyObZ4T
+yCR4zTxKqJ2OcaWFJ3awzbYoIacTxv+eC19bmxtoZTms09FDjy1xViPNxpeoLTa
yWQDOOgjGY60U4fHe2qE3sDn0EF04W3x+bmo3T+HLWRxF4M0heA4H2tO8iAEew3P
QWNS1Ljrcy+MaONpyTRG0s1Qwhh5jdJ+6WXgboGXlnc5fLxfNtmDA8loNfscnKv5
FnOxqV7sv3PTrAnpaogZVBMC/7yZakuxbZ2fiUKWzJ1XOOknm1EaNz0pHwIwV1mQ
kxjN96l5zYdoqo1AUTogMI+GgSCejA6ipMjW+rEVZP8m6JYEtJOw+PZaGnYZ2WpB
adxYBb5utfvOh3g+qo3jhSEkMRIRyaYn44ZxUeEtlV2esEhkAjY/OX7FvmDPqVPK
zIOIQqAyXkH2XGBhMMqfI0dteJvQaoHxI1XYqz5l2gr1gPt7+GaoRYVpwBRPq1re
Fy9lnn5t5iiE1/JvQ3v1EL7xHv68FbOaiLBP9xDbg2YWO5d5tlcFyk81LfIiObM5
jFCag+6gwULfsL508TQZwcacToF7SAFtd0hm0MCRjPjK4I4t0oBBCl37R9/CBiDR
Jhs1Uqn1IKkkoTq8LkNJ0tnUNlfeGqHCTvasIrCnt62/cSxY3u5d7usOLjyp+1oL
mVZjlXvyn0aSV71HtXyumDqo2EijVRWoShOLRGkp0G1IS0ll+NbEK2bvpQdFOplm
y1epb5hJF8Q2/dMQ4NyaE4hr5JqWm6Y5gPxybcO/rd6ZQ4rV6NLkUsgorg1dld6G
xncURW3W5fM6DbWz0b5De4fH+5nHEWl3S7F21dc0uO+5R22ykQaHqb9RoOEgUEDU
DteIPm3ssvuBMFoiwZ1/vyoj5nQECGXLV7YgXs8HiHykLySuzIwxpIb/sKcNXsHS
InZEMWy4nVO7vOY9niuT1sdbWdxRlaStYoQG5aD6L8fPva6pzKy8aszGeBDMJ6J9
K8pbJV5u6FCG7x6WPwSx7hLUo0w16aw2TsVuxXv3kEkHmT4WucI3+abfr1qoZeaE
g6+5nBnGONPs3DfRqgBAkt9LZujXevlSeQ/niQH2vMui7O+E3sfU1g7na93GSVWU
Vc3Jpwzx45z2iKNQ0hVQ9S1eekeLM8ODAokBkPRX1ZFr/NBCb+URh6xL7gEHRu8v
pNgCEBjbZZ3lmGnBJl5UnWdhUl4fA/J1xriePOcBzn7HnvFL2bB12lUBgqXgPAZF
OzNYserKqme2EFeboDqT6E73cBeZZiuS2eOciU6432hoqM+6fU5jAtitULCvSYWI
6EJg4dkf6Ep+sR6yvUSn3LZQMZXiiJDCMX7J6npgdag8eKFhQ9iclDty2WHOu6fU
2+4C2hkM16fZoWTgHUC1H+PJfwU6KeUVgbvIvH1qqzsXOaewBShlFQHpP27//kid
HHNkUEe1E6FNp9p3oGjLYcyqD3ONwOQ1LVvCzRwhEz4rwhxX3EVxg2AxntCtGV2P
ONqTlgiGcT0hg4djGnRQkMXylDn4lgzd+/vpbenaZlxCiNRFZENrPuiRsXlfH33v
Ti3SdWyfsgiQK2OhoXr8Xndin3JdF6IYkh0Lzf4h622fJJ09hDS3i4BJInkjrJJT
R8XRwpj71Z74VmsoVm+wj4JS1xQSUA5FIijiA7lcCPbpxDk4X+VI9BtH2VcsZ4cn
xa15DlBtA1kYezbIVbi/FkZz0MWcxdqG5vTXFkA9g10uCUVEaMeXrwvFdG/imxy1
3zShAdSZwan6fJmQ4DowqfGbxQLqJd2QIPSiX/MA+fF94Eqb7p/lV+KhbWXLY8WN
tm8C+FXiqMf8NJr9eYq9dmmrwbH01r7zDi0UYbAJOPwQmoCTeOSijbFcHck/3VOi
a36EUa+yiWRs4UouXQTNxZLzGzJ61SsGUNqGmSjtqEaV8KCxuFmEWdvJ2BYNI9EA
hNd9+l9LJxvI1xc8GDeYq3TN8ticNeeFpkRTX3DpSiQbd3P3eFhuFXVxtYdvmZhg
gKLVvtUFcAwsrlBJ4G0HOJsfoVyj+TcSMInMWA+rLnkLqpck88VACiMtcQXzeuKh
Mn5SJwMgAqwsy9IpwXCyOUFU5qyOmXYkXrxqaEysy2nb2UW5U4lgtMo6NINKAFPB
U9Ltylx8NRVDb666HjnzThzwN4Wpz4RbbsDTKQvkjKIBz+alGF2S0eLm61Ws2HSe
Zfl8mgVHrR7/uROsx13mGHy3mAysQmdU69S10IZ1DaDrRr6vdEuUY4uTHzIv5t6/
4+HZrhzQbnbQ2pwTxAKNS3/EDkE4d9P9Dto6CB6/wnL8wECSAPyDCfogFQz15v0m
Kl/wHyES0+CAHEIsiZZWOuNbqPfaLdi8grMTH3DbP9+27P8H/VZvILkXaDVRy+RV
AnyuuTcotHoaCuAe7fcnA94acUZQawFtlKyt3AL6GXxzxttoFysuPb26ooyoDttI
566+aQdPd/ol0EmBC2CoIDXnIUnH6+Hx0LuWMpyCZVuPe7mYB2K3dHxTjbab/Ed1
pIIEZVTQIIsEu6s65pGXsKo3GhD6cCBY873XIVjp0zzYr4TjiXPWB3G3/gVa8Jxn
O2Dngsi1H82O5eQJ7lYpHvPMzECp+BPLpOO7a8relqGyI/azuakGHPICXAFeiSUC
DwI9jBGu7iOo7rInOlIWwMzrhlKDxb0ONXs9mcnI4xAh+c4TmdaPYcENdC3PYrJ7
c8EuaNriQ+ipOlWisT63DNJg+NE6j+ruqA710XPw6HlbEri58erfZDQUftnkswj2
utvOQiF9/BWFtx9KR1e04kb0iqoFGizs/GC6Nha7k7x4dpy+Z2rcRgUW7umU3u3O
4B2mAEmq1rfH/31fUTemzb+IYGH/HzN8jx0czhqwRNmaDpFD0PraV1lhMcn6BY1j
cEXFv14VgIjypbsz/My/vpAXq5gfjpQgHAb+diwrh8ACAfDf9Q2SheAt1UFSXt+m
y0iJSeBjoUgPg0AOIdzLZ0xGvr5ekazs5+0fKE4oh+nnN7xdPn9i7yPzLmjf7n4X
9y/NO8FkNPbpfxI/zv+caHHJLlLwDDSABjVNsBN5cwvMA5blMRfJmDuV9QYIxCo4
dmfCJmo/EwkDeW5pVhi5IUcIII2a22YLjwiVdBHSZ5renIfBjv5F9dRH2DtyLpY3
HIRyJdVGlUk9vXX/KGxE6BVG2XuGa0ANkvUG4QAd6nZVSGj2dTMj0xGORFDeoRbS
2FVmQuQVSs1cRI1Ue45VSSTvZzZ1iaLqHC6cP4IfqHsUQnz//UNCBFWgO6j6aUZ4
gfmUNPu37fO3zrJKFHqSl74hF2YLnWK90aanCfx/WGSRL2z6zpP+R32GpuSNtolC
e2PdBycgvAuneAaXq9QaammSvsTxjKTgzK2wX2LVDi8PTWYmPHyOCop17kW2D/+J
WU/tSM75wLtaZQXVMCKhwLJUSpSw4obwAgXAUIOk/4HTI8w2IB6sebU90pBXvs6/
ozhGrYwG+O+hXiA9dQjPuHpQXETJ+ZRE1Te8MyDTvezHOdymd8OdPTZ4gs6XMpYG
`protect END_PROTECTED
