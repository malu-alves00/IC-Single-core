`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VPaVJoYN4toNp8P0+khDHMkutEb1pE4GZknZ/pljeCOEQdQCPXaoBLZaPVByhsph
oV5sY+PIKN5j0YffSSP8XVEWTi1UAA4nnc8NienO+oNxgEZ72MipRSS1qvSmJrym
1qUnefe7tJGj4c6WGm7qbknxUvfcE4mbXcYedXjNOfXphjucamrjo9Pnpxkw6J7Z
dVylEWoPn6OrUTOSV8VZfF5EKF5QMwfpJoycORCz+Eq8eusYwLZ6ner7DVQpEShw
/ifBCBc7+05qTF7/P0a3qZhs9P8MSP4wYWRhsIWui2g4jaLjFJ5VfGJiBjIQKk/6
Wtq47ThULfNoDEvNpYi0t/0bLwLAgI1I/UWEsq5lo3VmypK/ga72J1Ni1+yqpulN
RcKxopzGvk0e2MvSvBknQb9j4pU+6wescs4P65zNmpHW1KS8EBFvfNcj/xVeA0YN
NCA/yXAsrGwel1VCHKZEedYsTZIORtyYanxEM6Dnk74yTE/EKfcgTuPjzRy72NDC
zkArFZE/B4Cfq9qG2uL25FkRj1YLsIi/EIVdlK4HPy6ctBd7kDSuQKmEF0px7SpZ
9GQ4vw2ITeEh6iWnYS4Pbkh8D653P1yd2UG1kY6xEL1wcyqJmdYXut4pozyD7UZ4
YgmrSGhdCkkxVLCOOva8/p2dqmYsQN5hqyOQz+mIr9zBSFyWdDnauzvAwl/cxww8
sMy5tZcwwnvwP08lRv9mFZa/jFS3TIsMj736VM+nQ+hn4nOf3NqqXv6arWP68JxJ
k/eQcfO/X4nLDciAig0l81EcqasHH8LfjD/SJ1L2PTvvYVxaSHcWKANxuliKeR9K
nppVEgfvQ0QOxvj2KW9WpEWKavejHNFIKlulNJZNfrEZIxoIGxQFaKLCutBRN7Qr
J5JcnVKNwJji6hVyq0FgCM7H/XKDtKHNXVTwRUwuV74tWrloJ9xVnG1z9JfqlRKs
Z4Fd3jd/ShjSk/iIqHNA5/Ur1u+zWBrZOWiVNjhwVhzdMHTZuLX98w/JHuckDzaQ
9kp1KbYfpBVPeodyt7V7lnDcVE0Ektwmm7N4V8htVEkoc+diyIxg76tXwpGhJHma
p/t0xfqN63qbNcQ0k7QnTqYvxjkK/Pe0OMWz4ioOZUA5jEjbhPomOtcHK74zhwb9
Ir/SZizcdXWm1Dy+Lrx5LPiIKhrclx+uoF9JUoYE0G5975Opp04jFSstAuiH52Ha
Ck2s/ohiXSrPPG5eGlfGMsh3Vrn9XOrAChK2su6+M3fMmtWfO4YgOSQF+M1ofLmH
7XcVyXSTd7DCufotbaDzIJg/sTl8lu8TEnnJBWITRV7JugfavwNke/LLR14yqRk+
PyAHZesY7Ipv8wtET9DZEZ/5I6Zc750r/+McLIGcOI/tnNMgN9L5lx/yHFqiCK+1
qFVrjfTeyBL1UPR2KNJhcpIjj+09tZ9nbs0Wa4jup1PiAbkbNC3WYcMG0PSAFU9m
bLlWXpRpVzjg+3x7d3D1OF4vALG4dwZr3p7zULAwVZ+95b5m4X0Zi0qpaj80HuPj
FrQvlnQRGbSmFFWfekel4LLXvESyg1nOPh41NfIEtZNkrMMM/8CQiD8JrkyyB1CE
y8Ab708iYQygoM+J40hMuE6m6+Cvt0x+6d6Bh7A7vCSIBSYQDx0xfCZxZfmL3imE
Iiuh6xlsoYmUn6PHgOqcFyfoDkaTCTDNHbMcy/DjnhkHyLgjzls/+yXSLwieu2/Q
NuE6SmRwhH46hah+V7SveBtutPgJUro/6oGJZetYQGcMZnEwrrTLgqvplfjLQqPl
3/rlrll8qr3/64TAeyUgYBdBru6PDOwp0krZe9Awv5hiFMBfSgnR5gNhZwftFnIr
XmBDoqfBGbRBrMZ4LKGsJfO+HHF9j2i+7MPnalA9m+bd4cUUH72zkigJYilQvw7U
QB+BG3nWESPo7mssk6hwfnwgHiCIR5K7xNoVvH+WXFX5Rq2Pc4BCXuONqp2x5dNb
YdWHJoQeYnd0R7EYGfUJi/QGc10/2gRpKiZO5sBB53Q=
`protect END_PROTECTED
