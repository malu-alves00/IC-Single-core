`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XnYibuquq6WQOfloZr9Z+NupIvvdcTtdbyhO5OBglh/ZKzYX2mTGTzKSHAXwDaCw
wA9aSN59G2oUJ8HvpPs3QqznyMRTnDhQcTIx/98KGiSxYa7AKGMYE9V+lgDU9zZK
/3fd3FHlLX9JpOPJsPN6LTQAIfD2t+dQSOhEbV/dxcSCK1DZEclnNV/Nx7r4K9RI
h+HFWS/K5KXopFA49VvMiXuvilbP46p0e6GU2vSDP7OvtVKt4VhQvs6bcYQEb6AL
4JZ8DsIXY0aEUUTZTvAiE9o6x/Cq6h/RiN0lSEQp1QWhldqMbcawfZqfA2USRtIq
pY/EO70xdIHrIwUfhX6u3/Kv1KcBrj6nHAF8jAFCO6fLi2jV5gycK/EFmQj1uDpD
s2JlVePSMToJg1g6m0rkKaCXLcwyY84bqMUsxrrmLh7Mxbn1Di+mpCeutbDBKRzx
VPfiDtzoG0s1gQaiC15Lyx6tT0qZoKoamgGM4guT62u4R8ow0Zj+244LqZ7neiYh
Nv49wEbcFSFzpN6Pzz1y+UwOewip5Z573A5ZWqS+qFtDMCNaBqLWp/1/RIuOau5l
jzOkMiywkM43CkXHesP8Xj9oQ/RkVeJUeQNtG/MoGnz55X8hRb3vEmupjMJvEnVm
5sMTEr3QcxHJ5iVRlh50pVz1n++RpxJiiyBP+p6/EX7ikQlVItpN+WIADGvvewjS
BAqcQtQMD0JYCuyOf0+/5l5D7SnlitvncnEuntIwu8tlubBowI753iaf87AOiSNq
WUz9XURi4WlfNY4XuUGmv1AXpvR49O/1DoGIGb7j0XwV72A7czcGdP8HCDcswrVL
PKYXOnbEJauSWIcUGiyOzFFM/MKPfUP+e3cBKFjFtJaEFi3rbzmjxVi7B8DMPSli
IKIA3DuwpkAQGNzMTEfgOL13Gb1HM7v2vuIsiFo5+ao=
`protect END_PROTECTED
