`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Rl5fpoJiGKBaiygfKnkSoRBybtIodBtabNAsqVBeVbbC6GPFe+CEmeTycaOhhJ34
slJoUxxaTNq0Iev1grEM1SFt5j4TVX6M6cUtaZwj1OrXIicQxh3xDcMtyYg/ZtRn
DaZPcKtZvvnP6GG4oWGhVxS+p0xYdvpbPKcM4UBqihjkL+EVz6L3RopPfJA/BOfg
wXIaSwMYjM4T3u4GOLmy34SahZGn2osin9pTGEKa6M5EqsLEC/eCZ+15hOieoV0j
DAKyx7wzuJ+Czqieuszc/LcpZGC6jZM5/TL2PbUE7Y0HkCf0Qf4nnMhD0zRFNXcr
sAqwTgkSkLYYVzvCKIdluaPVKYAyb5KWWIEAGntX8scsG80OrtUXEXAa5o4KEmea
3+KEnXhzD0mapqBoMAgfiWXcSe21TnhtdQ9nTNYbSzB3dQWhW3ZjkQUEq4KZNzX3
78XXzj0V7Fk5j+h+T+mtpE3Tbsr1hS+/02ljuw5eHjS/YxvVfM3olQN/dt+82DHs
H/Tgi+XLBFVXMDQuDXiAd3D9wm+hQ/RQUxntJcYwRsh3uEnP/cIiUhdpzR6CUnB2
xc1g83nyHxoRffA6bPQejK66Oa3M1839+KoTpC/rWl2KXgbqtESXITBC+fXM2yUe
oZ/4hIapDEJhotJlDczcQDMWY42GjYlasDfSuFX19zjDFubrm/pRRiorALfTSYT+
Gryjw1Q7hDCyDrqYdfSjUqxRKC9OivDc7xOiSQii+OxLN7s1SWLFoWB7T1pLgyrg
1Ae7HFmJnP5hq13GFuHRG0IXuq2N/SmWrAk+4Ex4YtVGY/h2UfNKcP9WcK7o3+Vt
ACFGDqUF6sHn3gbwU+LIzA==
`protect END_PROTECTED
