`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Rm4A+M13gsu34E1Xsq7sPuuAgpFTyFHR++5NgUW3keL1h5bh+q8d1jJdDK5f02MP
s9L/Jl3KV750c+Y8XHsTchQfAiwbW8nkObkrD7U3IZueGGzZPAdx7QEY5YqjxS3S
bRHyE+UY311L8lqWIM7cW3Q+2eiaAMmcFGru5WunYdcX3TGeRuYk0kBTueY3j0MQ
StAow985RZLcb902bj7/n60dXNFYaBNx/n6clnmW6dFDPhXXJoE/LhM9aeS2Ucf/
IXAmOr79eEXLwQA3OiG5PbJoO8nUhsX8sxiFNy9quCL7w5MOtXQ3vQZ+MkKa4+lg
dREO767+aDveSQB1F8ZHN7nDbcHMG1trNYKDeVuVmsfwSSGJaFHKb4EId6jbQZpO
ul+y4TwApVfmomKhxMRv1l5bGdVw9ZFhu/gQFsaCZFb8fs6eiEPXzkw2a1VvLbzl
OUy7K6afc7AIC7fHTiyX3neuscH2rFUuYyMru4asioHUKJNPDBBrTZlXPgN+37iw
rmaSSJ/dv1TzHD/OjcmTdiHZSGMSQV640VzciPgxr3RPWzUeIoPr2+q1mEJJ0TZe
zFuKGPgom46CUIzvbfXywYFAMrqZC2U3aicPt45knH9F5OnLTZsG7Rl1z0PvRqoO
ueP6s6gpnEeGb2OxlmEPB0YAyFHFvtNdTZAvR9aGEPVe25CGfgxhxC5jf1rPCnW5
7nxB6y3HsRmNe2hWNlKviZ8ztHn6TnnCL9/92zDCHePVtL7T/sAnjHFCTHl6NgVf
ONr2D9+xAZWue+691T/oU3PxD5sXvqcyHpYE/VU4Uxeec92EIRp+2NXnTa1nUiRh
ZZYX3khQ3sz7UZluJgDW0W+RdOYAPWu0Y175gBkn+/vHeQDVgLiDq1uCvmD3QYHw
MzL7Thu7CWoOu+l14KMA+YoW2o8+UTiLXrUb0Jx/gROQtlEXt9B5fuiybngzWxgY
+PcqkF0EQT8JOIguVHjfp2iRW4rdywqSOjX64rBtM+9fYtR1x5ddc0HvheYVl6wi
BEa2T+JBhHm+9S8P0lV/O+Z/wVanrNFEvylp2wBRnTJmm09erw5DAtU45+iXbYqK
JvI6R+ZkA5FHWflIzQjju8R7als15/2qY2Yy/Snj6hJM2GEqLO8cVYEsy2NR4Jbk
WRQjbsrnVSPmVrGkYSHRLsZqPavde68bB0E9qw2v0PoxszPCwMOj25I+cbxS6lOT
79RczSta3O9cBgIGTM2Wz8oksBClYhomkGMUZbihjDIjSt+GF80MhsJRX0v96DIc
2TgdLD3BbZdge1Zb2hUlzitBUVveHhetduFdkic0YgA9x3o+5G2mfd6S1e/cnzkA
zMyCsvVL8FhE9uv8wPLc/smRwm3XHwDzsSznYe/6hT4m889GgRq423q21pgKe7OV
PK4Zz4ue7ChbWeULJpxGYV4GLRXTG2iQZzbXv13TdiiNByT1c9vvTdhBhNqcY1Wk
IvRmqv2lf/p0EAIDY1A1QPDJjt3DY3QpFYWR+dUWll6zFfraLCMLNsbQtT27P6GX
2mUHgrfgOxAGQPe90SOm2WhucrH55jb+lmD2YJvHPkEBlEXWONMEq6hiXOflEK8i
vIb1hdetX1foLoELsbo70DoA5p+EBAKsmm3qR+awfo5z9Kn/WMtVC1Vo1vasPY17
nuVaw/zmm3l+inZ7zE8ZX4WtyKCLU1sFXNqOfNkxjMzXIIO520v+xaRE3MWrUHHo
WmQiyZWLOA2tevdf5fmFsuVZXDny8l+mDEgjwKciUeO/c/4B2Y1Cj48ty8bX9rSk
biRSfNLrXzc8OaPDpzlPb2stxCz91ovnOYxHgZE9ZXCXMwhZshMlynJ4oqXXetPs
Hu6hLvVmiGgsaTossXpKjT2xO7eQye56Q3arFI2TKtYNB8lLK6V3WZ6CMcGEPVYD
P4dMEL42rE0Z06yyPzCVmr3jJmKHUSJw142O47WDRXz+WliT0BGY1dVELDgLFkJK
i8OCg9Gdk+IYVhFUfTVVdzjGyPTMQoCLNwVw6gGkPk0tsl1m8wF2VyWiA6fv6lsF
I2tZFlmk+j5kF/DmyXyhowENaroRpz+GqjBKBDomVYFUrqtH7WOlcGbUYRgozgLH
aBW5e0V7olsA33hmXHG1qcVzFhIIiw/83NuPiypqpdI=
`protect END_PROTECTED
