`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
y79KMpatDuZk/DqRPEhTBZ9ANRWkYBSrdVJZ7+X4Vz1GR6JdHLG9mCf38ze+yNG5
dISRs64AzFJ0k7orqS2phO0PgRAqZNdFFTP30o5p6o8mB++gHKyLUNMPV0KLDnLC
zHlHD8rNsINAS1BsXnSLAYFbqDDlInrnp0tGbj5EKAUV3jPzUfUYkEahbh+nPKVo
yXvw2ApvoDVLHPlzK4AVFPQgI09DkRbnVZmU9yRJAgaPfPaAmg26TkZgXraXcTNX
2U5JFRgNiVFDgKQ9Pz4TQtutb5IuSgGnnS7hSesoL1tl0/HsMSFoGlX95nRir6+6
SQpH/BZnCurPPdh5xhvYMH8Z+Gr5md6GkWlmTRSMYLOP0J0wuoG/nvl8qVcOQ9uq
86nfF4I1yuTsgrQ1FA9jQGYTvHEZnglvxMEqcbUolIhvfK380dQrVfSDjtFgD2WD
4M3WH/nc9efdeRQyzG2wop7aaBkV7e9TzT45nxCETw4qhk3nVKsTK+eKwNFYxNhy
uCxepjH/PJWZWU8CedPeEcym/C8zQ+YuzGoPubmTP94Ry6rEYTKoh9zhtjfyOS3o
R641BbPghZnIE1Ox/H9CrCEXWL62QJd3cEbd/SafwbGizB6Rh3Z9SxU8udOZLlFL
x2FUVa9wvNJ/DyBuF6aY9g==
`protect END_PROTECTED
