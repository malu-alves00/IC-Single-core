`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ldHLMgdCWnYTTpALjvQnVNUnApXu7UxXAk1o49li8QosGZGJ81hkna/BEbmbhxqE
dVrjAFeMaiCiPArAKqY+wNY7kuas8vA+oj9XQYPN7sWdVOBpKCNRKNnLisGiLp2q
bS9ychcli02pG4TQ5aK17ozILeK3+u58b1lQ5A020SBIjvPjCAkVguJGhaeQmSjE
LC1kQfoUoSeJWjLXX7uOabseRe942hY2uLrUMBrnsVIrNvPCUgC06r0/8fBUBuIx
0FFap76n8+Srttxns18bZt6Aoo+k5+05Th4F37aq6bxhSUBKRIwXTpTBwLNLQuMr
8VvKI6I+NJEBfybHyCd9bIgETF3pPfWYr/N8ifHtpSl79kAoBCY0hdltjXFFKOk9
xVPiu4zcTxuMgUm5xErUFgL8ZoTCQ1TvtdSAgjhN1emH3jWdeyEeDGlMxWZCCb5k
4g8JIaTyh0d4k0lc63DXCu23yZjcF8iFco8SmvzeYDBTtzndlw8UZwOB937PRXIn
S3ajADOHBWdBsfXaxmfWgvDmdcpctNgRFN04DdrUfC4Xu7XvgBcgyNuZrOHkwGrW
3IZgMP3DS258Hldd8nP5gG/ga1UQcj8me2xrcaJpzElse51iQ5Cvx1Q5UZgofZHi
hOth5vLyV4jVlJAJYuFeWq0Lj7+xYF2gfeldhDoP1vpiSZpbEYGB+cxssNZqMbMh
Po4hg/MIian011W1fL3EmwcQcXjujFH1ms2ZPfJwu8XfCb5oaKC1lpZ8LzkXa17V
Z+BcVu5icn2knHapmSjgBeJPAlfG0qDVzp0Cn1LhOQ+dHCfVdL09Q5LCEPX5AngW
v+hvFFdnpmclp0Ekstf/kgZ23RyQUVwNTPf1IAdIUv3mYAY8tGHIa9R2fdXSjYAs
vmdwZzzlkDruqjWukIneQq1Ofe4v4lRVrw94Ptvmx0y3OC0QDyF6BJfDKmR7nH1Z
w5zd4REFo2pEXnXHRkkaCvtMV34CHgnIM9kEsplG3bGnBLYoXk83ih1u60VMfJVd
sBpf/T9Z8CYXmsKkB2xotU6C31ey7OnUYb4DLu13UXFFl3aQBZyXk6GVGCC3HGot
J7j17B79wNDmWsbpmZVXfQRnypXv/A1Ut0aHEiqaf3O20mOoZ32pU5EX+wsLN/ne
RTYX7EqykNew8Y6aR/280vpathQYh0IOpSrJKk3sioHEtjmLvGNkhl6KaG8596NA
7ZENppGZ3RkQfvVu9mB5zgGtz77SneD35CMCCn0xA9eslcx4mS6wdZTvB9VBrkPs
tAGlrrEIgt+0v6UPm+ay7zp4J3C6M4EV+bxp3FixRTptFxGf6CcwUGEYYTieRb6r
oLePFeK3+1bDb8T4EnSVj5Ky07m1zYiZsMU+xjh0BLj0gAj3petRDTcY/K98zlLT
BP3IteXILEtZPCElBsyKX19f1YVsxuFk7AQ9lrvI1icqXTUZIpRmJwRSnX+2chLO
trOPM2ZyoG/LlrTOd7ha0rpW+pHd+va7QmswzlBuL0kNrYkoqmG2aMIziYgVFj2O
8KyJ11x1iE1rzLeFzgVTSozn1iDPW4EHSI9bafrP2V531lY6JIetlmcpbLOlFpNy
a5DOCmqryUiX8sD0wDSuurk/v1Af0MJah+CNclnoYp1fqjs/yFKg6sjzOwyqq9J+
PkTwUIfrBrx/Y/1u5sKHD8xEL7f6lb9ett/FmUlW2DDXX5jFhyPxRQtxMbQaOUyu
j/P+Q3cmByW3kLKdmo9T3ewd2UsNoQ7xH2pfK82jFigWSwGhTv+zhonRuR6DgmRi
R+rEyT97I/88B8mSmJ+OL7EDAuA9xmIROONRe6DYhH3CkprVu5ul2rVpt2EIcM4x
SI3Yjfml+ayrm2sdTOYbzKTzOvwjd+cvbAulNE0YUjANyfnUHm/zMJyo93a6CmP1
xXxROs4VOWYCcy7W/dVvtNShCnEVsMxZxOpL/xWxq2GeH+J1qQmwKdkJnDh7c7Gm
FMwL5ItSOztWEcONMrK/jOToDLnmWz+Nh2OJIv3IZSXBGGj56rofyrbgz+ZVE2N7
Tf/n++pVEkr2iBY+y/dEXNpMHwHjEMJEYRRY6QnxinNZGPr6s6Lx27LaP0Gu+/Ku
2M8aA8abianKFvOAIWOYi03SVoGq35BYq4QCV0//IUcyK30eeicL7SPT8UQnwLZ8
BLPUEs11nZIwdZvGfwdULU1BkoHS+RxstxyqTkxwIl3sl7DvAnIe5q2BuviTZC/X
sE06Opx1lPQmWUXGKzklbjD+gN2A262NYMboBPQ06hU9+PVbEkGD410/XQMoDlLs
hrmeyMLfg8/96C0uTzqXUf4kJuVnWvkmql+8bYZ8sMgbdzkCfWULK5yM3GXse7JG
94ArhiH+8IhsHQSgOdZ+D9C+0xUaVBVAOMKfnLR52LJr/FdRs6YKekN7CU2Pk+RU
FpT43PUdnxLim33lHJ6jZUAYISOpqQpSLyH96vtkCA0nifYvqiCMof3zk3aIqoEI
KyS6df13Yh5VhECBN3Y6b3xzsU77l2K7ixCKjA2Ndqor+FYkY+tNM01brHhrZtGz
gkvusw5jEzkAYSp2TMhJX6H/EWE5jBXc260H/Ud6+8fmMe56xjLFjJGZl3BuqCqq
THq+6i4MtUmDcmBqjVJbM3Kv+L5bJoqIUtKkFzpzhs7CvjkNXZZTtcV3St/QxSKw
OfMT8uI4JpRY84vGkSrXKkJeHau+6yAeeLwgMK6llM1RUnJDamFkTztDAwXPh2jc
5PNhsdqq45MrQsT3F3r4KG7N3X8ixbBY8lZVk1PfHkjk+PSDgsKS+IbYl8tki+bT
6GQNXZb11J0hEyXNPoh6pFvwfEi6gBt9lXCRi4MrK+5AcrrpsV7unZlRbJx2ftFc
SjTjV6lfPi76Il+i3ZSzVhBeLuW9oE40nwL20oaJ83b+xq1HsVCjEsA/AgmEa/3y
SQQPCpXvd7fjqB6aPoctwhRgE/oz5ZSqqAZWkIa9pUqeC5VS11nsYwziwhP0lSEj
1GiiamqpXrFkNwTi7YlrHrU56/CkZj3KhMsDuycFgxU/03N82NSMGdjJzxevidDd
lrnr105Mjf5TO5oFDpLfgNhLujZowGdBXvlovccmH4N3Ljfad6f0YfU6tU4jw5AQ
aYtEObWsGn/MnCw41qI4LZeGldV3jshINeEHMVeG5dbIROCatSoyj+RZXo4hRX/0
x5z1CunWjFlAbElsAXwxhLeIojJ9st3yaD2c/gbIXj/Xo+hPGN6Phu66OnmYUl9P
vb0AwNt7Yeeoc6gvaYFtcnnXKXJKLAQgtMcnDcEkVEPqtOVCqyp7dC5+WNeD5Xps
4GCzAhSkSV2X/4zcsSlzQOmtNAv5TH4zcXdHM8l/m7tX74j6lNa44yMSPDQvU3eX
+Eb2TuhBmdRDr77rDMJN4gQ5aCXa/XMMrumCV2lVtHw+Xo4miDcsS7PDRBwZCBl4
u6Au97bR4wasLyB3r8NvxhkXxfIRXkkzZKVpCBdnl9i1GeQ8i6jLmR3IpzvXSCv1
xDPFBJWQD9Tdt8gU26tkXAo1cFIUExXLmMeplYG7qDrjlq6M85Zq2fkSZnM3TVJX
PkDPcL3FYHuac+BjtBAbW+NKapUtDP4anMD/awY4LyUOd5SGP6ume8S/Nn8d91fS
igLADRmqWByxpu7p5/gu9TlPhiAEdgkWA5iXWUoLHFvq7HqRQvPJuxIwL3Ckcp1M
B4fu5eRrOPY2IkZVnXt/tT9qy5ZYzC9jwJ4ENf2WzM5FhAfdXYbZ3+sHxvXSgdDw
lPZVfwaYkZISyg2psnBFFN4bXx4MPYv7PiPYQftCXRaJQ0ZzaAUlLsvmU0KRo3xO
xUB8uEOgVv1UwMmvbyZnlyW5oEFFMYHUqY2fXQBOhhy/EMXFnFDAfa7jjPCXQHc8
a20P1LCPHGetYEq4rX/0RahCt0vK+19MbVRJhBdiJGfDCS6gJ6b0wUNm0GYZj7y5
pXispEvSfVrKUfcCPfsmM2NYA+p1UJnVhe98y/6zzTTG6D8D1kJ0puJ6/wKWLo6e
e8KED99YJWgYZ4lDXUVxVPDmipJeHqS6U//zDc30cHcHM1+FWz2achg2L1pFyHwu
0E+Gncd8vYCfUuxESl73VnJ2HsRrSLphwjK0U+RVS7u2OUaBe62EUsCdljR9saQD
7yU6YfHmQ0zswIWEHcSs0X+0ohUGKk66r7lSIa5WAYy7WLVdApYPLu1uK2DDpuvr
5Q6CqpveJEq2TJWNRVeJp4tzA3qUv9X75BYVS4a1MAu6n2TWY12HHtL2iWvfzSMh
GAe93A3/o0R8V8jXfpROK1Lnimew46h3Y76U9APPAnNMdJ9g8Xxpjg/p/M8WpQlb
rs9XSpsDB138f0iAMKogQoShJl96GRpdpzEnVGYosS4dAsQm1EKqrqX4qe4meS+S
WsrRUsmTLvOJVBuI0gRw9U/QG+wg3J0iSrGDYzL5A8VqycJlkcz/lw5RjQrE5J5U
BoiBRqRBt/AHA/LPcjt194h0qkNhmupMqZJZwp2+8Za34X4rPe1QqkqjXhZoBWyg
YDwSxdbMHhfBzrsLpr4if+QHH17wKYPm1ByWnQ2bR3WX3YdFynAjBHj0H9QfyEwO
eGVc+/qVFpZj+ZvOrB6UcnTIhCdbvM1Vn9By9lkpR2Tm5qluBCAyhcNIyS2xNNTB
jqHtOYxNjGq2LLYFb0ei15bn7+bI8t0eLiFdukQfQ+20BLgroC14760NlSfbKFBC
y+ekP18NRk0gfYLSd6m/YoaQ1QYtmhLbr8yYF1rz/+I7Yz1zM4xUzuc36mjBpard
37ONDUA5ofrllfDhJ3sXLLKHtNh4SFL2cWO6uGNezMFUG1uL01Yn9hxp74B4AqWI
rx60GtHyoxPmNloGok3JLzE46nyGzIYOTlaLah8M6OXsxDSKsPWehTBmsAoxx950
g00tyCUcFgP6B8DKWjV6D1klIMoF4hKXo7rrEGmjT09AJk4r7Jt+YEltEYFc+XLU
/7fGzKQ2ij2clhoTG7c3pqOBS3RmBjkLBTHC1SyCluTNpjQbTQ58MTqpeskBtRvF
`protect END_PROTECTED
