`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mCaSuDoZ/YQNqM02N//fOJnFn64nJUh6MU1rJT2HbTgGaCT1Vd3n45TW40mazSu4
kA5hWUpQNYdY10q41+JuMndCIToTkhZmEoNyte2PHTLHfM1q9dYaiSZcJqlMoL0c
CypknsuOpT2wSXIYSvOaZTOUmvYS+f3V3mCZ0gitnpo9jor8jIk212hkjmfF/wI6
JBKExDWta7pG1STq1BiKUDPgJ9bx0W7lrYHhIv18TtrlhMOwbMT1kCp+WqcGKD8/
9b4lcIuKD09tW7tC10kLvqQKPKgKDi/5X5FvQoonznFXO+VWWGGUwf2BfxiEODkT
aZNyJ5lt3xsYkrXGEKl7ZDfFU9WWiuUTu60u940+F19GItLstTA7wQGYJlVT/QXW
MiKJw2S6MM5iTe1OMWgAyCSP+mTxa1HamEzF6RVIE5f05ozUVywIQgG82vvbHC/b
+wAN2BXafFNFYD7YEzAXOiepSGAAFENlVMPl3MazJqexLekdzMmIE53d2bOsbxYa
hN+aFdrRxdYTKA2xSSMd+Aa+W35fzJsjvc14P9Avh7oo7Q2/YA3zg8KBp422EGPf
RiaYs7uKn0BHV+nnidzy0ruPJODsnVFFmwdaS364S/UsVgOsqpueuwT57q5k9lYh
o8ThPvqTMaS/FkdWJ7TX/n5UKSyHYZcwgeiDM4aOqRUe985ZmbSsMUyop2mfIDaY
E+aF6s6fZYhDw5BCGMxOiIes45uKf4uN6nSHnk1dQ4l37EttbiGTfXDXl5qiTURK
U3G9u338Aj3rraJS50ylZy+kT5A7IfI19MIXr6dV9GNXsVH39VAlqMN+QcxacYvQ
x/wD6tI4B7xWoTCUVwVnvmCXjGTheeItjx8NV9wZMLywXs/znikUni6kJZGrlVld
35JoVkSe+3U0CkTqRadXbORVEktkAlDuRPGtUDHNE3DFeoQTSypTMgen31a0F30q
gAFX8PUTWmvEwoZp1D8cyyn1pWYUCd2cnqkLuX6sMNgxhi6xykrK7DWI2dj0IAQN
8BTtGPZovoeJ0cFkCvtaxD5QSR1eBC3g+Jln7/k1ZcoCMtULwRUIrU8xWkWlm0Mb
NVlQ2x5+Uxof8l9BC23lZ3fyclLe09Gm70dCL518HVSekYNoZJh5CrN0rQFxyv3v
StDTGmSsOciMVtnWbz3VQTuasXEBhtDjLPibFlGDbAjPOkq2FDqntNf/vyLQJh5o
csreQ0U1Izyx/cOxYIFT88RR7sDYOs/QQrJM4uR/K9cnaIh7XE31swfZllmoyL28
ZAibJF8DfwFe8ADRkpAuurKIVY1W6fdUuDjNGuhOhYf5JSza0HoVsv2bV/iSZl71
8zCy4Lr0OnORtZ6VmWU7shIiPy2x7ng01K3nur750TbABercrB9mG+0CzaJyjAli
my0esuVWUgyJDEaxh6QIiNplwrvzSxAupZ5zfD9eqOTJsR0FwLFUItMufCNs1Ppl
THLJOeuKpScNzYZ4Bnna4QL2Wqo48pMuWcZOyEC+Zm0n5KGCFSiiR8z/LDH03NtS
fK3gBYnmA8OvuN0l0882UyoVO0ksXop7VkhDiKYDGD9TtGY9JSa59Ok8Dmwj3Fcq
fP5HAzHzYELuwSz/s0GTuX7tjd3KIEoQ9US+zAlOAyksEmQQ9ljQWBCDqLr1vr5X
SUxZhDeKCjvsi/8631U950FYSyYqYusQugtMD7GATv0uchXj1ofyb9ftFR6uB6zj
lG2B5lC/NaF3DnVBa8NkYf4ImofEQRDDfCwFNPG7VNH28j1AXyvYiU9nbOAO3hqJ
UcEttNOUFxvDfsxYR5nW0HQD7GmsBu8gyNhHT9asGiO2xpNZ/eFhvz/YJEqeEYRY
ctjm/Um+IB6XAOD6DWR2QX+8zmh6ttOG+5uuIoWbCuYHGk3jdBjxGo1o7kN4Z+HJ
r82uMmLW0nWo8Yo70diWUo6XTE4cWFZMgLqjlVt0SrztWXco+70rBiQEixBelIw/
XFwDBHQcRiFM2RfIBS34b07bov4ZcYtG2ETmf+mSHcz9mIJj6gNBK/qHJvyjyQ5y
yuAm0Bw9+qDGCKSdnYr+akob0ZdpCKQ49ttK7qNJ3RrajtvxG4l7e6h4Tajs4IAg
kWMJrZJbssCj1mNYHeC1VVmM5bci8xA8WmxWu/iVPn+Cuck2pPbC3YLQ64KsUhFT
gXDPjwh8U/ttfHDkiM0rDQiHufwiZ8KVJOjQDZUe5BCM0qsL1Fy3UXRjfX9xRhAo
p+Xrl3Bbv70SGBbRJk2NROE0zvLc0iMZRKs4LWiVqgrKJToNC/JBBeDpFpBqRJje
9rCL2M/j6i5L1uzpdUtJU7G5v6DKNCtv4LlaNX14UyfNlLE/myxf8P+0zTrL8GEu
qEYu3P8CLMXiJu77OUNDdReqnROERb2NC2ZErjrL66DXTw/I9XhhrTAOcSuzDMQW
7hiwSZlyifqVWLW64JlLhrtfBRq/PsmRD63OeV3haY6Y7QTUcs1QwnEtdiQEH3iE
kDrtPMVHsxK7tkPBLQQg7H00MB58kdxPDCBxWCGOwE2siSV5gS3D80kgxQ399ENv
LWJkKwSyeEAZpYBBIewDnjntR46zBRmJvldy9I0BujZjmD3TBuYB20Ivs5FkP3+G
4G5025Vz6b++if/jB+4Se2wKmzv4BfmOLyuzTFhGOqhG7IpW+ugInIUA8vwj2Bgi
XWaeuHlpSh0xGjBV9GFJCcaMCmkLb2Qm60MK+qg/H1nVul63gGh+lAgG+rptx+kq
GDmJrtEDmt5tu6BhqlnbvXW2mlFSSqxkmqze2462Oa5I1SQ4s59+gpZI/6zHiOZx
K71CX6oQaLDTec1/g5OaobUlk93uQX2dKeOu3kE49pgzfYb9RHaUZF+QNNh3Vkso
zbxuG55Z47xnJB2Ieda3xd0/8Kptg2+Vlcki8G1Jlqn4MjnAgodRLzj9uYQkcI8y
+0xelnjyIuwmF3vA4FPFU2pWC+IKmD9nLn+4JPn9oBY6x4IId8ramz2yXKXlzUo3
jBHY49bWqB/Wy4a6cO51G5vkRBn+IC7Wm3JHFAJ/NXr++fSPbIXvvVzrf0k0DDpP
SgHWXYLgEuQ1H25IVnU/QFBBfQb37hLynZn6AL4Sr7CwoDOt2NkcQZTQbADfAZpJ
iR6cK6OPaSK4pz8pt8uA68s7xxbInU3dA4TB8ciWdaDaTfuprHTYDQRqk0ZJx47Q
jkUUnuh+nnq5LY0mw0gN95f0d9Weo4kd1G7JBPOWRjn8y10W9jP5O1ogVoy1CRHR
dw2d0+kou+Mw1HzCz6TDBLgzn8iBKBfWruW26mIiwk4dPRTBoOIxekGqvshXX+Ev
CiIBYIgdAeD58B+brkO65Rv6c/mMjvURVfrYCjpdGdoDvgeSSrDCmiEYR7ziPoNV
22cklNx8drBurpyHWXkpX2pR8LgsT5jdmNqpInrrnc+nisQ6UmiQIIbjBCe+fuaa
tVayMN2b5KNKI2coGO7KsEi7ZQ4FPpPYSEIPm3LiuMZ6vZRYCntcdnBgLtCro93J
ni5VH+8QoWmkeG9FK1igXnz2lyC5MwL/0ZcphdepsYGjBLrS3Qpzl2QCyXFcI9mh
dbqNlOxc2uX3pMgyH+2ksNcfs2e9E1NAnLGW7Kprf8ScBBE8/VdEATpTbIeGxGwZ
JeerD0gDlXldCu0XvKOGGYLWKONRXd/wB8RP0u/F2oeXBrAJ1+evI6kxaNv7sJow
Dfhrj8xJD9CIvY97PR/4mFVLO2RyHpTgqm3H8ZpTLghamOFjOZu3cdXAcdjA3kJF
VnbwK4+4XJnGEqfP9KlGA2gJdIAW5DU+aU2JMDkkHGwTBteNjCx9BsX53Xt/ouAZ
QWRvt8vL8kVayJ0qUPNDYVkp+3mw1+6X9vYAuH/OVgGkJ83RNoM69h9N5ky44SYq
hX08nrKbbngCcXcm8ltDpMJN1qOIE5bAoZmJT4WxSF3B3qiKcjgz2vVlTerDxswM
HGs1hz93ctEPfiIBKsYp9+t1qsos0cX86vT+7Xv8+WFYDYC0uA9dYNWFjjpDF6On
6SQEEMxdB+5dDazznBfS6hefi4HCepMgMBR2d1/GbkKOTOGFnjn015Usn3rAsD60
0UqAc2hfzcFxZEG7afkw91uKTptCXIAPWyj137x3SHNxBd4J1oa3uYwHH6eRUzMi
v6WxYpd221gsVuqw47VusSORhnzJrWB83mt0YEbZpscTHHpC7XBnN1w0oBMJjAIm
UNNn1mrgwU2QHCyyR/mp/2n2F5h913oz6o5FdHpKWgk=
`protect END_PROTECTED
