`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9Y79r4pK7TrpnGtmzp5hGv1XHg9CItyM38P6Ltql+GhmnRtY5Hacs1+tgsI1qk15
W5gFqQ+jgpkX0m1PzxLn6mi4p32ZY4CAqIaqhutFxFtBNamzL8jqio9H54wQBKoL
KKloCqLJCfxf/ZSsw2SUDQamWAMunckIxSnHAR1jQljaEdsWtaEWgIRi/MXpcaoF
FMdOO7NbME1r98/qMgoENVUGDsnWICz3L+nRvLSLRuX8lte1KJTrp3LspRAqSqAU
bdDrpi5yAAoPs6l1qSepYSKc1OWbhmFXPt3Q9x5ByD7R9t5nEZQOSKfCJN3HHOLi
1UPqplQt+RR2YpWZiyJXowr4jp0BbL+4q7Dd7a8twz9wsz3sCpyi4uTV017psSkZ
rgqQ2llzuwVVOqXvQsNMp2QHzLfKoNHGedjtXVYcTk7bMR2bGJ+bbHgqp0RE9BSF
bdt5PbuDLxRAWi/XKPNrBswKaGftQ3R3gq6giDjWHTA+06K487vjT+UYuLassqCF
bHqV4D3XsjJ96kHTVIROSrNpPUueQolUY2D3qorv2LWcFiSnP8JcsYBNoAlIie83
aZxUxyhDXwrkXVj/t+EzEnrO47pUFaD2Bti5mN6VxQc=
`protect END_PROTECTED
