`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wzF2KXzfyMh0h7EcIKDSm1glAUCTc+x1aGDbcefqT6iOIL6ufsehe3cxQwUNr11R
sFTFdvXNteLEcMlDaadGUw0pw17rfMbZKkQ7BX7cdO12wqkPxr1SO20RR8hf9j1L
+QBm6NlR1fnh4ycEgSMT8fZCWRgieeO/w9ZklofTbn+VSSCECB1AjHVzfgZYJpze
Q5OguugnBYILFxnUZeihOm52AlNjqsuXmduWkFoYecSprpgC4v6DsN13KIBWUcZ1
OoPF2DtHGM4CmeoWmGk8m+NT0FpOnyOHldJuOqKi7c4JwppQcP0NOFyjh0aTAcOG
WF8f035jmSt/2iJBKnVagWZfPLjV5aGlHp+CiouYYA+Qf93zODLUPsNI21eVuMKc
M06CAKlV+9m8JgftvBLtqGM534n+H9ECH33XtrgYLrPCi5+IiMz7k/LWfawdI0dv
2iLC7y9WuD2WREuoaYtqwpYLZ01NLbAJscXSBsjTUY4mRiGo/5BROgRaSoVPVuJl
`protect END_PROTECTED
