`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JfrjvQhkGlvkuIFlLnxf5wNqf3JD67drNyvuc1NG5LmA/rMQLRp0lb5AysKzmNcY
gqletYbLsuy9ziD3Wl8dXyZJG+SQDMeAPqVFloJfrM1nGpkRQLMR5bncIdfEh/zL
kUNsRQBNisEzmBu/eqoqceYlNjf+ptR5XgfAcLT8C0cWRExtvPE/GSDmMwigNUbH
jAUBBZa9FMCAIj2LrLlCVUoHmekb2jFYYeYkbran2ekpLf2N9/ck7QrijLHkCZ2s
B0O+yrnWjoi5SwlH0KQYTx2mKamODjMx/UKHpyEEZ0m3Er4UA5PRPZgGWzjMRsBP
dLbpfgJXNbgmUHPvxA/q2g0LmQIUZMlJUcXQ3io38MmuVMp4Ryh+bf/94iawYUTD
1kaK33pt8GSKJ+FVS+OyvvspUyXuLlIcynWABAQecGpBAGXqjeh5b9vxWT8yTs+C
IgDcF6j0cdXTxj5sQefDvFLN8J8hawb1yaVLg1+6aYm+XWCfeMxCJIwCJ5TXetbi
a1KYeA47Do2oAuZGetKOd2nHOv9L/vH+Yfo1vgQamj8tm7M5eC8a9FBedJqjCXbM
f1Jllei8zGJ6NAhBID3lxU7CCQYK3dRpfj1fLNrKcmQD56nRqEsfIuVQplqtCmi2
soyRNXxvfgTz/qod3q3CF2l50FnZlpn5B6A+ytSefLfgni30iRPmyY8FuKaK9zhw
zMBO/yNAwPJWeNVv0C5ndn8JIxlr+HfBjuGQDL1Wt5M+Pncydz0YZ4XBsFhm+kG/
LQp2MsupxZWdzSiA/Za2Adb2W6Vn1sxJ96o6vqrDwuCMP1yX8Bxaak1CYME0DNR9
miEDmODuaUbjgFWPtP/zwrl0T9w+L2UbSx+rT6RHk+gh4LbYL21oVMhNyCVx5QVN
WAwBuIybGos8X8e0ZrSKkBRoLZYe5nHrCGgqqWvRKJVI6hmPYwCmUszKpZs9dSgs
i2ENvkEjX7IUVHAbLAwHFClLQTHmSJoCZFPXZgIAXC66Y5+QmA7djbXIj6jQZQ0Y
hhZOAqws81alD+OUgLO2X+mSs2YAKMwvZHbtI/IMCSOKaGPrTBg+D5s99tH7gQW0
uCRlp0HS1qwpUZiGYowHSienP+0HOxTEuib0BWUkJNPvc7uYyoFM5qbX5aBbjQlf
ZbNJFKXrIY4f/lJIhr/5SA==
`protect END_PROTECTED
