library verilog;
use verilog.vl_types.all;
entity cyclonev_hd_altpe2_hip_top is
    generic(
        func_mode       : string  := "disable";
        bonding_mode    : string  := "bond_disable";
        prot_mode       : string  := "disabled_prot_mode";
        pcie_spec_1p0_compliance: string  := "spec_1p1";
        vc_enable       : string  := "single_vc";
        enable_slot_register: string  := "false";
        pcie_mode       : string  := "shared_mode";
        multi_function  : string  := "one_fun";
        bypass_cdc      : string  := "false";
        cdc_clk_relation: string  := "plesiochronous";
        enable_rx_reordering: string  := "true";
        enable_rx_buffer_checking: string  := "false";
        single_rx_detect_data: vl_logic_vector(0 to 3) := (Hi0, Hi0, Hi0, Hi0);
        single_rx_detect: string  := "single_rx_detect";
        use_crc_forwarding: string  := "false";
        bypass_tl       : string  := "false";
        gen12_lane_rate_mode: string  := "gen1";
        lane_mask       : string  := "x4";
        disable_link_x2_support: string  := "false";
        national_inst_thru_enhance: string  := "true";
        disable_tag_check: string  := "enable";
        port_link_number_data: vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1);
        port_link_number: string  := "port_link_number";
        device_number_data: vl_logic_vector(0 to 4) := (Hi0, Hi0, Hi0, Hi0, Hi0);
        device_number   : string  := "device_number";
        bypass_clk_switch: string  := "false";
        core_clk_out_sel: string  := "div_1";
        core_clk_divider: string  := "div_1";
        core_clk_source : string  := "pll_fixed_clk";
        core_clk_sel    : string  := "pld_clk";
        disable_clk_switch: string  := "disable";
        core_clk_disable_clk_switch: string  := "pld_clk";
        slotclk_cfg     : string  := "dynamic_slotclkcfg";
        tx_swing_data   : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        tx_swing        : string  := "tx_swing";
        enable_ch0_pclk_out: string  := "pclk_ch01";
        enable_ch01_pclk_out: string  := "pclk_ch0";
        pipex1_debug_sel: string  := "disable";
        pclk_out_sel    : string  := "pclk";
        vendor_id_data_0: vl_logic_vector(0 to 15) := (Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi1, Hi0, Hi1, Hi1, Hi1, Hi0, Hi0, Hi1, Hi0);
        vendor_id_0     : string  := "vendor_id";
        device_id_data_0: vl_logic_vector(0 to 15) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1);
        device_id_0     : string  := "device_id";
        revision_id_data_0: vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1);
        revision_id_0   : string  := "revision_id";
        class_code_data_0: vl_logic_vector(0 to 23) := (Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        class_code_0    : string  := "class_code";
        subsystem_vendor_id_data_0: vl_logic_vector(0 to 15) := (Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi1, Hi0, Hi1, Hi1, Hi1, Hi0, Hi0, Hi1, Hi0);
        subsystem_vendor_id_0: string  := "subsystem_vendor_id";
        subsystem_device_id_data_0: vl_logic_vector(0 to 15) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1);
        subsystem_device_id_0: string  := "subsystem_device_id";
        no_soft_reset_0 : string  := "false";
        intel_id_access_0: string  := "false";
        device_specific_init_0: string  := "false";
        maximum_current_data_0: vl_logic_vector(0 to 2) := (Hi0, Hi0, Hi0);
        maximum_current_0: string  := "maximum_current";
        d1_support_0    : string  := "false";
        d2_support_0    : string  := "false";
        d0_pme_0        : string  := "false";
        d1_pme_0        : string  := "false";
        d2_pme_0        : string  := "false";
        d3_hot_pme_0    : string  := "false";
        d3_cold_pme_0   : string  := "false";
        use_aer_0       : string  := "false";
        low_priority_vc_0: string  := "single_vc";
        vc_arbitration_0: string  := "single_vc";
        disable_snoop_packet_0: string  := "false";
        max_payload_size_0: string  := "payload_512";
        surprise_down_error_support_0: string  := "false";
        dll_active_report_support_0: string  := "false";
        extend_tag_field_0: string  := "false";
        endpoint_l0_latency_data_0: vl_logic_vector(0 to 2) := (Hi0, Hi0, Hi0);
        endpoint_l0_latency_0: string  := "endpoint_l0_latency";
        endpoint_l1_latency_data_0: vl_logic_vector(0 to 2) := (Hi0, Hi0, Hi0);
        endpoint_l1_latency_0: string  := "endpoint_l1_latency";
        indicator_data_0: vl_logic_vector(0 to 2) := (Hi1, Hi1, Hi1);
        indicator_0     : string  := "indicator";
        role_based_error_reporting_0: string  := "false";
        slot_power_scale_data_0: vl_logic_vector(0 to 1) := (Hi0, Hi0);
        slot_power_scale_0: string  := "slot_power_scale";
        max_link_width_0: string  := "x4";
        enable_l1_aspm_0: string  := "false";
        enable_l0s_aspm_0: string  := "false";
        l1_exit_latency_sameclock_data_0: vl_logic_vector(0 to 2) := (Hi0, Hi0, Hi0);
        l1_exit_latency_sameclock_0: string  := "l1_exit_latency_sameclock";
        l1_exit_latency_diffclock_data_0: vl_logic_vector(0 to 2) := (Hi0, Hi0, Hi0);
        l1_exit_latency_diffclock_0: string  := "l1_exit_latency_diffclock";
        hot_plug_support_data_0: vl_logic_vector(0 to 6) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        hot_plug_support_0: string  := "hot_plug_support";
        slot_power_limit_data_0: vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        slot_power_limit_0: string  := "slot_power_limit";
        slot_number_data_0: vl_logic_vector(0 to 12) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        slot_number_0   : string  := "slot_number";
        diffclock_nfts_count_data_0: vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        diffclock_nfts_count_0: string  := "diffclock_nfts_count";
        sameclock_nfts_count_data_0: vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        sameclock_nfts_count_0: string  := "sameclock_nfts_count";
        completion_timeout_0: string  := "abcd";
        enable_completion_timeout_disable_0: string  := "true";
        extended_tag_reset_0: string  := "false";
        ecrc_check_capable_0: string  := "true";
        ecrc_gen_capable_0: string  := "true";
        no_command_completed_0: string  := "true";
        msi_multi_message_capable_0: string  := "count_4";
        msi_64bit_addressing_capable_0: string  := "true";
        msi_masking_capable_0: string  := "false";
        msi_support_0   : string  := "true";
        interrupt_pin_0 : string  := "inta";
        enable_function_msix_support_0: string  := "true";
        msix_table_size_data_0: vl_logic_vector(0 to 10) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        msix_table_size_0: string  := "msix_table_size";
        msix_table_bir_data_0: vl_logic_vector(0 to 2) := (Hi0, Hi0, Hi0);
        msix_table_bir_0: string  := "msix_table_bir";
        msix_table_offset_data_0: vl_logic_vector(0 to 28) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        msix_table_offset_0: string  := "msix_table_offset";
        msix_pba_bir_data_0: vl_logic_vector(0 to 2) := (Hi0, Hi0, Hi0);
        msix_pba_bir_0  : string  := "msix_pba_bir";
        msix_pba_offset_data_0: vl_logic_vector(0 to 28) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        msix_pba_offset_0: string  := "msix_pba_offset";
        bridge_port_vga_enable_0: string  := "false";
        bridge_port_ssid_support_0: string  := "false";
        ssvid_data_0    : vl_logic_vector(0 to 15) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        ssvid_0         : string  := "ssvid";
        ssid_data_0     : vl_logic_vector(0 to 15) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        ssid_0          : string  := "ssid";
        eie_before_nfts_count_data_0: vl_logic_vector(0 to 3) := (Hi0, Hi1, Hi0, Hi0);
        eie_before_nfts_count_0: string  := "eie_before_nfts_count";
        gen2_diffclock_nfts_count_data_0: vl_logic_vector(0 to 7) := (Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1);
        gen2_diffclock_nfts_count_0: string  := "gen2_diffclock_nfts_count";
        gen2_sameclock_nfts_count_data_0: vl_logic_vector(0 to 7) := (Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1);
        gen2_sameclock_nfts_count_0: string  := "gen2_sameclock_nfts_count";
        deemphasis_enable_0: string  := "false";
        pcie_spec_version_0: string  := "v2";
        l0_exit_latency_sameclock_data_0: vl_logic_vector(0 to 2) := (Hi1, Hi1, Hi0);
        l0_exit_latency_sameclock_0: string  := "l0_exit_latency_sameclock";
        l0_exit_latency_diffclock_data_0: vl_logic_vector(0 to 2) := (Hi1, Hi1, Hi0);
        l0_exit_latency_diffclock_0: string  := "l0_exit_latency_diffclock";
        rx_ei_l0s_0     : string  := "disable";
        l2_async_logic_0: string  := "enable";
        aspm_optionality_0: string  := "true";
        flr_capability_0: string  := "true";
        bar0_io_space_0 : string  := "false";
        bar0_64bit_mem_space_0: string  := "true";
        bar0_prefetchable_0: string  := "true";
        bar0_size_mask_data_0: vl_logic_vector(0 to 27) := (Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1);
        bar0_size_mask_0: string  := "bar0_size_mask";
        bar1_io_space_0 : string  := "false";
        bar1_64bit_mem_space_0: string  := "false";
        bar1_prefetchable_0: string  := "false";
        bar1_size_mask_data_0: vl_logic_vector(0 to 27) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        bar1_size_mask_0: string  := "bar1_size_mask";
        bar2_io_space_0 : string  := "false";
        bar2_64bit_mem_space_0: string  := "false";
        bar2_prefetchable_0: string  := "false";
        bar2_size_mask_data_0: vl_logic_vector(0 to 27) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        bar2_size_mask_0: string  := "bar2_size_mask";
        bar3_io_space_0 : string  := "false";
        bar3_64bit_mem_space_0: string  := "false";
        bar3_prefetchable_0: string  := "false";
        bar3_size_mask_data_0: vl_logic_vector(0 to 27) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        bar3_size_mask_0: string  := "bar3_size_mask";
        bar4_io_space_0 : string  := "false";
        bar4_64bit_mem_space_0: string  := "false";
        bar4_prefetchable_0: string  := "false";
        bar4_size_mask_data_0: vl_logic_vector(0 to 27) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        bar4_size_mask_0: string  := "bar4_size_mask";
        bar5_io_space_0 : string  := "false";
        bar5_64bit_mem_space_0: string  := "false";
        bar5_prefetchable_0: string  := "false";
        bar5_size_mask_data_0: vl_logic_vector(0 to 27) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        bar5_size_mask_0: string  := "bar5_size_mask";
        expansion_base_address_register_data_0: integer := 0;
        expansion_base_address_register_0: string  := "expansion_base_address_register";
        io_window_addr_width_0: string  := "window_32_bit";
        prefetchable_mem_window_addr_width_0: string  := "prefetch_32";
        vendor_id_data_1: vl_logic_vector(0 to 15) := (Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi1, Hi0, Hi1, Hi1, Hi1, Hi0, Hi0, Hi1, Hi0);
        vendor_id_1     : string  := "vendor_id";
        device_id_data_1: vl_logic_vector(0 to 15) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1);
        device_id_1     : string  := "device_id";
        revision_id_data_1: vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1);
        revision_id_1   : string  := "revision_id";
        class_code_data_1: vl_logic_vector(0 to 23) := (Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        class_code_1    : string  := "class_code";
        subsystem_vendor_id_data_1: vl_logic_vector(0 to 15) := (Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi1, Hi0, Hi1, Hi1, Hi1, Hi0, Hi0, Hi1, Hi0);
        subsystem_vendor_id_1: string  := "subsystem_vendor_id";
        subsystem_device_id_data_1: vl_logic_vector(0 to 15) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1);
        subsystem_device_id_1: string  := "subsystem_device_id";
        no_soft_reset_1 : string  := "false";
        intel_id_access_1: string  := "false";
        device_specific_init_1: string  := "false";
        maximum_current_data_1: vl_logic_vector(0 to 2) := (Hi0, Hi0, Hi0);
        maximum_current_1: string  := "maximum_current";
        d1_support_1    : string  := "false";
        d2_support_1    : string  := "false";
        d0_pme_1        : string  := "false";
        d1_pme_1        : string  := "false";
        d2_pme_1        : string  := "false";
        d3_hot_pme_1    : string  := "false";
        d3_cold_pme_1   : string  := "false";
        use_aer_1       : string  := "false";
        low_priority_vc_1: string  := "single_vc";
        vc_arbitration_1: string  := "single_vc";
        disable_snoop_packet_1: string  := "false";
        max_payload_size_1: string  := "payload_512";
        surprise_down_error_support_1: string  := "false";
        dll_active_report_support_1: string  := "false";
        extend_tag_field_1: string  := "false";
        endpoint_l0_latency_data_1: vl_logic_vector(0 to 2) := (Hi0, Hi0, Hi0);
        endpoint_l0_latency_1: string  := "endpoint_l0_latency";
        endpoint_l1_latency_data_1: vl_logic_vector(0 to 2) := (Hi0, Hi0, Hi0);
        endpoint_l1_latency_1: string  := "endpoint_l1_latency";
        indicator_data_1: vl_logic_vector(0 to 2) := (Hi1, Hi1, Hi1);
        indicator_1     : string  := "indicator";
        role_based_error_reporting_1: string  := "false";
        slot_power_scale_data_1: vl_logic_vector(0 to 1) := (Hi0, Hi0);
        slot_power_scale_1: string  := "slot_power_scale";
        max_link_width_1: string  := "x4";
        enable_l1_aspm_1: string  := "false";
        enable_l0s_aspm_1: string  := "false";
        l1_exit_latency_sameclock_data_1: vl_logic_vector(0 to 2) := (Hi0, Hi0, Hi0);
        l1_exit_latency_sameclock_1: string  := "l1_exit_latency_sameclock";
        l1_exit_latency_diffclock_data_1: vl_logic_vector(0 to 2) := (Hi0, Hi0, Hi0);
        l1_exit_latency_diffclock_1: string  := "l1_exit_latency_diffclock";
        hot_plug_support_data_1: vl_logic_vector(0 to 6) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        hot_plug_support_1: string  := "hot_plug_support";
        slot_power_limit_data_1: vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        slot_power_limit_1: string  := "slot_power_limit";
        slot_number_data_1: vl_logic_vector(0 to 12) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        slot_number_1   : string  := "slot_number";
        diffclock_nfts_count_data_1: vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        diffclock_nfts_count_1: string  := "diffclock_nfts_count";
        sameclock_nfts_count_data_1: vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        sameclock_nfts_count_1: string  := "sameclock_nfts_count";
        completion_timeout_1: string  := "abcd";
        enable_completion_timeout_disable_1: string  := "true";
        extended_tag_reset_1: string  := "false";
        ecrc_check_capable_1: string  := "true";
        ecrc_gen_capable_1: string  := "true";
        no_command_completed_1: string  := "true";
        msi_multi_message_capable_1: string  := "count_4";
        msi_64bit_addressing_capable_1: string  := "true";
        msi_masking_capable_1: string  := "false";
        msi_support_1   : string  := "true";
        interrupt_pin_1 : string  := "inta";
        enable_function_msix_support_1: string  := "true";
        msix_table_size_data_1: vl_logic_vector(0 to 10) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        msix_table_size_1: string  := "msix_table_size";
        msix_table_bir_data_1: vl_logic_vector(0 to 2) := (Hi0, Hi0, Hi0);
        msix_table_bir_1: string  := "msix_table_bir";
        msix_table_offset_data_1: vl_logic_vector(0 to 28) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        msix_table_offset_1: string  := "msix_table_offset";
        msix_pba_bir_data_1: vl_logic_vector(0 to 2) := (Hi0, Hi0, Hi0);
        msix_pba_bir_1  : string  := "msix_pba_bir";
        msix_pba_offset_data_1: vl_logic_vector(0 to 28) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        msix_pba_offset_1: string  := "msix_pba_offset";
        bridge_port_vga_enable_1: string  := "false";
        bridge_port_ssid_support_1: string  := "false";
        ssvid_data_1    : vl_logic_vector(0 to 15) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        ssvid_1         : string  := "ssvid";
        ssid_data_1     : vl_logic_vector(0 to 15) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        ssid_1          : string  := "ssid";
        eie_before_nfts_count_data_1: vl_logic_vector(0 to 3) := (Hi0, Hi1, Hi0, Hi0);
        eie_before_nfts_count_1: string  := "eie_before_nfts_count";
        gen2_diffclock_nfts_count_data_1: vl_logic_vector(0 to 7) := (Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1);
        gen2_diffclock_nfts_count_1: string  := "gen2_diffclock_nfts_count";
        gen2_sameclock_nfts_count_data_1: vl_logic_vector(0 to 7) := (Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1);
        gen2_sameclock_nfts_count_1: string  := "gen2_sameclock_nfts_count";
        deemphasis_enable_1: string  := "false";
        pcie_spec_version_1: string  := "v2";
        l0_exit_latency_sameclock_data_1: vl_logic_vector(0 to 2) := (Hi1, Hi1, Hi0);
        l0_exit_latency_sameclock_1: string  := "l0_exit_latency_sameclock";
        l0_exit_latency_diffclock_data_1: vl_logic_vector(0 to 2) := (Hi1, Hi1, Hi0);
        l0_exit_latency_diffclock_1: string  := "l0_exit_latency_diffclock";
        rx_ei_l0s_1     : string  := "disable";
        l2_async_logic_1: string  := "enable";
        aspm_optionality_1: string  := "true";
        flr_capability_1: string  := "true";
        bar0_io_space_1 : string  := "false";
        bar0_64bit_mem_space_1: string  := "true";
        bar0_prefetchable_1: string  := "true";
        bar0_size_mask_data_1: vl_logic_vector(0 to 27) := (Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1);
        bar0_size_mask_1: string  := "bar0_size_mask";
        bar1_io_space_1 : string  := "false";
        bar1_64bit_mem_space_1: string  := "false";
        bar1_prefetchable_1: string  := "false";
        bar1_size_mask_data_1: vl_logic_vector(0 to 27) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        bar1_size_mask_1: string  := "bar1_size_mask";
        bar2_io_space_1 : string  := "false";
        bar2_64bit_mem_space_1: string  := "false";
        bar2_prefetchable_1: string  := "false";
        bar2_size_mask_data_1: vl_logic_vector(0 to 27) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        bar2_size_mask_1: string  := "bar2_size_mask";
        bar3_io_space_1 : string  := "false";
        bar3_64bit_mem_space_1: string  := "false";
        bar3_prefetchable_1: string  := "false";
        bar3_size_mask_data_1: vl_logic_vector(0 to 27) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        bar3_size_mask_1: string  := "bar3_size_mask";
        bar4_io_space_1 : string  := "false";
        bar4_64bit_mem_space_1: string  := "false";
        bar4_prefetchable_1: string  := "false";
        bar4_size_mask_data_1: vl_logic_vector(0 to 27) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        bar4_size_mask_1: string  := "bar4_size_mask";
        bar5_io_space_1 : string  := "false";
        bar5_64bit_mem_space_1: string  := "false";
        bar5_prefetchable_1: string  := "false";
        bar5_size_mask_data_1: vl_logic_vector(0 to 27) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        bar5_size_mask_1: string  := "bar5_size_mask";
        expansion_base_address_register_data_1: integer := 0;
        expansion_base_address_register_1: string  := "expansion_base_address_register";
        io_window_addr_width_1: string  := "window_32_bit";
        prefetchable_mem_window_addr_width_1: string  := "prefetch_32";
        vendor_id_data_2: vl_logic_vector(0 to 15) := (Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi1, Hi0, Hi1, Hi1, Hi1, Hi0, Hi0, Hi1, Hi0);
        vendor_id_2     : string  := "vendor_id";
        device_id_data_2: vl_logic_vector(0 to 15) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1);
        device_id_2     : string  := "device_id";
        revision_id_data_2: vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1);
        revision_id_2   : string  := "revision_id";
        class_code_data_2: vl_logic_vector(0 to 23) := (Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        class_code_2    : string  := "class_code";
        subsystem_vendor_id_data_2: vl_logic_vector(0 to 15) := (Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi1, Hi0, Hi1, Hi1, Hi1, Hi0, Hi0, Hi1, Hi0);
        subsystem_vendor_id_2: string  := "subsystem_vendor_id";
        subsystem_device_id_data_2: vl_logic_vector(0 to 15) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1);
        subsystem_device_id_2: string  := "subsystem_device_id";
        no_soft_reset_2 : string  := "false";
        intel_id_access_2: string  := "false";
        device_specific_init_2: string  := "false";
        maximum_current_data_2: vl_logic_vector(0 to 2) := (Hi0, Hi0, Hi0);
        maximum_current_2: string  := "maximum_current";
        d1_support_2    : string  := "false";
        d2_support_2    : string  := "false";
        d0_pme_2        : string  := "false";
        d1_pme_2        : string  := "false";
        d2_pme_2        : string  := "false";
        d3_hot_pme_2    : string  := "false";
        d3_cold_pme_2   : string  := "false";
        use_aer_2       : string  := "false";
        low_priority_vc_2: string  := "single_vc";
        vc_arbitration_2: string  := "single_vc";
        disable_snoop_packet_2: string  := "false";
        max_payload_size_2: string  := "payload_512";
        surprise_down_error_support_2: string  := "false";
        dll_active_report_support_2: string  := "false";
        extend_tag_field_2: string  := "false";
        endpoint_l0_latency_data_2: vl_logic_vector(0 to 2) := (Hi0, Hi0, Hi0);
        endpoint_l0_latency_2: string  := "endpoint_l0_latency";
        endpoint_l1_latency_data_2: vl_logic_vector(0 to 2) := (Hi0, Hi0, Hi0);
        endpoint_l1_latency_2: string  := "endpoint_l1_latency";
        indicator_data_2: vl_logic_vector(0 to 2) := (Hi1, Hi1, Hi1);
        indicator_2     : string  := "indicator";
        role_based_error_reporting_2: string  := "false";
        slot_power_scale_data_2: vl_logic_vector(0 to 1) := (Hi0, Hi0);
        slot_power_scale_2: string  := "slot_power_scale";
        max_link_width_2: string  := "x4";
        enable_l1_aspm_2: string  := "false";
        enable_l0s_aspm_2: string  := "false";
        l1_exit_latency_sameclock_data_2: vl_logic_vector(0 to 2) := (Hi0, Hi0, Hi0);
        l1_exit_latency_sameclock_2: string  := "l1_exit_latency_sameclock";
        l1_exit_latency_diffclock_data_2: vl_logic_vector(0 to 2) := (Hi0, Hi0, Hi0);
        l1_exit_latency_diffclock_2: string  := "l1_exit_latency_diffclock";
        hot_plug_support_data_2: vl_logic_vector(0 to 6) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        hot_plug_support_2: string  := "hot_plug_support";
        slot_power_limit_data_2: vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        slot_power_limit_2: string  := "slot_power_limit";
        slot_number_data_2: vl_logic_vector(0 to 12) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        slot_number_2   : string  := "slot_number";
        diffclock_nfts_count_data_2: vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        diffclock_nfts_count_2: string  := "diffclock_nfts_count";
        sameclock_nfts_count_data_2: vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        sameclock_nfts_count_2: string  := "sameclock_nfts_count";
        completion_timeout_2: string  := "abcd";
        enable_completion_timeout_disable_2: string  := "true";
        extended_tag_reset_2: string  := "false";
        ecrc_check_capable_2: string  := "true";
        ecrc_gen_capable_2: string  := "true";
        no_command_completed_2: string  := "true";
        msi_multi_message_capable_2: string  := "count_4";
        msi_64bit_addressing_capable_2: string  := "true";
        msi_masking_capable_2: string  := "false";
        msi_support_2   : string  := "true";
        interrupt_pin_2 : string  := "inta";
        enable_function_msix_support_2: string  := "true";
        msix_table_size_data_2: vl_logic_vector(0 to 10) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        msix_table_size_2: string  := "msix_table_size";
        msix_table_bir_data_2: vl_logic_vector(0 to 2) := (Hi0, Hi0, Hi0);
        msix_table_bir_2: string  := "msix_table_bir";
        msix_table_offset_data_2: vl_logic_vector(0 to 28) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        msix_table_offset_2: string  := "msix_table_offset";
        msix_pba_bir_data_2: vl_logic_vector(0 to 2) := (Hi0, Hi0, Hi0);
        msix_pba_bir_2  : string  := "msix_pba_bir";
        msix_pba_offset_data_2: vl_logic_vector(0 to 28) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        msix_pba_offset_2: string  := "msix_pba_offset";
        bridge_port_vga_enable_2: string  := "false";
        bridge_port_ssid_support_2: string  := "false";
        ssvid_data_2    : vl_logic_vector(0 to 15) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        ssvid_2         : string  := "ssvid";
        ssid_data_2     : vl_logic_vector(0 to 15) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        ssid_2          : string  := "ssid";
        eie_before_nfts_count_data_2: vl_logic_vector(0 to 3) := (Hi0, Hi1, Hi0, Hi0);
        eie_before_nfts_count_2: string  := "eie_before_nfts_count";
        gen2_diffclock_nfts_count_data_2: vl_logic_vector(0 to 7) := (Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1);
        gen2_diffclock_nfts_count_2: string  := "gen2_diffclock_nfts_count";
        gen2_sameclock_nfts_count_data_2: vl_logic_vector(0 to 7) := (Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1);
        gen2_sameclock_nfts_count_2: string  := "gen2_sameclock_nfts_count";
        deemphasis_enable_2: string  := "false";
        pcie_spec_version_2: string  := "v2";
        l0_exit_latency_sameclock_data_2: vl_logic_vector(0 to 2) := (Hi1, Hi1, Hi0);
        l0_exit_latency_sameclock_2: string  := "l0_exit_latency_sameclock";
        l0_exit_latency_diffclock_data_2: vl_logic_vector(0 to 2) := (Hi1, Hi1, Hi0);
        l0_exit_latency_diffclock_2: string  := "l0_exit_latency_diffclock";
        rx_ei_l0s_2     : string  := "disable";
        l2_async_logic_2: string  := "enable";
        aspm_optionality_2: string  := "true";
        flr_capability_2: string  := "true";
        bar0_io_space_2 : string  := "false";
        bar0_64bit_mem_space_2: string  := "true";
        bar0_prefetchable_2: string  := "true";
        bar0_size_mask_data_2: vl_logic_vector(0 to 27) := (Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1);
        bar0_size_mask_2: string  := "bar0_size_mask";
        bar1_io_space_2 : string  := "false";
        bar1_64bit_mem_space_2: string  := "false";
        bar1_prefetchable_2: string  := "false";
        bar1_size_mask_data_2: vl_logic_vector(0 to 27) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        bar1_size_mask_2: string  := "bar1_size_mask";
        bar2_io_space_2 : string  := "false";
        bar2_64bit_mem_space_2: string  := "false";
        bar2_prefetchable_2: string  := "false";
        bar2_size_mask_data_2: vl_logic_vector(0 to 27) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        bar2_size_mask_2: string  := "bar2_size_mask";
        bar3_io_space_2 : string  := "false";
        bar3_64bit_mem_space_2: string  := "false";
        bar3_prefetchable_2: string  := "false";
        bar3_size_mask_data_2: vl_logic_vector(0 to 27) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        bar3_size_mask_2: string  := "bar3_size_mask";
        bar4_io_space_2 : string  := "false";
        bar4_64bit_mem_space_2: string  := "false";
        bar4_prefetchable_2: string  := "false";
        bar4_size_mask_data_2: vl_logic_vector(0 to 27) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        bar4_size_mask_2: string  := "bar4_size_mask";
        bar5_io_space_2 : string  := "false";
        bar5_64bit_mem_space_2: string  := "false";
        bar5_prefetchable_2: string  := "false";
        bar5_size_mask_data_2: vl_logic_vector(0 to 27) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        bar5_size_mask_2: string  := "bar5_size_mask";
        expansion_base_address_register_data_2: integer := 0;
        expansion_base_address_register_2: string  := "expansion_base_address_register";
        io_window_addr_width_2: string  := "window_32_bit";
        prefetchable_mem_window_addr_width_2: string  := "prefetch_32";
        vendor_id_data_3: vl_logic_vector(0 to 15) := (Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi1, Hi0, Hi1, Hi1, Hi1, Hi0, Hi0, Hi1, Hi0);
        vendor_id_3     : string  := "vendor_id";
        device_id_data_3: vl_logic_vector(0 to 15) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1);
        device_id_3     : string  := "device_id";
        revision_id_data_3: vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1);
        revision_id_3   : string  := "revision_id";
        class_code_data_3: vl_logic_vector(0 to 23) := (Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        class_code_3    : string  := "class_code";
        subsystem_vendor_id_data_3: vl_logic_vector(0 to 15) := (Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi1, Hi0, Hi1, Hi1, Hi1, Hi0, Hi0, Hi1, Hi0);
        subsystem_vendor_id_3: string  := "subsystem_vendor_id";
        subsystem_device_id_data_3: vl_logic_vector(0 to 15) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1);
        subsystem_device_id_3: string  := "subsystem_device_id";
        no_soft_reset_3 : string  := "false";
        intel_id_access_3: string  := "false";
        device_specific_init_3: string  := "false";
        maximum_current_data_3: vl_logic_vector(0 to 2) := (Hi0, Hi0, Hi0);
        maximum_current_3: string  := "maximum_current";
        d1_support_3    : string  := "false";
        d2_support_3    : string  := "false";
        d0_pme_3        : string  := "false";
        d1_pme_3        : string  := "false";
        d2_pme_3        : string  := "false";
        d3_hot_pme_3    : string  := "false";
        d3_cold_pme_3   : string  := "false";
        use_aer_3       : string  := "false";
        low_priority_vc_3: string  := "single_vc";
        vc_arbitration_3: string  := "single_vc";
        disable_snoop_packet_3: string  := "false";
        max_payload_size_3: string  := "payload_512";
        surprise_down_error_support_3: string  := "false";
        dll_active_report_support_3: string  := "false";
        extend_tag_field_3: string  := "false";
        endpoint_l0_latency_data_3: vl_logic_vector(0 to 2) := (Hi0, Hi0, Hi0);
        endpoint_l0_latency_3: string  := "endpoint_l0_latency";
        endpoint_l1_latency_data_3: vl_logic_vector(0 to 2) := (Hi0, Hi0, Hi0);
        endpoint_l1_latency_3: string  := "endpoint_l1_latency";
        indicator_data_3: vl_logic_vector(0 to 2) := (Hi1, Hi1, Hi1);
        indicator_3     : string  := "indicator";
        role_based_error_reporting_3: string  := "false";
        slot_power_scale_data_3: vl_logic_vector(0 to 1) := (Hi0, Hi0);
        slot_power_scale_3: string  := "slot_power_scale";
        max_link_width_3: string  := "x4";
        enable_l1_aspm_3: string  := "false";
        enable_l0s_aspm_3: string  := "false";
        l1_exit_latency_sameclock_data_3: vl_logic_vector(0 to 2) := (Hi0, Hi0, Hi0);
        l1_exit_latency_sameclock_3: string  := "l1_exit_latency_sameclock";
        l1_exit_latency_diffclock_data_3: vl_logic_vector(0 to 2) := (Hi0, Hi0, Hi0);
        l1_exit_latency_diffclock_3: string  := "l1_exit_latency_diffclock";
        hot_plug_support_data_3: vl_logic_vector(0 to 6) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        hot_plug_support_3: string  := "hot_plug_support";
        slot_power_limit_data_3: vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        slot_power_limit_3: string  := "slot_power_limit";
        slot_number_data_3: vl_logic_vector(0 to 12) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        slot_number_3   : string  := "slot_number";
        diffclock_nfts_count_data_3: vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        diffclock_nfts_count_3: string  := "diffclock_nfts_count";
        sameclock_nfts_count_data_3: vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        sameclock_nfts_count_3: string  := "sameclock_nfts_count";
        completion_timeout_3: string  := "abcd";
        enable_completion_timeout_disable_3: string  := "true";
        extended_tag_reset_3: string  := "false";
        ecrc_check_capable_3: string  := "true";
        ecrc_gen_capable_3: string  := "true";
        no_command_completed_3: string  := "true";
        msi_multi_message_capable_3: string  := "count_4";
        msi_64bit_addressing_capable_3: string  := "true";
        msi_masking_capable_3: string  := "false";
        msi_support_3   : string  := "true";
        interrupt_pin_3 : string  := "inta";
        enable_function_msix_support_3: string  := "true";
        msix_table_size_data_3: vl_logic_vector(0 to 10) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        msix_table_size_3: string  := "msix_table_size";
        msix_table_bir_data_3: vl_logic_vector(0 to 2) := (Hi0, Hi0, Hi0);
        msix_table_bir_3: string  := "msix_table_bir";
        msix_table_offset_data_3: vl_logic_vector(0 to 28) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        msix_table_offset_3: string  := "msix_table_offset";
        msix_pba_bir_data_3: vl_logic_vector(0 to 2) := (Hi0, Hi0, Hi0);
        msix_pba_bir_3  : string  := "msix_pba_bir";
        msix_pba_offset_data_3: vl_logic_vector(0 to 28) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        msix_pba_offset_3: string  := "msix_pba_offset";
        bridge_port_vga_enable_3: string  := "false";
        bridge_port_ssid_support_3: string  := "false";
        ssvid_data_3    : vl_logic_vector(0 to 15) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        ssvid_3         : string  := "ssvid";
        ssid_data_3     : vl_logic_vector(0 to 15) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        ssid_3          : string  := "ssid";
        eie_before_nfts_count_data_3: vl_logic_vector(0 to 3) := (Hi0, Hi1, Hi0, Hi0);
        eie_before_nfts_count_3: string  := "eie_before_nfts_count";
        gen2_diffclock_nfts_count_data_3: vl_logic_vector(0 to 7) := (Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1);
        gen2_diffclock_nfts_count_3: string  := "gen2_diffclock_nfts_count";
        gen2_sameclock_nfts_count_data_3: vl_logic_vector(0 to 7) := (Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1);
        gen2_sameclock_nfts_count_3: string  := "gen2_sameclock_nfts_count";
        deemphasis_enable_3: string  := "false";
        pcie_spec_version_3: string  := "v2";
        l0_exit_latency_sameclock_data_3: vl_logic_vector(0 to 2) := (Hi1, Hi1, Hi0);
        l0_exit_latency_sameclock_3: string  := "l0_exit_latency_sameclock";
        l0_exit_latency_diffclock_data_3: vl_logic_vector(0 to 2) := (Hi1, Hi1, Hi0);
        l0_exit_latency_diffclock_3: string  := "l0_exit_latency_diffclock";
        rx_ei_l0s_3     : string  := "disable";
        l2_async_logic_3: string  := "enable";
        aspm_optionality_3: string  := "true";
        flr_capability_3: string  := "true";
        bar0_io_space_3 : string  := "false";
        bar0_64bit_mem_space_3: string  := "true";
        bar0_prefetchable_3: string  := "true";
        bar0_size_mask_data_3: vl_logic_vector(0 to 27) := (Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1);
        bar0_size_mask_3: string  := "bar0_size_mask";
        bar1_io_space_3 : string  := "false";
        bar1_64bit_mem_space_3: string  := "false";
        bar1_prefetchable_3: string  := "false";
        bar1_size_mask_data_3: vl_logic_vector(0 to 27) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        bar1_size_mask_3: string  := "bar1_size_mask";
        bar2_io_space_3 : string  := "false";
        bar2_64bit_mem_space_3: string  := "false";
        bar2_prefetchable_3: string  := "false";
        bar2_size_mask_data_3: vl_logic_vector(0 to 27) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        bar2_size_mask_3: string  := "bar2_size_mask";
        bar3_io_space_3 : string  := "false";
        bar3_64bit_mem_space_3: string  := "false";
        bar3_prefetchable_3: string  := "false";
        bar3_size_mask_data_3: vl_logic_vector(0 to 27) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        bar3_size_mask_3: string  := "bar3_size_mask";
        bar4_io_space_3 : string  := "false";
        bar4_64bit_mem_space_3: string  := "false";
        bar4_prefetchable_3: string  := "false";
        bar4_size_mask_data_3: vl_logic_vector(0 to 27) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        bar4_size_mask_3: string  := "bar4_size_mask";
        bar5_io_space_3 : string  := "false";
        bar5_64bit_mem_space_3: string  := "false";
        bar5_prefetchable_3: string  := "false";
        bar5_size_mask_data_3: vl_logic_vector(0 to 27) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        bar5_size_mask_3: string  := "bar5_size_mask";
        expansion_base_address_register_data_3: integer := 0;
        expansion_base_address_register_3: string  := "expansion_base_address_register";
        io_window_addr_width_3: string  := "window_32_bit";
        prefetchable_mem_window_addr_width_3: string  := "prefetch_32";
        vendor_id_data_4: vl_logic_vector(0 to 15) := (Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi1, Hi0, Hi1, Hi1, Hi1, Hi0, Hi0, Hi1, Hi0);
        vendor_id_4     : string  := "vendor_id";
        device_id_data_4: vl_logic_vector(0 to 15) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1);
        device_id_4     : string  := "device_id";
        revision_id_data_4: vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1);
        revision_id_4   : string  := "revision_id";
        class_code_data_4: vl_logic_vector(0 to 23) := (Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        class_code_4    : string  := "class_code";
        subsystem_vendor_id_data_4: vl_logic_vector(0 to 15) := (Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi1, Hi0, Hi1, Hi1, Hi1, Hi0, Hi0, Hi1, Hi0);
        subsystem_vendor_id_4: string  := "subsystem_vendor_id";
        subsystem_device_id_data_4: vl_logic_vector(0 to 15) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1);
        subsystem_device_id_4: string  := "subsystem_device_id";
        no_soft_reset_4 : string  := "false";
        intel_id_access_4: string  := "false";
        device_specific_init_4: string  := "false";
        maximum_current_data_4: vl_logic_vector(0 to 2) := (Hi0, Hi0, Hi0);
        maximum_current_4: string  := "maximum_current";
        d1_support_4    : string  := "false";
        d2_support_4    : string  := "false";
        d0_pme_4        : string  := "false";
        d1_pme_4        : string  := "false";
        d2_pme_4        : string  := "false";
        d3_hot_pme_4    : string  := "false";
        d3_cold_pme_4   : string  := "false";
        use_aer_4       : string  := "false";
        low_priority_vc_4: string  := "single_vc";
        vc_arbitration_4: string  := "single_vc";
        disable_snoop_packet_4: string  := "false";
        max_payload_size_4: string  := "payload_512";
        surprise_down_error_support_4: string  := "false";
        dll_active_report_support_4: string  := "false";
        extend_tag_field_4: string  := "false";
        endpoint_l0_latency_data_4: vl_logic_vector(0 to 2) := (Hi0, Hi0, Hi0);
        endpoint_l0_latency_4: string  := "endpoint_l0_latency";
        endpoint_l1_latency_data_4: vl_logic_vector(0 to 2) := (Hi0, Hi0, Hi0);
        endpoint_l1_latency_4: string  := "endpoint_l1_latency";
        indicator_data_4: vl_logic_vector(0 to 2) := (Hi1, Hi1, Hi1);
        indicator_4     : string  := "indicator";
        role_based_error_reporting_4: string  := "false";
        slot_power_scale_data_4: vl_logic_vector(0 to 1) := (Hi0, Hi0);
        slot_power_scale_4: string  := "slot_power_scale";
        max_link_width_4: string  := "x4";
        enable_l1_aspm_4: string  := "false";
        enable_l0s_aspm_4: string  := "false";
        l1_exit_latency_sameclock_data_4: vl_logic_vector(0 to 2) := (Hi0, Hi0, Hi0);
        l1_exit_latency_sameclock_4: string  := "l1_exit_latency_sameclock";
        l1_exit_latency_diffclock_data_4: vl_logic_vector(0 to 2) := (Hi0, Hi0, Hi0);
        l1_exit_latency_diffclock_4: string  := "l1_exit_latency_diffclock";
        hot_plug_support_data_4: vl_logic_vector(0 to 6) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        hot_plug_support_4: string  := "hot_plug_support";
        slot_power_limit_data_4: vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        slot_power_limit_4: string  := "slot_power_limit";
        slot_number_data_4: vl_logic_vector(0 to 12) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        slot_number_4   : string  := "slot_number";
        diffclock_nfts_count_data_4: vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        diffclock_nfts_count_4: string  := "diffclock_nfts_count";
        sameclock_nfts_count_data_4: vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        sameclock_nfts_count_4: string  := "sameclock_nfts_count";
        completion_timeout_4: string  := "abcd";
        enable_completion_timeout_disable_4: string  := "true";
        extended_tag_reset_4: string  := "false";
        ecrc_check_capable_4: string  := "true";
        ecrc_gen_capable_4: string  := "true";
        no_command_completed_4: string  := "true";
        msi_multi_message_capable_4: string  := "count_4";
        msi_64bit_addressing_capable_4: string  := "true";
        msi_masking_capable_4: string  := "false";
        msi_support_4   : string  := "true";
        interrupt_pin_4 : string  := "inta";
        enable_function_msix_support_4: string  := "true";
        msix_table_size_data_4: vl_logic_vector(0 to 10) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        msix_table_size_4: string  := "msix_table_size";
        msix_table_bir_data_4: vl_logic_vector(0 to 2) := (Hi0, Hi0, Hi0);
        msix_table_bir_4: string  := "msix_table_bir";
        msix_table_offset_data_4: vl_logic_vector(0 to 28) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        msix_table_offset_4: string  := "msix_table_offset";
        msix_pba_bir_data_4: vl_logic_vector(0 to 2) := (Hi0, Hi0, Hi0);
        msix_pba_bir_4  : string  := "msix_pba_bir";
        msix_pba_offset_data_4: vl_logic_vector(0 to 28) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        msix_pba_offset_4: string  := "msix_pba_offset";
        bridge_port_vga_enable_4: string  := "false";
        bridge_port_ssid_support_4: string  := "false";
        ssvid_data_4    : vl_logic_vector(0 to 15) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        ssvid_4         : string  := "ssvid";
        ssid_data_4     : vl_logic_vector(0 to 15) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        ssid_4          : string  := "ssid";
        eie_before_nfts_count_data_4: vl_logic_vector(0 to 3) := (Hi0, Hi1, Hi0, Hi0);
        eie_before_nfts_count_4: string  := "eie_before_nfts_count";
        gen2_diffclock_nfts_count_data_4: vl_logic_vector(0 to 7) := (Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1);
        gen2_diffclock_nfts_count_4: string  := "gen2_diffclock_nfts_count";
        gen2_sameclock_nfts_count_data_4: vl_logic_vector(0 to 7) := (Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1);
        gen2_sameclock_nfts_count_4: string  := "gen2_sameclock_nfts_count";
        deemphasis_enable_4: string  := "false";
        pcie_spec_version_4: string  := "v2";
        l0_exit_latency_sameclock_data_4: vl_logic_vector(0 to 2) := (Hi1, Hi1, Hi0);
        l0_exit_latency_sameclock_4: string  := "l0_exit_latency_sameclock";
        l0_exit_latency_diffclock_data_4: vl_logic_vector(0 to 2) := (Hi1, Hi1, Hi0);
        l0_exit_latency_diffclock_4: string  := "l0_exit_latency_diffclock";
        rx_ei_l0s_4     : string  := "disable";
        l2_async_logic_4: string  := "enable";
        aspm_optionality_4: string  := "true";
        flr_capability_4: string  := "true";
        bar0_io_space_4 : string  := "false";
        bar0_64bit_mem_space_4: string  := "true";
        bar0_prefetchable_4: string  := "true";
        bar0_size_mask_data_4: vl_logic_vector(0 to 27) := (Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1);
        bar0_size_mask_4: string  := "bar0_size_mask";
        bar1_io_space_4 : string  := "false";
        bar1_64bit_mem_space_4: string  := "false";
        bar1_prefetchable_4: string  := "false";
        bar1_size_mask_data_4: vl_logic_vector(0 to 27) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        bar1_size_mask_4: string  := "bar1_size_mask";
        bar2_io_space_4 : string  := "false";
        bar2_64bit_mem_space_4: string  := "false";
        bar2_prefetchable_4: string  := "false";
        bar2_size_mask_data_4: vl_logic_vector(0 to 27) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        bar2_size_mask_4: string  := "bar2_size_mask";
        bar3_io_space_4 : string  := "false";
        bar3_64bit_mem_space_4: string  := "false";
        bar3_prefetchable_4: string  := "false";
        bar3_size_mask_data_4: vl_logic_vector(0 to 27) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        bar3_size_mask_4: string  := "bar3_size_mask";
        bar4_io_space_4 : string  := "false";
        bar4_64bit_mem_space_4: string  := "false";
        bar4_prefetchable_4: string  := "false";
        bar4_size_mask_data_4: vl_logic_vector(0 to 27) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        bar4_size_mask_4: string  := "bar4_size_mask";
        bar5_io_space_4 : string  := "false";
        bar5_64bit_mem_space_4: string  := "false";
        bar5_prefetchable_4: string  := "false";
        bar5_size_mask_data_4: vl_logic_vector(0 to 27) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        bar5_size_mask_4: string  := "bar5_size_mask";
        expansion_base_address_register_data_4: integer := 0;
        expansion_base_address_register_4: string  := "expansion_base_address_register";
        io_window_addr_width_4: string  := "window_32_bit";
        prefetchable_mem_window_addr_width_4: string  := "prefetch_32";
        vendor_id_data_5: vl_logic_vector(0 to 15) := (Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi1, Hi0, Hi1, Hi1, Hi1, Hi0, Hi0, Hi1, Hi0);
        vendor_id_5     : string  := "vendor_id";
        device_id_data_5: vl_logic_vector(0 to 15) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1);
        device_id_5     : string  := "device_id";
        revision_id_data_5: vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1);
        revision_id_5   : string  := "revision_id";
        class_code_data_5: vl_logic_vector(0 to 23) := (Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        class_code_5    : string  := "class_code";
        subsystem_vendor_id_data_5: vl_logic_vector(0 to 15) := (Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi1, Hi0, Hi1, Hi1, Hi1, Hi0, Hi0, Hi1, Hi0);
        subsystem_vendor_id_5: string  := "subsystem_vendor_id";
        subsystem_device_id_data_5: vl_logic_vector(0 to 15) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1);
        subsystem_device_id_5: string  := "subsystem_device_id";
        no_soft_reset_5 : string  := "false";
        intel_id_access_5: string  := "false";
        device_specific_init_5: string  := "false";
        maximum_current_data_5: vl_logic_vector(0 to 2) := (Hi0, Hi0, Hi0);
        maximum_current_5: string  := "maximum_current";
        d1_support_5    : string  := "false";
        d2_support_5    : string  := "false";
        d0_pme_5        : string  := "false";
        d1_pme_5        : string  := "false";
        d2_pme_5        : string  := "false";
        d3_hot_pme_5    : string  := "false";
        d3_cold_pme_5   : string  := "false";
        use_aer_5       : string  := "false";
        low_priority_vc_5: string  := "single_vc";
        vc_arbitration_5: string  := "single_vc";
        disable_snoop_packet_5: string  := "false";
        max_payload_size_5: string  := "payload_512";
        surprise_down_error_support_5: string  := "false";
        dll_active_report_support_5: string  := "false";
        extend_tag_field_5: string  := "false";
        endpoint_l0_latency_data_5: vl_logic_vector(0 to 2) := (Hi0, Hi0, Hi0);
        endpoint_l0_latency_5: string  := "endpoint_l0_latency";
        endpoint_l1_latency_data_5: vl_logic_vector(0 to 2) := (Hi0, Hi0, Hi0);
        endpoint_l1_latency_5: string  := "endpoint_l1_latency";
        indicator_data_5: vl_logic_vector(0 to 2) := (Hi1, Hi1, Hi1);
        indicator_5     : string  := "indicator";
        role_based_error_reporting_5: string  := "false";
        slot_power_scale_data_5: vl_logic_vector(0 to 1) := (Hi0, Hi0);
        slot_power_scale_5: string  := "slot_power_scale";
        max_link_width_5: string  := "x4";
        enable_l1_aspm_5: string  := "false";
        enable_l0s_aspm_5: string  := "false";
        l1_exit_latency_sameclock_data_5: vl_logic_vector(0 to 2) := (Hi0, Hi0, Hi0);
        l1_exit_latency_sameclock_5: string  := "l1_exit_latency_sameclock";
        l1_exit_latency_diffclock_data_5: vl_logic_vector(0 to 2) := (Hi0, Hi0, Hi0);
        l1_exit_latency_diffclock_5: string  := "l1_exit_latency_diffclock";
        hot_plug_support_data_5: vl_logic_vector(0 to 6) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        hot_plug_support_5: string  := "hot_plug_support";
        slot_power_limit_data_5: vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        slot_power_limit_5: string  := "slot_power_limit";
        slot_number_data_5: vl_logic_vector(0 to 12) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        slot_number_5   : string  := "slot_number";
        diffclock_nfts_count_data_5: vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        diffclock_nfts_count_5: string  := "diffclock_nfts_count";
        sameclock_nfts_count_data_5: vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        sameclock_nfts_count_5: string  := "sameclock_nfts_count";
        completion_timeout_5: string  := "abcd";
        enable_completion_timeout_disable_5: string  := "true";
        extended_tag_reset_5: string  := "false";
        ecrc_check_capable_5: string  := "true";
        ecrc_gen_capable_5: string  := "true";
        no_command_completed_5: string  := "true";
        msi_multi_message_capable_5: string  := "count_4";
        msi_64bit_addressing_capable_5: string  := "true";
        msi_masking_capable_5: string  := "false";
        msi_support_5   : string  := "true";
        interrupt_pin_5 : string  := "inta";
        enable_function_msix_support_5: string  := "true";
        msix_table_size_data_5: vl_logic_vector(0 to 10) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        msix_table_size_5: string  := "msix_table_size";
        msix_table_bir_data_5: vl_logic_vector(0 to 2) := (Hi0, Hi0, Hi0);
        msix_table_bir_5: string  := "msix_table_bir";
        msix_table_offset_data_5: vl_logic_vector(0 to 28) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        msix_table_offset_5: string  := "msix_table_offset";
        msix_pba_bir_data_5: vl_logic_vector(0 to 2) := (Hi0, Hi0, Hi0);
        msix_pba_bir_5  : string  := "msix_pba_bir";
        msix_pba_offset_data_5: vl_logic_vector(0 to 28) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        msix_pba_offset_5: string  := "msix_pba_offset";
        bridge_port_vga_enable_5: string  := "false";
        bridge_port_ssid_support_5: string  := "false";
        ssvid_data_5    : vl_logic_vector(0 to 15) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        ssvid_5         : string  := "ssvid";
        ssid_data_5     : vl_logic_vector(0 to 15) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        ssid_5          : string  := "ssid";
        eie_before_nfts_count_data_5: vl_logic_vector(0 to 3) := (Hi0, Hi1, Hi0, Hi0);
        eie_before_nfts_count_5: string  := "eie_before_nfts_count";
        gen2_diffclock_nfts_count_data_5: vl_logic_vector(0 to 7) := (Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1);
        gen2_diffclock_nfts_count_5: string  := "gen2_diffclock_nfts_count";
        gen2_sameclock_nfts_count_data_5: vl_logic_vector(0 to 7) := (Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1);
        gen2_sameclock_nfts_count_5: string  := "gen2_sameclock_nfts_count";
        deemphasis_enable_5: string  := "false";
        pcie_spec_version_5: string  := "v2";
        l0_exit_latency_sameclock_data_5: vl_logic_vector(0 to 2) := (Hi1, Hi1, Hi0);
        l0_exit_latency_sameclock_5: string  := "l0_exit_latency_sameclock";
        l0_exit_latency_diffclock_data_5: vl_logic_vector(0 to 2) := (Hi1, Hi1, Hi0);
        l0_exit_latency_diffclock_5: string  := "l0_exit_latency_diffclock";
        rx_ei_l0s_5     : string  := "disable";
        l2_async_logic_5: string  := "enable";
        aspm_optionality_5: string  := "true";
        flr_capability_5: string  := "true";
        bar0_io_space_5 : string  := "false";
        bar0_64bit_mem_space_5: string  := "true";
        bar0_prefetchable_5: string  := "true";
        bar0_size_mask_data_5: vl_logic_vector(0 to 27) := (Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1);
        bar0_size_mask_5: string  := "bar0_size_mask";
        bar1_io_space_5 : string  := "false";
        bar1_64bit_mem_space_5: string  := "false";
        bar1_prefetchable_5: string  := "false";
        bar1_size_mask_data_5: vl_logic_vector(0 to 27) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        bar1_size_mask_5: string  := "bar1_size_mask";
        bar2_io_space_5 : string  := "false";
        bar2_64bit_mem_space_5: string  := "false";
        bar2_prefetchable_5: string  := "false";
        bar2_size_mask_data_5: vl_logic_vector(0 to 27) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        bar2_size_mask_5: string  := "bar2_size_mask";
        bar3_io_space_5 : string  := "false";
        bar3_64bit_mem_space_5: string  := "false";
        bar3_prefetchable_5: string  := "false";
        bar3_size_mask_data_5: vl_logic_vector(0 to 27) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        bar3_size_mask_5: string  := "bar3_size_mask";
        bar4_io_space_5 : string  := "false";
        bar4_64bit_mem_space_5: string  := "false";
        bar4_prefetchable_5: string  := "false";
        bar4_size_mask_data_5: vl_logic_vector(0 to 27) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        bar4_size_mask_5: string  := "bar4_size_mask";
        bar5_io_space_5 : string  := "false";
        bar5_64bit_mem_space_5: string  := "false";
        bar5_prefetchable_5: string  := "false";
        bar5_size_mask_data_5: vl_logic_vector(0 to 27) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        bar5_size_mask_5: string  := "bar5_size_mask";
        expansion_base_address_register_data_5: integer := 0;
        expansion_base_address_register_5: string  := "expansion_base_address_register";
        io_window_addr_width_5: string  := "window_32_bit";
        prefetchable_mem_window_addr_width_5: string  := "prefetch_32";
        vendor_id_data_6: vl_logic_vector(0 to 15) := (Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi1, Hi0, Hi1, Hi1, Hi1, Hi0, Hi0, Hi1, Hi0);
        vendor_id_6     : string  := "vendor_id";
        device_id_data_6: vl_logic_vector(0 to 15) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1);
        device_id_6     : string  := "device_id";
        revision_id_data_6: vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1);
        revision_id_6   : string  := "revision_id";
        class_code_data_6: vl_logic_vector(0 to 23) := (Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        class_code_6    : string  := "class_code";
        subsystem_vendor_id_data_6: vl_logic_vector(0 to 15) := (Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi1, Hi0, Hi1, Hi1, Hi1, Hi0, Hi0, Hi1, Hi0);
        subsystem_vendor_id_6: string  := "subsystem_vendor_id";
        subsystem_device_id_data_6: vl_logic_vector(0 to 15) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1);
        subsystem_device_id_6: string  := "subsystem_device_id";
        no_soft_reset_6 : string  := "false";
        intel_id_access_6: string  := "false";
        device_specific_init_6: string  := "false";
        maximum_current_data_6: vl_logic_vector(0 to 2) := (Hi0, Hi0, Hi0);
        maximum_current_6: string  := "maximum_current";
        d1_support_6    : string  := "false";
        d2_support_6    : string  := "false";
        d0_pme_6        : string  := "false";
        d1_pme_6        : string  := "false";
        d2_pme_6        : string  := "false";
        d3_hot_pme_6    : string  := "false";
        d3_cold_pme_6   : string  := "false";
        use_aer_6       : string  := "false";
        low_priority_vc_6: string  := "single_vc";
        vc_arbitration_6: string  := "single_vc";
        disable_snoop_packet_6: string  := "false";
        max_payload_size_6: string  := "payload_512";
        surprise_down_error_support_6: string  := "false";
        dll_active_report_support_6: string  := "false";
        extend_tag_field_6: string  := "false";
        endpoint_l0_latency_data_6: vl_logic_vector(0 to 2) := (Hi0, Hi0, Hi0);
        endpoint_l0_latency_6: string  := "endpoint_l0_latency";
        endpoint_l1_latency_data_6: vl_logic_vector(0 to 2) := (Hi0, Hi0, Hi0);
        endpoint_l1_latency_6: string  := "endpoint_l1_latency";
        indicator_data_6: vl_logic_vector(0 to 2) := (Hi1, Hi1, Hi1);
        indicator_6     : string  := "indicator";
        role_based_error_reporting_6: string  := "false";
        slot_power_scale_data_6: vl_logic_vector(0 to 1) := (Hi0, Hi0);
        slot_power_scale_6: string  := "slot_power_scale";
        max_link_width_6: string  := "x4";
        enable_l1_aspm_6: string  := "false";
        enable_l0s_aspm_6: string  := "false";
        l1_exit_latency_sameclock_data_6: vl_logic_vector(0 to 2) := (Hi0, Hi0, Hi0);
        l1_exit_latency_sameclock_6: string  := "l1_exit_latency_sameclock";
        l1_exit_latency_diffclock_data_6: vl_logic_vector(0 to 2) := (Hi0, Hi0, Hi0);
        l1_exit_latency_diffclock_6: string  := "l1_exit_latency_diffclock";
        hot_plug_support_data_6: vl_logic_vector(0 to 6) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        hot_plug_support_6: string  := "hot_plug_support";
        slot_power_limit_data_6: vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        slot_power_limit_6: string  := "slot_power_limit";
        slot_number_data_6: vl_logic_vector(0 to 12) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        slot_number_6   : string  := "slot_number";
        diffclock_nfts_count_data_6: vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        diffclock_nfts_count_6: string  := "diffclock_nfts_count";
        sameclock_nfts_count_data_6: vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        sameclock_nfts_count_6: string  := "sameclock_nfts_count";
        completion_timeout_6: string  := "abcd";
        enable_completion_timeout_disable_6: string  := "true";
        extended_tag_reset_6: string  := "false";
        ecrc_check_capable_6: string  := "true";
        ecrc_gen_capable_6: string  := "true";
        no_command_completed_6: string  := "true";
        msi_multi_message_capable_6: string  := "count_4";
        msi_64bit_addressing_capable_6: string  := "true";
        msi_masking_capable_6: string  := "false";
        msi_support_6   : string  := "true";
        interrupt_pin_6 : string  := "inta";
        enable_function_msix_support_6: string  := "true";
        msix_table_size_data_6: vl_logic_vector(0 to 10) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        msix_table_size_6: string  := "msix_table_size";
        msix_table_bir_data_6: vl_logic_vector(0 to 2) := (Hi0, Hi0, Hi0);
        msix_table_bir_6: string  := "msix_table_bir";
        msix_table_offset_data_6: vl_logic_vector(0 to 28) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        msix_table_offset_6: string  := "msix_table_offset";
        msix_pba_bir_data_6: vl_logic_vector(0 to 2) := (Hi0, Hi0, Hi0);
        msix_pba_bir_6  : string  := "msix_pba_bir";
        msix_pba_offset_data_6: vl_logic_vector(0 to 28) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        msix_pba_offset_6: string  := "msix_pba_offset";
        bridge_port_vga_enable_6: string  := "false";
        bridge_port_ssid_support_6: string  := "false";
        ssvid_data_6    : vl_logic_vector(0 to 15) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        ssvid_6         : string  := "ssvid";
        ssid_data_6     : vl_logic_vector(0 to 15) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        ssid_6          : string  := "ssid";
        eie_before_nfts_count_data_6: vl_logic_vector(0 to 3) := (Hi0, Hi1, Hi0, Hi0);
        eie_before_nfts_count_6: string  := "eie_before_nfts_count";
        gen2_diffclock_nfts_count_data_6: vl_logic_vector(0 to 7) := (Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1);
        gen2_diffclock_nfts_count_6: string  := "gen2_diffclock_nfts_count";
        gen2_sameclock_nfts_count_data_6: vl_logic_vector(0 to 7) := (Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1);
        gen2_sameclock_nfts_count_6: string  := "gen2_sameclock_nfts_count";
        deemphasis_enable_6: string  := "false";
        pcie_spec_version_6: string  := "v2";
        l0_exit_latency_sameclock_data_6: vl_logic_vector(0 to 2) := (Hi1, Hi1, Hi0);
        l0_exit_latency_sameclock_6: string  := "l0_exit_latency_sameclock";
        l0_exit_latency_diffclock_data_6: vl_logic_vector(0 to 2) := (Hi1, Hi1, Hi0);
        l0_exit_latency_diffclock_6: string  := "l0_exit_latency_diffclock";
        rx_ei_l0s_6     : string  := "disable";
        l2_async_logic_6: string  := "enable";
        aspm_optionality_6: string  := "true";
        flr_capability_6: string  := "true";
        bar0_io_space_6 : string  := "false";
        bar0_64bit_mem_space_6: string  := "true";
        bar0_prefetchable_6: string  := "true";
        bar0_size_mask_data_6: vl_logic_vector(0 to 27) := (Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1);
        bar0_size_mask_6: string  := "bar0_size_mask";
        bar1_io_space_6 : string  := "false";
        bar1_64bit_mem_space_6: string  := "false";
        bar1_prefetchable_6: string  := "false";
        bar1_size_mask_data_6: vl_logic_vector(0 to 27) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        bar1_size_mask_6: string  := "bar1_size_mask";
        bar2_io_space_6 : string  := "false";
        bar2_64bit_mem_space_6: string  := "false";
        bar2_prefetchable_6: string  := "false";
        bar2_size_mask_data_6: vl_logic_vector(0 to 27) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        bar2_size_mask_6: string  := "bar2_size_mask";
        bar3_io_space_6 : string  := "false";
        bar3_64bit_mem_space_6: string  := "false";
        bar3_prefetchable_6: string  := "false";
        bar3_size_mask_data_6: vl_logic_vector(0 to 27) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        bar3_size_mask_6: string  := "bar3_size_mask";
        bar4_io_space_6 : string  := "false";
        bar4_64bit_mem_space_6: string  := "false";
        bar4_prefetchable_6: string  := "false";
        bar4_size_mask_data_6: vl_logic_vector(0 to 27) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        bar4_size_mask_6: string  := "bar4_size_mask";
        bar5_io_space_6 : string  := "false";
        bar5_64bit_mem_space_6: string  := "false";
        bar5_prefetchable_6: string  := "false";
        bar5_size_mask_data_6: vl_logic_vector(0 to 27) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        bar5_size_mask_6: string  := "bar5_size_mask";
        expansion_base_address_register_data_6: integer := 0;
        expansion_base_address_register_6: string  := "expansion_base_address_register";
        io_window_addr_width_6: string  := "window_32_bit";
        prefetchable_mem_window_addr_width_6: string  := "prefetch_32";
        vendor_id_data_7: vl_logic_vector(0 to 15) := (Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi1, Hi0, Hi1, Hi1, Hi1, Hi0, Hi0, Hi1, Hi0);
        vendor_id_7     : string  := "vendor_id";
        device_id_data_7: vl_logic_vector(0 to 15) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1);
        device_id_7     : string  := "device_id";
        revision_id_data_7: vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1);
        revision_id_7   : string  := "revision_id";
        class_code_data_7: vl_logic_vector(0 to 23) := (Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        class_code_7    : string  := "class_code";
        subsystem_vendor_id_data_7: vl_logic_vector(0 to 15) := (Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi1, Hi0, Hi1, Hi1, Hi1, Hi0, Hi0, Hi1, Hi0);
        subsystem_vendor_id_7: string  := "subsystem_vendor_id";
        subsystem_device_id_data_7: vl_logic_vector(0 to 15) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1);
        subsystem_device_id_7: string  := "subsystem_device_id";
        no_soft_reset_7 : string  := "false";
        intel_id_access_7: string  := "false";
        device_specific_init_7: string  := "false";
        maximum_current_data_7: vl_logic_vector(0 to 2) := (Hi0, Hi0, Hi0);
        maximum_current_7: string  := "maximum_current";
        d1_support_7    : string  := "false";
        d2_support_7    : string  := "false";
        d0_pme_7        : string  := "false";
        d1_pme_7        : string  := "false";
        d2_pme_7        : string  := "false";
        d3_hot_pme_7    : string  := "false";
        d3_cold_pme_7   : string  := "false";
        use_aer_7       : string  := "false";
        low_priority_vc_7: string  := "single_vc";
        vc_arbitration_7: string  := "single_vc";
        disable_snoop_packet_7: string  := "false";
        max_payload_size_7: string  := "payload_512";
        surprise_down_error_support_7: string  := "false";
        dll_active_report_support_7: string  := "false";
        extend_tag_field_7: string  := "false";
        endpoint_l0_latency_data_7: vl_logic_vector(0 to 2) := (Hi0, Hi0, Hi0);
        endpoint_l0_latency_7: string  := "endpoint_l0_latency";
        endpoint_l1_latency_data_7: vl_logic_vector(0 to 2) := (Hi0, Hi0, Hi0);
        endpoint_l1_latency_7: string  := "endpoint_l1_latency";
        indicator_data_7: vl_logic_vector(0 to 2) := (Hi1, Hi1, Hi1);
        indicator_7     : string  := "indicator";
        role_based_error_reporting_7: string  := "false";
        slot_power_scale_data_7: vl_logic_vector(0 to 1) := (Hi0, Hi0);
        slot_power_scale_7: string  := "slot_power_scale";
        max_link_width_7: string  := "x4";
        enable_l1_aspm_7: string  := "false";
        enable_l0s_aspm_7: string  := "false";
        l1_exit_latency_sameclock_data_7: vl_logic_vector(0 to 2) := (Hi0, Hi0, Hi0);
        l1_exit_latency_sameclock_7: string  := "l1_exit_latency_sameclock";
        l1_exit_latency_diffclock_data_7: vl_logic_vector(0 to 2) := (Hi0, Hi0, Hi0);
        l1_exit_latency_diffclock_7: string  := "l1_exit_latency_diffclock";
        hot_plug_support_data_7: vl_logic_vector(0 to 6) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        hot_plug_support_7: string  := "hot_plug_support";
        slot_power_limit_data_7: vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        slot_power_limit_7: string  := "slot_power_limit";
        slot_number_data_7: vl_logic_vector(0 to 12) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        slot_number_7   : string  := "slot_number";
        diffclock_nfts_count_data_7: vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        diffclock_nfts_count_7: string  := "diffclock_nfts_count";
        sameclock_nfts_count_data_7: vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        sameclock_nfts_count_7: string  := "sameclock_nfts_count";
        completion_timeout_7: string  := "abcd";
        enable_completion_timeout_disable_7: string  := "true";
        extended_tag_reset_7: string  := "false";
        ecrc_check_capable_7: string  := "true";
        ecrc_gen_capable_7: string  := "true";
        no_command_completed_7: string  := "true";
        msi_multi_message_capable_7: string  := "count_4";
        msi_64bit_addressing_capable_7: string  := "true";
        msi_masking_capable_7: string  := "false";
        msi_support_7   : string  := "true";
        interrupt_pin_7 : string  := "inta";
        enable_function_msix_support_7: string  := "true";
        msix_table_size_data_7: vl_logic_vector(0 to 10) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        msix_table_size_7: string  := "msix_table_size";
        msix_table_bir_data_7: vl_logic_vector(0 to 2) := (Hi0, Hi0, Hi0);
        msix_table_bir_7: string  := "msix_table_bir";
        msix_table_offset_data_7: vl_logic_vector(0 to 28) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        msix_table_offset_7: string  := "msix_table_offset";
        msix_pba_bir_data_7: vl_logic_vector(0 to 2) := (Hi0, Hi0, Hi0);
        msix_pba_bir_7  : string  := "msix_pba_bir";
        msix_pba_offset_data_7: vl_logic_vector(0 to 28) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        msix_pba_offset_7: string  := "msix_pba_offset";
        bridge_port_vga_enable_7: string  := "false";
        bridge_port_ssid_support_7: string  := "false";
        ssvid_data_7    : vl_logic_vector(0 to 15) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        ssvid_7         : string  := "ssvid";
        ssid_data_7     : vl_logic_vector(0 to 15) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        ssid_7          : string  := "ssid";
        eie_before_nfts_count_data_7: vl_logic_vector(0 to 3) := (Hi0, Hi1, Hi0, Hi0);
        eie_before_nfts_count_7: string  := "eie_before_nfts_count";
        gen2_diffclock_nfts_count_data_7: vl_logic_vector(0 to 7) := (Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1);
        gen2_diffclock_nfts_count_7: string  := "gen2_diffclock_nfts_count";
        gen2_sameclock_nfts_count_data_7: vl_logic_vector(0 to 7) := (Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1);
        gen2_sameclock_nfts_count_7: string  := "gen2_sameclock_nfts_count";
        deemphasis_enable_7: string  := "false";
        pcie_spec_version_7: string  := "v2";
        l0_exit_latency_sameclock_data_7: vl_logic_vector(0 to 2) := (Hi1, Hi1, Hi0);
        l0_exit_latency_sameclock_7: string  := "l0_exit_latency_sameclock";
        l0_exit_latency_diffclock_data_7: vl_logic_vector(0 to 2) := (Hi1, Hi1, Hi0);
        l0_exit_latency_diffclock_7: string  := "l0_exit_latency_diffclock";
        rx_ei_l0s_7     : string  := "disable";
        l2_async_logic_7: string  := "enable";
        aspm_optionality_7: string  := "true";
        flr_capability_7: string  := "true";
        bar0_io_space_7 : string  := "false";
        bar0_64bit_mem_space_7: string  := "true";
        bar0_prefetchable_7: string  := "true";
        bar0_size_mask_data_7: vl_logic_vector(0 to 27) := (Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1);
        bar0_size_mask_7: string  := "bar0_size_mask";
        bar1_io_space_7 : string  := "false";
        bar1_64bit_mem_space_7: string  := "false";
        bar1_prefetchable_7: string  := "false";
        bar1_size_mask_data_7: vl_logic_vector(0 to 27) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        bar1_size_mask_7: string  := "bar1_size_mask";
        bar2_io_space_7 : string  := "false";
        bar2_64bit_mem_space_7: string  := "false";
        bar2_prefetchable_7: string  := "false";
        bar2_size_mask_data_7: vl_logic_vector(0 to 27) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        bar2_size_mask_7: string  := "bar2_size_mask";
        bar3_io_space_7 : string  := "false";
        bar3_64bit_mem_space_7: string  := "false";
        bar3_prefetchable_7: string  := "false";
        bar3_size_mask_data_7: vl_logic_vector(0 to 27) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        bar3_size_mask_7: string  := "bar3_size_mask";
        bar4_io_space_7 : string  := "false";
        bar4_64bit_mem_space_7: string  := "false";
        bar4_prefetchable_7: string  := "false";
        bar4_size_mask_data_7: vl_logic_vector(0 to 27) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        bar4_size_mask_7: string  := "bar4_size_mask";
        bar5_io_space_7 : string  := "false";
        bar5_64bit_mem_space_7: string  := "false";
        bar5_prefetchable_7: string  := "false";
        bar5_size_mask_data_7: vl_logic_vector(0 to 27) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        bar5_size_mask_7: string  := "bar5_size_mask";
        expansion_base_address_register_data_7: integer := 0;
        expansion_base_address_register_7: string  := "expansion_base_address_register";
        io_window_addr_width_7: string  := "window_32_bit";
        prefetchable_mem_window_addr_width_7: string  := "prefetch_32";
        porttype_func0  : string  := "ep_native";
        porttype_func1  : string  := "ep_native";
        porttype_func2  : string  := "ep_native";
        porttype_func3  : string  := "ep_native";
        porttype_func4  : string  := "ep_native";
        porttype_func5  : string  := "ep_native";
        porttype_func6  : string  := "ep_native";
        porttype_func7  : string  := "ep_native";
        rxfreqlk_cnt_data: vl_logic_vector(0 to 19) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        rxfreqlk_cnt    : string  := "rxfreqlk_prog_cnt";
        rxfreqlk_cnt_en : string  := "true";
        testmode_control: string  := "disable";
        skp_insertion_control: string  := "disable";
        tx_l0s_adjust   : string  := "disable";
        rx_cdc_almost_full_data: vl_logic_vector(0 to 3) := (Hi0, Hi0, Hi0, Hi0);
        rx_cdc_almost_full: string  := "rx_cdc_almost_full";
        tx_cdc_almost_full_data: vl_logic_vector(0 to 3) := (Hi0, Hi0, Hi0, Hi0);
        tx_cdc_almost_full: string  := "tx_cdc_almost_full";
        rx_l0s_count_idl_data: vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        rx_l0s_count_idl: string  := "rx_l0s_count_idl";
        cdc_dummy_insert_limit_data: vl_logic_vector(0 to 3) := (Hi0, Hi0, Hi0, Hi0);
        cdc_dummy_insert_limit: string  := "cdc_dummy_insert_limit";
        ei_delay_powerdown_count_data: vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi1, Hi0);
        ei_delay_powerdown_count: string  := "ei_delay_powerdown_count";
        millisecond_cycle_count_data: vl_logic_vector(0 to 19) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        millisecond_cycle_count: string  := "millisecond_cycle_count";
        skp_os_schedule_count_data: vl_logic_vector(0 to 10) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        skp_os_schedule_count: string  := "skp_os_schedule_count";
        fc_init_timer_data: vl_logic_vector(0 to 10) := (Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        fc_init_timer   : string  := "fc_init_timer";
        l01_entry_latency_data: vl_logic_vector(0 to 4) := (Hi1, Hi1, Hi1, Hi1, Hi1);
        l01_entry_latency: string  := "l01_entry_latency";
        flow_control_update_count_data: vl_logic_vector(0 to 4) := (Hi1, Hi1, Hi1, Hi1, Hi0);
        flow_control_update_count: string  := "flow_control_update_count";
        flow_control_timeout_count_data: vl_logic_vector(0 to 7) := (Hi1, Hi1, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0);
        flow_control_timeout_count: string  := "flow_control_timeout_count";
        vc0_rx_flow_ctrl_posted_header_data: vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi1, Hi1, Hi0, Hi0, Hi1, Hi0);
        vc0_rx_flow_ctrl_posted_header: string  := "vc0_rx_flow_ctrl_posted_header";
        vc0_rx_flow_ctrl_posted_data_data: vl_logic_vector(0 to 11) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi1, Hi1, Hi1, Hi1, Hi0);
        vc0_rx_flow_ctrl_posted_data: string  := "vc0_rx_flow_ctrl_posted_data";
        vc0_rx_flow_ctrl_nonposted_header_data: vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0);
        vc0_rx_flow_ctrl_nonposted_header: string  := "vc0_rx_flow_ctrl_nonposted_header";
        vc0_rx_flow_ctrl_nonposted_data_data: vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        vc0_rx_flow_ctrl_nonposted_data: string  := "vc0_rx_flow_ctrl_nonposted_data";
        vc0_rx_flow_ctrl_compl_header_data: vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        vc0_rx_flow_ctrl_compl_header: string  := "vc0_rx_flow_ctrl_compl_header";
        vc0_rx_flow_ctrl_compl_data_data: vl_logic_vector(0 to 11) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        vc0_rx_flow_ctrl_compl_data: string  := "vc0_rx_flow_ctrl_compl_data";
        rx_ptr0_posted_dpram_min_data: vl_logic_vector(0 to 9) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        rx_ptr0_posted_dpram_min: string  := "rx_ptr0_posted_dpram_min";
        rx_ptr0_posted_dpram_max_data: vl_logic_vector(0 to 9) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        rx_ptr0_posted_dpram_max: string  := "rx_ptr0_posted_dpram_max";
        rx_ptr0_nonposted_dpram_min_data: vl_logic_vector(0 to 9) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        rx_ptr0_nonposted_dpram_min: string  := "rx_ptr0_nonposted_dpram_min";
        rx_ptr0_nonposted_dpram_max_data: vl_logic_vector(0 to 9) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        rx_ptr0_nonposted_dpram_max: string  := "rx_ptr0_nonposted_dpram_max";
        retry_buffer_last_active_address_data: vl_logic_vector(0 to 7) := (Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1);
        retry_buffer_memory_settings_data: vl_logic_vector(0 to 15) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi1, Hi0);
        retry_buffer_memory_settings: string  := "retry_buffer_memory_settings";
        vc0_rx_buffer_memory_settings_data: vl_logic_vector(0 to 15) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi1, Hi0);
        vc0_rx_buffer_memory_settings: string  := "vc0_rx_buffer_memory_settings";
        bist_memory_settings_data: vl_logic_vector(0 to 74) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        bist_memory_settings: string  := "bist_memory_settings";
        bridge_66mhzcap : string  := "true";
        fastb2bcap      : string  := "true";
        devseltim       : string  := "fast_devsel_decoding";
        memwrinv        : string  := "ro";
        credit_buffer_allocation_aux: string  := "balanced";
        enable_adapter_half_rate_mode: string  := "false";
        vc0_clk_enable  : string  := "true";
        vc1_clk_enable  : string  := "false";
        register_pipe_signals: string  := "false";
        iei_enable_settings: string  := "gen2_infei_infsd_gen1_infei_sd";
        lattim_ro_data  : vl_logic_vector(0 to 6) := (Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0);
        lattim          : string  := "ro";
        br_rcb          : string  := "ro";
        vsec_id_data    : vl_logic_vector(0 to 15) := (Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi1, Hi0, Hi1, Hi1, Hi1, Hi0, Hi0, Hi1, Hi0);
        vsec_id         : string  := "vsec_id";
        cvp_enable      : string  := "cvp_dis";
        cvp_rate_sel    : string  := "full_rate";
        hard_reset_bypass: string  := "false";
        cvp_data_compressed: string  := "false";
        cvp_data_encrypted: string  := "false";
        cvp_mode_reset  : string  := "false";
        cvp_clk_reset   : string  := "false";
        vsec_cap_data   : vl_logic_vector(0 to 3) := (Hi0, Hi0, Hi0, Hi0);
        vsec_cap        : string  := "vsec_cap";
        jtag_id_data    : vl_logic_vector(0 to 127) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        jtag_id         : string  := "jtag_id";
        user_id_data    : vl_logic_vector(0 to 15) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        user_id         : string  := "user_id";
        disable_auto_crs: string  := "disable";
        altpe2_hip_base_addr_1: integer := 0;
        altpe2_hip_base_addr_2: integer := 0;
        altpe2_hip_base_addr_3: integer := 0;
        altpe2_hip_base_addr_4: integer := 0;
        altpe2_hip_base_addr_5: integer := 0;
        altpe2_hip_base_addr_6: integer := 0;
        altpe2_hip_base_addr_user_1: vl_logic_vector(0 to 9) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        altpe2_hip_base_addr_user_2: vl_logic_vector(0 to 9) := (Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        altpe2_hip_base_addr_user_3: vl_logic_vector(0 to 9) := (Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        altpe2_hip_base_addr_user_4: vl_logic_vector(0 to 9) := (Hi0, Hi0, Hi1, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        altpe2_hip_base_addr_user_5: vl_logic_vector(0 to 9) := (Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        altpe2_hip_base_addr_user_6: vl_logic_vector(0 to 9) := (Hi0, Hi1, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        cvp_mdio_dis_csr_ctrl_1: string  := "mdio_dis_cvp_dis";
        cvp_mdio_dis_csr_ctrl_2: string  := "mdio_dis_cvp_dis";
        cvp_mdio_dis_csr_ctrl_3: string  := "mdio_dis_cvp_dis";
        cvp_mdio_dis_csr_ctrl_4: string  := "mdio_dis_cvp_dis";
        cvp_mdio_dis_csr_ctrl_5: string  := "mdio_dis_cvp_dis";
        cvp_mdio_dis_csr_ctrl_6: string  := "mdio_dis_cvp_dis";
        dft_broadcast_en_1: string  := "broadcast_dis";
        dft_broadcast_en_2: string  := "broadcast_dis";
        dft_broadcast_en_3: string  := "broadcast_dis";
        dft_broadcast_en_4: string  := "broadcast_dis";
        dft_broadcast_en_5: string  := "broadcast_dis";
        dft_broadcast_en_6: string  := "broadcast_dis";
        electromech_interlock_0: string  := "false";
        electromech_interlock_1: string  := "false";
        electromech_interlock_2: string  := "false";
        electromech_interlock_3: string  := "false";
        electromech_interlock_4: string  := "false";
        electromech_interlock_5: string  := "false";
        electromech_interlock_6: string  := "false";
        electromech_interlock_7: string  := "false";
        force_mdio_dis_csr_ctrl_1: string  := "mdio_dis_force_dis";
        force_mdio_dis_csr_ctrl_2: string  := "mdio_dis_force_dis";
        force_mdio_dis_csr_ctrl_3: string  := "mdio_dis_force_dis";
        force_mdio_dis_csr_ctrl_4: string  := "mdio_dis_force_dis";
        force_mdio_dis_csr_ctrl_5: string  := "mdio_dis_force_dis";
        force_mdio_dis_csr_ctrl_6: string  := "mdio_dis_force_dis";
        mdio_cb_opbit_enable: string  := "enable";
        plniotri_gate   : string  := "disable";
        power_isolation_en_1: string  := "power_isolation_dis";
        power_isolation_en_1_data: vl_logic := Hi0;
        power_isolation_en_2: string  := "power_isolation_dis";
        power_isolation_en_2_data: vl_logic := Hi0;
        power_isolation_en_3: string  := "power_isolation_dis";
        power_isolation_en_3_data: vl_logic := Hi0;
        power_isolation_en_4: string  := "power_isolation_dis";
        power_isolation_en_4_data: vl_logic := Hi0;
        power_isolation_en_5: string  := "power_isolation_dis";
        power_isolation_en_5_data: vl_logic := Hi0;
        power_isolation_en_6: string  := "power_isolation_dis";
        power_isolation_en_6_data: vl_logic := Hi0;
        retry_buffer_last_active_address: string  := "retry_buffer_last_active_address";
        sup_mode        : string  := "user_mode";
        hrdrstctrl_en   : string  := "hrdrstctrl_dis";
        rstctrl_pld_clr : string  := "false";
        rstctrl_debug_en: string  := "false";
        rstctrl_force_inactive_rst: string  := "false";
        rstctrl_perst_enable: string  := "level";
        rstctrl_hip_ep  : string  := "hip_ep";
        rstctrl_hard_block_enable: string  := "hard_rst_ctl";
        rstctrl_rx_pma_rstb_inv: string  := "false";
        rstctrl_tx_pma_rstb_inv: string  := "false";
        rstctrl_rx_pcs_rst_n_inv: string  := "false";
        rstctrl_tx_pcs_rst_n_inv: string  := "false";
        rstctrl_altpe2_crst_n_inv: string  := "false";
        rstctrl_altpe2_srst_n_inv: string  := "false";
        rstctrl_altpe2_rst_n_inv: string  := "false";
        rstctrl_tx_pma_syncp_inv: string  := "false";
        rstctrl_1us_count_fref_clk: string  := "rstctrl_1us_cnt";
        rstctrl_1us_count_fref_clk_value: vl_logic_vector(0 to 19) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1);
        rstctrl_1ms_count_fref_clk: string  := "rstctrl_1ms_cnt";
        rstctrl_1ms_count_fref_clk_value: vl_logic_vector(0 to 19) := (Hi0, Hi0, Hi0, Hi0, Hi1, Hi1, Hi1, Hi1, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi1, Hi0, Hi0);
        rstctrl_off_cal_done_select: string  := "not_active";
        rstctrl_rx_pma_rstb_cmu_select: string  := "not_active";
        rstctrl_rx_pma_rstb_select: string  := "not_active";
        rstctrl_rx_pll_freq_lock_select: string  := "not_active";
        rstctrl_mask_tx_pll_lock_select: string  := "not_active";
        rstctrl_rx_pll_lock_select: string  := "not_active";
        rstctrl_perstn_select: string  := "perstn_pin";
        rstctrl_tx_lc_pll_rstb_select: string  := "not_active";
        rstctrl_fref_clk_select: string  := "ch0_sel";
        rstctrl_off_cal_en_select: string  := "not_active";
        rstctrl_tx_pma_syncp_select: string  := "not_active";
        rstctrl_rx_pcs_rst_n_select: string  := "not_active";
        rstctrl_tx_cmu_pll_lock_select: string  := "not_active";
        rstctrl_tx_pcs_rst_n_select: string  := "not_active";
        rstctrl_tx_lc_pll_lock_select: string  := "not_active";
        rstctrl_timer_a : string  := "rstctrl_timer_a";
        rstctrl_timer_a_type: string  := "milli_secs";
        rstctrl_timer_a_value: vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi1, Hi0);
        rstctrl_timer_b : string  := "rstctrl_timer_b";
        rstctrl_timer_b_type: string  := "milli_secs";
        rstctrl_timer_b_value: vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi1, Hi0);
        rstctrl_timer_c : string  := "rstctrl_timer_c";
        rstctrl_timer_c_type: string  := "milli_secs";
        rstctrl_timer_c_value: vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi1, Hi0);
        rstctrl_timer_d : string  := "rstctrl_timer_d";
        rstctrl_timer_d_type: string  := "milli_secs";
        rstctrl_timer_d_value: vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi1, Hi0, Hi1, Hi0, Hi0);
        rstctrl_timer_e : string  := "rstctrl_timer_e";
        rstctrl_timer_e_type: string  := "milli_secs";
        rstctrl_timer_e_value: vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1);
        rstctrl_timer_f : string  := "rstctrl_timer_f";
        rstctrl_timer_f_type: string  := "milli_secs";
        rstctrl_timer_f_value: vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi1, Hi0);
        rstctrl_timer_g : string  := "rstctrl_timer_g";
        rstctrl_timer_g_type: string  := "milli_secs";
        rstctrl_timer_g_value: vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi1, Hi0);
        rstctrl_timer_h : string  := "rstctrl_timer_h";
        rstctrl_timer_h_type: string  := "milli_secs";
        rstctrl_timer_h_value: vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0);
        rstctrl_timer_i : string  := "rstctrl_timer_i";
        rstctrl_timer_i_type: string  := "milli_secs";
        rstctrl_timer_i_value: vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi1, Hi0, Hi1, Hi0, Hi0);
        rstctrl_timer_j : string  := "rstctrl_timer_j";
        rstctrl_timer_j_type: string  := "milli_secs";
        rstctrl_timer_j_value: vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi1, Hi0, Hi1, Hi0, Hi0);
        rstctrl_ltssm_disable: string  := "false";
        cvp_isolation   : string  := "enable"
    );
    port(
        usermode        : in     vl_logic;
        hippartialreconfign: in     vl_logic;
        csrclk          : in     vl_logic;
        csrin           : in     vl_logic;
        csren           : in     vl_logic;
        csrout          : out    vl_logic;
        csrcbdin        : in     vl_logic;
        csrtcsrin       : in     vl_logic;
        csrdin          : in     vl_logic;
        csrseg          : in     vl_logic;
        csrenscan       : in     vl_logic;
        csrtverify      : in     vl_logic;
        csrloadcsr      : in     vl_logic;
        csrpipein       : in     vl_logic;
        csrdout         : out    vl_logic;
        csrpipeout      : out    vl_logic;
        avmmrstn        : in     vl_logic;
        avmmclk         : in     vl_logic;
        avmmwrite       : in     vl_logic;
        avmmread        : in     vl_logic;
        avmmbyteen      : in     vl_logic_vector(1 downto 0);
        avmmaddress     : in     vl_logic_vector(9 downto 0);
        avmmwritedata   : in     vl_logic_vector(15 downto 0);
        sershiftload    : in     vl_logic;
        interfacesel    : in     vl_logic;
        avmmreaddata    : out    vl_logic_vector(15 downto 0);
        mdioclk         : in     vl_logic;
        mdioin          : in     vl_logic;
        cbhipmdioen     : in     vl_logic;
        mdiodevaddr     : in     vl_logic_vector(1 downto 0);
        mdioout         : out    vl_logic;
        mdiooenn        : out    vl_logic;
        lmidout         : out    vl_logic_vector(31 downto 0);
        lmiack          : out    vl_logic;
        lmirden         : in     vl_logic;
        lmiwren         : in     vl_logic;
        lmiaddr         : in     vl_logic_vector(14 downto 0);
        lmidin          : in     vl_logic_vector(31 downto 0);
        resetstatus     : out    vl_logic;
        l2exit          : out    vl_logic;
        hotrstexit      : out    vl_logic;
        dlupexit        : out    vl_logic;
        pldclk          : in     vl_logic;
        pldsrst         : in     vl_logic;
        pldrst          : in     vl_logic;
        phyrst          : in     vl_logic;
        physrst         : in     vl_logic;
        coreclkin       : in     vl_logic;
        coreclkout      : out    vl_logic;
        corerst         : in     vl_logic;
        corepor         : in     vl_logic;
        corecrst        : in     vl_logic;
        coresrst        : in     vl_logic;
        swdnwake        : out    vl_logic;
        swuphotrst      : out    vl_logic;
        swdnin          : in     vl_logic_vector(2 downto 0);
        swupin          : in     vl_logic_vector(6 downto 0);
        rxvalidvc0      : out    vl_logic;
        rxerrvc0        : out    vl_logic;
        rxbardecvc0     : out    vl_logic_vector(7 downto 0);
        rxsopvc00       : out    vl_logic;
        rxeopvc00       : out    vl_logic;
        rxdatavc00      : out    vl_logic_vector(63 downto 0);
        rxbevc00        : out    vl_logic_vector(7 downto 0);
        rxsopvc01       : out    vl_logic;
        rxeopvc01       : out    vl_logic;
        rxdatavc01      : out    vl_logic_vector(63 downto 0);
        rxbevc01        : out    vl_logic_vector(7 downto 0);
        rxfifofullvc0   : out    vl_logic;
        rxfifoemptyvc0  : out    vl_logic;
        rxfifowrpvc0    : out    vl_logic_vector(3 downto 0);
        rxfifordpvc0    : out    vl_logic_vector(3 downto 0);
        txcredvc0       : out    vl_logic_vector(35 downto 0);
        txreadyvc0      : out    vl_logic;
        txfifofullvc0   : out    vl_logic;
        txfifoemptyvc0  : out    vl_logic;
        txfifowrpvc0    : out    vl_logic_vector(3 downto 0);
        txfifordpvc0    : out    vl_logic_vector(3 downto 0);
        rxmaskvc0       : in     vl_logic;
        rxreadyvc0      : in     vl_logic;
        txvalidvc0      : in     vl_logic;
        txerrvc0        : in     vl_logic;
        txsopvc00       : in     vl_logic;
        txeopvc00       : in     vl_logic;
        txdatavc00      : in     vl_logic_vector(63 downto 0);
        txsopvc01       : in     vl_logic;
        txeopvc01       : in     vl_logic;
        txdatavc01      : in     vl_logic_vector(63 downto 0);
        tlpmetosr       : out    vl_logic;
        tlpmetocr       : in     vl_logic;
        tlpmevent       : in     vl_logic;
        tlpmdata        : in     vl_logic_vector(9 downto 0);
        tlpmauxpwr      : in     vl_logic;
        tlcfgsts        : out    vl_logic_vector(122 downto 0);
        tlcfgstswr      : out    vl_logic;
        tlcfgctl        : out    vl_logic_vector(31 downto 0);
        tlcfgctlwr      : out    vl_logic;
        tlcfgadd        : out    vl_logic_vector(6 downto 0);
        tlappintaack    : out    vl_logic;
        tlappmsiack     : out    vl_logic;
        intstatus       : out    vl_logic_vector(3 downto 0);
        tlappintasts    : in     vl_logic;
        tlappmsireq     : in     vl_logic;
        tlappmsitc      : in     vl_logic_vector(2 downto 0);
        tlappmsinum     : in     vl_logic_vector(4 downto 0);
        tlaermsinum     : in     vl_logic_vector(4 downto 0);
        tlpexmsinum     : in     vl_logic_vector(4 downto 0);
        tlhpgctrler     : in     vl_logic_vector(4 downto 0);
        laneact         : out    vl_logic_vector(3 downto 0);
        dlltssm         : out    vl_logic_vector(4 downto 0);
        clrrxpath       : out    vl_logic;
        dlcurrentspeed  : out    vl_logic_vector(1 downto 0);
        dlcomclkreg     : in     vl_logic;
        dlvcctrl        : in     vl_logic_vector(7 downto 0);
        dlctrllink2     : in     vl_logic_vector(12 downto 0);
        testouthip      : out    vl_logic_vector(63 downto 0);
        ev1us           : out    vl_logic;
        ev128ns         : out    vl_logic;
        wakeoen         : out    vl_logic;
        serrout         : out    vl_logic;
        tlslotclkcfg    : in     vl_logic;
        mode            : in     vl_logic_vector(1 downto 0);
        testinhip       : in     vl_logic_vector(39 downto 0);
        cplerr          : in     vl_logic_vector(6 downto 0);
        pcierr          : in     vl_logic_vector(15 downto 0);
        rate0           : out    vl_logic;
        rate1           : out    vl_logic;
        rate2           : out    vl_logic;
        rate3           : out    vl_logic;
        rate4           : out    vl_logic;
        rate5           : out    vl_logic;
        rate6           : out    vl_logic;
        rate7           : out    vl_logic;
        rate8           : out    vl_logic;
        eidleinfersel0  : out    vl_logic_vector(2 downto 0);
        txdeemph0       : out    vl_logic;
        txmargin0       : out    vl_logic_vector(2 downto 0);
        txdata0         : out    vl_logic_vector(7 downto 0);
        txdatak0        : out    vl_logic;
        txdetectrx0     : out    vl_logic;
        txelecidle0     : out    vl_logic;
        txcompl0        : out    vl_logic;
        rxpolarity0     : out    vl_logic;
        powerdown0      : out    vl_logic_vector(1 downto 0);
        rxdata0         : in     vl_logic_vector(7 downto 0);
        rxdatak0        : in     vl_logic;
        rxvalid0        : in     vl_logic;
        phystatus0      : in     vl_logic;
        rxelecidle0     : in     vl_logic;
        rxstatus0       : in     vl_logic_vector(2 downto 0);
        eidleinfersel1  : out    vl_logic_vector(2 downto 0);
        txdeemph1       : out    vl_logic;
        txmargin1       : out    vl_logic_vector(2 downto 0);
        txdata1         : out    vl_logic_vector(7 downto 0);
        txdatak1        : out    vl_logic;
        txdetectrx1     : out    vl_logic;
        txelecidle1     : out    vl_logic;
        txcompl1        : out    vl_logic;
        rxpolarity1     : out    vl_logic;
        powerdown1      : out    vl_logic_vector(1 downto 0);
        rxdata1         : in     vl_logic_vector(7 downto 0);
        rxdatak1        : in     vl_logic;
        rxvalid1        : in     vl_logic;
        phystatus1      : in     vl_logic;
        rxelecidle1     : in     vl_logic;
        rxstatus1       : in     vl_logic_vector(2 downto 0);
        eidleinfersel2  : out    vl_logic_vector(2 downto 0);
        txdeemph2       : out    vl_logic;
        txmargin2       : out    vl_logic_vector(2 downto 0);
        txdata2         : out    vl_logic_vector(7 downto 0);
        txdatak2        : out    vl_logic;
        txdetectrx2     : out    vl_logic;
        txelecidle2     : out    vl_logic;
        txcompl2        : out    vl_logic;
        rxpolarity2     : out    vl_logic;
        powerdown2      : out    vl_logic_vector(1 downto 0);
        rxdata2         : in     vl_logic_vector(7 downto 0);
        rxdatak2        : in     vl_logic;
        rxvalid2        : in     vl_logic;
        phystatus2      : in     vl_logic;
        rxelecidle2     : in     vl_logic;
        rxstatus2       : in     vl_logic_vector(2 downto 0);
        eidleinfersel3  : out    vl_logic_vector(2 downto 0);
        txdeemph3       : out    vl_logic;
        txmargin3       : out    vl_logic_vector(2 downto 0);
        txdata3         : out    vl_logic_vector(7 downto 0);
        txdatak3        : out    vl_logic;
        txdetectrx3     : out    vl_logic;
        txelecidle3     : out    vl_logic;
        txcompl3        : out    vl_logic;
        rxpolarity3     : out    vl_logic;
        powerdown3      : out    vl_logic_vector(1 downto 0);
        rxdata3         : in     vl_logic_vector(7 downto 0);
        rxdatak3        : in     vl_logic;
        rxvalid3        : in     vl_logic;
        phystatus3      : in     vl_logic;
        rxelecidle3     : in     vl_logic;
        rxstatus3       : in     vl_logic_vector(2 downto 0);
        eidleinfersel4  : out    vl_logic_vector(2 downto 0);
        txdeemph4       : out    vl_logic;
        txmargin4       : out    vl_logic_vector(2 downto 0);
        txdata4         : out    vl_logic_vector(7 downto 0);
        txdatak4        : out    vl_logic;
        txdetectrx4     : out    vl_logic;
        txelecidle4     : out    vl_logic;
        txcompl4        : out    vl_logic;
        rxpolarity4     : out    vl_logic;
        powerdown4      : out    vl_logic_vector(1 downto 0);
        rxdata4         : in     vl_logic_vector(7 downto 0);
        rxdatak4        : in     vl_logic;
        rxvalid4        : in     vl_logic;
        phystatus4      : in     vl_logic;
        rxelecidle4     : in     vl_logic;
        rxstatus4       : in     vl_logic_vector(2 downto 0);
        eidleinfersel5  : out    vl_logic_vector(2 downto 0);
        txdeemph5       : out    vl_logic;
        txmargin5       : out    vl_logic_vector(2 downto 0);
        txdata5         : out    vl_logic_vector(7 downto 0);
        txdatak5        : out    vl_logic;
        txdetectrx5     : out    vl_logic;
        txelecidle5     : out    vl_logic;
        txcompl5        : out    vl_logic;
        rxpolarity5     : out    vl_logic;
        powerdown5      : out    vl_logic_vector(1 downto 0);
        rxdata5         : in     vl_logic_vector(7 downto 0);
        rxdatak5        : in     vl_logic;
        rxvalid5        : in     vl_logic;
        phystatus5      : in     vl_logic;
        rxelecidle5     : in     vl_logic;
        rxstatus5       : in     vl_logic_vector(2 downto 0);
        eidleinfersel6  : out    vl_logic_vector(2 downto 0);
        txdeemph6       : out    vl_logic;
        txmargin6       : out    vl_logic_vector(2 downto 0);
        txdata6         : out    vl_logic_vector(7 downto 0);
        txdatak6        : out    vl_logic;
        txdetectrx6     : out    vl_logic;
        txelecidle6     : out    vl_logic;
        txcompl6        : out    vl_logic;
        rxpolarity6     : out    vl_logic;
        powerdown6      : out    vl_logic_vector(1 downto 0);
        rxdata6         : in     vl_logic_vector(7 downto 0);
        rxdatak6        : in     vl_logic;
        rxvalid6        : in     vl_logic;
        phystatus6      : in     vl_logic;
        rxelecidle6     : in     vl_logic;
        rxstatus6       : in     vl_logic_vector(2 downto 0);
        eidleinfersel7  : out    vl_logic_vector(2 downto 0);
        txdeemph7       : out    vl_logic;
        txmargin7       : out    vl_logic_vector(2 downto 0);
        txdata7         : out    vl_logic_vector(7 downto 0);
        txdatak7        : out    vl_logic;
        txdetectrx7     : out    vl_logic;
        txelecidle7     : out    vl_logic;
        txcompl7        : out    vl_logic;
        rxpolarity7     : out    vl_logic;
        powerdown7      : out    vl_logic_vector(1 downto 0);
        rxdata7         : in     vl_logic_vector(7 downto 0);
        rxdatak7        : in     vl_logic;
        rxvalid7        : in     vl_logic;
        phystatus7      : in     vl_logic;
        rxelecidle7     : in     vl_logic;
        rxstatus7       : in     vl_logic_vector(2 downto 0);
        ltssml0state    : out    vl_logic;
        bisttestenn     : in     vl_logic;
        bistscanin      : in     vl_logic;
        bistscanenn     : in     vl_logic;
        bistenn         : in     vl_logic;
        bistscanoutrpl  : out    vl_logic;
        bistscanoutrcv0 : out    vl_logic;
        bistscanoutrcv1 : out    vl_logic;
        bistdonearpl    : out    vl_logic;
        bistdonebrpl    : out    vl_logic;
        bistpassrpl     : out    vl_logic;
        derrrpl         : out    vl_logic;
        derrcorextrpl   : out    vl_logic;
        bistdonearcv0   : out    vl_logic;
        bistdonebrcv0   : out    vl_logic;
        bistpassrcv0    : out    vl_logic;
        derrcorextrcv0  : out    vl_logic;
        derrcorextrcv1  : out    vl_logic;
        bistdonearcv1   : out    vl_logic;
        bistdonebrcv1   : out    vl_logic;
        bistpassrcv1    : out    vl_logic;
        scanmoden       : in     vl_logic;
        scanenn         : in     vl_logic;
        dpriorefclkdig  : in     vl_logic;
        nfrzdrv         : in     vl_logic;
        frzreg          : in     vl_logic;
        frzlogic        : in     vl_logic;
        pinperstn       : in     vl_logic;
        pldperstn       : in     vl_logic;
        pldclrpmapcshipn: in     vl_logic;
        pldclrpcshipn   : in     vl_logic;
        pldclrhipn      : in     vl_logic;
        iocsrrdydly     : in     vl_logic;
        plniotri        : in     vl_logic;
        entest          : in     vl_logic;
        por             : in     vl_logic;
        frefclk0        : in     vl_logic;
        frefclk1        : in     vl_logic;
        frefclk2        : in     vl_logic;
        frefclk3        : in     vl_logic;
        frefclk4        : in     vl_logic;
        frefclk5        : in     vl_logic;
        frefclk6        : in     vl_logic;
        frefclk7        : in     vl_logic;
        frefclk8        : in     vl_logic;
        rxfreqtxcmuplllock0: in     vl_logic;
        rxfreqtxcmuplllock1: in     vl_logic;
        rxfreqtxcmuplllock2: in     vl_logic;
        rxfreqtxcmuplllock3: in     vl_logic;
        rxfreqtxcmuplllock4: in     vl_logic;
        rxfreqtxcmuplllock5: in     vl_logic;
        rxfreqtxcmuplllock6: in     vl_logic;
        rxfreqtxcmuplllock7: in     vl_logic;
        rxfreqtxcmuplllock8: in     vl_logic;
        rxpllphaselock0 : in     vl_logic;
        rxpllphaselock1 : in     vl_logic;
        rxpllphaselock2 : in     vl_logic;
        rxpllphaselock3 : in     vl_logic;
        rxpllphaselock4 : in     vl_logic;
        rxpllphaselock5 : in     vl_logic;
        rxpllphaselock6 : in     vl_logic;
        rxpllphaselock7 : in     vl_logic;
        rxpllphaselock8 : in     vl_logic;
        txpcsrstn0      : out    vl_logic;
        txpcsrstn1      : out    vl_logic;
        txpcsrstn2      : out    vl_logic;
        txpcsrstn3      : out    vl_logic;
        txpcsrstn4      : out    vl_logic;
        txpcsrstn5      : out    vl_logic;
        txpcsrstn6      : out    vl_logic;
        txpcsrstn7      : out    vl_logic;
        txpcsrstn8      : out    vl_logic;
        rxpcsrstn0      : out    vl_logic;
        rxpcsrstn1      : out    vl_logic;
        rxpcsrstn2      : out    vl_logic;
        rxpcsrstn3      : out    vl_logic;
        rxpcsrstn4      : out    vl_logic;
        rxpcsrstn5      : out    vl_logic;
        rxpcsrstn6      : out    vl_logic;
        rxpcsrstn7      : out    vl_logic;
        rxpcsrstn8      : out    vl_logic;
        txpmasyncp0     : out    vl_logic;
        txpmasyncp1     : out    vl_logic;
        txpmasyncp2     : out    vl_logic;
        txpmasyncp3     : out    vl_logic;
        txpmasyncp4     : out    vl_logic;
        txpmasyncp5     : out    vl_logic;
        txpmasyncp6     : out    vl_logic;
        txpmasyncp7     : out    vl_logic;
        txpmasyncp8     : out    vl_logic;
        rxpmarstb0      : out    vl_logic;
        rxpmarstb1      : out    vl_logic;
        rxpmarstb2      : out    vl_logic;
        rxpmarstb3      : out    vl_logic;
        rxpmarstb4      : out    vl_logic;
        rxpmarstb5      : out    vl_logic;
        rxpmarstb6      : out    vl_logic;
        rxpmarstb7      : out    vl_logic;
        rxpmarstb8      : out    vl_logic;
        rxbardecfuncnumvc0: out    vl_logic_vector(2 downto 0);
        tlpmeventfunc   : in     vl_logic_vector(2 downto 0);
        tlappintafuncnum: in     vl_logic_vector(2 downto 0);
        tlappintbsts    : in     vl_logic;
        tlappintbfuncnum: in     vl_logic_vector(2 downto 0);
        tlappintcsts    : in     vl_logic;
        tlappintcfuncnum: in     vl_logic_vector(2 downto 0);
        tlappintdsts    : in     vl_logic;
        tlappintdfuncnum: in     vl_logic_vector(2 downto 0);
        tlappmsifunc    : in     vl_logic_vector(2 downto 0);
        cplpending      : in     vl_logic_vector(7 downto 0);
        cplerrfunc      : in     vl_logic_vector(2 downto 0);
        flrreset        : in     vl_logic_vector(7 downto 0);
        cvpconfigready  : in     vl_logic;
        cvpen           : in     vl_logic;
        cvpconfigerror  : in     vl_logic;
        cvpconfigdone   : in     vl_logic;
        cvpclk          : out    vl_logic;
        cvpdata         : out    vl_logic_vector(31 downto 0);
        cvpstartxfer    : out    vl_logic;
        cvpconfig       : out    vl_logic;
        cvpfullconfig   : out    vl_logic;
        pclkch0         : in     vl_logic;
        pclkch1         : in     vl_logic;
        pclkcentral     : in     vl_logic;
        pllfixedclkch0  : in     vl_logic;
        pllfixedclkch1  : in     vl_logic;
        pllfixedclkcentral: in     vl_logic;
        tlappintback    : out    vl_logic;
        tlappintcack    : out    vl_logic;
        tlappintdack    : out    vl_logic;
        flrsts          : out    vl_logic_vector(7 downto 0);
        rxfreqlocked0   : in     vl_logic;
        rxfreqlocked1   : in     vl_logic;
        rxfreqlocked2   : in     vl_logic;
        rxfreqlocked3   : in     vl_logic;
        rxfreqlocked4   : in     vl_logic;
        rxfreqlocked5   : in     vl_logic;
        rxfreqlocked6   : in     vl_logic;
        rxfreqlocked7   : in     vl_logic;
        txswing0        : out    vl_logic;
        txswing1        : out    vl_logic;
        txswing2        : out    vl_logic;
        txswing3        : out    vl_logic;
        txswing4        : out    vl_logic;
        txswing5        : out    vl_logic;
        txswing6        : out    vl_logic;
        txswing7        : out    vl_logic;
        txcredfchipcons : out    vl_logic_vector(5 downto 0);
        txcredfcinfinite: out    vl_logic_vector(5 downto 0);
        txcredhdrfcp    : out    vl_logic_vector(7 downto 0);
        txcreddatafcp   : out    vl_logic_vector(11 downto 0);
        txcredhdrfcnp   : out    vl_logic_vector(7 downto 0);
        txcreddatafcnp  : out    vl_logic_vector(11 downto 0);
        txcredhdrfccp   : out    vl_logic_vector(7 downto 0);
        txcreddatafccp  : out    vl_logic_vector(11 downto 0);
        dbgpipex1rx     : in     vl_logic_vector(14 downto 0);
        vcc_hd          : in     vl_logic;
        vss_hd          : in     vl_logic;
        hipextrain      : in     vl_logic_vector(29 downto 0);
        hipextraclkin   : in     vl_logic_vector(1 downto 0);
        r2cerrext       : out    vl_logic;
        successfulspeednegotiationint: out    vl_logic;
        hipextraout     : out    vl_logic_vector(29 downto 0);
        hipextraclkout  : out    vl_logic_vector(1 downto 0);
        pldcoreready    : in     vl_logic;
        pldclkinuse     : out    vl_logic
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of func_mode : constant is 1;
    attribute mti_svvh_generic_type of bonding_mode : constant is 1;
    attribute mti_svvh_generic_type of prot_mode : constant is 1;
    attribute mti_svvh_generic_type of pcie_spec_1p0_compliance : constant is 1;
    attribute mti_svvh_generic_type of vc_enable : constant is 1;
    attribute mti_svvh_generic_type of enable_slot_register : constant is 1;
    attribute mti_svvh_generic_type of pcie_mode : constant is 1;
    attribute mti_svvh_generic_type of multi_function : constant is 1;
    attribute mti_svvh_generic_type of bypass_cdc : constant is 1;
    attribute mti_svvh_generic_type of cdc_clk_relation : constant is 1;
    attribute mti_svvh_generic_type of enable_rx_reordering : constant is 1;
    attribute mti_svvh_generic_type of enable_rx_buffer_checking : constant is 1;
    attribute mti_svvh_generic_type of single_rx_detect_data : constant is 1;
    attribute mti_svvh_generic_type of single_rx_detect : constant is 1;
    attribute mti_svvh_generic_type of use_crc_forwarding : constant is 1;
    attribute mti_svvh_generic_type of bypass_tl : constant is 1;
    attribute mti_svvh_generic_type of gen12_lane_rate_mode : constant is 1;
    attribute mti_svvh_generic_type of lane_mask : constant is 1;
    attribute mti_svvh_generic_type of disable_link_x2_support : constant is 1;
    attribute mti_svvh_generic_type of national_inst_thru_enhance : constant is 1;
    attribute mti_svvh_generic_type of disable_tag_check : constant is 1;
    attribute mti_svvh_generic_type of port_link_number_data : constant is 1;
    attribute mti_svvh_generic_type of port_link_number : constant is 1;
    attribute mti_svvh_generic_type of device_number_data : constant is 1;
    attribute mti_svvh_generic_type of device_number : constant is 1;
    attribute mti_svvh_generic_type of bypass_clk_switch : constant is 1;
    attribute mti_svvh_generic_type of core_clk_out_sel : constant is 1;
    attribute mti_svvh_generic_type of core_clk_divider : constant is 1;
    attribute mti_svvh_generic_type of core_clk_source : constant is 1;
    attribute mti_svvh_generic_type of core_clk_sel : constant is 1;
    attribute mti_svvh_generic_type of disable_clk_switch : constant is 1;
    attribute mti_svvh_generic_type of core_clk_disable_clk_switch : constant is 1;
    attribute mti_svvh_generic_type of slotclk_cfg : constant is 1;
    attribute mti_svvh_generic_type of tx_swing_data : constant is 1;
    attribute mti_svvh_generic_type of tx_swing : constant is 1;
    attribute mti_svvh_generic_type of enable_ch0_pclk_out : constant is 1;
    attribute mti_svvh_generic_type of enable_ch01_pclk_out : constant is 1;
    attribute mti_svvh_generic_type of pipex1_debug_sel : constant is 1;
    attribute mti_svvh_generic_type of pclk_out_sel : constant is 1;
    attribute mti_svvh_generic_type of vendor_id_data_0 : constant is 1;
    attribute mti_svvh_generic_type of vendor_id_0 : constant is 1;
    attribute mti_svvh_generic_type of device_id_data_0 : constant is 1;
    attribute mti_svvh_generic_type of device_id_0 : constant is 1;
    attribute mti_svvh_generic_type of revision_id_data_0 : constant is 1;
    attribute mti_svvh_generic_type of revision_id_0 : constant is 1;
    attribute mti_svvh_generic_type of class_code_data_0 : constant is 1;
    attribute mti_svvh_generic_type of class_code_0 : constant is 1;
    attribute mti_svvh_generic_type of subsystem_vendor_id_data_0 : constant is 1;
    attribute mti_svvh_generic_type of subsystem_vendor_id_0 : constant is 1;
    attribute mti_svvh_generic_type of subsystem_device_id_data_0 : constant is 1;
    attribute mti_svvh_generic_type of subsystem_device_id_0 : constant is 1;
    attribute mti_svvh_generic_type of no_soft_reset_0 : constant is 1;
    attribute mti_svvh_generic_type of intel_id_access_0 : constant is 1;
    attribute mti_svvh_generic_type of device_specific_init_0 : constant is 1;
    attribute mti_svvh_generic_type of maximum_current_data_0 : constant is 1;
    attribute mti_svvh_generic_type of maximum_current_0 : constant is 1;
    attribute mti_svvh_generic_type of d1_support_0 : constant is 1;
    attribute mti_svvh_generic_type of d2_support_0 : constant is 1;
    attribute mti_svvh_generic_type of d0_pme_0 : constant is 1;
    attribute mti_svvh_generic_type of d1_pme_0 : constant is 1;
    attribute mti_svvh_generic_type of d2_pme_0 : constant is 1;
    attribute mti_svvh_generic_type of d3_hot_pme_0 : constant is 1;
    attribute mti_svvh_generic_type of d3_cold_pme_0 : constant is 1;
    attribute mti_svvh_generic_type of use_aer_0 : constant is 1;
    attribute mti_svvh_generic_type of low_priority_vc_0 : constant is 1;
    attribute mti_svvh_generic_type of vc_arbitration_0 : constant is 1;
    attribute mti_svvh_generic_type of disable_snoop_packet_0 : constant is 1;
    attribute mti_svvh_generic_type of max_payload_size_0 : constant is 1;
    attribute mti_svvh_generic_type of surprise_down_error_support_0 : constant is 1;
    attribute mti_svvh_generic_type of dll_active_report_support_0 : constant is 1;
    attribute mti_svvh_generic_type of extend_tag_field_0 : constant is 1;
    attribute mti_svvh_generic_type of endpoint_l0_latency_data_0 : constant is 1;
    attribute mti_svvh_generic_type of endpoint_l0_latency_0 : constant is 1;
    attribute mti_svvh_generic_type of endpoint_l1_latency_data_0 : constant is 1;
    attribute mti_svvh_generic_type of endpoint_l1_latency_0 : constant is 1;
    attribute mti_svvh_generic_type of indicator_data_0 : constant is 1;
    attribute mti_svvh_generic_type of indicator_0 : constant is 1;
    attribute mti_svvh_generic_type of role_based_error_reporting_0 : constant is 1;
    attribute mti_svvh_generic_type of slot_power_scale_data_0 : constant is 1;
    attribute mti_svvh_generic_type of slot_power_scale_0 : constant is 1;
    attribute mti_svvh_generic_type of max_link_width_0 : constant is 1;
    attribute mti_svvh_generic_type of enable_l1_aspm_0 : constant is 1;
    attribute mti_svvh_generic_type of enable_l0s_aspm_0 : constant is 1;
    attribute mti_svvh_generic_type of l1_exit_latency_sameclock_data_0 : constant is 1;
    attribute mti_svvh_generic_type of l1_exit_latency_sameclock_0 : constant is 1;
    attribute mti_svvh_generic_type of l1_exit_latency_diffclock_data_0 : constant is 1;
    attribute mti_svvh_generic_type of l1_exit_latency_diffclock_0 : constant is 1;
    attribute mti_svvh_generic_type of hot_plug_support_data_0 : constant is 1;
    attribute mti_svvh_generic_type of hot_plug_support_0 : constant is 1;
    attribute mti_svvh_generic_type of slot_power_limit_data_0 : constant is 1;
    attribute mti_svvh_generic_type of slot_power_limit_0 : constant is 1;
    attribute mti_svvh_generic_type of slot_number_data_0 : constant is 1;
    attribute mti_svvh_generic_type of slot_number_0 : constant is 1;
    attribute mti_svvh_generic_type of diffclock_nfts_count_data_0 : constant is 1;
    attribute mti_svvh_generic_type of diffclock_nfts_count_0 : constant is 1;
    attribute mti_svvh_generic_type of sameclock_nfts_count_data_0 : constant is 1;
    attribute mti_svvh_generic_type of sameclock_nfts_count_0 : constant is 1;
    attribute mti_svvh_generic_type of completion_timeout_0 : constant is 1;
    attribute mti_svvh_generic_type of enable_completion_timeout_disable_0 : constant is 1;
    attribute mti_svvh_generic_type of extended_tag_reset_0 : constant is 1;
    attribute mti_svvh_generic_type of ecrc_check_capable_0 : constant is 1;
    attribute mti_svvh_generic_type of ecrc_gen_capable_0 : constant is 1;
    attribute mti_svvh_generic_type of no_command_completed_0 : constant is 1;
    attribute mti_svvh_generic_type of msi_multi_message_capable_0 : constant is 1;
    attribute mti_svvh_generic_type of msi_64bit_addressing_capable_0 : constant is 1;
    attribute mti_svvh_generic_type of msi_masking_capable_0 : constant is 1;
    attribute mti_svvh_generic_type of msi_support_0 : constant is 1;
    attribute mti_svvh_generic_type of interrupt_pin_0 : constant is 1;
    attribute mti_svvh_generic_type of enable_function_msix_support_0 : constant is 1;
    attribute mti_svvh_generic_type of msix_table_size_data_0 : constant is 1;
    attribute mti_svvh_generic_type of msix_table_size_0 : constant is 1;
    attribute mti_svvh_generic_type of msix_table_bir_data_0 : constant is 1;
    attribute mti_svvh_generic_type of msix_table_bir_0 : constant is 1;
    attribute mti_svvh_generic_type of msix_table_offset_data_0 : constant is 1;
    attribute mti_svvh_generic_type of msix_table_offset_0 : constant is 1;
    attribute mti_svvh_generic_type of msix_pba_bir_data_0 : constant is 1;
    attribute mti_svvh_generic_type of msix_pba_bir_0 : constant is 1;
    attribute mti_svvh_generic_type of msix_pba_offset_data_0 : constant is 1;
    attribute mti_svvh_generic_type of msix_pba_offset_0 : constant is 1;
    attribute mti_svvh_generic_type of bridge_port_vga_enable_0 : constant is 1;
    attribute mti_svvh_generic_type of bridge_port_ssid_support_0 : constant is 1;
    attribute mti_svvh_generic_type of ssvid_data_0 : constant is 1;
    attribute mti_svvh_generic_type of ssvid_0 : constant is 1;
    attribute mti_svvh_generic_type of ssid_data_0 : constant is 1;
    attribute mti_svvh_generic_type of ssid_0 : constant is 1;
    attribute mti_svvh_generic_type of eie_before_nfts_count_data_0 : constant is 1;
    attribute mti_svvh_generic_type of eie_before_nfts_count_0 : constant is 1;
    attribute mti_svvh_generic_type of gen2_diffclock_nfts_count_data_0 : constant is 1;
    attribute mti_svvh_generic_type of gen2_diffclock_nfts_count_0 : constant is 1;
    attribute mti_svvh_generic_type of gen2_sameclock_nfts_count_data_0 : constant is 1;
    attribute mti_svvh_generic_type of gen2_sameclock_nfts_count_0 : constant is 1;
    attribute mti_svvh_generic_type of deemphasis_enable_0 : constant is 1;
    attribute mti_svvh_generic_type of pcie_spec_version_0 : constant is 1;
    attribute mti_svvh_generic_type of l0_exit_latency_sameclock_data_0 : constant is 1;
    attribute mti_svvh_generic_type of l0_exit_latency_sameclock_0 : constant is 1;
    attribute mti_svvh_generic_type of l0_exit_latency_diffclock_data_0 : constant is 1;
    attribute mti_svvh_generic_type of l0_exit_latency_diffclock_0 : constant is 1;
    attribute mti_svvh_generic_type of rx_ei_l0s_0 : constant is 1;
    attribute mti_svvh_generic_type of l2_async_logic_0 : constant is 1;
    attribute mti_svvh_generic_type of aspm_optionality_0 : constant is 1;
    attribute mti_svvh_generic_type of flr_capability_0 : constant is 1;
    attribute mti_svvh_generic_type of bar0_io_space_0 : constant is 1;
    attribute mti_svvh_generic_type of bar0_64bit_mem_space_0 : constant is 1;
    attribute mti_svvh_generic_type of bar0_prefetchable_0 : constant is 1;
    attribute mti_svvh_generic_type of bar0_size_mask_data_0 : constant is 1;
    attribute mti_svvh_generic_type of bar0_size_mask_0 : constant is 1;
    attribute mti_svvh_generic_type of bar1_io_space_0 : constant is 1;
    attribute mti_svvh_generic_type of bar1_64bit_mem_space_0 : constant is 1;
    attribute mti_svvh_generic_type of bar1_prefetchable_0 : constant is 1;
    attribute mti_svvh_generic_type of bar1_size_mask_data_0 : constant is 1;
    attribute mti_svvh_generic_type of bar1_size_mask_0 : constant is 1;
    attribute mti_svvh_generic_type of bar2_io_space_0 : constant is 1;
    attribute mti_svvh_generic_type of bar2_64bit_mem_space_0 : constant is 1;
    attribute mti_svvh_generic_type of bar2_prefetchable_0 : constant is 1;
    attribute mti_svvh_generic_type of bar2_size_mask_data_0 : constant is 1;
    attribute mti_svvh_generic_type of bar2_size_mask_0 : constant is 1;
    attribute mti_svvh_generic_type of bar3_io_space_0 : constant is 1;
    attribute mti_svvh_generic_type of bar3_64bit_mem_space_0 : constant is 1;
    attribute mti_svvh_generic_type of bar3_prefetchable_0 : constant is 1;
    attribute mti_svvh_generic_type of bar3_size_mask_data_0 : constant is 1;
    attribute mti_svvh_generic_type of bar3_size_mask_0 : constant is 1;
    attribute mti_svvh_generic_type of bar4_io_space_0 : constant is 1;
    attribute mti_svvh_generic_type of bar4_64bit_mem_space_0 : constant is 1;
    attribute mti_svvh_generic_type of bar4_prefetchable_0 : constant is 1;
    attribute mti_svvh_generic_type of bar4_size_mask_data_0 : constant is 1;
    attribute mti_svvh_generic_type of bar4_size_mask_0 : constant is 1;
    attribute mti_svvh_generic_type of bar5_io_space_0 : constant is 1;
    attribute mti_svvh_generic_type of bar5_64bit_mem_space_0 : constant is 1;
    attribute mti_svvh_generic_type of bar5_prefetchable_0 : constant is 1;
    attribute mti_svvh_generic_type of bar5_size_mask_data_0 : constant is 1;
    attribute mti_svvh_generic_type of bar5_size_mask_0 : constant is 1;
    attribute mti_svvh_generic_type of expansion_base_address_register_data_0 : constant is 1;
    attribute mti_svvh_generic_type of expansion_base_address_register_0 : constant is 1;
    attribute mti_svvh_generic_type of io_window_addr_width_0 : constant is 1;
    attribute mti_svvh_generic_type of prefetchable_mem_window_addr_width_0 : constant is 1;
    attribute mti_svvh_generic_type of vendor_id_data_1 : constant is 1;
    attribute mti_svvh_generic_type of vendor_id_1 : constant is 1;
    attribute mti_svvh_generic_type of device_id_data_1 : constant is 1;
    attribute mti_svvh_generic_type of device_id_1 : constant is 1;
    attribute mti_svvh_generic_type of revision_id_data_1 : constant is 1;
    attribute mti_svvh_generic_type of revision_id_1 : constant is 1;
    attribute mti_svvh_generic_type of class_code_data_1 : constant is 1;
    attribute mti_svvh_generic_type of class_code_1 : constant is 1;
    attribute mti_svvh_generic_type of subsystem_vendor_id_data_1 : constant is 1;
    attribute mti_svvh_generic_type of subsystem_vendor_id_1 : constant is 1;
    attribute mti_svvh_generic_type of subsystem_device_id_data_1 : constant is 1;
    attribute mti_svvh_generic_type of subsystem_device_id_1 : constant is 1;
    attribute mti_svvh_generic_type of no_soft_reset_1 : constant is 1;
    attribute mti_svvh_generic_type of intel_id_access_1 : constant is 1;
    attribute mti_svvh_generic_type of device_specific_init_1 : constant is 1;
    attribute mti_svvh_generic_type of maximum_current_data_1 : constant is 1;
    attribute mti_svvh_generic_type of maximum_current_1 : constant is 1;
    attribute mti_svvh_generic_type of d1_support_1 : constant is 1;
    attribute mti_svvh_generic_type of d2_support_1 : constant is 1;
    attribute mti_svvh_generic_type of d0_pme_1 : constant is 1;
    attribute mti_svvh_generic_type of d1_pme_1 : constant is 1;
    attribute mti_svvh_generic_type of d2_pme_1 : constant is 1;
    attribute mti_svvh_generic_type of d3_hot_pme_1 : constant is 1;
    attribute mti_svvh_generic_type of d3_cold_pme_1 : constant is 1;
    attribute mti_svvh_generic_type of use_aer_1 : constant is 1;
    attribute mti_svvh_generic_type of low_priority_vc_1 : constant is 1;
    attribute mti_svvh_generic_type of vc_arbitration_1 : constant is 1;
    attribute mti_svvh_generic_type of disable_snoop_packet_1 : constant is 1;
    attribute mti_svvh_generic_type of max_payload_size_1 : constant is 1;
    attribute mti_svvh_generic_type of surprise_down_error_support_1 : constant is 1;
    attribute mti_svvh_generic_type of dll_active_report_support_1 : constant is 1;
    attribute mti_svvh_generic_type of extend_tag_field_1 : constant is 1;
    attribute mti_svvh_generic_type of endpoint_l0_latency_data_1 : constant is 1;
    attribute mti_svvh_generic_type of endpoint_l0_latency_1 : constant is 1;
    attribute mti_svvh_generic_type of endpoint_l1_latency_data_1 : constant is 1;
    attribute mti_svvh_generic_type of endpoint_l1_latency_1 : constant is 1;
    attribute mti_svvh_generic_type of indicator_data_1 : constant is 1;
    attribute mti_svvh_generic_type of indicator_1 : constant is 1;
    attribute mti_svvh_generic_type of role_based_error_reporting_1 : constant is 1;
    attribute mti_svvh_generic_type of slot_power_scale_data_1 : constant is 1;
    attribute mti_svvh_generic_type of slot_power_scale_1 : constant is 1;
    attribute mti_svvh_generic_type of max_link_width_1 : constant is 1;
    attribute mti_svvh_generic_type of enable_l1_aspm_1 : constant is 1;
    attribute mti_svvh_generic_type of enable_l0s_aspm_1 : constant is 1;
    attribute mti_svvh_generic_type of l1_exit_latency_sameclock_data_1 : constant is 1;
    attribute mti_svvh_generic_type of l1_exit_latency_sameclock_1 : constant is 1;
    attribute mti_svvh_generic_type of l1_exit_latency_diffclock_data_1 : constant is 1;
    attribute mti_svvh_generic_type of l1_exit_latency_diffclock_1 : constant is 1;
    attribute mti_svvh_generic_type of hot_plug_support_data_1 : constant is 1;
    attribute mti_svvh_generic_type of hot_plug_support_1 : constant is 1;
    attribute mti_svvh_generic_type of slot_power_limit_data_1 : constant is 1;
    attribute mti_svvh_generic_type of slot_power_limit_1 : constant is 1;
    attribute mti_svvh_generic_type of slot_number_data_1 : constant is 1;
    attribute mti_svvh_generic_type of slot_number_1 : constant is 1;
    attribute mti_svvh_generic_type of diffclock_nfts_count_data_1 : constant is 1;
    attribute mti_svvh_generic_type of diffclock_nfts_count_1 : constant is 1;
    attribute mti_svvh_generic_type of sameclock_nfts_count_data_1 : constant is 1;
    attribute mti_svvh_generic_type of sameclock_nfts_count_1 : constant is 1;
    attribute mti_svvh_generic_type of completion_timeout_1 : constant is 1;
    attribute mti_svvh_generic_type of enable_completion_timeout_disable_1 : constant is 1;
    attribute mti_svvh_generic_type of extended_tag_reset_1 : constant is 1;
    attribute mti_svvh_generic_type of ecrc_check_capable_1 : constant is 1;
    attribute mti_svvh_generic_type of ecrc_gen_capable_1 : constant is 1;
    attribute mti_svvh_generic_type of no_command_completed_1 : constant is 1;
    attribute mti_svvh_generic_type of msi_multi_message_capable_1 : constant is 1;
    attribute mti_svvh_generic_type of msi_64bit_addressing_capable_1 : constant is 1;
    attribute mti_svvh_generic_type of msi_masking_capable_1 : constant is 1;
    attribute mti_svvh_generic_type of msi_support_1 : constant is 1;
    attribute mti_svvh_generic_type of interrupt_pin_1 : constant is 1;
    attribute mti_svvh_generic_type of enable_function_msix_support_1 : constant is 1;
    attribute mti_svvh_generic_type of msix_table_size_data_1 : constant is 1;
    attribute mti_svvh_generic_type of msix_table_size_1 : constant is 1;
    attribute mti_svvh_generic_type of msix_table_bir_data_1 : constant is 1;
    attribute mti_svvh_generic_type of msix_table_bir_1 : constant is 1;
    attribute mti_svvh_generic_type of msix_table_offset_data_1 : constant is 1;
    attribute mti_svvh_generic_type of msix_table_offset_1 : constant is 1;
    attribute mti_svvh_generic_type of msix_pba_bir_data_1 : constant is 1;
    attribute mti_svvh_generic_type of msix_pba_bir_1 : constant is 1;
    attribute mti_svvh_generic_type of msix_pba_offset_data_1 : constant is 1;
    attribute mti_svvh_generic_type of msix_pba_offset_1 : constant is 1;
    attribute mti_svvh_generic_type of bridge_port_vga_enable_1 : constant is 1;
    attribute mti_svvh_generic_type of bridge_port_ssid_support_1 : constant is 1;
    attribute mti_svvh_generic_type of ssvid_data_1 : constant is 1;
    attribute mti_svvh_generic_type of ssvid_1 : constant is 1;
    attribute mti_svvh_generic_type of ssid_data_1 : constant is 1;
    attribute mti_svvh_generic_type of ssid_1 : constant is 1;
    attribute mti_svvh_generic_type of eie_before_nfts_count_data_1 : constant is 1;
    attribute mti_svvh_generic_type of eie_before_nfts_count_1 : constant is 1;
    attribute mti_svvh_generic_type of gen2_diffclock_nfts_count_data_1 : constant is 1;
    attribute mti_svvh_generic_type of gen2_diffclock_nfts_count_1 : constant is 1;
    attribute mti_svvh_generic_type of gen2_sameclock_nfts_count_data_1 : constant is 1;
    attribute mti_svvh_generic_type of gen2_sameclock_nfts_count_1 : constant is 1;
    attribute mti_svvh_generic_type of deemphasis_enable_1 : constant is 1;
    attribute mti_svvh_generic_type of pcie_spec_version_1 : constant is 1;
    attribute mti_svvh_generic_type of l0_exit_latency_sameclock_data_1 : constant is 1;
    attribute mti_svvh_generic_type of l0_exit_latency_sameclock_1 : constant is 1;
    attribute mti_svvh_generic_type of l0_exit_latency_diffclock_data_1 : constant is 1;
    attribute mti_svvh_generic_type of l0_exit_latency_diffclock_1 : constant is 1;
    attribute mti_svvh_generic_type of rx_ei_l0s_1 : constant is 1;
    attribute mti_svvh_generic_type of l2_async_logic_1 : constant is 1;
    attribute mti_svvh_generic_type of aspm_optionality_1 : constant is 1;
    attribute mti_svvh_generic_type of flr_capability_1 : constant is 1;
    attribute mti_svvh_generic_type of bar0_io_space_1 : constant is 1;
    attribute mti_svvh_generic_type of bar0_64bit_mem_space_1 : constant is 1;
    attribute mti_svvh_generic_type of bar0_prefetchable_1 : constant is 1;
    attribute mti_svvh_generic_type of bar0_size_mask_data_1 : constant is 1;
    attribute mti_svvh_generic_type of bar0_size_mask_1 : constant is 1;
    attribute mti_svvh_generic_type of bar1_io_space_1 : constant is 1;
    attribute mti_svvh_generic_type of bar1_64bit_mem_space_1 : constant is 1;
    attribute mti_svvh_generic_type of bar1_prefetchable_1 : constant is 1;
    attribute mti_svvh_generic_type of bar1_size_mask_data_1 : constant is 1;
    attribute mti_svvh_generic_type of bar1_size_mask_1 : constant is 1;
    attribute mti_svvh_generic_type of bar2_io_space_1 : constant is 1;
    attribute mti_svvh_generic_type of bar2_64bit_mem_space_1 : constant is 1;
    attribute mti_svvh_generic_type of bar2_prefetchable_1 : constant is 1;
    attribute mti_svvh_generic_type of bar2_size_mask_data_1 : constant is 1;
    attribute mti_svvh_generic_type of bar2_size_mask_1 : constant is 1;
    attribute mti_svvh_generic_type of bar3_io_space_1 : constant is 1;
    attribute mti_svvh_generic_type of bar3_64bit_mem_space_1 : constant is 1;
    attribute mti_svvh_generic_type of bar3_prefetchable_1 : constant is 1;
    attribute mti_svvh_generic_type of bar3_size_mask_data_1 : constant is 1;
    attribute mti_svvh_generic_type of bar3_size_mask_1 : constant is 1;
    attribute mti_svvh_generic_type of bar4_io_space_1 : constant is 1;
    attribute mti_svvh_generic_type of bar4_64bit_mem_space_1 : constant is 1;
    attribute mti_svvh_generic_type of bar4_prefetchable_1 : constant is 1;
    attribute mti_svvh_generic_type of bar4_size_mask_data_1 : constant is 1;
    attribute mti_svvh_generic_type of bar4_size_mask_1 : constant is 1;
    attribute mti_svvh_generic_type of bar5_io_space_1 : constant is 1;
    attribute mti_svvh_generic_type of bar5_64bit_mem_space_1 : constant is 1;
    attribute mti_svvh_generic_type of bar5_prefetchable_1 : constant is 1;
    attribute mti_svvh_generic_type of bar5_size_mask_data_1 : constant is 1;
    attribute mti_svvh_generic_type of bar5_size_mask_1 : constant is 1;
    attribute mti_svvh_generic_type of expansion_base_address_register_data_1 : constant is 1;
    attribute mti_svvh_generic_type of expansion_base_address_register_1 : constant is 1;
    attribute mti_svvh_generic_type of io_window_addr_width_1 : constant is 1;
    attribute mti_svvh_generic_type of prefetchable_mem_window_addr_width_1 : constant is 1;
    attribute mti_svvh_generic_type of vendor_id_data_2 : constant is 1;
    attribute mti_svvh_generic_type of vendor_id_2 : constant is 1;
    attribute mti_svvh_generic_type of device_id_data_2 : constant is 1;
    attribute mti_svvh_generic_type of device_id_2 : constant is 1;
    attribute mti_svvh_generic_type of revision_id_data_2 : constant is 1;
    attribute mti_svvh_generic_type of revision_id_2 : constant is 1;
    attribute mti_svvh_generic_type of class_code_data_2 : constant is 1;
    attribute mti_svvh_generic_type of class_code_2 : constant is 1;
    attribute mti_svvh_generic_type of subsystem_vendor_id_data_2 : constant is 1;
    attribute mti_svvh_generic_type of subsystem_vendor_id_2 : constant is 1;
    attribute mti_svvh_generic_type of subsystem_device_id_data_2 : constant is 1;
    attribute mti_svvh_generic_type of subsystem_device_id_2 : constant is 1;
    attribute mti_svvh_generic_type of no_soft_reset_2 : constant is 1;
    attribute mti_svvh_generic_type of intel_id_access_2 : constant is 1;
    attribute mti_svvh_generic_type of device_specific_init_2 : constant is 1;
    attribute mti_svvh_generic_type of maximum_current_data_2 : constant is 1;
    attribute mti_svvh_generic_type of maximum_current_2 : constant is 1;
    attribute mti_svvh_generic_type of d1_support_2 : constant is 1;
    attribute mti_svvh_generic_type of d2_support_2 : constant is 1;
    attribute mti_svvh_generic_type of d0_pme_2 : constant is 1;
    attribute mti_svvh_generic_type of d1_pme_2 : constant is 1;
    attribute mti_svvh_generic_type of d2_pme_2 : constant is 1;
    attribute mti_svvh_generic_type of d3_hot_pme_2 : constant is 1;
    attribute mti_svvh_generic_type of d3_cold_pme_2 : constant is 1;
    attribute mti_svvh_generic_type of use_aer_2 : constant is 1;
    attribute mti_svvh_generic_type of low_priority_vc_2 : constant is 1;
    attribute mti_svvh_generic_type of vc_arbitration_2 : constant is 1;
    attribute mti_svvh_generic_type of disable_snoop_packet_2 : constant is 1;
    attribute mti_svvh_generic_type of max_payload_size_2 : constant is 1;
    attribute mti_svvh_generic_type of surprise_down_error_support_2 : constant is 1;
    attribute mti_svvh_generic_type of dll_active_report_support_2 : constant is 1;
    attribute mti_svvh_generic_type of extend_tag_field_2 : constant is 1;
    attribute mti_svvh_generic_type of endpoint_l0_latency_data_2 : constant is 1;
    attribute mti_svvh_generic_type of endpoint_l0_latency_2 : constant is 1;
    attribute mti_svvh_generic_type of endpoint_l1_latency_data_2 : constant is 1;
    attribute mti_svvh_generic_type of endpoint_l1_latency_2 : constant is 1;
    attribute mti_svvh_generic_type of indicator_data_2 : constant is 1;
    attribute mti_svvh_generic_type of indicator_2 : constant is 1;
    attribute mti_svvh_generic_type of role_based_error_reporting_2 : constant is 1;
    attribute mti_svvh_generic_type of slot_power_scale_data_2 : constant is 1;
    attribute mti_svvh_generic_type of slot_power_scale_2 : constant is 1;
    attribute mti_svvh_generic_type of max_link_width_2 : constant is 1;
    attribute mti_svvh_generic_type of enable_l1_aspm_2 : constant is 1;
    attribute mti_svvh_generic_type of enable_l0s_aspm_2 : constant is 1;
    attribute mti_svvh_generic_type of l1_exit_latency_sameclock_data_2 : constant is 1;
    attribute mti_svvh_generic_type of l1_exit_latency_sameclock_2 : constant is 1;
    attribute mti_svvh_generic_type of l1_exit_latency_diffclock_data_2 : constant is 1;
    attribute mti_svvh_generic_type of l1_exit_latency_diffclock_2 : constant is 1;
    attribute mti_svvh_generic_type of hot_plug_support_data_2 : constant is 1;
    attribute mti_svvh_generic_type of hot_plug_support_2 : constant is 1;
    attribute mti_svvh_generic_type of slot_power_limit_data_2 : constant is 1;
    attribute mti_svvh_generic_type of slot_power_limit_2 : constant is 1;
    attribute mti_svvh_generic_type of slot_number_data_2 : constant is 1;
    attribute mti_svvh_generic_type of slot_number_2 : constant is 1;
    attribute mti_svvh_generic_type of diffclock_nfts_count_data_2 : constant is 1;
    attribute mti_svvh_generic_type of diffclock_nfts_count_2 : constant is 1;
    attribute mti_svvh_generic_type of sameclock_nfts_count_data_2 : constant is 1;
    attribute mti_svvh_generic_type of sameclock_nfts_count_2 : constant is 1;
    attribute mti_svvh_generic_type of completion_timeout_2 : constant is 1;
    attribute mti_svvh_generic_type of enable_completion_timeout_disable_2 : constant is 1;
    attribute mti_svvh_generic_type of extended_tag_reset_2 : constant is 1;
    attribute mti_svvh_generic_type of ecrc_check_capable_2 : constant is 1;
    attribute mti_svvh_generic_type of ecrc_gen_capable_2 : constant is 1;
    attribute mti_svvh_generic_type of no_command_completed_2 : constant is 1;
    attribute mti_svvh_generic_type of msi_multi_message_capable_2 : constant is 1;
    attribute mti_svvh_generic_type of msi_64bit_addressing_capable_2 : constant is 1;
    attribute mti_svvh_generic_type of msi_masking_capable_2 : constant is 1;
    attribute mti_svvh_generic_type of msi_support_2 : constant is 1;
    attribute mti_svvh_generic_type of interrupt_pin_2 : constant is 1;
    attribute mti_svvh_generic_type of enable_function_msix_support_2 : constant is 1;
    attribute mti_svvh_generic_type of msix_table_size_data_2 : constant is 1;
    attribute mti_svvh_generic_type of msix_table_size_2 : constant is 1;
    attribute mti_svvh_generic_type of msix_table_bir_data_2 : constant is 1;
    attribute mti_svvh_generic_type of msix_table_bir_2 : constant is 1;
    attribute mti_svvh_generic_type of msix_table_offset_data_2 : constant is 1;
    attribute mti_svvh_generic_type of msix_table_offset_2 : constant is 1;
    attribute mti_svvh_generic_type of msix_pba_bir_data_2 : constant is 1;
    attribute mti_svvh_generic_type of msix_pba_bir_2 : constant is 1;
    attribute mti_svvh_generic_type of msix_pba_offset_data_2 : constant is 1;
    attribute mti_svvh_generic_type of msix_pba_offset_2 : constant is 1;
    attribute mti_svvh_generic_type of bridge_port_vga_enable_2 : constant is 1;
    attribute mti_svvh_generic_type of bridge_port_ssid_support_2 : constant is 1;
    attribute mti_svvh_generic_type of ssvid_data_2 : constant is 1;
    attribute mti_svvh_generic_type of ssvid_2 : constant is 1;
    attribute mti_svvh_generic_type of ssid_data_2 : constant is 1;
    attribute mti_svvh_generic_type of ssid_2 : constant is 1;
    attribute mti_svvh_generic_type of eie_before_nfts_count_data_2 : constant is 1;
    attribute mti_svvh_generic_type of eie_before_nfts_count_2 : constant is 1;
    attribute mti_svvh_generic_type of gen2_diffclock_nfts_count_data_2 : constant is 1;
    attribute mti_svvh_generic_type of gen2_diffclock_nfts_count_2 : constant is 1;
    attribute mti_svvh_generic_type of gen2_sameclock_nfts_count_data_2 : constant is 1;
    attribute mti_svvh_generic_type of gen2_sameclock_nfts_count_2 : constant is 1;
    attribute mti_svvh_generic_type of deemphasis_enable_2 : constant is 1;
    attribute mti_svvh_generic_type of pcie_spec_version_2 : constant is 1;
    attribute mti_svvh_generic_type of l0_exit_latency_sameclock_data_2 : constant is 1;
    attribute mti_svvh_generic_type of l0_exit_latency_sameclock_2 : constant is 1;
    attribute mti_svvh_generic_type of l0_exit_latency_diffclock_data_2 : constant is 1;
    attribute mti_svvh_generic_type of l0_exit_latency_diffclock_2 : constant is 1;
    attribute mti_svvh_generic_type of rx_ei_l0s_2 : constant is 1;
    attribute mti_svvh_generic_type of l2_async_logic_2 : constant is 1;
    attribute mti_svvh_generic_type of aspm_optionality_2 : constant is 1;
    attribute mti_svvh_generic_type of flr_capability_2 : constant is 1;
    attribute mti_svvh_generic_type of bar0_io_space_2 : constant is 1;
    attribute mti_svvh_generic_type of bar0_64bit_mem_space_2 : constant is 1;
    attribute mti_svvh_generic_type of bar0_prefetchable_2 : constant is 1;
    attribute mti_svvh_generic_type of bar0_size_mask_data_2 : constant is 1;
    attribute mti_svvh_generic_type of bar0_size_mask_2 : constant is 1;
    attribute mti_svvh_generic_type of bar1_io_space_2 : constant is 1;
    attribute mti_svvh_generic_type of bar1_64bit_mem_space_2 : constant is 1;
    attribute mti_svvh_generic_type of bar1_prefetchable_2 : constant is 1;
    attribute mti_svvh_generic_type of bar1_size_mask_data_2 : constant is 1;
    attribute mti_svvh_generic_type of bar1_size_mask_2 : constant is 1;
    attribute mti_svvh_generic_type of bar2_io_space_2 : constant is 1;
    attribute mti_svvh_generic_type of bar2_64bit_mem_space_2 : constant is 1;
    attribute mti_svvh_generic_type of bar2_prefetchable_2 : constant is 1;
    attribute mti_svvh_generic_type of bar2_size_mask_data_2 : constant is 1;
    attribute mti_svvh_generic_type of bar2_size_mask_2 : constant is 1;
    attribute mti_svvh_generic_type of bar3_io_space_2 : constant is 1;
    attribute mti_svvh_generic_type of bar3_64bit_mem_space_2 : constant is 1;
    attribute mti_svvh_generic_type of bar3_prefetchable_2 : constant is 1;
    attribute mti_svvh_generic_type of bar3_size_mask_data_2 : constant is 1;
    attribute mti_svvh_generic_type of bar3_size_mask_2 : constant is 1;
    attribute mti_svvh_generic_type of bar4_io_space_2 : constant is 1;
    attribute mti_svvh_generic_type of bar4_64bit_mem_space_2 : constant is 1;
    attribute mti_svvh_generic_type of bar4_prefetchable_2 : constant is 1;
    attribute mti_svvh_generic_type of bar4_size_mask_data_2 : constant is 1;
    attribute mti_svvh_generic_type of bar4_size_mask_2 : constant is 1;
    attribute mti_svvh_generic_type of bar5_io_space_2 : constant is 1;
    attribute mti_svvh_generic_type of bar5_64bit_mem_space_2 : constant is 1;
    attribute mti_svvh_generic_type of bar5_prefetchable_2 : constant is 1;
    attribute mti_svvh_generic_type of bar5_size_mask_data_2 : constant is 1;
    attribute mti_svvh_generic_type of bar5_size_mask_2 : constant is 1;
    attribute mti_svvh_generic_type of expansion_base_address_register_data_2 : constant is 1;
    attribute mti_svvh_generic_type of expansion_base_address_register_2 : constant is 1;
    attribute mti_svvh_generic_type of io_window_addr_width_2 : constant is 1;
    attribute mti_svvh_generic_type of prefetchable_mem_window_addr_width_2 : constant is 1;
    attribute mti_svvh_generic_type of vendor_id_data_3 : constant is 1;
    attribute mti_svvh_generic_type of vendor_id_3 : constant is 1;
    attribute mti_svvh_generic_type of device_id_data_3 : constant is 1;
    attribute mti_svvh_generic_type of device_id_3 : constant is 1;
    attribute mti_svvh_generic_type of revision_id_data_3 : constant is 1;
    attribute mti_svvh_generic_type of revision_id_3 : constant is 1;
    attribute mti_svvh_generic_type of class_code_data_3 : constant is 1;
    attribute mti_svvh_generic_type of class_code_3 : constant is 1;
    attribute mti_svvh_generic_type of subsystem_vendor_id_data_3 : constant is 1;
    attribute mti_svvh_generic_type of subsystem_vendor_id_3 : constant is 1;
    attribute mti_svvh_generic_type of subsystem_device_id_data_3 : constant is 1;
    attribute mti_svvh_generic_type of subsystem_device_id_3 : constant is 1;
    attribute mti_svvh_generic_type of no_soft_reset_3 : constant is 1;
    attribute mti_svvh_generic_type of intel_id_access_3 : constant is 1;
    attribute mti_svvh_generic_type of device_specific_init_3 : constant is 1;
    attribute mti_svvh_generic_type of maximum_current_data_3 : constant is 1;
    attribute mti_svvh_generic_type of maximum_current_3 : constant is 1;
    attribute mti_svvh_generic_type of d1_support_3 : constant is 1;
    attribute mti_svvh_generic_type of d2_support_3 : constant is 1;
    attribute mti_svvh_generic_type of d0_pme_3 : constant is 1;
    attribute mti_svvh_generic_type of d1_pme_3 : constant is 1;
    attribute mti_svvh_generic_type of d2_pme_3 : constant is 1;
    attribute mti_svvh_generic_type of d3_hot_pme_3 : constant is 1;
    attribute mti_svvh_generic_type of d3_cold_pme_3 : constant is 1;
    attribute mti_svvh_generic_type of use_aer_3 : constant is 1;
    attribute mti_svvh_generic_type of low_priority_vc_3 : constant is 1;
    attribute mti_svvh_generic_type of vc_arbitration_3 : constant is 1;
    attribute mti_svvh_generic_type of disable_snoop_packet_3 : constant is 1;
    attribute mti_svvh_generic_type of max_payload_size_3 : constant is 1;
    attribute mti_svvh_generic_type of surprise_down_error_support_3 : constant is 1;
    attribute mti_svvh_generic_type of dll_active_report_support_3 : constant is 1;
    attribute mti_svvh_generic_type of extend_tag_field_3 : constant is 1;
    attribute mti_svvh_generic_type of endpoint_l0_latency_data_3 : constant is 1;
    attribute mti_svvh_generic_type of endpoint_l0_latency_3 : constant is 1;
    attribute mti_svvh_generic_type of endpoint_l1_latency_data_3 : constant is 1;
    attribute mti_svvh_generic_type of endpoint_l1_latency_3 : constant is 1;
    attribute mti_svvh_generic_type of indicator_data_3 : constant is 1;
    attribute mti_svvh_generic_type of indicator_3 : constant is 1;
    attribute mti_svvh_generic_type of role_based_error_reporting_3 : constant is 1;
    attribute mti_svvh_generic_type of slot_power_scale_data_3 : constant is 1;
    attribute mti_svvh_generic_type of slot_power_scale_3 : constant is 1;
    attribute mti_svvh_generic_type of max_link_width_3 : constant is 1;
    attribute mti_svvh_generic_type of enable_l1_aspm_3 : constant is 1;
    attribute mti_svvh_generic_type of enable_l0s_aspm_3 : constant is 1;
    attribute mti_svvh_generic_type of l1_exit_latency_sameclock_data_3 : constant is 1;
    attribute mti_svvh_generic_type of l1_exit_latency_sameclock_3 : constant is 1;
    attribute mti_svvh_generic_type of l1_exit_latency_diffclock_data_3 : constant is 1;
    attribute mti_svvh_generic_type of l1_exit_latency_diffclock_3 : constant is 1;
    attribute mti_svvh_generic_type of hot_plug_support_data_3 : constant is 1;
    attribute mti_svvh_generic_type of hot_plug_support_3 : constant is 1;
    attribute mti_svvh_generic_type of slot_power_limit_data_3 : constant is 1;
    attribute mti_svvh_generic_type of slot_power_limit_3 : constant is 1;
    attribute mti_svvh_generic_type of slot_number_data_3 : constant is 1;
    attribute mti_svvh_generic_type of slot_number_3 : constant is 1;
    attribute mti_svvh_generic_type of diffclock_nfts_count_data_3 : constant is 1;
    attribute mti_svvh_generic_type of diffclock_nfts_count_3 : constant is 1;
    attribute mti_svvh_generic_type of sameclock_nfts_count_data_3 : constant is 1;
    attribute mti_svvh_generic_type of sameclock_nfts_count_3 : constant is 1;
    attribute mti_svvh_generic_type of completion_timeout_3 : constant is 1;
    attribute mti_svvh_generic_type of enable_completion_timeout_disable_3 : constant is 1;
    attribute mti_svvh_generic_type of extended_tag_reset_3 : constant is 1;
    attribute mti_svvh_generic_type of ecrc_check_capable_3 : constant is 1;
    attribute mti_svvh_generic_type of ecrc_gen_capable_3 : constant is 1;
    attribute mti_svvh_generic_type of no_command_completed_3 : constant is 1;
    attribute mti_svvh_generic_type of msi_multi_message_capable_3 : constant is 1;
    attribute mti_svvh_generic_type of msi_64bit_addressing_capable_3 : constant is 1;
    attribute mti_svvh_generic_type of msi_masking_capable_3 : constant is 1;
    attribute mti_svvh_generic_type of msi_support_3 : constant is 1;
    attribute mti_svvh_generic_type of interrupt_pin_3 : constant is 1;
    attribute mti_svvh_generic_type of enable_function_msix_support_3 : constant is 1;
    attribute mti_svvh_generic_type of msix_table_size_data_3 : constant is 1;
    attribute mti_svvh_generic_type of msix_table_size_3 : constant is 1;
    attribute mti_svvh_generic_type of msix_table_bir_data_3 : constant is 1;
    attribute mti_svvh_generic_type of msix_table_bir_3 : constant is 1;
    attribute mti_svvh_generic_type of msix_table_offset_data_3 : constant is 1;
    attribute mti_svvh_generic_type of msix_table_offset_3 : constant is 1;
    attribute mti_svvh_generic_type of msix_pba_bir_data_3 : constant is 1;
    attribute mti_svvh_generic_type of msix_pba_bir_3 : constant is 1;
    attribute mti_svvh_generic_type of msix_pba_offset_data_3 : constant is 1;
    attribute mti_svvh_generic_type of msix_pba_offset_3 : constant is 1;
    attribute mti_svvh_generic_type of bridge_port_vga_enable_3 : constant is 1;
    attribute mti_svvh_generic_type of bridge_port_ssid_support_3 : constant is 1;
    attribute mti_svvh_generic_type of ssvid_data_3 : constant is 1;
    attribute mti_svvh_generic_type of ssvid_3 : constant is 1;
    attribute mti_svvh_generic_type of ssid_data_3 : constant is 1;
    attribute mti_svvh_generic_type of ssid_3 : constant is 1;
    attribute mti_svvh_generic_type of eie_before_nfts_count_data_3 : constant is 1;
    attribute mti_svvh_generic_type of eie_before_nfts_count_3 : constant is 1;
    attribute mti_svvh_generic_type of gen2_diffclock_nfts_count_data_3 : constant is 1;
    attribute mti_svvh_generic_type of gen2_diffclock_nfts_count_3 : constant is 1;
    attribute mti_svvh_generic_type of gen2_sameclock_nfts_count_data_3 : constant is 1;
    attribute mti_svvh_generic_type of gen2_sameclock_nfts_count_3 : constant is 1;
    attribute mti_svvh_generic_type of deemphasis_enable_3 : constant is 1;
    attribute mti_svvh_generic_type of pcie_spec_version_3 : constant is 1;
    attribute mti_svvh_generic_type of l0_exit_latency_sameclock_data_3 : constant is 1;
    attribute mti_svvh_generic_type of l0_exit_latency_sameclock_3 : constant is 1;
    attribute mti_svvh_generic_type of l0_exit_latency_diffclock_data_3 : constant is 1;
    attribute mti_svvh_generic_type of l0_exit_latency_diffclock_3 : constant is 1;
    attribute mti_svvh_generic_type of rx_ei_l0s_3 : constant is 1;
    attribute mti_svvh_generic_type of l2_async_logic_3 : constant is 1;
    attribute mti_svvh_generic_type of aspm_optionality_3 : constant is 1;
    attribute mti_svvh_generic_type of flr_capability_3 : constant is 1;
    attribute mti_svvh_generic_type of bar0_io_space_3 : constant is 1;
    attribute mti_svvh_generic_type of bar0_64bit_mem_space_3 : constant is 1;
    attribute mti_svvh_generic_type of bar0_prefetchable_3 : constant is 1;
    attribute mti_svvh_generic_type of bar0_size_mask_data_3 : constant is 1;
    attribute mti_svvh_generic_type of bar0_size_mask_3 : constant is 1;
    attribute mti_svvh_generic_type of bar1_io_space_3 : constant is 1;
    attribute mti_svvh_generic_type of bar1_64bit_mem_space_3 : constant is 1;
    attribute mti_svvh_generic_type of bar1_prefetchable_3 : constant is 1;
    attribute mti_svvh_generic_type of bar1_size_mask_data_3 : constant is 1;
    attribute mti_svvh_generic_type of bar1_size_mask_3 : constant is 1;
    attribute mti_svvh_generic_type of bar2_io_space_3 : constant is 1;
    attribute mti_svvh_generic_type of bar2_64bit_mem_space_3 : constant is 1;
    attribute mti_svvh_generic_type of bar2_prefetchable_3 : constant is 1;
    attribute mti_svvh_generic_type of bar2_size_mask_data_3 : constant is 1;
    attribute mti_svvh_generic_type of bar2_size_mask_3 : constant is 1;
    attribute mti_svvh_generic_type of bar3_io_space_3 : constant is 1;
    attribute mti_svvh_generic_type of bar3_64bit_mem_space_3 : constant is 1;
    attribute mti_svvh_generic_type of bar3_prefetchable_3 : constant is 1;
    attribute mti_svvh_generic_type of bar3_size_mask_data_3 : constant is 1;
    attribute mti_svvh_generic_type of bar3_size_mask_3 : constant is 1;
    attribute mti_svvh_generic_type of bar4_io_space_3 : constant is 1;
    attribute mti_svvh_generic_type of bar4_64bit_mem_space_3 : constant is 1;
    attribute mti_svvh_generic_type of bar4_prefetchable_3 : constant is 1;
    attribute mti_svvh_generic_type of bar4_size_mask_data_3 : constant is 1;
    attribute mti_svvh_generic_type of bar4_size_mask_3 : constant is 1;
    attribute mti_svvh_generic_type of bar5_io_space_3 : constant is 1;
    attribute mti_svvh_generic_type of bar5_64bit_mem_space_3 : constant is 1;
    attribute mti_svvh_generic_type of bar5_prefetchable_3 : constant is 1;
    attribute mti_svvh_generic_type of bar5_size_mask_data_3 : constant is 1;
    attribute mti_svvh_generic_type of bar5_size_mask_3 : constant is 1;
    attribute mti_svvh_generic_type of expansion_base_address_register_data_3 : constant is 1;
    attribute mti_svvh_generic_type of expansion_base_address_register_3 : constant is 1;
    attribute mti_svvh_generic_type of io_window_addr_width_3 : constant is 1;
    attribute mti_svvh_generic_type of prefetchable_mem_window_addr_width_3 : constant is 1;
    attribute mti_svvh_generic_type of vendor_id_data_4 : constant is 1;
    attribute mti_svvh_generic_type of vendor_id_4 : constant is 1;
    attribute mti_svvh_generic_type of device_id_data_4 : constant is 1;
    attribute mti_svvh_generic_type of device_id_4 : constant is 1;
    attribute mti_svvh_generic_type of revision_id_data_4 : constant is 1;
    attribute mti_svvh_generic_type of revision_id_4 : constant is 1;
    attribute mti_svvh_generic_type of class_code_data_4 : constant is 1;
    attribute mti_svvh_generic_type of class_code_4 : constant is 1;
    attribute mti_svvh_generic_type of subsystem_vendor_id_data_4 : constant is 1;
    attribute mti_svvh_generic_type of subsystem_vendor_id_4 : constant is 1;
    attribute mti_svvh_generic_type of subsystem_device_id_data_4 : constant is 1;
    attribute mti_svvh_generic_type of subsystem_device_id_4 : constant is 1;
    attribute mti_svvh_generic_type of no_soft_reset_4 : constant is 1;
    attribute mti_svvh_generic_type of intel_id_access_4 : constant is 1;
    attribute mti_svvh_generic_type of device_specific_init_4 : constant is 1;
    attribute mti_svvh_generic_type of maximum_current_data_4 : constant is 1;
    attribute mti_svvh_generic_type of maximum_current_4 : constant is 1;
    attribute mti_svvh_generic_type of d1_support_4 : constant is 1;
    attribute mti_svvh_generic_type of d2_support_4 : constant is 1;
    attribute mti_svvh_generic_type of d0_pme_4 : constant is 1;
    attribute mti_svvh_generic_type of d1_pme_4 : constant is 1;
    attribute mti_svvh_generic_type of d2_pme_4 : constant is 1;
    attribute mti_svvh_generic_type of d3_hot_pme_4 : constant is 1;
    attribute mti_svvh_generic_type of d3_cold_pme_4 : constant is 1;
    attribute mti_svvh_generic_type of use_aer_4 : constant is 1;
    attribute mti_svvh_generic_type of low_priority_vc_4 : constant is 1;
    attribute mti_svvh_generic_type of vc_arbitration_4 : constant is 1;
    attribute mti_svvh_generic_type of disable_snoop_packet_4 : constant is 1;
    attribute mti_svvh_generic_type of max_payload_size_4 : constant is 1;
    attribute mti_svvh_generic_type of surprise_down_error_support_4 : constant is 1;
    attribute mti_svvh_generic_type of dll_active_report_support_4 : constant is 1;
    attribute mti_svvh_generic_type of extend_tag_field_4 : constant is 1;
    attribute mti_svvh_generic_type of endpoint_l0_latency_data_4 : constant is 1;
    attribute mti_svvh_generic_type of endpoint_l0_latency_4 : constant is 1;
    attribute mti_svvh_generic_type of endpoint_l1_latency_data_4 : constant is 1;
    attribute mti_svvh_generic_type of endpoint_l1_latency_4 : constant is 1;
    attribute mti_svvh_generic_type of indicator_data_4 : constant is 1;
    attribute mti_svvh_generic_type of indicator_4 : constant is 1;
    attribute mti_svvh_generic_type of role_based_error_reporting_4 : constant is 1;
    attribute mti_svvh_generic_type of slot_power_scale_data_4 : constant is 1;
    attribute mti_svvh_generic_type of slot_power_scale_4 : constant is 1;
    attribute mti_svvh_generic_type of max_link_width_4 : constant is 1;
    attribute mti_svvh_generic_type of enable_l1_aspm_4 : constant is 1;
    attribute mti_svvh_generic_type of enable_l0s_aspm_4 : constant is 1;
    attribute mti_svvh_generic_type of l1_exit_latency_sameclock_data_4 : constant is 1;
    attribute mti_svvh_generic_type of l1_exit_latency_sameclock_4 : constant is 1;
    attribute mti_svvh_generic_type of l1_exit_latency_diffclock_data_4 : constant is 1;
    attribute mti_svvh_generic_type of l1_exit_latency_diffclock_4 : constant is 1;
    attribute mti_svvh_generic_type of hot_plug_support_data_4 : constant is 1;
    attribute mti_svvh_generic_type of hot_plug_support_4 : constant is 1;
    attribute mti_svvh_generic_type of slot_power_limit_data_4 : constant is 1;
    attribute mti_svvh_generic_type of slot_power_limit_4 : constant is 1;
    attribute mti_svvh_generic_type of slot_number_data_4 : constant is 1;
    attribute mti_svvh_generic_type of slot_number_4 : constant is 1;
    attribute mti_svvh_generic_type of diffclock_nfts_count_data_4 : constant is 1;
    attribute mti_svvh_generic_type of diffclock_nfts_count_4 : constant is 1;
    attribute mti_svvh_generic_type of sameclock_nfts_count_data_4 : constant is 1;
    attribute mti_svvh_generic_type of sameclock_nfts_count_4 : constant is 1;
    attribute mti_svvh_generic_type of completion_timeout_4 : constant is 1;
    attribute mti_svvh_generic_type of enable_completion_timeout_disable_4 : constant is 1;
    attribute mti_svvh_generic_type of extended_tag_reset_4 : constant is 1;
    attribute mti_svvh_generic_type of ecrc_check_capable_4 : constant is 1;
    attribute mti_svvh_generic_type of ecrc_gen_capable_4 : constant is 1;
    attribute mti_svvh_generic_type of no_command_completed_4 : constant is 1;
    attribute mti_svvh_generic_type of msi_multi_message_capable_4 : constant is 1;
    attribute mti_svvh_generic_type of msi_64bit_addressing_capable_4 : constant is 1;
    attribute mti_svvh_generic_type of msi_masking_capable_4 : constant is 1;
    attribute mti_svvh_generic_type of msi_support_4 : constant is 1;
    attribute mti_svvh_generic_type of interrupt_pin_4 : constant is 1;
    attribute mti_svvh_generic_type of enable_function_msix_support_4 : constant is 1;
    attribute mti_svvh_generic_type of msix_table_size_data_4 : constant is 1;
    attribute mti_svvh_generic_type of msix_table_size_4 : constant is 1;
    attribute mti_svvh_generic_type of msix_table_bir_data_4 : constant is 1;
    attribute mti_svvh_generic_type of msix_table_bir_4 : constant is 1;
    attribute mti_svvh_generic_type of msix_table_offset_data_4 : constant is 1;
    attribute mti_svvh_generic_type of msix_table_offset_4 : constant is 1;
    attribute mti_svvh_generic_type of msix_pba_bir_data_4 : constant is 1;
    attribute mti_svvh_generic_type of msix_pba_bir_4 : constant is 1;
    attribute mti_svvh_generic_type of msix_pba_offset_data_4 : constant is 1;
    attribute mti_svvh_generic_type of msix_pba_offset_4 : constant is 1;
    attribute mti_svvh_generic_type of bridge_port_vga_enable_4 : constant is 1;
    attribute mti_svvh_generic_type of bridge_port_ssid_support_4 : constant is 1;
    attribute mti_svvh_generic_type of ssvid_data_4 : constant is 1;
    attribute mti_svvh_generic_type of ssvid_4 : constant is 1;
    attribute mti_svvh_generic_type of ssid_data_4 : constant is 1;
    attribute mti_svvh_generic_type of ssid_4 : constant is 1;
    attribute mti_svvh_generic_type of eie_before_nfts_count_data_4 : constant is 1;
    attribute mti_svvh_generic_type of eie_before_nfts_count_4 : constant is 1;
    attribute mti_svvh_generic_type of gen2_diffclock_nfts_count_data_4 : constant is 1;
    attribute mti_svvh_generic_type of gen2_diffclock_nfts_count_4 : constant is 1;
    attribute mti_svvh_generic_type of gen2_sameclock_nfts_count_data_4 : constant is 1;
    attribute mti_svvh_generic_type of gen2_sameclock_nfts_count_4 : constant is 1;
    attribute mti_svvh_generic_type of deemphasis_enable_4 : constant is 1;
    attribute mti_svvh_generic_type of pcie_spec_version_4 : constant is 1;
    attribute mti_svvh_generic_type of l0_exit_latency_sameclock_data_4 : constant is 1;
    attribute mti_svvh_generic_type of l0_exit_latency_sameclock_4 : constant is 1;
    attribute mti_svvh_generic_type of l0_exit_latency_diffclock_data_4 : constant is 1;
    attribute mti_svvh_generic_type of l0_exit_latency_diffclock_4 : constant is 1;
    attribute mti_svvh_generic_type of rx_ei_l0s_4 : constant is 1;
    attribute mti_svvh_generic_type of l2_async_logic_4 : constant is 1;
    attribute mti_svvh_generic_type of aspm_optionality_4 : constant is 1;
    attribute mti_svvh_generic_type of flr_capability_4 : constant is 1;
    attribute mti_svvh_generic_type of bar0_io_space_4 : constant is 1;
    attribute mti_svvh_generic_type of bar0_64bit_mem_space_4 : constant is 1;
    attribute mti_svvh_generic_type of bar0_prefetchable_4 : constant is 1;
    attribute mti_svvh_generic_type of bar0_size_mask_data_4 : constant is 1;
    attribute mti_svvh_generic_type of bar0_size_mask_4 : constant is 1;
    attribute mti_svvh_generic_type of bar1_io_space_4 : constant is 1;
    attribute mti_svvh_generic_type of bar1_64bit_mem_space_4 : constant is 1;
    attribute mti_svvh_generic_type of bar1_prefetchable_4 : constant is 1;
    attribute mti_svvh_generic_type of bar1_size_mask_data_4 : constant is 1;
    attribute mti_svvh_generic_type of bar1_size_mask_4 : constant is 1;
    attribute mti_svvh_generic_type of bar2_io_space_4 : constant is 1;
    attribute mti_svvh_generic_type of bar2_64bit_mem_space_4 : constant is 1;
    attribute mti_svvh_generic_type of bar2_prefetchable_4 : constant is 1;
    attribute mti_svvh_generic_type of bar2_size_mask_data_4 : constant is 1;
    attribute mti_svvh_generic_type of bar2_size_mask_4 : constant is 1;
    attribute mti_svvh_generic_type of bar3_io_space_4 : constant is 1;
    attribute mti_svvh_generic_type of bar3_64bit_mem_space_4 : constant is 1;
    attribute mti_svvh_generic_type of bar3_prefetchable_4 : constant is 1;
    attribute mti_svvh_generic_type of bar3_size_mask_data_4 : constant is 1;
    attribute mti_svvh_generic_type of bar3_size_mask_4 : constant is 1;
    attribute mti_svvh_generic_type of bar4_io_space_4 : constant is 1;
    attribute mti_svvh_generic_type of bar4_64bit_mem_space_4 : constant is 1;
    attribute mti_svvh_generic_type of bar4_prefetchable_4 : constant is 1;
    attribute mti_svvh_generic_type of bar4_size_mask_data_4 : constant is 1;
    attribute mti_svvh_generic_type of bar4_size_mask_4 : constant is 1;
    attribute mti_svvh_generic_type of bar5_io_space_4 : constant is 1;
    attribute mti_svvh_generic_type of bar5_64bit_mem_space_4 : constant is 1;
    attribute mti_svvh_generic_type of bar5_prefetchable_4 : constant is 1;
    attribute mti_svvh_generic_type of bar5_size_mask_data_4 : constant is 1;
    attribute mti_svvh_generic_type of bar5_size_mask_4 : constant is 1;
    attribute mti_svvh_generic_type of expansion_base_address_register_data_4 : constant is 1;
    attribute mti_svvh_generic_type of expansion_base_address_register_4 : constant is 1;
    attribute mti_svvh_generic_type of io_window_addr_width_4 : constant is 1;
    attribute mti_svvh_generic_type of prefetchable_mem_window_addr_width_4 : constant is 1;
    attribute mti_svvh_generic_type of vendor_id_data_5 : constant is 1;
    attribute mti_svvh_generic_type of vendor_id_5 : constant is 1;
    attribute mti_svvh_generic_type of device_id_data_5 : constant is 1;
    attribute mti_svvh_generic_type of device_id_5 : constant is 1;
    attribute mti_svvh_generic_type of revision_id_data_5 : constant is 1;
    attribute mti_svvh_generic_type of revision_id_5 : constant is 1;
    attribute mti_svvh_generic_type of class_code_data_5 : constant is 1;
    attribute mti_svvh_generic_type of class_code_5 : constant is 1;
    attribute mti_svvh_generic_type of subsystem_vendor_id_data_5 : constant is 1;
    attribute mti_svvh_generic_type of subsystem_vendor_id_5 : constant is 1;
    attribute mti_svvh_generic_type of subsystem_device_id_data_5 : constant is 1;
    attribute mti_svvh_generic_type of subsystem_device_id_5 : constant is 1;
    attribute mti_svvh_generic_type of no_soft_reset_5 : constant is 1;
    attribute mti_svvh_generic_type of intel_id_access_5 : constant is 1;
    attribute mti_svvh_generic_type of device_specific_init_5 : constant is 1;
    attribute mti_svvh_generic_type of maximum_current_data_5 : constant is 1;
    attribute mti_svvh_generic_type of maximum_current_5 : constant is 1;
    attribute mti_svvh_generic_type of d1_support_5 : constant is 1;
    attribute mti_svvh_generic_type of d2_support_5 : constant is 1;
    attribute mti_svvh_generic_type of d0_pme_5 : constant is 1;
    attribute mti_svvh_generic_type of d1_pme_5 : constant is 1;
    attribute mti_svvh_generic_type of d2_pme_5 : constant is 1;
    attribute mti_svvh_generic_type of d3_hot_pme_5 : constant is 1;
    attribute mti_svvh_generic_type of d3_cold_pme_5 : constant is 1;
    attribute mti_svvh_generic_type of use_aer_5 : constant is 1;
    attribute mti_svvh_generic_type of low_priority_vc_5 : constant is 1;
    attribute mti_svvh_generic_type of vc_arbitration_5 : constant is 1;
    attribute mti_svvh_generic_type of disable_snoop_packet_5 : constant is 1;
    attribute mti_svvh_generic_type of max_payload_size_5 : constant is 1;
    attribute mti_svvh_generic_type of surprise_down_error_support_5 : constant is 1;
    attribute mti_svvh_generic_type of dll_active_report_support_5 : constant is 1;
    attribute mti_svvh_generic_type of extend_tag_field_5 : constant is 1;
    attribute mti_svvh_generic_type of endpoint_l0_latency_data_5 : constant is 1;
    attribute mti_svvh_generic_type of endpoint_l0_latency_5 : constant is 1;
    attribute mti_svvh_generic_type of endpoint_l1_latency_data_5 : constant is 1;
    attribute mti_svvh_generic_type of endpoint_l1_latency_5 : constant is 1;
    attribute mti_svvh_generic_type of indicator_data_5 : constant is 1;
    attribute mti_svvh_generic_type of indicator_5 : constant is 1;
    attribute mti_svvh_generic_type of role_based_error_reporting_5 : constant is 1;
    attribute mti_svvh_generic_type of slot_power_scale_data_5 : constant is 1;
    attribute mti_svvh_generic_type of slot_power_scale_5 : constant is 1;
    attribute mti_svvh_generic_type of max_link_width_5 : constant is 1;
    attribute mti_svvh_generic_type of enable_l1_aspm_5 : constant is 1;
    attribute mti_svvh_generic_type of enable_l0s_aspm_5 : constant is 1;
    attribute mti_svvh_generic_type of l1_exit_latency_sameclock_data_5 : constant is 1;
    attribute mti_svvh_generic_type of l1_exit_latency_sameclock_5 : constant is 1;
    attribute mti_svvh_generic_type of l1_exit_latency_diffclock_data_5 : constant is 1;
    attribute mti_svvh_generic_type of l1_exit_latency_diffclock_5 : constant is 1;
    attribute mti_svvh_generic_type of hot_plug_support_data_5 : constant is 1;
    attribute mti_svvh_generic_type of hot_plug_support_5 : constant is 1;
    attribute mti_svvh_generic_type of slot_power_limit_data_5 : constant is 1;
    attribute mti_svvh_generic_type of slot_power_limit_5 : constant is 1;
    attribute mti_svvh_generic_type of slot_number_data_5 : constant is 1;
    attribute mti_svvh_generic_type of slot_number_5 : constant is 1;
    attribute mti_svvh_generic_type of diffclock_nfts_count_data_5 : constant is 1;
    attribute mti_svvh_generic_type of diffclock_nfts_count_5 : constant is 1;
    attribute mti_svvh_generic_type of sameclock_nfts_count_data_5 : constant is 1;
    attribute mti_svvh_generic_type of sameclock_nfts_count_5 : constant is 1;
    attribute mti_svvh_generic_type of completion_timeout_5 : constant is 1;
    attribute mti_svvh_generic_type of enable_completion_timeout_disable_5 : constant is 1;
    attribute mti_svvh_generic_type of extended_tag_reset_5 : constant is 1;
    attribute mti_svvh_generic_type of ecrc_check_capable_5 : constant is 1;
    attribute mti_svvh_generic_type of ecrc_gen_capable_5 : constant is 1;
    attribute mti_svvh_generic_type of no_command_completed_5 : constant is 1;
    attribute mti_svvh_generic_type of msi_multi_message_capable_5 : constant is 1;
    attribute mti_svvh_generic_type of msi_64bit_addressing_capable_5 : constant is 1;
    attribute mti_svvh_generic_type of msi_masking_capable_5 : constant is 1;
    attribute mti_svvh_generic_type of msi_support_5 : constant is 1;
    attribute mti_svvh_generic_type of interrupt_pin_5 : constant is 1;
    attribute mti_svvh_generic_type of enable_function_msix_support_5 : constant is 1;
    attribute mti_svvh_generic_type of msix_table_size_data_5 : constant is 1;
    attribute mti_svvh_generic_type of msix_table_size_5 : constant is 1;
    attribute mti_svvh_generic_type of msix_table_bir_data_5 : constant is 1;
    attribute mti_svvh_generic_type of msix_table_bir_5 : constant is 1;
    attribute mti_svvh_generic_type of msix_table_offset_data_5 : constant is 1;
    attribute mti_svvh_generic_type of msix_table_offset_5 : constant is 1;
    attribute mti_svvh_generic_type of msix_pba_bir_data_5 : constant is 1;
    attribute mti_svvh_generic_type of msix_pba_bir_5 : constant is 1;
    attribute mti_svvh_generic_type of msix_pba_offset_data_5 : constant is 1;
    attribute mti_svvh_generic_type of msix_pba_offset_5 : constant is 1;
    attribute mti_svvh_generic_type of bridge_port_vga_enable_5 : constant is 1;
    attribute mti_svvh_generic_type of bridge_port_ssid_support_5 : constant is 1;
    attribute mti_svvh_generic_type of ssvid_data_5 : constant is 1;
    attribute mti_svvh_generic_type of ssvid_5 : constant is 1;
    attribute mti_svvh_generic_type of ssid_data_5 : constant is 1;
    attribute mti_svvh_generic_type of ssid_5 : constant is 1;
    attribute mti_svvh_generic_type of eie_before_nfts_count_data_5 : constant is 1;
    attribute mti_svvh_generic_type of eie_before_nfts_count_5 : constant is 1;
    attribute mti_svvh_generic_type of gen2_diffclock_nfts_count_data_5 : constant is 1;
    attribute mti_svvh_generic_type of gen2_diffclock_nfts_count_5 : constant is 1;
    attribute mti_svvh_generic_type of gen2_sameclock_nfts_count_data_5 : constant is 1;
    attribute mti_svvh_generic_type of gen2_sameclock_nfts_count_5 : constant is 1;
    attribute mti_svvh_generic_type of deemphasis_enable_5 : constant is 1;
    attribute mti_svvh_generic_type of pcie_spec_version_5 : constant is 1;
    attribute mti_svvh_generic_type of l0_exit_latency_sameclock_data_5 : constant is 1;
    attribute mti_svvh_generic_type of l0_exit_latency_sameclock_5 : constant is 1;
    attribute mti_svvh_generic_type of l0_exit_latency_diffclock_data_5 : constant is 1;
    attribute mti_svvh_generic_type of l0_exit_latency_diffclock_5 : constant is 1;
    attribute mti_svvh_generic_type of rx_ei_l0s_5 : constant is 1;
    attribute mti_svvh_generic_type of l2_async_logic_5 : constant is 1;
    attribute mti_svvh_generic_type of aspm_optionality_5 : constant is 1;
    attribute mti_svvh_generic_type of flr_capability_5 : constant is 1;
    attribute mti_svvh_generic_type of bar0_io_space_5 : constant is 1;
    attribute mti_svvh_generic_type of bar0_64bit_mem_space_5 : constant is 1;
    attribute mti_svvh_generic_type of bar0_prefetchable_5 : constant is 1;
    attribute mti_svvh_generic_type of bar0_size_mask_data_5 : constant is 1;
    attribute mti_svvh_generic_type of bar0_size_mask_5 : constant is 1;
    attribute mti_svvh_generic_type of bar1_io_space_5 : constant is 1;
    attribute mti_svvh_generic_type of bar1_64bit_mem_space_5 : constant is 1;
    attribute mti_svvh_generic_type of bar1_prefetchable_5 : constant is 1;
    attribute mti_svvh_generic_type of bar1_size_mask_data_5 : constant is 1;
    attribute mti_svvh_generic_type of bar1_size_mask_5 : constant is 1;
    attribute mti_svvh_generic_type of bar2_io_space_5 : constant is 1;
    attribute mti_svvh_generic_type of bar2_64bit_mem_space_5 : constant is 1;
    attribute mti_svvh_generic_type of bar2_prefetchable_5 : constant is 1;
    attribute mti_svvh_generic_type of bar2_size_mask_data_5 : constant is 1;
    attribute mti_svvh_generic_type of bar2_size_mask_5 : constant is 1;
    attribute mti_svvh_generic_type of bar3_io_space_5 : constant is 1;
    attribute mti_svvh_generic_type of bar3_64bit_mem_space_5 : constant is 1;
    attribute mti_svvh_generic_type of bar3_prefetchable_5 : constant is 1;
    attribute mti_svvh_generic_type of bar3_size_mask_data_5 : constant is 1;
    attribute mti_svvh_generic_type of bar3_size_mask_5 : constant is 1;
    attribute mti_svvh_generic_type of bar4_io_space_5 : constant is 1;
    attribute mti_svvh_generic_type of bar4_64bit_mem_space_5 : constant is 1;
    attribute mti_svvh_generic_type of bar4_prefetchable_5 : constant is 1;
    attribute mti_svvh_generic_type of bar4_size_mask_data_5 : constant is 1;
    attribute mti_svvh_generic_type of bar4_size_mask_5 : constant is 1;
    attribute mti_svvh_generic_type of bar5_io_space_5 : constant is 1;
    attribute mti_svvh_generic_type of bar5_64bit_mem_space_5 : constant is 1;
    attribute mti_svvh_generic_type of bar5_prefetchable_5 : constant is 1;
    attribute mti_svvh_generic_type of bar5_size_mask_data_5 : constant is 1;
    attribute mti_svvh_generic_type of bar5_size_mask_5 : constant is 1;
    attribute mti_svvh_generic_type of expansion_base_address_register_data_5 : constant is 1;
    attribute mti_svvh_generic_type of expansion_base_address_register_5 : constant is 1;
    attribute mti_svvh_generic_type of io_window_addr_width_5 : constant is 1;
    attribute mti_svvh_generic_type of prefetchable_mem_window_addr_width_5 : constant is 1;
    attribute mti_svvh_generic_type of vendor_id_data_6 : constant is 1;
    attribute mti_svvh_generic_type of vendor_id_6 : constant is 1;
    attribute mti_svvh_generic_type of device_id_data_6 : constant is 1;
    attribute mti_svvh_generic_type of device_id_6 : constant is 1;
    attribute mti_svvh_generic_type of revision_id_data_6 : constant is 1;
    attribute mti_svvh_generic_type of revision_id_6 : constant is 1;
    attribute mti_svvh_generic_type of class_code_data_6 : constant is 1;
    attribute mti_svvh_generic_type of class_code_6 : constant is 1;
    attribute mti_svvh_generic_type of subsystem_vendor_id_data_6 : constant is 1;
    attribute mti_svvh_generic_type of subsystem_vendor_id_6 : constant is 1;
    attribute mti_svvh_generic_type of subsystem_device_id_data_6 : constant is 1;
    attribute mti_svvh_generic_type of subsystem_device_id_6 : constant is 1;
    attribute mti_svvh_generic_type of no_soft_reset_6 : constant is 1;
    attribute mti_svvh_generic_type of intel_id_access_6 : constant is 1;
    attribute mti_svvh_generic_type of device_specific_init_6 : constant is 1;
    attribute mti_svvh_generic_type of maximum_current_data_6 : constant is 1;
    attribute mti_svvh_generic_type of maximum_current_6 : constant is 1;
    attribute mti_svvh_generic_type of d1_support_6 : constant is 1;
    attribute mti_svvh_generic_type of d2_support_6 : constant is 1;
    attribute mti_svvh_generic_type of d0_pme_6 : constant is 1;
    attribute mti_svvh_generic_type of d1_pme_6 : constant is 1;
    attribute mti_svvh_generic_type of d2_pme_6 : constant is 1;
    attribute mti_svvh_generic_type of d3_hot_pme_6 : constant is 1;
    attribute mti_svvh_generic_type of d3_cold_pme_6 : constant is 1;
    attribute mti_svvh_generic_type of use_aer_6 : constant is 1;
    attribute mti_svvh_generic_type of low_priority_vc_6 : constant is 1;
    attribute mti_svvh_generic_type of vc_arbitration_6 : constant is 1;
    attribute mti_svvh_generic_type of disable_snoop_packet_6 : constant is 1;
    attribute mti_svvh_generic_type of max_payload_size_6 : constant is 1;
    attribute mti_svvh_generic_type of surprise_down_error_support_6 : constant is 1;
    attribute mti_svvh_generic_type of dll_active_report_support_6 : constant is 1;
    attribute mti_svvh_generic_type of extend_tag_field_6 : constant is 1;
    attribute mti_svvh_generic_type of endpoint_l0_latency_data_6 : constant is 1;
    attribute mti_svvh_generic_type of endpoint_l0_latency_6 : constant is 1;
    attribute mti_svvh_generic_type of endpoint_l1_latency_data_6 : constant is 1;
    attribute mti_svvh_generic_type of endpoint_l1_latency_6 : constant is 1;
    attribute mti_svvh_generic_type of indicator_data_6 : constant is 1;
    attribute mti_svvh_generic_type of indicator_6 : constant is 1;
    attribute mti_svvh_generic_type of role_based_error_reporting_6 : constant is 1;
    attribute mti_svvh_generic_type of slot_power_scale_data_6 : constant is 1;
    attribute mti_svvh_generic_type of slot_power_scale_6 : constant is 1;
    attribute mti_svvh_generic_type of max_link_width_6 : constant is 1;
    attribute mti_svvh_generic_type of enable_l1_aspm_6 : constant is 1;
    attribute mti_svvh_generic_type of enable_l0s_aspm_6 : constant is 1;
    attribute mti_svvh_generic_type of l1_exit_latency_sameclock_data_6 : constant is 1;
    attribute mti_svvh_generic_type of l1_exit_latency_sameclock_6 : constant is 1;
    attribute mti_svvh_generic_type of l1_exit_latency_diffclock_data_6 : constant is 1;
    attribute mti_svvh_generic_type of l1_exit_latency_diffclock_6 : constant is 1;
    attribute mti_svvh_generic_type of hot_plug_support_data_6 : constant is 1;
    attribute mti_svvh_generic_type of hot_plug_support_6 : constant is 1;
    attribute mti_svvh_generic_type of slot_power_limit_data_6 : constant is 1;
    attribute mti_svvh_generic_type of slot_power_limit_6 : constant is 1;
    attribute mti_svvh_generic_type of slot_number_data_6 : constant is 1;
    attribute mti_svvh_generic_type of slot_number_6 : constant is 1;
    attribute mti_svvh_generic_type of diffclock_nfts_count_data_6 : constant is 1;
    attribute mti_svvh_generic_type of diffclock_nfts_count_6 : constant is 1;
    attribute mti_svvh_generic_type of sameclock_nfts_count_data_6 : constant is 1;
    attribute mti_svvh_generic_type of sameclock_nfts_count_6 : constant is 1;
    attribute mti_svvh_generic_type of completion_timeout_6 : constant is 1;
    attribute mti_svvh_generic_type of enable_completion_timeout_disable_6 : constant is 1;
    attribute mti_svvh_generic_type of extended_tag_reset_6 : constant is 1;
    attribute mti_svvh_generic_type of ecrc_check_capable_6 : constant is 1;
    attribute mti_svvh_generic_type of ecrc_gen_capable_6 : constant is 1;
    attribute mti_svvh_generic_type of no_command_completed_6 : constant is 1;
    attribute mti_svvh_generic_type of msi_multi_message_capable_6 : constant is 1;
    attribute mti_svvh_generic_type of msi_64bit_addressing_capable_6 : constant is 1;
    attribute mti_svvh_generic_type of msi_masking_capable_6 : constant is 1;
    attribute mti_svvh_generic_type of msi_support_6 : constant is 1;
    attribute mti_svvh_generic_type of interrupt_pin_6 : constant is 1;
    attribute mti_svvh_generic_type of enable_function_msix_support_6 : constant is 1;
    attribute mti_svvh_generic_type of msix_table_size_data_6 : constant is 1;
    attribute mti_svvh_generic_type of msix_table_size_6 : constant is 1;
    attribute mti_svvh_generic_type of msix_table_bir_data_6 : constant is 1;
    attribute mti_svvh_generic_type of msix_table_bir_6 : constant is 1;
    attribute mti_svvh_generic_type of msix_table_offset_data_6 : constant is 1;
    attribute mti_svvh_generic_type of msix_table_offset_6 : constant is 1;
    attribute mti_svvh_generic_type of msix_pba_bir_data_6 : constant is 1;
    attribute mti_svvh_generic_type of msix_pba_bir_6 : constant is 1;
    attribute mti_svvh_generic_type of msix_pba_offset_data_6 : constant is 1;
    attribute mti_svvh_generic_type of msix_pba_offset_6 : constant is 1;
    attribute mti_svvh_generic_type of bridge_port_vga_enable_6 : constant is 1;
    attribute mti_svvh_generic_type of bridge_port_ssid_support_6 : constant is 1;
    attribute mti_svvh_generic_type of ssvid_data_6 : constant is 1;
    attribute mti_svvh_generic_type of ssvid_6 : constant is 1;
    attribute mti_svvh_generic_type of ssid_data_6 : constant is 1;
    attribute mti_svvh_generic_type of ssid_6 : constant is 1;
    attribute mti_svvh_generic_type of eie_before_nfts_count_data_6 : constant is 1;
    attribute mti_svvh_generic_type of eie_before_nfts_count_6 : constant is 1;
    attribute mti_svvh_generic_type of gen2_diffclock_nfts_count_data_6 : constant is 1;
    attribute mti_svvh_generic_type of gen2_diffclock_nfts_count_6 : constant is 1;
    attribute mti_svvh_generic_type of gen2_sameclock_nfts_count_data_6 : constant is 1;
    attribute mti_svvh_generic_type of gen2_sameclock_nfts_count_6 : constant is 1;
    attribute mti_svvh_generic_type of deemphasis_enable_6 : constant is 1;
    attribute mti_svvh_generic_type of pcie_spec_version_6 : constant is 1;
    attribute mti_svvh_generic_type of l0_exit_latency_sameclock_data_6 : constant is 1;
    attribute mti_svvh_generic_type of l0_exit_latency_sameclock_6 : constant is 1;
    attribute mti_svvh_generic_type of l0_exit_latency_diffclock_data_6 : constant is 1;
    attribute mti_svvh_generic_type of l0_exit_latency_diffclock_6 : constant is 1;
    attribute mti_svvh_generic_type of rx_ei_l0s_6 : constant is 1;
    attribute mti_svvh_generic_type of l2_async_logic_6 : constant is 1;
    attribute mti_svvh_generic_type of aspm_optionality_6 : constant is 1;
    attribute mti_svvh_generic_type of flr_capability_6 : constant is 1;
    attribute mti_svvh_generic_type of bar0_io_space_6 : constant is 1;
    attribute mti_svvh_generic_type of bar0_64bit_mem_space_6 : constant is 1;
    attribute mti_svvh_generic_type of bar0_prefetchable_6 : constant is 1;
    attribute mti_svvh_generic_type of bar0_size_mask_data_6 : constant is 1;
    attribute mti_svvh_generic_type of bar0_size_mask_6 : constant is 1;
    attribute mti_svvh_generic_type of bar1_io_space_6 : constant is 1;
    attribute mti_svvh_generic_type of bar1_64bit_mem_space_6 : constant is 1;
    attribute mti_svvh_generic_type of bar1_prefetchable_6 : constant is 1;
    attribute mti_svvh_generic_type of bar1_size_mask_data_6 : constant is 1;
    attribute mti_svvh_generic_type of bar1_size_mask_6 : constant is 1;
    attribute mti_svvh_generic_type of bar2_io_space_6 : constant is 1;
    attribute mti_svvh_generic_type of bar2_64bit_mem_space_6 : constant is 1;
    attribute mti_svvh_generic_type of bar2_prefetchable_6 : constant is 1;
    attribute mti_svvh_generic_type of bar2_size_mask_data_6 : constant is 1;
    attribute mti_svvh_generic_type of bar2_size_mask_6 : constant is 1;
    attribute mti_svvh_generic_type of bar3_io_space_6 : constant is 1;
    attribute mti_svvh_generic_type of bar3_64bit_mem_space_6 : constant is 1;
    attribute mti_svvh_generic_type of bar3_prefetchable_6 : constant is 1;
    attribute mti_svvh_generic_type of bar3_size_mask_data_6 : constant is 1;
    attribute mti_svvh_generic_type of bar3_size_mask_6 : constant is 1;
    attribute mti_svvh_generic_type of bar4_io_space_6 : constant is 1;
    attribute mti_svvh_generic_type of bar4_64bit_mem_space_6 : constant is 1;
    attribute mti_svvh_generic_type of bar4_prefetchable_6 : constant is 1;
    attribute mti_svvh_generic_type of bar4_size_mask_data_6 : constant is 1;
    attribute mti_svvh_generic_type of bar4_size_mask_6 : constant is 1;
    attribute mti_svvh_generic_type of bar5_io_space_6 : constant is 1;
    attribute mti_svvh_generic_type of bar5_64bit_mem_space_6 : constant is 1;
    attribute mti_svvh_generic_type of bar5_prefetchable_6 : constant is 1;
    attribute mti_svvh_generic_type of bar5_size_mask_data_6 : constant is 1;
    attribute mti_svvh_generic_type of bar5_size_mask_6 : constant is 1;
    attribute mti_svvh_generic_type of expansion_base_address_register_data_6 : constant is 1;
    attribute mti_svvh_generic_type of expansion_base_address_register_6 : constant is 1;
    attribute mti_svvh_generic_type of io_window_addr_width_6 : constant is 1;
    attribute mti_svvh_generic_type of prefetchable_mem_window_addr_width_6 : constant is 1;
    attribute mti_svvh_generic_type of vendor_id_data_7 : constant is 1;
    attribute mti_svvh_generic_type of vendor_id_7 : constant is 1;
    attribute mti_svvh_generic_type of device_id_data_7 : constant is 1;
    attribute mti_svvh_generic_type of device_id_7 : constant is 1;
    attribute mti_svvh_generic_type of revision_id_data_7 : constant is 1;
    attribute mti_svvh_generic_type of revision_id_7 : constant is 1;
    attribute mti_svvh_generic_type of class_code_data_7 : constant is 1;
    attribute mti_svvh_generic_type of class_code_7 : constant is 1;
    attribute mti_svvh_generic_type of subsystem_vendor_id_data_7 : constant is 1;
    attribute mti_svvh_generic_type of subsystem_vendor_id_7 : constant is 1;
    attribute mti_svvh_generic_type of subsystem_device_id_data_7 : constant is 1;
    attribute mti_svvh_generic_type of subsystem_device_id_7 : constant is 1;
    attribute mti_svvh_generic_type of no_soft_reset_7 : constant is 1;
    attribute mti_svvh_generic_type of intel_id_access_7 : constant is 1;
    attribute mti_svvh_generic_type of device_specific_init_7 : constant is 1;
    attribute mti_svvh_generic_type of maximum_current_data_7 : constant is 1;
    attribute mti_svvh_generic_type of maximum_current_7 : constant is 1;
    attribute mti_svvh_generic_type of d1_support_7 : constant is 1;
    attribute mti_svvh_generic_type of d2_support_7 : constant is 1;
    attribute mti_svvh_generic_type of d0_pme_7 : constant is 1;
    attribute mti_svvh_generic_type of d1_pme_7 : constant is 1;
    attribute mti_svvh_generic_type of d2_pme_7 : constant is 1;
    attribute mti_svvh_generic_type of d3_hot_pme_7 : constant is 1;
    attribute mti_svvh_generic_type of d3_cold_pme_7 : constant is 1;
    attribute mti_svvh_generic_type of use_aer_7 : constant is 1;
    attribute mti_svvh_generic_type of low_priority_vc_7 : constant is 1;
    attribute mti_svvh_generic_type of vc_arbitration_7 : constant is 1;
    attribute mti_svvh_generic_type of disable_snoop_packet_7 : constant is 1;
    attribute mti_svvh_generic_type of max_payload_size_7 : constant is 1;
    attribute mti_svvh_generic_type of surprise_down_error_support_7 : constant is 1;
    attribute mti_svvh_generic_type of dll_active_report_support_7 : constant is 1;
    attribute mti_svvh_generic_type of extend_tag_field_7 : constant is 1;
    attribute mti_svvh_generic_type of endpoint_l0_latency_data_7 : constant is 1;
    attribute mti_svvh_generic_type of endpoint_l0_latency_7 : constant is 1;
    attribute mti_svvh_generic_type of endpoint_l1_latency_data_7 : constant is 1;
    attribute mti_svvh_generic_type of endpoint_l1_latency_7 : constant is 1;
    attribute mti_svvh_generic_type of indicator_data_7 : constant is 1;
    attribute mti_svvh_generic_type of indicator_7 : constant is 1;
    attribute mti_svvh_generic_type of role_based_error_reporting_7 : constant is 1;
    attribute mti_svvh_generic_type of slot_power_scale_data_7 : constant is 1;
    attribute mti_svvh_generic_type of slot_power_scale_7 : constant is 1;
    attribute mti_svvh_generic_type of max_link_width_7 : constant is 1;
    attribute mti_svvh_generic_type of enable_l1_aspm_7 : constant is 1;
    attribute mti_svvh_generic_type of enable_l0s_aspm_7 : constant is 1;
    attribute mti_svvh_generic_type of l1_exit_latency_sameclock_data_7 : constant is 1;
    attribute mti_svvh_generic_type of l1_exit_latency_sameclock_7 : constant is 1;
    attribute mti_svvh_generic_type of l1_exit_latency_diffclock_data_7 : constant is 1;
    attribute mti_svvh_generic_type of l1_exit_latency_diffclock_7 : constant is 1;
    attribute mti_svvh_generic_type of hot_plug_support_data_7 : constant is 1;
    attribute mti_svvh_generic_type of hot_plug_support_7 : constant is 1;
    attribute mti_svvh_generic_type of slot_power_limit_data_7 : constant is 1;
    attribute mti_svvh_generic_type of slot_power_limit_7 : constant is 1;
    attribute mti_svvh_generic_type of slot_number_data_7 : constant is 1;
    attribute mti_svvh_generic_type of slot_number_7 : constant is 1;
    attribute mti_svvh_generic_type of diffclock_nfts_count_data_7 : constant is 1;
    attribute mti_svvh_generic_type of diffclock_nfts_count_7 : constant is 1;
    attribute mti_svvh_generic_type of sameclock_nfts_count_data_7 : constant is 1;
    attribute mti_svvh_generic_type of sameclock_nfts_count_7 : constant is 1;
    attribute mti_svvh_generic_type of completion_timeout_7 : constant is 1;
    attribute mti_svvh_generic_type of enable_completion_timeout_disable_7 : constant is 1;
    attribute mti_svvh_generic_type of extended_tag_reset_7 : constant is 1;
    attribute mti_svvh_generic_type of ecrc_check_capable_7 : constant is 1;
    attribute mti_svvh_generic_type of ecrc_gen_capable_7 : constant is 1;
    attribute mti_svvh_generic_type of no_command_completed_7 : constant is 1;
    attribute mti_svvh_generic_type of msi_multi_message_capable_7 : constant is 1;
    attribute mti_svvh_generic_type of msi_64bit_addressing_capable_7 : constant is 1;
    attribute mti_svvh_generic_type of msi_masking_capable_7 : constant is 1;
    attribute mti_svvh_generic_type of msi_support_7 : constant is 1;
    attribute mti_svvh_generic_type of interrupt_pin_7 : constant is 1;
    attribute mti_svvh_generic_type of enable_function_msix_support_7 : constant is 1;
    attribute mti_svvh_generic_type of msix_table_size_data_7 : constant is 1;
    attribute mti_svvh_generic_type of msix_table_size_7 : constant is 1;
    attribute mti_svvh_generic_type of msix_table_bir_data_7 : constant is 1;
    attribute mti_svvh_generic_type of msix_table_bir_7 : constant is 1;
    attribute mti_svvh_generic_type of msix_table_offset_data_7 : constant is 1;
    attribute mti_svvh_generic_type of msix_table_offset_7 : constant is 1;
    attribute mti_svvh_generic_type of msix_pba_bir_data_7 : constant is 1;
    attribute mti_svvh_generic_type of msix_pba_bir_7 : constant is 1;
    attribute mti_svvh_generic_type of msix_pba_offset_data_7 : constant is 1;
    attribute mti_svvh_generic_type of msix_pba_offset_7 : constant is 1;
    attribute mti_svvh_generic_type of bridge_port_vga_enable_7 : constant is 1;
    attribute mti_svvh_generic_type of bridge_port_ssid_support_7 : constant is 1;
    attribute mti_svvh_generic_type of ssvid_data_7 : constant is 1;
    attribute mti_svvh_generic_type of ssvid_7 : constant is 1;
    attribute mti_svvh_generic_type of ssid_data_7 : constant is 1;
    attribute mti_svvh_generic_type of ssid_7 : constant is 1;
    attribute mti_svvh_generic_type of eie_before_nfts_count_data_7 : constant is 1;
    attribute mti_svvh_generic_type of eie_before_nfts_count_7 : constant is 1;
    attribute mti_svvh_generic_type of gen2_diffclock_nfts_count_data_7 : constant is 1;
    attribute mti_svvh_generic_type of gen2_diffclock_nfts_count_7 : constant is 1;
    attribute mti_svvh_generic_type of gen2_sameclock_nfts_count_data_7 : constant is 1;
    attribute mti_svvh_generic_type of gen2_sameclock_nfts_count_7 : constant is 1;
    attribute mti_svvh_generic_type of deemphasis_enable_7 : constant is 1;
    attribute mti_svvh_generic_type of pcie_spec_version_7 : constant is 1;
    attribute mti_svvh_generic_type of l0_exit_latency_sameclock_data_7 : constant is 1;
    attribute mti_svvh_generic_type of l0_exit_latency_sameclock_7 : constant is 1;
    attribute mti_svvh_generic_type of l0_exit_latency_diffclock_data_7 : constant is 1;
    attribute mti_svvh_generic_type of l0_exit_latency_diffclock_7 : constant is 1;
    attribute mti_svvh_generic_type of rx_ei_l0s_7 : constant is 1;
    attribute mti_svvh_generic_type of l2_async_logic_7 : constant is 1;
    attribute mti_svvh_generic_type of aspm_optionality_7 : constant is 1;
    attribute mti_svvh_generic_type of flr_capability_7 : constant is 1;
    attribute mti_svvh_generic_type of bar0_io_space_7 : constant is 1;
    attribute mti_svvh_generic_type of bar0_64bit_mem_space_7 : constant is 1;
    attribute mti_svvh_generic_type of bar0_prefetchable_7 : constant is 1;
    attribute mti_svvh_generic_type of bar0_size_mask_data_7 : constant is 1;
    attribute mti_svvh_generic_type of bar0_size_mask_7 : constant is 1;
    attribute mti_svvh_generic_type of bar1_io_space_7 : constant is 1;
    attribute mti_svvh_generic_type of bar1_64bit_mem_space_7 : constant is 1;
    attribute mti_svvh_generic_type of bar1_prefetchable_7 : constant is 1;
    attribute mti_svvh_generic_type of bar1_size_mask_data_7 : constant is 1;
    attribute mti_svvh_generic_type of bar1_size_mask_7 : constant is 1;
    attribute mti_svvh_generic_type of bar2_io_space_7 : constant is 1;
    attribute mti_svvh_generic_type of bar2_64bit_mem_space_7 : constant is 1;
    attribute mti_svvh_generic_type of bar2_prefetchable_7 : constant is 1;
    attribute mti_svvh_generic_type of bar2_size_mask_data_7 : constant is 1;
    attribute mti_svvh_generic_type of bar2_size_mask_7 : constant is 1;
    attribute mti_svvh_generic_type of bar3_io_space_7 : constant is 1;
    attribute mti_svvh_generic_type of bar3_64bit_mem_space_7 : constant is 1;
    attribute mti_svvh_generic_type of bar3_prefetchable_7 : constant is 1;
    attribute mti_svvh_generic_type of bar3_size_mask_data_7 : constant is 1;
    attribute mti_svvh_generic_type of bar3_size_mask_7 : constant is 1;
    attribute mti_svvh_generic_type of bar4_io_space_7 : constant is 1;
    attribute mti_svvh_generic_type of bar4_64bit_mem_space_7 : constant is 1;
    attribute mti_svvh_generic_type of bar4_prefetchable_7 : constant is 1;
    attribute mti_svvh_generic_type of bar4_size_mask_data_7 : constant is 1;
    attribute mti_svvh_generic_type of bar4_size_mask_7 : constant is 1;
    attribute mti_svvh_generic_type of bar5_io_space_7 : constant is 1;
    attribute mti_svvh_generic_type of bar5_64bit_mem_space_7 : constant is 1;
    attribute mti_svvh_generic_type of bar5_prefetchable_7 : constant is 1;
    attribute mti_svvh_generic_type of bar5_size_mask_data_7 : constant is 1;
    attribute mti_svvh_generic_type of bar5_size_mask_7 : constant is 1;
    attribute mti_svvh_generic_type of expansion_base_address_register_data_7 : constant is 1;
    attribute mti_svvh_generic_type of expansion_base_address_register_7 : constant is 1;
    attribute mti_svvh_generic_type of io_window_addr_width_7 : constant is 1;
    attribute mti_svvh_generic_type of prefetchable_mem_window_addr_width_7 : constant is 1;
    attribute mti_svvh_generic_type of porttype_func0 : constant is 1;
    attribute mti_svvh_generic_type of porttype_func1 : constant is 1;
    attribute mti_svvh_generic_type of porttype_func2 : constant is 1;
    attribute mti_svvh_generic_type of porttype_func3 : constant is 1;
    attribute mti_svvh_generic_type of porttype_func4 : constant is 1;
    attribute mti_svvh_generic_type of porttype_func5 : constant is 1;
    attribute mti_svvh_generic_type of porttype_func6 : constant is 1;
    attribute mti_svvh_generic_type of porttype_func7 : constant is 1;
    attribute mti_svvh_generic_type of rxfreqlk_cnt_data : constant is 1;
    attribute mti_svvh_generic_type of rxfreqlk_cnt : constant is 1;
    attribute mti_svvh_generic_type of rxfreqlk_cnt_en : constant is 1;
    attribute mti_svvh_generic_type of testmode_control : constant is 1;
    attribute mti_svvh_generic_type of skp_insertion_control : constant is 1;
    attribute mti_svvh_generic_type of tx_l0s_adjust : constant is 1;
    attribute mti_svvh_generic_type of rx_cdc_almost_full_data : constant is 1;
    attribute mti_svvh_generic_type of rx_cdc_almost_full : constant is 1;
    attribute mti_svvh_generic_type of tx_cdc_almost_full_data : constant is 1;
    attribute mti_svvh_generic_type of tx_cdc_almost_full : constant is 1;
    attribute mti_svvh_generic_type of rx_l0s_count_idl_data : constant is 1;
    attribute mti_svvh_generic_type of rx_l0s_count_idl : constant is 1;
    attribute mti_svvh_generic_type of cdc_dummy_insert_limit_data : constant is 1;
    attribute mti_svvh_generic_type of cdc_dummy_insert_limit : constant is 1;
    attribute mti_svvh_generic_type of ei_delay_powerdown_count_data : constant is 1;
    attribute mti_svvh_generic_type of ei_delay_powerdown_count : constant is 1;
    attribute mti_svvh_generic_type of millisecond_cycle_count_data : constant is 1;
    attribute mti_svvh_generic_type of millisecond_cycle_count : constant is 1;
    attribute mti_svvh_generic_type of skp_os_schedule_count_data : constant is 1;
    attribute mti_svvh_generic_type of skp_os_schedule_count : constant is 1;
    attribute mti_svvh_generic_type of fc_init_timer_data : constant is 1;
    attribute mti_svvh_generic_type of fc_init_timer : constant is 1;
    attribute mti_svvh_generic_type of l01_entry_latency_data : constant is 1;
    attribute mti_svvh_generic_type of l01_entry_latency : constant is 1;
    attribute mti_svvh_generic_type of flow_control_update_count_data : constant is 1;
    attribute mti_svvh_generic_type of flow_control_update_count : constant is 1;
    attribute mti_svvh_generic_type of flow_control_timeout_count_data : constant is 1;
    attribute mti_svvh_generic_type of flow_control_timeout_count : constant is 1;
    attribute mti_svvh_generic_type of vc0_rx_flow_ctrl_posted_header_data : constant is 1;
    attribute mti_svvh_generic_type of vc0_rx_flow_ctrl_posted_header : constant is 1;
    attribute mti_svvh_generic_type of vc0_rx_flow_ctrl_posted_data_data : constant is 1;
    attribute mti_svvh_generic_type of vc0_rx_flow_ctrl_posted_data : constant is 1;
    attribute mti_svvh_generic_type of vc0_rx_flow_ctrl_nonposted_header_data : constant is 1;
    attribute mti_svvh_generic_type of vc0_rx_flow_ctrl_nonposted_header : constant is 1;
    attribute mti_svvh_generic_type of vc0_rx_flow_ctrl_nonposted_data_data : constant is 1;
    attribute mti_svvh_generic_type of vc0_rx_flow_ctrl_nonposted_data : constant is 1;
    attribute mti_svvh_generic_type of vc0_rx_flow_ctrl_compl_header_data : constant is 1;
    attribute mti_svvh_generic_type of vc0_rx_flow_ctrl_compl_header : constant is 1;
    attribute mti_svvh_generic_type of vc0_rx_flow_ctrl_compl_data_data : constant is 1;
    attribute mti_svvh_generic_type of vc0_rx_flow_ctrl_compl_data : constant is 1;
    attribute mti_svvh_generic_type of rx_ptr0_posted_dpram_min_data : constant is 1;
    attribute mti_svvh_generic_type of rx_ptr0_posted_dpram_min : constant is 1;
    attribute mti_svvh_generic_type of rx_ptr0_posted_dpram_max_data : constant is 1;
    attribute mti_svvh_generic_type of rx_ptr0_posted_dpram_max : constant is 1;
    attribute mti_svvh_generic_type of rx_ptr0_nonposted_dpram_min_data : constant is 1;
    attribute mti_svvh_generic_type of rx_ptr0_nonposted_dpram_min : constant is 1;
    attribute mti_svvh_generic_type of rx_ptr0_nonposted_dpram_max_data : constant is 1;
    attribute mti_svvh_generic_type of rx_ptr0_nonposted_dpram_max : constant is 1;
    attribute mti_svvh_generic_type of retry_buffer_last_active_address_data : constant is 1;
    attribute mti_svvh_generic_type of retry_buffer_memory_settings_data : constant is 1;
    attribute mti_svvh_generic_type of retry_buffer_memory_settings : constant is 1;
    attribute mti_svvh_generic_type of vc0_rx_buffer_memory_settings_data : constant is 1;
    attribute mti_svvh_generic_type of vc0_rx_buffer_memory_settings : constant is 1;
    attribute mti_svvh_generic_type of bist_memory_settings_data : constant is 1;
    attribute mti_svvh_generic_type of bist_memory_settings : constant is 1;
    attribute mti_svvh_generic_type of bridge_66mhzcap : constant is 1;
    attribute mti_svvh_generic_type of fastb2bcap : constant is 1;
    attribute mti_svvh_generic_type of devseltim : constant is 1;
    attribute mti_svvh_generic_type of memwrinv : constant is 1;
    attribute mti_svvh_generic_type of credit_buffer_allocation_aux : constant is 1;
    attribute mti_svvh_generic_type of enable_adapter_half_rate_mode : constant is 1;
    attribute mti_svvh_generic_type of vc0_clk_enable : constant is 1;
    attribute mti_svvh_generic_type of vc1_clk_enable : constant is 1;
    attribute mti_svvh_generic_type of register_pipe_signals : constant is 1;
    attribute mti_svvh_generic_type of iei_enable_settings : constant is 1;
    attribute mti_svvh_generic_type of lattim_ro_data : constant is 1;
    attribute mti_svvh_generic_type of lattim : constant is 1;
    attribute mti_svvh_generic_type of br_rcb : constant is 1;
    attribute mti_svvh_generic_type of vsec_id_data : constant is 1;
    attribute mti_svvh_generic_type of vsec_id : constant is 1;
    attribute mti_svvh_generic_type of cvp_enable : constant is 1;
    attribute mti_svvh_generic_type of cvp_rate_sel : constant is 1;
    attribute mti_svvh_generic_type of hard_reset_bypass : constant is 1;
    attribute mti_svvh_generic_type of cvp_data_compressed : constant is 1;
    attribute mti_svvh_generic_type of cvp_data_encrypted : constant is 1;
    attribute mti_svvh_generic_type of cvp_mode_reset : constant is 1;
    attribute mti_svvh_generic_type of cvp_clk_reset : constant is 1;
    attribute mti_svvh_generic_type of vsec_cap_data : constant is 1;
    attribute mti_svvh_generic_type of vsec_cap : constant is 1;
    attribute mti_svvh_generic_type of jtag_id_data : constant is 1;
    attribute mti_svvh_generic_type of jtag_id : constant is 1;
    attribute mti_svvh_generic_type of user_id_data : constant is 1;
    attribute mti_svvh_generic_type of user_id : constant is 1;
    attribute mti_svvh_generic_type of disable_auto_crs : constant is 1;
    attribute mti_svvh_generic_type of altpe2_hip_base_addr_1 : constant is 1;
    attribute mti_svvh_generic_type of altpe2_hip_base_addr_2 : constant is 1;
    attribute mti_svvh_generic_type of altpe2_hip_base_addr_3 : constant is 1;
    attribute mti_svvh_generic_type of altpe2_hip_base_addr_4 : constant is 1;
    attribute mti_svvh_generic_type of altpe2_hip_base_addr_5 : constant is 1;
    attribute mti_svvh_generic_type of altpe2_hip_base_addr_6 : constant is 1;
    attribute mti_svvh_generic_type of altpe2_hip_base_addr_user_1 : constant is 1;
    attribute mti_svvh_generic_type of altpe2_hip_base_addr_user_2 : constant is 1;
    attribute mti_svvh_generic_type of altpe2_hip_base_addr_user_3 : constant is 1;
    attribute mti_svvh_generic_type of altpe2_hip_base_addr_user_4 : constant is 1;
    attribute mti_svvh_generic_type of altpe2_hip_base_addr_user_5 : constant is 1;
    attribute mti_svvh_generic_type of altpe2_hip_base_addr_user_6 : constant is 1;
    attribute mti_svvh_generic_type of cvp_mdio_dis_csr_ctrl_1 : constant is 1;
    attribute mti_svvh_generic_type of cvp_mdio_dis_csr_ctrl_2 : constant is 1;
    attribute mti_svvh_generic_type of cvp_mdio_dis_csr_ctrl_3 : constant is 1;
    attribute mti_svvh_generic_type of cvp_mdio_dis_csr_ctrl_4 : constant is 1;
    attribute mti_svvh_generic_type of cvp_mdio_dis_csr_ctrl_5 : constant is 1;
    attribute mti_svvh_generic_type of cvp_mdio_dis_csr_ctrl_6 : constant is 1;
    attribute mti_svvh_generic_type of dft_broadcast_en_1 : constant is 1;
    attribute mti_svvh_generic_type of dft_broadcast_en_2 : constant is 1;
    attribute mti_svvh_generic_type of dft_broadcast_en_3 : constant is 1;
    attribute mti_svvh_generic_type of dft_broadcast_en_4 : constant is 1;
    attribute mti_svvh_generic_type of dft_broadcast_en_5 : constant is 1;
    attribute mti_svvh_generic_type of dft_broadcast_en_6 : constant is 1;
    attribute mti_svvh_generic_type of electromech_interlock_0 : constant is 1;
    attribute mti_svvh_generic_type of electromech_interlock_1 : constant is 1;
    attribute mti_svvh_generic_type of electromech_interlock_2 : constant is 1;
    attribute mti_svvh_generic_type of electromech_interlock_3 : constant is 1;
    attribute mti_svvh_generic_type of electromech_interlock_4 : constant is 1;
    attribute mti_svvh_generic_type of electromech_interlock_5 : constant is 1;
    attribute mti_svvh_generic_type of electromech_interlock_6 : constant is 1;
    attribute mti_svvh_generic_type of electromech_interlock_7 : constant is 1;
    attribute mti_svvh_generic_type of force_mdio_dis_csr_ctrl_1 : constant is 1;
    attribute mti_svvh_generic_type of force_mdio_dis_csr_ctrl_2 : constant is 1;
    attribute mti_svvh_generic_type of force_mdio_dis_csr_ctrl_3 : constant is 1;
    attribute mti_svvh_generic_type of force_mdio_dis_csr_ctrl_4 : constant is 1;
    attribute mti_svvh_generic_type of force_mdio_dis_csr_ctrl_5 : constant is 1;
    attribute mti_svvh_generic_type of force_mdio_dis_csr_ctrl_6 : constant is 1;
    attribute mti_svvh_generic_type of mdio_cb_opbit_enable : constant is 1;
    attribute mti_svvh_generic_type of plniotri_gate : constant is 1;
    attribute mti_svvh_generic_type of power_isolation_en_1 : constant is 1;
    attribute mti_svvh_generic_type of power_isolation_en_1_data : constant is 1;
    attribute mti_svvh_generic_type of power_isolation_en_2 : constant is 1;
    attribute mti_svvh_generic_type of power_isolation_en_2_data : constant is 1;
    attribute mti_svvh_generic_type of power_isolation_en_3 : constant is 1;
    attribute mti_svvh_generic_type of power_isolation_en_3_data : constant is 1;
    attribute mti_svvh_generic_type of power_isolation_en_4 : constant is 1;
    attribute mti_svvh_generic_type of power_isolation_en_4_data : constant is 1;
    attribute mti_svvh_generic_type of power_isolation_en_5 : constant is 1;
    attribute mti_svvh_generic_type of power_isolation_en_5_data : constant is 1;
    attribute mti_svvh_generic_type of power_isolation_en_6 : constant is 1;
    attribute mti_svvh_generic_type of power_isolation_en_6_data : constant is 1;
    attribute mti_svvh_generic_type of retry_buffer_last_active_address : constant is 1;
    attribute mti_svvh_generic_type of sup_mode : constant is 1;
    attribute mti_svvh_generic_type of hrdrstctrl_en : constant is 1;
    attribute mti_svvh_generic_type of rstctrl_pld_clr : constant is 1;
    attribute mti_svvh_generic_type of rstctrl_debug_en : constant is 1;
    attribute mti_svvh_generic_type of rstctrl_force_inactive_rst : constant is 1;
    attribute mti_svvh_generic_type of rstctrl_perst_enable : constant is 1;
    attribute mti_svvh_generic_type of rstctrl_hip_ep : constant is 1;
    attribute mti_svvh_generic_type of rstctrl_hard_block_enable : constant is 1;
    attribute mti_svvh_generic_type of rstctrl_rx_pma_rstb_inv : constant is 1;
    attribute mti_svvh_generic_type of rstctrl_tx_pma_rstb_inv : constant is 1;
    attribute mti_svvh_generic_type of rstctrl_rx_pcs_rst_n_inv : constant is 1;
    attribute mti_svvh_generic_type of rstctrl_tx_pcs_rst_n_inv : constant is 1;
    attribute mti_svvh_generic_type of rstctrl_altpe2_crst_n_inv : constant is 1;
    attribute mti_svvh_generic_type of rstctrl_altpe2_srst_n_inv : constant is 1;
    attribute mti_svvh_generic_type of rstctrl_altpe2_rst_n_inv : constant is 1;
    attribute mti_svvh_generic_type of rstctrl_tx_pma_syncp_inv : constant is 1;
    attribute mti_svvh_generic_type of rstctrl_1us_count_fref_clk : constant is 1;
    attribute mti_svvh_generic_type of rstctrl_1us_count_fref_clk_value : constant is 1;
    attribute mti_svvh_generic_type of rstctrl_1ms_count_fref_clk : constant is 1;
    attribute mti_svvh_generic_type of rstctrl_1ms_count_fref_clk_value : constant is 1;
    attribute mti_svvh_generic_type of rstctrl_off_cal_done_select : constant is 1;
    attribute mti_svvh_generic_type of rstctrl_rx_pma_rstb_cmu_select : constant is 1;
    attribute mti_svvh_generic_type of rstctrl_rx_pma_rstb_select : constant is 1;
    attribute mti_svvh_generic_type of rstctrl_rx_pll_freq_lock_select : constant is 1;
    attribute mti_svvh_generic_type of rstctrl_mask_tx_pll_lock_select : constant is 1;
    attribute mti_svvh_generic_type of rstctrl_rx_pll_lock_select : constant is 1;
    attribute mti_svvh_generic_type of rstctrl_perstn_select : constant is 1;
    attribute mti_svvh_generic_type of rstctrl_tx_lc_pll_rstb_select : constant is 1;
    attribute mti_svvh_generic_type of rstctrl_fref_clk_select : constant is 1;
    attribute mti_svvh_generic_type of rstctrl_off_cal_en_select : constant is 1;
    attribute mti_svvh_generic_type of rstctrl_tx_pma_syncp_select : constant is 1;
    attribute mti_svvh_generic_type of rstctrl_rx_pcs_rst_n_select : constant is 1;
    attribute mti_svvh_generic_type of rstctrl_tx_cmu_pll_lock_select : constant is 1;
    attribute mti_svvh_generic_type of rstctrl_tx_pcs_rst_n_select : constant is 1;
    attribute mti_svvh_generic_type of rstctrl_tx_lc_pll_lock_select : constant is 1;
    attribute mti_svvh_generic_type of rstctrl_timer_a : constant is 1;
    attribute mti_svvh_generic_type of rstctrl_timer_a_type : constant is 1;
    attribute mti_svvh_generic_type of rstctrl_timer_a_value : constant is 1;
    attribute mti_svvh_generic_type of rstctrl_timer_b : constant is 1;
    attribute mti_svvh_generic_type of rstctrl_timer_b_type : constant is 1;
    attribute mti_svvh_generic_type of rstctrl_timer_b_value : constant is 1;
    attribute mti_svvh_generic_type of rstctrl_timer_c : constant is 1;
    attribute mti_svvh_generic_type of rstctrl_timer_c_type : constant is 1;
    attribute mti_svvh_generic_type of rstctrl_timer_c_value : constant is 1;
    attribute mti_svvh_generic_type of rstctrl_timer_d : constant is 1;
    attribute mti_svvh_generic_type of rstctrl_timer_d_type : constant is 1;
    attribute mti_svvh_generic_type of rstctrl_timer_d_value : constant is 1;
    attribute mti_svvh_generic_type of rstctrl_timer_e : constant is 1;
    attribute mti_svvh_generic_type of rstctrl_timer_e_type : constant is 1;
    attribute mti_svvh_generic_type of rstctrl_timer_e_value : constant is 1;
    attribute mti_svvh_generic_type of rstctrl_timer_f : constant is 1;
    attribute mti_svvh_generic_type of rstctrl_timer_f_type : constant is 1;
    attribute mti_svvh_generic_type of rstctrl_timer_f_value : constant is 1;
    attribute mti_svvh_generic_type of rstctrl_timer_g : constant is 1;
    attribute mti_svvh_generic_type of rstctrl_timer_g_type : constant is 1;
    attribute mti_svvh_generic_type of rstctrl_timer_g_value : constant is 1;
    attribute mti_svvh_generic_type of rstctrl_timer_h : constant is 1;
    attribute mti_svvh_generic_type of rstctrl_timer_h_type : constant is 1;
    attribute mti_svvh_generic_type of rstctrl_timer_h_value : constant is 1;
    attribute mti_svvh_generic_type of rstctrl_timer_i : constant is 1;
    attribute mti_svvh_generic_type of rstctrl_timer_i_type : constant is 1;
    attribute mti_svvh_generic_type of rstctrl_timer_i_value : constant is 1;
    attribute mti_svvh_generic_type of rstctrl_timer_j : constant is 1;
    attribute mti_svvh_generic_type of rstctrl_timer_j_type : constant is 1;
    attribute mti_svvh_generic_type of rstctrl_timer_j_value : constant is 1;
    attribute mti_svvh_generic_type of rstctrl_ltssm_disable : constant is 1;
    attribute mti_svvh_generic_type of cvp_isolation : constant is 1;
end cyclonev_hd_altpe2_hip_top;
