`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
u+2vWE0hvCLEdd1KCLErT/QAAmQkJ5WnVCf3Wk3V1iNKXbRDz/jE1iPM/7mWa+Y4
wl8bMys6LHCjcVXim6mKkxiqx35TlIRocPlEEL6JNvmAKTu4sk+dubLlM7y6sH1r
Nn7chH3jfSiToy1G3KR1PuXRDNirVOpLo6aAchA3MGp/nzf1kWeTuZFg5Y5UznFf
smmaJieXTsqy/HtP4q4Segxrh3Sy11OdPGuKnFn4BBaEoeaytFT1+YOE55m/3Wsw
CoFk2sVOXfzVaN9uhUxjXuThRuLYr0+YC1wYsY27BCaArgqk+AM+pYGeTCqiP+nI
eQsFKkoxrrDtLmjdwFPu/UhVIcadh0sLW/pvnHZukNOOqlbCrKu9CwWCDhp4hIxQ
2tuJCiTaIguYxSidLZ2AgdnipSrN5JmhvFU+Y/JC0A2ApiSb1boWEaA1QFHYPtao
YB8ppRNRfF5Dwc1qPI3JOGaT3X/bHusEf0s6H6E8Tg+wonzi04xjeK18F0o46tO6
fULSY9CWmy5Pmyge5AkObSRr5pdEKWHq4+UOxDfeDqfvagnzPgVXFvre46B+qEtN
dmNE0UBFUCUU1T97Rm5bQTMTLSury8LPe2VW4mgF+B3Qa4htXaRG9p7UrQeXQaAO
YVOAMZ5MEdirka2tNhUJo9zUGQu2Xa2DdBoo/pBggDf0slA6Oqk/gahGY+J8zLKn
ebnc/+w+EU/aOwRY/1tq90c1JqCgZHjA76DfCnFSquIz1MP2Gfj1liHTFl2e21oQ
RLhtQNywTxXblXiSSaK/MJ5EjHpnsCnM/XEE0mk7Ggz+l64CJ9mvAXAbmqVE33Gy
dA3wZsgFGVKHP4QPRpdBro+MUgBNMzIlmaGq7t8WRVqCAFzHvTWO4ZwruiaswEcJ
fxYD+eCQ2SMAS4TteaERtEhDoyF91mu6FHgX9YyaZJelmMCvOew98E2JJRBJ4/Mp
OKnmZNBaMT9HPNq/EgAz1JGBHHG2wnp8TxRyKYiqKB4qnpXGl6tbvFeWgVYDtm/N
BcXxYJoa7dBdywRarIcUlff7jLQvXSlQYx28eN5r3gskavqKfW2SvvR4OLrcRyIk
buNYzv5Y8UE4q7Aqtzhfq+pYtJB62VKbetW2ytGxH0PtN61KT/nP4cJ2/xd7+hAS
ofvFNKQU2ySpsUhWPmM0hSy72FtTUrSwPQ24xID3c8+1BHKwGS+A639m7I125Kqi
2Oc/LqMgrnPAF9+0NsAuMnuehkbKxJU6jiwxmbx3O9Nk6gjiyiDmaizuwjJrfB5x
bM579fwLP4rsAX4v3pT96MGp2NjFELMkWrf8ie31YB4vb6s93maepOC8s46JE916
AGqlc/dB2l0y2kzAzZFcIMU6YicfmccnAt4m80kZqsJYkruD7rj8huLRCrEHzVJ4
H9yy0LCYJAjTYkjQdxtcGB7rAz5c4gp5J4ZODPKZ32es5okU7ggjtvcBiZGLANHH
`protect END_PROTECTED
