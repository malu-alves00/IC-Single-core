`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0zyQrI7VCTX8Tl8wymfR1uFGES9YJgDOfpPrrSCn1sOaI5kcpahkK6y/g8paKoSP
VpI4ZxqvnXjsB3xLZFD7nKHlTG/ZU/nClqwt8ugBYwhjQ/1X6iDSwPSQyAJz/mDC
KaZQqSysVmda6dlkoCKNqHOHGE3j9rqZO9ZhZG/aKwKyxmThdeUptrzH4y85ugFM
kaoiANIQOGGwK8FM1XPqQpxU3085SPAjfZBzmGAJhKbAM83gznRH6/RwXsaud/mN
MuS0ZsfAr0c7jgoDeh0yJelAqk7FCTcKQDOk3k+sGoTuMR+WxEsRHNoZW7rIx78X
adK+QclZ8O5q/sPK1gOjrWDOXKEp6F5AhGngAke0TRaiM/eTf9OPAbxoiL7D4sVe
AIudXRW5ANZ5IBxPQQqu8+jHrYX2V5F/1KU44sayvWNy+FpzJLiBLjEdMEpPeOfN
vc2eFamRiK3ilu5xQjCroeMwHfrxQMUE25Z9L0ghXrHMA1GqOnLD5l9GhXkDCmPa
PCZOyRNwpVKjYNXRGlyUbc++mmtkW0OZB1YH6wTqklUgHQjTPDDF9r2lBt8iQd51
4aDfRGP0od4+WSCfLpTJlHS90iGyI3cANnLT1GSZVzyEwHT9xYsYGD9aI6kkf9PV
qows2F66Nki4TGmQKIc45/vMZT3PjM8L3yzlAjAjtI3Fx0S86zYRAOUB39J6wByu
J4LhtUiwM88JbNDpPINYEY6qwWjmxevIP71VO5/QIQCYIWRNBeeCuhKaD+CrDYuv
Fx0vqjKTsQPNfDg+YazhTXzc1qJC6nzxAfiOidDEtncHcFnPpddqzpNw8zUMvZo0
S9ysU3/dnlhlocfQ7BW8tSI/ML2+TLzw/eUNFbNV2E2tCY2kZXKR82+65IZ1OBQW
DsyvZ6jQQq+zG3eTavtrlreK3eyLTq4aaOFDkj8fKBDWolnu3dw87usygrjuGNtU
d12qz7XZY/GApNL39IuKa5LRWFad9HsWcvgFvr+nl6HfViVr3IUu7/Kv2aCEHYiQ
7jOCYO7fKS2wdIEdHWFNjoeLwkxco2cgxkGp/XXYLaoL+AJggssrGrFnsLauUTVE
PjbaT99gYzkmPLNppW7/VEIymedX1Caap/dAC6oYwEajfDzbRfmnSfsftPbJYsQy
p8J5PNY0vQiGYozS+X4YynWt81BgzMPNnAUpvNed3Z7y5qhekEgnh7PkOzF6Stmc
b5m7BqaAysODu2bQTbtUAutgpNicK3j+xma9wrJlneAI/INVeNT8ICX2RVvv2I/x
x4ctz+OFG7IWPWZ0JFjSNJEjw/Smh8SJt7tA7lqMWLyv4nAjR21OXjAGLEiNr0Gs
LZnKdH4aX9xvExECMwlA+N3ecKNAIGx2aoj4BgHaMJWSj5eLCiJXDGYkmUEjJamR
zuIBvuGB6zaqIsxtvBCJ9GGdEX+uDNC0RYSa8ouY6SBx1CD/Os7pWtl7HyM3SifY
d0QCHFISXSksBNFq6z7V4DmN9HyPW1b2yzYCr0F8rE40DNFFrOa0595nT5BJETYG
3XkyNHrpXnbn0NyS4M/4l1iuumexEFqVyX74T7nRLTilSAHGN0tsAWvP8sjfFwtr
rdI2ixpSnogBZpsIajdwlYMUK3LAVSBdPPUErfD7hIamAYQwoqAD2zgdba4yy2+u
r/Begnzr8TZhLk8EpvjM/YVnPMmS/qNppv8tuIeyGGBzCOZDP5XcUVXNTwqpz3rl
VB3Mvy6hjzunRwWlFzEyulYfjkzPNdzTw3A+4M9JZxrinJfDJYrsBQQKSqWtrTbA
xygSrmuBt0383FSU13GxCoaZZ3ZpEWL21Kp9IzNl3uZYm7FIF/SwgIjoq/LhlAtY
g6boMhtJcKMX6jF5JKLM3Bq1ocnGlN/Dz2JptjLG4rKfbfWGo3vYYrMVqV2S69m5
jTlW7a5UECnQlEzXNrEXX7eyb8TW0PFGNa6ILIAGFSCSEdh1XM8hL01JyenPBQaH
P3Inq3IyafY7KFx20kQ6p8vB7/5014s7CEfTdD5743+SFDHLJLYorXU0KHGjZDc1
49bxdTE89XVzp7svOq93/xeuKDxJ4TZcj1KoRwx0iQF7SW8Pu7UNrVzPbOQGqxuq
1xmSQYu7O7OcCvyQZAklJ4wK5VLd1wJNFZTXOOvNpUNIJ+jhJlpxvDHye5d+ZiRA
itzadupjxT0pWl0Md7LQ3zadjiKzAgSbZAp/p0PDsEy2ahmcbAFHCBv6sUguDTY8
CCttCnCmNC+XVB/2CtH+fkMcHrYSJ/X+48J9zyKLkD+0/YaeXWxMQyOmYxiYjxKE
qzdTRwryGIhk1hU4NukMX+zr8yzqdNsTDeZk1umqL66W9oMy65oa2oA3/xJwA0TS
z2eyKJHT1Ha+bC7EM1f01km7k+/E/REahnkT8JNceFKyP2r/Nltfsk883H8by6zb
7Oy+fm3dS2MfcTmSvubqK0gLo/LS7mtAuetz+z3pmGiAkgdwMTxtua7r/MWl7Tcc
T5TK5xSBVkWNEbe/Efy4NzJopPiUvrzFLCabfqr8JbbBXAdU3KLkrISU4TGe/xTb
O+/OITcpzNZ/KueeF4vogI3HwudFASaQrVbzBJcAadF+tKfve1ffaJKXfiY5hZJj
9qek/SgPQS8NFOpfKlFo6ry4rBwdd0az2K+dG76eOlNJBZoRB6QzHtI7JZVTc7za
oainvtP0/6pL+/Bvk+iW2mBd0HuvrAaGRepdkrlgUJToIqCdHFLU+IVENmqoiUNG
XCKqWmOW9hH3i+gLrSgoXi+uxixwp2IH+AGyyoH7yG8PywCTUELUEfwHeSitH8jM
hIQReJBshcjbBoqfTDyqsumHCpv9WLqY6qzzkE4FrkQdBhbX36f2On4ECHgsGAzl
ZKIWn8wSXMiiMNT906cJm3H0nDKRgHIpqXKdOhHHzRA+yQTPxpkAPMCFeQlrgR3Z
u4AlGIo8FnWKcAfFsK1G1NKliT0sean00ribKOsKYTfYw37JQQWOxsE5Q+H1JOOZ
6+AAZ62hW2oHg2ciUmyccg+PL8ZwhVcryaGbIMIdUTtHvSlomoWd3dUHf5NwVF1b
1+is/gzkdVQQgtjf32/px4lTJvoOP4WKIJPT5kt6vNSGpiO9L0Tt8hO4IsGcR/I7
R2Vzw/yb3+MB72t8l/LQrBuf5xwAj2No1kLOhZFSsXDtkrchg2LGQmWSgWRA9f8y
AESqhmc83+ET8Ur7TI6NbLcFoFwf/5w53P6YzQth6fBbD3UfUtuCjF9ENx34doJi
98wf4vrQ2p8l2RQgqsYMY5EVoiopyejM6LCfXy6Ttrnk0ux8hOqlJXAFlnNJSi2Q
f92YU4fneVkZr7IOalR0RqoY/5v+4jpx4WyIoD3/QZ03svx0eNVuRjDA26nEVn1q
lcwxQ6lPO6LZZ+fxYaiTw43q85L9OshXNarjr7iuWjNqXIKfP7UVfVwk1N2O8DIQ
Cydoyfpv8hi4vlWfhxZzfiRbvNFS8tWdDAf411QnETGvN7GyUuROsRmjjK7YhSHv
vetBa6V7GLM82iPdma+Vf0vOFii1imp6CF9ZQwfpwpWQ04D6YRyX8bJAbizzeCyh
iwIdTAyUi1O/XejX+Jv5s5Zo7iMxMT8D9JZtRR0ij+qJl6yVFGFOOC1TTJ4US4bS
e4tNaIxqPyihAD/CKwaSfvCjCMsGAghktV6GZC2TWBsaA6CDnDm+yRoLBHG5t0kQ
8+75Mr7Ygepolmsr1eYBzdvSyPt4BLANPTul/6RJ9ixtKGiPbJIaRCbjD1WNCD0u
5VJ5hMlZgNWSR/Kf+i2IQYhpzRz+fGr22JTpdOunPtYW6D6byH6OavNybIkjsca8
9aXJtJcv8yDfJ+VcHpjOEcNOyR5dyFyst+okk4AM0UVUsFywHeBowaIt5XXu5HNC
03OtcnV7wzpv4CMl4w7CvcguwadsUlSdRR4P5tELt1TUBzIeQpXDS2illtxmOKL+
5HWjFY7sYwkPmyvDbqf1ga+AFNZfzocB8dfhnbpNTkpyggOsOMcrGnic3EnlOlY6
DRge2K9cAjCzCQ/n0vfSlxAZnok3mybswE8SBOTp8zYfHGzuECAuHThWv6VP1gPZ
h1v347Zyot2na9Vogh8tGoGeyEfAYDmxidaDzsKesxDIV8TZukkFG3qq9gLE1hbL
WxImICI6iu0Vie5RUTgGuPBQAULQuifOMr3T3OLVjHHpQHmGnKrtq0/BgJZz6ja6
aIOGDbbtkpU2UzIDJpit+1sgtk8UuYCPUaodYM6SuvIbMoCBHK1WAbA/U0xNz4Y7
D0THzUEjXI+Y4nSzHEUXLwAFbnD3KahYtyw51lJxLW4qC9CV28gJ0Prs8LYqdb03
VN+LSdGfG/PRfwX86R2zk4LB1viQMpyeX0JkNnOluyaJa0JvIs7q3Kfofir8V0aK
N5YCo2t566vl/m6d49fWIoN6m2Xd2GwFZJffn3XzEYTMyNCMdCPopPLRNUI9TdBY
d9XJUhAKl/grDjwOgLt3RfjBrNnMcT5p9NyKpCskJRNkS+wW6ug8XYQLwoR+z+WI
bLJdwx9LsFAMq+CWxFHftjvAmSRTZatzXO6aQMYntSLgrRSift2gs9xiv/6cRD03
aHcjMKpEYCyZGXQORQWU0/U95/ImJVAmrDdbXNGGPkpzvOZsLqqpVHVdOfWSa/HA
F3Sx4oLRJONnSH+YmWPW4fmUzMtPBxIkTb1+m7YFjn8T/NO8KpdTdEK0KPF+PPhF
Ez3lDtWmMATIPXDmF3d6rJB/Vdesd7cKA7ePYOvBTa8scIvL4mBcw1H36IK16tAu
OD/zjjzzafCLAP6sNMBZHtuMvX52DZwTryl9kGOrIlax36P2jhpsUd9jvGErw/om
ibCjlnGhNwmnVIf+WomxMzr6P6YIdnDq26leFc9jIdMFdypGF8Jc7tzH5KBlmYGX
VhokG5eilTXr68yB3xaHbFLKii8VcNOy4KpMM0weeC9m47nGHPoH+pNGzK0zLROH
nMFTR7iDQx1u3jzeFDhITLXUfijbnj+ZJ1QVtxXf7EW0/FaDCaYbjb9W2R/uT3Mf
4VG31rRo8DzE/hn7HGa77eRUImFO1V8AT9Q40c/lASPnqiiFvQWjDmqp3reZ2cTw
zMetM9HGP+U/BVEDBL6p/3x5wgswSn2dtHP6JKPqEJ9VgNbRx91kL/7hn44kdzb0
z6EKXXu6jFi1MF8TVK9G2Hi3zoB8yKWGaVyrMKPAisTmqaRdAQH/+bBdT9BlUZCg
GokNjyyhw/kdD3MVL+mtn7wZZFNLVPT0HWRj+uKrROjjA3KfrmUSRRetlDbHaPj1
WVRJfLKyAkzwru55PwrGAuR0xNYk0k2vwj4R+E3RWVloKwUviL4PlZaVmtatK3ta
CMuk/jiAp/DPj4w1XSgrv8yS27RiaiqPJeMAMJPuvNzdeXHta9I+fnQMpOnQZb2G
PgEKF2DDEVsiRWW6BqRfKBfEtnI86RJYGrWi1X7mMAmuAF1v9xqimbXIyRO7XD14
souKuRf0gJEv9d1ZVpAbPlYknyU9pbG8ZL/cfYygVLyhWWsO5262w7V7vNcaecQC
lJxvUNu0VGGQOW6+pWDCEcOaSJmBje0vwpZsyTbkzBAKQlqEqn2f8SYqsjw7omZk
9IESNs0/a9TyLr3M2U45yZX7J3VFlg1tcN2cRUpbChxJtJB6izr0Dck8xPTlTRpK
HeEzZ1/0ZF04JGyC6b7w+0cF0PJGdnCdJUxDvJdWp6fVl0TpCeYrcN/ABYYL7AUc
4HdP2/33BxOATe1fTB4FIsE+zZtpjy+/JAR1EIRLciPGhdbRwu9APgTdKxzzn4V3
xTmTZjTjxjwnS/YKYdIh10350RkzhjpZPj3LDGGsh/5sIaexDIReabWQVUaiwNZq
dUcvyI7SW3RcPvxWK5d3yKqxNC8aYfHbviMyhinFc+I12GYKaVFZObPxNAzByLri
b1LSrU/AqkssrO816YtHM1XiQQoRU9Ut2mSWPKhEna9B9LKN3ydP4cw+hHhJkaTu
gb6Ch8X5+l/ul+NLJj6P8hmJExXqrL6OmzRcTzGPBuzOaok9s3rk5ovk/wlaSfv5
tqYMy+iw2xGiP4L2RoYx9ODwCYbR3anPh8D2RS5/pmPFxig9ys2KxhhYvR3Y3WqK
G3vVtX+Q7IPfKYC/vtiCEogUEy7Nuc8WXrTfvlESlUjkFriCYAb4PgsitkVWjGQQ
F+lBxR5JzSDhNS5YIcGbyhEabEdOEhqpVG8bnDkLrTFX8qQbDu2tk84xe5hMiqOq
1Ra4/ggJFLceQMzNo7C8Pmvx2bNjY0dr9nHuoCWA/881PSNaK9yuCFGT5CRIHhRX
Penf6M0m3IGBD95irX8NV91u8FKuum8oQ+dSBWxXsqPi09a/8V17UjaikWudY54/
U0iXeqTPtAOCxGe4+7VUP1sGtnNhhUGI1vkEIvgDF2jEbr0itVFPTE/mBev1xJxM
diDXWQi80CmZy7jwncW2kWhX5hUIgOWgrITDdtDkhwPlhGiKGpXfj40VQUF8aQLT
7KFFUS9wyBHvTiNXVVomqR5OExTJGXeI0LVJCWemQbncJNNBYOIQVcA6iwE7lQY0
R3RG9x9yiejrO2d7RmDOJuZCXpF79sAAPPmIyqPxS4QdxZ903aFSGBIejLeT2yVj
pD17BjXBKKmZc80J2/ng3rg7zB9mflmZBipBtaoxKK3xefLY3x3KXj8jfLofM18T
VKB6+8CvblPAqoC+dsfZYfyFuQiz4PJqeO8zLc8PS6g=
`protect END_PROTECTED
