`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rMzdXbYIssGcGN0BcfSBlQahnX+EogWiLnDHB+2SkgR3A6CmVJSM8h5xgFzUnrAx
1C0V+7LOzOfPN8tXeBCMATr5hklWZ0j2aUlNksyTjP3+KFyMDFSdFhxlA5xpD7G9
L1PFxGlGVKUX1izqgvNI0/Diw/B8/lL4GpM5Elim+U23xBcdrl5qVXUCLujiwfwg
O17ypC2DCBCJIJYwxfXocMjgNqpJwM0T9sJsrZPSKutm7aeWEVFjb4+oH+UZ8f3X
RrZ3SrnePnj0fgd+CQCrn1a+TDSxb6zYTJYjlklo2T90Bx7T0EBUxlal7I6v1Joa
EyJUyb2tRDkHcO620qo/WlRJD97/De443qGQvBtmS6Ht3bUzqKbZ2nTWkcgPRo+P
JWg28JzKXb3+6MzThTolxCDuAj9puKv0UNUrZYp6DjZlb9y2GQqZZpV+Soq0aLBC
pXegQxGy+VjChD4y93T1PpNAzH4QNn6H4XdTY4dfzxnUQoB6sbMJJ1FbZblNWRSw
ZWhLEXIrTn7nsyi3TOb7ikrw+8rYfnBd+8+c2Qu4BEh0lBLwkpwbWV/OrhIXbAjk
0ujRopswktpq1s8r1Kkv40nUioDGWwRZHfTkZfjQsVwKUBxXsE2kZwzpevFe0SY1
xa3jsA1WAr+bfws34fpAR8YBJ9PSmLw2RX5Bert7+Z2YCSLa0jqwnsETOzqbec54
mrLHlRcTZnlzYjXQ/N+lTsCDh0u6uX/ujLlaC2fwFAfQp6waIMBMXtB+fUb1jtJL
ZRfjug1ekaiWnu0iyHBOmKaCXrGlOXNlV3/0euiUkbDwOwB6zILopsJa23SuOOzS
dc7E1QOiIRNBfvSQ/DKJI2oB1FJyhSFC/yEi/W64pIXdWzzuoqfpWkWiM33Fzg6s
ETmVYUmddebr9JCovwX33nBEOR8Z5lpewg9FmaXGG4OZqIfO1CNAKDqKKh2kXNt8
Mq8UiUlVGkWDWk7bhVeXrCV/FG1US2Kb/r/0OJNdaItDn1gXMVYMgPT6lqqiWllR
ZTQkot4GQCyc+kLkhXPUG6wga0GaCskU9byrwYUWQELME1MNq5osK2QqPOb7qg55
vVhF2ADgugsXuLoViar32J7BQ0j4m4NC5F6HfPAzsvdORgTfGSKjEZ1eUqGfZlun
YRKorIc7i/WKUwIBydyxP7cWrJEVyL3xMflmK7OQLQezXRYPPVW+biA9Ck+v6kLC
/d8OYzCg0jO+gkWa2MfRUBKmAjRR6rqZiwDMhl3pKFyNtnc97hJzde0erpfQ1U7S
PfTGytCj/qN0ZDs3dswYyM9Ds2H+0/Juw1wSG6KsPl/75bBoYBd+jkdjSdjIMiGe
d/ZHd0ygw8RfJR70OF3bglf4XBw1bUdwBvgVuNuQvA9C9D0+6btVWSqHUp16rn47
+oA0KEL+8EaMKNKHUuEw/uYQj9OWDD0lo3K59/uHMFifrPmVo1/X3I7wYqrOczLH
8QpQPcwzB2F39vbnsqTm7FuKdj6nH2N1jY7yoRzC3A7JBMhbdJbE3ryzBkDfVJH/
Od8utg4c1MwlfZpfpIxU4vXoNjgU3zTrn/+PQYvpORAPtW361+K2ghW1cUx3XLa3
RcPeACKXeRVAsUR+BBSpShNV8MwfjwB75uIjpjc0O46RSuxsZvMxy9EBLBPhMdmU
BUVNeWWOJxi2aZaB6jSq5rq2FZ4tcoRa4B6vLbaPwd3Ru0DQUs+Jhit7VCGK6SpH
hUZmPbMs+M5DgIvv8hMjVixqHWWoM+eI5aiP7ypRBjdmJlAKO5vlnli59XnVQUtj
gy9kr9x7atUYci5fdcMwg3NqQqmxitKAbbQW+naRIFxnrqSz2parJttqQQBUiNXp
`protect END_PROTECTED
