`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HSTWzYPPr9AUkoknVcea9d2yRVsWNUuDlNvVUvkYh/U4XZDlM99colIV+P3E2ZY1
77Ue05F7CxEzd4IoCEmnC/R3vfdYppYT+Q39x8HMdlp++IyFuydd6lKRfLEcKaEP
F1GHhTMmF6Q+26DpF5hBLwljecdui5yjBry/KkgWNwuwZUeerwiDyQw2jsB6UJAo
buc2IKeUtkb4/Ta/+XomESF59X0+7YupUnIkehh1S+SjGZ/yqvbKFjKXSE66LkA+
ZDRN9QnahugZplzbAxyUM2kJjsmstX/NonPX6Rd5ZnWhNnTgpV6Qg+RdP/U0vtAV
+guLeOehfcjsYOV/Nr35nHU6GDVHZZbaPpmcwggQ3aJVHIClZ2gkd/hEh8eP/bVJ
yUHbAqdKE2Wv/s/6oQLhUGYGcD/Bc5Bi7do11Govwd0TBwuogvFiKh3EuA7bTgz1
uhXgnh+foUA2JgjtUOkfal+5tn6Mol+vh02FkG1jygFkPIS3Y1GE3EGzU5AHZcXt
Jc9o11SLNbZV6xeOVKcMDQ==
`protect END_PROTECTED
