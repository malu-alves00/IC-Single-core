`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DaQwJ/74Zwwd+ln/iy6sicABJ5JTMygmrtwGwYI67/tikrPN6LxBikh5sBB2tWNK
WaWen6cwHNy7NqwwR0yhY/BW9BWTbzXh++Ym+dVJ3uS//AHBBc1wJWzrbUh9Bcvo
vLyTMYZJ+7TXhtlSnjLk5DwZUDdg7tqzf8YRNwYdYSOIWuK0gkQft11OwAGDkUdc
9xfxOG3zu8dHAg/E4LuWSaUs7261J2kBaG/Qn97Og7e3YiU3M84w6bjfOMzNPwUW
TWWl/wH/kI/rkC1wZnrJhTWFPRpWDdNuxnm1Ing6VTtW2+O7uYrz75Ze9OdjkeoF
EuGinX9LYxCBiMCyAXVgs7/GWpFAqFRcvOFl9K3a713z/mgyWGN8AACTIdaNVUAw
zYxI3jnCxmdFzsOLPYZ0952iC+t7fPZD2AkulqUXq1o8hiuoFXuf3cg34UVqj+M1
NvamjTNsrErXaUTHC4j1YtsNb66STPGlN24eQVnMbTf2ASrqb+PCf+ieuv4xnhRP
+dF5wqFiEZO6mtgJU+Aehq4wQ+drP/sv60t3rGUWQDJx3U7JiDDRelLjHhPBbNsI
b4fpqREG47oikakxZd/5jTdlZTO8KzljSrSw+V+rFu6O2rVjcWM1pvcafw/4hBpG
DfuJNkWPy1yAmBCgAJOxXwStYg6wkOWZ8K3RdX7GranMYbYU+EVdL868F0BwDn7R
MlcEZm7mgSj0uSYevQi0bnsJRSnXTIbxkYMdwPCGArEM3PS+I6veQfRL5loLbHAs
YjR3gvBgNBitzFrlFFn+DoDpP7GOhILFNyrnW+F5c+STbbWfJ9J8PiPKJtY2Gnxt
mo+CR0Mn4T70+aDIvB/kMWNcgraWXtGMtr7bW6iOIV5G7lj1e4apwVG7+E24SVBL
9vwfQbw8YtR+lP6jQVOk/fR1ob76XKbxFHwWlwAT4DIQEPDOgE3RpyP12PQcCGzi
Yd+Xi8zWqJo8ZAQCNMc8v4e5r17C1E3j7l43UcE7JbByTVL/US4IQ/bAPvQnfacD
FlqMsm+dv9znZI3U9c+vBgaXrfyJoda+tHU4DPb7wM3zqk1fG0Nm0RlF4owKxuZj
QP1wY5rfFG3IdKLStEjDhhEQyhgQMnjkyv2qU8RJnO94j5HUYgl0kEi7xyaACBvL
gdKsSvOb+RDXwP/hUzuRb4NProqqj2iGaC24qmct81k6/L6UpckTHkpkwrxigT6X
m6NTL7lRL1UgAHkl36cx26NGHaKy8HYm7L4Ljb7bw09UtwezMdrlGKWF5H96SN9A
zZ/EJWT+xJMLpgzX26ijfpnvivWNwvahBLuINRWXlTpmop2SAkivwfajPSgLFk4e
7W25wcOEpr+l7augP2aX8uc6SUhKOpB89ISVwA8T91FfHc/TnOF1nMav/k2ZsUM2
nrObZoyAktYNtghEtGEE5aCKAYx68pqRN3u7XXaz6mgPaHuJgPAr/SS90XaTi5i4
2kMqthqieE6p4VgUGgzCWoGQ111z9IXdri2lN04qD2WlrkWj3OUDjY6suqAhrkVm
Zo4H3F423KqIBLXP7QZ2Euzl2wz8PHg9yvH0p4XINE8ubRC5r1owh/IYTNe3M7Xw
BQ6uUXyuoRJIDCtpaiQTwmYgkKZ2fprZd5ZQm1tK//fLGZ/TW1QSsblQvi0nC2tj
9Z0ltKo3x25UCnTlCuT2p6I4GWavhfaq/IaY9K9bfSv1N3qppRIX3R+TNse7kCtt
bbcIDsd8zWCUn91tpuwBQQJNVodhemDOFxudoLouKWOL/tJJEWE3wpXbNL4bZr5B
9MiW8My9lN+PDwv+lViw9hA9EB1DdAP2fP9MIhum9gcee8gc5ZpaWTm++mYWPJ1h
wLQ/1lqYw9h1hKT1ZRzazC4hIsvLiKkB/NdhEuUMqrc15J0UGaQYJi7pwUs+rRKp
mEAnDtdU4VDRfANPmBzgF9zLONIp3MYE9vP6tBUwItWEl42Ydr78Eu8PiTaihG5g
eD5pZkoGCzAJ4WVlFuQocWpXLZ98rs7T2S3E1am8XaSDClrkyNlfcck+0dLS9Vzf
innci8MZ75G599g4lcJkTGDcrTOfLHWtalDl+rZC7vazidAZA4ZTDaxDtzuseFsr
uJj/RH35ON8qAqgpEJCFj9FcGzJKjxM5QOzRCdyCUS0QCSp0HreSAL9ac69C8GNB
Nbvgm+3eDl60SH3JZ752rxALyrTmiRO7lZiDVunpH7u1WAsrCNDqGz/B7eAJZLrg
vcVS3+RKJYVOcvbJmVPq9DL/v9tP9LksYFmnnfMAEE7+HqOvEmaKvf5IEvE7FMRI
uoZ3+qOL5x6+yqXNeCWft9qmTpDdqFPpiCPNVIhYRc1CUJRBvlWhj93EazIAZocm
Iu6suezOde4LPJlcMqs8Ukb9XHTa7b7rBVBgCc8CPeqWtc22x7SCZQ+XlZOFalFM
Qx9iSZ4YLD+F3D1f0Mw9Zk5txuk3PDiH7c+FaS0urAFLN3iP1Pmaa1b5MMwukzhf
DTIfhmHqeLYLOFBKP7Pp9P6GJKkGhyXMdP2YYWJEtJ0IQ2NKhViET47vm6EyH3Bh
YY6JE4cSocTOkMkwAbtSQzvqVl0dPxBpqbhw6H9U7/X2iQVEi97Fkp9fj8VddJuY
LpjUAWudMOQPi3XC3UGQRFkAm7VaFWZObakTasR7cuAlEZBiU7HvaAzVKCXb7yyr
9K0eORWnceF7YeOe07LvTAYyNpXVqOWE7GTNQDVZqtb6Payk45kickWaa2ZsXyKx
`protect END_PROTECTED
