`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xDe4UslQlKBmrBuBnJSxsKLAcFdqJ7V318J2U1MqDFDiAzewel9/dkf53swYWo8c
yGLTuSiBc58lOv0q0bmOGiIKg8oUDA91B5KE2Cqeopsz4YCpUHdzvxtJGiM6WW7w
HQ2uFNi+k5C3nL7QN0286gImRnOYF7oTnV47wJf7yHlAX2FoNujXS1HeRwgmdQPx
woAufGV5zXEytlZm73iJ9EQ09jN/to6NarvEXyVuJ0aNHWflM1i2HWYnr1pax89R
mU4I6j0FubBW+kwmWePowFe5VURzbWRxI2IvharlF7c+fzhraa6El5iCkt5BWtss
Ff+Nc7uE7+2NZqBzTQFh0CnTcnzSt1apUg53NJntdNCzhKA308Bioy5VINtZJQjb
iYrnek653lFzTp4dTTtDACpphFZYZJ1Hxef8kVAXC195Ea1+JKgDyZhAAqdzmMtE
36emCSNT8C2e1m4X9G75Vqz4WTe67pOsZibyybMt82+9p1f92FKbefuDjhn5u4DK
UHpiLdJNkZuFV0dh8FA8Mo9iKca3pB9TAKuo49xiJs/g7lLeKIgDGNYe53fiaftI
EStqoWOe46aXCNYMFqZnCtqvy4r4gkYHZC0jrT3fyvIBYFbAROPoy0uk+zdsivj2
NDibww9WJ/cl8er6tLWtw3o9DS/AIr19Q3NotHkVq2qRUct0SRM91qKTtCtoXe8c
kF9n+ywRmudVn180jZOLgALxEXVhqY1KyIT/5vE44cYRE1Njsn6gt+Njn5SvtOGq
2As/f75NdS82DQFWJpTecB6mJpabHeiyL+G9Z8TP3hcKt4LibqaKILNq1x5wsNRO
XFh9+5VGyX4qF1O0EDioapsGASg2g5RVBKO6uKEJbE1B98crC47rMHQdssVSWpPD
xhWG1N570VGeaCPmIqKl2A==
`protect END_PROTECTED
