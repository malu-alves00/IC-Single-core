`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oAg+bW0OnaTPntOBYUYnH8vr44kjBI6cQrZ1rEw0HPG+UfbmHqBtQ+Dvirdz4H+W
dm/Ol9NyhP0avbOaCnIiJdXOBHjlLogLW24UqYVziWIvvzncIVfLei688m/lVgsx
7F39/WUTsGbPFovRH2Ka+5u0TQ03DxLrGmw1vh/wdfrhP5xLGqHWWTfnRfKPidva
n5+r8wu4RAFJye8IHWoLhcnyVZEX7w5Hm+Bo09E2w65UqXX3hxNjhmIOhAP3t+I0
Xxgdy5SyWdyBB0iRFrt1iYp2NYGg6uEEBebWRSQYOycDUk8wCaxmBOOqAQz65/LN
ISUvZu1LrtCKyCA2kgTrgRHupMuUT5XFIVMZa38EYME8uuxO9StN5CvdH0dnntCD
suEQLtrzLl9AWRwXRawKBmxD8cI57I41rILVDf+pKPwVPO+7Mpl6FD2COBgBX05a
OK4t+BIzNu2f84KFbuFCbyebHLJCqCiuW9HKpl9/3mvWPHuP0hBwToOSFJacMWG0
Nzpak2nAhg3laSdfOto5CP+q5Qgh4CHi3jHORCGlgb1/aNs0zvDWoqfcayTiuycr
a72BuzlrKRsHVoTlfS3GV1fvtPb6hTQmvMdSr9XFEIrFF6mOUlCgmI/5+uv9iOqO
6AAGA6kNh4mH2SnRaavfqfhpGI4zRMEgVzos2+WIki9FDAuLbHmPcpE6xbIO58EN
Z+A41/3BNJaUEt9hGbialwZUw8gYJrz2N+ngJThIUkQ=
`protect END_PROTECTED
