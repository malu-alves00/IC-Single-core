`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NEhKZ2F/Ie6Ts88BxPitzSy12Pkifaxr7FYkwNAuQ2xV1Bkl4suV70HdmosMdm6Q
IEAYeEETfYaOiVnr4McJ1OtIZ1r4hcHVl76Ketfx9e0+KtQbmoDf7aV9nHCsvcCE
zw3bnuHzsdfjXs5SvIkwFvwu7oI5oJrkhxFPtTvrSs8/QPWna+ZQmdF0Fe0B/koS
RZb0glhDr3pC2xGW4DkIFehHkJp9pZ9mtnhO7nuVQAjNemIq86CduxNZxzPIPAVM
DqobXv1IkMzd1IsHqkpvieVEvZUJNUNLrXh4SvgYVN/+RRhF4Q4NWMY/aUScbLtn
sPJF3lbcp48HI3bLGm9LmbgzBSxo/WCPOsz7R3G62oK2Bp5nv50JT3B2aBO39Gj6
lYIpn6w+5iXiIjYC/Pk/47dSd/9VnNM93uhNqPOE1gbWKDCo++1u2o83tKFIC1WC
jaXyPmQ7i1CgWCusQJskv/jMZDOWfKQc7mJAEMVrWgGQuaF6JHszzzPuvyUDmR6R
3KcpHR4HbSiPqqTYOh1OMLq6xIx8rIIelvCjEnYmUmx9Cq/Pw51dfsA5FZWF1l3t
lXaLPRr7ekO9IL0qLjzcpf1UrAjFxvbdcROOtsGxW3L5/zNZtSo8QPcAC13mD1m2
PiCZOj7ipe0PqcJVvvUrHKhF0idNmI5ddNPhpovmDX6h8LN68nbo2pDmTSmYZWDa
BPLvIOHg10in94AGKljut5/0FkVMiytAQDD+ORXJs2W71PhaRUCT8MTfsE7q2AJR
Yh7eBZ8UwSDaR1ScCu1bzPE7q7BfxLNjExM3+gcQCYpF19VBhxDYXL5189r9qCpR
GEkSbgpI+EkwwQEy/y2uudcsOe5+U/luLRYJwdfOerEhJhxOVBiih9iDzb/VGaky
t5MaSFo4ch3MwB+iQf2rF0itsfX8zJ8bUPgXRROePz/4v3VNvqAdpidk6tfoLlpE
Ijt89ioPdUkJyBtamlDYFI6fAGAh6g/HaafJTPzg55xDUu6sXQRtNtJPLFcYM8k0
6HULfjR5lRIxn/NrsgZ2hW039MamZr9jhqETkqE2wnlbf8JnMlZY1WZFH1KlnX1H
R+vvuH+Zp4FH4X9//Dp5gL7E3kDqlXw91MYmkcQhJlJ9wQ1m845nQkg9/kEs5BJX
NZxJomricW4T6T30tA9Jk0PW994Kvkw2ccP+gGZHUN9ZZnHY6MeOOAbZeUpUi0s3
fzueMSCY4IuXnIXyvqwy86qwPo2rhtp0aFCiHo9B6BYhnTqRbdKZXFMS9yiF6Tk1
LEx3sAqzSwGigRQ1tHXrrPgVkxKbkqTNYYccorADpK+GKTPLA0cNUQa+fyNpCoIR
r+CtWwstpl69ITi3UEkuVGb1Tl4TLKnc+9QJXss5eD2ltJR9kboytJ7ByUd5VtTP
ySkDBKSq2+nrKRtAVvDSHHeT/B6+UUqNCWZAmawpFll1xbggMZR4r2+wxzHtSDUZ
fRks08IEejLUUG9jVFtDcnPHE8oJEke99lD2VGyHqj76ugoeMeRDS/IMcunIpbiX
6MhTAESsf2hcIJV0TjUa7wDygoMflc++S15ZUvT1QJ9bcdawyJRLfc06O9YS72Pj
jhxe43Y/TpSWQzQmJAPR9hey/rjK4UnnL1toc1ENJco=
`protect END_PROTECTED
