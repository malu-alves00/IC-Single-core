`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2EqclHS1fqY0Qekt+NQjBnz7rajMQlgOxzJ4saVaPNdENn1DUgcJ1ZbuQexv8wcf
l4FWfoK7dRi0CXvLX8HLsqtqCmsPmi2hhJQSY5lWlH05oTuT7uJ3SALoHyi07/Fa
pRe2IISmj0o+mIwNVhwCjYRyaRUjnJGri2R7NY4f/njQyJ8Ibf9Nk7Yre6eJA6zP
zWMFs04P0wrqa3bJL/ODat6LJ+um0ndYJ0WztvEPN24zrF1T4VkzetdjlE7Vw92i
Bl4d0WCvvf6Sv8rcLH75ljLEZpZnSGq2UF54TgasgAW6qheOM+TNrAq8uKxtu65I
vqUDQGLjIq+00fLJZmrzi52wC68lqP95LC8TEWK5DexF0Hp4np96XzJf5AinC4V2
cBt1UOTYbfxDg3Z0aDt2g6EVpkUlhRgWRVQrATUyY2ZrWqyIp7MqYaPg52QvDaLa
8L6LaHQ/Xx58gnqqlTARDZk1HnebTTAo4rrtUlAZ5vm9c9LWMrJNLgfZ+oQTam/d
usrTNnl/g2gopKqb/pPcJDvb+QdI14h+OGcYnG1UwUepQ//hp/oiI05WL6Ac795S
OLe4zf4BdT5JcORmBDPviLUUBDwZnUqV+l+53azHsfSaat4E8A4EjY2uLPpt3wXN
rA2l8cSCb4a9oUHNeagphmvAOZ5gxoQjWjNkT+A7ctzhsZVmowxMMN3f9SdYTfdN
2txzdCBy/0JwyL8Jfh7hBVvldCas7e/sV4X9MJu6VVUQxVZlyJnhFchcI2b+rZ8t
G4SAH/ddqkW4rWpDE7ykgowOi8E3lRkWTL68o+OUCFA5NYH27322LgWiyaRjRm4P
aOJDoYmFdI3bPfz5FCUWnlcuIRE39AkBjzSKGh2HFIjYcY3OgIrhy8ZbXYD9SG7w
cFTPXESH2njWy8Y2pg+0odcwlmu3e7LEDgjp8YYcmc4=
`protect END_PROTECTED
