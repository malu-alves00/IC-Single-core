`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
H2I5bhZKqoj26Ljk3JpsghepMgPkdEQNm3HSEHdJYcHz/w49a/ny8Rv6d1NBRaC7
z0DyC1lSoKUQ1Bn7S3UysvtkgkCZk9awjA9zd1G1NQRklCv0/kiY19VvcM1+9Vym
G5MrSCxlXOzLtlmQNDCFzTcet7Ki4WVCl9JIjT7FK/r6hVClPZ6r7vzN/g/VncOm
mhwp9982sVJ2ktnnrUNPVlhZKaM4GRmRjdEow4CsAflsQnApu5mWNr5AjzRwWAF5
P8hT0+Xr9gsQDtP5Vunra0UsRcxF9wciZhjYfffh1Zh8uJ8u8i9Sd72CCxYHUdlt
dZ06ovznUKazRIg8xoLEH2ibs1aQ4xb6+aX+GRbOjq+Fn7XxH7XEFCWjHwspI2u2
ig14K8MqZqLY4IlESIWfswkT0CiVNizGUTqSeC/wZeSDn43nAKbXsQMl8n2eLjYo
IOkGWnqLoAgOvPOlm+7bCPh7ChREVnfgvi4djQkD+iCEkRmlexYUUtnBjPimNpQN
WPy52jcW19xQqw+j9TFnluc8txBlRfy5usnnUW2I4EvxYY3+8da4+n95HX929zP5
3397Qo9K5aQd8zjkIPjHCCffhRBZV914FPGgKehLsIm2xe83ZdRF3JaeqoANSUft
3Oj/2iO/GuT5l096jl6POrkt6q/mSZoV+ce9RplK3I4xPLJNm7Zj3CB08/8IHRZ0
x0CRXzjv7pD1BwzSRTrWvbW8COsffEwdEGyt/22+0ADOLoE0pKR8PYkJQdPdS6cB
kKRV3BEiHHjStgjAY5cAaiBUINmY3Dnb6a3wYLSbMyC89ObNo7eR6n+BvB2e4BjS
2POe9PI3cnVY0+Sl76rIMaaCdb6SsU3BJobNfZxqnzkEcKcAztzH83Kv1crciHIr
Nx8e8H6znO7o/sexuOvcTiPALKQZ1H9iiXB+KVeJws6MtmDkobdv40jQY5Ymc/nk
ojJGRsPhG+v+O9lXi1T9L8IOfi+rBJXzMTkuzfuDfLHkjZ4P0etsi0mqPiq+0wLo
+Jekg0YX8Ohnqt4+4fWUsIh8J0mQx5BLd9UjfSRyMLjVFRYrLoqmGz9y+oA4iSZR
tubRH6UoFINajOuwz3wEhQbpyplYBXUa+7T70/r/Szkagj8NgWAjoU/fRZs7ePRV
BetI9jrcgI9XrAvBVFh0UZjhScAHEn3B/cDp6Yg9gZk=
`protect END_PROTECTED
