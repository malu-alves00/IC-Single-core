`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5H0j2mbA/DUlZPfjhGEmXtXz84Srcryyk3OVuOWQrAUcwvpoOPqoTkHuvWq+IPNh
JqlT7VZQq+WMxnK+OHAEPGn/Sj3eBYvqq0ZxDvIdOTdUPSWKPEl/Y1F/WKq6kY71
Xb28h1eAHBjQiGXsIeQEkPDvpMo2eVMndZ8vWPPMywPFOxLUXayiAuT4JyNe20Gj
NBpGsT34x106xF2bfk9SipX1NgfbpLYznnajtKPu7X7d0sqnhhVZleKnAqQbuWs8
AficYSs5xsFRCboPUy+7Xh0OisA0Sntx04OylXZFWPVdWHmK+nuTTOaWfLtB8t5m
njjPi3CT57euR/SC+U91bnaa2QBPJ6+VlxGzxyIVv3lP5ZJhebXKyAO4nRBVpDsA
O7+7hvkj78a0WosRxQzUlyHxRaoXKAfu5baqHUMAqP7gCNrDLvlOi8NpZiU+UZU4
tEYVzPGraaGOJuz4PdkrTSE/QZKOLz4rpKlaBrE/lm/cl7hQG/NFx/Syv0Juvpg4
y8RCByXeZH3q4tzZAe3Ox1s7FbVANn0eytvx5BSkcHMN09rjp8feFMQT3sipyZBE
AYMGZkD1PFSjYQrbElR0Ts+fntCA6yr9tnuKfBx0A+5j+iZbQAJTsc7khPmnSPvY
xs0wXumjJhQN/K4fAdMiiBJHumN4S8iYlxHN8LMWy4uPMM6+bQFV9c3HjZerKaJ1
4bQYrlb8f/ZaMXZuC6PKk0tj6iqOo8hx3J6W/tF/k4vUQU0rML93T3Te3WSDglRn
asuxddTZXeUrL0KzlBW8pGwMcUgCczrEWxDQ6h/U27CuH942wadtd1RyYUBM+Bpf
pvv+DXgNNriwEcImAhRIJFPQypSheXWLoh65rX1bFsybEptOWrNLe9St4Er01cAf
bSJF4KrsDBiZmdnKB0w2bTTYD7ytqbASmUXeHLagUoIhmD80IgTMrqWr9orJFn32
EYy8fbSp7KPJ4L4+UmgLP1WgHXkx3KI4jJQsBCMhwtFAkTOozRluLUGJU853BpKE
XktVwVzUepJDI5+tSUIBZpPUzN3iZs2PTks3GAhhrZBHxH8FUGF4t0UjxSVbY0Xe
hdVRAdp5qlEzjI+LX1dSr/TqcbSPoaA9dX8gKS6BJWUxv/dabT/OX8xTR2jZ4Rxs
SkEMAQobxprHEvYeNlq8PFWcXoSwXL3MlLfda0kIiDuIbYUecoj6sboCzCRKmjPD
IG1eo8sqcMPcUXGuQ9Oi9a6LsSqQylofFTjl9zAbwFxOA5JZ4kW3Yr03KD7fAibU
RsVvSnPwXM0a2pI1Hser2I7ly3bhnuxChmZ5lVqRXDRFdfDcVuiDbIfjAGhoRc4n
WA7LDTiInQModuzEVcQQ+RlNsrxokahAXKb1I68BTrrHmdeL7HwjoD721Fo5EBR4
+B/uSA7LHnhG90HHmRC71+Lk9oagUBPPFWwOf2u7uOsoBbmgbeU7kXutB3josH3m
Up8zHuvCXnBwpZUiNcZjuZGqZrTOgxOZ7oZ42LZmzR/h+/vOpsp5C1dEQs5RUVRf
dHZCDr/Bx7qbaig6eeq37G956vBOpsz/RdKzM0KVy6wIjhv54WTlAhpxQGFAwVl2
coNwP7zyRd27NYYmvxQfznSxYjOL9HXMJKmkuS1c7lXr/yEQxePvvcnJKrgIBMuG
qBdeND0xAHjwyUmqo/zgEXy6kPWrxv6p7pVgv+Slh0oSUbGY5pikYwon1LSsE20E
eQh1Ky30jS+5tHm0CWFnIpGwcKZcDECSmTSpy2n5VcV49y3PJz5wb4aKpbZCnAO5
Y1/whz//wfbnpJahsElQNS05E/vcuWg3Rxc4theO44+JujFAcSdpXLp7rDFZvoLU
O/V6uTh/JIQYgwWjivsfcZIvjFZ3qHrwnaJovRRxCAnBj/+H3D+ov0ybE/zIaXtn
a/OCKNxbdEVAvlJGCY6C0HpAVBQrwWB4vnxYbVCSZNmh+6PLnRa2wVwHF/XFXHac
9MQmZET4b5ABAOSspOqKwL29Qx+n/b+X4l0SGgWTVryHxNtI2NLeWPcFjtgx78Ph
U3PY8oKNvTkQwQWL1Dp3epYD00Z0QwI31cO+IBHYYSRkGrLgHUHQ4HMUs8Fgp4LW
EIcflnFe4JIOTJoO112u5Cy1ti1KdS6fcFgz/yNg7x27n1REHNzmN8hAN/inMLAz
GE+eKkr4jyyavOJWH51XLosxEYq90FCiP5K9UFDM3E6cowp3k9I/77lGR375aMOl
TJ71d7nSZHxyes2XNfAa6C7Nc2fJNBjeWPftsCuNmxE511E563HSI44HHU717Zo4
W3ZVJl/iuLcjuCqRK9HvqgW0lNsNKfjzmkszGIqT9tfx5Xte8rDz1NXRoYpR3kbt
6kf4HLf/noSI7dsnL5riO0b8tnx9mqqvd2lUlB1PBRnRJqQvwAk8PgNBTbyU91e7
BnxhLYWj3a32BYjWfehtj+eSHg7RPvGJ8n9yRo0DLfN21k2QJCJND1dYZmWOjOPN
XJCFDo8vsNO5f42zAlF4U7PGyT5akdDPsMuTdHqWkcjAMc0MqDVw2IIt11ahVmiY
eInLtVb/8nq7rDpMbogJrRhDUVTwmL5p/XTJsb9nob/7RRvyZ0YAANPML4TjQX+8
Spiq7aRialI+M0gYqeqd53J7BzmF9twSKvEzDxzgrKoHcPkNWGyNdDxMMvbuk6Ly
K71dEn2jHvbl/DO/MetPz6XO/tbazSHC1fKdHFdxRLEvSwtCioLxTnxUjmyMVNQp
7MwYuRsjE7cEmM1U4s+E0gwvutl28qkyXp5k3yCiD7NMWTvRqrpNNYDi494VCLSW
6vtecua9MpWxPJNzpXb6ht85S4rDkzsY0RPyqz6hXIlMKsLyHgrkCClV8RdmEGfH
QTzmLPlHcPpFLSfpfi//Er0JhU9nMjYJ00nEo95t7Rcz2Q7WLDX+zIXdQBqmj1l0
L2/3Ne1XuVqVseUCZkFc1IBaPER95reIFpZ4x4n7B5MQjbKNc7Kf3uEQwkcujwjc
UpE52qYAwUuIErKzrV9ILMrvkzQj9Rot9RdYfsXWosFyngBq59wNsQoP21MKAZ95
HUloY2xQ5n9apUXNF3dpjvcXh3cYt1iGMwDzN5BYicb7PheYz2dLTVSXXa9yH7NF
V780zbZuZ9pH6oco4L/KBz//4x6AfaAwn4nr5LOaZlh3/rEbdZXbL63hpEuLg7iq
aGp3Fr32jiw90wPDDPXNmclUYYfKSfa6Xf0gQIjLgJbzH+wYShLezZnDtMYyuid5
b6TVQ77rDup/mzLEoyRSSO5qOHsoeTCM44/auUlqKn3Hx/iUXG8thedW0+jhSSYx
j9N5YtEk9rBJrY1x3HS3oKrTT0d4XQnpG5oRfXtUHtslJwtnTh0JxauTPzUbrYzM
g7oDaWivYaCtjCPXIj2jjE7NoViPZTUMWsURHul4q/+B/ETb4QlEPofjb9r8IAZW
FXmCGTybdeJtMOWgvpzqIarqZrGQkj/dqlAOt17k3AoLOp0j6fKoaO2GBV0xuGA7
v32xXOHIkYwMoEye5IeC3Tc0bhzyavzGJFQIjP/qYnnriKL0tE0Y//Im2rvSogJb
oguBM9ZG+4bX3mrbpk05t8Z9/nqLXWjHxkJAR8cPVRSzGp7uoPaEZLKQwawQqiel
MkyAt/9c2kpM9fxDo2czYSzqk6aAWwyzTxFzAqK6Y7QZWwpudop/wGtx7E52f7b2
m7nxOVubpyMwAWORuNL1i4sMFAlkrzTryQ71gy6kmIC0loLakA1X0gti71uSEDle
oC3nozlOclboSdyfpLhQm/rV4Tvk6w45GP4R+E+v8tRgkDUXsB1+kaCsOvtMGilr
YfdjULZZh2ylZGnT2Ku6Pt8HGJv2W1bf65XczreA+gHSytPkKpp0/W0MHOf6lFJl
7aBAhejbp3XcfM4IOBBd94ne1qpcKKSXh0pNPAtYwZRbEmFa0aBNFG+BnxkdqCzV
DD1ID0QxXPJshdnS78XApz4DJHPGXISm1zg/8k7YwDUcJr0O52DQW5IbWdCcfLuY
45D8shtCDFy1xLPU0mNEgL/PqUMPX1E9w6cPQr6z0d9l7/DzQ0vaEiyjmkBBw4Pc
VJLVvUq7o6DsyCDhimiz7HajYOGNWa2N8E6f0xdbRQqTBx7scQX9VtCfMGhynCEB
BI5yzhATQ+nucsRGWPfhHUqi/bX/UkwgZxCmMbpOyEwODAxlO0ZBiIvqHN+U06Qk
+OA2SvDX88TdaQN7AtPn9jyZhlhddrbMpFIGkYIYbLImt51IQ1CHebW2aCsDb5nA
PKOAVeCmTYhJPi3zgzlJbGQJVcKjwG15dh8fo59Tpt1nSl6G/IsoKlj8isyQaLr1
YmWfuwbkbAwBgq7S2wqGyWNUlMvG16fz/IQT7KSZtJwxBQ8RBuZId+s69zuhIti+
jin0IoHHUquoQpkCe2SCNFXf4ED8v5WkNSE7rQAfIySGHKTOevFNhbDAQArsGZBw
P4szMM06nY51rDrZu8PKx969e1EiN/MwusOJFoesRg+jXelAfb8qaWY2Fu56k08j
5CTFtXdUGq/usYszb5HYwAjtARRrGsiIuZ2IxbRT4bSzcMt+2jvhhXfPB19bhZvI
TDMOLvROk5/Fj8t6GxyEoRo4o4KRQ1Lc2js2x+zI+ONuFr9F5E3k97QfxR6kSH1S
n6TgCuEDC8GrAqCGEeCb+wXGI8iAKz/2wRh8kBRNHBTf6BDipyK0RW3S0KoUIWfh
CvYDkB46DMhkq1z+D+dIoT18+iT2R5J7RvpJNMYtaEQDUctwkOqVw+v2OQEPILgq
nIWNHR25pTx4m2ACJzd7bebYlEIy31zwLHFSIn5hj1ms183tGe+RXIzN2CyiNp9j
io+sMzM5sXJLbC3IAsp+rSuwN/MG6NHtCnHXu8S1QcWSRi9WXDf1OeQhojqsNLCg
ReF6lnUbKjywkwU63GKARmfwyFolnSlzMZb0gajO39P5/K3uqJm+VETvgS0CQeca
`protect END_PROTECTED
