`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cB5baGd11HwGwCWFRSFiEb+1QoJvO7wn/MRiQX3I6GqKnhc/OL5b2LY6k3ISXpFH
wJmlW46SY0OpICAwhwzMg35b7mWWpfvl01PgxiqoA5lJg+FCynLhj1nGHg3ZRzwi
YBJehKFBlmdQS2UeELgHbjDhgb5HfD01uaOLYGBfPJV/QcueBr00m86sH+wH0hT8
+hv8LvuEtJKxtnuz1ryFZ4nJOEvdLqMbh9zkeF0KMpUanryMx/BF57T2bL5oKmR/
wsqMWW1etrHphVF5gZTAaA+/MlzfA7qgC3E5ReFJ8WEcSYkpjWi3taBqkdQG3L03
dg5nySeKI6IGuR5HUz+BpQgzYd8fOLSm/o3OJRxG7jJ0G01Q9wp+j2uDsZRJNCpq
KEHwwcHcD74oKdW6UZmPm72LziviXG4y9oSfnscDlQBZTymrn8HQft4iWi8eeO1J
WdjTsfdLvaYSvhiToj2zJWm9SzLAbKKdA6YapQXjL4I/3CH42lo/W9vncW++OrCP
618DxIBkDs8U2KjzRT4g0F7iokdRq0iQOa0o3fV87UshGva/qdHGXXykkgeje9od
DXYExynn7L4OXNq+IYLn30C9GZDGxjXQAIGMAKIe02yXxVNSRmTUQnThDFDr7XsP
QBdatyuTt1m1Pfp+pfCNIDwhBRJbT9O+MtcfWhcd1niDuNh++zsSWz6ZxJEF1xIf
vIesH9wW4uHSNeKuoGkKDOHfAhwNNKs8R5my85V2aGHLG0ASBFPb8Pd6DXz/azSk
/XQBEy9MCDAYGm8TF9WJsm88VtC7dbrJlwWStTizRMLHBgwGEtIoLSmLRM0D+M0B
4Y0SddbccGoSSVP+2b+qqUawk7kFGNbsozfdDNs+uAqySHQOpjAI2YiV6b/3Jnf2
54M248OOM7iqNaOvVMnQULbWn76K875YZl9ls/1qBxBQ0g9LGllxoRc4WmTHLSos
Sdq6afqUUHGs4p3bobMJ2VE55FZ0qfnWPImMuHSnAb9FRQPBppcOChGGBaLTDN8k
AWJylxGLXmBG0PMvRBtGI1LphTtVisvrpW2ff8SzXA1eBjqDYz+dQzYZIaOrq40W
b7SEdSXTbbbiuaDAQC5vF2NPko0oI2CsI4QEDmcYVCIyD6Swrc3TzUtETVti9uTH
mxONlkmLZjq2dcysY1J+oPsQN8gh6Mmd4Vs2LkjXFp1el4ouFl6FluAoqQNYMUFz
mUZwcFb0waDsdnr0u5ayoOBotMz6UOO8/ptsQjm6TndZ6jvFXi+UsRbQJjwFyycG
nDe8LbU27spqfIpb9dR7KPnl3OqmSM5SWZZn7zjtLWHaPbv2ct2N8ciJJUEAOCjU
miCM40yLT87rT8eq8GB/uxL1XFylNVcw70vOuoajmBNq3vFAEbQJ1rewnKjEkL9/
z12lh6mlOgUGsnKzaVkBt5WG3dCZ9ATXvzotrk7P4dRQ1fsF8m8UJx9Q5h8XI7yS
0M65vN8aDPUwABa0vVASYVhnWHfyW+4w6ykKjw3ZXChuhHIlRCFapnV0AGOF2TcG
wF3yTHV/dP2homU6LFeDT2TAR6FYKPPq8k2FzZeSWJA2cuy5PkR00TlAfVUhGDDl
wiCcfqwlyMTOuK8ZxbgBWB+23Zc9FWlKFhZn7K8vCqacLwjCiUOPEy2f3hmR2igZ
Lbdoz61TVd5Q7y/Bxs53bHg0uWBbqrSG6ZXrM/d4YRiSVYcRkTLUKMKEayCnWudS
bDd+m8VZuFYDKzV6CQiROvHMmPiOhwNsNjCunFZ6JYmeRo7xk/rjHxJbEjv5uBQJ
bGrjD5yb7wW8UVoFDVGnPWR80rtU9gQmBmpqgiI0slIKf5sbaOg2v8Fqwuk6H/qQ
PtT8TkMu40jAWqgx5ShQyx0zirxE98kC/cSPvRpFgB21ro1ITbL4jBLWF2N1/VZ7
F+2NzjsgdvBZxIadvnAxzYeSzXKw71UNxEXf8IzWwuNtGIs4OHcqnK1eebIVlpri
VuX2i3x62XwCDmMqYG2AVhZAp6joSy1qXT8lN4lxa26c2IR0YcGtTkokyn/Of4iM
wZT3KTO+fOh3B6eQrIQJc5CxcWizoHpGLz4kq8Fe1dLoAOWJfgvUuK2C0v1Vz+Sf
zNgWBkFmcn1eaU8Aaq5SkuEvGr0mNr+r5NXUBdRgwPO8daRs8mr79FiQvdNIae7R
9SpP/TufoSBosDoWjMVB3voYurdJPkSH0VRy0kL+AeSL2nIMSV/WM8hNPfE6SFrI
tl+HPsjWC9bwK6yIo5oV07clafOJ2d4ol4uCBV0YYm9R8wYXTANkjjppSMKASPFP
1xRntoFzyvH/2i6sxfm0QvhGx/IJlVGrUJXVeNAR5z82o2zvYQvu+Q8pJM0gF+vP
XnYkdbU1DCDrwTiVS27qnUT3DdRm0HiJBFsZVgHkbVFqZ+/qSvcV/eVndyna0X1u
HW4xRK/dJ+W95a3TxyKSvzSQ+s01xvFwlDqvQ4w4nzLI/nYyU8D0kk8cjiRXUPVR
Qx96DBVsqgFZxSco5fUnBOFcv5DT/n67lIufNv9+FCE=
`protect END_PROTECTED
