`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
J8ytUs+R3PfB+kCDjf5p9ZssNC2riJlgBEGKP8ByvIjBShvz31mpwkFV/Z6L+2T5
NsIxFsH8ZKrLAJqNwvNWuEB9fwpQuMB6OHDrZVbepByCZUmbl4fC/uTIR+gT8vpT
YoPzdy/njVcp0Ytrr3VZVfqPWxZ2YQ5ivSp3WFD80UFNQlKdj4+QwBqyoJjhTfoy
L6uqcAAK6qj5iDRFMcn7+DIjwq6fHLd7J45TWDw9+I1Ic5VKOewCWwhB8IJ8Cyb2
Z/73O4fMp97vpCjSLFXf0LbVjiIvpnYwYT+Ikh6ghAldieJFz+0J1oj9CoTgRsYh
08pbeMrKbVPokdGrVB9TXGadFIYKA0kZIfEJfKwxxwdGFEi3ouhUpy+bretXtmVu
Q8286FsSggBU25LZ6Kt8MTU2f53hut1yYHpPXhXCZNIG+trVmb01ELPzW0PD+ybR
W8JtudYv0rF2z5/Dia1S/lDbuwL5HpSvkJlqnNFhyOzP4RihpygD/fXoW+Nf4kSy
JGWk0FfJoN1G8w51A8t9IttRqzY33bV2VsR052XW4qZ1nZGguxOVknqamVCcrnBd
9jUNdP0A/CyJ4Al5mXJC3Uqv/9QA587FfV+eAlIO9+cUrVO7Y52p9PxXeWSBa1j9
hkIB3Ef+IoxnSNzjtvxZ/ermau1lXi3VLekkLK9EJpWcpApWsCdIjZuvSQPqyC1p
mHqxUPpcYUcSoG6kjvIZvcEa4Ba1QG7GZO4bW2/ODJU723OQXisyUJi4zmO3T8il
l8v21+NfXh0rUjGMYdEcQ9a6ZpoGGZRPbzXL3uBzoipnjEY1IUGOsjtgSaVdooTm
1SfvUQOdUzLFcp6Uiqm23xdzC/Tu4Fws+FbRh6c/AZ9oaoHQSWFQFWpBLRsIDcNV
4ORPtQ/Bh9CfbbN6FapZSwTIjSgCZfoLnzVaRwmYNv1ajQLQVN49jnsPIRYNxZjd
QQcCH/KouusZ2ay0s2KR2IBh+RB9iUsBMbSvEkMRQUvbs6qK8hQOnNstv9/6EP19
Iy9dlZEdKnASqaOg6WNTSzChkLJUyYnD0JIcsTV4F93vU4kw5cb9P2f2fmfwqn1c
j/L7MBq3Uo+PPXPpWTYRUy2Rq+bUJsqMWyxPMznAxrazolEtkvqJ31KdlAVKEc3x
ryGvWcp6/1p4/7ufhJixPVekiEehYXPdNoP16Io4yzCldkIJUlFByC5SqfU0jB+t
ZGQYM6uqSWRxw8oUyM11DvrHN1GRHZD7cb5aGb5hf3vs7qzBTVPFdDk5O5eYbEx1
FW6y2JsCJaiuVoS9RBFzR+szKowkkruNMFvht14fRLlqT2RJdXKRoHAU9hnKlIEq
ChCdycueOMqVQT4qwHjkhVWBVMbBRNuCHt5L+7agyojZHNZEvGXlXQyQofhSgk9m
nN08yQRn8lcN2+W6aYIj+unfEAu5F3XQnwttGNGeUtTeUts2q72D6a66R04ibMtg
7z7eWzd8l4zclPa5/SROUBQzlnTGwnjiQz1UNS8mVCZEmaj4Ig5/Sn7GJzoeLLLz
2EY+8VfRUQyxsMYUo2mimvgl7d4PlaqDT8WsmXGoql0WKfX/ezNLwEu5Jis/C3FV
naeqeVdURwH1SQxhgI75Tl7NY4oK1Kyamsfq9YRTehk9WgpYwOwYgNrmXFKTCcaQ
KWM85f80cEt1ZFKiHdQPKZj2fSKjWzCLlBec2qoNPeL+4VhkeSart/30Df/uKFAe
kPZDghGva+2e4KKdMs4sZq+Jc1Wx0e7XM9SV+hhTlG8vdH7cstGXNahuSn/0G3c1
70IBd477ogUggIw2AXva109Vs+yPtS8/SnFD140arhPnqcf+s267S/C5mnkxzkBb
DCSkYhz+ZAEkNkZFcOrt+1oMXlKu4p1CYLX7d1aS6S25pZCsS4aI57e7wrDroXz/
pUtcpT6PWAqEv+vW7CSlBZDBTFjLHmQ4TyGg4XZXCdl7pVG1rzQWbLSrzwbj7HdK
/fKh/ig3GwSFuzVBD717FPkgfjz4sufMqLZ9bRL8yLk/Rl59WnxBAhnTREldTLZl
84zSCY0VzMjr9foMTyksF0Mgjqg2DzQ+CL5wrv39Uxs5HaC3MeVUI/QVnMR+OzSP
iS4BrdM6kX2nO2k1EDBRJL6RRH92fzuOTm6VaO/Tgv5WrQUCcmI9WpZUH3I4DC1W
n7zNSvHfA2GwBPLQ8YhA20pxWOfHS0o5VDy+DkO62UPwNYraxHXXWesaDWvUj8hr
bXoq637pW7ByeY7vEnO9Z6ASn7nJimuNw1iwInQV8nMmAXGI0JbYNJGNHsJEZXX2
bk/rB5v+x00fmbyqj/O1wQHhamVyQ00IlGT0OZ7E2iKlo8GfqomJYjkX5l8aZd2E
fyYaHhkvDd5QVZDmCm7+RHIJTHB6gunl9tlHxNM70zO1pfmahUtku0oBOQxTKZhn
LP8O7TP0ZgPGrdCDP4DK1dRzlRLFd80Jp4aqTRmkwWkSkwDu9KMClSI4sSgtjPuj
4ukHdeeBXGUVZTBeuW3/uQmn4DfMVB1/gJy/9GAtL4dKS8uqusxy5racxOgQbS+S
Mq5wguwj/Rgb0iAHrRmyzp+YfUQWWav5q4Z9ckJmZa0dYucJiuAlwVTIZ5nKk08x
uNATrRdUlG0s/5wbdE2Ds91wCLMDrmV32zd3VhfSPV0qZZEhcS9AiKXSHD+YgOZ9
LZgDwW9yECKD9pxLmFwl0wjZjFJSaHBO01ThJGP7jpPdyG4MbA06Z4tO25Xl+0Xp
VxD4Jnex3pyY1Pj9LrrgVaL22Y0fbdSagYkNGCp5qXzwvLEiLc0VbNTMc2fkOSas
730VlSfqcnHO2hRiV6pmVGQizgUwxRmRPEYcrhg28TVc9irVSFkz8GIKZ95xkDxy
hp6tnOhGnFOIxXoQSCX3Po6tjjSZJsk9eHLUvVKncXS4rNpDu+UwgRFw/WLxoUAH
Oli7cE+dkxY4yMVkX2Iu0ojOwYfXb8peBL4m+Sd7zDcWHxzyd0lCeXAVCbEhZiFv
75/QecCJqkY0DjWv+iG4GnB9rLPtqmFCDsJlMiPlN7ekC1MjgqIYrktnd81mNe0H
1NTfEvko1uHkyl7jAaWR7g7VWex5oh5xkhEnc2Cg4xdVGiSssEXVXSxMLnCWvjYq
Kvs3Rqfi8yhWYoQoTT6LaXc5FuSMwR8YOJ/VE/SNCIJkkjLTizqcKQGmu7v0JBno
9eziCAl0PGB/qZWYvQWCGmgBLR71Iah7COPDwB2YEHMkZtwTs7u543ztMTOul8YE
4P6i/ZaJ1HeM9UIjxhMYo02gcJpCFLW+NC8EyFsxFMQpEmKJq/BEYEq1sO8vZOQm
+eaC47SIAgdIXd6sQKLJHXqTYIF/G0cFfEa8Xh36DSE2V1DpnlXuw6CZGqmxaG9n
4IMdJ1liGFQypbkaGTXVnXFNt9mI8k/IlJWdpQ6QFZ5E66IfXkgHJE2uVQrghINj
1n+QI8BPL3lDf6UMrOqYEE/xaXCyp3UhFWvggKXV1l0ATacps4Cnki0B7w/il772
ySMNsna8/oFLKKCypqcphoLwZ4W9K1iNRnXA8zQql+XnG8J3TSlaJ9tpaKIW+bR6
AOqHPne1oaj4jApDHCGaErVXiQSPZ28efq2UVa8QcM2hVp7FDP+y52O1wNxnUg9K
yCPE3jUS29qg1iPVoFwjoa1808TUJbNcHLA6cL05BR9IgmF/BqSFpwt0+jQ/Q29q
yRkWDulV2+9rd169dHadjGd4xYGsSTFWkZsFm7xQaCmNs7hRU03ikf/KC4rXjzY1
ue7L8Fmb6spebUEDHf3yvc48CLcC9oKndUltn/Su26jJeGuTr5bf/xP5ptspR8mJ
bRKCxugfmgJZ3u5eIZLsPKCIFF8wLdbugAsOqkAXXzzZ/qo1CpZqxOVUNZgOCGW/
K8r5ssscD0+Y9l2zI85m8qZMual8VWuUhzELMvoC2BrMY5Rv/tySkJuQtfkl7pNe
Nl3Y3mi3X1Hr6TfALR/9y9a1EKftZWTpiK2bi4goEEF+4BB/bbAtXcSzMcjcxBTR
FTGKJtJSJdbWyPjZZHYxsA==
`protect END_PROTECTED
