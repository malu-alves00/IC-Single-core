`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gh96yv9UWW+yBCLU+lGnvfi4frL/9j/+HrxEpcxcfBKWiPPXN9UP6GrXp44likDJ
VJd1UvkAOL43e78lC13nZllohFMEZcCou5svmA5NZfMCe9Py1210RUqWm0MTVItd
XObk91in0kkwaOP+RctjD7N7I7I5DJ5HV35ypdRFnwd1GLMCXfb2K/9G84v2W98r
djuqnJqee0fk6VnKN/Ck5MYdw2i8c3BKfrwlpn+5rIa/wb0B032NErf+Ktgjrybb
/skUcHQGTqi6P2wZOklez+866amDxnocqWcFgKxhJK8ncAXpp6QRiGaRKIn8kVRh
JfqOX69VR+HYjitr1KTTAcL1busiK7Qgs50KktxXec0F+eWY8tn7y8I8YYHow8f/
arQbGEkZp41vkoFUW3MC/SftwtsBfHnJoNPigjh35pAvDms1nI8xbeKy7v/llxud
PbwRArCmjywbzMGmvSYE9WVxjMBzWyok6fK3BALWJF/7st+v81FoBAsh1PT7MvMM
sQUwTx7yaDyH9HtYT4PejUAvoyAhErQfSHs1/nVLBczXmz15PfIegTxMAMzedNVi
J3HrRGRe4ajvSVVXYJx3z+7LwMKtHT9+ec3b6tOuhffTGz6ZC6e27bvrWbtX1Slf
7GjKTRQLUJPEwaC4w6v5TZpeVPzO0XRu3G9pv8kdQb6VAAHUFC+Le9KYTXZwXB3Y
ZMK8uRYm/Snqn/ZUcg4M+L6Bi/3OBAQVRXlpdE10LWHsJ8OKyCfgh9Kb7+Isgp8F
7/aq3p8if1xS1mphPo2K8IbwJEZoH6tEVYdxgJBHgl4R3Ep2Brcr3vjT2CGKPM78
JFKbcj0+z9rW0q2bGbKEPvtFMvlvrOvShIwUob5xRzL9eu4u1k+gHTeaiVAlPutO
dHGKTpO0Jf+Akjxwmm5Wr9sloQ2xN7tmA2AL7BkxDBQpcVNHu4n55SbSwZfQaKYO
pU9b4sNf40wjHSB6d0XO+ueJ9bcC2RzfUzJBHNV/QDYnX/FUx+ebzhq0TDsDN2xW
bN+HBV1EkK5z00vxlNJ2vAPArqxSsUyRmpdIdPgCHqQEyjE+iii3LWnVmFMnpe2D
woo21UAXMQ/6GWSAmBy1vy2H7GQqeJagNLSo9VfDvVU=
`protect END_PROTECTED
