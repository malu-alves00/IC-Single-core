`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eDmLOWzUuGdrOniwKrRzIXDSRZlY74rDvY5QESNMRAm+1tVeLg2QaX/hmpJNh73N
KBG9YVF9hhuvr/Vn3LHAuM/8nJtKrstHENxZlt6HraXvIjm1sQdaE+gHm9ypDrvn
SaKw7HnOqu/buw+517MHxWUjBO7V2WOjyaQ0lPChkKyIYYwO6BCvnVO7jtwm0Lmk
JNjfpM0gKKktUeh20RxAA5jDx3eOvhp4LafPUSQxXcJbzRCQ1Qsfhnq+L1Ii3Z+R
7I3RXuGOy1Js3Q0Cv5E2paSHXjkcmwwWAu4XJCN1YSc+BVCKbMkUAIkly2meNeu3
FyRdOO5NYBV6b3Ii9PslQW1JVu962/jEbc3FsWA1F0ZK0EQUvC4cS7UKLZpEWGJ+
Y+Y5uoUBv3fyFieUBVHAaCS2zaMt+IlarHbVNZaXHPawS6rJmudic64P2cqT3lTr
zKtFfgxi/Pd+WBNxRwWjGBP976HgOzJ9cXliiZh+biR5GWAMh82P0y9Cbupc1bXO
zbyjWGPvx5777bfNSfIJu7PhiTTQym+eXaaKbyB2NmmD4331xWW3h8YWq60qYFGb
sR8uQ8DhLmBnVqvyyduRvpQAu1MBePUanF/JElpj+OltsWAjKX0k28W0vxRuXqNN
Dgh7vumzZ6ru/NpMM3lhVFiyy54L9InGFWjExCkfXSA6nKF7QOluqyCRlmXGgnVi
lzVL1HfoD9Xn4x/AWa60D+5CsrZHFqH2GlUNulzNe3qRZYdJ8fA2XTXZvr0PeBsN
c2ozvMFkCbp5UbhAlQGYPVsAs+1qQuWAuuR5mx9PUER2bG3u4JEoPcWZ3l8v8Hu2
D9some7XVlfVkjLsDBGyC1Wd/BPYeHg325XIvkGwrz/3mmn26rjmLOGLcKDx7hmn
MBga6mY8oJkhKdK4LXbggzXFPvMOPd02lpS+xKfnUdZ9tXvqQMOJEg+rH4q1pVvu
Ksg/cSrneyNeU1VCXz1V3DTCR/X69Et2CNZJycYOLnf8O1kIngmsCj0iB7hJhqQ1
SZj8whQte6GP2m2hNtGChDnDyoFKPbVF8aWH3l50vRavI56AsadIUcnyWVkmQCnU
3rKmyqG/lSccmVsT5G592aAF5z2iucOP/8N9ehxsHnbUqlFPcj2uYrbIDK7bGCBL
uF4BnadBUVXey3fkXMBdczGstDgPH7dVnCkvjPz2tAeOf2Pj5U/OYIp5pZfosenq
o/mU/8dOKsOUujiznWdHKu2hw1Kz1v6n8nY8Aau58eWNRtUKauEIF21+8vgeh7I0
tVgm7Jy58ncSqoBNLxHnAit9ByKFeBJs+LoO+oyvKu6Cw9+eJGcggWb57Ef57A3P
FchOrpSa+z17DX/t6sm4bSDLY8sUXK1d4K0TFr9ZZqEBPItCCO1BMP8vnX8SoSxz
fCo0AmpZCS2Jb8yPIMygPwVZkwgQ671XqCTW0DHb1HEDOmRw2MSN2++HoxHe8RTi
776zk9KPZiXbhilETfYqp63/7klJAicxeM0fvdpGe9H3Lj1nWb9heHAJuYYIMEqW
zGv0WFcGb2HGRqYGVD5QwJEU5bI8tbJWNQfWe3JKCE7T1+v19DmAIvYEWmG2MpdA
y0mNmY7wd8G5KcWLSlcxuNac9VR3QGY/QykAo9P/PuYYudMgoLQufRoZk/jRxL7f
fhwFJNKDuVmax1BkJhhbi7sKcPG/7tLXB8GmItHcrrir3Svt9k3tdIATfqKYeBzj
PvYXph2xC2mkBEcotRJLFOd2yJWUK2CzZp2rq7Hy/G02W2V6gOC4IOA5+o2omqle
+8qAZeaaawtve1qEcrMlVr2kCx3D3c1tBiWIve1U2W/P6nDw2Y1kLkj94WOCEA3O
o6DV8duVGpZ2/+olf25y1vBFerxI26GsnjYewfTnVj6HQfdp5a7Qc26tGNOq8ns7
iQMmfnjd36+ZJVqmxf1UoMjFkuOuQLU30gP1BxNGgDQYiljuXqKz7dg4qFTjt2yE
VLqY1+kDApGQFgkbAzEm2w/FWxDEP3JybtjfqGEiImdmqp54KrroyzH1WeIwvRhn
PhnsqHqUIVLS+F4tZX1Akw1W3AmpQYRPRPO8/EzK3+2/7Vs7B14EnuPxXdInoWrf
QYa5sFVghvLcHCcPgdBvrPBbL1sCZKGUmuecL9YwLf8DhvDvnZqpebFJULU2xG9s
BKUPO4F2hxIduDTL33TegwLOSZpNosmd1QbfIRfzAeBwz8HM7GrWuvRjMh95nZW6
KvB7QQ+DNw2It5OqP3/PEDGh8RB6Q5C/jS4LBC3vvRs/Cq71Umm8OA+CKmIbv0mw
F4ffBa1rEYazmpQI7KNgbCgnTkfJP6WYAw0288ZERJ98jIqM0FtDKkUZjcsAWsnP
GWkzjpSohl5Om4QEQzvgd4vdcGBL6bdGiNBRpEUft+dhV5ZRs/QkPboSBfqDZlFZ
e/epY3PdICKGun31GGnWdHRzMKfGsxSiYk5JE3pK7R46LH79dYNgdYNW7xwx1ktW
3hS4mPNB5WGWwKhAa3oZfys7tuZiJgEPdMqgChp/fg4npqvoTKv1BswlS5L3C9nV
4DAz+y/QQX0PIUiKLXi/JRO+02/rYSqS9qcfsKl6xw9p18nelZ3YSQzwzavoTlM1
T2fCeo+4FaSGJbjmh4RmYnJ2VUbQryWd2rAipiMq24ScjgUM/ExIwvWcoX/1LbS6
ZcjypuM/72YQY2sNdQWGWvynf/vpTYChcBknsmkiHPwW4upxw0Ns6fC/2AdWaI0d
THwwce9YT/Z0GtLwkzj3IvTcxBCEnzJfrb+awdcdZ+PHEogHwzaInsjClzFOuNtk
iUpfrEyGx7CfKcURn2gr7pb8cOGBB+2Sca8mWP7oFpfUpgS/yXEo8ygTC5IutCZB
JX2mFBLQ32oy7dk9N+XozavY8pTT/qOYVNWZb32Og33EV9U74heni4mBKRRrOT18
f2qPtV16sNk1OZnwubyfTKaRrEWaFcr0IyRMCwGp8keC66DHkQEuPGXp1zZdv13Q
5vcXxhW4fZFRrULIMcNdqKXGN+oYsTqrfeiaMqE54Et0aHP6lP79PQSqEEJsz6iP
O6Ki/ZqA05REg9OjgEbDfh/cOE7RZHokXfZdHoXnNeAHQcYThWr+5Ti5D5lLtoz1
tFplx0QQVw6wgemnuBzhuRvkaFhBADTOuxr58BmKBUcoEYChopzSgfDTvjxfYOlH
BeEgsXvkuMtCA06pq1iJvijCQ1npvE7WPazqXqp855tTJh3CVxdpJjUw9XUIJdu+
Rt3QfVjQAW2khDwmOMfzMv//dEsxuFGAXppePBllkcgANMiw8l4ceiXFo+0EdQUK
Ts8aBXAxZofB3mRBFHNqFEvdi3jfVfwfs9Bnenh/Hif+KSZac0ytIcCiOlIqkqR1
nEb64u02CWBhKoMd3Fru7rkU3+CGiRY4Wg+Si4aMkZw8vh/pqW/Jqh5McPumV7Sj
TCszmF/b0VY8o7z/8xwnqu7oHC5UOhbyy50PG7rmQa7zk0s9Lnc5bYEN+utilA9D
iQby6NBqN07UlT72q+fLURWODP3XSwbOWVCfeQhih6bJGVfOIQvedIMcoe/cw4Fo
vBBbI6gaL3JLQ64a0k3kSzVTyhqSTm+i0xnfNGtQ/xXFOgFARwjmBLo7lTAV4ki/
VeTliTCV/Z/e3jPG544jrfmAuPvNO9wx10vf7487RBK0FYUlFGXIfMdl3ZqKjXIV
FtObjhhZXwaIVZOxEwe3FOhyXOzCG6+UoFZC3TOSZk2zQ5ZNMMafiLpCMkm8KSH/
kZ9iabsiJdoX2VGNccV8wMXA3W/EFgYt0fqv9XjXRGbMgVj3qj4dI2VUzOxBOFjK
Ji+UIuSxlJhBfXeEqIYmXcHq20YCzArwE3IMFPrQf7NbophIq9p9gH7RxVxImTLo
yTpWws1J8tYB0hMQpNp1MKIC9xxpNtUJjlZAfbdOujgchzopQO8wTJli49kCnlgd
XOVVm+GI9f6pJ5Dm+eSyLpQv0qMHKz69j/fOTt1DThK6C8p5GDMq2PfUlQazQorR
1Ng7WlMgZ66HWsB+1CfpTTQENMNbvAbl8FeD6bxEX04=
`protect END_PROTECTED
