`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
viQaSfT5+j5geNeo4zflJc5OqV0OPdhPRlIJ3W24LVkZPJX6QuIRqPMAIgNmp6Uc
4Y+6eKY5aFCOfhZf0J9Vb0XNBKAS07zyOOO7OL9lWcQIQ0O1/7BF7YPppQ3XAs0i
6RSB/O/WRg4Hq0jgs1WVp3hvE2uKVxz27eZKoK6zdtIITUXlVd3ui1qG3m1wDd5F
HR+Cr6EoTfftqCquDFZGW+OvuIfB+Gmq/OnOHq7F2obZjDpcxr0petqDoC+cRKxR
ZFpMOG9B8lq42OJR4ru7lDRfXJHq2EFoMv2gA2d9lJrSUiZQXr/j0NUzPICxy+3E
scbQPBJQYwBfbZdvGAXneBgy33die8cEJ+X2nYlVSzaMJrQDcLSeuXIHQZCGfWR1
Wo4RpOcBCfkNB9HJ1G46fwCH4NBmW8DyzBCn3kCYNEayCJDvNDso1pGb7XAiX9Hy
zMbLneRiT1RRLtkIZd3u+z/dqwuB25I0Pe+lQ0GmcKCAfTS/StOZ2Q4TPdt1FVUy
ZOYYMDZ+xymDAFHTnGcDwtSnb/hxaP/sIH6PEMUg2Gx5SyxsIJQ9ZDY3kbZItNM7
Suusn9/0IRjQcFqswpAWjmT9Vhze8pjkbVhOISGfA7yBfNKg8TEtqAUmxXXmLr+W
U0ddNAkjoN82MaFehPCNiAiM4AZIafNZeKKPLUlh2H2OLELW6LqS1cogr5qTwoq7
fmURCKGZk2hIxB29mPWwfiKYMAOqJd96B7+JQJpNj1g+HStHwpzzaVlA3TTTGZ0U
JoJAHmkNDs7spSo3Cz007FAxnkFd6ZmZ0k7hfJEQs4/pBMSG1UYYlKnajePzeIRI
lz61QV40ixcXx9ovBVpBCYPCTy6wLwNrbwmnRj3Wg7LUCDzg1lptvJ40ZeU1XQ4E
DGbLEbru7SSY1Vyx6E5A+OENlIuH1pN4xxwL8IB6rVG78OC/hodPSCDjswX72ntK
DDAKdep/agU9Oe4vpKQMtFIYlx+V7dhP6wlA3uCce5P+GYb5jTprhIaxPOhqFrLF
2pdFBqiVgPC6V3pCOvRMjSLZfulY1XkmWRrZt/9kCjj0yGNxH4DJCyjoJPEkLZN/
tfvuTFtcxdhpSr9ZRVb8LO+Uh3W4UHqRfP7OTBrGAqIdRut1ugJO2UNIZHRJEGzM
pFG52KlJI5XFxuN9+VFxmJPfALvrLyLRRPf8szk9AvI/tspMpV2AuO4Js5lbyyFJ
5tssGLln1Y931kn5kl5u1V9SZ9KHgKQhIhrLRsW9WtA2JBTLjxlhPpk1Xv24cIL4
C0kzDc3g19vxIeQjEAPajrX8ITXHsJ6pnRPLYUf0woFnULsGcH3efEFgWGRCl0UI
8CygTBVCmYWi4jaIDGEKuJVmfVLQ5WUo3I0938kXQ7EmWRaNlGi6ZXWH6f9uP+5p
iUoU0cIOIfCW0x9STpqB/UKEyRw+1PyXpvRMsVyfhuTNE4aJ5vhkEJDsYomOVHpv
`protect END_PROTECTED
