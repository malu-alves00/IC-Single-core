`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
q+CMYMy3gnz+rc5KKuSFe1vX/rAuL5LGtxPTLC1qT/IedOrXWhddVI09jbNzTQDJ
osPzSB0rGTDivBRyxEOWXSTOpFRKkRxNIXbvBemS5bGLMTa6AIAGNb42BRF+Q/ZY
oEZUV+esoM/BzEILDMvnv67ndvxvSAp02YZzRIYuc+6b36aFTCHBrM5Us7ZXbY9V
hJwD70xy5dQqD29GIwk8PwA3jTlfF28WMajYHzHRAJa9wzSicJozCWLv1kc43l9Z
XRJeLsqJvgJSpIlQe01FkTw4LkW5Zi7krgA6JBchLM0Tql18wozvAJzF4NEfQxal
em/rfxWuqv/pVw/d4J+IF8+Y3mm1uD+R2aUO8lN4J5mn9RoaJv0GQKfIIfbvMcGh
wlaW2GpD4OlFw9vW/lVoD0LlKKqCnBUKkOlHf3rawS+dDEgJ+e6Xy5fUP0QcTAAr
WLRWZS/Uz/HnbE3l/BjP1rgCuRSuYn2k6MAq7ZapNqSTZ8ulVE4ffgZWveDUAj7m
ThEsPTUkgDfgi2aRgkreZ0lj1JPMKc36ONLy4zwdBMsrkeSi+Hm8ZDeOUrkTg8cL
WrWx7/p30s5+5Ol+3CcbxqbUI5IJQCOmFukcCof7cqtnlKDIWzRRBOnkRdfkkEwg
8s3xZERIKPs+Srdn8qBKX4ujuIf5cjQxyQ0H/qjMnQZLdgvzCPdm3AGi4zeD424A
TKv3ij5TqqlvDMA2zhsNQHucjg92/I7QQ21yBinO6+Cx9S8AzejIk/PablTHZZ9x
PH/MGtlQ/0WBXaZHxHzzyexsLKEpaR9eGkAnLGjkuX20kJFIKpCd+I4tqd1KtfyF
TkSED8K+KR7Fazvn34F/a07bEw5s9KQfbS4xlEAqcE+jBrc2kn88QoSFBBNGHW6I
I3yItCknv9sCORX28EO8ugHJszIfFPmv/fu3iSUWU97tRFEqWpIlHeaC4/hPnXMf
7p52+PF4MgjjUC5+whXAW+Oyd1vW3Nw2RPpHVt5BLaHVYfA61N+naFhrN3jSTaDI
BYdyJ7+F7TTvcjUu9GZ+kA==
`protect END_PROTECTED
