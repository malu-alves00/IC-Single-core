`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IsZUESXf4NMtED6wWVf5DUAuxjWEjAlK+8aRr7d+0hfXSXTlIieqY9dL77If6wPy
HdMMj5JL82B1jVshojPQdYSSabNT7bxcD/VmhOn/MPabWrvai/fGQg7gwSQDDKaC
/edARSM0lXonX3nfEyMcCw2wx5Rgsoh2XkoOdxlPUgwB4R4loVbv2lkr0RHbeiSu
GLFTC4cWQQjZGGCH/SCX5tHKK1LyBaHmBblXmzDiUVUNHEup1+/fZKBj1xzhd2NV
vr/Rd1bCY68XpF6QrlX/FeLlJbi9FYUNyH3S2zaUZmq2T3PcbBko3us3sknNW9ra
0uMdf6x4lpKfs6rzDc5F41gXeUs2nQGNeoVUuPCKmMpwV2xAnZDAp2ZumOMHhO2+
PTRGtz6EXMmLN1aX/0P06Ov9LoDnXwADoqg+AoFWnz13ZIeH6yu58Skd2t2EEhNy
9qv5oEv1U5XZMvNPaa08H0y+BwJtVQvdnNthkrKLL/kzNukZtPoglC+Z2hDFTSHg
3CNSG7gv/MosVd5t7xnue+4qz87lQmkbMeeyOg1pUYf2GSpg2kTdDrD94cVzdJYb
6LhWdONnK7+5lJXXIaq+GbNrDfXOHHWEelzLvZSyJOMEJSWhOiaPTCv+ecQw1SJ0
txdQ7iySPsCS4ttQRZO1DUPu6AedvgJcH4AEBnLYuhLebrJc/7mQ5C5ZC8uNSHPf
pGofD6NYBHj7uLKs88IPWoOtjSDn5vuBVKcgzDKOCTy8l+JzcBdDCzawFRvd/2Lb
kNSBJUaTGAg8b/ZDYkVwACRLpk1amiQrb5TM3tDWAhaYX8B+4V2na6NSjc/Fuj9I
4ASskPcjMe95FC8nh7DLL9xGBSq0PmB02M2Ow0JP8lA48QKGHRR9MqgKHGl+Pw4q
jDBnS0w9C719GSnA5zrpJV+MigDI6HFgh9MM0BzKaaQ=
`protect END_PROTECTED
