`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
A9rQK7ch4xNrynr2CgqtSFdwEsMoYCEF/B2VGNa23i6s4FVGF0B+aGyIzJtN2v48
HfS7V/9QsedwYSMAvdx/PTOXvW1XJnRl1TmYGcRcCWLXkE52PKXqS1mmCdlRX+V+
4CHd5/agRnAFNkSEvvFTzmR+NIINa43YklTumhCWmFBbX72N5K9gTj6Cp7CH9qdX
Zj+I0DtzMe0kJhsLWJwIe/7Q5iJ3YOD2Ew7w0v4yn5DCZOd11Yw9SXdI+V2yf6LL
TZ2YskqgeeQrBlsagVZXy+gvpxp+kw/3IErQhem6O14FeY/89TakpbEoMVatHs+T
RWwN8PpLJhDQhu+A12CkPhdZEB3Z+fqHFnOcLnUUR4Rt5XqjOpk1zl7BbyhYtKfu
Jyt7RUc5tTjVzlt779/l4HeypAcr7yppv/9epphcroNHQv1fXtdwQhreDyk6Ew0f
SIGIi5Hzvma9YRYDyadxOSgge2MOj76ghmRKZLYcXLWNPDZy/Cx8VQ0ERRQ2FqSI
CHOU+JXW+HZBHWfh2aOue8i1F95laKjCKi85ewF42l57HGRcLAJLlSVOA9zcPL5p
eOVsRtVA/8CzZs7a//SXEioRek1STQHsjxBiuZ1jvxW/eI/lQRFYsQJQSwhnfiRs
1x4g0zOGBqoQfh0hHLtD4COnIS7zCO3nhsMh/wjqFU12jRnTMZdZQYo3L23vL92q
DM4UhFQRgVhn95lM0dvygVJbVK4jqJNvGYJRkWHy0SMvfVfWgH9NfNNSZm0kteFc
wy0Am7AR7HgtgOsWzk0szVCHGrBymXIr1nsYDVunG02rc2qn/urelKFgwPnns/JY
nSjNHokpJq1MPUBNOcDmDBPzvOA9w1v7tUa52+uvx2m+AyU4AgNNyPN0MDA7i+50
0Lc6kEQThVDpGy1WzeW+ojYnoAoIho4YapJWr3JRNzHlJwDuEQzGESjXVafErKiB
LjLe/bOVTzwf+OwKCpX2Kk1vpZsif5VF4cnXimpFkgsqY7bcv8vyNsKB9Yz2hwHX
gu/X8Z+SX63YPlsy9MBd9F8W15qlo3ubrUmXJwupm5R0hnr5cwAp4YkYvMJDnLBn
0LCXIaEvTIcWIGPrnWZqX26c8ieLiRK6ztlUm0wpk6A+Bjzn6gu1Qxs4WmwGj5dk
YUyZA9kuCa6p8Ar1UkK/jkqaj+se9Yi7MsG8u9WTSEexD9zOAEnOP+GaXwA1ByD2
nS/lZ2GKyUGB9yds1RL9X53/OGGB3angO7AIkWJn78pWec3JhsXxlets00Xc3cPE
`protect END_PROTECTED
