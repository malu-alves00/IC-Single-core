`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MLvTHH0ts8Co3W79wC3fSZi61M0usCTUhri5tkrSdq2uIWzIVX4MThp7PT2vm+nn
h4JVv5K+5LQlNfEXJ1UnnyBrwZYfHyLa5KDhOb0LHZ11n4L/AJ+NYPfcGsOjLwYJ
CX17jzgQ9IzIYVOz5rj31hL2IoiRrFdglKiWcAH0BbF8jZhpd6DIt9Sx47RUVVP0
oSz2XVP/OkWVwxBONTTidCh8fMX3kL7Kctb3ZeZe7d31cUQPkY73Nc9xWfo1ybrR
9WLCiv58ZfqqYD0JZfWCiqcB9DbVHrEAl8oISr9DLWfAcWb8HYOo/xwfTRS6Zrrl
WieUCOX4QailgdbgrK4jsYcHH4DmeMz0jRuAVtzjxZgxTNtHUgVH6+I/wgx9yjqf
IZBEwRngij4TUKv+bf1ELUxY352Ti/88UFhAqOtBbwTbsIfduGFvmpHmIv/ADXzf
YXSF2gF/BTbFxCADHKxlBoBuVnnzneMya62La8MS10KwTM0j7f0NPXl5IaT4qKDk
Mc2J+Zx3KgUBmHQ/DcztiVK3E8MjA7bjaApLtGNuGfqJ+5Egmf+akbEE+P6BXj6a
4S4Hq+541NXT9mOsRI8nZPLEvKMgeFnkCUUjjG8PPFX/tbnvxOyUamDfv9w7yy76
ie3tJ3TvuNE9Pcs9MweEaiP0dDoK/GgxvlaAyEZxRTVufFYXlUzB/B+1LMU9gjjM
2iZ/LsY34QK+QinogOwsoRc1ltkRSknZ3hsnGP57EpDHC2BPTRT1eku5cDqPGCmI
Sb2Ccsgcet94G/7yYXiGZQENg3KML8HASkaSVzXReHN34iBDyPLdXtRSXLsPxnad
mDxB9bocBNR3tFEol3sj2M4/trdElfZopRv0lP7yeOMBny1Oayy8H0mr0axWH2dl
H9sqv0nQRIAzK17kI0dfK+kf5nMSpU+3sSSrP9Wpj7bstgyVrVhX00R/HodmXSBJ
gNnSOeD/hPeCQ+KtUbb7rZeDZ2bN9O+yLcTvmFh9P4+a9B1PP/8txvov48gt/AAI
XnOVdGcVqPidsvRX3tJFFP0vUyV9Bluj8UVS0iKKYw+oqzY0easFPuZkCwFq7/6p
nzIFMJUrKme3igPsfAOtavSU/wL7biCMdnLukCpSFixdCVBaRLNIQf3mM9e72VWL
vsySdrwm5IG5tdZaTk19cAAlel5zqqOB/2gso+W5AOU5C/UYOUr4P4nCWO/ZUC2K
IgI+L8og6EB6P6gMXDwAJ6aW0FR+SciGMa6hcsI33NEk6MIARLVpeYGIl7huK7WV
G58t9QnpG9gZDBtWXlWFnfsuEJj7ZCvDkVLRrPxDbxgL3FQrbdDMpBlmYs4iPU4I
8ciRlMukYiZ9QjItytCM4tO7bQA3pc1rsZE1q+yK8CURAPXeuwoo3MEB7W2w9LZs
eCrVjdku+H6e4A7udjoIIDrYLE+g6dujOetvpnX0l2afSKKoHa5DNhz+IVr4WQKP
icntgN3vJYs6LGPRVyZhApv51KXXQUJm0kI09O2iY50RuMC9xszcGsVAdlsL3jKP
DOPh/OLCcQIz/J1bl5OCqg/aI1ArsYhg56GRL8XwBdR8uHBRkMLgmZaWiY4CSREC
K5h3BLrTKCKqvT+cdx+7qPqxK6fNXW7dYMfXpfPPhFKYbiUvl/F6JdkJJPEpWNmm
`protect END_PROTECTED
