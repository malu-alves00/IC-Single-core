`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KDP01/53Ee6DuxDvv4y0ny9TUNZl/PO+Umivp3VxpbYG1cyJlM8NG0i+runUeyir
6TkU12DlgbyFKuRobVYMB9Ql7zP8nos2wv4IHCGrqg7z6gxSXPCV3o8pP+mTTAne
fCwQzkcL+K+jOHX4F3hUcqR1S1dgodG5enC+A2dqDrEsZ679bmCCt2/NNesAw3OQ
wiz2WSEBXmhRTUCDLPrWccoTRQFVegQgjYLHWWis1JZYiayxPd6dJiIQG8C2MbhK
NQL6g0l5CUfz7YAM/GWRUVc4Dcih44wy2f9Bvn4/Evx/z7DI5AUG4ECYXtTqHxEf
ZcIxMU5jrbp/x1k4u3AzCiBJMTdEYa0Si2eScpcx2xeyuTA4V0Ba2qH025WYfErj
cydcyWLWEy3UGkH6HA8gWSPQ4daz12u9BIuHSxxjNoz370wH4RsKyDnoQJiVyuvn
4+m/b+Han1uopPSLZfBA8LOzXeHeij2eQonMSjAAYs9erdOyQz9PhOBIsxKhjbXz
BGbrSQC9I1drr4eFyLkka1NNFbDZfb4j7/NE9GmXNHQUTE9vsJdqwtmGgh6KCJ7n
lnpfWxNpECj4PGMFWHCwx25lWDAtIQSZoti9Dt91KSAUOBlvfVvkW4ndR4uM7CBp
miNfsayhxek8nuKNzDmq05wgrztZPdMMWdWMLNoYvApIpyygAM5/IMZpe/1wvS0G
kuDDeju4anpBJTerdj47IObCTXW+jwbxvnZDNeqLWmoVAXk9+QL+B8vAvnu3EyEU
5wvG9nW+Fj9P6R0+gT025Wy0u2Mq0y43uOvKn9qSvYQsrEFao3JOIdXeNMtye8ar
edHSEU8DadfEra0xZqF0zeGbZMDuB84AgzFIdas71HGaH97kxfynmzQueUIcGAix
3PPtROmtj2/LBWvIyBjVPMdf4lwX6l8BtCJbJYp08N0FCwr+Fczf5IEqkztrYn05
hlv1Z6pjyGBA2bIARm7WjHGueCxE4jxgLELFLhkAzjOUz92xEgB1QVzBJyOarj54
gJJUihK3Q2n7duT4L29Vn/avZWk7sU5JKgck9TbRuFrXzmociuS8HYp29Ze2xNiM
/5yWhjN93jjew1QWwyjc6tWBDnLvCH7asNUDL7svWPAvM6wqK4ISV/F6lcIUalRp
9jnoEHU1FCIqP7gQ9oVnU8DYK8m6BMMSYXPTAP6JtCghAD1MowRcx33TkHDkgwXn
gg5rt9rZUPPga8yiXXgjgERMNNhpGKR2raNvO/y7r+zGM0VDqRumjfPSTGX4UF3x
WCIu6GwNGb944pO/zpFhTEXvJRycJ5Bg8+PB1jdsLm+tKQrnA1eJT9fSINReDRBp
NkqZCn30eGcGgI9qo3t+ljsI/HkJ2dW40yqI/NeyTAN3jPx2gTK2MXGNARgMWuik
E/ANutCTf6l+mGAbVA/z4FkTxIuffc7cEo9/npbmpspET6nxYTacdIrNLkN31K5n
ngPeyr+/4Mcj0FInbdzDyyf2QgKatQ1xOPLBYq8ZJqDx6eb2p5xiN0iJN6TSiehe
+TfsDk5aQfNBQUlJiRhxkuu+hoRmvBlkBhCISp+pGdez6HoQC9p9LeGVV/jRusky
sKEKEtn5ccH4WVZZoXClPMkqUyW3/LNztPVXtjAX50dEh0TogcuyedW4581ZkT0f
0p8f3C6GFpAR+D74JEVQqtGN87iJLClpMfMBmnHjo/U52FFITpz8WHSlzAID3QFs
huvx+W366DyGF5KYBjfO3mkgKdoSU6DBBsXcJOtNO61+jzJ/99Kpz1jq6D1TgzoV
Eny0ROhViix+qKvJP2jypyhpg/dOpVsYSJP9HRBBFOdcZGJdqyyKLJPVQp3ijGtm
1Jf3QEVz7CufzljxdF76QyWS+0CCa6zzgTfkCwGxJPiBU/q6q6Qic2/3XKL4BPhm
tv5MQiyoUJZ57ghSZDNy6l5CgdItTHIwF8UMziPS5TABjvPZ58kJy+7d58m3fK9P
i+rKgh34hoYdhAN8XvAbdu1E6OMrQS9w+GiG0IFnyPwvG8SMBItpraYSirCvMnJ+
xbTYGA6NCIPB/uahAidEpxcW2wlEnCFjOTJdMDWgPpnlCC26fi5Q6f2pMw7X/TUI
oYDxPb8J3vvYytpUQukQRKrzQDsZw6ZEffkhWi1m7xY307I4h/q7Ax5nD6UudYqo
95zM0KwJPXWKwCWxbcYwkxRNg89UBcS/0pLgMEc8XHp30LWUipXXQbw1MZdcpfes
Xg7qkylGwIEk8bWLtbPQEYFNjbiOE/yMrZloqjpEIYCSQ7x/Y4xhqo841ZcO1olQ
11dm/gNBCbeMVdjTOiU8S+Bm3cXRpCLygtdEiwt/0OWcj6Z+hVWL/eIH0TTvE3/8
AAZhDR//w/7+xoxnzVCwMkT1JU3CpVE2PUXhmDfkg//Alu5b1wqLgCofRXPS5pL7
a/wh8F3K8xQOyV/7/Qu4057okT/0o0OVUulK1jfgioTD+L+Ne19Nfh+8EjzHZWoo
aZg+SXmcba+g6tJuZtk+okEFBBtqYKodtDd+dfbwSqbuYc1oEXFM7N06KreJvsAW
bOo6RdFOgGqQlgR/kOLWxCy+Za4Sfb27xr+7cWHpbnFSoYttY5ztZ3aU4r1SMwW1
ARjjY5qPq5xLZfaZkG5EZ+TFtyNup1YqARV5/tXLCyyJp0zQ64vbPlGhnySAIdak
4fQqPukTZEEi7CVL8SahPfMlw4q/3gKo8fXCzOUw9D1YN0uhjMVmFF7vXmOVkaR2
wC0SycoVRfOEzCKvmZMqLwVJ/KYvF8qS9TsiOK/j1XCsZzBoHLB65YQ1OD/NRKSQ
+yQH6YysCxUHN07VgSI2V07VWsLS9NHe6XrDdyUrEdRp+cdmRAk1fyzfL6PCiVvQ
D+1wA5QY1NxoWmOAAyNH6414l3xPtgRVBY5rsdnBvUHpTLt2vDKqp7zT6rc/J/Ma
KUPuyr2X2kfrkmMBoXNPVjZ2TxRGdDks+xBvLPLR/m9345d/qDVsfRTtsWvGDaUt
n0bkDNTWkiv/H+ksW7C79Z+wNNjYSYNUVYYT4on+gSuTloxCTMDH7mljrvHmy3nL
MhR75x7sl3CZ8GosQthoTRE9U3YmrBeby93d41YFE98LvWOsLYSsP6qPXCZLjUf8
46EMYINt+qjpvqSJApYiqBTl6XIxBdEqcWVTAaY+SjNhIg6cnQcVvG8Cf2TRhg9p
i9mnopttOAJVJ4fEMISXbRDL8M1DpZox1rCpF13+SjoWPS/KVQQmoLJl1yiJZm9q
jbmBbkoYGgdAIVZppbNCKzaoNFHeMoii2dfK+8EIF9jc6iPOlGEGQB2Hb/sEHfnt
UfEV09AifOwamNO4IknCHgBHAi0EOjZHWTHi+YpSmA4OBNMCZVxbaaGRvJAfslv5
V/P+RKB53HuNhpNtmzLc3U27rOI42+twDkeEwZO0GGJqpg29uw2ZWxRkl4DPhCLC
UxtZDVSB3iu7gofo4MZfnC/SafX4POoqwFLj2zm3sjjpYr/U5XGsumM5abAiyWNV
GLJ/ayOPSG3oJuSlvtjAM4nwynakXRq66veb83gVrtZBswDc6duibL+po6lMQTJk
ZRK8qZmdmN2dqLvNc6iStYNq7MlpaDB7QqRUJHsac0xl2GqFREejqP+nNyHihWBg
PfTR1FHr6nDJyFVygQOPzDt+G5HQOcxqI/AtvBnWmc6hTm8PrBnmMtI87ohKHQgf
FVXhUcif3YTMIkvlM8vf5JfttdnNo1T9lT5aJ7obtT7YS4Uraw96XBaEDcG8tepv
rtD8xtb4gHKppGiKRvkAowBIBarZHXpuIqgtSpKN1x1cVFJAvCKqij4zreIeiTvz
lloiAFlgXU0q0YbrkZ7bxIaHgNpyxxA8xjfenKvCeZ1kUiqj3zi4crmP8RgYz+fn
7vW5zsXnlDeCRvNgPfq8uGeXk+e/XDdkT5V0Kek/rnh2am7VTv0cy+DFjQdduxPx
9pu/gaKz6FgTRke3U2TkPzEMtDBoQUO9oyVf0UyCgUhEnIDVWr2icczqFPgQkH+N
Ufh1Y4NrykpM2il6R5PNjrNOhyfBNAfk0wYgcwea4734v2r/rYQ68srrwGiT11bs
okO1Rrf7eqjK7SDgsocYK2R/kCi2uXf6R6t2J6EyvhV56+mgar5xPCKlHo+e0cL8
vNA2DAbDF5RBqyIgVNG5CRE40VVMaZh33R7aFPzcJYVgnk294LERxSTmTiJw0EDy
vh492jgrVLOIzsG7fODk0fnx4CeijdPMQ/8Xcy3LFbvxE8ktgvQG+HkONcC9VUNl
zz9sHr4nGIaL46jakhlyS+D2Fk5tAuNDB2Btz647BDE9UA7N5i1M1vDuIHEXAdsG
gkC0yewUedI0AZQC1L6UVJ8v9/O/T/fafpBMtur8pIs6epoQleIFiLCA+E7r92Dq
jOqA8MT4MJ+9gmmo9FFNh8ZkZovnaVCs3S44ZgLuPb/y6WNeL3qRLeOah1m/L2Pe
L6MIKe3k4b0pCsZ3JfZFM2c/Qwhsq3jJw3CgWHfc67Xkgzq5QJK6UzOqTJjFWzlU
M5k0puuoGPZjcqj8xlvYge0Rs1dtKyD6eoK0D9emfH/NC6VD15aE9RS9J4XpkQne
JvWHaITbYjEvQazcCtdd0dshZiv76yXxj2R4WhfWkVtduYmpvtCPkOc1eond/otQ
w8aJS0s03w4C6fbReGA6iQSTDKQ2ScmsV57z15vdKBTIwAy9o3uBl9jGAyQIMPeC
qw1pgBI0yKhVT8vBNEszWoy76mgyAM0xSaogrRThcwOgMoFEVLLkmux7Em8TEIBk
hnL6ISKOzyGusFddNYVBWCnkoUkTaroiBfhH+WBb35TrstqAaXF6TQ6/EdMg8H30
9lMl++bphaRXBAEnbkj/44Ni89gZQpyvA0kLjajf7HaNG5qf+e1GDhavwfNcTLKi
O9tLMI3f3LJWyoggdMiUJ/k2ltFDGnSugEwVyQEpyjVMMefTFQtw+c6l3qY34wGN
FnjBM7yYJBgxoT0dn/X9TwX9JEFlNUg9NJYddExfO9BwjnRzygidJhEvMp9eN17p
RIo/84pyDvlh8dV4/BzIMddO4YHJU2YKG7X5dfmUXJ4S8OyXZXwP9GWH3junsypH
9YrdL7C77xMUzAutKHrjyjXlX74mEyNDrnPYH7bkmInNeaFznO+6uZXYTKUArPFn
EsjL4p/knYgsyrdjG/aTJkrAFKuS3WQR5M00rNBcqyY8jVHfwjl6sCbXjOteP7CX
nFDGe0sffo0BAVApsAHO1TgBX7Giew4Q0KqrikQnYDUEkS1gF/aqeruJo+zdCNik
wFZWOk7aY5mwB3oN68QOWGS2W92kSmZeODmOxc6NJbreRUQITQkrWOyhez/0R+Hq
mfjBtmd9/VfTJGBKLT1pBTVY7hbrtbeBp3g0leP8Mjp1xCvgzv1IcOMa0lto0H8P
9rv13HXMZ9H1/OSOt0aOVnjowymiXFYnEovnoQi7Z5/rGEDylYkRFpSuZ2GDSbsJ
YNYxVixEqM9dJFl1+WZu9SnlYph4p9MBTeh6Sx8k3C8RLkzHUw1jTVOGRj5+uEZx
cDpGtXMsb2X+lM9Suwm4RFhBHU1W0vKRvFED+R72hZslT33Sse08kMGIlGfWdATY
5Rlz0MgP7XrceYs/6/3aWhO1p5aFGev+l8FwVPYIBGZNfpZqqoXL7rco3psKqfDa
iizG6MUSm1EnU5lXcq31CbXLgY1D07FbSC2gNCOHiAvr9diNI8Ofles0w0kYxjkT
/YLWq1XWhQD3zqaEUD6IuPL8x6KCh67CvX8drMOTenu36ZQBircukabOjp2iwdvD
Lt5oz/kahl+g1bQmzItiKod0dFv/kHt9glkN45nkNrDvmO7WAeid7CESV5/0YW+i
/AcbikFxqbiiuiNqgEEzmTWgGgXXzllV4w2d89d3Z1k+hRlFOKT3CDgMqHkWL5Cj
9ODtGCQGo1b2QswwmGx7GjSJ1M5bl2k6QaEummJ9m1daTC/Iu7yyAyPwgIlPRL43
VqySpvKYumX4SEJ1kSQ6zZO7lVhdak7DAgaZbvQz6RZTb9rUZUupS7z4hlDJAvWp
dtw9nmrTD0R2QPNWeyUXTknBDpB6k4415gJXpgOsS/wz01+U/5OAlYySGbYu5dnp
VPT+f2WUJaVA2mKgphVYY8P6MChMXyyrHmIwrHbFkMGzfab+yPidE+NUIX0R0sAw
MoJ7uVZnibcrM5X67SDO9ffsuyfmDbeWpYJf80XvZj5qbUIbtjiVm2v3mH5xpltP
k7nOfMLX5g7VZqTxc26Z5ghg49Z/w30e6bOp4KbPHcRudYNZI/1wSNWpyvNSF9m9
MxKirdaFi6A52Hfd/41phXIKbVBFxV4jW57AZ5vDKbbsBYasoME5E7KQwYo6X9tj
6aS7Zu7vkyqILFzIOZRhQhMCa/tvsa/XsZF+3g6K7vXTcfiekXD1Rx8Sm+CNgof+
vIPlIky0EVDyisga0aiG9RxyoLe4sVVX8KA5+7PsmSEwDJu3N+2+ig3rKKsY2Pdo
UGNnXlmZSe2/tpJlCVEVPC3vCYR/UYAPVzg+Ra0f2EaDDGzVwfqr54ggE7+j8F++
Uy+bjSe6SYKWf+/s1/UCFk5/bUpxmgkVK6nsI6R7o5OlUP4yMD/gKaLfJGKKsBiJ
3ZJQXs5K2MF9YzM6bq2/kU6JUN0cjcdNZnmaTkV21G9FkMbs7z+cSinLwfUI3i0V
PlyzBCQCHMcVPnzQB+XK2gSvE0jhYLKaWk/uTNStwmqfOqx0aPllOw1CZdk23BiE
dFh+ziwScdspsFhJf/Lb30BDFIvIGgRejjQo4q1f7iH45qVSshy4w7gVt15S8k+l
gKzXss5XEYuu817/HlEG8aO/DotZOtwvo6o8VN/Symh3xCqcJNlpck/Q7TgJlI1u
AaNu18xR5NXCj2vGbqU6SOqQHr6+69BWVws75o/dYpk0RF1bwpd5Ll9316fAauRj
4WVrfVa4Klx/E97zAvfAtSh5qfhj6MmtI9Oe030y78iVP4Wz/4fwKMsyL1AsH/Z/
PLI6kFJFWoo1khxqtqt8X4RNPhu24+B+oGe6NgFQQ0IT/DVQHA5WnXt+beRZa43/
c6EPa08al3mibMSYf3eKyqszpIiGoS8OJt8lWMWhnAJbNdV+jSj2uqtacaWRq6nx
cDIw8DjeLEJUdifuJedyPGRz4AZYrEPsuHsuoWVog6Lv35fmpXh98SvLnoZ4OpIx
ORe1MDEJb0piq3IHioNow/hdvXuwzjrFi4OMvFs9gYaxgiSX9PEpZRIwQRLASHg8
tobW01YTh0SX1fDM+UWOEVnX6AVVUa3XBIpOxvAHQZc7HJz/CzSPr+iY7yJmdrm7
nik8Hs0a8qCEtkfA80efoRV89KlSriXNe+w88XJeaFNEieS5/jSbNzClxmZo1iNZ
GZhXoAyLi2WYa/il5jyhLlDqd2WaSW9GFDcshxNv69bwW80ThLQJoeDmHc1HJHvy
+fW4hI+hs7imXETMuqXtql4qSLIt432Zyp2pw6cY7MyS9NppiIq1qxZNFfDETg8/
8KJdM3snJJhPtalP+wQoSEeGu56oX9zMrH074SGi+p1BqhZjRM8rvQA4HioogqPu
+agsbc7o561gdTD1mYhLs44GQDWU6/lhSWDVyvxtGzjzSgXBCW0Ifh+8OsYM6z5S
XK44AKqcG/ICHAGCaqHun9GAlrKDmaT2iJcHD7UesjgrFbdWcnn2jYZCXW4vK6s1
J2Jrt6kpjFT0a+h75R01vkM39XTq+5A4kfY9Fk/wQ+tlcOYop79q07z/ypyaFd6F
mP8tFPeMVDXPK1m4KkLal6GmRBJGtCA49+rxevEbfYVs/PPzn33+E0ldAG1oTUBl
a0jsvmrhvZ48ie1MS90keV2YLYEMpaCQwO1WznTboX5b53lK0CAboWmWpelU+9hA
sQpEpy2wkAiKqq+cLo6f+bRRH929KmUfKtwoi/bOvg7xabT6rh+hYI+Xn8MItHbX
jpxqideB9qplcGekoLAmy3FsV0EflldmeeKXG3NSzGvQL4J9/bpxHpuaWVBjNOwR
tmntMJ8FproXUXDcxZc6PnygahIeQtNFusK5kHAx/8cXQVarYGBp6dXY8od4GA6t
yq2VmwhRwA9LTs2b0tmJx9gXqyYF3zvqKSJ6U82rnGuqn8Ni/4C/0/3KOLi8eHfs
ckaTImG0KrDP7EyRB1ERr8W7YjEmbR7NqHPmCoyXlWI2lgUogdD38pizbU2mi+ag
g9SOtoDUy2nUTwrNYtZU4YUtfAJ3RUazhsUNjcdvnVZJmOEJUHs4p4d+vArZEeQf
vxZF8CORsMs979AJMO6HiBzl4Lz97ZeLrRKzjEr2aoSO9LP+r0OOsvBrEBh+IsvA
ha+mZUVQiuyclGNr65kRHMMgUJjmQ5Xb21LlDrAVw0FrTwXVz9tm7DJaUHJ58b/A
gfRr2zYaaVg6c+PBqEYHbsmasjr2vKxkKaV0xxFtGHgL+vY0VAK3zfOng4AUcfW+
2OWICc/Orn+2O2kjDlbSE8shqbRNwhozsLBNPbScCjLFTqawlHw5HZ0asJrbax/o
hHaxETYSGZZylgQotKcXvVrDf0SWQZ7XCWAYzDfX3gij0BmC+uYvRs6gMH+IIjCH
A2X233lAx+8aPq9qJnNMnP6c6XfKbXkN9IJC8NtnUNwoDX7J32VAHWI5Jkx9vz2x
MlP6VOcmTbQgD5jMouugAG3YKDhLUhEo5FJIK93hzUPJD6NBZHURFaOVSsJybhe6
JBJApAtay14Wp7jrm1pLRr96n54oRiYGjVmGWptQWMsYmTzZDtt/SHaI2sQLJYyy
fPOZuwwpKX7rbOzGk1LXPj3NyXGMiRXUi6ZHBzkFBFHv7UX28bbcmS/tAePJMreB
yYyiZqkJxzs54Hss5CInb1nOkMUiMEOgBOmZFyC5rGgSg8CLZ0JxTMotfKlLDpDi
mEodyvyJCsEgBQAxACZQZvustUsOOFWwDDyBEPoyuLcq9ZC/EWwVI6rwZeHS/x3V
Wgec0PZOlxKyUgkqxeBKjSanzBmCGpW8c4TZp4OOmDGyAEtRPAQd+cfgqaCfnCa/
RH8oUG62+FdI3abG1TZeAsxDPQ8J/2jM6ANyquiIQ65zmd4gNsaQ7W4Bg0deKj6A
wvhb8oV/H6d4sw4McC30WlHPApczr73kvsVx+l46c8kliUQR3ipjzxL9ou3DO/ln
Nz1ojy/ksx4cml5NBkb0fFFynVfVqbCZgIU4eLHxrs9TkZMj1uxYwxGjw3/k4gm2
OuCir+7M32+9CcA/xVC37ZT7O3kOMzAEjh4AIB/P3zmcJcJOzE3x22XEeq40JO4x
qLo3dmsqzpVuNtcBF6PSPznKixPFNHzj+pY7fLMldN8StmCPNzPPBE7c20EABUQL
aOkCnUmAVWdfJpTrGf5wa6WRsu5lzFqxOKFE21UB5fnN0ODAQWWtK3tD3MBWqNrs
oPYs9g85HU06WAP/LRzRrcA2uHsY/OQOn4c0Q3+HdXlTciKQ1pZEI2/ndmVF3sdX
FdZlhK8IfuUDBD9Z6VwzTDH641dU2jaRbrFtKc3HFHwy9W6aJ7TUdsBZf+J7hALx
x1YEP/NBbiMzOZMAn3aRMYlaU5Ba02Kohyh1DTnYHbj/ZVnpbay0n8PuJv6Im2Ft
V8VbMvBqwTM0AZ7TISk54eOXBzDw6fcgsf2giqUSmFWChxd2LcX4SbCYD5wbWyih
ixBDDze4wFV2CGYQ2m2+fO+ltsbjeT6Bwn/ZsfW2s2uKF3WkGtMrgoRRWgnk0LMC
vK8RNZvybwhekyCeTGMiBG3GQ+FdmPGKLlbe5IYYiKOo0nJfHdWd0rMDjNbOSL6g
cux1HYfU/+vSQeKvOntFux4AQEdVc7jmwM5izkbIUeg8ZyWUjhfD2Q1o+1auBq5q
cv+Wd7vsXewpIt4jeMg8N5Psu+Wd0MBJbgxtUxfDi4OdUmamGQXU/VGNZT3LSzAb
Y3adZD70cMJTmLKTyuWheP+fJT5nvct8muNIdBlSPhc/BvqvV1/CHYlBnOZTYLB5
/NS2tZWJggbeAATWUAOPHL6tt1+dd2+fk8eKMkGnRXCsCtOo6mjRlF//C+Z0GZkK
oe3iB4xIqXalmBXv9xdylCny9kDRgqlvZzGCk9WH+qIypwNZJTHAeLb3+ReowKvZ
4U8t+kdYh1RedlayS90Txa+gNvRzvZttMGtRQXvELOWjtISlcCeSqwqQ/JvYS4mP
zJwVXq/01aYrR40ywFmQ2KSMJRUbXfwjS5eppY/A0ICVkO7ez1dygBJxVv5fWR6f
wjInn3eV23dkzo+hgVCYzkFGKEuZCHsOXMDK89zaR3lj2zE4XR7U/ywTdbIidaIH
Kz7S7pEuQVFAOpuNWtDQy/PaLvOXYcmJoZ3RtAVtwlVGtohAQlphM4Lp/W/fMPt9
lH9NaylkH536YZIA9yPVqDRRrW4mVkBgoaRgi6myYY4PfFKzaeDWEtrYIGI5v9qs
SwP1cIzThPWBIetV7sce8kLxVqarRB7JFvuFzuIAD4N27R5ulwq/qDT5F7JxVWm0
AMoGRALsen/oXJx3RjYZJuMuL2vw06WGqmiFgrR30E9j2MlZ3IQNwqQEwh+V+NEt
zAlqX8oZs7SWdoshcGO8sHXEaK45M9e9QEUABQBPRQKnSxdL/DIvnZ6DjZSvpye8
ND9r8b6RX5gR7nNNEqVY2g==
`protect END_PROTECTED
