`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
btTm00TnfmRy4Lc/70RqeO2qN9CgVhHvwpa5gyXJgFNEVrqkDDB1k4NjAUsJRrb3
brNEM9qinPRaW4OHdGpZFx/9Xp4tPU65CWdeBheIkHSeSngLhJtUUDh8aCK8OZX4
o/ADS14aKjGNDu7KEAtDZcEsgcnsDm7wKFCgU3w/3+XOORZ0FidAvAZqNMFrkVls
2mBbB86njGS6NNQqQ6RRjSfgzwYxkmN0PUdG8+uMj/AdmIdk7HQPWtpRYr9QqBSw
Qj8ovsd7OsqmSvuIrcj3qBdkMyhYR+VpljaApf/FfcnGJhbtVkVrq0WU6iqv79PE
m62+oits2dpi0GwpufMTj8QjPgfqFGkdv6I94OS2yEWNs16nCPmlv4Gc4ViRV2sQ
PlTpJ1E/0TzvYaro8qKndwJ7ZZWmbiBElORmX8B0/b/HkWgZRZIa50phDCfKQKvb
4vSCI8vX+yhtO7tE/W2v7qLf8SQuCB/pDBTAYVKEgbJfiiWtSX2PiZmrJdC7xVRz
ViHRHH3T8yxYYZBrhM3/iFzVb0AAzJ6Q3XGFB8GhW8653Jc2DcItU0Le0YM4K0+N
nnek3bFZdLqpGF/3YXt3Ig==
`protect END_PROTECTED
