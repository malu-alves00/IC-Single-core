`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aK1dpZxgU+2wdOTwA37jeDL9C+5pR7w5e/ky9AzeKa3ajtmHzA5O9SZgbWnikFM7
NyQM1MdXSBsldznGmxj/LWijEf8KwYosXe+KlZxP1QzIYiNvRB1qzPaiwkb5fJgZ
Lg+ELwla319lIsCk/xVBryQmM+HHlY3lrHnTLOFzofZKieTc0vu/GztVp4E0ERla
pdrDFHU/1fVAs1yBEgjxZqngp2oP/w18fXSx7Ljey6SJRMtHJB19yu2D4dOHYEWq
vS06SabekPWVPQmQYZxeOV8ZF8ngk/VU0Y2iwDwPiK75+kC4Ux6hP2P3UQtBt5+q
Q0QCIJz2sPGA+yQ/HIyxpoLCrtih/SPzUBvBFe2TPcnfLCNXcSjAD0i6j6GBMz3n
hXgcNWhaJ2SJrFp1RNfz/6rj0wk4T7jE4E7iSEr8qjw3pptIH7Vxb1PTZe8UQAuU
qQEeYj0z2xXyhNrRtt+mxHET7M6U0fbEiQlsdtQnbkApFKMdrX9I4PdOJ0lz3c9J
IDgIhDNgmHfx4+QBMyEUYrBv6k+aDWR0Hj5rhni8VRUX83xUg6rUwnrEJEgI+fwH
tYQULG5aqdM8rFASkNACDWC1d9mRInHdoPDpe3veAb+kZRQEGAFNPQUypyA2QBwV
0Jk42/FLUZ0PNcg6MO69963fDnt0pJ2wa2j1wGrvOAXvWhqXSJDE+DXKDUxAH9Wk
Ws/4iCp1K0A7gcf8J/Ge2Ss2KnbyTYaiYuXNduLhf/U=
`protect END_PROTECTED
