`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RM6r6jDdvAojRYYcebyA3w6RvRJHK8vy0tM1zF8Tjcj82FfyL6I0nXrkmjdvyOSo
4LPA1evzyFbc+LqDONTyoM/8WgDXTduPIU1i3VSqwfHF4sZKev+PvTa+RR9NtPqN
QLKybH41EpqDNh8TkIUbqwJxbCNpQ067h3bBEVEWtPtM7GMAXTLvYYhmbaEF94hS
2jSPqSyunzN+q8Sbb0jtGt+GuspQPZHbuqrNrkKo+Jm6ZdwUhm9mLXXRLkqCYFfC
LxRQ9rje0i8RmaLGozr+sgGUn2NEouf/dAP8vdX4/0bZUwGIO7D/3cVNj8WHk4Yu
ibft4Axhjdr+vks3WZTybL06MCCLjgJ9ymLbb7R5GP2otgTsZoimGECr2m/UCsJv
oWoukL2BLp9PD+DueefxhIk5RsHngHBX7ILWUNAq3sVT/jNUl42OxdY59TcQNJiq
t0egra7e26jq4SIP2k8i3pbVL/78TaA8HZScE8QQd1H99ocR6DNuhhsVtvNeGCZy
8FdUZ3IcN1zm+wsQ7VAzPgn2097FNVv4C3CY9lx+6iXjRNnvMXVrD38qPNi/LWgY
1gqcoKu83rWPe29fDj9AduTtMXaxCFZ4KSOhvmp4id52HwtkBRuJxt8G72JWwVKT
Ee97PfjYLYloZN4NkDTdsBa2mO/sNBdp4IFYcuWPMxFVClr5RIvxE8qpjsamejy5
aKZF364xuEsLxiCfKH0vvE2R+aUQbivIpxu5FugyyJPaOgVEp78pPjZC0fvo0slF
mIEPibJ64JAA+Y6/b2rcwhqI5Cb6mUkbW1TYNYdx2GY2gW6QOzB3ZMs756IlI7mD
mZ1+ah99e0KFJlvhdnkSruACfi5hOraVZ2JYmGNOzL29DH682w+dSR94qU/SUTiL
bdixcOoj5tlsuW0OLRH9iD/yOqHQ3YoZd7YGIHE9IoHPyOP7v0AjKrp4rXiNh0Xq
6oMKbWe+cv9ahslE+XoWEFL746aLmqP1HK+4yh8ghyjztJeGMZB5+Bmcq5PCS3bA
6rmONQWzB0pI2SRGXxtkN7RG6Dj7+gvLgzQXGfu1tLj+Sorp8d6WTTnL1Iqksy6r
8x/s/uyjFFyIfNunzYkHIrdYgOlmAxH1FpK3yyCWBIw=
`protect END_PROTECTED
