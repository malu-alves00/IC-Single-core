`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xjQ4xf6t5j2TguRIbEhNtYmhsedN3TTdHqhjm6XRUSmV9fAx2wN8HUpSbKc2QYyv
ZpbhRx2oW9BlPRDI3d6bn1F+rc51wbmMFcqjTrITLYC6KCJ1GrMKIopLrExTVyIX
qSSCWsUnu71tbCEDFu14zzNMZgbyKeftYIgQ7w9u/F4xK5k6LsipMtnq0RL8i9mH
wvq+LkLSA6J0+gmGKpssQYE/VJY5WyzD/Y3B45U2QGpkMM8QWKRQuATL/F4tlRe7
7pzHKAgr+J1xD/GjTEhcbSGojj081t6m8uFPu1BAJ3yEQtQKSyR2WykNBuRRrMkd
prg6qMRtWgfksxS4YxfANtxAoWibIe1krzRMi0jMINEwqm2EZvh1L1FQMqdFAcba
nFXJiJZNPP2T2oib3VUuO6+dkj2bqTy3uIW6yjt7OQHnxOncBdMHWSF7uui8vgTk
Io8K8auWq/Y45eGmB+yMiA8dYQAHQtAXbSJMiW2O8tKVwYR7gPgUhO9P/Asg3r4N
zyop9QnY11WkilhEblOfz0RXupWgqNO8E1lmbmRuvSnCo+zxZSOcsQ7bxgvuK3K/
6Npu3yKa/Sw1cvU6XmhKs/PmOLBCA1RNv+aFQMN39mT+ch/hzVFD09xW7iXnEaR7
vVkO/M2NKuJK7Qhr7DEwKXEMvzTX+iNKLlCxea04pFRBwyPiUx3ope6NrlTmyDH+
fjsBFKB49cvnhfApF/OpFeqxzvYeSuW8huJgnIPyu540XuX6aoZVHjDOjKw8re+p
utv0aoqvHM7PE6T4f2AP5atGo9wretx7XF8YzFdernmDKZTSfOkqfEAAyCOLz1NI
aJxbu3/4qZUt3T7R0AYdojbDOzYXE9Kviqm1QTX+69jHv46bQTO+jTUbwKzBTvzo
LWdIz7Bay+tnL5yO9ThCLpEKzvBTffYx8Co3QOEKduqlEAhj9zv4jy15OiiM3061
rJk2iZHfgCOIz+ofS14SXOY0O5O8FdDUqSKCWZQx1RiYo1qIKhe0x0KQW4VAlOE9
Qg57QHQBS21WCm+fXpKFYYfwvAIcGn0jA7RySqr2jcKr9j6/J4NTi62CNy6Nipik
IIpxmsEqHwNWO4NIrT85yXt0oFuylgLeNDqU+eO5Gl1bThRZYDC4shBIP9sHVgia
WUWY8UgWS3WaCPH98pnVojoZyCw0bZ6fAhSZfeGDFVt5s+/bHfy3yCFpa48z/8Z4
OMWj8tKuSbyPVb1GD6ioSpuUCNKcOL6bUdEyOnL9BPiob3SLneh+6NO88940TwFv
/TBQW1Wqo1oS2do4pBecZ3VH+KYQEX1ajzyxPteUEF4=
`protect END_PROTECTED
