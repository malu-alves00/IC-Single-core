`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gDxeNhlfVTahAFTcCSlWfZSD8Z7yj0mb96yKVV2xBA1XHYl3cm2i6KVeRXEYCt/w
DHaaTjz4zdDL4efQrO711gBr1D0hTyTLmwl8iCdXqtBrt4musjU+HJNqzCfspy9f
6CIpu4/VtbD4MCT6wPaO5J5XFQEyO17d+RJhncDHcUNvu1PqP7jOYwn2KQ8jpVAi
fMlkT+cqb3mCP9abERwSnB0gORF2BMVcly9sB5dm+IPGPsUrkpU21sQCSwuP6OKW
6+Ma55ntqbzM4M2FuhryrODGr75bIaDkj36d8pNOX9C694tGCr+9LGPMkLePQndq
gecEBkybyG/1+HpM/JZnSBtBJG3OATxt4Ao+V1pLDTw1qQAOM8j/mDL4AkuZVTwa
zU7ZjKL/GGa9tnZcUl4xGbBMCTK5+HQTxZMge3vSRU6pCYJhHlCv+/DG9KwhpspG
`protect END_PROTECTED
