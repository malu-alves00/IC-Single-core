`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gvkw6kIM/vQZWCzAf9cpAAGMQYGBhYYUXWEnO6JCGlaGoyJTLCOnuhrW75zuA+oB
M9TN31o9HZd+QT7OoWIz+9SswUj+unN46kK+SshX9x31V28djhVlMgqSfZqXjSts
LE6ze+K1gNWOKheQXkBTddh+DhM4MnfbDDzwNGRvPj2Ih89oTHlujDXQv6Z1mdDj
GXuFZRGDMHIRI3tlfVAOYA51yY1zqobc7GSMfXyRsUja+So+qp0lprk89C6Worcs
2/ClFCeJyVyQYELEVkUTZuExEG96yjwWPZyc0rpw/vxe0DmR7rYq/Et/kGPw/yo8
HINF2wV6TLqhk5/ks7J7nd/glPtvAq/oODD3CSyrUzR4qIKrFlLihFlNLqvUk84s
550kzZeIt1p5nI3UXs2fyYzvXtFNK6bktYWELAoBrW+4bEJ6lShBRKdAn87pCUFp
9Tg+a0F8OdzIQEB4coPs8F/LQUL59OfdwA2rsuqasgJA71a7Jms3464cmrdfGxxK
wLX6tA1uysUKqWyXJdrhfCTSEBYZDaTnIY3Nb3G2HvCgLzrZjpmXNKP9TjA+MxPs
RQkCpDwy02/Q8IA8z5N9DNzzbph8cq6UNT9d6miggb58gmx++iOZl3YqU3H2iao0
FDkSZy8yIIE8xxHGoCDRr1EURSdqD/C2sFRRzPLZ3pa3r7nirwQrCUz/Btorjh1u
5eXUxotRegSWQK9ou2ZNjpaWn4kcsWOR5ya9ojfHvKIGBC5t8YWtqDTFohFlP/yX
peCpawCa3I+6HfK7o3+I5m+My1ASA/CnCpKoGgAqFmVA4RpW+5feLtwlCXFOHrAa
XoTa89niioPoJrHWgjACSd/IrdrjWPuyo9h+l9Cn0EP5KchMZkwAUEc+WqPa4cCM
jl7//aRTWwcWOxaYgUIlZjF4zBYzYt6Ot1aUfzjvzJk=
`protect END_PROTECTED
