`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MHyHl19+PQAtPXJPL8iSALWQ0O3VVkx/y2+M0vrj23kBbc98/5O6TXH6tcx6bpR7
MN7K6E4/lNQWLfRyyU1K/J6AS/54esIYtsSTVIH0d+TlI1uPb8yhhtR9j8FkFPOU
1HgriYfcgNp+H9qDRfv10CdSJqnW7ftyHmQMFXaQ7YOZGE9ztJPP6o2eKy3Ia0EE
VuVs8+HTbpjabC/yly81g+Om+O/GTyvgyfe1ayBtUBScMy6UdpPDOQfjNlfflMmd
q3g7bnGN+q0Xfh7j+Ju++UBdHmOc/6ELozXuoV5UhmDam/YBSUl+wvWXIDw8b7KY
2ei/DUjXr/tLroWp3O82xUpPJuUoS/79083lOFMPTLjPV2n+oCxGAju6br1rLhbi
+U1F0qfSQ/c1+/0BrDRL4nxWHytXuD9IP9TzzV4qW84xDsA65trW8ehP3X+K4Z0t
zwGzghSeZCuYIuCApcHz4hZJDQKbvqIch/D7Qf13jzFmGEuyZpkHhjeApZZeMUvp
ErRfqrnYAo/sqwuYYS3AgNGrZmevMZBjb4T9tmD/bkDsJaVEQLeozj2kTklxxXu7
/1XQ6sJSw7FJ4ynTvrnC9YMDx/WCliVP4eTZsJgoD2ZB9XyfR2Mus/eV3Av2ubVJ
GVWsM3hHccoaxNg46Ms0RdXsP/1GLyyDlYK9yjy5+U8odPD4QkYaG8eaU1uLZ2BZ
RecKe9dXZHS/ChNOUEd7hznDW+Huy0G8CBDeV5iaEllsxL0K3CbavxRFfEpNqkGV
hw0z5MH7dUrmPP42Ldo55W67y4aV0HWv/hb7Gcti0kNCSmLlNu7kV/n2H7xfdEhm
4YL4Mz0PEaAV4iP3ao/17QUWJ+3P97t+hctQ9Y3mfqW/WW0PUc2ylos2P3spn6Hq
0cvusnDpAOShTKbHRP+OVCEnkI6ptjtO5p14ls3UTnU7qS11qwiVW3CUlsCq3sj+
BXJsDRrlo5riSx0A+Vqa0P/Ifyrr5zE58W1sG2NEU3r0M7NbafO2uHoX/0MmfY1X
xhwyGsE7VZJFX9qXZRFg5+F6MWfbEHn98ocByqM6mSrIF47FXmvsaRuLaxRtp8Nl
ZsYOaKmqLqF42xWK8uMButydKVStl2YHG9k1vTckoWWPRXM5u0uDbK74+eZZJyKZ
iqA1CS+nkFfDCv0BC4H1JJ84+FAFBvLO1OJpXvaLZrmQhT+1o6RqletTUPO65HIO
2jKPeIQquLuDgDyC6R198pD6+yqm8/BTwOFucZHb3UF923grr6qwtmzpHyuXk1/K
3wG4PGO0mbbmKekBpt3P1WI9revQo+ix9vc+Fzdm/KGCZjk7Rk9Kubf/3yGKJP3o
8Xy5daGgGsK4G5iU64jEGjXPELnGiDGuHNsPZwXykp0srd19aFz7k/OnB+FWWJm9
5v1HJHjfy0EIBU2laobi0/UGtLx/KKvGga0PCuyr+HRlOlBuG6A9XaK0HSd6m3j8
soqZ1W8Xi6VO8spcnlNUBykligXBLOTxsz6wd3ELytvdNwG12LjNDqATnZcXWjLK
1+O/AORz1UAHonfVIPS05TbczCIzPA+q6WIAF28WAsQb8pyMF7tD10xwwEymsOQ9
UnDIScsOHQYuDpkG3L2mIYRAu5fZtVpQaWaKrbvr/IfRqIFYqErvnJDgow3vh+Ss
Z2ZAKW3bEAvwo/KEYgccPOtT022k+XFm4uJCjH1n9ACcEKkCkD6F2K8N2EAoutqw
XIiqvrxp89IU8BREUFiOfqH3KLA8p+8kETMPQBssSW+pCUf0mo2xaW/dhdvnkxD+
H41TZhj+0YgD+W8rVf4T27K5ZnmlczgEY5dnsmtEdf7y7RUykXBuqWoViHJkRX0W
BLWh72l9tPCb35mAFPv0Po/ICyoXSz6HrCIjzCNZvyaW/mazYWnQ2T96CIw0303D
d5fLEEjoq8Qdc/mGdbAFNFDfLMs4SVbX/BQmx3S6q7uAyuKHVBgRvSZ/fLs23Unl
GYsV0VJGWs2ojui+o9mJ48DiX3C2pz5cNkrhrlsECWTXTElkrL+zIlZmbK5kawOj
Hy5qMy09QLj6Cf0uOXoyrOU8gYT2lquXNMI4fNa2+n6wAT1Dpcusv56DSzba4tbp
V7rkrhRuYfBJWj6nChrxgSrX7x0Yn2ezWX9VIcqBzLRMRkS7qTpQt7pGXV9SKoUR
geNtakkOI5E6dNBrW311pkrt/sUdBHaj+APC+Kh4W3+XL56jBZxHRZsNE0c/YmMo
Cl+vq/7JXD4dBu//3kGT5cb8zTKHVTiEu0iUzBN4tZ1NMOSi6CosqjAnfC3NVXzq
jhjF37Qm/JY6snyvoNFNJIdh6DzoGdnFXLG3X1to84tv8OXaP2OXpGxjXerfrCnA
UEgH5bq29Mot5mrXM1mLqmXJTLTx9ZquUr4/UMtYZcinYOKtG+JRqpQJ3kSFkWVi
hAw0rYxYIK8vDvFQvvPizth/iXc/9D5Z8Qsf5A/y8PP/MYxYMQozXk2gAVlrPd9L
bmxJWZGpKmpYLoI7tBfEs5AeptY9Xust64CoeFLzFxDIUIo1S5Pv+PFz6d3KgMuH
D/NVpSNKlOEPgYCPRFObDT3iASt8ajyJwRyeMsjjBW0srIXLMFh35gpOLl1M7meb
dSy2gV+yWn+D/G4ylCyZ0DTRgdH424mM+7JZuQQPXEqnYDVRPxhZ0WNwwZpLzrdx
YOx6jLeMzURFkBBhKQDs3qZu4pf0YF+30iDXwo5ouNIpj6pSSaMS/cfR20fl5eQ+
h/DHLbtpcNyIvc1KI/OoJn5+8QJuWAU7WiAcqAB1n8yX+j1Id8sJl+70+dTyrCps
6Tb/oGwvPoGTQo0vp8VwKtcP8CdBrDCgHUxbOBu7/WKUWsam3yDUYYZY9sAA1z0I
H3BPcnFoOFnrtYcjQbSg3FsyB0p+Y2V5AJI5obHdPD1LTiNT1x3eSHe5g75M/Bek
dY5wDXGYhUjrO5ZqNvqfAA==
`protect END_PROTECTED
