`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3QAgU/lD57hG9FNCi2UQkk8I3F8N6c/C97ma3nUnRq4XFrVj0KkWh/fmeUfDewWx
9LMjpY6d4pzBvryofETKE4eeM89AMWFtYQBr8347JMMlPz5zjqvNKKiBPgE6rdw1
7OST9zVixSFk2eKakkTIV0ce5q49rVcTa/N2McHOakhwTSmpL4N8h3VMbQ5Fns7T
I6U4/A5eWAXbpQMUOKy+L7Wt8HP8LXIoAWWIi1QgYvoF++H29BXNxzu2ZAS6tTFy
YWLfxZr9hNBnMH/1qCq64rZTz1gujhDaoPPTfjgUyfDtsQ/hIaWMuK0ZRCaTtcck
P2tLLNXhmgYBBz7ygqKOmcjACHdAyd56tMKUwqxQWVDOoqMmgMCaQlzmA1QzaGu5
Psrn8hiRttqQKX5hdeMGxg2DFJLzcyAjUXRNAWNnrzjEdZKL0Rbwyd7/5xxjqXa8
R14Rc+ET/E2eFG8zAC3TZP/ctiW4NBoI/tCsT0InTwLu5SCUlFFHc/aEUq83w/3l
NcaRCGgOWV7S3432HqpgVE0qHZNxHXlpSbkDISldkorlMP6CMr2rWStPMG//ekFS
hIqXeE/J1O7zwhiCNhGqD9UsfZIiPuASJjU4Mva2H/NJWEIv/5xPOGAVIEm57MWs
5rMr/bOa6PB5wXfnuthWv8CnGCsfnMQCr/8Ck+1LRjw500MoDNWefkdRKYQF80/7
X12AA99r2YKrlrkHPQZ14hBJ24cXpJcPLDoAQ1RATZpUNBnZHy1p3FiqIEDqza4C
5bbSlloJl2+tIFMupV0pHXRWJDxvwI7nkiSyw0c/KeW1eDvwPd5CezQTExEwoS9j
6zTlwsRBqbAoQ885Djotb/K8k6YF0S+Jaix4Lqp94Nb65tt9HGVdxPCn89QO1+3N
VPQiVtZ+IL5Kak9W/FeZMrd2JnOA6zAXP2Z5HA6wRNaeETdF6nBCWsuwafxgJiyw
wDA4Yrl1/ljUqmnbsNqGHZ7V2Xg65lM+tcVQHfLPP+UWksi26CzksKsCY9g3j+hA
k4lRzRSHR8F/GeY5w4WBJfDNwymjLcYk6XshFoKW2iu2QDeUat+myKn5LoOOLDpl
UIs2CS8Wp5bohEli7XZleudFNm8pdS91ojnOmG7jPqY0Lm3rGSdH3/87Mu7iFduq
qL/MK8eBvRR3XLYceD1Gsh21+2r1RW1DituDyKFYlQCSJWacn+envzKbhx2cdihd
DBOO089xURxcY3y7oAddbOjfe64d/Bfidn9puZUWafROzRUjT5VYOwGifbzSwc8L
N7MWtC5TY8sav4FBGwXufsG1NXPq8up4qwb8pFY8VVsoGbwtJ1I+0do4mILQ1Cr3
aBdZ52ci4ijy/7D33vFZ5JLqOoo8lf1K9Y2tyI0TIzKHJGYCdFjZ+z+eOMG0tcbB
ijrzPva07rxydHMVtLic29G/Cy3I1LWu4FdCRRKVeLL4+NlPIO5gv4OrxAg9kknB
9bDl84LKRd5rES0iTd7CMnmvqh+FBEBCDaaC5TCo3nOFwAPlJFzDqGjlOwyoODJL
9221WyOlzgmoYNdeiEzZUhZcPA85p2WgjlMZcNLsFIHbUfNIYBHqNOcVg3gQBgqY
Q5XVxhq5OKf8O7suAPehnVLeFPjlGPNAOppR4T2jGd77Ez9UxLk+zLhtOBmbW+7c
/nE3JtQwuMxz99+ktnOPntcbAs2C38NQ0o0Z2gEAYA3fuUCawr2GxGM1fXAOD/hD
8o60S97jQBzq4PZiCmmeAemvn5XE44QfbM2jAgyEufBAx7y//UKd6xO1ATZWxsuf
RDuXXXv4sWwT8gZhj0VyoDQS+mnciZ1vAxzeYMgxspYYsnBmAxiLsArbbpIoMXNx
UGq+fA+nne97+4JEVw8GZj0WPegkUlaCuXRXVE00VyekYZC6HAmH5txeloFHk4OU
vkbZBfKGKX3qE9A3yl4NU8S/A+v/qpctFs6M5lcaY6+FBf2oszmIwkZyeokK+0st
1YPBB4IGv9GKJy7zu5ZGL7ZbBvOnosoyRku8EkAA1Pv2nZwq+f8zvRej6b3p+Kan
Mvyqonks89BurdfMnNBePaGSwQZ4yOEZdHPLGjjO6twhFxqAtwKUH6sVDH6TBRb5
xP5mzas/T0PM0Jz9XkBesKo1q8zAPqEC8cB7/Vlp6uC4JVYRQBiLTI2wvbXGfsTE
EG5SSUqEwwpPnGPFaLlomyqrNvDaOG/aIPb/tAcsf/tpy78ke1WPwvoaLpOWIprw
JJr+r/kgLpHoMyl+vUSluT7sJAg5dOkNllrjcI1RUGozax3RNQ4roOKdtijZ2NHj
/ggbFDW84bFrCjKH9rhy2Ql1FbL3ge43DqzdFxFSisHICK+0WD6WByXVRSpTO94X
+fq58rVQRYCrHCKuuV4ceT6nIk0WnN8fG7jKfjq3eoA077QP3X9WDwVS55u229u5
sDx3wCMYLo3r082y3oNLJjLCUw/kN4S5fqsTkxM1gEc0RFsHa+2Tnvi154cbCKn0
zuBgtMf3v1Cj2aj8Es71D8Wj/cq/5Zw605LiZh7UmgOg8E3bg2xF4EbximQTsczl
96QvPESy+eS9Dtm50q1QLoX4bRm6dtvp+9An0J0lzq6zsvnOJ1xwlpAc3sncVqR1
C9jlFeXZfh6Pk9yVhkbyCOa69ASc/kfaSdtoBq5UuWCCGMo362tuiVtus2ZjSNBw
eDXBqHFFUIUhzEiVCMHy2ez3KpsSZOYVE6yjbaOdDKjRlYjSZOAC9Txj8G/QhR+m
QEH8aFQvJlCdDj0LXkO11qBBDBi5cKM2i0DkLlU3i/T+ICkfjmZ17UPGp/D7DfoB
jqrroYGLE/aeP9/x3DMON1kgEMdlHHHqEHukNmtxFCQQtmFts3H3zjfsDC8HChUD
tFhRdiJjiTSr9Cbdj3zEruIm13/+eYLg/OgSxPCgfVtt6ieIXFKZFbrw0Ll1fO5g
BotJtJiGYCB2x2ytV1tF9sxfF5E4NhX7Qz5ON2n7z65piGjCcTwZjcovwSqCQmqM
Mc1PHAwI06m+hNvfO4HccBiZu10B93RPmO2lm/jIqELGRnKBy26ZHIHL8nisd1nX
sIEZo1HNT+9afRV9wkqR/B079RkaDgZPySwh4/BHOMJ9FGdxWtYsB+Acy5wZUODY
eoPSfAIOH3XmDNNCXrNLzr+rhTEUTdVOtsyLzdaso5Exbw36Z84sH6J/E7mStx4X
y6LtxcH7Js8r6HTFtSfAGBIbqUZq8E1j7S3pyJadvoUesgfvfuhyNCTikDonAdtO
DXTOhGmjqtkfp/QnGZ0GrHgPHOdXsr3NdwzaPpWztxtvHDhuB3ZVi337/EnjYK3P
8fcIqKROQrnheCg9KRs5NPCK9FQqYS9pfDxYdbqc1Gb8WwPb3Oudx02ixFzbvx/g
k9XM7FUYVp5Wst5YihLmIWnKWHewkSVz1RYHXvsVABv9G+jQGvtf+negmX1tRB7+
JmF6lb1iV+SVqp2tdug+ZFoby/CjL4T6xdoVmkokV5YXLFcWsxUUEEmuU8WFZx1b
2MMM/CbiUUGZ01EGszLlWKdjtG5R7PF7zTyptnJKDqwTaiAIR2hmuZAp7uLqG2ad
z+wrmvfKfzJ88wJuKfEkpG4fr1uTpe9kfBMLiCXX0zQ7tUItUwbXGoU3w1JijoAi
bnsibeLTLG509m9sMSVbVd/B8rgDTs8Vmgz+6xfoWNxfWPuvTS4LtcwdXTeX2taV
17w4k+scAZkoKrNpTJjS/mWbMoj9h1LKjlTwaGTBdALblSCCEYKOUn+WLZC+Mn0b
rhq99pmE79Eu6ew+2+UB6O23TDcW+Sr/5C8jbNCuVG4SY2QxJ7jggd7URXWQg43u
90hzHXvbjVjPf+XctcPxND/HKhNk6PwmuacuKHLceZ+sWtn0T319201E+wZCLgKu
bxYwESvWYmSLhrjSif84vcSbNScgIruyba3Jolh8e3LB94jGBMT6MB2HcxSME8/Q
7sl/8LtN0VBtIgwVJu89ZHSRtVbeyJrKh3bx2NvmdOXBNugOt8ykAO5/E7Cp9TRS
0vWUHieL2akVGEX48ZDu3SP6xw036H7izYbJ5gjJOsRccLFvmW05jHksN/tmeW67
AC61OhYC8uThB6tDCTrZnt2Zt4LzSx6I48y/AlTw2/8QG3mPo7/n2VCEDWPo6i9+
9NKTAtNQWUni1q4C11mHwrL4M2ugo1vqCWcRU2SKtM2zgO32ytLaWNEsDG9GSzjL
W6J+S5eZTOMLLFM45lscboVJdVxUHWDrhiY+WPSQHz12RfNgQpi5Y3N4ztoB3VtL
mwRJUCct/ZK+gDhFWUkr1xMHuVIaauhDSofHxoMzEkMc+qpKYluDAuBWzJ3AN+Tg
TBR1G+65ECNsn7INnefYeU5TGcucZSH7HuLKxIFaq2YopLs9W14jFUKw3xDki9Yp
HsaVvZASFRmRd64ZKfQwkPT2hZ+IdHLFG/YE4MGwyRPUOicFV+2gm7WM+kxOjYA6
jbybkGv43Vf9N7yh9w7RP5Bsz72fGzl44zxwha4gzN6zjLqMi2JvjUX9nvq8Wsj2
lP4ewlT6kYOsTfOrPjZaqjhUPkql2LS/wleaxxVgVyPMbBfgRgOHXIcQVf95tSwn
T5JRPqteyTLBLrtilDf/KQro3YU4vV7IjLKcOTTKNqBeac5zzalC7nrWEWDjw3oa
wqaLH/RxsPssgdJ7qAvAuZsSE+DlukmoY6+aSXqIb71D/MhjlvtRs4bgPSizpGRs
jtbwnD2qRt6V2J8uVnKB+qlfjLdyShJ7pZNsfzP4UnglyA32hfcN5bs2+gH+RBQI
JpUwOAWQsSWjh5TPERpw42si//2BMLqJ6wbCv0oKfJvkL0QT8JPaZN5IfsC7s1Po
BOIOIGRsZjxaAK77mhv008StCbDuGJBeElmFNB5CYo9kL0JnqBcT9gxI+L0wSBCm
YWsTFE0npRa4uD+o4ixMXO9u2wPGq+g5Iv9gLaAafJpRCPax3/JQeRjWXWZX8n4L
dDMcspluYAcFCohw5i3NwXjwAeqaUHFr0E15wzHNIP5gViJVPRKfpaeA6SrFJVnB
TX6Qh7CBzb5r2mCuxyr8FztCAHgS9CGMfeTHfmpRclbyVuqAKXfT3XpLux8qV+HS
z569QHWfPb+AMwyPD/uYgyytTrcmnAiERwJkX4JjrIikRYSA2B0QgaIpUPD0aeCj
S7wIgAgxQ4/2J0AnZhIJLGiSbMIzY9HRINzGPM3rqBWrF31FOEcT1CXn/BU7PLC6
PsbKoqIJjGhtlyVgtDeL+h9QfHU1b2ktbx32kNidg4s/h41H/bwpgdmfK+JmDstr
olQkpZ7WMly3vW7yfIZnBQHvfndrwVXZWhCDD2CjNgfNJn3GzBuaClWtSaInBF/X
D+EG4u8+JFORFrFD6tucJMsWud9Ok6uFYINmxVCocFn+1smA3LgQLK+iSrgbbJIL
jw6nxzwQKecaDeiOSph3f1w4kjSKmgDswLiHT1ZpSF1+/OFGfwFvdPATJW6LJFZZ
JQRAd9FRK+AHj5hwnHQZHjEerIREBp2jIGHy0VYf8IwOKgmpOFK7TL3o+sKRE4WS
1yZ1KuiFW2lVV29CszWkJ3vHH+Iyzqda4VrxJwiz3KDNmmDOIAUI20b6yWZYY2MF
+W8xDjO16uA8/peBNHpoDlS/bT13FCG+9ujh0z3Dv0k5irD8Eg7pH3x/4FPoWeP9
csF5OO0xv2Tss8HfZVXt8VpAt07C7W7ofGYWnmgWaPdTMGlAqVKUyxKs6YDT7H6c
CjRruB2mZ+NJ8PPyDlvayzXsAsDuQOrTmhibEKokDgmHXoK9ubYRkuADq7jHUJqD
+THPUvwpr/eEVYpnbmklOAauh0L+9qp3PlQHxER5k20Er8QHJwbHmbIKNtHPw1Ab
oAz/RG4GhDckK9FmZwU6OVuFDTNP3Q/13xdHOWPPSyB6cbbdFoyWHbKtI1FJciDx
l6hNnmBUgHAqYUxB1QUBDGTfrLM4QqgknySVN5Oq6YakmUlp1Sx+wK1qOTLLgqol
ymByfpEfK3aKTQkahjctHkx4+/YXnKJh5BfnZutm/YfRNr/+JrhKjO7+H7z8xX/C
vC1amxO6WW/y6MmIpK1JF/HdQKlEIJe1ikQW8hPP6qh1Xd6+ijiZ6yAUzGr+dODr
Brcjb+4jD3aCo931CBEs+jDS+tGPI8yKRy+7IZOgQIlU56HNHFc5TbFljKdKLOpl
JV1Zi+cTpOIoTeiQx1vBZVGCDQw23cFXtb8Bk6jYsSqigTjpQRx6sXHpcu5Mk1Ya
LxdlAoNfF5+8lKd0ON7GQfg7w6GbzfCNcVxh4EooClU2oRxL7gHHjXTBS97tajDd
P8ROX8FvNqXNQDlGExhKb7chJ3yO8TEyK3LaTgnwDkhfjCGWwD85tuQooHBFcvXk
o1UWZU3svAuxkb+n8C+VCUQ4iScVgEQzTDKO86wuZICG6IS+9qb0qaKvQEkcfIA+
dkZ8ARzNWeXnTioS36eydys70JMlM2iZ28vFPTrkyECoi7ASxm/d58mx8xPHjox/
CmpjLr/fuKJewCGay9acEGS2T+AT4mN8MYWzNtoujkZNNOebw5+GnbSy0RGCTqOs
VVeoi1Qnf/qcr8WycLbpYIXB3tCRtxd4EHypZRPq57oOha6oSdsHg+gUk0J23lB0
kvnexwMJ01QQZigsGumGkCYm72q3Oy7kXfylzH+VdKRUydFJGxeYDiEmJgdRWm8Q
2NSaTExkZ8X7eXOGIzBohO+ho63b4PVzJL0UOWO6wgB31nPfgF18V5ezbjE2Ka2p
TQOUKKXeKoEH+KhSUSlzwnfv1Ebdvh1RoV4gIV93+NzRiwDxXmpCyoUGM4cb20Kp
DKWhfY+RYAWtWgYwuk9xZjjxlFtGaTUZjZPJJ7R2T1XUPVysJSmZG7ITY0g+wNBY
MsIMma1d6X6Y3yJ9TPWtcAAzWFaYTyErUpEVNvqz34zpFg2g/iOizvx01KNBDzRV
xvqLYjnW8ltsu9Qn2cuuuS5WcLOVKW2B8XORi6yNz4wARlcEy3WYn30iNvwlbLF4
wkXVXXZc3QJJ/BLt2vCvJFHXbePnycpI5NbmAX2mXESqinYKiYCWZeXywCKuJFs9
kbYSnrBoB8WbzFPuUeVDT3Zds0cjTwnwZ4hvsSeSgnTVvm8roW1xYVDMMsdlcE7w
EiICfc+Gz8vHxBBqY28IVlYG+rlx8x/dDmPEpSXFSK1Pf4kzJ1QnBh9qEhj0Mm5x
5xtY+G7EXcoG9HjCWS35pA3zi2axZlqWIIZ6w0vk+nMBhx9oKKXkvJhiO2FgvIIM
vVSF3U2Y8R1kRTzmmfsTJX6Phln1oCJF8QxCjS2CGd1tMSX/ESe8PfYeVngiT/Ae
ADmc3N5wJmsoXjk/2+gcdwioT1RBFdG8KLAAVi0no54OYgPbgsJQxQgfSjTiB/F7
3TAbdH+0xp+AEHbpssE3xzYqGwFh94w21stWuKQOIcxAXMTWBZwRnRvf9Y31JO9u
tfdWBqR2O39E7wnjCMD5+PXTBJ7qaymlnXGWWH9EbdQPj8DypE4zyC+wPeMnyDH2
CEcRwqk+S8ryWom9gl77rryRI/2E1K6rZz7X/p4GkMl/A0QFF4AERw7PCVj8C61i
ioZxvnWjrKN+EongtiS4HyVcFZEMe15Jrti+zBZyb5fr8Bmk8A3Y+dzFKf3kcI1F
c/8bDtoXfpE1VGKcJbKSQy+QtSEiic3rqlsS6ab+CE+YuVwNAdkQBOpdFcl1Tfqz
7K/IdH5Tx1N4/CqetmKnnJPf16qhsF/svbkBo8Kjn63r21+DbPe9zYzf1+t2M/id
u1SwRf9N82Kuuim8uyUdVTGerXRgAuEG9T2oOk5Or5qHQql7bCOdi6af+W6qlBUr
uN/2QZAOCuO6vfjcN/ytHOcNy9lrczTqCVIIAZz59EVOG/LrqecZeWhmdSRwu26r
hQRcbAHRwwYEQA6UtdFqz/lHqpLGE7yXuLXeo1LvJUiML1T1ssuIBm4x6iP7CPsT
JoUvkXa4CGDys3E+P8QvNsuRhiMsGVwY4FgVycVEXzhTO04SgzDkHEmReMvhZemB
nDZ/duZoZn5cFbU44pnNpP8/euH6bbxULF/J9BYiCwkQaZS2snGZ2aW/Vjq4PcBO
8Dhzm/7KjTBPGs8kx9HmZQSlg6SFdt4rxZ53misd9aXbgz8xfdd1/D7ebobwGxgL
XrEPj0BYJ9r3N8gtR2p5cRJ5QNghwNynhbV7/hND/bX0yY20hnMmio45PG9rfvKo
t17dC0smyys0Pi92m+dhYPC5or22gCGYZJgw3U9SgiPHDzr8dd1pG0mJf4LGKiOC
kLVpkagpIdFTDl+usIS8NiLvugPpb0BTc7H+Jh9ESykG6ng4/uCqryennpvaWKJl
EuiIOLISLhPEuV2wiHVOyB5BdQL1wbxQsAJZferY9tgGzJ9acsQIbgQwzyzo5c8I
j1OsI6MZef6Q0xg/Y72s4jPto9xxc6sgBqRejK+2Gdd8gVpKAEj8JZErKGCtAeSr
1Aiqg9bgeUDyZjmAygJL7PoYh7KQg7hlAQqyMlNRWydhvJxYlxL9qUi1BmgB4L6l
+WdkMSL646Ec2A67eIGhLlfa1emJYKNwFPKPRP52daJ+YC/NHh+SGheJg21xr/1O
9Cex6N3s8kD4u5NmZRG0lNaL1YTi07S2gy+2mJa6Qc90iIXeix2+2/XNHrhw14k5
n2A6zcnBxq2N5IWbEQgBOApwJASMEl6546NMIv7MnaWhYXQkEr0YZ55cRhXOHFmd
Oc4TEwCa0e8dWcCMhCKKpsBbpjxn95xOxB9pXOpqGwf6zKbb/zVIFIc4RsYqHdjI
Yu1ky7+W7mHU+bL1FDl4eCXXYOzsf4eB31IOK6H1CTsdK99rE7bM7Ks2BnPDqjBA
e4kIz11XsM4NUcxExov7S7Woy0AUoQjc5tDavX7Xb3c3VjlZWf5Is2dlc4+stOG4
m8GJEZyfU75foQn5Fyz1f8aF+kXvCwjfBteg6qTKAy3CshunPKYjjuEXCx/2meaQ
lhkjIzaA9kLUMA5eX6ItExFjMGnVjRlC/Udi7MO9nJLuu7z4IAJYUVOJ4AELIaof
EcWwl7eBhRbxgoCXbVagwVQB49epxc9l+jp9QgCFjRfzc23P01w1BMr0taX0e2qj
bMa3KJLb7QHQ7pBEk7UFCfaawKwwiG4kmerhWO+8gFVxF3Hc8oOEabfgL6Pulr7N
gBotp02dFrM2UqI8Uv6skph7x0DPeoTweszPwhMQ08cnZSoQvFoxuUzagOONSPt7
zObRHlBKaPMMwCKOYWWzxs9Za3zGM4hCONhSBfzmuNczb6mgvgRlVbqfqPOpxkjG
0ulgVrxmHide3MoGh8tY22CWDdQVBu3jOO4Lzn5cNb3HWLLOomCUXirMP8AzaJXn
vcCJsTXsJJ/Q2AfD+HQ8EEBSRBvhOe2k7sPIBQpxPfGuRrOd/9Tw+L0ipFh3hbIa
uRSFBAaDWU/l4bozZNkFpfO15KzMuMVOILZxDh+4mPGMbLWflGJtUGu7HBbaA7RZ
8IIqwaqIQoSgBvVcH+Of+UbXFzSSqsVbXEGOA9Kh49xM/oTNvhI1BtEZNwkDambw
gXFa+HPejuhCn1ZaWxqyDK0ybRnsqMHugmGDM2Al4ZrlE9IKQ+DmschWxp6bmHLL
2R2eK20C7CdyC4Wsl1uKlUuBrUAq66vBGh/Zqm0FEMh4HLfcYQUtTkEi8nBLpJl7
zdPYviySYBAxLom8VFjtnHP+/XSW/z8Nqp2E3023hZ2LVQ/YpNEvKW32WFCo36/h
j5PakeiAVpCb2X8QyoTPka1F3QDM44lgH2wNARsD3CDR6nQxPrfOtcSGMXCzj+B5
ScOfq10BtHVz21yY6WTVYHntu0zW5ciZioTQWuvPkRRb5LbTbnuLHVLGnt8YryTy
kDEeoeqKdlkLK6nuhfp95QvzOyaSFM76oYrQ30lGCeBxkfJp9oaCcCmJrA0zwkU1
vcWeBvUyycuWxzoT6cERxBWh9cNUFH/6UYIEsEC8ZBRZuCyLLA94BV3wgaNGFDtq
XFeNIuA6BNDuaij/z9ZDnG8Ry/Tk9iS4G958mna+yr3NAmHAsFWrH1ctgfVawL49
b2eAYKl2fj164FSG2vaKwaBT42m8OQq5udoN1yZh5hQrFORJwDRX9ZF6wxxbtqtA
tIqM7/LnGabklpg0Jq8W0EsBuIv3zp5SKkCTy87QIvPqFrivKoYt8Hqg3FMlfBEP
mTucvJS/hCiYBXUiYKt7KLVkYxVwC37CjWj3pmv7UjNucHAcBm9x4WsEhx2pgDhI
GfzZTi0p6HsaNpRW4+jfpLLL49QPhciMZdAnMaGrmdp77sjbUu0HtDU9emFmVm4n
ojWDWtJEn2o06+aunkSnloguLXi30JhV7jzZ01YUacFwfxZ8mQIdfIIGpAlu4mwq
nKciregK92c3eGcJq8mtLHifsYH83g2gvyA+sJMsoxAKySgm6apmUq+yjxVP86jf
DV3kyqjBA9TU5S9u6jC3Vy2eEC7JvWBWykdIlnac1KUrCky5NbcMZ1QW1KbJ4IQG
tcrgBFhIbETSi0GV3WfMcUSTyhM+tN3cBPbn6SpJCKikfH3OxBie7nWPL/A6mFpJ
C/Fcy6s0EI/0rx9n6U9z29FjdyHD827ZPvMFONAmqYg3wcY0MEF28bcSWYONZxkL
m9cqKN8NrdDeKuznP3vG2WGKXshTQ+DvTvDtDHlR+Ng/Cp7CN0CcYtn/2zvIoUsi
g4+M1KxtkLNPEQqFlEoMRGEY38WClhYqrDBwraSmdttFGw8JMPXK0vyL3QC8MEHD
RuSYuOblL08woORTBYPFpypR2qJQbZgJKd6XOaI8PuktTbqxphpiykLWcSiBssNv
i6B99b19qn/jetXs5lOwlIaCjlamN9scnqX/zfO80h0SiiBz7Fg5b1XOhzKt2AWB
v2YEhaoNewUucTRbr+3ySxkf5LVVKU7hnM9jA7lCYDLzkTK2WbiYHXoAsUGxJoYi
b8YJV2eZD4FqPb/1FRPvV5SrQ6mhqZMfaAQ61p4q0uPjGPpBzQWHFPIqei2gFoPD
Y8L+x4SXNFdM+ftFISvseyNVBVDLauS6cL5vIw2SKyhJhkw8zATG3FAkr5/ZhS74
2ebgFsPBJdm8nWFKAi8Ol7/1Iqhr6gOErGV3OSuyHeHsvBn+YRxqBnYSLa1O1sVz
dw9rFpjXU9pp5zJeqM4fzf5F066VXbGGapvRbgvSteWExCT1o0hXqFSpq6+aSHSA
E9nUr9xu0X2dld5VKKMnwCcqU9mOd5Cm1DWhrThT3RFgCaASPg7lhra1hiyEQ4Hv
8kDXFrajAsCmz7iHvl/gDwZxnQ7BkImm1OKhuGozlDbbd4SI9oqWaImdXZhXng4Z
e9a3pUfRP6zYaYRQZJKYZxZDewKELL/GQ111RpX5iKsZUKG7Q/DxxxV0SzSyXljV
S7hGFeK+2xsfDU1mx2TYB36VLvv9DsI0i8TWga9AIoijVyeKHauCP3ctKMYy28fA
2fYIO7Vuri+TeNABS/IjZyedIqf4Y5sh4IKQyDdgZ8Qu9/ZN0ob+NTkI9cLLPcx7
WkifhpoNmjR4etW8jfHQoMWCTtKi0Bmk9yv3G3Aqkx0Id89LOcPr26LdlcZTtPc0
J5IUppQwZxP6exbSaylBU5X3pSIlyERYXTeFnfeJuWFIXDSkfgHuwMKp/OLHHacK
eMKRZw7iv0nYVcADonYTCu5EjIIWQQ+9imQuHMqQmx/ABUbnqu/44AFRZTtaw78t
i9FL0SJRG1XoTTi4ZARlucE1rlsl/Qh4EauDHaWeu9h2F28seLmdRToJ7HwgAEuH
1OfmtTM21kp1iP+w/k0ktkchlEAOwQC8xAW3ktS6L5sgOzxfvPdlfPxivx8lFS+5
530hL7rSIlBM3FB3m4tbrm6KAB1RhvEL3zjSXBsjSYAlEOYuLCkvnq8SaJcqLGoi
7T6BJ6aYck2hZQuRhAmyy4g+A/e2JgVCyWVXbsnORZrg15cDaeihkMsJLxCo7U2K
B75nGoKkNwkMDtomrFBFKhaDQ/K0kgACh9EFFDz6WyP/bAShRGeI/oDl5Y9NLft4
KAdPsUPqgnCjsbECh2cg0r/LLovdHiAsGWL5nktMKo2ryNgwD5WMi9Dd1yDfbCsf
JmcqLbc9DXNskW9P830j/eGN/aKwR78ZcoRs5v3nLnw1vMVLVquKyoTgzcxtxiXx
Ut+6UrfGCBS/FzQAuHrY360ezL+vSWqxOLWM4pEzoG7+VhX9K2pyPC5cuwueSEBX
+KM5myjiKGusTSY80miAzoF+dOkBHegFlAtQer7ViCzb1+MErjKYkzInRy34I7h8
t3e3MKnd65qjPHSJAMnvoz6Jpk+v4DMUQeh5GK2evLmsIjuyN6bWhtQt+8juL3fK
KR5Yn+irHWopwj7ahKVOMkD5JmFwRDhilTkiSZzikaTIW6y0z4h3fPBe7GU6dqwn
IfFKwi2zcndBRhtLeqa8WWH/BfIAb3rpsWhHZSvj0PfZ4r42XFQpB8V+fQjtTkm+
VoehvvveRs4Wd/ip5m9cLM/B4xKLi0SHichNshApvJgxitDCBychQDNQXb13F5k4
XaJaknFQ13HHPyM56n48px5QXmze699GZ0OV2zq5/SOF4z7aZjBRtPh2qn7Ka34W
gYeBoaSt6OXXFOwWAlSGYXV0cWUDcKO5LkWUBEBkkS5Di0GdCNID0bemI+AwDURK
N91kwgopdopVljpTs+UsEinRSTblsQkI0H5wsc5aW7+7M8sBeUJmDrDr/z5Md+hL
XXA+QVGbSgmtwRqwI7IXJEag+9uAs6XI+WKseCab1Zqxm6laRDsYCBBUAkt/kmm4
wOW+fElx7uAASoksdNuiGbDZnQQRhKruzURmJ0BawCcCz1OLPn4H5mYYqbGOOw7J
FtqRBYsgogoNrCj6kO2qxuqRpQBqvceFf00f0+zG6m8gqhZcupOhaFsffSK/H6gV
8vhd/fGA5OktNRUPVBktLxKdS9QhF2uFxy8X8t4WWRTyR+LeaRbhT/SHny8i90Jy
PJRvq3pX2aKe1dDkIZmSQMDHPUP1nmT+6FWluwF0KQC8ZEjNUpflqaHH+36byIP3
zI648wnBQDBFm3ROh1jYYm1c8juFbNu6tmvGx62fpi4STiri2QGnod8vxqe0CTHJ
YJxcm9pRi1WhsaMDWoqBxqnu8INd5SU25gqVy+gMzAp2crNoxCTSHbMPlXSFQlXD
7l8r9SCbYPFs3srSK4JCgEVn6lfH2WK8bXw7dd7scW773sf5Fu88oiwqAIVHsOUG
wShns7K7KIqCbrVzorS8t3WkzyyqBsQmUNz04Y9PVMLqGGDsDnbfeFk4zCNTMi1F
utzFbxlpRmc8ExAvR8gPvJNbTTOmzV35cVE/PHFq3sPbeWhZbNlVtUka1Nx1QykS
+OXId0c5tEvmEzMLKSFG1ZQryzho41FB+bamVLxEcythY4HM9owzH4N9vgC5uoZu
fmVXRUmFkLB2PySMDaLgygE7MZDTNpX87E9BwVktUggFo3ZXnx+s5kAWHDCgDxMX
NsDrGw5keEgnE7cemipIg2+ayi5+TTR5aPwPVP6PhXObjzBf7SL29u0j+RbioQUS
O3r/XBLWkY1eEoh0XIfGfwkkKiRTMPeIpjLeOMhblN79Pv/fxpWw72AEjwZ9hq1t
c6BSdpqSK/yTD2+GbE9tppAU0Jk7yqghNVZDQyazK91dEEFtfJKbcV1R2IEN/WWV
5+HVSbyFfPbxe8S/8VJrZxtVEWAO43RZ1L7WfYqpqWBxTY11FTVjBmxmmp3miXqJ
GIwnxQToFTfMEqvHcPh8GW7qujrG/Arc23/krgxAVKTyHhiS+XlJk6TA5M3n4Q6Z
5lnmFB6GKZMsyupKmrEdCFfFGXkSKM+kUEIxPITXK776o1nxlR8QzIXlPUKShpPK
0yJOU7mpRFX8NRrImtaIc4WVfCVp9649xPZhX/QHc3zR92FwoJBsShxLkFbSS4GH
ln3PSAXc4SUqhchCy2/Tx+jMKdo1EudE4g52Gx+6uoA+7i5W//r0UToHbtLQe7vd
SKL2CXw5MbvVdrWUtEbEQjpgaBfbqMNkzZ9qee+SFDIBQEzoHM+jbpjdqASYe/wS
+DDbonWTzdjOSrjeLnVhUQhmKdCH674NZKk7HErJDBegJEuopaFJVKKLMMVv9kmU
FLzUvHufLnA6yHPQOkklD7FDRr0WWGjJGp3sU0aSPgSk0PWH5IYKM0s3QJriSYnt
ASmzVxgTuq3Kg0qbM84HpZdyU9vtQDnR72VaapdOwPhDZRzVOZgpRxIDMmHD3QRK
CGLtwkM/OVS0HwrM5x3MOdTxpOh0uN0wER0sXRXPcdcKLHCkqNypZcEDrNfs+cSF
CxwrHJOlUtkaAinktO/1WusP2r/X0gmhLuroajyWNZ+rYugv4GFtQzAbfwxXjiQe
nO1gr7waxH+Y20JX82b0oD4wQCTW5NQ0d4+hIMdMztizpk5pQ4zXwF8YwmHNIqZ6
LMvSkvv27yG6f+Jcib2d8aP1mnRIFUNNwEpa8gL+hHYd+1DyLgNy6V35nkk1AnnG
32zhynbyyzeffpvPNQcOzjLLugPzITfPP/xCw5Pb73RkvcqtRhNEMqpPPwhW3D/l
K2oOYZDeHPvziYOoIq6Uw3AWSdm1mFJqjp/iQhOhevYCuUfE43h5uG+mH3sqCobh
zWjh5/aoQhW9gxcfSI3OK8aqUDQzha3rIJgugnNPhwaaGLJjrC9ZLuhFLxC7sm6Z
nBvI9pNdosAtdWjjDuUssUc8TsMMNpMrQkHEg0lLN5kIapzJWTx43W4HA0cuKIOp
t1pPHM37Nck2NukC8ZP8yoXyAy9gltfz346llz0MaW7OyGBVxp1Wz8OYvibELJN4
7m4hxuBnA9DJ7EApUjZKezgBzpgGd/quLcDWfD8Pm1HBS+WOSlX7JcekYceljZJm
Nf9QKXcBawgyVRGyoR7l/8saONNue+6T6KILJeXTZRmBVMwpJHah5T7buWwtYeZ/
7dcTo+e3+GbRzj0BwTEu860XJ1BjfvSaeJV1x/ZtKUhL1VFkVbpX+1yaZ4M5H/4N
RLIllqNalrgEY12jtgTrZGN49JyuQkVm6i12aAeQGTHH2OxgWd+iDW3dTKHekF90
9nAOHe4hoFW6Cln/q5tanadYN3OaW+v5d/CJzb8kXiUG93zYzeK2yUg0Wqq0Zzc2
WkhDSdLDvQaannsngvEyymQ8hBnQE5WsKFOJu607j7ViLLf+e6E7eRHyZEemphnT
s/sCqqtk09Hiezy5yuQjjvwMc0PPKXJdkL1DiSYu9bV92kx/3nW5be0vNomEVJBB
ZFOLX/npKW85R4/29GC8DYYQVAG5D/cNf2W6BQr5j6CCZeFiPzzyRG6wXPFyi+ie
qRMSCRQwASf1rr2shLPm+gMZoT8M+AYqDoJzq89WMJL4e6dPl/tqzVGZfUWvuhnH
krwQznRPTQDSAAzJWoy57Xurpy4+QbzOSkPd31ILpAeexQvRFDd4wnbSBMU4WcCo
UU5moglKW/lGl6dpdNSuJDPRgWFoz+jnOw4/Yb4l1EKSHkTd/9ZtilHTGYTURtLr
Hsp28+erFkuo+TfR1tRSsqeRzrmpM0+jtDJC7X7zpZyZHFOrSQHUbhUolO+ZlJB4
ZLO00CZEHvFp+NoMw2tS59zVfKm+yvFiXuYmS8Y0LJIa81myR13Xxh+SV39jzuI5
iQEM8HOGs5Xr93PKDF+UBl4MlU/4yPx9A82zhwZruJqIQBWt4PwL9C7G4ydklc1d
pcZKmx/eYBgsf+xMn1YXD8nyPyxYToC4MIcS0CQhHSzQ38HE5+Wg3W1s5nvaILss
NlY0wzZWn/ji6sVOkJX75OOkcbfuCUtyTI0ct//3QHpxqMHJVQl1uZo7ZDgTCsnB
xlUHJ3njotVgGHNGcYkbiQsiz26VWSgpJnih+y3EfnCrCP8gI67r7FiIsrGTUW30
5IA98OwTD8+CxkRX7XFL+FUhjPMaRbJ2yrbnm2hzE0F7HwG7LvWr3eKb+fU7JqBN
naRboL5chGb5bUlmWyVUFWnWuZQWXvhQhCmmyew2SYEG7BZ8JJ2luhPN5D+IF/tN
jTsbm52YH7hucIfTsc37J28bTYPUNfWlOHXeBz+ANbFrUYAEfqPBZvNeuiwoBqeZ
aluDGKnlVha1IackI813VsLgsU96HlTrrPzlY5HWPKObGL4QXmzKyFQOsNVwMPFk
bUChdm9bx0e2ieKOqq9+DT7imgNCI3L43BoVzTS9KBBAt/BX2na46aeSXa6M1e49
Eramu3oyNRDbvIJmERx7FUEEeIkmxK1TdMIOwdwS9NVZ1xEtsJ2EtbVYLE+VuiLs
H/36XvDj4ua4hAXMjjkrw6KW83aYQwUGuNEqAGCnIfvfiLEMguF1bofg7A6rNp2r
hhTxHIQZ4TT2SDr0E2it1O0A2LFhyc+vZdtA6KIlIFhenxl6d4jRzLZeRdNJWlFc
Giy8MlMXA+07M9NWusGDv3Nw5b4g2uN671QiEZIHRJ9xOxpPuETWABUvxDc45YEM
98y7c2TC00UU6aF0z+xjMFY67MA0DLBpjyKxY8Uths6u1BUIUEqcpTVwoQmMh+kX
hZQZwgenwmOSgOt/1IB1Aoafh3yf5uzNuSrnfyPeIFzOPo/ciK0XEsyCWkLeq8Xt
jE3k8toARTx9/AqMPO8enu18IphIWbGlFOCMwQWSkKHfzX0bABh7JPV1pMXXQLBk
a25LXVJ76yoOzx4mdNYgb0sRBP0J3O6MJFvzaxJ7vf9hrvjLMFKCyrGBoXFJwqSi
V2DJ2DLXUdXoKJlKfbQ3/3KU8x6LSygaFh3VOjmqjgoibkxlMeUSbQVoOdlOsw/t
NmN/3aZm0iU5ZUZqi71u81uSleNplvpDu2KYnplHSH43IxnTyIFIu/ipx60GHg5x
81Jczoe/gr12VOuRd3yEetzYf6juqDcAXkkWZfYcfXDLYjC+xMlJ8jsJE0jRTV4i
EE4xfsu0BjAYgB5r2oDPmHoNZpN/rKET1wvXxOmI0TBMI2d7Ep2/WoTY2G+fSx00
vpDiFKDH80abruE1S2JWQM0RcELxZbNJ+5idn52aUaVw2XLfPe4eaAXW6+vRiiRP
1toFnE79erCJnkZw432dOFoMD73r8krKdE0ktp4PB41CjW0awel/exJzxBVXiCSa
FDAZAD2OiJPRlpXiNckfODFL88fU+cLXeFjYleBCzGkIsOvUrUF+fQPqH4Y6xkXx
A+uS1Q8qWyO4W+psGb2zQpuvdSIafQIhXDQdL8F6D9CXif5Fy2jAfmB91tAhvQJT
QnqX5ejG9lDJhfuqdV7lSATXiUmCabP3MJSqxqFedXYrpv9FClEKIcFoUOoZNY0/
+KlcnfdIuBlBmkTgiMY+hnwXALhvKohkfNsW8BJsFNrFbFdw4K/NxuUgbDhkjA+k
FVVePggRpaTkxsncFCHL82+oU7IeIIj9vyfI7crr8KpcXso/+TCGU4zjQWBMJsRz
Ox37S0ivIA1zvZpeIK+Kh1FYFz129rbDyaW4/IyQ9BnFkgG3m2m0uQUCJ6FpubDY
Lo0yWSZBrIL8MXlduj6kc+Xv8TzvzYC6mJYc1Xgt5Xgu9eA0yfsfODSqnhnksAHw
AdPuwFj2eYHDYtCna+Wcs5so2C8gdolyEP3TJl8AQ+2seQJZSsC1dDBCJI0hNqnf
n9T/VRvLrR6B0ZIzfNcxCJJKnDM+ht1afsWfdhrwGl0QcLKnAs1mcN+J6ZSXPp4A
x5Tz1URSisdWV+n+WKeJXN1Zv/KfYlzFAHiiwlmrCEZl654Ra5PZw8N+XaSzR2zK
2Vcw/h2JS6pdw6AKAipeCBM1JBg4BxnyIdxMo++XpK567opSB65Te5VDd/IA68B4
VtYkXv/xa9n4+Z52C82HC60gk8w1FirTTjRS4lydeb2WGLc5uDSOawcF2mpI9PGC
PXTvLRUZ9N+bvzqUZxZfJPs4EVaJnZvf9lfj/NfKGI55NUj+ksz1K8laRpWozFBS
VeYT6ruvSAR4Ob5qoqT7YWFkmlpOXhm64Eyi86/avdiAA+NR0a46IMCsJh59SZ7o
fP0lMglf3ZcMkzMws+WTo+TSJwN6043S+KlQcydudEYSKZzECh2+ythPk14Ef9AV
m72yBZfx6YElBM/IfjgT24aGMcYDRIITegUaQbyBRW5Xh2S9m6sU9EWXVHZjNdPe
y4TBH0K3j+iwsCvpiBPNppsWfeXLWzsd81tJ9xG/75JqU0kgVQVUUGACqu9mKARk
AEoQ4BMT4Gf6iYO9YUH71RZ1uRJ2gMk+otQ3qdlGQtRY42g7yCacZAQeQYuGj39w
A27/fyQ4aE5cfwnVLs61DO5U4WZSc9DIVyBd5szltahix4ymSiX1wtHSwF99q9r+
4BwyR7Rcs76RcN5db6sz0KSB5V2j2G2AO8gjKC9YV0pb7hbDXT7EHOq0XNcQtlKQ
ZN0wvrlkdzThF5c0WqNMTvUSFaAtrNpi6t++G7nHujl8m24LZgtXiIHSMXS4KrFE
G2dS8wl46snvWZ1FCYBq1zc9CHBDlQoW/OqgcXBvNwSSeepSE5LFxV+BsVhXSuIS
FebzmTScEI0CNN7TfNMhRPWC8XeA3eQI8RO9BOBjnzE3cBvoEvu2vTXhulNAOaGd
ZH217xxlu3OkqNPTMUXYEJjQQD+KI2fm8937k06xipAPLOWidL6RFJZNSGft2hpX
I6g8CeYIxtmxywvIwCl4slK/xj62sel9xrh/9YXetM3d7M3+jc5/DD4uE/CYOz7h
9kTajhQKceX+gE0X3RYnAtayoFx/4Ml+DG+daNlVVpOXneo/EPPMwV7AgxNQpZ6+
sY/X2k1H6JW4K0TDb09FvKdqUBur8UXta2HZGyaSKjdS4O7ZikW306ePMAnHW9qx
OCHDk09VMdVFmiiHMbSbLg/f1K2uc98ux6myIM5+NqR+gn8bPtyMtO2YGQctOx2D
TojHex9FWl3FfbVV+xmIV6c9P7fgeUhpCBtXIz4EKBB7bQiHb2r+6V6/IS/bvmPZ
Ofj39nN7R5pIeadF7pOmouOkqIpcPRad4h1R7GrS2DnGv/SeuAf+C2DNAvhTn3UZ
TYZpW5Dvqa5IwBET19Tqph50NXYUpW6W4qw0Je53qWkokAqfkJ1aV1lj5shPy4sl
ElPyAc+IFCOFNkd4zs7cdds92NE3lpLENCy1PzWOD6gBxlhqdnvv+Vxj8LrSfT+e
RG21XoEbqeo435Cf+95x0sqvWv/MxAgBVu6mWKykMyZMm7J9j8H8ZuNAaqBv8IRN
G9t5VzcZju31IqQTRZ1vnLQZgd5vhHGeYgOeYjJTzyfM2QlyDM8j6NBXN593s+Cs
Ob88Ilwq9Bmkiz6GCpORsm24nANzsP4Gk/uwnCxQqMC2fZEhDuxBabOOwIJnbu98
9/vrqFx4vzwSCCURFt+aRNstmGfGvSkiTLAlFEPIaGtMqWetmLT0xE918MbL5j/D
l/pdO7JZ/t7KSpPhZXlgBEoDtqXhwZI4UvjHR65KFirnWQbgcZU45BGO0SjGYYKM
W+by2g4C+44cDDe3282FH63jYjg47PWzOvI7xgBJwo7/9z+uxCZAvEIrBWHSpePV
1Lm79zvz/ftZzl7Kj6fnXma1VotrPpwY3A9y/MLunRLP8x7o6M6+6cdzBeZAU/PH
nwZPbE8c2bfS079DVbHX9+4DZnCNhlQ48Q3a2/HHoAj8TQJddkVSyMtlDDDOc6rO
6uftr8nsLa3NIr1iQm9Ja3zn2pQv8XUiNdwbfJplwwt2RsRRFyOzFDN2Mx26FFiS
kSibr3g3st1GICsx/WzjPdw5jtzVasQLy9jy1isevSta6sddV4gPjzuXmDJL5DOp
yc/1yQK0TEHgMFm6YhwPNfcPnJV05jPp0tBuG0xyqweyVWdb7lHoZA7rgsBSoYqR
2T1oV2vGH1m47qpT99mAtbe+8IcpQalhX6WjqiZpC+t4wugXGvs2JvmHKgDGzaiH
/HWRbVFQ4fJMpUR1X1IXScWK5WSleV2alJzsvPb2kZRuZt41ZIX10nLnLQTiG6Ll
7kkfxtNMv9J1YNmgJ7XeuB8yuNcc8XRf/m5qk/kcxzrDctkXDt4fUfRJa+1U3MVH
cMaOOD1VZ8k65rLcVpkP53B728RXoPR4ry9GhL0q8OgOVAXcCV95kNvH5ofK6fq7
yGFY2b5SKnltcKKdVJcNgTF9E5SYmLTmDpC3Z2x1dEGCvXGBnIQwe+RVpUCoKrbu
YNB9S573tcWgUaXST4cirBaebYrtcN6WI0iPmu9vws8tZ0AYE8tu5FTlUrCLWouE
vguHTlkxWZFVGjDBENI+7oFXY4rTgzVL996up5OwJ8TUX6kqOCVFfci1LipF9s5x
X50nFfYjNR629brqAGaHK3px7FxFqoP3QMRKLGDkbRQQR9FDCEpBXW1QgPu/aMvR
BiKu2ACCY+rPns+9a54Ki2gn+u3FzsN7VCl9jEXGDqn289D5MJu80Lx/QHDjuu4g
rN2ThejwT9FGxpos4pSzm7m8DJseTVfWAA2xl+JDbC9qVrEu4CJqW5XHQxOOO+Cy
Xyu0PgFwGivZdUdW2T3/oJcB6vNOqJ9g3QhDypzrw1vTmUDLdcLh9/3jnSG/SIFe
jTJIFZitmQfPeoCXDvvpodp3k/pMazs8sL/yyqHf5/AGr+p6eqQaksV/kCFc/eTJ
ke2TsG/a8mkKXOCql4AT1qoVSAJFWG36UGVINKShbEDvx6HDxsmh2hIQuPEOl5vW
fNcOHg4C7ip04LQDjjDki/cJnzigh0fKGrcIGIQ2HjKHdfhnR6290Z4fxES+vDHr
AIzqHVDpOjDR2GYrCOkiK/Thlfg7Py2sFGd27oU8ntKDwD5wzZ7dom5LgyYIlapu
XGePHqYwrsTaKoNGm+m69LeIm8Q5Ar/y4jXGqCLb4O6rcHGsG+Wp+xZ7m33PRqrp
9DyWRg9+xSlYHuPCOa/4GbYSqV2/Wnj3oTI62VG7iGZLTP7kvkEzWgNjsRF4ZoLA
KW4id7969swxXWFIjWlCla2qVZoXiWKphFEo4SrhCvIbumWPAP1xRD2veT0YNrKH
1G5hqkC0MnqyMU6PIdwvBR+qDx5l39YkFblbjJUG3iydbJBeVzEJzdWWhv8WE67p
lSAvt2vPpJqigSBCzVYlJ/G4TlYkYVbekZEjXq5b13kbv3ampxDQlo8jDJx2OxGP
BeFY1No82P1jWGDyPdcB0aT38TNv6ckDxNSQHesiHnRJA0RsozGc2yXEnT7jcY8N
YdMzxY6ksScgzu4eJRSt1vbrtnxQIi36De+AKNND2j8QmFGfJuORkC4zjpqc9k5u
cQhEVHp3Rw8iZ8QYOtk3r4unoRYwhf/tD5el+SLmmmpLjaBF5Ju1Tkga4ZMaineC
hlYWJjiqedN+ItYRIpb9fo2hwbiTenmWz1rIcVe4b36kzF7Eu5OMKOkhEnTZTyAd
lY7W6wi9uveVxbedTlRwuBqPdF5Nb3EHBC9lWcs53+UyLxqOfYgx81yiO9c4mZOd
dwOWnltR8/BKvlfzKzhPB+mcWYzbUjJ8cc+Jh/ir+Rg1SBA+V+vWKeV+6fY0SfZV
eppZ397rSgPy2UIAT5ReHy6gT58n+7p/RoqGtQO/W4GuXlZ1H72E3KiiwqUByrFg
CkZn8jhsBn5hI9Yz5Kf/q/myuw7BJyXkWasOmqV9wBavsiUpQNS0N6SmYfxruavV
M6SQZvUxhbJILMU3zkhDClRcCJV1L17l2AJgrZ3MKNpBS2ebcWIWDf8yiuvozOWS
3gnu6nIpO7NKrnQa64yPMNmp8JMh0USV7Aws7RtPzhiQVywH8tf3mGEhDu1cMUaS
q1nBT9FpC5aDB8cBUjbTH2HPpezdLoKUfEjwfro7WOR+uTwprCbnhv/DRGyeEEHz
PQXbWiNsAGihbpu522upAVYKxXbPkW/vlpgI/0IF9KGc82lcyZJAAYGHrhn3ZSHj
Smq5B8m53/ZvUom29KRaoyyyf+RUse56G4m9Gl2ckUZkGTERyHWEC5eAdhpqx7Mr
CCU3nGFx6hztI1iFxqgsnUxaiqG2t+ikzLAM6qCH4m1QW/CCEZeFzrcbBSWHTqo/
6ANCHnL58qaGX+s2IWW4rw3halOUDiDwwzgOuyBEGfE8UhbKzwRMqizkuhneUui2
o8wK+7XU/PT/hNDW0UXsUNIDyhEF77UNIXVhPoYUNVNQj8Mg5sqUj+tdS8kgsLAy
TKqBvOs7gUyXba3k9DUlsijJBU5KzftSrTJee35DGKugd1OJqsHAZL3oCjoND8fM
kNHCNMYnWxh4rvwU9Q8BP522bgtoQZ6HcCras5Y2b10/wv4n8iUPI2hfQQXl2bni
+agZbtWHMf5SiHqWKL0b9D988JPexfAOET7SI0ZBd/wu9AsinwOqF4fC3GOAw2uq
ljivMKhfptR1/5y1reaTQr1JvAGzKYZGl7Kj5U68PKUep+GzikGVFmEzuU0mNjBy
tg1ATNdz4H8r2DkjGHMMEXFK5iLBuNJTwnJWle0Y36791E6dp1A4uGurWLthBTSt
VNEaOHC4a+OGLSO60HLMOGlOmfDAmp/5lxJu3Oy4XJyn7SsYdPUT183NA1Ltwbbo
sAiZaZRRm5QQDCv1mu6I01RMt47JfyiltPGytPLK5oCzxbB8oPibtbwV/YjnKEmL
eBm+HOLaQ3mfzzAakLobNaOS5ElTw+WkL0XLawJcrL14A2G9lCwQFnzRTe2nGxmy
p8xfKjlXkNuJsljBGYhiZGJmaac8b5VrFM1qaQSYRFywgXIw7LilfeU5H03H+pHq
m6uQw+rtze2ziRZJ5omY6hTWaXEbEHAhfqcAhstHDsD9vzfIbUvCscgnSdQ5VuHs
kDqgI0K4jJ8evQAriZACUFfNY1A+W9WHLlbKen9XE3Alpu4mk9YHexiwgFeDMNwN
+CHjyTVSxVqjND1yPcZVJ2c48+glE1HyEG+h4NZxuIPCEFGH7UYWbjlzh2Jp6itz
03a2v/NmzoXn7JppGj63Lry77+nZBa4qlJsCyjDcNCIX/+qfpBvSSnrb6Fh9kJ7V
cMBoUr+aTRpkR7b+pJlE7xNiqe2t12Uv9y8FNc4DmWjP9oo1M4UJygEVplIW2LhY
G5wVKA/j0xukv55grpVcwr5HReLstPQikewzMh7Ix7v7A5duhZsnyvmfFtUDG5Oy
9CtSkTU0do+PZgospbDYGC9tGbpm4ffcb2WS8FCjidWN/zFtjFuHAXPMZZcLN5Rw
jJtfazZcpdeOFsxL9PjsujogV/QHfpnxR7RB4/UrYMhJM16McGW37MNbGETBfvv5
NwTi4fdZsebwmtfbZJNrlcW7PpmTn9ZUmNyExsKhHoIUPR3rzJSPOE7Z1LU0VONC
88ElJ+5cZYHtx/KWwqo5YMBCx/Kv4WAzoUS8fWV1SzLCCPYRHAz8NSz/llv8I+3r
GJC0rnxx8zhuVMZDXDsKhloHqmI7aPqolrxHks5hKQTRlZfvszdVgDtajropxijE
99Ws2nD1uRJzg5bOyG2rSlYF4vLVATIfrdVckJJpFv0qNuWb8WzSN87hyMmuIgwi
GnJMxiDPt1WtAsQdYBU3cA32bs37N0p0ePbadQ3cFeHZmutXZ3vsNhSmOmQbLPkV
rwrV/7qxa0rcZP4eQ+69nyItZ8KwgC5SZ/SugUr0zcoWYzRotHuT5RPJGse0YeJJ
Txunrgb4ZjzfUDkF9Pcmd3nJBEuHvfvcTV0BBGgWbzHRleDHoJvK7IwBleSXHTRF
zOmh8Xs7jgsbF9PtKUfXetI6fcXHhC/gtaLepsfaxzgrdOHugDT+wi4eJEUYknyw
yDDsEzmGrePr6zIiwEkJV62+cC1SfAKU05yFI9cMYvhVdTEgSTknZLk5AC3AnV0V
tVipX2+dSbZuySDPItZQkDzHX/+tYr19eJlh9ZVBAzRH3b3yKbaLvhwLCt7W59je
v//HKhHJg2Y5n7ctRa0wiEJCTlnYgOcCit44Wlf29+Vr3ckmzHzZFEZzdfEcCUYL
cbr3oGHKbuOo2TJJqmS9jS9lyhBgV3cBYgMbqbqSSF/dvQm4A+JRU1AKy+z5xtbk
CaJD9oVjHZMrs3ZRyaarq7bL8e0eLnk1P6KuHFiFJbex92QxAwrto6r2mSu9e5oS
Utrz0YQ/n0/E+WilIQUWxMu4MfkHzeal9rBITsMHHUHjVqiVKtXevIE4N7ZXY9Vz
UQ3RhRoiv7fh+AMI2UmeJGUdkSNWYFLWZos52ph3xZwUxdyQtT31d5ID7Wjs9rUV
AoBSlbAP3BwScHHh+nk5EedHcnAZUnqzdbTvqs0Bjf8xU+IRlnVPx5HKFHXSix63
ps33C4SJ6AmVun8t/3Jhj/Jj7DwA85o6x5R02k2pqVB8SMnXxHRWMyOg09Q0QjO9
6Z0HiWMJLYk5pCslp74gc0VIssN4oc1KAIwrrP9fvso8B+9ygq0TDQGI37tgQW8O
SMuCqWknuXEujWdmFheBOz+4tCnLC7iFe//YgGNk3W0JgT81M5eD99TjbDazXSs3
n6F0+y0uSKJ+ZeKYbbvhebT5+uEojn+ElD86/enidXloEBkkkMNDuWGAgn/QASAg
P/4wbnbW4eHCcWL9Z2Do7WuWDvzv2AtOW8UEWkV4GBMqEpW7FYJFTsGFtAB34OaX
JRuOnwA+sly8OQL3XCdu9k/1dBXg/RqZK6yhfcN/efs9r8qB5snF6gV20X8QawQ7
OVlZtpu1kvpxtwpSVoKVnspDPI2TvW8MMNl8uXR/cQG0k0hISRzqmVCIOiXRQybB
3/avDBI+4PjoIX0I+Wf2R62k9MgrNisTCuv2OxLli0+CzNCS6zln/Oyp2rjjLq18
zX8dYkYd6tBSnox1NiwTfKZlQncmiDmaR05VO82x2d6YrddNM7k0nraOq/IoZEKk
kah6TxJ2JsvIJbSzidpmX2dO/KMMkK+WYWlwqF4booPA1yJhxuIdwQ0RDCO+p5y+
a/Gg4oVEBh2GB5A0BsEtfwTWqxxW9yYysOO5SCZySWFdTJR2b3LJMM/tc64VMBv+
07/VNNMFB3cuicy1Xulkq1pTUMYTUvl51n4K2DJ7SDGI5ekjiJGmBoMOEZQHLPUT
fIVVzoriIPWjWSiOegbudDG4PsEPM91adqp9tvvPdBGL6sew4zWaMByMZnEPTtDb
gAwILBJFtC5X9Ok4/BpJG0OuaBKSsa+s3lCMauzB3J/c+OVMFKDI5V1q/NAgXzxW
Pc7bUe/3Fz5wJg+ZUSEwh21+tqk66hAMuw/tD0aa6GXpLiAL/kTU3kcyBS/zY6al
zQfl8aDsEz2r/QZAzdPEr3twq0dUOqt5QxAfnKcWPfkDr2mfIeqF+C4QN+7POl1c
mPs9C9ZrPYpqke3pascP2S65odt2Y+0RavRt/76aBieGIkkYAL5a+5VhkN/9KEGk
jnPF8pqtAVjC8fH+rDjPbQmAQiFjIfPDI11i6TaOWFAMDu5NE9O6qe9rOfdiFmiW
RdnvY7KQjo3I4t2NV1LRJdktyYxIPGOds40vRXkqgf+0grJ+pAiultudl+zPEnAt
ChmwSHUbzTJdaDYY1ngguW2lt/Gh9t0izoFbZQVrylBoJ5MNG3W7rO0Bdqyu8yj2
0qrEmBfHaedkLKOT4v2TRtlSP+qjy1X4gSGzqqCCWL9GEKOZnuM7DKAMTtm01MdG
Dz9vBtZ4V1akVMC3kDC6eGCVwhGNejA4oUy3ZgvtbfnTT8Jl0m1iJHoKtxhDAakI
22stAd3l5PXL2bRhKMFOc5Ot7xFIXzdG63oJz0dsLH12PO42LNtNJkgI6AKbiGOS
4Q2Yx5eClsNIQi6X5glU9sJBsofYXDb3u/XGi0pXvcG3RU+GWKB5qOM3xZ+G1csJ
XuaPG1xD8vs5FBVb6VarfpfXgSB3HZLMgxr4qZgB2QExVLvq24ORYbS5zE8v67oW
HCLsDmhBNI/Qu9cQxQm4HIM4BV3xu+waZTpLr07u2gLDVBeMrwEaz4PNwsAE6ykn
g30iSs7Ji8fXAThhlYbVV390C270mmKgsQWwOZEU0N24RShyCRQQGtvQ+ce113Ah
pp9GcGH+a3pk8RYUH/Szhcm0nEUSII8XPzeBdwSLqDsG2/KN4sJhCS9eH4JQLISR
MiILIYvD5Vr4vDKrcKGpddxn7Hjz/7IxlJUCdM2bsk7kiHwe9l8gu2Q8VglWJERh
UUDi8eBgtOmyDBjzTWVOBVsaSRRuzc3LlV8rtSa4iWUoHW6WnEC0GRO+tAPFyVwz
sPJ1Px/jQYx2NFun32gxpw+iorc7CYuyuH5UysUM0pPz7gTL4toeR5Si5suCDc4d
1V6/w0vpXa6dF2Ax73mHX9CSb4ntZUYiIZfb76K+6ZRS0t+rWFy7zx5aNs11PHEm
7JNh4PcFXrsnRA9Ygp3nmzYFK0OghdVTl+HDc8BYqE3SjrfJqCbW4na1WF1gfikx
cViMbSt0vIMSdGU/3VWhooZsTcR5j1T5wZzyp7qB9Fp8YdX9SFCh2/hXKPYuTpvY
9462TXxMPntE7yv/qjBcmDyHzyciqxLnzvfy6r5eEud0cLNJSvCh5X9YBIWdTsfT
WGHAug6+V81VkQqVgbeg7LWWEON7nZ1jrzE0WZMolG7tZwJH2QbAWe+nOYbbFW5k
FHWv0VNxXWH4ri5ImMr5xh0MB6W0yCw7XWze23zJgQ7gxqu6K4a4K2T/lysam8HH
VRX3S8VS4n7a/MqoUioAX4EdBXQk7ZuuGa663S7VjqliU1jomH9DuZ6v9c2iip8w
K4FxUXHj06ggwG96Z46sYLZWXFd3pN6ts5IWWmbMUspsIrbNbPkrgmRGXAnvAWS7
ZpBVZoFyrhMMQbD7Z7lPgQ+aKgfFTLhQemvd1R2n8a8uE8eCT+qbScQ5H7C/MtB1
jweWpksi/dJHpz6nlhPkY9aFVMGQwuNPMesUHFxAAKplikdoiEmli5gQAGgS0vX/
5xo8bMM+Zan99eaq032Cp8+5wRt4f0ZTVih5wRbQegdKdNbwf6Ec41BlKaLPnqMZ
Ln7YreqdRsU6G0oLrIDn5MYVX4DgucYwRC1aOdGMg9cg4g4BP2vezHyPbRqckQfs
l9HUCSfa9gkEkj5LuFX/F4Vn26Lh4qsSb1u7i+Z+djSHaquLknff5jFybIv0P3Q3
Rdm5EYkmZ1kx1L/3JDKIVpdH8teF6JRwd2+35CV451TRfn9ufHnbB0WPGzTs9J7k
7eXUSaD7xqYTysjD5emlvhla70sPhA6ubqQsoEafpRj+1Cu5Q7tXSi+A0wCX86FP
T/Gbl0rJYgz0SV19WLOIrQwgi7sMLLiobND6CyzYTidSyZQ3G/Op9wxa+EcFBl5z
HY6KlNEhWGi7Xn9KHDXz5ik3DHClEW4gqq1iHauNk1sUfzofEYnD2NMxhcdpRFG8
yaNI+v0ihsBq3uQUcipR2TFpQle1GMrIm3uiXNaoVbA99ExYXjPTqP1mqtjpZ+eJ
dNqwWr5aLrUv5SteboW73ZUBDtk0OM946caSnn+/rQ2xnFtDp2PrSxEbknVpnDpl
1X63If4ucuPuZGiA8iMtKj2VzhBk0EqYaRS+HxmVUBGrobptEznJ+HUMZBtaUFs7
TIxgUXL2bwzeUrSO014082D7UfBMl9jTkFv70qeCIPpF3sDyqbBESFjLwdXikVNm
jIVQH9AQvA0VdZz8q92KsdM2pCNk4Vcbb29woghHR/KG+HQBZM9bj5jD0Dsyww6V
+BRSSPGQ/MEiAOwKcYpeNjZUIebPa1EGIAGjKnky25XPD1uBtwlHoxFnOprF49Gw
DVkf40lmvzBmcgI8ZHnleVm3lwepTBPl/ILey2BJvgkkO0q99UcfxuLoIfLvCZP5
cbgGKMFLPurUG0ATechCvrH/uq1yhjfv9I4hrSuFqTcgSobWWZCer6U7mSlKwiZF
aijP52wKRHfZRliFge1QM6KpVb8zNAc7oMRQ/FCv9UtfNsmYjJE65g5JZUweDEIH
jN01ahlQEHfKzjbjQsGYbPq04gys2I0ij5j4Q8klQYOTlfgGsiBnmq6GQeRS5CJR
c+JZZ1UR2uJp5rS8JLNPJQYayEH0VUbEb5U9V/dtxuapKShWgaqjgabbHE8VYQm1
QHwPW8L2gCJIlXPGcWMcq0FYVJF0vzXGSfb/oSHhWIogInk3X4AadliZhcGrf2Bx
lwT3JYKigQFNfR5ZRLCyDKalFkYCyBfq0rj4BJkM5UBQHCudoSnERIgtck84U//Z
vErpMuft0/C29IG636ALTdRwAAKob1g34jaJvEBSoaHZYWtC4yZkwTdfxwPv54kq
VPmt6WLHkr2Ss0GPpgN2dUxI8OOnDxAZ2Qnid0ObDtyQVK/XmUsACSXVF2AzeezC
htRDmxHpmk+d386Wi5MK7nVSz4i3VUhPJc1eZ0ouDavJr4IDLn609zk8edBC2vYk
qdkcCQU1kicOlVTbduNu0ug2CcsfBgizM4RkgN973QD0nFn2HyhUxg27riQCqsNs
wp5GxNwdPDHVrir0At8pSuyk9gX9LFdejUB8pyXnp+WZxMlr/PjsAZTyYnBzO0Oa
pQ5+oY5C+KhUS2F2ckDuLQQzzBEeC5Hk1B9MJ9UlGGBUFu6tzzmBfu4UqC9ERMuh
cXY4dWEDu5y9b/I5AG1zRuIyohyVJwnCjDc7fkc+xomABIUcD93v/0ChM1sykmPM
pC4oz65oPdFBQqEWVMz51TJDtWClPrjBRGNFtUl0aZmINuCuY0lBfci3bW6WbVOr
zSFmxeyxyNQS7jZPCRzWoSvG7xfisn1CjAjcfsMF+cDSbCM0WWbZMxTarAVLf1Tb
l6iUR129TqpVCCO9h1C+IMtlSOBbTJiI0tPQseoQomIDFd4vYMJosSMBMiJLCiZK
0wihBZlcncxF8JMgxp6DPUX0+vABx+s7D9bnUwoIW13iNUzakQQrnoul5zWZA4H4
JwVydI7D8NlWHwBtCPoTD9Yu2qkXMUaifPVGizyYHaLqlJcNczzVhLFWxpRTSeMA
CGYvKtlAe+BmLtz8oM/07SZeP8ZTGYlERTHEtJasEqzK1VmS0u0N62QpPjaIOp5T
YxteFbMscYx5zVrDa++rASKUa67p8IEGE1i17SOla13mJJRYLFJOsj6j4IgnuHuh
vSo+RoFM9d/gwpvxoVr/A0XK3cIsbQbXwpZfo7dPGjM09uDgowHwD2TxnSNr5fo0
caxwxyQRqEA5wLEk4o00wgn/k88+F6+lcGqtbI12PWaM4BG3E9R4h2JyegtaC92L
zGC0Bm1IElRob34ZKvsVBZ99M7iISDDNjqC4bad5ccC0pg+Fpy01staUZbGdesxJ
rlebyBDxZCm8RlaLg9WkBp3w1PKRHH+HDQ7Juth9nwD2TCJ46ZNgFzqMzI2tk0fp
r3Aifk+t+jv2AZ959DuagrwfunmwQkXLQyXlKO8ZlJ9sRQgw/OeyVZ1quNYywp2F
QSTSPba9Hu1G9dgqC1NDSE0CGzCQz9gDpA99X4jHdRuXdNr+e+GL0E+FKA2ZADDA
NyDa0hhs3Cxuipsqu6UqnBmBrWzzD7U0oUE7K7viHe90sqGcmufbVzjyXQyavMY2
uzU07SueC5T7xHCl0u4A5biHhcHb7fBZsyVYFac2jRavqPVamONuZaSf4iG6CUGT
MZCTvQKQ8FzKGxZMsWyiPvyM2S9pt2hhBXnm4YVKqql4tbaYPoyOGfzhO1Ht6SPc
KsS7glL3qmFgE4CZOb2zn7WifSdDJLBlg7AkKHGbe6i6ahqf/oUGpMDrr8obZCWq
q2SNAcL3Meaki+e7WKP3slflZT63F8k6nhpCyun69FMWbnfSSt7SArQwBYR2kHs0
2ZQ8kzKrxsTdXpb+abC80ADM21thiuGGeTwzxnDuqFu+l/UdCtGbjwHnAn0x8sh6
LzOKAj+Uvpc75PPvB1GZfyq7GjaEptEXTWD8F0cHdwDd0gV3zrnufgepFz8OetMW
FdEzJoLyCBy1cQLZBR/A+MdeJ7iqiy6xJ8ECi0RzQB+Q6xgMD5+Q9rEkp7tM9ooq
3B2uRFWkaI3/+euTJh9ksVIZmv6xM0WvrJ5E41W5tgkeS7X6MOMJAkcX/hUagTwE
tkz+RFoEoKdeVUU4ah5kjI90LrW7mFXxPM3YXuKdMvTT6qhUP8am+J33zKtq00wk
IGAl1P1w/i09pI3+q43fPGJ0bDPPoZE6SDMYgYKfDoOrBUH2azV/8bVQGZOCNApg
FKHE0No9MGsR6CKVMsCSGvNdo88W1vM/jgM6grrpUq6c4UdBvJjXxbA8mqg1+Bv+
XC4/+Nh4/gTFbIPnVqqoHKsgKav8H0o/PI3F2fQCwbg/Btp+Wq0DTk1aEeMU1oVd
gMzhF6dGe71+3M1wtbsnF6olDsOoyZdmFocIYbQr3VzT66V17ySCvnAe8meDFiXG
X2RSWN85xo5DYGy4KxrhTkvToNaytV6IxKQcLMNf0iwZ6IMKWz/KVROUWXMIp4wC
/ODW3acNfApkvrlQipF8slXQ5UgnImwvLfubbSTZh+tGLssj4r773pnilUKplb84
l/an4puPCHR31N1O/BIiqS6mqRwVKxVT6mobkuU6M8av21+ZalsemmBI+JalnY1i
PvS4+VYf9bSvf1QPpKR7eaJYB8sJCyECwk348nc5hTcjH+Jo5JnHrAJfyi7Y/m+z
PLOkSq1sZbkxDKUT38690gbL0nrZE7r6kMMgQkU4rusKNoIHk1eLjnxIl954ZVHW
/c9LNUbrV1y/lsx/ntPKG/UE5bLZbvNF117Npofy095bVYX2u+nWB2RANEs6Ccr/
mG+JkuQA+Ll4pR5l9LzuVfKbuAz0QmPZgJPbtUFYc1oiVFBx/50bcCP3L35A+YhH
gpkKS0rtahlJn5Qz3Rm79edkGnnuuekyCyAtqS5XHLWXwaYXqmcgC+euWQt/Luzi
NypzEC9qegPC20iZUTvQxnCPUJTw1OYSjp3Dhe4QuKnReeZbaHzYlOY/nDGs0KGA
r8Xqc3U3tib18dm6kJE5SPx8ckJ+hOI2rPrzIFGx/oS5DqSkERPWgFuZr3ilevJh
VSJsS9NvfkXgOzhgc7Qj194KmBoaqSdHGrZxM8fv1XCEOk3V85mM/mamJmcukbWN
ud7VWrcIfr9uV5ktFQGAVxU2hCaBzBtzEUIaLJ8bGP/1zyBLFTN7s0kBPrifWTOi
1+a3IkWgrfxZmS+UEhiYOJbE8lnvFVhR4U2AvEYwpNvGyiFPM3gsfV7R2BuCVbQT
Nnl6JPyefFafebkgXm54W6+iunkgvOdeFkI4vCXtie5bKEbEG38FLJBu8xt6sQOh
VGD4Paq7AvWJtE9/ItRcPtGd/hbgWHJEDHd4tqi2SGzxRcEZvUSLnMhAC3/80YdS
cYsDIFGnLCvtqSXHFZD91+V8+pyiJCYxsAc7tJYGegibqzf2/25BMPJiLXTFi6nG
iwKGcqlzAftfhDPs1ehaZ3bT6JTGG/kOCFyvyjAP7eSBgPhjRE3B4WDPAlgN0DIG
KWk72In3vu4wMJOpo1vbWYNqemO6R2cMh2O2ydACXMOsss1DbYKUNqO0rrwBQdvS
NrtjCX1AfGHJG52qa2J64GBYZ9hDu39SYKjxbVv+XFdO2J0A1YfDSr0LJTdNUqXc
vKQS8xNNE8ep4r8vwfoOMEDt6GtaOFVpB0WLTYkFUmJqtT30vYlPg7q4RtdM7H/f
BmeK1PhlqgziMD4oqnW0G5OEovDZio1ilP094HHhx7bhS/MpmW4WWV42j9/Fp/lk
GTYctby0YDpJPv0diX+M+5SCEPKUdfOw9f0UYwrvLCGnFv2+SxfAm+WvM0zd6gZN
KMfOB4aqHcD2KgL39ac2iFBd+GoM59XaKVQx6eir9F64LpPX08ordhQQDnKES9T4
Uh1RAaegha9daif4kOYK0vOq65aSccSgJdc5dUBz8FhAcOQEA9MZFx6U+K6bqusK
ytJMkJl/yStKzwx0HMtdwjillbvfSVrLIfiKzhvPPXyk4faU53GflFwGV+l97OBz
LiqAzFBb0N1elpG7P7t3ggL91v3djs6zAwCJuWbEj2Hh7lUa784YaASaoB8ixwS9
iEWsF+DNgovOC02X5fEsm4uEeU1Osmr+EMySpZnAOjbU7PK/HDWKKz6NK7oV2uzN
OvulZXnXBzBF2bkBDmeAFw1w+E7C948iJKj0ixteugJRh8A0Aq3F+5eqoDC40SA2
nGa6jEWCKqFgvLAIYk2SElN0jIC4yrTBygrZxnotVxptK2dzhyXvmia2RxQJWe3h
KtBPoblmy2UK/Q25AHXt8Q9DwKp3/3+5Y1W4vGjhYJlpWbUGa3G1Q42cm4Jeo7q3
IgaaKZZ43f+HGeOjnPLwRwvFzw11LILj8h6/Xxp9EqPL6H0D7xCrldox1dEaOADt
bdxDw2TxFhGNWnDD3Qctx5SwzQi/2nGc9qeBu4uNqoai/joGtTMSC8+ZcHEpUgOQ
cGmjAL7LQ8M20bpSeac5lDQ2fXJcBsO613xhVid5MXFcY4XbwFIrqB/u0UHYH7SJ
j90dMVEXKNqkwiLcP/uLZVxoCXzvJYLX8Rk3t+x/45HlznA2RAt0FBjpE/ifczDd
I7ZpqggNp6lJeJjJSi7qK489tqa8ACX0BW1kUmil5SvsdG/cXkBo9XT87w6UHWBc
W/P1LiiPv0qF1lEeIL+0lRhJKT3O77/3H68IM1d+V3nKZkNjt+4gCxPyrJwpxvXY
6FzwQ3v0f2TRi8S2xSMKgDdcB6JAV1Aa2CjDENzxhB8RCSY4LJwHvsqswGeOh34+
evYZTQHhjXSzGZkIQxcaummd3DFpYMRqT2laC4V8AJmeAupP9LLbnmja2jVvI0Nt
tH+h6C7pqAzWggvKD+Kl8WgvTlp+rZIlAoOgSodc0wXh9posBSkZcnaGF1ZvgWjs
fk2wynHES+MBZ66Nvaj9j14fWTQzVaw4Xaw1M9j6AWrEBbXYdQTkCC51v0Oel4w3
nqPagz/NCTUfFnXd92nZHytZY/bZu2Dop2lV587ElgLMyMjyiu4Bf3jP6IkWC/TS
PFWkf0Nj/2uwsxoHDFriFTnohnF00PKkFYdulq/B09NElcLR8kQTjLBqPckjzOlL
P8mHLJfiIO9c4YRuUdh0wotQzlm/YErqnY2UKNtBwrywwo0+hgHPH2znU91ZSDeM
8NVV80HeXn2plx1W3M3BdBQ64Jcaejfhv11j/RMs5Usw/kpPDAfWRMccUI+wbcL4
yGEQyw1MLMjJJTLn9WVoKjG47q/txAb87Eg1NkoPpV6K1uhZeF+KYmISWbsZGFed
UGleTb7uN2vNICSYA/odXqqp1dtln/jEAOOex+SNPfXNeAiNuYGitcA7Z/g8O/sX
Zay8PcO6zky9PzqFoeHaMWbUvCG/zcClyqJpil0VkO3fzJoFUv/rkk7cVMYOJFHB
wjkXMee0MNfRVMCwNPnQ8gRryZS8IF8sUzyPrhBR//8U7WUSKZn75yW+GZfrbKn6
jc2qef6W9ofpyQ3daxeFhNLfi6pjyPZ2CqC2gHzgSUXlKNKdmWGjx0rdEiNTJRH9
aZNCHbI1Jc46ekAmCW2QDtWeLcHRN9m03l4hRLE6NtHQ8sPbrZtyNvuPckGrXHVb
5Ygqtn3jna9Sp306sg8/CumYYHv+HCzm7dvpYFK5TJ/Cg9Qese2jNTns6T88TM45
/k2ZJiZebiGS9RJhqTgTVdzbi3OfRcBOWPFVLL33l+Qlz4w/bhXB3x1af7O/HYLU
/CouDOJNBFsnWkhLvcrXAD6pNe9MIE7sVcSuzMm7Celm2/qzw5aHgulUrkjdCRFK
tyVAoxVbU3x2xaz55IKVRzywTTgDSpmUwpgnR/10He/EjydIx4fnpcc859IZzwt3
WjHRQWBnQcQZaxus6QSLpNRbYQmzDF74uYZN7LwhQDZXT+ZVon2wNSbAhX1veUZH
KhwZgOllBG0mOpwZ6CxjgYESCNTba1vHsTor4B9jc0wvXUWrgPsx5xw+gPkCqAlt
sV1LQnUpF6tS6VZqST86YNA8jSnkhxX+dmmgbMqOl+RHMuQDWo8lfk227Bvl5Xs+
L1XW5TiWHS9IwBcoXi5wbqTGCkvykn9tKh/hj22Uoa7OR/cwT8qL9e4VvlfG0AHW
eMk+6TQ/Y5uIJRRsPfc0/fd8CzZQ1oVMaFsndDh6NzKyfqbdE6RkPyGPHEd9eTrP
Cg7PtHAgMt6c4CTx3mwxHFAWTMBjVx1xRUBkNVZMJ+UBLiGoVp7J+xOWpJmMG926
qwI4CWDufOI3FdwC6OJP2YCAbUkNtpq7BbClAO4NuwRIBhNY9tTa0iGOrgpiqOwm
k7z0FveCHtWBv4LcFkYXbaMgEJ2U14WVOcNnb7IYI0b2oHFUtNDAarGtexJgWdxP
7GtqWIxOfZtbhXY2sUmtrgbLd+fkGh2bPW/qXxMFdvIYqIZV/f0UR79m08G8Ik78
h0symf9eNtr2RJ1r1+RKpycHs1Gkfs+Hnu1p13JK/x3ztG4kKg23pEIiyDvw+zYn
nCnX8cHIeq0RIcNbx0hykgXHUlCkgHhiedERKOCD4Bud43eL4om3i1iuNbi2uojc
5+fx6qRYI1kuijTR1AgGwO0C4SDI8tHLdtzwwdGvvoPlN07lR7iDwnmWN6p6rAMh
itLpa7uBmxr2z73Pfcr6PVTga1hEEb04R0TZ4cxs5QHa+fyTSt6F64zvZVdcIq94
gJ2EVhk5PpqLj9BHU/ys4Rq7ktcqzmQHKLYaCi7DoyTa3p6Jn8gOe7euQCUO4/pA
+aE03LYyV8JaWppJzhePZbO7LHPijHtXwK9rsfEQXBadYV0pG/43TFAOZoeNuY+T
vD+T5AMsSREiYzxPSjylC/rSjFu6MM3oeCaWXSLVwbwtj25xiJAgEd12tglqG/We
7kejf4XFDT64yo8S4mJCJVjjlfY87uBNq9VG+QHi87zyES+Cj/zyQS0W5Evu6arp
wPx2uMYcMqmVv6KZgggcwNtM+fcJ5evyORdlvemkazinhiYq7M24IFOrJpzgfZH2
AmpONkkR9I5XWlXOs5v+wcszGz2yI5ms6EGrwCRQaW8cdlSHFvRwS9qTUZ0+r2JX
TlnF6DjnoNY8CGWTGTZRUjION6MKwS34mLc+EqU25jmyUwJzt1cBUrP76j9TYJ2d
wSugFSA2wVYw/VnbpjHefCz8qr7oRw7BpbXa7HJX3sLIZYaSAlHvjE4vdo+H3JXw
sEb2qoOGRQvW5BRDfplUZ6Kaw8SXiZLOjeY0TNxDGZVQCDF1oIuO2ShpjBy5ZwvI
Kcj2sc3rOZE2CvXE7uOZeCOeWzS3zwTIzqdiJ+p6nYPmQs3As3xjutwr8bjUYiwO
j0oSSuGryGNC8mZUq22N8LWvofgNwX91S1eqjYjPvzYxbli5Z/dg7gJhz2LI2Okz
J8te8mmvnT/hB4pueF4dj+qMgtQjJylxnvNSIgeANWeCpmM5YNoIpQ0m8Dc96KgS
wwT9nYIwr/NMKzMxjA1Ph2Py09MOH1kwitBiA+VT3iShy941pGyx2whtEEYjZJuk
wnP1U3YzjdLo/CVTD0Saevy71NBiLOHztWoiaSq8cvDHUy4UNN/je6Ex/PZg0HGJ
FScf81FhSUokjQ+DpzFt2pwwhB5pQZ94URT7EpUFy1RnOxNXb+S8WFXGm9pbRS5s
WIXrIxuKhIPN8sjEGLhfx9dNTyRURoFGzf5TeQT2JeNHoTm/JRxTt3mW4d60FInH
QbzL2xXg/fUcEXkYc8B2jc5c0RUxoFtQDPTvIfrlLBZbE/XrNc/g+9lllmbTcd5y
JZYLB+ZmpUe2GyGSHkArAh5RZha6zzxYJASgETsP1cVRSAyrTVnTvY+hxxB5QA0k
rVAViR3UrNhtqCfKbPN4X1cTdIOWWrYFrZeomtOfBSXd/oIndt7Ol412GNPYALw2
/Wksxumaw/UlVnMESilNedyznPXWlay3gFS4y7MsVzhUbzySIRh60o5wMo4kwtXK
oU0BwJYjFKaUeMok0BS2bUyGOTAyYp6HMUTr/54ej3cmnOLn3A+lRaZh1c/68GjD
qZVpihsU8OunFhPxWVVHE7+6n44JlS6Qv3o3krPoPoL/1SVa1Xrlu2HLLfdcSztQ
J8Q/zcTdNqDHqobGfQW/vmseqC6DPwk7tHP7rdkLWVqIUdVEIZpgj8AL8DqapaGY
joXROoi217EXs4mDZiA3mVzCht/72tqNHNVdLdMAYbXnraGU4ghX1HYVBUM0ujRe
GKnEV01niAkUkIpMDvq7Fm3pvPDA/kdaTJVoLnnbTHqoIp/5k0XmHb6dB30d0FXi
lZNwkGQuxDtnXIgCS+5Ba5dqBlvZbka896HSOhclPifT28qIhsf9BT+ih1qZPpAb
QdyJbs/DxhzLLh3BdFPSDSL8CP4h5Y6/1PSrxHvUuRImsAKnRin6vEs9oB7EVjcI
1NjtnNPST+E58gpoxwCGrHlvyEA1FSBri0kc+jzzJUWNfKmT0GzXqMjuYnPEWgIo
KB7TcmChXnUJzN1ig6TvI+FW/qwk/8lE4tBlRooN04tafPWEurzjp3IQQffTNoCF
3XHtXitDpB+A77jy2QFCz4Hwu3yFC484ZmG9xIKxWsMQD85fcf/LLB/x09rg1VuD
VSSlMFvmsQ6aDX/PJbzSiRr3/wPmoQYMzs/1A/TALuU9uhrnooghUs4WIP+XHQrR
O5xyOWhyFc7K/tlLmY2fuYeyKd2mbIeooyG786g/mgwH70tzYSXDMEtrG+Xnb0ce
+x+WMuV/ac2W3rUxp0ztuIud5AmsEcNfwq5nNgYw2VbKeOi1UIwlSscSI4jGVFN2
2FgluHPOEpyiDjFl5npyWCLo7Dv9siH2NGo7j/d4qg5I7jop+XH86jw/5G1hDMp+
hVpw1/dC7tidxWDBme547yCuoXU0WIvGG9qV3qD0v7cOOK/cYB4SC6udkVNr6df6
m9z5AE0gI1LRIL5jS6NC/qZQq1c/gNExgyuAswvy1q1AIfs0dNyomzXmBMQ4ZzPW
kB3Lr1nbQZho4jDsVNE1uEwue0rFI1tsjMbR5otJd4F5sF+xr1NJe8JxqsK9KYPL
2MjUpI+QkcXTZuLtLWB46yIKnfWfnjhsSN4riuCq1z8GXXXltzXTZSkbDwzoeKJZ
dBviTTWPCC2ZoK1o3LvkPnmGVov7ZSgglK61N3bwfqH/hnyv3FJkIfOTzpOqoAkm
dXg/VLb8CVxirLwzPEs5Gz5ZgEszBhETbfJ8Bt9zuDVqSb+07JIhXb9kpoKo132C
A3br+M9qsg8AE0bCzpZOy71P5uHaO866EdFbp0M7wmSy34iJQ8pzFungwq32u0ou
e/U3CLGkNbqcDzR71pGSMUMiuwvih1eYf1ZAXgRYM8d2G1Yz4w6G7FXKRmhWQeX9
EPTAe42so2P9TQkyFN85V9yrVMvoYzQZotoGuVUNh+Xl7euGDnLPL/5PXT+Vmw8j
mtN6ZotIC81HLcVvDLy4y1+K2ebyJtPeUow5Bz/7c84vES3soiBN/ly+pGWA/6tJ
b3ab8rls8Q5YUfMUxFU7IQSpP2oDp8/OnRpWLXH4Hyt1eVirJWjbpE4/U8Kzu8XO
foHSQ/vgVk4e+sNdbQwjmRXu8f101WeBDmELQbuvBn+3YPDyt0qlxv5D3En+4oi5
bDQLw8zp+NZ9sqgtEecAZJkShgEZcJ7F4Nlc47OAgH/oH7dr5pPNB75/E4zkN30a
reViURQjSzytsQM4ZFQJfuCh4p7CYnb8/WnQtuoIxrCcGioSldE7O/UmVNB71EJ0
kRVAX19VYB4NFgBDGwysOKRdm2DUqTA6fwPoDyq74TgFpmlL4eMngTbCTANEN0eK
cQ7aFx0bq/R1DaofojvZDwaV+eYOe6pncz4Bg1AxWmABo4RVtlEzEBVG52wHIo7f
5sPodl5gIOllFPcdOhRq2i+UUTqmAAkz0aqAL69ttUQ0+ozBgbl1HjCadyXMzVd6
P1ObvBRxau7BaNwJfiVS4nfXv919dX933PTa8Dc5ukMV6FbKgw4EwHvnh98lU6SM
pQl7xJCLpbLaFMI7Kb9VLB9C9y+4KYXDoqMT0GrRwj1vnct6rMwnhkytX4VSFDAQ
Jgu0c9+5LrFZ6GsS3v/eCV5DIsccXFNyR3gfluhhxc8bOs6tNfMPS75TsJbGZl/4
I2XZCpelUkAfkwdCjvdPHZnOTabowxOZG2Q1Tp3lf1YjziZhR1WYJGhZTOWkCTw9
8RG6eEf7wcTeqpySk1Pawxn0ksJFQgvr8q24FYt2bnlXRmpIF3KJn4ZquW+HprJD
s1h00uSxdqoN+c/MNU+pu3L02wiLy/x4FPfl7yvlLjcXBxWqBe0nOPBg+cEvoCCK
O2nhFF7e5Y4dqgidiUemCCmdZwQWf4x5+qqGVN/oJFeMcwfa3Xf4iAslsrgYRT6o
seAhA6iaaQykMoJm1G02Q39aOFx1fQzOiB10rL2+CWOqeZ4NjgC7qvwmFhGGHCyd
6DV2jSXqOrdF+jPGC/O14zWf1VThSmiPjUSAGdn21PXtGkPXzVbMw+3mR8vXoOrT
vhFIg2LC8A2c5bJQBn/rGU42DIpiz60rPlI6Ci194ZJm5d5P1we4SZYYRKFzzWsX
lO9jqG+KKGgA4jcRFTxicPPfCfJlLhJ3MnneiPyNJALco1sMImoYQRtDEcrp9YDq
RXafsUiwFD9Twe/iwKcvn6k9e1j14k6BMsrPe7HRYPyoXl5nx+P32FSRx0WLk7sx
bzrKBMNEuWW8UM//bC38TsVWSEiqghsu+YI2stblKrlN/O0DtYGoDMMQ/V1kNdtg
mzn5GOmQA4EMoeYnCKwUwpM3mwHamZr/8AMhEDjLVqO5jHwusfv/m/v6MMLGziUQ
h1ErwvxksLVcGcNslN5t2eue9ByGDLBeI4j0WWqqAYrA700RZUWAfa8sT134X/1Q
AWtpOHrGDB+tjMYbrhmVmkuVht6RoFQX8BG8wAJyzQ9Tlnl6PZLcbG4p6KrFp6gw
V82GnBd+fqlEMJO8de8Jx+cRcgsnzMno2p1bvxgSBMj5G9p1xIPq+lKHcafNH0Nf
V/77MplLx8kCcIdXFiUGM31nAMyLYakxLVHIMh7OGyBTYG3CeFubszt/pPm8Rj+u
b560foYzWSmq5Qe9Nc8P6zr9KCR2Y7ejPaFMLduPJMYbHgob30oe6if9U9tRqskA
9mshDdP+7yaY5rcHQm9BUjevmykY4lEG3SsPRLQHimkknPKhVvs83x5BV3C+M8Gx
jQeZNajxcPozzGmG7zr01tBc6DDcNgGin0eUL4Nd35OC3rqXnrZz5Tr3QcNGgCTD
mBvo0Du54ac8LxvB0UFn/1P1QXmZ0EbN4ysJkMimhf3Y6kq9DRA6GYT4zfHFn3rv
gr7fSRhDvCA0GmTAFvZmd/EZHiXvcNRnBmJxMsH2zO8KJf6szo7hQxd2ZdjUQ6vW
Ek6myXu5GubB3VPX/7eNgx4Erh+hWN2WF6zesv5tto6GsgSmOUuTnvqT5s7zJcyk
jiez+KFNrk02/u0FgOP9C/bpDBHk7+hLOKrvYCn1e0XvdXD3Q0swRPMAWxO8pJkJ
f6Gvjni9Zftw1pIWjaufx/UxQxx/rjTb4cKy63Mlpsnj+sqliuiatREG7CsHkoFH
VM4UUsjaY9lObmsTFZ/EVv1N4ae1o6x2ixgwwiEuc1fLAsgcjeDfKvVMNEaU3w3C
eh0FzHQthfblwO/y5/AWwq3I7MrHbcsp+/eXxPTa3zE3zvXK69gJMuWCyclyY0aC
ICdMLxqc2WODzXaYsDqmvwhJ5S5ptn7UT3jpNQo5IHrhVQxb7qk7qGAvmlE8ZQ/i
6nNmYtf2SHmTeZ+2DyeZ6OsJpm1chNVI2QiTW4tJtqNey4I440MKi9VJXu8hwP+T
bi6HMzAA7Hhiyg82ONdyeMY0OVdqf3O+2SJJK/xcm26Of18Ds7stU4AZ/yGisl/c
1liMpIVEXpJEOp3aIYjdGzHMSWtfe5OgmRhfaezPKAi/zVaFOJUBQyza22cdVEmT
Rh5Ya2U244pEJr/TbHCWrB1FlPwNaVNljDdCG+vLRVJuGhmXoM3DA6r/Y6lCXIha
Dx1qMUMWPP9rSTbrSFj/sOl22nEcL0vLRhllP+WgK9KF1iQg3tTpc4RGjFD/dC7H
HONKA1s6xqX/yqdJsr0snQBb9tM+aff0MqvJS71hmb4haer/b9TFaqSvF3ZA8uRF
quG0bI+FAWkH0W0cYzfPPEAk72noFjfbPiSlB9p/zbVBH+coAD0riYrx3rtlFqig
3DcALfK+nUg2RiobrJcSu3xUWBTfxkMrotKvJn5p4j/vdJjMZEoACuJf/Gi99H5y
3qTXEZH1zXkbXPL4SnC0SYkzOHhoAPqZWf2k5cHYzMIuIpaL3AYiXexub7+VpGet
SomgB9z5QLvznPRJe8ujj0gOYaUMj5LHhunm6QUKYgQB0IEEwTK2eJ8LBQoR9m2k
J5OAAOXkmYAkGRBeYHEqLhm6EMZiiQTMcpXNbLcS/wngVIbGKrhLxIy1xwWk3LTr
CO8k7nTdSoP9+b+u8Nr6HeHEWkBA60tz7moQ+mCirny39hzc0o28Uv0TrYYBB4tb
7iBLTmj2kNmmFvepmcklXwjhNRFamuJ/R8IDqzZUY5Wx43/8/0YmAIu/eroygVuj
1eY3k7DX0cZJQLkYoOpuI9gw7JMwVRxpttxCpaM6S7MeUFYkJQ1bVHdJT38q4aV9
VqCcVCfusKRk8+VLN8GwJW6MmTcqiXIJwJ/B+v4DshkK6gWE832a8gKatAWPsVPP
yhqIPqnO1R0BDJhcKt2EOSf/JCm03A6z4TqUgccVyWzE2nwxpnI/+0Hzt4JuOhUU
CmsiMEi/faFYrDy0OieEb4OilJsH+Slw2IHeuAKckIq5jn9+GnSRbQuW1xKcVc4n
Sll30VO4NzDc5wuUEcOfV7t3zGS4E7p8NSS4pDak04OsDUPK9pfHWaEVWeLNHEWQ
KkIg8KZ0LTn1H7T5UpcEs5/yZTt3laL1YR3XVMo8sBOkt0aQDwO7S7eZieu5Y7cN
oMt2ITGQR5+SFRDi4A2XmeRO4xhyLD++Q+vBBMC6os/FvJErGLeM5uZjcGsnbcaS
F2fqoLTPUTkai27IlACCtoT3bEu1sQXdxU8PMNcQPHHd894vtZdQVzt5rmS1NIA7
0F30ZTvlxQwI6fHGxi/0r+CRGDBBRqeL9W0WDDGzG3QfFZ5O1kWUHEzS+AGz08F2
GngB8/2wEK+UCpUnUoXDxTu7LSUmMIwMaSyjN1eW/l18N/c/X0zQBXlzWx+hq4fU
15nUo4EWOVOs+huLTgCsVXD3Gs6kXfpELgnyOo4UkCSXV+PR+KVLnf3k+u+hyvN2
RqCz1o6PnKOsnJfb/t3w6+YUT0IGm+rgUKBTrp1/XeLBByuHdI08VC1MZs0i4g9T
v1+ioZCBWfrPYMPYEDslXwwt/OQ/Uocw7OhxVLp37V+kPcqapeAOtTVd2Y4lGgQq
ggcW8wsxCM1l/DAxcGJwczayyB49HSN0sM9eV0AH0IG137xIp1fYsx7Wscn2veGF
V1G9usR4qVPx0H8BatZY1hqYfuhFQwL0tQaW7oukUEgNMt9FsZfgg4A/1IZ3uEnS
HloJnsdXWFCpaOxFCQV1boh86yQ1DctE9RRI7Qi6Chelvm7U7FQqysPMYddOG329
UN8VpBTwaBJi9RhqNBU7fTbZEPEkxXpuDAPvVQAyMRCmdEiMS250xarCHA2EvISz
WlLxLxv5Sdi4ec9Rrr19TnW3nIuHb5pROomn6yvYiMob4ijiGNkfnWg/gthwgYDL
nGTVszHHbYD5hujaVqaTSnuQwNy+r+UPYZXowyEzFkqmG6LCh8o4Itt5U9WLYMOx
TjllVlopYXNe0qB9AtgsysRB+skWNsB5nOQ5XgTtJxZXsgYf45EN7kK9DDAklVaQ
LOGKi2DWVtcccWjRUL5gQHknRwLkc4D6qt8y6jATUIxVZfhKo/XG0kQM+P85Qzze
dQs9v67WsYyXizqb9qkTAUa1AnmWlbNAKZVoQccLWzHdJxRgq+j6oHU/WViJY683
2TIr6jOIGmQ0RQcC4V2waO0ErQ2lMs8a3zYyxPeP55GCFgGmmhUemqNqon6eY1eX
x68nxTP3pJxCmDgfw4g6V1xNdgexxf1VpO+Cks5ptDbQCNlq0OH6sbRymC1fF6Fz
3tryq6mUhn4N8SGc3f8H0zemZg+LHdR3STHP2C52NZnQhVZjP+uNGWUMzdp6r7xf
dDk6rIVddR3oOXP1rlfEtF6+n3gW5cUbaOMMkDDA5NQr4o0tVZGdPTffBj9flMoK
hMuA0f6bp7ujq1o/9eSJdYleTLvd4YA7e8lNyfqkpSZKNolVKwNRj/ApCC5XqVQP
9qxpwLY/a/CZ8cVT5kk9zyZ5gOsSx5jZi4Pd2m/urCSGRxCvzm86efwuxOe3+/Q0
4xTaltOe0t+mfKDKEc8SY2qFuU/MJ7B4FcFSQ4rRm58SfbxY6V3QUZP0lVgOQ8ZJ
eBSfGCk2z8er5e0rQM+V9OGXG2W3poxqCzHrRDgXxUWKsGN0eJgihR0eeI1VNBBL
d61watDT++PB4L1aHLutY4kUDEm+BOv33NIO5QNvwiiN2eMCQNRYjiOe9rsg5yg/
D5EgbW+tBxYuqfaz+m5IS+/YSh+Pn0gDr79P9jDLEDkOxwJ/KnND3r0JlZKQM0bg
Ubic/EL9YGGjp/FEIGChIJcULoSIbaGFXNlkGfzSeV3VW2F7rSVIvCAv0fosEfjC
feBqR4Hi4Nok5wAY/jqnE7nRrrz9dcU7BDtgpcwq7uSa1Gd+Fl5iMg/KKIx6o4Nr
VNUPvB/Tl51vHTX/niJisBkLQqqtHI5hlcFMwsZ1aanTsJRVuI0z42v87KlHuSrK
SPyJv/I7UjoSRR0J6Z0kAFj/V07zyA37U5v0Re33aZlR9/z6N8o8u0veKZSIxEZA
qxwK4upbI3XaWf7Ix9gfBTpJQUE1YwG0OIPHswo6f0kKEO2hvI9NQw+3nI9HPWwC
I+itfBnN1bHvcRpJM4JEr/ba9JhRTaHC6SittyWO/MfTNdj4ta31P6Y772+sWoGr
7tFxJVMWxy1KtYhLec6yeZuxqWxAM9Jl6z6kHiI1ThyxMh8vZcyFW3dkHW21dc0P
KUM184LWoxGkBUmNvr1RCwShoXxGClXlAiXtXaTo1O+ePHxIXaLNtSNyUfLlIK0n
TgfjjoVb/tCJF7EcL7DJsYrhnXnlxv4z24Gc0yYPI2n3FoAtZFnRLy1ekQZ3UQBW
GhFHg0KSKGmjRdP4cLBROrTdYq/UksXYHHzzdxLQCwPhf/EGBvHneZgNfoMnIqZR
Ea6MAkdcJZAIg59nMuEc3d8kf6PyhPDCCOAY+L/Uu/un8N62YLkP3QsefUbap4cb
p6g6RHvunaz+YrpKCWn9iDOFqMW+jNh33HsK9SyXeIdYbwp+fnScm9c6EnYNrOzs
NBUknqkhN7BSFmq/yWayeAlZVkk3UDKrLj2hOcyOZXSgmqkGC8hFcN/y9D8fRYvb
Euos0MA6Mqs+JfxbtVqtMNv+O15POFR99GZPQznPo3APmoJWzKjuPbR1jq6j6wMs
HSESM3hwUZuOEyg2XAHLZxITzvxI96i6l0jAkIVHfSGXq/KRPRGZklr+Z3GfPE0g
r/kX97Im3PVXhblgdQSbEKsL0AUMfNkfhaYRGwTSKGDR+wpaDwU0okFDW2wOnzgd
YRxLkxthiDHJ5/uUSplp+/5ULJqDEzhcmy2/alVN2wcj0vss3PZXZ9Ezvjg5SfZd
N+Pf5Q5gFp6+WCuh9GRnKQAuhPf6ISk4hbnsGtA2/77y2ExpMrg93iZA8SMTIkT1
xUgMdH8mmwDIfjc5Wdjv4QxTwMDdJae2NntzjUyY3lVo6kDuezNE5jq3COgxV1F6
niTBLL7cQRmQU4P3HrxlSoFOr4BfTnnqVVaNEjIM+aqabVGwcnKjyV2nely1MlPd
0OZGM0m2tNs33AhwFfTEee3q7oNbNWLt4EB1Pg9xBgPcsVMj+GWH2QTSbe+Rihx3
hqlhDkUrWCz4svDi81socuULIui7SxNe78PcvjoA88ipxwCUtHhNdeXMGfk/t7Zl
6fDFVMRzssPrJVPCkgnFbg04QQS4ozvqqyRKwvRnlIi8ZPL8EBbDjUhwZWs8r1e2
8fqbJFoT3PnWw4/bh4Nh8Bh81yd2mYgYnt3GAm+gcv1TqotO84Xo4cyUcWhYj9x8
7c938kDSJ67eBpNCeyD0dWnV54Uuap3tLfWVsKjX+D8DEu9dEAbaRi5fBlR5VcXv
QQUQLdcWPfjbitAa2gsljb33kQv3BNQdsiwhEQYry3m9SJfgMZui6SWAT9N00hfw
1KYiF7OSCgbhpVDZ+ySJx5SZw25v9Wju1cEy0B6LWyZIsHh72W0nI9FuZB/SjqL8
oXyhq1Q5IOl1dlAJYHIK4QMaZFgI4VsiPzNZS0zUcW63YTBFMQLYGTyrIoKftr8F
reFO2h2WNe8UfGnHU6prdSZMztmdnos514xQhOcARqPA/p3+pvunqv9D1+eAi0Ii
kk+WoYUhOYss90W4Edlrdl/asZJIbbDEsvHtPPx7jVA5sUPyNaxZNZfR1cGs2nod
r7jYb0vPzslEH2OnfNa6uCd65NqvueiUBC3BmS5s6jZs2hTViDl/jC8F8pjwSn12
Rfa85i2utOmZULBQFDr9kQtHa/NxJVX8Oaw+7WOc/CpjUXC/RC7zBoFbxvWo+VXO
/njT+FVnUKiN2DPjz9m3s95f3Xh1XT6jLgA/CioAsMgwmqMSYp1BEKWnJ+7PhzAX
GNRVrwWeKG4ACHgjrHBS/87FAQ+3nw2TmB8q02RhmR3Vrr76ccZc2tF+AjeSS/WI
iSiyEa5AIoaGDOQcVzPZe18n2neaw+U88fktCpjeHUIkobSQkYbk1v8gSeCeo1ej
zb6vBm9AOFenWq6ksqWfZfSPINVnMUtbabtsqCge9ZXU/q+X20S40m2XDdFrpADi
3zb3rD4GORQgTlRfXC3TuGbPT8RwgwrN6GfnKfioh/1qNLaK/xK0oyrmUKOYMRT+
xDI01A47fmHIBAL5gjvh7FnqJhMxBDbFHHrdBkpkBFVl6GpYf+lBMgHJC/TOsj06
T7FoNnh2AK2Zt5EwjkDTYURUnvjAiY4xkB4eAsM4aNEWmu1qV8tcxI6nqLhkFDo4
0UDWoMUkMuwaZsdtCns3xAv98SR4j5OqNX/MHSxceIOkt8Mva4NbmqDvn+5Z9CPT
ib7FwzrHtvawPehDJvUik/QkJ04tucCY4PxxudoPM8F4wbhLb3E0UZ2r0Wv/YHdJ
XzJsY9smlEGDOkS8wdY+tiKnlPrWryubzlaf3aG3bV/faTZhRg38TciWkVBfZj3G
2+FoaWnRZi6OBll8+RPm3v8XlY5iEap39es5EYRFwRAJwm1lTzXBKs/AbgLvR4R5
vSaV9eZkcbae3m6PTosTjTrDwYKgCllYMtmFmABNNqwMlsOqd4teektvI/52pt7q
2bmNNXc5DnKPBJCLWDZXzyTHVeQfLoP2ZSQ+oEyISJ4c28vA3AqtwcPGRbimBzbn
rIjUF3GggR3Nq9/rdGBlzcq/InEoa2csj8oBI2lR0LrY0K+6eVOKcRZj+eaPUuTw
0MsjV5quaru0dquPlLJKs3c/Ilb7eEAyUyxesbtXM31TyBjjdmJWbHQP8fHEVLME
gARyTu8lFwIVUl87329SuLuVDlSJRaS6XpkmZzf6XMQsd/GUNv9xfiarAiom9mSI
yZniNsuTXauA/XKHVUpnCepO9jWw9Um2AIfRcIPqRWw+CH81/e48oGcMz9cOczsu
5/3+DJlKLJnYNSL3/2Qz3pgVZJMQ1joDqDYw3W+9GM/vz0twlOfHR9U4/ab2alz8
ia0U4JPDmGqzjmy1Y7JpQzENNgzvjxQkaJUwWDzTWv/JMN5bdPZFYY6k9ofVcJbE
NTFti1IN0iOQvJWcg7dJZPPE85Q3vldzRDvSc+/RZvSqbgr2O2VFEHH+uh9xk5Zu
Rm0x/yeuvuTXV7L/Tqw2m1JRlyT1YIs2pihMarn0Mzp4i+ex7+0vpAq2FD8Cy5zv
miIA2kEFxGCoAcui33MhtLBvUzbGa1VUVGv43mDZGeEKmb3jLyROeAuifjEhJ44f
5z2ofBwhx5a/HfhqSQ8gp0F9T0z6/dFrXwkjqOzne5ZbRgbnnVwJpTTjMoZPtVbN
Is+EoozeG9/7h+hnD9y4xn8toTDNm3XWWEQj9O40uzK9A8B/2m/tk8StSrggnvRx
lFcffKwk9hPZC2GjKXis4TTyfNn/eJ2eyhzrJujypwGeKocrZLNaNu3WYc94982O
4XvsDa6Ot0kWA9fx9ydbHeDjx2KsXlte3MevFCpodFbQ3ZDuS1n2TJbOW+T2Czgf
P0Mnf9sJVi5XNAyY8QL1RJcABil37CPiPQlZHBvgA0Yp9OaSvTeRNZCiShx/vjeH
WGiblxTLu8mUY1Pv7cc2K2pINUwzxzjGXR+1DE79wBOiR+32YtxJavTe/4SKpJG0
r+/JVM/CpdhMwyL9prOwr4xZ/fdhr8jTLaoQodgwTK34MFwxbRmNrEtr8YJ1XCXz
IjV9MN/ZU5fSq3jGnLPrOPVHEkstHfpjpO8xytdu/UHrPx5aFaE/bgxgp4D82MlS
Y6YiEywyU0RpaQUIAfesuMdwcdEewq6/lwzjfqR3437xv9EjksGxck9dAhpUyHxb
TfX4cWHe6t68qet4GAurXV8zA724/TYO+R19M/omOY++paigoa6nUYD3ktldAa7r
EekLQzA05j/9bMX4LDLpJlaJQkke18v9v5fJw87w0HQ3V+cTAJwfTK8K6GL0EegE
YBooq+HJOBdhbXPztEyyEzPLCAh2gppz3nJfsCrTpcYNjz0hTKT+zXUpSWSfZkVt
Y/K+iAdAzawTYLHRLSGkpdXZdt1rNnsEiUUkqivT/T0ITowt0D19zt/4oIhwSftt
jb35hz2/7pHNKZzDTIkte18iDPdGbLa8pdaUglNIuYcHztki3VZxHS14G/oCrc0C
tsPFklHn0tNsDWwTiIsjoVVYCBFS4fjfMA0CkfmewwCl0r20809rDAbsRPFPjzFW
fbPF9KyfX4WQNJVFub15zYy9BEjOpVYhT2h2KIpuy+K7y1B4g0Fs6uMcXFzZStpw
xF1B2+fOtfMmeWVFHvd7dZZCBXFQP2PwTCI6MpoBg0HyZ2cWgIbdWNaE3RtD6Wdq
aBkaVCZTSjjUH1SpLVwyh3g5Hg/d6ZE0ht/+pae1otjk124X5LQi1QSkhDZFC3mN
oI8qHdhKOgbx+8NPjHbl5ITekMdqZnUW3tS05JiDNDVms4PkYTHZz53acsvgDVy/
Ot7VXlOhfVZkTvly9otwtvYxMh7pyEcdNpcYuOc0Dy9yS25LtpeawCSThXJhwRKL
qV/RAE4v33M7eaSrQS7LsxIugIUizaE5cLS9Hhob8f/RMpX/bTENe46UVON+y8cf
0XITA2zIF5JiOSTcw9r4th4gU8gsS8LbVdUMZGqSOsao1PimhzE9LgXc3KW5UHGv
3uQHYNcN+ReB8ufiO0a99bKhnmxsKOx/dtnCofLITYLnD1eMSCnqc/oT45I6cHbP
etR7QQ8FR8DcVDTyAcIhWbIwCM1XiqX2CodirsE2ZqZV+YciKVEW9S4/jdgjSXqA
D+FnGELzzZbeK17iAPqQXzhGWYn7XC0N+ZYMK8rbsbU4OkNBqQtNcixmNl8JEWnU
84d98CQKysl/7LZ14RfG7NCKadtZai1hvAOsBCaFJuodqb8SwoVsUDRdQ0dutv6j
l/rfTQTGCoOEIn1WUD6C393pEw7VI04Dk048GpM0YH/F0lnfPL1DoksBakRbAKkQ
S6ZQsG5RVT20RR7IWglE24LFWP0az8/SJv7I/eUf+9fAHnNrLWnnljqAbl3mAGlT
Xdy4M+/AHiCIE1vB7S4iMVSRKCwXNkSG4Ds6Hr2cOuNT9m57CZaO3f3cz1j8jTpx
FnrpED4NwsAZGf9b5na3kk4Zdwv8CkB1df/fccM4OzxX8amNa5fYv2tIpdhfcmno
a6xpUGhaaHYBOZKPauqXvt0E30a7wGYrMABsXJrclAoOAKStRJSp5wwkYlHYCZMv
4lGpfqjK4IvQ3YrrKwqkPNhFIdOZkEZb1X7JKi7qfiTkNKWml3Zj1d8r2X56d0WP
s5GAImbxoi5vf9HA26/E5PCDncK81CVHQ5r90o3xBQFZfsoXk9OUFelI27JaqASJ
BH8uN3pBYYDcQom3kc9xcIvM0F0gONFbGtLsxOt9d3GRrMZ94AnjjvCRj+iq4Trk
pmwwsK/iNAoMh5aH7Ht+17H2TS+FIId3chK24D/PdoPKS+lzMlRa7Fk5AHpR9ePN
zd6W4kDe2NnFArF/LkaG9YqSrZqQC7yxLSS+eiCq2yH9G07DPc9VlOe+PnpBCdba
BoA2kNP1HgClmchWAPX7MjHEA7Yb5QUrk+3RhMWTO7lIzsb1f8kiuMvwsYVEHJLC
fr1TwuulrbXM4GaFIyvFurcAh1d1lrsPc6pGq0ISoEx7KIhEzMC19AdasNE2Vz8O
UIIiGEvYlrUv66zm3CuLxkEUFgTTfk+I7yfhyM2qgPjHbw/cnKbKpmQluAVW6VO+
3WVJC6WOao/BkGcidwGUbzpQaMTus2+eD9lGbNyyjMn9Q3tBw18zqJCMjIO8BuXq
IRXyDKIUOi7VrZqrPQIvBZ6mlrI+EBh76pbmkXzUxugA5124YFRhuDP0yYWyZKAT
AvhRNkX5tNvyOdnjNhuR5BaQzgzoTBY+WDxVz3qxmhRAg0PPD0u13l8qaPahnL+3
vPLon55wFWJ9n9r122Qa5wNx/LOmDCUipwhil0dx6dy3Tec9pWLtcHH4eZW5sWob
4hh9lA4CtiQ4GrxI6X4I84N/N3GQm4rL8ylFkGBKJFxA9hGYmvKjOcE3sKfMptZg
CJb8qUInQc/vv1skcEVpUZulfYE2WMwZwA8HfpMqN98sB4aISFfSFdM/QvM7jNFq
SIPTyl8U6lXaBZwrozHadYRNz55HR6ZsKpz+37RP+L/4coZGlFQIkmhpp/2RBS1s
micYeF3/421HA0dJ6vOsIokxFhwz2Wopah4MBmHGz8wdwKNdXcFMc1yRbbFyKNpm
y6nkdYqgggvSBylWU/cH6yVkzNR8IvNVMDMvajCH+YZF/m6MVups+cavUsOXriak
PCQIvp7q0N+p6LqV+M+3H/LXYT5x3dQaQ5O81i2mPtVkZMyfrxMS7b4ON8b+ckb8
i1pD83pset9LBgT/FFRE8V0flG+jZ33I4A0f+CbtLFS4PGD9EmhUSutuNX5MIuEA
UwgbPwFkBdgzl4A+csuqFNN1jbYwhu0UNSVadMO649yR+M4wMmWwYXeHC/6QKpJL
QMSeC0G3dCZNbDkzJGOp84DfdtKWRHEizhWakJbmQql1CcmdpRz6jgtjlSF8q6tA
VEr1D/LCiyvB7Z4fp8Yb2RJVZ3JXGH4vrHT9my8oT1KnRDrVLgi1gl65apxI7f/X
NMiTT06XeHWkLxv+L4NXpAbc8RRFfpv+yHbPZzJcPg4tyJ6kvcAY9HJ5hrQEp0RX
7QbCSrGgYRfFUVC8+Lw3ua1hlRAok+K2aEK447gn6e70Lh203SIagjDq9PrHZ15u
DvKZ2sQwXWZtk3zY/VHzuubBjkgMBzFVNpvPjZcc8dqi+icvenYYYqxbf35a15Xg
MtingkzWGIUdpU8/PX17D8uSv3GajvNc2XpQ+ljpN5FyzSmGklK9rummogkCzUQi
Ikt5VQ7zTNhnXF3Qs/a1uACFnShWnL/gvAmCEB0YV6F6w+gLH69sQYltQyIu1zpq
ktXk0toH3dhdDzwU2h3jj0bkXZB8Q1h9wIqSJ8hlO4uJZYc5hyzUKvtAj87kt+7R
jezNrerib5dJpj5tv/VU7aZiDbbQkcuNL3tCFAH7FKfiqavI26Qm3h62hYWcmkam
ZnJet1A33zABqf+HFiRKZnyd/+2c9FtX6w8RRs+gzqOCFI8HECIu9/MUX2GIzkn3
47XmeCtDCvVacOAaxOHKVbwBV0QGfFxaWaT+DkbNIi/zL9TUzz08aCsNF5C94QES
4IREpklbykAf00/fd4hiNwyWvotqE1uQmQgCIbIsYPdzRQKyySLrXgrSTTXPdscy
gAi8WzDXdO8KIWQ/BMm2v1nDHPnUHEk+n3wFlQ9qq09wPiiQI2lsxj9aHsNN6UeX
QrcwdRqUd4R6xjRzwQfwR86jBGq/rTdldTgHL4U7LWcUbHARfBPZS2LR2EXEt8hm
dM3yKmIGw7AEuP62FnANE+wM5LWn6GKJD7XujzbVjgA0wSgXXGgQJuBynkFTUzAX
Abi26CPuN1RvcRr1+WQgQQy6Pzkb1RpgTkPiMBH30Jj5M5sNYAzHhHMjLimh9QyN
Owrw8v9Qq1BLFSgQo4O4jGFz7FQEF/khyg5Xp4mrdriRO/+dwyeCRKQ617xRP08Z
NgDO8U7OkEWtaQCrPGaEAOWPbUe15Yp1yHfSYOp8hVb4v0bx1i7ZdYShNHVibNq6
TQl7AsEaAyJ4GNyYkZm9+SeZuw9he7tpVp5dKrNrc3Uf9LZoYAqWoMGMKnU/kcfx
M9W872I9YFHQS8P2JQ+ycnwS/gsI+sfp1VF2hk3snh7OnX1MGz/Zfz9arZTov2bu
Jz5zudF/pgAIKhsQXvql2cQr7srMyo9qS2Aq80gxeLm2hRMLPZAVfesOmvOvKAPy
fJ+siT/HNJPocF9beCAZGlAZeMgTkZocbxLn0OX6wA5nChF/cS5sE59BYQg6iFmQ
mu5K71Fc5VtAnZVtl9aCH+duPnIItq34Rjp4K0mCGwbLzbNbYF+vlxZU9vblM1bL
AQui9tPcSvB/wcOl+KF/uOmT3lBznxCxRRh+o9Yw7s9Hc1Mlpe3VX+qTG/Szm6Wa
XMqdk94TmhwhKw4l9U2sE8nCKNBghn+eWeBkjTazawa9RJAplQauFdprCDBqlO9N
ec6Kw10L0qHqlTs5mf/m+AI34LJVk/kRsyK0OIdewbvNmWsSywOOwdLSKy+yTM0A
IMoIi4rq4tdJLQVc3Hw8o260JByMhmkYf2qgLRzrAVht/QYbOYzIydbhX26vGWSj
MJa8Z10oPAQLY7AkuWFH+o4vI6efg8WjNzGqn5hOpON3e6SL8YYw/uYAu60Nmb2d
lfwf0CMyHg/i4dCCzcj5jrEW7CYUvrJxHDGO8Ekw00erPoLko7dRX/0qWbojTSut
72H3saVXelwFwDLqO5J3Oi3GRjvt610zuo+5wko9BNq7ZVc93WUxnQmRz7fsX9th
OaKDcdLQMXePObaSLIiTdl4qdHsmRHog1R03N65Mt3A3w+hayC/WmG66OzLcr6LP
Kk4A/0v4gX8spbbFnemJZoMXkDYtVrLxWbl9KybEjEP22T2JN+d3CFZTI+jTe4Rh
d5yC1fGEdRQJ/tNRM83NAyLJ/sVtXQsqf9Q/RzUB10Oe2eLmAIsCVyec0Nlp9cv6
/TUQvrtEE7mAjDrG1oiFYDM3k8A/3WCUdMu7gqkYPcxAoGyBzMCLLcX9LUultJCb
VqaHypuO0Ak+H84++5wb/wzPy10+dy/pk4c/btxGwWHoqhdwG+YuMXH7PJG+YGuw
e8P26KN1hTDMy1/WNckvZXk6Vt+rr35xLHhbMfrLebhkrvPyedCUkkgGaiyCsvuh
ScnGxguula9BqNxfy3DJ1mCv93qbgSoUpQKGRiigDvb0VoRSyqbwzXDBXUgDzXKh
eK1MV7lF6a461areqf8m/d6xz/pxoE8JL2HAbN/MRpWuH5tECmlTx9FytTCmMXC2
va8pbhngQIOXQfwtZN5Bi7g+i94wnD2G9eEF3ew1fJSJjPyw9/dMQiEJ5iPLc5xu
rYGteNKIwv+Zn19Mf7kBxwB1PJG0g/tTMbWXEBy48Wj9suubWN+33q+6dslyEHiG
+RawxQmC4f5C4Skqw6KSgbiFrkBQH0DdSN9/xZbN5eQyHQ2wSnAHLSwkraqS6ZW0
BMN4x1TirUBjBJdKXKaFfvOKeFBHFmASAhu1NzEC8BUBVT1AUraip7Vb8DyWVFwH
2DE4nZ3x8viojwEaVi0bO1piljBX29I4xjzN56aJayhV9zmDzEZnwyoZYjY1zwW3
aFr9T8TrUZ8NaAZS0WtzcLr4Fcg/BnCuNPqLYmFcYn7zywbJacfNxRqy1oxAT0OW
GeBW/osH9ZUOT6ayaE//FxkpntJwf6x2S5i2Sy69sjoXxHIQl1siH2jv2ye95rlR
Joz6G4SEp6HLcdm5UFfQYwPPRuHTnnuJpRGjKQlu810LCxbsr+pMZu6ZNC025bP9
pk8cbXJscbDnljPrjTuhBvCgysYQdOJJYdWxhfNkcG/mVTHLnAvkb4tIsry2MWVu
AM03No2dmHI4vBhg6eH6oaWXEJKZikzO0YnCPNHLDHYNxTbwcEUx8KkUXOiaHGgV
XqQU9CbmLHVv/QzDA/6icGLJze7X36VvGrP0fyqPgtibpXUWLgxr3hZpLamKJ012
CDYwp6wB1uy6T9hY1kXxCd14OO/+lFfSpa431f2c8+G8ZZaVjyGO7gpVaiPcfzBy
Tscp5lB6wGzyJMrGtmjMBxWH8yl8MpFh3POJ9GBCKuNddk3kmdqNgW5dhMD/TPa5
A+DJu5hbZ13j9FenX6EHW3brkQbNnrdt8G0DFyw34NgYyBqCRKDYy8ndlrm7dQxr
5/nMAfI2Sqpt70UWLLCC9TIqgEDGQxBHtu/mvCXAiuXXS2uAc+Z/VCiiEGBjwA8t
Cnv+/EH/op7V1fm14JlnxRuanw7UqcWbq3sdOtN/M2jIKfxxDA2c+QyyY+/AoRXp
QnxuKdLW7F+QJiXdbOcq/aGjKWRbgHbdkT/+tRn+iilobmJ/p4tV6nloL8mtZsBx
2+mSBAUw8RUKNtKd5FrYPOmcXerEfhbOorL5G8dSRulh4PNQOGtRRmpRDdlNrRg6
GlqDfRPHQI+nQw+EEsNCHph/csum8lJG8md3FmuVuBWhTs7uXr+MyihQ3/2/3zqZ
qGSAorsfupHm+st+YhskMM7SE48eV+Tx9v3DOTbszzaMPH7vSxdlUOjQTEUFsXBv
Av9eGpHyt0ABzXFY62ISzz1KOUviMtlPHvka3TowvnAZ4dQ/8kt4e+WpWXjMERtJ
8sIL9s7bWGF7RPW1YMKIdEpuMBQ95JpZrQb42sq/wKS8tvb3RJKDQcxF9Q9C2Nva
F0sEGSBh1tEnYT3ZhrB6cjW84PebVSDmXGgbE21dhklBZSA+J9kqNknzGz+Rm7WD
ycZlcT5pNEL74rroGcx8xXvM4Rq0kkW8PRstAKvbgGsxmPFC1r5Qry+H4Batz2vI
kLBk9SRueb4GiHSFpZFQGLS71czbW40bo9CE8Lq5fivlrBaRiQdW7prnwyG+uu1X
guY1CYmTCaRQ0dBCeAInO2OOHLgazlLnnINwD3dnMttZ9sB3jrJRFR4ipOQ793Ed
ir/tUJX3whvvBDXCeRXgdHKGtlaYksxsiqYRq71WpQwGkBWlaZsE4HiKDzz16Gsk
S7zfGqami13dhvWWF3DIRlD3CfkRGl2aBgiG9ZUIPYvLtDzUPWUw2Jx+3p9JS47g
vBvjLBXIJi2a2hKoyw48AX/E+ofaZQ0KvZgbm/zV5xnDQoHzqkCnnEK8tklWSlJa
ek8I65zCHKNWJbyUFY+YU9VHKxHzkh/OGePe4DpnjCJd07qatAYHiuGdFV/j5LI1
/Jlz3RnwAgUKPM7f0DKdTFNwIjQQRhRLtgCednEMEVwy1W2HkxuBl8A0Nkvk+bT6
1WNzvgr1f1VpmccpWopxNkNEWba0yvhOtN5GLzf0VjD1fOCGq+GsOVe/cwxu32RJ
RcYI6AeNa5Uoo55IDXuaYhB5qAZyCI+bGlnhL2zEovjB+iWCZpvI7DhMwjyfqXOp
eZWaKv0koCNdEgtkzeX7XvuG9NOrEzf6XGjTzv5qqduy6gn2ifZ8XFMuc0JtgHwS
qwutmpUaSUrmt4uHtLrPQhEfZV1BZFf2BZ52tJP+rtZEIOqXA2cutjWRCNdnqIDM
rx8GGsoiszxysgzlcMolPShozkCP5+/ulhW8gZUEXqazI+TY1x+r6voQlREzEmiO
Fy7u+oZ70p0q2/cSDhGowj8N5S22tdgMbfWK3SNGD8aR1Cyb7kOKFhGrXlK+T8nH
aodeKSo8MODtMrEFVqBPbk3fK4skd+Ivpu7GGroPFjDjp6Yh3DG/dmeXOC6p1hpk
`protect END_PROTECTED
