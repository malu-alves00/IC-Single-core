`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
f8LHa2JOqaU03LJZvmJg0Bnv6ZXcIblfFORZABOYA7XbQv7aXJgs8KEjg0WpJMV4
OsRYIOdBpYx+8G/duQGOx1b8IZU/XTvfLFmNjgqsTqCu52/SupM+l/Ke6uw30ZSZ
jUsG+c/JShk0f4ZvGZNUquJqRPOergp3XG0tlAR6ShHb6p36VyhvZpIBbpdIh0l9
2iR6lny7i2zVROjSfAC4AVDTUgz+leLMyVaar0xbYwfW/X8GiffDhJwDO+1j6Wz3
4RYFg6ymV8gy3As0K6kIouLntTt78QefRAUubw7WLBp/hnXpMUjHTcbVUiL7Y3Io
6jY0VIPq0LNBLemRYTB0SozKM3IQk2vhTn7S31MQxMxzqERJcXk3nfLiIQcl+ECI
OVjcd38FyGCMnu1XYL+qIeOtkt0O0hm5mtzw+fpw/qpHQRkIaI/VhEOXgLq+CPEp
28PnEKL6RQ3toKO6+DVWNhrytcxiFRq5q8g5hm7S0z5tgBoYfwcvKfE5DmjQ+lr4
0hdwtzix0yFZrSP6kpI3fhdRrMKk9CrsrAGZIDv3Zr8vlM9fyMLfxIZaYP/UTfzw
pG01L4fz63EUKM8cJ/jpbr6EWPpWNuTNj0JebXcFAHIXSQFOoRp7bxWhNCbNlCum
U17Hn7pg3c51ST/otmSueEnJMdZ9tGCBAjdEPSR3nW6sxf8jziwTtJ23PzJpSuMc
yL/vPIrlNru/QLfuo0Zp9iQ7D/5+SA2axJ3lkKeS8aggLJQaUspi/6UpyfCwVDZ+
QtDlgTKdIWySM1GsfClS06UzkCG9nly9Oj68jxPyvgRqBZBl7Uq0/xSZ8m0jdPij
wJlSYJ8H2ANw1H8CE5E7BAZHIv2U7QRqE3DR1fnRiMIkJGYDDvqZQHmP0nBQTmQ+
51WsuhakhN1po9u6H9YNIFoJ9plpwYOwOV+pvdQCxyWLCoevKMV+YNPIXuqOzuwp
oVuO9VECkWSyP9uHqr+57dGz/MNZ4yBy2dF37/XigHst1BxHEpVw/UlP6Hv7wYVj
P9Mo0SjNZMZH7ev8UasLrRMtF4nFevBZBiR5sD+1RX7PQoy3ljltMp4w5KpDrq5G
obhlhHZnGSKvtYjoq0Pjs9yAVPwz5Q4b+yQrDTh3ORx5INnXFjIr/aLOJ9PuimJ2
AePI7cF1lhHwd8gbA81QHqkxttdk5M++J9lfzj9dp9QZToC1aHbTlNDVsrl2gA9H
Yzk+HzYfHen8NVIraMKfOF+LPjfdmJDzZNXiV2PTWgRkuL8uIPBNJfvRBUdTQbkZ
VahhtSNytJoulH0ldoe1F2bAdamVty1iu1kMA9Wu5Tr7iArhL3EL4nEAfvhhesBw
dCrl8SMhDbpo9/UpCiE2MIu7N78cvDYFvvjkEmgtoWGJg5BO/7/+9GfglqcfTQMG
/Eeo2/COpjiZN+bXnEWmcLIbHyVhBYzxBHPHtsyk0hAVXAGV+rL/p8o0Wb2KAum8
TzfnKHmoBPsLEDYSD5/t0hKgtIrpXKcYKX2h/fi0Rt/d7tovj9banuPhIZB3LMj1
8s8HJJVRyS2bsph47h9zI00u0soY8Bg/9+48dqDBdfHkanHQ5CGewuh9pAT/xJKo
iRNuKLV79DZ50oJ2t1Vyb1Y3A6189LrqmYDze4cAAQkVsTTM0RyR1COnH3CvzS0w
45Vvd4vv2w+68FaAiD1N3Hk2x8XgBLtJyaHQ2sYVNnMOGgqHZfphLwm5fVl/9nA0
psR/G1+EPCKJQJklURo8NxwEg31NT3G50GfpGuzIpH+5dI0BLTgdqsbyAUeqSscJ
5La/i88uy4BBVaXerpg5Sy5b9H69nN+ZW5auD28v0pKStV3gHAJ0wIqOcdrVT7ck
gvr91rjYz4vRDDQ6qUx9Jg/mRoe+dPdCwcSmbk4CrE+orpZk5tgSgPP2NtTY5H++
KuXybhC5TU55RiDD8Sp6QEVsojwG+ZcvNB6QbaKId99kLBE9WPJhEwarEzovrq7S
rD/AdOW92frRMJbKOls1QOA0TxpmoimBqOW9u1o9f4AwAC106fR8nnXsuMzXr17y
K+nGqfyUtEaT3uzdRc9bGMTmjeLgbVZAk2ECbWHwnOch7ujNAAZroiPrYFY5413W
GpUAWAjxd5417nFAlLTLdom52ETLwWjWMO+qFS3P0p0t1EFpRzWHhlc8kqf8+0sJ
AEeK9GMo4HmHz/EFS32E+nxHARaTPLpDwvaM0q3jAZZeS0a/abBho7rUj5oOAlcN
+jdSR1A0wkNB99Jf6GFRmdn38j19pTYH8h0qNx1XBUYBM7sQ2uxiG0oeyyerUPux
VLEIlzfba6IV5GJfk2Zm/qIbvEHuISxla3Qb8MCJr+shG5nMd/Ol+6ZOwCqJZmp1
fVevB/xC5NZBmqcYXqio66+3V0fK1fp1/xMBtXTVyZ1tU9bX+LuzSf2D/Ny+lU2K
`protect END_PROTECTED
