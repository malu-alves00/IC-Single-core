`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eG4is/m5qyk4e1QgiWOK3ZuxuG7B2rs9cq/Paq8OjaU4Fy8nH3KyV1hrBo8QUMAu
3MjwFfc8eSJN6rg2XMu4vIag6CXKfiQfBpP23kl8xT0m32Kpn4wVTZNl1xvSwwmU
OhGEucBWTltrSWwEmPPaHq+4UqznyvI/z8VC3DSSyyaqeR+J62b7ZZz2bbfWjv8o
5/TYeQIUvs/eAZOHoJjBz/17TPil7PJrGrz4+W1rW4hj3YT2u/W+9rmxXwztc3G8
SaxG7Rkan8UAyBawzkd79Ax2rm1KFj8h59lIbNKqQg2n6kSYqWRyJrBhCKTbgTnQ
kkcwY/zyO5pbN1Cg/7tb6OOYXGBXexWLmI46973DvRlk1EjpPY/7fc7v9yE3hSGr
zBZKoLNoc/SHgHOkyyJta3c8AvX+WGGZAKLl3Ufo910BcoEic0FiAVAVZtekoj3M
dEni65X/aibiavC4ZXgkH7Q37bguUTFxEZ3ScwUanYdZOqgc29o6sqkrf4AlTPWp
eulvsU0Zkuj7vjWNvRUzazYG7g7uEHyUx0O20GR0CMDmml2kBeot71pYfNY8LYxl
2bs22vRWSZHFoogLqxCtuSrDCEYDMg+Y8V9JXbRSIHt7enfFG2KSeATfqVkpVEp6
33mzrkGafPN81QMB7AlxOLJfg8th+rg19jvEDcQhUMAGwZ/PKbcLsSl0+M00q5TV
oY88T/32f7M4KdsfmHNEZ6dT15i1EsBJ0jYNTx/Bv8OilJ0pA2YHs484eo90P9v7
vAaooSkHaH6h1rGc+7VQgXW58qJ7x64HmqUp41E5B4zztwCx5bCdTwcMcI29/O94
2U3Syfr2Q0dxIaTe38w5oQxsJnNKd2uAqPE+kkqASRgz6h9A9I8I8yoBIpgz3wW+
AyvjdKeqqaB3yr3TXgrcv0HDKPnsnzNWrbGUEK9wFdlrNYQ2G9635oC5E71N6vYB
FZ0sXhCoyOtXP/wPTbAMSFrKTjElteekYDP6vIagWqh3gyMckEggR1CT6jnArGd3
XpxBN4gVIzX/m+d265RseG50w/+LiE2oMgmtyUNrdY7g4LeQwq6SaHZ/DjjI5e6E
yRowBD/hSPWT3bXymUSBUPfHRX7gi199pAc+bQtInVtfS5sise4wcBFwEL1MCdig
GKx6YhrD7zwNKqUsyCRKH61KncqVRDDzuJ++noNnW+bVJ0LtVqV7ikgXFpnxyW/2
mICLOZTjJv2Xu+k39sfW/Tisk2QY+kQWk8VyQ3ViDtYXRExMlYEyR89tL4Jtmlx5
xlfijzPMwgmg0O/mLqk7LdarFapJTsekrsxu5pxBDcY/YSrdjhm9yObfBUfYVG6M
prltEpruO9H+a/sj6EOKLS4lqvat40IoUEUR77iNu44xorYrppkST9w16JBX7xyT
wL2J1CMza3TRdFYEXhuh8huPgQBbQ+rrSzbLMe3VgBM8AvJrrKGQ/zThsP1KNtnH
0C4nc5ouwKqngWMMDBgsgAfb+QIs4DDC4WY36Gdup09SRJ3BziWwfMB9gGqsiS2O
rKuOA89O1p//v4VZPjt4NvL/huKbxgbjzuPVs7t1781agaP0OTtvYcZv272Ewlj1
1Y58/X/jYIpJOU7x80mfTIR+K4sNWV5CqfozSkOjp0Cu/7P7MXCCI3rlrvqVjGIJ
RfIqcs2nn8aLKQGfhMrLa223G9s0f+0X6ViYJ4XBXHprj5Ai8lTOFvCU3Sc366Q2
g7M/3/CI0q/4fjlVCtEyg3a3ZUmb4gJwL+1t171rbWsKgPi9B1lpFkyoYGSqBDaf
uST615iIjZu52w1EgbGtxywFGPEDrgv0xqOrN5Xcm2PN39ivGMV191gvHWtHtH8y
/m4Y7l54AkNgkkTgtwScFgxK9pbp/T+G3yByt/P7ZGLjrqPXO5uofjcHVHHzieSK
6Dcdlv8gCqUy9iXCwzpgxPb/LAJqODqtXdi95ypki+DkwpJ6nog0xDNDsJPRXhLt
nrovgXJ/yaagX2my74y2KVreExm8VwqZVwrHRT+3JyImYDbDzcupHH803ytDB7pY
1bNqqmYaFU/bddrHEwpSwobdRe+eMa2Z/NsC8nmZ8d0kQx6TNoGwUbztPDV9RE61
2Oyj3V9wEH9DyfDWH6/V71CYieavANiLFKidT6pY0QTg9xiENaDyT9kUH0TkDuZg
aQ3I7ZMno4GQjJlbM5uVIFf2/8ut0oln/1AYVPt18jXgERilsKuaTEqNuCIQjjc6
RCP5IiNoChjhQnZghzY3hnGKaKrzHUxAUB9lARK0+tn7o097ul0Yn+DnRHbGp3/F
digG/7egMeBalyqTuANOn5pRjAG77LDmG+O67ya55M6ypW//CPT7DfxGnHC02Y4B
t+/+JtWQIVAoe/AuoaN+d7MA841mTAZx+H8wzBZAO04/WJuiQuoSIGf4lHXe6jg/
0kApJc6S8u1dX4ybWu+tbK0yEdx4qkc6Ma2U0kbgklm0Z0uIhtLq+y8M+D65Cmf4
4oGutksfu20dbMX+F8ElVucfvWt8YRmXF0bgi27mn9NzTbXAmJn+42+t8lMzunls
eoANzvw2PC4qwYurM4f1kkNloVB10GYfUOsSkNBlxsq2AijOQBCY/CBNlbuZ5yaX
LFp/XTM3gi5ALvPbqWWi5kwS9ME0IfX8uVq5ELcWJU8oD02KZjEFQNopcXp1fzot
b+IqrJ+u46AakXi/MxVdH8h/qKHsGsrTb0pBrdcQpGGRbRQJbgHH7Kz3tevuCxjT
ZMP+MZkx++CgmOC0jshDGF01FajFxPQgfvmPXvl+7Yhfmqw2H//dINa7X7E5IT1O
HzPC/WTjyS+lGt1IXQe3bcc0yltd93i0Byc2fkxWlXEyVhoKXVJ5bmxNFB0fvcaP
G4tF7ekzDBoWWm1BEYA64wKUnOhGyH8joTh9nNnX42AGrnoSTKCjMN5RR3IyfbKF
PZgkQrM2kZLt6AE3OoAgSXRfLuyBmKv07YFsSJcLozE9zy4aQ3U2ASQlPRTJf7EA
lm2Git7be6NA6omEniI0sx17rEb74uVQ0nRcGgcFHG62JHn++Z8J+zVse/UB4hXY
2XpRlpHavWBgogWFeXle8azMsbOhGM+GGIGaRiZTL82bsK9AWzKalFY4bSUllQoV
6tHOLweE7+h282OuQvT65o0vYbM1unUK4r4hYtToXpf5ECpwpozOWzWfXbAhnDCd
eKoocYg2J2EFYpUlFAibSshBb11mzjXWDfY4tz1cARD9UKLDRDqEXAHqN9BOXMLs
Ts78P6K402+KFWfhjsfPf5sIsT7AJZYaeth1BfXwqYTEQm0dAPh+A1CcXfC6gEHM
gzqRFBBA1XstLfi0HKgnESBnH32QAY/lGXbEtBcbs8ipfeGpb4epyFUdVZHApu0e
bg9kARCHs9F3Hx96pmTEE/NCulEako+bMvpeye9aQD3nU8L6wjlMxQj+qBdrSHmV
5g6o3O72m83VQR10R0rPnRjuWQakTsFU5w0ZSMlhzwDCz0rZ9no6kPj1dry7Hm7H
2yzY3tMBCPY4F4RZvGsphCFPh0ZNFA8Y+kIKO4xbcuru2WELgo6CQFUwQOZT/1eg
2Syf/A/Sztval6VI2erPqYDjpBtX6HcxSaZCsFbDenjI9GR8v5j8Mf36mDRiVwBv
+F+g45dp0OmzBjejy+bbbiZ9y563aYDYRLXqnJnKdTL4hp5kUs+Hj6rdKpgeUTcW
PZ0rsKVg1WhqGLjwA4S6T3FUv9FA2K9tDp1z5u9n3kV+0KqMyVcTSlcySvzpfSdf
cA+VbXE3LCIwn3wkpKBabTNpohqr9aQhJ5rFO/UsUwvvgiFmfpFeXLbEhImPipBx
XoeF7hPEg/4uQZ2bwXYZ3dauictaAhCif2B0DNz7kdKFegsKkyLCd/S+P8Nj+JqZ
dvRs+7sksn52FWzk7aTv2Wp8wOgwiYt3uqUUDNy133sU4SsbfVG5rkOGD7hQgPXi
jfvU/nzwUuzZ2CtrFL3DFV6nxjlIhzdWyZAmYIBjhDiHYty+AEC3xd+D317u4zAV
lb/f6luhbwZjcy52viOGHW3G8Bp08eOLI4YuO9Ea2L6UJq2cFJ8m/8YFgD6vDNkZ
Z9+7cKlX86VzUiXZ5T/gSXQpgowOyUmUHGCmWWrFSQY0z9k5l9PekNToVzoMUBmt
aZ3GQzoMpE1GZk95N06BAw9L6oxSCb7Wikq+Ae8PMc5Tv4F4XkzUee1ca6e+59EU
/KAS8jQ/uBPBTTCwT4LEBNZRsrEcYkWllDoe/OP4QlrokjhkmAXjetGDQaYIi1Wr
ZPEYiEjbdraxmY+SEGQIayumLubxWa7h9s1Um9Ki5/M37IEcYabZ2w61FTItN0Nf
1rsmA1Ui+Cm2uLhdfv4OjgZbtqnjv9CpxpudmPvnpkjjVBMZ8bcSmsEjIEqT4dT/
gw4z5i+kZaIPxIo5BeJhcBooGitV5tfjenNeYCKESCh1W9GfZTz0FTs2mZD8MJ0R
65cQyBkt+E5k8q9qzb2KUh38b1Q3xB4puOWw2jZaK+Vl/SuDdISahANzoYkJMHtL
0Qenw1PLShRWObS03bNk/0EH5Th9b6kTsixAjdXsrYRXTWq3yIXAzS5uDZEdmq3z
mjoK/dkSI2U7zlwRPt5eH0DYuKLEZc0YWfg7EhA7z8dbsSbe4dbGNg2qRHou7IDs
ueToCA4G2SE5hfAbDDOWAokC6iHDQ/40H0OXQuykURpBUA7WXTWprEzMO8RhdXzP
GG6FHLslaFR2i2ekO+git25VCMk3nu7Tg9kesAr477QJ06wlSec4oEkA3H2BGZ7w
TPV4zmrF5C4N95uJEPCnpzaQmKiB3blXBlSnyYxzwBLCTm/UQlEsMSoVmnz7ntAk
Ru44gQOtLoilN3Ou+hCq2IkdZZI5LpkXJhDaVtyah6MAzlig6+qbctQ4c0ZbTw/P
1YyNuY7G1jAECrwHLgbdGK49N/dvjaNWEZ1g4musE87cSYHLnCLYZ7f3QA6QDPr4
74vC2+sWbPH/RVahm3yT84LZe0BX1VLmqKinBoSIkxqr/YAaKXuf+STD1+ReamdQ
BXWWzwdqHiNs0EeDjo7ce2qNaG4Hbsedt/01PFDYcTrZ/HYAw1BldO/13h2q5dVX
ZvRXqURTzDr3FkxjlWqbeKWQo9dL1CIiTQYHVOCm4aUANoT2OfAisoLP6eSnmXAu
E5SneSWTL9zO2tULPGqCmL1VSeQHmth7pBnkBCroh3Cx/4jRT+4muLyHZBDNXuo5
bCdGnGgExgTFD4ouRGo5CrGXAXxYYmKB60uRP/6kLaR3uwHSieRNhdv9UqL2Ibma
vz46ZrG8E0FVH0YX/hspGboP4gz7E+4eloIWCL+n7z5FkGngd6Fzf+sxTRw30pDF
0nboFWEmSIMkTaC4pSX05+kh380HgAORWIxjSihN+RUTKdjahOSKFXM6pYhjo53T
XeUkSSpG1u/xROkixJNtHRbHqkTJROeElfY1dfnAMHR2chAaHMSiGYueYK7OzFMx
Gf6hAjP1+EwJnz6ukrjDFiW2dFFI/b/fNiAn0u0Nk1hV8rg4Roq+YkQQ/cQeVACW
NzL7PBeLm2YktMBHf5vnQ0XieNrBNP+o0koBC7lT2NCtP7PcxsubIal4NJBeJWrI
HXMiPvXuY9polXX+37GOioq962qgvr2PwWCnLUjnB2EImD1pnWOT7aSNWsKAbOLi
SljK2XLK4VcmUdD89WpOFvyYAjF+N9HB1hKju9c1/UNsQoFniKghWKAjfuCGGH0w
SMwv9QJ49ToEKr5zASUulJ26fcQOC8HR9aNiMsXHSceVKiwpT81dIwVcdU66T+b+
U1dGdNY/i9J2OVmQPTQGPphJwrt8rMDvVZSjJ5svoXfP050waN0mqw4UOq7q+XFD
4myxUlYefCwL2J2X09IXecq7h8hekAUgSWG+a0ojiqbV3AzBX3WQHQj6RcwxvJjY
ZRaEDZwAO9KCpN1c4u9dip//50GnG9h9irPVmL4km2saZZM9Ay/x2fINBxRK8ktl
YX/0Xj8Jxn+UdRLi/MS7R7Ih8W1jRZdr3RaaDSQdcfA=
`protect END_PROTECTED
