`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nTO8N077Cs58tBxasJWFvaVZju53gTcS8A3RMjR3QPWsWGD2f6Pum9yyi6SK4Fue
3gGOZt4NUsa74uuc+qoircYC8OKQX7QC3TOb5NsPao63Qti7Q4zaC7qReRIJfx+q
+nWKHMNcTXeGbUokVFQfxOIHnLeq8HLhMWLCuM4L1eAk5PhvdS/9HG0XdiOHH7qG
H2Z1E89PUDGYssDOXxcg+HM5v1hwjXRkb69QVaw6u/cd62qS/Hfa9evsL15Ct+A1
ryIgmE+gC4IJU1OSRwJB9uS8DxvdszY2fimBd33Rm/CCspyyJ+EniOI31fPN/7qp
/m6ph0+AkYEjCsw9wvK3Xpwwiagc1AIJkk08W6UdOUVWcbjkWaoCxQ5lMmnWvLXf
hv5Saye22aW/HVz1zc3fihSZIY2g9114YJ2bi7CyOCWpXijjwilnqTDwEDgK8qcC
`protect END_PROTECTED
