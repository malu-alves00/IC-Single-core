`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
G9BcafRZufyW0Zx20ZERWMDu4vJkEhXA2seVphzzxj11WpCJWAOwv1zzVooe3j3W
avr+wu7dRVLCp8Vo8De7K46235lxyhIpmu2dwPesIyUspHUXXdplI19ZufXb24oY
2HxInrNYrlzCZ/nFZ5TZQzZONqA/S97Tx7X5lAfd+DrVaOOX1H6c1dFHBEOoT/n7
1OKD5VxNc+MVa1k+EqNhWpZjvXPtd9oCdRnf/hWinLb+kMRUD/uj8ZWeMsS3vRlT
QJrgInz61XzNNUhAvROMIW4KrEw5CTcntoIbsWQSrhzB8yMWdzT+TfJeU1Bq2Qcy
r9rgZW1EZI34f7Hxyc2/5bZeLVouuMaDFgEod2H9GelQSzD1y/eSLLUabsRKH8Df
QhzmVpqOdRztArq621C0ky6d+I1R1BoD4T/bWuUFcuOWz0zxKYrGDHEfgJwqb44s
crCZI0/8+uiUEDp/n7mMBUndPxp9ecKjB9RKaK4Nb0EoW13O5fbjrTEnuLyvRmsB
keRU9+DZCyGuj9a6lXEAB4HtpaCCcn+0DZtAklF0f3NZXRiqJHlGA9tkIibN+GP+
QcbEeDKA+QALKpFJujUEV/BVZea0YzmOjy/3wIioo1qWQUlpruEFAg6MGSqoZXpS
kwsmH7hgpu5aD0JSQVkAqVh9Ja40XzRB8c/oJkPxZJwE+83+mzvS5epPoWGny9up
0Gxg7Tobkx/ZeFcmXto+Twq0xQVkPQORfUrY7ps2r/Kj9+fVbvzQeJHX633AhPZo
Q52tYae2hwsxqpvAUHiGy2r7/l5jU7HzQ2fMADklbPib2m9jm9e51hopAcyTQU8y
GRXC6BUZhAimHiRKqo+VcmALNvxdUjf9wcv3Z/yoE0xqa+RIiwkIEoMIQXH8d+EJ
lCVSB6xTfqUwZkeaUifRXa+82xLLFzykAYIDiQfAY2T9N+PhChEw4gs3sSUSK0dp
6S23bQRHd2pv2E2DOZMY5gSmcCF/sCJecwwlqingD2MZeDj9ayBmbrf2b9/pTVQf
AORLFXE5KGa1Ltq+QNjuzKZl4IxHX74pMbf8SSgI6OCTObvnXoHysxVXsvYu96QX
7sPyk2RPKyy+OVOOwGv1sFiAuCd8ZRA2EWMAyT1imZhqVZRS5bXDOfHX8mjY//fD
NvFwLZFjNZtFT27YiL/TWfp2IszxJghrxkmCffXdiguk5QhawbjF1psEW18nYBAB
VikvQg5Y9QMxqWRH+lWmD5swox10fUDhqlJ3vg8KckG9F6bLxdw77hRQzTlWuW7n
S4IH/Nnlm+uIQ9bMNeOTQiT6o876AGYEOAi1DL0DNsfC6sFSswlp5xcYLjfG6Zgj
ABn0yq0yzRlNZ5GZ4PPrhoAn4ksGGqcOPQr6iXcYe9vME55ThknnlmoAARxpnYEU
Y7GgFIKvaTDsu9VxSZtqclk58mGVZgYRb9FZsaUwMw7j1wstcmwSuZVbuh9vMJ2O
uEOp4RSL1J3Zd90uDKcX432Jd7/vF0U5ntfiMmDHoUva/6lKQjMThm5y1m+FPKpp
bXUiqCChtJccbcXjaR/B2nimvG90dDqmTy462wP72msOH9q0x4CEzX3Rjg+A1kTE
OHqJdpcvYyUsG5Y07XvM43vrqiqR1tETayRK1yGEtFaYAuB9lXKnnHeDu86Oq75J
/lHx0qB6AZyDl/Ve19hFn1y82SoWN6N8VeQnaO6EgfgjbVPJgREb5c+7VXhrP67F
r9FVs5M9EyGnU27ebprbKtofwRO0yfE0cSe/E/UWWI8D5YPng0g8E6FwL9J7m6YE
jL5rVRgKK6NaAnoJeqztpoJx+5ZAFNgkjLAW3yh6gpRQ1Lc0J9QYIljW2aCvJvia
T2ck5ufLNs4Fj81s8CKHVMy4lngziDV6x7HqZQyWuD/iPRwyAVeA3s+0VzWyaurg
kivthGMGcreqGqg7YoVyrG/1Fk3uFPd9mlNuhOKUt573y9xvhFqZH8EJ+xVN+TwD
vXg8ZWNYkeVU7Ur2ykNG2QKhIxnYN4dvaJc2lBeGL4M2opfHtRmc6QCTTzQ9iQzD
k1H301DitB8xVwnH0NZEZNtJCXZPIW8tv6ZVMBCBaMiNKzZkWwyye+CO2Z+IjPjQ
bbX/URJ9dQ17P7756dMihCyNUUsj7qpm6uMFahrXL60d8pp6sJbzBnJneA7V+wl5
Wf6+GKF8bDWgLh4hxUEtE2kVDqJVlqboR7Ahtzic56andzC5Kv32EL6T7yK1R8qy
IzB9OXr+j23s+ylBU7EkJ9xc+Q9XxBodREJXOTe7cnjggfDw0EKY8hdOd/hDpB7Z
i8J6E3TLkCdptT/foWxChXmNoljpE3aF5QSZKaZ7HEaPe1oxn8mTWo+rBSl4vmKs
/1Lgdd19uLAaTvwZbWKcv5rnsdf9gd2Qgi8gPVvo1rAdghJlGu5awybYcz2fcvC6
Bd1amA4btLA6OPaJCVtVBJURFzdSwMPRhOWjSAB/BsmLHkpGKJIMEYJgQx0oFfzb
wH60U+2eIDrSj1T5pMe+FMyRHtPVlv2KHYg96Emxod0KHBkoaBphCyb20qlajuXh
UHGXfEGqE9sVekcSwx4qt9c5lbGwRhQ/mSDc03GveAST2lKvemOThk6e51/JkvN4
3XkLh4Dy1X8Tr6/XRucJblLJGN5jlniEytdIyCCTJ23yJ98U5YXmhQrkrBD7Lmy3
/5vEpySbmMMOXRJbB0T68CZGD4w4W+F914kjdAQJNNIdLURCApVQbXmopoP1nxvA
A7K74IvWyi+Ag6h/8M3XlQ==
`protect END_PROTECTED
