`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
d9LYooQlvBk3dVWXdJbxgSxDyTJtAr+TOG7tergX9P713BaUr9fo3lhymSz3LK/N
iaAtkdXsnSXOHaFMU8TOkX2xKqaUsLk0R69usVMW5ZvS5UO9yVwFiIhYyyl6ZWSv
xbNnXqOP0FE4yoY9V1xtT7Epu0REbjNhwBgRzd8XR7q6zQayXTemgzAWGCHOK2OX
YfMskYlpJeBIQ6LWXNeDgZVzh4FBpPTXWZ7suu81UvYNMwx3/o5dQ3yM05eoi9+9
Ydzw2lTWNpHYzRCdDDNDjaH6gE8A847uZK/+EdrfjkHg/X6eAy8vVM94BuM7NsJ4
8HVxmWGUT3ipJ53yoHdx8DCXmvvPEGrJnv5ZD88vNskDr/Fj8Jymb1rwNPZmyqZ1
1honIStnV8LnMpNjOS0G89rZnq8GRzLnMIEi5moYpCUrrPm5yBAB3TjZbDtXi2pY
nJ6yyCA6mg/rdJ4dkRX5mu0KG8IabkD3nSpsq8I2UMHWFQDyjRh6wJxz4wDeki0a
074/yyvJ7qoZv7z2aljIhd3/veMHBzGnPm1xbEdr+w0=
`protect END_PROTECTED
