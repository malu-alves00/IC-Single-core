`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
S3yx1Q28CqJbppcJ5dXtMmLTncHYKIjUJIpFECtwdjeBUeM99AdOFTye36vwU3n6
dFo2R2snTdnw254H7mXuHgKqbOXC2hltwTAJg6O0doSVToCCI8gzvrL5Ue+m20XS
b/iP7y8mycOfPhkjZ/nD9BnQxtQ7/zxoUNozxv9FH/RGLSorhIO1xVlSw/LhXraF
cHCtEXh8T7Rgb+tIP658WQZg/KdRk9EQcV8XidTidNiv4aViFzVFs3350JrRT3KK
Ns3fEcDml5q/VPXDDG1YxFOYOIU2hpycYRHp9H/ISNYjidK1NqaEMD/+lTbNoR6P
hIcOoFTmxHvb8RDrIq9bn5N41lMhvj0ynItZ2brElvd4nk9w/cRQOPktNjWbQlpR
GdxCpgO8p6MvPSDqED39RU6xS9+yHg20S2kJlCr8kYX1ldMLgHZdH4kJRCsgtUMe
viie2cjIIoqnHI+X6KoEFj2OIxxz4Nn2HknNk9yimekhMoYpz0U6+rkjWcAgnh6j
AZp10Zks6tatYjyAxH+Y5DTi269E+QIOdpQT4AbKtvPDcAVp2Y+5KpOneFeAGUsa
TKNBZj2zJO61Tkbu/vtDArYImwu58ohN9Y3yfR5GHfMfgH1jG1/rwWhboSiey6dm
je0TVjINaMdxDOVxzQvk2wFEUPpwGMUgcF3GjIyICIoKv2LwYMCcgmWQslUN/PQG
o01fImG3TrNeop+R5043eBaH4ht4CylWNLLn56f/SeQoAbGKjVeCF9+R/TLmLwH1
kx++oFABLPyCCZsgVDK7zDLh9UPQ5E9qr2sP9/C/guJBw7+VEBApali3RvCdk/TL
Z7hs37JfiuERbZ5CGXS0PFOV4b8aGQPnA163vP7OcqlYYaqPjfo6tCl0o6c8wNoY
75+YtrAKXpVIn0JKbMFYpiqp9Qw16CkSLDYHAv908r8UzJJ2lKT7OBOQguWhWAv5
eJl13vs9LN38e+GfqBNWBEJm0ohzvyw+IATjVtnKZ9bA7PrHkCwwmM959QEYZgQa
/cERwA+bdXHz5l3HhtLAcCEd/cOncrznn2x7CN6u96orOzbhFQk6rGyr9AN3RzF6
HHs55u3ukZQuhHMa3tTlQj/i4QDwuTM79nL7hnljY/cfEw6gD8jeP1+SoHhJM46X
RqR4cVy/ieONfCtt/SIyfijYy9LQVZLVfgKE0RkKHp08gz4gYcFBeXyoP6xUbVV6
uzCYVK7fVK9lBCTaisSG0QrUY3fINMZbRDSX+aHnwvOTdmJOKdTMPIOGG1BgK218
mT99dwt+YkhO5PqoMW+C2i2yXmvCuPDSM51baGz8sEjNqo64KZPryrb+dzWDu3sP
dH+e+hUuxmSJm7Z8LvZ3/XGAc563QAv8MyuQTJVMzQXHkQuJI0wkTw6cyzmqlefJ
TH9GzbytTmzwg8cM5fxtRwMO5m1Dn284WrQnzgAeBE6C+YMEn5Arz2+AMW2kZwAo
ff/8G9e5ll7IYAXdEMjkFd7XlIDlcqJzp6rjTpA90HdA7PnS0/DijeupU7BdAru/
ZqQ+/M+2+gVJWjSKyAXXZX3xUlCk3ytD0yKLXTDLLjM9MMLWdHHxeorq1TGblHYR
LJuRUpet4Ap0e3ioRD8/aKtp7mhEH2CysG229xrJLD7gZASm4Oiiu383Gr0wRwj9
7n9DpsU42Ea0EyD24L/JHmzQ17+uUg68IlfFxT4DIXeWMpt61VtWlL/9HTgZt6yx
O4EOCetfoFBA7M7M2TCPUs9IE6kRf0swqq+gEXFHeX8PB5GoW2JK1oafMCJkU0zQ
ARxViOrFgm+HW3gogfBR6VQUeJuWLLvcHUhj86xJRLgiWlAxFJRmJcfuqU1lYmJG
kZcMPnmKGo0jhGMquIRKuObJiEfenn+oX1OkOZHhSO7oBaP79sG86uY+PMuopn/J
Rjpw0ehXXQdCrm+RzGzair6ZP3PAU/vHVXal1UQEeGy2f3cx9XtgSl8Msmlrbfx9
wft4+tCJtyRV4zhE04byMazh4BRickOUgNvl/TUOCQrG17s7o8l4ILlTNYqNekrk
B7H7MaCmujEQfgbA7NR+ahBpmpE6UsBD5abB/9wBLeGwrXvnI5bcGBngq6n2Vm8n
ro8yxkojlIQoy7Kfz8I7nLlOcv1uNDofnPtXtENxGDUf4HJ2ZTkCUycI66rbMdb/
7pnmP/BlELiFc5oQlKbTOspJmRcNYX18X9Kt3wJBeuKFEzxdD9vS5xXkz5MWNNuC
Xqzb5A4UyssZjzg8nrFUi08DBuElWM+u/wxGcALuosDZjsmdQ/OeUoITC9ZZxx74
oZ+xZhE7Tc4bnH0Rj5q6NNVGUYPONuwgAiZC3KxkiW2UHnzNxu5+JXNcOljRyS1S
YHzyte26e1mi+sDvluHfFXaRtxjsJc7hzWSbuudivODWLGXJVrracMv+Cmrz9oly
AjRKrcFETIQd/K76o98UPBveTtXYDUnSJhobLMtEkN0gs01QzTP5PhKK2o4PRUtH
vs24wV6BVhVBUNlS5ErC/JWX4o8GguM2DSdXWdMah0/c5OLhqsLHx06eo+Uq9EtS
PNAnxTFtC+iZTg/JTnXRVVQXEnfIIlOlJiZYSoJITnc6wZ0b8yyxDCby+1oiQL4g
Y14q7KSEsGLWn6P6afngrg==
`protect END_PROTECTED
