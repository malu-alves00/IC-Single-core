`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
adjU40QQiRXndMzeUna2TKRJMlZFMpO+sWbIhePX71uypcy/P9ejQkUG+twC5osx
TFE8FYpPrhlCWgMKeoV6yQzzDlUuQXaOEyTljHeSGlqmkvyGev/uTaWTABP/o9BV
bclgoDBT3LkLo184zKpQ8X/Z/UoWAY2bt6nMNsaLilUnavJGeSiztfo54djTNCcu
/rJAstl+Ms6eDElSuX8OXQasZrUwOT3x99wKh7Vkj97+mXYrwBCyZrIoTEQL7Bk7
xfJfTrCA29QPOTGcvsbBDz/objk8ISE8FCvf1ssfXm+FA83/OXLExsImILXuGApn
zeQSGYwV3uxDy4j5qtNM470B6YctZmi1hyF/pwyTP/kIST0rVmLeQac+fLJc+yyy
u2QsFjXo9W0rtigLYrtpioACSv6Wou+wHhR+ejPrDCbz4OEWIgWIb2CgUMyrfTzC
9CyGWwHeVm3BmX8MUK+tmeUM9YANoIAv/tRHFmA6uMrNSbq/wxa/C07FiprB61MM
TLiftL2usq8TlolCAnpiRsC177L/HzoVhbcvNwcxmhXx0/jSrjSxVt3IaCFqyVVY
GDxmV72r5kmeXnfUXJ4nNjt5Vt1ws688Guc0kZt7iL8PqSbxO+fvb4ntf5dpHuC+
/dWHYLJn+M6efmzyfaZRA8ARec09K4XvQ4ezbH1p3fLmjJk96R/mrqBb35x7QyuV
UMGCobGQlI1firq7T4PaiQFQlgXbFRdYnSOKuUKx09QNf3Ip5P3XaJetuAZ7n3qU
ONTAhJulkANIJjv0ENNPwJucHZuNl04GOaq0Sk5yqUvDykCMmKJ0W7t4MtMHPkCh
Z/eP++VC80ycC0QcKqCzTYEMMqr5xTOHD0IdDQmIg7D9snRa/EUZWpPPz07uSxiG
1mJAKnpXkaxcDliRP+9HF23khgM2YH2HYXEM8smySm4OKeqgnczcrughQld4iSaA
wtispmr/3mbrf55FHScm/5Zm5ADYnUqf993ZS/uOnPDQ/roCHmFQGCMONbm0u201
R98Nb01ISB4QHdiBftVGf0A9zvETQTyV94v1hT7kAtE6990Qy9SHeFSoGwkH68r1
Ia727mhAaf6ipdkGARZV7fcFBk24RlL4qpM4+Z1pFccneTjYQaaNxBHrZ6LKKjm5
Y6byAHxmwCrf84WJNDnuFqwsgdg8e5SesKZTtJSFhorxDE7g8leIK83q9zUxWzdV
r9iLRFT73AJYAqQiVPweF6+EwD3ZC5JPeiODcbYm24sazEe4ume40o0u8oKbHuXs
INaOrix363+QT+zqVYi4PQnOVS/C9loMKQKt/yv8u05+RSsGHKk25kvKAZUjfmxY
NPqzB0hX0i5Pyo8XKOtzULBqErSX53ZCuoGoYbb5+OYXX8sP1zWGPC36ShdDhXdC
Jem1Z93tGL49d137cMdQ65RR1MIQ6vPZvhgd4C1nfIadEFLV9pY+S+0hPw7bBCvY
dChOXoKiNVhBwpsgaM687181poMsHjj3yexfHlNUEO4=
`protect END_PROTECTED
