`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DtsEfWLKX9fu/fO9MbGW2pItm9cxXl1Fjalq+cv+JAOBVKGgeSJHSCQkh0i0s7V4
WYg9dy+GMUm/1eVyRNH8baS72iTfzwW2/mLtKxCsa38biOWvED0IwQO5qYDkcnkk
zLHtVCNmOG6UpJeu8GJtJiwBrjbMnTcoQ/SqDdeLPTsrUPWEkskdIttGoRk/EBlb
IRlt02nUGU6cvcJ+WKt6IlVUadM23H6pgKfdTx7IWMN/bESk3IH0viClMSlY/4Eh
NUAQ6xrW82qAiEHENRUiKIaytPWoTT9ehADDYQjFWLSc26A6RKJDdrCeynr3G34Y
057hvZn35SjhJodYx8oQIzrC1x1aYNHXNNSNiuzCK9fmgc3smiurP/geSDFbhR/s
CAEKqzASyzd7uUEc46s4hdpCjbVrNRts9qXQThE7vKAgkUJPoC6+9iyHlkfwm/MC
mByBJUkMako6h7ukm9hkZz7YcXvdHXdtCr6le/3IoxS/Awua+ZVF9gR63PYId1rk
fIKtknbhvxjSXsYD9kEN3qhPQ+Y6CCcumZGdGFX/pwxH3UG1Jey1vk5WYmekIjga
bobYVi8T7m+7NbxFvLapRo62sjcbTkgTsYmOnvo/o2E/e7HFsizboEKWT2KnF1Sc
MdWqJZoIIdFbjzguWKMGbXU9QVcpajiX2rsRaKLmDlv25x/AWSCqhPu9gYlEKyl3
`protect END_PROTECTED
