`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EqbKz5Ws9X8osWfdJ/hTzZ+vFU2lfATmuBR/LbRdetLlBvNwUQUgu4PdvmI9DFd2
ShYHYfx9Z/1C8SvajyXD24HUXLbxYt2UyPH76R7YOcXqMNJADybL7NCJr1K7WzLg
/VjTkhgg2wtWEzQzmNqwTv79c3+xQneLSNw2W/1kySghZ/1vtIJUcv9fw9Z8GNYu
ur7Ssc8GcRIRxdKM/thkPDpjxOSYqVy/iK4Y0Rajfd997iYouql7kpbajig0zTSd
xzUx+GRxfWp6Pgm396gPfzUrvij1KlvG22uhjVilmseDPS8MeJ+sa3EZxBo1FXWm
Gsw4NSoeS5nYiDHe/Asq3PsY7lS5aR301PSCN5RQlzxfs3DzBu3QJv1eWZl3lIxJ
faEwTe9yQMLUSIOeRebxUYvd4IIR2csCgHI5gKWttvOtI9c9Y3jHTVtvmLfKAfF4
0OUyKHAyAbQzEllbfrhXvsMwMAughyJ6hggMii4N+R6qGLuXotARXtr/DHbpgmRi
0OkVDFUS0JxwJTaC6pyZ6/cSC5RqKM5tQZLXEIPzoQaSG5g9L4aHjSHWPyI0H6/P
gMju0Afm8RSYtIMWaDF5CYIKxHmLp0FpT8TModkUTivtqdSUR7LPPHgbfble01jJ
Pr2lhJX2RSNyWnP1nQDfPpijQOqV9qwwKukm5m5meUhybBnsLRrKVZTQxK5PYdMt
Oflpf51rXPPmGg8qbHa+hHI73EnPTv5I9HULGHLfeM+Z2OqXL5+DybotGL4umaF6
AJxUuPir8+OKgsbKz5D15c7X8krCiYlBxfrhstLQ6iM=
`protect END_PROTECTED
