`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3hSrv79z0sNdwiB2jLA9/3S4Zc0uk9SHuREFYx+SbSUVy2K3t7b1IngQpn7SD1gH
RaLSGRHAuzlGw0+2uWBbKP0qoLnD5qOrGUttOH/5iYkuNJzEOf5LpWdztOIts4Q+
6xOfNs+xsjsdQvF1PzvIE4RcuqxqMd0pcTd6H6KQcnQAbr0CbmoWNxuqKGq3tkI6
earcyaJkLB178t8yZDcgTw2BV1kWmSkvWV6a3D00A2imk47J8ar0CsFKtIwDW2ID
r7+AkjHwrY5LZ8bxE7ylid2DVNsfNJHDoVEz3YNtOQ7ss59ivEbyOQX3E/zi0AL2
O5l54Na+x5WClExlaPhUAINGROVl+T9s0SMzJ12vqEC1oOhliKh/aWRYqgzlVeGQ
MDFTSlCV9wecMMujnUpKzW3RcC4jIeoxgjMTfzynICCUHpSsw9Ss2NFdDhH5F8Wg
QjqneuHQHwTm4jl/ihQlYIclyCZwmXi9yIHa+ER53/LXbmJeZS2REhd8ix5CFpvw
64bUvJ79PLYSTEenyG59fnkcUkfPCep4GFRUJ/aRKW6acQ9Q903ziP4ElrMZGhqX
G1UXGxYghavzTjkU1FhVcbLlBU+WbeHwHmGzO+E6FIxthMg6Omagbw3HIzMG5QbB
sBRQhNYVDhU5nwkKXJ4jRUCXM89W9AdAX62R3dZ4PFIIIfq4U339UjMmQNB/hYW9
0R14OYDnUfbYnbh8mPDxVkkYfyXMkZcRHmPdau5SNl8cVy0FlJvjGSyEx+DXUkXU
ww9zv+wuN5v/NIStuW9HvGye3HooLzW+xzx/4rtkva9mUmrt+jb5pSDpjPZpDU4W
vmV83Pl3M8vQT1/l+NWKDCzYkQRPBjG27zwEJEXK1YSICAgvz8NeOSeaAfQ1W0OU
KKYlnr8CwzU5DyZ8xpGhHUQRBfYCNUllHhpe1SMpH9POKLdv/QnJ8lbdAE95DP1b
l5mrOcxcU8diNsJFRTHQHHPt/iLhithUyv4+xIv0SKBL/tPWULGwGEXrm4xG1NhA
fEZVDLFSvxI2vRfao4VLgiXu13yQYz8UwkqVUsYzleGFH1lEDYkk0His0E9ew5kx
hgWiuzvsZlNl53qUijWj4hYtxJ4/IVe+EtQjAp8udKWefp3X+tSAh+Vqrfr/dsMY
8SzXg1JmKohJA2E7UepoTXbTWbHdkbes3tb9FdbNzVby78v7qN6IvHJ2xSvB8GYn
NnzTmSjED4ekK6iSDbEk7NDIF+qwc0BZlhLWsA1uUBOTnf1XaMysZMy98dH6vkVM
G1oWD3aRyEq3xWzV2pM/hiA5SeH6D8qQ3U95mcJ1qHm6E4glLfxD4bu2Dqf3yoB1
Tlk4vlM+eC0aPkBZdm0P0M+32ybVkDMQOnfNXF8KrzKrX7rxZxXRJ5X74Uvekcm+
Vs22BRRCt24JqTTEtU71jzoca5LWLWPSKc5FyCF3Nts=
`protect END_PROTECTED
