`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XIy3yubRxBpvZpn3c23Rj3QQdYyV21v1stHWJ2SWcAzX5xJHvuvn8vbb2whseK57
Qge4FsaQd12o1h1Sni6RCFUc/aioKv4+MRdvcPl97sRCr90hhE1qtS6H032CTs/L
Jcks9g5y2TPag3kMvUnjDFNKbi7zNih0lOJWiltzN2NQyW3La4yoy9mj+fqR7jq8
wpPXnc4ByBgOGyrUIbVJK6kT+puC+fb1NLwAU4lWvzM1a3cJcoZDjys4s+he/vwc
yQP+EJrJmMT64u4Dl+mFwvcUYCbMGbjCxUKwl8knV394DT34MRIDMOg00NBmltaY
BdEFKbhE+AUg3L9tCRikxig0Pm69w3RhvI0bsdkgIbFtxC6jm5+Zxch3fiBapxjY
yoP+kmtT10TRwv9GjgLx99Dr9YyDGwLkEwkbHQ/+AET/o1u8ZRf0eatwkTRNvZEt
1b3dmdYBzFJcQ+4O1dqUlHBWE00RBasroKJqHdqp5imT3UAZxc9h9tQWcPlKjzbM
g6RYCEvT4JKlFs4XeRvqYfMaYAtdtkND9xVxky3j8XAH4c72Byb/RXMSXlTAzT9q
qITZudFot/nJppbMGki7DSFcqPbCQhD+oyhILH/cV2zPP3TLtnh0meWAYnD5lvtr
Qi0y2YkIRDSfIsQrzePzdq2MKApASPdoKlYAnJ+FL7di5Ujm1IZ+2tkSleFFnkQM
r0EM+gcr0SminhCHuI400qRUjVWQE5vY6yMKb9zEJju5KDBIA9xNjdWF18Sh7gJX
EIFJqcdPcRFBJta6gvMFpkHWtu1ED9vcoOY2h2lUZwXEWcqcBFyvPmKOWFkjolq3
iy86B8OMP0/kyHfS3UB0eUlObDOseA8eQnT8CFfTE+Q2c9TLyYd1VujTsp4ngJRJ
S2aCyr/pqcx1Rkr90be71rZhOso6HcU7iHjJxS51k5/Q1qx3lNQmf3QJbwafULfc
it1Uh/05pwXOmZgHrt3kdD9DmJrUxhYn/dtTRx2CLqR3YRHUodeb1ltKuP08e4Jq
PpbZuFiQo5g098qySee3qkm8RxEkxYoA1yfseKygnL9B9XPu0DRCRQ0/VXxx5Vdj
Oud5VGjQ4V5r9xKRNaNM5cBu9FBjRFHd/5ygFYTissGWzzksZLscenAm12U1QIJx
HOeqO5Jk4IXSA++l/PASr4cgpV388ul6KL4PO5lcQAVKHG6i3zXSCtYs4trK8dka
cpOTsHs/Zrlo/QnJVhjPewJ3xErNQ01P9f7dCyc6X8nKpfCq4inKOgYfmGigSPo9
esvtazm9EyMHpLkjNxF+szSNhTgLHlS1OqWbsQY4X1yltkMR7E5x/eTggPwhyWoI
MB8i7Us+o41z5HtJ0abXT8B84cEznlpcmherJlActfU=
`protect END_PROTECTED
