`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2lV5GhgYndPdqeKmDNZkVl5k7UYAD0myxHNYpJMMePC+AjnHL4A8jFJtfITvrKfI
gT5/R04fAVQtinAPcy+XmNRtxp01XACLFc79KlU/z1y5Ev3fOR0KEr1iW+I51LsL
FxIyglKgPXN254npTwUAWz8ukWAuHfqbxR8ULV5xr15zr5oEy7gbBSzNhRhZV59P
6EX953dPnZ6PhgrQhTIFkh/7PKH0LN5MNbWZ8GFPkKRdQgO+hOEx8mFKkO2rhtpf
kAnIGuHrgLl0rXo1Rxx9VEcf3LSRJLq2iqCbDFjiC0HypyM3M9ZAhc4iDWQ1d0Xc
BGfkucpYrSIVIeC8hMC5SyAMNDJ8IHa4eiHoV7eiVRcY9+XL2xkJIi9Rod6Mvxjm
aMiXImEnW1L58okR9T8DafsMDWBQ5DyZh0yJYDUUJrtV1TGMSjKm+LFYAhTGeNja
jBRgB11fLVtyvuUUzZh+7ROxNDLq5S4JvbE3C/89V6ZN+1OwgVQV5MhLODnuGL9X
GbvIEC8kzpjacZz7I8VrZsWUhca/GCc7FsTAedbCb3S+s1yX5FMZeGyTwuqM9ZGO
zMV0a5ljYdaICNwRK49GBhyDjY12EzWxWTkNWt14MGvMti5n3fYMka0Mb5nVtXgD
+Wb4Q5l3LAvtOU431qb2oBXJfqP7/sehqkRyPxRfoHw02BnjHOZBP0ABHNNDrfyI
nPHbrAnK6oTYR6NNmw5+QVppOdlVT7y4FQz+pbRtDi53ysk2XEIFgwqZYytv3Iyi
Nm6FHHo9AZbSHHfgDoIjetFMPu+TESwsNmefEWnXRmOA0nejnaYCfvgSdrRTWpv0
E0Vg7ycPkPt3XbMAm10jaxKGtfhTw3UsoHAZNxnNttMd+teVUcQBZxTCNDhCpGgK
wIiU6LlEFtne+K3GxxbxyskCPRxgDjs/XitMxN2qKFAdMpoWxOWIpOCqU5SYW2iG
w4lZZo2nL2iSuTXjn7hXNKs8ibs/NuoZ7tNJmZobYNXjHQQJ4tLiVYdbd/U7R5uv
zP+otmDdnkN+ZbAcfXHwsQ==
`protect END_PROTECTED
