`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Z4RpDNB+hNTIhH4Kn84N7hTfpPqsg9cJy/zSgYDZVnB3YrcajJ5JETHRpuU+ERgp
2qhSgDVdLeFncTPuhxfpDphS4skGslX0pSfezirlWYjmNk9h7OhSdrWLITXmoJnT
VLssvO6PJNxHrm0w7XYGCi34TwZH9nW7eEjnqt+Q3QqnN33ivheZcwXBv8wKA7sL
dCqA/swCfqHLFRGxMXfw7QDBk2kzmtLH1GMghUjsqjQ8+fT11c79jc9JI7v02Z1s
CEk+qxjx+BnzjP/wII9SVTRkMA9A/HqdVGBoQavwdxBB+VzEzl//huCnu1rfQBW5
s0nKqgEPLs2Y4KX0llyMSDq33LDCWHJ1Le7g2oe//wvaF5oRYQqs4XTYHtQyjfz3
nfpFKGD68dbNOH+ga3sfmiEfhtkWSPi7fUJcMPwMXG7xV0eqtNBilJOqm1sycKy0
ygVTTzS6BLeAZSvabciXLtSYqAKwwNXWEzbTUQo9e51qghDoYbf3aF17fsK+9MQI
0EeTgcTKAtSOuEeb1JmWgp8DuMDshIk4niyIp6fhVt2a5mPx4GETJTZ9EzQlo7Hw
SPkFoXWhPjpNKSzOypyJKqt9/4xS6huyjfVbVXK31u6z+pJI4Gknb9feN07f5spc
7vgqgiyg9nZPmrg+Z0okN7DzdEUyAErz2VM6oMgAvj2jcqRcTz2gVcs5j9uVyM3u
Bgypfzbw+KXzCB6d9YyCKl8oEWZOk9QSwh00nlFv6oiFQue/BtRo/DvuLza7i4Ee
OirCgpKg/KlAKWHL1eg8r2QIO/r+IdPxsVEnoEOJAR85lkRk6gDBTJKU0CVbsg1Z
BqGcdPnNyHHUl4KnMWfLXExarPJBQBqdbi0eyDmkgBS5ZdqdmhgrMnKhrhb7Lood
gQtVBmcTHpGeTVii3tIe8Bivgqku0ZX9t1T8dk/oAAUctroKf/YE7PkoxEkIG5IS
3sXd9ytrjLzQRmj0Vac/BKR3B7p9d27hWU1yvwJu73A0tu+FYstaNV0ZOolgNJmH
3St/P3bueEp9fbZZOWKviceRloQ6qSlwtfnFQfIYIU7OhKBCSpSm5+ZpNJgC5x5o
1mt4cA5mNXeIwpbIdlOY0Iga6gJXvux//F2w7w2rPujo2DUemPUqB0uE/mlrJTg9
61ReUtFlP/E7pTwDWHjDk2q/8YBj6oYD+uzKSLAX9o2v2JvxyFEJ4NTQ7XtEnLZ7
4aEPbekDdDXLh7XtrgDePfBhefZSTul8FvuGeho9vKedTSesx25gSJAlr9XBX2Ph
7jWop8a7k85hvQE4XveHd7wD4Ja7J34Sr8cI2t5KqSB2KWynJiMUesIbnStYwAcm
znujWQjf1ugwJMPX+jCrTL2K4lR0LhaWXOzBpwCG8+Q6jNstknPWxFfNcz2fR3PA
//YVCUHhOy45bHlvqwtXXVnN7YifFFwin8emlieQJCMMIo5zWV2xnVUADHcII9yZ
3lE4qLvPQj7T39yYx+or7yqb0gqoRclW7g2ywJ9rT5S9GfxG/H7lZsYoI10d2I0B
sFvT6isAazbF/Cvk2Uv9bGvKGZEzDD/gB05Oe4+oLpHMC7dw/0YdcUFIaRRrA3QJ
`protect END_PROTECTED
