`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kpygmRdYyglxAUtSUi2j+tS3sGv+uxIB+ug/rQaGbraCggv/nv10hqYBn7bsI93r
evqbR/6BOT7WhMM6jhYzD5+esGGBE5CJ7ArGBO3HcVPSmhi4TkPT+WqAi54r9NqJ
A2/rP59y1tZwf7p1RxetDJP6BGSt3qk5MXsOk2S2hABN/GDN3BbU1dQ1yvcX2Dod
wR4gCOOSCo/+06sx4zThmi9CF2EmRwytUHZWG0iFez2Q4AT/0aSkN/wwYuTTGKx2
qsAUaL6+CzGJI368AteymIlwusI5Rz7t/nnFTQBVeA/ecXl2TN6ZeCoqvwL/KVvi
XZfsD++fRX4wvzTjNB3ZkPQreJm/89uz689BVcOE/lBFtJVPMKIhm+FtEmex/Nic
Vl3hc63HmMyWJV329mfO+TVvjwbKFr7YSXJdzjSoleF/kTAPNIaeJDTFglyP4Xcn
UVL2uP3a2dMuVOGStqbZa1cBwf707FVfyaI4cBx95vSvkSf/D7vhp4y4lqAorkoo
X6HMK2a8UZsUbEp9q76uQaXyX7zYYBBq6UvC+N5ZsiJanyhZWqf+yV7AfmWOCeXs
evfCJfIEjeL6L9xwWLJi6fYWzKYrlOoGp8vTlVHf30XGLqGg9/MODFrA5n+qjqch
iINbQNQyVGDo5ERMgBmqThnAdb02wlnQNWduF3ZpZbWSC3jekpSIZ6mWauiNPn5s
77FFKu9VnFDpE7vzaaxsITXJDA/beIxTEari1ZUW7i74RK7sPlDUCcxfw48spnsP
VVwPzXbILX8zxO4xMsdNCu8YvSF1m5iA16O6IuN8YhrsmtOX1YwV/zHRTGHaaF4p
`protect END_PROTECTED
