`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iT7b58XBQIdtebmXAyj6ZNXbaBv/cRzGs4FJkZ9TMQsZsCRa4O/VzPrVm/Yk/j+5
72rQFRpymzGDd6HtAgcZpJTddrP72CoDWB/Gc+39VUp6UE4iajNZdhy/9VGi0K0X
kSIGh1EYSOwcF6OsdUbMyPhhPPV1Bm4ds0Qwm1e+H0DFOD9k3Z9TC4wJ73YVxQXA
V/UMdJrwlgNhfKzB4Zc3sqtMYtITQqIWiTF6wRNXlqbd0gQPI6zVjL/KSIxUSobx
0NJ5FmageoA3ixF8RMPxrs5AEW/G0VfYATlJ98/x9iyfsU2oG3LxuFqWCMw7sxzL
GI/3+gMZ7ia6ycySBOoVOJ3EwqC6zjQG0BYMRf/VGvvkWoZUts5D1/8Rrs1lQBPK
Cf5YoEqOiysaEdRUIrYNaRAtqLxpBeVPn+8oKgm5NIZueboYe6nRHL8hoe1/y/Xz
oFpnIpeezrCoNLDQzBbvT/Im7PHe/zUTNzYuYiGIFSW0VThub4fkd1eGVUYrMX4V
pWbOT/nuYq0fiXz6l22Aembo4A0TqYWWb3xZI6Cke4oN1Zcjqc1jgUjDRmD/bYF5
UQL8R81JMcvGTLXMYHQRj3svhXeaTbdTF1f2PnCYPHKpVYUCcH5LOcYGAtNjjYpz
3STY3BpcrkSquCQnNr1JeHSoT3tleE3KWNmHtXw8LTOEFQasR3l3TgL5e3HR/olg
bXJiEaqv5IYobdqkF/ZM3oiQ0A1bLYloeHGpPzxFvXLhJ+CuwP4/DU5Y+Edbrgj3
iAQ6Ueklh6iL/fgPP7EJ8Ypz+gqGzOYsREgHIfBIEkw=
`protect END_PROTECTED
