`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
POROf2cxcqFeg1fwy1pJFNkea3eXn2JlNsoaIN2XeEh2LY0wkiBLrrvvBuqcwYW4
pKpkYy3KmFrfAU9eExTjAWOH1ZT/gYaqFoNZ88bhwmCoUE3DvHh8XQRBxp7H6EIu
pxj55Vx+bmGVy9/b83lO3vUXNNCsbCwWXkRQ0eoTW3KuCQHMg+ekzh22j4yAugoJ
qkqdwb5MBZ8E/SsMaEYQmGwj6bIInSBOYcjyk9bCF6kFOQWijtBUKjMdxnSIFTUU
/dyctigk4vnoQUP94/d4z4fQ7mFOI1IbZgSmsLcCwgGf/dVQry+P2FLIbyPmcsEZ
9eHADZ+X0TpW911XBG0Xh5dFyjXjEK2ewKsuLoE62Jn2Jc4uqH6WWijHEvgy9ugB
vk9aw+nJlITwVTsw/DofY1MCrOa4cyi2KuHW9NMBP6K9v1PG3pqBQ2fvxrtH1At1
vDx/nnvuhVXqSMr4i2sgh0cZLVf9knrs63AW/7Ek8UbdACPPt5YQOqZTaPG5tbsz
JGK/deY47LNrLfGvMgSRaX5vQpZwMa7vULIhK4R4hZiVU+/75WK610t/vmW1NwX4
7p5LKtP+VfeoRCfrEGXScPYZhVhCIBxcBOtGYj2+miTr4IR9lRO0FQugADI0FRME
FpO2ypN1/bRljCmyuANkgfJhX4LipEgLadJRJgwHivSYCduFaOnP2LDGM/GOBVrm
Kk842XP9fWnADfg0tgv6Bf0bVlvMmq+VFGRXpW1rApOpA+qr/+xVO9CiKGZgPjKP
5Q99tqNGAFiHy9grWFan4kfIBie9Ly//Rwg32Kjq9LUXV7wcgvuj+nXA1biGcs6w
YMBoHJ8gNZ259OpdTaQwXE3lKhBv7JYvk/LYWxDeXVH0LJTJvTN8zUgEKXaEkr6n
rvoSyHYYVm3+OK4sQnR64exCbeqFfKtIuehFnAgQW1hJEslurYBj0ViETQfvxLL+
52GP2aVIxvFnuDd49fJTOSDSDpy+jED0k8XkSr+1Xv2X8WZACUrYX4fqBtR5bOlK
nehmjKzREDarBh0vjDNx5l7b1s0AmwlczRnft0hcl8YaI4ByeT07khCZAzrmYTbQ
iMpvc94lQURKwprPbsGEcaZK6jBgBuqnMgyl2WnWny3dm4LjpakmP/qYKll/tBiZ
VnJc1STIlDRUNPo5H1PJcZ9pvv3d6OQmR2KEaiIVyEZTGNnx5IYcSDgvwQ2hfaZt
sxbzI3x5Co17VgKtus9RsqgVy4892KnHiaIzm30yc0sBPoH8C7aIYx2bkgV8SzjE
knD1c2jrtyHCs00LTCCyxQ67sn1N/b0uzEi7d0lNJgwhsTvu9SprmQbpOQ0wzQwQ
4ZnvQHyTq4dGyCnKjQbgOIQHVDnQ/jQ8zI4UQTDc2hrjD7GzTf79VXTOPPkfK7x9
6WnoQ8pQri2/SYjmiSSTgtDA3t3mO8tKtbBcdz+e/1iDyq5XNHpMKUH7tPbjwvk/
KIGh5UMq6hFu6KTBa3DfOvJNc/XiuG0CHOWvcSDGGzckWAGkvc1x6iiqudlJtkVC
MzsnWB1qPNZN1SwZXFZXDCy2mVSPWeIYmpTWpmgdIGpbM0FyXJuLJpWbqni4NsUJ
6CcSu7LT82CzBFype64JuhvAlaCxrFvuUrhvzetKkA9B5tR9RWLdDeXEIlPqu4ro
0n6iLbvcrLVmGyW7WEJTWJUBz1ASoM4cpwXYWP6KmtiCwr6/i7Kc8svDHScEmQO3
L7ywjhbc6nI7aqJ87PsMoLv975IJs/YqBbZOv5c+geXszDjMpl+kIApgmeotcYAe
U3wm9nch5nU9ASozxb3ftclL1RuZVsCGrZKLFMNqdMgEiwtkvXqsAUqYL6m0bImJ
nhyeQzgqiQOiAWEQ9fwIfXAXMEqfHJHIzFSvJd5rce9VpW61wYdEPlku33Qb7C3d
OI79k+Df0t7+EZK14XM76cp3+F2vrVPTB+mzTo/WornQpaoULRBebjyCNRulBtn6
slLBeb1KhaqH0lZRAvcBKeba741bRyX1+YxUY2bhau44s90gvUYON5hyogOFnJ56
rxggBOauP75XAWGgoeEMETZYkGRJvHHBKh91SEniRoEGLw26Iu0UDrYFDCJdWrdF
1ykXFfqm5tS2ZS3xdpy7/VjX5dCjVxT2DWKHVjQyHoW9QsWNUbqr0lmgH7eUw6ag
OloCQt8FakKxn4wQSH0XJq6PICU5s31NihMpE8l0YfCMhzXQ7byUdlZ5b8pmvOPC
g79VzX5T717xqW7Ru6skO+BrQJXQZVcRr424NlNwC3FfwAUldp7I19Q0+IVXT9by
1oeUMayQYhyFm5z35TkJymBbBY30JN2yK01/bS+3lMfJooKLPxTkn3leaX25SpxZ
qYrpxrjwEIir5j7/9AsG4+JuwgzBhxugoiaZMwrRRu3UZthKqO4n2qQJuwJlrjKd
VtrhGigUGcSTwnkmBD7uWdHlpKN45hJf5vsyWQpZq93/KWrik0txjksezlYUaiOc
MyoPvYC8qKaTEC+fRT2JSp9+4sNMs4RaXztdMZ5C9b3lD5veaiw+oLdOm4/SQ3oN
qqbwT4+DbNvU2MVMODl8L32JVsNX/v/gpEu/ZD2dnM6HRQbiBfwB9AfZuhf1vpma
0yfGUK0pfB6fH07r4sDH4j4TiOjPs2Q1/qmee1R0o/CfP8YpCyd+Wu2fCrkoIbDe
E8zWzn4VHaGQ8Zov2AemLvdDM4O6UL1niuKXnzeUSJRp6/MOvV8N4pLVH3IPlSeY
3TDH9QctN7x2ApkV36BKOG+N4AWl8X/eg9yjSRZ04nMDCm53c+RzALYYu6GWtTCi
BZQOMt5VDE18bkraMq6sSS+ep//ExCZKOU+m5NCVrw0x5YtwYHuWj4EB11BYZNsl
Ixl2alPzZKjMMcLKeAh0Ea76K8HQ6AvXESwOch8ub65QImyMi7aZTqKHDcCIGKJE
WTMkFVxj3XJBvGJiOmvBXeY+JNEAcMVzoKxf2DDq6kH+kdGYEBkwmR1z66BjsaaE
iZkDp9P7YOuf9vSaIEQ0sjOilIJMIKtFi0ykgqT431d3IzTtDVtlTr8zOReW0/FK
H/FWf+6Ao98E42P7PsFYIXfwNOk9VoWB+DB1VcNztbgCgAriHu9GZTPjTwI8hxUH
VAtNfUMy6i3r5oA5EOH+HA47UycVEEMjfZCTXkRuxCOcz4XLEVXtqAUPwdOMQ/Z4
bFGH4xEdDL+jtK8+VnCB+phMSjH8BVWPFWUqvOZG1dxsAjFuqRd0lmrXqTQRG5YU
pl+A1+Pt7dMqqOxAFcAS6lCYHNOV/e/QM79CBEvP/iA=
`protect END_PROTECTED
