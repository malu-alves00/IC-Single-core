`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uiYyBzx78Sg4JLk0EV4NX0NFcyGJ0IdcfTllTDa/Ba+W6nEaHGIfwxOIXa9TGx52
/o9AqJ2x9NhfPDSGpH2mOL6/1AhHTsS0vOL/+/Cu8vNERCvaNtuc8SmQHZ2YrB28
0ypSSvbVtU8VQsIxQtLlYz4lTZM7Pgq2TjcSJIP4Hpw6KTP26+wFhzNb5fQeTyzM
IumGOzy2Hv57Gn6kCVNRtzHNEkV8+M8E1jhSVF5/0ESlgEa+c4M6pvaVq140ota5
W6OGLRhVjbhW8Sfhm5klbngoLlFJX8z541C2HB2bF0iyXd/KDVu/5xVTNwTz+3/N
N53IjOeM+5qjvywp3cYc3yS+mr3UeZ2y2W6luyIpAAachQ29fZgn4WFDTDCYkWuc
tfOCJE+cfRo8E4h9yOVABA==
`protect END_PROTECTED
