`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WpL7hP3MtDr3+5vUHuciqfjbozpUhAHz/PNm6bsypaTgyXUn3EHIvPLSYNRyQ2Zn
cy8GGt4Rb7y96eLblla/CymTCNoficG57O0JSGxESQ2aZ2ucc3masiHrijb+YL1X
C0iGli1ivSpfdu7+oYTwu6Nxyv8/Vy/vFglKG9sgf0Jx/zAe+E/phyaF7fvxIPiU
k7gg5DG2zDVE5BMYSqA62nN2SXfI/Sd5ic4/rROiD0WNsuejX5ChoGS2V+bLVfAq
DRt3FxbpRvJQOcLQ1ghnxVjHeMXX6NDSzqh7oYxit/9iC2lbglIdmbJvMMVm9vXj
yYMQetTz/ZCSXTcDCi9/diFefkYrj96wexNI0btCzTbsKnuKozcvfLTFvuXVVzB5
XHokf7uFQdb9pwmuKVcKBIawSLoaqSTVJe4TdfMtb1BC6yaHd2zVlIHGaT4TIU/9
+ZGkPExacOWufp9untlamqIQvwfzGN3BMUa+MdC9FBtBAXW0+3H8a0SHrHzGivV2
TaZXfoIo1IswL8jXpFgNzQn8zFXVCdLPlkocg9FN4kB3gzmqjV681KxDx79qDejP
7ZSu2k+GGrbh6jtGuwFqb4JBvecARHVChnATTBvhSwTxTY85+Z27ypIBik9/Akx4
pvK9ySoR1lQeiNJstnf8HoMFNJfw9n+q0us+xdIw1rTYgVSfpVJgaphmgeY9eqnK
j/1ZwegOjRSKHtNGaABK/VacG5C6lhFflvdGgj/cl/o7jyOR/SLll+ivqXU0bNJv
oALTwWdXPljW4xcZw56JcA==
`protect END_PROTECTED
