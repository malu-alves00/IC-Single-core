`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PUN/9xcwWTUCuLQHsGqBLmzSAL+Q4YDr9UHWF/xwlwHVjxgJaxBBizZc4jX5KcG8
blLQZn2k+hvCHA4v0wVnymh0gSjwsKAI9ffX+aOUDa4suoTkvKm5O6wgDWLkEhdG
MZI/8gSE1Q3VKDIEWfyQxOTvz73Y+igb80SbQTpI0UVIzWYCPIHC6agCODxeuYiV
CqTTyMsrgByQ42mhdoti6N2lU8etVwf4b/KVINM2peKdZ9xAK69nRJ8LdyiKK2uF
BAwpmmYXnJlmAGSYr2YBVCcSODixQ7eEbl3EMbTTF7QEDY5G+WNBIjwGUSYVNsUF
wZpPBTevcF+ca/tQCjANHVtebuwQZ3q9oYm1Maf73nd+MP74Z6sW3PvbcGDtqJsD
QolkoBLOUNlVDcno5Erj7z13Gt8BqsV5wNZy/OyhpMva9W9ClQfNBFFqU6Dg7PUd
KIbMSHz4CIme7Ts3fovcRqnOzVO+O07TCDxxdosQECoKhm1mPg664St/HrbCvenv
eaWX000YfWeVzjFFECAyaPsMR1R1C+3soGs3j8eSmOoQnTyPDB741Mi0AscG0glo
D9+8yBbX+yFQuHckwtFPcicXfwHpdlFgHjdiY0h5kDWz/0EAmWqh25NHWXiFZUZ9
HK8ytsJ73ujiTcX0cHeAWeVWM9jnxdCVTgX+fVJS6z5599Q1E/iGzpYKPJtu2slQ
8JN2xCXRyX+2SdBIANFY9kZSpwqXlPt2d+7LB5IfzNidkRkc/zwhrAWQDi8TlxBi
f1Cb12OTzqn9/B61YGwX80bRoJA/PBjHCbotPPFLMvs633gwRA98eY4zEic+JmnW
feRyw1sD0g91+27TY8O+bnpGaneos6ZIkVzXJZrGlWhdZGfttNFm8n50iLPXZOjZ
1jk4hXM8LvOAUH9/h5q+aYjIZ0mlr/Up936L+S9/NdtViDLZtwxtcAbHkD4Sny3Y
yoQmr/BU+lp4Q2xsxZ56Na9rcajN3U1ogKozF6uMg1dAZIIojkIS9u/Ajo1MbzVS
JPyJD9fh3zRbhhroFWR+90/uhWAoXGyOveQV50tXhFE73ULnm67i1AOi95akFTT3
sYmqETMVgiFowN2fs0eCmKLW5+SNX8GFEV+L+aMIVvGRhphP/Qmw202mFsv6UMab
WhZCDmtqfyi0Sy9E6evQE+Uo9xaFfZmNXZ8Bb4rRMy3clIdM0EBqUehs9VI/SqPO
JSB84dWg+33JsS9JDRzqDOIxlEv1p0/UZp8Dw2h02UrjBR0giwm8pZ2iAzbThPcY
xc/FcVOQv4ysnBPDv12smpNFC1D/wqG3iN3X0YSEsOy9IOHD9cOQDbJlYbe2i6XV
MWlFi8f/7f/5ocZqqxxHCLvLJmEpeUTmsbqvu5eUxdNKNGDnuT7z7HcCuGaN1SoE
eJqnO1durbGxe5AD0iUWprJSrgRyensrPs5Z161t38W+SO5AP81IzBKk4rF8efXi
lpbHUw+btBKDLIQYTZCcSOBPuoeMoYoknlC0YzI9Kn3BJrypu5DS6HGlqFL9dLlQ
En4mfokRRDwddG+FlGr15oPMcmnNOxAgsP25Z7P7b1PxZiTSjfukQ+1hIqee4QWb
n3KQYs5GgEr8bEb2I+QCLNf5nq7qcqvJ9Olj0lQa1wfANMdOd8gqE9weuKRRlCtM
+NeKQ05ZGbQvISqA1TZC+CwKAZGTQryC11TMlyzdPoXKXW47gOOoTYobnWbm2eaE
JtXe5qeSuCNDjbJ5bg5MEt/oejRxz2jAAI55W4R2SJDqZck9OvgX88EaiQuFNSJu
fvqvtA4+Wm+G6BG34Gv8v4kDUZHMJuoEHdboNdC3mqgzZWkxMGUiRDYSVNp2cFs8
a1ujGZZSHt8x3kNVN4zWeCmCfX4vlj1hcKh/dW2pSSPMQqIbiGlvpgJ6kbmLNSZ4
rDHWFjElurKIvyk3ahYCJ3PISpIhqCSviDN4FkUq8SGDHomrhtUUkwzXuDZxwb1+
cupY2g96lDuIq8wtljZqCSprO2RIf168dusRPlbIZZ5wT/f1cCyliz0nMHyQRnpv
1QejeNV74ioSMrjOjlYM8EFWqNmVfAQT2vRcRVgL+2OduttVrquHERGFHj2BQcKJ
GTGr2DVPMjfZrc88pNtqm2L3I3a5dx7OAek5qZWPu8/RhSkLsf1nUvEi7sx7JrFC
HPyOv6skFYCWVYJNJiytTWUtjIEITHQpohwmp0vVGEeifHXII5Iwh8kyuP5hC8fq
LDlVoadteE+IhWTujKc5KkLMJLulktUjZIEZTa4DQ5K2v2qH18Rv8apqlw63dPTY
ss0y7QoK2H/xeZ14BKd6S1qypRPVvsn4IUQjhS/3xEC4CBuDSa8mCPgrvBAvhKWp
65NLL/2koWVizWN5D8VKV3gAT3AUpAUTGUKiE7LZmQFEHQKcYWov399ZyFBbwR1R
QlbynBPT/gT/H7WS/lpysYHA7c3xwZmhzpwSGBeKP9Md4r3PIlDGGqEj11DVcbT0
8hFzQwQN4dJB9KNkziy2ZkxiGQuVn/sCIeNRpfXE53dvNGyt6UtHuB1umqxQ4nWP
vpSEMySomSPep11/aJW+Mkym9V9g2Axbm3WIGwPV0Cmmn25cLtKKXRrqG3POaZMx
KwA7LDxP40q8E/lrwNK0NWUofH0i1+eCJ6W6C9OHtR83qweQYE6eFi0tX//d/+2w
q8voV7lRQGHaQc32iAeNt5IHamP26FEIfDSJY3vH/ToLuWt0H7nl0DP27ixVMe7v
Jp4UTsbPma0H+OmH4whtZ5eqOuTgMxzeKPoHcPH6Wr+aabs+0DEMocL8cRU9n6GH
9jswwHyKl0NaaW0W4pz/mUK/df+ApGIsDe8M57v3NZKKvJYvJHwSg3RK/6Ym2KsC
PloolP9hwoLZfqVJSAk6FhejcagPqxpzTtRUqpAJG7gDBboO+ScKLlT0x771ETyM
0c7HCveP6YlPIJEUUQcA6Gi9IVjCTcWd5NwJZJixc7L6mBLCc48wYBjGpqIZgD6s
suY4RDpx0znsy5ZYkeBypdN9oEyZOEXgyJLqSPrVyZNylKyYvTu2Lop7YVvSOowJ
oqSJOToMzBcgf/td7+2KrgDXL2sN2Kmq7fIyPEBcRPailn4dSUPtpXfn3etgl5/C
2tMh4GV3kcAu1ymSbBTXlVvEEwYLfH5Jec7+A4E3dBI35orxhPQLQpr1yO7YM9if
4IVwv7neZkJ9j2ha0PAME6p7wh0VuOaeU3zpw75H6Ua/UhHk53UklJv6IIRnFbld
pdjFIllOJLVyVdEKlbkmipKn8h89tmTnwRY+kwkXCFde1p5W4lzPe+tAbQv8G3BP
vhSQjdMIFlid6HKeedjKW3X+/AsFtQ6eycbUrNKmlb9BepW7J8oNjPKBQfKjWew1
l4Jqpec3fwBv5UmHE0rdz0PrPHukMW0IZxYHx5xRYi6T+7iWymzeozJRSKp7zY78
bjLXJXSTLIjelCa7po85emvDHAU/6se7aD/Drr7DTo0//OqBqJa95Wi59cEkNsgY
jQ0w26YbbUOS9w3w3bO72Qynoa2R2ytjoVwTlhyN2RMfRBSPgg4aNFlLmHqOW+wN
wDjyh9vLHS9yUCf+0S2h+69ltBUrXrILCWYIW/14lvC4nKruP3Mlc9fq4ftGyEAl
SCy25t9yBPOY0/H8YmrG1S2aqA1WZQyuK4PCyPTnvnuzZAUYLliCv4ihQvy+Pw+K
E5Odb3HNfk9UnipmcN/3ZR9N7XX+gUK0qX0Rwnn2livNa86QVYY1UMYz1k8ZnSoj
4K7ufzOxxnfxDbHBFTZlPdfIymCMHaVAl2Jni9Djy6+rswr1xy7byqfXMF0KoO1Z
FfZ2p80Db9eQArLEVaYBqs6EZnYXXg/Ut8PclLxY6rnBspu1yS9VGCcynhcntXqD
TTsb0JlsvwogcXXEtqNGMaiyz7/uIkVOqj27GCjQzC8fPUh/0+ng6b4M4euplx5b
ESX2qLeH8tUxNLxP9ivK/Fcn9U57h2JjWVoFFehzJPyLbFpy/YGHfmPtZhn/Uknx
nYGDTRw0lUhpXmpA5EeK17FL/B50caAIUYcwgliCSyWoGi70j/ySlz/p+5dvCMt2
OR9fKilMzyaV1YonzIn0qFKvYZeR1aVJTX4GOUdAvGkZZrlQN/XVEX/mr7i5n5Yq
b3K7qiUhswSNS7e/1XFvrHY0Nn+ZDm2GmZmnp2MEKVzebQ3XMC5aCGwZvQbYAsAc
dfHpJTpcGLMd6wEy7t36prx88Hi7hksJb7L/8XJ/QRI3RA7de61syvey73k4+qlo
TIXrYPW5vZ5M3WDdrsIzMYzHzoOkzDjAoL+CDy/Ntyu6uBDIHiKF9elwtl4CP3nt
3hLkLWLUHYxLfgJeeO/LhxWB5SNR89AuZGFJVN9/wJkKYeB7SGWwL56eqe5pU6gT
vkmUWRW4ew3XagkwrnegWLT8FSmsUCAyITVmxorULSWMr+uM2hQFBh/vQj2NosJq
6axQ2UK7Jd8uSF7WcRyH5BK5VtbAS3WD3Y4qujtZhD5gMN4FIpo3/MO4sZHKGxHG
2D/scxS0Dbno5iX/ntI+ugzoOJrMF3lGuuFWcKskmSyvzn/ni6kjywgFq8llHQ4E
h1N1BPJmSLyNJkBmqHc9wHtsKjqZoeurPcMCUUHT/wl1BrsaZj3Tavpf3UMgelPc
9iF+Tdx/dtMz3/amoQtejGjc59acZl41yoRU7JFNzJZtQG3ED1DN2lmf8pkMo2Mj
LHPb7UwGjqrQ3EXSMHaF2UhiV/YAH9iBZMjzDs/eV03sgjRE0n9qAWc5TBoFo+/l
jp5YhAv08JS/MF9hXbHaacQVKDt0vQcMkR97mi0SCE81e4rZMrbTsoVPWac/vUEG
icMkKpqytgQQZx6wArM0zDyKbe900iEfm/14alV4K7WTuAuINNZkTIk08m0yX600
ZUz3Aqk0A+U9miSD9kEfnKJse07exVOEMMohDWUk+Edu0lpIjHCfNeeZf6NHtVHY
Eh6C44Mc7KT7YKX1DRkTCPPb/VXeMqWSbi/ZBRgG1SBBp/7XqRgZX4gXXj9ndMfn
WbeOEtJNC5o0Zoc3Z+vHfRX9o+pTUbVLk3Q3MoZs9NfLPJNEhx2gqydOWurFI3aT
x408x+c/8svmuKfYzpqkoxpemUQV9kiT00p+/RUFtJA0u+G+AiTkllQk+616eKW1
OEaFyCfmzZ+bZ8ouYGlImefYS8e41es0uGTJiAcJhz6SaUh+0Mj+IRwNzK8JAiuw
jopae94272GISghzLXnzaOK571wEv2ndaPsIw2vSSaDiqaJjLh42/fc+h9q1OoIt
V2ERUQehO95vtQjuOIJ77h0Rt5ZaSCNBrlZvVlhkSS4B4aC7wbDEImt8y0aLmneG
eLkQgJT8rBkBAy99v1o8Xg98q1lVWB7U8GLsHWXuyl4+J4bW+4kgIyVymPC3kz/y
PzMrRBGLnUt2fVrBUCARzLWbyXgLip1yp3KQIxyegLMSoUty8/iCTKjhKMNqxeQy
yrAvLvsQ8m72zEwtpkZ4LNW4Zld7cA/T4D/uON4t3a5VK+wvcgBNLumBabWtd06U
k9yBcoHBGPDpFodlrfvFs0nuI4QxzY6kfxFXO52nDgfGWCWD0VORhW96+No6t+Aa
UwDrp0Rhzym/h/mi6qKPtLiycyMHXiJJnFEuBOeGKwBG//PZegBCYF2sFqK+Hbqv
/xfStsSna11QV5qDp4LJB6qAfRVDt6Nh+4+BvDt7aTEIw+7ODUIJBCVdIOi19ovR
l5QdMa3vjRAORcwZpW3CZBgF3ifYwqQ/mRuw2AQaqiDG9wtnBSpbilc3jM5oxUgq
/GQQ7lewRGAG+L/xXryiFVXqqiuhb64EL9Tj1ZmtT7QKgz96UWzjetToGkRK+ocO
wuXL6+7wAoH7aFdCufb7XsocYk+Q5MOVpQ6pjH02yzlT401mtqkRcP3GAgOfOYu4
gi/xDr4CErS4ONGLyIMmDIajTodYbqtK/+G7nql1su6Oav01GCgI07xeprf14F0B
s6mJKlzGx6EeMEUykL1jTWHTb1bSel26vHbsNPKHzT6t+aay8mP3RHtDKU53QgfX
9z9FyS+Gp8+rj0ZEMu8/qp2iXmoNoZnUC/Ch+vZJOlUdhoKgypgigSbg/Cdat7Hj
AGLrjbSM7EphURkGXB8RxlpBPU0ZiNXnWJQnOZsI201Xug8A5A41ILxDXvF6JHIQ
mINIE6Np/IV4MjEaXOAbEKmcJr9JU4zwGVcEMW2tgn7SUUoGhEsqGDpKpENcBcnY
jTiqLi61xCwBUXhquU0VgwRciIKL/5EXVA+mVEHrkC9d2MxRvkivrRxw3RX5zyOB
Fao3rfj4tZQE7LZ4SI1Vy/tIAsZ/ADvMnYzImV5tKxNmsz97oROO2iv6iWqsHMgD
kOqSKG9yFP+73IaEAXfw9CFObWr//JXUvq2yLRydARrPNrLg0iPg0DJZbM864Nx1
oVFldaoKz0QJnElvcrRnL7fpjt2OSMLQEDQJUzVndY+FrEKp8BehxBzGvNoSCpkh
GPzG8oceGiP7PqgcLKTj8rUZSIUApJuKkFRC10oMatBKy1QulHUlA4Wkt6ySwUgs
JQ1jZdxU7BL+yBwUedeTH1B6Wl0E+yXmxdTRZTlfLZFcEzPIsD4eO1Gf4lm8Yuly
jwSXBrkWWt9V4AVz9o23DwhRP3dTOm8D7Fif0UPvSY80Y24pKzd/hnYGLZGFBVpH
fv7chU4bD9a3pwAvY8Z7O2CmKqN8gp/oE9aWCZVM/N/pJ2xFn3RnbGI3Bb9wh6po
GZw/vVG/7HYTi3gJTSJ9QCsGsh48d+K++Jnf7lEJi3vhnOkuOXGd1CQbuU+i/00e
KBiD1JoQctDizI01Bh1tOsz5a6hZf3YSfKUvnmjY0oU5Ric+mS/yJ206YRg1TW/M
KJ6PlZq48R1Yms489GFtq4F5RU8mz2UEa/zG9+vC2kudBItXe9WgfLiGBD2R/Olm
9G+koKhckt8pVFWiW9X08S3j8pdlSrq20h+WVEgE3phMN55h23ioSDJZuvIu3RIT
NNJm0esDDmPl2x1nw6PAFIQLopH8IZ/OvOYnE3cQEDrGFxwp9LsrHjDSSM3HK2Gh
SwOnf4yrTNEyHo7KvKl2ZIM24Kkvus9UC6DQ5cWV5FNg2QlT8xjIij8vViM3t3bu
yJHuqRZ6m57nMbroCwc/r4JNfxkD3HiVj+OKZ7X7BWx7p0NCox9NaUeCFzHtIbEW
sbh4jmbsUNvDErFIljvCCL+ZbKCIu28HXxT+RtVYKpn2DlRxmJduCx80Ob0TWFut
e7pmvXjJluq7m6u+zipqRHcW+R/Fi+CY6eXfbCT/YAxNZcVYkE7ZUQX55KZ7488a
S4tAyOn3MDP0ULTxL4z57iSd+tplT3v5QsbtrmQqp3hu9gTy6IIlojQdb90V/o9Z
l48R5DxY4fCemiX5l3a7C2jp885XTFifoNhooHmW7+8rKcorwneFW01uFNCx6oEJ
5/BU+QXRQoPtisl1+dw1qreDDaZRdnivP4GKxBF9+WzOb8eNKCHjwENBRCyDnNyk
drfGUCYta47nUIw3vqtRzYAVBQm/jZB1eqdZkSjlpmXoFEFibDEnoBlc69KbdU2f
tJ3MY6jevR7Xn2lUDZITKXb5QH3t5yaVGCs/tL9UBjSIxgrsGNFTHPeqwEK5cfaO
Fis5wEXIMzvDTVI12UMoMnpboSMk2Q6esYXAUM4481gsrcjIXLxTn1JVXMGna2U+
qR+n9CAV6bm7v+VvYOLdQ6WKikF3089kmANwO5/uircGEx8gqodYv3jul0orbR5n
uQtns8t+qtdgtLOJY7Ex+SwTsRyxyyycnCE0fd9P0OyMmIR7KGcmBXf5F7oeF5Bs
B1h+gCZnRSGSIkTx6AoClNookJPzogiJ5gw7a8/KlMMxl0klhnBQshAHPfHYqfye
O94OJaDLK7A6oonQHnGOFx3qJZK3plw5uHX69hSVjQQvu6Q+EYhKCA7AFZ637YI5
4VAYN4zwkwo6vS9YPxtzaW8TI0voaEK6F5bjcRc8lcPoL9A2hB8LMbf56kDw5b29
S33jKUMehrpmzY33qaVxw1PWd3Rk/t4E+fLYV4XAk3+0igmmgHH1EFs8Fs5PPO8Y
Zsy8ldoMBfK84sMlcLBZNOaHPDHBR5B7Sq8FTs0WUtDs4CnrAd8d/E4JttizyCwd
RfHz5k9CTfmAjJyfrZZ9FnOJ6lnkNbcHkCQnjIhTIYRZy9o0SLASNbY4Khgc7d+C
18cS4M3zM+iwlwSHjKpLb7bDjmFyK7lKIPTb7SL1kJdGeDQVzrq77KFqatF6Mrxr
e4N3YwolcBfNOPySkqCyqtgNPTklFHNNtGC3lctlVjjqurbhxUj2AMPsqXeySF2r
ItNFc7rxrAsXBDhc310NGW2HbysulDmTil0WlkLjJSthSaTyeCx5SOe5fMwxKiXs
mOKBCZCvquhg+bXYTIDN/CSCMvuGNffNknllhtY8qn1uHwNckIqrK36byS0IZ8TF
Ocx0mIjPd29qxFMzIPW1ik/Ip1cv+31BEZV6YbkWmDYescrVw63WV/6G1R4R6J5b
1HgVssKiptiDMrrpcpZMku2fKbaoH671CNRhbUkwhbYtk3/JRrxzWc/xRY8ujltl
cmW3djQNBKKYI79hZB7fBTkCsxlmBb+c29ivdtFUWtE0ijslPSexDkU9VGQDT/0E
LMJyI38gWzbfzBTuyfsR1pKz/QnfLOGV6t6VKRHqDX87yASsAGdht2bdr0GvzXYM
c1OKVgOmvVnOuuSSohlpCdhLKyqVqYiLW72EifosxGz0KqTUg8QdEe7rD7/EaydQ
df9Iclz5pZ7vxKNWwMQL5UMbbqL4nIvaKUQsaq36QM80TbA7SxgRdHc21eFDfmPx
FLEfpUrZ312O7cRRDTrVBMLxbvfAQxrc7h4Jeb0r0Xqr799pZVMIIi8t6MzN6uEq
a65Cps2ijUdccwvyKmJ7ZkIuNXhFsd+XhShRYU4vfd5j+I+1rLOFyM72sjQ7EAJ1
8b9JKh9BRUGgkFLwT/SjhTKKhiJUALd9a7Uqj/GxKRzGXytyuuAXNhkWBPJyf/Zh
vFwvsBSywkvR+PqhjzHijvTFzDZqdKHpR134V6o9pUqa9apcMYHev2eftyNSVv8P
LOjKR3+joAO6NjiG2JVBnIIS+6Kz654uKlc9R3ibkGtqEqBEuP2931OkmqnXkzT0
th2MQUyVMlUA1C9v8SVDneNBncGPDOWgqwVut0nDQktx/o95vyYElL8dRWvdL0Oj
vJfNFvn829oTvPHrUPCkvAiPFgTWqReGVkV7M1fE3YMkRzRgPln3zjJfmtTmmkMb
0weA6pITTtGmPw393o2XejpSUM9rfOOaI4GXLOtcME95dbBXZMWerUsT8WsKEDx2
1C/OR7KGVkfkEXIwElEMFTgoX5dNea7sfN8x92m6OrNNJlY4dCrl4v9iqfhH15vV
bnvO/rPDI7rSoeru6pp/uG/cMvWOQqLbqMta6TN4I/i0wQHw46XsmKpBjHsVY96/
mqmQgD6tfLDw0SDoKdSW8IZAhY+Z5MIF4ICJxOIffybX5r9Vvlg8dDs1WjgkkeuI
kaRgloZONurR3DVSt6CfxVqav2ueLy1LqC8Idwpur8Oyfe/kKgm0LtbR/5bOLEiW
z4kvy86tli5xKJCb0tyZrZjaSJqfyNH3a8+C4KgDE+i6dlzmOLJFlQNjfiFoTzgA
0urwTdBozuoTz+ijInUC6tv9+Uw0iGQPkMt/aixQsIK4plix3wdG7SQrWhqWHo7B
xV8Mm59DTzoTOVrIDmU1VuWk44U0ad+Z2vb6mlW4/Xc0sElHf647UcB+hL82TADK
mpJc5Lj2L1hsG59ovwmAfEAPf/xyBnklwnhFgVwKVRoCCJfftvGDkUCWLl488Hyl
H41Qzbw8iu6CAoCEPnxZYaaATeRiAZX0RI/TVLxvaaSynQ/fzSLprVZhM0nDN7pi
W25WR5oEz7s6n4cKzCbjhJD9dCS2lmEThcEKAeHl3PPS/28rEBgUU8ydoVo66cI7
NocqYkb+GA8pJNGyR/hFTOrHAvjUK8BalNBOhvU6qg9Msp+/txD2CqUaT8TR3GXS
A+WN+035adao8UrmZbdcsRtEvhBFenhD0YbdxKwx1c5Vx+G5HBPlZ1F6vsdDnDVu
dhiv17Rh1pS86a9qUx1n0t17bv9aYV+T5QsETwZZRN8sTPrFciOLlCweQpajzALw
6YT2eKNEA9JZk1Z40cBbPt0VNQWPtnHMzOqERpQa0fa8vrY75w+8CAkoayiIufII
vNDqVQzhvHco6qfUrwa2P2Bv4qv0z+uFQ2QVbrJTPSOL+vQjU4g23PXwqqV3egkD
AZMUBOwZ1Y+5iRJFfW7a2hfcU07hYOepZLCUwBv4FA98nFHA7NkAL6oT71g2iegd
uATsx+eeyOJ/aKSYN8r8W4kJ5lHjKRn9hzmdQlKtxQmWBiNeGJruMrOXEVVZvtfT
DKxdlzFxDr7ylwBgyuH2jyxY+qvZqy518DHh1zz+GM2IXlYx1WIKY5JE4lXsiYVz
4Y5zwxyAyJCuOLi7nZ1PDEPHJ9s9snrWciopSZdKPNSGwZbraIPKXsbFPOubzxpm
vn2TCp1j77AedHQmmMwZMjKlFdC7aAAmi73RCQbI+nqazo+mbdTHhul6ODrXm0Lm
1zeKUrC1umb/uoASS2JSz2AlL4X4HMSt1MjAJlgFb46DAH+cabprXj5GOnR4HZoo
cROyfqEozvkEhyBf6MZ+YFeevzURFjhy/ue9Uk8HScnFv/CRzvIDOsivXNRxgOyw
UVihMeyjegqH2d8VSPuHLAixYCyGOJdkOSoEv3RFV8GQsScneyxSPcneBrDT5UpU
CIthJpdcMZ0fcOKgmTziX7vVQTCtAHzv1+YFoY75/zYwGakFjFLCrHRNXSEHnNYk
MrDDTykZNG1/+ZcOvFLP8+dxHnCmbwcS8NmmS8+sJkC4tj4KFTLvB32aQGvRbF9a
QTPsduFu2XRg3ZNFqTOYr9Vq7RlGz7imDJna+fg+b5E4WOVWdKZbyM51i0s8BKX5
ALSziYRVLq8R6XP7mXLIjwZ27oooMXZIg21dEKUrSRIK35Ro3pW30X9vP86xtEHo
ApIq9XNJh5+naIk9gctOMhSW7ry1G2TqW2YcbHThXnFKwsp/DrtFvwKJ2UJD8BSu
95vWLh3UfrpCWHJOUyzPNLV42EXAyUh3WIxWmmR2pU7FU4Akz/lG0/sNv/9Bvc6B
5woRrKRmtjuREqzFfBKkPA==
`protect END_PROTECTED
