`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Sn+gBM1mp48lrbMN5sS5tJUdM0Tl65TaYqdQxTfzH4Zi+fHzJ74xzL6XUefKf0xT
94CZvBa6oT57eaDseh7dGt9ixl7Rpg4Cuz3d7STuw8zBAoSYcef4r3I5x06I1/CF
hO1tPaiNszQDwQvyDAXer4+i7JIaV9ccFL+qQjCtcQiYRAsH95kmygn/dF+5ckFg
GsI9F0izj6TFJQ4jPjwJKGpi2pEJIL3HUZWcyljLpkPYl6WGmwxclU4YPLOgrDlP
Htx3I5nYIqhPEq3MCeXe4m3EyLX3zz1wLzEukgB72qQdUqRnvkH7xsp/ykaG7DfF
XmxOw4pUzyzN4AZ5VcsLvxSurLZj+dEHICHbwznSlJaohlVkAQkhTBFmVK6/J7fS
RIqFafPR6rx5aoyxXf34aCfgyWuWToRgK2IeRfFlHhM2rotxkqvuP9MpUcqY3reR
UVOmXug4WU4uY8Yr4mTnxtmc2Y30y+GH1k+TU9FIr46aCJXUBkike5oOHpVqe2FI
WwuMpLo/nN5P4f/qfPEPh09UMe2Klr9HC4CmJG1Cv6U9Dzyl3Use15Ty5h+ntf0h
qGZ1xctZuE5ErWAxjKn1w/LMMXpFkAEY5GIZqnq81hHEYHCEkXDp9IEQuBYEaief
YUAO1sGaw0qdfB9G4Us7aVs5hC32mz1KBjiVTG2O+CKDf8pmcXMKEbfL07fxwwUS
KCGYZssfF6s78YUOij6GX/r/7cOQVC17Zl3qjWBuQpAvRagnOeoWDK34D61IftWI
ERG9PUmgBEbC60abJDCLwha2LdOJOLKdPLhbQvYqIyQs/WN+HBrj46eJNkJ6SndX
LAVP5zcFjP9CBHPXjiTZlyiBzlS8pQ0sxWeZQw3To/lB8qMK8B047XINfrtmZfGW
Dm4c0gpTFkORqFCO1GDE9GV4S+9NzT3VY2tG/y28WiDvK7qJLNVfLezrfCnPh3PT
NwACPLXymxmtZ54BlLJLY/QfblteKyiWwEXmGdlBLTKYfGlNHVcoZFZ1XkRiUP/8
GiBf7i4YlVMw9QHkMTcth4O/RTJPdQdkCB2bdqlj538U8BPEBmN4F1xLAsuEmtmR
vxgHiUpQf4zBr0S9JaiX0NDZ+BaP+AMANlu71XHq3kQBOxVs5r33ZNnztxUeHV4R
jgs9fRRA8bgUNRpkAfYjuR+XwNcxsTYS5jQ7dTE0xNBjy2LP94V+vRsX3OqMJ6Ms
zOr55e4bIe9GRicc9X3xNqualR8qf2PTiaxNayCsNarUyV2+xNyU28L93sn38Av5
ezUrSp9OVfuG4sCaFh6mDbN0TtA0QGaHMzbmRazym1gzNhDWjx6R/ir0rrjt3UNt
cd6rMQ7G85Tq/mlfRUq9jcpsahZRp4wFpaWCgQ50HIqjVZbLymwB81XqKRC0DQpD
uJiwTcH1LK2MowcuVauVMWl+0Q86QWCXoPTAtki9/fuTyMEgz+32A/9YbIqeFZS3
kNSSyUACZntqko1ITfTY3TCZ/oHwwNDqAcbDbcR8Fj2ggj5xsQVqzsriEbxLHk1B
GRHDtU7/8XJeOLClp52km6XrdiR7MCMBFkCs8U0hgjIe3GR0qcr5ayq6cdPWaCFQ
0bQ6QFQSSDT+j/CYBQ2ChwISOiE26260DC0I7WngXCPgro6av7j+w1aCecei+jve
NH1k9b2al8iLCqgiQqRv+gboTUA79c85GSnfZJi8jjhstP/7dStjQ8ORgfkTWqgY
84/FzmyN4CPmU2O47j68VlwoCOh/+nA4N/B7GP18IpNY57jlPt+avgf4RY4fypmf
DDvVXoTy3UOvIeJq1UV06ExyirGNCUOMRD8T5sPgUKNfp4Ua4EXsC+54izn1gQg1
Kh7GPJ/26oXCtj4iDQc3+p+hQ4oI0DSbUL1SqkSGVzMg4aZwpv6c0dK/CFs/sNLN
Tz56dWzt2KO9fAbJVOSrQxlpBHv3FrFc+W2bCoTrfE461EuxcH4C0aNnkQcmTEEn
+7XRO1b3nTwRQMcv01Z1/FsZvRFH7DlEV5pv5iZsGEDxniKeP1AevAHa4vMmqi1r
Zi24mJpMBt7yDmR80urJX2zRjbVdwwug8gG6lE1WVWG0drRaM1/7FTiZHGnBLXOm
UR/ixWRaQOBsolFGSXamuc2tb9JtYAwTmJTqH8BFZ143UP42D8zwDd5XZb7hrCGb
LAzZdF/16rc7/S+pDCSQo9bNucP2S4oiEbkNB8lJRIYFG4TMbSbDnmpXk3Qn5bRO
KDmIVZJPj56/0I363IhC0fHn0FQd22o9IVdw9EJhmPWZbKJBqLt9e+ryT4V1BrMV
D1FP5xmNQg/8cHkFPtD/VX2ejQphD5I79emhXd74WK72sT9xx8RGn2mjP6VP+7vB
Y+/1kTG8RHGZwKL9fwVBdRlGODWHm4ZZweiCrzBzH/JVa6jRn0d+NSEjOfl7hHAW
QdGV9ck7xC/kddmq0v6iYh0IUcjdi5j7rXnHhmTTAbuDft3xXN5oQmY5dNZSX68M
8yYqo7sMgkJD5eJ/YlwDSDNNXoPCaTJ+w0y/2sceVBLmY2RB3CvxvizQSY3mcANA
nuNmd7KRDWGGO2DSuMLrLr9IRzE1qG30JqCox5NuQ8QM8+Qn0OXiMZx4IkaUGyGn
uX6WI5zNiENzkHQtJHB2th4B6/z34JQg67S06v9tCklli3Y3zInUoZc53/7Lv3YZ
`protect END_PROTECTED
