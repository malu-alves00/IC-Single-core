`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xNPQEIysCuJZarN57ewCsdxmGP99ytuUx8ZNZHPGoOWhXlCFbZw/Z7idB+kudGWj
XrC8j5VSgDxbZVWVV+ed3at6p6hkGS2lg0v12kjaa4p9S5B0uvDjj5JUdiJTO/3V
9W6uyRRd01RH/MiS14l8tP9iMDwp1nIRWAY/cNdo/sHZXA9Vqwyul5sq+BeNz9zr
1b+6tctafRf+sO9bMykQEkKuNU8MyG8lXhjATZfWHA2Po0XEoaq2Oeq/TtxD4+R/
8GdITDLxPZ1McxcFnu6hTcUd1Ki0NxpwwogrloPq0ncydt/HbKN0nsZlhh5BEki9
60e0/LvWpdBvlWbsBMFwugPGLWKjqEKgWi2/Dzxkk6xWb5KPAiLP/5RNZNtuCX4A
xSx9LhsNYN0F6RKUN9DyW4+B2lcpEPR4fXyFL654SrPIYn/UkBPF0QAR5v8Vo1w0
KhxSlPc2+4uKKKloifH/FB33N/b3AwuXBbNwEJeVZ0rteuFKIJNAJFllQ1g5KOK2
kYdj/H+2nZdf8MvX9OdgyRvw7q/OMiXbbVDVQCzd04ifdcQpDh7YMhqtwBTVz2+Q
+v/8gvD9uB1QwjuFmfdOlFRtLQZDs85xgN8p0S62Dkk3ZikqBTQa20QrLQ+sd1Ip
pwe2rxCui6ZVWahQcCFyynlQvSiKxQxdSqwzdjt/cvzeRLqg68+5VUeFWxo1NKj9
eRJ4vh79Qwx0asswP5OTy2cqar0kn1zE9pEjGkpiMH6/LRlrNXYRPSX85Gwt3RF5
CwZvjh4O9Lg+eJB7qpm4z7DmWMGyzUa3a07UnmNcP1suh6QLJ7tc5YbyCVTAYKuE
RYTx2/96zXs4vcQwHnvvcMJEhjHHLW/jFjejmzPVFVHerxEEjPGMN/AOs2xwFbed
E0ArrdyVEcCQJHIz7EMRbKC+3zVK/3/A6gHdtsEZ62JGNs6XCngVHp4Tzc+AMSNh
/2ZP5CWSij+f9aWgkrwqpXpy0Vhoh5nKvh0bmhc/4zzpM9kNzF7rPaUI7u96MI6Q
bDeA99uTqVxnITZeyDD9PnXmGxmBQeoOgpCPra+RNfM4zyVw9IE4zbb1Aa3j8/3K
XL9zSEd2GEQTUxI6gBg6py8wMLCyEVT82Ql/4h6TyLOEkaPtzM2w0UBf2KSD4j4I
7UI+8KrPreUNWg15orB7GcWvox8DK62exauFZODH0rQ6TgiqlyIVzvfRHWGCU+kN
f/tv/foKiZIM7LwtPUfSHSMSjYHfN8QJChKmt5F8wyMAurClnffuYPNn2nEDHFFd
KqNx+AFFdhNNC5YOiDMQlfOwjTBQ9XTTx39JGHC/qLGKHndTOU6yZh7B+/UcoPU3
4f1gUpD1X9eSFPssSROdVhNWUXzsN8d4nlQleEFPdYowSmhSg5O8ztIgIOQTRV/J
5AIEV10Ukx82w+/57dHC0sgoBrbHo1z6u3mkpc2fI9QwiSAaBmXSuBHXrqHC8tfs
ereBpbQrsWXSwtqj1M1AnQ/O4CCFdlHFth22N6rxcmalql5/wgehnFbRPLrr5587
VPCpZqf4mcPQhmEOU1LqsNl+zKGjsIQGQf3fheBukCP8NQuWiTP0gnZKEUlgHOG9
3J3mmMaJLH5x7INxU8pXqc1982Y4A1/VOUjgs0RfoLj2VW1Bi8VmIjmBN6Wumwqw
hD6KTKQVCE4jsyf/MJLqkT7nuo0lkvNRMdUWuSr4uaHNvLEEPL9V7lZfJRqWXAYl
4ON+0i6albrZz8vfGlPoGlLk475Afk1cqZIaewuqVRG9LyVuBFq+esQoeFAFWyfP
3RHsKGxCYkOWOG6icpaW31CoPL/4mxOvHngaZ3v9lxe9qk7yddSdHMvyT1pL2RI9
YyK9iKiKlKZhsg29qLkPX6WfvHx9/bXM+4XZPF1DE3zEN3FOiNPdjEq2oJ+VJrQg
oSIfEVmQKta/l/E9FV5JUhyycvGeHcBxEjR2OP+zqlrxIlySMaZ1eNP9zuPsWulx
wj+de81ZxNCBCKpAINmjpIC07F0LJwJt3v2tnrIiw11KQOkiwgg5iOg6ehoBfWfO
0hl9RJ/kUANKQ3Vn5XLjygbODw6FtNA1qLgXoD+rHbLxyV5WpPdfdApkjZPnXH/q
yTJuQEnF3eAwMb3lwHuWmdBm4bUr3jkVhxtLjqzb6gazXf1H/+W6OeLuYTLFioru
H4wdhNWG8VzL1zQ9bQQgRcHeSvrd6JPHXICMg3TJ3Fzrt5mn36ABQyHFT+XG3f9z
D6Y05ISttf1/tkaz+JRku1s8LpBQUswq4D/8exqGHx/Rj8mIncVIkwb25wUKctim
hIAIoa5mQ6GoVVjeKfwD9to86DIFjXB9sgsk0o5XWxlY4IOR3XPoOY+TmF0Cy8B/
5Od5Z8pA1kWwo6D8X8dPawGKg/IPcGBDuhKsRpjiUNlcWLgJ6zRNrRd/UcIFgWdI
ODrEjoQudfZylwRZolA58XfvqQAunrrHgHDMcOEc6B851WDeiwkgE0ZzC845iOsU
n0HL60fk3UdooUEOQU9DG+Y482f99VfPlwXib3IvX0PZgqitVAfp6ZwEYEMPX0oE
zgWYPdfXJvM4i/y7WCiyrNR0a3M6r3gjWehDc1AJ+6PrZSHNdCIIEriM7hBzqKZo
JDFPPICaQcHKr0QXyV+FrsjqmlzOuuGyGpkM58wGMU9XIGeitUvkvkz39OoSUGtZ
BUC7erzcRK2bhoRxCF2sqa1hyTR9TmdMMCnuqF+ziMAn+TmoOQunRDEU1GlkDSsl
+4D/hIigaIdgnZ07uRO6q9h59qHhkLaI18Kclj/bjtZn0fQ3UOcN5Pnhg09IomqR
ZStW24kXLBOIaf6kaQDBU00Wt28j6sJ3j1Kq5xB6/Fi94Z5yvMg8OGo6fApS7ltD
lqsWBUaTOD7N5ii3DMGJhC7q2QGSAIuWJSr1MH5N7V8s6P++AxyfI9jrC6PlDWZB
Iqr2EgBDKw5FWlY0JTVl9rhgw1x/j2zAFN1vwH5PL3w4D98rJv54zzla4BqIPSJY
mDq0GZO8MaEoV2jHGfhwpNCMLRaFJGlVTwAdoVnvQLZZNubw6T2DGp2iezfNjyUL
6ExoWLCyu+Kma8diqdpfGsN01T+vcpjUjOATtRp/QWX1dR4viKkXeMDqDKP20ESr
/Oyaqz+VVs2o+cRyBVnJr42zOMKvb7wInV1Q2h8voWRFBcwHNEzxKXQqw3neaU+n
M8VQyWP6JgmXpf+zZii/ItEu6nS+U/rYyw9QHOPG5alt1S1gOdkE5meFt5G9Q4oo
Ui7PBcWr9ID6XI3n5jxUV9+3LBM4KbCgNr5goVRi/XF1tD4BGmwzD/LiarcH+GV/
KaEeKmEMjXRBvQSM1RTgZ2wp646YS8TtR/BFYbo6bEvSGkg5l1JJe6Xky3INOxOn
o/A/SHH8UwErIiksp/67rgQWF2+9RkfsJ/1IXV0mvvLfYzbwXWYbNL1DaTLA1yKm
lepwqfCp0QMd023qTolCKN+sirA0TK/PHou2g0Ww362ZUUPh8icFs/KqKFC7ufIj
Lf7zdi3uvQQy8W9DA6aIA8GtlVyGxU6E+yBvN67RENxhTxVbrSym8PKTT00iGwXj
Bcjup+yyD+fIjuQA4Cb7MokQS1dILCiZGNSOM7uhGPIXmGPK4uFH2ROF6M61pErf
PmXf2SObg6Ac9MlHnu5YmijxRq8pRRk43SWY0bLm6aISb3SB/kTMDDigQAim+pH9
2h3ekHwqppYai5EogcNglpB0z+saWealVwXEwv1x2AkYgHazrNgxZHzbQZMgvSUz
guRrhDpvdMHCa5JrdQBmqtGxx3sMVljN1Z3ikySYBxKNr+zDzPC/ntbWxuWcrtyh
faDcPoDXyjITizrrtFZq24WpCdO6TCCfWSKaH4LITseXwHyZfGJAiCBd6Ii/huYK
SSpEKNNAhnrkDEpBxo+4rfkT8d8/F03GevbCpL6W266+r2nH/mVc6XU7YZpIrXzR
HsGyubQIb8Qg67nnjKkWD2Vh5A/L45FPAp85ZXiqvYMGn7gSg3wnUNQx2knLMA6D
zM2EAHXVV4DzyEVhueiwQ5w0hMlL1t93O0jHPscI4Qs9/oOdShaUKSCeiDgVptJH
CQJYQHkexNrdc5smnLK8QeZ/vJYZ5z48RJimW8Ba8kRSZjsWCbWZMZmRljWDAD5i
5eJiLZXlDCeFELzr7y5TrkCsNzhxDud8hwlmljVIXjlQD9tnciV+t4XqmMv8uBqI
e+lLxCwppSzFU/Dzc5kgxawevzkyB42l5WTFVZg1QyBXclfk957lxw0rSWLgmA/N
8HKkYUJ5C728xOpXSHv7KBNC3PsIhre3tV19dvjVwjiAFWCaKM7gG44obD8YFtYq
8n+IRoLgsVqLgeCKPW1cC+md2TduV9GjbS9TP/gdgP/aEoac0Y55/Ia2K1Q+rbSS
JBkcDSBS7Zf6KN8PFr/tEEdnTa3cFHI0/JjvIJ6YNBkps84I4ILszqsROR/2sEzG
ib2WZrnSMaIqiRwj/TUGU45xEbMb/ES0fviZ2LCnioY0RNItI/KjQ0Hh1GGz9TFq
X1BWXNOS+C79cAI4mtCseApc4ozgguS6WgIHnomrdDHwrRcb6XELv8HgEGvpAXBJ
osveMoFAOLqfXjvNN0ZBUfAllDU6bFtIZ1gm3wB8ru+JgSgyJHkqKdXAPosAlpXF
O89XMiyZmlLUkuU7uMdWqbrDP90O++ILVGcxhgRHF8ZTJELmuj/rzCF3AW+NHsYv
6TSqKr8pi0b5L1h+Pwnlrhv1CkJosaEWFKgtGPnqcvE5eBgvhrM1iRPO+I0SoOxx
7pi2JBwHnknoLo1yKyg8NGKFGHLCWG7AYleuGO8FeyHgk9DAoZi+a6aV5kMr8mzu
VIZ6AhUOOd2N0grNrJxqkUPYaESlBtLSDewUf3Lu3F3uEjB+Kd4HIBaoEG/+IxwD
I79YWvr7HFDJqvWY2H2BY3mTQZJ3LkwAyHFnFdLbjwnl5wF9zUj+bHG9PbbAlClj
2FCA150jIlDo7iPtIRFjybkTsW7x0Zcserz4HNaHheR6l0mDIb9NeumHh+fenPAu
VgdjZzkys9YYsG4Vbv3SoPkKpt0dZocP6XKNo8KtTeXl2RVx9bg2i6HyviyY7ncs
xyjn6numS9pQO8uUzkNQyAj2g8rH8STBMW/QUs6TAsVcbEQxAHgH48A1R3Yu+p4I
CUqAK7N8ti33ncnDWMnr8/yJVMOtPos6RgpSucugSnQBx5wCw9uuSb7L+L/7xvuI
lEUEJlKcjDZTMzGiys5acNKrDsCZv6TYIKFUldsX+TWesKU+hc6isNQE9Z9H9zFg
ZH3XRDAsyHsP24dkrCWBoBqEdc4PhVlvtlCJNQdWEAnNEHuPIv3hYYNizCvejd6V
WHEsg78l9MC+WH62nKqbIRnks6RNzIaGmC72NSxaCdMPXJfaG5F3tR2jpyYQThZX
t+hfCd0vDIzyPLeVSc+m7WclJi9E6WQ+u9jUBMXLCKucHugoTYE4oawLqRpEMNhF
25wq3S6dEWENbkN5wQSKexQ63o/RKhq0zRNVNn7Qf3ogOybVe6CUjvjgsybpw2vD
jtOlasJIbr8SZdwEkHJjSpE9oiPJu1hucne/gaeKd26uWqQj8oF+vx6BLFvGcHof
kAUmH0dLajqj7CltDids+KRtDffEWE9qDt+daPs0c8VUaJ5Rz6oJAjqVSj7H6o+o
d+wZkt7E6LGE2agGfCRPKOcAxWfCME4w/TSTAJuJLW/LWx38QMIffu/KuXFrdSSR
4vKaXf636VvUaj6x2t/cfQnn7X9J+TQ3OfUkxNz/jT9lQdm8cxDuVYzgOeLs7fWL
RFS26TxnH0yUQ7gofp1VQF7+y3Z7tQ/Y6AECOOLWELBPt+4+Ztf3tHxACMIARkE/
PqJcHst7iWHbFdGgmwPtJ2sh+O9Yqw8TV8aP0bIEa0VmLc9srPtSpeerV5Za47CR
bmkuB5EiqblXMTE1XgZAajd4Od0weqNHSk2g+wceaX48KCrdsLir8MEPber/Hf+c
WXckmGbMZ0qrHhk6TOf1HDNDESmjDKcj+9W/s+8NbFUJN3dly/KMMS+XIVp7oMB7
mR/CrO9Ac5VzkuueMj0ITry1vcxfIjSGZAo388KrNFSfQXav6+ty/jpRakp6Ybav
CI9SMXFfy39rgrNprgYMQhKh8pbV69wwANZZf7TliEqI+3JzPZAdnfkN8/692mAW
MzwDWYD4IxZoubbwKUVIgsjvuxApOWMBYKJ7Y+nnrclHdU5gl4SZXO/n4oZ18vMM
4bCp/TUFwygtyE9eNiIvAufDtVtQjyinY1whkuPNcxibqiK1Ov1wLujzK1rLzpMQ
dM3jHPKUN/pqg8MLBxvT6sl04h5P1/Mm6b6Kuk68+83os8ByT16dWX8ebKLtJ72l
xze7hrseEKM2UuvUu57y/Vy7TtSrjI/z06/1H4Cg7epgmfjsm4hY1CjCA3Y0Iy0f
JbmUhsk8xIG+utZkaf2bx1sAuR8okT2WCu7KdrY8C9qFMdybZURu9WTpBHKrgt4h
gkobda+5wstZeM+vkdvtEBI4sQljxM7H1WOj39Cpi7KbAD00rxHi/HGPDRTJwySk
AUbXPuWElpVNhvj93WMKEd05y5QXKmZinQ1dF2QTOyCWbI3m0Wr/oMQVrEUE9uuO
FFw6Rcv9gq+ie2hTgdjEJVxhMWOJ0ccS4MjE4BDJwOnWH/+UwpOhRSw4lD2CE1y9
Bf3vRZlZbrvhOvnvelnGD/IXKGr9yRAybAmAlhNN99LuRoHYh4BpYAcL+OQ/uW57
zLFh+GxBdqmhXurzkqDZOnUd71DemChv7Y7Ni2FXtyyxluRHBHC39GEF0Wa9xj8W
6CFE12qSfrE5SBZTDawVOaYVPy4iJ4Jj7+NBbcviR9eDUDglgsvRhZCPzYNddM4C
7OaHT74CXiy6fpWl8sisBNuVqcXf+zWG4/6t+5n4ZXMXZXtxSDfCrboWRrPLc1DS
qlsttj15EsPd8RFyWoNdVsbuRKbdX46Z9Wli6lq9F1k2Z0MEl3LJFq70iXGsk8v2
L7NrtGBO2dHOpnFnxT8zQZoPv8Esx6PnDmxSCXUKDerCNnZkvaFRTa/ipHIUX++0
ZrfVET1ddIi86zrc5UQfdg9xsiywQGZI1yOENRUHMdCHD2S1huVM8IJYyqDkghpm
KBZYtQWoQtPpdpcPOL4AYZXKaF36hoEwZRHJlBTu9WVWLORnlBdil2FetHn/A5c2
Oe5mcADIxKZVBdMERkmt8pEijyUo2DapEapFHV2/XnbYsYiqGJe/XjnYpksHZ/Jb
P1OpSG7/vCjeMATkxLxapGFTpiHSgbiVYZhPbcS2SVosQ8AqZbHB2eATmXsSaND9
gjb0AhLnDYK6rsPROJ+lOKiAeGrv7gwAzcMCeuLtNArqFv7J48W/GGW+FPj+D0wy
w9sRFQrnYMBv6pBJNKC7H54PcmkIQoA3oTvtcEO9hR+JyHsHAy+PDo0v8teszpSX
OX5gbT8VO8StpkzsSANoZUHizl9rm8BM0qYYXsPca3ZDFZrtCX1SMdvK+F+y9ONV
OJWUEMDM6GYMJd6x0sBTGNfUUhRB+hULPILGOZ5CWIRWo4bQfJaWbTUlIDbuApSw
6R76jxP35qtFPvBwpU0k5Fpu/l2EATrfj/kCWtP4lizfaB6x5hCFOFjmWlVvdazq
II5uExnE8RyyZC9F0FEcFoipQ5PoMAldIfiBqvVKGhGYtnlkGTN0DYKb04fPogbd
5wL9ryFUoumq2q+dV734Top8ylMQk5Bx7fhI0gwkZ/WiQ4eceg/n0zRu8ovug9/d
A4M5NtQqOPPOShSrh+aPNdw+PdU1t+FOJXSqENEhTVrpZHWYLfKcEpiy2R8+sN0H
8ytdUD6jVnf3NzMxm5ePWSJkq25GzhhVDg34v3+27UvWHL6U/8bMLXfsYQpSo+de
GWXvirMV4JW4fXfZmHRecDKJjncjwiZHwFa94wr1RK2ZJHVR0hEM28YqL2RcG68P
s9KG0QTQRa/zXL465hyOPNl+eDYlUI1XDcP/QIU8Lf1ejJzFqQ+vFpYBNMWxeE0V
Zz53FhuvouHsLqooI8PPZKUmMIP+CAnp3n//N3Ee52INb36SllvJHCmDZtET9kZG
RSzeylVElqE1lHiQcTjwiSEjFwLwLmOJjVkSPBV9/7ZDI8DeC3pm2nORU7zQVLUg
3YSiBaMRZVermszVrNR98f3wTTnqH/WdIKwRcwrA5i08Lf+VSDUN8F3E6vbOxJGa
zCNfIUaomd5c5boYgItBFbuIRufBSzuJVOii/2JSnl7Yg2Qo8DycR9zMcEDUBsdV
aDNUSdGYGeKGqhM8hjaTLRjTgEuKtbkZpFUwBES1dNP8jzyCDJbo/wOIahcsJEM/
7tjkNQGBwjGoVG5nkS5L1X74FK6pO7amKpBH9ZDmmiKT2eN7optN9lqdVoTB+G4U
QI41Hitilud26tGvZIYhS2t88j5OenPGzgtZP/MGrYEWXBaUi22LAYgzKPFg8ESC
dndSN5fcZkb6Svc4cLu6NswRknWNjn/ehy68MImYGBNW4D8sNIJKW1tjF/O54t5q
WGjNJHQZDpfIXnmhbt72eUJ3qfY5F972YSsTx4HIJvb/MRHh1H/T28YYdPLpNAnW
WZq/6HbW21sLjIH41IkutoVpdSxV9HU25JQOMQIvXcyO3CCzUyz7rcjP0x2xF9wa
rx1kSDxIgMJeRLH4Xw8C0aOTnW6EK+cFuilHDnn/5wJ2VyU9KLY0v4D99/jtsiJt
EmIDIPpuKVnCRGk7i9t/XSe8j2qJ2GAKLAJO87pdTI0engpF4w+fewTUMzTbNiFL
NKIKIGh08YcgwQpt32ts2Qgni7Q0IXPPR7nkh5r1wknIOecMITfUNpHK7I0gHqCo
+G3z/CeMAnMZpEJA+KKJ+frUOtSW3sFB6WIZetL7RTxu//OsQfl+pqjwMJyfa/on
E/So6AR79L0vovaYUUCJ7NfmPWkLgiIfOm7CbLm2CCNvHIujokQ9cRBcRa0M1Uq+
14PepfDp4/ETms4rYSbz2qntUPQ+w05neAu2WvFSGNdrkTi5rSIVLc7dyTtK0nmH
Vm7XywHfsSJs0SalUc6XoA5o/KLj6kTQIWHGnkjY/5KvT1teTiStch3mbDiRYTFy
NnZSatJb91MV8lRCuSTJxUgjtTmfCFduBrN5gP0kKxM60sKtwa1ji7rYugJ/fou2
DprExYVRzP3xYbJv1mIM3eAise3Pzwsy3AZh5y5tiFRSB2u9kNW0fNAhJWiPbi+B
YJHEzuMyv3NxU7MaJ1b/ExwcTbxOIIA5eb4nYSszeX4VARe+4RWme4GsqN/JFnSU
Tsgwp+DHrYQjpKv2v9rHlpov0n9TucwGVjGBNQbzDlinexOKnR+wQcZsqG69kEL7
j9SSCGUcNZTTc1BEgpN/Le181tCPS7HWW93ZCW0F8wvoXD9fbopAarQ9NVsBbAx4
RlenHzgPqSbKebClLQ34eTYiI+p6NVQfyys5032+rWFD2Wbd7C2v5Jaw8JUjAyHl
VrxNgJXvaRBylF+HPkXNr1qfUFLwBQxdSF8JFHdYKko4TM0YROyqwulz7/JlqoeC
Tb6dXI7D3gtVJ9Dnq1dhgAuaiqOL707xTa5hnM3Crj233qCU/PIvUl8Bkntjlu3B
YbI5aBgS5WjZchueDmALq+mJiXl1Ap6159jINuoaw1uYKQO4ujoEKPtkg6YxMtav
R2noWv+9iHPCDAMyEPnsR8mQd+/3GX3euUBHtNQ3QI/lat80f5usKh91nwzPGBcw
orXRJqISWh3P7xXj1r8NZrDGZ4vmkgam06qfYDUNVusQjSThaNWqtzd4hW9GInRN
RjoDLRLwTL1Lstc+SY/I0yvto2VlfGYCAYtUjs0uqSXouxvbdW5RXweeZrXjCB+E
pzA1czBODynZY/7sRdSdbrM87m7M7X/+V1otCH5rMwR+CU5veoZBXgGwp7BMqZuH
Lo/QmXjryekYQhVRImpnbK20Sc6q5CK5WtMiaOYDiSANBZAb8S3yGCU/fJKsJAhG
YSboVpiEjsQTG/lFxPYVYHx6T4k2PSMns8cd05SDy8eFkqZOBh2o8Is1SiA6WZTF
czNPxgBMW5T0bHRORepOeym/0QeHp98Co6cKmFHfsKUfmHLizIB8qwPvIn4F1Oxv
IIMoqbLqMS03IrfeqFVnYt3z18xbC5HQyDWC7R4GFaENtmeTyb2P4as+h9Ts0+Ij
d6igDGRXUoX2zhtS+xuqnrq6er1aaxn16tMHRozljfPYxiUoBDsEGz0ocw8l6RqN
UE2PTnK8pVfuR6xPeUQaQWlrABQKxGFoVoHPnmTTx7zScKic9rLGaXist5Zqdn5N
w77Lymiqyrz/LXRunctq931Bb51Ejgmj2BY3do7GFhJtZHzIPB7KBvW8lTMhIV5p
2MkruXpHzn+3cOmwD2QY6qODmnjxGGSfj/iPJLJIfhs1v4gRTuAqxQmBqTzLOz/X
jpJRNJsttNJUkCSAOKI9oS0jqHHzhhqP7ikEl02UBGsgBpxW9dh+UzZrI97x1mGp
fBQH8VygaJo0G0Fm2peHAyjXCd11fRgFt8Af7H+wibFSfA4kLP9lnXlJfXWoRPP0
KK4PxFgjX5zYurIq87MKtdzSi2PXQHBBNBu6Am+L6T+xcYqLsjo3iH5raVLm5ISy
c4pZuDk3d9M/gCgfFytT4OkhJyewDB4LSKmzZcsyxxWix/zonHrqhL8O5PT4Ju5p
Dmfo0bU5xlK8uBnuTx9GHO3iQPRtMINr7J3d2H8kwj1GNLJUtERzeHkodkt38FtL
8oVi/XB98j+Bt0rcQJ8hHdfHzWjcq4OJxczPbqII/X2Ul0GjobNceKYOQx+7JAq/
i/ZXX7ZvShNfCR+B8QJzar7t+/L5a+yIHUJ4Vq/I358PdSR78TM4dnIKlxUziDX/
jrSDky4J8ZVbg7YjwaANBot7/NL+3fQKD0f/fD+lLNdzrjM9lHvsvuGPMZlWGVax
mgBT4RHzQr+Cn1yVSTf4BntfPcRNOYrkF5UxYUZRD/qDM8dbmjoF5ihN7xpCfhXl
PnIzID21NVDPpjk4sCOb8gX+TaHaY6LOuMUVjMs0lFEj7pmf6ZSnz2zOFAmd4fZu
MWjhiYso/ctimHHxWrt/nvLWlloRNfPn2vCX/v/BFIKqg7+zKKi9iB3qsmWqYiyt
THi4Y+ky5JPHR07BV8gzBIWJUAwoHvddj6st07YwIMv0aBUOXbOfXES0s+XFSuCv
3HVAtpJ0GNo8YVVi1fOBqv+QANqALRP5kauYuoUzKm1shv+PmTLpwaCp7iRHUYoY
q0Psckuuksfd/j4yWSB8nWKoVso75QOEwJzGOsQ5Hvm2IfFnYXhXaGmiPcyx9T2S
x+o0JgIXJB4UxLQoOO/YiWtQkJM1vg2Xkh9+qa9lgFy3uEaN5ngGyqFoR8Buhr6U
cuVxrvtmkYetSQaJ612Y6IXi4JF8mVh5ip2ckLjGam9qeyPJlt3w2CoPVxMRhnzb
8gKkrgij8vggec3FMil5BB2wZOa2EAbGEbzOzTMiAAdGurNepi9vjzrc8w6Tm4wq
v3QTA7ikrgQAgOwnfnHwY69wm2KyQwqL5GtkiYDF1FeY1LX//HuR1a+rCEVqVeG+
JjrdSkwj3vqKbB1C5bHHFVGdQtBknbWq2X9tBPMqEVdPrHN3ERBveCWN4QHuimPE
zVn6WiwCflqoojkZmH0dl31D3PEn7/fcz+UStYQgBOHy6fR5F/jliZDxuTS/B/e/
Gzv7IGmHEguxNgy99IZhmOPzRTrMYxRP30LY6ifLUobv2/+hQ+x6inOjWRrdrTCC
9ADBpToiZ6KluB8CjuCMXUkalgR/AR2y9Bn5stKUz80d2rVFRjM1WrdzOGw8+26Z
6hiqz5kfc52S6YDQjPBTJAHBxGTZIxxZZiU5ZWKfh2j7+weHyW4du0fAXdW047vg
hkFql3HuBFpuXi5MeNyv2DL0i8nYJRrsAYDGpTtj72JmPEHJIlqc5j4/70kHvAkX
tR82BKwLOJ4JwvJC/SdVXCO2WA6nqaxz4E9xtBHWL9DzrXsZw/6lWSxVQUcswAbw
g2VOc1K8/g4pa8oXLc5R7TwGpbAcJZH9LCXRM3kVB6kRENXb9sRq9arDDr8IqNGw
WqhSbzXDSWnTndkRHdLlYfzNidl3Tal1VOcLH7M/wqn2UE1/Hc8ZyeFdqIpYtYf/
yp4vpC9FZmMB/E3sFD2ubzt/9qXQZsElxoyt6ws6JOWnVExNjIXDhs/ZXjTeUvJD
5zvldPeCPAroLVD1CimdWpzXaCXDZwStjemOXg72LIvdUjZaMAKJa4EaBtRX0YvS
5H3qPH7sxMKOExL2vwqYV6RspZA/zoItNAATEEYGsX7L+5CoQvQsPXC+T9JUncd/
utDhOUpSVAH3dhFu/VRnffMiQFHn9zQpxUtieLJf7MiEdAGt/kW+Li8102WYNYwU
pNVwaNdC3KWr5Hgr6i505X+dQC+soNeQVi54XnrieF3sEgRxF8GIisgaQF9W7BtT
TRVSCUY+U5c53RoQ6S/1F74KO6KEyXTMmFKdiWOA3GQnBMrr5kh2nfiR4ftnv3lt
K+yemG4V9R02OZvfp7cvYI1+6I9cwOh7SjOiwm6eoa6Brr36wIk1Xoj0FNQGMrSF
UsBPNq3sf49ALzTRwP5m1lexwimszkuDvOxAErPA1+Kn0LeZmtjEga0tCd2iJTII
J5JI9CTnFadOIP8rSRNSozOMg2m0fB29H2/bWxtCKxSfCfL+hSLdMt28JACoTylC
/MqAq1wExy+xNgkevV57nOlmA7/pNeMiMmEekc7HKGzFRbKxIwdlKBCv+jZmTTM1
y65UgjB/o0OCzH26entqzANgmuB4UQ7AucCdX5eZ1HGVxkzVr+lX/YPB97PZMaqL
2Z1yQ8UlXgOcLEkG3Po4BQe5fIVNpGo3l5FqYEeCwrTRwiIfMGZi9R6PFG3c1+Dg
6ZL6nADbYaoscgOfFoh1sXFcL85QtrT96lwdrCx7pQ0R01di0KUIpTE3TWFsSKeE
J9sxgtnSdyBGJItkLO3kQdlyTzxcf5F9xDOUoObyBm2POtje5RKQuisiwW+mwM0J
5GIzw4EBYMkytXfs9mcWablC5chdOxHScvU1C44VmLoLtjGiUIRxc831MjoKMQ4+
dWn3EKlNXQvZ1PZYGJe4hYw2ZHEkS+MZ86Pk8bYcRInkyIaGzdiFgkOjktLD+lpD
+YqHpzMwMBe7YYTmfKEbTQwyo3FLkVXUxyDzhU6LjiK5MbAk23MuXYY7BattmyQk
nplTgzrTEg2jv/CnBvPNi+mF8JlOljNbNS+hW8dHt7kvHQ373yxxpFJhDqi4ppBj
yshhfiJFLEw/QC4ar36QDRZ4ed0Vrveg4JDtexVGtg3c+ROf04WPk88XaOm5lFKz
04CCt5jefmJ7WoVDqIEpNTDlkQVBsjRyiVnZO2dT8gkgy4d95Ez3S3tDImtEFExg
L9Nv88CEEEOfrpM22vWGYEJJYf761kNQu+OEPy+VKajBSP87Okuz58k8p7Na9X38
ZiDuHO1joINlrZWwijDmdeO+10Y0bz/p7XSPA94SGgDXPlKF2ll9ES1reGVrSZAI
9pzGzQ2seIjGpPheNYYI2cajbdq88lDNEyWlWkoBVWqCi9cZ/M7pwPhJPCWEywTy
B5OOcIaI9IaI13nGXUHoHvVnU8fFqOxvDTONoIrQtJvIMci2exfpeZUIOmHvCqkB
Z6no2dW6pL04DRo2EawsOkudI0hjqcVRBQUk650zecb6Dskaz0+bNhhkTG0esV2r
W4++SITgOvdOTSB/ZA5Y3RNFg5/c3LE1R0ZMO/O24a8CAX6uLGJlMPML7yjKba1v
+4/mpWcVrj5ald8sGuGkcJBSFBuZjjH11ltpOXIi3H+zhLp+68hMxOmC0CsD9Ci9
MnW9a5wsxUvbAZdLyQFqA7+VV93U6VLn5dFEo3Rgi87NdqNcyAAz3YL9davM+4tS
8cHx0brj4JOLNirAouQ+0UGeouINoGluVBEpZn9bDVH8ipaLFPG3GlIWslKyJO96
4q5e61LmEyTH0iIJmYJ0EohxfNBYmMwI7tIGsXAt5h2f7garqR47jE54Je3/MN8g
/OjF1DlZwgIlSheJK5QEl+7aTQFU0N09IW5k/Gq0QNchedHLBuo7wBVcB4jjhRaL
35hYAB0JruUNdZy/eaBRJQ2PA6X7RNWNicXfgRxtEcqZ8yNbx0kHfgHt8yARiqhv
xO7bScV+63yru5WZMhwg+4J2FoutQBeRXD4ezT//SxigBAUmkvgGbz9ZUMGsi969
nbkM6gDwdyrCSlviNq5AUI/uOcskaotvJmnIlowDznrBEeFEE1Krisj49K4MldTo
PIDOEtBotPG2s5MnG3NX5iKD8BFKmWB0z6NItbYnQkvJpI33hEE9RKRU+vRmFlr3
ddmdM8qm39XF0RKtarC8Gv5TX0nV49Gf1/apqnFkdp6iPlV5CrY7br2WtdB6sey3
Q3UA9JRHOBeSLdTvmRPXwgam1yHR+8ZDRQNIJ81F9M9QyBh3xDP+ubXelsIPNOyB
yYzS0Nm2RObIacb2oMhnQHu6Gf+bw2Y1vIHy2xld+4qDUvx7QwdjTRS8WGdM42Li
OTYYxnwbJ+pCasi+/Vn14eDV/uLZZHuEGAjA/G5DTjGkopZ/PlSmRcWDL4bfqK0z
AcSInlB4/iP30ddSXRQHtzEEpRfjgGo1Zj4fZGVr9Ow9R9i+GwOQdkTc7q8jkr1J
gMy94Bi2OLgfOM9T47PYzhwWRqvNqP+05dd6GdfXX8rh8M0TfiKTrwyXTrAilaQ8
Y5i4D1y6eXG33uxjbEtetnKly4JI4MLh1h8wyNu4AphKIWeGF639PXmj+PE5Hom3
86cjf+otn6oBpGresxxNWyVdKZF+lrlx6yQlJ/VYR7U2fbRJussZZr6DgYIFMIl1
9cczPA+g09I21p4j5Y96e7HFyGBxas5FTaggkeBgZDrj8j3S7meTfD+JpCIyGh4Z
6kOa1/gTFBcmLJ/Z7pdM0320z3YPWnZlVBnhLWs8xg+xA934nTleoQK3wUxUp7wD
9w9KrIqcernt8bL394auAbT7oQtqL7cJFmMG9g0OEaPY5g6wEtPE5Je5r7G7zQKD
tiIDVYpm9n0hHoJuNB0NPhk44mD+V8ix8qvitA5FLbWjCs8lbWBEDix4tP9V/8Ba
Hr6Qj/hZhv5zTVD6dEAQUaEME369DfG/JLTabz4AJcri0pA1wWVLM6hvhV9CVVdJ
PFxUSLrAgTk03bdUGcRbEYmM/9/ZApYPGrsfT99LHlzub0NWiYZ8kw7hOW6z2RCh
G/TBwQF6LvkmlCvRpaDsPJrKKW5AlcqdZj930miptE78gvqCC7Fl1g4QCTtybzvW
0RBP+GPVnww0bLDqAham61+NbEmn5jBV3Yzw/aFHT6r0+cAYDNzWed4LO6L19Cp9
B772z2Vb3Luo66HYtS2G1ujuvnG7nq7xYG1hbd615VP+QEnqgLxZ8/eKByEOBDDB
rtLKU8ccadAJOsAU9VVvS5cSzbNBtOfwX6CN9O9ExGM0K7yQ821csFlTKus8/dwQ
yC1lqx9eDqfD+FQXi36saUCm16CXYfiyJ3wvjwmRRzgVvkzqYK0ZSa8RubHr8gOk
U25M572S3UXDbtwmgMxZlZbt0fuwvcPPC7xx6UCNjC6lU+Fr4j63CQrbpTn3DKgs
zGI12FkZwK5YvN7GKsVjh1zLLubYrKDfnZHPrTFPycSZ79geAYc7jsk+QjMcYhNu
ROXlKQ7TMCyz5j9mN9+Z36tUmbAXnSxJEsa9jgRiZV1hmhRHhIAQCtrgw1zsloqb
nV1oYaS2OMpsj0LvEHNsz9HLoPFCrnCTyMMe6sA8svzTpFFDKBLHNUShGFda7QuA
ECowDo8eR6CHvi9/GNXQHS1v8+y9Dtj82iuWB0+Y3NxA/5cZtNneDoVBHaNbW1pW
/ri6Kb8NegsTUamP6a2/N0sBZp+fUA2Uxhvnse0ubAw9B982R6IVLCrco96cQ7t4
59mAUr7QGudjaNzkBb+Xe3G3p0B6AaRFkA2eZo3ir/7SuF+sKIGCfsHLIna1NqXB
i5ay8TnbVnVOrBkfg7WZx4BwplRFU5pbXfJor++fdGaxHkyJPWETHkHRmusbx7MO
4GEKRnqWD7eoB2s9O2A9y7uefhye+y7UrXCH/nCFGdYIuNByBV9Y1C1YEedqju80
vJ3Ll37w60pZmgfSqBPzfwJYI1pDG9wZJzCBZwNLlg5eGDNYPEWZtGdpT9j61/Gr
yghPe2qFhmHMzb1nfQzfXvNJ2XLuPjZUT5AoS/pFNuyxejPyiDVXtJZ4aE2gWd1A
Z0bi5PekvWsBL98CoY8KOkZRsKn0Dzhc0YbcY5xQcnxqXZz6cA8pzWf3uZkFZihZ
YrDcPeOO1lTwydKTA1/GF236xUBFAh3CKYS0zw6tVsrA9S7lOsa+m4W4JrV+E2m+
Ls/9Wk3Muvfg740ZMin8ZbUt2Jeyn7ihdMMWadyUA2CRJPKDpL+AtMXpWr8ohARF
/E8jg1FMzjyVB0t6zzdbs5DT1pfXyK7mdfq10tQNJgxvG0/khdd6/GWBrVP7txCu
zQyFZcX9aT/rQb8SoChqcOBfquWAuIYSq7ebtB89rcGPW5YZ0PuiZ53r9byATDnR
u0DJSvuMifP2GWa41kF2YkMj7/OTvdkaKnBKPkUSfDaqup4D4tgu1MStbLMhz5so
vbr8R4npG3BOAr149Ovj3BG2vBRpQn5xAZeCIyFxS2WGLEoJF4/NIAKMbgGG3Yzi
uqrZe75mnnnyliLLmmJDjWx5gAhNjIJEGqrAbQxO0hJYh3+uXsHRg6lxvQYqmowE
uptwYd9MiZ8+oQ12NsTGypA5K5BDCJIIHvsGHkznAJ+NXhfpbSqBJiuo/8fM6I58
DLgFjb9GlRMqhnMbcqXr37nVZSFOeXp5/L5XEBNgHN4yiilkfhg8UNPOv2+xaSPT
7+QpEC3ly69Kg+LCNa6prB/AzcWG8M6KxIWubFK+BLqQxGAEmJQ/rbV/T6HhQquZ
FmKrDTQnBXs9hBnG5CqtR74Hr0N7jF7of3OOGFIo7elWS3gF4xzAjy04Efh/Z/Qb
CXePz9nQ7wDP07cpOmf2jhKGZUX862o+sK+xzHO5NuZdm3J8vG2nfwkmobbk3DKC
DjPYjj1bIwt2nvW6wa3QGFf9VUT8c8lqrvXg09dXwBJPsMFu6EnAFnqr3TR7WVXj
bNxvhfMvmpLPdW6JB71kBFDFtyjXE3DpnXFjKp7OcPf4gRLKwnnG+3p6KU9kZV4L
VhSdaj1Evgo0vI2+JrYs8s+lOfsXKgn+feodSrYMLinj1zCFHS7yopb11VOTo0/6
QKWg1JtUW/ryANUMrpmiB9fGmgOIkiCyYvTWU2NGnmN7vqMv96L6l64iO/ALmxw9
EeFR6/8tBIN3JpXqam0KpfD5efhdJzZbEG0Hvefwe4/8QFg4cjMS8Gitxjp16P2t
ftsz+3S0iE7nSLnb3/IA5aEWPbd2X0p/eTEQ1qVkOA3tBJVV9v1qOykY0CauXR59
UnheM3GW7WGMHh+XfuiUrHlRkufeYLeNDXochy7maMFE2qEjbxJlhqAY9sQqE8Pl
Hf3wtQrpTk/RB4IFtgZ62+yAPXSmDLi8HjDKedxiIa0R7SU6guNkCUcqtn/liD+3
WUaBoAERtbuvg+8Ei68e9uMYiq9WkxIhKqqTJdvmuwz9ISzQ/v002q551m8lHg/r
L202cYOsxb7VGclF5UDeZSonW9S4ZGhw7XkvhoIKfqVg5D5jFlAkINkVC/baM2q9
KOhTUtDFnfHS5BPIaS6qfX/AeK1mZPVqzxYaj0BrP/I5fAxwNdm+YcPAh+94BjSb
imIN38nXOND9zYKcqib0ahAoSGg3g/MDlf/nK9cYasLDaFeOrtfLE8e4GKqOKHr2
Hww7Ja0Z/gQT6vmmTuIg2MU+aBvxMw5ZM9ROhbor/eL9R7j7i0W/oBuUUVBypTHa
gNNYDJ7/482ExZWs9horOBMwsE/3GYtLxyRO8B3Lfx2ESkBOymlUszfrtFs/tbok
7ePH/gvy3PopN71OgCnfDHd/0T1fCRR5ZbB1CdawU7ZbSJzan3CLE+xG4VzNQpVU
y2bc3SSldStHoomMwX4wMultVBNI9Kszdh7IBF7+rK18KaHv3Mxacx8WjqVuhtPT
yqng5HmInoPoEpBnnLBtfdpP3sG8HCQqZKOYstPXpIkN6nZrjmsVG6aq0VzdqWya
xgJsiGdtYjb6WJs1Fy3dTDf6UC6bilrlq/zjUrRAB9AKzat/wBAj0naNX5WLvhbh
7i09BuDUTuh4gCi1tQeN5V6KnsphrjaUynudRNoLtZ6xUwic4Td5897peqaBuzez
ignjSQkxYR9hEp4KVVnxMY2jnROj3Js76k9CZMcSg4oOsuG8RkZyiMvhTgsEJHBM
NakaJTuF4WIGNN1fzg/EeC4LjOi4XaFbDTu9SX7QaQ7R3sQkxUi3TyLOqEV8p9j1
1qImhvDeuuZV5ULy3Y3l1vNw/waOKvfoTgMfzQj+S4aFmpXGk5HejYHjwB4Gp/m+
HlqpeirK+TkyGM7py5Bzgka/lV44D2ev61go1VzqOfUn7G/dDsbxRwTism4/xYoO
Et3+4yAELrFtTDGYnEmreP6iuOdOa9nIDXUY/9DA46CbARYnQhkH2Qn72pY/Q2nj
5YZeMfWDxIw/Z4OwHyxseJKhUPWU6jhJsuabMbf0Qr1nrr/b6oUDoH5DhzYV75W6
pwR1xzlDczgPbZabRXWjsmE4kF6AsQETHIUy6v60CcuEspOexH6+behczRyT8y1u
CsKxAL6aXcjbIU8o4ETpHd1tdXJDzmhhDMUvAimS0kKljTnkmdTrwtQecIzpy1Wf
5ca01sbZvbXD3/ubhOJ6KFbGxQyGYBT++vG5dvAOwt/PmoNaXsQ1wbJJqret9lcK
yKgDrPhBsazoj/ua22jAGwPl6HiZhWD9wGk5pQK7VYoJ3Qsw4Fi38/f1szeHBvt7
jihHpzPE+BOAJF5JdggCecVaIbcVxleyYsakqWw/2fliJsfNfDccSmOKzCKR+sTN
Vw6+AgHqj1HbTPIMAgOiNo3yF58hMwHk+0mK6wNjaTPazT8kAznut9VoTVcWU6on
PsBY8Twvm3rjKSIn7R+/joqUZjy9ZVFJ0eIUUMxG2TNKyHPa0SLbQTtRyyZT6F1v
66ZqN0yGBtUCOfDPk+lkxXPjvDqef5rqp0jiR8XVncCqvaogEEw8xCmiAdAwN5+Y
nJv7IJuXiJ5PPR/vZ9lI3TjALE+UbX4CRzjZ/BdvnOxWL4JEttxY1d4dkaJi1g11
kdpnEqte908geOxSstNBW/abtBlvUT+KFNYSDJx7sFeNj/5lQymzMlJ0r2GwurSB
BnWCWxaOx8P98J7xrbWPuCSAw4854PzlBUZczh/qvIP4QITY7gy8RTdZoI48rWAZ
Inf2/umm6Ua9H5T+k92v/Vm23qWllwRMPNNEWrKUaV18x/4MEpMEAgCI227mneL8
OPGF/439JFfGxNAg8HuUjFta8qPe7nWgRZQPOg5SinDWN3ficUa+N1rLkCjUi71p
qi3DYzZ7VYfndGC3WcbvDZCHG6L/phs7w3A0DkK3Y0YTUlWHPcxDg7Lk3qJRp3VU
eYhbG75BZLzJ0+tSwDev4cxFv4fgi+eHJ4DWnchAHYehyDuo+AutqXQBSPOTgeo0
GvDk1DWRnN7Qq6+2obaTWF0aEMHvirLX5O5h6Lh4gWPzE4jttlP5wYbXo9BG/p6P
o1AjZQR6+JBY+OrLb0l1k+zJ0b9IDXUwhXwlaWt/tOC+AedKepiBFsKWvbQKYizr
itsS9RUo47GwrtfTU929KVxyO3UaCctbtosYgaPdwHhdVAFvHVgotFezUdnSOOir
eBxi5/XXv1JXSpkzWe42ZnUX3qzeO8gMDytfxik5+fDN68q/VyvMY6/h6QQ7QpwE
GwrwPj8YKXagvTXRPqsHs5yJGSgbC0jSVXm516yv2KBLjAsJ77T5s1zMcV0XNW6z
FA7czLKJKnKU+G/ME+G+wYGcTRmDt+alW0yugQkC8vKUTvCWmhBC1QcugvFn3Bes
kPGWlUXpcBnoeS7FoYAoUSzZRiUSByK87iAqJipyRZ3zJL04jL72oPuHpx8kwbAj
ppCcJQiT5J3dCg1SHE8+NTZmFlYsyVcz3BxHad1e4evK3oP97sT6S8LjYMu/XRVl
BUO8Vw0jAJ3B8R5uK7htoV2RaTq/k9Le8rP6FqT0Ks6OObmRw/v/2H+fLocpz1p/
abIFl3owAeyKi/sK2fuxfGnatrGNmzvLjB3JCh94LFdBghUoVu4O3xkz75WJn9vX
vlLXX7sDV1pG5ENiw67CzfsunB4D5ufPePKPJr10zqOjIUr3Kski80EFUQZbrRjR
G5jhVGidpthT0Uihgf7IA0iupknV6Wbq3eZQw3/pbNhcI+47iUBYTWgHk3Y7rm52
nMkzhWoOrjeM46DtWt4AFgmxlyV7rEnKBIBnbGjrSA1yKI450K0uVaaonHyvYzds
ka7kwgEg0FLYXYqlilRPbJ7rjJFI3wQQYiLR0qmBTyorUNyESyp77ivfJeDMRXy4
MbWX+uN1qaCUnkaatViBg8R9sGnoobmVByDkd/3HU0jblUBWbgb7Z3Qo/PFB3iQM
y6JPPHDPpnpvRzb34thwDyQeg+38fFm8c0paOzQlz8Jjvv0ey485gBvkz1qCqtpP
UHfgXsgPxA+Ls+RJdQjMN6kjg5O9Xx/Uh+96XlgDt5fi1AbRExnt2eUUr+71cliI
kMNTH16++soMDGAmGUKznhksNlzQhFmD7L1ZJLCWp5bjqB5l6cLoo2npDq26TE9k
riSo5ifAENMdDVCwr64MtD/NtLxYxGZfyfWNKnngUmEtP74ZmLxpB5/ik9Eo00+z
99pt3QA1cqGQfVysaLGNQbGwZuQfPyghUojN+rYLLBXZ29ngqLgWNstQhxraevmX
nhoWoHJFuCAb8pzMMtafjWpCwGHFRXmYP1ESsx0U2/oLD1RWQvJJYzm+euMJqtA8
14v1lCnE45soMIKfIsg8+p8R9/E83OZzd9ixHG1U07RAHdtLn9p1eEL51Z/1sN0d
ewyaYiY++yUiVDMJXwGVfqmeKkT/iaHEHZ8O7idpE3j4m6t9C0bEeAO1B8BUwDEJ
Ic5WhkJR9nZ4A+OLKYLxdVHHspx1yEePlCeDFtFQL9wdvg5Fw8L2GvMouLpU6JWM
mVIULzfxDhmldjZjmou7NlwOKVpUnfgqnsEjQ8eEArUHPjYrjAwty+1WCbZfxuHX
OYVNGw8LlPwkYmpT4EEw99han9ou5EN3gL66AMYqjaYwD4ADkH5K9o/pkcXJCDDI
RRGs+FmZ3BUWf35vJmYDRfHkhpconNca/8FG/XNlSFDVcbjKaOsSKVI4622P5cYE
cUht+JGvplZ4mxhMgxVtcf59QQpa4Bm/3xmQN5STKaP2u0wnvKgtVwA5UJ6GXkiR
AbADkJ8MaIG+WG5R8+OF2bdaK295r0A6EI1LvwCfKCFNv6CLAiTC/2ABFsDl9a76
N4Sp6ly81jecEDJpkWiI39UqXzmY6bfBylWjiNs2bch6ffoTGyPuJDHMKBYb3dMa
4W4HjgupUF5PQCpoMkKgu/SqnyFXYfaIa1Cuk8skdEwTYbvrQDP4gx3crG8H0hr8
pF0YIwu2MuPtl0WnzaR7/NuiqixbnHxLJQzJ37QI33WXAxZmHj2NemckLd6p320T
p9liJBbeNdQwjVuScaxMfR5IC7LC3Pa2SE4DWarngqTkuyquq0oErzbKFMOf9GAg
XCfpeg+HE57NoR2KArKzvUTuHsLqf/sQqavXU9ZIPlESKMTQFw+zZ1GBlXCvKmXi
ypH0nInSBQVHjW7sP7/XSJqlMKLDib6BREDlHIxuD8wSbMqI2FD7br6IeWYLHtkJ
sf0y8x4ZRRzc5UhlIjbO23Ta1kuZ3v15IfhSgpNuWPJSQa0HgQsLQ19GhnaOqGOi
jnnc25X+D0co9Tbrlti/id/c8iZ/pn9MnizK3Di+8g2i1Ej6pGbVLtm0FKSKv/zL
F7uoWRmFt+FAlszh5Lhmbi+jzqqAGO8lzCma3X7jrEearDlgVUcpGeq8IQmcnc9r
rJM5pcb9JOxkBFiQvFF1sZ0hmHZqKL0QFN+gINstBJVbJ1kpsDa0zQPe2tNkHcOX
sJ0jAFaSP4lGNW8gIlZ8+sLAfE75x6yo3R/eUzJ6/bWBRkF0aXQ4/KJ5kDuoJB6D
uuXXBABDVn9usRtTXsHupyDNJ5I8W19I/6OLVy2v4fBkyvr1bMO6VQ5iFXD/0dCO
plSWjNa8ITKE1iyJHCOOADdsnrOeJnpUacXKgtjJa8wdvsWWvdVRsvsL0qIsBcDq
5nsBMgw9H3pb4w/3qqUjTkpgwGO0DV1Z1z9LkidHjzRi31bo+UTdpJScrTcmpmom
Qcak0JTWFCxOY72unu+oZmzTwl9g4XpFqUbL4lOBj4GFm9ajwhC77yjpW9ZH2Uvx
F5Yot9fEnop5z9sBj153bXfoNIFpFAPduyVwuAjz0NUAXv+0uPpAbYntm4y00g5X
2C5JKfGtFy/CFrYH/elwh7819DSmFMB0hqI7FMShAbhSJlt/jp+rVmmB672IxP2Q
t4gPCZLC310GrZK+quagSiFtqHite6I/WjSxOa9OCCHYcO2yOttebUFzJ/Mya1x6
J965HWI+99V2v2ZdDxBfkcbInS3XTJb3vPMGIGQ85cEG2242BJ/hD1MHXVOk0Geg
aIeRL4bKtz7MQEaEuWBIRUB4/LF291KVJgQnWXNbScfpqGW0KS1MpzYhzxAJnvq0
s1SPPSjkia9DTjVjWorp4GS9dvFubKd7OWQYtmog5h+fr8r3C1CjgGjcDf5VWQqG
gmUoK/+lVHPKJGMjOgSwxIcQmbaLmNFk0kVZIbE9a6PjHYg9nwxoYMlf+o8OO29T
oOaJC4UzA3EN58Mf94zegQBf/tkv1dKO91kt+PD91GXzeYYw71osNo3WVOOiaJy1
rBeD3tUAhz/hRaTZPV9tssGDWRSgBOwGXi0e9w8TSwqcsfyxVW2fDVYy1A5CJ9Ry
sp2u7deFWjVjfuinmxYyPZA+A8+BJh+WPcERSAPUWHUtAY+EUGaGhM5sXS+SSr+t
bmvRAJOfXHa2cyMIz5GZEOVAsI6D/lD5joh8R8O4CmEdfsAoCg0ieIJ8yYTXSQ4q
dDGz8J/79ZN7AY3q0unUvZHGKQlI3/dvsvRI10pfqBpmFR+402OlopBktM55jqqk
FrMsj1s6tzJOHM0jFe4McmWk3zAfU9jonMHjIp3EkyHxzhyLD4rGkJKaTP/vutfY
odvR//EEGOGhriHZNZrm5q2tQ0n5iHFfACEa8YbplA+Jehm6bqN03F8sZzPJNsmo
VqLZ/9ZB52Dgpbh5qkG+pel72+ElXiupzTq48hGNZEu74Ec7dKaRSTWsXandImHf
PB28ZHW8SiWmsesxHsVfdPJU62hpIHFxxoe/po29/2KlxXMd8FWJ2yAFQW3CRq06
rfSphPhAlYGH1L7oPWcoOc68azhLWQkCdAbbw7bXVcykDT7kLeo08cVsTE0fAtbz
CXY7d4gvqmRl4+NuTqTi4EvczUcLZCm7/0c4lRzwamSQUy39CcUFzjdw7lDpSbC5
GTNF2EIu1Ytst9/oAH2vqhmQzGN6w+vWTU/su4n8Z4FUJpJFpZLqlUqNwpH6Dunb
VJWpLkBcovZtcIntX1s0VTpxs8GP2YDwoD/qToLfC+OPM2hVg7ilKaAwRGn1TBOd
FhnWenm9B2XMWgEdjUbsA/LFPzp3ybIPaIfSy4k9xec1y0jtFMLaD1ois09PbR/w
62RFarmJ6kITkOuYHMw1g9TfQwmklW+8k7VYQzmBtnX+O7wvUPowIpm4nV1YrLYv
IaiZHzDnmGnT+a6f9934046rVxsQ7kAnvVBvIAYBBym68SL/eOGlwQvttRMasx/V
980T8CmzCMuhrjmJIAyFkHj10zwQo3heY+ZxwzbQMuWcOA99a/oOxbj+J227QvMK
+WaNL5/dIwB7Cd+hQhHCX+NneNd01NLW6mTP+8WrF2D/3l3eXLB35YwXCjTjJKin
Cr3ntu9TvliVa3ngqMiA5TuFRmPdweuYiWxNa0xE1QYwp6MNCxsDiwev1c2v+qcx
/K0a/nA3wXL/NMftcWuampTV0+DojSMpPm1Geybv0kLlI1jQo0Q5c3RrNfxNRY8W
ECXzEeV6I9j+wTukTI0JcUzPoPMJ1yX3OUXwmQT56qhdmJt8N946iyDC6WCnqMGl
35WZf32QnVGVAcv9Z7T1ss2Vdn2cfKTN6vw0tgtHMUgaoJSWB+NS+C96LTY5blgs
GAimZK+nVC0+dWILPRzdX3K7A5DajU7cTnKkNehs/IEabOoB23zDyP3/6BrGdmbS
ybFZ+3I4tv0f8YldIyEEf/X9JnuAcBEqsstYYthoDv8bya0anPjfyLj1wWGD/xd0
nRU4YwQPw6j+MWiO0z3vTGRId3Gxx+HPSdCxi7w31jckEAvZdlbV0spSXJYQ4dlO
J7IA9XGBOlCF36zMipQi8K+iIqJPEEPOGltKzxn3qSzcanVZpSNfP86AAQqv0XdJ
Z7IWZAwqzpKpSG6fWLxpO2DRXxX6N7Lm3ehu+4SREWjB6fHi1ltDRbRFazggICVo
GUfxjjUcj1j0tpLryCkSFQ83RQr2z6cj/nQXuK5VGyxi07nqIh7t6tNIukQXZZBW
ZoA0VQpHuRBb8hQDDDzBXDNrD1PX3SdO45Td6q1XeKni87OV++COrp3M3HdC2La5
E7nwQaxp4rI/7H/7Sw2sO+Yatml6abHMCvLZGT0akrUvoY0o00271cYgAb0f0ezV
MN8dUO7IBuVa9M3rXRJJ4KNvbIsClp8QQ1WgiO5cZceVmv+MkR4148gWYABhSewU
puurOROuvU9N60KyvQkrZGTkc+SQSPoGSE/aqrLn6cOZuzr/BnVTaHIivDQweYc3
KYSeBenKKuI6NTa7GDdT/BVjq5uGhvy97g9sNSXzuF5TaQ6i+XFM8cP9inpbGJgX
RdESEhrcnZ/GqCfRl6xxlpBjibJTHNVkZluQRz/lM8VE2O6idRhZkvaVUTYoYCzT
26Yu6GFFYPLjgrI+H2T6gCEuEQWievaUnIAwyh/r8Qy+tbbaJaTNp4nm0LMzWE5X
ALhJcs7R4Cl/RibFGZhWyZQ6yk0+k3xk6pnpbCO1R/JYNT/20zX72kKkwuo8G0cf
/Yvmau+iEDUXX3fXkMBtDAX80W5699oEwXDcrvGEsROXUVDcqDfxbIh0+5ndI6iF
ZaFzAAYC3A4iizpdxskbycHsV/cTXjOhY/w/XoYA540Y4CagXKX96gbzKOIBKjhI
FN+vjiw0Yuya/1RkxlYtNLJJ+sxFu4lb/NYqhrX7eaVvz/bf02q08SEdLrMyMaY/
XFHEpyd7Etp4+3IODlWXLdUWv4f2y5UpBn9a8dPkVFpAILgOJCXeWNIvMuaw3K4i
bGAG+ZGg8SYc+2qfZyTudSUUipJRoHeTq9BobGYjcJdA2eK/MDx2UBsni0jjrhFr
PLsTRvF9sNer3idPWHFySnk/oHPlYy229KNuhhOZTWPPpRiqMtt3bkIXBZNQH8tw
cIC8n4Ad2TBx8a2K4Ri/9b3M9CoEojqwh6cl/Y4MHWJwXSBL/wlNTjCyqWbn/Hg4
TwUJuKUEcnVzg8f2NPjuURj5Xl0DyS3bZOcSugX1qiQEp9cOCBSVA4pD5Ch5Y/hV
LX/rVLDEBu3LhoUz5FQr5m+5KDOXnxt+q9GG8xB2+dWXcWnlbPVTFGI6XE7tc8jN
+M+ujRpOv5WRSmqlJIrh46QOXy48TY3rg69ke+Dkv1tkfBzcaEh/2oRY7kXcDJSy
ISfPNrvFjdvadeD/ZUaYyW8MUBKcEQ462zgYCrJzXpSU4USNlnWQyCjvk0aKs8Y5
1y+J2nPm8rAvBCSfU7JGgkv5RUpHKlPbVNNiua7jBD7bmLUdt/Et74D9JNwXe160
byCi2ox9tdp3hoFQebk7O/qwhpY5EqB3HV9CfQ3x+h5AGyElQtyYU0O6oNWwN+WQ
O+H/8EAeauXUdmYE57dcAR1QMjopWW6Bj9PEjNO4TbuVibszOZXndGNB2qXQJsQM
8UT6ucdssY4MQNbDL0l9UfV0NchfH6u8/cdpkzHMkHspBgq5PGXaN4woSGGOMhkm
dYsUIIHPSxqLssJBtJTGOU2E5286q8cE13+0cahvAUMMpSyq9Bo0TMJ3dPTdX5oL
VOJdOl3jFCrnkPcBEv65GNDDkMkUX7nJ3csnNMFB4p/kIXM1kCk2Hq5iVucPp1Oa
ESnYosTVbOVnqf0f0mqlBaeRU6pFQw9pjRY7Lcn2EtM4Gkb1UN4HjCBJfL9E67IR
QdNfLQyQAdulqILD3fA1P5WkK8nWtthmrGdIkcK5VpjHBwAAD18mwLsC1SG0wbw6
luYxoLWEokC4pt04PNWEr5CjGrPUw1ipQ7NbDTGag1fUviqUC+Idu5/cyXr+5xNi
oftm5WuLfczggq5dVVjA+s4/9HtynjiUxrt67bignnNjAiIQn52xZ+IHwEdWck0M
4IOr4HdYDs8LZPrsfGJHMErEYXvuekrdcmAhCa8gGte5p5EadNp9AUH/40WAvTK5
iwFJQcOI+Vogo+jGqUslX5NyGdSQWcGngBZ1ht8yU31wrW+2PVnPd02HC41UoNK0
QVGxsExKsVk864Jv29L5dcMM+cI6GoqVTcx1rwRC5EMzKGoKMHsP6nAL79FcOART
N9dC3vRPBIo1JXD0i3UeeyYK2AOMYpe/d1BwMG65TTnrr9bNh1Wc65pAT1da5k9H
9bBmmczf2O6drLjINRf/nSjiXWN5p9fnCfRuiSkbpiT0+OCHHgPhONdd8yDzVNHJ
up4uoD5GSaN6czWmRo0XSazrT3Vr5Sx8jVqxx9WuaoKxIe7dU7DHmed0WTRwCT/P
tbiFYPAhLAcDK+ixnq4XoqqXaf2PYXpREeRjkrWHBiID0rZSaUQM4ZrsEqDLGwtq
B1IW+OzEqylAMjZZE+iZyFBmyUHtow3QpXXNseCgsFP4ZqKGNSdOH9/bfX29hepz
86qfnMA0X2pzHA+IOiLdIHGVAZlI1kjoaI6kyPrJd9cc3uKvrh0tP7MZvjPyaRhx
81o27LH1j0dXQGQ51D4XSIv+BowEsKF6aqERvTtfNulXOJ3JMsE+Dz75iQyS1R5Q
ZqiX1JUk9/OzAirQgwQGC+1Dju6hkm1kQY+2H8krWWp6tkLDcQfXdH9z/qvfuZSu
RrSrknCglOSerY/3WJC1QNSMi2alsg9ASkvtOY4IIPeunz0dVjzO+5Xeh7RSl4fh
hZtdLWXli/m5hPeKXm8NKy0CPZhBkPVRvAFm++uLMFODx+W7D02u+++PRL/AfFfk
XjVOw9ZyL7ze4/KC5APhUyJt/YwfqywNoJIPVupxXIMYLGvT9k+6WX9L2BBiUXiZ
NwosULCJvsOySdopPPCvTc2qFkX2QxTU121vCECxkJLhp2G3n7S4LdjpHYDq9GPM
DP7VpG4nFnuviAGQSydXr3d93OGmICyA/6H+fyKiby4th2/UlfVtMbKr5syCfeeG
hh3O6VPh9hpwHHEqyrZIsIVFEZXNOKLllWMj2BdbjBugW36g99mpMkjJdVFMWfTL
8yL92HcCx4PX86keAxA7ID77VTL6y5ojWqv37ACzFlpX7khsEzH/B1Tf+EQZkw5S
/PlNIrJH+GW4DZJsbCTtd5LSe42kBfCl0naPA51H5Ux2xZAf+7/LH3qNGAGbyLfg
JMCSm3lW43pYhBiXqb/745wH0ip6LPzpSaec+nU7dOuRkJ73dRU3gjQrQ8t6nezs
62PH/qgylNriRAJ0/MDxvOA/hHgSuAEuaZehZMClsLXcnqJFhqTiNDUUxgMdF7OV
nuBlMHqnMBSto2AntfZEuFU19ipGvDN1HgPvHs6+5hW03lUIp/ZTBzAKL0M8JxgQ
Bj9j9MNw2Xc1U3RyyqlooWc3p0kpM0X2QRb4ToRUsFQeQJeFM4LFyAm4aCxJqoof
FPi0A5UGJwwiGDn109wMBhoGMIU3BXRLq4GICDCf/fAAgsvDA3SZSjEOiIy2/Dtc
ttDvVlRPSIVo5xr3WNOVYg8KtbZ70POwv65bIDTSqQ4EMkVbmO25EidfQAx/tLgK
h/4IHz205yR1PYes6r9LnMDpu1cH687k5rYTl9Mgn/izTD73PU8RmXT9wb7BbBYb
DmWMvkWTIoSzhtNsKJ0bXzIbOubi4eBPC3Kgsdzo+zn2kqfzDxKkAXNvMaqjM/5h
hSCOJXRy7LENP/We5lAAGiJwgT+1KjZC1hv1KgehsKSAZfs7UVw0Ru6Zo6L+1OVV
MuwQgElqZPhsBFLVvVum2IAgCvk8d/TUQn34SVUYzY2JsQ34K8J9+OsPDr4ZL++X
9joxdD50uNYHe2ablpQTBN46a9noLbi53ATcrwady2+hjowgBC9SwK24qN6YbpI1
r5qTBWvJNqX0wKxvdXwMzGCYlXL30bpz96FubZGGtpaybhIqHPkwRCyUYeutVK1W
mmrJsDu8x5IRxgVc14WzvIqwU4PU+qJdXpl57BRRmFooId1O+VnUaS2vbp8uAKD3
KX4wY86OCQIkHE3goJklEr58NPwdiNbiFDFkZh0/2YcRqHiGjfVEVjIzLG4QoRsp
RlXBfrNT54hhc3wFHsqKGKL6HGSVcxlonfJlq2553nrScyissgKcm9ADMaCpEa57
Mvnwu4a+YESj2IbAq84YOZQ+3BnFz0TGCfuvpuJr0mHbUF2wrF9YIwj1WWyy/vPc
s7TZAfSKW6U5E7HDUUCxzBtzz+NmRHlwjWPu8QPoBt8WRHn7UUqGVgZFUmbG09N/
UA0yp7mt6TzzXXCB+jySbb5lXsXdw6LhtoIB6uhlDzrbibHB0X9D8NQnk9ia/jSl
x6mhoOpw9hDIng/eqVMcR3fmrr6P6ej6wzm9d01k/5KFb6Ng7NvvviMG0cilkj7a
UHn1dVZQyHASyKp8WTu69AjnFUlnHvdj0WAiyWEWaqGW4JrPCOURz176xaMBBin6
XhXvLq7RNMVXV+L9mjBG2xic67CoIZQWGhVbzwv8NsH7lW91rC7Suc+PrXwkmFbI
jcXbge+NA5fCGlBMBnxfl8KeSh6YiexW5J1n99nqA6ss3z3QGeQ8wxVWcvHSQ31z
V2DqjeFweZlybhvHJ/bGeUdb06Mi6pe9wR1er8zL6c3iVztllS4t7C5Zk7ineoC2
/gZR2hOsIdM8Zr5Uj0rqqf3KKSIOtwoI+bN7q7eLgEP1gNwt37XjLT6Ed+PKbypR
w1QHt7X49/TaJpR8ZtlLOUd43i0EB/Mx/rXlLputLEONSJPgfSWq07lNSKlrOHmY
o3EPu5vXeRl4cCw6gW0gbPZMWXD14uIfHUZlArcIZkYCJUNfUDLm83Th0Kvk1AJU
FB0bwOMRVC6uqxIB2GTYtA4S0ID0YC2NUzE6a9UOzncAbpubeDQeg03M2RmebNvg
GYqBJzW0K7wv2KBMd1aC9EUo8USBKMcdm5BewY5tWCuxBPCLTT+8lY2e/ofWVHui
nDeoUrdLmi6+4GomdSDEWQSWxsyhic0x5QssBqVgCPRg4oa7QHT+68Sse5ICjAC1
2CEvcmoPVAwJoamkvJnSpMO2uPxu1pg4+BO4RSEZBYJfOGtoW5occ8WINOgDGnH1
UYe6dF5AIMpNXwspuI7RlyWAq/D6QhMfRQ3GlcGlchNHYoxqe1nqW+wWiGmCxI8i
pfiL9K1rwk2DBgmcsq56YT3adxBfKI7yD9n64xMw2UKywpBYtDW1VFSgQm8U1MUh
61kp0gwVHh8jnpNeybVXijfgM+0bwANWHjuYpkDpLJqXB7L387LH7bqslfTEzYuB
+Ji72T+aafwGmPoef6qeFbw6IQ7owjWevA4H+YY+ytMg/gQY1jT10bDhpEcflXKN
mahm5yb9lKyhwSTyw86IVaEgxwADp0et0/pzq1OMm45gibpUl8mGPQ3vzyP/lu5J
YScGCDItnXtsjJQnuNq8OhXvhxe0OLpcFIfmhE2OcI0RPgBnz9dt1+i5duQpO5Xp
02p2p4g7NB/aPiCWlJuW3YWmWNIMbMHkVdFCvuikf6ox7/4FQ3Y2X/+xIbx5ltg4
T8P/WXHH3p1ceScZANj0HyaF0fy100VlnMk+ygEgk/XkithM+A8uwJa/zSUxMXIN
lFBnLgKvPUSZ9GSr4TPEo2vaXNXhD7zK6yuIK84UbMhxGJLC6/NKmGKJCdDE/Uv6
ZmChRShLPMGx3A9kZMEqZ2gQs4AL5PUtdSqUOuDiGrhhNH82Q9X+xCEA+QPo/Lpd
9M2HykhCxorXMX5zCbelq51wIb3hVsL0/QlR/mrkyUE8sAsJK9i75EXxi05HuC9o
Zq1FN4MKON/M3z8rSex/WXEb2c/aDuzn5M/5IboVyHJUIOGHWc8jxpYT8W/DdMIp
+RcjdQCRnIohn7Qa5Sq2t5GCxWrNJkiCaUA2z1NfmGuyQC5CZghOGlSvq3Jrfm1c
9yASRbU4GZhQJet7F7zC0RbTk2qmYXM8cAbPC+th3z6hh9WNB4SV7MS+6OI2cV67
zZsOoDdn5Nub07y0NKJRw7i6xTWA1gzs5o5a1R/0n7Wxa1ZoOHEBSzNSpjfZfNud
hT/xQv3L3ubdTUaUyXS1XTeA6vQlxtg7zRKPNepjxJ23uVo9UlX0gdoY837Bq9wz
lJ1iQqmPlwLrmYksbEzcVLcTX+ny4QwsLLknAAKQzVc4M7IYNwsldkhiztWrCCeR
euQ4BsIaomGUpTW0D6K+ViLZcQk+iyLUJvPc0Eywphx8KxRaYxrTHuNcasW6r9rf
zZVmHaryq+5tFMKPuAdQVFjOPksTPXXCroL8e1OGhXsjTT5QEOHU7CEZyybYqx3Z
iqg2U0peB/3UX9dHXoxmta1JzHOpYeCG+khLPef2nbUp4XSEqXNVWU3skNMTk2bU
a5mSqXK3euKbwos3IlPvkceGLZuUy6FQoGlkYSbLPSxgkJaVOz3eneRpLbpyJbV2
Uplt/Z+JQa5XiSOngnEL4MgupO8on5wXApZJaVBaA9swA5M4N2AljfP6IzHPE2rT
7B2VPOhuEcr4QXsBoPSIeA4Y/KtOp8vgUWg0a8Al15ZoIp56oK1mjTO1Nk15bR4B
PW3rijBJPgVjCYB2EVwAbqKiojbTZ/Ku0BdtSXEGLEVHsFJYj9uraL267hEXrbql
OKdz8YSoK4CrLhpyxrfSoA5DrGb+DyQg3Nxcs3Mem5zfyDejFNJmcI5W1NR+alEI
t8yGbnqSefNCBMrAQVQKmCkmqfZRoOu/u3xDlGl5R0lZA2rb1NXDFLjc4OHFhdml
8nnOaVHx5bltmWoeo5NW1BD/BBIL04U1F4yw2nG8+QyMhA/5UoS+88NQeJK0ah4e
5TQTECQxjF7cTQf7UQuxxLm0Rk/G4SWC23bmTczIMrs7y/xTsJVPH7f5ZgQPutlY
/UEnCiIi6i4oZFayw8UlK4whqEbjM0h15QLy2KKx2io3rmHYp03pYj2AoE9jBdc1
v+GSW9PSw6cTj1Hdt6UzbDsBTOp0cZTCgeYvXaaoEwHpFiX2GnKV7feujah0nkuz
nYcyfelxsIAuPwEOYE/P+JKAr90YvjJboIgtUTf7UNaY6qMOSeFF5DRdyybM1gOD
cotUStHK4JR8ebbWjfZ3PGUlh9mUmCk7hE9h236aXiJEtEAzgKFXLy/V3wg9buGJ
Guiq7kY6srQjH96N0Z4VDebFo60Szwh2qxTeYqDE5DV3084lrE3kKuBrcqzDvbIv
5gmYJtDtUaG5KQZz7tgJFlq6iMImDNTVIMyrHFzbf71qPZ75cUwI2DEAKuCi24f+
abZcVOEplc0L/d83312XQiUjAbUDrkNrBb63aJWriK1WhgflJgVkeaasd7N/rkn3
btsTaH1dOoJ+dmVrlTWAMbyqIgEh/fMcHqizZSZBQTWxEb9bcv4kbt6nlR35uSFI
C1OK4t8POeu3Bla/lJuv7niXtaJeu4gDiXcgdtBmVRyX2Ou+aknnLJD8YqinEDd0
i29/mbLua/sZyqbPJWqgIh7aueDH05BgU5OWyJ3sPARi/kaSQg6TQ6sZOEpBetR1
MeFH4WZNA5Ne05lGLUBPK9onq8+Hz219xuBl0J5/tToyM3IhY63Ps1BPLh05tpQv
/j828GvkVT4QNFxGx3gOPyO65XllXuOGHYtNT3CScm2fIN38PBgcbL5wGxiGJgVD
QNimxYJvnY8HeeS3aw8OsCZb1ki+HkVIAOzljb/Fl1BlhH+gz6hSExBfdDphFTgi
CA3d5ZHBt6UY5mAX4dFlkAUKjSRjX1TCMQ9m18lEeifuIcVaDlhCWRSsSeJtMZ5I
Mw8DaltPCjvvnni23W8hqAz/u+ayS/e0A9KggaTrZDKmKP6xX91oxOAr+SR+ba2A
t6wNpqxIFeE4CiVWu83HDs857rL3LGdAl1hvV5UynxeCZ3V85DHm9x6nGcSd+15X
Pl27CTRPvwelwLP4ECg5WYG0uy38dJlyBizBTOCJYkIMAAZOq0VLGUjhtNS9VuKM
cATm5fOEUr4808eHcsynu+NeddtqYQYAptkQpqFM8AaJwMmbp7y8/KEZsP4xLjvJ
AHngo8dnTE0yafFyo7Rr/iJhamyL6s3Bph1Hl8/W3YFTYgGQ6GgCAx0letd2D+aH
aIGpxGiT6p3P91YMk7OmD4sE5UwenIBm2KCj1F61N3UMYyv1rPWNozrgrvGG84Es
sdJdn1Wcyz8v907cRHN+5+i5xx/kzXmJAtN5iA8WJCfItZTTo+j6TQybFiLu46yl
fB0HcBglkAJmLKVD+p3uzZr6eAlJ6luOTg+nuivD3usQ12kbotbynJu7t5dzmJg8
8kY7MUfrYOD/+mWl6mMUnuhadvrEX2EeY1tiBTH5akSTXv2Erc/VLbkIxoZPD1JR
LhLBincNUlkKF4wfQNl9Hir/rZSmcT/Fjxq50+MKwtg=
`protect END_PROTECTED
