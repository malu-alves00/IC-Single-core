`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TUbiS/8pRbme5cFUsvrjREETQhkLfpkSGlJK74vL1dBxsPFYt25Y8k52d+b0TS6g
8lYawRoFCuCY1neo4deYSVEuqVtWY3qAVOcTl/uXCwy4rGk69rDPxD8giK4IztXk
hOJ+n6aD5JhDcJ3hFlss8NxPTUZD3ht4IW+J9HAyikFdPUxHYnfuml5ICCQ6fSpI
z5nw8vtHayJg/sMprVCCatYjaRO4s2PjEwY+pO85IjvSUlPzlutQW6K0IAh53eTM
nsPeRtAB069nXPxhf8/91omomPG2tHfaO70KcnHN6Ooc5Q3MUptnU5ACwp3oxl+D
xAe6al7kyy2B8eTdItq+EcE/GqCsrI13h70Wj2d1OndmwX16HGcfqsJo8gnPjxDm
5KMTwWW8VuiHFwNArau/01qwO5d6JMOzx9cfBkYgQDbHkvxkC3Am85Iww6Sk8v3R
JxNa13Ilo5qaNBaMeybKC8KbNKCgCA2R4b9svuXdIoLYNVDevKr6ajur4+vW291Q
2ZnYgWcNX1WxU0GForcRjQ==
`protect END_PROTECTED
