`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iweHVh+aB2rJhiVsnsMh6gGBE5hngPCCYypQI2WgSNazDMwepzyTpsEYLiMng8SQ
zaSlZUCAAjA5GF0gmYNeaixZzixfIJsfvymJ62Z2hI93FLSjM4vzd5FAv0IPLi7+
2acAOH4VXIR6naT0BsUvL8gmT32MYKbUxp3v2p5RRCrE18hFejr3n6AtBfSTr2Al
ZuJkj0RD9p3M0AUAYVaSIC5j14+J+SObIUcGzJJma+wPROcc8VuLsgf3Ghjdmb7c
9ZiNhx3GYjNudnOsgsGmh6wAVYQTTvYFo98nwC82GFyErvBcY7St1XmeSpd6wY0a
8XtxmDLOu9g43l8df4V6stI8Sf9aLLO5dXYafPepWU/S+TRn5DNZryNdmWjX5oJe
mV3aT/DggJmDQ7WuW5Oxxiv3dzNp28kk50BQMW1JODe0/ccCKdEbXRioYD9//ilU
O2taxaaPy9Gl6wCWh1rXQzuZl2I0EBJz7X8jmyH+X5tbXPz9tqKUOFGC+WUoBRNw
frts0lnarYKxZ9zXnHctqcG7QE+WraBLu5wNsxjHzZ/HWCkcFBfvK3DS31rG7swD
+tJN8w5T8NuH88bJXIbsv8h9SYGR//NDObQR/CoKil3y63A7ubgCGCRP4HW+ruQn
ybrmcp/CQKd5nssDTeFRHRbfCJ2DjeIyo+elKqhHfWL3O6N9VdO8ehaXbfnNqAu4
+BcZJc621vrHhRmKv35XaeNWaoUefI9pP8vcdr+HwRE/xIwu6fqcYXKev+3dK2wV
kEEcWRNE0hDyY0rzAoJsUA==
`protect END_PROTECTED
