`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iDpPbr6r9x3Dfp0TP9SOMwBLcuIYG8H59RG3jap6SksZ7jVuurVhoEFtv1kH0vor
mYIrIdHB0NENvNF9/iCXF3JtujOoo1AV7Yol8LOyOaP/KXcjl87wwDdP/nvgW27v
kP6zm3GWnOK0nm9jufI5JggYsg3RMUSlI3VwqKxeZcpROH0yKw6meFHCq5/LvCD0
sjkWMeieemWSKREG5owB2WBpHL6vHnurms8OwbZxSKvqZcszivy0z+Bnuk7BFv/u
HTZntPez9InujasH71dcjGNIKskDGdR2mmJPCuF20ef4wQPIQQewM/3rAuy+E7RA
fztnMTH3VCTn1azFSIsyzXVNaDimMZoayz4SxSU8jZ6CW28isbgy0byV9O1rsX38
iblVhgUvV19BztoYL6k4/tlIyQiuNIuyBMS4L2xPBD5+vZPkUumjESRg9XTC2rIp
hq5VZqr5uRYri4EZat2OTUcA+IoXBiDrGyFNN+3vUEuGlPZuP4aLPgZgXYApxL4z
SD+vaUlGaePZlTxYKBjv172sTRF7B4MuQFOwfJ/Lxnxd4+aYwmLFomoVDn5hr6G6
WyStWZ3en//2Wj2SMM/ocKj28vIZIJS4vbKCptNwDmdNT95gVjjhzqGPGesWqcTc
A4m+ktpjf6HbI+HgmqyA5UDKAkd7B2zmV3cgYge8Mnq/zUiN42LaoSpjaQs8Ggbv
ycmTQ3TmNVOhXLn0zbzTxNPef1xTeoFbYLAWSeeT2oyD8V7hVspFBmCbW7VCBzTk
KaTLrJtEsJPfB2elhMXX//wPdxgWILFvXaLvOHEfap0sf/XPuVyrN7PT6KUci6QW
Z6QhaaSihL4X850dpIhM8SCStBQaelMvwN3y8vdkEu2CWFx5KS75N8vkhy82PFAh
wlEwtOUJs5YMB7Hbu7fZzOoJbvHWfULVTm46I854cXH01eo1+KAckne0QsSpvjrE
sSr/KwSOJeffVWwMY0s/DwLkA+iDTNpdDY1iQScsquRMnjy0MiMRNVei58ULBoyt
/VfgvwXv6lzl5c6qVqmWWkuVKfHL0XcGePP09NQs6IxXdIezdEvLDTEkfMb7hgYE
YaOIwMfJ5sSMS+qFlkIZPWlMTt7+n8l2/CkytbH8xXZVKvfl83/aOIW7f6nlH06z
c//K4Tc0FNGtYFvFPRJ+bNAprSP8+zQ+tAUBfSdE5F/8vm87WGF9perw1BBmlKWS
DGVWydFh+3EP/LK5H3d2Fa4REMsTSX9uEqi9Poh9/xMBut89GnHxOEryKC/Rltjb
iKorlLucJe/NkuHFPW0Pt7SyoI30YjRwMs4j9wIj7TtSc/wKVjDzIV0//tqw5Ws6
sV8cQ67Ond0YBhFvpZp7CfDrPTr4BjDsXyrGrHexdBKYuo3yapkItKLsV9hO58Ce
l765jKtiGpd6f8YeIxPIWnLY9rcMwdKykL1YU63BUdpDGNh2n0mGhort+1h9lNXM
p2eOjsssvHivUkfNIFDZ6mzTSel4Wi6CmlA+BSH4sP84ELqgC3MY3SvujenCOvEz
FJmSPWQ9jN5pR3lokVsndOQzqcAGwrRLNgR38s22KWNg7+fjpB0KSwisHu6XtVvp
bas7rFYza5p/dxdTDLFq0Si6ZsWOQ5bc7oHgrxa0QNaVazwKNedn/c6HU48Z3+BH
0k1H196MYyO72ucFZbmn+Udau2Dcc+XAXkfrKLeJLkdTk5Whahx6O860NfGwuRs+
OGqwkXik8myu0njHxQ3/gZchs65yyBAnuhhbyHEWLZ3SPEK2WYfJAa5qHRHLDZwx
ggZHJoJjrY6J0F+MSjrom1AGR0jnlTRHjiJyG9YRt5GWwnpK4SyJ1Aa5n2zPzm4+
h1z4rVvXNjFElRmU1flaFspu+0mfrOMt229VIfscQ4H3pX0DVAq1FNK8EHFXnOnB
66ojfg1cTW/rqvCdoHiraCSILw/H35dR+U2K1Zws3otgpKoGXrJl0eaEoIBzxZj8
DzebELRZLnDfpiPVIuVQRSbzKD07u33yU4k7WNDpcgKEw5nonaU7ZdJ/LmE0G6Fs
ZIyvEpg/u7HxBPzwLtaciaJ0nYtRaHotYzFv3CjRk+PIGKvx4KBeR8NwpyTF2kKO
eWg1QLsTWwXwyxDf7rgOW9CeTKvxWj94PqsH3XMotagZeEngjHpH7NSHqKt3r/Wd
oeAHoLTs7aZjUzTRXCJTjt+hqSwXhtkuulbYpipZEX7N4TSpFDfKc8Xsu/6UAcdr
YV5AsrWck78V4G0ZgAbxYHK2IsQTGRvV6OqwfPwlcdHO5+JY7yx3wbKvofxhZFOk
Sv38QhbfBI1B5gCadSSJjyEHXyy2r3CzUA/VVpJknZOI3PXkl0+8PbRRTYhfr89D
oOI39rvf2sHKbuYbPnbbm4AhRxMO9knnuDu7b7FTPkWKuAJmq8oi7dFJ2yoiKcHn
+4Yq2dwh587VXH+AmmcLPYl/EcGi+tJxB58N/MN/nZZQsF3O2d4xLWI5zYT5nVY6
97sF4Vte6hs3abVk2fHoRdIiYC2vxPzYxo5Shxd5UF15UXiu54bN2sBEtKR6SxyG
DVrnpCn8WPlZTraTFOwyvDZRUIaaCHUvgEbXX2ukgUJqOTZJeyVyJHP5J5TNMDg3
Ts/7GhrsECnVvTHTONvpuJFsghggT/FSidI4DV4NaDOcYpmbBYqaa23fCmELYMGm
yWd4YCuzaGbIjqfrZ4MPYEqGJfid3gucHxCWNjJBblXJTmW9q28a20c5YCYdHWJK
MOaGVKe0umTA/NHBKXv4s+EvqFZlPgpKbI02dUz4z2j2qEaBjodLRn+4Af30W16A
Z+JmIetTxuwZ97ZEpZTMd93FJqdwU7qkUvbKrjvl1fxnjsqk+VObw1d+gF67A2LG
0qmahKAqPADBZj6m0+vbjh0J8bGtZJlT5hy5FtY8kJsWEEEWelw3F65+CDYpqNGE
WxbzVqVWEyS5qcHNBeqA0mHqYk4mv0P/ByBmw8wK1F4KVy4T2qGcLduRsNKXM5Go
vCBQtzbMbC/cZhoQD0LbKsmyIzhMBrk1w9/5W8slAKs=
`protect END_PROTECTED
