`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0UsT4nCbG+z/cUnkvEEjRYzMWMUNx0K6uF+FdKAhrUF1jrhJ4Ac71nQMEn5GU80y
WPe9LmWv23n6KkBnbYRSD/W0S5y86AvR7GmvvjAZKbt3bbbXB2RdJKJh0wbdtKVs
m2S+ZLpd99g4Q8kYlYtgDDSCJf+tixWHH1jcU/2wKNyNU//iOrGS5Y2SvK6u31RH
HY/fZI0d5eC5QE5suFJeqJiMycMzLVntshwCNdyJL285wHMpudrKFhf0QuXlA11T
tkyodwMQgGqmDKFuImlSrdW6+Cj/pxvybvIshOW3YwTU4rYVJATQtxmIqJd4ljfs
++JKIpH5j7GXVO5whlBDo33EL5UMFoz/QhmTMUwxzkODy0n+FXonwUVhUSiG71pU
oi3KyxEbvTFxcHDEa6gP0IruphkLjwk9TcxfK/TeWIcXMe0RsYnIs76vAgOZw8Ai
6jqD5WfpEe18i3ufZ3q7JxT+bO2TemG05uDf0xo6SPIsehmVSxxKJL+yV6secW1k
bPrKuEdMFlrd6DO60HAoxf2D30yDWDZQc4+h2InCQtaUx5lmPEZH/Iaj9oHJ1OLj
s2/xbWcoMYJ9HiXPvwQf0E3ft9NwNc18aMjfRHmbtT8J5TR2oSJpBGOPdAEnAbwt
3koNIIAvuu6yDHQJEB/cpUQuE9YT7+ORQ142h1x5qutZzXyIJSfbK1kjhOHtUM22
lKGpE5uKKuuZFFT5LeKFJ7Ric46m16Fca2Af230Ahq4=
`protect END_PROTECTED
