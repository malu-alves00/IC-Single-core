`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jLZf5Y2OsEd1sd3LrXjx8t1QFxX2d5DNf/Bp7uOP8w4KlZBJLLA1Bz8+ZVy5uft5
i1KiY32ki6tQDTCKXFxPwOIPeMn8ddZbOGvuWFqINBUGLVH/GgsxIA195rZmAvWr
GDZZIch19WlVe2um4IBAJgckdXh8moYw0pu/HB11vQvyk2S7XMBEnLISabdgMiMb
eUt6EVGfyTUxmtZZtzUWJN06ALW+/H1OzmCMnM0/Tkh7NNXjWanFU5+KWuuI6iIC
Drc7PepaZ6+C7yBXQXAOa0VVfMMyYXkrhWfOhLtG2CvLRkgqpqcqOqqax7/vIaK3
KzO9OTt7K0dP9Gh0eYdb6JVWSs3zj96Os09t6tN42C+R9tsaTSihpQgUCgOiWroD
HpmEt1FMZBnaH0Eq/lgnT+tNpRK3D5ZN1cLf9iq5x+2N+Zkz4j35OLwHDYWcJRXl
j8vfRl4zm+2h3yj3IfvpbbwEmXiszIXU4WMN62DXIQON+O4dCIaueI6ZDs9eKvGu
xIeIQHT34XJ0V+k+XgVDOeANt3x3m/uKwiBNfE/MnUd5t/SVbnyAgEP1+gwmhwTC
YtSMHgvYyGX58VNnUz/gSAVJEBTGAlUzq0BeHOuSP7Qy7wNMYSz11ulHmQtQaMFq
IwojU6C8qN+1gYGIHDHtziohcd1QpEvZRZ/yS6cm++Aajwlb8DUzFh9xNerFe/wU
tnD0hWT9238KJzyNKrG7TLXqSf+RXVJaN+6VVNjenMPkBunspR8LzJ902rZWBUoV
lKJ5Tgd9zsSf0M3IgHzCyfRVnQ6y9Fvhl+AsSw5QoH1H/w/1XGUOqC3hncayvrUj
zngk5ew6HuA7EyyyZFxPVEfYeCV4EWCp3lAntAlRvXqLA8MWx2PbRwz8zExIsU1K
64WjKV3Q3lVKiAKAQS7ILvEPDsLPQ66KP2k4ciJplwXes05j071gJcNl9n4HDLmJ
P6impQH1JSTzJlAWAocBT3bjtR6i/9rg+LPlFsIX34Er/Iu8rzRR/azoP6YEx+7z
ADBFteSUQKs6wEnIoeutldrF5JENq5f3DIwcPWUTLBuuyCCdLNQnM0UlMES6Z3HU
po3Uqpa+2Ej6kUxuElRqnTYiDwpmGWouUO/tcDiiDx7dqnonTz3Ab8166/7egwy1
d2JuAwWRSwLBPtq/y+A4C/Brk64RUEeFxXlzqtumh/9hEjOHOOjEOCO5s4ch2TsC
7fu+RBzrmzypMFezvmQAjsAyzE3Lo8V9Z95VFg6T9ljVKU9WefDHF9097os+uCbs
53HuMVertZe3sKsGs0CfdBzACyXjqVqxa75p5aipVblr5X416dMWxoPPPxg1TcqT
e7Imtu7NzjEQ0tvLjXelnQ==
`protect END_PROTECTED
