`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
m9sFWXTLPpq96C9i7BzyPxkCUIbFT7DglWy9OSON2e/Apfbd7oJFdeGuuyJeeeaW
AYGTI+FfiRZTtyLc+p+mwpr+5/YsTvXxLvVc/L6sRV7+GbVotVbr/8j7wWurD0pC
jTGRUKTEUPRPGiUTA9NGTxbOzwK9szKdbsxUguQKXmip/VTHd8L5XhRGll2w6xJf
T748fdBnujSASR5grfPQV8uvKGlutRJ9w/HiJUZg6T3zGkK+3ogo6NO4u5uc4H+r
OXji9n0/UdhCySZzAoUHYNo8s7ZHkXmLapV8NpyHnLjz3F5JvSpucmrFzzSDFGC6
83+EbWBSgSbOfpz1SH3eEpzOw7K/6vrX0upR4kh34g1bx5YQpgsFR5PyaqWGyJs7
CVmsf0sV0R0UZQ3LW2Cisz7MImsCyphQh4e/LQWOTbG653XlNoHTozLJWRqnZuWn
/Ecdoo1d9gyijtR5duEmIgGxt2w2lJTuQW8NidcB3lDYnzqvdfCFI0yLjcSyDHgW
zPYKo5cwg/Wy39x2ZSoGj/w6MF1gB9crTGNJHIC/rnyVZUCWkNawIzxZ3zuAeOmQ
xDsYv21fj9ndxBd50+caBzf2KGV9kj3nXXJ+HawxqZs88uP+TMAUUZIDEg8RBGEV
dj5qA62+LozZjILNIGD7EUr7fIWCEGIzW0CJuNV2BekKa3ZoishAYIaLNSw/B+CK
ur7ELo7knnCItqu6tRSM6ok8ugCAnNXVOmXKRx089JRllOOYWch+gZPzDTn1FG5g
zqZVT8KlYBVgM2RTza66W8Y05MNYnZCW3N8zQD+/sRCOAcJXNP1mgeoBdy4MnWWa
lOiocs7SQ+ul2TR4w2YVzboDBjuHKT8wcLkYkXFL6Vgir0ar4zCLbbbe8+dPAV8D
bcpBO/A7RQpJ6YopUagaDUas5V2fK5i+ZHFvKew6FLsvpY3aBh01Q17ktV281nZ3
0teow591ufPx46VgPHypzJjuBVTIm5d5xPsGq/BFLV2y+1sa8aeMVIZNt5lPA61W
dr41k2IfUCJ25kvFGn5loaco8CRc17at9yfN7I0SsaVaVo2KyLXWYbo6mpieT0as
I1jv3a1TjdbayhGGuH8ywuZd7jxZtl+0f3vq9W0BtlBwoiqZjiLIIz0mphUFz3w/
+t01h7QQZr84OcgNU9dWF0FizXjszGaK1TwgROojS8hBZfrrieu6vl7pJNUr/nL8
Fipm3uxRI81ssVFroMsftnT+vvhSoMItHgsZaa0zPLXyE5gaNfXNqSKoQ33/hlcJ
J1t8jnWrD7wFXEhT9NXKilAUtdibwUlaJkQKNahzz05Wa9Av056TJ/DrUtMzfdWf
JlNkeooEXsebJ+DMPK3L339UiOVfy0moF4nhP0x1/YsWozhZoFNlEAsB6xaPxp+C
xGYKj2/b4a6GsLSk8FL5sy6H0hYqRnkBnnQOa6ZzCkxgimJ7FDhwNpDyrLq4PrcF
WFeZdrVJ6LAP52udqzI1LP2XVex7x8XCFsDOaWAO34M6KnJ6DxBP9nQaV3MdrnEp
OsYAfhGFRSgwXDnZntqkh6X824r7x7EEujiKaAeBmMkKPA/RiS3XnxfASxpMN0+n
91POyb7WVhpfCCiTHuRaMNN1o85OsQ+EIM1kkrQgOUmmFDIUjAhFYSy/yLBmd1nL
05cy4jzUgkR2VQVBTR1XdCQykW2+6yGvWodV3pHsFdhCyanGpZKMvOsp7A46quEI
7HIz8LNe3+Loi6zQRkcDnuX9PPZEbikzqvrsVZ0uYSXvTBrnOVlIHjnwlQlT1v8n
guPzQvpktBIWsvZ4QXcrDLj63eUILrSGaBuI/SXqAFRilBvlyqmi6f4AoS56BTM8
W+3daTxGy4/fRmqMRIdN4/azqNc950/5dwb1CtSE8VoQEZD1udKpAORncYsz1PF5
ymrpbxjU62VGGgt4l2xbwg/fx5B69x8eT8U2P/3P/uVQFL/9Iel8FoqJynncJssA
+XeQQ57iBpQA0aOctvKi9JDyK8vX9DRpmlYZV38N6+19CeRt9s4cTQ4sygWMADQg
tP852gtvQ9HxEBcIHrrvmmto5b/2kc6uxTUahIzqZQD7irZ91WJhYxPzF/izdMKX
a3awapOQGc947ws+B1jodmOe4IQyCHL411bSgPWSz+blc7biR6f+i6j6sSICjjdB
2A54a+iWIrdQL6ZwKyL0ZahAjQSs+/Re7bzJRHr40xNGGnReYYI7K4Twj9IRJZeg
Qv98aD1MwbTjjEVYovJ/XoX/ji2CFUUW/Sx0GlQKGtrRzFB5O0W/nsyASI44uM0U
sY/sP3FYLHd54WNRgGEKLtWq+/Xbo4ZPXDZgeEa3ESYpAvvjAn922nduVx7rqtbP
vEjxuiYvzPn3wPQmoKGJRTFcfiXm6IXwiWu+uwgTiO8kn+jpx5jlPDi/SeRsw+J3
MemiBdImS9/XAS4RC9QJ17xye9bIanUu3ngBCfSSghuLlFsBLg9eWsHnbgCTlmNF
aNDvRfrbYs3SwRiJM3hsTkHGpnY4j/MginorhlYnmFSjqPnNjyGsXSfcqLELLtlP
WLXlW65JjXDDByvT0q3cBg==
`protect END_PROTECTED
