`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HmQ3otYo7YvLlFuvvobGo2F/OVQpF7T8baZVbxF9Cmk0pGMazky5cr5kev/ZD3Ud
y3wzttitMcnFcnmkjoXndLJH5LuZc8CAcn/wPZBqMXp8wjfXMyXJ6cWvyB6WVSVk
rJEl/lasARr9iKAv9gDUJ7cRhZZHgkUWOLTuQlpPF4ZzxXa05/oqsdUEJqur00nP
MzhhLpPVQUJebssiD/mj48nf18b0bK4650CTkWdtsQxNZX3lwmLB9deCgz2FdQ2M
xySsFrNk56T7NhIzXZIHq5DxZrCiYn3ATvtHHf1V7doawFpHvPZtZAjhHuuK3Hyy
I8zQilX2qrCRY/n8yHr/BPfQt90HovB+U0DjZ4csj25MZKQzGzxg+IweJBYz3xeF
idZRKd552KY8H3nWoKiNQ/ErYf2WQ+URe2x4ypm4QbNph+dt2O1kWDCnLBasX0dH
GeurJpgKKuVPBwwwR15XL1HldBiGVvLpK+YMNZGgorTPuvlajECY3exqQ5mus0Ra
BS03IHxCdHNvzTI3RkOM6E8NudJvdxFqUF3Bxoaok0ZyQxBQMcSgKPaoLcwRIUZh
MTQpn/4YdLx+Q3T2qZQF4+E4JFXcL8EhyJBvF7p5ffJIqkEATpvBn9c/mMjh5dmT
L4oaAUS5QnVH9mNrHzKGncXeXHh8N5WDIlPeLXvkKl4BFxzKfkfVWJw75VpmRLY3
9sR05lihFkOHYwb1GLFUI/VQ9B/hbg8Uoh5ayFR9Va0JS5XisAzlzq3J4L+TvIeK
xmNbTJ4fGYB5y/7G6SMNZFtITSumCIcbNYxxLZnaLZmuDbbscVS9hGKbPMCvM6Oc
u+Yl2lxOBp96qcr15kCHwKXMKbzMIDCeTo7id5JhPH8T4hNLG0GTOsM1E2ykrR3S
qVbgTUZDA0VLpCr+ORfQzL+gK/TC2ijEmJ8R1vidxDBxO0PRDQbvhMMmteJC+I21
WOUBWVPksTRl63MSEV3MbWVHbIBY0mEzOJYfOI2AApg=
`protect END_PROTECTED
