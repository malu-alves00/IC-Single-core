`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pOIeyu91xpHlIp/ok6JvbABpgiBKF9V3WrQ2d74IN7DKCVyQJDUZLloXCezLeOLU
UZnjuYH0qw1zt05K9vAxMLvW66EfJHejF/jSyF7FbYIcNk8DhzP2wlF199bU27yf
oYTmtttE546Kdm11FNNzYecgHyssspzqDU+FUXaYMLiXdbhRlwCzyC2WFbUAIGBl
Jufb13qyBlMAH9Q/9IoBcAr2qy41qTiociEx9F7gh2TBs5+3Z4E2a5l4V2UNZf9j
fywKrafkeJRHoHS6OHX/oIdg7+nb4nz3we8r19vcydlTMt39WXbRHGslkaZkOm+I
Hfu/+ChgjMoMXE+EKS10lkTL80T46EKnCd6BlC2WA183iu1/42PboDTFy/k+BWQ7
Hcrh+2nU5pGgQY5misGiy6FnXx3N2hup57OxBOAsI7+hDe4FuFD+bQmRAvilGsKr
DOmrr2Kb0xLu70hku1EB23gOM7A4rmLRkO19WyCpc75yElYOHKPsjDt8dp4yci1j
iX3pnqAMnS3B5T1jS9589hG9Xeztpt8plFMCqyz7T/gUv7gIudUfE4EsecXNf+AV
ftGg73pt8t2NOPhGE4FoD8kOquLpMzfyisQC76evsfY+nYxBNoqD/biRcO01w1SG
ia2uzQjWnkymYhWecmVvVG06dIH5D+DgaULQ8QnX+rFCgubjSwQwp9RJHRBScjBf
6IGMUb+nW2oa/FcqgW4WgIHfMiimPIUSu9vThHhX2Kc3vl696UuCDLNmWJ0YWhVJ
MLoMV25oqC326B5CXLWlKAys9qDSDgIpcnqO+9m4qhXC0Vf1sHFsxcJ3C0dXrYSa
i6fqdPqoumKGbCBpJTP8ln9FG3pGOCdyt9P27nagUUtms4tcOtiqn5Yv/UV8Dpb5
9hMMRkXuE3KXuILgVaQYoQdOZhh6ltTPqvqoDvS6hVGk0Z2/C75M1ymt2lnVt5Ol
9VC0498yxnxGSLWZgSJojfe/yOR8D2kViSewIW/CQvlGMf16DsdBgWA5Y4l9twWt
0/ZjX9YOq8REFErBdi1RYUBFq0wjMtye2Dx93L6XyDvcOAVuaHRe2yukefRVXhM0
AKljjQn8cL9n6FR5td3mmGYpz117itN937VFNNc7wgNcAu9aja00wsEiPTgzs2yj
I4EFQnVOvA9YWvrAxTCRXEoiJLzif8AW/0FLoiRZffBbqBqf4zd7QgxVTOgzCqut
go449dS3TwRg/dYUWT531y4S7oJYi584vR969jVSaA/BP58Pi9aKqsJOgvGxWol5
Qe3m/QM+K4wSe8/WbQ8cMYt2pJKqIF9Bm1xjh1VnPb2z0HtpDOaz/dWdI2v7a5Ij
e/y80gVmyJRNr7MJECnl3wYevgI4UFyprzcYvhijmGN90KzXbcOi8eI6AWQsaG0q
aFx1nfht/ONbeF0j7qbObV89ovq7YjiCOSEH8lpZIJVfwf0+BXcUmtG1Lk12oC+g
TiZUp3ApnsEmtJWvE0DJ7f1/dZLVGHmIAzkSXvOC3J3YoyN/6Bkmmcd06PVxU076
8zkpz3CTACDn5O5LcN9g1TG19S35S6fZ75kU2x4obk2LywO3nTDxA/5MQXVgHpfl
SW/hfPQ2iVSjoKQOywo54JGgdNA4SRu1cGlq1FalDm2FGLTh+CmyeyY4ogfoUMX3
XkpJlPNItuGZM2KQDYzK9dG8xpOxa3180sIkJe+EjDnK99xUZ1UHopRF1Pxm3qyZ
a1BKB6v5q3PHyNhsKRSX9A8gvFuUqnas311b1lfT+G43bNbg0IAi+pxGODjse8wZ
6Tqg5cTI+sn9tc4TladHcNR3zEdqVOIdzQlOwSTiJcNK8mpLj/IlsxoE2FTMGyxU
R0es+PTwD7gbZWVBZ41KLrN6fazZWTxY0lPPTEdml/sUyNXSanKaRrFPVKI+AF0Q
oe4Z9ztdI6PpqwgLdctn5TS6YXzq53QbgnX1lL0m3ztTMGeley6n9V6zQyHVgznh
SRlgkyFovh+H8UNkS4Wmr/8PLa4noKMKmF344UFIDaenGe1lSo4AAAFBlspXkVqj
WVsvXBjhDR4MBrIU83BbMOQkqJfBiQyehU8P07eMYeWAdIP4TLHIOBGD1dDDSkM/
L392asthVJycMEiYopJQVE+rqIP50Z0twhsRKrqFNKPlBI+jkibjB8xDGvutRzzK
NsxXM73fpnu6cJMTKbj7PK8DpaGbtSJgrFOs7Z9Zatmzk8/isyuvcZ+ibAGTmEBO
uPy8x8hK60gAXiNjz9qcUXbF4JvUx78Ptnpp9kn7L4EukBMgw9NMpwc4Ma/TcUTk
+r+SfZyKXYaMGF709h7PDGf9i0d9/qabHoTFXhbxqHHX0rNkAbZ9juKWKtfEAAep
Q6cA8gFg0UMNv5DpzPwJ0Oc5+6SagMchGqSHVOPY4/cFa5GEFTfcivratNs4GZRJ
qEShRMEGsCobBYo77yXlTT7D+hakqA0Vo+U0tDbZrcelIbnj6GAhlVDN8NsuqkpG
BxqiZKt3rbIx3/SLRZ0DJOcpLwAkXDqZxddUovPiQiU=
`protect END_PROTECTED
