`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
u94ozrVgvE2f35bUefRbZT+k+lqaJ/SSjuYn8ZVzrvBW3bfatCBfvvLdxDAp7lrH
e0+TeHlTFAnaRomcYkrpT/ceFXcgakmYh/DNOJGKlqQO8YHLOiGxTf6nOYdAXzv8
7kFwIWXQN0mVgZ+PbYuvI6tRnMyAlrCOHL6ZyoTWjEiBtlW5jEUJL5u6sD+y62vr
ObREVMKR+zTSj/ba5nUETc8r+r5Lp3dpKOrFaMD0MU6NdNfWpFpltm/imyAUBO4+
6i2swHchyB78upzMO1kVHRdtluIpuNHf0TjN44lS29FgRoegwu6MMy/pTQ+530Yr
H00EU70WkQn624dAJCQ+o3MR4zMGlbXCCr3ftvi8I85uVH6nUIOp6w5PbQUEbBbD
ErY7/xo6xnUE/eH6siTyk9WzUINKuIGZs3x37V9qwofU+b6OJNgExKPrNmsvJ29R
u5M0oQYuZ6cq4KOV1jmg62Ex3NjF0RhBT5wVAX05GOnwVxR/coWCIqzdr98quJFY
oyqdrthOK8xwov34jxbu+fGu2iyxUfr3Hiuct+/5BOAMWqPewzOBw/lh0YT6fjIL
p4WdvOkEPKnxR0xZms0bIEgY6JJbku5J9JFDqw6YDVCJ5S7vz861VjCBah4TmS5v
9IZo4RuRvij/ZB91RD/wbz+GiVhQ2/Q0K/xQjkqEpCO42iEgx8wV5gS/NtE+zy68
/7Ds/HkzxYFSNbCMUQTozDaRfN1dpTYwIgwSwhSRQaKOQXwL+BIgdpJP2MFsuBJM
tD8qvGYi6YTHNeduFfDqKm4+hq5ay7tMw+c0Qrpvy+beBH2vAzP1ZuADDMnIt+db
j/jIewm6OQgME/0vOAOtxV+RSxtXri9Wk7fZ7kFPrTNmnAj78miWQnX/MfgdhGsk
gyfcAIaN8M5xH1qS3tZKRXZKkzDDrNEp5u4K7r6fhnHYGaT/8tMWhgygsk0U+wQZ
UPjrLxCdwdc4sstGOe43+M8aEWnOJQ55vKKLBfSnaKPZNnEnsGbvMpbP1dobCwyA
fkePNL5M7g8COoFyWEE3hDMye9Go6Rl7/jKAnFA3O3ozBpCmmWUIXk8o/Dbtqm8g
4zejT3i2Cq0V5okZCVVhjj5KuTwM23x1buKxZEqatw+n0h02oB5uvboZcQ1Fxa96
HEIFOcH31/62Z4PUxxqPDHsX0f+5xoLJ2nG9eGBZAao=
`protect END_PROTECTED
