`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uHuo18y+mQAzxhcwFWgu33h+sTQrDSpsP4/budwp5lFPOWa/kt2BmpL3g6GbVpDk
A/DCD8wcLZ1MhBscN6gyRrjcl4AV2s3e5QNdd7IVNiaBH63IkKs0AaLt6rFn0kOA
1LyugHOJmGcdxpDVnogGKWQGA1yKC0jQ3oNP9VxMaIvhduJEswCKJFSHDLZUZ7XJ
4isj9F4A5HC9h41ZA+Ydac4WW9FDFap1KjKa89UNg2TfAZimNGOWhU82ETNMf3r5
OgyrDRI59aThry7cMTpLjLf+TdxFqnwbVYhemP2jNHXGoj7aVSft3Jt8fk0YZ30L
KYKrRxEZMp+aJoYeAoFhVvHAJaiHAC5YqcsTcDCJBtMG9VCY6K55Nz0R34/xTzGW
5ufoFzBMh7ejs88AZnu7g8PHp8xbSRuHYnbtH63QZy+7vcaymSs8R7CfEsj9zxYy
Ls1/x8oCFFK7QLYrdqql10RvzvkYiZ1a4dmFya5GDKwwOy9SqgGC+/218HbzfV0q
mSNUzv6DyXAb3JwpPodIuou9u6kGeNmDWPNXmQYxzoxCWzJ4d1QosSytrQgMuI/w
98C0QoyiIwxnByuGHsUzVk2+2pevz5mlceUslw+ySc7CBUKFEbSy9EUWXU7v64hg
0Y38STWserCmZH+dLgEas2YujpRVT5FQR+kPH27a49AsOoD0k4pxO/R5YDtnj2eU
w/OjdNr6tYQKTSW4MJrxNrR1TlUJl2IfG7kfewgwW1j5ylsGr/isjeCuf1hEdbjY
i2/0JI+oVvQgDR3omaxGSQpY099l+yQ5Be1X0UeIUpJ0tcr6sHOGOyEQ0h8860IZ
h7tprVraEUCF3d2gUUVPwSF1fov/0a6gvVeMrPBxScRYCs6l0sGaFtSK917VCMG1
UamuXwXedQyoNbwVWAHUobnvRIi29Dd/w59SvLip97sOk7k+ld+4NaDjm/MB13sI
RjAY/9dxgVkja4CmAxSxuU/NxcbAvX/npgTHsajVbdIyXxbzQFTXTdxjqmnbbVvq
KpjjK3hoYZqjZ3p5yy2S6Ef/0qipE2fUBz2YjrXoIXeKpa7cEFzAsuziymmb7p0M
4WRtud9pkOVMKYY5/N4Yy0g304FkKdIxvPTMO6+U4Y57Oi+uhNmX6k3Z+iu9cjbJ
zVTRP2NluCvJJsRfbr10NTLwUZOixPB8dpT5oKDqgCm6yt4eUGLMvicNWjpp8vUI
LeGf0UzKOy9BXpSXroCshTaUgn6qdASzAxnje2z49ZroqmNrhR5QTcdyL94tt+3U
DvApUPda7o4VTRhw2/0Y/U68zlsG8X42LPT4TXzHW83NOCXke3ZnxoREt1dkaALf
7DhqDfG8tpwoUW9Amar30EQBqQwEE6X7QiLcZB5XPIUhrNgUoDlBu/sCGkNk56Gc
5H3gwrPFN2RC6f9bXZbgRmDakozoHlF8FXMH4phcOMMCeQ5n+ZRi5kxhqQEVHMS9
wqdoen5e8m8I6cTlGm4AB2a3D5R3ZGzM4uyEzeCkIZjAc6KXuNFA5JS4Sgrrfb6v
Wrzk+OtQq3GLGhIvZhd/SNw5e0+1AF5KCumNWuS2ZmpauNSUoNyb+SmLxp9RY3rz
WdzoqUuBL2C+mpNOOEGjBZ/abMSwoUOpCQQehOCh/5Ub6Py6c3P6uUqHGW+hq3xT
ztL0wVetXhp/0Cs3OpRJK6bqPH5VyZopGra8XI03M4occGYheTxfOg6O89egGrpV
FnhKOmpS/CFNHFF1P2GCYawIOdOcOeh4Eevu8XFMIT6NTuXb9brCM15vMD5l9/cB
T5UfJMcHAdrOqlHbEdHFduykmSKKEDm3nCTnAhO40CP67dAuHI0b0GDxXcP5owo3
aBL6FOZmCqBt3pHP0KznpKm8PwpAhxa33GWcE8BKWLhKVC+7QzzlcVGjr+nI7xxq
I02REzOna9GT4Iky32Uvu1um5CFNMEamEJ1UGBorcVdLFl9sFWrZTo7fgJQDnRDG
I2tLAAng22dlTQ7OjRacwoaB6KGFIpL/Cx+6nu6Hfy0i2JK03DKdaXi4YNLIbREe
DTNSjNhLLFFeF1h+Jrcp2u1oqW88ooYOCOIHrthRctNaWa1GrUACSVmuvAW7IIbR
9cq5QHKpxHBlpIkif/pYQJAT+6Tnm3WPTXIpo/MPt1p/zH5ECc6o/eT50ROMiyoU
6GLwO6VdavwYID+v+L7Sdm8sWLoCbniyRzLWjtiNQlh5BM6MN7VxVUFbSDQNTkVD
S57x7jptTuoMznXt9g7thEWW+zbYbyavds/w8R8XhhkdPcHSKPgXjfrHGHZnjSQe
t2QZ03gHRPcQ5T4lSyPoOW1oF2Bxg8eITaRWtR/SdgxUHNZiN++u2RaSsUK9kKLy
PngUDj/0cMSvpZ1hz2ppDK7/ClVYot6xirEkykBCVnQ5u8oSTFSamaQbXG0wgfeg
KBdbla4sPQs06qAnZaIquv8V5/Kt8WSg7bVtXIjDJdq4ijoup2pBw2psvyN6Fa5r
TyT/9UeA/VhJcdyY8izm462QTXro2n0RHPCmorJj5Q9wftKFhvpRNJmC4xUR+fFx
2YrZmYSpWAe+xchCfS5Ddg==
`protect END_PROTECTED
