`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aNPCsl0w7RJcqAIot7k4mjz5LfX9hMBcgWJvmse4/Ku+YM9PWJEKNqDeUUkjy1z9
Gricy1Xnqg+MBfrykPS9BNP0QkC5UYP3pzNi2UHHYbTCHbOL4q6Ww/fINKplbZC6
mA4PJGAQdhB+PmVJV5DK8YTRPhLH397MxbH6ggfxIv/iij4rqCdfDxcD1X6BZSJc
NScS+JoPiokBfHxbcCWtutyMk+knV2hG98hzXJbALGMjhDL8gHX3sqqRTBLOyBVq
G6MZEAFI7PAfSOoDpJ8OZ3m92wJ4FOYc5XQfpf6DMJx6uco6TM3HPPfwAFC1rqmw
OYoiPSW1ZITqfL+Svn+L0vObAo9aI/Y+NxeTq9jpuhtID0/2ufMmHvKI7rpe11rg
8khpkVfvdMXm7/YxhzfDKoI86FTKVa/K0WKuBfQVETrH8lk2aAnv/WD76ovePrQP
5CMit8PRNM7JeyxupRzoDT9+MgZlWVUgSipFnT7MBxii+1btLIRTEtbDDMznyl+q
eSR5yEqLqbXhc/7gjZWDdMugtpbN9RzSVWdtn6+DAlNlRTuZ94DEVzA/kJuzYMQ5
DKKifbA+QjWqXYyhfEkAWCWKcFmGfYVD0vf+JNlA62sanR8U7A66hCmCqUiAsVvL
TSK4sRqgEE9dcTSxKGUjmYp+bcTHq6DwFgQxjNttHwVMHfpGxPvle1Qbsg83ksXY
HGEzRbdVYJO5W526qNsrTdwJEooio1iMR1oSy2j3CIRlsmRFB87lDxTqAdjXaJLd
7JZDRyI26Ma/JQ6+vtMR3smbTpZ/tXuX2+FgFeiVjhdhW0JUl32OcA/ncyNA6OZj
/5n18HqnZkPyUhcYP7l9UA7l8vuVcRjX+TH6btV51feQjgft4RkDQAVCZEItE8q1
4kAAvZYKRqunvLqE/wa/tQo4NFatgAYZPaGuBxtt03zwWEk5ic8P+apqlznRUGNX
+VxvvpzNtAi0VGi19PQx4wHxnH3TjA0xteLg0Kh3FOyCEknzU65H4o4wU/85Beoj
nB14hZloZ4wT+2yti90LnsAkSGz85fmgb03zCS1UkiJgI8UJdeis0S8EAzEIpwSS
hsP9MEzPn8GY9+XYZBoSg68Dn6b/MBeQrwwqeL8b19n9zsM1QThaWnoObLGsdt0y
n6yViU7mZsRnXSiu0T4ZItC0SLA7pwqCmbctI/cz5p9MqDVq01qfqTlO4cgBW8K8
Rk8v2npbPkqoz3sgCn0rsApWVvm4aY9WnWk6wWFp7NV0BIRnjqJGRlpLcOth6Bs5
Kv++ktZz+A8cUlOyEJlmpUp9refMO/5jEqG2GrUZE1XaCdrmso2KY37pEWeZc/A7
fTVsys0D8ZwoB3BqsN9328VLH2UY6jK6K6plDb3qzdFnN+ewpO6zWVbDqa2oewev
nodkIELBUUQJyC3iFUGKK5m8k360AfkuU5IyyORNc7hO+nC0bWzGZxc6ewEL9wrv
3wADBXCjpmNDLr/MWZzpM0VpZxNsijRi2KWVG8vjTPzMl69LjvWAdWBW39U41LYG
ItyMY6jyKehH3V6Qhs2W79Yzy4SSq95Y0191vd96NNcZjtNCyprPqHwx3uAoC+LH
pCEZgLvdSoOfT0qbhBOTGmuGz22LhAZEERNUS/ryNBpnLHHi8GVUtt5o0zZHcgwO
ufOQdHXgsLDa9wrdglZ+DyLK6phTI1drgFz7Nq/xa9SuK1fuiIB/rNn3J+D9HDey
By64xkAo/r2ygI//OUOW1PPfPPle1d87nNY9IjP/JylGrQpEnNOlkujOkvRdHxf6
ZUeAnWLxyAPJ+GVHWgkIEQ6O+v5NTpud4lEMHvuqzs9Tlyz7lSrqOin0IHNtV26N
BgLXSBCQOes+Ej2sQCOlp3G/W+Rt+O+HZLtamwsFiZLJ50ZLdGhBnEUpwL4aWkER
dSfMhswJtEWTjhFXLZbattLbqef0QZODBZCNE4xaxIyfwvFy6fxVHNUJRmspqqM2
UP4VmGAHsn89MQkeC9qlqNxweFmcBJSjMDVra2/W3+POpXlBR4ZyDv1f4Ltexfys
6436Pw4YyWc/i4eNFP6EzmU7qM4CEmg2TMj6laLpkS6o09BI7bMfRvLhqdidihyX
1u5AAw3/LLXeaMatxZDhSsb1hYce16L6ciXP6NNB52UGRKsum6wo0IPGiPWWvZUT
PCFKCTa2ha1Ja07/VPj21UM1YQC1I74n/BB5Skje+nq6SFqxGqXls1Tyv9h0JCe2
+J4kvsf9d00ajzPD9XMWRv3r+uGGRx7GddJw2UZQQSqATWXUzN7fQ6H22Xg751sk
g4HXGSXzmFyuGana/+VbA2YtsnUbh4hdd32fsJgfIrwnBCx1hqQS2wD3pcWHeMz+
588pCUomWVXocAytgZ9bypusjTFMVIkJ8UrBGm9eGdHU7Vd3c0tduVBWe8rrb8D8
CqvaLefzlmT/3HkAAIyd9Opi/NRZgdgBpPIm9khnG+A8TCFxy0MVgsHiLuviey2V
gCNHnSzOeRbs2gWAEcHs/GHNOhxQAGDzo/hP83e9Dtz312FyiTiYPFfGjvDBPgmT
7S6U+M8uRaxmOvyY33EkaiEfyEehb0YeBbOvztn6lX1zrY97PYWXptWTdeTEs0dd
3Nuzof0L4Rf+IeZatYt31RHRsly2EoguI/7kQDk2txUWH4S5j0OUhtWXZKK5LNR6
VqkD6C0WLg4kqqHfhHqJO1+VKqvjdhWqrdvZi7zoCzl/byd0cVBDUxG9VDZhQgAx
SIEJIWRUZaZD7r1YaC9vU/u/fLJ7tr27kckXZy1xPmdT7XfMjKXj71Cka8bJlDqD
cotHLspjZdNEZuD5jZSXnCCzJR7jwqsjZmpNPGmTfBtiO0Rrk7XcluDqLK90FiQR
Rhbi++fLSaCBBkgG+E161tZXzrLYqTACwHJd8d4/uGcGk4hniaYaV6+mtsFkD+g4
WldlLtpnO/rcim14ZaDXbO3Zmi9oUEO+9jU/Ds96ambFIpLIU+WW2RNDonr/0K+P
8Sj0mXJFLNlhe8P86iRPl46ZWqznAaz1TUso3/BfpRJVjUsF/GObaVkMfHEPs/a4
gER+bPaLCdmmXdPyMAxOzroxsOICDCaThHflQs0XCIuJQxlKd82sjNOJCTdazbZv
hDCI4qzxVA3vC54msEwdoy7i1vuLH7kMis3OPPX+Ua9fRdV558+QBYgtGmPKRrcv
uTMoZOc9SBoRP5aIzYeAIVT3upjcsq83UHoOlDklRpSPXYx7CMn45+ljO1dLdgj7
5gTxwBGjdT0/rJi9k1UZVzIqcHinIt0lNv1zPDx1Z0r5gqnxw6rS7nw5fELWg/5T
u35hVGQgVaWPWWbfIqQHGxZ+UnRAb/lG3e7go4+0xip6vZ5PSNdLuPQQw9inoPQ+
PdqfXbNhZmIJTtzC5VpcDvIiqGbdgCoXeVZj8vcDqT0ddPyQJ0+6jXOJFBjmW24I
5lxEECU97e9VqMGq5nINbv9uerFur8LcDW4/PQVv+mUJ7p9tG5xyM+tO/a7ItbGd
xVgId4qPwaFGEauR26vRp84zTi7iE9R+roU8r7ShACa64qaTj46w2d2+5iHLjh52
N3+rQWi1shc7SGT+RxxkWR87oyfpv3tIxqn/ECtnx4882kqRfVOk+9ZtKiHQnNDc
UpZz9J47GncsYr5iPXyftrqlnbtz0swn16K3x3ulPAPhiNpTxGjCOxNPRETPNB1+
/R03o8nXrUhyUQaHpOfWDNSD4QSW/8IXGLanhFG+nRtXs4ODy1j9x8wTC2c0Z1qO
LRd/WPG4IQPAMHfcK7DyHE1JSQumzJQAFKbg6i75s3e3e3slOOuI1sC78I3ZjV6S
ciSYtLzSRLVMDEtkRYEzqSp1VgKUyU9gZXyCOTIWvLDV+7lfsYryL/uOGSpFIxyT
/EYpl+QvLQnBHoELuAJInzF33ZehNqeE+7A27sp6bgrWecFhXiaH3EgsWrpTx4iE
mvQLfEXMU5LbQfGs/RL0mFNGHtzelyaPw0RoiKyvqbPsKw1OB9FmX36aHYTPbAGu
Lob6UpJovYJ74JmyAvzpEebwIRE5InrdSvzcODJ4mXgEkONvuSSmhkDfpoFKRg2J
Qku5Hm69LWe69sebfKO7rBcvfytdf56C62b43ZRhQiM4Tkxmpk65SdeQ/xnCM3lM
tHqkUaQILRKYNXEZ8VVJoJDJhsBam5iW3NDDp0j7/TwsmSsZFGkLWkU7YNSktai8
nSTaBshj3qP4HnIXnPNcclKejT0OWEdWWLIktHgceBhml40B9hLr82VPicihsrfT
n0L80eD5mvzvuJSMOwpu03+qOPS+fMqtPOFg60Y5G7svQ76GD/uElZmshuAtc9IT
/tfKB8zLas718S2+984nZ5Qx7gH6I5zHnBSFX1fUpd0iX+mAruB41NS7gK2V/zny
TRvVRcz4wNubn/5kfOFsOPYzUdxEQm7NXmx9aqHzWV+nxbg2ifYthjzScYVoNRsK
75+vdfktpzwH7LAQetZLdtfNHPIXwmc9Tw5JKn3gPbA3NaGJU0M8LYjnabtzQy85
n3HqdkXWpuSq/Kn3CQmiHF2/2XmWqMO2h/sRyS5sq5LDRyF+gFcI59LtVLBgjqNi
exYTQHJOWuXeueJs3jxj3lk91nU8jJer+an9Mx8aTgw0lFv1edTKQ5pk2QJKjhpQ
xq0Zp1abBoTP6KqiAkpuvY5Ip9lrNXWNz535S0dcdtQPlFgM6dSHFbHth+2ROOIR
UzAm8Fea0L07upbTLfBqwPxwka3zxKULOq2/415hMh9r56J/LEcHcRlLUK7J4YjW
JiXRqEWi/eP/MWHQvEFIXuM76WSZQq2VSUaRMDPlF2bg7odrTN36RZsXpGS5sNrN
cS9jWVSiHRNZwFKI2ml9QSW22LwW9YJYF0LUiKMRxMCQ4ygboHqqZcdeB6iQgylH
fPVANQch3FMAL2Fm1tJlyTXsAM0Det1eCZl3QJC8+fP6rVuDCc+/bE/uzjmGSnve
93xZDp0zoH0O9xTZJAzPsFpZILxi2igJcNTwm0zPqporcpvJ02PAzNNVswQ7TwVU
GtCxBlQoS3mRLr7S92vQ3CUZHw13hN8mlNAkuHIrGP4tHC4QP1lJEEujcw+1VI/g
3VNrxPGCni8W7FPoJ555b0qmewpt9+COHouMFOhGP8HUqesnn+NtkPl96RZVLrP4
iotraTr4u69Xru1etDwv0Zxf+4pegiD08W7DIh1gk/mom3eVfDF6EkXYXt6YY+Yb
I2gdz6vAiM69/6VeMAt896dwzbNvHeb0NC81JWGv5RRN5qU8TgKXNGe2vELgV+im
9Fq8Xp6oe8NPWoYoqSyRJOvxBERzhxCn7Ixpm/71/5uH7pgEXhuJLHilYOwOkdvi
YjsMDhM3zYesWHldsZrMJPvCM2WbIftretql7I2kH0oAkfeQytd0qMQ1KhOKS9ri
Ft3blCJSLqqHZB+Tdf44XgTmjihzi3PVS7UysS/g14OgXmM+U22UKH86CMrfwxyE
nXy7wOOloKcStP7a9zocz45zoCxt6yM1djkn/92Ak1ntYU+E6K0ooWhlJm42qfbx
pPKRpC4zKZOvUOsOGsDc2K6jOOJHsfbGev15r+iTdDzoMVvKqXSqaHL6EMTN0127
emhjZRAgnuIUx4xoxgfh5vgOk5R5A/Ds58D5qPn7UB0tK4WvfBIEhSfH1kf4sGzw
6EmdMmXqyiGjbZ3wR53STtO0R8o9l9PnHHVPypzFj207ligszuP/HIgyV89Hqzkt
C5LUdb8OhwODA0g67O+HkhbB3EA6rgRppg42XG7iyBhjk3F0ozJ3hctwtck2R9NJ
F71DuYh1KIEu8Yy5I2uJGQWP1ta3G3B0zOQo7QThr1Qd3QWPDm0N9ZiVvSzLrAp1
8NUlsh2/1adebhnkoePlpC/tq2hXHjfsZ1cXQP2573a3umKr9+tGxzuPqfOJ1+rX
6tfY6RztEJtKIu35Uf2CcCnQlm5EjaHU38LOSSpji63pBNNvScpfKToEWKoRCcCK
OTGgj/7eyMlZziPhHWR8IVYLn6lnRmflrAFOtjPXb1bi8awfscusMiayLF/gLVdN
PQNaHiurCSapmx5FpMqK2i4j1NAvj4+5e/EturZPXa/7EWp++Gz02BWUZUCqFbmb
6wwM9Gf6Tm1bHpxRKaetcCRTrdauk6q2d3gMFoQGa+ala5X3L4oU/x3vJWYcTKvu
zZAuqwEALJn4MME+y3owddwB8j9ELHN3Ur4X2WUrwhI28JHVR6P3wGhgjqgixhPR
A152f0nAuQYNCVikZCWgwekqAKKeMF9JJn3tUEU+DXdAYQl+sZ0/k+6Lxsksw59n
OlV+qyAo6vw9dIFGNUnM82FDsPBjHK0ilmfRBybzmdbbVgn9J0UfH+R8aXlwaPBG
F46/ANyWkpT08ILU/ZzREroCPU+I3P/A/qp8Xrf/GdCZY3nUe//i3d3bI1kJnqe/
K6JbI+x2FF31r5ZUQOVM3WkKz75SpjlPoHc4JBvzWHcX1pouBSWAuyneaey23rkH
EDS4o3C39hCCC6jPO9Kf9597KBawPHPMRHzK8GbqPMglyLdYKSI1C3wNpZj0rM0t
sTx7k+2fPx4RkDyLBndZRfIaxr27O1mJAoWh6rp/X2OPqklC3/XKWVw72o7xkNGb
HV4BouxbQsPga8PYtWeCx3DsjCOchyDx1H8Wyj1RcuHsmpv85Cm5dzlJLPbZ3T85
vIETXTF+ZGYhoTqZZS410+XgmExBuI4VZHPpQSMUiRUCgxR0U7uW5pIIEE46UWJt
mSV0zFNd4HcxpVnUnfIQ/K/L3lC1yBQBlWsu3AtXe6Cx2kBAleqRC4DQiyicHBTm
tZN+JZpN0021vIrSztrEYQ67zacCRjWSURi/i31NfVM3MjnuMOcAoYcH9YQzIyS5
zfUxYiee4UkNV2SCn2dmCml0rNIFcwKlfhUisoXVKnyhUl+kN//0LuoS6mb02ii5
+og+F87e9uF2/J6TTqwZE5lrmczTe9vUJgbWbsfOPzBgVmSY2Ermg2K/anXCYP1k
6G4kYt0sdn1iI3H5CW/xOr231JUBt2nHRNzvPLUlb7nj8gRzdluLuOWyTB2rRFgC
Ceig8Yw8992dfX2UD0Cdmq7yGBGYo2XwNzfRQXaBR7xpm6Q55sH+Milick0okwQX
ldS/hLe4ZocyZRPalsZv1Sp8Q/YnkK6iOA3eoyG65Zrv4RNaolBve4DseUP8bikB
vXCOLrBPgr+qvrkp9bb/fQe4tb09QFL6XtLYyw5JUI/JHO3c8n7MsCK2/AhN0lXR
0EiL+l7VRbPwPk7hRWwyaa9FaQ2393MnADsU4YNlWX55Y0/8VM3u0GRO0bHQHu+7
1uILGuJXqAT5qBjQxoublDYgGGGLCrVj9Tv2QzooLczSceRAnPTiKbqEFJOEaV1Z
Iff+20v4btxXZi9IHUS/0EQ+ecCJnqzV/rqxBfC4HBuGWrbhcvgH4Q0wtgnIRS1M
6DokwZuYKMr5eLxR4y2gThEr9J2R2Xlz7ar3hv6ZvezqTDv67rBn0MkuuHr2uNCl
ipzhocKJC3gb0EStlBvKIMh6q/cyFkBCQ+7qzGiU0LCmrqL8F6MZ/zy4ap4uaStz
Gt2FIXrujWSUzOu65LDOHDyv7pBgbJ1j1DMkcyDljxA32gwAc6sxDFENpBVoX9oi
M23pLO2Wh1GrXGZxeY+9UR8724MorEvAfJ66R6Krjg+cpQoxSTHHDO/x5rtei2wz
fYKAb1GRB3VnFdr7Un6d4gBVClK1I4QZ64C6HiCx1an1lweYa7/1u+aVcbowZu2o
ymzcY2YMbj+e0skHXOpvGWVNrluzF0IlLliDF/7tcVF5quYQZ6XrSCORx+cNt9Sb
Q3X+d7soaOAPVPmuKIG7XI/JvlDIZinToBOmfLHgJtY48/1k8xurZq/gdb1Ww/Si
Y4tI2/jcvqe4FKmZscAhgs7qr+2flc3yw7aoYkghPHnS2TLGxqDBqxHW7+hRnvrI
HKZnyDtuuVQGq+YDnuLSA1SadYLHrdIuyC7KbpyiGk72zvnuTogl9o+sq7PvluVr
ze653H/J9Y1YUIlnMeFyq3+FcQycD5O2TGX/Ld6L90HQ9j23Cmvzno9D0Nmo0i7R
uWdt7+FIJYLsyiyfsadTzIAHsETMjBMn8AjGrkAOOIkTzKaL9x3pM4DeLCKkQdWR
kapmG+iZjkZ0MJbNbiBlS37TfsxMxUeJ9x9al+b1TR/ZcTJdiORmY9wCqhJ9cuxd
YOBNScHPB7LcpYD9niYaClxVk6EegqGIcJXAFLj2WwelqDgGXJ/4dFK31vtsFW1w
xTBx1bjqfFrpfUCEuBg1xQkEMV4owSUNzv6Zk6qNCxZ0deURYItIT/WHRowEZiS8
7h01b9QUvvmmhoxewiSifjM38TfhTxcfywnSZkMtumhdHtIs9H19dVvbUJ9yNejU
hxFzCsJ48SkK9++V7bgv2I1/lk05OIymOrUC52sE7tfG/2B5MhJcqLkNh6SXUIVP
XxWkDj0l/XCUy1Fw988F/XahTC7h687oatATAgom46sjJZjxmE3ZhrLkgNNYPUd0
V74UVfKejVe5WosQC9AN68KkPaE3McnztE30jmACC4v/rwGNpkr1+eRF37ZYqinw
vNB175RFAARXUwyiLm1JlL/nSHPvWpvjaBepMeuYBSVP5YVtsNtr1oviKdg+B9M6
xMlRzHXpVBv6UTo//3tCfm27/tLtufL7IjCO6Z19G7x7PaNLsmn6hW/m55nSXnE2
ySOCucVihVeveeCBWyxbDeIIJatdz+F8/3YSFBAquChB7z25b52sCofnlYsuUFog
gd7BcQFhgeB0xXDhkCbF27TnKZPO8DaKuIOeoGa+4EqqyihDrwxlu8huA9FCksFP
s0xm5Jrqcz3twQcYx6euWfArg/iMkTrRMhzi9cfE0G4QN63do6JgLEIe42gmURh7
njJ7KJx6ECkHfvZ5aVxvrqU/gY8hIkeDTjFDLJ6tXirfXzrKj9J40jwEdXboUqdt
F4aKIXiktmnjOxBEYJ7JOuCt/yhyF20Oiz95yYhEOq7EnRG2hsh2zF2KwZqvigkU
gCo+1mD/yxelfAWu94lciViFBJemohg8ONf/l7ZUZTZHLpwj6dzo5y9SQNya+4h0
SLl1bLlVlAO1srRO8IsMEo89OZBqRYQ1DARtNQ2P+OCH4a7skOfLqx7JF9WIX5ld
xj6ge5Dj4JB/8HAfpHA2Rj4rvm9VkrP6e/M5wj/CCMY0JUORBIDyiu0FOc31a11U
pySe9ZPFnJggx+cPYMYdXpLYjjAp56IPMFJ371ltnjqmihtWNFMOWPQmkLS0pJb0
lKg1kkvtcW972UrwgtJ7NiLduNz/fde57UaNaWPw/jUN0cr2uqSs5gPOQrJ9ze1q
RBJHtdrHhpRzMeUbzIgJckHzj8X8mRt2Ii8hvzSqkopY1S5ujPMYFkSQadMSd83R
HpoJzorMEEJ5GEDBjm+6iC8yzEByVcrZ4LW7cMmWM2rkVNSqdu87KVEDvhOSTgrT
3hxUeMPT/mDDLMpEuvpAtlwW2vi2gwJGrE0DeS6hWvhbCkNTZ+nS3X7IbSkOHGZj
/BoSj8stheJd4oNHa0LH747nZqSyTqT0XWHEFlrHlnPM5nRQiuBqMAaQdR5BwpQq
hOCPNY1OE5jCYLHUae5rmtQogyhPgA/Oat0zlJTEFTxl64P9i2oB3BNjDzy5AJNi
cqa5L+GGJ/H/cDGHilC7Nf3TxtleWv0/S3AQshfDAzxJQHTrzgB8t0PIlxiUhQj9
gajCaUtYzGgMge+8yZjqbbSQa4RubRygL+llwaanxTmFEOt0Kb1FbpB3Hgh6jUY6
DwDIXoqn7IP6nH47N4+EjYobi1KowLO+OKPTem2zaFjTYGqIycoKU+R51/Zw1YFp
XkDl1aCzlCGhvURXXVc62ENWDr1w74bxK9L2yYOrrxq/kqXJtLPyUatV1bvFMMBp
+GyiwcRD1vip+KvpThAzsaw17K2Gf8eI71dmZGf1iCFpo2O0wTzbkht03WiJKewB
w1NE6N0euW85ODlDzllYCbpB1U+AooyLU9i+pdRJBm2gCiDDwmtmV36utX/fjBmp
GESOwL+vDDRoqk3RVC78RXks3OEaCDiGnguEV6lAs3zSgZNSF6Uajb34WRstvnRx
dgpNlxb7v860Sj2vCFzrbx6w8nZVnuICr/yafVlbBZpikWU81kTHdFHDPggicx7h
BIdJc8+BvkqS1XUNxwmWAiazjwG/IC5f6QJXYmDDtEmshOMvjzad/WDjEAiLxz3Q
Z/3DCSLp+UpJTDQ4C2w/5oennFMBkKcTo4UfNxs9gAiMqRgrRV6zmFuwRjMBrxno
5VAWIUhIyVmbkhdl2BFW1lBvE+6qVJyVxRahyFTkaeCYUN65lAz7ul9WQN+x5mrs
wAYYN0LZO0oopmC5ruJO9ap67CQEn+Mgj9nPs89v3x5KB2RkpVDKcE218DJNOfWp
QeFOfAo5RwSs0K1COMXlDHhDGutaDXdKnlsp2AWQ8xY06oNUeu2U/O7BNAc8UsYz
oNzkKDbyWes+sY8mSafYQaxAy3tqUSBadLdiH/SbCwplfCHRZGGv8eFb294QWH2q
oHxqQnCt7z9idcP2eNL/DptrVpwFe0DFOCiBFWinoIFgGw3DIgYU4/fiKBbFwJOo
5O4SPNgCI4At7uY1L/MD+F+LO/Iev92Q/s5HHw82deLSqZ1ZzjK411GFlJke3Nn7
gL4ctaYpGQd0OFgrlZR7AdhjD+5DAOlRUCpbzedkb0gbebyr3NXMFWbWKiDU0YjS
exLUdR8Cw+Q+BPoqsl1x876Dzj0qgyqEM0j9aLQn+2DnoRBtDSiGiYMPhRLPHuY4
UCPX7GlQfiBo1NWOFsKAdgTsR3XTEaga14HZqPuCsiWIKVRvNx5uI/zVBsvWPcHJ
hIpf6riitBn9DKTxkhPxenmgjnLosfaXb/fjiT5+ebjecm3dk4q4z/+YS19TbCDu
uGC3VfAIueW/OH/ozrmH0E2aW55RFVUnu9U44VX8GvV2rnSaJ4IdgPvvhYSL/HuB
MFwjcAglJ0ompJGOE8wXhCrWa0udwGtct2olTVaiMbC12w4XNi7kMNm8E7GqebnL
VHnDzttPKbJIE+zBOVNSH0WlqS+OjfutJzem/jzEcCj3k0w/YLDn2gGtR7EsvsUR
pbe5AplmA2K7263VpcT25NBLwMPlZdUTeQWCB7kpUqtf4UwLb5+HdUW+ZYdH0R8I
0gcWao2Nt3VT7Tgc2XRxldwaQOUC9GAcCosMUj0MfAaejk4NeR7mkZQs+uHsfHmu
B/VujVeneEPqQ386Cn2QlsxeuXXm4Zjjd1RdIlUlf47uwLzF5anPdzl2km2d6Q9L
XODPM4dB8y78Q55qQUQ7oeU7tqo0UoHSvfADroUONMEScBN1BzUJKkeKXmu3QKpL
Vdk5NjcT2wG50FYFY/CP7ozF+pcUh/T/DjDkHERp9I5gXb7Kzz6K3HYX8m0L3z+Z
Yf9btzBxjYieXoTjh9B5pg/AM+EeNu++HR+3c9rOdvnN5p2L/+STDBV0n/sJ/XPt
zemWca2k/fGwmXnEe4B0TZvvNAkv6iF7EkXVvCTiZloeXVpPSnzXEhOZ4gXzsvdU
7qa2HzYIJXnKVLoWDSxwIdHXvL17HHZ/UHz27UlrDeYo5mnywz0+V3iY0sWzrYzd
eblfEWsno/3b2DEmOsoLfTs4M5hWFu3RX7tR6jwunCYH3NumJ2fDKr2HWZAp1fSL
jOQRkjCrpiOXfiHLynKBloFzlN+KCOLBmibB0Xw85ed7VhcEHs8oU5im0OPQ2kXV
xYdKJ3g/9vr58o8a2rG3WmGxlNtad6X12As6ag9ceIErgBzqgLEoeuSmL5ONtPuP
H1+b0Z61rCfb5LW9PmVGqk7eRWWzWoPPZJ820HqDX+VOHih+QslKuYoocAFGMkbV
80hS3X80ysBhqrzj6XdyLE/NxKyPdTnYGUjkdt4pPdV1UqGBI9rYdzIZVx4iEwVN
1EqCpP40gi5EEz0FIEx3du6wi41VcQMro8mgVo1E59nOMC5J0LJnavoacG3+XHmk
iSu3Ng46RBugZ8GHwOnm50/LRAoSpWV+cz1NXEqiSEgLmgKnwgWzWiXva2/gUImx
NSA0iVwMA1wfF+7s3TayZziqfE2ZJgRZeIUUO4ndJjUjERzJQqeAP93docy/Ka/U
WPhUnKvZ8vi0OHQy4Xxl2L8WgyXi75wjcH4U4IsUgLlc7GQ6JXRpEPTV9cfB4YNW
y7w25hqq2GV2pZLxnVy5oq3EonPaI5uoSxyA8KddciXynx5NPyvrjELB5nM9+qKF
2yBZ2APU2vuPV99wK+kHWFoeHQ2nmK+LU2sJJiVYci7MVslt3j8bicNB1ImOyrRY
MdQPBHElDkZVmsKSqFR0QSiCmry0H1U+GZepb9NN8aWdtdwLjlhVXRZBipe5AUXx
NDsd0wHx9jr3BxECYhu8RAfxg0elhQyC40lmF+a3EhQUN+A4SZrLjt9LLKSyr259
vYmnITaEaJ3VcTuxrOeesAdWhgEsCkJdDc/xZNCKGBlqjJlTKgbKVTwpydsVLL/U
rEMg0bEh4593P1+g/V0sIuHEoAKW2B+QLjMvwAmUCbPGZ2+SIlfdGFU5K3/S3yh/
ig1XHq6dPJOkbjb8d2TXyLyRw7x5JukGVi0KTvRRexVJxlGXv+8cygEuyFGkwFES
hVmheds+r7Nv5ivMqUzUGSOUlEH/na7+sTQdHo6QjQUTm/Vr/4YmGKuPEOGK7X/q
DYxxar5eaZf5o+4W/E0o/dwe4hyyo237sSae0F1NkNTHXhHn9DYEGNiDTtPPusl4
cQf/NwDaEXUVdENjlnq19Dr7JHHzG64i27CSDo4PsGaUs8NVf4gIo/dEz/T/saGE
P29jtKGIUaqMkfYJ4TKpTbqgYOolLGyYurrqXBCz+0lS946rFuznZCeRvccu+uxf
WcYOetsw0HesZT1/XiUIyvoUcAUnBEA+4aOf1MCFXnXCcreT0Xs2/GuKbClyFRKh
djhUC1+BrJ+6LJTZ3cSUSzX3lmAts3dQ/YJlfijdRcm3obfoO8DgV/ep0nizcpZ4
Afw2740LZYw5Fz9aVzy1JBY7tVd6+aa2maZWfAa/V/LRpDNGHdsnUh24epDAsPzp
UsaoJRcMEPdKEOOvKPA9hjL5FB1ern0ZuxKV5TEU1cM4ZLxtqPuRRpQdZb/dQmkt
sJTXk/fvg45QvQtW5duZNof7FjhRw4Ya4vo8Nh9fSGbW5bx8cJ2MvtTbhLWgFzMQ
R/Iv5sXr2wgnpuX36gCHJN68+lhnY4XbLhRZC+jHCToU2YGW4A3kkUksF0M1Ofh5
/dV4N4/lTr32pXWn+QlJsDZ0Y7ymxFVjDSfa59CYpuTSTxFd3BpcCbHPQi4JniVZ
zS/n0E2F1ER0erivPVqUhhfSKsokkfxTBti0kHjRTM9AmaO+AEjsCtAkOi6JGrvP
OeH11QnHsLWVCDPj9iVOgbYpjjcBP0jvSF11ckeSCdK16sjTZt8ZK1sJr9aMYNuw
RWPfuK13ZPnh0tabHc6liA7Ddtc0tR7NZX9bHJMoUcBg+tnv2tvffodZGiqLIwPx
klZaTpV9HyXk60nT0gg/274pNr9jbKxwv1OtR79a+pncVlleeYJ4Wq8yRgVTreBy
xHHw59UxdyoE/A8j0ZM1po1YTCEMgC5ivUN3ll0jFqTHqy6zodypynZNreqJg/Kk
kEE+rKOI7UGpbup0JwJEGA970MVZSm8IaR38S53AvzU=
`protect END_PROTECTED
