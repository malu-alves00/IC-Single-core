`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SO5btojaSMoBsOavBfo4x9vpz1qkO5L/vpOJ4LWhtFRHx9ziu1uhtXfvKXb9r1KB
DgZgS1tBuxlrbtoVCJ5bynqFUurbcXFj+bwv2/O8U/iIbp3xBHVmzrPYA+9BUonv
UtVhXV0LfzJW1VTdUKWlcREs5NOWDdkh8+Dhtz6PYjMCQMFG/0M0zUkBnxEz/c/z
q9SLDCaKnl4aPNRo8nUiKCvUTWHHzMjJRPqEIJa+sd/lumwIbr5OKWJUsky1/8ps
ZoyNypuDsD9AaC0TzNLSFFsrHIuN4EL9I45eeG2Eyt4oWWAAX/6FNTtaiyn1ylKK
sSM45OhEPYL+hkODJv8HcZVg2GwLWhY0U4lnHXZD638Bprzjp0Y4o/4MYW6akoQ0
X1VLHYXdEVkb7AYELTmgfpkODN+upI8q8R9vrL0ghOVC3fIV4LnSe5pyvZGpiC3U
J6LeWj6eIR9qwgtEjDlWay2u28YYguG5PJh8T42kIqx/Xm5ltJn4sK0apOfwA6BS
iPURkvsaLy90i+ekwnAlDTH9vP3483Po1fXY+x6TmqEkhnTOyE5tCSbVUV/T56Wb
1pRFkf4P9BkaVtH0Q1PmblqxxClORpCdyxY3GEXVrG1BMlGj35Nn+oe5hQeTdAYL
XDMJiDwLQ86UIt0Vo1xvFmu41cDVCxEpgHcKR+zfwLNUBfW8WQaD+IR1GaCqhmsE
Quw2Kb8kka+NO9o3s49WxfHM6NYtxKpvI99t5F99rGyBhiwvfBtYm9zgFHbJLyy5
hhT5FqRnvltjJBilIuMt9T7pWjYPyRt1mUK6/ujnjfpm0s83NzJAiE7xZntJcB3j
qkZSML70x+EcbZpA0KPMtHgBjhjb/YR6QSPT+5pScHmNhVwDgmjXTmjeAYnwP/Oz
MGdzhXwiUt/DUcRqHvHDkYY4BWpgbx9ASvztIWUmmN6E/BRo3qGQAdEzKw+DlMBi
o52xxX5iddeLziHEwXLS5nbsREFXxliYcJWp5ORtNZWAVUvqEtcAY3ocnkGilb7a
fX2PfYqrdhexxOhwuQ5Uwg04W/zsCNwucVKRhl6h0uUJVo3OcN1xKZx+WTR0iNp9
z815XP0vqDVbER0AooBpI1hm/MNqH7wEKwpiFsG/eIG67X5S89O4u+b+QvVNdKro
ZnGyXtNGq3BlefDg22YTAhgfjZA0d3L+1b4ypMrhj5jxSVcfQK7EIAiPnRWqz4wo
gnbG6dNBEhDSo2kLbNntsZMKenToAOARfaX/VVjIw5WsNSLVEzKfAvHxc30CZQ38
vCT646ixm4jNJzX97hiFCQPJ3f/a3KFcwrMGIyfta2tgnAUEHqiiK9yX743NE5vy
R97qciLiG21Yyj2XBRhbX94PHCX3eYOWm/yvkdR6DKsmDN20bH7cDSPRclXAudie
jCNEvnlEsEZb/3oSc7GrwMMaR4EDBDBX/xaiCSRK2YXjUJtFbso6eSCEU7Wgh+XA
NFW8l53QLZicXmXJJ4uDhcRrk6c3Gqbq8ZjuPfuOvkpL9YltpT3ab1e9MpwQ3dxb
kUmsQx5mBZ865JNENzrRvPUIDbMUji5iyrW1bC8FW71Qm/7y5BwmqwWpGigeqPi+
w/s8GkK45vUiytHxGi8rJvSsuasBXE6hQbJXgoJD++rlYDarHYv1QTV9RKoRrcMI
gKqIUOPNdLuHAv3i90qrXjYT22K9SJfzzveiEpTcM4+BdbufKLOKDusg+hqGqqHK
q302Z8OcWu3sTrOssQpvCzXAC5L5RmpD53QPLMnNvE+ajSZSY4bx6Z3hqYMAJfAw
D3NyRLShQ2QSLAKLkRysIGZ9PUlmBlyDA+WcxSL7P6wRzd/4cbCz/9+040FUeYLa
nEnLtTpyO9V0xZk1Yfg6K+BZGMhaVoMp4yzSQHz95Sa6MqcHUmjRLzp2Alg4igos
`protect END_PROTECTED
