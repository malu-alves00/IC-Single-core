`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NqiaGNiUBpE1/ZUMRwn5dNYiT0YyQ/Axiwc+9CaB8E3baQUV11kiZy/s2+4rTRN3
vb/6RFKeoCkcZhgEJoRoEECV7pRyOlmUbnoZJowWjMXT3USDwDg1c4DTrNC2FjqO
fPCANmzsjpsQ7PPapJe6ij1OMSWrYrO83UVZLZ6X4m24oHuPn3XapwASUoHcvoE8
q9KVKyNBvXUI7IuYViL8U5yjBWaVU/M34Aro/yZNiG4JA1uPtXEaWmxrrBMKf1RT
gFUkr3yYHpL98f/XW2wXxmXvG15fn5OOEN80s5LVkGCrmEgfwEau6y9PQSJvg+ns
7dkUpFqMU1GJ01y0uF5+HiFTbIw6OJMWLBA8wZjREyq2/2gVYyn1nOjsqRTC56cx
ALz9hjdMuzNTKFIarU2KMNxdT6LiRfSArpT4hikgblFJi0N4jHwZq1oc6D2/IuPt
BsEnI1aD8/qwTKFsUiZ3ofTck2sDXlzlp/l77MMb/1Vmv2u6uJa8uqOonSX6Jqoo
uSmxgLhB3G09LqSeShJrkm3iwpQSPDhkMCQA2/y61/dBV8DWwDq3utcgbe7wSqR4
zRbq2HEaGMKWSf6z0dJT2dKXRfkPK+khEfbrNbFY3g5AfywH5plJ+FBkFio81wGh
8DnMJx/yakwVgjvvbdgpJARKgkphP+10YGmPQ8/RD7Kgdbt23ecKXAeJ6A3c4KJD
cu7Dzg3T188fNAttR4jE9ZP6TVq184iVneQsasqdd2UPRAIwX3oFvicjZs8zlUFj
jMvv+auA2LYWcAEH0vhJXXJipTjVmSM+2stSaQfguP+2jDfkYqgA315Y9cIvmA+t
HJIlOmIK12jRlvnQ+tIIokCHOWJmLof3sGcxSMwk/ewJ6A5ALTZeFu34roNTkyQK
ZCTwNt+q36IV8iDejYLuFh5NBQLn1ASsnSKo91pOAtYnT+I8u7SPnXKylCafs3Tx
v9A2NiOeCD8SAofLR/9YyAExEj0QvKJOCoo+Ovm2twWMfMXADdN6pgFGd5MpZP+6
NSFfqqwG1qi+VznLAZBdjmFhthu93KQgBIXsYhAxTMOrarwtF4PUoJ/l3sPXbGZg
tluCnfyJNXocO1qjC7SuThGxeI3M+Vs3TAc8quGdlO3FxtPCum7WlFTXOvrn8bDu
Gs9YkBSLqhdydBQlusRHibzsnWeTt5bPjs43GuQgWt20BD68vExN5LEDKVarhqBK
Lq+nPhXInnVNZapMlyZmz2XOoYX85NqFtgykcVwILImHatkrXo2qR3LFBkYvuFpi
P0wsXABGyVV6XCr5f201a9jp9IH2ldOYX2kJIJxBF5u2Ln4Py0aDHbN+YAVeLmHa
Qmx2PoFjfcSoLpGeZ9pNqcaZs3KUacOO43y/dYFnZ+nAREOc3f/mqboUipfiATI+
Eo3TIul7XIh2fDCAj2f/UPVoGc2u7i4W9nECrw8EhU5VHLKKdDl7+uFVeDpYnsIY
cJUanoWbtGarNdKGO+mnZnUjjI6XB29Tz8Q/RW0SOLDrgThbxeO501dsADCWji7m
vqK1qQUL0NUG7ZPXygCdUrUBeF40wqYSAuhYQbcRUUCx5UVNwMhBlVryyZ+sxUkf
WGgdOsGoyS7DFfze49hczNxstV05m/TjjAGR64lF6XQIgQbYN8jOi0X/T368dMtP
JbZWzqGR7X20QkWcKqA7HDaCBew5C54r8JbWLM9yFP/IaOrPbqNuj4p+WiP8cznb
My7S1S/hG8QlDdASLyfbPpkZMGvpV7thjXJxiYKerE335WeJSYTS0GIbBgZPzq6v
bUCH63SOW9O4HTAUKU7e1Wqvikt8sG0GTZyTyOPpxpVHSL55UXbv9NWhgzdpZsUu
FtJP1NklEv5/oEjNaL1+fgxsEvSolOrvz/IFvlrH4NPhTkb/1XlZ3eY46aWjx0Jw
1WgSHOIbsGOOlZyG3UFPRXz3et9tBf3LXI2wnLPSFzpNDKRSZ0qDbcEi2Nr520+c
1wlu8g0ghk8hYIavtAwyqROGuHSEm+6fXwLe7sb107JHSg7Lsu71uhOkU2alOyl3
ne8lOiwqXN+H9+IZWF9UTUYLk1KM8jyC8Jz+/VFkXs/1s5KzB+G69NmGpp4iqnRW
xlGvAVI+pTu9LvPTBfAiVh6imhFxRz7y77HNpajgvN71cP+U/gZWQ6V3A92OU8dI
9s5zepLm0vt/UGgeRrAzFzgu1S6nT6y/xIwGeAq5/lghI9IuX5zhIOF45mtUfjn1
sNDOS0c2iT8RI1cbUs0K5foNyKxmZ2rigSc6isloWnXCqJQamoglYHs1nkOqSLbw
0WcX5B4eVxWjvDn2ZSkHQ4MVQJLHl06pBqme7BtgPrKInpBju6T94ABvfFdOUzzf
EuI8DfrXAjPGJ5NveYWm7UCWqh0sdOVhqzAnAsW8WNT2hvoogvkbWW7fecHReY2M
xBttKKN/+J2nreBtDBAhJKeMkQSPpUSusg0bZXRiARh0UNiqTeRbKhDlfdQd5pHs
vxZyzia+T5A/bS9JAPOzNw==
`protect END_PROTECTED
