`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HjrFpiXzhTWyElSSxSiRYE9n3x94GC3bwoGqWaAFRgJFxA5hWxn8GZXPzRSFCvRf
RYl3jCCNTlpyBbddmWqrXw8EL4K3SI2PACcZvwHbjGpOFRntsov8xshpDxQwlja6
2sQBDhDPen9s1jb1g70FnBVQDwpa+9f17UOdBHmt3Cv/qRwI6s0d3OZTTy0BrIcZ
bmUa5wjgTCKdA/SA4A6cZ8X5h8jtHOcRrDIJo7rGagpLhW74WOc9J/k65oXVIKkd
QPOOn5OO8puGoiG+vx0doVwSFEDDyD9t+yrcBNK8XMCf1hMF44I4GyQUAuCEaUB3
/ym5r2K9QP3fB3sCUDI+LOjL2+ln6+iY6Ac74I/BUUB66nlzDu5u1kY7dYkuXbG6
KvT8tLUBkCAt5gZERkPsu0qbtSoFZEtVDIK7FnATOUZ6B+lNd/1BuLbT2JqjOGaK
N989P7MLm1RuokQlntloGq0dxdTTUeDyqNuZrbLFmj0uUnzdGdWHG8H7Ylk/YJKg
HhMPXSwhk7QPY9MOXQv65bpRBwKrDfjE1QuE+n60XXLAluXnOFc0FMBfgz2TWGzn
6UuTc8cYEIHvAgX5ecI17dF6HExBXlr8d3iKcOgeZLwBKNMhv9SkMHRw4GMN+tYj
V0JSdFXZQMG/+4zZpR23/bKDrl/+3APqgurKG1HmPcGMONdiDKh54w5kZEBF+z3I
076ExHgNYt8MmaAuEDam0ZisBiNpbaMyaLsP5ld43084DBOarfYSu1Ys9tkFn/A1
yL+cc6+CEvf+f3WnPy7E9Mmhrj9/sAHhBz5S4AMHUD63CSnokDTBLy0IVC84mr07
peS8n1X/0hOW6Gw++RGM//1S7tG9bYNOf3d/5Mn5aRJsbEnt7EfcDznz5NBpyWR2
8Evbx5vGFGgyqlt6oebOTu2Gj/+wAQTzj7a7hh56SD2kJQYhSq5bfjRXIN19JgaG
jEOIhS6GpJh2odXs4hzqKxPsHr1Lmoj2AMVP21aYuJUZPd0PKA1AYPCZEiCg0RFJ
HgV1lS+2BguNyHMMsj4AoRrkolZRulH8rkr7xnO+m7lgRn7yX6GD7c8vpNbhoOIC
4zg+DvcQ2mXy0TPBWZYWXxr8rk8uihiYMH5RPJbY3GxIm24T8bZcYi4AIA1gGDOD
UFtkFcV7XSSOgphmEOnVV0+PlwWudmYLccmjL7ieB5wDS8Am9e7VOelvzctpiCM7
14ZjgWY965X6THDEupXpB8bB3ITPb0G+QnTNRgC+7lRw4L7MAtThuCI99v86A5eP
YASNxSQ3HZtqeglYO2n526Y92XTYO4SaHHpdqSIIqgRyIm2jPaxK8+q/dv+xExia
C53AwIZL2SJh7CD97cPv7+8K6UundG0ZN/g//KoTCSm2jv9N2QP6YF3nc7S9gU+W
WhZgDF7m2qvrfJSz334pheuR8tmiJV9SjCfEoRVjhYJWtbH1lVyK7cA66VjKa1IX
IBH/d18eKvyHACHEgbcJ1qzy1g3y4a8uHxhcERYC5LAjv+50GsWjVmvNJCpznmRp
Xx7/A6XtIUmd/BYgAVyI0TxIWcllXjDe/uMldKJWEQ8PzEoSy9mcZ7oFXbN92eXu
TCDyJLLGE2Q1xed23VVY6IzIP8Qm1yRERGjCZkHlu4eodWm5SrRqgnrujJFsxNQ3
viPgx+26a6OG04GMP8RQlqdsPkwWN9CBvDu1A4Ym9TjOnPcvLQkOu6kw5/SIT4yl
4eslmTaCXdIzwDsNKKQ78a6lWdjyT43tbDDMMgxrE8L7ywt8kUcPjKp9hQhyfJpR
xqjiYqFI4yM6mxMgg92WZno8CHWH3qIb8U6Ow6OOABXpb66LNaPzut45whJxG1lJ
osZirlJ54pakDjjx5aQ4fJoBUpSkXAFUvQt6mnjbgp0fm+Ul7u6dNXu1/6fOYLdA
r2/xbCYnmsyZetH5xxZLBh35zcf1+YiTBecuCh9x2+GzOchVt//nUpPt9OZXFJn7
Syc6Vn5zsjXHYcUC0dJjfqYK0zT4f8hlg62Wgtmw8ph4y29Lo5czuBtMXrmTrgkC
Yq1onnPrEdEYk60Xc+Dr/p04SHEE0X+9yPmn+NbMdztdgQwRg4xzvioiIKP5LV4j
3icDUJDnb5l+aU7/JBrNRYVQy9QxM7/aJLRmR9cC+od82GSxEas+eldZ7LmiPlwG
7s0Fjvc3F5cErUjRdJiXzeJxmXRdGN4nyr0g8DljfnhvqxQakpETzSy/msAslRg7
c0zrTpPkST8xvWQDydBJsLgwpwU00wtUiGmkUSlKjpO1Avjh/TilCiPkhgbtl2Rn
elGZL6nzsAqtdIt/NpMHIGovpVRf8iBX1p/2ee0soEVKQ4/Xzf+7GQmqtw+VQ87b
sI2yp6v/H2kl/d7MfHYMHNZYxnlN02NjypMMG3n6sZTmITPMzXRiDo9EzjSANNEm
z5WBqaRFQtirgF8//7Wm12Yz18u7910x5uHNi6Z1pyXz8xD8Q0bAm18zgqAzxiqe
uDD4K45GkvVPufGyYY6GBg==
`protect END_PROTECTED
