`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/vvGK9kTSqZM/7LjSCqSm7xy3WoCT1lzpuxT0XdSfad59P8zya9thwhP9dce/Uyh
Tkt5UTusHv6QlB3BcC8R83S6ZSXgNwwLYpC2O/YdjF7SpzBCzDuDAWQAm5ddFurI
XY0iCBhVe/WOcQtJIgY1Y35PNFzhJfIUtJosrJqssi3b/SYbqR+dwZGAuiBEcPrU
9wQy0j1AcirJ2e5eiKEotaL/kdQ9MCtwMNY91jwRAWSClOsxUiQZA5qbWhXR7aGH
7koqusqz1Jj2djMZ7D6ZgCzgGD4wljPe/TM+HwBMqV1Ci94yug0F3/jNZ2sj/E+N
Eb+wAqEj/kwY0r2qrITLeq30K2ujVDn94/sLiQZLkwmQbSYv5w3qjOlXTnei8e1v
iKJg6GLlLTDFXnSqEjTHty1a/H+ocT+1Qsmtz5bIPLnq+ZyYjkUIWYIbYL8T/BrV
k3zL1dAoHWabdS3JjlD/eD/lAv7EjHOq517HJftTWdMLzIvt6HemNcoUmux6in3u
0c2sKufJ/OagOHKWFvBdeHpbAw/lvpn211pOubmictfNYfDYRnGpFeJoHW+AvCOJ
TdYOfi/IeSJUeP+lYkOJJHArynBSebW1R/dcAXDmr07ZyDkdyAkpK+PLhVqdfuYP
pDqDPWZVFybyWRg8lFCZR/4K+qn21m3etfaKXMLYNzjVPsfaXcerJyUBMMa9WqUf
fPcTdgY6spOr+ergkxkDR+UX43RvlcemzbVIgVAye+B4IIWn3g6dVdKFLXupyoVN
K6q5uRPuXz9UG3setWkmhyM0cNMNLO72aVeQHq8EXduAC1G7r9dlJTCmojykuCoH
aUWao4sWVtuGfdmKv70Jj2RzsdGYm00oFxKHD/OLUcaCK7H2FDhHOjvlrSjpD4WY
a5ijUp9R8wIDQHS3nacwv65RF14ivy1kCSk1nxmNr0L2wsgtqwMKuI6p/+6zcQzA
gQDtSRwcmw+/c+tM3T3h4QUyUjoHC03va47/AEC5BFEuZZNBWgtEphBlrZ19xALm
Wcmiw1tq3xM0xygonx/upDSxYEAEdV2g3Waod50cLf+3epMwn6Omwb14uAN/BsA6
mKaTVEu7p5kAcYbdwZrbc/OJw3htXgJlWiWGpE9Zi8idO0eqEzeZuWtdeg2xhVBL
SV7bHjCCbXRSz7to2FXIFllc1r52Fuuu0M0s6TJAlnt8LiEwuaDYxa4I6OpwuYT3
o3yq8dDaYcK77hVZUGFjnDikb6AEn3lFy8xJRu3jr2iDbPuusUEnDc5CP2oAS0h/
+JnsQY4bDYMhGW/VsKrs7MdpOcTkw2OoL5ZQBoj++V60DeVtw/rdjHQ3tt4GIAXP
OwGpMvFuooiUymW1vfbrNCl08v1Ax2ubr66VYTDM56TJBRgvFNYfr3t+mym5Fkdl
ob6PoHgUNEFThN/IDhOVkgYH7VMlLBQ4qBPo41idhr/plqeb9PkA190hx7OAQWVu
Mgq/oxqJ8l3PQWpu8zpJsoUBZ9yGOrYEeDV1nO96KDqtdKpu0oh6XZpWzCw75gU8
cd+OyN/F0m71NUkJzx+9k3sZpnBYPtqXzyK0PZ5fV2XT0OGI7eA3znX3/N6wEIJO
sS2VTpWPfWgCu163ZQ/CzhQR/FVHlQhkBBvrFAVMPG8EZuAYF2is8bt2FYIn88RL
bgxQufCZ/SKPZnigqbDe+4z07DjhijmRHsUywaR1jIypKj6VpV2ndXUnHAZj5/29
cG5/InD5XdonxEBLUI9x5Q80rC6R5lWA9cH6gpwzHN3PBPgcflcpex0OdOqWvnnn
q3KqIAv97xnjzjkdUpUaHZx+m6lHr1xhGoS7lkAqfavvE5c3gTCjETQfn7IvHeL0
a29178sutP7G0jpXhJl/imY/A+FZqZft0S8FOQt73l/W28hJ7+9Tm3U4kjlGA2WI
Do5LGAojoST2/W+iw5cjiwcbZIFhi8Cj0Zl2ae4RoqLiqh1aExl2SATyA/T18DEb
WY/k4p/CsyzAGvEvtIbOZZ+F/8wK+7lQ+A3+O7n43xK+1lH+5wBXanpMz7uPlYOL
ID7cbnEz+9t1COxLBW/G84XOmGya5nf6YTEIW0PyikdE3y3CMF8sllzlTQUbINzy
0rPrfHJTaDlN0lAj3wWo3r68/RtFDpMJdiEi51L8bNJKYQaa3pBNDBRLanSgFvSL
tDoq2c5u4tv/w1miuDj27KVOvr27v522UzCcM/G739vQmD03/isHmk0cO83l13P2
9YzhSAvclGfN/K6T1TCFJxEN1zMJNFQ/3U9LBgkuPArzqDzgBkszbiYTn3NRvKbV
9C1pVTZ/nMpDugP77KBqpCyKdd7nRSRLTXDzddJZRBV9qMrxPXr+lGJA9Camv0ha
jF/3bo1tZ4OtaXOBJtZxQHQiFY/r6YWdRlv8MLyeRypFNJjTEYEAyHlKUHqBC/Hg
WNfydfSrQ4Bt9EDgu8gc+z7Z7HXG6n1iwqMpYP3vUCjJtmXiziX71e3vucyI5qnJ
lcb8xSqEhbof/kewDoxy/GkeLczfT0fztjHCZ07RfYsigFSRqgxANNV4Wr4eM8WL
yWc8RXZkRlm+DBQNt9p318VBHlNrA/VhzgUia6RjS/Vm3hpLr0s8jXPjWw6f6pxy
yZSd47WNtOrW3aCrOf9IpUxMwwgOjj2ntIsVTXk6mV/1GKfQRcxkavcqYUqly5fd
C2zXOPl4VelQPTw6i1NVLcCHfpp3U0MeqwpQB5OBupijgGZR+sHFCJ2WX57m+bvV
y8QwsIAXkxlbi25Ea1w57jgxWKg+myfzGUiFGbzV/aRxWvDacanbbGS0Oy0K5po3
nEAaNllFYdyYmTb7UFwRp7DJ20E6ym2MR17yIsRxSqAj2Nl14eOIi0osyqqJdbql
RK2wtx41tvKH8azY4m5xyGeqAjQm9vVYaAYH0ju8sqmjpS1HmaXvTIXnfNYV53pK
qKkDZVIC0T+AyEjknSIEc+6DfGxxfZZ/g/JG0oKsr4a/qgvnrKYTDKXSmYb2aB1T
D68kvNxHezNZ3GYIIJU8OKotWRchqHaijb8z+lKHAlVYc5J3fmVSbCDjXI0xIT56
vm8RndxA8PvgA1OmT5eEAOV1juvrtoStL4slKjjDD39sclImyusXt7f+OYMFI40+
z/MAMv+lppgedDeO8z/6vy0ca5F9tI7PMKsYB5TZDhZDMMQdWj7sODQ6CLKybL1b
k9nb59ru0bsMSmhCvuZ+UN9/VqCZqKxIZMT6s9ltk5VRHL3okCW0ZfLma9y2QROw
1+ywCFwzU0tejwNlAxM4IwmHASDIh4FCD1hgeSgpzFjaszXXFxewo22Djm1eIhAB
gLg/Z5//HpCJHWwo6ppeDh6Gr0fuWPCGRE2YrXEetxKnKciHQAEVlLBXTyD+1iV+
ANYeNnxEPnudjhWxbIq801RbdxjBnaj/LcFX5m3QhSXemoh0q5efHr/a9Dze37L6
QiG8091eWhFN+nVuT/3xIxATuV85Qo88rXE8o1xyv2A=
`protect END_PROTECTED
