`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/OeufWA6yjwf68bhInVw4IMNnYPLZpFlF7Hx+SgcW3sAI0s/8ZyKho0OKVxftDZA
am9jMJ/fTefy/aQy3RWSQa67jKkekEtZ6NMB4CZnccSAERN/hhSs0aou5SFy8gdI
WbmpSuSYE8/QpVv1nhYI3YepvAsFtNroNRoPZgCap1TzqIZuiYqP4Sj/ZFK9blqz
JIp8/nVlLdQAS/r+qbIFE5Ss5q+TYO5WYWnGj/sBsdlj9hG5lY+IIlSpky0vjqvm
iz/vCyWvaEoYa7QOXQ/r1yZ/hhgLYJTP7HzxLzuLKfIweK/mFCY4IgL6QcW+uG2F
4iB6767HblC7ziAos4mkwlDp2cE/A3idXUwiuCOHIRgr2GcPs9H3HuOoUGN4994W
flJwTVuZjfjmj8O6NXZKjVel6j1hLr1LHB8q97qo17ujA5Q/CxtdUDAxsuK/M6Yd
LOdjRAajmC4wJ/Cj0XFybg6EsZijR5N8PLZVf3Act4dHvIP0gMp87Nyf8XSV0eo4
lM/07O7Xyo/G1CRfldxGNek9OAXCNrIx8AuNaeD5v3815NQtKvjVZQM2W1ME84zB
m/cWwmWjLbECtBFoTIG5Fu2IuEbIX9aKA18wc84z1lnJLytVxs8g60F0tPKk7/Pb
9M7x1W686oQYZv2seZsaHM0GD7MzkBYeu+YJJ+x8QFcmrHL3M46G62i0OjdV2Q+p
QawRwNCyYAlmqEzP/IsBaPuckGVhVQfCUu8KHLILIstH0afMZd1fbKhc84CflRPr
XxEpBE3F+ySMWYa678hofdvjsZ0ZwoK/6M0wGUp5TybknY3soitTyL2iu+JU/aiN
+KK9nF0gAjH63vwZU8vskoKLv2M/XmC1E8/0Swuj7Kjxe0G+WKvCw1hqYcKIQHPr
6A9/V9rRAHXp06bNMMMcZ7ujAZcWoN/Q1hRgiHTmyA/i7xb547u/VRMK0lFEwYml
Tj7HMlWzOwdoJQ5+qCama88d7s9rv1+l5A4LKz69JuvzEh8AuGHCHB/tOJLfC7qA
ch7tvN8RXQ2jz/CLDYpetMWRIJNJc/7fHgOWBkh25LZVu4C4k0fq4ee9T/IRsp7c
0wYyaTtZyDAgNCcBQV7bqDWVttYIQ82LxCdZspffXvDHwdKV7z7wtaSMJWQrBMgy
PzGgu/TQ8I77lnbX3mTqDueMTQvo3EQ15oqP2viHhPR4dj7BamC70g+3kY7wVYdP
ABDEJLjkVZPxbqPbG2p8n31FkL11NEJKPhVr7cmfZ2BmOhQ5o6YA6FdMPncR4Q2i
8k0emAxWWLgeEJ3e3LZ0KhWD41gCDLBn1sGJItrG7hliVXhP6Eciss1Grgfk4780
m3Y5ue91glKq9EvW8ZS2Yfzgnz/Ow/PaYieXnIwDvrH/8yc/i5TJwRoDVZmSA6xz
PnxSKLJbgsIuAyPvy+/uc/4OTWG0Ch+cRytWkO8oDZSzynS8FEBmKKXTtVXro9ks
YRSgMzy1YyMEFxSx3XPAkDems60W4EoaYB3ZhVcLdqaVRF4iv4Mfy05XJpb8Hn0i
510gzMkFdc0zYusOaNEDh7fuZtUwOARtMbnb9uUZ8nN7KLqUY65cI3Rd+AH6h5Mb
lmniFxhKouRKPftfCZRrSV010rE0TtH4mBlPipRFXrXUHrnTFVInCV2AIkslSXKM
znyl2rl/FXcpOjpKwlPUJrJiq3yg8T8KaJWN3E5goG2rrYbOHjie6/cj6LAxFcsh
/6acsbigmQFctSEwnzdXATklQbChd3G66M+VC5oCiFtABCHPLxDSFNK+nyQ1y7cY
3kecOFG4YkpS2vN1pHpaWLUHtH9U7FsVn9Se17JbtTVGryl/su7ha09YZWUnSpVf
+YB2Tya0h66Y3hV52fnsEetwUa8niF4FOPsDybgrpYzvViHHSVnOaL23pRNBcQZr
PyW+ftPqBhvvAE+GJK7DZVaapSUUxWnWtrVJPq5sQcBbg6H0WuRdOch4X4UjErA5
QUUe5kSTcWu/4qv2C6sZUb76rmELAfjKZW9IWOnPJJ5yNzgjyFcQ9j8HE0lIEMnB
Kg35VIEtYANbMQvH/CJTQZKaVT8sx59jO2FmR6v96eRT5hdT1u0Tkj/fJl8NMgie
ppAvNda+3KyQN+pXgc+xpcCTvIL/BJte1RwLxIp63xrHSIFAWp+PNrFsf2nY7MO9
dNICATbOCHQw5n8WQe5UluuAjS11MVnpG4Eu13aG2xmnPQ7tYiOyHfM9ANLtHJjT
rH2rVH2FSBv0P/WBaGi+6buaHb50XmwmcobCPFO+0r3Tr9bqkV4/IJ6CC42AXGQx
sPUtOfaEDWs6aL1B5irH3OumTowwE5wMZoFavkvSGHIQzrAT6Hlstnaw9fwaou5B
VNBknagRX7HiG5g00E6xCV0AcULRKlsdAn8EsrhadEHs3SEdjXiQxjaJQqkI3pzx
5TVLL48+3yrR0+6ydD3EnCwIdF/4HUrPEP/xSoDEIdEQgw1ST93YG5UORDIxybmZ
qlLUOAvXMRwbNdWknc7uULHiXROYPqYJg/U80ZGxIOQ7wYtA25HFgrDevYfa08Vu
Prn5XGgsp6rl6YkmHCA6owVuAXdwATwisHz0ZKp4a8t/nE4fHlUqD2qZVzTs9r/b
Mhpi+vpyK50hZrZnrMBpUVksi2xLVb+amKc4uF6VOPcyn8Lv7id8LnulYvubPAEW
WYrnT8H2b4P3crr2c+j02aM62Axf3L9g83N4IVFU4kPWn2U383emYPXc3m/IiPlK
9IOESdKyWsA8UAM3XtjCoWJiDlIrJ6zhEJaV+0ykkZ01nH0pmm6spBQ1mcJHPIQy
XHnUsO9g8/sKhr3ww2zB2aPH9YKyJbHiStq3noxo/CWdtnGZbwf4eO537mImGSj6
NopPCoDjphjBgXhZSoImKJoOxMUtNNo1EP9+ncQbbzMmjvtbxUJQrnfQUFYwDtc8
PERlHf+t8J3W6/Q7MsQZu1jbc05h3P4BL81vx37tgXSBSpTLJ3lNWKR8UEeOVX+w
stCtqoOBrc0Ea/VVogwgMeJrqpc9fJaSXF32JPho5jXxtRgWnMVEB1Nh57zjMZXW
4HsMlUcbK+3FjKukmjAMdtBoiOBoHipGnB5Qhv5dIEAlHw0sRVZpc+rFrMLhmimq
IUVIwkRlpDVb6cBspuq+FT2S8E8L4VpkEHIkLJgxPfl8MSX80H5852PKOIPD+bCp
Neb3AI/lhyckJnq9ONAX6pwAKtzWG0rDgfdEXwKvt965U4SqQJHioSh+fsyINJUM
I2VRc2bqnFm0wRPO8UtmOrkQb6xGAsL9h6MiWPHf5yQwpWD8ZDlsB69O4E78cCpd
1M68gCVQDeIvG6NltTqQlqxx9Cpl7HLVa0C4lmJxdGOzA0VLXTbkg0FutnMZDpRI
bduB2zptvTOZfOLeNj6g9NHCuZc2GEFV9b5fYEFJTI1hG0DodS0QxgKoDHAN1qsx
xVrKwK3fFvlKpiNgpCAC9BrHJDtp9NwtUgbudxpoCaS8zcSBzcESb6sFYVkpuvjo
/sLuHfZWk+fs91EW1hAgpch07YY6Aqe1LNXcuFuLqTU2bfcvtO3OuqERzi4omFZl
QXD9GQ2YU08nMblQY34KRPMhXQ3NA/jyw3f7E8zirzM6iXABUmRPe+VjqqLDPP8A
A447yBQ5zGnRcMbdgBDC0B3V9KAJ0NHouNZ4VSO6aTY5VaZVtjrYoNF1PteOH/xx
25Rpb5ztdle+zEkQq0/Nakj4BROZ/PVv/4PljxK7N4BI476daxgMHTxUL1VkIu8n
QEW2P/4sR2VpMc0WQJIereRmA1I0FtcmIRXb5jpiFRx2d+jjBhG857eR8kLW00UT
a4PYLVkX1hjwlD8yabL8JPFH3cUq3uboc73zfk22RhUUXNRhUSpiv+cljTuid4Lh
NHe/cvcdxujjYavAJ7+wncLaBvPr6QIZtVkdxLcQYjPAa+gI6TygfbPMgka/7VP8
lVLOumHzSKu7SJN0bjlZtJ+HG/1khsdi9p5gDd0pbCuis8GdRj/wxViTi+mjcUiM
GZrdhmjR3jkveEdVv4zO5kUl73ogxSOPYKCqEt4DEFrKRFNUNhxv6UxayBoPyNvB
ipIqzux0Nd6gi8L4esf4nav96N3raNOL03gKfrwnl3b+GF3UNNJrRNB28XTSHpsQ
EaRl4PdoDLa1A5nJwWXIU0QduKpndfC5n68W415R9c1zmJRgNXNpvPkHxwDI72TL
S+anDxaRnYnQL/SsmZmHt3H2gwgKxXwsk0xQLzGmAsxcP+3HVJY0s6WIw0nk4L/5
BiEAGZCLcr03BPnHFeR6q0fQSWtAffuIFhcBTXvd/fM4iNhWJAP4etkhgG+al5tA
Nx22ssyH7uLQ6V06mDwednadRAz6mxuz2c8CCs9IRp4Qrc6rwGeFex3wAB1ixMZv
Uu2WscH5pPuf3FkPGFBZXCymmXfeOoUe6JS3sEXggUbKK6+a/QvP2M+5qDJ68YiP
0zFuP1sjPcNhYpjFNKGEH9y4vIdHJTcsa681k72TMRZ4WUdwO9JZk+D0Izbb+BN0
nfXzvCvofkRD/I/9bHEKUgD32WThi8ky9N4RYicdshe0BtP2obEhRCE19SOsfoMq
9WnOEaxtafXB3OM4OTjabEUznDZUcTclkVBEJ3LBMdPPT4CenApXWj4uC5ZUk7iR
ww+Bg4IB4yKy25X7DGVT/NypxoLNq5uZ+646Uf5VFkJG9DkhLtp/yPrBaDcjPZx1
92Nan18/JHYw4PqNs1kPdvw3JZO49zlbymgpMLPLz89NhZbtFPhD2QgL2BPWUSy+
b52sE9D0ZiZ2WMzBvElzmrn6Qjr8pJAqFKhp/V8q9je7w/+1qDQeXDs0VLBbkNMN
7TcMZS+iS7bOMtyWF8TDThl+gcQHj6i0iyYTtSupYfMQm6tp++vLfqJrSfFeDaRU
m+UC/AHjNfW4EPlcPzMrnIsg+vTGNdEHFzSQ97gLuJoKXuqkQuaR3cRieogQaW5j
bHC1+LvS+MHrx3Lj9v3TMamMeq0UZPsbXkBjju7MtW6iIjUUXm2d0cV9K7rALsLE
b4jw9uJgUZiwxhT9CJEBmjQpKXUE8Ox9BY6s3Q+sbKY4qYYdPOLg0J2NIi77txlz
1ipoNbL5TzNUc6k+qXcIUhOIbFJiEwB3jRJFjdYYjtG3BwjR+SfnBRWWIFIPh2Th
4eNmwD72GmujVGYsRQjrUft0KuP5Qw/FkVZ34aXPa5s11qAEJ7bXovxMLBVps8C+
wuh+x72vdsATOPr4dW60rFe7UsVL5EmiBBjaJbXP7TsIQ3F/ZaxxkzvsU/NJQo20
GdqivgX6av4TcpN1t20j0uW5SdTmmHlK2gNEsvBuLZ1SE3oIThBR3XtmNHjVFZdd
rbzMqjIWK9gJlsRU5tI5I4clpuhp3acv1PPqpBEr9GrmuwGeVcGr32MXqc6Tsq8O
GpOiH1+YMAgEpJbEMePQj48Yiqthg5oRp4tkmoukbp9wphd3H6rafmbT3VVnYCjD
K7w3LOGEV1jX6IxScVuLXt/qI3AZPDZ3WTnX5EgTFsgJy/HZ2AGyEI3KiLxkQm/u
gXT/p3gDgRogGIdklwGYcKgY4nXFIOhqIzZua1nKxuaMlKZAmMvq8bQ6zy+6/7nq
A1vSCU4v2sx7Dv1AFKeLdc1ubUVuTWUxOZxYUEOO92BfVPgdJi5l2dYCSzt+4ISc
nD6M6IHmK0zs/d7C8kO+Uf80aBn0ozPhxZujRM+Qn09P3mWxKU26IfbNcJSdohmj
fWmR90aJErAAucMGe9tPZ1YxDnhBDXvwATO+118o5zpalDjpBbrknsj/B/ubljed
yOMTjRzqjN3FmHd7xIXN6Wal6JHzeECFkcFN9jZZIrckKDEcoCOqaPGshGUha+WX
09tWftoTFg2BdHaQhgHEgU8P7NK/a1ExnYMVBIVvAydjqP5sBP9D8CTLxK5b6Tgm
PZfZ5ELc7VAmu76ZLNPYzGG9iUQ2UkkEh52uGPJS95cJjJr0ykPfgAVqYfPE7rAs
i8Nl83uSwzGqCPD+VADiJN7dnNdvPcA3ZKLRb8kvosBsB36S+VlqoNjqIJDsj1tt
gXyBVBo97uFon1Ey82QrcMe6eTu8gaA3U1w1CgndWw0ODWs2RHcCgjQiX6VPGg6O
6U5dJ1ECazo2z8nrvF114+xqyBhsL7Tu72JKHcZjxgRlw4QJy3pb05A7q3DGnLIK
qMO7+GlHte+Bj67eexgnVCs5G4W+QbYDAMfu/I/tgCJ8CpyBK3ziwibDbvjqo8gu
hVn0iavj7olpunGNZIK72/9nxienWmLIhSc4LDpE7yRPoK6o33i/ob6cVZnUuRev
kYsL1kiow3OipeH8SpTMOOcJYmLCr/fLFsjTjGB3CyYYSDFeTBQAeAcUkkbp/ujb
MB1AuhjiJ3SmoiaffRaXZOPf4dAfrdu4LVRq0X5iBjb4HHBAJmyiJq3T4yvQzfpS
P+fBYarJ2DKNr2dvP8FskkIqhxWWnMQn68TYRj58U5naTWsiA847cK8dXqmOv3hM
HITal+bRh2pzI5twFDlrW2VuPnuXGRnRT7nkus0PZRwOEKlXuBEOGPhIF7vKON+t
2u4DGTgkzHG5Tv7JowjP0xBkCOq9sYHJ+zsBEtKxmcoDYEFg0nEcd4+/0OZ9lL6s
yKKQWVHFvEv54ZORzG35z/8NPxgeIWTXD7d8YF1vtuHkcNPbfnxL7/rDVULzSGxX
st9UIcjz4GG6JkQIH1XUddCCByOOvXJOLtxmnmmQYHTmWFvCaMV6GVAUQo2NEXwo
Hg6Y/rO19VvIFbZGHhNoaoPLANLEnzY4LtaEVCoASLmQYomizCXt+BVkBauk3rct
PrBmvMqQ2QBb91MFLd8hpM1fmu3TFCNzqen2Z1jtFHWm6W1ViI0dmAvG+ApKwigf
GLzKGDxHsRkrkzocb56HsU5lLE/F56iwAtVa4gGq/v6bUfQtMLuOnHsYVSe0M1Pc
X5pXtYIoKiLIcz4HoN8tmGG3t32zSFa6cm3UlzRmjnynoZIfmw9h6wLrD5EgdRZQ
j4dkF5+f3+s9XdgDvBC1o0KVZbEAPCpG2dzYNi3cY+4pEy+wBFXHYbIOuqo7jEnl
HhTSGTlNraR4bzIC7ZzsZM3tRujROU2TvtNg51vvV3XWUtUFcV5njgNKl3OwJt2E
gfG7cAtD9mhUeGmmyQMHoICnPItvJ6yUr9F7viyf4/YOa6RmbYCwsbfUW7FJ+ZSi
j2FjkQ2z53qrFMCNcN0hIBnToug/xJdOGODSm18/UCUgXVSk+NUzAZ4nPTC/qH7s
vU2jVr58PYZDFqWmvKLY/mw9JrDX8kuqFDWLB2xleFH51ZwklEbQ+4HEu8ThTBVJ
oHcYIeaqBt9t4KT9io1+mKqOt9zKXUBY6H2/Nh2MKwde9JdAmCsXKwZCbb0r2H1c
wxedKbmbU+aPJPSRruIrVVFEMMKq6QHe4oZ6gg39kP1CkYaopoQJyNnTEp9fM3P2
HaE92AjPMpDaD7Uh0Pz6yHLaUK3bl1Pa/IO/F/VsKujj7INKKX+MUaO3RZbceX9T
meU89shWeA7m8zf7zjUsgFXNO/OQi4OwTTeYU2jR428Fex5b3ERBMkxXj4oGp5Pt
N0SY+ihhSF08W1WPC5o3GE+U1H3dOZcmq+uO011hcFHBn7IQdmHocR6rtjYijrQB
DpRXqnxw/oVZWh8kAwjLG/I6TB3pUFts/geRAtXzsxijEJI8UpmsK96oKV6hbeZK
hOC8iS4AijIIZOc2ruhjKv9riZUAyBwtY7sYPVBX4Zn/KqlQe724M9V9RxTFVeRQ
OPDigGT0g3Y8BWyCsbrN9thzI7EjSWHZ7IqNSprMU20LbuiPC2eiMDtzQhP0xn/n
FH6eh0EF1cDvTdVKlw8grG2QBfDV43GgB9d2KoAb6JkYJS4ywahwLW6wyyhflCp6
0Cv2Z2oNkR+q3+BtxPAG3AjHN/Ngf2QItnu48WDHyKr2kemvgHLadJhwBCSfkKi5
1A7W5gzvLEG08sCcNMUD+SE/V19+N6dI1D/LT1OXvhVgOiakQOx3H0Lrfx6ClBj3
fQuNiquKseOE0RFvAWhb8hDV8XjvcqxumYOl77YLCvojnuUWLogNyeSTmPwI1Ovk
cMDrtl0Hc/+IZgMD7XE3v6h5QPjIdL+QgzYbVGT2R90wNcpGDxlLfxh2UbzHyj4p
zSawyKL8a658GAsqYJG0uR0EE30+G0awL8OnH+cVC5NVJrtQq117HnVgCLLgzcVQ
fCuq5P3lmfs/Ke4/SOV59Ag+ZmbpgsbXt0SzMEfejtg2bqbRNEdriaCyQXsmG2I+
0IlNvtZMVLoO2NQ01qfpfLozNBdH/imW3nVv4+pi2V7M/TXtf/+BSI+IpPkt0BxU
afV+m2vHDhwhWtRJXWvO5CKpYWopDoztC+2M49W4lTZyx3MU9xA72qFKnL3ya2IU
G+q9gdmYXCrQez2G9a8JdGHH7h73n61h8X+qj+2BBSFZBifGoP2rDSt+ydtf/GYV
bC6jZWChuqqYVstdIQd/exiz2KQsqU9xqbtwOCNwj4MJIagbJ7Kub3/estlYv/dt
kGvLW071msZlvr5pTDSbSgLiC9dyaaBsOn0sDIIvtzCzk13AxMkiFz+rLP3Wdozz
2JZNTELstxCZp5X9GxFdjivPhSK6rZJaIcuXjyYZBTXTGWMj6fM4XJ9KvpzyjW+r
ANUnB8Qgs57eg2Qo7gHagWyG0PSIrDZTzmqnq7mX+D4asD1kE4hH9qz6zanpMt83
BMWQW2dBTpIjSZVb3v1pinZGVXPbVVE2ikJYg2sH9WvpMra1lL0W7pB3PBHeza6f
7nilOnCVegh4ThfzGyLhIw8aPk6kNftZ/6+kkACDAypScFqfzEdTX+mxJLPLjVEa
9ZxbH26ldrkbCP7hNMNNJfuq6DWTfPDuYnogPrFCK6QsG4sWt883NdFLzJPgEWx3
BnHruh6SJZ5fkycGjN4CxrsfRddKYEIgEZfUrmZh9ZNNErrNk+Tnrsa4T4gfdb3u
6fzd5fLn1jSwvirb2L2VWX291Un+pZXGoGZFP7yKEvwZfrzEBYngQVNBa8PWPUTC
SBLOv6K8sPptVCt1SQtbPP9YYvbpynaz9cGkUpXIcO/aPblzqFCJZzlhSF6B0zfz
FqHrkidvRYVsyFtrOSndR8M7iMxF3BXBF3EcAbNE3BgWperDRiSYnAlFwJuz1dp/
LIbxqd7qi95Csv103oSRdvcRCeW/hx+15sKTkF75ugdTF8aVi8dolExsJkMvBNtJ
hwvQ//29BqF5VVvjAZy4+egmoEJXsKQHPjiKKCgdcVowGX9aeNt4dN/MOtQ/RWHp
4t5weIcfWN2cZsKOOdedIroPiZ/63/OGYt58Y+qzfcTBNWsowBJwExlad8kXkgp0
heUt0rWLiLUooDrT4bFtPOLLJ/J7vljRdQtfNgm65dvIDzYc6TwmKW6hy+iNQg45
mtM/PYdrf+L7XoNkRudMgh+z0Qw0TMXncbskOX+s20GZEMDnYoblPUs5bRWRZJTg
ahnZC7E3tpprJkow8IhPJr45Z3POrLCjxIJXz8lEHGmi0eC8wZy1qhboJxGK3Kt6
0KuOqg5bNWjyNEb7O8r9ud9zE/rgZuU6nfu5QES/BtqoQ1qM6Zb2BC4HT2YbEhE1
qeEyc6OpmJn4g74sSpxVl/mSsO0Mi2/PPcLpMECN8hE+ezp8SpbZ2govY8z6ABjK
txXixvsHwnqr0Ul1fQsm7a3KgYxfUPa//AJv6W0zsMQRHsu6ejBawrFivR4S25C3
GNkNRLJWdVOLMKPn6iZWEdFUDoq/62RDZhdYcgpz6HdRZPuX5l92ddbqMSRfvU0J
me/Z6rBlx0uHzf9PldnNv7d5GEqYhNgD7XlmOm7Wv+A0sYoiS+WsYs3SuW0R8/Gv
NgiL89lBNcL/XIkKdn9jKvI/VNajxSpB4Dnw8vbUa+rhat49/XUS/ZGwfhQTDERc
fwbeHwn/Dll0u/qqCvFrMepgb1iWPc5o5a726fLBvilCZ7r/Y1mArxERx7DOYNf2
cM/IPOgOSRmUBDXAXA7TpVE+TnKfFNJf1XRloGA4NVjIfus2K2Q+XgJTWjKWYopd
Ze1X8/Hk9MSIWXxZW88L4aYapnYYGKzShGV5zHW0GYKMRTkTW9G9tQfI+PtCm4FD
n8MHiNICDwokdpbGg8SDf/4vO85hjMs0uesdllYgdH/OuPj0YZWs5Asq3UZNGiFo
nAkI/WWhNybafgJ4rbkqnSkJ8uCPVuH2u/uGXRyOUlvF1iuXii3vNd2MHgR2/2v8
HbJpaSr8K0zETtnTHjS7/6kpX1XerpU+jcTt5V5Bq9gGK0SDTcTkgqRbmCTI6YgK
8Smd4uDioGdqbg/LOyzOBWKyYyAXfoWN/uy6vXVQ87I8/Jer1Ve6V17nRxPfx7PN
LOIUnwjQa2ccbGn7Qk3Td4oHrh9nr8kgbz/JGXLE+enDu8xTFZHYTrFCBX+eUcO/
0yiJiAQR+E+izXWebiENpEa32F1EmrhFdYrCd9iHdV2XULs7dbLF8s/4+XtTcq/z
zO4TAUh9xWQtMhloRaZW6lCd/K2wTMMbkWkGF3GdEOQWfDdVRbk6aZYd+QxWdeUf
SzYpm4lzLFcBnY/soBmbhulLvMh6IwjGy7u9SqZXyTzOUI5B6sL8lwe8Mx0CwIAx
z5B4FUZOHu0xab5URchWWmc2W/Bazt6v9mPXi/2r+EiiRmw3bKYGrZd1bHCZkuvQ
98SDngfBeaxjKNraqfZ6cTp3S9CE+56fy22psFjF3i82tyrY1e8dwQHJo/1DxfQa
/miCH3VPcn905XszaqH57ERx8HXbVKjMMdONA2E7ea644+juN2CwZ2wiVeh3KuQe
7diZlwjXlBJmQdRm29tsodwgN/6SKTdxEqGaP9jJOHMrfwjZa0IlpEJ7tpE1px7e
LyiQrWW6fz640DHOhBWFiPtwtU9RjqT6PbTwl5RtNovAJISSj1JACKctu99Ruw5b
TqXYg+4EwqBA8Qm/ce5kXWdhY/1FCN7ebFAIT+yIY6pCmUyowzEK86Y6qZmQWZbC
dpOZrUYAUlUi6GLswlGK5krBg7Xyt/gdrZdio2Yinb3cAllknKvb7mD4gbxtJo1E
J2aKVsO6mFJcAmk5CG8XhuZf76QLIMcJuwRJIf0sfxpPIPEZ0O6kVS6W3hvskp+k
m1KWpT8kSLgDG12At162JxFnq/KTPgYd7Nafk7bPcwtsv5C3EEiobyPlHPXHsGYd
LAvPon7lXYqDnwZYC7fdtnZVXTpG7BuSajV2y0NrxejLocseaTCXBGWDWHoqSaN8
x+nqJQJlK4mNDpwPuJ8OjIAS/5840rmkl8H8zl5NchNckeJM/rDiOMSJDXawgBwI
eK2czwMe5NoPKuWrhuexi8WxlCjsa/9XR9Lpd/Nmy1diMqDMDObv5nWTVqw69TLO
fPSpjrchh2Ee3GghzOpOn9X9IOi8r4QI6JBXMMwJNk8l7ThkE8rXCccBn2De/6LQ
Y2HOHkuSNTsn8GzYCCI+S5t8iekxn7HBemsnmumt5CDiplyh7ayUtYDunwlj0G/a
HVDd66oYRWf4qSHTwWjZZ9ZhKaLT4ToTZKwyM7T9OuZfxVz0QBPEgd6VBS7Dz7O4
Y1ac1qUEOHkX1Pq9ChZP4aQFFqGjAJ+/U7XweTjGt7NKHCx8+HfKrkr8I6Nrc8X1
qgZAp9N0iij9PLGhm0QtVclLCwSe4S/gvlbqLGneNf7fYER6rxP1074+pCRfsoVT
zOgAbHTl8PZ525Tr1nbNuQOjPOOgO3hKQpO+eLIM0+c3BMcQHPbnhk7dtSkVV3za
LMQoiRlmv30DrXMAs8oKEYqZkOcgfQ4FRg7q+3yBZdgoJGOxRRKuvCZiLjOMzZ6c
UvsA476TIP3gyzSmwdvzDhpz8uS8YgH2FtDE09Au34o6tEWLJU6ukjeb7R/gzI+M
WiTW8aVODlQP4+u95f6nuIZVbTQVUpA7jinif1lBIPw7L5Ae5Mw7znHA2G4gsG6J
q9YWlCoWD1mqCWwx48c8jlavVZmubknPNFdbAgljQukyV+5VPc8LFcnwOM6E776D
lyJE/N7q31vK3JrdcoP2kB6wN/mLzCoIB1Pft0CmsuZBpFFrg5meRVRTLCF6btEu
jBUiJqqY5fphTAbb8T4Mivh9vgo1qGiBcoK2SZxhbjmf5DEiTavAvKTMhjG9Pia5
3CDzswy/GzL/EopLJcQ2EeeKQKh5CEYy8BRfA5a2evIFhskLfy+UJdhy58na6Keq
80CfDIO4Z5Y1SejVMfvOBRXLGT42G8UtTdZApbuersDpPxs7mAtDjAdrtpOY+8Go
k5r7QEYxX7NbYWGkqjJixSzD1xhaowCjxs1Gvm5YAe8IxHntesCpSEmBTjyd2V+r
XhAYm+zjIDtxWa/Lsyg/fYtO+xUNAS+5Vwwa2mu4//9i58Wq23c0JdjErGXDGA/z
OOlr3XYNHLM1Nf874nu1YEfUXCqsxklgeSbvxPhC1W/Eeg2SWvPzVThZdklyXAJy
oP0as96ZthODvafNE78LVBRjH8tRyB9DLsSplFJKvwsIay1W3dxqmJUoZ3KybAnT
VoLhO3EjC7jhi/CZ4tOUDJOKdeImvNo/FOUqFUSUKZxDtP1ATx1cKH2G+jNZHpOF
EVgZeAhBoBoW9MFVvOXMnxs6NtEWyPsSo/KhgbFakvVtOgLMihQpoDLFsoXD8mw8
p6wtKfGkNXipI/BLPyfq+/TIfPK+c1irE4CyjW8xRicT3xO6SXG6kztEZM4Yohfq
++8U8MVHYmnKP/WGe7HeF+DXoEBOCQq/CzC1Rokpa7Vxxb6eC0A2MWmokx9I8BRM
3yWCpN3JF+2LLtHkS1jwwgjBsabxs9OO3v8nr2p2pmtsZl4SE871IrnzOLd16f4o
U/4tRB22EhMcRep4/L5YTsqkj2xyBqdm1KxKpXsr1oXHD1oBSiz6McY1PjV/7Khn
y8hLrrWJxfOi00zRw/auftdkQGEQkCIcyQ8/U2EkC+eyOeoXNO9B6Tx4cMc7JjmQ
5tiw2WoD78DhOXIBBkHSTMo4BtYAkOzLrLoXLTOw9Mz+AzOuh3eiAQ/ZB38Ypmdu
+B0s1T0Y5E4KDXD5YnuLuliZIVfdpswGnOqCkIO50UneXITET9o7dzj1sgvJl73p
0yHPgKpqvPccsy4uWfTbw/tkn+jKgRxEacQ3s1xcKMH5TCOL2J7roke9zjPfEghe
fhAa59HB8CnFU/pVNUi+4Nf2FYUpVNX+4qzrrDQoIcdlkizrGsMsOxA0xrREe1JG
Yh5Aixo/P0BP85HK8zHsuVMOAp7F9iIpIIOgFfvWbbhQlmQlrshHSlPHuJpPOXtt
RkYNeTjVpHAKqeRbN3Zgep/bCtmadcWIe2Bnd4RqHRCKsHDmqq9N1NKJZXHRcG0Z
f6V8Kq++/vJNlsCtPILqWeTO2L2T8dBdUWlohl6L9GCjWttyXhXaA9y4hwkYzuwA
kHdOgkt6lhQMKaUltwg5NMsBCWGpmyMEP7jFUCxZDDmvcKz/NmKC7iOXXUIIH5hu
51Yp51jrwckdfCWa8lWIgCN2maBd2ZwgGv4PFspXRcUr4vt9itR/lGt4v2zgwy85
TQ3X8h7hWBi4ucPZ1Y9w1lbyenPPdHRj6DE8qzAw2LDo4RH5N+b58HUpdbx1eN2V
ib6eLKVRtkXws63yCPi+LOwzgjLFjAtleP2EI6U9tC3T90HuEkpaqmny4ASZ37h5
QVpMOxTEYbPiYh6wjSkI0eJBJyb2OxZ6mMzK15FoRF3/Fx50NdnJC35rbhTLDO8W
+LFFYSV7zRBfuFHYKfKmT+TMrw8S8KvIS+Zda3mngOQ5cTtM6FvueJfEX1zccAQX
c33hlNirt4D1NH2ZRe/4b6Tr3ceDweZXyPLmq2Z318rQe8+G5/19o1LRqUO+fAxJ
DCwVdN1KIWsNy+COw1O+hozvIv0Oxm87g4x3/z0KE28ln9i/PMwnU7OaSL+bmV3c
kohmZ2AHteDU2LLu6hkcZUeAgmakCTjMTaWCz15CkAcXqwTEdM35MTVkhsrNM6/S
Fb/BPAb7Nvq0KJVirKdUktmGtMbsHvb3F6s6H3XupAAy5wTjq74mu+YNReL58EFg
aBkIVSHbpdrGkE13LVnQTAwPYpyuY1q3L0IlgPHN35PfW+q2xdFEK3ywHDZAGuAc
ps1VG1aWhaq2KZ+VWlmjLee1A6jMarbH6sP7iDuA2BW1F35tzwVX3cCNiFth8ngl
0Wj00+sFP5sJIjUxHzQd1PdUprRisyz7E2+juVJi9wd64AQhhqXDHbFH2Iw4lM24
2/hGBwXoFpDgeKRtzvMILmiHlGbX89LeCevYNYpxJYYIzPRTTE02Ymy4CuKCwsPT
LM1eDVlVG2CMuXXDkRQ+3b4ylG2eLlM/lCiy7Vw7eJ5St6mjbgHtY7rLcuJHkhES
TfnI0rNfnEEizcsJzW1lewzLhrpMq9xov9Wlp6ryxhIdDhdM+j23A5+cBBdfFxa6
bDYQw5KmrhyO3Ndbj7sIYhpKcvjnTF0Mch/lGzcBH4IRQ+sd6mhzCdXbr2fcd2dz
cSrHW2LK77W4t6fWNiaomcES8rjsJ4ruWAbRBHIQGPoEHIyBJPvWR60TGPFmyVzB
H2wCTAIG5W6ANZwyD6T6DlYsbgpoV7qM4CdfWKcvu3k0z8WyqIDfamtUJpFjRw+K
cvm+r0qLg4Y30Cf6TQYe8+PotIGfAIro5ZFHA3mtSX8JsIUEcEE2KKSKwrf3tcGJ
dfaatP0LGmn6tE4AU4QPsjSQuUI7DTrBZkxoQCn1mVr09PXGH3AdbHOUITLOplpy
z7pwbycoOqyyyGODe/9KGUh+AdXqItNFFZd1OMUt7rzFuGblIOYhVHFpG09vpSzG
nWvQ1EgISoe3VmpuN3xmwjnOtsL91x3u7M1SZRukd+P4sKuqDFM8O+FYIdgJrtj+
EJih2l60hP/E9JayxTSRQNVJYecfdLLkpkWEuEvEHghnURwVXHte+clNj2V5lKiM
DLtqEdM1VbPWnt5+FjFlL1IHOSQHByE6HaTBDcMd9k/tshzmkFMr4vyrp9cO0sbR
Y+G5m6GdcMZaMicDDWwp/Xsoqh+bW6IFfCdZE3pT5Zeh+qwJAdzDWUkZp97uB5t3
0RTDM7hSoBmvdKG5jcoXUiryt1ROm5zr853bgdHmYArqmGIeRqbofw/EQ2DitznV
Roum8Rrew4Q++8MuQKNEXPqkoyllPmB+u6/nHGLt1XtAixrLE2ew4f0GCfIcDtOf
q3BeIOoIEitoX5fYtclg/SrYOSyhFz71gumaM9WsaA1wt48XTGs8Kz+RVPrL92Ev
DjWsOjnuBrXmB/zceJs271GSex9ehmLXfW7vQ8tg5Tat4Jwc9IrmBXKiZxTQZbaR
P7+dgIoZl6aT/E4m9N0pbboAoYUpRMQKI6OhFgx5nPChUyvykdxULV7JBKRKt25b
ifPlg6VreCfEud93X9rcHADwowT3WHrw0HwFF0dchbhtcP27EmvCKH8yNxr+H+AE
bdnW5DKlxEtPIbz/lHEIPtYpSr3G2s3a6zsXp1IxHyKNqM1C2NbTJqsScdx9SNfg
LAKYARPQ6IOY/3Fq96npAGIni452qbMdtAHitnCnMz16a9zG09Dxaw/aIEUcuGLe
er9f5MFquSRkhQaUxV9DxTWBmuC9k+VwKeOJIyumcNgMn57YmZlQ9UI7w73mHjUr
tvAQmR2QolLh0A1dS6jM4hRgRsdH0NhvTsqywSAKwdPKi9rmDe+zygpfpY9PnS81
ESZi1vGGAK47ncqSanGybViOkRL/V2ZEkPHsInNRagmcdSWa3691ltKoIXnG3SB0
yGZ/wNX23RCD+6vqYJJ962M3KzPdWcM+1P3fgY/zTyXTqYRTrrdi4Nmq5KKso+ye
JdDhtDsjNyEOOpcQls3tRwB8RwCFasCI/M9cBOprNsSPZFpBKdcuLFNr5SA1ZH43
YK19FyOxRR7V0YYwfwpq/wVKCOOD1JeXwdTGJIUbNEDFlYjd3qvdIdo52Dd4Xz7L
3kA15wyaN6vf0AuM2DGg8c57shjk7hH7TgTSdCtiIa/mxZ4xbPjM00RqRF/tW1QB
e1tpRNTp417E/sTEoWH05awjAy+v+5U+u58+CsmGHGf5mBN8RMcmIcG0547bA3k0
vSUqDgsES57V9C4wXA2qqla6QE8XsAUgIIBUofdKV2pqwvxznbTLa7NSGyMKWuM4
jIGDRxbvC/1esNbFeoNqCmgkZmEbXyRUl+gsRehrE/kYUOKeEXJNNckmab4KKtLU
tLiIODlXCzAwEvIBBCPwSXFilU8q2x+FtQIJ/b/yKpdhYYflicYa3r/dsbyuBJKV
kVTd/3Dm+2vRSnnwKI0tedwUuj//FkErPeSasmttXjL0ZdKcBZL40Vilpax9jyER
ztwJTIwqaP06hZm+wC5WT/so6NhHt0PzItUfTXbTLSJtBWYUBoaY6sYi7JJKSqHF
2tPmzYCcKnMjXzilUuzAPlLv/a8hoLE5LNEVJpG/xYSFWLPZq8isQv+DJxkTnUWK
CYERya6e0jzmx1hEE8r7fXsL0StAEUJbzzuI8joJ0Q9GKf6xKp8I+7d6qf2vUjEU
iVr6S4ZuZ1/h7872OqOETowpTWugQP9o7ORIfAxvmQSl+6P8gOfqvuUo3tFFKYnY
Dn++UtI+wqoEhoZV1KuAsveMUxllFOZL8RGtUFvrcqOwHhENF0BiK/xNbrQq5Nle
y3xaRrarXIbioSuB7WosmgZFltbtGwFJdlABuJocwFgUc+1wlBepcdfJlvnBZCOV
jTLbx4PW3+mq+bp59I2VkH18VmIvv326abPJBvLNxiVujDFSZY9F7568zB5NUrm6
kmLLE+oU8TbsDNGrcz9aXWX36QgHRlZZwhIOwXe3S+h18s1vGXfseJyMMdL1xyh0
rSMfLffZsD9HhpRTUpCg0flpuWaAgSrjabrc/YTLCkA4CY5ngwlBAX+s5VTp2y1o
+F0Q9ZJ/ZK3XmWCbwy00yNBHxEV0LihmFayytNlbtVl0W+Gd3XRlZsQJJdZuTmhS
n9qLxMu8DbRbhv9GWRtjgmSObDGWtkujpN2A5W5iJy2K6Jy0WJq9HueqNv4rgZm6
7734ssAMrp23/2Zg58Ki1awyFlTEsTdaJZmE5aLNgIdSUH5/ffmH3+wUv8yGIMJE
LT13tmM9vaLDcuEDVA/Ww51Z5Y9driuJwfEj5aD1l+uom3uU56wGX4UAasz/0b6J
bOz96cY5Vp+y+I/QDmJY/IoQ/b04n/a/DftLCwmdv0IWhRYrh6psTUQquryupfnY
0C3/HmxIie6vd+ZbnrVGb71GAP2mrEcFkdtSON9lmaMSX7xXcicRxMyfNfI2EMT7
cP1B6ljJ80A686Gx62pvy3z/3hWTYg6XZ5dSP2NaSd06OOnzOYkOSx5LEpsUTRUr
J8d2i2a08E2bapkLJlC4aE6RwoHHRvmYYVaYhberPUQR9oAlV2mVqk/HBIpWHpr1
AHLtDayocw9ESlRGoVPf9SNaAG8LNvL6mn4aHLXMDc0FPf4fKbdMuTv9KwmnrpXn
KVstiKLnZKm/4tdF0nMjT1BF5zD+uFMUs2iRBRYk2ACR8pmNujG2sD9OiP9ts0Wq
O8pNg6YMRiMuSYdYWc99muRZwrxk3/YQtVMPJB57HM+2s92b+sEW714lGehPL3WU
QsDu2yEmoRCCg4vqWdaVvn8HMZQIDsmwVHNC7CSEmtZ/gecpjNJBygLAKEIgdl+T
0iRjHPcrcCsyuPV4+ZBBtpHS4F9hfNFYC/0wp9/6N+8eQ/NMUo6WxXfAwS8DtILw
GgC/+o3iUWR33TBIZGZ/RooKKCgtA41jBvfxKBwnANrxRkQ+2O8Wmq3W+BSwvwTL
L+jIdqbxoA4Q2BkQv09szwaz7Y6DD6aQhhOc+tqWZn0eOEz2vWJ7EbQopS2eJCU9
BE+TRnvR7aPZvSu5UzbV9XJ0FwRutYaB2rd+TfQTBxJdihOpeedQp25Rr6Tksm0N
oafEvP8a9ze7vyGTnI8c/HlyqLmQB06NFqIroxEwiJ8rgHc5QvV9OOb8yHxglKAd
rAUWedUd1gM95I2y5f+pouPXMnyHXeNpMcnTcGZSmd37FYF4ejqtVbTTOfKB4aRz
oMmhqZU7sWmtxAEK+zF5uaBra4LO9d5jeG8XVx+ulAlzreaqh21VSL0NM6Z1YGFB
cF7Tv9pj69ZZ4HBLPCpf15qDGq2txWwFQgAbDRh1H+ZzeARDC/Ss+EavFUEWqGXm
+tZ1RVDP5SRuL2p7ETN0LyO0CzkJcz7nq4+6fGzfrZQYZBhYUUIaKtMjIZuwG4VZ
bJmLCAJ4+esIGOG5JrFrKGw6245LPtLKSn0sIn8jx9SchLLZ9Rqvy25UZrttPZ0p
pW5ZJGisqbwsRwUqeTz7AAHtt7k7PbzTKVWXfCID6qdkOgGtX3Y72MRfRwu4OBjC
doGCG+aLLWyZZgy+E9h/1CoH9Du/kUmCcUwYRAOb0EnIw2fxbHHPddmy7QFTcS5R
dwVH+3ONTQe5SZv1Zbz5/idL8jM3VlNRBO/7TmbRQibKn1tEb8mrsQmcZraVxhk7
XS8Gd12w0pVWcl4++oFxPlvAA+a/7dzfZ/rYrhG8KtB4CnbSO3v56yICi6QqT05W
16XZr0gVm63v7tx+AncycbwstC9A/78+MZcXwOypY2TLiSnRAxkd/Cf7GVLDHngb
WmOQ1piAG+wc5xRa81qIPFUHBLDf2iGEpAYIZxha+6DaFoRTdaseMZg9OOEICCQk
nGkEcWxJ4BREDqRyChBDE2jaXT/N98n8isH0DI95DSqUOY+OTAUxmIWfXtatwpZ5
RupDfp2qz1nvHTx1QpgyRWivX7rR7AqE86k1kM9sOspmK6u6y4aoLUp6h8jcF/kw
MxD4ICxm2jTmFqhpuntGBjl6r4RLunXWcqSaIeh7HYBdIjdWXZyiLxJUseF6vyUl
O26O0mjb0D7O3N6BqXH+zi4Sf6xfl0cfOUiWOD45xvU1CfNsSlvDn3dBamuV0sjS
Nu5yU+vXDZzFAgJR1C2sNtonTH7nzjei66xcnsr34PGzUI8mUcyuPmI2kWSneArR
ErKrE2nAqDG+clh3wdAG7cNiPc4nJqtcNVxtW2/xTLXWiIt7LSRCCSMD7fObXuFT
c4mFXC6qRjYG4Dhn4zGgRXKyMySW72QqOrSAfz4PQEP5LuFuhMF/k5OZvFKdoWcw
/hmK13Wb5Qf1V7ZY/Vk8Evd6u1YpwDV5KzIxWCPplA3bwIvtEKqcycqIEbeMuRYq
CHB468K41ndLKAOm8C0kknohM1kr5T09tjDQ1mECFGmVcHofbHu5FB1t4OCU6hKW
NmRaS7oH6TBzY6Tp1lSFKTvdfxOihAkN/J3M6GssTwr9XfGhe8MEAV4z2YGDv0C4
l3gqxEBWiEClW624ghWGLbHU5GNPq8db13FERczepK6r7MkVEbDP8gwFz9HwJ774
0bbW3OTRXbRvrFsUI7MedgUBIaeS6auskqREk6kpz3X77hGTIjdansked/MrSvdJ
KZWMZ4pH/rI8d813wtG5nZWnzA3NtmtXwcY4Ga5f6Z4gq9fqpS3Zl5Fg4OaLCg5N
YZXws0mxif2eYnxHvPb8EXOKUFgKPzR/c060iSO7e1EnA3+uySJ2p1514GvpHJmQ
XQXk+44G1p2RqkBQlwQAHWZ31Q11wJxBmrlKaRAtVYnAo7W/GAxIasiZYy/ux7WK
aPdS2og0kw8LDLQR/54pPldyLbwTtdun0c8al71WRM02gbRra++KUgdytFAAiJ1K
jHR971tFXUYYbKtaPI+5NQ4gp68xoDlXgSIwigSwNV0KTvJ1Gj9dmfarJdUf2Rcv
ElLp82Pl34b8di/HYIHHjJ6RQe0qLLCXttEJGke7VDNWDej/8SvWY+OX/GM5fZsc
8vZUj5vCDQwXtngKReK0JeCBsaBnDGewpDHWQqcYrLc2TWSI/5sigZjmHYNVeEhH
hR1hPHa09cmBlRLbmwHpdvXBqeNW5pWfVP+HPh7zSz4jzVcwrUd3a0rNLGiqoVII
N8mixiCHXKTjD6aU3w1kYIi6A0vxT00yqz5Z3C4ZjmHAnsqk+9U6QWa4buloFiz7
XvOoc9lLuhI8KTm8V6snJrK2XQmenPvN4rpXfmIvbmIeY1mZs1UNkyeg4FWbRTq/
qlg0zt+SKhdH3eQSjbP0I7HgZoLADDRW/0Qfz/D7xNcdcXVpe67axdXfn8vbxAfd
HerHqctxOIMRHqrHcRdv5sjFlGGgLmHLEObArxQRc62a5xMd+wzViPCQOGRBSxYu
Gd6QHJAV3qgPb4IqKZ3a21p0Pke/ysVoSy4uSFRf4Mp4mR19DJCcjqZFKcQ7DQGz
x0p/ZzM/Bdma/C1xJ6726N9ekLt4W266tFF2Rt7LmfnaIMmpFj9hhyXcstF+rseb
Ao1qQvwuzjW2UDJWE2pOYvsn40IJKRLkKvMwwviRUdQ+Ii58iMS8/5+gXEoGO5qv
hn79LnYuyPPRLXZ8rBhu9cOm3Ttb5lGEKmEJ+G1sMnHsuQTbIJHZP19mPcmkFG39
NMzhBSrgH1JisxSesnZGlvRV4vUjj4EqpuHMkonSlKD+G5dAgV63bQbN8nhiCU04
1Guc8jJLX9yKTAXJum/YnufYDORSd+4CvAzfJBZG8DTOLS8OjX7LWENglAuKyD+K
zjrDRIOmiWTzdFpB9j5aG4bVXhcZg5b1sx0cXOjjXAyyKlC/ewFqhowN9rSmPpfd
WpVQ7KWYsdMRpvSBPJaCTA2WZfJ4GmsnT91PRMd970yeb3NqPqOhrQSL+vkjW8rg
nohYBR5RtNYTu5M8L8zeIZBfDuTrzJ3jI1FkUEpnHYLrlndNc3xyYMArouE9VkCn
wMoc6EJ682ivSGco5CQhfUlYwymvYhg7ilv6sQqkIYVbMQkavKCPgGotqZ6SYi66
3BuX2mAdpsLpseS6hD+fb4M6oGKmw5U5sjzsxqAvbuokN6DkR5cVI0XS0r56IBcy
4m9SiCNVkRosOyEvXffvqdDba6WXhqWRE5PY+i+S0uztkN+RjYG1/qTZUNqql6e9
815sI3fYZiBRXUIc06ydjIdDCIMYe4JkgC+57xA0eRQ9lAQcbwHDYRRSWv/G6Toc
VFvC6spPpWLOLk7xR6JKWnkW43Qz/bA0cgeVye6Crxzy2SuIqPDZGeHmCsCuWq0w
fr5hnJM7daAaxjmyqyH+0c5CNCkvq6gjpih6boJ+m/YkSEeui1Eecyh/jq4uMihw
sHSquVBRAylwv0VYwrp71d06BqxdVTbw9kLpUZqSn2B+B0czeBXhTmgkQwBk9OBF
WvoNoBU2yW8AFZ7Sg30/rroSFWGfWPjkYjCEPGliBA+D9bowvu4UpCnJEkxOC2NP
lkr3Ksu0kRRO+OMqRYMKOznwBbxvZMuqXNW1kpdA5tR05TyuBvWYIUARLJ9I5csI
GpOZjOTEVc/U5JQ4ySHD/Rqj+h0BQJ0Y08or8Du3/TbSWPFPoSYngBhxsTgGI5kH
wj/dNz7dBOeUuCyZRvn4gOyjVtQU9BMGjPryzdElsMX+bt7HL/JadRFhmErHVDqV
iiAlYKAlPsco48wn/NrcWRQTCEWQJLdLPQNhlKGbkeSd9hNBclycOV81F6kemESg
a7HDeEUHhZOvJUpl6iuZeIbRmsYHi30V6ajM/m7LNwtCWHlcHOrOJKI6bU9Fcfef
LhrRZxpw1kyKnF2nfUvlPoLSY2eeXMY3x6/46M9TAWhnIYNe0NkTnJ94tMg/D+M+
jYK0AZifvcmGjl6pA1X5+j0eDfNOGuf39r3RJH3v3KC3qqZmQvkwXfaSLEp4Ok2r
s8ZR4Ag4vNztgWkEqoHutQWfBUPiOZdIwed/KX+G545C1+SyiVnlwruGgXVvyoDR
b2zLza0fi2LkyucV9+4Oh1VShBr/Qrflbi6VbI7SWJppNYYGXUleD6/9SB/i257H
8bC/tUiWRxQ/TQ+7Oue0Xb/5KRTLVTeRWg3L8A4IHwuV+aGuNA/meNr3hWSDX86/
GkrkxAEVxhTmpCG20DVic1jS3vYI3JehSolKoWejObF925VegMkFVDvYSe1mjy1+
nzpm3vzjFBm9qpkqJC2X2TWtj/it3Fkd5TEMU3kQQBAU3JMeLr5q9xghp1IbaZqB
WAyzIpJ9ifzrDs5PRvFw3tyZN2FuhYt51L+WRg1yrmO47bRvBYjFBEb21bEfx4cD
GZ6/ltpWEvZbhi030c/Kl7WqxkZCmiNfmtbLjoalOxI/OovtOwBCm8A52sE+1ZZI
sdsqNQrDn4vIBFacOy29vaSlgyZ5Im5NCdj7yxe0PRgAqAoEbU4tUXdFVikrMuW4
282BO0IW1SF8Vttw+gIZIdvGd/2UmfCacxpAxdU51ZgA8Z+0M5QKYp9XJYE4eQhm
ohdRTuRVoMYoSjSp6bivFqkMJFJKKTL5+IYZ/6e0q8OYwMEbVRo7FdrpzrbfRYDV
KJGWWdqEP8MKXB8q0l/L5PqNwrdJlJ+LjbHsofJ0xgP67e15+wWOMa1Shv6me2dv
CBA7AoWRrBtXw11VRjU41jgRaMxD2OAnlXJLrFobKsMa0TPTOgERveTujt908Q6J
+oM3ENQSez5BtGCoyd/0ApSvJXbxYE2X03m91Qi/4P5cS4IFj0vt3r3hV/DbWukL
UahMN1yloPAXNtpaJsHU55gF5R0qT4XJtbRklKoOu77KAvYTvrP/uCKUbJkgziKa
bbx9AQG1j95RqiDzEayPiKUNgU6rYgmHOcOOLIgg5zygckIMunEGcsG095WQ1ha7
9lfy/wMZ4j9QUJqSE0P0ct5A5q62Y7+WpZ/FmnULar0cED5LX8m2gljaybH+ufih
7KcQY+Hqa9E3nJJsHqtJsBhsdyePodb0drIA0skNbktHaXgdnwTfTeduzDHQNrGz
ZbCEKgqjZkWiW1T1fABbS0EwLd4w1hYAJJ+JD1OPvFB040HwEv87y5j17JcRFNGK
KGDbAqp5sytFT5150aSZKGgjd4iRV6j3IEz5+BQcDUgsxlsvJsCXQU4J1BLLxH2W
RvtuVTQF63Ca87UU4nHvYM/ydS55sYetwP2Jv37+AMyTafRSzQtVQdUvLDJSe51q
p8JcXhysqRJPGgU9zdlGSIDMA4WI7rHac4JZ9NhaeHg2momziaUatr2RoWu0C0UF
0srI62DVHECFV1fKoZejjTRuGjfaoqhKLkhrT87odFViaZ/QwoOJJXGzaIhKl8tq
ongTDLBfIP4ilNqA5DC/iErFP6ZQ3fk/RD7kSnbZLSZYvBH/fmQBVTowFFoUs/X7
DiqgLzxFN+B8i2jzZSmKH34NFyPswD1AEPhaf7NzRsUTjmv8m0tavW1y3xTOyx+e
zX/86hK8hLy+nv9fSzZZQTQ6ZH6Fexts7fGXVxscBx90FyM5P/KUO9RHA8r1N1Uc
WppMOEUPm11gaF7Grp/5JS7eYwGnuMEA6I9AhxG18QAS5ken30xu66z/i5eLfBUC
gb3u7JAH5Vm3J8vQkORb9tQxQ1uYrf8bm2ggDzKQyafHfD0BVvXU7wfQ67yDpIKq
HFWXe4/s85zLcZ12uGKS5czvijtdaqI3UTS2RBO2OywxJw3mwzcW39fK60rursEL
U2IEp0mIyv0fD9/IvmNv9TuE1NYkNGZvwFBv4qYkwsrVUByTTmg1UaIA15rAtccQ
VvTNOVi3cDMnxO+j8w6BWeSFhU7A0ivPyG9NRb1v8wG1ESllEJgZov6Bqh3OetFb
aHSjoVulXj/qE8aK6n7KzFsALmZ8s25AHbFbh+pzgsu4vb2lZ2EHIsON+kdy3/iF
srHoVJcmZXv4SigNJYLRJ8dy7G0bT3hj2gY1y73B9nSYNt40LJQ/lY/TS7URItzp
S/c56qr7u/+BfUH95jk4b5rHAVzsQtAuDEJqEvrH5aYTvin/yEPJziFtX7+25WaC
2LAVkjKgn7MWgg3rsvbWzdYuus1ZfvUi7i3kc/NWaxxN1uie9xMZL3Jeto8LUFkH
YbZMuGhiaCVKeAGGc2g5gkyriZMa8yvMyhw5D4D4RnAl92Zb9Vu/PGX1j94qn3wL
RIqNmlnTYmFxM78E44qbAgD/Y6SBjEAKAORU3NNrPkjvBBE7aLswl1APxNvycBaL
U0ygvYd3gd2OrICBg1eY218Wnr9FKOlwr2XqSX6I0qbEFVun2PQQcEWcXybxl0WD
IlzaOpvK0YtZ1S3em/og1v99hLihqiQtv7TNqxHxo8AcMjKwRtSw45JZHhT6d0ki
vgqYYFm9+tmbKXJskwcz6Q2C00PXlNip7leZNCrhyTDllsZTwv+eWWE5W10oXVK1
F/2Iz+qHSsr8SobvQVd5jpbsDNJ700L4HrV0ClWxw6Kg4AQGutp7u3Ec3raD41dm
vQtiaWjTb8xBgO8+LtUkdSugZdF16gCMJzGosAf5tE0NGME9vfvtGhamYRC9Rp2L
KQG0WS7uKGCJ72m7fElyk8Hn2XFoMfvllSAuKjtvJgpRNSZ8oeaW7OxP4A1GwQMX
dYwOj86yDyBZMpkoE3jAVSzp22Y/qQnW1GqeVFDaz1uUhSWCR1XcV3+1P0X5ENTw
5j6mc9bpQ5S9nvh0OSVB4/cbIP29oQrDk04UgpPRTymBknLd5IyPgamUg17m8C3W
a0PAjlrt3f6A6sp+8pW2ueArh/DElqQWJReC5Tbtg5q1JkrYV7dyQLYJ8bkobMHC
VOntSb5CY8OGI+HSJ3cMpWxP76bry//md28HrEo1AFyYMHbhfIc9pyOOgkbfhUVJ
3VvvtZg8iPfWEBRB3N6ShKz0IVnCyKgHsIPnFg8p7gnLsfYDty34sl93TzxCZNAq
5Chv4rH22T59WME4tejbnGG+QUpETBHdBJ4UwGkK/XwqyLobgppRightg/QslB7K
+DLMV0WEsiefj0ZxuE/Xgfnx7PCgN0wSfLvm4zV5+1uOQF3Zu2566qSPjDZyKgK8
sELj3gQB/zZWUWnH96os7WX34oiBKn4yyrGNv4TftLciCke/Y1aNo22yJqPeW0dV
lt1pwGGYqKiWOGvQAn6rcLWYCLsJhkIy9QsCvUOWlm3ff3l5jhOQ8wKncp5XIpmE
OuX5eH9msIvEuTRyz/1zEqeshqjWBcOhgZcqb1DrFGBrBuxYerCuDkswPxzfcxpT
MKEKooPL3uHU7tpddws5rnmW3J3iMoFueIZo04OzNtLkinO8wNKu3dhITH4/P9m0
lbiY+lg/h0DzfMdMsV+JWx42/CQm3GjKtHtV0yQze/2k2qB/0qg/giFOu42FkPpE
4OisYfIUzFM2F+18jihtCgOY/d9ZSqHc1rAlhaOHXFXDTVomihfD5trWkn8SjZGi
R+rWVFAgfxoEcNm2ZBmT1CztDKI1GYQ66OdfqBEGSnhK+08BwJ1CfWrk62tob+pt
7V19EEL+WlFp2AXHdAS12igxGhmbDyc0SrVnaMDJ1arFgJwJTdFVEvufRQ7GGhz/
TCLJkHUuyPk/dk9Nt803GqREnubJoKya1wxXcQnprNh18eb56Z4bY4SZ5CMb+C0z
lObhrFNdaNJ02XxQFRRUF6izH47AdfhCpQMEWa+zkMqx6ycgUkeHIO6Ky/NuY0sf
B+qm01FvGg7HDANhrWwBqugUIb9Sm7hQvmI0aGBVn1lTGelTlAUei6h0QUhma/Mk
BcmR56mJtY7l1KAiuVg9FID9AcD7mgMrUJgXxrVWF2jrlttXLLPfHnHt+X7r5IDe
9U9qRiWbuj8l3iN6HRWS5AkwQcWDQ42CCf919r0hxcTqxfX0q2tQWDvCCFIsVgeu
ujvAduqj6WWihThVjSoGen5xRzN2FDTg4m7/f2otOnwZGXtzmydCOOvZsfbKxS+r
JiA1juHUuh6c1dmDFHXSL0Aj+YtRcveD043YYxzsfZbVZXWEGHNiQN25P+GLN93o
J2PmVd6XMr5q1lE8gGtCYPHSn+HkScamHiNi/tJ1N2mkyaJjLLH25qAxUcGTGVef
F9/I8LeGOlYJdVBMLseKZYBkZQsESCsvbkCTG4DQzNUuBbbTpsqo5KLvQ4S0kwVJ
5a2vsADli4KAfxI+0uEYMhmuFRt8GMEfUnF9BjNjR/CfYMTcwb9AT40rWicaP/ZF
zuN+8q/2Me3A79fDCAbKlCZmY+aowDD2ADs/9OUJdZCUI7nXVioRdVlLverN6eeP
54iNvgMOngdRJdrt16wZ54IkEYoUT2u41ZJOsPTARzyyLSzQoaAT2YSKjrAShJrf
zRYvjpSXFg5sJwS4WCQIKor/QkTFLh2xtJcmPko6kyA45nNAEpwcfwDd5Ygv43Y8
jo+6dSZGYKADkcT2mQrYa2p3Rdf61uzeClig0zteLoM4sy2W0LLLee0obO66Abhk
32uFxjytPC+DZq6JEMzLDkqY69yB0333FAxytD/fcCzcyj6ZBQamOpBBwJrtTWZo
hGi5z72+JdUwWhuCnIULgM7yVe4vRuKaRw1bb5rzfzav2BrPlT9yuVibhriic30c
QUttbijLQuD4PLm2RKZo1xc+YT5UP2F/WBpIcYhXf5/VlfGIulw2oqH9teDbsmFR
ARnWpaRzbUWQpd5RMULru9bR71SqotMCEPD2YiI/gfxwq0Xa92YAqcKXNg3FHVp9
t8Nwqeg+YuyrlnZzS3yH2DThD/1GhAYqVWdYGfnuj92lpWEritrnFoGNufpETOke
y+4CXjrfvH/Gr8a+Eii6l+o9JJCV0a9nLjoSaA0GfTVcDTiQFlQ84IyguL2AObJI
QcNOB6y2QD5/l8rOyRmZGE1SmmV5Vwko29U6P3tkPf6mANEyKTRtltX6sIA+FWvi
HfDqLfE+JDO8H9U6DboldoTo04pZuhkvXeXXZ2PgJM1m2WSkORLU084AT3psWN2Q
75KIP8TPONKd6mydve3oCmtxi7sJseb4GyRLz/P/S8VWC65HdY8LqfO7vI1xnrTC
mEkr4++RdQEA6Xq5jPgrNpSu1asr2J11vWRWT4cJzq8FHSslut3bO4RDiIswQD2c
UPHubO3XgFIFXtKYdcWKwt/ekDGqSZP/DL3HnMX5Svgxs5oUr4KgZy7eNj4u/ADP
455l6UPwWOiVjPauqdA4qNCMhRkoUHoXsUjCQmpdhPxZtBy2zOT9BVOdLEYwCFLM
HBQ00C6HaI0//maD1U4AGdoR5OFhoVlLjT6i6elQVW7KAYsinsc9K2pFdBeuHDwc
6Wv6JbHwKiEEf7l2M2eK/ov2K+BW3BXcUZnvPIpnJZOutf366UiKxYMbdRqDmCd4
W8MLwMxbWVpiye/SLKFLZw/Qv3OCLoJp6j26DNW0PyRLsoFB5O2+VF+rcZllDPDq
XEdrF1g3XVEngUUUMubRbaNLC7wxHfdoiP4+QpnkBql9+lxPN3YN7qiLuuPEG3v6
Q1O4cs2a3MWV837iDam9BsGSqFl6cEUtZdEop7wHpmSu7cyq7hLnKECxzKtqDHtG
fE6kWbtxO9mP4/5878DBEgT3BY2l2H5zqtpC4XbdGHd+T4UBVIeQRHkJovvL/JiQ
FxUrGbSM5RTeaAszGstwl1anjb9l5dH5UwQ7HNuyjRIWvXjL4O0C2Xd2NEZgpXgH
2gajZ6erg/GZg6rWSPDkxUXgXEvEw2kW2ilUMi8f5CQM+mo0Cz32+QNA+ifgMkcm
Lnib/7hktfDdUL6cOm393WKzZm3TW09iE+ypTlQrVTrwSWGbn6bVyNHk3DHK6swj
9iWXGfCGCGfJBRqKjirOYIaU43Ox4eImGy8nrUAz6N40AsSEZhzeiugglwilzWpI
bIudtcE38FQhsKsSsJXWhRmrlceL4uI6a9lc6rLsZKKPJ397EufACXOPAz3vy7gg
5bIMRAKbxue8YaHZ1ESKAMdlS6ssQ6OY80VmrTQtCl1yd+wSCSQCx0kjoz59BXoT
VZledWeSNhtb2o9SYtf+8lwEL6JjhWQNWfTmDYys3vYk5vpZTHrHSteMKHE1zOK6
0tYZgQHTurnByvyqqoyii/5GcG9sR+OxMYP9C45HraZULSHUeZy3N35OqyDur35D
c96/buz09/ERo5tAEGHQx2E8eTRlCI7oRP1lXGuR14Mf3UAbK4IeOE3t6qKXCH4Y
+yPCwKhgpRLZ8l5D260LSZfpcvKCaox33nLMZfyiln5gO9650ULlcWLkIaHwN+Kd
IxA43RGNS39XCGDLM/zhLmXSbCnBykvr05ZbjV0V0p5rIZERsQi1AiaiN4PYKJAx
dAQuy2NeR986a/GdXBWe/AHuvfSQTgzC3FSLajJMO7EhGKHe7QSMu2v3zk3IZcDI
+HBa5a9llWUw9L2Pdl6/aS6QmdzaILVpKbYGsI/XKyErA5RNM/sARc6wkc6xPjcL
3MyxosaQMfCz4Yv730Y5/qDPfhP7GEFGxy1K45j/Gecg1+XWMPCx/FTOq8JcsKEB
zBXm5LUn/WptR0mmgEqCjJ9WJAuyqGjbvKSdiNu/QIhCHf3kcxVrkcDBmaSu5mKK
kVoQWXEOd+ppFjuIyhqUUAo9sy5OjXHmjeseS65WhVLQBESKy2zdQgDjfRpuKiBX
88DnYSTFhv9dM6nSo0tfMSO9s66C0rx4wbGb69fBdT2lRepH5ITJ31Muf45r+fGp
ExiAthY1O2iGjo1qYCXlzKueTjozt3MEbwAD3MSXMP7pL98ncpzRVBgiPeU0tWxH
+5wHHk+npp3rOUeQDhn/E8N3Urs9Wm07y29wTJucQzD5bRWbdWAxq3VFZb2/0q6j
cYS3+CdXL5wdi3EtZbToC3CRa93Qnk5CV2lfIgNtcLUBCMakWQ97LigxRGIGA+Dv
mwApu9QMrsOxs8yGaZTV7Xv0ElM7sfT3qDJk1PKpf0a5kQPKGejtWgjsyR+pFZJl
z0VTuwjEOCYiQ38ldhiX4KKttNgpnfYyTWryjtolrcyeVSMg0kaLVpiK5JchgaiZ
XUhFQ4IIh93wBkFyx86tLyR99pUShysafwxMY6O0yYZNMHztvWr7hczye6x1lCq3
KYcGcIhQ9NuyPOKL2br2gT5t33op/dzQLbX7rUi9UTkymu24J51ByYhslK33zPrA
x2CUmxSRftnq8JAKb1R433bCog/aAicf/M++jF8NZwjraPxEpxhQYmp5HU5fBZfd
JoP0RJvY1mnX6+KM07tOJxYaLZQVIPT0vinNCGmLBGRZyHAqxt4ZbiwtQbcV3O0x
knM6z5QvcaC1d9qS5HqvxCxaVjwuXdkLts7gUcSvcvY4fQGNhwU7w2SuYlGHavVE
FEJ+/ua8bAl6+DpxB20RNoZE1RsUc0zdhRKOqBGk/xsDmdSukyB5gqx9BKhAlU1K
vbiG9S+wbbU7xmcPZEfDaMw2607qzN9DzHzYGhBMZWzNgCMdpSR43NTcPe8fBtng
MW+OfyJ3TrRDQtisNArwdyVRwY6cO04rTIgTrNtTJYD8aG3uccd1bP+vbPkb0cKB
qJoadzo6nQioH420TBY7CIA/m4rf96jsrCXATg5aZBndvOeEwq8ew6dU2OkFvYmT
/39G5C9rwtQlrrA/f6B6yfKzfRajpUKptzuDCvD+m9VVtv9yZi8DGjIg5FD+OkDg
nlSaul0uFGUHLNuDnWbdEe294yUTJt9ahZVfjJZswLNzodhNYoG01fuWxQNEx7qz
BIjixCgTUTvH6dIpLD4wE0QGZPUwxAzAj3VyYj8ldCpSGF1VrkINWkFhF1q2abet
YYFVyk4p4vXuxP2m/gkk9QUlURKuvWmILa+0NLB0S0j8xvHhfmSAi34K/U9hDS7n
viUeE/beuh4+NeSlVg6ddyKroZa35uDBp6jVj+gdnYICSIQPkEzCQvC8mBaD8J2Z
mVgVxLAyMzJsTG3whrRSM26sL+x1IyKZx12GTTqNHxoZqZ6UVc/Uvib0iushxTAk
ke6CmIeGFGBivubzZ+UlICsO+6xubTHVJJO2LK89JS2SZSwPgIpO91fWdvqVkfsT
KHiGU7zB3Mz62u/lq93pf2aa2djfaA9pMZwJAbJ/MuAZa9fZivZg1TBV4l8oXIZX
E3AAdtM5XOivhcWZlV6cQldxFNHvIXMqXFP+2MsL8yD3WQGgNJncEGjrWglzLxmn
X3Ty4w7VVJEwdwT3O2+3BKHe+E9Xk2aGigS6oN2/oGFY54GhUVduz4ks9A7cyoP4
lHwR96k7OYILVesCK4a1Pe6Dv2xyohFklqNugs0CkwxAXR4uII2kjVtltVpiiLAU
f6jEuAHBNREBWsREab2QT6vQhnf+exTNOiO/OlQY3K+1LC9m1feHY+v9e19GllGu
Qso0NhRSoXWmx77CgT0urdTEdnxHqBWpHfLQvNp8Brk7gIS8OyWmSxhJrOovGll2
4lo+mLuUfhknFIupKf+m4w14F4WfdyC8CJddK0bNhHISbJvZ5nKkmUmInp3CZNMW
aRCXPt67yNSaAmULf/UU7iLamsopJK9X7PGHNdVoHNofGUM0oE9ZAD+Q6uDK+Sqy
L88SdSXJsIYCIOa7ImUgdHqZsRZ90fyCBZZuMxfDfOgOldI/FW7eHBSQ+5ik5frz
Ta50hQTMCb1DfzcOC8TTzRF9xpR/LD1rQI0103XQhqEmVX4vM+c9kjrSMn+fSLP9
iNcx2hvj9aM+/xDpRunnVETtlQgPwxrFTgAvA5n0VU6T5Bhc6DjFyZD9dOfCwwdA
nrI1rA3kcuiXE6hoNzpwha7vhO0m7xMu2yD+ZNbBSeN0J6/otcBp2GTnLY+iDouM
Dckr8RLaW1zGd8dCd11ZMFZUvE4Yfv4C5xV+1SMnE6dUeFITMpesn+rN2eaWzpBi
ActJSsAVIfr2X6u/JKc+Wvp/ygGu3MMnzhcWA+uD81b/ozWiFVBbm7y+hNVJJY0z
qXU9Uqt+fK1gSyklCwckrOxd3B687ryEgMX/XG4D+FMvcRBZRKXvrLKQ0XHSXTaB
Y0QFnTkBzjRNZhxQewo7n3VpWrbHMXC5JAHd9lc5hO3bUg+PaqlWERUkvZPKNHwN
LsSG6wOH8dCD5l1riAuXcYA8ACvmk9vqcBvaPajoQ1DiKPYBTZAZZ0pYjmqjIch5
RnkjcugXeQYij1gud+Pz8lgeQIuYNH0LwLOAW5ha/cTXMG75BIMMkHCvc+THe2np
c0MJR9EWgbEfH6ZE5PEmt0PVEoBYqpcp7i4Ld2KW8bsVzS+CMiJoTPP/4OP3XvzV
Rmo/MGSpL/wg1Aosz0rwJcwC9+xSPB71LX5S77Y2bgPhBzFU1eVkikUlPEII4io2
7wDwEOcRFg7VdYP7D29cXjBESy5xuDRwG8sSSmTfT144gIK/Y5OKjLCsHcZY4m4s
EeHzoEpK/juKPgb6HxBOhC5iyKxkoWQnGHFDUtd5ljS5Nwigt9XpZzr0kl6x4IWv
aZ2hwZbVpMI5F3II7H+JIyhELJInZhdUp81thL1OaYRu9G0Y0iYaIA/F2btU/nYZ
/ehc+BE28/8vy6nma6Faxkr/+5qK0Nrr7z1bKQyw+PPGQnKNIlhPkhsxEo5LylUN
PUVdxomGJsUb7T9xLaWs5WRTxeSittKaPGSvqQrApdo0SXhq9rbnc6RvUGD5r01Q
v258NCYs170zPSTxXmKziuFcdrxB0J7leJV7utoWFFxG+iToy5bRPmvQZE96gQV5
p7eCKfTvIMwtJ+SbVYtMYDQxtAqA8tRQxZ1DsAV3bW/gaKKbUllgwqTJCVZJRfci
BtDQ2klkVi1ZLVrusotwaLHFtNchwkwSxn8gViMOVlgQMsM+0THdp8qBTvNYR4f4
+N0Vx8Himn94yNfvo3N/DJzX5q09Ak8lAEkya9P2QmXhYpTQ/JEGJHGzc6TgaagM
nS1n/JncYbQkwCDdFVVJo85SstfNYhFeg/PrHoA9GsiubpoOqUbPmDmhXTm7fp8X
1eaSQK0amqmOLbTwYnwZoi6Bt0MZ/kc9Y2wIdOs1Gth4sdO2FaZIkKY9AxcsiP95
nFPKjLXHk7UhY/aOHLnYilxgNobLzFO97QV4WoIVn9Mx2MRrTZHUqZPTpRvjkkOj
Dj+W/eEsWZz14phF2SS0jjkbEefWK+Nh2fyIqap2n+gD1xUr2QrAs9MapPLrzA0P
NeZ2Xi71F0tLbeSUYfox+70rIhSrXf52XxfnrEeDm9SkLNh6vmEdGGnPB1/s0dVv
UlP+z7bgwfF8bS7377PAweq5oDQYo3fxYctYr0R9yn6V+XpWQIgMsOGlxa4inq+L
1q4KNZYvcUhibUht2m1im7nPhIb+eTWLBuOo2gdOymZExcBQZIa2bT5Hbbcl9jdY
4s9UHQMUW6qDf6aIQJzPKUsaCjWE8Tw8dGbdbKgwALg75IdZg23A9e0BprWO0x3+
9RrCutMbPVhClulfHTCtk9kV3UDH6vvu1cRRso/aXR2uv6PUxyquazRNbKg1XXXd
r4DCFxKbpbtPlIfzmdy2BmM8bn+vFfpJOKiP5956W3E/Mh37F17aVUJqB5nkP/a/
mYVm13jivKPSXp0dJmisst9cmzHleSe4FCI641U/McAf/ZNbhxYvZ6Ymw1cVjJby
MUb5oxqS/S9/z0Y3XymUAllncHVd9jJQnWAY6Icdv9uEwx9U98v8ZUpR+Ls17kED
+fWFBjCEex06UMzODCL4ekLO/+CkMdfN+4GGiybDdEoC6tKC8/zw1myFe29zjK0c
m9XxZhcDchOOXkKBRqrtQ2itvhCfP0FTtQKqjl5jWszB2u/SfJkr0470BHsrq5yM
2eLpRV4Sq9jrYITy/Hn5gBj9HNH701V0J2aMNe7/AVZ4NhqtMujLbaDnKMTbmmK5
s2aLe0ZteerRgrQTZdpRgcrjPW/2Ka461Y8g86mEUwzkvEppDRA5hu7sPVVdupie
gji6YlGk+SaCp0U3IpZRp9P4K79h/RZmkTcipkSQ/DzHK7G9z6tjAOkMOW7rv0l4
qJjW1pqpwh3QsTX5qObd9m1dPGy4LtkIFbG579ZPqu2Y2tc0sNq3EFOyrOrUkepZ
ZzYrWaN9ZcImV3fBF5PABw/+3VR3JmH9QLmawMFV1A221h8t+MOMqI1t7IegmZll
L+UgFkPg9yFwg2Y1v6ibUUXIRk8LyWfYqTU1fgYf3oBpp1HpdRFHAIUouAyshERf
QWMuDg7sdAkVcP6mwWwcswWm+sh7EkGGuVkDnOf5aVJcjfMsldLt9EqChEPHXhYE
H0R8+P+F+LWdbXToaaP7GrYBMhn/qGjs5wRJwobudxSFja0RGfR/Eznzmo8xCdUM
S+zelRrtehDB25cMeleGvVYMisOsD9cYkdmXUMdcbWGdtouVMEzGuOVPZL6Mcb/j
Fqae6oTqJkFeUTsUOPwciF1fHNQKSoBvVJCWNcJXydncTy0KGQvhqhxXjwP0Ldmz
Yhv9SOsJWaiZJJ5NrHHINiLXq18qACwOPQZY46fdzlnEVo/lkG4nxa0P7fSRyquB
cQr6awr1ellExYwHmA+iel6HiMdYcR5Z1oWPIeJ3SwKjlk+Htz6XlxlQ05hFzK9L
iEHQE61L0a/STuhtYJtHskDpe6WGO3qUi6uJ6iVz5wRcqKNz3ae/RFrSsXuZdrw0
E+mJsRwMZPcpZjK45p+d1q1E642i8UV1KlbVZTOazcwzpH47iSw3QS1ReCEQaHTV
XbSzSZzmak2KiQQdxyePdWyfunXn3aRpgS1LU3EDCes+SeLsX9epbW4fBTcIVGl7
5e2UuGhtEw4w4w9/YE6TOWysAxRWlPbDz65tBD0GutBzjAtx+CIj/uzE9H6S+WWU
3BawTkhy/CZAm/49cYCq9HuBxa83dgXC8Pbghk1YjqJyUW3jAJ8yKVpEK9bFqXOg
Wnaol9z+Z66Buud7HSTktNnZbgIvo3DaoeJmUV9z7sKu7j0JqWeD15DKZBas5LQ9
+ETT7m+RL120mn7cpD13mpsGFdvHEhusfjUFDZ0ssFlWTNET7r2TNuZitwnh7XKQ
NSqMZaBHg2QX0pQI9snxCVoBijTiVFOij83ntU9nGFxGggoMWl0UAM3SvSVhN1Wh
LFAR7RX9/eLfhuaDWmpY6bJeuryTknUoGYorfKZW4FRLqrNVtcijk6XNtun8m2j5
J4ZEwPVGdXewUj0mNy0wVAaahUdGtukBJn57P1MzJEn536TQAD96ZWucV0ifohsN
JEx/UB+pxyczjeywWCsrXcQIGyGMkccl/rdVt+LlubpXwzHKNtdJW53rQV8b5cG1
JGfcpbze1qcAK7TqSasL5OnZ3+fq9HdlYIuSQNpwvijVQg5uPjpp/U0QCcwsrnpH
zmc9MGB+T41H4QJiboNefl8WsESDqE8Z4eqY3ihwgrg5jHEwZsU9xG73SpJMHZHc
MN8szvq8kLHkKa2TlRJ0/wWbO9PBESfKLPltxDpUjBj/2FiEiSyQuwGGF/6viFCD
744GeC75efFfUCeMDd0bVy23f/7TvU7gncxM7F6A2TNyAta5Jy+50I3WGK2WCC6s
DZivgUE37v7cLFlXomSgdIvyw/cAyswv7dD9sl1I7w+1R7hGFZ2IBt5r5MHMZbXE
c945hpWqkCCgNnx9xhYtnknYa+4uvsZLrwlya2TLfKEY49dc4E1LmXWSiwmhuchP
eR2uvcAKQissYG7oWe9676mI9xBjqA1PXFrRV8YTPsNWgf/GM6vKNK/t+RKJzcMC
ahPJyvNHjO/byuX84Ap1elRNrgUWFkXI3s/IGbEu0UksFP8UfjH92V3NTvOiXeMz
P6sf3+oIIIVw5LZIp6rTUUEjb/l0R9yW4UDgaeRTtObHCLLgMjlcve8joXrHLW4M
qgcDmRWyJmYk1CFGzV380TaJKppf+a5SGkd8jqSc/HMQbZ+jUi1VSsZvFaNeHt1O
9mO6W4dyHMxrKE7N/IfeFDH/8K8Qdyl08iU+I5SyPh74s6pLY9si7awtdNBs4gk5
RCa+ii5QiEjABwHajwtiwd9ZWqSx5GOnQvCQIx/fpsaO/OZ+g751aS3nMxsAA8dO
X6QOFnguljDSfYiAijuUXNUrq9Le1lnCJueo9yll/c88WlkfDYpS+mZ07Mvq7Ynz
c6OnpmfV1ic2pU5eApA/PDCiUbnvzi76imaR65bJmRp7sHCAmnurJfMaoygHALHg
cGLItVEccQ3oHSYdp0YvOMVrV51ywg8Au4VwjQ5iBxmVQayCBkjFMfPOqpbIdA4n
bbZfZionh3GKJXxO8LvgOmnmbEFp4dQkNH45cPX6JpGoRURZhHmn9Uwtl1in71+o
Qi/YhEPL6256Gc07kv+NIIlTsSYVizdEwCECaR/k67vT6bfVKPoPvVH++CTqbAnR
1zCrnqSRUh9HsLCxrpm4I50RE4Sj4efQyMCG1XkVcCOK0z31hwTboE74exgdqv5h
ws0SFf7j0lvGx49UNJPt7IOXdwWwg/WnVnNqHRxCiG2y4F3eV3gcKZb4FmUrtIdi
1ISPDtYrRa9qshkBiwnAd3+4KySlO2tfKan5aEop6cl/6EkMt+Krb/ghaR6JROrK
eMdEKQpPDZ7+e2HYoYlkaMeZXni66RG5HddEtgzr68RjrDB3QTU4jCxpR0VpE7SE
Lc4FeikvRERL3XSQ0SoVHp/E88K91s2XvRSNURbU13afb0iqs4Y7tNNv+oSWZJny
u0743XbWkMKdHz5aO+1ro1+U0OqXSF71pDnAdVj0hQZt6QiPh/YUfL+TQ5Bbhp/P
Yrthfo2RNJzz1RQeXGPWB++cZ0Eu145eZtCKRwGGTiTqQGDCp36H6lHnSDTbVakL
WUaDrdx4Tmvr8Ha0VU8AlXcnLIWWCRN5UxGgmHdFbqZvzr4Foy47OXGV2HN+KH6c
7hmuRtoGo0darfHKh0YDRPonjiTCrLHtRz8oIPEXrdyxsV5G4v6UtvQ9nl3WshpU
tLhXWL9AJAppPMeswQe/JK6WTyJeu+S0wx4FKx97ddadkWc0MVEGl7zp+j9cn+kW
lhyaApMlvB0bSEAkoPEU4L80bKbu2WFAmTq+f7iu8EBfECrqe76ZYf+7Nd7tNI06
Fd8dJI/FlXiPWPHUqlBoQqMGztYmakY+VVmWO5nx8s7C/k0z77hEtH6dgjwpwNUT
uU76kmGEAd268MEFjVh8CZePoziBHNoDXx1yNxZJ0qPFQtTH97UwYExbiNXcjhzi
wYHb6cAdG7hXMn3cipQqH7pMblGuVcTFg4aT1rKQNQOOSx7Uzzl/6U4nO+QB79eX
l3dhTc2XNiAtMZe2sNaoYqaGo5V4BofLb7AGF3ugOMDhs/lUOlhYGudMbEDXbNkI
5gl/DvmWUM+neg4W4nzn4zxojmh2LEkDHQO2DxYtBnE1yp/B8kEqBZ8IitDTOuYO
IBOvUU8HRTB868ULjGJIkkkyD0IyVsjD5TAGM1Q7kaxTqXn26jKeaj7GCd1xuBis
2cN4K0fVfz+YVhBeQ8Fl43hAIAHQgo1FJf0WhzZS/IXNJNLfj6REZez6zvpvWS5v
YOxbrZOJOf/t6m5cGe/0N23JFhF9f76yKO86dUtXrkx0PjQwlSJ+6ftmlNvFT7AT
0iY51sAWrKcdOebe4MmTSSsaVBk//N9EeCoxmPuKgQ6ra9fRLbSjGS/4sMYJcs3u
VZp0jCTFtK0WW9UQ2rgLUVq4DOz0zd5PR9aBEzA6roSMrxZ9yTvpxvSmTR6FFy7U
91mnos1obf4dL54+4FjWmzlAwrDZ7tLfwOdbiMVQwVFjYfSQXehcVyLNUgOhl0iJ
EO8DlzET28tvmHKuolrH6i5p9VlD+zd1XgQtljBN8M2lkODpUbOCMTjqnwCuj2/v
j8zfm3RgTIz2roRSii286U4uWjifoTyt2oynWzHx9ws=
`protect END_PROTECTED
