`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pZwCY6M7aAM20uJNx3mag7/f1hyS7GVD9UNpO7j0CjDCH4S60YNj63QMH7YTlVO0
swpk3+12EXUXX3pTKQKltJ6beX3LeR6BqJO0iGW+0bqTHUHklzmj6YGiNdXoqPWK
mCfdUNJrmtHGslQ90LM/65OkRwZE1xRTMpBaYMQLzyj8c9PsBi8Vd9M9oI80fAUG
eAdPMZa45lhGOuk+uf2lTVYowsrprwo66RBTyUKxUcSqZeDKHuQUcJGFKkMp/T/Z
VZVNfpDSj8GjwqP0RIKMQ3Uu2uUaI6LoDhyPLUlj0e+pg/b6Ty0INk2buVz6r+ZW
2hNW1KNhXILx3q8aBFrzN4dWvhGJh4Ab1M54gMnht3EqyukpnlnJceMuKbm7lfHI
mp/qVdQoCyOx+qCvA1EUBYv8qrFf1fFQ+OvSpL8mSPKux+EKi0yECDPWgVwfrkOb
AxgPxSdlb1FKzpSRbQLfve9qF/dDcTwcieOFRKRw0oDxCQk/1BFCAG54oMc3xKC6
LdQFGGOYmCDY6IajK8F6/pGyrY4QNZGh4CkrkvQYj6BiWoLhVJZm6Qd/mc4oX5nU
5mh9k0wyEh1keWn1B71txtMd1b3kMUpTAk4KTe0HOS5WMKWkSmNK3Z1g7sFOK3Ae
X29ZgcQlq22LQXqJDp4xWEXvKKKCDZPL5PN8NGZdOaGBebykHaAF00XEE+LgaXZR
2JZDyP9c6IgIJCpyVP+zNRKyQTbOWPjg3pS5c1WJHd533GFOr9Sx+xN+9Uz7lEZK
6keGSd3TEd2bNml50cS/YxPpJs+AMu82WNj5/7ZnSG1RdCuCaPTCchT+jj5OpoS+
i6JkS7c1XYtyOJp2bdRecOxWT1H74OqvdFXb8YeI8WRTwUG5BXz/iadi23YCXZhF
50yjrHGHVeeTqbMKSq9sagH/7TtuEBpnRkaSeXCfghYlyUGFXIEtezi/XZWGgvXe
m4gkpmsU0RgGlnoHS27qCdP4Y7fPRDq0tNLkCvb1GEB05SeqwixUUoZ3A/RPWHwX
nWSg9GL8L+uwu6Ve2S7HPmbgzMnjZm737ADEMaBTmwjVWEAbEb42Eak2jChZp17Y
Ynk96FAL6yANUiRuFiLcYhfSO2JpX8HiINTjFnbsDJqdJfQ3g/Cc3+9P53LNARjn
iLa2hseDKH/iQ1PJB3wWkVxSBZqHEfOr7ZDE9RlVnqs+/chAxvhwPesAsiFQtitm
INn8dTRro7f6d9vr+2GIpoFS6/v7EpmeKXUx8BgCqctY6AISUvQiMUOFffTrVyB1
xcKI87yUTH00Xr2u/ZV0oQshRoId64Tsu7yBey6SYis+cdaaEDJzEUP587G0hNZB
8oaaw5zM65U/TFk3phtFcL8YwzPK4sc+ccWYnJVI2RDZq/Uyn8fCfsn7b5jeDfCS
4ELhs3ZBCz9su3So6Eom0AM4lssQTE3gzrTzdLL+v3UmUKOFioSfKNfbvq+3ceKn
GZPZjG/+H+A2qFPJ1/8QOSTK9YgJS1pxB1AenkBQuNWtaPWh/RlkWytijnpH+Na/
zSKiZCUXx9DZOxiZnOsDO2r01I0q3w0C5TfO6PNPPgH3vEs/MA92yZ7XRaC8Ms5R
FLEjo8sGDWkd1TZ8fXKleF4sSzgStMVP3bNUsWbvClLjapKauR/IT7aXdzn+56FQ
6p2wlNfr55Ml3Cmgc+/kHcmuNeRHkdAoZqCQnX63yibawa76YEGcf4e6ob9sCV5K
TsQRcX9OGBF5WH1+19ZkGcGhFlPYtv2xFPWjAa3Ci5b0RnUk2n/u5VLnrio+/fOU
xMLforwUM1YumYcxRmJR7+SxQ3AglibsfjK1ze6LeTXVSpc6LI4ZhknKJLZGax3l
UkyDmzeoYzMX+lSBq/kmOxvXHZyivSFBwS3wndIDrHt3278rTDZ5kVlqAK8uQTKw
qI8mvbt+oudAONKiEtJcrHwmj0+5ei5fiZK1TytNymkY4bC9nOXjISHRX4w1941w
vHTbgcFErgYyIEYHKzY5ht8TOg1w2C11opU0/Ly14fA8FBaA3q/Va0M/wUFG8rpY
8EE3j8oLYDA/p4zul3n/hSZPdBm7WcIhRDo9LmdIqmqmXGNR83a7UAw7rEDFaptP
khLKpGUaZ6R7R+XuwzcrDzgY5uAoRl5KLgWw9mHUB3lXcnNAp+9AQk/RzG7c2CSb
+TUuRKS+oe/7dPTdaPDjGqtr1S4K93a5aBP1Q0X5l1hhdfSjeo5Iwoh3SgYwN3s8
qDCQk81/EO3ZIODVwyxhs/FXq4qLZctzHIJTGnuC0AiVM/Py09WeVZ4UqEQ+vP4X
3zr3quf3f0Mljk8/hv6eiWb18PeF0sFF5V3KUDLN7GLHVyuSSpT5UhsIS1z4dArf
KmQJj32lgMPQohy/HfTRsmDOIaPlYU5a2iqv/7iiLWirLTaXqZbcMUGnZUnJpQfH
Jgq0PkZiNS4MlGPWUG1/mT+jrEnvm8tPGSCPLL+ABeby7ss7p4hVvA0H94W7KV0/
oLJjEifxBbXYKswPnnQ1ec3QQ9hRArdzx8rmwkAx8oXR5EfBMcyqLHPFYZzR0Pdn
wA7IEBIS9d5L04IkMMn6pB+/Uu5n1UlT/lRrhyz76XNrgzYHP/xDoHYB3ApQd02u
2uw0R0XmthzfIJv0cpAkgvKP4iw9g8CYLK1R1DyS514yd+muhI07OpFXIjF4Zi7e
+PyjUYfQDJTw9zQLsb6UGaX3C8wbu7zm5hwCS4FL8BMX9IlDWXOgrq/UK1/kinN0
dii5i2/OiiOAF7kCbUnZGmzLePurGpyszo6/OPRJ2yixxfmSEMqH2W81lV0qLjoM
2EAl486ps/jnN0G10cSqXy3yHp9X0m6MhT46szGZlqEn9kelwRY3wCpjEci94duG
EXuWc6GzeSx4bEDO2VW9SliP0lxOx0Vr+bmqqqweu46q/+BbLFUC208Yt5HWRzJU
s4LaoqXNI++H6mal6aQPJe3N8PZnvMJRKc3XK4r/lLA7hsWHpslAy3JElu1q/qFR
DoxtlQVJXyf+6MP79bgEu2qrsgiwsNXL2HtdoUUcc4YLWEQCjrS9BVzBpEdqskgF
eVMBKMi1/sd/fWFm7u8VgY5eV1axPnWk31c3b2PrgFepE/go2aw83OCrQGVuZMyO
qh3b0BvmwG0FvqooQhAEWg7cMibPEQlcBVjY04/95bDjcQHGuXiGyVUj4y91GFvx
FE+pEO9NsdyodXgveWxH1qP7iQvKQ/3UIvjHsib4M9iLi1P6hA0urfe97SQNOgal
ujY6axCLi+2VSFp3B2mBU4UXGcQVq5ZH1nRCNtkQe17zC/MEa5Kw1Esxr/QtPXwg
v60CvHScR+DCODJ7f0Tk35znQexzcb6IzY6dm0di6cCg+sOBNIVRABtrXy1s6Zhg
`protect END_PROTECTED
