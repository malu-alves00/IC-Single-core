`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
an8gliiPiwYPo0pSf6ObwrlDgCTfOdBbAYA7qeaZtpcGYHvBAHCPyq+2HJtNCvJM
BtO8jrLcxocFESDfuJgm/4rD2ODsr/NgqrA8J53Ve0edRD+HKbc0D542Gl+gHmzJ
X4Dq+YtfitIh+2yIjPlPSKqBrGRTVg8hZFB4hs75F+CUP69yGu7ZSekHAmF63Ijt
XlQIFL+VIn/CcEsS25amlg6yC0CUeNCtDdOzJpBD+p/rWIMaLIJsg5/HGJfiqorR
wvb7IpR1AA+HNd0/Q8LmUWTgcKSTmMxoRSo8hID1yp+TNFjU/KZ5wBMkWTP+Y/lZ
MhQgtTqMsDZm2yis+O4F3bZthjKLqqPMhkwC/d5GNwwMTOqr0YCKmrYsOeIHeKV0
8pqgmOtNyUMWBiBa0BsEaHAJN3AJDBua0B3Xs/1M0rXqeL+rfLGKcccK9wN22vxG
peDZak+pJMSCljOjAM4I7Uk/ja5kymv1/kVsSLG30Yu3va/a2IBa7Dyi1kdvqvcP
j91sCs7UhlJql+9l8me5ho1l5b8DFdlQEsPE/X/vYu4V0kynPpvOugw8iBeB/U9e
JlmV61CRvuFRNnOyBX9ahakduBwesvpVKIflgws+P0flhFlhEiquAqq2EBdcnIua
drsLH6woK/Bp7NzDCcBOK+fXB/RkGI5IenbvsjFPr4Um8kCGznzoNQc5n7RcFPlk
oeCXvJdZna/PXanph6Z7JcRs3/a7pBZkS7U4pzEjQV//cKofihxl6g8+LFwJ/HCx
sMOg4cihgbR3Sch5qvye6J9SKp/7P4YwZdmPL5lH8DzjZJSvdBwQXNgIJ/m/HjrZ
XGwoGvSpyDECQsLRN3iP6m4LHvoJqVifwVonQbkMjfN7R94tY4N365tFt/WX5VFo
Adu/6/N2blRDfckHPl7zA95mRhoou2ldqBjB5PqttSA1RhGjBrdmPn42KUuxGioD
9rHmwraDWYWq0BHuCzetXp+edGE7rRbsrh7MGKScGSYFzyeHQaQ3YLhxnklhcaDk
PV/0ZabPWhcm5hGKuriv7esDHUHjN9lt73TcR/8RyHD3lyNJabiPszDKIUTeU0XC
EBv5WE9M3vfSFJtKUJzFbkpaYsrDARJDSP9QaTe0BOYMXHEBhcGdsiU3a9S97EF9
jUhIePy59a7tRenzTkCFCj9Zkk8eqfc8agkNwTpGIrozoVA70ERfgY4INIWgccsr
zl85+yXdCvAlRqjkEiLi4AJWKpoLbYzvcSLfS2YmJal2lzqrd8JJZRO1RKW8+p09
xs50FWfhJcrFDk1r5BF5xffg9bPkL0qNG/fDuzhgncxFA3WXfZPpuYIzX5rbxzby
Gm5rnylaSVwt442GxDe4lI9iabG7L5aHj2ox+EcGvcUPCMwDaLZLB450d+v2sh43
cPFPaPhQp+4tH+IKpi47LZAM4D1W6M2CpMgE25MnJp97NsTnSKrU7xxYKkmlVU7b
dcQIdYENeqtk31yfxz+xncIeLfR4PKNCy6+HXo94JMY75Ti8NIg6z5sqzpXqvMLQ
tMgsYbsIFvt7vs+TyUj0OHMLOHbylFEf1UWPBw8EQYVaSO+zzu71Ay9AjGEAZm+m
`protect END_PROTECTED
