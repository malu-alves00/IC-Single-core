`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
58CqWVX1wglbXcxcYu5gVhlJq519kBj7TPoiiv48nnXshPOuR7radcgL6Gq5tmJc
KGFVaE/SZ1Wf6Yz6/vl3fXP1U5Xh5+/fNI0xYHR93R5V/KBHjOyrql72bIdrH0dU
zOCnmGiwI8C9+6BFERAXbdbOT3ZFAP46HJMCKdkcQVrRaVkVM0QCvtWhYhoVK2CZ
780CTPT+/9pZvwQFAPXw4elbWSKMvYpHGPPNy0X73datPA6UGrS/VyfyoaaU/c0C
1r1egfa1cxZsi+ngtDbauf62akkdUJNp9AiUrfAbThxXXynYEkcRlqnVyXgFcvzB
Agjy8vCIoszAQIp0CZ6wXDY66Doh0AV7uPYjWlD/AogOOjww8KHoXwWZ4xLzMbM1
gqndG/rUM6Dy4znGI3N9kIGye4NKUWWzG8s8d4bz9CjJW2HnUXee3VF5zcHg9gNO
Q4ginKMhTZJV4UreOhScE0E30MnqCImtQgWJpP/ft2k5vXqQH9bXz/CaIlID98NE
rCBSZl9toyOIbiOpC3gosPObNqlppPBLklFJGRaukd8MHvtPZpkDY4Fm9oJjz6hr
Z8H+wrD+HonGalQqoyCTfdQ6h32denCAp4qlSaQLsdfeoGXhcf3r4Pymqf4KULPo
PmGHKZ9WNeij5+qTa7aOl9tfys9Db/oEcPpBzxcjWQCmcuhHWNQsofV21JdsK1BL
/xqmr47sa8yoQxUvgaJb3rEi6WfMM1/GgQCqsm+XHIhrnB8Gqf7ICwFJmOZPQznJ
K1nE/YILilidUPy5E6Mjv1Tk4Y7zY/DjAldT9xfnBr1mOYoN0iLDGuCtAvM4RTVh
5O3hbUUeTde/4SrFoZIUmK8369fsZaNSpd20KznAnHsXFGI6pBzUP2EImLQjp6t3
hrfKsiid0wIPMZvZBgI+Zm+OmbASQc82Y51YlveDhtw7G6ejnOa78wHFgXJN6bhO
E4zC6meFUQrk3vKp9nycvUShqXIl2KCIy9cD9xUqJZTvLl+RLOI/EeiiiPjpcQTY
mQv0FgPww7oZ5WOc5aeRXYMm8BAcrtYsqw20+cs59RdjI0ix+Lz42QyBLiZdWG0C
k9lU2HgiwfrfhhATYNtECdGZeNkRIu5udmNPx5d2p/nRl3zv2oQXUhaZw9D9fQZG
1CaM6lSIPU5cUVxzC8+snrh7u6rCFwj3rMTsKqRyru4dS5h5rUvuemLb03vVy+y8
mTZmh8Aog2YQEKly/cpx7jzdMHzzwYXpFUArMlzA+N9WgGyrYBnWYH1j2rA8VtxO
UniaF1nykeW60tsUTT2romEkJKCcK8vL0ZNtWNFvrhjmU03OuGDj1phH/NzntfuA
kROju4eBHudGatlXoRCFmn8RhqrOHTUJ6pvptZtni9AY2qY5/DVVB/9TjtDch86N
+y3gBH1cwTomwlRTr40MrmYJRWexCwAXCDmlrU5nLEVIvQ6Lb4hsLuhxb5KSStQg
JEouinxbL/AbM8yzueg+w8weoSac19bv+OWgxdexMyfGRTbhC0+T++e1soxsOw5z
2YwOwoWMBAzcDf+764sKaFdLqVYotfbwneiJ0aOIxnZGB7TWCUmeyke3xrhGhaMQ
xCjwbadqnPdrBec4FlRFoJyW/Ni3n3cVgNYRBsWPfroTBk+3yy0rEAplvSO5dpoL
gbNI7dd5ViLyyikzIHmcmgV+v5y9Os89j2jyac7Le02DDYac6zhva3LF2v8LE9D1
EGbpUGkry3AScqHfT4trgysgXxve+kUztzQOHm9HE5jIZSADUGgEzkZoP3PAagZJ
oNtQ9r+1kzO2gCipms5PHl8KR3IzDRDxwaDQVPiqJfpuDOWt9NPX09RXUE8xFPPE
6uTbk6PTVyjezgqJleyf0uOGNSlBp1vJcxRlplQ6Bf37dX4EluGSEO9h0Qk/xcLp
U9+pem59C9GapN4jTiz22w==
`protect END_PROTECTED
