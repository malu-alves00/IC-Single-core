`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zgDT5Su0PPknXDF/bb98+EFsGiQ+8tjfs1g4FBUhosMOoQZNBKvuQJ1NHb11WmiA
DR55X/aeAlpCLybFtlxT3ty19fSReb5TlHkL7dvEfKUvZ1cLGmbV3skxnc7kVE6k
FMzI3VzXsgabOaTbPi4GtVWPrf7OBrFvVShwl0kKGPLL6hVFepJLaR2btFxt1i+n
2SNIHYVDePjxxslw9LyRbcd3CRHPJ3jJ3tz6eFQmmszR+tWl9HpiJeb6u/3haIoN
KTJYNZA2kSXpwnaoJi2gIyJf/P0nbmgMR37sPfDlDyxIw5j61pZHBLrLtNl9Df1f
DCtcMgfFVPGlB82wYiltysxbSFSx9NOZGHmN+Aw9pAKzD5fwKuH2mCEUcl6iPhak
qjYQm+udhJdxb22WHVFfKkRENX0jLFUzSQhYKlmCIcDe4TwGjfd6vnWNBuu7C1hA
3M3MI++Rch53c6ikKGo/LuZHA8T9kGbUE7owGsqFxkRvSoIN2wBzC5Wu2oBWDXmo
LoIs4Y+mdtbaTxdbuwfkC+o20A1MwHSMZCC2uRmjBGba58oTZgkp7Pp5PtKeFyte
Lco7MmtSxAyot4wqCCHHU5ZISTNLRFoaxTmWBfLq+DojEj0a+rE5Bh/OEXp5izAh
eFsh774IQHV8qXdBvkCbS2fPL7kXVfbI4RLu/4YZ/2NLqG+L+Kl8HKq/HuJcFBSi
Xsw5eDytAzMWptZDYlq8uaXhSW/xWU/1vNrLQj1MWoRmsX2t4FWG/fu0ed8moKoW
wW2uXRGVrz3Dw0l8MFsH+gi2XmPYB6Xx1rDWOZHSWPNpByZFfbHQZYm8L1UoGBPX
wSW85FJJmwnDRa7rkTDQLqAivcuu9HuyDk96KOc/zxrRddZTJS6t/oyTiTOf6QCI
kYsAcZI2YVTkRr1hup88S8qJ378nIRUz1zl2/nekJYK4EVGX8YPjpQkydqlc+5bE
yyrorU/Xb8VeEgLHuLXfRIodqmlrlktzyifYfPcel7DvxuqtjW1KDE/NfKEQ+n0m
TcbKcyFv5+mn/NosA8SIPGb9xIJwusYjwMxJnGIJA32Q0+7QAv1ir98Kf+/EeHhj
thinyIFy3Upcck2GHyY3hHcnux7y/Grm0OZx7DDrjt2RV4N+Kg5GxWBz/GF7LBB6
B1oAXrEV2Nwap+2DNQySs3896tPxgVVbBJhC32HCXWopNf0odu/MqQetOImBYLPn
0h54Rz8vNOVDK51OzWP9EcZVx5pBsd3f63Gdeka0aEslZhtCgYvDyOmc1mEwJ5kv
dgpSpdxHSTlx8MJ++sOn48p7FXdYDs3ReXjH8hFXOA1scgLyYDufRZ9G7M3qJ/xT
zgwcJvb+6IIC+2kvq0PxvLiJSfmj1TJrd4NeaCQ3onYbdF/vt8OvoxBAjXFWEV8p
Yt9cMxrJVZdBu5OhXv9GHd1V8pfcRAqLb1KzYvCCg3d7bwLF2nvFSnYQtSLIF2cx
Z0xdFgTrDswOkXwFJDCuR8AIOjcXGuyvc3UEQZdPQyFZsjIH8dq34jFBiFpsZm9X
4L7lpfVUMSdGdK06wWxjxFVnHKXb7epJUyWeOuZeX7PEAdmioQcv1u5z7CRFQ9qu
P1k1TTOviCLGRHB/WRBFPB0KzibbZCaoVUtfrRTJAvsy2cDgapCIdn7Y6hKcFDUa
3mKXWZufaQ2uFFoBrcujJUU5cm8yBwIknRBZCIb4oau29Cl3Q0BhAbVDGyFpSPEU
wjymKj6XPBMQEWoCHyHpVwm5EBmAGQA7onSM84XARdo=
`protect END_PROTECTED
