`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RgpcZYWVF2XuDmtwt+4l3qqrvvkNdHvWHxsTqLg5MJ5fddXwjDmRb30x8tCiPbIo
8NLPPf0fgL1gBc57WNmOhq36QdGXSGiTlgMNYj/nqBoLcwEibAdONrYeyWK84sW3
qRvEUXyOgaKIE2DzCgP/H9pp173KW1PQKcZTXzliEH2OFrSbkMDsvNZ8LUK4MEXk
XZbYc9WC/jOCWbbFXTIwVn4LR2QHRbiXRxkFAtHIoOoclw/7vRwWaD1SUOi+SExM
PYdHmnpP96E+9sAhPHnrTRdgq1SEAJvFaM88tQEWFViEXjvOcdwxTv8Oyq8h/Xpy
yG06ULk+0yumwTs9gnEexDgiAARlzIlj1HHl9D/RkI+UexMjyhcXzh1Ikk9vJjAG
g0uTA84xT55/S9jRtaRfSbbY01TdT2FYcRiZKzTwSGjuCtrFY5tFIeglW4D6AVdl
cJHo60sJPHsmF6/XmAV2wi7drMjBZRy5NbPwYwGWFGB1Jht7qCLQHTQeqoYJYd1P
MuxBC0jCRTzoi3XlOocDF8JHWMGqiyjU8j688gi9/9DS+Piavw1hdNbBaM1gND4s
gM2nlxg3h0M5hVwhV7lDyy/j+7BdlQSTH5updMA+eD6011d6qOayHxfMdx584DBP
Kj6CLRquVyncp1v+yoNxifcsmiyK0I/wnCAdrH3InCkLlE0tPtUAXWpki9Pgo1kA
Le+CFkaEy2dvatC8nT/ujnLpb5nx7oO2gmGElrcjAtTQfL4ub3pG+p5E+2ilnrFm
ePhAuN6sMgKccd0DoKdj0wvi1WOJl9xp7+UEVM/TPfuRSqUIUjlUbR8IK/rQi9DJ
VTEMrMFG7jq8rW4547749JoGF5CCn8F6EhotHFhYLScPnaFFon7Hrd65GsPMsqzq
gRsEBSSCGUj3CH7VmuXEQl55jnD+3fUrwcSakHDVuuTu72UTV8En9MEQA1lEh+lD
FLW3AiDn2cu/LfD93gKZOZD/wWdzwwGfK2k+soMu22AcUW9/EYj8zqWS69CJmc80
58mViyaZcH/FA7FqxZsOCiiMG6fJeZ0NnQPPcf6i9s/skjPP16cR9UydYDH+RXDI
9pjkISqNBsbIX3RBTrkKlkh1ZZpKT+u1bOEHPp6s9Rvp5jGSZr3/uOfiHeO3rvSy
i/nK8G6fz0sn2jgEnbOISsRZMOro9GT7hLooK80WrLzWh1s6zhA58fzXoWjNr+xv
0LHXN+T644NgcNExgUVuvV1MLaCopFayn8zz3BvxntHAi7vCrKOI4yh2GZG4X5uD
CfiLIw+Z/Otx0X/1sERCbwItPgIpRqn8cYmvzfm8xptm6Y3+wNxo5DN+42dtx6dZ
CNMEmidzfWAEneZFv3xnpPX2QdzXfbxlbEyGlckcHSCWqqIbSoLlqegK5hOU9n9S
NSSWorWsGnHG4Y5cukpJFu+VvvaXgs7GHQIG2wkkLJx57lnneI3PVRV6+XwZBGpr
oejFYJxgLYtb/hS0gNUuk9qA2TuQT1TYxqmBX3kp1W8oANB8B7kOHtEdFu3vj4cZ
ptuLaev/AE+OuQggibpsUEAFcqS1NRNAgip/mwqiji5EOdY8Uie/YcvXVmz6JU9Z
yRVQpoO8p8rbDWrd5eoWrhdaqUPk7ppDj4lBw71lXAghaL2Xh1DqzdUqWbZ3apKn
Cki9/Otz/YoeArZ1OCc+KG2p/LvoebxMg6DHtsNxK/Wvs2obGTHoWyE2nLHzpK3V
vHKuA003MeRb5Bza6OC5/khxPVrCbBME34AKAZu9mSUhaizbbCPOAq20jNcJrs/8
t+M8vMYqAWgIwwUL9JLbqGLYsKcGmcSE3ctvHdF7rCD+mm1818jWezADN/XHWFcX
cU4D+aYCNUZldLMklqE6UkTUJYOkl9Wx+iNIGJ5D8CSZT7KRa3pJSO1s+wPD+sGc
5KObyZrtXyaOxJDnx44HklBrekpRsZpVYqrjmb1Tw54KsvKvdMRECBBW95i49oPS
cmmPrP5P2dR4ewSzK5bwseZPuBcC3Vo1wpLkYIgw4y4HG/0NB3p4JtMiIuuRZFIo
2SoSLYHIfQW70QB3JBlsIFz9+3jJnbRMwGG/uJMQbNdcGvKWIn1whhuAvbriogSW
BdqZFADmLjx7TRlBW9nkZPoVHFDR7EXZUx6K5MKw05vO/BTOXd06MtR4iYSFxA9C
nlVbVxmEQsYw4K5EadDzjeD2WJHfq6jvwVd5NkjNw0VHnU+ncEmT/TuyED/IerVV
D5Hn8MD+P6glsADxhkFZ0a2hTNavzlbfD7VN9mn6dARz5LRrS3yGB7w0S4uK/s2m
sP4rbFtronJBVzMRFzZpK8eylVXb5BLH+rdWIVRIjB55JQCL+biFD83CKzcfJ0cu
RKY/O2/TZEPdRrmhleiA2TdlKy5slqmsDrOx/8CQeYI3AhVwnLv410dPIkqtwJJN
/Jaag6t+EC6NDPrSpfcpXqkKfrMPF5zYhQBbpZZMc4JM4149G0Pdm0DJujeDL4c+
FXY9orH4+F3xdfQJUBzfUZnSkkFAvstjMeTaoqteR9L/T3wUitikoBIxfXAj0Sc7
B24JPzXd/wOI8WblKfSELb/ALwMtfoEPz1Eqgh3dkwluErmPucmkim8qmA60DAZP
uFmXoKrpmfQO+ccYKyyPZSMRjwCcptg5JaJehy5/LaV5/Kbfp53R9I/8omcTHzlN
ce9lR40EHD+7dhT7OOI9RIyfJDE4SjxMeZxhFe3DSHWsOc/TwGmIbtSFDYI+ri2H
QIgTGopIx7bVaM0p+rOJAmK4hTSFedfQYWjj/s0MNxxEEyJBmAZRUv2xLOS0OAkJ
EVhARw/viW+4+iHsbA5uX7gDg/15uLrf56Mm4osqyv4F6roE85v0sHpWPYWZK8wW
ygEJUqPSxKZ/SaxeBBxCMOu7iF/0hK5RpwOsBoVl5dI0qaEKjQiFw7kNzVrn3vdg
af4187UuUHW18yLGXSjz7EGPTIA8MjVNvlZ+X0zWodc3NWg17Fg/lnRLINtdabH4
8a0YPadaTA3+xyw1ZmWxtLX+laiT/Tkz4wBBeMR4rMzP+XGoBKDrGG3d9qbybPgf
KVBkYyGrJLOVNUuJ5G/43JnXjcG8l83Rg1P14dpXNeOziMkA6aBU4Zg/kmht6iXx
BdfHtP8dYRCmwCjl/1XRuEOATePtw9xIiShrXPmppqjB+Z/P1aEIrOMZeatAtznu
jqgVk5OVhu2omEBXNxJZCnkEgKkilKzAhYV+/FGWpXlKLD770wz/iRd7s3Wq/xRs
wKeTa0I0KSlYGEZ7z7iH+JqA8pBo1yIqUPP5X2Q5OdUP1yYOmnsTkXfc11Cfu5L5
5HrelaRLZOb271K/qTAIB3hdWuBErmZXUSt757rQlC0Oho0dx7VMZPYY1hqBQF72
TipSuBLdr72OgLHU4Y62fEAjJ49DZQ5tup7QS/C8pnOwFlfOpkYlt5LG3Ls0N3VT
R/AwP7NaylEfFbi0hMDPS9c3Vmyjmai+0V1hfJfUGVQ1GVL6N+PyyDw+4emVnK+K
OnUabMaD0ia36DsnVeZEZfmRSD4FzHT1gflrIhDi2aVrJS+1n+FWl+LBB+4/dn2y
BxE3aakRzoeaxBQhJx4/yX9zJQ7aBWApZxNqY0SfI9Fj0KRhrWR6nDrwHExgdO72
IAddcwzmdRBxDDfY6sJ5PiFdtF26fZb2g+Sx7XySBrq9WW5MJdiKMkmNFG/gakO6
P5v1AIxodZe83yKNrCI8SA==
`protect END_PROTECTED
