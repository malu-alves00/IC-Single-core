`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ohniei6BwObgaujw8Nb9Bh1cHE7UDFOE0SVuUZ2+r91J0rJOHPhQxbR2yoQ6d9vC
xOoHoehNVj09DHrtinYhIi/5HsTRX74liNzZTh6k+iWuHly3KeeCCzEqszGSZYJl
qDEJ6E0TLBuh2R9U5l0tbTRXuyiUrspsVAyAXU/2O6bXlySh3J11gf6oXYR/nPW4
vwVAkAMzqzVoOCsIlCtVIF/J0uNB/4VkK+ww+dv7ECJ/lBotG+hw8wpZflPPiyqL
tkTPsxlJTr06xkifMYEdQuy8ZMxsxmHhEMAUwmDacN2qdK2Stv0Lrogujv6KBvhD
B6+jGFW6d9uyd/Gyx5qpTHHpbQep/fQPcL+ziXC4SPBQHFPgMkFr8UBH1sDe4e/S
3zfpIhzgoqgLcj7dOOh5lflVsmk8sG7dG7jeWq+2hlNfgteZR1cq9pxjuZjp8Q1X
pWm0InWn3n3sbt9lOcSMLioFE0o4q1U5nq3BU6p4GmnD0sXAPMssAarA2WnA5BnT
oCam3ZF2Kpgt+ROlY4UeNyGahlrXeB6LtF1iPTTvDkE=
`protect END_PROTECTED
