`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jm49bkLdAPoOkNzV3MsZHWuSC2pGkBBE6XBJMv270G2ClIh7/rGdriBRLQRYTmA2
JI7tUYvKD62J6TzA0CXDM6EOP3LW8XMcdBmLG3jrtR+3X15LPmOeAaHl/7er6IYI
ILC/rlaFGX5Ez+vRuJdNHA8epi6MOLtCy/0fVrEE5y5jEsgOaRxkXaxV2FLIIIFn
BjfQz7mGs7ePtAwA+ylsIXdzeFMa0nLF30eytfNENy2r79Ojh7K0km+exT/Oq5wi
zLfvOEWg2GXCDdT6RdGzITd1mIuNmqEdc2GW/QPvNKPLiiJ8IIFLfLQGMezYaGQ5
lmswi4TkncmaW93OE9omJzyHLfqoweu4VoBWrSaYGnGyAGPgAPSRUaSg2J/B/aIr
sxJfdMYiwktM54zxFYnFY/PR0kpELAcUay8pdpc7rkaGv1mOCapBQFpxXUDfGno+
O6fVWh+cZxwcC2QVJqpDmcWXx88bsIBnb0QlSmwVb1+VunXLq+7qhmVuLGHglvSK
iUrQgR1DU02ASAYfueKBS8wFOCPcKNc+sLEii8ddDnk78Vf+PG/c3tgSwau3OItr
9aP1+pzt0ArrcLsRTEmeaPkgw96yqEzQ4FQwCWnIqgu4NM8oHX2v823CrXDYt9mo
SnLUuCwcqGNfKjAIKcug3CADdxZSyvEEJBgJXfGkTWYBybzjGEKz4/oUB4U38fZF
aLx7NaGD/1Q4VGUAqJ3aU9CcI0+7/UbLRh131sXRZz93eHZYwtFkcjAA4sMn9vcS
7bAL1VU8dQ4k4VHgSHyWx2/g/L+uQpuL3hf1IUBEAU1z3CKKsv0Sq/x8bRwjY//w
tn7AscnZsa6IXYah7LQbkzEfTipriBQ5hHZU6U+C5KijXvOVTC8kCQL4AAGCQc8X
lagig35mTOt1UfEDKqeEDXxb5yo8iH/8u+z5dbuKM52e5JIAV9nGWtL+jkRaGEhZ
kfm29hNR/aMt2hg0xJCkH2Hhhm7TQHZBWk1gyq4SEbCT/aAtTqFLeLgrC5NTLlws
kE9ezmaRdbJKDwFIDRg7+jiRwaPzpTGdGNrBcHgtNcr2WLzx9kAJqEdHSE6P1mtW
n0/vJQR1XI8AH3SsJySa3teRZkAI/SoyzO4S4JoOQfiEMZTEhyPfzLG/IKS2rqNJ
qbBjB+eCSujDU69LfuPZHEOU9Enq5A0uoy0JTqhu9hFDW7CoMOVI0SxU1as4C+Tv
3p6WkFqm+6iLfo04aJxthF1tGzA3aTJfFdMW6LNQVUK597V94ZmzA/ClhphfQ4Sr
QeOZGN5j9n593P7knb3wlzkCyfAQV33OSolcndYRx91/S/Babgi2VQGq4QpqgAYd
RGd0RbqWmOIGgrWnx2XRKoY5yA2f/XohDN1SIiV/IJhbzkTBR8MJanaBlf+vNjMy
pWy8uL52P5CpMVZbTTfa6zWNqedKdqMTXVHA5oLEY+DzkaKKpefXoBOcXplKmGu2
ckfJCARaAMX543RR68/8V0YJ0PutSSIHKSa93sO3DTcBD+ep7Dh2uqbxKp3YSt6R
5tLLmkOpT76oHT0nK9jmR9Ap8B6lHLv621YgOls0bKb908q6l4mfQbpkjHFybxO9
IaJ19RgtRmfjxrMBwAOrvKyAgDwAGeEKNM+38KYPEifC9e3JFmpSqjQTiu7bNOWR
UHXuppM2FuWsKHH08OmVwz6X+FEgFjunClgtvQYvDIEy2PSuBXEjWS/KBwMqXsaQ
r43TQaj/4dGE4kO4as0o8o0BcfodqDHUK9ZzrqjowTelb3Xpd0ZgVY8MCAXxqpDp
0IG1vks550+qnIfQtBqUispPuP4U70dqIQHE/3NF9jt5vRmJi361wKPUnW00Svjc
YSVnDtWl1TgDNvTMcK3Tz790tiIfS0mNklBXW0lKxbpuEff5aTDCujol2vuzqwe/
MMrDubO6dWYVvkcbM+P53PQ9LIArb4gB1mYjQsxTNZUR7m6v12mfe+4zleXt21Hy
oT3sQrgUDF4GOJIREvWHts7Sb+nZf9UJeV4B2B3HIG3jJLDjXjUHCqVKX5J3TwDd
sf7LrhE20p1sGP8WwUEcZfE3ububPuKxughLFOrjU5qjcJns8m0wEfEhbXogwVHT
jME7ElXdl+GjqDDjhwWSZHPmJldp9AX5g0K+WhUJEeKxzJKMJfoz9BUiZBDp+cqV
KdF4jGNUDTpD7y3fUimULWhrFnvEGmlU8joMBHet9V9jxvT21DCCYnnum3vFya4j
+i6fqWqjX6VnLCVl0VQ3C0zb0fca1+6HzC20oMB/3qpADZhexI4xQeyJGWYrMhQZ
oAN+AJk+FRLG+U66IN5pJnNrb3pAvXa2y8O7IMQtBFYXNJcNyLsiB6CptkiqpF/s
uGmyGOr9WD4HJRKBMbWvKiEXYr8m1pCGht5ZPmBzXqUx3QI+mt5gsUgoEQCtNpyS
QpBBuQd+vWHgmRAzE9FcbapAXZaQsJi0oMhIR72Ghg1inxPf6Q3F8ydbC0b14mYs
4oAZo/z4Y5xleT4KNkyXuzovq8nfRj+PaAyYJqPGvmSUpkeCLuDOxDVeQUGFuNCs
JN5oWp0roJKvPTFWkw+bum/Ctyl8pLIhMIdkWV5DcMZNWYeHVrtE3/lIFoJ7TS11
yrZuuyyewNQOrUu9O/bDPtL439nFmjH7rDhnYhdQaHqGR94WiQXPTJ7px/FrBbW2
aHZGd8ZUODQJ7SC/jxidDtV/3jr/WhBKqfIwsWxEdLXQql/uSjeodBtLk9+XmV5C
RDM2hQAvup3gx5NuM+YFoLTwe8OXhC82TQT6uZfKG/p5TCcZ6t2ydUHRQa9vnLI6
3hw9QIUDK2WO5q11lznrq/2dL134/0KDrcQtcprwyOE0tbIsEYgwH30Y5QrsrhcS
HSJWXWQGxQnJyt12tjJrnoLv7T+sluijDIeUtDkFMqMtYSN/liTl6x78B7m0jS/Q
YIR8/1tbCSn+EDk5uItnuJCY13KYgfMidILULwzx8HCXI+u7e78N92VPZHpaYbop
wHLKKhgINlYnyIGI29btu0V6zt8W49w2bROxjsTp1/IbEcFnhYtvE7wUaGizC4pb
r31sc4UaVbJ40s0Fw6xOjpZhnAYYe6Eo7V+VO5iPMy0eoiVfhPxpeR/WgcCLya+6
HXT3m4HAdkhwJhd1Z4czWVYOfpdgZhyJcwA8GhGIfZutskHCG4KAVx8BElplMkMu
EN9WmJHq5IoMaAb300Zz1ueH8hefwxhGJnLzCYiGAver4Yak7oipxEcIJpq2w36d
w6+or7D5PKpEW2V2OiT2Bb+lPdVAOiNJtrnEfvnT8nEAOPQBLvG9lRcQ5LZW4pya
j4qh8cXFojUqujevxaL5xA3bK5rsxU4LBlj0v1xhe6bq74DBS2PA0UXvf5cyuqU+
jLBXdc7YVUxuL8aEEJDfHrE/DtCJJa+KOjvF9uA5Re8+99pc4PUdtvmP6D+dNSt/
Q2JU47IAeGmLiVNJzPP1n63AeE7eidgGV3KOTgQMpmFauJori/G27ioOry9cerXI
R+RMO6egeUp3fopUrYtTZ7piXHTJ9c2OsEMbw04UZSlfVGBvNU4vilBMSV1AwixF
4YcLDZN4kt3q07N5fcw2K8MfkvnQjTbSvycynrlOGoo6VVjvmP62GPXa3BKx1pem
X7O1J66wcUjbHXi30XZc8WTkLRZrZjWzH2G1OvOW6lhuZn0sCjQqJ8yFJgo1jLX6
YBwIlqg+V7gfeZ/ITqalVUKjyD4vfwEg1IayFw4WReJNoJDz0xKE6znNl+tYXvGI
NWtJycCPniMVZxehxytWk2W2rjrpoFytzOffo6j4PSLn9pnctzrfOAnkZBFW4z3N
Di0s/5ZSjCX41NysHypGfiJZH/mFEoGZKESM5d6KKO2vALZJL2aKsQgvFs09WoFJ
16dqAJ+x4Z0aehrY2Hz1wkdYVBxRoOz4eDg4eGWhzffjIKzXHaGnQhjxYHuab/co
7dB+iJQTrCOJPXJrEiLM9Q53vwOpQfRkFsDbgZP3WLyXfNsgyo2tF8jf1NfA0NZx
HZ80CCguVivlgUdbkB9IuZOmx9JxxyikeX0CHjBnEvhU7a34c/ptxjRIG72YYs/5
VaiC4OboztwmayZ/V1CCRR6iKXDVEYWp7xgmQfmWMHyxg5Hm9b98Ebie0QfdXDJJ
xGcusSAV1YsVKeRId8Hw9Z70PZJnP4QTerfgx8JzFhS4ExyU5evpVG9GMjc5/Q3I
5dLnd8fC1cdeUEFxRlnDnQDKdbvJXaJC9TYR0Q42VoVNZ1VG+gR1o9uP8HBLHJt4
Uyjd/ow6dQlSm0ncKSgMTiRqmZcpFF8Eo3Ei0QcTi4Wm+3ZqgFHJYyvHh6Ex19rY
UyjEVyc30xwbX03P+be4oPp8hmIIAw9hamWv1FU4nr+5Ea7yQ4WnqMRK54ueYPwh
vFLBeyt1eBdNceKlfJWBsCD7Kis518Br9hmuJaYlG025xw+KhCk4xXytG+f2Sfg0
EfLVoj/pJ1IuupnLFW77YvsIJ1iJ193djFzsQK0MLVUsQbMGHT4laXe2Kabf4wNT
yfX8cE7aWp98rB6VxTk3hoe9lhQ0F01Km3cHs/2nQM7QiAJ+/uJ89Os7ovP8i4Kw
/odM6qbUk+eFPsF9Zr1qydM8CcjIawLiSpzcB5F8l7I07Kj9hu7fGkt2XBeMpfB7
5jtXUudtqsXeuKNVDMcImG+ezONMULj+XpBMT9oiKdhw24YDSzQ8o3CAb44KP7DK
gZyUpOIFtlaI3vI5SSqoL7BkB4+CKlHfKrvbDqwI99p2Xj3MEmp57/DFJ6PSKK4j
Wy5aCPXr7Zli7NgCyNgJGt5DteycFqf57s1OFRt/Rf+lcjUrQtwy/1/v0t/V5v9A
mJ+KFnD+haYoEXvX8sGyXikLFFmvk+Xp6elFkNpWoldFGJeZfMNiUrZdPFuX7WhV
/ErbiEvlo9mGc5MV9JQBG1tt54wNNhcU+lRSJih5am0Fychw++W+VrqCd0yhx8sC
ZuKXYcIyxWam1+AkgUTBci19MQxBDIphEcZMJqknNtD5O2Pt7lufIgP9XbcxFP9M
8luJ9pRduVaiGIFcBS108rMM1f7HBjjW4hpAIV3XrmFZtpR8xurPwpWIhNrblNEG
/yAV3tVpRosrlMWeso4i3PlBHITUF64b4Jk7mf4Lve019DiBM9Od6c0p8UDoifu3
0VUBHQShM/U5wcX0uyEXHkFBIxJpCEfM2luW472BmF+WkILxtqgjGERrP/9LTsub
gOnDMvGX1bthPDtVSf6/IM7TtFpHLFtiP+E5bDOE1CQIXFeLSi4EaWgr977grXQb
k0huwsRqrTF9dauWzQSIfuv4dn+SlKbXYJIvoUglL6OIlcprzeabDPgPkOZ3YS4s
ekWqO/XsohsWk/Rn88MNElGOxaERBX/dUqVqasv9LTUk9n1VSVYmklgH7tLCb34o
mp2kzjX3VB4Q9UkTNbWP2qd9HMqi90TChXGs220Is8dXdbhqHlXm4IFAsEHGxk7s
1Bsv5mtC/2ObkyNPyXutoL9rPaIesL7tUU7Fg4+SJttCZETpnvZZ9LdxFLArPnFE
bxfyVB5XLULCTbM/JojMWO9n4JOZ1Xo+q4W/OJKDrdffbjaDgrQjZbCu2jzkrGIw
6WryCt2CM3ogix67Wi7VaA==
`protect END_PROTECTED
