`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
M9rxU8dB4whVbLSpcZDRH51T+SVHx3n1fddgYmt6EiQsrpYNaxz9rN/pxeNKL6N0
a3Sis9Ttj1tZIB4PRwFxzLq+1PWRMwoaQlui4Nj8F4WSRiwFKegw+IH3G2QJ023y
lhitlwwkZGKBRrG7X+rKZQhTLrlksj5GMUSJgRbzK8ngL7zht8bZZT6hWWcxbLpL
xcOREFq0DP4OFIgURRFlxYVTYb1TjGpJywyjGpRKLvdYSl+a6a3t0F2Hxas1Zy6f
SzfhJFbB42NZK+J4CKoe6iPtXlFN6gnDUCJXrl0KDwImOUm16ETXAxa0/kvwyf6n
6Pv8HaojMPGKgSztS8ZVHArmXErT8Sh5GrNWn7PqXxjgnzNQizXzxFjtJE1o06MZ
5vn2RolpqWX67irHcuUPVa50JkRwI67MHc8ct7D7mjZYo/0YL5+BVru8sgsv3XPR
wdF96Hm96U6tRGlxUKubZfPxrgy8RvljfpTmePXEZpN839k1eXqNtX9IF71TVGEo
8UjTQyN2Bnm2lMKLVeKshczoNK8BkPbWTuVAHuMuEeqyZORjUkTUPEANJwYOxFDV
FyYGo1+AYrV+SVt/i2Qq7D7RdPydLM9I7ik5lq98/uNTOVplOdYhfkoBw7ncgVFd
k6H197wd4fyMRtqXVsGkB2qU/y8bH/s8GTkHW/9tmIi5nA4NEbuxots8z98yIWv4
a2c6ZlaN81rS/bWWVl9iMQPkqjN8+8CCZj6BOer6mxSwoynPundl2wDLhMVmzr6e
7oWrKp239urvwi55Lv4ZhSnkEyB53DtNS9rsw05qrE7cV93ooX/xDH+DWMQB4+8S
uE+dE2nn3xkShH1o7CbzNj/sBOHs/u+IfKYrirBlUwdFIH4Iu6wIbhNZMIBPb8Ru
ESxnL902MiOPRveD3MT66FFvwhwjhIx7CVJxTpGD6ZoVIktSNmMxluwi4X44bUhd
P/qX7hi2ypCm5IFgJ85hC3W0NxRlgFKbJV6Dofncp1EQdnKJmeqsNFF2tSlGuUzv
qMqvmv/mEgz3EA1fFwUDhkCkZ04cEElhStxwQYJmGKJrrL+fFmIJo3NY1pmHWp5S
as4Ct1Btk4oZQQ1jMBuY5Q3Mb3CNExKryo7wRj7GW4oRvqia/LZMtp8FjdqQ0Y8V
oGm+W64nQR63+vbEY9aslVsr8onjLWx5dwlOYERmrrjCj5VJ7eVyypiQOBEKs2ae
xMcXx/Y0jExPusNF1fTnsMlmvXAMIVy8RSUkSdLgPOM5kgsW9Cr8AvaSt2QfnzU3
ffdUHLVqXIrdZK6vPArAbgir2Qh3YC29JHhz0Ye7h+CnFja0clMLgn6o6cAHBcxm
APjBGKSyT6BqDie5LIva5DzOYybvTLc6IWGvV3TtjPH24yrqmWdMGhpQnoPvpa9q
3H9LUYAP2wLtgkmOGRAyyPMvlP448XXEQWabIssXUXYaUTb/+F5fWljoIioEftWa
whXnam5hDZKWIBdd3CwV9zvIFsPdLNsUd+Q99EljaxOzXFIfIMGF3kGRmbzhvzAD
XJ8W3oBkTThcst4ZrrV0zGGxeg59GXzCN6xMbKzIpMOGaIj+0fNhjJE3cP4q3RYB
FJBLirFbzPMpmpOFOkYUK0btAoZUk6LDC34RbIFmGkg0oiok4Q0Ib77cGQULcpAc
LXZyt33G3Zuetwb5v4DM2J8zulLrbidCZOI36b/FWlqopRH6vjXNOSvhnjBV9Eyq
MkXHiyVD01OGyQ/6zddC76ROOuUevmFPpRfmPAvVUyll0ddGVNWrQjNUPX8oCNMx
IkIQUpudkle0Wy4rK24wIGa6ZiPT3MwTlNhMibkpsPw=
`protect END_PROTECTED
