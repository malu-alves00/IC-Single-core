`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
t+tHod14J3d2U8ivbHlPNPJDo/licgeHXjj4bK/bp+1gpQWIrRCj6Wb8QRacOI5V
hZuV+rF4J5OTPzAirhcgQ4iLH+yordoSV1sKeZ+8heYwM7OlHzf7ULI8lHQTuJdV
Egc1dtGX5Gr1Nzos0NbuVqbcJllfSDm15ryEaKt6FRUlkZYN4k83/Nevr/ytY/jz
NROXKaSAD5SgoM/0AKCOUNfdBEXwX90U4azGZXMkefAYb/E8evWW1KnZlhNCMRuP
ogB8MpJPMvmnHHDDIVxZ07mHEaeIhkJz+Y0dyAvd+VXsBWHlKs4pCTjP17/Rc6uU
HvM8dxqsMCIoO1uPO1NLRgrvZt6QotosgyIUAsW59FP26J3WdoDQkvzrKMKzPcLb
Yx1lNqbQfWkvPrgyPqurkUTO+7B0rdIZOK9u/CEJUeziWWEFzsJOp4jnXE/3i6oQ
gLLECstciYE3bBzhvEpTPlnVvCVlGCoaa420xKbNaexvTjty+ivY5hJAd0cJBFK1
NGtJWFa6KvtteOjziyLZ1hxFGr9P3GH1Z1ZsL9M3XfNXeeJb8Wbc6mNsUT1iD9LT
GSrYXoUuRdyPOt0s7SeGxVsfXHNZaIxLgBDvLpQCCa/MzpczN7vkcp7OvUoM5JnG
OiP1DZ1NX9iNT52/PNZ/DQHMtU1a/sDidv1M7EBTCQYiYaaSRFC5aEMuY3K2AiSm
OhoX2N5TxaYDnrb/+FVN7uB/BBPTMOIVITWWDQp3nZlLnrmotIWkCbIecDQzXdSM
T3xjYLTKdS4ryCwxGizezU1RwdkKrQf+QMAEj/Dd7dHgYLywHiIdadDXHsINjdik
8t/nrTw8i+4eXgAQrKEaUgARub/YqfWnT5LhPXSFaqtX7NzS8Gou4KWL0OZ2NLF5
d/x8nXWW9yhwbBdJZ76wCo5gxn+K71RmB0+0nr0QXMSWvueCX5eRtVSB/ya5R+/e
VANHXUyZuAS3ceHai+gd++93CQZUrrl+megDoTd3x7BNzQNU8FsjSJ6Xbt/H+mwh
n4IrPPqV4qyjCFgk29FM5fsio07eLZNPhi8lNVpbyWkuj219zV+o+EN4CDiexGAr
NAo2acidunX1yGNCN10nSIoa5/dhgeLGBqeCZooWiRScqonVcyiATgv1hLmOGjvf
afj7dbH3jEYIyCaTQW0M0r/L3ml+pi/RPcqyyhqbnEdNaibfIYG1tmfiCBzMW1rA
VZ9GXw6jT0xus5ccrAGTr+hEzMQZIWowmYQ8LvVPIQrFAD3jeMrSAGuC9foTryv/
zPe0zH1oQyjr/JJ0J2maNZFrl5yYT3fljT4l3GTfmBWQl0DW37qvK2dinTtlnDMm
3cC9Ob9RfRPkjXrvevPBYMYcMMjGprmwTZAeer9ru/lpkITY/6682JLHnuK9Aj7J
jUWHmNjXDx6SVu3wJBiWWcBQbfKv4jeatD++tqFeCShDbWFCG+QRz+lGPrFFllvt
OguGYZHWsPtNodJTrWwvxwQGpKESYojknb3xWo0MyCcZgq9CZ8sOCudxYDyo5aGO
3t9w9h0S0eJOwFWt21+sgyHdHKyA/nNDNzH4VVszINEjLElQ+ln5OdA90mAN3Q6B
7EzOWSE8IL6PciufqbQ7gX88EJZY+THmWk38tPmR0d/0pcBgof5p6PKBlWvrEFga
VVpAz4wEYXf/xWuxffN/sQ2ee/nS+EzenekPtullgQKJjmY3N86pcsg9buut+1oA
pHyN7JQmKVYkKdIqkuqJtFjlcdJ7pNo//cmQuzafON4znhNgHOSksHD2907auBcI
fPZKk4iuFhglKrvd8Qn3Mj5TK6cI6MUD3veqxhkZpVN0jtxLVAGKhISMj+Ij0Y3m
Wd9ZMql5KoW8L6zj7B4qRv/7os4y0Rrbd2gfp0nZLAru271Oap0aZjwDQAjQ2t+4
7/nX/293DJlzzH/mEKT2D4dg1Jt0Ytq1KHout4JZALrZilHm2DhF298zQUaOlJnq
2z4HLwCbbNT4cs/jQzMLLLMPdBNVntBkV+emyuYvof41nOoDdmLOtNEZnpqpr4bW
FhP0TdmYWPYWsCnAk1B4e3kDzUE/Ll8LZ/mOqKXeAR0gM/SIk9IzpiT9ZFJIwbnV
sr/eQB4+GSck/yStjc4DI0zCs4hprHFDJIyGYyygjPq9+cud1cxBkQ3bm0ZpbxJT
0dk/odblnSW8Iu4GNPOkvxfnBN/cpjBTvzmlHhpphQJS+tZkMcWSwdshoHAxGvTS
Za0QBLjYWPcFb+ohR4AwHv6XIV7ncEM+qjWMX5QbbLjSfsDVxP0r1KyDOIES9fBg
ZnFp0fiWfSkksIIGifYchAwa9/KGepSHPwIBObj/YL4rxoCs7JTB1m81aXDGb/Sg
urDVNDgUEtFbzpyDNsUuwpA99s/J7WNkaXEhMMFJ/BmL7uxBFC6GY/y8Jv2UhUpS
9sW3l/Y9+HPb/EjDt++eXUbciXgFHhN14ihE4B7EmzCMoiGGoznRC5C5m+Jol48Q
vb4AJf8UUuf2+7/xU+n7z2dKJIjTrRkrOd4XU8uXNEYeBG9cJKa7RbRCRvcGpZaE
RRK5O4x+GvEEMMRixpiwT/DWWIIW3IG3lR8fXUfhqwSDWzbRn5OxX2d4iQ8GFFFc
2T0/Y6IlggXx/gtsF1BQFxawUzcKHnkmLmNmWZu6Q3h4zbXtLFIqWzD3b3q5Wz65
A9+HWvlmu5c/bKZ1uSyIq20/uPFkNLXonbDT93p64bPQ3gPSOX7tY5v8MG8JpUCp
tGT7HxQVxrGSlX9DVI2/B/4AEQKe46i84S9EKcD3CUDnl9leq9BgvXGFPdFk9nok
0BZk2eDVpnKtE3tqU++TNrkbhQUsBpKj43JH6jgJqOyoLhTUpCs45opbXClEA8wi
bcfzSV72nTHjiyqz0dKqLVHRp5H8+PXzkB+Kq6OOp0mR0xhk3kHgrcghu74i8JgP
3/ml+JjbpIcXeK0Gj4HxcCwNSXkgGgKG/YZGe+fpZ8fJWe5Z139n+6VQQw4rHeer
XDYZ+DzrfOOM6kTnwoJxjRoGHpsmX+QhUgkcvTCkxvIKtPKplmjmVkXLOxuh68X5
w3p6+jZwf7COXmvbU9DotcZ/bmwci1my5o0yvq6XhgsEwRNDG8UO3bKzr9B4m2Pf
PvV7hYIMmZTxJgo5pjQ6+a9J4b9m1cJCTDhvNroiangK93txsef5J4MzbMJA/sb7
fmdrQeDpiPZFMhLi2DegY/4Lp0q8n2I/dnIUkiyxlGrT3lUyh2ioFaOqQCjP/Rhp
dDcfmod7B+/hjaVriTPAqzetBnoSyC4dSZoXIAyx9BDQAFsRSJeYEYBK528u+0so
kQaC/ab7L2Wynuh+W7BTt7pmFPxN+Q+MgBPmNcJzHguW0Ts451MQVOUHYsI6gDBY
SjCmV3fZfxXcj4lq8fShx4XJQxYsA8nFP6ueFCOq63b9KuIAHo9PZa+AE2RhhGr2
I3yVHV9fKFVqtW3y2jONYbwUfdXzrVUI3hDpVmvxZhKRzkyG7YJy5JxELWYKL32x
EvizNEa12PQ28cWV4Ex+KYI1r/W9Khfgv2FnVXaYYRT7TF4Rpwd9KCBcLHd+sN2P
0RkiJqKn7u7KUMhOoqVDJzHvNLkeucaGhaDn+C02+fMvHP3GvxbizpzKmYZKP4Xa
L2uS/QOXFHmpyYW4a6FtPKd50/6nersaNax50m4lX6j8fj26BfxAr58pN6jFrJvE
I7Z0L5hd0hiTr9v/zrnqBRcmh5/nwPOizfO5j6WwvVufb9ce3rYeOy8IhwZdRJ85
ECVMd5PA2wvyE55xsmN5Qss6otNF1tXRzqfvrkhPMTT4//8rIviLnwlq6xCtjU6i
XibmdNuBx83RCIH1RF8pBRQ6xhh1i1BfnYNiOmDRJQeVI1rCvFg4vBHwd9PMACKd
1RuABipTXCXbAGrkaBIhBWGJ/WJyzyu4whQPiQwNUtcMhwlP3KEd56HuKkyLTLEt
vhA3mR7aoUH5S3vZDrKbUZYHh2yEpD/B07mRLMwLk2RBHTiVnLlRMy+5LOpVFFWB
43TIY4Rnw/im1l08+4yaMik6ZL3mN4i9MR89rojxqK75HgctRYF9ZVxC85WDV0x6
hwBYO+Xlngv+7tUEl8STf0Rr5OjSZpT8mIn5AP9PlDz4hPlJe+M9xmn/WZghQkJn
EJhP/ZHG3+uyJoKph+EMN/d55+aCIGddkU9cjaL7+IREtSwDqTm8YXuzG7WHeI1z
rz5Px2eJBBAKTIUHVxRdwTa281KBB/ATM4wk7k/EDrKonGWXDniEKv0zn1QEAwqg
Tg61rO4zVvL/VMRACMSJwLQEfJsv+V3f99oYuRlk/X50oQXS/n7yD2kyvLk+UxH0
zeYeInGVypfCepIm1EpIQtcSds2pzPljWVRTDtXBacxdJtvyx7+k+PJCeZHQf/OB
fqaQGyEj0ujTw6GbTSPhdsDMLGQA64zu8XDCDoQ6X2HzudphRO4czROu1MhTh6Ra
Xi6UVZiM58yDPv//ELUah8FEtifsqRbNVZmLHslj/V+w0djet/q6R6FQbntLMvIP
h+RH0Ah9d5vL2RbHUR1bDjrTD1u4ybhYzieQifB41HZgIGTj31yj2fBW0SJewquy
of1N20YcJuhLS3QXFNbh6azzo9VAwTKxDWJLc9nBipFDCcLH4p9n1Lhup7M7k5hw
9lhq+PLvXe+ZXLnF1FC4R/cM9g4pAeHPRWMtRgigjB8vItndnFaWG+YM2+R8b5hf
eN5bCHV0kpSkoEnCkEL4GoOMGJ35Ec8G7+LDAF0R4lSDNqjzlOqhBPD27ZdABNbk
2p91T5Jer+K9iT1iNApUTcmhXkp/onK8CY0h7IMoVgQ5JTF0xKo9rujhInJ92OaC
SwUiS79AE774eCXImuNhaQ/N9PGYSHYNjxtpywhTXEffg/MpYKczi5tLdABAoU7S
gWOhB4bTtpM/JfDuf18VgJ9TwYLQa4Mhbo8aUT6f3BjOyVJWgowAcYTmyhBmM/ai
2N+FShNsGWvo+rcSSJS8bGQxVjLVhYryKunS6nkyQPEkxDa4rsiVQo9/EPTPpOxf
oyBUiXA9l9QVv3gu35/uZn6TKl93JAo1f7C1OyEjq1NTW1WfRbn1iUnXbzlYuME8
pBW+WW9Y5FpRUNjdmusMIITCrjuL4iKLfwKGxubFouFKfl56cX2ZHaP8MwWiO9vi
y8BLD6iuaCytYwK+kxKPkctiAJ5WhbQwCOKKDiH6OXBIfhFGMSjBaNwKOaoF2DAA
KKgoUG6wGSu6Ag9mVl5Y+N4NeInIzop6lG0TyrBeXFE0lyTO+SBcFJRYLLLVdxtu
/viHh+OL8kiYkXicTQAKGEOnkZDyeugxj/WcJjspXsa/CMogrTFe9c3LL5P8WIwJ
XqyrFhPmhtyUmGudfTO4Zt/nr7tabNTI1na96/WDS/seMXdGjXBYp5UikYuCqtbe
1NIzMQcyB2SIskhxa7QNu6LgHt1LdPSOuypW0kFS3ero7b27734rqBPxPciFE7XH
cWLCqqJcAPBosHobUtBNPjzaioRBctuiy2ayWt7UP06sspBiE0oUvDQxajXjTqb3
iQErzpjjiRXOxODl1f2avycgyTx8Oz06Zli1lPIVx6vuo9ujnBjkIgHbnbX+n4TH
N7zeCkQrqFa94lSIIKAf4yS4ZNpe6OPsT6TyxMYaPMSzKotkSLilWD89VtxgNvwZ
7pQihFpwmFDXSaKYaeEWVP4IC31+F8qAdYLc8SQVKC6AqojkPpio8aYhAok2Uyj+
ZN4RJyU7t/yUh92X/BuwwcGUohLaaqCvBKroy7fMqv5Ql0/ZPiCpk3OoexObyHOO
QKoKxNpRfecuLQj8nqW3APjbeFpJev9wacHdSL7WlgtpM04ipKIP2q+Px/8C2fI/
seKj75hMFhBSd1o6upEyqm5RxiOj9kMlqfruXMV0uIsRU8LjQkStKfRAnQMenwvt
qwSss8Xq4t45NMff19mQdj6w7IM88hVJU8T3J9LAk8zZjhxVadoe+MdWGrL8pL0a
8j4/hQQtnznyKuSpA64V/94zXvREDVaICRd7/RG3e6gTl+BV0IlPAkrokE9KHq6A
+DgKKK6ChHMlOhNoaWE4BNYMIhqXC2o8YCWH8354WVDcvsKJhOaHvWcqMRp6Zzpz
9knQgBy+d2BkHS3YQDiU3BtMPKllC+r+YZjBFz02Fyan5JHikscJ0walAH0Rhf9F
UmEWJ91QhZrdWRhDotP3fAbY67o4C1/AlBLvJbAkbCJTp/Xx1QbR9K4hZOkvPgCY
aK/hTiI7tnNNLVoZZuIbMN9R6VmaEiIWcjQ5GIzZKD6vJLhNiTv3IfHeJqT3HOl6
lE+0APHsVwmF+3vSX3Qy9+0pJjU5pKoXXc6pBDFrwRatP/pV2PLdgGf0C3y1JvIX
CNSUecB+tVEBhyrr0qomvvH3OB31MPh0dO0S5t23CBm52muDlComvMr0V2VlfVUP
JA4CFXkWIUVj7dDQBaXHShUOqqj731EZfmskkRaytfTifaEy15Rgjv631O1kllf7
0CQY8A3J1xJPs+KmG05Gf2Q/h7dVtgjaRMgoLZgy+MvMCBpR6h0kGd5wuHAGmzKZ
f3pu/78rnVTXjv3cislmQc4drNjfaaS/PIA9SGMpN52Dz73R0T2UyJRvqYkkiMPL
yoQbcid/5FNZOTGg3zyPAa+TTcE8yO113KH+ESsUAQF1qdHSKse1Zi8PB4WBfAOL
AdV7U/6yhJw6M4ghcbAfSO/tBvX8h3uHyYhQ9p86dOgYY8VNI/vPuqKeauxlxBt+
HRmStE/pZFQSXZI6XzWRHn7our0DTdCDTnjqDv0t+KlHmUX9xoHSDGcorB/Mz5MY
WOSpZpctkJJODbRkDShihmxfKkMgB6V1rcjs5rB5QT+sui9sbdynmeHKSBGiEkjw
wLrBPldQ5mxUq7rkXU9t9LCEzI5B4ByGV/Z6PLa2KoxfJXiIkdds6D8rYlq2012m
xSwqitO341u+JysSJ4DpYF2Y5fo6AH7QzvoJvkwbuwhXRfLWvvfB7Bv+N+ja1luu
ajTGWMHy9mg7On8a7MLL5DqRPEclQT2KYdDPGqVYxURoc09lYgE3m6Evhq/hKT2b
qAjm6iTTfN1BPWeWKg4z1/3TaEIEzwpJV3TOYGfoPyqHAUfseqiFiOqiFqsZ/9wC
IH2SHPsSuH2s3tDvS+wOc2UUPuuK/suJ3ukF1NNzvVjCLhglWsFejf1lowzuUmGC
BOKcn+e70RbK4Wtk2GZgVBjE/qFRX72SR7VuOlS1N8P+mJbenzsEmZCBs0rQ26dG
JCp+DsZ8EOF7Kd27WDASaakH07+bCQ3b3Iq2DXhDjN1/UnRzvDRKk8KLNfAw8KEM
iLZwzgzixP0XzjehbanEWdwP6njKbwXAnX3PlX5196tXLHdDRqrsXcivdTIkAMKY
wTaRRyZB4rE5tSP7Zzb1HE7LHtSIA8ENX1fuwmeNCbLlsSwakGLpQP+aegqjZD3T
vFZ69m1J07cScNmzdlG8grJhDcw78p+M1mE8FqlzgyTaMVq3Z/0jNzPxk5JEN8oE
3OEcILHkOGPriLdvrCDX4ACTvYtP1fWFWos5NEqDRKt+hCcYmL+S/YsynmTdHEVE
wx9VFecV5aXIRCwHC8LKRF15+b7q+UY2JQJgjxE4ZgWFpQQq+StVaHaUD8KDBaMV
f1a9U5C29MwPBtz1uT5V54QFzz1LWeBogR58UXzzMXrPp1MG9SJH7TBpXdrXnAIU
cUbduhEWVbo67tIBjONFEMKy5c5sG8IGveEg2QxZ/hRAdpU0FpuhQ6pwGOZV68lK
jBb3umDY4UIV4sn3xTVOX6MAFw1aIfW7tXxTbJ3y2uSo2wMAHGKoq5YgNg844Fzi
jKcfl2XJE5X3CZ318NQAfnADz4LREXS6I0j2VugPeca/pizCzwVU/En7A5ed1g17
8DMgDnTgs+woBP+eFySALg==
`protect END_PROTECTED
