`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VPIg5IFAc2ckn/IYLegsqUVcHrPN1+IO0uPDK9KvK4MANHJYkjBVGc8wn3jBLQ7R
qhYsakQt3XJ13JAAeMXxvxDbtdaZhCE22DexTvLWXxZwMSP/dwEj0doUbdD3xelB
YrycCSOWGW5AVWQvkWb9asYKxUPWNKWJAlixoCj6H1QnDYtiPDY74e7viDOmiDN5
CFJqkVMuPQukcrFcfNhEHtKVuaYldhC5kOvAE6G+X62p+wGWl36fcX5Eh7lXRUZh
m4ZuGV3vYrmHXiBXcJ17CHoch9B7EfxeCn4dOBAshEsJUnMQe0jXe00d6a8GRAPc
FQgsrsmAy+33MwdO0rSFccVrppC3sv2QGpclEijXrD0r9EwyZXknnNJC27iYihr+
rKlPnrg4maGTrZun//huka8P44TD38u2+dV0koNyDA6dfb+Qtdaxk1LLU7cdmEss
567nPH/3k22/DTvH+D9Y+yxUtXmjufRlk4nfE0bs4jLn5BkL43JBwBuNouw8OUIo
IZyhkHI0PZotqVIN6VYix2ee50eMchV1IiCSeFX/4Es2ZkD2QRcBBFJ62VYyMhB7
IYN9fU58ol9MTen0qjZC3rwu/QCOx1xGZpzTgs0FoA7X/btoCfjexjQhDQsRtaf0
ZRd5oAwkHg2jvzV+Hfru8S4Ydy0X2OWcSw8dejQ8cFqofTp5JVwI/JJaSbm/q4k2
3Q3BGyuovwpc+ZcjWUlhKN6QOUTSEQYgrIwMR9W0XI4BMnsz0Aqu3LtEilOWLDLn
1sYVrz7461e7+BHXQX42ebOV2MpuYZJJwERt5QI/VtW/tMLD8cM8jnOl7CHIevZT
GifE48+7geTTLUooJi/lhB+Iz1GnmZyGumv+xM3VGZxSAL2f5ukdLecgTukvUlk9
C7H+Ig/exL+OL6Rfs1kCKho9Hxs2X4xNcaMGpIxnc+0odQPZXK2XRYuDbYzVl4mE
wn3llX0N+dhZ7PlIz1IdwwqzppiI+3De134IqFc4LQphhe4UDlQG29v4Sq9pPh44
r2Pgrg8be0iZKQOWgP1CkMlnfaJ9oj27XUXutDlRfwafD84DkDnltSeNP9SE7khg
LTHAJ6ULCeqrQFUdXiDNJjtJEFo+Qr+MGXuypRoxazp6ejESToVqeu2eeWRnU53r
rcXveHfoR7Y1bDrERSXabeijb8Ns56AwOtmGmy7gfriaw9IsD2+KfBRu3YTGebWg
GAe6DSTR9jClmCDcsqmRk8WPjO1f91rtTtufyXLIMqGWQgu59F18RaIKBQ/tjYzZ
tEzuUxoQY81if6qYDjl4+GmHtPT19YZQ5tDxp2qSwEOlU0ojXZndRMipBT1aWrDS
vbGYcotekWiUesDKJ+J5zkRz2Jf2V8b3FQVg7bqr/sFt8goIkifh+pmArGc8DOrA
5ATuQkV8VFAMMz/jtw+J4agbju27Iy8IjQ5hESdNP/3IagaFtT/nmOKEd7517ZIN
vszAygH+9LwJSz6uggWGnBcAca6TlnwwVunnOUs7XnelkOVgkIc9S8wsVz5bcm6X
B5ilYfDe8aWL0myoZ3x6C8gasSNdTphhiN+b2NZtN8g+hkMqm+9AUwm8G0mr5o10
hPcmDmXqIaduDbV1hkuyoDTDdkdVy5IDhfXWFXL0OdJefAViLfOkJ9/IaJQ93GtL
eq/urVKVsqU63XWWyV9PULaZK1jMcMk/wr05uxep+f3TW54n0VxUqsk8haZu5JG9
+mXg5koaaHhgh1m19/wOqRWZiPHBEQre3pkkDrWgl1OAxfcdiQSnUq1DYTQrhznK
wYUfeNgU9lhcBXgcHli7+mT4Phv3FEcIlhAE7pLiWgWL7aOsEfS4pzcEdD7LtV/x
77KKzd137hRXl04Mjwh5GTdh4uur7OCK5GpqO5lCGd27U/7bUU9TNmdHO6B4JgHl
K6UYd6vt6zF9jltRAprH4ouH2FOe3nVB2JV2q5yfYlaIoPOFVc8sO+MKZZdQ1E8E
msS1LVAt5iTXb53FG/BKJhj70eTzoo1Hjp//5C9p8eTLkMmPSzyusv351oXGRQfI
v7hPniJW4kRj0ZFZesNwah/Gw56gr56vGZqURg0NiuqG48oj2bwlZhjPuDZnJnq3
GxjVvFxH5UgX0PV9LC0Xp75qvxnZ5w2SJKLEGsIuji7C3lI1SAukYvwoSjDwZkYg
g8ZEbhNhlNKHP0Cy5vbqBTc8nrJXDuJkGcgS61aRYbd1I/LA2v4ZG/ZISX7LQpUm
CXCQV+xKNaqmFsihXNppvsjjiu85qHHrpcbcLmpfmmmilgFtZauT+JVVof008UnY
wRvT9BJwcL1bqrp1icFWVesd8Bno5k6rgyvrZm5CDZ5JZ4Dll2SmmJO11xCXDPry
tGz0n5MPZv3lQbBXY7LmSCYghC1dU2LK70XO5w/c4TkE3qzWAmtzurYWCNeW/Qa+
OTwx1tYgiTvjxoL3wzf1IR3MhrBP1SQ+3okZRZu9q2WV0VJDJL/r26D07e9Er9mM
EbWQFjAVMS6Gd0oOVc5Vg+TNCfz0YnUjKtq4j357U9W6L+AA8nnmytvRk2mDmbim
zXSRPzwHhrMrntlhbaxowIEofvLNFUpsj59x27Hu4JmBqnsA4t0xHUZRyOtzXd+I
nOwyG+uikCkF/JK7p6PsfVVDN1xFXppZj7otUYCamMAKVBCgnlWnFhjhXyoXYL4j
VhUUrQa8OWdaqniPirp43bYmNI4W7ri70hNi7PDiXMnCOOOAEivyxxJAD+Jd0TFd
MaaEAO7ZoeOVLhnI9inZwJQ14/jd2aFmYCvwsQjSsIuUJ7BW66CofTDyVGbuuFHx
6N/YcZXCOcYMkVeS1aPCaud8bxGnDdL5aDqGB9wJynRV/z4VDu0CGUsB7sVby1jK
2e05rN0EjZR75fQ0UYE7aJHp0SnBz06Ahb7jiFyaQ316aI1J7fchTwN/V4f9SCzp
Kfrg2KDPcPmTqFSS4F7DeH2VqOQ7RPUodivMRyg401f6irP3oa4Zk4lJCfhS6fDV
p4DjeyLTbGRPN3QqEKF6kiVI5U60rLjHrksK+oqwDAs3Od9z6PtlCQaP2E01vK2w
1XlPh02qAF+knxJCcfT/BqE6Qs2ODgRAgfQg20FnnjZzrr8VzNwVyfGdsEotEpuD
TLTm2lHFWwb2mJZfDWeEl8y/MZpUGeCqsg1YHv8oWNzVDhIOv1Dd/TEhCPEdpXoH
wexN2A961/+jvrmhG07cmtn5aI6I8Wv9jRO09dPS7IleG5BIcQOQeeugmqGchDSt
bdevNa6kh641KgBZaRVj6ftKZKHqYmH0aDQJAr19twSR+zBKLllDsumofCbk5HG7
TbYEggqB5S6covk9MPdKkNi5rjsjxTFIID2cQ1hBR4Czd5LTyfTnyARL4WkjbMba
IE/wMpyObgZTanoWX1M64oecUi2fp8PVLX1uuSeqpBw0OAYuzAJRT3ijCGuF6F9U
8OrRlsC15OR9Pbre2KZHP9PWKR9UzR7sUOO0qHGbn/uTWWdugyk5F9TBir5BFPF0
nI1X58oLhKwDHwITkaGd1FguAACNVhCHPb3vyVO0Z4K/4kTX9aYSlxdLqAt5+ogq
cflSwu5gISB/OTwhxZOeIx+lsWK8Opf1J4WOrzTvkuZYvpgCK+qN39yfRhvuKXBv
i+7sSD20mU2EUflxEoAoDpVgTlWLEUcErShQFrZBcIyMZw/hRbv2vtNTV8TM42Fy
hfl8cXEm/wWEepxb/C621cOF2bq7tCCXK9gIOPVfYcbdsxb4suNCyiosSObGbWr1
Nj/9mlbooiQ09fP5qUHz3VXvwPuDsqO7RnIEv9ktXUNeWvLq4Y7r+QCCGcqKhyjp
dWdmUcOk1PufqPpsx37Bz8c5DkG1V1EEUIMdzTUmtACEx4GOxLR7cvgPUwQO1mIh
buGKoDXpgAhnYeHulC8WWKPyx1aR1mMnLZrg6BdigD/PXR5vEHmdlVx3oGazf1fY
U2EF7izsxHdfBga2C5WQs9C8wFFvSExF+kA7j69dnAnfXtMvJRFNLNcQapdUw4ZT
kmflTgH74X16ZJkPkn+SD+gVrMbLzNE+p8Vqiz9i20VFERqAO+b8DdpnSQ5xKQSH
N3eW1Tm+JqQ4ga6KVpep5uwCjkxP5gkR6MghIbEus3vGui5ChRsQKjf4eVH8RRQW
73xrWrBHj7eFsSPNhXN0sFIzphk0D3CEvWSxZqeu/XgmpxH7AruKjC23vrPeZlnM
dfcYbH3nP58lhSH8OOaFPsaOHgzO26ysJZnZsovQ1LEtPhT05bSl+g9JQT1VVt8o
zZE7dqzMJGj+aNb6LvgFbAsGDlrPKrwQ4h6sx7ewXlR5m0GX/kve3zxxKHxDXq4s
TbxR0sHtNx9C29QjeTUyLEuTUfdLhcd0K8konTTUaqckxJ/cfuv4DwykLnzooA9M
FkdBwH49yrPkXPO+modHY8Qn9GDgTPJA1/+xMm/EI/HBzmYaycg+G6WDcQvJK3hc
c88gu21hwzhJnnxOZ13d9s3mqj6DMeQpWIYpMh4OBPw0QM+xoQj4rRb5CzQCwR3m
/04ZDXS91bd+5AMka6PR5TNFwMqOrvFyZBF/Jh4K4Fpazy0usUphxhB7Hwvv7R09
acyA05olGkCW1P4EvIMsbox7zuiwMyPjNAKacIn0+k+Z95wkObLcHbkBiNXgAJyy
Nka1gZpaYkXzUAxAeWq+I5J6j33VtBzWiqgR1YcG5e2CJAowS7TEDl9+PQmKb9iW
IWZzm04dOrWzfELxngSet/HPwrxMCIVmlMK6RJ1EnZHWOEZc5lD17liXhvlbaqsa
jtGVQXEUMHMakVJIPzIFLYWF9dX0eVeNAFNLKO5xqoODEyLzx8ZfRafPEJwM2lEg
7Ie6Aklpw/YPHb6cAK3PLW9FtET/DpRJVfQGVKJYG9rcYeRIH7WH8fhhg7T7WVgU
5bBuNnxwCuxPuuNBGgl+XiPXiy+C7SIu2CCR0ElHxwnIXdezTFY1BrYDaI/LiWPX
2aQQtpV/Sr9/2wYRlpSGUrMb0J2ca5r+WMO+cdap+nvnHY7oUPFkP8i+O375nRhb
AOTZWA+DRfAKjv5e3tFZfJKCJhJKLel/ISu5tkxBu5YvMcXNj/2Cv2pYOC0dJYyM
G5cnhZ07aojEtyZiy1LfFhmfc4+5tmEMyTcre13gzz7sZp0w0Dt5MkEdvcAEoK7g
978r71pQGJdnhaoMbnNx1rJxvx8lv62jKKMI6FdkzxIhchEA65jmjdMhwM5qFOEm
lUGAkxfVmybxoAkBkDIMegrdUhqsGzeG8YA6mbTfwu5lrSslm8yGcGtzHYiftlNh
SzNJVjGrbnJVLay+FbHsDlmFaZLFUYsvr7UaKdZfnJCItR8KvQhlAJwBgSRNes1Y
5Ot+zHXZgAx1z+xVtDAmwu0Mtw6tj07cXX9iIJg+j/9wU8/FDXTw7lZv+pbgtz0t
aonbxSPNxsSgOUPsJdPE13XbOSPmSUtFFPu+rZ+rpjIClxVgsly/4i3BuV/NZ/Qp
9ooN2ZE5y0NVilApA7D6RQez3gd9pJWs9a3D6U38m9QnXwYyPFko7dXb0YyOJSbq
8dinSuQ1WyVxCIrK/ZM3cTD3ueCezkY2dpGlWDRu/lKCI87AIsS/Hlrnj5BkLFFe
ZNI1ZPpOvzmaAEEkclWtPETkHT8/S5c6uCTIkDon9Fe3cSk1ifH6O0BJ+9/zqs0r
wez0YpTeZNb98ZzZwnHPbhk6fpo191HFn89F15FOBqBzmL41XrteoaOGUOB4ncLd
s+F+Z1ZKdYpVwxc3i+I1eA8g4zah/+fGl8VrAD5ZOzs40Q0AWJ6+Jbb/mULDH8sR
x8jPGG1WwzlgWfX/4AEbj4y5yCiJBVnnnMuv2qUnf8WCZtwC9Uy+JRdLfnybXBlV
i+9ZsqcWzsHEjNCpaS69UUiu2rYM8V/nBso8KpZ6nNB4d0JKDsgmePggFaBjk3gr
04zyrgsV5PSMEkOSCjpOFi3BYpPHIzjz4OZ2ZznyVV2QAxtjt3gU8tzvfCOp5WCm
k0O7kYnbYdraW6e8iPLkekUuGTcmEl9ztxeDaZf1FXy4NW6jKQs3hP/toIfxba+K
MSkuZ7XSM3QBAlBLUxu60qQEUgxcjaQwRSM8QfLv4Z2Rh8E5kc1DkP8eeUn6rYSX
L7uiu3tDOj4WBYVv5cuKilLMDyR1xMbhD9cE9wjogTjDvOl0YiCPAutOS/Mu/D50
8Ys9yImegNg6pBm2WEtZ2Et5/hxbXvArCLRuWQ9IDIHHSWI9Zwti/ZD1dabnC9vv
rtxIxxUzcgrE5wvRFl19PoDK9fDQihC/FQ+jd9segxlWQhtw1D6Qoxk+ACWbD6Yq
KADByN/tkJlIQP7/Y0BYigGo+DxIrrYg9R7zy9w0fR4K6394Y3k8DQtHdwpbd6qj
str/e4rLn98qeWC/IzQVAlNGOwLDvefIfxTSM+vMf3Tn5uDX9/LNvEbIY2XOvges
1yW+hq18dRWQ/i5LExMnhAZMj96mSNcoZNA+hK4RgoiKrwxQwVLEF7ObDGt0xDas
84RXLyhsFrjoRUTDGnNBcc0V4OdyS16dumnEQdGCF5V5FNyFkYNIbAzY3xq2qf9O
tvgXdYRutdSDium+f336i1pD7JV8fUV15ukHctGZGFiRqM27xagZ7p8xWlYG4FVR
sZMcGEdZBCPl5XuEYMgaTo22Lh88X7uUvkDV8WIUKcsmgQqyKVXVE6rMn07EYzC3
vho25YoG7iSXK9RSu9svunJusVXBJ9dI1fVFcmZUu+9F0efftmdgPGXsb9E+Wl9o
ms/5T8m15mwvBUIGxijx738s7AGsEmgUYa58zHjTqSmT4GlkGO1Sm3jTe6rx3Ifl
KWpjQiwO4ex0Nivy7GADj7TeG6SNf0KSWW29TBJVsDWAxS1UOsB8KNZbpMOW8/5+
+YoEJ/TchKB19+2iNuw7Msk7fws19k7GvTwnofDQ+9JRntGovhpyBBpW652R1jIw
/AljP25Whp6RerUwjvcWjD4xpCXSP6U61zFv+Eopo7PlKslLRHgm6U3y+oCjzMbk
8M5M9JHnq1uxQTECvR2pcWd7JASFmtDCvXoQSye9wzjeN5eZQaKy6t3thgWs6qZi
MqYR5Z5JhsnQZTcF1Drf9umXkaMslnGMrp+t2z+HbbJUNhZdv91ZPqP/iyh0HepP
HFQeGKMbobBoRbaOOy5HpFcWzILBF01vGKC8XGR06jPfrtnNenNRim0LPcRYDeSp
+hnzyQfj47n8N0r3gJTw2UWlXz5jtQFZi5FFGoNM3iSDsr9/vY8mGzw8FAkBxzBe
1J0MFheJ5fKCnpm/E4p0hC/vQlJemlMlACDthR7b9LEh8B9GFXiY9QJBZYcRnvmE
SfK8IG0X6gdFV7/8K6JZDrDmrTzOwLa8wBfss2mC1P6nMDqoBsQ1kVVZ13LZfLhT
ozzM2mW0baM/5KOUxpPcPVpnxStxRYudoNZU0e9f1TKxaP1wHlilCPupvjO4Qip+
jV7pP6Tkaa6WbTMxeM47TEh4k2RYr6gykZ9i05JTduSrP4OsIeOr9dhIZBwj93yB
+AKCntTPlLficaYpJgCU6NzYd4tP7xAlupRtEu8juNZxPX8eQ4Z1S9TtoPc3ar6W
418uCyfMnwpdtzo1ImN5FxqaKYVQUKGeQdzAt0Yg/V0HjLMd7dYiVn9Zi/IkMyFp
7Ee9SA2okR99kBQwcxST/h2v4uIP759Aydkc7vX0TXkQVX2BcASgovj+OXlkKlx1
taKLv6uKptdXPQTmzJWkGtAjJbDp0iiSYdqdmZrZlPhZ4pe5FBEk609cwZVQUqx8
6UsuNqwlkSZmDtirNzOCZCkMHeATl/g8M3iqa4GkjzidoR/wUAW3WM9zGY4Bvpsd
VWEdezn8FsZmc8d4GpZxCFmhbcstTIN0KChIST2QNjz53HbmdGgU/8HA9DY4Lt+f
jAJc9NYwyFwFcpfP/hPTTV/2cz8nh9IcFOlRVLXJmPkJC4xy9IuNDeYCZoFNraKx
hAYREawFPRflIXAmNs2R6SK1WIdFeEhojpNBYvl0rH3bOwtRr/Dzu0/QRwh16xRP
vk+BuNgv5o9nHwX1ePRHCVKvzdBiUl5X3w3VqMjr+iKHNiKmieITCGiAltTtBPGh
MwPZm8Nje+1e71EnvZsy/d8DJ7ovp5bNEFYppV078MWTQ6t8pW0DFjQYW7KlgTk+
PqUkRJJN7cQmF/iC4yARHd/EAszQcFrinCa5VGBRb5o=
`protect END_PROTECTED
