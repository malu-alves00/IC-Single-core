`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qFnL/1RQcP5iMFvIGPlFgcS7rZFx8rZYJ4oneQ1kiXBrGAboXjIgDcPO8NcMnbZc
XU1Dejhtt8wo/kn4gI0EsSgm8XkMRmSTK1GVIqVDuhWP6oS7hI0hFcA6CyWebFpH
xRk+AC09300tC/98FPcWL+w9yul72FT2yzpfzsHy0OUWaw31N7a5LW7OwOdeM6ll
0NE/Fmv9vlGG9XEL9CLAw4vKr4lUX8TnMbBQLKab8xd7+IVPg7x1nWXWdMdvCiJb
RsHAmIyBr96T3EKDwOYTbHgkOHb9rEUInyn2eIwCdWAATIPrOGziGFcCppJmkUVX
Ge2htaib9YZxSwv7ja7eRnrIld0rN4ehXShdDardl8QAVQ+/450spbJi0IL2EIdQ
U8aR8J3z47VMKrGTM2duYlCxQS8dnmSk9Y/9+eTUUDOdVNj5DGJRmwCjoHW6wAl5
bR3emD2nHTxN9HRdrVCiQDKWILeuxyR3c3Xo+/hcR5PMshrbx7c+p3150j/fgVWL
Cdqw0pV42IqrQF8IVGVcKzuhE70JzkmTdPP7++C8m3IgcRVw1vmLN67WOjmLmVsY
eAKKipQZB023tad0pDbbnrOXIBdJ+1yPeCiymdoD6SQwQUPqqRbmPVq3o+qtvSUS
8rhzSB3lOoTtrG8061zoj2o8Ksf0U1+PysYxdg/cxkVc4YLjd0PJvFb8SYsaWe6/
fJjW0/30RxrmxBiDluOLcu1mhIZB2kuIIAQm8L+cEJ7SG0PIKec+8NMZsisT2P2u
mq7tf8cO0FbLZXFFyYlIaH2euVqP5LKvAK9IRcR4IqnTykTtFxrtjNz/EckpK3zw
lJyzx62YkvHSqVVn3GjbiT6R6gwChYnPfEoNPWQGXseemiK9+2cMBl/Gm36gt2fz
VbpY6eptXUU+6I1bO4lBJCoJP7QJtog0s+j9XYUiw0qMQXHBHB/bglgkWxlJOQ6b
4oZ+aVHbMl9UyB8S2+J8oVuphJWqDdxSgSnPgo0jLRx0rfldsvOgVDJYY7RQizAv
ULXgoiq7UdhIwNMTFFi2cn61DrIKx+I2Lai//IThyZKKSFxd42Is4guvFISkOnRt
YhP6KKHVbBEfg2f4epCRZ09QEhy7Bv8P32YglqUfA+9a505bo56VXXcy4/y/aRlm
jVoGe3TK3gnW0DFbubdQnMXhlPYFttNYDjzK5EKaGZQwS+FHk2CLUFnMO0fvzEEn
krhy2V2LoVgjX7Hd3fC6g8pN20tVOy9nL8eYDwGSN+FJw3gGgih0JQBu8ohBAnHL
3fS7MXt6Wcjiqy+LAoiA2xd3DqvGV9Rel1jCO4BX790oA/FVOGWQTyeZNLo9Tbyn
SInaMlQCcVoNx0Dm8KSY0A==
`protect END_PROTECTED
