`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dDfuPAhynZtK6IEbZ6abNUKZ7hfvje98hduZLV9JiXUo7e6Gm4toCOhUF3Jg6/am
MDnGAevMPsQ43KL+KP38mlCGiP2oczOVLm7PWhA1RdjksAxOfQ47xrXkw1ueUPYB
HYnBSgHastG2V3X4E4jaIFFJSi2wV4UtGEWw42wo/evgDzkSkJVspMkzaLa9Ljt6
Rw1lkOySrCUAPLq5K0AZEJj1KR/m47pSTLrIVY+ZpbSUm24X2AKzYmREnPagiGJ4
14JdgDlxXPbEQ76pyPa8xHz5nDqKzZOIgsTZKuN0K621FbLSs7EImDw68aTFQnRY
hXrHfhvWtBIvoYILcB4MGvVOcpBq/iTTv+sCnCKwsOHgdqRosKqNYSIUfSn5TyD/
zafhbmP+x6wkreQxyUo1j6V9KGgto9USizSSA9NfeaiTx3AgrCAQ/QQvMXst47dV
6yYNL07UNZsJ4OWdFEQhFNzxre2Rf1h2RJZsmQoaW/GbX72TsPfBC9SD+r+kUWb2
u1tBin/57cEZIX4Ss7Fs4a98FVWDfNp7dVyVSOp94zH6AtPglp2PeUMfZm6/AfiA
j7CNlmBRoQ1uR39hH9JYBC73UqL2knJDhKU8prg3ib6QgdmGgZtSX6ECB9XSllnT
EmXqCpu8mqi/vheUAd/HBiZIqYgjLnaVcoW4nHj+gGdfb/O/DixtnUq5PLoViHzY
Q7iVU7dcmulbqgIauD9FBpSxR2qGeWpRGHqZ63BfmiceJr6JBf7grjvCHJGk1vT7
BojzTgafgUVx3qCjycxPJn3RzKzP1xqd7/Cd0w74rwtHNU9s/XrbEDDH1I2xZQce
YtVfkjb8/Ra0ngiBKLROrHONdv4QklyxPwQV1vCxCwTxuhFLsHg6Q8JW+j5156wY
/yBR14eJ9IZoftRHYLh/zwjdaDmnhqAnuiVxHVcUh2wcjUaCiucwrRud+LDH/Bxb
wrl+q62aFAs11o010BVNwT6n+3IlGx7tFy1RfjTkly4IMwUUnoGnOVO8SoctH+ax
zA+TNY4B9Lj+3xcmNJH+4o/ggx6VSIqbvRlDc75kzSIr5jDTt6rczos4pb9bm1Ig
WKQrrWq7AHrJUnsHO9ovR94EEL+3Cm9D3ELZrs0vzogXPv4saFW6Q/ItgwzGFj6O
KZOke93eFdavX8t7RnSjCo3sqGtobn3BFEri0Q4PnOGojxQSqfRP6hYFp1vBz40K
4mEuKml1m2Tw8WOr0eX5QzfcV1/dX+wksWwGykI0eZJSxnM4s5QScAd1k6NDgVFF
VD2CJuKL4pd/XRpb0lxc7fLc2JFcxs4kn0iQ5O6gs30X+TjcFM16NPb195RdzaNi
EekOTdG7M/vviuMBX2McDqfBI+xGHxaJRPKZfc4a2DbpA5EU77lM7h2Yx682hINq
6yB8jffsvIL0e8fzS4mhbD44Qiwv5MquiMdjFwvbQn1aqTmxLIt+71/sBX6Kz7A9
VtCohz9TqTI9PECf/WSWUSwpexFnEhM/dRUiYGA5GoLuJrPnQ3qaJXYbCKoqliYO
0YL5W5UPf8xU5VnP+Hwiy490hCR6vM+g8U87MLk6TytVcr7j7gvbRiG8l06gj6e2
39em7BoHBnNRypxLWHb422hFxh2ASAH3wdQscMQKGwtXTJrLMiohlfyzXrFYE/0a
T5HvVA3k3VBU5GUQIBRBLXuTZt0VPFLZh7Fcs4Z3AkgmY5CgwJqJlqwB0OoUS32s
KWK7KgnD0gZvXsZt5ZCwnu+9Ataz5uAUtRCfTzYqyOwk/uofK07mWPm+uM8k7pGQ
rtxR0Mvg7ID5FGuvvnZQsT8mXmGvzcDmhzS6EpFhOrsVcogDVuGff2LPC/ljJQVz
BLv8w/ImNnMjK0E8DoI3yTM4YkTaIzCZ71IKGn61MByWNc4h8oz5JSvlSfuq6cq3
3PjLDsJPXM2WctcKBGROKU2rUX33mYgKsgFcNB43Pqw5wxJ0jxDXuBsMyur1tQkA
DS+/dPHFEKPy5XcN4gvWWH+Ys+hw06g+UFWRvaC++OHNF3JYgvH5+Ou5mqZlY23z
+gU1Azi0RZfPvsneXY9IhUMnwsGTRKpcV4sMlU8T2wnwVhDCxQ10LEl1PYjHOlgu
RqWxzC5lFN8x6r4eA8Usvv205Vuxto967tJAwVlhR4fnOdYpeNf1lNPOUr3zZRzW
TOdYYosv1UfMSRqbikXa47mtWnZXKvTMe+ErvalhqPENAU+BheEZARdO7iFx0MFp
u1y/LLW+W9HwlINS2Cb/t/ccLSDObd9UblI4pOfOw6F1DO1Px2KJxeEIcEXHaW1W
y9xvEL/aWa1HCQaNDRVamMf8c4rt9ic65dRKMmDwSj+B3JWcNV9LkXyL3hG8hIm+
3e5U67EePO6wLsOmz17C8PF5FEAy5yWx/Z6fi3nO4FojOq+8/uCVRZ6mNZ2cp7dH
YrYGr+2c+Si5tC5frfg3RmLs08VFopR1dQDFVewIXM/vrZdWQg9QWUyETN3SLkXX
95HmeDGqbhZS1V1bi0p1kdpBmBjDUeRBuSNmr3BbDLV0KFIxaBAhQ4jbMGxptLOx
lLZNYJL526/KZvtFGk2yHg==
`protect END_PROTECTED
