`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
owOrIQW/dnP+jDG7EYhQbZYU76zUUmPzzfmST4rHjFCcZO9xYXocRZVaOggpAzej
z5zxo9/xwClrkdSZe4wz/4bTn4H3xVNi2RSdma2bJ8MO5UBdCCn1ORtqaKm/aMCR
nAR/23qg1rOkRujXiUYWvN050IswbuYEW5Ex0kIeqaIRreWLnf91FW759VDTx47m
R6MgAxqp865lbIZxFe/r31T/uPEGwiK2j2zyBuyTH0onViXE9supsOPyOqBEs6TO
pkfHIXQDKWrMWxDHwRD1ZvIZ58La2fg7NWGJRqbOuKN3W7t/V1c5bMcA58h3tobl
2MXfUrC+8NUWPjjUfoXpaTGVx+XOGZWUtjv5EVj//9GXg/2W7OImEtxJIdjZ1/U7
mhl3EremARuUHrLXXORjZ7LrKKmRsbDzkV1jtJpwXBG7SfSnCYsfWNJpkCohe70K
cutKhBvekv1PZ/7qk2It22ukmUf7/mKOqknhxuI5zBt9hkoBNhFvbAClIOucghpD
hvrEcn3G+jdlIkrWCIQj2gO2+mHPoCzFvhKTv37ss28md5nio1uA95H0H3MQzuWw
KwKRF/+dKb7RHRiEI/sKZxjD+GitlxqdVpBSNUTTXy0=
`protect END_PROTECTED
