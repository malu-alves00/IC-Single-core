`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xkFJxd5UfN/vNxictn8uffldaD9tokofVMdEr+dbbF99kbnp9LtwMngv20FKFd+j
91h43Vqt5Hc27SuBO1+dItaVDqkm4bn7Mx5YLqy0iFA5rIlG2dnaP72hYzpxCO33
xqs27z9wpkQSepawswHGz5guSsm0T4c1fZ70kaOKqkJi4RpQDeTAzwNdS2po+Fc6
ARzMIm3nlo6nox7XD4P1RUCv8HsgnW73eGZ9msSM1RaNjKBVB/QrIjV3BYmkpsZk
TciHNyE6T7KHyLUMAkMBQW46ZGGhMZIqu67hG+6XPPoNQB8i+KJhoKuCYtADxMQ7
0CGORLpGPh03Gm81fRblbt3LJ9+HwPWj5w0H+BeM387tPYEJR2ZEfNDXyfHc/I6K
yuxDudFG25NVYVjjcj/CQQO8Dfe70E1M0sv49yoWQc/vKi8EvRiyk+CSE1CIQcMJ
Jq3Do3KU0H++FBtr7o1X4j/DItQQaCem+oVSjGXsifv9OU74M8Nj0GmvEW7oRaYq
pDNIaAMMpEXWovbotc8l9Mg4ohT1RYhZwxRJdzyk4KcT+lJ+NmqK0nIIRX/JSUJy
hAMdJCQYkgaOHBxDnCXWMRlmE/x7uqcUJe7jO1Y0Ff2ATO/XjEDt7rNxVFqCWB01
sI96jAfLbA2nncXD0do/B6J2/EE0a/jE2zuwo4lFBs3nsQWBT3KGQGhOiNiA/7aA
r6zaOihMIPALCWcAf8eneTxXpt3qZNwB4nRscShG83laGZbuqXAsbBUKcTYkTyAr
ku5GurzVHNWFi1MfUeJh6enhNXIOpY6TvoW4k5EHAjUG6sCjHS8frCoh5NQE9Nen
Yg93vrH7EzY9dHsqCWA+uarOmGbRrlZMJayv8g02Ce0oEWRsfzOt7FmIU200aaha
1YrXScyWlYbP/2/g2CsJUYOmg5cHE0MibMndv+rUcbByS0kcp4hht2OtBooYi3MA
uNAgR47d9WoXcKaWJtOLaoGlO1cqOJlgFk9o6WtKqu39te4qSNn5BjzGOhw+3K6s
V6NUPmSRdv9GDHvlk1GlGKXNs25yphvkNBDmmkfk2Vpl/A7k9doSwFOmSHsYRymi
dbfsyQberVDeaRnXsMOotSr+MHJVxo4FHReSgqmMNhzSukr1YhTA9tk7HhL/yNYr
/qaliJINnerWlDfawRPDhCMXDaYIyPwQtJwaKVAkiot0t9SydMOdKzfii4PauODT
CG/ojTNRczdB6ePO/gqbzvTOkQgz6HN9dTWrcKucB0wIumBRNSkLuf1HRUV/Tn48
2wB6qjrcgSHkDm0VXkhpVdmUuTMJsWdaRUGFUJIvrFvZA/Cq5LG2s5UuUY6xQmdj
6cKRMqXE6WnTqKMEED4cikDYgCP3zi8unDeuHw/vyj7pFOY7oOoCpIV9MlqvC1Zi
`protect END_PROTECTED
