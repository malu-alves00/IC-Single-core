`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6xoWm9Z8e5U8Mh0TSP1A2aT1893cDmz8JmrPy2wI+0MqGYS/luVzkyhHPqLJWQ09
AVdFQA92uw4vlJYU9cRAWB+sHTTm1Bj9O0pnqXngvNejozJhuHIdn4I3Mew5g7zq
Ys6sNN2qz42e2FCdTeSnz6AjKEFqIKKw5rG22IXdqGuZxxfWgWWH4PGUFFDdkWJL
egujvIc/XtNG1jY7Jw7X8lihyYGbGCvfiCjhrv4hMMpenNvBL6PY/T6vsMda8Poc
t/wpEn/UQntHuxtTa1smqu9Yht3XrhaZ2hmCYIMtfTLiRnUdRmdKejt6eCoo0GlP
0qehR1CaLO/mIiwlBrgIVgSu1MWFPSgfjuiWglcvKLABw2rwq8JLWP7b6NnnAQGQ
PtbQ/BbnuAatELfeZKVJ2Tut/bpSqDq2nxZiSpH+7uBagNoM2QVovgo1M8Rd3FQ3
ntL64RrHq2S5JoFS9ndj8xqYCOmTRRqX2q+zV6H+ozwKU3ETZH9TvDPXxbM+zVVI
c+3tYhiNeLVJokw4KT9zNVg3movB8m04OM+lpQH3q6RESCKKj/DscrRbx2OIzb7f
RiEpd2obMNZyOyXLtCDyqxk9YYE9YREt32K3extTPw91dYfQrzonRJvl+xN4Wjct
GbI30rV6xkoPDuUhYLs9SpUFlTC/wOn1xldEibUlXSFi7pozgO0XRTz144cWEQbE
HjHYvAlKiTaQaCEdidE7eITX/PW1nd2G3olgDT2sZl3uWnIpC8XgTdnzPpVhuOC8
jH7G5PPD33DCcP/ER+25nqFQGYnhylBQfto+VNhQ1XOSYun9J1ESAeMLTvOZn431
KJHANhJQEuI3BQUgH0dEApvbYs07KOux2rYrIFPELGUuMzjQAYCEi/gCKN7/uGpq
SU0cO96zGnCAu6peK3g6FKCc1MxMu7YxF64oa2EBvFESO+mMFbwUlQiWbPz4y36N
SjefWGvkdNv7aBAf/c8hDjePtCwu6fZZGQr+bnmQvqp6JY9jLc3mLenX9317tPwH
dxN+M6cmFxO19Dqt/IsAzykmTIGreKn9ID81ZCv8aLUp8fOzPRe5UKgU8WUIac3K
3js/e/llJrzsykr9vHH9MTuZQfDawwGAdX21BqovkM+Wy7SMx90xlLDBbN0Qpf5d
F1swzSzMnfT0EIG7k0Jg1QVgRnNFk25Q6n5t1Y0HA1ggVp2LgcMoAE0Z6XCWFhFa
tnNcVmrvkUDhqq/wO9QuWW123EaBRFZHAPKqv2xa6p+9jo5UYpmnBjPltzL4dNUU
tnIr2yUNfls8SpQSoiWiAxEe6dNRAxqAaRQZr5eHDZ85k2nLW8uBOcDK5q7+7XD6
HBkq0MvwBBwmD5rBrI7e8iFDCS8WvKe7qDxU6xKBy2TEzuo1ZepnjDq7Ovb4+CUc
6osrRVyavD/TmRLnLnHm2PINyQu/k0zNQpxNgHI6o8VQlZlpWrliqwEQoSxw3xfe
Wscd1J/f2H2DPegqLpSwigCMfq4FoeNDnufeh5Idsz5XJ0NQVByBn0h2wv3n5EKQ
CnvNK2kUvYnZLVdoa/ScGMUXKuB4CMrZC0nU8ZqDFPpKvwx7hf6mq/bd9ay1TllN
XGiyxsNkbNEilvV+d+p9dOXZQ6kq01uv9IQqZabvWv8DYEJWZsOs8QTH1SgoKEXN
gUSsQdSQVGUoIBC5qi7ATmwcAdtZ5E3vGwg9/h+qpD2pY25Z7Y9mnoCC0Ry1cSre
ZNi9Bx4yp+IizI1Aj9hyhtEn/c9xPm+pPQcHb9WP29Cejyl7qJOTxnJsSfigPVUG
uLB0G7d3etbTqap8f+abu38jAZqAQjE5fjD1H+q2+tFctr51hw0RAXej/EvCyDZG
m2NBKTjpwrsUBE6ECAOFLrpq9wVWs5YpNPlH+48WVHnuZ8sSMzGMntbhKhjGZ7Rn
LdxVPp5AS84zQyNmu4Jv3crqHDMg44vvUoux8GyUP15Z1EDqqGViZv4kTccbrzkQ
le+VuLzGiNFFwgTDkJI3wF0kIiptgoBOa18vC+0fAYUllWqehUOVq12TvOPRXLew
ZbZOndvP/W6Xx/c5CBboIdc+WIzYcW1zoQBfi/Lrv1mKGLMmcROvWxnz12HOa0OS
PizPexcBcdkwbWpWnVw7SKCYkKdChk8/1OnuGxHUcUY0gPNfWQ4esSzjT/AmtxsG
fLUnaJa7p5JvwC3KerV1ehFgPNWNu/3LqiPxEgOwurFjnWIUBU/3voZDEBcpZ562
me+8yN48/2aXtJUZdrkVmf3NyT5MGgZXeLL9XCjN7xERdllb6D2H8L7L1VVHPSZP
QgHsANR5wgWMu5iZhQ1z5g8snKJTPt1zuu5P5quPCY7uAkIg1wirM+K8HQ61iiWo
9xlBMv/2BB+0EgxMotVQhOV7SjADeDG+6Z6B1SffKzjbUf+96ZS9wqYLqBVE5g16
pytbjeJOFqNReq/otT/4D28CAaIJJ7wUzGtftnVajXV5V+O1S/g9gsq5Ru8tKOO4
eR2zdJw8QB0P1XSSUjXV6FsDpuzL/rofP9deaAUFcPDX4Zq0WamNVpb9teq9RtR+
Nvm3Kl0eYtngnubnOYZoZCNvupc0V9bU6canOqV20fJYQZavldwc8MIf9BJ50/B2
84Ay00WrCUNIT2pTV/UAldrXc+iJe3XAQd3XBMjZUoC3WdZb2eZAn6sjvV7SBbuK
q/YkcFBOEVLjhCr5UJFFUa1rXVLXxWsKwgYoJ+exqdMgxx/9h6CsZyC5CoY+2Rrs
NuYE+cHo6/pmqB0X9GY0eSEPAOgG3NbQNyMSuxnHy97tVloo1dm6lNCMyTVyawf3
Yssk1UUmc+Z0+UFjYdNlVcyFaYUYe0Ku4Rz53VklVNZ+RnITDyg0GlAXS2LDtS7y
vb2qMxS/VSFdS/Zof0iUJf5TGHZnmLAQvumXycCFUb2uDQBFUXZjEqVcnEfckEgQ
4pBZSYS0nzluVbPgFtqs6qIVU3Qr3CZvW3ZTVi2ZHuPa9bOS0kY/FYjMT3SiMHMj
2qf8/64Y54Yd6f2P6USo8Ljw/jenDvK/ZJ3o4X/5ftRUf879YDZc7KVX0ulhqovW
3Lh7izVu5q/IGL/ewSHpMp5N7RZGP7habWWR7W1cwe1Jib57gOVnFv26z8KDqdNy
hXbRpbuZb9232h3c0fw3Pv4GaBNSTrNsZEmJJdP+nefYvH7fmNCvFAnZW+ehyCO/
upeybLHGFpXa7GLKpVSAC3FwL6EnGy76IUGebvEJHSBjiJ1KZxLHHV+rmtLvfmsA
1FhrdSA9tNiw1BbaNOcfCZnvynVCtHVgD+fMSCJptcJ0ufCD2NnehCscYsHI9Bif
qARuwEKhijVxTFnbsOKgeRU7H5s8G6DyTQ3bAiwWq/UidoPm0d/ma4qpsBTJAKLD
NEOWmXFcc9KB1OWjAsHeizEN2yn1ykNTB16g4AI1AK7x1omRV/fhw+tTcuxmi+hf
yOvsnkeAGDttswm0c2iKF2RmJtq+4cXmkBdsvpbUScBcWTmT9WUfis4wVrU2zShw
jytmrBuP4J6jshhu4PRbWyZQHlHubPGu4FIerOA1Nh+4XVOprjwRM55UKh0LR//I
kJpcE+dZXjMMy9QiTs34iDCe2XDYI1G1hpceyU9HxMxMYWxoHkjVAF7sINnulUFI
GZCIZhWX2qyhs6SK5gKNgxvfkA6dJe+SCpGIgmkLExXb5K0csBspIhBdnMnMCM5x
V0PZ7FeQJdSKEhxtOZ+DP97Z5Y7ZfbTRGuvQdlIMIVNLyCKlUJtOd9m3PGypizPy
IdMJBPbFVxElUxgxE5qm0dQ7scT4k8kw6x6NrPVgsq4FYdHYGK+dnrPtsCfcFSm7
0630KDYqMdX2qFOcGceosiBKHFNvZBD2fHGsWK+03WU0wUoPBTEoX4N2fHXnITdK
gDszKI1psXORkgWx2HFhgFBoCv/Y5PdA57CIB0p0xEVuMa0ihw10oZa269DrgIyT
dPGwOoFjsPkjqN+HdRwOigu5rD9UdpFCM3MTtSiRFwCh5gi/HQqJ7RRD4z9lomic
xOrTfRLYhlmPj8KCy4IZ+AjiXoXnPbcyHXaEB9MxWSasnyC7JfCEueW5tgZCjdHY
8/tKWSftPj2NWGvuGd8KNpI70k0s1yOGXNKYSmslOLn3bheLFlK4A1waQLYLoMSQ
nutL+IQNt1j4VgCgwBNtcuZ19CmmPORnPF7JL38UlEE2MjHDusjpPKgseWbJnduR
qQHBPDwZmsyBVGUbzpZsfRTunj51DKxO7aDFRVVspGFLlisQcjpc1oPByQ2lhntQ
pvsMje3c5BUDYreCmSvIFflS3UOoELIgaISP1qooPHh7n9Kee5XMNh0XkdtxpctW
bChjBCMraUXSsowQGKFgelA4jF87u7PQ8+EvgkQjjqJpv+QBzJtMWu+5kHLzE2Uo
zP+DR/cNHkqHBoruAyzallPXd77wwlN6vWrrn8Y+A6pxVRFKbVr3SjB1KKUOIvnY
i2fd61/4bYq40BZdCLLv2uTQbpkTeQH9JzepADnJSObhShS3fbK/uplvqUe3tRwt
bVcZHgoYQwTLYqVhPY4uReI83ra3bgpLnTeiE4elPRbgpqAjNFjDVECyleHFqohX
nAXg+GyHuUfaNpXmdz8IIfyNkgUF1JWt2Mhzu0byKQTIUj1CPGjbR8ncPhrBPyRc
mwiaJFZQy4+YlPvzvYm4BmAOneoLEokL1Sa9k9hSIxrbDjpvUNvzEANSnAcCZRyQ
vCnA6YpuSzvC7Ir1rhA8Ddn/Sn3LcF5zNYCPNZhuviX9nbOAVm37I+Qj0lgiCyRS
w5kwwr+FZqLvZHkdUL7Q9UXbXQrxU597xg/BhLWh6ASqvuJzIgODdX1qtr/Ee4lg
bSWrDyFChrLCVgufyM7JyH4kuENxlpdL+aJc0vZe9Za3iRDFSkIrl4sL17I11RhA
55tAnCWOEEL0xzGtN/cZPn7OeOZ71HaMwurN3iNVz++HUOTaFuD1nmrG7oLL17SE
Rv/HlILVtvXEoSF3RiIxMaqLSEngeyFOy79hJO/njAKGtG7X8o95JFL3lzpNOCHt
YI0WGRgYocKhzc4/2Y3cJMKQZ5XxhYhuPm+gGSRTIwlXWYdWhKAGlUglbNVALSbz
pLlbhQ7H4hv3QEnmRrzHrljxf+aD0HTRyU6XFB6j41SxTfZy3Tn11o4EKo9F3Gzm
YD4p8WDB6eZ5I+0ENAdAOVEOWhagRloNWI39rRXAwYQRANeDrrVAaaGaSfl/3D3R
AuJEYft9wqPOPqKKGJqqDim+HU3R+GSPgsLLVS5bgcLOinenFBG774d2eX8icB7C
YKV5MDyItNhKHDrxKox3swnhR0/JXLSYwU7wknWvbYcc+HbKWuOC9lcKdtSbHLFo
KY7EOvOJY7Nl3MU7EzUDBC0AFVw5lWKlxKlemuwnvR2+JU1Cdu9oxBjDCKl5EPGP
UaPUSYV07/xVz7QXrLRr1DvfZFXCdT3zCKKuSjcNbF1b+zv/zBkGi0yOvhgcKrk4
UAlPyP1N/lw02aBunfgkx1Js5skY8FiPHX98KopklaQ56lmjkKWp7zkaf5M+vO62
NpZyARtV3/f0muzusphH7ISuLeAthrwBCALMNeEj3/0euCgcbw4tS/+ffpRHU7pk
3wK7iZViVQZSnur/3p8jzkxXzUnDF43Q+h2Dkt7e8QJV4/lix4P5hrmFTPyjUAXz
1r2T0eNttEHOJqgwBvg8ZoPLE+UpDTBrPJAyCtpMvL7S5vTlJqwkqQbbX7LbL4Od
7Qqb56CLQS5xIOU7Q7jqrtVW2yZ6fmF+68z+Q0xcbJU9SGAfxufbLhJUMhICRrXd
+SEBpeyZ3ZZ5fRsaq00MU+zLMDwcM2o1+0VYGQYnUYWS/ewl4DjnlLY1HwmqRX7d
kmeoOkQu0pA01Qqs+bQ4IhgItkzS5cJwz7qDOQNXqY81DuN1WI5OgC1TpESjlN/h
lrWX8/jTO0EsiQAvYZimjO1iFXkH6Nd3JuD7FXdw3BZrlddHWOneOyzZoVJpbYUm
kDbmTcE1MnwCPZHQKFQ4J9Rn8Q6ixZUK7I7RIq0yxDPELNg8+Hba4bCK8JMbEFGC
4KJlgIrn5wPamaV2CE5rm4HEw1i0a4cHN8OlRw7gSc+igCGgWUoRM1JPpFH+We2+
Y91QaVGEhvUDRGB1ueJNyi1zigGV4qBkiEYhU4WkPFHd6z56B/UOtwVb2FMYX3tz
34+zHvndZ6v8yn2qvKCQovtBypgpnfnIqP5eEBI4cHQUw+Ym2Toe93SbKdlAixbm
bh9rrmPOe9xgwQR1tV1YYlRQXXx11XJjmXEsGTVoRgc3NoIdkzTL5F7OjI79E/2T
5aqPB18oiN0YMhItgah5e6wIHqosrV5s50/MRZbZuhRoCajVbkcxLfSwUTcbJjLU
/sraZN3FCex8U/l4BNuETbc2iZUlBTzH0giGyrgsMoEPtgZXgzzPbcDynZXLzSyI
U3YNZQMbD0ciSsuq5X1X3oiIRveZ5PjJwus17C9Ndud3y8/Kr1Zg4yVsY42yGO03
QT3tfLQ4j1lp2niKsk3VS5MQlE2jQ1xViejMoeTFIDx3JDEWH03R0ji4AGyD0CG5
qvCgvqIAMkCxP8MG+OXrjWRSbpel2UGXUxUgiQGf337q2fHxBTaLrx40Izcvn4bH
Os4t52RfVPuxcZS+2ffgf9Me+uYTFh+nN8VEkSFggII1YND6ASqpRrwOl0AhmifY
CzAlaqQi66M1PYKWtnNa881ArhphxtGL6xxSfpUDmy2okjowxGNvzZ0ACn8fo4sB
5NThW4Paxpviv6D4YDr409QgTdXaTBiXAR39P+IvAch9K3CEbixXdyQM8AbeSil5
WACPlXCCCeIITpY1pQyo6PhIwRrSLYcYZ2hUGvWhNHWvBojsJUpOtJ26a6ORv6ic
yXGswfq1Z5knfCBN5OYaXGS3AgfPn1LFyxMoQdvjvqIJZSbevksa50HQ9xX6GA7F
aDYxE1Zyo2aj1PpSyFZolsWz8IIXevPtYRJJr6R8rzgDK89tKI2M2MlemdyqS0Sr
7FBlgVzLk+Toqfzisxw/dpd55FCI6QhOMuMJB140KydqbGb4MgJKT81I7QrVLJLY
PhfH/fV7GOATY+TNkf9avhKQ6xgVgtzPjn2Mt8cMKLzn8rzrDfX5fJ/obH40rWkU
y5laXXq4cp7SnsFXlveNc2d87xHy3CuG+mVdbGBL8e61aIncbRFNGTPMe1GOxfSK
TMilFDbx1UXFXwmWdVyT/gPn9WM4knI8VtcfL3KixAw4B2bOtvHIKQFh7mM4xmm8
aDXV62TWMEV6Bvu35tHwe581gsJAV3Fd50W5shfa/jO416D4Gveof0FitlZAmNoa
FHOJ6Os38J+the1OCu73Sd1Yul1Z4cRmRDW45MDUA7ti6vCtoMmtBUEDPenpQxpp
Y8zezbgFdJ29j2gVelIVn8sJLjcwytt9Vj+AZ0epz1Ocg9b0fNDwrS8iB5QQPo7P
RbhPcwQaEIu2Q9G1kDX2L8Ci5syj1ENmd3KML3UiwbwzJk1nQ5ND7v+PhPX5E6+r
hnW2SU3ABJUqprXLqTSJ+/lCwGMsHmV8fECkwDrQ1HsHcfpF4TZy+8dNng4slPcB
SrqmgAlGClEWRNCVODSVYR/RwnwU2evTdgHbRS0yXJdGuJ2o0f18sAqJ0kRHI6i4
3UQd0EFvCxYgceidh2TzqwJR2B0+mJprR2MaSMLo3d/CB+muuE6DFHQQWF3bgdHS
PRMvNzQ00LRzdsVgl4U0dnFgEtm0Vd2CabsrcZfn0rg=
`protect END_PROTECTED
