`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bzwIfn0TL7rf607YDcGd0MU/2bqpKcS7VDEK/SiV5k3LDZquopHtSRI+pokTn866
0NW8LS+0+Vpp0hm8SxsESy06QRi10SoluBlNwQ+Fj6F9nPUQlETa66KZXYYtJ9tY
KN7kV80bfFu/U8W7rS7BFCwqVo88xK/WC/DuBBYgnJTKk6Ac5XTvd1quuSt0ZDI8
6KywvccNubB7M3iJBUJAPsJXH9v/oDLTqCb/5U3Q/wR2qpVcIseYHddGOfWkySvw
bZO2+lmSwGAQTYZUyF2wBqH4VZPfblNE+LIRPrDVmHwX5/oLawfdyaTbC5kFrE5e
Ws9EuRk0BI1qYvgxrd94J/Det4uW4klp5/5j5xohTH+BUDp+8Zkg29pgr+BtC5Lm
ctG/HHOY0aSu6FkePo2RcN9xNpMlwbaWCZL1FqaBvHXVToFx2eNbIWsURapgZnp7
jIDn9FEEuLh43tOS+lT9hLuo10+4sD+YfbxivkU+1GmamRmxKz0gzeQ4wPHMKuU/
6cQTglv1146mQKYjbhGCK610BK6gzbGNlRaKCf8q13nj3JI+hPU/Zr7kazAGK0dF
jocwMOqMBiL3fyCt4VwnPA==
`protect END_PROTECTED
