`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nxS0eBLyKAnrJSmxkaiVXN7YAvwQqflaRPqt1oVQsN3KHAlTKwRNJwDOYP7Av0da
ZO5BOzJ3d4snL548Ul+WbThi/0xwdzpXQSNgTArHpcLy6I1Agn+hlPlaguOv+Wjv
s3P1HhS5RJZZS1+13+ha4ojB48ODST5hixUetGQ6QjQ0VEznYBd2/KqKCmhMjTdG
+E0O2ZD85p+VNI+rop5gCtj0P0JC0sdtr9PO39BWFmDHVgdxk4Cfh1BRIDSmfGZc
dyj0BAvej8WQDuNW7WwwpVeqKQEo7oadosfWd2dvx4WWWwMZn+GN5qk14O0twFY0
dazM3/N10fW5Inl197yDY/Pn3xepIT5dp+t0zwJPUlkzKFzGqdOOxLj2mTskMMPr
ISr3zEjYXMd173J5BmujYoJ8f3pn3bOf/HZKt/K3hDT3twFBjUkKODE02RPfXLCl
QWiLbv5gDG6n5SNT3BufA4mNS7NJVDSefqKYAaYLrZ28h+t6D3b711lO8tWdcjQT
Sy4/XaAsZWQcqO3Mx2IOkobDXbvjvMVGwpwTTiCIUNKZwfhwnsGdAufH8Uj7WIxm
ZXJJ0O0uqelq6TvxKPii+mlJZw9EAeyGgAP1TkAwB2FDT4ykJ/WNI7Yx1BtEpddE
hER2mMDgVRhapgqCYKjTwwJPvVuN2qzPJUbTR9oLhMxLjmXfs+tO7CBlF5DCwTPR
447QBCuqhZMcyoSCym37MpHSqwGwrX8BG1milvmVYPESUxcOY4IGC0u77IYlk7JQ
4CdAm+e3QUOehP0PQn0zKg==
`protect END_PROTECTED
