`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lATAVD4EJHhctrY2QN2d4Mb+GeWEDywPKJYR8924yRQSe57HS0ytzwMhNH1b+Bcx
sOexswKJBjttRQZtZTqru4HSrrnKLGwrjzvAjp+jqlw6L7VeGA2jrwMEAabXm/0l
3c2CrvouU9oCnFWsdRrENcIzphJzvoFT8ABSvRQwtiS2kb7EAQWcLSlZaOx/euwh
JkZt1y80z3pBysFhH85SX8b8WQh8IPSeOxzzrkmPjvvnDePPbYw1gAW3ScsTmwP6
KQcjAdNaWh8HXJ9FK/uSaj293koT107QtE8tdlVjL2YAskXFn4uzQhPfqzepUhza
XR9orxTC5hHe1Ky9+spHhcswGxo/CKDscMJF909AWRS3oEWkUIfNeK8VhtyZ0vxy
ZPx+3js9RrUuYizABBlZ0qNyy0G3rqcOxjhSpROQhaUB+YqRlMnuwFEoeanK96eq
zBSz95F7+ef2vsQcx+T6TEQeg7ePHkdkNDTPYkyX4JMHhcd+ZGhWDX8Nt12eyeki
GPi+DPGpBn7NwnyZTtN+zUE+Q1WFOFRcsQHUghmAgY1UCPdjDOOvFGwsHYbYnSgI
oGmE6pzK/XDHQHqV9jWWNDkwDsWMXNs1nS/b38GMkpMG4GZvvjSbfSYPK0u0FFyX
IsuNwwwk/cqIC0PHgVrc5ISOFltxV7WLZE/+rKvjE5l7cLJCTgUwM904sH5X89Nn
`protect END_PROTECTED
