`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qdQEh/eduh0m2GhJuS4p+A+aWQWd1YeMnVxN7XDqbAq0GtbgESHd+Z4ZW84hwGmv
Fu9oA9OsFwbo9//ULjIxwLI22hAgwCYYjYKjaeL7O2kZZ718PW0WWGSlOR2LpILI
FtckTuTZG3NUZRhCeDASwwIJtx50IJ8md0gDxdFzNJjN/4KtUFkgR5pYTE3RvEIt
zhtAY0gKNL91cmt71c7g8UYLCzPmayH3wReA6AZF/RE+fUxpN9weHvMWZw03DzbU
diEgdBrf2wMMg5aQCGKMJpce92MQHW+wOII+VwaigS+8XOraNvklJ5c9WX/g9ity
mnJPWX8N04mEedN6SevAbU9kIHH/rgduFHRD35EuAAeLwRWKFDVgvpFNPVTusU/K
4LCxrRj1lz1jCqBcPqSitVF4oSpVc/ELwvIUlEhKAcqTqwP/8dL+rk7rkjzxjRVe
vB9WogryftWPhQ34sya/pICdFtK3t23zW2U4Oy86s1Pe7jL2JpPeU0TDqET5RRqi
b2r8vv8GtOkkR82X5PJlsVz8EFcancbY9kp8vPN/Qs9urpDbn3q7yYZja6aQ5+0a
AJA2crZmJV/r/SYMCdggwPd1PcYdCH2nhScnoOh7Gg8cRBd+0z2Reb7pw+aodY1n
UO4XWudT1bbjzT4R/Z/skH+l/W4bDIyyc9Z78LImn/TQXznahirj8T3A5Pes7hcG
k9Xd5o5ueo+aOoerTc2sxo72oTyShwa7yB96UpOOLjEkPTeVD49TxSmIKwcgbIUT
XU7BHJ7U1edmKURm0jmljpnbE5lf60uN/OarXyv+lHDBh9VBxE5l2dSPyg+wwrvW
hx9PaKAKS1yzxMJOXhxaI83WzHjicCO1E8/NlOa0Trs1AaMK7ShPDTGTwShdj5Z2
BCWEUO7/wrVju2xDlSQJbfwPw/81PEQpnajhEQB4WX4lXIXb0syc/IiQKYukM1LF
jIi8m2zfsHOi4FKzII+d7VzJRgVuZMeue6HI9A8sBZBcDI6pU9b7d8eB05Xy3Fyl
h0GO0c7tHUeOc5mfOumrmkri/khahlbEdjwf+SLxblaUuNL7q/5kOXWDCxXZwKk1
NiesokinsE6CpsaiOk3iFX/1DRiY+sPu0aVl/STRtuNlJch3H3IHXQ3BQ9zmM2Ea
TvfKulSuCUQKQlF0tsG4LJ7b/PACQoJ1WD2PdBgKLodg1PbS71vPxNuMftmWQrVW
67warU1bwqtG3vqpVTCMUBgDxWMDNfCb5vSXjbGzcF8=
`protect END_PROTECTED
