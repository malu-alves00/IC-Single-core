`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sNqgaeZ7NiNNauY8J9uW5lBYNtag8Rfq+2A2IY/HP738U7ALVGTyafIrIM9XBGS5
jIZKhmdzLv3ZnNE75VNG+LKQgBVtypBWeEyqEY3ksyWyOqzqqeuBhg/Hbsh0BM4N
tnWtM5zeGLZlukooE7pHTWmCtMkJiImxTZhI40EluTKdzNBSy6do/THbdSCpFuUD
fLeYxGE8P/uGNXtSldSePIZXNi6JSWgWiRDKorFUp//kuT/n5X7rm9j88sRRNw3Z
CGxBFWG6PkuOx8Yw/qNjAHEMYY4LYGUkbBO8MVt+aq964FPxYqUqxeZDWmh9Efhi
OGHhYM/BF3kKDF10oMM/pnBjjqv9nTKs8mAB/mKZXFz4v5OXOaPQTne3kIzlJaeh
GnS1cCtVULyZGW/4NlfS0SDtgkzADc/x81d0fXS7XtEvxi7sQ8Mz0VRclolXVC07
dPQAN9nVFU6kvjQ4Pmjj6Piz0s04GZzsxA33mT/WEpzLsXm16ibIz509J0UXGV4x
7l3KXguYgPm3ZCYUgBFReOILkAMhT3oUgqc/9XpcgJbUiHcUo4x/55Z2tMGm1LxD
CZ66+7uVKbgIer0YWee8I83bCh2LZ6LKl8HKaqjrh5G7TxIMcpE7oK9/iuH3y7By
RqUN4BvlpKp0xdINugwkCgE6mg+NkT6y0w+b1VecmKsvP/vqqTxHgZF3kkBZlpPc
if5XdeDkPZNAvSykFbcAZ0LYzMjZBpXVT9aKzD+FRuShGGuHSdP005FHSGVP3JAE
P2OZCID9snjQTHy/p00uf3AB3Rw+tb4cshiW8gXO01OGmIUja95usohVgrNt2rQK
CeVqn3WSvRO8itZQ4swRZnzB9z9nxhiSXCRo8aqTWfFgippnCY6wTQr5ap/iACxn
vC3GxgiV6z2Mr6zmNk39jQyr/pH+e/2mJT8J7qZzmNf7epdjiLfhW2LEFSkpoqBX
mAQPJwZIZGRTOX46C8x+feZn62pbf5tYzixxRnpeROY4k1sEMG65D9KiP9MM0gFm
gsfBCpYUyYEjmEP5gBkdl9vJMZVFGCkRDB9Qe5+1fHP5dZ/ID5iolg6IxuXkf8h6
Lyv6b/ydaIZYCUoql/tJbQo4gEt0gzfMKIrz7FFmjMXtCSukrAyRZh0EjKu8FUfo
jbCTOsDW1h5Fqetzx5pmKsH09kfIPzJgAd4KvN1W0Hm0XnJMto+2ABfng2BwlHNJ
+gk3SZCxa9fPAl+mvNTcCBEYPCL/VVLaottJDkCRjAIZswKH0/cVrsVv2hZAmlRX
KD/jjhM55OE5Zxj8q/A069W+6ECb78fuZyfsvykpdXzlCeJvE8LTiB3y3dE5kSUX
eqW9zMUjldIKRTuZZX8m/RbyEk6QRPcKPHN2pwATXaHyNS6bsTVTPGyJ7AKVcHQV
5v1DjOljW1F/dBBaqLMHRrECDAxj88UnaKvOYkZhSYhqnHeLZJCNUQS8qf3OECAp
lKCbJcEeoo/xkIsvvdMVgA==
`protect END_PROTECTED
