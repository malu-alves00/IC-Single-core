`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
glRLOCiZC4gzw5x14RTrIh/dvMUFA/UR8wQ36+sa3uzPmS1VxK4TeZAwgapYKyBJ
aeMHvWV6W3r2A/8pC5tMtOoXMMR2wIxw3stiAMbux8O8wchSFT6Kc0de62Jc7i1q
fr2CPFHgC33Ha/CvMyJua0BYmqhoK9p62sjNmXBIhVNqytgI05VCKVgJKt6Xxvsw
UFt+yzSNvb8LYIWDND0yR2p+y9ptI8yGgrcSuyJ0L+/NZwT3B4nQStICqcb+vpv1
UzbdK4cwUpKSFLqAQVJ9ZrNWB1t0GwGmp1Y0mqBY3NLHjZ+dtx3e1HdlOSILtkcx
S9G2gghNTv03PiXr7dUMVf070c4AlNksilj4pIpn+8wQxUHB9Jo2L+Cr9GLOLgGN
wXzUPOQVUNMc3ldyn9FwJmdH4p86QyTZOfdmUYxQo+vGsvKXzhnx86TkDCq5Q8Ea
2puG2QdRJADQGoEgXPK/fIGJkcqV66zy/edBL5vaHMUu+cIvbW4+IdcwExZ5Jp2C
FA0EQRP/w313q1DrIqfdx6ss24aM6jQ7n3a/+x6Wuqc=
`protect END_PROTECTED
