`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rSpuaajs3DnUzi2pHFdAWC81SILnPanV8SozztvEi8RZOCYqrCKwYkh68haPQ93n
D44881O2Kok0FZ8JDZtfUeWupELKD8ZghJKPlPTLmZd4E715dbETem9V3xpJgLih
8ci+Q1J2q4Q1AwZkPCnx220uJPjMxQv5gsUadQ9QPVNlz8zYGYBlFezNSW7czO3s
fXMtS0CMmcHo2UYz94LyLMdrKjCqnNwR/Kyog3frEgypw7P5gil+Fdv5a5BmjEJ3
2RqCIYkVggzrXTZCabiWbTe/HENQR9o2jD9S3EA8baKH/YScDi+V59nmSwSdAhO1
Io2s/7MlqE6WRmg1wpLS61KOoVJ4tS9F5tMr30Ycdk0=
`protect END_PROTECTED
