`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
M1ds11eaOHEzrY048+Pa5bZrus4INW9cDaiH1Kip8WiNUPxN7DlBxOXSzLpadGos
+5aMDwhqf8hu5vnwNIGwBwLcHKq+8D60AeuaY/9cPK/64UPBws4nPUz+S349vSm6
zyykWK2nn8as5SSYJ2PyWjoKsKBSSJdLdh662/sq7vrFwvyagF0ExpSETjDHqM6R
n8mWSe/WW5a3/Y029J0UhNMYutJCk7gBrZPWK2lYBJ9u9kVOowOm7WYkWCydalqO
HEmiewFM/kcMv4O9+LuvEWkXmsBzzFxadzP3enoxxvq3G8qEYVGTYHVRwFaO5lGe
GtVpUADuNNEozKeupOCxxOTKryzEhUr5D7XWZZmCJpayLyAxSY/ql0C+HEVAoUK5
exWwj8zqVkV+Gv9IvF+bz2yrv7CAu+8x4MDZhiJwThGcUG6Jyy6Xk9GzCxvykZLY
lwMeQnBTLQodSmAejiEFIA==
`protect END_PROTECTED
