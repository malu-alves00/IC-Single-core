`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wrPsh/QZj3SBSu4SdrpXhgWdjLXJFKcTlOmvcIzwAd5GNsDksaa6YFfvzXM57sfl
UXW2aTPNS9Yah0ZgIYFYnas4/X4DhhInH2q4AnoyyJbCWxmMdbgnW8UMdw/zjgD+
6whnYXfcm5Q+5uWgqeF0rZZwUXcezKz80ou3Jojjibl6EuXw/oyMtoDfJiFvSbqW
tMjbUGXKrIdPgf/mfs5CezCq/V5M+f8sHZeC3UPWJoGFezB+Dktd2yrPWqSHrcIa
tIwFEQP2z8+g62pqtQjYf7kBuU1HW01H82FAFmSXQO2EwUlzinrX4CIfO2wu/inY
JT25tIhKIYfaU5SaGSX+vzNCC+DvzkPBeaDVLho7tnFk6IsKeYZh1kfkkHRwSRP1
pOaD+OGR8rIhxgaQyRZf9bxMoRdBDq76A9digjGVvQj0I0EBiR6g7G3CQMUTk+FP
ZgycyYY9viuLg3kPM9f0wUp7YkZ1yAboJL+365hSRf9MI/dU8zw123oHOzF665WX
20FGJJ3iPmh7xSh7pgSZMTn+BuX2aaloGssfedWKMhFfRTPhs13kyv4KAQZFsHZb
8sxFijDKjtdvpgzTwyBRWtk7W/4WmprszdSX0poPCwmxZUbPh4lviurJdD9zScyL
gJYen1z2OrrzYq56nY4qN6Z+wc7FInfSUayOam/WHBME2RILDFm4qAd5bQhh/JPa
Lzn/pD7l7uLI75ra/tnk/5Q+asQ7/1U5o3+1/GdNRP0Wk88a2jYvQ7D7I3R8SDwx
IQ3vvdMM61jFc+T3HBVX6Dm0hP2OwbbfNaHZ4f2huAJAuFNRn3G3j2zCA/luGwh8
jmqz//BUpVKa/DzSZjhz6zeIKOxs1ZcKJtIJN9qk5F0B85p09xa12ppGyC8KMG86
cprqGDAQaJCsBhRfD+VCyb+xI/Ef3tlHDYS8ReCL2NKb+dlJhtAs/rq2J7hXvhez
Ts50HF0MM1rs/sl2tzkystf6pBBGkqD1kB74Yla06Qth2DQQRr95QyPViZXXGOBx
stpsRVym2QKAphSS/7zjByEOJTmRCPC41stCPQUtsAOym2goCyc5OiKHXLHLe250
GOIP6AVy4yWfPadaKV2H99v4Hiqzn5egrBVAyxncHKHWsvhmLPd3lEMSWjguFutg
i01J8sxIjZ8yAKJiE13pNPFLfttOZRyYwMy64yblHbbRWk6khZEif3uGdbFp1fwa
8IucvLBQVD4U9JRKxo9q8BHCuNt1Wu/vQZx9TKY/ZZLDWREWKcYyK3J4lb05uniy
Rf+PPjJJqaL/UTAIviPnZoNyMKKeWj5vyMIoAIzfJlDR7Ol/i6AG1CfI1poE8r4h
n8YcoMl3tLxumtfXtZXSElZI85p37sFUuc2f5j3zHBEP+AvZmzRcMw+zjqfZSD4c
c/q2fBYHeKjzPdArLj9GwllvO6LG8ZcUxCVL1yQm9qo3Qaam8Qs4AhBdO16wzQMy
`protect END_PROTECTED
