`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MHAu+C8jL7RzTskFvR0kzIdATu+MO8Uf4fqh7eidtexRKXBrEW6YFZDLOBEcdJJG
CnB1+e2dgxyLliFt2Ifz712BO/cYbrvWLyKw0qsBkVIEWE+MATiiN2a4odLNfdtX
uSj0ljl4djHsKhX+V9UIf9fKYhdtMdSPZmtonAyfD/YXniWI6WIpH11VgKnZM5tT
EEbh9i5BrUbyUzWh+H+wEw7ML2JvUW2EfSweivo2S/HFpse0nkJ09ZGJ6dvdwXp9
r+ucb95Qeg33Pz/bGMHQBRWGLoF30rhnJEImrwbbRCzTfvnZ+V85+NoAf6HepkYe
62TL4RaAQAp3UHVQG3pTVmv26WLeebAdNfJ74lKCGjwN/99KsLQ+A0O/9OvU+93N
m/hdmgLqEnjYoUX9G+KGrEq0IStYuac7xBQuvlzp5HEHYnv6dbkWfcc9zLEHuZxO
0ty5BxwR5luxI9Knke547bCT8n2tlGYL8sjWGjihERwQLiDwYgvUGzYYfTK2LNKW
f2eqjt2U0ji3qN8WG0F2xvAjILX26XR+3YxnMFnO5tIS0kVCYLwAFr0fX/Y9Id2D
+bt8Et4pqzGGJopnNbkZzI3bDfRuNC4AYCJps2yd37bbUHW+uSD76BGPuTgvcFPd
KzPmKColSYb/k7kIYmx5+w==
`protect END_PROTECTED
