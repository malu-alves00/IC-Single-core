`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iarNAhvNmzRpG9kh2TqDa69BvdDpzra4Vl1C9AQrpc5mWYzO4Hw/+KVKgT6jsxDD
zdoQdEPcOdoZ+pY5tpUDnaGCJJeyEH7ZNjQc8OTOxfdN85u21+4cQwLVK6aCWlKu
K1hx6bHZVfS7rLBerxLptZ5WawixgjFPbfrqH1DkI6zUzC87D3WixUeKUZT8v1eS
ALid6CcomIvRRA4qoIUneeFQzAMOA3yLaaTp1pMs76vQmDH+Wbxc7lmtnLUVi4um
AsYhPYFljI3kCi2+lcQCA1+taUMG6d7t0F+B5GFGAFioSixn1YPnd0b3cg7FxV0X
32BfWbxobgQHWhCFNzUhL6Hjd4ULUBPwfmSjMHtL2NpisWeMU5yPZJUelZPhvv96
7rVBIoj7o7u+hu1w23hbz4+pldp5Z6UlqO6zTExiOG8nRLays1vM7M78ov2GDwhq
qVNylS0xXcC/VBhFJao3ZT0KhG/wBbJMJfzXBCN478zMvggvvvVwxvgolUo4WK3B
heY6x7MoYo/6YE4Ip/nEV05VCXyd7MaTh3kavBsDb/ekJPuUWJXuF/3vIBtORxR1
eG7rhEIeNN4gmDwnqoAMW3L70KUtnYenpOpJoQNWlC0ct4JkQrM7S8wTWe3N8xZ0
DoguMS0FUwa2CfTRzIpNuu0FODZtibiiuLV9TUBzQ77IPNG+9NmOo6ZI92nQQWMG
1sHe1Kx36Yw08MOpLCcpmXUNv5RiQafMQCIc9qfIK5tL2n2QZDxbjVJanumdFAuE
UbVCMwai00deaqxz1DO/IHGVhR+psgJYIailtPeOnpa11J66LlutLmfS9Fr0lrix
KOL0LClS6volr7oed2OGb6QuOABHUXwhk5p5jvSABJp8kbV1uKPdcyEkGje6pfRO
S5ORDrQSdrwM55JvvlO9jhel2Z1xB2WAed2fJ7QAz+H9H6SUeIGmKxVPdfjahMlg
NTxZQnM43UyOjD5EpuV3kxozHP0dm4lf+9x49YzQ6AHwP4ZO5TQJHjv69McJM81j
3LBqqiFkf/o3vPZ5rzd0VxldntamOvzFVT2XmApU7WGXuozqDzbkC3tz79FNxoIX
GKXb8Cjp/dTAO4qxN5TWxLqo2hQrpOedh7+jjQ4ch5285+bwHwRYeDzt7FEtOLH3
FOYVJZJPgNLOXAh3quYsOT5h/SUH4OZygdlAZW3G+Qa+5keIDqIVQKWrol3qTSt+
xhwd4LVw3kGuLR8nozeuoNK/QJCMGiumv5dVk/Hg8LKL2192WyQBxfEJUtbXoXlk
FHgoF97tuAy6OBKEVBt3t1Q0YrmtMjkzUZI+z1EFdii3z1f7kT9UwNIhpYxQnlrg
B12xcYNI9vwj+14yqOVSBHAOOXys/CGqEQ1nNNigl6hLwQbmILjcqgtP+F+Hx69n
4HzxIwyctdqNEyYPJT+r5xatg2ruNJyZUc8T7Rm6DxIQ03ZIJ01iq8k+B7ElQ8l6
8aHyKsbAxLCGCLXy3yBwsVUq2+EKYXCb3vJlbhXTUmibaoCQxQpnDPtM1pVXNxhN
`protect END_PROTECTED
