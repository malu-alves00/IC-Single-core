`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1crdmITD31BHAIlFAnLNUvMaFOQq0a7HLJ2qDRh+tOtxbzzXnLboM8Lw6EWhcHLR
LybIHNPiFP6LijDOj9vqEamc3jJ9I0z6AF5gKe9/PKoYvgQF6VUAbiwhp84j4Byn
qw7XYr19l/lwE37RbLd/kQZCAjvp0nNG/XCdaR5TBHyedi+3QWjcGFX8R20Q+3e0
h9KDi9yg7+WoBX02UGOWNmZvhXA4gKm0UiuzNgl+WmFNY6YNZkZgu9kmFsRjOzXn
dK+PS4SxOo3kFhSm11HXnNzUKdcX9FmZPbZdG8agkkv/+7Ak5n3hnHqOnM+DNeT+
N2L3YP9fXkO/8Yx33g+Pz2iORM5jQqIoPY9ToWaB5d8mAvDYDTGI5WEpeP4Rmtju
YcaaGpj5gkVo7eWbKki4M10tFbW06GyYFHdqw7NBLj1v64eZOPMn5u4L9mcLWi6R
xJxyawJdJW4fOsT9GhU229vkPhgUjQpzLmFN9sWe+M9KeX9Y57xzXrrJY2lg025T
VeIuxWzUZsJZZ5B9QrZpowYKjl7NmoVE2IbRAdA0cmKS//bwRJgCoFetB16v0MAn
GslYW2GychSuA9JcxiV29YWrTTuLEvpOr9uSAGu4HUlY0ij984BId9kKBhUicxxz
Xbs/h2DS7QnbaVAhSMZ05pO5tAGCykZSNFbF9aP/L0EkU3fNxnuCZeZpK2AoLrMm
aByTlGiK344UQ6ihpVGpVeyAZKQGl9hKGc+ZJuPgx0OIidmXAaIteho5jsq9FBz4
YdSZDwpcwzB0uRLYPKEYgiWloXvQEmq+b6Y8rSq9MvbcM4JptjKIA8zK/5YFLRB/
ppR4M2HyU3mdN8lvRNg4Kcy14zNN65pcQEsYlL5l9fxuyzkxSIIWfwlanHrsGcfy
s6t9jnjSV8pG9J+S2CYv+R/VIpECflKdrf4EPDqbHnch4IWLvtJa9+Gzan5BQFmS
oebUMIu7eSbJh+TT3MwBpOHgcQEVO6K0Wrrul6Z8HJX2BIClsd4mzvKcOHejbkqF
fehOaACf4s2BqHqBVQI/f7X0nVUNl05L2NXeqyGrNBS1EKdaRRluzM8L+ovHFexx
fc8C2Bps9HgfdXufZsEJ+bUVnJ6gbfoZZK8LyfMMwzs=
`protect END_PROTECTED
