`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jjpAlrb+E8n9dD1Wtx7XSFnQ/iPFrbajVP2jJ1+Rc5e4StPfsLCuj8jl0bWDdUtg
G7W1dwE9Dwta5Cz1bGyEWQ3FRa12XATIWtizUpD8ePtuMXLlUz3kgwfQvlfHai/G
2GLzuGZ+lZiQBSyz3lJNPBYZHsZEI/tfS7chAiidVhVzjvGu1EwzSJlndPW1uFJb
kdEaZj9uwXOdLsQVOcvdI529z6SGgtYwVVb1o6Ktu/uXA/c7Zd+UqMovctPgB7Pm
v61vNcvdybrg82od4kxBfJ/5wFpEBSzRDyiiHV2bek2EUIAeXw1gBnr7XL9JpC2x
de+G07ntdR09rukZCGElTiqchrjHZm+mmNJmhcJZyC9S5cu9ONUa6NnePV79ddE4
WpoYc08xYkrXp8ol4qbOeT2iXGNEabF+90v2gvgFiwjgYxJLfJCHpAoo1QroVD66
09V/0WuQ4Llj3vpsU048g02HBVCUo7Rvd7+gekH9i4Ilem7XjlDDx0N7gz8RfsRT
udKbxMOFZgigqYQNqmh9vgm6/WXa8UC7W9RgIPQ9FBKRODW0EO2nTJKcwdJqk0O7
APuZjMlb2WRo79U4ukXk90s/84LtvZqEdgAcgK2vJUlq41wKzZ13c5bQW3yGhbiM
AmdziKYnkSnbFSuwzLgcMr+h/cEmrbwl3ammSiXWlBViWFkycIejFPmK1wGLeHAI
mtqMa9DC5RwLH+IyfCBd9h1ZeIU5xNRZLtzJ9emD77GvRZwCAx3imKS8/EZutueZ
FROijZ583VqTmIs/PI3E4B2mlUjLu8yIGdf31vh6Fcg+XwCVaK5NbU/pidQv+SFc
WOCsWI40EScPvGvxI7IP+7YYgDcb8fPMI/BKCbhnfdoIZ//6n6vi9dth99W4BPO9
dW52iOKclG83/xV0ZZnPc2kVDM9q8utSUpKvooQKjRM1P+4wNxYn5wjrDVclkAx+
g5UA/ZZFpwtMUDq6g4ChN0G6scEf3aCbOYcbtHaNuofXcfxU1jlWyxmjiqSmSqJx
uwdW/UCgl3aVELGAR2GRRWcTsWnkPRF+VZ3iwXveiWzqwG2pERdZzoKqxgF+cc8I
E+9MV6OWyN5KpZGbhINgcSMHzBM9M3Cho15TfzGObndWFzKMvgUrONbi/x/iCEXn
VXaUaE37xmHrApbQfn4w2f/XrCLbmYS6BOpwp65GVg5pNHM/484YDbMCQ0uSD5rw
FzKiTLJGuSVFse/xEh6dUv1iNVjVuv0MCZ50VvfwoNCkgH3jpkWNZaEsrwgod2BX
oDPH3iZiU+fnZomwKtmIZ6pa5xwMnCls3hXRG+J09XNgbSBbgCUoPCeDIATGw5fX
Ckh42eJ0oJM5y5JQl5SB5Dmtyod96EFETi/9BD4xkvf0Ly1PYJYcQ0VMdQWxuJFz
Td//cQKveuQfW05xsTYlwNTq9FDlymjzvJYRye0Y7QdpHWeVVoAQIqBo194gRxJS
25A7csJjU23VpX6sKG0Z8zr3Ot6ghFbRBBxF6eIQnI2YmULujISHIIlsSUgsOzta
FIMvZHCBNV8+aToom6l84v46G5fc1FtzXW0ZbxSyOCwBYI50nbCNZSkl95F906bp
0qsCoWIyHu6zdlV2boQOFTuXcsxp6hJ/ltxzlRwD+tTCWvMSAhopBelIXiqyK3M6
1a6hFb1it/juaZ0h8P01S1/kAxlaizE0VzwXSjwVTwYHH+Bop5VQs5eTdF5b5GDP
6V6AmLOynKR50aV0ZaTWEf8ouPJqUersFuFQ9YLNJl7g7wyUlqZlnKmAYmwe6sue
0SoU2mbEfJayKBj2Kie5nHtoWphhoIbW5CqXgo/5NnN67U1CEkEwDujnjZVNniIK
M7LVBh1KtCTFsKBwMihfqe4Q807VEA2Od6ic5DNzdxJGCpmFGdy/VMso5NVkC/OF
jvjvSwxP0+F2bnCgmHPqqd2sl6h++mApZ+vrqG6mbiw8yJHqrE+m189zfn0Fv2fi
M27/K3XJk8nUyci2B1gVyS6S18+Sb5Cq0POY03QMAFMPnmA6oG8H1HFS6Tzk4vwu
hOvvxLFoaoR8sgAtZswWTeCnFie1kABIFmSiTrfJ2/RlR6MY92jCfiOab04fav+4
+UHtsXFyC/csRF8fxGJlB+ulUWHKQPMnvKUxCZqwz97LeuD5FNQfBx1CpjAUqGId
or2jdiaY0huMnUx+o9EQpjwd1EoEL4g3+N/EJ50leLFRccMIVTPTPTKnkEwX3TAa
kqLPTLN4fduEZzx1NZIatHCortphCm7Fb5t84C1UOBBbsIqfoSmlvVwAuDfs0t93
CyZGrixy9akWFsNPS+/fUJXIkFTP92xrbFFs9vdbSVu7dVkpFed3TNhcOuLBh6xi
c9gy63oqZkW/uFeL61EyrdboptNtFkI41omaK5aHSHmmO3te+VhRGJW93I1zQIvT
yTm02II/0AEV7VOFx3HpO9/oWEFyxPGOYVHOOix+grsExmGIN7ROizmdInm0ly1N
K4A07elhvSb4L7mWQ/L3rbE3zCwM9Xj9mpxPmHcAzuZf33vpDGmOaifyHtBngeNo
lYkhDpbvU9oopn4AtrtKNDkg6knUKxL2hoQwRtAo/Mslysf5JTqrkqW1tbL4xflP
oTJQFT/G679fgEOS1ZUh08R8YUId/hyt4ISj4Su23bwAUp1eKyOMa76tdBoFZs+Z
rcd4BWeUTEH29EbrDq2erpxe4uVpG9WhmVJugpnk6R6JGu13cqYk5HmAxFgZ0xfP
BpMzpo44d6DlXPQKI31iK13dvNOOyudCDxnwyU4MSLBx9HMC8ClG76mpJPvF8NSJ
cmgq14R1Sc2nJLgDzUa9s2zdANM5rhxZAXzydhQq2MPxBxfBqCxo49b+movDQ/nt
alJcYAGxI/r9F+c328tONBN4yOREJ++zfvs9lnYsQ7Qa5beT+61g7V2KLH2Asyo6
TVw8TFywFjmh+g1qaHD1nvCAyn8/jSIYRFsRJaD89jmQMbg4P/p7NATDnJd3qPK/
Q0L84oiHFbjPOXBnxsV3k+u9TvRwQQQ1me8K4LIlRqr0ub/CLUJ0KvCKvCe4Ewwg
v+YoKk3tMTIgazuyUfNEEuByJn0j1SyYzTeA576BPr7h0tUXadN70Daw0mTCzv6H
IDIdxrifrjdTPBY1soCQrL6ASgMP+DkENzgi6AQG/P74Wi8Mdt13/1PhIRIP5C6f
cM6txpqF4FAofPxXTdq3PdmmebU4Yb04uMAcFvSpdKZuF2eIYD7BJjP/UZDxqiLp
J8ixHgaCPwwFltT/OckhKLja50JQgv5CwkzduC6AuxnxOhPH/m2iePTDGY9pQwJw
6UQqLXGO1lgl/29yg8BZoe5/ho/cViDKGaXu2osmMxhD0yytHErIPJrbmm1Lu98i
JQpIKWpT7pxsPjq/S2IdOa7Pj2mZ0ButBV/YWa2Q+YRMU55/bDZRX9vhLdJd9QkG
16Utlm9bOwUwqx9SKa5d1TGsDZcQBReUBJBcb+rx57Ph03LQ7YuBlcymNlBo9n7b
WmMOQq2tpg5efbnYoNjglbEsOyB9Y1rSxN8dkx76k8C57PYk7judncJihWAR6cBJ
VYHTrcFclFeLrk+WcpsXqcHBkzD8wpNmT3jOhLPbPEXsk8i0dUQKOPV0qYBnTw0i
/wiAiTEVLMNePEN4PpzkKlC6vXesQR62IuyqGBa6nW7JBb5jOyjmOmgqxn22lwXj
RMnftaWzKdhjx619D4wC0PV2xEP2xeGdjAdgGRWVu5zpXrGQLxRUEPoCwpBavN3Q
65ujX+rnrMlDDYbCxNDhXxXxdzMSA9jNy6ByBXg7aFAYpm87GbCFMwlxi4gStARu
Yf6q6lD7AKi7sZhWBpgPmFnYVTyxy+7xs//YQIJVXxkUhVWW6rDktY6VorxAKbxl
T/oUJ7QGYBAb7Ms4/XlSaKDn5xea3b44x+6wkxiJAoLjknDeWN7DhbXcwidProYo
4AH85edVBUDh5h3Xf5qCv5vgOdwB/MjIHcMYQ/HZUZK87jTpUNhXkOUeLidy0IzC
NP8vKXFhNz235XnnfbCYJmeVxz95vEfwg3ojwstZNmJrx/ZFdnO7iuFJlXzQAPk+
yTiASo4yrFCL20LtA4F16+GlNndIGSnz1EEYBX5JXMEedydWORn6/3IePlXNQvdx
Mtrk7Zu6JdWNP+3T3Me79/lopr0lereLV8Y6325z6gb0p9eTgBuwSQSSjNUkxLom
cnxTkX5umk9x745Z6iJyT/h/zFbIV6OUek3n9njBLXuD9hBx7IsDaRe+SScHF+lF
u2fzeBpEVAAK4FkzvGlFwHEApN0N6+0KcGtuwUL9VTC4cF/jSq53QNlPAz82M1jI
rBmIjQiL+E19zp28YtzgkV01968Y67A+XW5rVrqECDa/+FZihjqQwTiat23wNJDk
Cfm4jNwWGVWzC0YTGluVlDAWQuUIgLDEayXmim9deRAwGxNJFH7pkThyWCXnnaom
eSwllAlG/Xwx/t02ajlAHQhwcLQL7C/olXJYVH3DiqjWeNbe40f+ujHjZt7AZQPU
LIygEihkwo1G/iKPoYkSCvkWucgff3Ln1sR07NT/ipmW/P+MqDGCzo0SXGYUR8+X
f28laOfDmNqUuXJDDrt2WSatCP4f7uwHtB0AeHwvFH0CztPCt69R8grzQN8uMVYA
JZA29a0luiQCLljxMm1QfxHcL61YU2u2KhWeiL4Kcf0yay/fsNxlVprKOrc/Z72L
obsDVMMATW4tE21WtvbDet+0B4W/ddmKUWDhLWig/Ip60fZKffFdPRi+4JHTFCQl
XX21WJkHI0BXmcELRyojVT9n8YAtj5h/fNKEYwOW1rRdCk0dLD9CDchIxXKCLWGG
vLI6PznOD0oSFy3JnGodLTkM1rOcq/aFcf1Pn/YHqkNvukVHAo0tVAtNjrB2gMOd
pOVJS9sm2Kk5ciB76LftKnHLiXFA+DZz3vdgs37h5kL7RHCr20GO8xqVQG7pXQTr
ESRO0mNiQYAyKYyJaSwO4z0o+e1EfqeIg19h3ZI4/+dsM/fk4oSgWRs3eEt/mMhB
Dmf3l/UHVcGfuzp8/Qzt46uPow/XQ50AYjzkkoL4BSYGHF0yRCh9/xwbZG7LyQyE
gnLj9wWwoN0i2AXwdl8MZtLOOIeiMZyAjM1XMiDhWcJQOpt/Z8l5/odp6I2vt679
Z0lDMXeuUNie4SJEYJfs+haJwXeaZg40eoTQon+6kP5l8aZt4/7KmFMKBrUde9jK
fQM8AIWApDUebH6NpiPKWyyb3c34XH0gTAuY78svKjVluqv+kDJiKsnooLAxnYE+
feRpt4LSBtfdwXt3fLNNEowSt+AJLvkwNTPsOxa9oJ2RTMt2WX9kGGGsPQTnl/NC
Odjkj+/xelpJyyY2Aep1aAGJm8WdcdUduZrjSc/dyxLDcjnfk8Blz+A8XiMG2zbz
ncaD7zxAHnWpuVa7bwk5qHVw7eR3y9gqp9AGX/5gkhfgNkzlP+e1sxwYfWHvJNsy
itvw2m8Z/VneoCCN1v1XRZtuQpGyUuTp7JTnCKT4ERdIQqY0sIWWo2CQmks/+ZOH
oKiysFld+VprwMMs3XLLJYQA5fJeIQHdmrut4M/NW7bM7kepe/T17LD4fn2PdfHJ
ae86oQp/ndfDvCJre2/5osJu1EpkxpKsoY50kY4YkORIVQotxmMrdLLsYwn0H5X1
8Y/vzuLto/syTexMwxDfhDV6cY8iMLgTzH/9jjz9jzsYJdduAmsfELkyf4Drk5wM
t3VvucXILRYaPJlpXhvJYxfk724H2O2EOaGSbtRjA5cl24bQy3qD6vubumRyPJLp
rDz14qr1VONUnPpncBqtO7snFkJS/YfVH8TF6kNIeIJK00k+TRExFPM3eD6J6x1r
RoQspMH9tR+Q6fovzWxeukzcdbjd0kP2P6gvoEvstkBL6YNXEu+33vZUqWM5c3aa
xVlr7PAcTEqJw6QpfrrNfZSDtifQyMnS1MXzRSvwhwp42MImJfuP6RXZW97rNxHm
hZ0l8wSgYqCjGjs4m+wY8QjHAjjaV8TdBs2JKy8PWxq6d2nqyMgnNF62Sz1zN3GO
Y4l6M5hoBYKjhgG2T42x+mmjEa7jagRZJMj1xSr4XlMmQ2IBg7pac8ezbvEbumsU
fg4FQIu+PPOgAbMrGknOx71/bgqi9uuX41kGW1aWCvz30HMPHtPD3XoNp8ByYdCh
9dRtPApVQBUOZ0Mtu8PNU1RJOCui0NcIwATFH3VU+sg1jc0PwcfIReW0udxJyuyF
e1zXS/c6V1S02dMCPGOqch/QxTwGol/hxdZecwugasu6E4xb91tt5wWDAAItuYmS
qaojLmS4Gy/vvh5WpEPQoImwgc74d6QgH/bLdw4e6ZNWVMYvVNoRoEJYGjttUnez
j+kmYBF/nkJdrrjWqrPNkLbFZKwuk1HWGENRxNT+lkZ8/iofH6UT1CgafgruL+Cd
9oP+wYXbf/j4oj+HBShfluxYqvr/Ms4O7vO7jWG05DjKDCSq37ix2dx/U79JklNz
rXUgzweYpw7pLhZ07nQSD110pX4koeijWo8TYIIV8Pef+a3iX9Q0O8SvGYFaf3wb
BSc6rJIvnBsk3Ecd7UXQhUhhAjsI/iWcekd61CbaBZDlZWNkP0AlbirkJU045AAF
evggwXZWRjzIcsoIBO0KhK+A3GoB4qoL//ZnEdBXvBmRuRUUJELsq6WgSDeWTHy8
uFHoPVUtRf6++Q9LXEn8ccGi11D65SyWF07xelbykoxm3/0CJ0zrZ1yx2rqvYZbK
Z2zm0gkTlEI1FZ1vb1WLzNBGEQSbac/Ks7YPTB66BgGVywpwQ2CvIpLrJBTCv1TB
+AvgIjcmPVf76bawdi6JM3SgcqVia3c/a+NiMl89xBb/KXxCUP6D3l6mWckcJUUg
XR98RTLeDU0c/YUl5FT5n3NK1aNJf5hZW6CqjJOUzmSMkpObSSAdtA9TY+2skHLv
Ln4zTQw0QUZkmOwDhqelA34G6yrODx0SB3JbCYsy/KAIn4CAjE2ZYS5Eji0uB1yR
nAubohm6pcjtlvG8K7Rq4ze1iQzHmYSne6T1V7Wh0HNtOw21PgP/sHCvlcDA5p8Z
oQpJy7BwgSDwbhy7PVpLMT8xVT0Z12l92NPT4Zeh0LdDMNDolk0MedL4VHfXkNFs
XI0ZJeUTVwDPgjuRJCgdd5uekVmW10Lz8yf80NEvp3MnuBKnOLyNi28YKV0h5D1Z
w/ErJb21E6psHEVxr+YKRFjC116wS/KSrs+WbXe4YJWMAU/pvaHT8KeMdIJIM2fK
Hpw+vLIQRHMJJlP36C0biT9sx5OoOTud3ad8jIpMU10MOcYQUyRNIOK5AVvHEt6a
lnPn5mgA6avjbqNcGVe/kXdl2wevCXHIRdc7eScYZSXph7oiQkmmUSC/omugSjG2
a+2fwJAla6BypWgob+acXP/RrQZ33v5DnqfN5lXMjbPga2NhVzcCbhQvHA56FR9u
JteatTOKHUygiZD6ukFQt6XSvH+IDkVvAC2hhsInwi/IURKFNiuG/eT14TFJZmxJ
ov1WYjfuK2MuNdXxht2EbXPgrr7VN72QgwvDLPIgzUHQxMJuFSr92GnrzcOegusR
lbZ31pGutIeT3ByfwvAnTX1Up0LX+1X+06o2HW/5elt0DvJetemP9ewN/DGAk3gY
edF95m7FJvgLMFHGErcmElbhUdIdnIv6tfQnGz5x1lq8dPOr1Ir+J4YVhb9y8oXW
Ovk0asH4btcKNyN+o9eNYsMlQUTzIeoInvvLNm6Q8xsQdsP3rmEVyXhX2ZyDa9su
G7kbA1pOY6a4U/ls2Nw7sBc7YBUk7R/bXyXNaK9Fo2q4y0/yTrEE3W6leGQTlyLj
rCv3xwTRBIJc5mc8BGB34gjaxHailt0Jp2VCBKe62q9LhB0z+vL7nEH6lq4dUPg8
CJtqXXYUwiLLTk1yOh0gq76jGpUEzlAYFeNuS2mAftqi3doxyWx3OCk759n4hB8J
jBjlEUpaSiZbk235K3966/vJckVU+m9Ymkj5REjmStJrQZEHF25aULH8nzScSfqU
YV9dkYwoJYO9XUwCgbRrUY9FT/c98a9kInc/LqudzGxQUlfSDCG/ne1MLXvna001
NHbWuA0fsUZZ+rzO2lx2gBZe5ZR+YiN9VjwCXamyBWHBeUYl7mbziNUYsV3Fo6yL
5L8RYVccPjWqIgyZ5tbFD//Okt8S1hmwcp2jKMKnn4tJjQIp3VmoIfM2d62u+egb
JM+J5JRa5t/D+d9aBJtONBILlf/uNclHR1H5gIRXyeCuP1sUHm+LYlRaYqnYIuXm
fl3xf5oJqoHxEXYEOuIUdDTOEtHuvl9DUdkPfmc+0+O0LUD6xX2qFspPKxmFjlB+
6K20e15t7YaCNa89y/u0PLUWYyTBHRg5WZvfzDkiMIlr146Qur0sbKp06KtiuL6i
EvYmiyuNJ2C5wkhvyXZju67y8SMcoyLRF/UF7msM22apMFrgk6+6QCnLYW3Fo8CG
ZqKT4sZOTTksOM1TruyoHchhoJcDD5aRbeJgTBFq4qlsalvmwOQ5XV8eGrsHeMfC
DldpK0Mp0hEdbIJkGiBOMljBLM/f9wZIOocMoZiLF0mA/Io//QSmcxrtBM4Raf4H
CyJlmaRfOAWMzT20+SUZs3zn6EwOoXSwiCmBTInMOdbs9pDFabgAz8wr72jS/sil
v8zTQugMrzR9m4QNqdxXQy9qhC2oukonQ3qtY4yHt+ldVP5UaIjrZT3pZY8dLh/e
RqUf7xPW62hKnqmjOn2jXYAdS/LKUJ6X9X1cABedLsX5z2hqVKtQdzE/VG/r3lTs
HCtrc+/iRPiUV7ZYdidjQ5gpLX6BPFUKdYDS/yWmie0rtQAEkUOdPoIM9YQOQ6co
GgSdAobFNv3nku6WQpLiizrFlV0XM0T3H8GXqESMrmzM1ovMMinp4YtMmYa42DfA
f6yidikEVguo8sXJwx69U0Rsoc1xJVWjIAoLcXDtrz292ySe8TrFCRGSyePbdVRw
LPPbvHTI9foVJh68OZ6mPEaQhJFoBKmrTF1ETyHMazojPrGOc0OYKAaLCl643Van
23+RC7BDzTBSns3Wj+2uLxAwjh0USBsNp4xcnCFDuFOKJDjgV367zFcP7maXqAL9
auXeztWjk39pOqRtCJEe+FCKZQskHixBhRvMvchkUhuUM4QBUPfy2/aDUI69OPAO
NtG2XJJmGscfUqnku/HW53KgKSleZPiUXqMKfLkHVwIgU10aCbSsvzrtASPgbzwi
8qM2S439FUhaxr3gCkxTd7cue/UQenZe4v/kN94/9kODItBrEGyw/5lP2FsEWmeJ
H79z355s8ROHFFV3wjz9r2PtdyOCXXIKc53nfiWh4QWdxrpDXMSfZprBcCEw+VSC
aBpa/PTzH57K31ynDbDQ9wdnpFvF/hcAjgw4q8YFjAcfe2p5cVDCNiWqpRTMhwsD
jxrmjCOdRrMfLRR1PSZdQi4ZTq28Z0K1VTpRCx7BDFij0LLHvRdbvxfr0mzlJGqS
W843UmQf6VwOuDoE4OyZAHwZ+sM6TR+qiW+zAinNCPqRmbuY/BiadQTcVbzBUaQi
zS7ZA7j0cJ55jrrEpNRa8/KeQYQWIZePYx5NgODmS006sKfJHNameB/FKVfF3DEE
rTCFR+6Ov6Pc+MkRxEVHBvxBje14o0O5tpsmqXEmv2Wv/25L12ahtdaTsf93Mv1k
ky/mPn8cI/Bh37RjCMqmSQrGMASgWAi/K7aqajVMn917zozyX9Jg9w1WQxplEG/3
TTO8vXGkvsPHnaIkcgC1MHuGcQfuaoekx2Z0WFK8h1r/7DiBQSslKYdWfSw1wBDh
QMwF+G2cEUOZKkKm0FT+lydTxmpb2q+9ekrJe4cRF3smPQ6Q1vpkl4F4LsZqqSZk
ZsT6HFkjtQccdezdDk5MNc/RcEMfTNEbIz38ReepEeWhec5gyZWw9+9gf9s4Erj5
oEvA+IYM5PjTwuvOBhQTkUMQeYzmq8r8Xa/k8b1s8L6OLudRXIQ7+OHHTHcIWF0l
0KRSmIvqI1yxzLa0KBcQoblzPu6P9cZdW0uEuiyf+uMAWSpLeWdXkNc0kODJl3uN
tIlMpVadHscnknyIRE5vD73D46iWaeJ2I5khL+CPIssCf28j17SoH+0rkU4WzN3l
KMwOsspDn1umAynbzaoLJ81Z438dTJDHNIVOLQu5ih3QB+YHOsF1G1LGRN5c3/IJ
E+lOd8cwzYjph1QrHyLyjEbuysJLqoPhhd/FSZWov5Uh9nomujosc2+Wi5gcTrVQ
b4ouXSYnkwYu+EN0Y1M0AfX09HvqWJhwaOTFOkbBMURcVdsK3w7yXfF7FF7YISGV
oDev1bvlgP0ZXya6hYscUFnY7X84sj0+7I35E0NpeHFZboY8xSfS9GqJ3ygFqcgL
ZkrZrIZ2mbQZQF9lGKkBFuafyM1+sFL9/kWmOusSkeUmI+lHhrPJEK53nWPqWG6E
OTRZSnP1qzuSpSQ3mpNpMWefCExE9hVf+mNlXk5kxt3Ha7NijclYhsVBZp+GgVeG
WgoT8MsoGEJjGueZ/aeZveux0wRYpNxPVPEkdvnkCVu+gMXLdfyj2g+OSzFCN+jw
/AEezDwV4DWgG80Mq+Boa7EldG3m5oT+oUBBtA1LUzjaVW3iI3IhCMLLwFSfesk/
viA6n4KPxmdgVzR9yGXJGj5ZINIyeUlQYnyBZifJ52muBS3uqcjBClVqnLmm3jY7
utDk9zQfJEhohUFuDSb79/TVsSR/1WMhkQZDN6nK+vx5oHpaLj7YGExWstaJsOMY
zLTcnEIN/shqw9zTfcF2naki4rDzd5kfCy0IujQbx0L/9UT1ERmEtPNon0A5X4SU
Yh/HId5xNqWiclRZS80fXNh8yXAOH22znCK/AYwrerSYTmxfzrhtCP91SPDR1HmC
M+gRNfO02S7g5afyFWMb77J1BERV82whxarzrOOQMR4tlVcBLq3iW+bHZZIu0c6g
Rrtko3njxI0h0uEtfBEqblvU2xjQlDeEK2LxOIFBEq+OCaYwtd+f5XPUv2SAVXsn
vdKtAyUPL/WFUpMB84Fv9YXbfzMbX5RTQHpvjL/iDNmvAE9nPefKgjVOTnqnUYw+
ZXrmym6Ol8/XS1H66Ba1Ew78riL5gluy/pf0geFF4QVeep/HDtmzxNHtO7Mxnig6
0OpAnDSOCYc95eQkj9PDK0NrBz7najBZmGo94VhHyUAww2v3sZYNS1ZTDSlUx7TI
CwjQILtc+odgF7djVcOuLlZkxXmBN0NYXKn5Q1cyIJerL6pKsoBSlBgr9CCSb3K4
tg8RlG9v+cnx+ddbcQAh2dEle/dXMxPtPfoxbU0EG2iHQYEzPDV/wXv8U9Sqq8Kk
6W5MlbAdlXk/udWjLNUh2al2tBmlp18JwS1LrPCPUh4JFcGxdIdDLAKpkWCRYSBM
J/m6RKDrJiTWKjBTdokHGYvXaGwY0dmsasedwgevTIISo2p6xm2av9VyuKoTPiBj
oYZ2jpKtP4mnxmsVEfK1L8dAs7WpsIas0hjPu8WybgVArfEmu6ihyFuGqB1xdgUS
Grrnzd15k7Al+Sxbz/xsWMGyroH2cWax7ZDd102wxFn8tB5HmZYeZa044Sd9z+48
qA6MTFAiTRCjg8lDhUtSGiaE7FgsR2J7WXBT9vLy55XWrexASvmCmuAKzPe69M+m
sEjqOADkq4H7ehIFs6hVedLieqxUg6wYogmme71zF5CS+U1+/LOO8Z4g2VjC7QEa
fK6fIfQiUo2Y6v2YGo2MD8pMjNI1xjNkJdAuEEfxmPY9SdkAd8tnlInJPQScjU2Q
sW5SN2nGxMOyK58gt/gOrsyQE04XmS6hWDmYvMaNx6BjQZDUmyGnoMxL56lOGSdE
qa1G4yl+vEHAg2ZmFDm1f/otiRsyTHV+UfSTU3RLYVPtjQRprmHh8VcuKRIBh3n3
ckmouv1fqtY2EteKp3d47Nj8/10vUaLJ7dhw8tJv+xfc3AquS0tKaLdGePFIJF1r
cmEJzxP1LBXtCKWJXF3D6y9jILsXY+2c/vX0+Vhu5b1r3Zma5LpzHJ8KZdrAPhIf
ZHHUGYpJO4ltGXcULURfuNp/5k0leYyVli8Dbtbty/Hs+OmYmVqbzgO6jMYVM60J
hnmwVcc+pGkl5EhCbqf6I6aSfxbKoDfX2ngj3PJXEinC3cRPCdZBQc8WY6P3BxdB
EoZPnSZDjvpXachVecjlqhEhaswh5Oirqb65uU0a+kV2ilo+nU734Acdq+y7sxta
yd3V94yH88uEUsFYbnRs18yxfasEH00+QchgpdAO4xkhxvmF1MWLm3oZPXzfHRut
GwWGv8xQzoESomJRTBYY/NhD8LHh285h2KZRrPzB3qwunmkaqfJiRQCH51BhqZyO
Z/vQJ7LdDi4jC0psDPhWcnA/3XNNppXvlWOsOWDtweQuAwlmCS1z/V+25Sayo3bU
Enq8VjBuXN8w7Oiev78v/r36/5L29ZCS/yXpuFi1g2llJnyGbuU+/FGiCbTJ9N8H
BII7vnSVjBfuUJB6kcwMQyGNej/djgylUN1/1Dkhjeo+hC50xtMtH/FBgNGTJ58u
dFJncj+dSKCpKCeukFEhml5q536sZjCum7/H16y0lGJd4zUG1joCENNLypZV65Du
H/O+f9ehtpnCVKkmFjoaqeUkMXtROkM9qHixiNsCMBSM5mKh66q0viM3qiPsmrMI
6iDiCKXD9zwnDDdHXi+x8joKbVxevBSgxdh0rj3JH+UWvs/DHGqPeHkUPbeU9cnt
UbfdNuQaPuCIq8EIdGMZJwaE7pCI2PgjIfm/C+RJEsaupnEcU/2aP8lVHn7WbN0p
KAzYgrNoir6XntjkTD7VCEo/lNYAN9coiDizhSbSU/g0d9MONTOHyxiuGhNU+m1h
CODsKL1wMTSQSJYu+pLjlTod20G8i/82PrpR/F9EhKQxqyCWbP0+MJCbzLWQyR5R
5Az1ZfJmkgWC37FeBIj7GAHxxscpmL0h2FN64cZEBOudeuU61a8FycXcZgRyGTSf
Fti4mSBhRLbqIb+yvnQo71HxAEWSSTntiC6tFuCknKj1zEGCvH74gI09S2rCidIS
75ESWKUiKRXXhR39U/MmL6p+TdmOxc73fUFHxhkS37jV7/b6RxkXOfzEKb9h0heg
yBkydEEZiXDg3Dh2gn5RxDgFSfJdi5XCDN76k1iQDUQHloXOEn944LUxmXbWXQzd
6vvoh1ySuHA//syI/alk0GiuMZoNC6GI58oN0qMowO+SaZf3nF7f5GRdOydzhIvA
fRo3SXhS6sSWffWDQTXHmxfR9Yvw9qu/T4+ykTDG744xBoCECNru4YNhOuMQyidy
YVPbCuAQF7g1nQeR7KNp8wUZgntSVIYWlyV5+DxOh6Ycz3Yl7hgDQchIxMvtR4fz
gTFYJZQK/ZdKMKgt0GFVw/4kPkpZBhykdMOxRscpe6JKYCgzA6EoPQLtZrukjPyV
FBJF++yfKlq6aNevgVq/DSnFUiGe6I6YAfUL6eUC1w0ZywzzZ+PdaBNB/sLIM9Nr
HKUoJ3i7ronLXbr/LznIjOi7+dMoVGWdpiaubnMG+cIPdePg6ynrSo6rRVKC/r40
CI1UzFY+dtLGBoxzOG2PSgYLQaidF/LrU3GiNro6Lu2RdIvsZ+izq9awX4ykjws6
pySlknZLfxQlzHbIJMfwQ7zYTEJNFvPSX93GzTfbSYhgnUmuuqexa4Qy/+x5mlJw
NRbewWYNXpGMNEmvTlg6mVCrGovumGeZr6EMdABksD27v74d0nFQWdtb9ARaA8Vl
zkbz+5Cc9gl9Z5OswasP6sqBDD8Otb4BlsCqkdykll5qS1g4lCmHmyUe6fQziAhi
jm9kbOK1XaaKrEln4ErGpXTW5F1qhD2h6vcmmL17/da33G7yX0FCLaIPxm6nrn+I
UW7gqlU5cRngfI2eOkIQ/oKqUz0SRn8zVBWr9GRSEuuuRxtZeRUhLZ2LXDnDftUw
QttmV3GBkJQWwigXFtFBlfTUwb3hINNmMXER7i3CCBG2jKWmNpbTDm/+1CjAy+Mk
2jNmCbk9ALPLXeoyQ8g4d+8J1gZb2IYYA1oIdzp6iqE0xly4y+kT+S4M+eAjliAo
3/hTl6l0j89qv0rL4Wp9P4XpROETADrbMu4RHCeFvU48SRC8DeERwg4xuMSyo+g1
BioUWUocHaHWNJ+m8njrUiz2CvG9lUzooQ0rpWajoSYw9jm1CuoI74U4nQdDnXM2
`protect END_PROTECTED
