`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0c9bKC4zrc7diWoT26nGgJSmc2sPT18vaB/Bc8mxbQoyyUV982IqJyJMaE186ZMB
cLKtxDyaoKHEVtzh2JUfwUKstn84q0RY+0o7mYr8cCWMYgS1n/Q2dgx86Czt3kZu
TDS+E5qhycr9QgPn80dPZ/uUxc2JFFsCo637ldu2fGaGnO9jDuYazHP+RAZm24UU
odJ9dWoWYKb0F+lyiGGV+vna3MNjzIrqnvaesVcbTzKpZBj1aXuDTlagy6TRoIf5
Dm561eO6YgH9HaDp8pOTcVlK5xCatGPLKvra34QGovWOFdU8h38vthU5PSwC5ahT
hT9ieffvMQbg38B8Dcx9+mnToSARIzeCZP2x6OjLpU8QO+ODECdTlFW97AAWPW5b
d717KNp4nwf5mszqJJadiyTnnuM2jkHnalGARPa+Nab1G4JX0zd+FAbGMreDG9A/
4gTK93FqFfKhyJw+tqgiPwDNEh2Wrli7YXBTNHZ4xlN9MJx8y0Kt/fb8h+1vP2vG
KGsqHgb24QejpG6TTJRQOqtMDjYv8/xiklKtwvB1nC2XmDS73vkp7IZrH26RuVTH
XD7cyfr0haZ7DJ5tVvqZoTQI3frU5Du28xa/CQD7NQDcCwOb44HAy6LK4JMsFSTJ
zPTrHiViQlPNURkZZcRp9BsZPbmkBO4nP+aGX5T26f/oTjeuOf7oY6yzMjK2uV17
hpQmv31fPDVU99jge5o+bmKae2gQ//Vk2F3xpxrH2yIw5O/SiaHpXVKmTne+Zdmz
slYIu1UAzdGbVPsSWbKI4oiJV9upJOnEkDVVTc9Iw2Bqb6RN7+as/iAkdE09A+KD
ZMzmrNbLLS2bs1ag4ZMb1sCVHa6EwyVqEtBARBrPLJHROAYHoKgF8qP5pa9+Vkzc
D9wv2Hda1lp5K1+3c1Irgg==
`protect END_PROTECTED
