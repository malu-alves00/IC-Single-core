`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pPfzp3TG8l4hxLLZ6ADW8Vt15XAIVSkoF51v2crzoqffc25DQ5pEy5/RTuaK/j4d
vTch1B5gKiO46A6xvkuajRxokuV8y4aarWqWyjkfvZqL5v9WWB30zTrGUCJwzPSc
FRQ5CzK2lhJDxbfCEx1NYApG/pJPh1YEG6W7Ef2CMyQudDlXsMMeStzsioX1UMnz
szRh9U6uExGDTEazWSbPLgjFQ4OBUmflehtfVRHs8pKlzVuIwo09smRYJg/n+D5q
DlRqXrJV5CWkcp15PBC2NV5brd/eLiQQp0OXYm00jo5Z7OmBw7xS8YFtNV2TPTwr
QYkGciRnYgBrn5LO0A3h+4qxaRxOWZg9Z6oD02gRTienOZaYIcTAS48HiFMCnUwo
J3e+Cd0ELcVn/Msh66ul6aJZVoPceaeDL3gLNmugk3mTOFw+K4x4efq4bPPKRxHP
agbFkqWLeHKUbfOsM/m/DUHjV/AfSsch9kHYVrNQnz416pNYRKKbPdgAjKQJp560
vc/G0itgQy0rhh0VUsuvH/7m/l648lf0FBUS58vjMIlWcaZMc7nFs0Siq2x9/GnS
JSfcYGRHNKRQcarh0WcfrSEs3HNQdT6+ADOGOhhIh6lnjj9yRu1hpYD8Ag+9/Dhj
swt+YmeobwFUGPd+IkmtTBJNVNj7ITEyNypgnIM9wfomUeFmH/CjjQmLwqvVTCDv
KysPi7MIPGfod8X4bZTvvOVyBAcQAsl2dLvLmUflr9c8M15JmcykN7KCQUaTHjnM
pqKxv9V8I9GvtYLhSpHTWSoW+TQ4CpzlQKlszN+OEWL7JQvg10k9W4TXWb1U0tlJ
Mx4ytDgtfengsBIpRMrO+HS0iMRyNHQE1mU1UZW7oPVVp5nGixaG4PdqsFpmC+Go
i0hYXApsbk8MOR3r/7sgzwz+pR1fBxSnvo2F5vRYgc9xpGya7UuQWm6SnfgqV5Qs
Qaj43YD6bgK1l/Zsg5jle8VhADzmQjQ8Kuu85RVL1WytYXIc7ELujWfW7yPw1XNa
b6yFAqXtEXltp27TrYQL2NXt7AND6LEj3R3fAjXcL++QeyDwqMi/JFeSXjqWqUo7
U3Xv9NXWwpf3VWoNVSngtqAhJ3TC39TEwLXUWZaM/x2SYFElRmQ1xqL7q4NtTkBD
YCnRHg7Ljfcx+CPj6ZaGYsszVNM7ejc9DVZes5yx1DKuDdA5Dpn+KxDr15bLv3Le
swVvQ4zVzN9BCaks45nR3/BGVKdtDihoQzj+51BXMIcrBIzY9B3nMBf1mmL3pJYJ
l9OaHpz06WxNtWZNolmnYoGtEjwu7ZaCcB2kLl9zfYOaP+OhLKNKU2hGI1KKiNzs
qSC7I0058FgBKbWRHOEJHHeKLTA5/Iurf+/laeH/Wth8C7io5acme2gb4z4ejXq8
gWtvXnupq/txgBBCpCmWpygxqzN9sSUwsingiU3BPFWP6+o+XBAehAxf62nYCxma
PE2Seo6W1sVZnj791EkK10jpmxaH7wv93szarxRVj1LFYxmE3pqWeyjU9/+iReXn
setsZoyAcQAlU4da69l6zDLrQwgm9+XJbu8mBw/VD0sJER6yUxSPgaPG867MCxb2
HzyTSm3kLdZdjPwrNJXJOWe+GcHz4OeeSblS/qiGkXYnwgPNiUnUv/vqJEit/Mtm
4jCVcOEs71UJ1nA2le/oUjomfZCgL6Q4e0bPg2n4xNG51ubRIJRzWCMpc2f2xqYt
yIu+bs6wn2zxD0x3Mp70NQglcMMY800nyyCVtpUM+jOB4sPZAyszp4tmat1Qlo5F
SDuDIRU/s+icpA1DMh9F3uPn1YcWcmrlehrWTdpvu4KEsZ1FgsWVYYwdj+7JSMnO
+hxbzUKCT6kugmnx4IiJPO/zVfeyzxDW9ScAkxfVfaFvrg2dgwerX8TcqgCdgzDr
ugcYrF8kPG3tAxGMX9mkx2+B68CfeGkLi5kD7kRpfxIJi2GvkCyPVWrD4GjcTU0e
EGFGEJEy/mGTTSmP2Q5m7NbJU7ylPZtO6/ipTLglF7a3BJTieFh07jhedIeobjex
BG0TGRDhgse8+LRdzOwu/isKyTYYht3Pn3gcGAG7N2c7/oSqWXstar6GTBkFbdt9
0U1qmwK5+KV8eakVCpNkrca4lso5x66PnEGjffwJyEBwWuEf78v12FksyW+sjipj
OWxmAmHPm6niLnqbYhqEus43RFbRKqdhHx80RRv92lN36TZfjljLCGfep/2IrWUO
syjEQDFAbu/ApnM7SNqWeejz8DitIFwcetx1Hz8OrF1fhzv3MkDuNiUILaj+OYS4
mL0G3TsI9KnXBP2FJPf2r1Sfvn1GOz9XP3jy+DqUEHalG3nLwkMP3rA0gvUdKa1o
tq/zo3Bs2JEk/9UvoXKGhm2WUD0a2sySqdSafTkENPN+vzBkgFoh+68VFgvTtJND
zrB6wYByjiOFYZ8oLqpGR3Z9quKH9DJeVUOA7bsLRZGqfgJnVYUiVjUb5RbtVSRb
ZJuV2hh9TF0Qh/FwzS8IyRY3jKIhUn9nQdzouo1jDmIcEu+foun0OlbzHQxFKBQc
KhT7JnHOq9EhKhd3GoG8hiSUW/48hOWgk/Atwp60x7x2mHypx/CpE83FfCu9++1A
HRlHkjK28/zyvCVEk23KkdDdQYbsOl3G/0/aSbaC80A2TddLXh7T7fdJ9z8SQX/x
vUnNMzWrqRmf+D29WMD/WceRjC3HjnDITuidnVMaE+JLdqTuM3H97wdlci5YSHtC
lvLEtAofCXJ/Af4Ej7bwITDGC02J23tabHKegzwVM5tdXyDb6CScfx5OqYadnq0Q
/FUVDsqe7huy+5zomVRCzV+TdEqyNacvORzqF/6Wc+MnRrjH7jEAB36rYUcBQbky
n6rXx34aSW9N/TDI1fDldGH8KLuLDSdiCEPsxZsdfJB7VL8PN+9cH4tqwn2YUWNF
dNG0k1kaiAMNeNfRuM09sC47/ON0x3PIf2rF3WoONuZ6bYhO6R/Kt6big4SW+ZcR
sInMimHvl1YgmU4t+j2F/V4mFAWq4wbbeD+kAl1SYjggraa46AvyvI51V9IMti76
jmFv9BCVEKuE0/YkgnEdUp79Hg1dJv84BxGaLzM0SxI0bosEbcX0rQocoB262tVc
AQz9908cJPDlw5PHWwmGX4FqxLt7cjlru8F5o3IlGobLxVmW17Kl8iJLQvC4ZUE+
uVkxmeH1h0HjKy8dpK9vjrd0tjFSCMVGfyRGn+y6NBZAtapJy7l5vpG/ABZAiWVU
dYWehEsNvJav1n9qSQhOh4z6nQe/IDko5Zw0Ik5Lie9bitSOT74cba0XrG9vSJrK
elStPyZOoxkcG7SLcRtMXJZM7b2PSomC/oLfogVc0ubl0q/cHM4Y+AnX7CTIQ1qK
7K5Iiow8K1f7RUPk2KfIy6k6xh/Jhcjta5ArO0gKCOJqWccTUpqPBEyoJ9p8Az3f
vhlvAdlZbqz7E6yF+pgVJWAbD5b/c7l6xwyv86XjfjFfq5JZnQsnPe4tRcIxnKt1
+7nIkoTvOrbQBJRoE3iVzF50TCU/pYBIHkqmK9I3pXsY+5dzeLyAECphV6/yc+BF
Hoc6w/DpiOqv3z3s5r9UGXx5wfMWMZz2TjfrlKpvF2fhbri308gI2g7tIvE8FyGE
GH49QSfOgkyex7fS47viNpk9Nj5hZs+xkdLOi/GTbeNp19gSDyeHC6IGK4WZxnAd
yH3KLkWyyjWunzgEdZdKy/cPUApHgxd0fW9yvJ9n2xOqvD1F4nf3/4+sBKxd5GVu
tUBhmLAyE/llAvuxljSNYC5Cfa+Nqia7/eLpAUHVFHSgAuZB2OOpYTb/pN11R8jG
oht/wvLsrRvzyaIqiySlWkeu/RtdW6u8afL4eZNekLlW0AiwMqYgaWpzk3giGVdx
aIjpaFK4KggSXwL7BesLJZCrXszA9Y9QkjSM1duP6YsFFOOA7kcy+0ldnFzk6hrM
ejO4nQelRRSVVITTe+NLU7PCm8vaIUfn84UbfBKDwYv7T2a0tSLPBE5syPriNpjN
4uOY76vPIC6Ahs6YzTc4QBXZIyS4syQDGOnk/gK/6mGD7Ww7D5rXLpc1KajIqqEo
`protect END_PROTECTED
