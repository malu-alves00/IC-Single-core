`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7YGfssyyeli4O586aemLa9q38ZCgydN+fhuqZ3R/53sdKg2vDHuZ5mwzvZ0HXkJa
NBGHOQivZrT7DvzYaqVcLsYP1s/yR7c7Dxpo9tJQ+Tp8Wb+5MDaliQqkJNUfJPXS
fdkOObN9p6OmIY4WkwLA78HsD4XrC4Hk/5dH2SaNQXF5WqqlaHqfH7GQT2izHioB
a6OxisRZQFDfSGwhQBsszIocCTDwP4Ic4d4sn2kqjqcX+uaWwsU5VgwmjDuIH2Ql
WDwflCgcjLdl2OKsIMjFIblXRlaypayNfU7uNIqALDuIK+S/kIUewgeti2kqjAy1
R3HxnRyc/JZcFtxAQuDdsy2/wHUu3+v93PTyIXw2TYxyvCQK0JZbhGhbRhqNvnjl
X/zrQAYEeHcmrTCDPEPdbF0SptewmjMz0FrAFbax9zzicHl9zT2yoU85C2/3B8Qw
tRRR10FjmhK82FHb8S9axEuM2dAqrGfe66CeZnLUBP2hd/qQcBV1sRLo0SBchEj7
kQpOTJxHwtNSCzVC2ss/gmVY2bQbkLmRChQFuJuw81t6iH4qsG00znMbio9lkJVn
OkSnPinhRDrFX3se/a1y6Omc/FNvUUfGLndeiRV2KH/3DWyTuvlGpghRAHLOvqt4
Nc2dFxWmbJwM88OvoTiasfPBVtOsPO4L3ql/dczzpkgZLlaZJYjIWSLH1ySCM9bg
KbMLJlMtd6uMYz1969ozCvFhxX4VTPk0KKr7TLMPLNNZfiX256eMghNZEAdTWFfo
GtGjnd17usyMpjLyC6WZcK4QSqf0dR1LhfM91G58/RZfw0zn2zD/g2T9AFBxSjjd
qqwxQ0Iwf/82bAdMMxOohx0S1/uZ+pyZRsOEWsf5WQyzsaDHVuIn81kI/cwvAh9j
7ye5tg6G8MnlwE2ec9OU1kN1YUUgqJ1Ju+bC7ihK0eNINfdcdNP1ZAJiv4F4mgAc
MEZBKIqgoqm4MRcN5/LzLlSNMeb8Y3cWe2G1JBKcQhO5WHF2QA8y6IQU8BziNuKm
te0tw0ZSbi44CSYyyLKXcRlMW4E0YejNq/fln+B+OftHfLIelYwsvmCAtGzaLkEI
pSSnlQ9fCCiyR8OLolfo3HCwFQ4PPYTnwz6qYdBZIMYLGATzvHhSe9hzFzzE1MwW
UU2C9x1OZ6K2TWInGTcJJ8+d84zBqhZUKYhYoZfe3u/xEhol/laZbRB5VfH6ZTqO
rnJSHpZUhuC3uLlA2l6NRnHL0Ee2SAij+Bdy3dKYmgKo4mpSBvX35QTlorrMJz/q
3/IZE9Q5qika5IGPJwnhLK122oEYDlrRkSwD4WEUQKg4Sjzidw7qfZ0pX2UB841h
z25J3ZdMf9YBwYi97mSZFaSlYO3YQHSD7ipA5rt05d3vU3HKOGjZ3e4QVLLzGTzG
ElI2+r+qZokkIrVDeDiy118O/SMPJn+AltxRZracJrFfPUPjZquc6WJIX7eIEo1S
`protect END_PROTECTED
