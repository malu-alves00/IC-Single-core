`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DqF6fsxo2MBcr1sUukO3pSmHoTZGWhrZfmSweU7iZaOmpERLPftq9JBIYE8blfzo
7h5LqT2b2nwV7TC6j4CQtBV5eqZJTYODgKiwoAiB4A0zY7605mTFbD6VBSuUYbCM
sxfopSVYm1iNgkSvG+yczbVV8lYcozmU1NB4c2vX1L3AWQcL7e+nexBjBU7qcUom
A45AytWiwxZGTAWY3eQUWExXAThSJLFcXUd8ZDw2doHYU/LcUyi0j01D+bHaDjL3
ls95izg5EYnt63WWb6Rpaauwchdc21wQVwFpAyDJMjCmT1NyxqLo8BCaIFuhr9I4
Am0pJ3ppmLWKqRwRktGbTOK65UdheyYOUuSQLY99pCV4n4KfaRznZaBpF4u9z40n
6eueRqY41c+AFSwrF1ZxS3hL3bmaDxPY8RsPiOhsgCy+L6SHci7YoWItuMSCsFtS
zI/zICGkG5o0FbbKWmaUbhlvsaMlaluyNFHlTFe9ZB1O/KB1z4VnmI26YNuTkotI
eMfJPdI59cxcmyU3EExeiQ7T60w4b3gwAOOTLwuAVA6bwlvRg2uDJnzOgCD7n1iM
zdakPHR6TsMAwkupOYNciIvu4roMkMDdA720NTGjEHB9m0gSBz/d25uTBLxknbJD
fNDBNagQjCxHCka6tAjYVNvxWl6MzCg0w7Si6F4piIzzcL6psDHJRQgvtkfqm+rH
r/llK+wXjccO0ANZsXzXHka0kjd9T7Sgz454eWCAeXPpaLMjNnnW4cCkZ8fcL0CA
OJlMl15Q8bP/naLtd5YPf4uq7pEqaeUJ58W/OoVgNnKJVo2pdYrjnm0vdqbQXiYy
BQ/0s4asMndnzC2Paz16WSu7Qq1ix2KDLmZbLLJGTQGRsU1U03DSWliewVCB6GTS
N3VIs4LW9n1cHZ9IaW48O5kvpBiS5oE5OZTbCzQ8H6K4czGU7lIvLls75Q+owZWY
tw6A6BkOwI3wakVgy4uX+9nbTczsCPiBQSjVPGAJPCK9mULDJBxA3jxMZUdnvqE1
EgA+yLwayJ3xM+lCN1leNfBebxNlzm0DQe84cnyf9WHPSVSjjeVYEWh30YiBDeUL
zSAIjFFpZ/9Tm/MqmQ0C0cR0oDhJqVpCP6XN0JMOlBer8M/f+Y4dqzFquPyzAe5F
6m7+SjTh6ndQGO8u+QkA0LQaqYlS2X+9tQM/By9s6aZc5ONXL43UAUqo0kkR3Yd2
AS/BItHXAPUYNQFfD4ISGpqqFHiW88LA374RrC+fifLCFWaxcij9JX6T2PhJjzgy
GO0eLvTcSY1RTngUb13WXpU9MZ6AIyRVfXBdoXx6d1c71KI1vbKDjEwPv2GA+WBF
p7izyu2xeFkhXbiYDba+780KRJ6h6luRW7UVrEOz8vebvQwrd3Kmx4x04EfeFSHA
HcojWMRKc35xIj7UAIJybeEvrXtZvfRqkjqA0TjDWJeBjnsGnaTknXiGxWTwg9Er
yYG913UK8Or8BVLnO5EEAapvQ4CyLP+wo9MKI6tjTl30wHnaHG33L+2vurOOgpjN
hq4pXftNIFEiACCeKrz6UIhn7gD9FSUwLfPtRWekMEOuJPETbijpPT6qo1rKCZWn
Z4kzYolTLL+HVakC8k0Wxw==
`protect END_PROTECTED
