`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sPui/NO9I9CMPjZIuOfEsUgxejFt//z6kxzmcNIwUYzFwxCVSj4Ifx4rKKWD1dJL
cItX5Nj/d7QvmtLqqXj1/GnN3aYESeLAhPZ8jvIuI88TdhMXohlVIRFKTrB7ATIw
mtYwRw+uo4MKLgJwT2I3GttmnoxarT3+GfnPCqrZmF3THRyN9Sjnps4c59WycN7A
SbaiP/pISRU7t2cEnDPRAxC/HR/OsMrC9iZLsI2g6tRAGhz3RTnibtIEDpElIyaz
OcCuEKwcnYzQVu46RFoYQCk4ix7V2+BhWEgmOQpO3clcCYkndtpaK0g+22kPipV0
wvBcflFWDr/O5QB3zBhNgAtSNSRlhIdmHU5YEZooUb9w5KYrxxKbBa0IiQggVhid
6MdMj5dtBFn/vSpgFtQgKsfk/59AObgNRQsSQbDX1z/p8XG70gjEzC8tTchLT9oV
+r5wJ97ijrpYMF1nWAFPbFUpwlXfkLEMc/iLUfiTmyGklVyTaenBhZj5E8cGUfwK
U3udD7uUfXd34GAzSF8tROjwAPrTjB4gtpBLqUVWDfZw1Jo997y4wej3VWPvRM6M
Y4iWIs6LaDW5TR91IzXVE9FiEWT1ytJ5WrQ3LbvLEBambH1+WKmmyEEsu+HWuhzw
8kijCPsS+6Hu/AIWF+BAMAUb1kmjJj5cqKEYIZS+3OcN4Fdh0t5Ms/L4HlZLu5KQ
3KqO0gED3Qqvki8Hj6LiCse7qub7LvAMksTWUBvWNFjHT2rlzW7UdFYBs5W8BIY4
LIp0VNrcOoy0rq2G527m1EApgW9KdEadAPu3YO3qPgPXWPvaq6LFU7XJFD7qWnSJ
ZUT4FR8jiEgKwvdkWCMDG6GaBhsX6KLaNSfl3TKXZNKpZfHh/a/sfxwXnWwkJtdY
v4fneFb2nZ0aPn7ps1X+anlNMX4njZGe203dOgJBdlsS/nSuF0nXxg47sukxeCXk
upwB0KivZoA2MuEoNIACz1gFv751n9DenOH5wRQvH3Bibl9mFtKyTAzhRcEU5Bmd
/svZ+j2UwItM2J2I8kFcpW/Y971LnmcUJPwRiZMakUGTkjoYZypRCQxddSMVYAnz
lTu5S5iKlsUD3MBVYk4i6YwB+OZVI79wondXJUqaDhrtOwbVWi/4I+oGOzbbSH3N
pjRaJnPWzdUA+G8KlIasrs3pYD/gAz1J+dIq3Lp6TUgE8yuFgDhpYdFV0kREx0jE
fakTpVdPKQ6RQqhsV6v1cspdS/rOzJhKZpSlVhEjJTxqp0GSyc2vhkST5b1u+4v5
/esqbYINMxAm6er0VTdziYNETu7yn+h//g9PTqlMZDPrYhEgWTmvJtZvKADfdt7h
GDpQPQKRrnECfMWJsEVzogT1c8WDVrELgYUKKzLUnL+/0EDsJOSN7wNTZPMoxc2x
pm9t+uGA2c9FNIYZuHaxxcHorSeP8AHPXcMq4I4ir/c=
`protect END_PROTECTED
