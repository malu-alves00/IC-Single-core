`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BxWKCo5yxtWP4xjZz0tlw2bKoNQEUrzO0Y9a4gcj6WONJZvQQ7J+qed9KH7UBsb5
9yENCB2qe7dOiyIZ71gkMSlgpDyQfTWDV+k5CNoDjd/sen1otYx4TBcFHScf4qYc
RCtYKEwGEcaWrCThHYx61SMo0mzqR8S2aLHKX0Py5dWGfSueqR5o/g21/dZPtq0s
JiFlrb8jlyxIJ9hAVPq08pmFoxncTio++rZXgee59q33RC8qzJnMq0a050jJAMt6
lE9OsvMLFb3F2ybcDW2aiBIM/AT3lX94z9Sg0sV5G6ZsxrpKW/be94xXOetihCNe
gzEmdLOmba20PnR6yQoXtdaaox2g4AzAC6cFHImdNom2sqK7ZV1qcUxfyTX5Z01t
RiEGvJtdLDc1OPgAhNKh4ucvbuY6sOKkZlSdvyM2cfjuHrl6xySWQswdvf9L6+65
2Bzpqd8f8nfM1gHdUqvUOOJ9wJMPKywhV8Qwy6a/Nsh0Jc2uTvTwYDAa3jRb5l08
zM3DzZw5vw+7ZpvbX8yvu8MJqOumD8X3dWWb0a1xPTuJFoBW4CimIs6q1Pok6WLo
V1VtIJyL+YrLg1wZJ9KKNCWah664tDO4YCqWf3OETI6Rrm3d1klBbPc7I25YioSZ
ILvxhOSoX/Cr6Ht4LCe84R5hkDO1JVgWklfAGSDyFTg1J9cC8C4Lk4CXnjmL7v17
hIhGDfmzfQNMZRgeU0oJkYgjDrOYK4g4iCxvnXJTalk=
`protect END_PROTECTED
