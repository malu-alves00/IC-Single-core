`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oSxm1kK/d88c8+Oxz7raMivIdEXERSRXVRBuHWjpRVEidK7Jne40Ao1LxkiZ8RJq
vxlunxNu5Lev/zbwxmNUIsgsyR+rak10g82VUlTobGklB6RCD76mSx/9cIHdOyAm
8GTLiZhoi07M15N5KHXmSNBnsLT4zSynq5O9WBCVaQQsuJmA31hgpqGh/DkQVlOj
T/iM4gFJCrJqWzVXRqi/U+ehATQPjwI/AfpVJXAQ2rVhM4xETsRN5VrT2daTWE1h
1Kq2+7p/3dsiBWwrFdl4eUpUwdOphi8PUecb7DfjcxaLdG1MyNgotZY4KezLWOt7
66N9Re9mH/eDt/8lbgcdM9d7o3HIOGbh1iHLMVfSfCmdRmTrZlanhVS0lWDpwnkB
XagEeRg30mFL97TTKQjJZ83uGDOucOKUiiYktwt4wrJB1bHVwDDsTCMCRNFrtbGg
fnTQMqPL8j9bW4MxMRDkTWguJdzQQcmCxAY4jpj1uuVmhuxiiZGxbBxImHxCQ3Ir
9Z3MTS1Esj36/t3dOjoPeHZPckuTaMQ9y6XMvnyHdggX68mGvq6As0NqR0c/foOX
hPoFQcIij97hP/1L/TvrT297RvKUb4KDcVHg3Zx16ZRXLLEwqGLtPEpT8BGeimDo
ae/DFOn5os3tVphviFcGrA5QtUyi4/daheotJHzFPRBy0ZE1oEF3mrpydu/rKUwD
VUsYLuAVqFw5LruDukCd07Fy+bZo7jn08rsoO0/tSHIwpBos5BEqLVUDOGfgDy8W
VW/6iYW9dOs2JluOdmVZmOoKWPP3G67xSXGGEzj4f7ESXgK/EGUN1q63x/pFZjn/
Q8iw4urOJnM2U+DJrwmntpuTjL/+T+gnuTvFdRD+6zPYz0k85skvfHrZvt/y06FM
`protect END_PROTECTED
