`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PxZcDtrF6vSW50jal5+G8QRDz8QIHlm/Art0t0XT86PXrRmjq4bijbPS+9zZTzDC
JDKVeMB2hzqBsOdfqAgfm/KEjTJabi2FieKGZjPbV5z8tgJ9qlO5kXSoi77GLbtK
AI6EHEuuyptP/gaQN2wqKqUs23qxHwgvxX71HIqfSzGLXEc/sds61guRrQ4LqSIw
cTvTZM1kUk6ZR4Y4gm5WMsDo1FGK7z80aXp5L7JQHwrvTqoRtF8MrYsSW2WPj3dr
Cz/cL7gQ4z7jLNsyaeNlqud/u1aKsU8MVARn9HxFNep0qKEenG4S5VfVQCquTms/
LxecV6UKptj8/G3oGoW1cz7UCd7/Ofouq7aYc8CSLa+TWvm6WpAkx4Hfv7aDeCMn
bKWsi3dDSMD+OHFcF98US9UcBtnTnVNLjWRn6v+M/tdAMmBJ3mgW4q3gGHC++n99
OXVW7WvsxZyWtV4OnYF7l/l8wWGox6TuRxze5CUBEwAGB66hU/0gI9FpmxUXRduh
6cgDpm3Ic1bHWKwQBWH3Hd0G/lDxwkJR6Rw+W/F8LpQEDPLf0xtpTe0dg06R6vQg
8lQMYZVhqjjDQI/kPQ/0qa1KB65YD5aG7MqpcLOi0UkSDDhJHmS9DI+xwrgVKAYj
pIDn0uLbv5HqvrwHSYB0B538F9jjXAoQoYQwJBpOjAipvMGl+qtb5+lxHchqjg6r
Xl4fMZZd4H4b+uUu2o2B9NF0mhUH14UOyCnOqAP9C9UuzknxDoz1tXSBuT5jkRRp
zC7jtN49/WKBK44f9vYbRjqxGsPVrK4YBN5oY3XelsYIy3x5JPo+9lBVFzYzMWC3
f5bKOVNpzRHfzzeNxI0N2+1tkHUE/CF5FasVIzvi2LnyZ2CTN5Vg90j+z9CZ6yf8
WF3OiOi2a7Pe8eHSXuWGpD8Rk0DfmMO7PiBg5MDKBCcQYbWJXwMyn1AFoxcgwROh
`protect END_PROTECTED
