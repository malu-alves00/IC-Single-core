`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/4RIY+62/JGo/h3lJae5Wr/Tu2noqdCYlnVkgqNdvvbPLW3+dlmyVBVTjHnhYyCe
k7CeEwj7bp0m8qJI90AWN6XejIAQXqSNF/tOjgsWDMfxW4RW2goNNBr8KFz+kBve
9guGTKzSxxqIh5fUaSWSNaLxdeoUt0yRD9bfolYLLL5WdMNBfHabyM9OevyAhSs1
ON4da7X24EL9w5leqBuvNzoU5Uigy7UYT5yjBSZrfotgW2u5xkT/UIud6BqKRyKH
RfOtOak9sRXkJMNwflt3G48K2NKdMes2GuWED/2Av181nWkrZNm/jCFi9GOJT32H
bk3yP1DTHjxzVHmN2uvJhIH2iZv2tmD5oY7bvvMr95st1S1q7iaYlSr5ezXuiQiC
+FdkxXYy76oaeJytmn3ovjLsXJ0UYpX9ChRBgPVcq3r847zCB230PFvHMTM2WSXJ
MvThRNyK5Svc1ttzo4vt01XwvDzlNcenOsK5/4k6YEY=
`protect END_PROTECTED
