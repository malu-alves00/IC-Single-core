`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FEfZpjHUfbY3wCAWnTtEhfO0QTnc9O39U6ef2FVL37oTLFU8wSxTT/XS6LjTVh1q
Y2LdOvmhjPaic4ZwUez8wum+up8F0G6Quo0PKEVRpNMP6PiJMMBKQmM4aemHGzqE
GhZr9JeNOXv4q5UjT9+IPUhCsRpGLlFqKTEGOUb8bUecti99hIMyrPBrUYeh4ern
p9uY2ak3j9LzsmdA93yv3EOVKyRw7+baT8l2NRI8QjZfInZ1upQ9tA/nZxVVL1qf
z2LhgVW4bn8q3oQKx6MjgLndE9KGPEi6yPHbEf8XXLj3TuSwdv1dIAi2fS/V4uXo
SQiIQACvf+4erIoLAcZu8A1GuxydqEt0Z+2zB2fr/NA4G60k/Oz8Hc/yvW1t0dk4
K+LaHw7EonkXCxxCwJkeOwjQDuQaVVhCDo2P0ExUkwaIIH7xsxxx3spB/fIEWlJU
e65ZqnTM8V7je9+r0nB09QKeQDomwsFb0t1a1ijtC490FjhBIDentTcbSFFSLVpO
mRbexZRt0jMGgYEk0pnzMg==
`protect END_PROTECTED
