`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
spSQw42M2v4LdGAHXZzr5z3LMzdupfMoQxbbK1Ap6867LgFkYfc57z2DcaoKGOcL
d1FZYoslcOcnN7UNkuE8hJWu0JL3qLgMxlytOFR+gp31Iu5x1Nrs33gQ5XQADE5h
utHLwfpjq6v00GiupLN7g0RfGOxdssLlgXJxt0kXlASWRyJHvSBciqcR7Ajxg87w
m46zZM2yUt0CLD8Gl01HjNA0lZRGxJ+IzHTEG5Vs7ea4FL4UNMsEDhK3UQR1Y1VG
iQyK5ReD/qxrCjAVpzQcLQEWWd0cEfI3F5CL+BRnNPDRmQEaMXdGg+FDRCnAA+p7
1vTvxAQsL+WnuHLs8W//YePS58Zu3L2NdF1S45zIhY+TvjahO09qyA+D6YoQK4OP
DJL6ZKm9mIDtsa/gCKMMBJVfd3lI0zSCj8fwAVV3Q/ewlF1qE/RHEkFFH1yyGOxa
SVBJvYA6BYKISkel0vibozK7kHnkpHhtNVFDmTh7zeMIBbu4DACbII4Yg2jYAlSY
AORa+v0CaME/Dtcff7VEOBEAw4ZWisglFnmDw60YFPJVw2HeazI3JC170XqmOb9I
5jjjVTAJIwLYDkV9QBZtvYDiOfgm02nSGpqQnohSbPUqIOi++rrsP25FaRHmdKqW
Y057xJtLIkcp0v3mCKARlApgWvVqqS44vb5/0D7g8SOJadjD88KWkBhJmLlC6wWz
HHh2dgBNozyQ+pEBF5RVTpvNYuUbHJjEF+qfcPp1dGoZwXNzNtB3VR6J90El3Edu
9lzu9CB5ovIQK/c/GQaJ/RlvmbeaGM/4UmKgrojhFVjV8PIXQS+ebBxNut0BQvzZ
kO9L03Imoflhpn/eWQE5W02N15cun+wfwkkgs+/P131jOJRDuOdwX3Sh8SRHoQUA
I3lqX95YRRcOyxVXe73nLNdORIWRT0YGy6M9qYUh5XtMwGbREWPpyDnu0BKYV/BQ
h4OqY+oQaSJve8dYljsf4mK3n9rkEiGCNy/TXE3oqsZ9hZBLVWm29byPI/35NtE5
WQ3AkJv+QK8ur//xpJFlAldS/o1IWHFAa0ntcdYpfwq4jnCTbSkH90KezTvxMzOl
WlzKptjn6DjIDnWlNko0/UN5GpZ/FRUPRyRwF748wYX6Z6t1uFnn1TsxsI8QUBaw
gUEEqecYiXuM+wOtJ7NM2vCGtCkka0VNbXmZZ+6faTbcw7jZKCKpIxdcX2BnRaDh
rVsJCvPzquJyRTabQ/eJIQ6ysKd5zOyunnJiALuKj7j5+5xVPxarJgbCjL7W3ygZ
hA6vcOy1QBXUcKXjqDELns1J0B0GYcbsHkvEc+0FG5ZiZJQQMV99wXNQGWEPx31y
WVyDSfVcIb+j30WBpCu1LA==
`protect END_PROTECTED
