`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9x9BM2GYrX6uNN9zVR9ruxRRsd+gva2rcu+tkFCmpAKoBF5P/1BJhU3xSBsFuvCp
dmZQQI/RoQKiJ+afPIX0V6/LktbVgO5ZwVijWRpccfzMLuMGbe0ZxnUbaMfK+yZq
zJKV5ls6L+QjEKkHxGuMGQEnmb+WSu2TwkJ8a9DZqShcPpI3iqPjv9JSfzixt1ab
dfs3S/QCwsfHPGsPeShjzXzvYj76uB3ZKma80UjiJ3DAJyEKCJhzXvNjyiOitu4+
N3XCMCbC21GXwvFAq5sz7JCUeE6dHXvJCZ6ocPeMnYzwWO2ALUaub8CSz+pdBcX/
vrl+X6pE+vocaX01fAci3qa1ydG3a6qoiVklpfURN663IO2JNUax8u2hcIm4x7Ub
QAPblMwI/zJ3rkaozs9I0hc7RJHxWDFvzBPd7tSMWyV1IfpP7zcOgdion+RV8T3P
wrWk5z22WSRPbNdsO4P7b5pIEeJqheGUhCZmcSYSsGi8ild58cYPWrdCqjMZd4rl
rqru5nnhAku+3uVYoLKvGYwJUPP8bUVmGx2VfpE7k2XyigBMclCthgHPpx0adW+A
gWJJhc3Y7V3VDXHrWI0ESIf6KQhJwG58ENWvKauI0XSDXz0xnVVXkGdZhHuRO4+o
2/Cvax04jiZopPO0k64sVrIHEvYGaiqAcXpS4EaJRRc=
`protect END_PROTECTED
