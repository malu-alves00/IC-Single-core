`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UGW2Z6D/qDZL4y0W6eZbeKxSiAWjtEg0V+WkCLwU3QtQL/p2MnP+CqNt+uuYQft7
cG1cSeRHBWorro0O5fxR5flM11fTnFwjSrh+/gzZTRV91hIGxgCyjRWw1If/DF9m
KHlgW67U2KO6htg4qpq4YQ15+VBlNO+c1JtGyuu1OgczweAbzBT9mpeAcoP4nVFk
7WOJ4f0ULaDzC1emzs0DOu3UhSGo255Djlt2Zvk57ARS5cPfSqGSf2QUBbFnbdKW
ABeJ8/JVf5j2um45gnr8yZuAxRctf2p2hTeJTO76a4tLK6m7Tpdhyha4UfnyIYxl
EjN6mQ6bW2TnJBqqIaGzPC0FLStLkOjl+rdS2UtnAx887J2TBZ/Y7nE+t6y9S4SG
u2wCb/EmyLNViPGywK59y6WxRyLnsVeH70kCGP9KJfEfg1IcBKOrM55G4ESjvvPB
0OfYeEiSliITrPqL4DyWCYQnJQEIw4dDG72LmLIVOLFu2eCOI/gpX3loZwvtuCw3
BxBeFO/929h6sBPToBR2iezSALl/EopT6Sta7CwX3JaIJlLo2Orf9/LBYjRXlLmy
PoHDweQN8gAFO9Kn3kpx6GVJFGVzqRhJaISfQ4hlwcbHdeXK1Tb37EKxPGqnusTA
FhrEbTGW2CFOhwQ5/CJFvGe6WGm7+i4tqpB72BMfyJ3eVEAzmj3n1Ar3lbYPMkgB
+QdSrgZSc9wMH1f9YOL6gWMD2RjeTSeoOG5+SG1H/9qfjji/JIpUfoEplt+WIOIJ
f3SrwnYaQmueYHkxQWfL4tlHlub5srKbzO3I1mZnW2b8Cz/XCC7LK81d5kDbrEWM
4k12OJ8pUpJSzO6BHyPCTA1Mr8eETMYGlpL3gx4kKVCzEwv8qV9WmhUG+qa66qH1
IssGB1OQ34iKsauIjtqvqFAyhznJdjUeLbuPxihY0Y8Ur1WZn7JHLn4vhZ5TIjeE
cXoPX7DqOt0MaAquN6XwfPXanZzZZfVH7g7dW3VSRtOLHxGwpcqm4fl5zF/wOAn5
CYMXoIjIrD2fnsK79ozVQ3bP6E4BCKxZ+MLOW9Q4xyNP03UgLTpxtxEdJjWZ4upQ
Oa8TNv0gOhk/Sgf8E1fd63AoD0qjCZZz9zFRlKFq+nBlivClQiMl0uM8aTsV/HMd
nNav0o8m0CZTpQETcw2ftj44DsGoLruSREujjkkZMQeLkpfeft4nuaMl2GiAZD/A
a744j8TJnlf1XEFlJKWx53Z7g8Rlz38LSfAqi/T9Jh+JsDs2hH3HwYYJlHjigO1D
aii5L+8u9weRpkbkGUhKje6l8SsycPNiR4nczwHd99/4+V36O4Rxryx6Eo3EACci
K2r+dp/yPRuT7V2ulhkXfwJo2y6oGXTF6Ije9gnYVrn1dL6/Bwr+/MhHSHvgeWcF
0JWkS6efyyAe83cJAVCM1lM+UMxq2LUhTvMtXLhI8SXHN6RedJYeBRILn+oxZK9O
pNr92srmSNGnTI2a1iM+8Taz7VMfdRI4n/KzKgyMuuXCwQN2JlGC4wlSRMW8PTqO
AhLhCVGsLAd9LMmqmE1wWWTIXCEuf7gvrjcf7W9z0eaI8/PF2i9BHITJ9vl6NRYQ
Dkoi/8hsHNeCz9sWCiAk/+1JEIEvhmAa3D9EF7iThB4zYIqmBsvD4WqIT+7m6d1i
ugzhpPxETE92Mz3is7jEH4PfeFSsh4vtap91g3MbzQQ/M/SVOA85RFa8fRCFYr5e
gPfJ8CrXOEfV1lmh7V67DfRR1vGGCsdHx5eIRllNvtmSopMaF0dC2ErTG4PsLJ+y
EU/5rubLWO2oGNhAwTe6OJmxfkgwVeJsz5ZWI7lcmZWEceu0OD+RzkgSPCDrKR5R
EtM4z3v7roMu8YJD+eeqie8693rr4DfVM8kBbhvrQj9jNQDNiLghOLnlEF5Xkzuz
kHUTess5e5FBCAKJjQ/5c+M5LY3aDHpQIBB5G5bWG8Ew6b78+wFfxln/lW6Wpmud
2E33kNodrFPPvMgGiqtLArL4wmf4mjJbs5v6fQ5mNg90Ybca8Ds+ELeR7/6F7aFa
OF6jWSFOKAggMAzfeQNjHkRNNFR8OspZzo8CvJHIeU1+kij/99uDrXG0COQfIT4f
TDqJFRTvhRMMe0hk11c1yUAQpEq1buot+G3jQTuWLXNIDpPkHdWDqrwUSUlO9e5x
7oDGC/NPZP3Iy7PfZAjpteq9JsZbU5hagrDDKSQbYupa5WUmEgEl124t44AXtyed
Dxv9hNXCQTJbxeDGdsxrDs7FkFFfXSRd6QTF9zhKolkolWBy1mXzWoZH5xnZdd4i
EGs5OiWpTVoLy0AdY9G988rL+G7pAOUV6Ng3mO+C42v2hPrBNRD7uUYcmt3lKvGx
I9h3JS29QTkd98XLlBVZLbocNR6zvDCmsThjIY9gnOm5s5UrfSc/COjWbLQNpieH
gDMNWDCjxcSkIUMQl2H5K4EJAV8JtssuCB13P4oRDgz+QQaHqtYNe+ZcUybIxSz2
DkCWieaFlZWNK2d6oDAITvxvZYDQdBACopnxOpgSZqf/nCBQya3IMTqYpmeIjZud
QncjmBGdRFsh8/qPAyIvmFpecWu0FLZHJK8ilA8/5OOHXzGpKZKfIy/ossPjjrG8
Occi0Pb+4oQDgiptMH5HE+AHoYDZ0Ldx3212dpcXBaVeEMedDQw3bkWncqHOmdXf
Sxhq3rhguUpHPfFrNO3XXvcRL8fYn+zj/srXWym1i6jA24TZOb+3DIjureq9A6e4
zEvr6ygZ0mDTl3flK5vr+tlhQLj6ZqTiPO/xycjfGsVYEuXVx2Ob/tcGE25TOsxo
6qogDJWHirwycExjPm6oIdaURrRSuQRred56QemBRi0HyDX3ReaV6qP4LN2gyt6S
hTxK9AkI4vdgTDVefSx1zaKqHDk5nhj1sMgLgrZvrGiKgpnulBPZmOhsttohGWhD
NcNGHyAKVH/dwKjvt3OP+RWuSs/Jyl9GZGgJxCVHJOvrkMo6SwQaEY/pX1upHoO2
yW6UoPbNSfYRqta2jCwbEOyQUcEMHnfB5spHTMAod3EBzHl1VDIFqsPCKAkD5ap2
b9+UqqUCQzJWXf4B23MtHoWtkT1YqHpEVvBoGd5QZeEDOxShWgZ0+E0s+Gk1lRjz
ISIF+7DWdJkQ3DUQXaGCFm+Vkd3qkbPAvXZXyVzYqSDhPoUJlWBYNkJ/3tJHvgEy
qiMo90j5qpYM6E6emyp5CEfdKl5MuMyfKdTmEdLUtVW8Kw8mMhlvEFI4eAbBQDq0
OfPRGU4p1cDag53LBWP9pkm3TaLo0djJCPylY5827znJ8gVcr0Q9xulItCDaA6gv
1E+U8oE/14hXq72v7C2QxxWk4lplp9rT9JIXOlKjJqlNCdFW7BOMgeYZhas87jt+
mEzJHiBwc1Sx1g/li0J8Qpy1jyXz4XpUHNTFaipKo9pXWaNUHrkqPOXGn+YG4Dkf
7U9hFyjLAtcv8kq8OinpGv3W5wY5yJiJrva+H05VNn01N3RzxNr1igyvZx3ZtYhT
bqdtHmoEjQESAc1I1SbbTSDaa6jqSY2Re40el/g8iQkAN3BHZAsaZtBxTgnYqF/F
Cz/ZBEpE49++C68NVFOXUtWCZ+UMX3gCOoXVdfFyS3yY0R/oNJUSre2k+IO52GjH
GQ79uBXfm7Zkz/hFTiNpvchsbEup+/kNJx8E9sc8ciU=
`protect END_PROTECTED
