`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7HAUyGJrwOBDnRYuZZMeVm4yo89WBKRvZnDhP2nMvsWUlEK+9xWSD/vcISkxGOun
/cCaNRmJO59ICwZ2elQqoLMTVudrrD/pR2vhPiBI36e/kb8oPJwZgWwS0VXZ6AoQ
dek92T+FdYFiWHhLXFlxR6x6JnnT4Jg/FR1AyFhJ7xEUUChUMpJJBs90j6VLM4SQ
MF/bsCqYteSjX9R73iLWfR3DE1J2pXuiXqYqsJ2wGQqT9ygV7w8TWA5fHtiORl2q
I5Q/xGK0M2VkwMtOp+ylClDeCKUG+tOyJc4oUCzbERyuO3JG5ZMyIUSuR1kMWBcj
LQ3QOXG3Cdx19RkkwGK5/EREsExXfEjkyhhP1ojis71OOFbaaYtXH0iISpS8RmEN
DwVKHPupwRnJjGrA3uxWucMFy043Al5R/eVIGIdwpSjwjeIXKHZGbJKrAmTuwLTW
LUEI7sON8udJHg+NpcZGn0OxI1UlfyI+UhxWrgim2AmR23nq806MVLlx1cTyaYAm
JR+jvftIiZJrpQwzEiGWOimt3N8MJNslUss89YEDrgemZJOxRrQk5LgD49k8ZTkL
dMkHQkHNpx9+eKBD8lfKnfk0RFSfB5hspR6acDGA03/1g3hjg7Juu2n3ZGc8jBwS
LUGvGYIeo1Mi2LHJZP2wbxA8KNne3wZzmxcfbNHX8HTKIwvRS+8YDuwWpBufpydn
tlirINrl3eWl5rRHOqkHVNtjFYCNKEA+apwRTEwtEIiadwb7Po0Pxnrg6O0hyIZU
bUipJPkuSE6dvWQEgXnMYfcVY8+jQjUFoh6lYQdc+5tHHopfPeTyyh3Q8aY5xBUi
21b1TKWcHm6lS8/WdZL/A0mRuLTO6oIM0s6UgCpnRcjVqx+EXT24d+KS6MRhRVZQ
Jo9SB8GLQ4ISMzE+fFY5vsn8U6c5P7EVaqsHpLiC1610JtArrT/I4cY207FpODEf
+QqiZatmhOMcDSdH+HeibTYCwpvTtb1/TKyGPZfI5Ht1fPu3gydvJWKXTcOxoboo
i9fF3EfpoqPfA8d7QE8Y9gKAQJsre83QuifXYa5MR4m1vEHzT/n8dBDfOVbb84YG
enPe7hHxfahf83vZnpt5TlpjccQWJ1+c5Rr0Vxu1StjlCIvb1bHcBeAAUmUh0G6C
BY4TMh/+7fsYJEdIE5SnYJONDB+F+7YIGXQe7nYcRU2uViGusSC5+NQDRFNRnSqM
lujr4EbrRrq8wEdo/Cj0X1L2gzN52XKRVXiEy6QQwYO2pz7iJYc+AaxeB/2/oOHH
hOwBgkAAM5UxB07h3mjm6ZL/F/9+WCkT6dPD+sjYh44TFUHpmfv3adczSZWexTaC
j55AHAnKW0dvw0cv9KaWjhjSYqUVxDHYv1zyLPj+7bPvB6iWxh2k5BB4YPdCisar
CDSK7dSnrlfPHQfN6zQUT7zLCMOwJY6IFXC4Nv18Wy873lK5xEm1ZZXJfSJkTEi8
tebQkbYOjwZI0+1J21/6t1fajNyOTRKLClbzYSNTDYZgZFgqTgivJhdT+BemHNog
k5Y2tJZ0p1efq35Rgxd0yzhTepMtxHmkncZnF71keMg0LEfJfZFyJWLuUHbTh8Z4
Gwtt+hwdZ/Vm3sdo4V2CpnG+lvC27TYG85xnECuMlKJF6CgR5CVslUOUt9TtOp6l
uSsOALYzI4xVCCH6dQ9Izo8/dg8J+5mxKVa47DzSdJpbBdYlbSqEwVIOi97VRLv2
jcgRhhkLPDegLdsNZUJQMhYBTc+ZsMKM+5lA4zdBsNoE8831ziBe2mPUTZMijzi/
lSDq9V7HU/BfYYA0aExrXo8GVk56ZHHDB8meZ9uB3ne0igHxjPH7CYxZSrAmYVoF
U+ri5dF26l59+TOH8yDxShDzj6NygPc0dN8jX1ZvY9Lzkz2XGqwRjuiIRuOQsE/N
5Uwaip1HqC6kvPxHov+baM/Dx5x2sDfb50g2pGDTNEiiaH1f+DIyj/+IbFFMDCW/
5WHvzDeVLbWX/6d1ymq/w3+n8hpJFDcPwkfq+e0QiOK/5mHCPhZsIi/WINVum+uY
pQc4oFVafC5zGZZs/GOF0Wl0+PZUGs80ZIJfuDmQHWhLl9WsMsv3K+Dl0TcNePzl
dxkcs/htXc2GHmVjNbUnRtzjonFqb5HI/2l5/F8sgIylPivAw55J5exViggouR1r
coNwerurmltS1m2SPivHE14gQuq0HGTsK7rgyN9CgHGoeF4u2glXIH/2s2Or2LYq
zjc5T/jRNge5kxpn3DB0JrH3Y8pgCmy2yUKN7xgkqjvuy1YkGflOPollEBhxXIHU
fiaH2CWqLlNzZ+e54LPmqpxmWleNYdzUBEq6gOYS+sxiS115fGQ7dxzCtXb+3U2T
X7oo5Xwpki6gY8FQ/ogJVdE9GOY0N/E//gJhAaAhTU54fAQjthRPKGjLpQ29JwME
`protect END_PROTECTED
