`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dMor5vss3bkyvu95YATWeBRAtH8gkRDcZ+j9AlvKvq6RTO8VdAXokxTZc7xsLKec
bdhLRIay4zzFkpulZM3wcG1iIpC9P2bH8zU5hEyCrsoj+8dWenL2NdCv3sVW/If5
kjnwkj2YY9skiB6+a6W4+6QOJO1Q4MIgQT7xTsIWuG3iybjLv4hMxjJElwhIkRzd
3/mXiHM4K1R/ONwHUGLkFoPvmCEEUG1Ghva8sAHsz6EZLpN3P2PVj/8bcUrXsvdO
ZuKSZqV4dgAWGzyZvGlH1CRB9e4VHpKvDf21GDyq9LhpR1gX0Ijd+gAeTD91rSKF
Kb2ii/y+DM36d+iB24Xj15inIhdLXnnduRViGaCg6TZGIjdjQiF2ecwDNfXGCmU7
K6AVVCubHCMtjiYupCB7FxDZqS980dzzMWmIEo+gDCI4uq0lIIQRPzF58EzacJHG
oAr6Un+YgTC6Bq+bWH4ZW+i5SlrXxUeSZpcfRgKpaQADReSrmSTwHKACfmoC/wgl
Ep7e7z7Q8eInMAZQOATL5ZE4ZcCMMbchfh/vxT7teaY/24DA2s/NPnFRZGZG/qCF
Abr5RP5f+6jfHXSMpAZH3cqAuF/MQUJKRzllZhSOvyLwRzIDQlp2+obI/MiT4tDZ
7nKRXasvYakrcR4AifCjTLfy4kTme2bE1q/h2G75USLh0s9xg5IxznuXMBinRFG/
HCalJElhqAKTQ81fIDN0OSCLa4q+wJkthJvTvUIzC1S7k1O+MCEZVEC1mtt2TflU
ssFRff2VmarGrWwAD7WryHtqtv88lwOf7wy+ATcm2fJcV6BO+BhGrQdgUGfD7OKB
iefvrjerXtvPz8mhnW2tlxT7EJ59XGPW+OhgiDoOoXdGT5mYj1uA4fIUgdPYu90Y
3jZn+M5BCnKgKOX9uFtWuRKLUkox1sEXplM6JwFoIBJrttzpjM7/TtmvTXIhVCq4
PxrewWxzHT9c8xSTchNeG9fzu6YdsLygSJnWPoGiLm5rCb6g2hP4QeDJ9Xl1NiiX
Rnmza+hBJJklywMrjdaXNjQaM9fUW2r+SZBn5ZnEWFEmXWekgPPhF2J/ro8EfGtf
xKGsjNhkXz1CY/n+9GhmWAKIOpmQDV/mXWFQ3ua5U5Wak8pXHxWw9Z8vmi4AMqC1
rLbv5BQNYI8QNFr7EXoxs36gI2KXDXrf/PSYtfCuzZCNYzx9i6wP+8gvh+0Q1I4j
eU6AUKpiJSRo+PlHLZSKXM+d8Yv5bOneeLdX3vPBWO3h7zRpMhTx4Opwpa87DdK4
4TvZX2QJKgJEztwx4PxtxdwlM0Jb7NKJA4VyouVqS6nc5zrzFNHE1S/xhBUCAAJd
Yx8Nqhk1pJ3eJ3Pl8zlZHQhVmVEhHOEivFvEBjfXKYltx7LUWP1ud+b7fHoFDCzo
+Fl/ZOXyj7LXsYM5UJP7eCU3XvgwongDTbk5U+Yfd0fvdkIjmv7w0Bw4569JRIBy
QdyATcY95zQfPnHay/peQoCvuCaiPwL4exiCg5/WK2LhQeNKmtpsSXtELkuTRLfw
ihmf2EweLbp/qxQ7x5HYEc0T7X9ty/FjK0Fo5X1zpsEWqz77E96MPKlo6rxrYctv
vOrZrSwhGwUGGtc4dZ8ME79/YojFJC9o5gYN+2t1pRdy0Z6oQ4BUo8jn8KAFia7c
cAyrGMdQsnd48W8YzuH4hsERZEErwCZqEekzTQrTPYAnhWltMukb6fk43/XGnEGr
imb1fMmzNUTbK89yAZacyhb1ElR2OJAeqbk7PzHH8ZK8S8YOVbMYJ4SKKpJIXP5W
RKN/VptoCpLMm1XkN8INZnGp9hGjaF0tnAreyigYAjKR4Zxm30mWVGKA4w7yrLgw
Iz7J3FHgZWQ22UT7w46JAozB0miZU22OO4mfzAU5it3WyLNbkybl0Q4beDabRJXn
LdCMbvGTzNAaB4ki/KO0m3dePlaQQDC4g/5glLJCK4idAHEFfnX8EUIbnhhbsaPC
AjDUmrnRGcpIKRtK5giuQ/rt+mUOMXrfuJZSAgXh+Dzq4aci2pAhMzrXncWusbGt
vLglJDnYeLBjsYO+TQw0B//kCYFO2i+kji8WGW+t1jjTZETjk+iDXZ7Calg+fpsQ
LZfA7MKwNjt48wNxYYNlWHy8CoxiD9txJWIkv3SJLOBLJRPuGEBT2W/JbCbkZp8W
zIKxBOPF2vrLcaCSs1pR7qe8R9RJYDhMNK6HMIYpJt+3K/aFzJv/ZXJg1ZSqybBU
h85ZVZ7nqnNNOzPT7J9fjm0DJT05Swy2DKoDW8VNfoGF7Hla32t6HVz1/wZm+0wF
XA6+mnRLiW0pI4l1rl/0KAfyOPlKQKLMeE/EM+QOspQBuluKMKAEHm6DlFtuf4PB
ZcNcm727xwYomeYoKhwfd8oPzko9oNyGeqXC+xY7h3ePCYM1x94t2I0DekcFs78M
qdQhS9m4dennkaq0D76d6gmQ9Tns5ZXvw/fHL8lKIcPKKTJdHOzfGjZE0xz9X1bD
g2Uy7ZCItnpRSgDpaMBRluD9VQt9lo65C79EpQoWgT6MjFVOhcr1Wt/IVnfTlNNX
506jB+aylCA5f9h46YkX2BY2KlEiYP0UBnNiC8tjsW5yi9IfBK7M+pkhWDO4Rq+a
tCjqjkTALRbvXr2tLHl5zc+4EQdHFqTuAJRwa5E4CcGKsEgHsh327DDBP3YnQt3Q
ygVHuijysQY0pBp9lcqE2i7KWabVuC0uimZY95IRisCGrIyDgkgfMPtLSQsYlGjZ
DNxmH1zVgyx6aFpwHZaFOIQlJBvoZQlSZ20Ks0CiS2TDY8IATaIo6mzmjJJE2mwc
fgfHWYZMzMcuuhn0aq6eJBAn/lzonlwIExcn0WhHyKd6+KOS/V0i5CVqvIuDXPJX
WSPFTLJoFWYDGcHg6ebQJlVB6Qog0Y6pyQV7c6+MUa3GeSfIWY7WRbnCpEx1+AEg
d3CFyv7goa9xeSuXO2Kw7VuR0vi4io5e2QyqsKzm9WLyMwmGBt6crweXEPu8KT1T
WsYfw3qdyYpkm/KlyL100ThuTEeKJcuJeZfERHO5nrmYvGMJCvzX1+Jho6ws6nzY
eXIBWinLv4lwqko+IaAkemJu7dkmhLOhDypvyjJrx+FbYxlqz6Tr7Exq/CI/dtXw
sQBdzFQADQlDgogTghj7qtUiDKFvIZYuItq7RyOJNnW4h7xnIw+acJaHbmzcwb03
gsHlnzjYkSjOulpL7IDC4P5DQWIgn99ocFFtMPBiEsLzPB1Ix3HWJWMcT60EPybX
y7wf6mHCLonvacPnM2d7BUstBKHPWkrdOiP5bUopgLJfz2HkC4/QU5SARnrwgfDB
tE3wSXumNrxX44G/2AMYhhLA2JMLj9fQB5wYMWYrqiontWvvQ/AzFfkUCQeuPteI
XM7eCam5PF/CZDGOkT/BnhS3qD8zqEXQoW11UyjXpLY4WWuCoYy5oWy18vgT6qzM
K4N5WopxWMgreEIcCelpMHzPura3qlT8mf/zpe8wzr7CHaykrgnnOU5a+bJ8XqBM
kVnMO0k8zWULF39KE4zbLQX97FiAd1q0KfL6eJhHe+un6A2xhc4RLzG3jxjk7cez
vSGEtKrtre0yeXEyOAAeWUxfipPvOr/jraOZueEbWgSWeEP9nOfM2v/FvVKKrWob
ZzcZwVVoi7FPR34G648zGyb5jfRhiWDcmMxXROGMMVY+xdRf3P2K6PijaIemCtkc
R885NitEb/HNTxN1YGaHO70U3mkpCtTtAmEtTCLay/PkHEsOy6OnLWa/crit4m+u
M+HL01VcADLCIQeOb2h0REZNzx3fcMI0UMdRrpFizkXRkuWe4uC6B3ij1j4ITvoe
91ena6bPeUZ1PZxiRrE59UBsUJyYTQdFtIdL/YKZRc1GZilaqcH08lzTQCjVUJSH
T71WHasnq2KT86vo2HOalopjNkgauFZeOTm2wM1Drzi9eBe/ofr0HIMeGc0nBd4H
xNyQPyDpNBtxgOO9Na+WPVyhXYm7Ss89GoySwP8ErQYh631WuzEB07+7SuKgbFZu
Nc4DsMsPhdX5sY8ABEGLwrsquTPx7jncNp26PGMjvGvLpLShGGuw2pzqvFLXT5Ul
+cFCQs8FROVXiSpHNTn6pPiUxpgJ5pUwoTfVkTfR+kL6yZ4o6WmdqSrm8SLZzIkg
bzpbNlP4O7IiSrm7xwCviUdViYP54RM4C0mfc4Gzn2WqcO2OhNXsn8PGiHE86iWp
h4qlqpP3dFg+wsne1iKv8IvqDer2LKnJj4mmyCSMsPdwuLdgeIdGXZrgz0rS0ffQ
eumYCT/pWaC+JM/3/3PGZduAx64f/6H8I9DG7iLsTvzPmJapK8sk+vguhh1YZizX
7DSIxagloFsFGERTe5db2tSgMSbQUiMMt9aUZs2nG1DbkHuul/s0DpDD06Gq6GZ2
A9BDQ/6bh+MTCwsWD26dBEpi1UlspXG4vpHPzw7bEpvN7pf4am/Yfd1EfT2YRn5c
MdGCevuHIocdzngi3ws9F9BMYah82X27iJQTfln/tqVBq0J8wFQLIMD8PkVkaQL1
MSyrNb5IJy6tPT5TuuZB3PSpDdJSJy+9YpAc2ttxzVK20dqcv7XxR584vCrY8T+U
vtxo4WOzv2iLo2aYXm2I/l7t5xDlAbATN974O/aeyGo3R8x0H936aYjc6s6DGnEN
jnkaRifvGCvqw/NBUnpTBLA7SGeSJn6gO+6Z5PFXj6dHg4Em+KRz0ASTy8zRAgaH
OUxrLt+2lhGmkd47T/gaSraRoQtKWtYYGX4UufQKzgU/b0yLJoNefFXJB5qi1Err
8L+NrTV8Pi4YiSdFjiyph1fn2W1DauF2TI/YrPBJW8N6EyptKcMo+Yddzv+4sR28
/ZgtJPbM9v6gBETve8LlA2eYUUkvmgSgssPYYm5XepDBGYAbuYjX0gmdvaqClB/l
zMXTEuR+D5JuMKIfYXnsGWcsRy/fr3Dbx/jZBiTT0YiY1uuqag2ucQbgagdNCo/1
PCfEsKzYovPYZdM0/+XfxEuncqVMGz9gm7uY6KafKB4UC8njMdLiTIZ1RbGs5vDi
nOLTCq1aITUHGoU5VXdGQUGAngSZUX3HAtcQ+QWHJwVljYFp1idPyKJkFQJWI/1R
38ZRGmuWJ+NUvC/4qJ6jI51+C2/OndMSQOtySlhqq8lovp61ZpVlMg6j5wdnESxv
pZah6y4CgWGYa5QsSCvwBNzcR9HnGE/76TVA1pPfhxW02JiaO67IAS2gU0YR8Koc
S9iA889La9+UwBxHxENRF5GJJQmkBO+nEQJKvosJoDA4fGA7gl/GAFQaP2FMTWIx
WXMrHH3dFtfcyQLPEFW//IMVsW+2HdHiydiWUdW1lUhV0oxaBxe4J6lWeTTRQcSL
zoXDq4XzL7WLoog+BkDcDJVZdRlZ+ovRvzpDqydQpvi6eI2ZkGmKf8GeLwKu2Ze0
ztW1JOb9juHSfscPj7vLh4W9iFtXBP1LddYgoRZhfk4Pwvq5etOigEcGCcwJWeWN
smC2ZQhyp0orT+JSbWUI1BfFwFHPjbVu6aSoc2atkB/Rdi5hN+Ak35Wq7OPRx53J
Ah4gO0Dl04IkuMnhsKbhtdqYxEzSmwz9s7zjxrkpVr25MmNKHZwcND8rAltWpffT
qxiOi/RCq4WBk/tqy2ZGQv9/VHP3TL/gYn9faX6v2cs0CR5LEiUNnr9JYyPZWzWM
yM03XdROX2+LDrdg78G/9iH3TxdYAlq6b9fDafM8Qx1uGGB1M+8oLa7wBg3vQ96V
K7GoqPPkbggQtVFzMxLBTz5rvpra+yXGIjB3dTCPdoZvfjHnI/ow29t/dxFcgQto
gGSSV8b9g3TAihMvoNhvD3GLVmtGdh8e5PTy0q/VmEqyTg6V2Qf7q9J3dO84IkuC
XzSCi4eWAv9aZJoK946ko1PE1yDLGn6/YZqUXIYAyppg7Q4wVTgOrqquz/A9Oe2C
BK4eXcC06GZjZ7rwpfUOQVgGTRk9LztX8Tbl9CyZEwGWhXmwInADA8dFHH05csr+
WKrH2Wrw8xa1ykEcXdr/1SJg7dxnIehsAFn/JV9tfID0bTekBkk5mNWiafS16TZX
su3l9fmrRrgv5Ld2RoxnROtbBrPS/+whSkUUTJuayKShyxSM468ataYyCeto3zoc
ThlgNBVLVP49ZRJFBHuGlfrZL4OCmF2Vc5P879zguFIjvwBpPigwT/tyaD2AN9Cy
n20HZH5Sk1Y1e/aBCjgxsuoq1F1Qti0JLlIX69CkGxhGnzUqbEyTPudK8RYyXdL7
Z6LYDLtaxU3NVY7mUkX5q1TJ2WJJ+JdTeNTF+aJm/ax2zm6fpK5czXYZUr7xwyCE
KuKVW0EGOz6khL1fqWjqVZ9TAiPThiqIA+I05119YsJTmHGi2NZSqiHC+xo0EmDP
x6KWAxqfDn7m4LVb6lJopL/z1DI1kMlLnvRW/iktj97EaIVGxGAEWjb+AqVDZgBa
zcgzYDa3VIzC5tHt+GJS3a6BPRYAkY2ZbB/gdxuVKtsCBteQAAXa2xt9rP/ZR4fI
RbLJzTItzJozJRwqdbVudizccte0Zr2x04JqVF3qOtkRhD7TNN3KKSrvbE+Fwts9
2WfxV2Au7BvR+bRZ4Le3MYg2OAQGc9IRW57Qp96VgyHWJSIXHM68rEzZ6avRlTP2
M9v6ll02IhqFjyoRfZSlknlCYuGP374G5aN1M8fiZE5Bdxgrx2Hhhi6l9Cbzcme9
bjqHej3vhqIrST86I5vTi8wzAIPPt7shednwarj/RMrvQyNwIFWrFMeCBqzqgrUg
N/Htl839QMwTYTIqZu9Lxrhuxq4Fpo7GL6wLRzxHosKk3D1etBELT1NffBm9rM3L
RQRvVP0cnhWgDrP0pmVapQ/OPxF1kl2dbS+651Kgk3ifA1esTSIlVSkIrJvzRYDe
xHZR14iB6gwjpNOEQNCNQRZsP/1v/5LVKGeH6zC0VtlHueCEXAWhEGjMjreTux1m
6xG4MH53tPMNUsFhzTOmpzW5UDqZiUCval0L/ZjZBzkG0oFeWiC69vSlJuynvYC8
XUjEO1AJjwxa9sU92Fz0qxg3tngt9e+jMjTezyJYGt0tYy68B1pI+86zslRqAcVl
PYgoeFNweU/nu9oJ4C+tSXnfm7D7RDQdJ1a3etA7kRdZ9Myr6AJIUUtR9ADpwfuX
wUSp+DkUvtjKwq1Ggg1hodx4B6r5Kw8lUB/Xu76TFKrIjh37pazwFDGZsmD3IMc8
LIxnszSE49bSw9qzc6bX/625elRb5RaWmsWCfcCHHcp/nuCXg8Tj7orC/OjI76gV
q07VDM4SYuiJPwZyk1sOD/PI57CIHD2fZu6tz2QpKUPDB3CFJ0vOCdAL74BLZbuF
q8j3AArZnxhLo3d9m+Q38RtMY61r5cX6xAKuC/kctYgq6uZ4vLCpdKEAFAp2mZZv
ZhyQytWLOe0SR0+lFASt8IkOd1bgfAM0XJbr5RNF7i4zehxTf+P4yws5SUY/Ga5Y
IZcHKX7y9+9zyuAm8afIkIjjsxyS+PrM5wv7XMX4CypuZ2rWHMKWrcb8UwmFwvs1
Aq9CDe+kCQkZuQVtQYpmyzlvWowH3d1kORjzPUMnJHGpqIw8hPjeX9Eb+iVpttzw
EGFtYOAB01gj2/Tqbb3aKa6DqUSNAUQBNW+DKExyock5hix0rxAVg1edc2Ec08qO
jyPLfc3kGkfCrcTmnjSN0PPROYjrZWlgREIfh6CXmib3cnKBj9dHcFwKkZVVex81
8KdrlsLwX211ElXWBUCzWARA0B8Whm43JnTJRzZ14qdMb7BNG/SPk4vuidLyNKDf
Ul3taOJqM18t22BQnacjUmiYpmaYzVQJg/9JJL8fw4T83zpylnKpoDeAgbtMsNsN
LswgXxfHUFPh5FqUazcqeVcLPbQUXyUlQqgW88pDZ9YaLoBRQVorAWd7BLcpOgaz
NJsB6w1uyD8Z3YzNmu71QWJ6hX6zO/36kTnqNg8VNmZ+jXXaanNJi/u05FzgGI2T
GlGhJ2lEUf4H4n2DjKrOYMWKOFPDzJHt6kXZiM9E8kxH7CF9FKhl8Ce4e0pRVMuF
MZUsgQ/88xMsRKkAgPhWVnRr5DnUbz5Vfu8Jg+VYoeYGh6UdTtOlDdiUsEeXYGwJ
6xKY2/H0Zn3BkZySdj9+jq0qWnTJrdTnhe9CQ0gtebKOLn4zjsWG6gH8u8dn/CwN
Y3pDi8wd6KmgYis88O4h0yUYRKQsawJok56M9002wTeMf+A7a61TKy+32kwBsOLc
JDGY5dqavEJQnS5cdcq54G8FvmBPD0M5lTm5ArQA8v7xQp0coTiIY0ree4xAG8Ze
89ucwQZ+Tt3VNQBE6DJsymi9LfY43vbzKSHIKC7b7xsiNIX8WVsdg1pDHFUVw05V
hwo110aVjIyuNH9Z4Anp6tL54TWu/ljCZObK8Wfeb3R++L5GZnHsV9RkhFHUctzY
FB5nnrri3oUTcrFXy+HcKygU32PkCaeyfa3MgsYIb6NLTnpm0v4w5R5fpw4y7oku
EJTh5/LHeLcFsVVzRihqnRCj8pX4KzJYaE4CDmjF3BdjjRyvBWCwvXRyVgb4b46X
q7xgxx4hbeqkXW1TVMw2ynagaTaKXjOX+RPqboHSms/hYcqGztgfQw16eowfuJ08
65zjT2+lWflgckTgKj+AWcoowmKCt/s9EhDjVgwlIkXPiO02OlmIdplSipng54wZ
VKrjUIxosPNqGwTYkyzJCx7rAsJwydn7Ay9pZ/HXgb+D9QLrNUgDiIAIGG9DjTi5
PR+jtQQ+IRWqLPC4jxh+GSGP313tmuYpwUqNrz12HaUKN816e/nE4ky92TExrTgA
b7atgCQsp/c9O5RufZIyDAgQO5W9PHZ/8zgN1UWrMdyECO0LFwsDC0D4QKG3lb/b
FJRJWaWSTXFVj878DoYnPbH5MR/dGseExe2KrsZmHIV4hIm1d2RN9SKU9iotsOi0
CMZ/J8DmYOSb4Le4391smboB71zf/G9x2uCSVJYJHvxuaW0dXspQ1Jo0v+0ORv/H
oZlNYTekGcU+aqjEGMK81yLfo5q739NXVyel6BBz5GN/lBqg2YZujU0+6zNhDUBf
UlJkvEQ7XML7OExuMDXgIaKHbBOhBpXqbKOVqANBvxG532sSMAU0W5AlR/K1/6Er
iCiQMEloqAgq/uXRpxFW9tXJVLbGJ1Ci3PAm2ogZ/+y+oqPoJGdwQdluHB6NfOqZ
N273bEeAD249Xd54gCD5WTKRxvQfE7NCEdKZX948I3c4tVB7YeTTeib38g3Yc5kP
PZk/TokXxx0T69HNJ0SPk/Hjmcl8D0DNb1fPZ/MERz31FS2W/Iur5q15u2X5yZZX
4uvfDFSWnW/vzumXQRuL3lwMKQh38RCibmhvBIIBuzDCuKrzaXhKcKCKGhy0Sa+q
jKespdiEpgwKshKr1fJLRCj238Ir+QWvmZ4FVd21hpUmdQ9m31Gd8t0gPgyZLiRD
/lWYe3ACJC42kIY103LAFDj+6o0gMAcAaXksyACaRwk6yvva0uSHhR4QeWkYwzI6
I1pBZtmD9Q0jHH6VpUoDXI/XBOKxVQ1vDOU+XryA6cVrt29mKIEcpJAnOA5XT1nI
PbD9t1/t+mU3IDHv3rZRxqhB47qAjrXsPrBPb0ngBAD1BJ1wyH2EzR5iQhifiBuH
59GgWGHIKDcB+c1bZAmbqwoSiQeCFmkM9xP7fkH7tk29vX1zfh/UpIECB14sCyRj
4aWgdoM8YA0pUaINQqxr4vnrrEKtg5FQOQV5eQcEn2IPPpgghZzzdHdMcxU0Zmeo
xY1jZqi9k7TfMBDZ+Xb/KkkSAo/sbNAxdb+S1VeXF7/ow3QtFHx/BiD8KEy+XIus
BrHWNvILRlY2cFxioN29gPkaRsCuWkspqm9trMfKzj7kOocwQyiaEFQl/E8J1dM0
Uj6q258CGbhboZJBH1JgjMmpSIm6P/SJy5/mlEDga7N5FXghlanO90n9TGMSpInR
htKD+Y9xuwmSt8Nlkq08s7QDva6pQ6V33ctcXO7cvtPJgRyTIUMLVcmY3R1IGNj9
bwRYohRggSEPAN/40gsaRbwsrCvjZe417I0wcB++8njiK+byOHkNggi9bcS76tv9
fMjATeBkn8sgFmN0cznurmzTQLbI+X1lu10YVqVE5a5O5Q/+nmhHvsagaa/BTAyK
eJdoT1Wno0+IR75dQGx8rvVs5KFWsheXygEXv5mAI5SGn6vjSkeywQ5CikCGXXHC
/6m7bxW44YeNexmAiuGqNeDCO2Qid+9IuAmXBCzMXFCTvG1KLltbJ94Jspg3JUuk
zMzBEIO/Aa5HyFwJLT2V625/pdMlidnwC+CTW/QLZHVby6bbuJ1kPWyXqryOB37y
R+1ipmtVE9pG1QxAfs75vAFLpz0PBu2mKHUrbjv10YjogYNxovfCexhbwjNiXqNb
I8NyNHOcEVfB2C6MIE/vmJycjNbY2f114cgJOfpW2QIrESlSfExYbZ/Ua2teVamK
lSBcWzWpq75Zq9Ehrb0fJalCbJ+2YXLdfzWIJJbE2DW1umo7xeVon0+7BL1v6Y88
fem6IDsQXN70/FFJSw8tsgSv7WQLV7FkZnrHW+W8qBDDix8PRlMXgtRQBG2wmkoD
KlSLXRbLP/221Mcb5QTHuFnsGe4Dd7/5oDjYzugYw1FnHYheQx++NkPXAQhrSoak
U4a0vHBcFySJ14GzWdhJ/5jJgdp0M8oP9Qce9cKXSkIcLCPECm9me8tRkoM4uU2R
RzfDTg539WWyaQjohs69dv3QZtSuC69EXZ1wMaxzSfl5WYtd0l3Myc0Nz0NN8DDp
e/OmDx9s3uErkoPR2EAJUM4Q36sj0argvZMbwW7bXQJHyo1qVtEbU7VFXLsugaiD
viLnMjRL6N/fgTDSwimCxZuCTwpe4YmjvyT7h3XJDZMAdIdgzTU4QPJ5782yy86l
hfzJ3orBVAJN23eWxbDMw+yR7b6E7c9jFSPvHlBlUKFWZ6UYS9lfCbw81Ohz9fpt
b0Tv7na78eaC/nz0vFej7RLyKnVicZeoYMpJy/IgJg01zkZtxrMEV3CQws+Rdcf5
j+jOsaB57UiP17KfLxvSSFgxZqLNsXxuQ55j06mADxyTJggiJzIwhzJw09jvGL1a
exulqqGcxW455tiYGuQYIscfRFEIdyaVtS8z0isRd4QGTZnJNaAnCb6PAYSpA3so
4rsnY1sLd5+M0aYWjrF7tnKy9EeGZNtcbBG29Skv9WJWfN889lPhbjucTPIOV6eD
YJisa4r4yhYdsRrnz1kyt6yk2/qpKBxsiDM7j7TQDwfzr7IuPItmdGDry9zLEJS4
KRbOBseIEC7j29aWedVurbwx8DNsXrcWqmnoKAtcXOPa+k907E7YmIt+rWnu8ocQ
8so7XUsQQnLLoxeW5VCm0XMfyWOG6irVnmg/bMgUIjRVz+PEbp2+ttlKUo7Fywvw
UdiHds/mYT7Vi/O63EkXzGfzCGnxAwoSj0wgoCfec8gOqxQ793BD8+3FU27xCsVl
fnMWG9WtXKKVJpGPaocBMXI84rffbXV3x5qsoyuDm7NgfnkdwsHLCJbp2VfqBpcA
9Wz7IFkX/D/bCsmKl1IFZ+haTahMw7avcMhcEv3SxX5Ulj/1AEkRAS3eb4eFitcN
bsUyRn03U9IfVitC0n3XiVUeBqV7/8hGFXWkPpaCHmEswtNyDvxq+tbrLnL6nLbm
jmboVuMsNz12FyYuDios1HDrztfGzEw31Y3rFMrOzQE2mDpDHq5E1bF2rnfJgffa
kutucXDbtdgYEk2DO06kDytPTYZtqMi3l8UFNmn8XKfUynW5BrBZ7M7yP/jC6sR3
WVPXvfDn8zdzmWaZTm+6N4zYsGAywvhpHv68P/193D5GSOCM5pCpjI53Ma0If247
szw/5DdIAC8wuTg3ITiRV/etHPqlFBNN/1aXAhVEExaLCdMDY1oIeRuHz5+EErLH
VvdkcZ6QnaUpfIId8+j+t1Cro8vcwNHJ59fu/6BK0kwIoEtW8m7Vp0K8vAstd55K
bNqfX8PEaYjcHIowEX9sPbdE44EKgt6/QFYIXYd/NcL2JtwVyVGES5vL5/WHdrQi
BOTnK+5sUYNGT/1zXQgpqgjx9Ci4FzBKYMUHYrDeZSFsZfOzSUYteF0G9dp3XT+W
XVNbs1jY4rGwyEl7iRWTs60YYKhuMpvnRNTCJYeB/0MmmGaU1si12hPmWfYRoXMq
h2cQK//+MagyoXukny6CXhZufgxuDR9pV3694ti/UCWbyA5yrwR/sxLtkxW3977I
gShclGRMFZF8B9JJ7cEpm+MIow1T614Q9KFF+vVfJuzxW8Cw2XyZ8PLoTx+1Ff2H
x6/m8teyIs/9j8ZEGhjKBQWiTWxrCuej+3E6wJK4bp+xPCcaQPLA9a/rQH7CCmc2
tCCoxnL9+0k3sUEculis4aIXdrJ9Bn+IMTDbpCeOCNSOkfo9xLP6lCP4aa5S8MEK
tQSR89S8USohvZuEkZK7mT7d3HKNsIphBGcV20Z0kh2X/O53TrZZWyD3+1eoEG5X
Q/kPJ9XFyEdX+6SodfHkidij7CpfO4N25+fbunRp1+uqf5c00jzz6AwT0kj8wp8O
p/VtUF8ToDNmZfC8j7AmzpKgAsSzhAOVsKhm+mfiDOR1o/23YBk4HooqifDLEGLn
kP0zPip9KHKQOSI3ePxCJbxj8DBCG/+T660a5TxoWt/UDMn6JXZ98AE2Af92BQEP
AUu2q1eyhY2SJffl/JiVWzyLEx3yFu4bGtO5PWtxttFhl+pU/AiE8J/dzVAZ00ms
g8OJRbGEvi14WTXq4OOVDy/3Z8q5WYqMoCu3XPHZ8nrgM+cZ4zLLazo8s1lL2ox+
1AW03VgypjdLzKZlo19v3c8xfzbfdxjAB8LBcwoq98g/0NFYEE1O8i4xGT/W1W1C
tiXw6e4ucXxma2pUcF+zYfv24S4oJ7ZwJdHYulpi1QfW7UwJ7JwZMZ7AFFoUJRvT
ftseU2yt+ivfS26lFvKwghh+eFDpaCwLxLrckviLvux6rciJUOsZO/K9v2sChdCl
xgXv8BRjdtd6htQWf7ECz59MeprGXU8Xc+kZBV9W8rkZ4ErR/E1jxQPU3k2l4r4O
cDRjqVuF+DjfBSMmS06ArPPvuLsyXQ8dZysYimXTbUObVW3QOPWUv3vB9HbqsddQ
T4T4Ee91v3MUvTwOBkGveaor+oh1teB8gH14HVumgrcldw+BX/ZKLh04GAEWIMdp
84TkKmhc36rIqpj3h/L62TuO2blcGfKOrw1WK64b3UBwl45Da2wvfC+YRG9HkOmg
2sj08BjWBtfGRIFa8KUfPDtTcX347Bbem3DIHCwGy7TBgtw/Eq1mZFsNG+AP2DhE
8KYirtLNu/+lLpLpjNPCn8ynzQteMNRNrCsExJjlsjqzF4tM3E+JLyceMZ/LrRlI
z2djTcZKEWWmFumo/IsX4UYLzCq4u03IScn7jh/nG1mpnbxFsygVisvKIHG/E7Wm
Bcz8VzJt4GComs5GHkuecpfFGkIn/Gpp68lH27bqlLDvFXFxuNr3o1KIEg1CtEyb
XZ1IMtuNsC6ox3Xvg4Pv/cny8EvK84KDAwEwhLUrXikMvXfdneYOIzuxBvaKUX0F
USTV5VQmXC2AHGmoKZTUkXYy4X3HDMaeaqvo/B3WBA8TtVDwCqWydgjFjPgXmoFf
ZksDEU/EjyWv97Flnh4D6T4Iz0ettqgbeL9QPGohKJ7HVRQF6QVXvZFSbuBT/PUB
BRMOCIgszirYZNrqPyY+K9N9Vr/p/sNkO+DN9D0usT9pTgS+uBVCE09Bqgr8wtrd
BY1TrgWG57yTVRnvMRbt2suIJVhsKtJcXqQL9bToUCZ3xVHqyXFmxlV1maRYOiAm
Ab7RIcu8IG0fEvvdKHs0U4Z1BY5S0/k4uMEhf8VrwIq4qUXwPxAr1E8ck/rcjJGz
aLhRyl0fJhOlpJ20vvI5kBuGVXX4ZpqSK7gN1us+6zb3aZL7TNKyyyhZMOTprchJ
ZuTAPdx0vE6/wceQzVgyrfxvPi7AO1Z0RCAjKWpSP4x47KXoyq/Pq7/zpKAalwk5
J3IHcEWXWdPWwuIFh5y4VJZpoEJchUNugwhVQ+N3BQ30CiOxg8Tso9H7Ms5CQAxD
nhYQOssdRhYKPHcni0Jsr4roElioK0K2s9CM++BP9BaOgRGKEe2GBiI9BHAC+oHy
Zt4NrLEy2GZnqgblW/QqduNybgvuY3Dt+vZRqlqxqRDA8avJeuk4AlkeLHRQqAGe
wMWmESH96egH7hUMn87nPxt93w4FrK5P6NUzosceYjkZqOFt6NYUDZwxtTbgGb56
q4o0eX9qaw4VmF3fcqoQK046aNYbXTuV7ItxCZIzqZE0c6yA2fLFs2uy4RUBmCRo
1RMAF1xro6OlLISftg6MjMbmmUxJ0T6jE0sGlunxca57U3SHL7quEzdfFDa5D4gR
NK/0oR4pHB4UkgNHEbl/FJRufZxqJs6FTkmCsjI4P48Goxqq9r/HGIgOGHEYM656
ZKhUeCjKvUBmRJ9TDTFLC/Fdb5WIYoVOMphgjpWswjEPgKbqLc6FoTDFA9uLFkS+
LQFoz096a7cDTAWR98ubdnJK847CnU7SZwpRWn/UDRTeYle7CJhkF0UwOwYU9WgX
8/P9GDtbaakDL7STOhQUNFFL6wNJ7laQfTI8KbmZxKbad1rVKX642NB3Iu40LAX5
nVOjpENoKjTH7fdKD3yYGMiCo0zF9Rnn1+BGn2/TiMsNkPlqLAw8/qKSNpOlycjN
wCggjuvUzEl1CkZPszVWgte0I3O2YFDVur6K9+nxbvxDVBvBQOYhtijVBxOhPvhx
oXxIjLYmvMWwIMVpEt5rMF+yXpsJpiyLqMKknqDKqoJ7PQwNXALS7p+8B3PuSmp4
+1OKus6P/fZOZbMygXtQq4/dVVMpUHd5LKlW3mtnskDYnBwl9IkVFMXKrx8eWjNm
uBdDiz6FxH4xB1ZSD+225zQttDnO6iGGaQiCM2HbICKLcFCS4kZO7lXkeGSIRRLT
6mNSdU96EmutsIyhHerbcGHGjvLqUyHOp24toHURS2oNe0We54DavajY0nJfPhbA
6HokLEwuzD795nS4XB0D55u7kKqdVwUfVK+4yx3Qb3uOIlqmpJKj7y2LmBiVQLTa
O6oTVeZ9zkbce4Gsi3jw3XgMiiH/uSlHfac2bZdIwYaGZfyrwgdoOomjQB2un0e0
PhXa1cSLvxMi+KuIaIO/D6OQyNYjfjRAKjhJckHzfhHpjk5a79FwX0Bo4bpAPyJ8
KAoD+yO51PfG+BU1EAy48UfcgiAmY3h4LfCCn0ZVyYwpefoav4nWfjYJcprAHTlm
T6iSUIqysL989tE/KpZa4bfgZXJCVqn7aGT8CURpun3+WFURH8Wr8PupOPFbpYJE
mrpZPNmPjDidHYdEnMU9CH+0vSjpTM8ejoRWN9sMVqk9aOJnif6Jr2WNq+OSma4H
2FSgU8OHGsnHxAQEWlzIwPIxyQWVKH+PsZGhzyWgZQX1/R0M8BX3FaV0x3UR3sNl
CIBkfyS+ATgRKoF1Xij0eThGguEDipIsqaOw8DUqOw/q2DUEebbOQN/8jJ1RwTg0
bo9stLYpF1xN46Z5TTHHlXPGo3b1KhY5b4QwrHHx1tVb7zZT4A8MxdgWWdGg2ZOR
x9GSWjJSS+p7TF8kC5d+xqvOO1xeJP7N34ZUULvY5T2fuuuEySXyMHXtVNeXXd2l
DFvEE4S/br2ca9J6gYUgr9wOXPHVw7wxcZ3B24beTzc/ZRhwdOLQ2Ac07H2m6NlZ
K+olVWMLMKBOnlnq7YmxN3315PVzgmuE8naMSpIfSV/cpJbI3YNbY3DBaBrrdjc+
Ew8dyGCWGVxmStJEgGK7Y2VjRb6AYEX/L/6uAR9XQEKi2WItPSpCeKirlJTC5Ev5
XPi4lq+VpIflE7I23tI7g+81cJ4OTvG27V36nGUqV/QG/WYCaI8F4zQbmjHsC8w5
lUoP9x+0uFlnt6DzZJqrbqnhyznD8/CbD2JJwZiRx7yRF5sk7ZuSaFEzVORsTTI4
/BEBwvDgLjGkvovnV+fsaZnrk7pQiieSJlaBzQtWDVEixlGXe065jURCC98nT3vG
nj36Z5GrXDIm7ai49F2uQhm2PuG2E3B2fjaEoa/ghwwvXJQKiDzWdMdIgFKWBxy4
TJkwYHrVJ3ofRDHDep+D2JQCCJ4ndH5vbJreXWskxsxUQfAvJLSVHlNhEcU0294N
ib0EtwqkIR/t6pRSOS9d0M4d1k/4joKEAyZOJyKjKFZkOf+6rVfaNfp80QUF2oVT
7ko5yNCLw8fh0Ib71tmt3zwYPLiEfAZCqzYW7pZf55M9HIo2SFTpcihXIBUYrV+C
40x9FtB3dbg1Lmr07txSf6kfbcsCb+air3r0u5mJtSs25x9S5mUFuyGH068MrSVM
61FUcZ3ByQwABeiQ7JpqjTy08yQKu147yUoELKGvasZTvwrQDEdx7FY8j1PkuF9y
LytqHUmcszRemh8wuGkB0+yZEO65ENnhwgKMNcDjp15awGVhF5lkVqhrKo0nd+B3
zFAHmz2rx+ZzWbDd3W4l1V+dYai98QPTKmrCgfo0dr+27e/4OmdiofKcD8ywy2jU
NIYd1uFyNUKoYFYlFMEM6MN2pR4ZRZZe3EQqiSbsPQY=
`protect END_PROTECTED
