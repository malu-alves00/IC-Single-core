`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EX2ike4n1nfwA3IKmYB9PqOPrBsvm1hp8WtU1cOuFBo/MrP80XToZ4JBOZMoyzB8
kr/45cyT0eHz4AOxqcm2pBXBHTmH47q1pnLoxzX9OKyrMb3BesOUlV2/CzzqPeyX
JsVjdLrYt+NE9BfPk1GT5eZgKKwiF4DfR5V2WT49tvO3q6mc3ocdztPRlrnQ19iw
GR5CLDsMrcoLywdVIoAI8fq95Xeuj5E2Bkr7HYV+Hb7+bs/iT792KlWWPfelYK/6
Ir0caGp+Cde46fzzQ8uJKAqvQ4Paei07kVy2it9EPVOgwZj4EOYtk7hACQFb69qg
CssOPqezb5Ic0Feb+4YL9HfCgXNk74vi+cwTPIrAisVS6qg5+nJCxNxu7MAiI+8s
Zbcb+DoHTp1xFph6PrnROMau+WhN+dxgPt70duIutE9grQXkT3VezdIrtTmrYPIk
LJqtrUgtKiH6Ha11YrPc52+zDNU6G8Tk+taEthkZcPRDyFKusvh8ksfcPAcnKiHq
0eOklb09SVAzOeQcpLWOZG+/fcN7I8T/GPQqqWbKLscBZ1Em07Us7rZKGewoJ61I
x0rHga53hro8igaHho17Q+2wjFPoXsPtJG/PHFWxo0v5FMNTHMc2BQkgD+F/rapn
KY1ff1y83Z34iXiB8i3cwWHEQAP8STP/OTmYOomrCnILkVcTI1s/B2ftEpqe+i54
rExsY4Ite/wLFm1VbE24CMkGEZXJDdhIejayI3qFcriqxR2cipTqX6C5UdFBbaM+
sQEJb6sY0MIBxw6v7GEWUKrEUJfsZKjM+phS0fbVTLT118tl1QnZiz9ebnbgj1oA
XAIfST1PjDjktOhSSHYHtIDGWr8wKKVl/Dw34N2y/XiAdxYicVBHAh7xaBXQbNBT
+4PgAX4g1CFGEvtmkE0qPJBk/VsE4toPJ5LGBovR1muPsKCzVVu78u3r9N1gB7cH
2xlKyrp9nQH/OlrG98MeUM/jFKFQom4paonz7zMzuYRkzImze62Ey/tPjVOfr4XU
uNhDXkUB9stH/MTM8/YsVYG+MzcLbsNVuGgQZ832hpDYIIzG8sctgqIPaHMZWRPR
b+bUGE13MTZzMr5QZE0GZSlNdBFEx+VWNeE89ZsPIorEFMObvwZYImrwUKGsfE98
5wYBvQmsK9PP8vPLwGyCI8FbTRww/BjiNdeWbAMcLkBxQx8Y5KpRr+QXqrj4L0sW
6io35wETaqG5NWXpsU29kln7BeR4966Q8wJvmsVr/Hv6hjzTUcgJQaVhpTwLHkxO
iqKNzkOSedzgNSYsYdO3p62YDAiAtwR0tUhxMHdVkXRZiJ4PzcNhXwTaiVCXwoYq
cZVefpFNca8Ndi4oQ7RUFZwDQRs6h146EaBXvh7QARf0OQqrqlCwrLeaOcCOio5N
jh/OrQn6O6kmt7tYLDW0XZTTr677XPk8U2gm8g87/JSmaYmeUIDOos7jPeTIQtRV
EJm8z5XY8uSgNRhg1Bb2tmKBiX5nZHzF6caEFj3vYqGO7qc9+nqX2kaCMskOVvsV
Fapv5yk7/ioaiM+os4PSnG3CohkFjgeofsHcBnrcNleLu7dqj4oDfmlRGvNH4pJM
jrXMVVbxgOBaRUUoDu61tfQpEq07LDY4CsWZi8q1TnkrNeWXKMla32ifRNBBJrOn
89nngHqnT1bZn25mHoSp78f4wMwTNiBR5DIisGfnJ6NS+A32hIEs78Lnfncegpj2
Qf0/Vk55mKSwyCq7xXrDo3d9a43SlThniYnjmXxM+DXpkQrTcvfHEpic5iWhSgVq
V1FfT0MLcT2ELd/xwmbXP5LNHPq+ik4clRtLi0euSO85cDyfQqRb8TiFPQzrqsRJ
/G0DtLIN2pN75v2lug9aDwkuiskKLGVfEch+XfTYswaDfmvXOn4ila/JFHZTTlx6
CAVXyvwC5sNQJtWtI9qs+Mx/7/r8cy+PVCYrhaPjD/24Aw5ZjlgJ63bSeJuu1htS
OA59Um83+p6wv/Jo3gHDC+dvY/guzByT0gthDfPxFhaiFgPUMwjWeZ+IKj8oanAM
omEIJMq+bqLjoKFrbXK9/ZhNA+eOqADMhH/sArO4edMF1m6haFpNL3OveTiHYSrE
`protect END_PROTECTED
