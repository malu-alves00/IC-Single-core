`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pAlNRpK2Tbx8dEq0RN8ZF6GlL36QLeO+TLz0IvTJYtV/SWXuxzp9yf193jtFThB+
32tVmN/YSGHrccciHSRbCUQgjivRCuVn3bi8f28PhTZTfPJ/W49NTROvATUYgKbQ
+wi9FKwdMLqN5oS5ZhlNCHWerROSIw0CKhB2H7BFw+gXe1RuqYBxlOHg3+kvSOKy
aDqLR9VlLYcs+61b5/irUAJJcvbX/CICFTzco1qt4rt50Ognp0koNz+FVolyVYWx
OCwW8N9p9UBfO0KJZHca011SrpER8b04VWVAdPPx7+hgJAKJBNJhV3Ebv0souXBH
WSoujomGEVElsD/FowhCXemAF2ZA4jqY6E4ayx2z7Kkw6x6Jdfue2ImQtsCE6evL
2Z/70Cje7KJc4rNLVxQYHvyHIoOyD0eR9Pi0gFL+0KWXwT2HmbiI6/IFaenFokMH
qAvsV4Bhvlxru8UjarLNVcEUnp7ZqgBXM2OYw5IE/05RkjCJj3GLpWme0Q4+zLwz
K5A/j1L0gxpDpYB7wUGTQitSnNh65/xgtg2B9sU+vs2+CRxsuFjQyTEE2a33gg8g
JK/zR3vNcD5tOuW3iO4AzN278AfXXL2oBjJQiCOOWgZPZKYHDLYLfrUERd182QU3
ANqI5JA4IjuRQiZ4KnoFjZisYUwAZfTYSDoMwAap/MTHpPcjRXpv4dw7kblgZqTj
z3DoeQe+dJRwKKO2n9FrXAqHLrI8xvOwfdym+CvLQpFM/fg6tEu9LDh5+G3fyHd6
tzh+tW/3DDP2gF431QugAeQkts+H0KfEK2FowV3GLXp3TUc/JzgmbWuDBP/cV+e0
qTGS3DUFZJMRHX3Wk1TAC3MAtQlsvBaOtQrnW6R2uS5rI8AN3I4HuFNG85K2GUdw
OPiejnG3KcHFF/g85MJBv0ovZMC9B1/ltE4g+VctlCk3nu5tqP/y8S79T8yk7UDJ
j8op2mrsW6fLYna2i7bt2JLHbDctmpKxC3y74ThMg77xTwHEPCwKWQHJPXwa930W
lNsS4xiJ9cgg7a8+yqfnvR08MBaqQM9jvdaKIOXy1SrvdR18mJG6KL7IGlRx5peL
zb+nHW1UW4LSWkdAK9YLBgZlWnfZN0l7MW0fOH0Xs7UOGQRrANwsznIiPgPm4fiT
+P0+ukzcdz3XjIY+TwW/CBhqUeg0CEBlwNLvl723Ev3ifnDORDlxQyh4N1KxPK9G
e8y1Pe8JmALxCUbrr0gu9gMsTQPwofc+s42cIuc75GQmsCUwwHiGHDs+yTVsx4UU
F/AXloBApWY9hV06HHd4b4uvwjCh25gmFkF//Zad+elTiy3YobCe1r43iStAmNyO
+jYuO1F9Eh7QceRIsiJbfFWrDQz7BW/RuYLhjQ8KDvwrg4t/a8j/uoaC52VRU6KY
pyp1Pa4qZp0KdIyNeUj3/PX9LDAPwTcSBDnYYxPkl2tVGVgq8wfmcGphZ71EiH/i
3FIWEwMl4ziSE33UoQnWhfpRcbCCg1qVu+xSZ2PnOyMHSYFmdxq8V5uIX4ZRN/g9
uVTTGQ8RRCbyoPvU4K54IbMP3ORts8jBAFSD+oocjNtHg/ZNWvpswQUf7NdRxkO1
TMJSAkVdEGXClDDb86IEqYDu+lpBSjSneLMM8gPy7t9568Rdg+rCAhg9PLE9TfiT
5FBjE//CiTbYA1A8zLJBQUmJebyEPu1YSl/Va3BZ9QDAPTctojHKCxRTjlM1ueg9
paAd6Q0Vwp44Q4h7QCxFE1rgk+DvRO+to+QOl8bMGLlxQ6qo3M8tWNcBDINV8vlM
xWJNJlxkVdzLezG4ZlmtjjleOKXZGyFm8Li/Zt6otouSELYBWQ4C5KZnaldI5RSX
XvVfLRwEfTbMOm1sKlceUC/lJsJ/VMs8eOCblhEXUt4GJG7rIhUXHcO2lypgmS96
4uPOLRzk4qFWrzgOmN/b5Fh9JmyOdiUZ3RvupPDnJ1hVg/JEx3bV/yO2C/d9IW0l
4SDz1s8OqmS8T23c/Oqg2mkuQ+GhD9ehbDO3mFtGs88Mc8mgOaZk08/QmUngSH6T
eBFAh2SSGSZ/mwm9/wC0I6UKZ1Q7tL4PQMmgq2KPVtnxEkqmCDjAESRnfCQaA8Zg
2l615ySX2b6Hjn7Il1OUi51BLDR3ZBhqUkMP8kafaeSB//Zc4/2sR2yKELzXxP5S
cfe5FO4gTwNUmFAKzdI/SXBMgkpbKXGk13XY6T1+UJ4BlOiSfJ5bjgXV7HgR/Ki0
NyYvegAASVLzocBw4d/J+E3DvybmUb5kaqPsfBs1Nu1rnpwqlBShegkGdwE0LLGF
22q2av9haEUFMuAi69a1VL0vpI6k7Xcq0GZ5vg6pnQDk73zJrrLyXfisEYg2xyPm
yopXNEwwUcnhbollDpFfrxT0bzuRIunp4zJuh9Qmjc5+u7JRzBR/aH8JEgvSlKSU
dIXK62UDF8233J4CPq6jBQQ/axMJ8nERVAGTyc8/WQ1UkrDQvA0fM6DCMVXizaU6
VkJ9X9bNJrWmz0NlrNEtC9SUPC0RTTHot3gqPFldpasdB4MeL9EeJYlZeJ24GyZz
XEMffxHJshY2X/kWi0qfdmJfJOd3vl7z1XI/XifyF48bkNG3cko1QJxe/vThL6ck
v6GoZRKr6HM9Pu+hz2ILlKBu2xB9pZSSfNxjFrMDHW5gT8x3UH0sadgT+rEgSMtx
cr/eG+cj4crJK7MtOjju/1MFg/H40M/uI147wnZ8OWDCLZJWFyA7AYqTS2cS9a7t
VPt2AB2iTlZhnZF/3BqrKIVNnGaYCn5QEXhlsoM2BsSi1/BeEzHPfTzCQEQMZ5Hy
Dha1QIhyLXAvVKh5dIkYaf5Gzkw965oVN421Hxtn5xsQOfRsPlED3UoraRI5ygP5
zvRMHdY9l713R2UxTyvXzbZ7wHRMFPNbT7RP8V8GbIJVmhVIhGYwTLc/tqycRlxG
Xi1ZGgOdpN+ZJV9kZrjoxPbWGKCLQnPB2svINApuG1CXedPpret4ZlmxvvKzKdc0
4muhAp9n3CqPfOiigsyQeQjvRSqRfuCUkn95gRTmHySM+SGFRkvHyymbqws/sCiC
lBbh5whUx3seNJXHpz+bmgCshED/XEsuBiAp78MMj1nopjUocrr93dYt1k1swWjZ
QDEPiejfXW1IW02/ojub5gig+YEzqrC+T5+hzpGkHOhbX4MHwrifHUkwdBXuS/Dp
4vzDPItOdXP20mbNde/d+VVqub2BDhKtJ0H17Z+TlNcP155/GC03A33fhVIM4WSi
VgjcD3/jSOODyK4o7dxnhW2LnR6JWdPOhVZAkhCex0Z95iSCMZkiIM64pc0NLJS8
7t2DazkG3fv0bMvhq9lV0IBD5SZuZNrPfT9mRwqKkjZapuHQ2DtwWRgzhrD15+HX
6jtJhQ40o8+nWFMU76n/oLiLIB99VaBMYN3tNSpSE4QlgElR0LNl5BUq744Xd4e4
YagwG3IgKHrJOvf7nxQM7dW97WZTymXlelrg7bh8Va+Nrg1OgwdB6uLdxRLTXOKM
IwazP5hDaN0oZwtTLS4sNbpQegaPmF+Q3Orq5ID4gbZF3GAeqA7dLzQMC/qhb/Fb
+P3kvQvPI02l3uvjb4dsUsTmrmvd3i8vOsrDWSiP/r/qsnS825k6vKKvrgSaJOiK
nGH8RqTMYtzOH+oBl8E9chIZXOGXoO3i198gyNjZ+TxUZR0Xlo1d0tmW7HI+ocWs
AMwo7DWIXSWguE1XEFJJkjRerUlaJtxcqY3ZR+fILMqAo7TnidvS/A477LlGW7DQ
RX9J++HtFtucEtffDd5U6gaAG+QacUhnrI+vOYbYudkjfoGA7a8Ehx7zcW7A90f6
d0Ac5qvbYA5W9I7q2Rgqqx1kp79FYwLwxmQGVrKJeTDkOn81AuvmS0h/1yqi5Pvq
ZBWEF3ngsGMHFmmsIa+hFrpjbVYc+xaeDyXu4Q4gTnE5yEvDLTLfapzRzXzo2vhI
K6xhezlu50OQho+cPIOEYs3w9VHCIFODDI5pcQglx1OdBCVdL7HayOZjE7Kt1g1n
ERHBzZz9HR0xQJUWReMGqYSv3cRUn1vDfcdYWjMy4H4+i6xsheVxT2srQETynch+
L34AaXgZVIDL6mj9OF79OnsDXaT9JEZPqT/NXCMZ7p/G0Y1uWdqzZXB07YCQ0Qix
NjQWDKjobEDL9dRaELWTRnvL5O6uhupkbvbmcQP5Uo9TTttkqLUe1Ff2mhisuf7G
ZOrOqpU/PC3VcOthzQ5XC5Yo39PxNsriHJCWpy3/39JxQ+GLX1qugDtf7KzQLFI8
YqbSle61T4ITm/eb59uA1qOEaoeJmkuAmx0KlGX5rbECbo/1h67I/2xOTcg/LKfD
jy5uibNotgFKyx+ZhOMvWBYXhomdDJ9nHSJm8qHvCWit0Mp/vsyqXlaRc+9dw1Z8
kbFPjhwSz2EJEMm0Vk+cvxJXQ12T+FYXgXvqEmlVrTCDBpxQ6gZ4KvzF3yEKDQqk
ya0zFY1LX8aCUVfC7maYUZ1gJLT864B7Sf66rEPaVuRv3BqEaAe3hc20QGc0sRZy
0meLzk9aV8Iyg/3IzM1x8I1rID3y1KK8xlMOqhE7zXHFHNjepwY5W2swhr5NqnG0
WIYijkH+DzKjOkGH8i77wAcAG4j4QbAK9xjVURgAmS82gf5DmjYpZanJPVMGvB4q
XIj+1PFDOsZYhBUjE4nG4sG6qfFjZoLHHjoOYkenv2g8mrRfoE2QCdjJ4VkFulYW
IrgV2rDwlCqXe9VY8QqkL8qjBGoU+qTL79LsEOtU6vVYAeXo/QdiVEWreCXIiNz0
Ey3E/MdH95xJ1K8nLW+sRuoYacpgbOs23WDyzdIflA+2RJxDYffC+opf9TAiaUuB
wR4VlimAtExA3mwULp66hDGzqArRqMgI+GGuVZLgvzR1wFles9Ni2b6T9nje9O3p
WPOCSjGM981IU02M+M78E5Ztzybha7izaeugKpyBW39ME2TktmqzSvYlOU01zzLG
Fp3Lcxd50BbVEV7EyIl8HGXAE9uPBG8QwbU6fBo7O+CGMyEOc6hNQlwr3IxJEXEI
mG9bOh4IL3b7kHsVjidrRJz7eipKsbA/9RB1xURmBFojbKBCJKIBWOOnMfHkiNaj
WXIw5izq5u/nZlRcjgaGmTAz/kOx9T3Opf6YHnOSBCym+20U36aqWGGN6XS1Jpae
nsXGZ8B3r1gDOklKl7c0AGqUXiaH+ZteuMzWAy9nhzKeDlgKe1oAsXBATn7Yj1c0
ifE1I4fDk/Hl/lE8MUSMt7UVB82OvNTSUC9xm/if2bhYsV3S4qMuGngVe859gwXW
CfbYpsf+1BNQoFudxvyxSdpVhmPP/lFCJFkT05vZJ4B5uOf21FER2my2JunxjEOl
BKjfbJ2+dq6BU+LVx9P+hLk8vxBNFhkXUDphNWwqfc4aMSUmBnFRm2Qn1vtv0E4a
BXX97g/Zt9hUYYp87eVezaAQSXsZzGWq3dQwWltkSec3RFqaqO6DLSAvE9OkI3Kd
mj704onltXmMAIwcYXjFjC+L4fb3Cep7tNXRwF16z+bfYtcbqSJHDcqAQ1yEc+8V
0pHj0CyeMkhYaVxSbyZcx6vzYI4O0sM+SgAirBWqow+nQboM6rYPyKpqGVT8pns0
YoQ1LnFiLEWBAgSvJCZ4oUePPbd9+Ob4cEwDwdpxQerf0HjlulI7KgLCGCTEdqmV
ATqmfls3hfQIQT5KpaLNcXGSa9rclHDNUyJQ7/rl3j6J0pcXLV4NfGd7QzJHLYXk
4NMDvYJZL2fs43Id4pg25x2K4rxt2xoefV5dB0z7+3U18fsb8lUwGRILshUJOkm4
9QXPiDHhK9aJktmZImr8UqwcTms6Eut9EZ1YT1mc3GpTSWE5GoIOSL+6o4jOMnbL
iH6otcgcLineTCj3CJ1Iw0952z6Wqv4nyjK/InSM+B+xnVWXIyILnL+ub3x5JV3j
ddsoXmTqrm31K3lP/Rqt/pe+Ne9wiCQ0tl1kL8McIcXuJDKYmP0/dy/a8Vda/DCZ
x1loa4t2m2AMeABtLKxpmAdquM62c87VeZ8rn36wQftmG+pJ1UZg5pfozu90foMJ
w251E8wiip8VrI0NW5QlXrE79SQ/kwW476maNMbNjFcdwtlZtJBaNVHDLR3eg10Q
eKPCKQxnjCgx0QCTQw3cCe6k2rNTkdzfWMdwMzzU2fivtwh70lPFBfYkKX4OtBeq
ktZcNSDrBTzI71cA2j7W0UEIWBhIT7ESiAKhD+qIJ+hxSMfbuh9kJo9QariW7f81
yt0HvVktsjeyiHrVPtrVLMPfGhW8yCIKTAMEhlP+8cSoYqvlHw35qYA+/kFJzkT2
1wMzdj9h1EbEslX4AdH/LSN57s3Ud2rL0skoB98M1njTQ8M9SboRTdFxWjPQTDeQ
nEBkzOq+1TwWR0YLAFYkupb26r8e3bZt2Fk+YerEsdphk6cLEBZHyZAFun46LEU/
3Up8UT/UcNvrGnOUzF4fpWyAy0Tzt/4QzyAprg/SDSoz4BK+AUc2n7SuUtNqmYSk
A603zidNpocoO4NuVbIijlZshAqs5p07+nAMdxVm2yMoHNXM31dL/UybZTGlWkAN
zgueDCYxaj3Mg65gixgHqw633fMvBpILxnV0qXs3tjox9FWHnZY7gpv8OrAHy0XX
4KtpfbyzBxVhoRqro3mRq9KHjzHwWXrFOoVTRYdta+s8ouTnfBKh9gAB8Ul/DhRa
ETeYXLF7rVJbvcaqJ4ilJMcByPO2u4eqTU2LvN7VxRkCdhwCU3eAzjZZQdC18GRV
9nKt2g/AIhIDbMQ6O0DFtghb4DuVuvIRv7+KeQC9KmCXFxDsW2LHVhENEe0tJIbM
ot+SVlQvhkQAo/dFZXyv1jCBLvmKTyT2EC4WZ/A5fyGEAgtvkS+8DN8fdKa2Zmk4
5bpskhLykozUs3zbWR8+UyFB5mzT8oKOIoyR7bC1K9+AXAFEGJkHIahCIAw9EFXQ
7k5fjB+DY6HbmbSo0e/rT03BXKjKZlgitpxFX+Iu0MQR2IaehOtq56WZzqQSa6iq
6FIu/SCkGKiLECQkKfPTy8xJ81QW/2dBW75rQuaY9PFN5N+fZ8xf03qiAzI6g6u2
jhLMaL4sbAhJ+jRL3HV4/a//hy3VeBLG+Zm31cimnTKnwMgTVYt+FHfmltIVwTk3
N23q3kudOn07/mTYlVud3KQo+kKJB0ftUlZOBoPgKcG2R+C9PkeitWl/KEPJgyyc
79YXYQKouTD63VcCN5OdwyYT7xi+Xm4DFNj6CFLsSCiY/2Q9cUL1vbAVVS1EoIpV
WK4H8DX8QK9krdi6sPMbWSkXZhJ09R/zdkHiCre9OfAmDIkkyEnps+Zgv6JS7esx
e1/W4nrw1Hgjmn5JhAUuMtv9w/wL++WH10leH+rJ8V/yKeXJjXsD70ildQx5GGRX
19C3g3ukkvAi2nul+dNZIOvG3LHJktuBNxKUiXAvIttiM0zBDpIHA5wP7MBnFG7j
+SMhRN9wWkSDJGdd4aUTtU2D8BSfvdB38TRH5Z8KjWKZDjwVz86t2cX0X+47Y4M/
AB/jOd07o+5u1GxaRcggOZwVy0vi0tNHQLYuRFgIgUV/D+vIFGlvCmRHDiyMahe8
ZeRBL7aa9cxjp/f7Jjg4Iq+Pa+j3OlZfja+Td+Y05w+vNZm26d2jI3ZbnidGRKzv
tpTa2XVJXRSHGAFcFHAL9BpA8C35+4m3Vz7yO50+w8/wMLW1zJQsvcPkadMc2Xcq
cBOjNbHt1A3EbH26IGQ1MEMjQLq5YoQw3eYsglqLprdvPnLawxa70Tl/P24SJCU0
mi8BVELDWBCDyOlgTKditRfwKBKF0YKWZePlofKiqlmqiFBv2WsFRYF4/ei2P7Lx
enX0sBEl3ddmdmbKdyVJbMgqUp2gVvIVQsQBPHH9p4uhYU/sRBffMjc+VbVZV4hc
JTxPlUQYVRNoJ1CNxdU9pVsxrKMXq6K8oI9EAZ4vLNfHZAZSGAthq7sO8ycX9H1J
45LOgtszVLKOd2rL6NHlxzNb23xrUPVVK1L4X6hUAty4LU7cLODn0dm78Qz7IjmU
tpyLTSz4ITyOgLUpfV3MF0VdHv9xwRlU9HMwDzB3kMPuTg5nKd+0QSIhDTSUkx+R
yZsjDRl0OUjZj3rnf4t3NUaBo6mjs8chr3HiQBpUw132ZcXjNnmgKu3k2J3rmJfY
F0/mmxSYxw0rkAz2vtd8i4ZDiscrFxro8JzahHVwFk7xXcn4UKsVSRkLxazA8eRQ
vAZFzSXetssqvektbwI80zzK/E/PPlQC6ssYZYxz/7TLxXnWxne/p3KwKh+WfC6r
6wvrBgty77oEmvqj6vuGLZVBtGuPb4iH0iHgWs5ufL9PxP3zR/1sxu9ynzUEGiaQ
Sf/BLw+DbuvytdtoA1iWRcE9jcfZLx8hgSzN3UPvC+VxLWZAvTNijgfSmzTMMNtz
N7k0GskZ/omvu57Z4Xo9f96e7oqa8WsN73wnUJuIeGASoEFwKpmJ8TqvvO5PGvEc
/nCCWfxPyqTvJ02cwVBRlLry6AmsksdRabdt44g4rYxBS/6OMbVj1bxC9Tq9bOit
K5vCWoYACoIUQ65ursh2pQT0a/oQtYuPQ2G3AG4cmupWt/uxib6cAvX1/OK9W6e+
t02VCiASt9tLb0aiVckjRSJJ268BZm/ubaE9BOCI5xTw+YBMvWBnBAVWUr53m2hK
WCtp1NW00XWLPkBkLjMmp4qOv3Ke6rtY3iBT8/ZAy3+8g7SSqZQm1lH2SxETU/XK
TbNFQZw5LcsuFeKqlc0QsZUSZCtLNnRpq5Nj+OCPTJGKar8eRZWja93t1RUOA3vX
4g9BaLznkqNrKftQYpX8YPto2KDJO8QUV5by2WC34XM=
`protect END_PROTECTED
