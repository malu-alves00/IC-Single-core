`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5GysiCIHLyg6SNCn6LH7c3HqIcITLUN1QVlsTrioDHYuQb+6pEgOK3bDBFNwvhg3
QEQHGYj07MoA8QZe8PZuwHVZbKgSuImUhZwPCZbYseasPsIUWT/pQNjhiI3TmR4D
wJGPzNSmtyuF5RmY6tgxqpERmRROP4kFFW+kb0UZ3goyJGTWF/uHubahvfKhlYXt
ufUOLc8KIVOrVKOvkIRbEhAk2cV2BQyQsUTH1cZDV3f2jXTtccIjfdDBQQfUc7Ls
NPOwIeJPraKzjZ7lzd9eWmN52gaY0MeJf1f1kSz6EY/9DAidC8Dwn/GDNYSimfAg
LPOobYYU2uPgyP3sueE6GqQr09FnMkZ22/TbSnEFYYoV9WkcV4R79iiT9y5VCtvA
8Bw8X96FLzrwLyAAmdUO5UggIBKyF5xTek/sOpxlOAoZBBqkypPEjsJCHeLYcO3y
puQsVE7FIJLE+6u8bDSegLTfZfvc2dbcDL5dpfBOTw9JnrcaF6Py467T59gReRWw
Ztf5+kKMOJiGH0762SR3AvdZ+AfAysceDnakRXrubi5dq2Z9fy35OqwVNP9WXPSo
OZkov7O21z+hZcv4nMRRTTDalDrjt1dfMJ72oakw76Bj7RFMmAWYIoy3RhWAywdX
9hX4fzErdv2Sa8kBg+o8wKwFCWBk1t1eMN2BNWcJ3md1giAXMaHLn83vzKM9HucI
5JDvWbYh9sT+QTqcKC6CFuRy3D3Y9wtyDKoKx8dEBBnZKOYalNTzMk3z8wZTOqg9
LZb8+TmSK+JoT1WZ0x1FzvOL/iv5FaO98HR+iBa+69SPPo5Irxb4p5CdFTyTvpXH
WlYkyYc9P8C9hUVgH6iiA8M/ejtAGWaVlzKrQ7kByevoopYR279Va0WMxKnXp3au
2WxbEtRZIdS5DL7sNe3zfD8Hqiy9Fp/HYw3wDfLnLdNka1gSt2H/ecksddbHRYTn
2hS1TPFbcQu/dZozAApKeDcWwFjgSGJJyXoHIq7vzO0qC3TEJddpsW03szBs+2iC
gO/S9gWTsAwP/x9ikxehTaRHzv8Jwy8LQMHGG2bHg4aWYs+Pp1ni95LJ53QOobDG
grH5/6aFYlFlJxES3K09NT1gJgusgmXpIJ4XJNfSpc+iG9r1RE4816Ol2JDSrNr+
/8LROdQPYtjL6qcoQWK/lc4U2Mb4JnVK8NKmZgHqJrIxEI8lAWhi1yhiub5aahwL
Dfa+CsEEYy8Rhm+gSHGcWKK9HUwiko3L4QSoNZIZQViL5IUaVY1zo/DQgtVqCEpE
0kapOZWEkgQhKeJ0Zlo9gJi0jnFCW4IZw7lfSJP8FFA//1hWD495aSWGcOmqaHfd
2o0HU3Ra2LfCk1ffdSsOwixrPz7kJX1x+KbAiDSKyymSy3fLL0PeU4+nftjYwNSX
DVRK3saNbH/g8HrVBsJajLnOdScR2ywIQe3pXSKJJ7uXd/LiJ0+G0MW2qjfPiozi
APm8B+GJs7rgGUuxZwSRij89KRHJXPeMLVUex5TcaOqilHFxvzFcCD61QHM+0Sbp
nyVRZlOUD4QTEy4uub0bN3VEZiIKIQa8p6FMvXvDSzLxzMRNnxwDY5pTrsCgYECw
JH8OTs0oPuZA2z4PKh41TRTjj3f5ywA4qwzpashaun+oEKxUuSWWg+OziUcgPXnZ
beuLGPafOtV26QcbnqJTmgQUUzVb3526j3RVZ3dSmsgyYadJ4emeYyeFsYsEAG9C
F18MeWVfjdJyubMOmhCrECKuZhpeDrpiZM8VQek5yX/L7Srhd5WLK+mXyuICVWQ4
1DiGzAx0EGYaHEwjrme12wRpUjk+nUTnixNezpnNxhk17i1lY/k9Q5oKTLq/QntC
vYAQKOjc79nVGkPwXWUSjF4qD9oOyBeE656kXPuBdkN/5c93pzV+NPtFnrO4tyHR
38re4eajjO92ceJCbo21ilC2Rl/KhPKNYq4Vmmn8YrkjuqlJ2kKWJL950jsJGKwB
tBBlOlk3QuBe5FZdgJ43IX4vSYguYngWjGBpnJddGiyWLH7WKG/v3C6SV9YVhFLM
mDG+2jakEtHbNGYIRWMk3D+ysze3MRWVCZeVPQHMqr7CwmdLwkqFz2h/9wkC4Uc/
RpoeoEwstM+tiY2P4yZTocpcfjq8ILg8JTA7Z+0AHdZeGGiCEYXFlaOESI7tm0m6
8a8tFl1uICwsmmBx7VJU5EsQUPpg1oQsIIfwjJwFaGLPi6xpV+w8oJlYHfqFplu1
5L0U/TRsQUDxd5cVsKlTqAqpLWh+g39r1JS+BkwaoBdThBwU4RZ1aBLN6zCHLuBm
cb1A8/2wZxmMTp2bdsKuMhh+OjlpUS+pEhy1ExVdcKcWfIRjuEhv2Wts7N3z6kyZ
0uOtoTLVN2fWon/f9hrz+DmI3Mv9n8knTHICnFJA0dq7vYFhkDF/lL/jLk//dSL6
gCALB5upTEDEpaUYvXuDhXlybaxIpty8LYD5z0SQCqzJdQXukTIzjOeh1B7eSKhY
Ya2U3AsXZA3UquyJMvxoZiStPKxXccCpocaxHFik0NGMsKhIh9C2D1N4yZDxx3K/
2v5+fwRIigZO+XWxtbLe8rVBBjgR+2Kqc1KlclxOW75u2ffeLcOPAbrOSdDd5Jy0
qVCa2mtR0c6RXc5uU/0AcHi/0t3DIxjz9LsuzLCKTS3CivwwSGrUmNdYb/i/H2/g
P5p6u2DdVZaF3fl+52LN2YbWYONjb6/JP3rlrAKzNPXkUqjn1xTpeSAZ/BzBq8jm
avNr83pj+SCw/5UixlOkLrGRnDVDOKci0EhK7RpN3b+UvtHNE/Buw8cgj58YcwpG
AsXIobuDtMxMogX/Q1nyGkaXMmupb24RiW2j5iW2RuoTHkrPh5fsOlOHGNNTtXvb
suhgVJduYhRmgQxBw27RaNYgMqF9VpFtvyoxEtZGBmyO+vA+cezVo7ckY6lOs/nT
+wvw/Zf2E5oEoXIGVUJ6sF3it+94QQQSFal6wbRV1c6MsDgvOHYc9OAM+uYWFZbE
cSU/HMGGwiydWHtpvu56pVPImR3gcPJthPbx+lyNJis7EO9S+pkjZexgaHbankzB
yUYNWH0dz6XO8zJASEsq3R0lrJaHWGY9vEfy55fkl2idcwDqG+wxkRTY3TFZwHiA
p+970xF7sWdfZ+ut+evVGTqEC84NpOHz+Pgzqz9wzduUZhjG+8GNIc8Lxj+WtmFh
qIiEnm3CJoSpg5142nuAVtawQjghaDOEwKwvmbXgN/uwPXRE+2pbT1w3rLlhp7mD
c3N04RWIXY2iaJI1RNZsGwirGtaGaAVRqN9c5lJF7VMaqWk+5e2yHzIJuVYQaGVB
Jj1v4bn51zT5R5aeDBlmHyWEW7dqjwOTAf+xR+oZ01O6ENf7PHly3nqQNfKNds1n
2QkO0kce6QIHkiyqfcvZSl2OQndT5+ywmSMUiNhBTv+jRbWvGRGRTIx1NAqYXfvp
YQsPEp++9BppA60USrAWT8qNNfM9v3CCtWv0u8K2AGg4Lfyww/3H3i99zbgvVqWD
yCKfChQP4Wf1Fz0wvPrFuhYNmcy8Iq0dcApxwmMxu5DVXZn4kAod8BiStUct4xwU
uJlbeY+fRy9xLaSfSArCt9L4NMdoC/REnZ1p6ejwAgnuCpca1zKcraaOu8pInTdY
9pePl+1Mvdv5hqi79+nHnvptmuZ93CCv7Dmll4QEcKXmE2YzdpD4B2IC69uSNG/t
zIF9yC5EXV9q8+Xi8rbiUGJGkIdElryDWwtCSODSaQobD9iWWIpEEEIVcDg/5/ni
mVOin7Bd/rUKmweptUYzuBkiEx5BLjj9YRBWuYxpuMbRe+cNgs7ssaTNVJ/o+d+t
zv3koLS03B/IqP1aF61rNO4rxdjGooGVgEdh4axWtAPDVynbMqD6gljDabvK9sNz
pSvpK6DZsIre9cJlS4SvvR8qHfINvkGfiag/+oOiGcyuP+wLhiQu+DGmNcJcOI3A
tjZVjHAZYLnMWmS0LdUMK6Z0bVoeS61KnZasP9UucakInayF5ypY5Y/kXNM3wKuH
MMjbtn3vdQMdnhCrWYm4G8QhFOUA68P4HaPQhYBsk55qHe9qp+Q0QlUBFax9ektd
i9Pln9hd8DSG5wTfQdU3suPYVYJt4qlQS1OFL3t90mwHaMQTwUBP26dwF9rVTOL1
2Bjj5ZGhOyAg7hFvsdPbS64Id8GHkubTnWXoGRXuSpbLlEXy6A+N08WsjGl4aK7G
JsJ5El7OKTahbDywtfrow0pVkqjcBqrVi4q+UhMM4E7YaaB+bwn77UWYEKQfe1S3
puuPTMVOkYbwLGWADfCIq2GfPGsABSquxPONAgwoisJD3zb/ed84WomyHFjDYxDm
utgEIR4FO7lFpzV5MJ7d6gkqtsISRX/QTdDa2OtfRUBbXTtJuT7HKqbcr4f86j1C
+KmnEIaDZED6NF826UmetRTkTU67Dur2asGhVDOWxf7hQaMtt0rdCOL0eJIRJ0vR
sO9//0UzSIXFtZTBNsb12x9VemSsh3sl+jMj65el8SFjMIeUotOuBtqGakqLvmiP
IeICW0an/d1Moih8J4n7TfWorxT9DQZLiO/6NMbrm7mlqEhSHVUJL1XzYBMdB3fm
LYmG9nzrNF5+OeNZhxuE6fi7qpDiLZ1F4SazrtHdWXsqoLFUcI5gzmoYuULEDMLj
wsb4HmKvQzjBo07sImQPYXOzbGGjhed5ch/gi+PXUKL4jcfmTzN+MyL1bwq8S1TY
l/JYGuzS0wsEZSUQI5AHfYNleK99+Wd0jFb9Ya/S9R9xkN3ijEy9y6gVSerJg6uq
Ymhsk3Fj1BIOw7u0XQ+KzPXeKYBvWbWfrL2u93HZOz4EX99hJoUPfWV2ObsYTxdf
0JkUzmrRPLIS4NSAeGNJ+20TMkOSV1oFQnq6CbbSVDgUJBV7Pplkq9iXFSqPi/OS
ttjpHgBojRrkcLXBhNcMI6/kNxAAb01q1+lI+Hi5kgjepYB1doEVapMarkCRD9xo
K22u8O3UF4SvIcmDMtLRhL+5EgqEz9OIhIS4B9ajgmya8PfSJOiOYGBgWn65HRGW
WB4+VoKXN8Dv02NSKNh/Q3QtJISWidMwRhB2/JOF3ZOlF5aEIEgTcnbO0K/DdpAg
tCJV1ZU/ZeptsuQ9oxP/Gv1Egj85Qvc8+8epeX0FtNBqTkWQpZ7jOzjscdQwApb8
M2ycAcwugDe0/9zwWdMNwwfgKgwhlCkhnbjIsoTSHo9Z/hfTHy3MbAJKn6W8ARxR
HWZ0xQUByx669WYNAyFW7zwGt8SCCY+TIuXt3FETESA2GqV5ujNQpJXcK6cg6pQV
aXACs3j9NYANX0dickvXcTzn9NkkVULPfT7r01hfBXUmbYq3SMTERHLoslJe83UP
rWNjDY95gPrLQ3zqvv+Z3qJsVmygg1JU8NbVUwmf3Zg/HNIqiah86jAeNSh6maux
B1fjRQrMwJlMMaO4Y2cFczzs6OFxaSAaA61wFzpK6nScjjX6K2tQUMg5wySTPFTY
JeM/ctBqmY+Z0bOpikzp1OwxPX030Zlqg4tmCFBjdXQ+5DQyd5bK18H1iYuTxg2b
T9AI1SwzcOwfgTHKyWK9YZFE9I1htBuiBri6hgK9rAhoBwEcCSmKKSMZktNtnAIY
1f2UK8b/oB2BWFIYAyYBOOcPMNHRO2arqV1Ox+6A2rluQXOUNFpg4YjhH0nDniON
Xip3/rkAUSbqQ4aQz/7+72vY55SWnXRzqBgYHnPrd+sZJoafP9hsqC12IxdQnW8o
IfbQwHAtSTh8syQD/lQzEnXrxJLGS6kXoOSCfRP+QBK21nRI01ZdfF7JkYz7t1UY
do6q3q5turNgD2xRaizC2qY9984V7S3S+00hkQgXL6dffA97Cij4K7J/yzwZuZfx
5SJ+Jd7lZd8MqsdD78rwjZK2u8cx1XZdE6wJ0abSFVihfb8aB5r4DqwQ7NiXHnkL
PpleKz3bmOx82pUK6fNaXcZjEs7glIAv6ueS1lD2loYUa7VoFmBgM+cT6qjiy3uv
6Tdpm6z019lnMAhJXMxomX2c1wjgxyWVUWLbaJB/j5f68mbddtA28XaVCMUuXwvG
SsWcRYeAB59nV28q8IexbVciCeGUvc7hcwLf8+Kagur50shRJs+QvxcpeVnnouB+
KjIREZhPnKNQUwft3LBcNnSmtP4eaeq0OjV7lX27f3dstp6qFjgUanyfC7lrJZj4
xpsdsVN1yumI+KGF8oOu5G19FAKHSBLDplSSO+SZVGPyWFm/L7RKGDOUCrNFmAY3
knNPUALeWNCx/EP/VkfiULK5X9YaF1FWg8J8lMgcEmh1eHjHfiZPC6pdb70Oyw0L
cGdmLyuqCo+w7LYH00KWi6IVUhYg/EnXOc7Ivw/5DdJmqH1qgaUO7hhPKlQC7jaX
oOryuzHkvC/yplfO+b1B09dc6crlh0oYXwGBGP4mKipQDIxKl0YyQRH4bEg13LXw
iC7K9Up9tNiHUOkdw5BA1JkmrhvcoquRT70eXtSY65b2r6ssznRRwWhkPj52wSBR
zzvvD6ERwDsRJqH7MCsYrzaS6s29GKJcHfg0BjdRmcRw1CHVxmfnWmtv5Pqy4fSe
p0cKk55ssiMwhB4ziOLS587qL2cjDdjKYo+iYxT3R+IKKSKCZPA0hhjHidvHy5LE
+QMCo4JcJQxMeN+78qXkCpn1AP9kBE08MuQOCnCugDnucEa+135SGGp3eEFj6FR2
jmNI+tAr7K5FBH2afQzYCEAJKQniyzcIfYNgriQRHXdrkN9NACR+rm+0N4XLaOyG
hvNXtsgd3avUh3nZ83+5U7GU/vR/2awflpaqPrhCjzOpCClMX7zE56QOfw3IOuS/
nlgkW+PRYqXkMCTqYTaTS8SimvWKwtufFN4t03jZFG8=
`protect END_PROTECTED
