`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
t95slHk9XMeTHbckg6nAVMeitjq0+PSVgQFpjF5qHJLS+nNi3q1aOY/10MSpD8l7
Rzcs54xiCfI4aE1g5eqvJE6msHKyqBwKJ5okIDD5chXVngcMxVaPfc5PwpbQ+ztt
2VTMg6tpVAb1bycL00M5rZ73jeyiQxRaigJW9rV8V8Jllvk9J6bd1EqEmuBvuS28
82aglyiZKz3JebxtaqnJ74C0qvSL5TrXFbo9A0jTRDwfma+Y5+A18xeiInUEG6rF
JjDfKE7Ug9n2PZFXeBHm+w8eQ6gQ6/qrNWXxlCUk5TGzUlfkiFFotZRJz65Rrg7X
w8JvBp5p5HLRqg6MLL2QHyJr04EgFDFpq7ctQDuUXXSSxFeyyRnj1tzpyEwgfKzA
ao6VPYQLX4xuFGk2VE3Rq3KaMaX4lXkpyzDzSRimLUNA2zeoCtso3ufbJgY9GG8l
PINTUffBMPO7MpR5ArtIjzUPwofQs0fbrh4w4tEj5BDbDKFyX5PKvG3qOEeoMZUO
1xRHkCUltxQMuKZOuZ/MFxkc/t99gvBabyLUxgT9HWH8me5PiWTsyc90p/8/PIOX
/RR46TXjDdEWNFl4zS2WTGlxxFgsyYwFj+tkPzSpeTy+wLswfpixJRdvf/t8D+uW
9gHT2nTnFbmJdRafjwn7JyoSk4acpIBYVWhSJ9yengGH69UclFyZJT/+7ZmoLYP4
JkrtZXPgUObA5OPLHYfrE1CYgrkV3QEvYNMM+ikVq5J8RRQVjiyukxN5CG39zmSH
v0DdDvf/7B5e6z2tfeITBoL147d/EGGjH3mTDk3ys7HqIfewIMkEf91HMmPu7zuW
mxAGFn72JeontDpbVr4scEU7BAMlRy+gH+qn3uYuxpaXBwspSAJhZzz0Rj1btOok
96kNYW00y8mDT8gZnaMlwqA3Rus60+BlgaOlmhQB3weZEPj+NvRHgtpqKQzCXLmh
0R3wozLlJ0psFCCnDbkOKrOe9hYP6tkcRmYIEkLKpTg4PGubuHr0H+Avq7JpfT84
lcinfVQX36YJbZqFnozz7qUGC3bXhiOeX/zqBFKlJidYggKokiCcABIBOrTDYyfF
dCi5j2G4Xg1tf4mNZJS1oEZNSknr6PJXw4hmzjGAtrqYcydxh3Co4E55t4JHGGVx
FnI1+sRxbUSJfqkHbr4WdJbdbDaRiBOmdSQQ5vsiZ5XfLCV0I2HzTaG00CEggGqe
Wd6lRFBMNwR6IhZ2XWh0u/hkALg6pXIK5ov7Ba329pyWRUNj/yj5TFry2BZ4hjef
rmTaujangjwgwIewrsC24y9yhezjhT1+BBzzZsfkJ+dy+fDsfSaZArSd80nv5+kC
UG8344FuOQkjxmHIGiDOkklj5dnDGeBkVCD9EGHJ19FJ8cnUAEXel1gZaQFzaJFB
uIGUJXElMdTex26OH+gAzAzKRIItNn19DeuDxX99EowNr8axPH83PpgDmnZtRypm
AgMgphLhwWsJU3OvKkah8jqCBu+kf+23nHYFdINugQDsrcuygAaKlOTjU3/Hul/h
bxm7fS+nO0v+s4ZG0rmtTT1bvWA7GmwcCw912MA9yab+qi7NXXIFDd8jB797nhw7
tm2bBkeekvJp9HnL8Zds1bqln2jgvXGFO4QblDxNgsWoOVujSEGw4f4dhVy6SSr1
/3xc7d/rrOVFlLR5muC2M5Yc1qrP1aWYz78T2fkuuAD+JO54vx7X0L30g3yS/r7c
XFJf9JAih+Yqg8vVmsDNDqLINCEVkkaEKvBcNdgV+9QIt7rzEl9E0G+y2vtt3kyC
`protect END_PROTECTED
