`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NdHrKXeGhyIU7ReVPWs+luHjOuceapffbtp8C3tlxaoIs/NA01gkKigw+7lj4ChA
F2airmrLh85cqAvo7jVrwOKaONqO8YYeqtSVBkNv1kAEezga/0MhEj2+1vxxKPb9
YtqQBFtvs2n9Cchw1sk8pdpN0RIuN5IxoPt9NK/VmE4lOoqfE7LX3hpixHQquXOq
T70cDoXeZN8JBgd/QcXJdCYDiTW3TcIW+tZqrp1lZ6jwD8+OxO0WW4cqntXudB7f
NGZoFO3yGaRFKsYJp4X7hhewkWKIi/0/RArt0OHEYtwoMhbkJ5DiFxTvYkqVuoqG
4y9vZsMsk0/f80TbeqKrOK0Lw3KNqfj8oytmVYZhHeDF//jUcdhKgf5SFbleCwxt
nbRNh6uRv/j+cu+dp4e4Wv6qeLeB14beNwPxqt691D8n0Tn4VAXlUrKO1PckiEfe
gqKPdVl6dPJOVL2tXDKy3L15pw2EPHZ966Sm25YN+4fwQhOZ5kw1nmnNAgv7hphx
9leD64+IyIyr5jGu0lo4Kq0F0T/Jxl4C3zwu6NcDFrvI82B6h+WnA7B39WaFNvac
SP0W+PocOAIcNdHzW3qfEXHN7xH7gsGrI3GTVoIVus+DpSGdBY9ZxSPXOTLNd0ua
TwH83dFtC7CBm5j80jiA4aKEoNvgh4UhQA+C62AosyskcVwm5tg4IKrzTcy1YsOy
B+Gs43zy8k7cdNP0qa+3DYpS4HWB527u35xLhtg/ffzWzzW26v/gqiEHotPFUlWt
gATQvY5RSXyVfpmvkUU0aoSF/FthsbjKwKONTNuU8BjIK8i5OASreVcv+b2dM1jb
p/OGH7OSXq0lJ65+tm1jg0GS9DOn82YMrp/41x0sLc0/wuwnXO42kW+8KQJsf+tP
yI7kzNmKJoEyj0e7N6m7VvTgQyBnvNmAaEUG8fipYHK7v1OvshZNueS757uey+TH
kol89TRD8KH2tBA04mf/sv+Mj/3EymXQjtPvV40ZZV7vAdeO6xqFm2vyGUxvCt1s
86DlJ0Y/MMN62Ec51uIAb0/XlEElyCCNeJy6EdtROb45rxNvwxqd945TRXwKN3Er
W0qvqOLcy7oGvT+hoW7trqwjWBIhWmocRHzG9oFOR72DsDdhehuGzy3oil1acov+
bUANyPTiSabB/AU39Bz77ZLUhAENe1i+r95lfnEt6TVlGMTlONHLRYytuJ98yiw6
5yqH8ouTNQzDaUg/VhaigwNn6GDbyOBEEdbDl6z6OOnhly8rRN3tr40X1Gmse4fw
NKn5w/prado/pKjCxmLCKzBaXUYzowSFDYy3qnanD4fFBEV5t5LrOCALO+vC68n3
05jfzhOyoykJ19dsMrzD+8G9yq+G4GbmasxZJcaOqhdQbF0N5yEqw7MNfi3Z6b66
B81U1ank9rlzbwAPK39higxsbXvR3DVpmpqLXYm2aQyhrxcNTt9GzhNnj1HpUnSw
N/JJ68lpzwPv7xBMtO2su9jyXxro+qfuzrv7SGFBfcJGjsu997oYt0Q/8d9yhH1N
/l0ro2DrfzHrBXhFGsz8IlA07Uh2FIZaVNl8rPawFOkgKs2nteKOStju/LfP0mMF
qbysPlYcbd/OQuLjRhezWULgL8S1aVd6bGIC7yTfVWkEN5LHYFtr9ld8Z48FhIOV
iFp7cEN7+lDrS0df9cdIXR6spc1Z97bYdi9z2vT+C/U7GDnWhC8a7d99a1YNG1eC
fRzLoXwpxdEv93kF2rXyuzqexuyllxlDFuAQ1EEBZ2evUZravb7NIf+KmEvk5m8L
EfAq0ufuDL+fEmz7xUfdZtMk1frGlvB0rghAHONol9XDDYKqY//9gA+qUfOMfO5e
XvzuNoKM241UEaZx+7/zpXSSjgKh8+PrRHxr/BbqdzPcO2HwNDh9qBc3IR+T6jiC
UNSwtK7vlA8blZ3gKi0Bvl3ZrjC/5HM6rkORRM78QqF8tpS3JhyG8pY6W/aVmxml
hYEaw1w10QhxnUUP+rK98FRIl+FRO6bzyBTVG2M46bKdqMD1q/FDnh3784rTH8TA
AXSs/nKdBB0fRX4drW6TVGFXAndFca2gtElthyObc6Zhn/iyqgf4z06eUffHgBOX
EK3PjkPnlMuWRVQQcJWVXSC1O4SsCsZ09wCFvrzI6iv6tOLXup6twbH66oTKSltX
7qLRXKYh8SS0UqDUhMOKHDyaVFts6fGiRyiNIj+3BGeE3X+bh82Jm3+FdUPXRFd9
TDR1C/I80+Pppzs+qmoCGNFtLNcK5MN9P9kxD0VRvVjI7qZfp/zjOUxx7G0i0/my
Bf36T4EQS2Dm3v1DKGkYt3vTm8Jq3iVy88pZGQS5bC5+InUNOXjMU1msWSBvg08S
0+xVVs8l+5Pg4OvqsbZY6gmtX/s4Nk/9Mxrj8B6tp1FDrAKT9Vt60OLHFv1GaCuA
BUAO/uidAtBP1qIEq9UN7mTS+sdJ9Iwjn+v/Q47w6XA3mvWjdQY9ycdiGxF716ck
LY+j3Qf7LtVmBjhZYcKK6iULBLJMfHR7LmeShiYtYctRyqt4DQ8monBS6ZNJkZyU
fAcWDnrD83ttqRTdTuzS9dwyuRc1YoE5Q16ouVKs1YK8q6mgCWp66e/uznR9Mxpx
2FvuHdUjZusHVAxN3+54N6v6P2BNQozGDVY8XmWKJcceRwpcVdOL70Mn7B0xSjuK
9Lw5FB+PXrnKdE+vU1WHDZMgQbbTQMAKqKt/LjFoyscaflTnZAp/b+XDQGhsa0zi
f4qBNscyk/MHZqD8GL41fSvk9YB/DSEx/i65+WaFvgGFKRAe5cN8C97iv05osIwa
8qmZCg81aTOdQoN9KNdGmdAr+hjxX7OCsU1YuwOS8Ibp8bX6WF0hz8cJcybp6y6u
7IoGEPft9LkouGJH8AfYC11ycxwZT69eNjPJOSf5Uapu6mtu4y4YDu62U/hmzBaF
YH/i5sC2yGVEkhaI2+dhM9SYaZnnCHzCajguIICgK9TqCjmWHo56kAtbNAIhIwN1
spOy1VhFtRgX0r4KE3vSaugOjZSRHbNU7001FulEpguVIm+1gYzvXEQw5dh60Dz4
9xgsI/+vnPxuT40rZhtQ1TK8H5vRle+ebiC5enkmlwKEry0tj9bHld5Jw80XxciS
Nc32r69BiS+JoD5oqMqQk2Kp5ZkeCyihv+FG8JbNksEvrgYTWJyIkx9BPTfey4li
T+jTter05wTWM9X+9tZ4UhikdPNtaybzLMFejXZe74J18K3N9mGf0yNk6BrEGjpY
aHgWspZru+NpKJHpg9oV49FtnJEO3srpITSw3OTEaWNJeWI1b1xsJtRtBQhnxkhl
Br1DmqXJ5gdN1PIqg/AfEHPDvayc8SlHKExm6ORGRDI1km02qNpJsJMkT+Br2UXn
aWka5yqGtypoXy5heMD+Z3Q0ZCd2Ap+yon2M8xiyvV38UotaDHOMTwTIpg0OhwWy
efPhwCfsjLLFWf+o1kuykGzVcYy2hylCN5FVWmKsk0t4Z9HPc78qzabPHaCp0g15
6r48Mt/3uX5iXDDsKG9HaAfbwbgXFj8M1xX5chqxDHfzYkKBgNZwaAM6fEmPx9nd
MPAXGURChOZl3ET+ubNirJ4hKtJngYH+y8k0Yp3RLvt9YcBL8ao4uDI0ZRJtc4Td
loufT8mG7oEz5ozmCcMlAP6iLX3R2XjZP3RT+2ZZC1L7GIAVu2t5LeXMpXAfdvSj
sw5rvuUc+kBOIifpMKX8g7XkMUOrpOeH1LHuS6oZnfNUj25NARWaWV1O9rkiFCTT
aQmS6BpvkaU4m3PvsUxVAPD9x9cQbaNsN3ORmt72EAXzfBck6DwzMLyFl4PHLkk/
4Eu51QA7ec57tjvD561WM/lFssEBvCOhYyqrRt5v2A8GajTDN+vvm03NMfgNlkK/
oET/ImfCBMVye4oA3VmqYWyFp1Y+SiMDXgutpGnImtJ/x7plEBOFeesRuArZmO2o
79KeVuBoaiHaPye9gW3HZahVY5BuJHVg7/s18pkqGi8BYN9dE5H5yTI18uuBDvB2
LH6s2FJMDw45i8t0VET3kGF3RK8cCHdKcGsTrbS4qWsb2cHhan6SGE7tXzprdP/m
DSzfOUPqgROz5IEM3oJHjOwkHUT+JdUBVINwO4gqi5/D0ZAMpTSkJVlGfpCD3CbT
dcOMKzPOrnIoJblltZQJ5TWM0SqlAZEuw7wBBBG/6gcKdh/5psUS50QfZL2v++tE
54RDs5i/bgrPPoX/Ezk2sgfZv+YL4PNiOMM112ld1jj9Zz2fRRaqOl4cbUK5hs1t
`protect END_PROTECTED
