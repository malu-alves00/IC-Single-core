`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xTHTBZVNans6Rb8gSE5ZF57NtkRgYEDKUxguAvkpDfijCQt5LKi8tw/dY68u5viQ
ria9uVfSgMhOU8i0sYYeVbcCRQBcm7w/S6j/or/wd5PIThM9BkMwIgdHXaymag51
zw+P/LN8+MtJhApyZDhj5gwLZVNCLJ64XLSdDF7Fc2vI4YQgmo3a3R3IMNWsZ2ba
gjNbAF95GedAJ8oR9AMMW+LwHYW6FgM0scNugAg5JvPDy2EwOEfdjGDE9u5HUcF7
c3u3H2EGB9e/aKXYPMuGZ+KCvWnzcgt3CuBh4HLuarK/UAHuuHQ07IleRU7qEAQB
JRxuM5qutISRBuE9FS1TzKYMFmCcOSYIfRFoENzwRJYkK664Ph2/P5DZGiiy591p
8q5UPLrQTTfTGT8OTDWb1OnF2Jy3L+jqIABw3X5HJP1I6OpIp9r69eg5kycnoV9E
LE+i3IDitQcg8YybYi+nK1uz6eFaM6vtbqvL+pTf4Ys9Y3fbF14aLPc6gSzOQY8a
2Jt9d/lP4mvwkpMoqbmWZeQOXdPfdDx2I+xg2EnnK/cxs/maN8jpmy10PAz9spRj
bnSR73vUeIK+1kztXCBlV7TOlBMKiEFTIssl0DnjSm/Xj6YVQKq0JJo642aLCZof
p5nlVmDyB5ciOaJZea/3q4r+Sb/30rI3kuQPtcSXikA27D8kzOzJwVwpD01UQpOI
0rlPi2kwFglmj7G0tlmhgwk5PEfSmFg0SqTCcK597jHRv07iFCwk6VYTTqxUY3vD
Sn2+pzcIKl+u+QM48n/ljZFqR60fAXKC3nRbDrOzLTqFNoxR9fWmSO344qrzPOYW
5BwOe8DNZYHMmum62x29XlBlusDNC8KLkCi6eT+cGg5Cv2y8HZ3+E60njvcJNlgG
4QppogylJLqlrR7pxbq7uOf50t2EfXtMpUvek7y0QLFIPlZWnPvdbOOjmDlcnqcW
IO16xNpNkv+zmgt3wF13xkOsl0sY9joET229lZAlJg1tH1AqBq/FM9oXeRK79FHV
atKhchy6QOWuL9WBraXhpyoftRLaRsa+8o9GKi6ifood8U+zkmiGwI/OvPHCsBnd
lqEX6moc1xOcg2zRyHsIFjbyZaybdtpU18MIMc5U53R2sW2rMfUV0rnyzmXBFqhr
d1sDx1oYCjI6OQrFmHlX9ZFwo9i5emgL+ruOF3x8EPgQ8e4AfY5n3P6B/wdLW5ya
y9ijlsy1S9cWKFpZPbtCz5ONYIETlLJ084VYxMznmwuCl1nnbDdOpjlKgkwElkDG
gWtJaibi8T82bAQW8dEKtNoxv8f6zRNRUoJjQKF20h3t0TcxYFIcpqME5krHx1sO
Sfx3yiWhK1rf2gT5mYmL4Ld3+3ZHr9GtL+fpgueI8JKKqEWqpHgxhxEUg7NWjoev
IttG5rA0S/+dbntsgbOXriAhxNaTAbEkbmA69hXHqKHrTvofhmGZoE0p8mut+vb0
9OYl/f4mwSHtZMqAqWjtdaN/U4hDMvUrYnN0FlcGWKwZuJi3ABBFgGIA0oQBnZFw
+veMg1OnEl5G4LidhmmiUQ7ut1ZSGJmVKZbnrRkiBSeksrae/wQI25ku1iJIIhDz
5T1r4RkwnqA3bsaU0++muNfrN9q21P/sTETsuZq4nRq3KiLfBaTVEi+wdTiGwvyq
8Y2kLMPdSNsM5/LSzUICDcggbDq1gtuEwibiQrM/PyzvRdtxI7hNfaTlNAexJWuG
M1GjtaSyLuaDna9vxfqf6APDYc7SnRh175Uirg8lkJGn4u7MAYGIYx/N5igdivNd
ejC8J4jTn4jbU+VqEWi273s7POsT/Zf73QgO1hr1H/ZaC4bI5AV6jlojSS1n12Qm
RHGMCH73crELE5ZdASoZ/mZoXj/878BJ1N2iIGVafoyOySrX/fk3CDz1Agc0VJJU
1yOnJl5Z1wzimV8X+R9pYEEELQIjFITqNchNtYS7m0r4/CDv43YD1lxJfZIMXZfT
tnf9icguObKsMtXA3U6EGK2Y7L7t5XFhrMaMQFBtywoKcQxHQUTQ3ltoOpBJmFrt
a37A4F9DlSgE8w/89sVMllOFDI+MNTEyQmfLOrbFuHu1raIuUJtiApvshPPBp55l
BXJk90T2GXUTaIs0CTCcltw58osSsHG7W2MW0isiRXC/TXkGKGf+BoU+yMDLOe6P
8smjf8Kc3LAbVxDHBiy24BasZRCTIzwo6ezoeIAZv1bJY/Ct/tkxoDkHdv5Xo/jR
buj65sleRwM2jXf+A5qXWah7Z1ZL0K6NyWLYneRPC8bObfkYGZV67Mf17uR8Jemw
7D3HMrhJxB1TPUhythqLyvZF56N7adezj/wd+coyOvlwkn/DAu9MhJqRg9kqCjDW
qJ0G2GrB5F+W4ALNbFqufiPcPsweRVhuhXNx5iT1sognro0GKztJEZWMwdJnPxqA
iHapge8fWcXHT3Pm2B/EH40573W/8hdVSe41pt56bfWGsOnQWjH1gbzvLhqQaijX
oC/dbWEnUmRmNrlkdM1U2q3ntCeK8+z/ErrHqt8WB/ZSf44mcf7Sy+TpINEkYsUv
9JIid7p3kMZipDuSGPvN82m/pp+EF06k7HhpaoZO4Dk7CQhSFW7FMFuG5wKyK2gP
K8D40m+UGZPIcFKZL0aGDtuKzc8ZyXr+rkbDbrZ16XwtwCE02P3ddrA4GGadwtdn
0IwB1J9G5HY9ZfVZu/kXnxlk+bIRcz0cz16s8AUaujl/o7s2+vUgxY3Lw68qeU6l
6OxrCuQ3N5shIJK8Iv13czvBEji5tPX27aA0KKqpiayVmclWHNfZERhoWQsB88dm
3HrfrYC5h2UzpD5Ba63mKm8mjRMbtrp4zhdYsII80x7zs6ZYT1M4oaOJ+uawijX9
MmbxsmJYi0HRDzmV+UVRHmdhupwalk1LSKdWHCha41CEjmJlPPL74xW67p547trT
TYOpZ11yWUC6EQgovQV7f/OSJYOjgdiY8ZQx+XrWnoWCCFQBX2BUyEM2BqgI+oTz
NkqgoV8D48EqsnTrPJIV8ILv7ufCLf8YLp66ptywdqoefO3+4ksZifrnrSG74HjI
kAQwe2Cph19reZph7eNs9itVGu5qNqhElG1nJTj1ER18vMGnp9bv0DgMdK2spDat
loGz5kKDz+5tfQ6hSFEtTSHfHY65dgAm2kRLX4xaq3xUS3+Lq14i7vXU9C46Gkpu
8BaAL7cgXgtvkEAK4e7U3b91wuQDS0Ppc0sava0HlHkQOa1KNY5W1sJbRMq7s4NO
+OUTSQ4bP0WTcsIyI2179csrVwUPkgr9dIV6QDagz7k0iCJMsivEeKKN4FWswNol
d1wWCwU4/cK05rJaKAKvmA==
`protect END_PROTECTED
