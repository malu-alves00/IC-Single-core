library verilog;
use verilog.vl_types.all;
entity main_decoder_vlg_vec_tst is
end main_decoder_vlg_vec_tst;
