`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Q7aolL1xn12W/JcRp89UV7IAbeMI3OVuCuHMMDobPEtjSIy3qywQQzAIwyw68ImQ
I/vJQPUuysf3euqn1TRcVv4BCnSxHM48iSyKSnpIGiLtTsEhhnTouetU6c9tdEeo
eqFtItFtuW1g/oDQpyPADTj4KYC+Q0tzxNDyhJeYJL0jqhXOF8pfIwnzCqV0ToKE
L0WGYgrWJBDBQNPg206gzppAANSZ9EUAbDTfp+fTgVhzDvsrJSwNmpejU6e0IPUZ
BYVkhQ22puhDVuew8RROUJCtk9j/D+U56Dj77ryn7rvN0yQaAlwOPlOQZb2/PePP
B2xPyprrJGmQN18BjpoODQOekZ87YnClqd63axO5EBnu4QrKD+vfRn57QNRiZvzN
T+M0YdA+zYJRAueLRl3HsmYgQ8COcIvPHQ8mzeOW6GCF+XmPBXWRmlnI5y9HCjuI
m0PzY6xuJUCdcjuoBYjMtJsii4l+TW4UjR3wUlHSWzde79ig4vwmvoV6WMQxSo8P
7PMKJpG0ZPhJfGDEGGAT+6kXzX6B2v/k6Azw9O8Ekl+f9NfSKuL8gAW3mTA/s3RB
nSqTKKnEcdKGW3/usO/ZPphhziQvvDQV8Xcgqcw8CWQOW9NGd8qwqE5ldX7zfFgI
ZLjwKw6rlUmPKLQIIJ+qjqJAidV3TE0PrunXOPLxUa3P9aO3mjI5fK3jPbOOjT9t
ggkW0/BvsKGSTCqSwk6ov3X5uvVQCzlkjpmasCY8KxWfVYcu1XTnEi1Qs1Z2RAQ8
Za8ohCFNb29kE3h/hkf2Q8t2CQf3L0M2qazXykblPsLBAm6sUlJSKdq80gm7SKKU
OSeqV9utk8KGlqJe7gEcuPT6QrCog7KmrHI1hjbdV9VOpWTUbbZ39OkrmG+FKWo7
j1s4/GqWpyynmglQfO2ayyQi864leFx6c87mZ39hyFm3Ju3SgzJ3XISYqND6BYdx
sqLHU4U1dsYAbX/2QHfbgAEw6qO1RyFcr1ddgzNvFAaAbMMwFFGJCMt7Xq16L1w7
g6LQTLfpr5vZ0N62U48m2qN7+bBGG/FyHo+XpgsY/BzUCCD5o09VoKi/wsTM6FH0
fBpJg61Jc3lpAER6Dbt+8A==
`protect END_PROTECTED
