`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
L6/U6tpFFnWCzgo7VOy2WdkYRFMZdF0DeJK0TTqv+yMAFU64H5XJUfu+j73PekHN
JAvJd0hauPR0Yk9QDwxHDDyL/9qWYeJLXlWbt2hoBqmYD4uZV2eynZhd/yxRbCUy
qnwzAxT83pVB3acj/p6XK8t8wJzxronJP5sy9lAIMNPuMptdoqoHVeEUV3SNO93i
FTR/f4RrPm2ot4G/rMC3KELqoUZRAP00uAYXQTaLvJEgec3JmmJKWGq/3kty3oGZ
cvFMA//jzP0SmtUNAs/ZAkVJ5hO5vqPCUvCLRehsGJlxSFu7EjzwWemTMaJ3bSXF
0Rp6eVnQ5Pi6qUAosiwblUw6flEUOtwqGeziytzky2l4zZlZchkxp/wdhLLVI4Ae
f/ja9L3t8KAbjESBKe6pZcx6Yxek63n6sVUdDLT1zSyvpNu6VRWrQcFlPvqUV99t
wK+hVPy8VXeYqDRD/eMHQE0WFL85xMIuxxO2YiGcx3rLwrc/oe7qsumEB1lkcwkk
HLSKbM6t70GNvs5fK/qi3KZ2/WMotwSZBrXGxbsaGbHxY9Dr5mScPcdG4miZnlrx
amPYkDaSfCU55wWlPphDkKNiltHelhFu3LUIml3anBCjvJ+F+jI1RGVZvvFAICbQ
nUHTNb1eCMv3I2ZydcM0fjXD8X8pBnzMm3WqLHROo66Gyc4Yx37mYZBfV+Zafhz3
lc6vTXNee3oQtV3rwiFW1VfnKMgHTfPvapsWNKogIgKoQ57PVXyoKD6y33jWtilI
ho4921tidd2XC2mz+L77VaZwEjrd9Ua1D2IQ4Q10QwsNclTGQRd6Dr1aQi9BK3EA
si5ciiEVcKbLwAbfPk6nd6TCarBch1dwU+OcQi3Su2WfxQnsqqxOxl+iQv/5nwWJ
ZxA2L2D6b2+IiFnd8pX40EhF5hbOOvc+iqENBnM6iKSlfyF/GXecDFSm9RPodZPG
BaysA89eGPT4uzDCzoIReYqDXP59MK+CcktyEovH1CX63eFUD1ol3p7ZCdFfpL4z
U2HSc3HMNymxJ2Nmk3ZVOqExEo6cfEHaZI/RB0lwVuEyPcplr/I8dVNn5EQ3KGZD
mlRFTnlJxf4F+7az5E5icRli8o5lNmpdW0ipLbdlmEgQ9zSzlqelqJtFuTdih5XN
n2Rqe6TthaTz2Ollx9sCblNL8c6Fko9RZKQGFhPm8LESPImMo+fWtx4gcS/gYG36
QjA3l/UeOzxFUwNBMztym9Yp6dmauD9eyiiw6v+2zq7/fFIH8N0AgOke/g+t8eQf
rh2MMUViS9+GcU5poxxIlnJjqk7EjhAaRILTriMxJtPYKNuAts5iElHm2qUA8eNu
7t2kFpPpF6gbCSQi6EPFew69XmdFwgZbRxlPL9QmBP01bmmEYYbZerrOtx3ya9NV
J60GMB1I9BAI4FEtg1FSWJYKJ5XcMKG0GL72oj0FSCUTukUAv2Pyw/aAmO+xeVxr
yr8AQIW7bJ941vNGoKrGVEZXqKOxxHOBE9AtSe1QzJJpAjI/Tw9jph/c/v262Q4i
puoCfexd+MivAfv3s9Jc8d0xMjUvOh70arGMW2sXfDxzAlESS34A3ZIUNLdXAptE
1OTdi9vMIn60znS07EHofHDg855ckWUY0rUdg08EEQZvYNU3X6Wk7/8+5bAaHPgX
jF0Rh1oFAaxQjrk0xKlh1uOoRBvSKThOufGHcchditz5qB8uyEOS1bJaWAZL2WV9
xhJMcjOEEOWlgPnpGUW+8oQ9t6246zJ/GfggbydsyFjtnyjN17UioiJ97KjIR8kh
tWc4Zywoc3GrTduQKOck99KiLiOPKpM2S8J+lo4cxt6fNpDMIZgJk3xk33VFW3BW
rT9BR9/3OcWMw5r8wk9m9NiPej4avhhyjqVG0h4GRkabM5rUe9jgDh4er0ciDeSg
FytR/wR3eA+6Ayn0QpfYGc8o6/1pgg9Ca9aX9ARzsxFdg5sdFygbCpvhXa59E3vW
4Gd9vjtpaP/vTZi6VbkdHauoxvkpxDhisZYKOLwLAVImFyJ4eBdtkMIWFrdWcrTK
65qYiTsoI+K5BQhnaEJriMZ2Nnm11Hy2TQx4F+tBvtInrnSdf0Io49gAxc40e7WI
LHdY7lnzzgTY1AC4++q2xeJIkp7ht0uaGT3UICO/oBbfloQ3JA+93xdbblhwr+J+
lY4Tf1DEDwRUyik97wrAeNuTBQO5PHWVUNVqV4I4YHAH4QoIBunTanyj6ZfcPoS1
4dey8dtsalV5xIKXunWTeNUun0Yd8tRSAdBopMhKswh3WeIpn+7DuvUQ6c01ZAOG
X5wNQi2MJpdPaaN4m4NK4ocIIVsbs3otwhcOw6OgEPosNot3f62Cfgpd7+fyv0et
Uq1Fy/FQ8EYaZP8Bzld/kPAG0H7Rt3+mB+l0DJpcDBG7eEtmkUbFi7nMTPTfkgxa
/kl1wHM6h/ygfRUiC121ahACzOhewbAUiqaMqsihLndtERAeRMK1/APT2Wy68p+H
1PIB7uQlSI99fYm+bPtkklXF1q+nhj3NAKghk3cdIuBQZa/vcFvadfvWNYcmFF4c
0WW+Ni97nH3M4jsPY1yBR9wgGXxJCNqI9oEaJnyY0cqYQyOSA+T65d81fO/jlwFY
5r+8s1sn6P0/r3aMdgI2YBHu0PV/h+IY8s+tX8K6mlivlb32ckGAPe7ww36akoyh
krLrFy/NlAVXlbaba7XEjfMuUMKyOHzSlcdY7lVP8GvP1IH3faM+lfgEEfJ/vxBl
NsZmpPbngVUF2lOZTkFo7rpUzgxeSfEb9qpbU9UGufR6x/KFW7nOt/fOEJlUSf0m
tLTG299xEhhKYGg6ufogPkHtQi33xdjecfZAtcSvH9zEq4woNN9gp1njiqMyCKaI
FVH91TC4L6F76beuxvI2R1Oe8k46uyVcMyvj28TfUgtyLXsEenpaNc/q+G9a1j93
lLd3G2TUJZTAF8K3e3FSqpFdm8k4HJVuynTx+R9wY5OldbCWAG2okXMYvjHmuoPJ
EX0zEeaf2wcAn3Q3jIeLNeSDgRBcibX41jS9Q0G0LCVUBLTE3ZSUu2CjNbNhmc/N
Rp/5+R4wMw5sP6+nsdmArpXVSoNy/U4YU3px9vQGxt1u+Tm57EmJuBgoPFI8UCy1
vjmaKYt2gbTcOzlEG8dBA4lsor2lX7Qpjwkh9388nfaAXopg+ePyxo54xahjUz68
rbpicyd6xcDILKVlhMdSzSzy+xpvuY2zVTgDG4UXK0Zr+lmaucAMt/5hQIcE/5nD
NsXNCvxV7ikba57shKnyEUNLS2JJRpkdRX22Z+WrUAC5MGpB2ltp8WxzKqoxja6a
amhV/ofXo80WBNIovLO2dkxlQWTJmaCc/61deQ8KfYwKeRcTksGgoyQhbTEVC0xS
b4tnNtRytUB8eB/uQ9f/SZDkOimkhbbF780BfID5I+omODqeFYmrKzZHjTCw+2TL
`protect END_PROTECTED
