`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IvLuVciqbr/zW+eKxPXPwcebjvDNo+Un+mL9sxBzm/9pckSfI2G7Jq7SKzRwUfX2
YTdCwrRjmMqasXc+eor/Gq77YZgnQvyHOHpZmjFRkE6D0CI3tr/+kZ9Y0VaFQZej
UTA6RwFcLBgevhnwwY/vW8+tsouWEEyg8qr8Ks+f+3Wi/Z2jn4HzzRLRXoZzWXyB
mjesT6E2fpxtYjhJDti1k5uR2iqe3lfc26YEavxYfUK5R+4CI+UeqWP/B3TS8H/R
6zKEpqeDfxMQMPaZOOLkHZaSIMWyI/uhCCtJvmE1IbvOBSS5UgNsS+7CmW3lwdIl
PWTkSsFUpsnYtLzslTePZIArbQ8EQWzaXVX6Qb51F15FvymqL4X8HQq1CXhmoheR
r7sGP7+7lR9rbUP1NSllBJWUA9xRa2LZL5PjuRiNlejRWK0pH367WFdDu+s8kOXS
frv+NaUA9785G9ilnWJ95xPmkIqTtcNnp1I+hLFFr+j53p2u2sqa197US2YpQDU+
E5QTX+SGhuSPUnjvflzrYo79+n43PqKQbIyg3H6A0NayIIG7JamFO1u0BdV88qlW
84CjBGfJXpDGZw07fEJmPBja8xOzNMh4HpFfPfe9GpX/0A/GUnodiyHAtRkAZnng
p9D2vAubpflQme/2RcJ824lvvU0EFA+jWlrNY4W0Are9hDfxMXOnEGFT+7IxidgY
xnWukuaq9jwJiiUUbszgR+ARsm6OoHKMuDyk95IYroRN9vy2nbtl1aYGIHCnDxFh
q+dpAZWoBXbIOwIMwTdWX8ZYJQDT/tCf995CImeFe4xCbPv+YXyOz+uVBHiYqmuK
EC14emqlAcavcOhr2DVkg2P9hmR4844ZxGxGIRoLKNsvyL2Zff+zfUmMYpD2igz2
Jxgn7WKHNP1R9m7gLErb8hzXrE18KgTpK1Xn5YGt315z0DzQG+dfF7nZeR5uHl/p
4C/I5ry3xsieFft9zoDMMr9KDXjZbtcW58g0uPVKe3YS9YKOx/k9DlGKZMdei69e
GgRHnxFSiSeUz0+C3oYmyb5hozrFWYctuOxRm5KA7SyHTC8fhdkYF8z7KLE5o3ZO
Uq8Ab4z0e5GadGly5ZWvHzKHjPd/iEiJyrwGLGrSBqlu53y1A3U7AxxZBy7h/krh
MPlC/5Tz48qgIkFF9z+GrZ+tbt0UuHw/+ZIBFDFH/lirA9XoVJvDVhjx3e05WFEv
fEDTio+EHZwbj1V0Lx0X0yID/clW1lNSMuariOgYqE8sxHerWhaxs2Tuz3mLrekA
K67g2xYSG2ZVXqe+g/FvlmRiCp8k2K/BFyM7UOc4d8F2ptBUKiweDUgRJSYppem0
lVE98vew1VkHb6mEEm79eqHMnmxENQy+t4H28yAepmvO+PjgqN5nSBPKXlfGpxr5
Ngxl8e2z7+AGVxLNzznL5bbhm3bDz07no0vBX6d9PdaA8S0xYvhBEkY9JLoc689x
qmuIbftj/zUtr4PUFUmVa1/cwQx4bFFntPYAohc5Jz75GMtNq41SXLnqYrN8QwOq
DMov4tejhjxkDAEtnMqPy0Yy8+zAzsQurT1JuOF4EYHcaZEuT00DZB5CGerZ9AgR
b383acYeWJ/CxfACXFPFCaya3ISRBxDnp0KbDjp92EXqANVA7iRs5P5CQgP69c5l
PmnQ4MYmiCS/HZik75NFuR1zW0nqQDQVNMbkvwjyGuSrywGWlIqtG08hwqveC8t3
keaTTuM7aSbhSaUBViOJDyB5lNBi1UCRqX360cnVIPi8gO1fgDw0PVec0oeEdj34
aDID33mJc5+tmfCnGBP3P2VscYd4XJi2KI5hh2v5Mhwh5ULuG6MmTdXwfadGF4ZN
xtyoPpqyWVRpyYH+76q6ZfGlF++ckSezlVJ2DskYkrLTSLDyJUY852lFfoCBdeG9
`protect END_PROTECTED
