`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6KUFftsiyFpTqVKvOC/4er8LS8eTurx63TgzhLVStM/dmYYnp0TdY3dJE3cV23Hp
VL0/P+12ffGAeBc4HZbpgfNRUeRRNMBu8YR09r/qXN3leemGcr8AvxzXF+s0OuPy
VeUSIKRz1Kh11WyuO8DNeCZOAAZODgRgmteT4RjSGnal94dZU9ycKrzJfvVKrQpc
obRgpFSBScGYRuRMBggymj5GgHH7OXBvBKj7Lqp3IlTm85eAMwn80NwduPheTlcQ
0lY0j8KqCK4Mn8zdGxF5D9pHq4Ln+bXlwlIwyLiTv6lN7+FfkDwyPxEldFhhTPzT
EEt5JTF6XOQ2ONYp3QlYiqZ3m0Ko8cE0c7lV18WLD4Umyz+mM5oUjYh4wtdrn7wD
YIobuRVamuEs/H7v1R8Pxi5sz5xENbBqujd9ekosVo8YAtQ82MHUm2/xSvKHNPwR
Ru5oCcA06pjkrN/dGkAj7llkoALX8TIjqiyBjhrnTtibeA45hSvnA532ldaoG+Qb
XxtbKVw8Rqpe9KznYbkdk4hv+KRhnMjUvWfep6qxJIZqnV7msTuGh5I61qcVOpCK
0nr2mFYVXRrKroFKSHMX+P5C5lqOKqhN6YJuyD+A1SQg1mpT0tuWX6o/Lz9cFkhJ
G/anp1DsC/98uplhCHhlukYdeDmn5FmBh/HWMY9758zNVg2WaM2p1E3uX1TIcVAK
AMlPLTo6/PP+avyrVIv4vvP6VkumyN5xHwP9/El2Id6iuhTqRtWG1dzBjPk+JNiN
ebUHoqHFTwZxS5gWgqP3ifrrCew03ekLK547VopCE4t7WgsnMkhKF/nZe7ZFIv/M
Ip6iCi0/jysw6Mv03s2uxE00/l14CyYpoKsZMPgt15RfcN7O2h7O24NldaW/e7Ln
Ayt8LgSizBXXFlf3M2zOVO43qAhA8HCzk5GlO6JdG8my6dPTaCb8dwc7inXJ/xEL
Kyrhg8TI510Tv70EsevXx95bFbYmyoQwoRW2cRyH/BrTtmzP5YdxDbBeqS2vJYZ8
PTSxHX/J+rBoVR8xWfXRHA/efBTcUKwj1vljcDHXxOOPF1oDGGstDOhTp/9JcCQD
RrBBqdCPA+n/tjl4zYwQ1cWJtGFxB+ZVu4j254IVAXw44MfKLTafhHKGenms7GYN
k1LcFjA09G7dVDXPPWnMc5+UY4OnQAsspNb8cmsT7bk0jbvy/FZf6hSz2URXoGg2
/s1DuOIorexEMGoFb9udyxBMnorPyv3v/eqigckEXUwzTQUNRAHTnrp/h/oxf79j
hsI+AAPAZRC9fOZCxlUMzGHaw2WAC1uXshBfZ4r5RJxW+KR8z+E3jsyyI4Pf6Ta/
CALVnXSpbyIZWUvRAkxK7CL4IV3llJXeMFTCT9b1/amNjEFc2v+8KbXHvxKqlh+b
RDrEX6FW3J7otgao/d3kKuAAhXkn8HIdcL+52at+cJjH75KahSJH2DEjGrThvoL1
2IpCE3xmfUj/+i1C7r+7y7aoHCtxL9wcK+GquAqQIsYlm6uC1IHEsdubcmRGWJbe
bpfko/SsEG2aGJ00s2Ny/4oz9qtBB4bnP02Njb0myYslv7JTSCHkkh227Y3KPBmr
RB5dYPSL8vjjsYn2hsELMcmWXe3umVbMcEQf8T1tt0Saww745QLM3kESl14E7oFR
5uSb7nsYvKmaQzs+MPbYvP/0ILmnxc6YIWQ4Ld4qq/CqgRUb4WTrzngoav7t1smV
7XTMZkxAifmaRrNZgM/ckw==
`protect END_PROTECTED
