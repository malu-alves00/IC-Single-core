`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1tWWaryPNDjb1gRLwJKeUSprdIFHPEFuEpKAZNWQWFaqAREDv/nVyGXmQCF67Hht
dUBxk8F4GXhpUb0HXUj79i7PWR4kaBJrPDCez31c1xTq6sTIC0WS+KfMGsOrpKbA
3CxilOTXuLlqf4RefiKHaqDbNcmrLlZ/4ZYRVtNaMnNXQlxSajCiOZmwrqVzXLoU
3qpvwhDo+j5Z94tzNRSryrn5uabqKoaDYqtAz+IZS9b9m6SQ+ERV9w6nU6S/awV3
ZW98+vVjsYlM264JpR1jw2HQhmHm2lTe26GROddnGceuoI/CU2ty1SV2jJ0p9oLb
Xtm8Yh6b+THwZwQhMuqVaEn9FN+1nzzeOIi1Iy0ifdSu32nzMzcImk48OplRkWDC
CeCFAT89mm13Me8bLR4p8at/twu4HPz3gnWjS+Uu7PLgxKRcYd8GmEnjL4sG/CTl
+XHfZ0royyMDyQsNlamdq+kEh+QaYBd7DvFMa4I8Fuj2u1uJO9+BbFLxREce6SbS
cXrFKNWTgJ9gHaulhHWvZQMf3mVXVi39qgdijES4G8kV51UaUwwD0VhggL5r4hON
3jzN31a+RVI19aAh8XCuzI0PTKhdX6eCYLTdsn08xboWcrUMmZwf3lyUScsgL2ds
/1RudMzSlYsC+T9WZsqOIPo2gNuV10SZxYyI7SJXJjnqz3y+L1gWuKf7Mbl6Abma
MjPeJe8tmsF1dZ04lrCLGIuI0fR84H8oEeCJAU6HCTqVuegmqz3xwlBRyXks4w1F
4mb8c6ixkD1lA/62Ha6psdeoJfLRXjhy+29RLb+Sy59UkGMoh5V8D+fJivpX8+n1
T0FGueFnCsjSjTC12MDepiwujpTcWID/CZxaOZSGbm28zzosWLlAcWmT3eDr5M/x
9yg04m6Gjx2ZnyFy0QhlUMCjHlX3thCiZ/BV8eDFnSqWinxgazyYhUYQ6qiQUSqJ
pfySTDFH9j75wmuTpah7xi+Kd1UPqJFmxSu+n7lYhIL4F6Vk2aoFC5sqVAQHg+2N
rMDXOeZtGDw1VWKg+7726GwN4BcL31l+yTqXo1jtfTmhhjFOkCY17AZMOJKsFL48
FMkOBaAgBBxquLTbRLZxeJgWxzOP+SxWHNLQtUBRTGo5rrgqCXRfqNidx0R5fk3n
Ud4mIcMvzkfdko+ZLdX1WAecEna3Sg08xmXbzZeHhJuosSSBGurkmsRYFScqB5RX
Niq3sFvDmsjv6LdEqjReoV8bK8gUVzXIf9r+c/fKjHrfyxPDNt3haTP8RPLg/cyO
M/fXMkoBtzDO1jvAs3WykWKlvLb1xe0hXVs2Petfue3gIl4XUUJKNdXUgbUvPEvo
QEBvtKrXr6fVFTq0Dc9y/cmLyAAzcBPhqXm+mWjgtiM8dcg79HHsmaHEYOrvkwCy
gH7cxBPcbfyUF7cvd61RA8XZZxMgP8OH85sjj1+pW0CWPXP73YOBKT1c3HyEJTso
KGF9HIk0kymJKZ0NVH2R8A336+HRPSTr0r9qaIPipNKSWZhWxQYkAKDdAhdizxJw
eiFMxTw+EVSjFeMCvZUQNzKV8pLUKhgnRj2yd/8i/JvkNfMXoFNmU+A23dNLkUhF
yf3AQSpD+Kun9ZbSmaeZimErvDwk+yu8mBcE7nuaK1s=
`protect END_PROTECTED
