`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PPEIW2MfLAfHhYTG6RZ131cDScnR//1qIWoY4MFd4ZIKJpw+XW5JmxMvU0QeupIw
nQ7GlocI2hbWaoHYrR53k5CuX8UaBK8aOIVjmdJSxqmqqJ4RwUGvUpaJD1sI7bKQ
QfnrUqvDzp6dhj4k6meTt6Yhc0B0fwL0kXxgZ3w8eraWq5a3k2ZG5KRhmFcE3EyA
I/pRwI7+w+Gp1/h1SNfGLTq1u7WzCRAh2eGX63Myf6bTKZy/1Bbvw56lnOMX8m+J
r17yY74nluUfeixiIsdvu/ldrP3MjbQ4Wg4wyWdGMj0QUbtrKsCW2mtdUVcZPjAv
0F+SUiLiYeh91X6YmYlHV67EhPW4E3ItBIV8kC6TMmRexD89Y02cuDebcGlnZVrP
skFebhs/KMau2PwXiXjnLTG+yjyo+bTMDQDqa5n4qWeA1eenDXzIlpP7UpXUKuTF
ylLEoaDUzHUz2A3Liqbbq/ZMQ4F69zzPs5aZA5Okyan2pe9LzTYHqeCNu/fqsbKt
5eW4hqX41YSEJwQFtLzdSdrsMJlVmVOWsWBN9Yc5OQGvvZrijex3MGjrJ7RCZ/b6
iG2KsADuDgwCD3ZBPZkuAyBpQWBfK+xL+IRhXeHqMFMjZ2WZelRfSJXEgID0sMXm
C/u5fV6PUMKwO0AJesLmnk/IAXHMJvbTKDChOvAai1LV2x7ZUh0+aPzRPPo6htkq
u2PdSAMALCxPwUhB2AUML3xfVGGJrShk/kd7l4xvtxL9/8EhbjLiXq8onPV/GnTe
mtt2Ij4OgqkCaZPkGGQITFsBPzQyt+t9Sq0s8TPcNpiQwkBF8Ub3hexEYlxTrDup
OJR6pFNonHBoCLEp5KUuuno+N/wuNtBaVcQGKisTRj9xnDLHWJintr4JAEdMDYAz
LPblc87RLt4tqf2howlkhsz9c6f98+FL4m0TN5uc2IBNrYV2mG1rtO4Ir75amQ46
f7wC6d/cTOzF8s4TolWqA9LEtJmjhzvdZ5AE+tyeHoh5mqYVSy8AxhZrJBxWqW/M
dyAjNikf46sYFfLAclje/IkC28rDLHHHtftwB077dj97iT1jhSgwN9sCBVHrmmwc
6YlMJfv/hgNdxz1hkbPMnM8Q2VLPmz7IAmLRYVFFsQIho6cxsFF6as1EaatlhLE7
Mlc6ixQ0jVintS1E5xwJb3Y/gHGrwj0e8Ai5M8/KC1jY3zKRyd0Ae3PHqeOgypsq
3U7ehGEqqMdt/XDgdxbt02sBhZVmfruC1XHNugSHDwQYKgOaDA190tXHAzfB5oPZ
Y0PzhdJBGOVNdH/0RYRKrj9ZE5DTLTZJvH9yEqdOgeEHeW/qRGd/zEv8doyn3DeG
kKcBg6TWUWdE00PaCF1b6o4Ha3ctK5ryDQgZHD7cPd4PnmZlY5d2dIjm4U9hBl5w
gWj4ojJzhd0MBJ7AQFEs5na/s0t12x+ZQMmPgz+PQ97h1k+WDBq4HPuMi7bTmkLh
vM5/r5Z2Kgb1aB5C27GNG34OHan3KUyGzFOpXYJFOi1lekIc2J8J93AmZqJqJGlD
C7bhI1RGVGMmDvkqM2pJK6uALo7hvwhvc8UkdYku5djL4IukDmxNbynKO7Hy3brr
i1uXqORuINqxBbHBscFttw==
`protect END_PROTECTED
