`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wDihOJy/t7aCYoai2Mi+gM0qMWotUkablwqwAubKQOAqXRpALEsBbN8qMvWD8CNq
KQH9FAxQiSsTP5R0RGcSfNTEErBo5jezynnyv2n6z9HL2O3TyEat3dnopaZ2kOjZ
A8szLlTx3OC6c6b/3Fww0L6v1z33yuSJJneejmL47/5mIvjvwxqyQKc3OElYaQ2z
7GSjNMLtqvfkGNflNNwqlVeT4rA8QzJESOhwjHJIgnsxochIwNydvFwymQ1eBzVK
Ope+IiRRfO4GpgdW7UdyqtJj7VJahjRGXv+GkqM9op4+3Mmbu1t8IQpN9BINM7dw
FiLkXcABJ3tRjvpmqQZKhEGoBvWzEjQiatd8j3AIwjdRyeBhnZmLj9su6D6RD4Lx
HdV0oDUh5WT6EZpaHyy9ATUduOQlpp7cTCIgloQ13sO6Nqt7iyBTq8kuvvXCzjBS
9X3Akg8zeOvBHvC9xkOHvPTzthejnRJZocbzTNUMuZ3xXqiPn1ZyqIMmb7KHfbgt
CUyBIZatLw+7jE6X4MjqXTOlmvIdcHoXqCLypBvUmaIx6PBiY0ZxJfbvpabCmEiG
QoYVNA+VZni8FWH9kZ07WVO/cki7cC+lRHqdc4gf7gLIBJ6iKc087sjkcUQrK7FO
6MJTe4nDoT1K4sYhlMsVZFv0MnsbVC4kMODOHjnL9pCvTQ6nf2PLJq0KiE2N8Anw
XIpIFqTKQ4ANboI0eAhX+2Khppx+NDWl/tdMZt0iekOTqYZdz592O5iwCHBlXusj
xiw9jTETF3A99XUBPxjLcR+Y+sfP9SoizmckhwnowCE8cHhi12vGgOpOJVM2f5Uz
5VKUgwNm2SrKDkKe/hlIwvR9D2a6OcdHP3mdJ6slelZYvCSg1BdVGNN9X0jMIq0W
eoknsfjf8LdcI9/E2AfSQK8IOzp+A4XUh9OcjQqaMMDkTl8MrIsfr3QtbPH6UkwV
cyo0SK1lIB8ibMnfqOen0xFCEtZFci84xQhWlsnJEY0EpbZY6s5McIh8uL8rPraj
m89GsjoZ8K9XVn0BNfZ68cd2ietzVPhndDGa/ZjC7kipVSzWhgo7eE6UukZxOqOq
paYquVTR0NYE5XJsb84vO5aW/E8UbWJ22xFxdPSyEK6ldVUcUUcEoYKqgs8H/eoL
QIUxsR8clvuGRlApHwcB0fJCPlOj3By5t5BlSUSsGeQsfhvw5C2t9VRCOoGF1q58
HwHg7YYJiDww/bGrn4WOQW20qIJomCUStSHGoWSAyBfeTA/xMjPLpEZWMrOYl0lB
4faInZlDoZLSZTaJIaA8GY0C7tntqz/UpXtb9U9y09Aypnkxpk5ccs7WHgYIAMmY
J91ELpBtIuk1WjR8+tHfZ7TLMwlDwS1JTTKDWk9CX6OFPsjeZ9eWrlvB1DhvHVFN
W83JEkUHtvEm9+Xt6WL93+S7ndFDa9g2MXzkFTNZFeRLlgMf7egxO/Q6pqvOwBxW
e8AxDR8660um53xDojqSj/qae+EGWtg7L7IXaZMtrQ7SMxVNK4giZ0zCLyGy9bEo
JxA24Un9losujHAx19mw6PrPpk58P8NgZFq2wXMLroWRd8NSGKb2B9hvUTjq8L8U
X48s+fYczB7JJ7wRCqXTmIw2QeMbFyQBemN6yVCbs4a2ktQMb45iVdGYjqTB/V1t
BimysoT6cNyhp2Z5Eo0Gz6L6c/GeH9IRwJzV+NY9ISeu3Og2/3zUhYhYJ4KuH/vA
qLeWXXVzwsrPNhEqT2YypOHE2m/HmQThE1virxAsB9uYcALvJaqNrjp7PVK0e2E4
rTtdZGREmrcAeQ1jFYoiOp6uA1JA85Rv8t/K5+XY4bH1MhuPDmBtTkdQwwP29YLM
IqlWGVP/k4p5C96T88h3B3JLdO7VhlUJ8Ctc7N4LgWdl2GxUHL8cKVDbujHAXlx6
PuxtDzjN8ea+NrN5Pz8onrCRIG+zwYMwb3bGwpZFLHJw1OGquuhCOhFEQbqsdrjM
NwAybZ6OQ3hcjckbY24oejpF2ZIIJruCkZPiliWaSlDvR06i2a1py5FAHwrCKVDD
R1mYKLNfWV2MJ/Dm88jcQDSX8fnYM9TsxllT2cvbWqxSKyD5RDyD/yN4plcX9zbJ
IbWF7Ovk+qjhkvTtG/NjBW9SW8q9q5QjxsRmSxuH5UOKmKCf6clyKh5klYTgQeEx
HPvpYX2xQt3Y1KRud0m1eiw8/br5IPhAlepIjEbZGME7hcQYWrUDGxDVUwxbhBGP
c7EQ2UxTYtiSLWhjFEhvJLai2qOJjhvoaB1sg5aWr6JPAnTGqJX7eScNQecUHLFO
rgR7stk5MaRpeV5yadK7ZGSdLlUyBUAGlvIM2ocb2ikeEbghU8k1I9vXVhFCfXNu
X5w7C3e+BPBEyHdWgXPVQ8Y/iplRSueM0c6bLdXiwe9ovICKJq1rq/kZZ+4AVUZ7
Qkx955LMDtlmxmhsy8ZCn04k+t2HyouiC88Ht721jADISTv9wB1L+9WCGmMXos+9
hWkClqrDiEKBTBzLY3UaZiwJORUon7+FkIDP92EyzBtc61/tRu7QW8PnotVPykSM
qubFRTsXJPYmHI0dTjeEIZNPj+imEtMlzwBs3upJDwHzs2FCwigbb2kskXYkU7pB
rLDtI+tsDDZpYhRBKeHBcOZ4sanMXPdVU72/9vtQso8UF03derRTCuXUdXfQHcVl
9imwPyuFe6vHIus0guLnLQ/gem6prxgqXWntIiDQYPBQ6URkc9QCArTHLcUj4oof
mDP5JMKjr1XnMoos/27ZRG86b+ZZ0qxVnyfG+tdawiaX/Tp2uO3V512fKZnzjYnu
XlGoU06t4LQidJzm6eYqAkWpGzxjKmAcS8Mxyjs0pUEmeD2FgrR6XkJvqYITGK44
ofPHHYr4k1cpDqbPkQr3q9zUDaW+pKJG8W4Rv+nQizwAgPqDglJ11ROhDqdH/Tat
isLhrea4LvHldqX7t8imy6rlRyRBFSZN7uVSH6rHzw0o/xTk+ZpT5N5tBNk8cETC
qbAezHc0zIb24AUioHc33pAg6SKiznxjKDjXLIM6kj8PnGmGptMNKAIJGhrJOHoY
2DKw1ZGxp9REW1R34I7nZ8yEcr5PR1+twN4+O2LiXgqeff1cQVymlTDiXqxKojB9
KkKYGBg3Sge8FLgVsP10r46rvlijZP3UfkxVfAuew3yOnGjEwP11JBVX9kXlSpA0
6t6Rt0pBR3OQ2k2WUVZ1/6sI3/3EOIrfstgb1pY7t9J2O2H4UI4CHQuZq74Rl+6l
Dwcnn3PcApR+st+ib6pVbd2ThKY0uLJa6zZpIG82g0F+zl5lF+OjxSlc1YK0UYst
e1rgCSHbhPSjIsFcLGoM3DoUybB9GXhdTuSlzpTi6oJHmB1uRw4/gpq3uIcwHZrO
QqmydHw+kxV1BIDOzQp8VwMpDSBrApLwsbcG/MeGfmTqceYhMGmxdldSSwFXccZC
i9wQSpdd1LBXf0IX5yOZc2LdJl6J9eAyxijo0Lxsavl65kjrDjHQrZsWdgvYR/eC
/5o3bJfzaw17H75QAX++9KDIyNPLtVs3N/FXc3zU6JS7DXp/1NGE38xl/t/iZurP
XfOfI7sRg6IR0kGJNOZK3jy+nPPRW9AYoBnOBVSLDvuduqeNCwsljYXaCaB7IA4j
ByAxXxvg0qmZYM3bR+1vrQ2u6o3cWoQHQc+qXAIvHQlpheH2uP3Ge9cbciu0UHXD
F9rLsViHBl2RCf6P8QVa4vgPGPC61KgISk0PB7Pb2B0dIECJB6xM33S+473/EeBm
uC0U/ERoFr1OvPm9f6JxBIS0K7y2yfzOwmyt2suZz7KyV8z24T17M3Kyw937nYV0
/kbx6xtIAfurKuw3bbu1l4xnt3R/P8auXtrqhu15u++2L5cei7+0N2nn27Z2VQqA
R5aUpcY6MmxqA4UbV876eULbLAylNGZYi1dTjvWDyqvWTX7Jmm9ZUOGBLzRLTQl6
sUrEU0O197uNJbmWX/NuXNU5SaGpa+Gez75znDxwziZObh4FkEwb6kgdwdXeU1MM
j9nDBV/v+sYZlXdl2qfwnAsar2RfoSDdYWIbRqpnhP4LVvQZzf6GZtqfgREUuG3a
ly9KPbcnycRkMK1+GAUtGm2pVhUWn0BYywmiRGGf/u9FruS1b7IcDOEwyZYVNi8C
qYV5llRgewHov8bvrEHrUkPhgdqkIBwCDdgt1eaaq+DqaiPGpO7ZcoNG0CoHB6nm
tNFlWXSsszF5QkwNaPLFwqKaQjDz3qYjTL+Img3af6Te4tLlty6Ux9RRWda/rCjr
AupiCcCGojyNpF9RO0NdFOuN1DdCzHEdFlhqpo3ei/iJzJGX9CHiA5Wg4zcEvWP8
Ig5L3gHNf6JPQxVNg8RyezRYqqmivP7dDkLs7Mcy1zc8H/V3fiinsEmaaX03xLdI
uE+AoLJKO7hWThbkeiLdgQ9fYDUrz+IDyyBu3PAPs1s49iQj2XCVOARlxWnjrHAI
iwvmwS582FnnFAAaf91P3OY0l9GV66ArYcvnWVfy5W1c07g47o2lsFoHuyVvx+xF
0/fnfl32qPMu3dDG4IGbZhKLJ3Lnfz6JYeNswowm/jVbm3+RdW3YLt59C3FL10+k
4AKG2x1zAlpGDUOI4Bsm69jT+hrslXYSRCLb5eaaka/goOl0/U5HPdc2PWjqMrNQ
WLrtRn/7YMh0lUMCb/YkXaysYufKp4adxFPlcLiEwsn5vPRszeoZgZsB4J6Zlvo1
ousVo7+kaWw/p+vbTkmfUrXagJvmZY8nTyzdcyUebWmlnJePclu9n6tFo/HPvgzS
o+WLTgDuCyqwJEznfzGhWGK+hcrSVvprOwagq5eXpnwUWfrufpXWhtDOFnHO8FR/
71YZLmLUToVduVV++3mAs6zRzlQWiSGacyCiVfKwFkZoCAshkdicUzAl6g5KriGX
2mt17MkngUuFVgEI8OrZmwtlMpXajZUtNQ0hIX3Vl/4lVJCrx65pHJaS5cvSLPgW
WmkUGUbKeyPVesnVTZvGy4jMaMC5d8UP7sebcHsLNfUHZXZrXTh7UpboRhNsZX5O
p1qpWEjdyOICDmtEa5yx7GrGulSU8DGTGtVet554niUd6rOuTUNni/GMhvXCwY9y
VYFJ24MuQfETem7x8Tvml1Ovs0Yy2BgPU/dthJwuN0wAcKKVAn8NjN/QG/1TVT+1
sSqBGveaAwHew4JMsuN+jOwFjRUjcGIzubxRr0YU41at6uMHvxgSWFVHtW5Vf+9B
XHfkntsHqLbPA1EoBtPF+9MMIi6ZJBP+KxURrekm/fW4BCkV5bK6i48ilrHsyPOO
nmR0lZqyYIhfE3cQr2lSqjYi1D5Glz+Cs0QzaZyHBK5UkWRx92gRDdUE0BWkZasK
gHIzKCYxodyuLQqWfgY+x/FNLygbenbFZ6cwu4WddQfl8ymOK1CwiwjX8bjh1t8c
wgyXTfw5jcGfM/K8rNHU1xE2KV4vW9ZyV7n14RSLxvREc1S1ca3+KLJ87F8LfDuw
fCiCnlOtIU01qhgCVnbIxnAdUHPVOUcP/OwUYbO5dUS9VRp6/hkIEIZLoHVHXdgR
JwfVwLTdLzHlfg2DUjq65Pcl/61WinEBW6JXHQ9lZ9f0OBys5EFvGoOPU86Wvdf4
kgKt6xHby78ycSLOmjENrRb2aa3zUgMGaC9/8x04e+aDTN08qxxx7YGAhObnygXu
5uQLEPkO4/EVtX+EUh6YzsI+9X3UlLQK7XibuAATAFfsUVsTWB/P43bux884CLk2
RChRKu4naIYcTyQR4cc15mE7bCken505Bqk7yrIfi/YpX7K9gIULoi1QmbgXx5Sf
YiVXkc9KiZIgsflMatGMKmhg6LFKWI+FtqdQ5ITgy2+1fKbDsj6ZvI2Hnz+HuHgt
G9ibdREmczhr5RIkXQZ4InrvfANqlyoShJSUvHY6OOG25iAAEdkuT6iFq1HT3MwL
4vYt88wjXSz6HTllYU954ZVNI2KKE2VEyMQ24wtCaK8EgDPo1y67gdvsSJqc88eO
TDjGNXY6DHB9l8ZarDIQgGTXO8wTac92eRM0xHWNjBQenzHhvftcekSXQcNR7X+L
OAe4cmA2rp3VQ6LfGAVQVPsh5BnW74+KuBDLjaAFUsPo6q93ynt6tc+hitu8sAYg
2WfgV3oLB2uDHUn2+DlT8VCytQ6WktHsRwLZSfbz18FpgbMxTRgD9zlywp2rpluF
aohXOgC/Ma6ayAxnNX2KOKRGRi4UiK4Ye1zervLMZFQjmBVQPuPdKe0RsOfHis/k
aim1iAv4NmdrS1tIoIOQFNWiG3BPLLLVU4sPUlzZoN4kA1CuaHCqOg2JfwhWSfwi
2sF/aBC+6ktbKyYdecWTQ6U6DB2p5wm3JKBsHPpLOMjftfs6jBBMV9DiPEQl4AWe
zuvxfYI4SvBjv2M1xQGRMtyE1ZiEoH8ryOZJfTL81rJN9mU1mmr/qcRjuaM3P5ZG
dhDhN/NNZ16c+Gvclkk7CdDdEBL5/FTAbR7zR3OzFXgtjd2iSOp1ddxgwTLqETJO
szhseeerdYjJmoOIi6H/prWioOGy4biE+vQyB8JtV+e1jz5y9dMdiOTdhT9LQtJs
DOMg9wUSdKaMoDuFjwg9CvXyl7wcLpNO65umEqckC0T47Ue/DWz8lhxgRpysZ9F4
h0s9v5p01LiwLWrMyAtC14dmn6VBhzvSmRoXRYr4Iyc8xmWGtPB8lToJDb2vLhAD
IkuRYkLjEuaNH018iHgE9I19cdS3rQQffNZJBmgKmMDH53+jmknviFAo26fwtZoL
6J5IUmAlG6hbb/kvCmGNOtgDFypUYEzG6rIhnDsQmJwavi/KKnjttkCJobEb3v1L
SY6fdX7CqmQbN9bKkTFYvjE9+g8zmgWB5sT5gNu+BtDzJAZgw2QM9UL9/BGA7B02
TKiqUPFA2LZwMHMz+I8/SvMyPRmdWvrzCE5DMZWl23jONu1HELIobEEJL/pXcDiM
DDGVWup9u7FnAS/ntP5Th/B05zXcQ6/yLDQXE9sYNzLtQvnZfZBm+mhE266GuaPO
90qk5Gs3n2KV0dxg8mJPpboUrEeWMhGPSFXGRKUGx+kyjx+n2mxdIA4G/QaNVs+Z
CuR74kQFx1kOD4chIK47GVHhZ+zxMOIAaae6qCdTEmC+5BD+gdWWDYQ2pcjf3nf5
i8zSsrhKKO4A8KfmSZwpdUL/WBzRTidXir9aJSen43pZraLCJFQ2DvA4nmd4QmWc
FO9sDoVtKnGaKk76aoHTXVRToQOd7hCSd0l1FnpebWu8Frz+gDU9PuHB4cGjEqlO
hd/WDs/A07bgeh3SbCRGEJ31Ihsg3br6M8jwhTwve90BM999kjYMkJQyZjyBPIpo
tY9HllU/7GbHd0dzwB9rwPb2mzKcnb7XWXvkw25xL9b9klay7hhB5zNCJU96urAj
1LQybSbBDYsZtOQgvz3dCkvjwGTzzQh+4xsYM0EiLlMapSFSXB89Ebmh6Xz9oxJt
CsKIz+MB2pJZrd0Uw+txgIEY00oCuy1weNt2DbyM7UR3zE7w0rlXxmoiEZs+UDwj
JEYQIBnZoT8w5iFZJj+azakZqhxKTh97o/e61dUj4QDwgM8DPOUmRfWhkwKbt1xK
scb09BZwH8SkvZEeEe0S6S7INGELlra9WKg+wZT8pt8u5l6slmkvLtoZhrs6tvqT
UnNXn0RDcHHxNkQxzQ9CH23tp+pztFXyN0Am6RuHpv+PCA8AWNBT3W3YSiONwAtG
SvHTNMuo7c9IWx/PjSSka0ANIxdXB9axOgrpBIdrsKToGw2osDa9yfGDxrxu4YkC
0Xg0+kBTCCCZ9WB3HNFVKF09dZcbEhXFqUU+MMZ/8vnoDz71MxM87yTDikMkZknI
SaPleZRX9u+DlEEnT6U2yABxuMrIQ78DbUWlpbUqgeeshISExZdvlEPFagT60jxz
YwL72rBLCaFQabyljv/QI0EwJQQfNd32ufhRIgvenJHl/L4qeJOfsTKtQR5vkoQ7
HE2H3iLhytRhONH/dgIFvJc7lHB59qjmnPzLmLejtQkSfxPY8lHv3hwKFEwStLOk
MQ8LW8OQUpNccWFq/CZQMGhc7jY3RAMcYiLblhu5HDV99goSkBTinAEdEbBagO/E
1DU4m+86QEOv/+0JtzpoXpzOYrZlEtfYv0tBXbQbrg4CMouTNT4GkqTan1PuwLsv
+i2TQHW3AYfLdWgJ80kS2y0bellDsK89YB4u6yNmulUfWO9kLbLe3sCXWlSTnCr/
svhrFF10PjdMe//dCPSEq/X75M7/luJCjGvzNAZRhpU4JZE8GGP6M5cQ6VCGsntB
31FjHRXVeJrLicJD9GVQKn6IUUzyfbetWfAM6UEV2QVsdn3bLuxYqHdGSmmxKFm2
ixFPw5pgoxnPd9EGgK5QLiAfxVDzjXtrRqpiBewwY6VCStzSdvULOw1vsQNfqjp5
qdOAa8LEMpaT4dIVFI07dNZkA5mVQSyEYOMfx0D7kXl6uJoBEKplwzMwb1ZjkJzG
9rUq2NgKJrSUEaf3afgzimWwazNv2lBSJPEgV7mjdcalhG17s+2Ipe0I2E4fO4Xq
GlfkdBiQR4U+byP45cgdNgSoRANWczB27EYoF47FNFesQ6k2GQ/FNXkec+HbUorQ
9x4lrd39S9dAy2w0f7zQdpwrDASv4FDUA8tclCWYMMOro4lxBEQd4lNMbvZhY1we
q6AyMUftpRImpjDQ2UxQQsQMNzoAJF7o+pTdgxt2MqosqwNTAt9lo9V/HA82+ouO
tRPuzD2hEVpMZWeZ2iGswLK3DAy8IZKgh7IXziM85CNBN9KOUaEPQFlsm87/9Nqh
j0cjiGAoJUhsymjMmJJZesfL8/nzAGwBaItlin09Ww/n1gXmT6kyphGLNTMFavBi
Mg0WZz5qDmlYa1Bfesl4XfWV1I1spn5AEsLFj1Vf79Z81inDWoW6hlyvFVXry0DS
C2O2ntzSGJb/HgTBraD+vf5ntCOdjnmL/9A9W4QO4fsf8IbsTseIq5v5jbmcDYiR
GCl8tkfzIXJLVRTttC2nqzlDdZdA8p7itHS9gJPHNRic3RPzFnfmA08wdJ2RErHy
43MHqqLTeLpElCHs/x0zR5NV3lOa9/3GZ+MjkqD1sM/IA4MXRz1+P9kdAVciQQ1C
RRefMt5XtJqifSxPg99y+gbs2Ty+gWBimuc2ypwcPDrs0CE3nlOR4lWTyEHQSKiK
sDGW9q7FX9rd7WImOe3AqzTa4Mv40hVGfhz68NsjP18wMvoSCWeTG8UfozsvVVPI
2VUCZ5VTDMgB/voOdaIywa0vWRWhjJCl9NH4g7h8aBdk/y64iP9oz8dHUEceHzzr
5aQeC41kNVJEn4tAGcBBpxg72Bdc26E3wfR01V6fOEMqzPrM1xGbGeSn9XbdidA8
C59gZgOTtWpfXTl4UMSqPjF4lxqGXoAv0uK9LcpCa2ZdteNBXMpPuRrZRDDq9gcH
tWlvhTFcdKDHmoYqhv9jh1VOoE8dYvPXGbCSNxD5lT2jDs4Ls/Fn4hcVREG08TO2
cVcOos3JOZbu/nWRCNdvueGp9QQAAC+AWyowfITcIbFx89KN/nB7ZM8C1blZ5Zaz
SprRYwHbwXoRcetYrLmyWH1syoKwua3/OemcWqqzmQlIkc5TqQBiRirWavonIWqS
blE+4tMmcGoQBQeXGTYY0kzv2k8EsuOQ7LDk2PxbXk1WZDhEHsBP5Dec1sPrD9gx
UMRULnKbFR6Ycvp8h7sXhzVC9axIXTN39VtTtvjUdTTDxRzPetvjXtaDVD/9ZGT3
dZAUiYAb4qYsNAWTzm+Naqu3XHnb4jSpt4+h6dbUfcdRQ4ipKcPObUPjfbvelNU9
JkcUYLw12vVzW1pSKcGWWoVyQytFrjkNB9ykxn/9igOWqXbon1y8VQudYKAOnMMK
mJLtfOcB9nb8SdImx3Dm0heN4R/TEgBDD7PwBvMmFiL04ce5lpKZEbn7A+0PB1JZ
ePhpdAKj2GZRxOJ/BX+K6oGCCsvi7yFM2RDtdoRDJ3WEHNJ0B0yITMMVnhf8r8MD
pMxdipczRkO8MbUKD8wJN5MtxvikduggVub422JLQoF16XlkarWCKfxNejFAot7U
b568x1TPmOXdBjV8jCM6ERmoCcvkugDlN3MPVAJ03Pf1QAVaM+gQlm1gY5+3xYBY
94oGFdwWWua1cos7UzsPzpT7vsAzQB0DheLXdJ9UuV6dfWIC3WbWPJh6rgRDRn7N
6X7L5QAl/RoF6ETQ0SdGs4Ukpkzv6sd7qh6X2pXQiNn8o6CUDI+5RQ6IMQwNHqcK
C/OpIBslWYJfN6RsAaAWiYHwW0IxRyG55Aeztv6ktcmkRMnsO96whl6gYwNGPrjy
zLpHF0C1FpTgwVQpcAjDLIJVvRRbE0WTcvimfYr3IL+XTibrWyjzmu5sLMex+wzi
AFcDMgikPtjpdHI7+ZxaEJVLwUlqirmkU75aMlr7tTiJHaczFhHVSm6o0AoTu1iD
4463C92rXUBjoe1UWg22Ldv3qcc7x9qnvIZdmeZAtKWcnfjE8oUIazhxdcpJRve5
44BuZ522S2YFmJ6DATnctAJ7kzo0jFMz1xccRyhxzP4wRGz+uPVxi/dCRfP/xtOO
1UAsmPsZ+D4gaUTDfO0bHFfNpwNepU0W9lyJ1PjM74+DH3gnhpW2OfmVL08yHQFf
a+CuvPsibCaJIhK3y+ia/0q5I7XNjh8Hat0BPAz2QlMYd/6Kbg2uZSLN6gbwtJDM
ouo87M2XsIVC/PO4rnAO9hWVuiKZ4b2vLIOSA0L5NDrbZjayPySNDXbkDwfoEZxu
bXgtoQ+vfSvrcJw9T4qazZ3/ehFIls6zu3vRQ+3dSn7U3Ugj4XA6sAsRkl1ouZRu
Yov5or6UVQUxSVsiJMv6+Q2yZvacwzrXtB+d+cURpHD29DpX4IxQ0gk1OP/B5qwR
wgxo1ieALvSbLlx9xCbAOcop7+/rOhrpH3k9aiEuRSpY3MaKHxC8bhqn+YjwM8Ft
aYmO7lfcS+sUTL740DYi1D9s4iCXMGeAnK0D/fOknozK00QQ+J64O/nRHA/+Jf9z
8L41gXOhNSX3wKazRwHNvb49r6QHLVme85reprEC2FUdWllpaNHsF812IVtcrEwn
JZOhI9AaJXsOA69EfiDnZxnZXTa/qx7nMCLecrNZRfbe4TTRsY9+EJrfEEgMcgO5
xkykEeOksjwuXTrMJLG2hxH1ZTs/Nih7LC2N383Amrvk6j5toXJZlZGazvCLIT3J
eDPTYHUnPSvv0VpRCcMDhW1hRXytUK1tBvhyrvN9PToahZFxa8jIqS8L4aqOofYj
oiYyckpV0NlgGCWEBNy0DuebkJBWK2lLuF+yt2LNSgLsMrQdhJNRGOrqryfu0O6F
MRGZ/mL/HIhQ8eVvnFQccd7d7K0oLnnUwPX/XXj4kROz7E4fsP/yJHCLVJ5CWqSL
Zql8Da3fMXmRt8naf8DsiFwS+y1KqG8WRqvmJk3TbhvMcGXXFhGCn0uyRIuZaCzZ
VMi/X2MKZ/oKZuzTZlULRwzbUMeogNhMHy76F7U2m69VGYDzlXvSapVJ/ddV2mcs
b2OWQQELnddinn3X0wFPcAfhJWDB3WcARR7biS0yJgt5XePJ5n7l+WCKYob7mRUB
mqidn0/Clb0XaNcZQhUg5RLZYPUSmgGMRp5byKoMKFXRlXUiQ6CH6GbL4dgFeHUV
VwX/n+25mfbMr2oBaHHhybOjmZn2ZrazExdW5s7YvilBjvsdqCFPNF2hvkF1nREp
qZxjyUZ9A5SNrmc/X/z/zBR64wsbY70xiXRURQa03tybcP+Fd6Z68TlZ6SOOZuba
PGluhRsRWbYUnQ9oTrgAYn4RQz089XnGfipHJAZq3rcd77iSUvUuqm7pP8Ad76Vt
4ZoGCGtslxbhEIPosJ81Mw9ymvxRfUlZgyn5Eb2qZ7cY4F1PNYR7uelmF5E0J/kA
UEm8vDQkxOEmMtDMOJROyvFyvJutsIYXbd0Ha1PST0gE5C8W0LQzz1Xu+YNS/unP
7rIuamNu8I4JDD/HyF0Y42XhKBExuZfPHpFQtvcuXyOGYcggD+NGNxuguyfd34Kh
dnAbezjaNjCrsb5/aQM/STK8vggIpcfKQ9yc850csxA+cLgL8Dn3F281deSTfown
EzZj//+PCeAV+9a7SBVhSDjzsEycSngVY1coXwhI0qwV1O/594NR7KEf+H5yFAfp
XS2C6q/FMxYXbe2GNz53DsHXEaHtUMJPL5tnGfk8z0NuhequAErPBA8dBgVK7Rry
36CokK3pBfqG53y52vFSTezMqlnIpVplpHND1c6/AyxPL8GDfvoBBsdlsPzfqKDT
qlCIzEoNwfuhr0zge5+4uM9j7UzbNQqKnf6jMdsLJHctbULCP+PwtnctmbfmuTRR
CBsRBV1yr7EcNmF2CEfyleFYrpsytzMJWHYwTKKy6NzeBq37LNCvfESTjqn89nvd
yqB3FVPkNasuOBHRTof6oV8KH17q2MSWKx/YKZzs/+90Daxif0YRtQQZ8tN40cfP
JQvzMCaOcyRPScjxOlXdwyRw1ASTxq7fmf6K2o4iVYteV9hwjBP3ZJAkrUEH00aA
OhEqDsJimp6VDS51eQlfKdw0RkJiKpPZNKJOIzi7c6C79d0I5WOYgTT+FOC9jTba
W2AAag1cQ8VVBtLDYbZq6++P6H94Jd4U/SUZ3pSlBO+PexwwBeb18+0w9g2k5x+G
cyIehhu/4y0jzxElmJ6i3MtyFw3agfxQxnh5k+vF390z+jLtlObWAH4UX37fRlYp
kU0BEc+3X3KoXDb69RqSk9Pozv2Htkb0I5c4mx+fzaFph58b6cNzWxXW5XPjf2yC
iyrdPEiTeopAzuBc2fFktaflcQHZbESCuAtmrDrluAouyKQZdeQ0sT+pPGSIyjNE
e6+VvZB3GZHw3KlWloD7viVYsRVUKjdG3ghUlt5g2SVUJ0rT4SUlSEcyoqkYPnvX
CsKhfNTJnrXPH4qo8DkPq1oFyVV4nggFgghcyZSbAw12XQzCF2s6k70tQXrt2/s2
3UNF1SC3dZMSQy/gTMA6qtKsTbrbyixqQSQHgIM7gKvpp2MdcA4NxZgES1SbJu3u
2n2WQ5/kfnsFS73ZbyKTEWFvm35lrY3JuSDaRDGY7vlRWAhldUvLWV3m8xQpCSEP
V2fJVBJ1z4cnp0Bx158hULOhGiFwwBwo/OoZPrvXU7fzbxYguHmQZZ8MEIKGgO1w
ezkJOXizJZ2lkLGbOr3HNhelTh+vyKU52MKw7qy2zPxcFHczfzV3aUEh8L+vQu1w
8nh539yxTCy3xOuNoCYexn9glFPHkzwJxEwT9QGLE8GQtUewh2HZI3OS2Da1rBVX
hGvEWNFU+0js585e9qSS0Ejztm+WHJrBOW8sej2Ur3N03bS1ZB/12WUpiDa+ppMw
X38qopNay+Q8N0t90ixcVwtvZSmQp1wcJI1zy2wCkpuUraBmOeXdWuQtxpcvOaol
KJpg7ogOyJMfJhC2eux5MfkTTpx+RzVgyCZnYgzCSNY8RkCNAexlSdfSxt3Qbaq4
WwVW3CxbuvUR2labxeE4mAiWpXidgWwftAqmP3YmTQBp5cSy9XTw60p+LcsevMKI
4M6Ls+G2/G5LPtzj7rQr3QKOJUB/VXEAadfo6CcGi86Ebi1aJdkdbsiZ75J920U1
f21W/dzKzH17GdbJmMvMXQ3H9zQTJWIm564Xm+iVt9oGBtdRHwy1zzEAZ9DdO/vT
ybY5IBm6kk/m57Kskx/hEeeoanbG+l8TIglfbiRrc1dOLwHLJ0lff6wABBJGoEWs
oiFmYZlFRUvNf9OouUpdbzfyM5aAIYBPrLixXG8bOqE5TMSxmnAyDhKsK690h01I
02Zhmbmm094Iddem7bR1dvjC2P9YWxb0qXZC7WfFa51DliKB8mcy4Tt6c1HRgUbj
31HDYjfOYq0f9rAvTdQEgi40txsW96B30MH1B780uDez0r8e7vX5Id/jl++LOtfq
Sn91W7NKAQ2XjVeoNW9ua8l8tu/9o3Mugg2uaY3MgKal4qH5JY1iyyh85K+rIS2Y
Ux6EF/R2YbOt+5WTDOH7xEtjYq9pkiHPLNiMw6ANvLFHC4CIHxavKNofiv20WKWw
8cV7+K1URX1sxGeaNZ4O8EE2Hh3n8Bf4k3YBU93RwHFVJFKKOEujWzJu5P4u9pbj
5aIZNfrSDv7sqhL6nM5+Q+7iLQVBn44yyaEJn70Wiw/8F9gwD8TPXPsZeByKyC6h
f9YQvxRn590GB8+YvhrjX3mipUCleZXLy1p37uLGC6DCtH6FSfrauhGUT28poySv
WAFvEiC2xYY28sOYyEab0cJ8JEZVwP1BSdPq+pPvK9CIHVFs1ROhQgaJ9uIT/s8A
LQO9D7NsdJhvb+S7CmfZq4uS2Xk+Vv572YoM76692bwjyCa3A5DrvKYeqX0zGq9l
t2pd8100KbDIX1npfx4OvNw3d14k8brjvJwm77244udP1yDGexP+tDhHoRuRcg6E
/eW683t0/y9nfqt6IZRd0MYHb3AOAxnQI979i0SkTZQLinqiLvcXBI80OI11q0rk
cHXwGxIqRkOt1u4B/KLwKCe0ndDEo8VSF+8UDRQ4kpak03wqjWuvr3n5PLWZVN7h
XkYWAWVbQISykiqlhuC8Z9qIWSJTYS70Pby60QdKsgEv74H15avm97ECkdht5/av
HBWVkfC+BWfzB6SNeI01JpWwI/3w08w5v32NJ6PNZLUzPvl8W6ZS9d5yzXDtC9o8
F5oxJmbaO6KQ98Z0sKY7isVMsjFvq6/HSOPdIe2fQdol28bxjhdeOCqFDT6Rn7Od
lu/IG+ggP2XNfyX2av3m7l1K1ZZ4+YkejpEUNNyhkpCN5O8/wh94v6cDXrFfkSTy
wSPGcQnb8v/+oNAIEiaTVDpWm7AtPesxcJUPa+oMxvcQk9VhJSh+yuEHaJTCTsbK
zh98EsksOHGf/F3ivlsW+YQQTI0EYXrSSd3boA5eWX1HXcLn5b6kKZFSqsq9CSiP
qawV3Jolgh/kdjIa+w4r+UTve7LdPqnmhKxlWucWIwgHHSkH3zmB1kpdYQ0L6NTT
sAHbZ+rzgDq+GYIVFNbVRUTqTXlEDK/7mOWGpjrFR5Snew5YZD7cyiRjLd8RCe+r
PMVizjm+Ai7cdSlrXCq6NW2ylog0XBeiuvIOLRuD1zhRjB/ZZzQ9baRXhVBWi5jS
dj7u85TuUhyHcxtub0kGgqUQubw1fFGlFgu3F/sg2muJcSL34IccLT/RF6qfDajy
JEZVHaqRJykNPC8iGuDMlepMHBGscdfALK1sjQE0b+fo8Ga4yAoDe6RcVdUhbHMu
wQWbFbCHkEoYljYEvRUaoT9fI6oKJDxcVVSOgExAYDbc/43WT5GFlssXpV3LTLX4
qLmVT7t3jRBwZAcQpx6ZyuQt0L2qENawhkvXwKMTpWE3m3CeMlsNjqw0tTIACzow
eI/hmTF25pBAV2Bi+OKbvZt9FwBJJcLyLJ1b6mRf/+FxpwK3L4zwl/MjNjCXrItB
Bre68Cml7WlfgJ3yAcOvajFV6XTx7N4GF2FMrjwtQCo/fpsnC5KbWCx+1u1W4jDs
WA+N6cHnCq1Nnm173V7qesBzNyc1l3xbz9W/N2I4PCmxkeXN2MNGw48cUT0XmNRA
uu4Cl4n4RFZeODwj0OAdxZiZzmMkqsYKgUBAL2+x3W6Ebj8Fi+2lpuJSdYZvkKWV
epAC0uOBimBDMfbr3N7K9HQIXVDzXZKe3FQoB2Y9aencs7d+ie+OLeD/UcJIxx2H
K+9ErSqjmyvDHSUsUdcIBCZUqS/JTZdXcFHN9YGDI8qtjymbF1uI+aabsc/DxrCe
SDl740D6rmKrbYtAh5c5z5b7MUK8WrMEPGs38EV5OHtEaiKiK/foBxJRd+UAZ5fU
GPHy9ytfD8clo4v+xxcxqkkXtjZtTpaHE3RbZmhdwAiRve6XSmUVaEv5wxlTvEw6
uxMXl3X2kvIw1e405WfTCOwT3cpuMrkeUBOcSFu45qWVto5hFMgPpaR1Q9P15tDi
C0c0/lGta+TJyODrwU162GebyOnFwin4h21ZAoRMdRHVQx3sSrsb9RHsQJbRldbL
4nIRq2hdgcBXmG+xWAvmK8TgI9rsQhqRNioMx7vPu0nuxBKr3oPpH2XUDiJqnPDm
LldpDHUZpOxFFKr41nroN6Aw6fK0roiMI4tyB/gfL2ypEfj+7Ons/NjGOqLJAo8Q
Bl+evKCOP5keu8IzFsZ7nyNc8Lt57+XIZL7hZhtlqEWAa3S8X4Lha3l8+1Gfskh3
GDC9LsGCf9QXNFufTrOLfEzgvRCGDCQVUJge6xZDyfLf9XQZvvPVgUtV7KArNA6A
rGR7hCUKlXXJunGGqDcFmu0akw0GEmZZR7ik6VuzXyg1ODtJUcdyH5btKvR8QRfg
cfPUJGCnsxSuu8kLHgJ19Ty3or/5k6k1Tlchh9vH8Xg5sUCxaZR11CYEjFPpeaP6
/PxwciGb5NS0tNjU0dbM963v//VaTS1zPB3uJYYRpV4bYMEqFbSzvUcrLuU8xjD0
Z76yB6w0EbUfbcsrkUdPFBNe02mtkNR72GfgSEs5NMvEyT35Hb26ghXPG8tTojRC
TXsJNpoIjN3NGL0ZHaFjbQPi7v5EjhlKlfH9XdIiN1MbkqJwFvHQPVdG8jiXe4hP
cjg/V1hx1BmMA3lTT9fj4tKcWpEjPX5rAWyej4vUUdT3iPdGxaWKtWOeZxPNyG4j
+ISlKnrDbCheoxr8T830C0ej6MGvWP/hLbTmM2mTHifTeINL0ofFhT7dtmwmOhpb
TGyv8PCazrPJgOzWdeNn6q1fxIWJqjm0f4w5VLW63JeChms1Se2029Iuf27WM34J
UNuW5V+r47Yd/378CjNHKS2D6FQtH/dzv2xuRDkE7627ZJxWKjOmYMT/S+XegC6K
dibqvZU0MsHCIiOClfnkt6kc4YlyCj5FarDZBGmU92WFZgS04z4K6+l+c29hx5MX
J+AZm/MFMZzA+wPtA2yLGAtJXKOv62dRr1quE9swCb1rtHO6afAOuIoCjucywhP+
AACtKV7lDxXfcJ2Ckj028Mr2ZBfrVl8LgSksVsAOZmTPbihhlnWHV/BoN4wERy8/
GDA0wv/BsJ83A1gARVcbXeSF+PlScFoEqP5nsgPBXOeiIsxWE2p2v8kV5lTlEKSf
qtgFOaI4+KSfsI7A03HZK/zIFBOQE8ajZdXXTsgcYM0Q7Mrih/aRSl2J0IxqPaaT
3ALoaeBOhgFofkLz1WkmEAR9CNnnUt2VemaU3LE5XG4Dgc70Wropp7HvW54umLHg
Qq9Ag3UpowfqJv2feKQaEV/uGkljlSEOgNr+U7qxfwz2IJ+cTwX3wtYgyDKTEoX6
6anxuEKcnYq/uyla41PS6h4B1QSQNHjAiRNsAbHsHYwiqego7zZIdW4k7S8+ZyoA
NkxaMFWoE9ItVoZ3q4JMQi6BCw2Y5hnbbpBR/1Bjp/mvNkriBx9QjxR+FsqC0sia
uajPxD/yCgz1/Zb+anAXHOaUojjvp3W5C7CypRvReTEkdIqjKrJfpI4Uyh6Iny04
GqwOpsZ6+7oGAUve3j8AkTNJVF7dELzCQEU+6MqZP/p6CLxCrEDyC7wQKv/PpA9e
3wzfs20HXRKRwnIhEmENjIGImDnz0jHi7YWf9Z5wMgTj+mdHpcDxhsr3ApCnYCEL
p1BdQ1sc6XQqvwuPzNwYWlH4tKRU0a2t1R6yYM6sjxpy1KzkUAmrBwzs2DOQk5od
KRrF+oPz8WoTtp7b8WuKxxjNf8R/VV2BAATSjSfmmjf/jyxl415ITN51r2Wz02sn
t4V8da5eHQGEcyGpfO0LR/dEXgeh3nIFjH7Ca+v5+uiZxTYFLHR586dWuwHBJUJv
sZ5IkbYrc2wprhCOEPscmnVyqPkWVDLxso5x2d4X/g/J6vsybjKUL1wFu8BViAnJ
g4YFVrfKsKBL7N3brri9sQJ3aK0b+YlTTxm0UeQpY4bC63pKE66+dBR4P9z9YMlV
ciodw339tjeK/KdaE+p92MPgP5F9xz8LDhdzh7YNgbcV+Gh4ANWYCXlB7Sl3uUS+
rw2k7fyRUUXJxCVAtZtJGZHJw/0mwYq+agR5cTDBjM7lu+xr4HgNq3oJpLn8geOz
3ixVJo373m4BNiLx0LRlO2j4QpNwp9DiWRzzUIKcJiozjkl9VJRtmfX6hc7QvWfW
2o9WuIUBgxMGFj4U1iCf4KoHXYHwRXiFrFhiPLdDJlULbo2TipllXbR1BpQM1JKD
0VlfvENc9/lBKxswc93e3R+cQaTiDh4Jik6DkfcOQ3oAOeuhhRQ6Ny+FMHKcrifT
mGAb8ycs7d8+HPdu07RHliQc3sDDJ6+/QbJyw6518O+zaF+ufIFY8lrrAIRC+Z47
pNyd2agr7+4tbBcGd80DdeEHqwRfdLuC1bvwudZO+4THBCHxrdfwZkC/Oz3sFF6P
afOo2u7KhSzjC4V8t7b/Ir8AdITEbYJ0Y9ouKcmS8ERcT1Q0CC3uYI/LiGONVf4B
Xo4bcOUtVqwmnXZrj4WltSCsnl4C9bTwPtYUbm9csDGwF2j/mDGIAUqpnb5lrEBz
yTTwKf1VdRwf0fqJtXBbWywtqvumIuFLaigHmGUjgbPziMmtxrMrEg7oYqpi0+OR
MjZg8lBS6NAsuKBM+gADqb5vj3Xw4z2r2TJefK9Q8pCn7/qjvwynAmJqtsmlEwUE
bjyJTaSE58zORMNPPaB3QP5PFWqV5IKgAKK3TeKT6SfIiencniSESnJ8wDPPMLon
/AJi43+7VyMkXhJyTJ0rKwKfoY+9LEj/fva6sYuzGBLjbbcitLq1jbNUiKiA66bI
uBtRjyVjXKIiIyWRG4DBMOXKohdviLHAB1plP8l70FMOW/R9eUmF3dv9pF0Memy6
qZU23QhJUEAJxQG6a7Lk5O3qqdZgn6He6w9zPr6PqiUZsDq7Eiv+2DIrR1JVR2PC
wVP5r3iCLnXg5sJcgR9ccXv91kLXWPykn56+0/XGe6O7HtGIrsIk2BMpUqh+0ZXA
87yYlSsEmbvuQANSEcNgq48RdSp+qjI+Ru1CK36GJAk8bcB+PbVG1iLRvitclx5W
nFAYv9h8SONDY2CLlHPbYrneJDNMlETGG95B5DS19UhMXPceql5VL9zA8YDhO2E5
Z+RjYfZCkM6tZn8Mh21P8ryixpdHqp9shYbBFKEcClgRpsMVNFzPg1O9fACe0KDB
b1462EA5uehenlPCJQ7m3bMEpRsyhH6Y1LDi5LjK+j34jsZSWAdDfvSoO9RlPMOx
xcoqBnYUzLMi4lTMRWcHEhX1pH1LBc3hjWh5g+1lAOFhHDzQLP5VaynefJpu2HHm
2en7AisSODHFwd/PL89+cCaFCF/wzvCYt+GdkZOpD4+XeHY3h6bRlPQZP/8YpqSh
1VgwjZNhkBqF6bHE2w1vduLALb5hr/aV3H55Jq8jzzn+9+mTc4RiLMhO+WC9L2Nd
qcRZ9b2LuPecx2x4zA4fgg3b0NCovhRbynUAvYiQqh+9V19dS8KCRmi4vcShLy4z
KqRricZWR076HiPKwgRr0RG9U+4h5zVPexm7I7825IsTn38Npwuv3ZFMJYQu0b0O
RJV7vnRUNsGeE3PfzfiQFxzT/E9yxrooXO9hlTSRuot24WyVG/kshlhrDbTi+P3k
D4eTMmd2n84Z8F0yPfUb1CWiB577XpQ1HCGzG1f+HYstxUGo9MQAMKn/KkVxlnC1
VQskkNMndGB16ezHxQhSCM+pPKIYGWrz3lGSum3wsNH+1x2Ib+bEPDOD5MpnnL3H
fUKexqB+Cq8/M0IL1sn/X9wasRIqxGa96H8DI1HNtZaqIYvnjoO4uL+q2rR7gjLK
qcBFCr9DHqX9HVYLcTZ65+iT0EAlRqTQ/Kx/LjZ4zqQNdg3udqsAZLCcT38XgkLK
uWrS01akCZrpPnRAwrJX21IjHII/g5rUKVBEN/MCXjxPBfs5L6SFVHAVO9rE7IEa
kyi1mzN6z3gZAMbtiLchIwY2Vo2p03fCsbHipja6V9TwJmltWSrza2Pag+tiFt+0
HzmSY04zpfvaRs9+pc77QLTj0UdpR5/zuXqqQY44v855Gdehr9Sz8zMgb+AyFS4i
gBPFd0AY4foOZYRTgQ7gqcvtXDrUv1yUPMIyU5RwO/T/f1oErVeyU9SHX7tAhJkr
tFQj0X2mF/vTdWHfW+RzR4NNwwTo97+56dXxvzDe/zniLzMMoQkBNep7Y6PJVGUi
wddhTW1njK6ylAKBh4Ygm8I4A6XPfhk1pcqB7NNb6N6O7VfTb8L7/2xL6YHjbmCO
0NXZIsvPd0wkA2/o22gPc2SiClDOxTgeGG6ZxFVD1ZA+wW8X57BZ41BzgXZUjQad
QUjKA12cjo2hF0jGj6Ti7bO/CQEjAzAC1CDat9i2GHgDgQCniBfpVVbCrKuIqBKy
Y42LUtpmOXcd0W822tlbs1IFb/Kotoo1Xe11djPoVCxuFdhOdw1m/Wo7m3IzUwNh
NBXrBdJ22+xBwjesfjY8ALZ0q1ikN+zKP0HT5aVuMUYXqCFryxEye08WD1yBSY02
9ybBiFqtBpYNRMyTckC+0cd1YsrUXar5pZFKA4P63dPolh0eak/yWyRKqdQWdOHs
v17aA9AxtzEynHpSuUsMGsse21AgnjFi1vjnqjSt8aQckvRrRCOQFffbPyKr0GC1
WXVGcabgpO+H00vp9Iqe/jYFdEaIo+4Vc2Kg9CCmlb553mg36bRO+x4vCY2yjUpn
N2ml6TNwK0D01Bm0Pk46z3ITE+Z3jK+2H1bpTAcFsbMWP1DwSIun9Ilsb0eB1DKw
fCS0GswTzK6xMO7593RShFOhnh8fk3aI8UENBBjj+MK430OxQAaxt8f396ExVI5p
2X/ZA/WzWOYQ73Fl29IaIZHC/lNeCLZWBV1nOtXnRYd3FGXagPzaPXtqjqgrxCF/
6wK2KT/J/PLm4ht6HmdtlEGW3yMl38NJ4eZLX37lERvl9mbD+sdu28AWIFg4IgNN
RLLbsc716jd2tKrRIdwFJ726ATvTSq0qsZCPlT/72ZAd4yTPK1mvn0OVTdPoUgz8
YaTEIoIW87pjfizTkXnLagiKrE9Z2t9VBFJj1J9d3gOcBUGJ6laCRoBQkWIKMz13
fKgtR3YloDdqkXmOnp4xvq1PlS1XA09O+y+ihIF2KEIwqYcXo8shxVxPR1hig5ps
MhB1UIpCsWA+9+3AULaWKNDkVsEyDh4RNr+C2b2WPpc5X7FMXq4qX6YdeuL1f3kG
x0/K5uMZm0egQ3Y2zJ9JrKqpdbGhQLXlBdRu8FCcq8DQotT+qphcBvmJHSaPA3DS
ybTD8ghCB1VhgzZXS4r78WpTbAU2WYxHeXqHotq7tu37MPSiGWba7ZewGzJO9+qW
iHN8BCWbIyCWWRkhAr1jvny1p3B2ehBa/V+lo7ne7ilA8FuVPw/VQ56EFlSJz24C
NIah8OCuyTpgq0MNxG5iAnTinZSfta8jePrSHctmrgXWDcJuk9ZjjEpvLRu3YvRQ
dpAJYe4yAs2Q6xWrX8JP8UDZXNlvdvNJqbbev7/Bbo9bt3B9JTTK2DSix+Sm6eQV
cMf2/j5CKG1jAyFRaR7852ZH/2s+B2bfuz0iqxcNV8/Ad9uzBQnZvEqt+ycjWzIJ
7txyfcvGGcWLFnvw5uP0DjAdG6mS4rDVi+r/30cBp8ESAZG92s/WXa2FdwXN5WQU
nJUX5ZS00xfJnxRVhxxKMXmoa7EAh8ob7fNHjzXDlsTd72cZUYZrfMeOl29RA4rM
WryD8kV4R608y4/jF54NSIrgHOByQM5IQ0tBBluYxs0Ymqbzd4W3SojiwXoWvrJg
6eu5Y7rYmcEtE8l1stAaK+J0fnrrAXlK3cDXhRdfUTdV5QHce0qSGEnMBSwQoKRM
V4nVO7ZvpcgUxUWY5U5h75JUFMOEy6x5Uk3303yzHDLfXxxfMirqI+cZh/IK43Rf
hMBDbjSKejqWA93dPKKrD8hE3+GitMRnEPtCuttVltMhL9wn5GbMOP+HAq4NNmXk
+53an/zJp0e4fQAuwqS/K2foD3D2q4WedRwtrCgBoKpRurlDbsgXDwpzqbcxUck9
KOA6sDj/vLlfuJlxo/i5a9JVZH8aESTJWXcrkQX76pb0uduXDfO3AJMorumaAa2m
sLTMQotpkdQu+ZIWq0XfPaK/++mC4WNu9FSCBSnRgjDCrnqrhir23WAHJfB9GWjH
23N2DSPHdITl8zadl3o/xnvhOSZeHHs4X6eMJsL40YwEBR2XBnHPnHynboPAWYo6
oqhliEJPMRbfX0MNOnf2pOGnGKGknXRDMWztc+qUzjOubNvgSANBzm2bmqgTVh65
8ktFp6k/Sy5gPeOsAw5OJYuLWZJUFzNvJcsuPN2DRBj2pQi8G3cZK73/MuBag8eQ
ysnHLLG0fol6PK5XJjR7uFBNvHBjMswEcFKgbdv4tM56o2s7Es0oZVtxVFvxK6e9
6yOgsCSpU32jyQFxYyemrZ5P8opmpdjLPCzi8o3CxgkCeVojgEyg19IUsWuDgUAs
qxS175fLrqLHQv95R7PFCfQF7RQT9BK/JekatIDDDYh3A4m7yF5eRBo0s+bGGDuR
x7uiK9DfyMx9wylehKGQziFyd+spvNPOgJuJ4YELOuJ4RiBDTH9BrjiNKIAjcDab
NQd4MVOUSfiJziP7xcU1FKmel1pnqdZ+DaYo/iu3hZpsD3v+Pgp94lWDV5aT+093
igwAHf3tRJ8LkapvV3gqZqsgDIlyiqCgYAlz8oot36edZ6vMlTxeYq8Sp5t2WDay
wm8mIhvzdqaGQgspETzDVZhZbzNTpoxQlzqbkvwF9z/E3Ax9aIYh3e7xR8szd6Qo
jvrPADUJTrgmW4XGUGUeATRZUqYZf5GuQGFN3A46e3AZcvKQteZnDBMW1FkgMlfn
ibeY/oKClhhgBxc+xKt4RokGYaU6opsDyWOZ3TlcxPmmyt4XhNwk7p0IYn0/8WvC
aIbJ/TdeQK7sKZKr3awpuPDfnGQP+yYIW0SsQ5AxbtTMFbua0xrMZoqi5l8b16jA
e9ND1LIddnpqA9CvVUq6ocQdicCp9/Vdy7VJj9RXxC42DnTsVGu+ylf1+cwpJ4eO
aoimzXINs3wKKCT4VOFrnLcRfPOHlGJRauAi8XRM/kcc9/VP9TPs3VgSgS9W8PTe
zGO+c4M5hkzD8fmJquVoeF0jGidZwRLhzviz1tcH5qzcQfr0jpgl9O2/fkGy2C3r
Wm2RZddE4bxiAuOi7oREDgcFs0OadRfnVRTCsLF/bOFomthW7y9iIaEUwOPTUH/H
i2Pf12r66UkSBFqPfYYF0KhWpBU2nP8jvbcQPI+mnQIHozmasEsvEF2lqCeUZouA
/Jmab2tjStU+amwjtsBC0J7vs3/sigxMRKd3ZxwgFsr7WSqR8Hq8V1iNYc7LwXBr
xEpMCg4S4HAd28YZRgFzZ8xFmfBqj2+GhvBSTU/oqi4G7pXnysJR3NFYlfJybm66
jgWv5OEz4UTUzFN7oKvXDtoWmlN1WwoT5CkUWQQn2FOneXoCs+dgTRV/nU44Ooc6
LPJ6PKFsncxHFd/gtxY0qc2vZU8umx6GZ1kz8nqzPvzab6AHPWHCM4iB+JeWwBTG
YQtS9VeW8yQo67wReunr7ji/FCzO0s04mQqpcELAL6Hg5Wb1klxuJ46SD0GTmjfi
GTM9AGnX8gL5zwZ5XruxZNmrkxnONcjVrZ4t0b2LLded3aPY7uKk1Cn4Q9VJmO+I
E4xtbbRXtxzrLZ6sxFt2VfJH2CGi6tnxAJCzBVs2CJTCyQm7NI2wu02M+MC99p2b
ZUFX4lDyKDoPGXAeEGjb8IWdqmIvX1wgbyWvPW9uCS99b6VSjuM1L8Icabua/Mwg
AgLYxPY9MwDVvYYS9FQrYSZAaqjg3TnEvbZSn4LO2PSKdg9DZB1pLD05SgOWjUdc
KkVvuDMBl+8n1c+JcjEnfZge9tLiVqFUThAoHUvkqMNbK4UtVY1M2tUSubRUSwmH
h/qN+/W9U+3vrrct9ca9VLAQYLv+9PRGNIa4ceBJw5/v3reXZQWJLoZovdy/pbk7
Hl+G9/Qf8bdGbpSwSG7kUWuV4955jWc1C6Rro/OBPKrwaTUdtS+8ze7khRLCKg01
anyihUgwQ8tSVepKi1wd19efvNR2z01Y9fYhspJOZlFjQRHx59kmMv2CViGFu+cX
uyVQYhikSeSwA82LaHeppOPMs+jih3u/kjd2Ii84nVpowo8uzA41+oqpFWrUU1/n
Zjn783XPEsh4wdkclJ9i3Veg7Duq/eklS5xBKLqE/Rgdsk3b9+NoswPCWPacXn6q
dZOyjDZiwdRHAyoWfXme3KMsfQ4vu/PcvIsVSZ6/IdGrBWM+tzN4iJm5ZajShVZy
VxHMSBKdcKMfL/PPsG1+Z2gLqd39OppB1xd4cmkD/xRnUL9UlbaUUVYAiAUJHGmG
66aCrid2aY9LSBJz9TJZzheHjthdgPOohPh8YrPZ1lH6wb4KOTotYSWOny20cT/b
Kmiw7CXk3hwJvzTqED+Sm9GANDR7yDvsPCoAtCr44sxoC4GXKa8+2kbALRc2A9lO
hhMVKAtsv6d/q6tm9PQ56qVbn/TvEoHum/fbnfahbVCLKZ+6TmryTpYEbBjX53Gj
8pNFm0opoxgmU+vsBG4/ZgvEpUHVLZz8P+CPg87GCvIwWr0q+Qc+1j+HlakZfpfO
zwIOkGVt1L/PpvNjTZRDS/J0W1ikRr7OoOYdKmiyjbZndzj7VTOqP4y7QstmAqq6
yJWGp+AiWL0aYOAY++ClDORUcX8h6BAH5jGj8b5RYVrwBRPPvWy5dmtsCsFmT+1X
3F5vEdtsJy+SORgGkPjyC2VB7ghvme8PZ5Gcv/Z1XMLv3/IvK9nQSd+BUg585twz
R9q244imPZwZSMYIJT/cQf+0CO0ZHSR+u7EsnJMAsPRnGV+Jq0OZTedYSJt2v+iE
L4dIuATJXWdATkfrKyqbnEj2bd5maNs6C37qwMoEPMo8imzi5qpBm6HdG16oPpgU
v+GaBrKzG81pyYEy0TXbg/9cUoloq7515PxcIm3qUZK4Ggq19RoRvlFLPgoYBddy
zehtolzTxDJc3fFbzFVvntY7cTwj/1Ephi4ySxGE5ipn0rKmoWjFWQTiVfHKdVVz
ajyliuxF7JhY8q3kFH9e7WyXCaIbTeDJoVJC+WyUcJqXO48/16VuHlIzxl9umfZy
Ndfd1MyPPQwuIEXa1g336inGEQOBR1AjTCq186liesAg/422ior4INhnw0US+okm
grIHadexWHQBKHmz5peD34nxHTrilZb0CNgBHrpufoakP2hOcyOeWXL7VHI7w/kc
ZmQv5pVa2UgrHtbfZtvHS9oKWLn9XhypGTWZtuoCy1Y4o03BNwwlVKRR2LeZGjhZ
K5r3uxxczj+KZWBTh/YFJExxlkPtNY8NEslwyq68BV11AKl7cc4JDPAgVkRXMxq8
NlsMC+n5edBXlvy/o34jfXeR5dhzzaNFNi56ssDMIPknBrY8cSYHsxv7YdsNYsHU
BO2eY/og69ayR/nbH4vm1QbacUCWv4bpuW+tsshQu6Q6GZWzqDn9DgGuTHn/Egnj
ItRXEYSYRXy+Wj1XN3Q1JeJAvjNk3BMIEMdEZXnyh6Vu+ZB4fh6lFaMd5w1vP0Dk
VJ4pcCMrhwwZdS3xKHdCu0SmTzDOnpJRokP0aPNWdL+qjBajNq+skzdNdhAWm4ps
LCtseBC0uTiMJ1YNihe0UdyvUKGfBRLA6FwutqR5iLLP+uKAP7OlOIljfyPJbUY1
0rJVDDfaKymHvL7CodUb/u3+V/yyMWbC3ZCU+mTkoNN/OHgFT1I2MBA+96NWtsOU
rdpMmtDHzcA8s+bGR9MYKjJGifIlZBE/dH24DjTCPsLe/4OAv5ZsDtaLjoEwCG0O
OwcmUrht4ICQM9I9Ran9vjG7IM+FblP28If4/RUYHnYctAWIlmeD5h78smmVZ8to
k4aZcK1C+l3CariA2pu0dKuirxuVWb1rcRxPnQbsWOmEk2pFmMybTS0ESEXBbaXL
FTFhRIWAYglQalHRuOQICtUZwi7liFkOkHrUK3bV0NQkOrvweufTRteBT6ViUuL7
L/CrEAS0CQSGcaweM+/93Yiv/wmGhXdV7o+s3vADxKJBNXIdOGecjn78z7Lrrxlp
9ZGBBmiQU9e46RZVaguIHXBTsAsTrsiL3irCe8RqQcyELItxe75NOsm8HNk0iaxf
RV+o0XUe41t+gai7QZfmb4ttjuYoULdh3WtKkNn8mTWMUJrj3rxJ+lmbhkVZ65x8
pMugpQHr7KxWcQeOLYs1p1z0C3d0WSrXqxm9IVOh7QhB5ZAP+GHc3Ydbl/LWzV3A
xfD7I/5eLRit5xVBxT0Ob4BmCK609OecY9oeBLOxpmFxafIglrhRuYiRhGVI16yR
TXF0HDGHCXTYoO6Dx5Xa/DROl/BAC1Kb2a+q4ztLmgEyA1MN+TNmS0nGWkLeinYK
jGyLZxyD1mEPJ9yJDuvsQ/i6XwbTi8Gt+wcAF2Oqp7bWu0XyanOrCO4qknl4Es3c
0BimoWkQEbYTF/6mddcbUDW8uRhwM14f2UNpzctM3kkMtWwE5YVcwsPL8cVijFHr
nMg98qxKydt+/1lUdNxQQGrb+pmz9e+3sEbV+ZengV1RySoqmklQnzNafXlchLwK
Pg3eSfeRqvRHvqaAdwNGlIrFGKEsiFzZ4lHl5I1EzO6AjZeYoBsYyAoFMeJN2tqN
X+uTo9NuFMbJu77FDSzFY476uNCgNK9iQ3q2BQz11eXvmwZrEGHa/fY4uces6jyq
nwGBOIJTnJTf1bzE5GLwsjFJENFMp5eNrfPnX3979D7qqtd1nKtCe2YP8D1ZUPBM
j9hmAExcrWkh7bk4EaP183P0kZIIkQYF/MLd5cHjxUgESZcjHhUjph0OCxrivMpl
E1ryuZEEWJRsQhIlW+RMfvCOs0SC+EDR+cV6TO/r2Tt+3yD+JqzUEj5pgH0yClLG
KOj8UNzDq3ODPoQDyZsFIzhr9PxbDxOGnjC8OlZigsUJop5XFzoCsS/dX8VyVsRk
5Y4fsbrOYAxhojmKn9oUUzheqiqQg067YTOqDiJ3clpEq4nItqkaE5d93ERzE8Km
yINP2zWg1rRS9TYdpYksnQuAgunKwJnSzLNv5HtJPs25hPmK7MNy0NX4a5XTSLVq
u9CBB6txPQijxsX2Bk1nU1b9LbbLg76Kpu5Hbe31rh38T5w4p3+fAGAZUikQ2Gl3
xrNh9Gfki8Hq+UdIVrq867afjqO7HaehAg+lTNCuGuGlQSkBuwqyK1DoDKNshMcY
Nc7htzheIqx5RcVLXEcUsAA5Is4fqH0AlGu1fUV6N2YVO2igerLjx2xhyLf99Hv+
KhreSeV2q01ptHwofKKjZHuKSBQlLMcCrrBbSp/o6OVuqnx/RYbIUKTc8afS8Cmc
FcUytnPKCoX4GAJgnsFf3nm6gwoDIKXO6R9QueDjlu4uWHUV3dcAnD0fmE9vdRhH
iWoGUXBLbNBNG4QtmRABFz8Xkl+Pl56iHmVtIdVdUZ0Q6KdUlwc/UyKfPSd0YA/7
lSawMoT2chB+MhKjME8VPyJn9W4iWVL19tRLHi8SM6mFBfe4yUYfGYJCN2K/b/yE
ahM/Kaxb/0CqYWyyyorCi5LuTNRuzzx9lRy7bkqTkIswy3LYWdPouOsy5gsCEqP5
IuMQl9L2t0XeJ3iJBpT+u03c+xFaGOZGTC5k7nPOPawjpz5GuZMypRTQxQs1nrJW
teqBBtA5FCDIZ5zMcAcQrJzIVraBGzlUO7ZcOHn00IDX7lJb6H0LTUcYHOQN5OHj
Oou95ei1QQCudY9QZhUvXS/RjsIfw7pZEubj4qPm+mg3jjTrjaBzg9iGyx2A2XSw
XOAf6SlVFdYZb5+BHLd3GiV9zFPs2qG4JdIDMl+eQYOaB5HLVnb6FqsuNA/0LX37
7ETlXRyhdvz87MEspvYIWCUzAETIU7lz7ohJkvV+dQWfIH2rj7xNvbJrKtyeCdca
yhPSqWS+jVYOXeX9zqO2QDUoijQRMqIxGcuLxC67wREoaYWshG89fYGj+mdQbjGQ
le9IEA/OQKikTwaUuUIjxkoU6nji5E4UwXtrA08DcFJjo7DJL1cJyhyPKuN72bI/
a/NYzIqspXGNFzFX0wQq0TKfLATWxHd0uz9JP4WVv4OZ+Cy/BpFyf2NvBQ2r148g
8e6cpSFguD6Sbk+Rev+XkQ5vlInJMpU56p7OplIWmj+yGLgcgw+GQui+Ct5edBlD
zwNwObCjIK1XelaWwgcvv35lUKeb+y7g0wqCw2YGWkZhK36nK9PwsEgJrQVTTP0v
xvJK4YoOxmFkrgdJGdHBbtf8S3E+o61hggi6yytzShiKArNb+qbeCY1Cuq9KEoib
xm9MqJk0eQoF118PovEuzuzPOwl4CfpCx9BGB27oDCSbnO7wbVCuPZM97rxnCVng
vRM9ezFFdNNbloaytADWebr0+lj0XcztQONn5q/SrZRZNUWFb8jqoi4SDFJyLlZ3
A6P4KVRRTxLG1uhlfm3EuT88l3SIWIktTDvAkC015RiU6K90IWx6JeqqGwf/sQ2U
5ArAp12cuJnPr49VGagmK89sHB0i2WRR0wynlRE7ApTd2WWNQ+ZF2E34noHkX+9S
4/5BcH1ahzzkEBe3wFNX56fQJzFMLt5Ru8AVZYCj+cNtF4Bu8IM7FsGI+1easry2
AiNRZLcbQ49yXAluaxDPv2g9EB1VyG5mNk6bdMMukQLb91O44tnYGbrKUfE5IMf6
TpMt8z6etZIaE9ggyO2jSyKKO2SlYJNB2qQtvgvxi20DrLFrcGeJcfqnuNb/Zb9l
uJgZZE6Q7V4xiWctuaxkdnW9j1OIKNtaf6OP84d9lJc5FzzlaE/dlazDyIbzfXoo
lP+9sHCUzpoRTlnZhbeKK6GcPNqDAQ8z+D7ENNI94U9epfm4UW8Pqx3WR5J2W2fr
bmaFUTjbqPAWHu4HVyxSn2PPEYwApwBBvc0pRs+065GXqecPFs6R5oBnSmYjQmJl
g0d2rZfjzR4JWepoxF7FmTGVUSn15vrrl2M6ui5Nzj0XTR/dJFB5+2n/EIxi7gCc
uc9HA5n9uXOFCfxUV6j3uPiHLOr5SCbud2+3cNstO4iGbwyJ0YqBc0ZFFuJMODCz
3WpyCM3DWv3AEA9G+85+wsrlG3ZbgrGLHe9LSqGudb27X7zrwSgxIIcBVBbzHZOw
2aiL8ZAEtecBBpM/UzaGjW+OO0Np1XXcMpZIN7vhWRRQWS/6d37Ku/urZ0kHDWYx
Hjd4yRF/1xkn9sP/HnOo6Usb3O+w4ll+P4BD2slpA2nJbEyDQ1dvge+4uRBXpwao
/tLrs1sMvsok8IiMF9VyqNNFKEEPHSZwJ4QX1KLg38lZ/tn+kp2ytUF/zgo7St+H
FqnblIeB7EMoeF7Ytr0UguAueVNrclOxkWKcBeQd1YkPQgsLQgpKYAEdkbHVsyiY
TSrE0+eytsdkvyGH5GH/vzu2nLh9/kKUrImPYH/tsYx1aIhJ4dJXM6r1iZFMZqbd
xAVBDG1aoa+unT0LVpAEZpVxF/giAnhsY4nBMOdJPinyAIPbSf0D5ztMClKwV2sh
ruwHc9JXbVLyH9wPmGUqbbgpC/sIOfg8Dmiruur4vZMt2tFMMOBKyvzgnfFtXFGI
X9i/h0lUJKrUxr456KxJm9YiC8X57ca4AMWUPktzaMhBBqlgy7PTf9oYFRh5ZZw/
bpDLbQ/YfUYk+vsarfxxTxTJXspXrCB+CUzMARIyV/BaI+qkLwhjaxpnUHtbxGRD
RgYRGCUlvRx4N8C3VkNUd/KmFWF2KCNibuG7Rs8Z21z30uDCc653SyNuAg1PlRV2
ZiXgFmCguzU4OhE2PmijqevXy8Q+tilYLqROr3ZAWhwg+EGN7h5SX6U8GYDaVpff
tH1wR4MZ+OY1RrC/x3tc291Dr8Gz8TGy5ekfLWI7duaIPOtsS3gbUQTtJWvYtcFV
t3U3HCZ2aSGJ8/HzHeWR6FQfm+ajsSwHmdAIEgJWceUnysZ6LbGrxWhkRKRdaZzp
mVzmsghYl0sb8h1dRix0D9+tB9eITED+T2314wzja5ht5GWkAaTVDfHMl+Opyhwe
gC/AudGYSLdLWG4/PvIeyp/dN3+JYIV70BWw+LbcJpOiAxcfJs2fcYtS+LvNaFmT
+o90ddUhwjsYFKE1gv6AROkd/AQ/CpL5kfxy70Jc2/76xKF4vpkgqvpzb0c90ymQ
6NxQkMtlVqq9FoNGLpJlMHua6Cse37GyU9SYpJerTWBCxGQVosuxL75CBFfhfCnY
Sy0KOXObdclsKI28ZigQv7BWXCdwDCDvco5PNMKGfu8PSR353JO6jBygME4oqMSg
UQxKEY01j9nYSUhGqWgrvimCz0KnKFagcz86gSG46zVWaEpx20OziL+1ucZbFMh8
XpVHxfyecuCkE5yCX/a63wVZ9GqiFRO+8PESsFijZpCB2nv9oWnkXPcfyFDnCVv0
dvDlFtNCLPPeoqzTMnIudDOsQXNjAgkbrVtP7C4z6JC9439XUTjsuatLVHxLDIXk
/4bNl0nzTYbIUEl0ZL3KACkoyqOJMt05vaEeEEf0JqMpyyp+LDodqljXWRK8LlV0
Z4ffUG08oyHgK00VS2UPHOcDv8jHWu34s0kRZDPrNbFhVctZxfTpdYbD1GnY5Gqu
DjS6MT4XuL2qHkEJdp57yz4QUsgCdpdK7SOuiZqgIkR3+pajet9WwIxZHaaM6J8R
F2QC8Bc9fzp1k1vKDpl634CEarKyeKpYO/MYrW++yFrKjbPVbZmgUJGLTIEyxrFx
glGIvMaZtKy9/te5HPq8oQiZJvoUl/UsjIOvNozynnL63aTjFWZngucC0+s/E6QA
wm+0MgJ1iqVip/Fbt1UAXiaCgqk6jSiNfsClbY2mW+7h22qq0+B+85EYJZ101FsF
eoPh6VQjByPv2cDi39wAV01UmbajFF2J3LCEpDzLClrwQ5sU2Ra4Kme6E3g02PJ6
LM5vD2hus4HVje0Iw/OuZlzjaJsBMecI8WACcxmqXLnGiOdOvsxf/4bNuzD6DsCS
1zghW8qTpZqyTuoyGvimX7SsV0hf8enr1vTG1e3E9puWQGX1ePScT3feYLIVisM0
Ok7LMg/0ZEbNKMuhYNr5ASrjDc7bQG5CRib/fq+ecBwYabuSymGYjNO+eG5Uv92t
UGjhcAN1d0PB0XmFPn4tqv8FDAjpyrXBVrK5D7E2Uc7+UavnySuJJM7wjo9yVcAY
XhpeT6Wcts25xU3ZUIq/G6s7ba2XW8IA+to6MUP/i7AOpS8u69e+A++1aY+IB2AO
sZ+W/qKBk6g2ONd+htdlClwrHjHqsyDhfxiqKcjv77K8Zwdd3TRw1hNok8plcp40
mqdHt7Y70srEitCqjmqThnhRgWyKnC5va9/Qn4ct8EU7S5um7TP1OI/8aLNeCH/d
UmM96jpOX44OKIkpoxC+Te7bNOtnm2exDY+btL5endXgL7PYfZ0A+mXT9kty5DVA
uuYu3p+SIZmOclORt3mgiHANLdj9tmFoGqKxQOi5e3WZ9SCacyucofY7MJjYWQYY
6tHsN4wpa1/o62HIBUAKpdCA8HdH6mMb3JdABO1No9MUbpyXqSaBJSe8kfqyRWGG
ZSOqaVdqZ+bYFtTy/zk0s5xNA/7mPJhlxGhFKtir1rMh48CQLYDV0wcj8IFyVk+U
0pjCcQjzV4nZoJyIlGVna1aWQ92UkAPXV2w3nZgpvNtzg6OoutCgf7tRcMWFRRA4
YxLsb55mqJLHPATS4SRQKUB8p98hrsVKyqKFFVbZegQ=
`protect END_PROTECTED
