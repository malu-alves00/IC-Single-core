`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KTyGZIVQeo49yNQp9tLOaNt60RiOeNLBFnXixrAMLKHA2rzcPABzDZ2VT4HLGhWs
ixQrlN7IOGzLVY4j7MJtzx8qAXDn4kRBs9kXA/YzgLWl7whuzpYgIMsHEqNb2EW3
73rLi0He15NFCfYLgoOF1u6RRCrutv82I99oTxV1upjvPGpaTVGOuWsuIrOCc2ci
20F2PRemcqTEejR1nCAC8SO1fp2MNr1Vbf5/PpXqzdLlHvA7gbTxrCG25mC21H6d
QbxjTHQkZ8PPRaGgYqQJ/g==
`protect END_PROTECTED
