`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cDTJqUhYVF763NuVLE/dAjGcR0/+3mv5tiWV9lcLQCuIczmj+zLPZ6z1YhbYy/AX
AiTEWro6KLTtW98fr/v/sKAVe6Fz2bsJ7xvLl9v7U/e8FGKB+RCW40I+W2HK/gw/
WbI9/P9u4SCDFGykI0AGxZDze2CyzhwCtv1e9+j+TdkNu0f/t6Rl15OGfuHR8fQt
LyJRPiNkVZ1HsX9nkSg/rGWyyyRDi/SdDHgaalasIab+bAtPcuT5gsFSA4nKvMRh
BBjxoeETlkQjl8lsVKuyBJx1wWyzH0znZzJryR9bjYDHT4Lxr+LPgRA2JiXDBi6B
mGtlNSsSTRGZGUkCV2CD26OrFegO7QJ094Nee2Bwmsa8Hir6xHlAvCHeLVAQ4rhT
Uo2t7nhkL4V9Vd1mwlxbKZ+qYvJuu6O5PdY+X+KkXy0TQ4qFDR6QCiL5VGJm98GD
iGbF7DRdg0JDsQSXeKMb2wxniSx1k6M6MatM91lbaNfZkwCpwmdypnLb+TXWwKmN
Rc2J79W21+XfTFlslg3uBWhI1ouaHumN5DfWaP3p7YkHEtenwIUXofCTs591t85V
S3Es8lJuVeh5Iu/pKL07a5EB+ABLDy70zqHy/kq82RGXbj0tmfXEXfi3jgv1fB7M
ZGhOds0gD1TRwNx3aYJwtGxI0y+RYHcVGVfEfyPg8K2ynOeXjKq9n3vXj9lA5Yo1
yDybRqLWIPSTeWO1sJJnoU8jnTvhc2aU4WrkBCBwDiRFed6SmUenmYzuqzQmFK5P
wgZrcdC0vvSL86CkQ0gycGxn0oTK3TQZ0kuE6E3+UAaC0ZZzi7SWiKIuONNVMfno
FwgrMUwMz6OKzSYfSPn7Bb7rRIvrjTvHQG/Z9fK5acAEgwLdvTxJXZmtdjj2GVrl
mL4xtmaMdH3hzv/dXC3RDhHoNq2I6gv4/vbB6LPiyon/m4tDjflg2uQQ91HX/N8Q
`protect END_PROTECTED
