`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bLI7OfvmlUbdn0KFTN5i5e7GMFh+uyQ5EPEkWfliXr38PAGMXU//5W1wkd62n9FA
ydlH2r4ke/1S0YawCWSQmcdGueHO39sUnhLMIv6k0EFsPMqRZDwZpljinddzIjQH
Tw/ISzlrHtlMVY/tA5fl6LFhrA1DPrwC4jAxbX78b8ZTI0svcDDmQJEMkJYp73QX
l5xKF9SCK6xn1sjQaffp4k+qffdJV7DGKtYKPPizHuX5l5vXYMqCuE2OZ10P6NgM
U/ilQprm3hcUaQvBU5SGqdl8xssBerv8RaW2wCdhk5N+FfFhUc/ll/zkRwbX/4HW
ljVzfms9UGflbpZrLzATsnCpfS9QM8suD2qnjcxx/Pxl0DRNwwyaqwlOCqppK15E
x4QObmY5Lc0OhYlpIpqfSxGtkioTFlKwk4tkrGOThN2NA6HW16bfHT3id/jvi4NP
kabw03Z1lsn03BFru9YQix5hpU9g4B5jOMEv76vW0zIk6Z+bAdVBiTrXz0u1ZF8j
oR00mekzun6I9kF6w8/ZRQmyiB5FqQOfH+am/r/oL8n+vQp5tnJGD8SVX8W8kuun
6+GC9zIO3H9YQ357u04ray6q4+OEHszHNPK+1PlsRPlwyWLR8Q++3N5I1HC54wYi
5+6h57d4V6N5SC8MIchxriDXqHp2PX3TnRSe1uuLnrFrkppmiereq3jPmovDibxK
aeLBrrA95/pyCSUtCg48PRZKXF3Hr+erVuS0+3zsn4Wfm0YEt8CfBIElqgil4juY
ceytKe1io4IdAj+fnjVl7hKH8ZBmsSWG2wDxjzUe6fxuZWnMKmnUZQOKyOMDoADL
SED1VoU1IaTeEMBcfdZtwvfjVA3K24TFSkkc+m8neJofL5sw6RdLyE+fb9gIgD/b
vDNdtwzIZPeJ4RJBWy140vfGX6Qm9Uv1Vx4DFoZ2t88qrtBN0f7wTjXGGyRP00W0
+Y3DNlsBaKTzKaN5EkJqEcWChnDUcr28tbEYMFKbLMSorBl6UXfV48lXzJmXBRSO
rnQmzzO1i22Gq5f6p4Cojh73qhR33KBTFVqoNIEld1/YttVZIZNCeGhJPGjY8Xun
lZ0911467eUwz/rRlWkgcBkcAoBEVMwcs2eOyAXA7uGND0en9cOB7JzlnofPniYk
EMc+RIgOoZPaVzQ53Ed+Z9eXQroJ5FRcHfsQVZ+aPbYF6imeJFwn4rsrzo55/cYR
qPCSnwqE3CrEHfUUR6wA4me59ViersBq81NNcGf4nLTsNAI/q/LCvvRj2fSLmgsJ
Kvuej/oLxwBlgH9R5LcaCSck9SkVP8ELMF5LVwlLYVUIRxLuafYgM5K/wGTl3ZSL
84UfNVehMVSpusBkDTbHejN36pcrKLZ2Rsbr53mXVqpitjQu43U72JRSzy5BQiX0
v/FWnH0Ct/+tAhqKrH+ZoqfA2ooorACAilPSwXYoUx/qmhCbWs+YOUXoeYQZpbNb
seD8aLAMR8CLk/AnyDEPz7TgSlNBkoqEr5ToCRk/XChFkIC5NEA1AQJlY0J9sf9b
B2LiTpLiMAsCL3bLbeHIKoYMw5hIxPfsRa3KLLx76mhrw7shMsz/7KPUgz7KsEiG
L5Djw90bpgUbcrUdILV5wlxtVCeTnP0Ldppf2I2Tyv4ItcXUI0hLSeiAJcRvD7Ox
BUBmsNMpPVlm91yW9Org2INsM9N+nQ+KmafM1hEes81gHcFAYQt+W3X8sRygX6lo
tTkAslJBPmEx6TalPKOI8UAtvrgEqzhX5k2tQXe4rt4ARanVp9gtPWBrP3sfW7rJ
j3LJ9LGMFD6DZ3+qNR44AN0q7tp1p0Tj3pVc/WaCd7ouGMnq88YL7DDYxu4wcpIu
Prj4U36CRWnqVtI5DPK7w4MDyVmaqRohjFtUASrBWrJsei5KYgTwf9wntdIFkaT1
pPIbbhltrDZ6Ab+T/jleCwOr0KMFR10K+Xg1EbiXokrsYC0D1R4ztPaPjzUTvNe/
aAyFWUn6mqZ44ZR/U6YvFoYKLhIMsFyjPNYSEx0tEReiwECoT5IeuEhMuLAcV0Es
UaoZXhFWgAuCMeBGWso+A5KzZ0H0SxR5nLlERKiVctAnfqzrkU4YtsJ9ksuBYT6C
Yvxo5s/oBYYlhEWI6fVd2GkP7jDVg4xJ+iHN/1JB16VuQlfZ6u+YsqvS4Ryd8s2c
151SQWi+TSebzv4loAbB46bXdAKnvtb1UXKiTknit6iZmSSImmHsdweu05XpkoT4
RQd1/sHKP117kab7nG3/GAhtQfeGs684fnI/ZdbuQYzunVsPQeVbT3ufAv90h7Nj
pvT2HW9iiaLjN3Jn+pyudjkA51NLX7FMZt2L5YbluSW1M3BjE3lNl9ny+HItL/+f
jMMI75166Il1osphUa0nVM1NrMAvrAZshOkGiEVQa4ibR8mqnNU9YfO5kEipACuP
UjyIkc8G/tD4pO5VaUhFiZc2rPUmdIKFcGTndc+0W0ca/8RVj5F6TxnV0Clf1svo
Xx6tD63TpW5LcdD/hgs7EHvUSCO5yU0wJQ08FgcmwS6bFV74TrXidRjwfjHcNzso
u/RxRJSdug7YTQ1/ygY3V+RDP3B/eyqGDX1t5PvD3wsTe4fDciEl7G5UnWvQX87s
SGOWeq1h3iMtQSScH5v8Lm1O8t9EitsLM+h6jd7+tcYOO/geYAvuLUgWyRROO3Ka
wqxpGoP5TsfSdlwvZpSHPr8CUwpAaEk3SEcdPFuACFmZcy4AyLYfj55Uzk5pJKIX
2lwPkiVbK0l2hmlsO0LTkGq5uuYEDZXyH/+MJfwkYJ06hrWYq/IVlkJGxP38AHdO
u2CVajBAlQMhiD1w0E/bu2rDXRfR4My07Cc39j28vCNvUBgSCm/tJyy13jsZ+VIP
P69lKsviVLDSrPWg1xaaHeJYf9LUD9NvVc+Z0RK2qOnmYrkTu4BVYJ7P0Hek/BnG
MjTJ4UhW8z2bYRHW1vDgyXbr+bLVqSudLlWn/epEak3ebJBFb7MpBEsHBr1G/miE
nwtN9IMVo+oLob9rCJUXEt4rmwg8Dz5BZ64+eRX7tLh7Kco0Fh+5kr4uOjRmnmn0
0DXS+VvKn9zF3P/q6IW6PN8jOKUBlrAaVx1MHxBQL0g6tCLJgxUL6gjcu9gzadM6
yCwoAygfsbn/Mn5BP4M1v4MgcB849puzbE+RlNa8Yyf/ZcX4tmqMap5V/u0zcTrp
97GYtqJc5xGCB8uyeEfErvzp/o8CMYi61lnaSH9pTuR1uYAxCEa6pyZgd3gpMNWR
6M4JWMh/mAON6iXO/kKXQr2AlMZJUJiDCC0EooSIDYt5sgRZOJiZzhN3plfj8HDq
/IH67zFtzGBp3PrYMM3TSyuTK2b8lmyqF+gBEIT2ZwQUCryj4NE2xgO1ypthnQLE
9shvWJBwxvR/EuPTP2VGmQTHhxLYuPuiXRjqRg7BL4SP9VD+GDewFhfwry6l5akZ
ACdtSRH0O3iyoHG7/9N2nUD5k+S2IWrrJSxYSWsMiSKm+nfjo7haWP9o5eKznmay
//2olrYkA+1OTB9bXK84xRH9Y11uy0E3b7qUQgJK3y77xcfW/NZPv7kG/P/WDNR8
FZu1N50LpGzVOQgM4scWYGwYhyqx96ZHXoqnqt7TOjlkSbuGNnTQVdIzeHt6c6Jx
rz/Cv6XVs7FDtPPNcbSzXbNbHachrOA1zxanqi0xIF+1Mqb3p6CLmSIWqVxxC5bW
qZJSEHiNYvpfw9JW5+X5Ip6a1w2w9s85qoHnx0FZ270cqHRW3KJqk1rYOMuJ2mAZ
vC6T86iHntJj8w5hIyH/l9SIV34lDgHFIVXtdko8wyqXmnQvhKsuDTvQKkD3gl9m
L8Og2FxKlZXnE4heWcsr8OkQVlO0oTttvZu5qRh5JBZtNiQwDX98OMFReKCAci6C
dloKZmVL7tS/GIfHjEhs5aekLDcoPPpMMwvXVHY9UvtytEIFthRsGf++iYJ4H13u
myZiQFwZnKrACV5L1m4HTE9B5nny6PQT4lNqL2JmWjiIwdoY71y3oZ6HF6adeDrZ
V1tlbW5LABCwxBYrMUr5W2HBUnC3y/M8oM4MUAIRAJjHMCvse3IsXPvwMNQRTdBG
ErJ/bZSKtQBSPIgpaS6mTJ7IuheB72wcyrFgXvwNV95VsmPwRQMjkQAMOkuY7k3j
bUz2oHNgEkMaFze3hC58n0yOOGiQ3SrbpE/ZpLX6bNEMejICA7Kv13nU3+yFCqy3
cmj99Kq3QilCXDeLKGhsIPQ0SvOfU5hvBM8tnXYoQ7aCwO16iKn1tQnP6AkZlTML
`protect END_PROTECTED
