`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pDRlSjQEsWXaOg057OVC80yoXqTZcrVLDzKZLaJxKefq8ee8NIwEKtZpqh9R2Gss
wqTfopF5pnlBCcpAn0mb3FsVTpytzpy+PUAURf2mlVanOouMIdOrVYlFylFNkzTW
AWljW3mIZMSPZ/4ksVsU+CAmNmHO7wvA6YgOb2tMvCUMqnTXFHLJIbmtlaPIGB9y
tRY4LwB70s96pKlwtPYOQUj1urPwVc8FYqQRcfwKelw4ThuTFahjqVEKJQVtxuUv
jDI0p5Rq7RKCDwvPwr0OkkHIVh2JIsGCb73KYZ3CoJ7v0Zd/KS75PdP/WBuddK2/
P2CbcOu5Q+ErXEPtb99pslq3ILc56CHTkpNU1+Z/NdKsj1EvfKF+k5RvXWyPPUQo
5zn2BGLnrFWNNV78JarhKiny41SMy9K3ukscs4sg0XFOuAXjdeUoscpIEmRUhro6
43dh9TNfp0QTG3KwGUqVeTsljlbyk79bJWDA3Du+IgJv7iI2LcgIiQuT2xY1LjTX
q1uyZSnla7mmCKnOi76npb/WTmtnsVAdrCzWr0CtV4fXioADpjafG65UyMW23B/c
97CzL3Df1r759LuZbngP6oCdXOITD3DYmxYkJslnARDZGlfPKi8o5lQ3sTw1qOnF
XYa0k8UtjPnHUFVhYGKcacqY37JJlWwI9X2H8a53ZOsDmlwlpsgwu1BKdmgnb7lI
+yx2P0ZMkD+5JEUaKli9sTs3DJMLxCv2SM1Tuqsd7o147TZRQmO+qsW1ZDMIqVqt
66yPygksq8WX5WGqK45tWiWcECg9rYEUr7WgkDS7FuC7ZeOo6uc9BGT4pEI/M7Fv
1kKDFzbsL0MVxn2tmIBspZPAbRFE95j+P5xNxrM0XGwLkYsGBQ7La3Tj0XRnp3bt
+ZimymemwN0TUd1cYGU5ZQNAPD7Ym0hK3InblxknJ0HVUBNCVOJc3yGmoKKaetOK
r+Elt/oNcQyTHGZ1PdPvSWoBCvHf0Ludwef+5Irx0U1emZ7hMiyBHiqmQqp1RZM6
8B0sTNGqFQeEkw7TPr+4XxaeCtmjZaCZq/WSgyAOxVlQykHgYzLWxA/KBuAqUjJR
gvSg/s8bhhwENlJPVzQXmu+NTwzD+U73HwRno+DTaSvp5T3hXP1N1u7SgWf4RDn2
EHRJdukoxuHJVbBsf6ku1jzfRjVr652iKBDugkB1vXmBL1FnXiaWAaDlEEzWRSZx
PlBgR3xU//1Q6BhEVXHI9DwYfRFwKLdP86+Xi2T+TixjR7b+nebjl4spFC5T6wA7
`protect END_PROTECTED
