`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FbFXeaL1NloGNwz55mvWq9c4plX161S8E7Nj9tKDv0nelsR4LNrnBtrnuzgJo9fh
hLjVDAUU3GzvhND0qogAYcGYDe/x5X0jp2MLjTJ6rtvTa/lGl4We1de9+sjbMYM+
L2DiD66tpcanEi6prwelLNZZYemenUi7Pn5a5XTxwTuSrZ8qGeUmnOwrjRYKMK3+
li2ikeQowwnaEMtmGwStsaNl6WKrl/2bqhGfhCS8hw6//LElYuCoS2S4RXEu5zho
DOoZOw+ZxMKH7N5Tfu84gmjWWLiCQoRnrNx9nU1M07Lqdjg4CsZy2wKXJ6/Q3r1l
C9eNqUtH9K2KKedMfJyFXdT0lfrFVnRb+PbQgCTWBlSnB/Jyj7vA1PxNcjC43ImR
tFHtocIOhJvv31C/QTpdw93QwtbQ4x3450eMA2xq6r4YK5OPutUn48J7lxwCaShm
UMXHLGQvlr3hEYCgbhAqsJV8UWkj1hxHB7qAswxCt/dj+HotjxoMktvLFvvTadwj
31tdpGM3AHhNBamDYhpO3CdEzAhv3a0KyuAZr92UufzgjHYFZG0KkBVgfUWk0R9x
vzXA9TO+y8Ejjp9Fbt7YsPj+80NoWxPqLpNXkewfVrKM4jvc8HL3FKOn1Pw9/sKL
W94OyAqArDIzCx8oefBNf0pzpeL+nhqI0KaU3ZGZsnktpnLx3TU1Fayhf6kKclUS
3rXdkq4dG/vkqf4DT0tP6g7gRnRSNEwPfL1QTJHwWlJANPHJKeCkTJ26dYd1vgJ8
wM8Ka+uzlUs88nQBrkXjiIGoACKfejyFS1gImyn28ds=
`protect END_PROTECTED
