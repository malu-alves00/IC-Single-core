`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
htv8AEa/l5pCs8Y8onWWuf+jKxHzhOBSnl/2pR+BAB5C/LBe2PZrZp3OnXD7x4rx
QITnAbUR863h1dBkhJKDUbLMHl7vazQ7ReGN/P3gkFLwS5mUd6AGuTLQA2CaKKmJ
0a+0M3nXKeX4OB2jBsFVkjOuZK+iqdH2oMCjT7Zf922DqqDE2LBM9IRY5kLRV75l
WQN0xmzVNGzKnkLv/kl+L43BkO6wBgDN8NuxUTLgCG+J4XZXEljmsT+xLUsyYnIn
Uu413UxbTzaz8oQwjAaHiu8QLiziOhK3aZ3Zs5f/XMIL2XIvNuYtiCtGKcRAbl8K
jNyC4hjZpwai5R4HnNKD/2/UgCxoGTyaet/wOBnn9exl89eNBIPF0qvB7+OiKcta
QGaudMmCt8NvdWrUOBwoKw7B/tCui3BgjM8E6jFQ52M7roCm79alEhM1u7+h/nAA
5+lTK+QPAgHFkWBdYeR23BfaBlim8gNyLHOrFH3uzEZJh/xcTEMw5pvxYAGVh0ux
nGLeRLBHjQlX1ZVmw5USoZNzzz0G/jEdSZpRe+NbCjeNgXw3zmRmwC1vVVmZ9iDr
CtWO7/b+42m2O2gt25I5Lj764zXS0DRfMVXZfh5LF+zFcGdwkpfZyF1TgmguiUfp
Avr4Jbfpo5VxftXavmAgiHQw36EHbNdj6SlY1G6sr0drJEt+l2Y8DjcY+YKSaqOS
Sb93UZqESl5E2SQVrUhz72Id2eXUMrU/vjj2il5pqQj3Kdtfz9W2AXpmmmX/0Wwl
j5hUPE5B+f0+w1jcC+z21gmqVHWmSbTzuF3fP2LrS3ouChCDTigjfZozAoATiAnY
wjK6y9xv78fmTCKTAZS+AHEwX5+Mp51i0GLRH5FCtPJv5AxXhCU6y8eaDnAlUgur
9CYCmW3begHoHedS9ZuAa20hgHyMUN3OyKsxp70gTEuIqm4emsu1lBfA7RH5Dg85
BiLXvlypdS9lAzR5D1faQTyFPnmpDIDXIN+xBQ618G2Xy06tfZN6GqjPuHV/biD6
msPCuCAYY87uoDyz3T74W/N1TyKDv9dNqLZP5/q3gU0xPJxwdVTzzHRbKLtEgHRE
4af04KyH2p0wjcfNZp7mUXobHiKfjfM+B7o/9ilenV8i+mPYGR7aI0iz2SsxhouR
Ds9iVV/u2XKr0X/OcBZ33FyiEvAlfP0+Ss56b6x9nLgfbB2JEDn9EQwCp24SnbDH
`protect END_PROTECTED
