`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7N31xGXXdfxlNpP6aQ/mkzwKAoQOJ/pD0UxE4L3rs13KkQZS6oxdekQjTOtuXQcy
ajDmCgwlEcdCW2JlBEn1owX3H9e+PNgb1fDcK74IyDl6LDvzO5TPV5KdsfIwgBae
6WAdVV5G4dSCRRtSyPXq4OjLRPbgbaamjMrMf/9dukXq8HDGXbTQj8EIIsnCHhsN
kmAwmqVGLe7vIu3BsT8ri5b6oC38cE2yLPlFgGe+ap5vO+xfHkgFl8EJfE7j4gKP
bPWDKeG/mQGzggF9ta6pSzxkxzLhNJbLTDWN7drnjc5OYbDlcShBzxiYM9DF+ac8
M/hHxzf7rP2ZkYpkMpuJNwa6DXExhw+HKzq+Dhi62R1aJh1orkLwSs9my4rE611G
XAMwkoG+O8Qp3tjGMQcKw/BBaawtWWvm77p7eP6xjouWxYDi/8pPq631hMq6tioK
pllpginhB29GqsUl+l9V73+aNaXvnazLNmFwvSEE/nLTvkd2dWViDhldB0dqwYL8
S72+hgpvIoyK9qNO/JZu9Z+1pVUKYqd1m5SA8jwq3m6aSyNVQxMVpvUA5XnqgAnw
FM1rb62BewJvefuY7Mg4TxJE3GP+KnVAFRRlXE8XwhAod3cxngPfI8QugIDkQSr1
8UAmRfm9mfu4+gvvuseTmMH1GvgekGPkf88qqAGqvDMipv5+mZ8mBOrl9kcujMBr
OZKZTQ+GM7qqG0/06Vpj1RBRe3tetugnBGipilxSFd8SMBfLRo7QlNL23ckQ/kcw
4bkoYJhNvrnH4SVFjsOWiBYH95u+AOcxulT44FVH5PFskUWLiyJw7au/VUlRtp/Y
MyzI1d+JeBiDZm9ejUFcCLoSPIHflfLtgt9f24GnY6OO3W9uN4F9C7WINVM+AcD+
PbF9QjF8WKWGgDeXTf9ZJeTkvJfCtDI+JQlHUzvwlbo62yFGp5t01UqsSIBISxZ9
STUDGaWC5i4rT3ExS8gESE9SBa0B3vcpLlFSvM37nGcHMs5rs8YG4YgtrEY/xqql
2c5XXj8Qhlre3HDjlMKBuO8NsyoNfh5IPadGQ7YaJrqErCD18qirNsc+ektXxITA
fER/4dsD/FeY8jjPsGneno16UY5Xx76fepnnxOZKhUcYggltvs1Ao3fAac7J35+w
kdojkvgjkTGAESQ9rgZdkMpYFV2EzLAHyd2yc6wZIbSyc0WJ+6gz1vT7McXDI1cR
NB/skZObYVtkEXMbObniOIU6plEfEG6Exqj0rdsH3SNTjKZjl0GgtovGiFmqp2xj
rdKZyAkGv8rzFoMO4YOrjlDfnxbzpZooAaPlqEZpCTEvqHYwM7XOEpV02ty5VLLK
pDCoD2u0iHsCOmM1DL3LDNb4sDFFGdlLW52xDEb4JxTKr+S1Cf5vwf26uK7zpsZy
Dqs7KAnJFw48hfgGCcWmKi4hh+SxZRaALzK1hTH9LGi8JIPluarLW2IiVklH64mP
LX9UJEO08ijo0nCJpFm0H/hxi+C33jSAoIih61Fg942BlRfdOVadfaqLJLsUSPl6
MS7Dst8xehuP9r3TQvbh1HHvSqfUhC5HHhV1+1FpPuzQeS6Y7HYZRu0Ji43tdK+y
6izKQZzVPH3QpIKmeqivPU6tOBa81a8Nhfd2oPSCDTUAqIaM7qQaVNbZPGMWnJkH
WfLLEHMhL0MhEeR41Dt4juav1ki7TyIGKGs4PxBpsKV80ONbDYSaCJyYtgVDEIaJ
FgvXsvkOeoTjyEeU5GFQse8icrJZsStmIPYoxqogI9awLQlfYmTjgiy1N8bHkML0
GhIjQY+uRRJmuWw3QFBk0WvarBIabu4P11Ewbho8gCaRlSHJdtgdYnMht2787taz
+x4677WG8DFVbtAtIJVTamk4XEHMN8htIv932vX/hBApzFBTPRfkuXR69kTSyT5b
ooWzhxFxXqnUh1ooVl0zekeA43TSyosRicFKdCnuFt3Zw7DAPjNteZd+ueF90U7A
yI7pbxy6dVVoiw0/gkcL4iHebsfZGlk15fQlAMiR7c31g83p7ApU2zNhd2K/3zSV
9C+EN9G9mIF98JL52Y/kaBXy7SnjMoXbzU4XxL8fs0ejqfWSpoimzVaGbsI0Q21R
po9ljH8ulXS+758sBddEv6+CzZRt9J58WXRRMqVrAcA5xQ56hER4OLYShwfenWph
Cjzf9jfGMy/eZtfmmff9PH6jV5GHNssnH4l48w0Foq8uoL2ddPeph21e+py/6tOL
jQ6Gc8KOKVXHbLG7LHzSwT/HWvPlhZnAyMQKv8ak3hzCSj3/wmEa89T5++8ftL9L
uOZRMfkQXsNR9LbW1bdGqOqvirchPzuynKToD1siynuJzC432DL2+YbR1DaVpOD2
t/yoD/SB5+lGd9F7RJ7GhX0hw4+PnXKFS5DXK1MW93HzHqZ+tJ1GWflRjiZvVHuj
vRZZtM4RIDqTAX/P6RffueYqxl5zXZ8ai6HqKH4sRAxfIftfGFTiZWYivUHqviCB
Fi3S20UwcjP5L1D4ZOihwaQX0SvbhXKDMVFQjmWUR/YpZ5e+hUb2tybHPTJcxwND
r0nWZpy8V4KJEli3HBEvBENPnnAHE18qsVmHarLi5/Tz4bsHB0AgyjE6RMDd9hNu
2bCcRSvsfT1RcK+Acl0o94/x4sdsU3uO1hDqDRMRP9uf2cTpw/hqHRwOWJOUxxHo
aBYe1WHvu9Lzzm7SpEqS/S1v+3/ulUZCRZ9/NQXpbqOOonY83yKvBa2XzJ1ZOqDr
PsmCAiMn4PyLlzcc5urJifjh/k2po5xoxwBQKux0olkPNPs9Ce8PLPTX3w+XcwTx
C56++RC3zJ/wT/b3Araho5dZK28Sl8EQPeFPIgNjHhBiOQuBAgjKNX7qF1PVeG/2
df23B5NaCrNVkMX2JeNP3OTfvmmBtmrhZBSWiuS/5U7zsilllEe7DOPFGvXHclD0
KhmhbJtke8z/3EVQUrNc9xMuT1wZs98tpAOtNvNTzt4kBTE1GZU1YyIkfP59RGsH
mGNhNQEC4BAlEnqo0b0iydAtMA7I6NmuV5f1VFfUA6EnjWUD4U6D0mAbRyk4mobH
NG3592jc5U/fSMGh8hX1E4bRQZ2OEybyww2+j5xNNWp8w0BF6nwr6ZA7nOzUToiS
65fibCb4d1e/SBu0Jbau0Vwys89JEt+qTk0cVI2Gd0mmWxRCoAogMiTlL+XLLPAM
gubS4nZKI5Gos0Fl0iDOCeGZwNRIGnT2sc9fZRqri1cUbKhXIMISk/1xAAUsmMug
luZ4Br13RdSHzko+fxpPgagAGBiwBvTcgO4ibOQ2W5F/2i/7mL9YPN3SzDZDkgW2
YjvvWWth2CKekyWzbo7O3tpxsbWCJxE+zzb+SqqhQHgXVPHaELU1bgluHffU+OFE
XIO7OqoChcpl0kY02siS63Ye3bvWLmugY2eDlvfUD9PfgsDM4Rb5vRY3W3Mtbker
igCKXtbNTdnu1Jw+Ke9fqEMipEYdvUpjm1U3HJs03Z43Qo4HVBTeXGozOwNmyRNg
UhkFDIPlitqlzlonLbz+5Qf8ACLvJP7pV5BTHaCr65pttBRV3+9P9LwvfRtMUGKS
Ix9XGU1WqPa9BO6Y1YtCMeLS+mTLsw+U3t5OZEpEpMFTJNnCnkipoqHHmule1o2h
bPxf+sHc+QZxKtlaQOEcoUEWTcnH+ww6wclndcFxMsxDrnzpH1O5P15FiLNDiUz3
XwkXQvY4kTmTZEjbbtcmSlCYhGNDGH9PNXlf4sqXusvvrcJFpXgLRl8Rokg1mEt5
zzp/0sOkKIXSyU/l1mZ3mvNXzVKmg43vO1y6kd7CNrKwaQ2GXFaRsruagv/DmZiy
lYQZz57N/kjxeHbL3iesZD99pYbpzhTkzdqMPgm+LrdXGs4O/sMYXIEuW62DloYL
Ke4tfMY+B0s7zyH0swacHsglrekZe9kpPVPmobUpb80sOfWdfG/IsX40vxHgbwB0
h6wIMwqD/83sdbEuaUHkVUWAgdvoHpKrKzF4ruFpsnqTXwIERWSeE/ExffOUPXVN
iC5Nqp4Ac3u+NHr8IgDb8nDGXFmNJyvlhlWyLrjtE4VNHwPimn1zzrM2gMdvY8c3
vnzE1PG5bajKfGYDX6GwP77KzVzdc0zJeGwakNlKmCJChzNtVVaMIi76NA2nQtfr
G/Izf/j5pYGZv3BL6Y9xZJgfv2cwLNkUsCwfrD7GVxtm2eB3PdgY9ymx2BD6L5oG
UciFDCSNCEuNwWW1mH0dKwZhYCdChEYxNnpme2CHf1mDhMwxNgNJCQLaUoQkHhXR
1TrpyAWvllPpUFmf04ks+N07LeZLhm3Ehn+WukbLadkm3n3LaLpA7IvDDwx+0lS2
VhQ1RAk3NYczdFTVvSnPxer13nZDSf9WuE/3kdz33B87/wBgUCnoJE3Qh3+umN/A
5NHXmpQkc0fVoToGgl0DwqYLiHZ1N758f7nAI2OwlAN9lvC50W4teoP3mluueRdt
tr4SUum6lTuc6I1NVNzlDOcVJCp3G+M1L4//4GJFpn9IJQzWNx5jlzjtk+1oWuib
EZxI569lBU6DBaOFu13P85zHNkLwk49htFeNRCiyVuFyukaVlYE5/x/vpQdCL/ef
n/1mr90NhU44cCYAz4uMgyZ7OZnTa05oxNURPMGcx5hJ1l0+oE6NW1KRVZna3QFs
c+1M0MbsD4+HubQobe25Qe2TXbwv4r+mylBiMkyFLt7JFVe4oDQhgQoG3QFHfKcX
ySDirzodztA0PIMBvqawxaGcIS/1Y4m8Tv2copaZOSvCLseJVu5OtJys3EvrVHFN
`protect END_PROTECTED
