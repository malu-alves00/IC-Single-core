`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mE83n67pAkIEz6DoLRjMrwvaPrghhFglLYyQB5PCx4mzbRdx5QgCDti0odTwPws+
b6nPdX5CbF7Tcp/CwboaR1hQsQtlN1AdmS5yRJGziXjyj5t3QeliCMMn4NxeUshe
qwLqS9DrY3HCqHMKgHYlx7bXbWnXKNXhrGAxrIQiaiCGIqYzzM2vmcm/5jYRHugg
AqbsVlwcFe3KVb+hZ/xRuFB445cfr11XU4uWWeBH8FrOIFUoXA2NX5BkfAIQhEyr
rJGoCL5BZ4siUI5qnv6NZhSayVx+F2G2PSnIJSr2xMlfc0v1GRHyNOtuF8+v49Ls
+Yh6VtNuzJjHFa8zKbgVosaLYU2tSLjLupWq6wJKr4JmuciX/KFbX8qCBD/XcMC/
FgR0rU9Md+3yPwo1qsWPoIgSJdBl24NzagF7p8MovkYBmW7epciycwcxRGJvkLQ5
G4S6gPIXIYrOT+gNYHUKv1L69gU+p9MwsiAHtaIZa1k=
`protect END_PROTECTED
