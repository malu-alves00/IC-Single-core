`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aAllIyK2yB57KP9oMLtpAcBAL6Vy2MboZwSAj/smxfAY98vmcLsztDHGIkyw0kFh
S4/Fuw7ggOCgadF00CEGZ8JlePK0Jks29BahgEk0Xt0Ub5bGiDvhm+F23iWlTdK5
xm8464uTtSwhKGl5A6+zOVL9w4YwE1mKEmGuHVW8mirakGkA61VAun0U7u1qqyYg
FbrSf2ecx8gOl964ikOi5QAjH4TrEphDejh92xeTtA0537JytCGArjo/8IOADd8X
ZzWr7H7SfZIKkrMtq5rX6Jun7oWrx5dq6WNCCEkv2f5HeZ+x+1RVeCrFEZCRzlXX
OBR1rxlo5SEzCv3uHtXfyrz8XSyJsB+UG2XkJPjnsaz9KZQhnzw9e+4xOUo26Hio
bO9ygBFAwrSZJuTMRJd1/PBVEB3HJq0cD7/6YchLLzM2sWKqdvWEtXl7/gVvca0p
Ex92Nt416OcpotL9DoJCV/EGqN7PKNzZeHzPd3EmeLiTmySkMnrAOsfYiJW+5/2w
QcWm5p2v2qabHTgK9NsBeJLT5IcGmY+wQtv+jM0pvmjTNr8+yotCdg9j3KVrect7
iaTQMkFrBp15J8R82TB3KOf8ADhtXRYIV9MhP0+HtXkhMtWYxQDeoYnfxH1ovxLn
Ex77SqdG3+K1PMieFdRdtMNSEzSs5se3lLaSUMlkQ3ee28YqDoSH0dM+gvV8zdQh
ZWA3cn4vD/kpk1tuQl8VNB2VMZptfrrKfNDkUo+oUaQu4VMsYo3xKVMF/QXkWta/
UZ0zx+AOwVonp4IUdMUA4a63smEeiF0fomRsu0uapIhTuTZBiRxVPo5syQ1J1lkE
Bou3RbxV4wpGVNfgFKjbxxwFCdhCOx6aBfjG/A0Wya2QrH4EotJEHDEf0eEi1nhh
KGkBp9rE0Z4fN12c1TIGyLZVF1jOVa5vduNDZvYyjKqJbvVvpKied0nwYU7TW2P3
XFIkUs2cYRyj9X5dMFJ3wFX01G3f7PF04hcnpaQNzaTmmkJxmTT6Qn2Ccb25+rRo
IQ2YlpATwdIfdvOerJB4CM8qwQv+Xkh6l21HSyYrCSJkA18qxhPICh/o0xlbfO8z
Q8VJBrzNGeU0L+q7d0vwg28x0uvLgln5LSh3Ip0+20mZVBc9yYlvCWREPdtMfest
NAuNpPDLModTQDp6HJLzn+Y99R62ylN827YKt4ydkf+UknpKJQmUHqB58T9T3S/d
OWYOq6IC6gQ6ygar7HaF5lA+pA5FGZGoP3nOdFmgRPu9C/vuQfTNrK/5OlcvEgQ2
sxEGy3nh5362DFCP4+3M/Z81DKIz7mD7uIwfE9OA2Q9vTvYpU8T4QoqadcQHLOcH
On6iGwxIjXFgU51+mQo0Av1Xc6Tj22pc5ilFic/yB0MWrbLpsd0zrvL995Txt3LO
HNHQ2UJCbd/L8IOQuXHmv0IF97sYwR5Pbo+13Kc636F3Mr3SmNOiCvHxPR6zjeVf
caLyCYFZdGWtWkizBaXskYdxdAcqz+a6bV3mClrqyBE9t1k9UXBiyUkc1bkmAUXc
B1xXzT9ubjfq9fxWZoOBY+c4JJunJrBPmHv/dXgXxg8uTvRFHbIXw9UNW35m/aRa
D6ree+f/rmcfe88lvjS2AXzoPolWvw8FTGz3AYHbcYJQhusIa+SPVqk0NTToGlS/
GWqyYd+JjVibLAZmEPvW60G1VfoRFrCEk4xieXCYWKTPeCowcLXCsL352dJOpc7E
WY/IBZyrZ779giPO8GhxvYfftoPUUT9eli/32Quo0kncFLmL10D0QUOq3bnzaXtt
/xSWCdTcgmy2P5K0bMvvNe9mN72IeZy9nFWOYOUZPEaydhaskR9DkxzEGQv/icyu
u9Bg1R4FDUxTs5PXo1HQQCjOI8YGuVtlfXCAtVolDQgDJjHGTvpHBNOibx2Vlko/
cX116TgwrWwZfPzYVpOHALd8+eeAXp87dnpV82M7M+rIFO4EOAttXxOVfAJr1DTP
+3/y3c41gO/ZaN6fZrr+a88JrqE6HJ4OLdUMI5ULFdMn0p7Vvg7xc+6X56LZC5lz
rWTwg4wwAX3z73Tvf/5/XQ24i5A69Yu48G2c1X801Q5idDPsGuI93nPqexXTgjrJ
xfYwf/3rYqDoWNHcN8EG8nSw2Y1iaOyuZX0zsZQCySsdEavFLj0b6rUtPna8Mwt1
g1vsaWmduMKc4seP9zWolgmvcifsTzG7JHvm0DkGYer741jcNxt8Syn7ulpRIddd
IbEu/6qyBTGMPieSRPIhDFmeLIaSTr3LTvmRIhAPormGMWl5G7k5nP7NALe9nF3z
LfnA5tIzUMFKC66h4o2/KFKEWLMUatqtaf523l/Wn9PGVk77N+CVWPTOhSfR09wR
hoc/i4gw1hE+ICBHJbrEjGIh3HFuzobAxu4IMTdoN0dIc0LFewGx9LYT1TyMHfrR
VylOSRwXYcGGBfwnVkZRTH3dmdJAB/6Ji8+MaQnYsv9MDuamzNL01EXlm8gc9k1Q
XGWpnjG4nux8c396MX3JAhsCcP8vZ4key1gc70Wym26xoZLxQ04KIs4VPxKkdRIL
JnTNG38HsFF2R9tFWnyGIMeZZugK/3osjB4X5JmjYY07JRRyuJHeGktu9bH6CACC
Q+w02Ev0jYAWaExFTdltn7Bt//B9Ljk8OvPpmKGFObW4D1GxEUKiQDbLTnlKcgk8
5zUPDLNiEdzuTPXqg6IsBx/el9qyYT/sWLl7WGWiTloWXos5jmLLlUaUAH/Kl/nL
cSzFJtQG8r0h97ZHcZITi4rO50t6sQ0UD8/cSuVVCb3Z4ZKChXkGGz00NwfGLCLP
evinmxoby6nGDHoXbe7jJ8HrriUvSSglIlreWSgXSmRqnuiJq42XeO/i8lW+46Av
j0MXwnyufzkHPfWVWCsG/Ud4t6sZZuujQ7voqwt/oSoP/BQeKtqwHCsg2MlcZ7A+
mTCTIPX4U6uFpzPdvCrOHAfowqFeEuhiFahtI/pc9A+Jal+8CwQCOQpPeYwGSBtk
lQqYnAPt2GcglnhHd6nGSZNayIW45C3enH/Rm0v6BORPCxoPiBlhv+bJQ94wxh4o
MFHe4w3KyOUt4cd1yzsuG9R+EA4eHbeCydkkzGi7ZFOhtYnoXPUSVGf9UxknZSA2
IzEAspMNp9oOBg1H1myucKXq7GtMcLNBQr0XCSwf3w1EQ6Oj5EQwmVkINWGkdqWH
uCeFV4Yh5vasyLnz9WdVZMJA4WgGF3VfhaFFBj2ZejNofT+N6d7wN/TQsTbDYUBO
s2S3hbNAEtvUT8Qxp6bUFRxZRtx5juYqzzOpQIKE2wgHSIhA/ySSzxSw0paJzxn1
ZNujQdX4En7n4GxpA49dEK5/X2jORgwHO1hN0r2PQ0HvkWrq/LmdPiJi2qfwKha9
wg8SlEkAQpet1rqDskHE5Y9p60IocNOv50j654DirGRkpiwCdXBVGWlUcHfrBzvP
/U0wNfuPkAD4T727byUVBbst96O64wOkTo9M68upI9VNaqiE7PZ57GeqZbsjA4JD
o85yxl0hE3EV+nI3/Dq7VdJmqIXKGiPYRnTaPSqiPORJPm30XjVYBS5jZQq0LaV5
gTTtZwZf/JbJUpU9YBVZc1HcPdhoH2cN0dmHwzU1xUkdwelK4uygb/OXCWBjWWIk
ifLMFZwczyVZSSgsqzzrfArbUQNoiJd8QSnWefiiSGUliFRkke9tCS2goFk0/daX
CW3MxaDiIpTFaRUcCxDIKk4wSrYKQcZlLhAILEfEoEhx0z+ThHRakHVuDPWsiY1A
JZbqznrLxax3SMOXIL2KSrdiZ1zNndLhuRVkkfta0wJJ1T9+LXUmAMdtLqmyVYm/
lo1/s8CMFWRtDTnTN09vhU3ZRtT5gj0YEZOSYQ19LvA2i/UNtidxizhfhXSoH+LK
kxBYgpPBE+7Qzj3bcUMpTi4+Jcnl/+1mF0bwj6cvWQqAhqrrx1I3a4kzcx9JN0BN
caSh65xhHQvLqhbSCkg3zY8DlxEmYaMC+dhkxoOLUo5N6cxR3conWqlBxLehdqhS
AvIGbiH16UZMvrKAoNUp5A2SITBDs864cawfW4mEqm2AcsS9/5V/2pgepN/KKciK
A5GW8ZYwbfFeeBFGD4iNW5ifJcfIqfxNtf95cGo92MLzRSr7twJ8l3Ja5m9OZuo3
YsVwMmKa9fkSJG1U09Mb3B6s2i8rlNOJqHNjbKa9HfCywRP9hxXPnA9qC+6K0oNO
0eqgm+GfBYLNBw/swNE/C6Dd/uvl9U95MuTIpCNbGiZwf6h/DSSBCfAQxGb3vKDV
4sEIxg0IGpZo6N5RElYldDEq28aHDNEXqhAWt+iJCKDBq1QsvD15IARBkwcF0KtI
YB1qy9uvoUzOs5si2fkfaUNgxi0i0Kl7vjDZNqrzVQA2HejSI7qmoZPCQj91nmRv
QzdbIpUaFzwlL7jInL+qHRwYHIvkj5y25/GjNpVm06dSpE8oBefop8a45Q8BUXlP
9B5OOp3Vtemgm2QppOIjnoR1kLYV3pnlrBEHS3JbCivU1SrBlANbDLzeCH9+51Dy
ZdtfnCBjTNULPBRyDLpB9Bn/BmXZU6GD0eiSZkdDq6xtCj3pAPy2OieDAUHad7L8
hrWQHBs2I2Rzi1/muB/UqxoTprbbIjXLTLy48AKYYHLd5YOJCPRd0ju7F2CICL3H
Ul8IoW3+AQ/20ttN1UARqW/T4Tzh4YQW4JmJceLFabK+Zvyj1WyQ9MagDyzvi7B7
ATXdcjJlx6QCKUo6mcpQCEMS4hyinfsELNlXZptCfgyCPFdAP6UvBKCgmdLQWklu
u0e2gAYLm3+FWAmTNpR/lLW+i8hg7PvhYf+tn/5M0jahMZFi4ykxS3TLZJjQKoSv
elp+9JEllFphiYmYEuyygqqgj7WXaOSeoLCa4KfKKk4uXJKw8mVTolcZZRn9HU9D
`protect END_PROTECTED
