`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+j7cefWexBIVWouKiAW+Rw/NE6Gwq9FkU2+cXgeRY0ri0SLQS0eMJuEIoZZDOWKk
TTMGAJbMYd70pgVN5IZpiZs5SgYKZs1TiO6IqNc0kmt8hSHpXqmPzGOdNZTXHd3h
O7pvlidIp1IVGYILKeo+bSP5gwslAHyyx153M71yfzTBhqN9c0XxBqdAa0ST/X27
b1lHBua8haEhpT4RJITf5uyIPctf5TX/dXSKvRzK7h9tC0zRbMVw32tkbA+PzSbQ
MCnFgguyHkI7jAWMGDddiDD31d8Xbp/4koOrjZ2sLojAyN4HrX2fb5Vn/Gwrgifj
D/zQaiCSgqpFO4YSlRZx9pIVvi9yRo+26WNwPT3sjtCz80oTuV+X5zsBmrFyKp0q
L32+lzpk1BahMcKk8f8bwCIb9aoG1tZeerbSElpci2fDG2Y9CpKixZoS066DT8jY
zubmZU7leKHj7YzOVSKWQwEf1e5CyTRXhajvd6RJh9TOTc+OrYejBMevGCQpvNPz
dqBw1sZPrdCc7oKzcggaK2LAiF/FpPAEuAUloZHtsi8Qbq7Q4zsB3D/z4s8lwHZZ
HPBUked+OybQa6s4JYwoC+p88lBzpqNvqb9geswwT7ymxYc4wh6AnPOiXYrXKkmz
b2iGeQx2qP6kbMX9a4f/SIcKsrAR1GX11Wo5Dp8oiwFjmNlUluhP/nBedA+7/4AX
z1K0yd88/iCcWRug8M868iVY27EH0ZtlYJgysvsyjNg/OX1bYu29/NkrbDbNfD6N
goOwyqxsAHDZ7fG7N4NoYmzA1wBpZyW0mwscNw+/FYvnei5AxVKaEZtEFgMwHCQa
VkjVU07d8hU+JOMflf2+y29uUlLYM4yh1sjBhGvnQZX+E6HYnwbcEazzotJYFVyA
khSOJKc1Mtq1fmgVV5MHbQhem7Yb9YE21IUbuYOv8eL4b8xgmEcymPHHsUbMx2/z
zEDPWWsa/2WfiletfF7NrP91JILgV4WByYJ0JPf7uMw3PbWmW1vezmbHmapYB+gT
6PZGcWEAH02RmOy6u6NGrtyBgtsnSVGwB+WHWfrO/UhdqOF3fmsBFdBppqvgFynW
zO6NmERJh3KakYh7eVnzgO/Mpyj3tTjBDJCxtB0SKARo5WF5aJpk2o7lljfWSy6T
fddpWGhycFX1o4kURbnlpnTRXlRE4o+4j5lapsdslUiOBJHNDJY8CoyXSAo2wDoh
OvqGbNsIj3tAu8fX8mddUkFptsEpnf2mZtF1yNMmGz30szZMAVzvw4WqWNSfPkbI
1b55PykRzQEOpPbn/6Dg2arN7+exvIyVEYS+D3oVf1WbyqJFtcB5jZ0/yNL2pwou
s/cDz8IQB2D11G3HNOASXZ9TyveIHCdzghVk8EJlotKHUqa8geBQNeHVpuPWM9Jk
GGbHkxI3JQQk06LjwYujy9dhlSLiVDo8gXm2MiAG3sVPrsLGYO0u0/rORMDbldOY
7Y8UeDtiuS5YlNAXQcmOBHMrYLKDQrydFG09GPK4itG1MKliWQORJE7SsESYHjr0
JIinxZMZahAF4IxsM19vQxVyzad44ytS8U2IHy9ieYOnPsJ/wxd08J5w5flgsJzD
veaOchritwWuWws2nmu1i3RGfzzSl7XPtyZgz335OW9hModJB0hF0sZ1JtBRj4MF
byMoRMdURcZkTyu5ZSeXx3nP4FHpiZ8PNWOraC28zYusbe3HyXy5QKClhPNHEOul
LvMc7UGWDMjplnZDUuAjujyciWtjeapBJxHxlTPgMn0mn7z7fObr7++M3jPp6zEw
u07oRX7qjzEDVNZwMxzhG4nt3YHNnaKVPiDRZPRvMe8+38Da86wMcokbxSQGzEon
5t8YpQI8tzlLVojsjM/m0WAjrA2juiG14BAamY8DnNCChfMPzkYJMFx+NrKuZHKQ
bEfrcJxmtU7u8n+EXYa4NEPzky42IcDERjtmRLcKOFRfZX+nHDv8z1QqDZfq3rQ5
AOqKpz9NfAhYREfkOpmwz1Uf0V9kXejltfEc02noHMsockI5OgtH5iksM9WmhNwc
e9WlsHvZU9M9kgcAAz+RX5zNIu/QgLvgcvje2BkvdfBv7B+mgPpiJ30aOn38z0rG
wmBNLp9IUYG/tVp8zUu4AUr0hYmbEMHqoHeRHw449DM8oNHXXGDSBAt1tGFVnCvc
zo27bs6OqIG42iekWCBVvKJ+JMPBtxNFMZ9VTPghPfdg6ej/EpeQjdaGKaIxowic
4L8GJsow3yhXGyWOrENp+gywB5vW2+JsA1R3cAIM+YefvZuRJoaY+dsyIWreIPol
owXFvu4UYNjda5Mbff8+QDZQiL0KszcgUDpv0Gs8EEBvWV7p5oGQjPKwqIcrt5mt
sGDJ528SSAgOMJzsNyvbdvfjIp9CzMaCOB8TMgkLj4HwGFeCnFeQjVc74rNGoeWI
yqFgsCvN20jd8N8lxmcR3VCzjtvRVye3mqH68Zqljt3lpnfEXB/Fqn6H8UQ7hGHN
NZLo2MNn8YvAdPcThH34mDu5jEff3d4z47d02Xx95G+Z5EKp47+K2yP4n57xtPk4
pWFfmcZc0yEZhq51G4GxlVOGP6SjZ1yfc8ZtWNNbfVBl00koz1Y1RPllvykrPwNy
ZPRZ4VxyanouNk2FrOOEzo3RkKDVTClrI8APylhVuquHB/YDuzYj7g2DLiCkH3gk
COc9evp1i/UGhkd/CnkIiYClnyieyFaKLvf/Ci3axt7GFXYgjxZmduT1Z2YqywTu
2RPZ8ywqMEC2HSw/QAL9Suxkyq0s18xqLaCgNz635Te5HWimANJfpiuPI5ecY9SC
SL8J7U5RghzmCFZjyfK1pQcrh/sz7jwtR82F1JeuHogDt8XISWhwr+DD7iaCuvM9
Zfotsi0261SY86CwKPsfueNsG615hsoQ4/E54z0VmNurf8KoVmYzbyUX+rraob6J
5BZQfuSm2eRUw/gMeaSxOtO6oLC1yeDzr1e1GmbGTroAZaWgaaJ3fGcCY3zqu079
KWii1RyuxcozALeIcixTYNbyIu0vFrHZ/gx/mbfNaMbSOPYfHW8fbnzxkTXy9IEd
BzlCxv6dx4i7ZdpjymqyEW4ldNj/dvu8tbWRgmLTCdoYFFKmbmO59AsMLuHzcklc
eZ/6CULUL6yoT+8CshugvK4m7yflGfX8v8c5DzjbvwcvC+eHyS2Dtmn7m6TfjHSX
4LeTka9MaR8NDg2mGA1spoa3BCsb710VJvbbDLYaz/rX3F7MLXZBbo1xdo4hg7fq
r4ZRGSeoTrIPUDSZtWWOcs0595r6Tsn/w9JfwsXDptvSZqduBX2RNFbytwk4FtIF
mlIoZznpV/M111kDGuf3kjzDIbJzo1shE0zewnxA42QrUe3B8SicyYnzIc/rG/9F
uy+IWQx1V4kYJAOKMQaTJ2UYOKsU/0rrXCzAMb6FK6wBUDI7u214xdOT+ypcixea
1672iN/rEbXGwUmkRMT7ZlNNQ0kwlyOH1+P/fNyj/urX4YnUf7HXZxcTyXU3aCy9
/90C+ecvx8m2UgaHF+ma1hYHOPXAXvvQwMwJCqBgPGJHNu11BejzuDWz/BPeJDAS
bX8DqTnV9yB78TQdLE1mttGNd22FKt4pz0DIK0pToz3sx01daHrKmKfv948kfev6
UeNXP7Rm19iyi3l+rAGEhxAyB0prTlp/GWxYyC1k0kUM7F43o1OGzG6z3CItY3KB
XQtwig8NSHtE9pVUlFYQPMx/Y2e+JTKGpF+3fljpoTeaXZ1fpQheWppAqU5sX+LL
shhnvd2qt0Tw3UX14ME88FjyQRGwutIf6nXKvKtk99hQzQJzZKnujyl1+ILv3uDw
0uX7i6d66YclfclZWaGX+ritXrvXGOnWqvRBVuVoiHZG8pJM4VRrdbh94lAo48dg
rSUNlOn0P0Rb+8Vzt61DozxghSoRozS74wTwx4snMo3xhDMw73pva0hoVN/h5oCm
`protect END_PROTECTED
