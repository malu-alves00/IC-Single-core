`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7fDoMgOqkXDbiaUeza/xMaIHiPpBeWPJF1WwLQ31GDQcAijN46GmS2VhiH0iHgIq
ZkOhQQT5FT3drMt4W9vzHJ47AB9A+XUbe6DbiUBM7PWjsnkCOPp//Iu+i6lD9nLS
OW0FCSwg7p9XADrh6gqvvWqi+sERWTqjz6muUN+m760n8agRvDXPWQ7sUUriiE+c
5+Ezf4JIxxNCfCXARKgmGUptrsYBF7eg4K0VyjpR347O9R05guH/rYSP6J+4m2VR
2kgZZjFlrdXkGosvSuPIoFveb1mequxxasdXor/oMeq/p+e2H5jd9bxCFeKrEQNg
EoIiuyJ92IIf1cZO+qNPFm6Pg2gRsFAf9Ry7+ewgsW7JzbXX4FCnuFXKmEcqYgtd
W2IdYRK/n0QnIN31KIabbAcs82Uw4Ka3tTQLG0HZNsrx+KJDMOvFrn/5ZgSjdQWK
RO+EThvP4bHT7AKjfY5jN0cSsVfUWemvjU4je5JxVXic1V/pP97Ns96r2+4JuMKz
viHM4QSDBNNqSn/d2E+vIVteYo+jrdf8rivF6u2kjrwU6K89lcMaIup1ZFDZuOv4
TtDU8tMguHhqRZtT41FwJxGBFHTBH5dIjlSffAICPgwozu0klvyK2Im+u+3RIv4S
og8/wcL6RbK4+ALdizIJbf3NzI2ZPbAMfUjik6Uq1m0xKt1h9W0zboz+CQ0ABOYU
YtrgK2eIJ/uFcJlHC3SGvTfnf7hclP2kknzTQ/LyCbmttqWgh1vWsDHvGc9BbsL2
mq1YuIwnkVxs3RUxIfnuoKctyofpOdA6B0s1iw73tkSYUUFg+jxmLwluOz8fumUz
Uay6Da0LIFnxENcmrPyy9x/w6J5YM0qdSrOiEPDce3geh7MrYupZJE8NwkyPcpGu
x1aplgg1O2CazmMZo2U9vCU41fNW39DdetWjHcn01zXex3oeL0bsIa4L6ZZFEhdB
3vc5EvPLfSa3yG7XHXRBvcMzp6xvVy9mNndTkrSDvI8K3ySccyR+0f3MQHDU9uJJ
C6sg/LmeQDWsWx2gDPsIT+jbfH0nabJG5XfTxpOZ/zpRhRmwEIqgYgeZMvg0e8lg
25Cf8pO0XREwk2km/sG+gVKJrWwv3uFlzJf+mw6rl/cQp4jwujOqqKuOqAGZpnTP
QNOuAZXtv5TEZQN/3TRRnm5HhZyNa9iZLRnjbTpI/gvS5+5UbUA9wEmmVHDjzdFs
EzIjOKuwVHBL2JPVRWablPZ3ItZHLUuwE+BDmD9d4nbyW9gVFtOdHDN5ActoSqnI
51dHcmEDiyvoMxuKuNapKdF9iVkKZysoQVuosm3lpC225RJ5mB1BVDaQfymF09zs
WilOSGkGXX5bRl9PovR0dXhrnXkB7FDv4162puo8fNK1kf0BqGqdvXcQR8PpdcaG
8Z0+ni2xjA/LUKK0bcBWpj2jcQVvf5NqfavvBrZNaMFqNNLNqUjRSh5zjn1Euczj
Ggi9hd2yMFSEOWd4oqglg6CwzweR+6s2Fzedmu3gnuY7JmA/8w4kD+5Yfb+YnUfC
HfqKu41TjLlVYssVup5jcJMGvxqKJ7cI9frPBbQkvz50JHg1xlRzH2NrnSLlFibQ
jytptkqygHgdEWnbj6pRnIxPra+5pkXOIFJVI0BHDuLl4kjgscOF1uLdRAenEDzs
qX7ytQtUCN9thHScjZKnd0KozVEe9LJ6/p53ZwGlfoutzhpcrH+40zI/pz0anIH7
oc71NHjgIZiS2wwU/j4YizNhXvK1+eYI2cfscu4u1PahIYiAWzXefWDL1/zYKMhx
DFOtyRlf/9nhSEl6H0CMQhZ9TIo/8ZNtAyItXUzz+H97Gsyj2U8jO70W2Um/XXzP
XygHz0Os9JaEKoT8MDQJUKu2EG7K3LTFs47nbiqwj5JVik5o9j8YNF+Op/aXge+D
pNh/kjhLZAVTNL8SzUKfU3r3kaixlorijICNPs6doIt0iA5o9kcfP7kTpWTD5fuT
aYLrhkcILLZiEHhIPIfnUcmECafefyDa+e2KZlA3SoUloRAGDRRnEhTXTcKlCHUU
gpPakgH+pDnLbaGGkiZ+b0OBYIgPSFy9N8Fes54hTbQ5ULg+Y1K2YlJcAVJ7NtnN
l0saIPPui5a7W2rP2VSxQbMkal6VRNCkdBGto2wiSKWVQvI/zi2JqnkaAk0y+6Z/
uDhKSNrbtvFKUZL+0GVYOV1wcKFnZqXwtmV0VepDYiFk5yP6qwno55wyYDJ6AksO
QtSrMu6m8p8LiOoKGuHxitGj9uzj9r/PDEjKLR+Ajo1fZB98/2EpdlAXKW6eUYIi
RLARd8pAQrBK7PmsK8HQEzTLFPEbqoh9SK9lezjTktQUjknqiF2+OVxnNerW6oAa
YarNJk5PDRQ/LlIY/sl6hAzcUhMzt8HUKuXe3Zdv8PXFTIS6XryOBcjvWwKA32dn
tdKG4Z6/Us21qv9qwmzIckwmB5nZZrMaQmEx3pBRgmIdELJsK87k/ppuRSMzgDIT
QleRpm5TdWcs20djSqRamaQX7tjMC9LwukOojaYCOlJ7ad1OcKl/jHA3FzF9lsqk
cQNs1WKFx9/dhZuQ4CDfiyh4bZSv8gSVY23uLZFwZQft7Ox5VwZXuoRrHQztNtAT
P7ZwR3XPeN6g3uMPH0XQmldRU9Z/X63aiHsfIRsiM0eXxVaWzQqgwtF56HBdQ4iV
l8XU+DY8j+dNcX9Rt84e0LVgY96xMXpHf4tWFpzm8yRF29ohX67wz8H7NeIKhVEo
V6gpvhEy+mz4MJUyPsstJnyAECgHKPG1BPrnQXgCyNoICbzPqieVYMrGDmhxfsnT
91uMfM6USJbjjChvaeuvFLvCG9YlOq8esZOXqMrukz7el+dzW9zarub8jQJTGg0m
+mKU6oDAEFr7370S3+j7G8e0i/WhAOnUHJk+/MEvX8m1Iivj2TyrafH/57BPHPkB
Kw9nXUlVzVLI5LjDisZEt/3fDw5u+Nr/wg9ZbZGg19RrOvwX5NOZsTWXVkpBT0CY
rNZiOOVXM/fd7j9x9Q2mjy7jOeJlkeGe07Zbs6+OBpllqP7NjD0Da0bIE/2XgPgr
xubftlbmwaXJLjYmlclbLUPnVzMwxXhw+rp+3t1iz+Dzp8fYCaWrH6Wfyl1GMqF/
Vo2YxFaEhy4wQ62bHIF5AotQeWGveYvV4w2tCJiVBSyEy3ZoMY4eQZaw4EYvvURh
uKTz0TfLEdWJDx0uRbXexaVbiUnpZx4o/XuO7VPZDjqeOiSQiqxFewZVkw+zFnFj
Cl6A9QqukDCHgCRGCOXBxkkHzVEJ6LuXLC5R57oeybWI67t9KQuMFV2bECKYnqsV
L97wOB5wOqGGHB77cG3kjd6Air/pgpM9Lw275McJbfG8s+aF1KxGtKLPvsUvwkM4
b1YS0E1hzgnNtEtGnudPvt1Tq3uqq57PZmlKeqkMeTUioZGs2SLt9mCgMW4w4iZ/
k/6kydEiaATMqMC++4+XmTDvXSImLaCMxAnwcJc3nu5cS7wu0QKZoiXqQr1a1M80
u3RgRRi5fAMoQKi+mX1yyn2/7GC86uRkMek6uDti/WsCVvgl1LqZ6b374XiMDgNl
r0xi03ngOCF+Dfhx3YB38ez2NbIT5ldO/vnA5GU0+a/jyejKOpVFaOVPNVjcqebv
DmAvkxkK8VzHfB3RnfE3hS/CYftIDwcKbfZjCFsFkqpT31E0BMFQj5imC6B0mETT
V4df5cmugGdHw0tAKJ4L7pNhlmynWIa/jOuP2d2vBW7WuvLbHPH06VFYYU97Rzj4
ffTXdav7xQzm3KxNbqsmYMFQtuJm6a3vTCf6C7H/TcsgZwkqeHsFlv9H2yEXvkEw
FCfbZxEQ4aw0Iykhb2ukMrM486gBThlJfgK0TiMJj7mzLv+Xc2eRU9xm15/ON1Mq
EV4FV+mVORXFYXSkKWmmR2TrnjLVzQMM0nB78zYUwrxN14jPyofl2+FGmDn7lEau
Nl2OxtFb2qbUFNk5L2BZvLtUYuPkaNfRPUCXQp0Xj6pjD+fceE+RyfCvyThf6c7g
1gRXCCLqGDxRICftJ2fT0oOyqKA9Ecy2og+DlFkSkd2ol8B67DLLheMeQc54nhI5
ThDa0aV6NG64ld4xz/+b6RR6DHpRxlUZRNPeCpslhQjDoP+3fEn4ixKkB2p8pppp
xJaYI76AR7/Mnm72C/lF34KgRgq3QmkqyoTfkCNR4VxGCus9IjpsJGYJ36cBmvew
atIZPAlN2erkk3CUNDbi00OC+1qpERvwKM+4z3sKEJOuK8dpojLn9bTEacr+n4fa
M4/KsvsRVql6lguodgf77ql4Cr4Znsfk3mSgqDGEVlYlJ/O9Pbj32gWVeWZbw3yY
RD6OfndVSrAdIGsYi/6Npl7j71xDR70zK01FTS2n4YR1PfLfn8W5pB4Mbj8Lj7fY
sz4KaBNsJ7WrVsRKSDgA2hxngJ/yg4xwSvM4V1t1HdERc6GxyDa7+V3p1kO0Ueec
SNgjoLhwVXDW3CMKre7Dgr1NqN11RA9nmp1Fxa8tjWGgxqYJqlZVXmYybk9s6di8
aaYIGkzxxTQ2gwqh/ckGp8o2KSLQ8GffAYziREtecP5P/42CkiLEu7fBkesu/oRa
HLONWXv0GUHP9HCXjWt8kJXmrp/J9uaDJWAg0wwI/7NdDBf4hE1igEETxjb6Bh4j
JrSetTM8X3KwUjiUm6R9fMyYDlhlrEB9T7Jp+n/xq5PgiWiIj7Kg+69LJ78rFWxm
4hA1KmsWCelD2buwYDwGyqsycEVj+ATqjXYJ/5duSlnmGtpX9FtLkS9ZUSFnRlHo
I/hy68L8UTJigqTasVcu5xpc6bimxWArceHPPFiQ65YumdGnEUwRyfWR4hn1JWZr
O+FBhKyAg7FSX/P+6FyDKPEUvl+w3Yeea51rMJ7b3+Cq9PaoCFgLqGFNgwMcv2EH
5zfDAI2FcusBbompztinPQ6bLsANkUJ08N/8xlSKqB6PHlBS+H6smDXUSjsgGgIP
F4+CMGQFU+Q4x93W4SCEex2og0U7fW+AeEm+e6HwKmIl3382dONvwCCGDOxHdyT5
ZfitzrHWg0ok9XntTp8mSP9KcES1niOkE4TeU/wHNoS3SZqQH+GWGt9fb/OzNR1q
M8vHaoyXprmMKMcT/doU2irlwOSjTXaneOMvoqRDyc1z02+M7keEP/qCTiApUkCt
H3mGSL9+vRdKl4nqybgQmeCngO0NZ7qzr1cVx0bw+IhUYRobIvm7o8oKDMOjiVIO
u6bRfZYvLXl2ZZfe5vbqnNxA6LZ4JngBTV5rijsPaeDtw3G0f4x8IkCCyjbKlwtO
S853HCbKCdY6uSK7pvwg+DbNjlYYkrQr0yW1nhU8Jm1dUmA4m+O7XH02SKdl1ejw
I5PDT5F0C0VsJna54IuMF7kM/KKPRllzfg95Ji7Yc9Z72UMPnJ8DNqsNS/UdYqm8
wd8Yu+0LYwZkSqb6Tw8HviflBXyuD7zJbWd4ePMc58FHYi02gAJRAT9lmUJ6tsV8
4WkCz1C1zWgo1MIAX1pVvU1tILHBVEGSzP9nLRwcETWGLzrBVqtayya2g17hn17o
qGswjbMB9ceehW+c+itXQoAvHBTWSteIRwXm1Rw7FtXfxV2l8sdZsmxXvwPdGNuz
cnEcHwAgZnvWG7kKC6M2Q+YR6dpubNPJqN9pwN8MFhBuGLdxV3UP//nFcUsQq9ER
HOb1OMhWzgV6B96AeiCqlTncLp8M73cMfvKxPyR8mTdbNlzgjJ+9uWnY1wsYO+QZ
L08fyeJ6AUNGUycwCd8lLKy4fISt0rgMKZmOHchkKXDU1R/IOldiumP9XsQeVt0+
R5GsikPfp6ThtxW1Z65toojOcM64VIJ8rmwh7s7kNJCnTpkYHmiSSu5DZ6nB8vYK
kacuQ1wpNpAMoE0/qdWrllcsgGA3TYKVnLdsOnyeddTkDIPaWhMwfAENDGApucBS
AZwyYPRWUGAKP64JSDM6/HevXL4sWoXaFwhx4sqz0z+vdUNsgELAhK+pyR2Ld9Gv
UXgGS2NzcyNNxrPfMKzrxSuz5EasKRyKfcPEYs4X6og=
`protect END_PROTECTED
