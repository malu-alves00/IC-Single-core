`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/V1zotBLQDvv5IhH8omaWWZmzk2N5oQKUx3kv91vHCvwwlfji18wi+om/a0Nv8q7
J8kH4jf4Rbm1nFi97kaFapnWb+o3lU5VNGHtFfjECVbHRnmDtLOY7OeN0Ui9aoqr
fZGGSXY/9oN+ICWMSKkNJ3ZEt1YadjHtO8icTD1SJyrLGxCKbIVPtYz+8vWWB8os
57/uSmjCcy3Bu8hghyaJSEHrgUA0jghZ5S4F1Y4zZWB1umB1/OosJuVF0mWSV8nN
ZHqh+u2EhkHpUnozlCTHOVGJl1+AVXeImDeP7dZVLRK5Q2CDenRdYOAjb1F4OEUr
MjW+i/ehAoXYdTS29xJJNphr+tIEcIuJTIPZjSkw/vHXcFUhz0TCGqqVGBWnYoYJ
NG2EzAbZojj9BhdRRDuCQHkgFLSg6AHqWXYtU1XE400Kczk/8EY3RV8TRWyGUnFE
vcrr4OazyKeWGNKcxX2UauA644cEVfmnqEP5J7VIdOKwHchOF/G5KQPAQpD8dsqV
XG1ipdXkbb6CMDj2mO5DgqFpXs7p0ArxAoSvOFDMauR7p/fcbhgpmCQqI6eNVRS8
Kwgy4L3TR10l2ERgmIoa8KoHJ4Y6oOjFSfOac/V5Flrw5OJ3y2YbCxp8Zh6jNQic
kJTRsxk2y6P/TdOg/Wxctk5OUJ0SxYbgQoNFxVCJ2kLXacdCwgA+Ucft+BUDayOQ
9MMH6YTrY3GS3DlX8vW2PJZWHp3d4EZJKpttMO2MLUIOKrz0kuQayokDpVyBV0d5
oXUESfIOXNAusIUmWKZEO3XwMpivo1S5GXM1mLAGUIgJJZonRZiugo7c+UfazRN7
8tjuoTlXJBLXw3BArRbSq0EyefWmPaa4rlByA/6r68VDBfFsE7FQpHE2JSSLvT1T
pM+y9msm47Q9tAH/KoX+5Ko3gZV0g23OFL82nrz/meoWZg9ckncrThxkANoeq5xR
p6lI24VQHmAfVYKRazV8UV7EG/VHkyFl9fC26LHgdeuW/aMS7qBy1zx4qo1NQw1l
8ZER/JF86Re98DMCxJ12QQFZcjbsapUNN60Vb7JT3HEd6HqGFJbncLhr2fVOpldy
alzrI5QQldPrqjr792ETTC9muciR7iXxBBYf+W1bKHjDa8rgqBYedKiLhIxCHIJU
UAmYQA0d4k1yTmVyzISmF6maikUo7JNAUuVzvbHjtjqiPVTuMl/h4rme9dsujpYS
2Lf3yPWcCFZR/t3BMFNr+x7BieYnxV1CAe7yGP4CnLlZikV8hoOlSt4fy55M4YrK
4Id8CDltYeWPACURGcT1GVidXXrgLX73IDxHgHhAecscyZB+VWZmH1jsGTPmPo0G
9O23+TPbY3/F51FAaRuT2u6kpQQ4ckZJxcbkqJekHB/as7ZyqkwGJT7+LyginjVd
8St9lqYTAJ64mp4HMeCR1ezbh4qdYXUdawUn5N78rKuL+Z19n5zkRnr9zEY2e0pw
`protect END_PROTECTED
