`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lPQBUg4+JOeBrg4OSq7HuPlmhMCkC65fk9joyarY2BquierxSeot82yP1m7poH1D
XVvvzQtWU/DVlhRB/ZazHLrjYWbVONORGBa7waqkbW89+F2xV1jVLGxrCcT8ChHc
Kk8BHlPXisuKD4uCZweMkaLQC5uPxb4Vc8ALw7R3fRFLa0d8CvlBNgEmYtogPmJi
MblfVCAu/vd94RYRrerQUz7szyHfkYkC1roYI7WtQuNSPrNcigvi+nlJQlqO+SMi
L0m5FNucIQ94L3ucy0SXCrStsH2Bmv+uD19smx8SYTVrqcYUdrNpSfZRvYms7eWF
wE9Pn6xwHIaGB8T5WDe7rMXcZaBHf8GXorWVy1CPRneDAUFvxl87ibvfe9xXqIBB
tPOlxIoZRN0Ht47sJaTJECfOsA5zYmL641r8Ud5+Iz21Eu2gJjsFXFiTCnOxRBE9
rFCxq0shgCOCG9h5cSA5E+3gs4syENlxlCYD4l6Px/H5DoPDyS8LaRZu5r6greqc
qMjSl+om9bLfBTeVEtpHQ3s1X4qeGAcRodfogrdUSUUkGmRyh0fUV+nxMo9RHlFg
p36RnNoSP7y+lL35We+OS4ZKYEuqlubqgHZzWQjw+NureWi6t6R10CEUtzGxeAwx
3G1aIxYjRfuQ/IiPjo4Ge+St78/rzpUXnUkXY9+hPbsemAGIfnQGopyUJ0mlnoiq
CTVJt427XH497x6U1MaanuMJLvO6ZvVCr1DRCQz2kiNo4/uB4EeO3w9FenArE9Xh
BBB5ZL4BiXy1pB9ruWYXwSC5XQC+Go+Ha6U8pU37dMPCPkuz2X0V+RVjwZE8qV90
PXur9E+51JUrYA2r2TW3ZWzMzD6l+Al4vuSquurcouT9dSE9h/ZHPzC1TLxeLuRe
v6QfCzBrJb+na0tI1ggLso091gqxAZS5+gKVFYJs6OOdc1VeJq4Wl6a20pKVkOen
QQArAqUrb9S02E6c0JEoQK+ZhfUfBeyh5WT+gq2WaF6zapyWHYljLKfEgAAO/5ZY
i9OM3sEr6E8erOi5M9l9XnoVcep2e+1YOjCq5fOJtRp93d3UyUDpV2siuMhodCCd
rNoM0T8hb8rSP0GA2Icohe0NUo+Cwib8v8bUCTbaV72kM04cNT3zWYmV8Q13mOUF
LNnxrjRcHcDSZDRDWeA3NB/lHQKpRLUP5H5dVE9hEnB9Nmn7NLikU8VXbGFNcuXp
vTF1teo7h00T24lmHkHsr8sgWyNynWmOffxVtZCF+zPEgAHhGFD+m2LCO1Z+CnIB
XnOjibiHlCT1g1WiNkiYGJHeYQSRRmOZmHx5bxRwvUfuPD/mqu5qbdqzWtozbNoY
ip6vxY9fzTWQhIWprS8BZs9wSGyTz8IoQ1HMZV2M85D0mHNw2K1Bf8jdg7B2YJ2m
EzMqAY0c5CoDde1jQeSsYmMhrtPX5iNO45If6QvBhVNZ1phT2Vyi3zPAZS3XefXn
X77CqYcSS6Gxpitb3WcneXcnfI+uDTIoGKxyot20rEFBby/3l6zrUn9jhlZYZSRX
UDXHs9h6kQDUqSlW9+19ibWc2HuCYTtcRFjRKsym5TBe3x3IEmTzQ1S2I//pU/bZ
iSf3x13OPh/EEeC97dHEcTbNkxdeaQKXbdqw6hSJm99fSWrLnIDbZwRhn9iwVpBc
fAsEGf3PRIuwmwhp3qds5CP6yCxTSFVEeo4luDmdz3LiPmfUEO2j86sh4m25DvDm
lDGUyYmdN72MEn/f7X/tdtB8rr2JhP1vXyE6LH3lETP3HHNybQOsG0ciOy7Ac5Sh
NhGINSj2G4yPGsoqwQ+lKmKrE+7Javv9aaQro9CPZfdYR2R5FljgjAOO3cTtGr8+
nlLNJd6odhGqGJUsKG1Gbxkaf+DZJN1iPqDKEXLFvobMrB39zi7Ihzp+syz/GY43
ArJl/FSdO61sJKQ/yrXDr/dHbgS9o5HBSM6xaxejvFk4SNkkR1lPUVNqKCuJnho8
qUn6BQQQELfitDyV90QpOCgVwExtjAm/e3R29nx0zjQvpDay2uihLxN5ski/B0en
dh8Q59O381yplv2XcR/sOXFHZHLKj2E3yZPuQ4/BNBzzIlNkoFIW8GbrqS4bf8s8
QOSSSPoUtY4Vbm6zY6cn5/WHfLAOuZcMZ6bU8JQFGk2z9DbCFIVoBs9xUeuGPDbE
gzGPYxIIHzy80FNWmxa4qX+6ZJHCMPopY4B9gFQeNhAqUWZcaz6WxYy8C9IvS6Vu
q+R4nsWve4spuilxkhyl9lZ2zCsKGPBSBiVaw6qUbW6ZwpEos54+YcAGq/l8QfHX
8BH0nPQurSdgVkStNyZ6rJkD1fwKXMbGwGUx7QdwA3mBTOsfqDyB8BjN172XbmbQ
X7ZWmPLqc+eXGzv4Abbrmnwf6vUjypvCm+aTdUve7SOxQWcKsZ3xS9PppCHJmhtM
6zf1yfx0dJjbP9rzeQLzDLxIJWDOPzUpFUHWRTUmwjHme6VQezNYJF+XnRmXYxse
WVc5OgNRNWeka+7orIwG5iZIpRCg0tlQfxr3T8XR7YoONsb5fbdVTb+pGP57mY4l
EUhRrACxbDukp1sCWla+e5sNi1jtYCdivI0YRaMxQqj/fzcK+trAkK2632Hb3zIv
OIjK9///E50KiQ8rIJ8AjawNr2osN93p44fEKzNIq7U6qFlHR/uK0IdAU0Q2EvSG
P7XxQWLBWdDlmZU/081weHJmnc9+9JylXPXOIc3nTO/x7c86LxOR3CMWZDVjTzlT
6KdsmtPHa9x99JpQAPzj49rbxVdSXsrxhXtw49PmQ8vsrqEtxDkzVP9qFyHnlU9T
yuHK03ec2sY+z5TPeJeo6icQMd1lyZDn/qwDJK2lPZyhg0u53T+vDTqCfBTldRwC
CIlkXmcegnlk96GvrPCOkzP0S0eD5+BphbCB8kzv7fagGAGTHXsZFbjCMjjobSkI
IK3ME2NCE0WxxYKX/vYJlczoYezOi9fU/ybV5Ad+6GIRykZydByA84q0xjtno+vM
yjbtdbTqkjYRcdlDEmy5UTJP9/Axh8kOrMBKQ8M9qawJQLzqtDcXwgRL/RQXkxWc
bw9rNYEhzwSjboxQfLRBOqmZhdtPZksvGAmbIv1Woi2kHdTGXd4cUm5E1RdLJ/Cc
S7W22Ko+6ST9/LqVsF5uc/CYmrSBw/L+/IvXwZfR3Cqrgz1kc2BvBLGsXsX8uV+O
ZXAZAnQdjjs3HVMsoZS9gUVteI0mFIJ56N7/3SDBweco/p0IWkoUwKBdh1qLq4Lp
gavbSC3OWa/LKf3KRZDA5g==
`protect END_PROTECTED
