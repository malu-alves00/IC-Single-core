`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dKIkynt4l3J/e1BWlrr4r0y5w65PT4R5DUVE1aFtOL3aB8Pl7I1HyD4Ie+AnGkVf
YXKULUrsB1orGnDQE8oKT1nIttffFY0RHgQG7LTcuB+1IXiLhb59FYTMBnsWgqxu
KKS6j/KdosU5MCtC2QK3wrwwInzqEYFZpF81giwaKNDsRoIklhwitid9Y0OY430K
wUY0UEEuTuRff9ZKCSOsIydEYwdBdfEQZ/tw4KTuvTh9UAJwfu07JJObvx2sdE5A
Jv2SYoIa2OOQSZt7MBUMH1v8FRxZEzCWT3AJCGJhLfywbrVvUPg0LF/MNltQnulr
8ovw/cemLZt4IR3J3TaBki/pHuDyj5aqUOl+uL0tIOgMqgLXb7L+lDZG8xHH021K
EzVPnQkmsZexbscEmLd93KPIUa9MdJ4rsbbjF0ms4oBguDc0XbwDucXEo89RJl9e
ERFRPRvJHtsWmRu4Um48mBSwqSAZ99HGLmdMPacx0NJgsdAd1vAoIYZnXl8a+6JB
hzS/BFOhJampQjZpx2GnRTBBXQTDZbxtzW/Id6+3eDJx6KsQ3mJr21XYAKae0AnL
DwoZvlAjzPQ5HEjZFfgz7qf+Re5T1EWSsUTWRxyFaQHWI0DfPnCDzBjpjJc+4ZiF
FTX0iSgaWwXzfmalsPJ+rgkMNXNvRywp4cKil3mZwdWY6jPPwVxlrTzFYKPj6dpr
rOHEMemFohgIjzrfBrmRm99UGTYhwxf9c3dtXEWu01gbk2PirZTyG1Ymlpn5Wf8q
sygojjLxFPcvyl5Kzmru9Dr0IjQEW4vk1gcgO/rPSPzzCmrZJGdT5N6P521+SI8f
1Od6hTnt1gPmN8jsremPGFn3PPIpDWveb4MLrvc/OxJwa8me2S0zRY2mi/Sh0R1F
psQhUGBmN3/f3ZvxdzRFYr6663KmmzcvH72CSKNgCM3/JM8JIjNj/3stYvRoKxZi
jvScj43i2DqqTGy7Ftf5uUDFNXaLKV5p2gHxHWZ1Ow8+MK9gnR74pNoAhi3/+Jvn
3wq5OVVL7aBONjWUx/KLH6camTa3ByxNm02zaxOsR51OwTS4uLZdFDyUMVpEF9n7
BRDTqv7//J6FbSH92Wors6dxLPb1y1qAznIHNlQqry/jJoFWaQg7CTDdY9NfUnN8
+vscxrPqSBcNlX6wQfhFLMFSOjpvezIyVHa6yJ+gh4RHV2fkhpwBWy+J2SNrlyrs
BN7KZNOMkBMz2F9RXD4oQGzO4evte0m9NFjSdWl7exRuE8kYmHqR+Xi/3l1Vm2sg
rUq/6PwdTxawjo+oZVKN/Xy65R/i5nexDPREcV7DwWYQGHGbNXsp4N/GqpgVCEEC
Sz+gFK1GFgAPB8RGLRRXSVgP1zhXfOz/j7QnOevTxiegEZEm7zpKg+yMfN5iZ0kv
0D++Zp9d+ts96ESYtMgU3ONrzWgQCySVvke55C95cL6/c4G39QKDC7cD3Elp0f/a
nARFOzDbQXOFId3yplrWqspCJSTF3zCdxB8FobywzIJ6gCyG4rVYkCEbziQKq4Pe
0IzEoZHm21Xpf5DZlSWRCa1PVp552VCOznMapAs95W2x1zV3lyDrgyDYEFalc6+u
Ksuis+1HqA9KnMYe0LHt5ieLJcj3O0qj21Xb1WaD9EdxdXSXtG0G/1hMjhOePGDV
Alwvf6RU2VtLxgmYiurpkrQrcZT/4WHnv6Hcfxg3Edtv4AOwkO168kX33x0578qY
1D2aS7z64z9BkQhWnEbtcG4fTF/RVbPG0oC7eXHYukvY/neTaLn67cCtvey7fYzg
+ij3eGYJQrkjg4zW+5GVA3AKr2MpEX2Hdx4ouHBb+RuxAJ7MtB+b7GpY0W5hsBFQ
NS7aIaEBaYFV3S7CX+lV6ODf1dSlxA3owMh8OMzy+Vt74n4rU42Fj9g7ZchzQull
KLhCQXfKslogilQFi9mdwFJE+ZZHGdfDp3WcIiHMwE4Y0U0ErrzlrmLMXeBfNteH
uY3EdHxB1VyWItGMl8u+zL1ucOsd6NP+aXHsF0XINtvGdPnISsfI13BT8TBqLvNH
vERaurlGoOfKmfrOMrYLoz5ca7LkJOSDcEUxRwCaIBcpOPrwoC+qHCa7ScrSLCCJ
5APJC2F4jnja9CpCLqiuefXwT6eukYOn9Cga1CRydRfvIEQ8YnqMAG3928+vx39t
xv5FkQvcssaRmfL/9jkXdeAtaN1FCw3gEuryargQq+g4VuxCTRVB/9N/aKHcEQ5P
0/as+iZaIR8z5HqRmpJaWQrcakjl6ebgW+B9Kk5/K1Ho4DcPQuuJ+O8wwlLQ9gmH
S+WU7r6ZRv36r6VhM7W9xd/w1hQUwzxaD0cUFwdYpoRKTnGiULpMM40/KaqYI+Yj
ijV39R29A8B/F5qhV6G337gdmE3VZYEgsOUwyhj4YMyfSqM2AsVUZh1ITGxVUUik
zAhW19Aavt8mMyh3kWPPJF0aMtvJab35p1WDXPFvzF70ukr8Y34DRV/qWOM1sfC+
Jqs0XuMxEyZYzLY7miydhJ34H/0INv7NmGl65fqAPyLh3Zu2f3kLHk3pjSOmjmAt
9sy8LmuTQRGHXVPOxpc+OhpJteuycPNb0Xm6ThqH2hnEctcxeu3dUtEVPm9E2VSf
hRavxWGXWrks7pFDjJGF7ZxdNgaZlHPb0f/1OiYdNbyXqSTnWoWhk8Mbhv5k1AgK
IOdCM3VIzIW90znIItVvwUbDRKtjmavVuaohCd+iGWXGqKquOCYoB+jDcRBO6gan
fTomruooSW4L+KBxjvFJvNEa6RfNWt+EDqmt57XGRKixS9SspDrfO7mlSZgpzCB/
CzNjFDK82Wf+2HYkaggQ+m20QYR9R9MlhygQbVNZmI+vjnljVm8r1kEqyvV8D4d4
zOnJ9FH/nPxlv4vpJDhrDuUTWMbqBfqgTE2tsJpE8wLsQDOOBGcvdtgcjFG3KOjL
SHDtYZaCZNtVyEKLV0lPSG5M80JDg+on1phRD3MohpKPctjbE0+aTZMRwKR7GxWa
0ZgCUO9OKkDDcdKLWhWeihhfkD9QlycBWrmsgscbRpXeevzHE8YlbzA4j8fl5dyk
KYviMTOuJDdOF4o1oq0Y+3Jqxa44OFmtar1ZbSZdjSQb+j6oLO2fk8I7namRD5j/
qmIIVMnXrsPmmldtyJgucBGvj9N30eZJo/ZFlZBSIoEdbBy+awzPfnnrHY5ADYEX
WM89XUebvpSt10q16hb+QuTr/vxJXi2D7zMQTNwpSsG0JKfdab+VWtzczUp2TM7y
sFRlIfgqLvyLGR/LmpB1wae3J3vm0DR1VOCqnUbqzC041dac0yQOXGyGPQsZXxuI
/tzazXib4dMiG2LSdmKh8H4IlldXbxf1NdXt9gIotgvOMf6B1gmCEKnobsuJu0pd
0u1HZNpqIa8MGePM/4njFnqcOaxHBJ6j/af4veTXUo1roINMGowchzyRo1Dd2rxv
H/mICbWqIiOqZYqYhqT/IQdGyRPcL0ee1HVgDsGJw/oz3gB3/Pa76f8Nqyl7KZv3
G8ysT0wHXRW0v6Lx29ORcYtPG2mOm7i7nz2vZW2RM9IvfiminK/ypnqFA5lIxzt1
g37riZYNjrKiSuc7mRtUMgoau9m/Sr2GY+/lILoFf4suzt8f3cs0qbqXeA129lEE
kltvaruKsK9yXBoxjyGjt6De162BHtDs0EOZbapOaO5BKfm7arHeej58oHUFdHEH
lP/xRYUlu5dIKxuBgCnD64vZ5Cf1Cbax82WKne44UgEmD3I71PpaFrLPTTd8jSYt
Sh35Nmm43G8xdZeVaQmuFv9nbkDMIG3BoZzO0V4wIWCmCZG0T8qOR0ZcUKn/mVIv
IhvJ0PdvJXe2NLwVESa3Ro6HlB6kfSvLIdfZZhPeA5X+kfAt+SJlIc5TQN/XdRE8
u0HddzNiVbVPJkQEsLWJF6Q5/kgHOBgCaS3zwbrVoVrQWuijqBjwZKd8alUgVcYJ
qYdfHsJZwfB8Q3pjvYgIyza/4F/aVP9J0nbsxdvk8TJAng/rVWw9aiRPREsZmSe6
MWKFiHmZ6Wj/YAWO+1sLKfOS0QfK0EgLusKX1YM0Zs9OVqHrdKagVNudcCp54PKi
QP8N0jffnI2P8N6c/+rDhQFzO9CRO0ERwbHfAOYlVWEdZsvrfZcaDNmlcec/oEBW
gnL/ZBdo2caV6jG91rolIk/OOs2FUi6zVevgdUzOReNsLi3vxFngxhhybYBV9l+o
rUGu+5sHQKX7U0vtdT6RLBZrMQNUozWdF4uD5Gm4PG8C/Kryyzk7xK9wHmrpsSLN
DsNtp2ByEDI/F3bt6NcDFjgOHZtkKKZ1MPbpdw1mjeHbNOXb9GFlOh+Rmdo04lhd
bhZDK9XeQbbvsrtE1EM8wK97Gq0gpBf32nvpOC/lCYIj1o2ChfZJoMDu2xqYqmA9
/B6pgqoIREfcPsFg2QROMOsTsTH8Vft7nwlyT1FGXjFRIXEzTxfkeA7CGtGCThPO
C1BOjPHTp/ArkKCmAkNN1h5pRXAQs81r1sI5kqrPiocp1XqhcAm5de/D3hB/BD6y
LcMpBuNpI7jwt2eYcMQT0V0n9rqa2db6asBZ8O5Q1By7o2Nux6iiekw6ZH0GeJNp
4tGGKn7xxRUL8eZ4GTNyhs9zm/DTVAI+KarnQrHfiWPXa0OFKFpO4avSyBP9C/gF
mb0sxsF97XsOE74Mxm/P3VN/MvVFEH/EOLe2HKebmTM=
`protect END_PROTECTED
