`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zXV0n+laBm4z23Vh4KcVWvXyNiqmGAIRWwIAU4gCxi3O6FOgF7Q0eT+bDf0r2rBl
Qy1myMEojdtJxbBtZc/YbfkQ215k2GjW3uGlHnkuC3ZcH5JPZQejmKl5WsaNP+RH
NQgD60mhYtosH8hOBxeRTR7mm4kwwME+buqBvkpQ4HRe49rH76TYVtl0pWm6UwMy
WT/AyU70APfovM0eI1rgAkL6rQ55huUG02YeV53jdDH7G6dRRuwOIWFO2x6V62zd
QwRXKl7G0FR3ZZoKNQfAg5oD3wUJHUQ7uTu3kZDB193KMZf0vrt5bVzaObjlCz3m
9DkhGzxpHKTQgrfPywKOE7t2CGs0NrhPLZ6OWDB37jXRps202vRiGJywkvPx0vnY
`protect END_PROTECTED
