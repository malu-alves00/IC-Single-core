`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5ZkcujTiOL+bcETXGryKyc4OAC+zOvARgEcLxMxzUYtPtCi0MlD3b4o0sW205YQ1
iJBJPagPooz/Z2a+khRXPc7PNlocmtD/NMjP1G8k2yd6KkvUzAmgu0m8xpiSHq8J
GFgL3WqNvjRq8sGgRcmJr0KtB01yyC7Tzw50D8d7r8g0w/GwvIhgfYyaJ9RP3W7w
F+PcJ/S5za9ewZkVMWKgb83TjrKYByLkXYaK62vtrLVipfWDQE7Hy1p94jKSZeqI
rr0HGBN7l2ObmA/a2G6NCslwnj7VVOB4TDqVhOnFICmNUZ1bsZEiUFgC6lSdpgIj
IaLQDig/c96wlgc66gmXTvIC6iEp0H0ar5GYoq2XCuL/gdmXkTq2z8ucoOIbFs+Z
SNjhP6aVeenMuerMMU1ZiK8Nu+PRso8jR3WBxV9fAtUh4S1mi3MG5Baa/G0ov4NY
DD/NIPOkAok3IkXNmMUOtenVejAHzOyUXHN2rpo3/M2QKpBrcxSTGfrQ6ANeS4Ps
bJV/IIZyXf3QrgnRmixPtpjuA2vW8LPprrD9LkaLmrGBrLDa4CJQcym7Afqq4Iyj
BEExJm04bDQFL2Tc+XV4mYvY3+g8O+wHqrZO26GN+LyBX2v/p/Kjh0ibQY7Yjb6Q
MY259UZ3TSGx1v7EPJLUmxyrPelQ5XTrupQOHuX17xslDqiU4tsEJFx/Fq820+3C
o9JbWhEmQPERcYGm573GRJK+HJn4C/jmXxzumCzchCOY224G/h0Avsra3kGi3mXy
YfAkBLPe92vQpOtKw7ZSpvzwQItPhHORgRaPbkDXwCjejHXNr5yXGIpzwMyk0bDM
cdLogQQmNjob84e2G5rSLQrgHZ/8fT0vizKR/ljrXo3OMQUozJ1xNF43j8CfB9WT
1d2awW0aQ+4viCH0DdKzigeAJMnNjCMKmFBCp6TWTudAAT7UfN2B9ty3bNZp0hjd
yxYmv8IDEbn7zXI67E7yG/0Dkosc4FHa2eIf7P6pjy5VvyAxIHaewe4A3UoNb+8I
89Pa6MTg1QuMSNP7ZTKNw7YtGRNXuydSmixvrkvvKIbu1GagWPfU2Fbm8AYyyhhA
7DGOY7P+lfmjqXJpZax9g9j+oGl2Lq0sDC0RUaAkzAnEQNGm/iutHmkQC444+Cew
pr/vZoNMVRkaiO/dS2n8wncv5ENeW61w7mQ4/UBzj2zRLEmokwZXuCTfQFlJBcXs
vTzmQTHwFxBHck8kb1NhndL/jRj7V1EX+ra+BtOGhmbEDWmeKbvRIBIlDvMiqpms
9W2N0n2oI4P/LMCJS0ztnWYVVD4h+Kp4ZqvG3RqKWUU8jKL/h1AuPsBP2mvpvEcB
nSyxkf4UMQYdfbylzizO+c2xPensbFUu8JFG0eNq1KA1iHwwTK21EXX+869NNCjs
6suzQRSMw7GpMyuq0hjirOvtkowdgE9/tO6rAtirdUIp7o1z3CuETFACWS65npK/
TlnI93joXQ+upKVUmajijWIcLg92gJ/vfcWEZejw2UGqEThos+eoh1OoFJN6HTsP
EHvjrgRfLE4XI15SzQgn9XUxKi/3bIYcXrzFRhg2IzBnYsTggSjAhZtZZY68BnKI
JrxzXi9AhI60kjMbQ6az23G5mpYetaN1krD66msUnZ8bXArrhYcooGL5xd5dnQSd
ZS5qxkHA0C2GDmeMC/RM9oG2CxMxm4QxC5A5ORvGtUjtSJE1hVvKnyCooGt6dFRl
xVmKdPlRnA1LlXkrYw3F+diUAFV5KHCVP6HJbq1/Bu/3fMt+Sl8EerkQaAJoh0ib
oqFnCaEwbw90dVDhwcviVuFRT5WPKZwTIWIP9m4d/oQXMXunZGgpt26b9gflYtUE
Mn6q5wuVaCbJpzkM5oqZDD1fTNNKEzeF5wn/HaMuEicZD4dGl/jIV6ltVkBZs9of
EL+VtyLiMYTjpCrRi8cxXHuyoHGNAQklrsefmxyjVKPosKvAy8q2GYVu3AjwSqrp
LXaq8MW8jy2RF7oY4q8kVRkvhpI51siuf0e8BVqjRe6FdofcAV3roZocaeenbV0W
O7wJiba/GEr25fnwQ7RJkcIZQQJivKCONwd5ZyBzm+kFTfjjr+za9+kQe4xeQJZZ
BT32+ZXFrG2upRp1QyVmWiwrlWeniLNs845fZioulAJ81DqZSfx4HelLv4U40rkS
pr8R86NT3KVgj5yXLrLbgNxHXRcR9/q6IMpmhsqyEfotRIb67tT7t1p8pOJgbddj
gVuwSOjdUlJghQSi891XnI6ij+8zh7llO3kAJ3kmy6SDSHz/8d77dtrY0ABop1ae
QxTss2OUovW7ycdHrfr7cz2c8tao47WROfRJj6lwt1Pa3GglOpG4liU6SdvC/gyO
Dr2O0EEbTIvlb4FfwTFIPMc1r6rZh4bHHs7kmWDuTRGQXxQ6ABzmhlTs/auVA2iH
VkwVpgLCTYXekgCQgr56vfoyh4sVj29MedxbDpDE/YGu6Q3RC1lJqn7ePVIu/yab
GuSp+9Nby8RWz+HlC1YekfumxdE0OfhXd4eDmAMRcD9VynwVgxYlnjXOz5Hu1TPM
GrUDMjTYNyUMxotvN1SpwOYhgQ0pa1f51rCqM8W1cxBNOddeuZwVRuFfDk9lT8Xv
FVyi5rwLMvkmXpoKrQbdbfc+d4LaxVYAvmhtFxZ5h3/VSeAnijz9rDbxxoG4hd88
FyrG5d3vaZoI/ll15/f9sCPWO8RSZ9wurCf6K7J+6xyNhb8ANqHVEK1ICaJF93h0
0Uu44+jZs4TO8yZHBnroT8r0T7ZaVE0rCnQNWkD9U/yf1cO+aF9r7WtL39ggecM9
qIz8M1DxbMf8y2nxDWVMHs4xzDMQV1AprhkJa3L4GnwQvUO8xngThrAKOdvZG/08
oSXGGg1z+Lle9ldgHiG0CpP5ie3qfcpzU1ESF6TNA78dYFGwnByOz5ko4nx+CDaT
2Elsb0MhgoQnxx1RAvQmZJ9VN+PRRiYzPC0P4bTSNCBF7zg70mFrHMcE+8P/K4/M
YA1K8jxkEQk/jaA0V1siICYIW2dupQGZJ7ho0P9KbuKEVeuZH3Xt7dtnk0UN9Mxf
RvVMeJyUWEfuGEVFvZKomUIuucLAzIiw8rkZfz8pyARKTpA+tRkreI5Iw05kS1pM
ljGQpUy+vik3UABgJea5a54fE7USc0dy1Qp+JiG3bvcM/H/c2TI7WtVEIMBxTo19
pgoFIsfNw5kw5mB85BHHhOQ/j7bjoSwwbwSKLX/pj3ZOE0dvobDxtwwwNwh1c8HG
lVZDv6CVAfWu3Hxegi7sIuquT66fwArJNk6p5wgtq+gr7RVGRyoZgnt35zgcTh5g
/KUX/6+rVRxPAdtsmS3b9KkEi6mooNYZPqrc34QL6QAAl7SYtAFn/7UvlCrGlp7V
De4tCKGBqXarpu6sy2yHp0bV+uuYemVpSioRjyD8ABpkA/jvOb6OGMTouA6O9/e9
8C7Yf5a3X+KMSUnoFkQwYheG7ZeHaQKFMwz6q9/rtFKX44t3HDAqTs0plykO2QlH
KkCaFkRmBz2D4X3waRf+AXeKJzS09syKQwiiTPOezMv1WRTV67oWwIPF92tA61hC
GM0DHjBO1GwpPho3DAqXfALQlkt2nizC2gw6qa7Jud99kqWHU9js8TsSXPd5UOnq
7CgFZDHyyy6eJrHBzkMcWikudV5so5mRVyHhd3m6+gY6LTmsARZPrvgNmiDHxRwy
86+8qEioxXYbXdN7OTMsZ2nHPF7O5Z5Q9Llq9jUZ//47xuxb1Zd8KQoLQaD/AYQt
smRNre7J9hWMRON6LxI42JtAyTtYKh5AXe8529Ht63lLrrM2SmpH4i3pJ7XM5E1O
GZr8MMDL4t3/lcZaWLNcampH4L0mImOIdSEki+5rpMiAbY+tK857vmfs8bunSMNh
l7xGKffaV1H2DQX7Ztzm4aESU3RthFmzUUxOE1FNSXwW6JOHEDgGNGOEvQ6XGNOq
+aId9zw7KTbEobpiv4rkCvQOgYuwINesVWCcNE7dfJT3P29lK3OP24dYUMz+roi7
f601+m7ViZsXTZWvwW0P7E3/zhaPj6V2/uspHngxD4M5TICxOUPPsnPddiqrXCAK
SBgT4iGH36rD+xsStFLRYJFAaQs3gLzMDzbac9IkQwcegESmqn47LUZagsMgL0Ua
Ps5j6ta5Dpr4nhoQE6ZG/lbOV5MNDZEV7FVTvqUjIz/TZOVCSAYbVOHPtqqmqH0h
lXh/2z5/oDbRNRVctTupcCS506jnjfIQML2xHJ68ofPy01a6m/PTWq2k70iL9O7d
3gpMOkZXHuTGzFI2oAXrDsO3B/coa+XT6lJhiVYLynrkgTIZ2o/joJw2fK6zyDGN
E8Xc3pZRA3Mzk9A+TWO8eyRkHzp1UXD90l6R0KZ8vy/E9VlWFvLJYEpMXG35eI/f
EvxisSSYfQKfvTdyzyPfFPsjTpFk5nEC2nnXOTiVWWQBtyVrhSbab7I/6biTmHgr
Vn5gdMI53ygNtCQraDiDSZNDaXw/D6XooG/DVF50tXCQCcOvFNJLC0GHcFEoMnZf
tp+kkRY5SJxY1i1d9LPQpzJ8/drjkMgviu/91V/onBHtKqmKKhUatG1UT3ZZC3Ol
CNXpEsekIRdffWeNzpU/x6bxMEefiniKYlqb4UyrZTFR9dah6P1wq3W6oeBQNHu1
HVufFBdzeMmC0AON5/Mh4Sj+VmOzLa8KKez4K4kz+e0Dcw5CPmH76Unj+D8hbjF8
vtoFBQWDCfEBmfIlkOpwtvNN4JPSBRRG2ghCxewNsWa7Xxu5ll8yup4u6Gpq4OEy
WjmHBAGZGUwrYiU0Ib9yLkIpKncEcxGYs+Pc/KvOq/5Ig2of1hgZwA/kM0VcPsr9
kht6orWlHfMIxXBuDPKTvOPANAxdKwwlnay36cc7ZH+ZW3Guz5IVphTIJ3+iZ4dI
Avtedu5kNZgxbpEvb7Ueb+KgbbF8wU56aIIqdxF+Mlk4SfholiOISE3s3PW/sANQ
t4yM/pqbGJUiGaYOOlRgmpAJfF3P0QfCEUeLvCSKrbea9zE+RCZ3mCfW3RPWx8mC
ebz7GrAyX8+j6B6iWTxRCaWyaXA+pMopHxYcu9X68thdyHW7WO52cbGnsl2UK0Nb
jMEKH7Q47MFrXLuk1LIqcAB1w1oFUjiCNQi8UCWwmatpblRAIH5MwQto7m6NJ+wP
2nPRY+eLQGhYw1Dcz7Zk43YiijR60WGY5P9tdm0qvoDplf9VLEMIZlyjlQcLJ29w
KJcJhjA2e64g54BWbK3f8YQxM4pDwkU+RQgU1D7Wrlck+JY/uV4Ar1VFYZRnr/Bd
etWpRnH8hLdMWLUmMZ2jaBjAn4aKSk+M/90RSnrOQ6Sch002JJoFL422LwiNr11v
B97UrMEqsgETmyKO+13Ox9gKmMcJf5nHp/Z4BFMFd+uUmY37EmmF12Mz8VF+tykt
rQJgmDHTo1OjyPJhxwGhyXiUYpnPrsCKQuJH2MIoCzGNcbzFHSmm8Z4lvO5dGFKd
lEeR1ISnLOC2BUjVkVxt04VqB3PKR25Kq4AxTOlfvob+V8iGhHHoDDPuo2tVb9Dp
M7zmC9ko2fy2asbvZKwYr5lcSCTBhHnEcFUG224NWZHW8szGvMqBnKyNbnqEcSg6
Daj3FHQv8TAvHD+HKYPpvqp+nB5hVP8vpkdHDTEJ14CmAYvC4PR3uqQtiq8wt69H
I5qA/jyQx/h21dqjrsUVbJSpMV9/VjG7FNZcOV+4APIkUqrWKd/0Om2iHz5fpCgo
ZVukyZCQ44VKooyYFmBqYlnq2wzQDhc6Bz0TUNzKh5idsLNKGMwmcvMr7i0JJR7O
1gvuEuaVPHH3mSOk9tHAr1kmFKSgKLn5mA1D2Q5/1OKg0YKzNld4Z2i33u6Oomom
PBzEaiA7bNR5tKXhIvENMwQnizCojgTXW8Og6K+vx10QVhQ5/J5QUcfp+VOVwjPl
sJ624+JxdJESk7qiiC++ZPRtzWOYdhU+lDAolcY9KE9I/jQYUZJVB+AyC0sYOgba
774G1sr3b/ZfV9ln4ovgYqPDTivsmPnxZdfXHdFpItnVlYErbkyVnVz3YKDc1ziZ
O9+MXHHmFlCV44MJAEuHO0lKgjghSChF1OlgY4NDS4OVWuqQdrWJEGG27y+Nty9z
sHvD3v0Y+na9hdaox+AD6bwS5Cn4Fc9rL1VfvVfnQffAmWOhDYdOwDqA2A2pahi3
igZXkZPUHsbIgo53GgPAAPNlf+x+ErNjJOEuoyzo8mkh4QsJ62qMOsASnpkBkk9V
wAqQ8MP3ncfJyjhbkxXujMDTr0mPzhUMhY8JmJHU97ryHd/4Ipagx86q6iEgzGp8
WL1dpGZKSTIIfqGAR6ycITRIRkSs2hWCH/s32CpAlMLHWzXrqMc1K39rxz3fY9/H
a2mNXGFVCuJ3yIso21zNHAdHY8NI6THcL08gmUHek4gBiRsJvRUCHqUNU9H1VttB
FWfIVD8pGnwMmr3MIe8dcXgmPELbChnWxXtemhk3kPjW55NaemKirY5mNTPy5LD/
VxR7doyq/FlWaKgyO9HiJi7yUAJsKm8QH10B1u/TIsplkKs0gCGinoctiovqcq3P
HNdmu5VTYV8PUpouVlo2Y6+8kwC3WxnG3SSAvHh9PLq9DRtwrPs/GBseu4wjJ4WR
x2HJRTdrgdQqk/urrbk/RbSK0pCMLA4HiapXFk08YrXwy1cgpNB7s92HKwqcmvq2
D9lZRMbAzqlF0rnUl06vBu6LmAQI8p04JgnLS/ptgxJHBnDr1FdaWKN0ZDSZlTSe
vdUuA7fpqjToolNGu7V/NzQZ8R9DVjNU8j7sIe6JrM3RFk3xegaPBOlZ8dUQorGk
jCjDtYNHm/f/s/yDwfQ60BuvXLelKoJaX6PJ0aD3cWDC3v6PYLUW0iDfknLTLUWi
dTpY99/55UXdGsk32tGKBIhinGmmWAYlgNOJdDdHluaSZzzVnn+hgkI8qLK8mJQh
IyXyrCznyVHWpm65np9EcjdV8iAPA/V64cqaMW/0wnJuR8BbWESlRTYOSjs7dRU0
2sorF3ylc8a3RvMr4KecTcVVp76eO/iQR9TR3umbTKwrsrQwe6EvU9W2LVNZTfa5
Cp932i7lJc/5TKMuV9Urcc4HulHeF1VX0hFn0YBj5JnhuIxxIw8kOP8Ceiz577PR
ed3mD61EdoHVPRIG0arulrA09lCtUHaZLSbykKqR9HCQcrC+SPRqKrmqUUfz4bnk
etUmMQlPiAS1emNHf7z9tQXwq4L+eyTXq0L0P3QkjhpNbc1D6FZNNKbyPT6cYGWk
tIp2yKLonMSG8JKTzi6m0G8CsNoE9mMtIgZdlbYNibdo4ftvnOUYa1eXRpIWyGU4
thZuK7wFe8TLnk3tEXE+iGuAGhIICHWv05kgJNTkqBwK0rUrhRa1bhBEHemM4uRp
PsGAtH9FS0PBSCR4Oc6yISVtY1Oz4FogxbVatIULzMhGRRuktGRPFPY9qmY9qsIJ
v1f+UCE9Xii9KHNsRWWy4Tl53GsP3VCMbUWC2gZnvpN6eDQHlgSyJc7fINb8jKxI
N7pCfwF+FoZw815xLQHedMBQtMixTVQmEzbBIe96jZK82Swj+FHK9bUAjhl37OfJ
ZBR60tThOaL4ZJsR1+BGEoD4kdgTzV9KkiBV1TVLtUwtnfuUwzNoMbzmJV47q5JD
uofQiSZIDkU3RGrP7/+RXZBXVExB/n9Azx6S4Bx45r/1x5SV5wBk6kp0J+EqGIrB
td6cPVrLgYIVd8ZwLvYi+9ES7vdZUkaQ87d6FN3Jj85t7VFG+giJWZUzinikjgSC
9JSjhiNPGX7R1+jSvohQI9FYGRvEBmdZmAxIcBzntxN0b53TUAWzu10aJ0eoz1jM
EEFEREY5x3vnOS2ogqTgaixrJi+cAGY7JLfEfpXpAexDeCwxGJ7GyuyfPliUqAHf
/pkLPrZDo+zAEpYvJVJGBIc9ZfzfhVkj9dLraTTY3t2kI7dGUQa/R/ady7Dr9o8F
5A3aYneUgQJJs1B9gzIxj10c739YFMT/l/G75I15MJx+5aEXVCZJ+ryq5wWGf1FG
sdEZQjqKehYQrCjr232enCFhhDK84EuFAD7FpP0xp6r7dVU3J2KCfckd3KDdGozN
TMbGGslOWygTiQEFYTIWi7X7QWUi/tADwPNwfIFdeV+DdbuaGzc0cfgFRyHT69n0
zAu6FwpV32l3z/yHA6fjrV2Og6VaxdaD2Y/MGnnMTh7JxHBiHt6L1rqRT+p+r6Lg
dkz3CvvsQyAiQIAxBw2uMtTJpnY8LrSEwzTQBg35HVTIfE2p1WB2udVDidddO3q2
e1GjCK95mP3KQFWECeM4GlqNpOMXOKUIjQvIxB4FtK++6dwxvmWE3dl5bWbR0tny
y8WRIxIRbCL3Jal9oK0W/+nFNYjzWjFiV0sQK9e1RBLBbwi5KmS238iwzunssDt6
HPvtRjUWgYPPTjQEF2xrd1Dk8JUAyPyVBRC8cw3MbWHl/8OZlQe7dZoPSw/U0dH7
ssMPW5S3OyiuVqfmYxW/1NtGdhABOY9bHIcjhj0gIaqw2eebqiMgkfHnLXXl+3L1
KmvhDYLfSAI0XO/qfQ7JMDNxDwY0AnEMzhVYJHllf5hqnXKzgdpRXFz6Y0Ui0Kq6
ibR/C2dGqNRXGaE3WtwNdQLkWH+z14hkLBwOrMHtAXsvdLG+JALJdk79HKM+X3Y6
hDHJcS6sCMznIpeGiV15jg7UtsIjm9/l+J8LNLBxSE1ZgPVrfAuETnSKCxt9bPKj
iwB0WG0AC3QVIW2HVIx3b4jUgXplcUA5aMKFFxP/IVKopgvgae394z+sPPUqHBo2
YKYmPHFasHHx9ArIyzgDthDUEXXRWgbUL0ljWYY9/WG83TVAxZ0OCmBidcMjLLkU
wo6cg83/nhyMl0lVLxdHDcjFoBZ9hsH3vcwUoRkfKomqqJ6Ze24JQaii0tNTnIio
Es544laKPuAc9YKdOwM2oOHVYHisQQXN2T3Zz2DLspKyHOn/r8etz6eDSYnYeLXN
9xjWH+doAf/+0zfG2llCP9sxZbs6qCrHjJIEHuO8dxkuuEniawz7/kWqHD23X37l
zGCfsn7pSu8wPcrhJAMITVuZcCfsRpAd19uW4ORmAVrrLUnp5GJWcvrl+I2AuxpS
WgAQM935v1AOHdgj+wuuB8EukpJSzdRn5bExckj9+a9fZkkhdEONrJTJtn4xmDW9
QrX757bDBv5cddYCyyKRSTQgEBNuua95/OBo1clHyHqtSB87FVMq0Aov5nnF4Wrs
nBKnjsJYfY0vLQlJYAFUob6wN1xj1W2mFrZA4zO48HQlnzK2kwtbJoqodqa+A9Za
WOJVHoStLJhv6pFgW9t9+nw62M2YM49jsawY1ruGjVekhJ0qVCPxe6W5CYKcDyL0
G4+53ci7Q8x9UjpHdKjzyJ36rtxl84A7khv+Xr5Lc1/Mpv2WNXY6M5VnCLYZ8hnt
RTfnDDfThcmXOZRdMphOYfuSNOzfxXy3sjX7ezUAZiEUpQJMoc4N5wA4X9xiod4I
cNUJ3z2QlOfl3r/O3pWAU7IeLBmNmle6seN7Ca91Z7D3qLt+TwvqUVR2zrxkzeaj
Tng0wZMlIFUFveXkYmsXEUb57Jyqiiv1EDgKcaCMUhJrPVXHJ3R6FpuFE7j4d7ih
dnt8q4P04XSsPQP6r3qpot+p0WBQFEtG5cmZjBc0Yb+c6boOrkxaLsesGeEXR7Ta
i0GyroYY4ipdTxc4BNJkER00viB7rr3uedbXYe6M09H6n63ToQDkmEePmhTdY74Z
forJ9RlPaggVeT1zSEPoGhEPiMxGMCFioY5SBWqeSXOfM08cs1qsmcibJwRv6Zjq
ETazUyYu+H5ucipx1R6yTL3v069ImMKbFgNRF2twMNos8yxmY9kJLupBUq+Jv6Fw
1Pl7ZzrkSKhKnTmIzANOaxrYbVg21FZC3HyR81cwwya7NinD3I9ls1lbF0sDu4iW
TLh/yP6jOtQ3WXriAyitsMUGAt/PSXuGlit9akAdw5D8IbZ4y+Q7oMcGukI4TlHF
b4rDQIL6ilOEyjemXQsuiHYpEE8PnrIIRNUXyPYHOaTn5mRLTv8CLxYdBprH+8de
xfi1H94rm804Gq1U51vhhMi5Qb7W/LGUz6oIJ8zmGQRqqdA6eDXZzbjMk3I7IvUW
qMyWuQC65T+oYiZt9QxhMAAOveCMRIU4BPVRv1T9qHPkMaX0kATG248UomJ8XuSF
KkjP+tPkDECk/Nw8VWPcG5t0ZI0nMi/rVi60BOy1TDFNNEBB1wCqmYqVdKS+T4ew
Mfi+L8MwxWqOz2TFzUim1vm8JVBMCwGJCOvQPnCgsIU48vt4Uw299d0ORxv3XLlX
ZYJWvlfQVWjKErQvG4z2LJgLiYrZwNk0DXuWXyLr0oWjd73oNrI7gcEmHcA7XIuE
PaIdYFgJR+U3kFW6GvQ9Zp1M0jw/SKFYOPGvP3L2N0yPas1HaT6PN3hRK/VUXUTs
YkFe19o9nM2wtzy+gxwyhaxsxB75HBwRVN77ZToSvGK0UCKag5kX4IbqQSwAKSfR
OMDU9nzx+cVl/xWWqLAkrcZPWgJMzQp9nezkbn3nfXqtpZOFao7q6LzgcqSxPT6x
dXoPUWFjruib5ejVcr22kGseg6R4Y8TWXM42inpFGSJ7/4ZtLzTMnUSHBbFsqrvj
QgcPKGayqdNuw6HQwNlq7sSZolwHeYBJrfVfjrAYIdlnTLXWLKkyYzolWaFYQTSC
6JRVbh7P6JfKo2EVaGWP5SZAxc1MPM1uS4hET+Q2Fw7BdWhf0xBFzIgj5V8oOFTP
yq2i0jryWsgQ9CfQ6PDEmyOVu7t/RZC9gJd1QNHg7cmFTTrXWdyWSEoffy0YrCRF
WndKmEQx3PbzQUPheqDuyq8kmTDjPXZe49hgyqA0ahm3A7Pwwy/OAopmuHHmePye
muplxCUNXhwadEh51Ies/i/7j3RobYe9mDeurB4eiOo2m47yddmjx4vxcP/gIFjE
iMdWp+ftrWlahKBdcbWnd0yhCvAtl3Ece5HQPBSTdFgsxwVZLuhdEl/tW8lqnG1W
9ZazYJwCbIfYar7BukssrpRwnPOPVgAvOBBu7umQGTsbfDKbxaK5yJ+kAvh5PThI
PNJVOdHIGSeU+h+DOLL0+8d0Ws1uUwmUFB8KoTf1YCxN/E4L0bEtfeRJyxhsHj5d
cYkuQ4JemmlXmiNsLd4MLqEHjBcVxa1smfwWcaER6qxViaO0e5S146WsVe/FLUIi
XARuu7JXqsmzceprABvIH6agUhuSytN3tBO65m9tDd+RrPxNbqrpv4uVmKsInZ7/
5CZbwfeVr6ktYQ/JviambLy0tgiffyA19sWZmtgIVCliFbAx2g0r9t06RaLjC33y
FR6gG08Kf4mv7u/yukAsuxzgeNizZ9znRzT7I/QfyeKPm/22kkxzO+1STiUXWSov
+X2vnoCrwfbii2sSQaXIDU8vt7scLxU+JWAJvfdwIQBdYtePNIs0vFRBOrg0ugrk
13lnf0eT4108/capTNkuGPUbLNmHNldbtix32iahd/Qzy4lRChzYaUIvtW9THV3V
4hlcOK+TLav7Ahr86wpPzEU1fQT2V5CeTwyxtcdiUMKsHUuksIgmNlGj3qg07+Ca
z0jPAhh2cuKygFgP1T6uSM/rzUiCHFTC2uISxcckTNPTwd3cW/XWNlrAh9Mlnbaa
ZPstEmoX4XohkOkPQF0TpUpgDHUM+P7J4BbNp26omDHdzQI7WfnID5ptf1x1AVfe
fUyUuTGEBveM8+c4Qbq4b54XKAMXqO7HaFPt97WmB0R8DEZ+e+aMLatiHu5QWebd
p4ehFU5qdd2OFKPgF6O5KSGCO36gq65VexJEczazHc9gXGb5KmA1FgfsQIuTe9Fc
1Dxz00JpJFnv69eNT/0DeqYXXXKiC0yyxt01nzrBy4KPQzCUtIlwLw6oFI+5I+E/
m20Z2DoptPrVWZeJ33gSqEaSnE/yoU1CIJhj4Xi0rWu+0gxr9Lcre/JRliji/Db8
yNbg+WJk58KqKlZAAPTUIsQE4Gqo8WZUrd6/93088gAlwa6JciIBw8eu9ecqUBvk
0cEQDA7DdO50YcCL83V4t8FweJ4K36cayIhv3lwm4/3vd69K2NghMis4IrDJOU/J
O8E6Hveu6wzMfMz2Yg018jCnZZmugKviha3b7NW3PJX7YoooqkpjOFr5JDGzxkA7
8uDT0wYbwMY6oHEW/n1C7uzdAR3yMN9KcMr83vtxkImJd5vIOp0VknTb4wlReHRk
5b1zdaDkL7gmF0Sqf60o80ccSGakw0gshGmJ4W04JTnB4/J36WIR9tvoSGZNLLzH
YTv7Q9wfx0TBYWlJkJv2ij85bkPVEaat7i4EDVlzhhARldz4beWCI7J/xrH/VhJV
68+ByX+yjMhkMNBb7NdAlIYHghf60W+v2f3nrY7MwjLPcYgY1soJU+eLoLGKejsI
hN2eUSh+dVHgRNzbjMtvGpr3bccA26NDmJlT+Mq46KwKWiCRIJukTn45lgWvmxSj
s9d0v4S4Ycyzl5Ack+tq+V395DitxxsBcEcx1gmRFEok0RSo5KzS0pwkP4Aa+8+f
DGW0jRAKxgSwxIBa4FC7t+Omt4jPI6eb5/v3vL/Sw6wKUj7f6TkICvNBmZoqu4kB
emUKPlhnMnQLkM5U0nCHZEVXP2+3tbCLp/MvQYmCBUOqG1cncofu21MmUSDoW10Y
HF2XmHtqeneeS2HmXfpTLQqDVtQqarDz/XkXlWBHI8oSqQuQLQREWkMxS/sDuz2q
3MDh/dRPJkX2VE/noo5jueX8zhCleHNDnE3TSMHVgnPGNPp5vMQCda1TZSh+mtuV
H1tllIliGT0so+GWHz6XYJYzFQhwRz9+8uup7DhzNrpeqRNM8uOzNlfbVyB+lUec
ywVME2Q0UkiEJLy9XNb4wbdzDnI2ah+OdYFlu5OgbwgW95kuqohcmSQUMmEqlk1l
emb96sWAXfQH+RZ2C4KiatHENOzI+K0PmwBWGPkVgWA5+oFecis/XeVivELYzCXD
O9Dept03YwBJLgicqCJhE+zybAxs5A0BaA4dKB8dUrv05WUxiV7D2t1vjxuqTAHy
yCW3z/NgqrmMniXnO0q8abqUwilfF17n13WxkkxmB3sxObz5lwHgjCshJA2S40Pp
DJ3Cj3BBolhagDxqYnqfYoNU8lRMAH2SZeMQol8dA8uQIuaSaMUd3b2muzrv+2g9
3Y5ktPxea5aCp1Cdqk9qiFjRAeX4OHontVN7QDyY3muh8EiJBSICXiskx2ELZmXx
`protect END_PROTECTED
