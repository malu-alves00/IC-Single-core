`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5sbOf5Uha3dtey26xRpenDXgPV1gy6KtMflcJR3tguZXejvb5n/Mb94yh/fRXIME
RsoBWl8nOO36x/hxi+ZIbfmijKNp42+O7lGEV5lTA6KHVf1LFRICGlpfcg31TF+d
AfBCCxAq2IIJGifuR6AgOXozKb7tTXhJ4vBfWdcC7F7T7YwwKzurX46tfxmaWaJo
gJ24x+isbm8DENkP5ZXCb2sz2WbS4wlJW9ddaTqOFn6nihf0frHP9qLbFPdbQQbA
xQCLiCOsoxpYYf9BTfeAc7Iook4KF5VIMw0Vj9bNv1NW7nTMQpFGFVEiZ9Q4iwRH
9Vm1iPldFLHmbNeQBiJ2YiKi0Ea/609u0hmEHaI43VOOcFd/fP/0GUMSpjkS3u0P
Ft7a+yR/csW+UPXZz9vKLndwiN7ycBFOezLsHaiWP4KUBz4mKVFc8UCQxYksnnfS
fmrJ0UpjJhMgn1iH0+rXLFUSY1Hr2nhEDsLGoazWA2OVqJwzUWm5s9DCoXI415cI
2L0qBpMIp8rfVGy56kZyMINBbWp9FeudxmBUqUFAYv1RYwoQ8cWmF0zs2uzDalXm
mJuQIfXpNEClUxclLM8wb8UZ3ZDy14/HbrG/Oo4VrdfW5EL+EbHkdvpmZGiguW3D
i6YWqug8aHNGhgi8/WeB5p2Tj5PREcXFItjo+djqAAtgmT4554a69ILFUki6mES7
ajr1esXdd4s7NH3t5/o0Jl/XBtrTuF4dLadeNTwnCQRkPp3Uu+F0bXq6rB6e3Uss
M2euRew1veFEajR3Geijwml/hEsKZ2sb887Wv4LKk5h/BnjrTK6t8QaI/CFUvVWn
o6ySUTAjObQrLBL2tmPnQikML4Njjg+5gyod4MQyBsKbQuL/05dMWZdfhw4WNIbD
LHBGJPNZWi8+c1MmeDdmyuTqOfYu53dSA2o81DdxzLvFrmXxsi5vxc7QioupUCP7
uZmnWbr0CvVKSSWe+TBqWyzCx2WAGmBOFxLlCiXo7yFwcvaYf2EoHPuFby/9SQYl
DYdKcBaK+Zm8LUAN0Ym7ezml6uhU0HcndTB94XYC+MacaxnpONb8b9IJygWqKMGv
OA4fQcS/nZAGWIgNAw5DHP1BRD5+TUVl5AxVH+9yfKjtvIwB6NfNTOL//052O+t/
rfNKdamsL9OvfNQaGBBnaNuxhHXIeG5Jadx/Wq7ajMuY5lRn8DpYItAqnCUukfgs
GA3SbiYiFpuHbGjbiGqHsZOiA9cJoM1oQ7igpUlpzyzaccgpdTNjhNcFWdCZm7Q5
fm71mgFqp1GgFFudzZ1aFYA4IvbPdvE5zujyrkphQ2WE/ouahBjAf/kKt7y9IeUm
GKCHrqe30/VH9iV4YXi16mIZ1x3xZexYXWNQvBwNfjbY9rd6Kn5vJ1XmclBA2ePK
AbpWtCok1qRmTYc1HDjvGX/mvYW4SZ6ghxVaexVgsQ8Kyx18v5Wg5p0jaW205MsY
oJW+aGoiQRMcrFKFbYgziNNF9O2PVdL9Y8J7afN7CfU=
`protect END_PROTECTED
