`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JpCglh53gW4x2naec1qdWr/8U2PbRDoh0b/0QKQ6lJnG7rUFdJlTVpSG3iINa+nX
aD5Hpru7RSrycQH6c7gk5T+jUYCloQBCQB1YNOjksR3X9xAjVgdHo6fKM5yrZ8Te
/V8R8b6hncLFidMBGOhvABg0lOSj9jAdx79DGasOO2Lg4hBYbZjo4x6OysTE7wB8
wacMdM8BQpn1fDpfqGXMJm5cblaLZyKp3IdPdYiVFPqWT/P38B2kgK/72ubieXEJ
EP8+T6cq9treRAJTVVgZB1QbXtSWSF1jJsCjucbInIw03WxIbi/pGF4h5hSYii7j
oquqbFWJAs0CEBM6b04zNA2FJ/J3my4DuA1CWKZvrLgKAENqAcDcahOjZjfk7vzK
plEbhGm8wi9aLC3ro/FGsnvdofbEyxxGzLghX7wHohP2nhXoO9/1lw3agWjcr1AK
tNCWffTMfVtK5u+lMQigdDoXiYr76K4hII2/773DfdM6xtfatJqy5HKmvYUHVrYg
hczxsr9hMixoET0Mv3KVNYeawpbUJhgcmmUkBrOd95dqZsqy6iJ4/yooM+tmcpSZ
jxDxC5ZQF5AZ0ocIinwFCOcuUcrr+ubWI/WklYPTLAPbW1trz2rmMyAFpDRINgzH
OWPz038FaNPYFeVMJRV9/ANWKQhuvOvqxS7A/ZIdItS2F4lE/wUY0T+UiM+S/tRG
TMRykUfRFlCHDTLYhME3C0FDybrzDiAV85tQDfTpwliX48HijE2NSKDZ+ioSY0YS
xK808NYaoqoXXAUsonM6xgGWVk9HRllfD9vXDp5AfFzZPqUdDxez9pwJNB6+BB87
JN1FBGwZeSBF7vE+7FlB0uY/3EE0cFdFmfUCRu0+D02i7dGMtPb6H0TxMdd72DwZ
otkFZRPmT8zVuDch5iKZptqlqurVOeRwP2rl4LZ1PDQtXlJxaRidytLPrT1LnB2h
biwSfkx2t8UeJptKVhId1//SuLA/yqjifFI9dqbQbEOfPiyqt1MN4jV+eBjshq3o
ya4/UANLltV+vDVbazcicpb1SR6YQVWBvi8JspcI/gVubqxaekJq8MNASSLYALlh
BDxNpAbgE1mzBV/bdCWp3uf0fz0ZErzgdzJE6viJd/yP55cEdfr5jKh0i4eDgD/x
+MAkqIKdDi5QmO7iOopnr7ZyTuUwwIKu+Sdb1uhAgSS76cDBVbVuOlwenq/DQUZ4
FuPYRn6JgwXhEzjrE4WagPkmh3j8/Z749s4Oz0O4FTcupknbKQfRLxaAI8e2M0m0
rbf4MSnRCemJk+32dx2wKY0suubzc505DVS6V2ihunnSPjYE8yjCFSqXy+anwDTF
N9AUjuTuYe3x9tSmiljjqVNISh4NHi+QSquAFK+EG0ogS3xqZRHD30jpmyjDahBd
rUiXLB43vwFhFPJKdAxt7MDJLxZ36Q1KEnIcLwhUfArOueCe6Egz7DaTSQ1xzP7I
dDehdPpVLF/WI1xzCq9vxaDkV8ifelazUvsrenFxfEaulyX8bMjAzvU45aU/lj+t
e6vZMV7AdJpoUF0kVK3KWUBMMq4T9IuAoKghfuynm1VSiMw2mcDSjn7wf152BPfw
mfOayR3AV2/oRCTWs/EWWdYB+FWJftZAnlmA6LtaqHW3tkfgg01/WKNAMyRhodSK
vdI3ogNxHF43w5tBesDDkEDgLI3MYbhFAtcvEzFmhuF0I3pXC5v7gIZ0hEX9u9fn
YteIYa9qLBeWeDbWu9sURBoq5zZ2kl8p9TdYSojx04tYIRnIVALY98cxBQYw1cjK
P4kXpJC2oaVkcmh9xkWSgAt4I56UvYI4XWPvzSpUzvP8FmYCP7o7YESsAUV4QsUD
LGa9VdxJYdiFD3icqU6nUc+T2O3gwHg5EUtVHgSHaM2HkhUoKLpzNxPdla5SY1+A
1YqmrHbmlpOHf2EM4n7dkI6VG0GrXuJ+lUjlrB/TZ+Jq5TqTsp/bQxoOZK9zCVG3
mldQvhqWbHDK3btkmn7LAC76U57yvqmyBph1SVacRl0A0V+vrgvqk2kG4OTesPwm
J08dxDyuLbOQtGuzV9/wKNVhw08CPAxFAm5QzqwVJYWf+0KlJIMH6UlMQvH7AKCi
y7XfvX4GdC+NDmfnddng9+HprDGzZA/x8BZj4mN0t9IIuMiJHiuGjBjMp0Y0HQR8
zygpWgn+eyWT2BUqmC1D1UwE+j7qOPDag7heCgO+cO5UOlPLdLVeBRD0+bqEKfiQ
DuLLYuCyQ4UTk5REBzQ1Q3m7fdl4H13psEfuko4Qblfc//1sjIlvCuSdZIah56+p
WRPKDIRlMe3+EKmZbc80WP3y69RzGNzeUiZhTtsMk+obBTD6OPVe/IaB5AMsa97R
z90BxjWaccBLnC6sPnLJyBFicGPKK0qo1z/IEoAAFj0QbXnkFbmBQ1w5uZpMlqbe
R4BhLUWbl6RWNX7ad6YRB3++HF59nzsxwoftkspU0IU2yurJI5jvsx4uug6Ffpsi
d3QFm4lIjuXc2rS6WI95Ll/WQpisDKkPsHzA9WYKpaMJzOM0MSstpH9FnYEVbAcI
vX58S402Y61fCNzKLSoRrOxezQ+uEm279PPN39yTCYHLqlmmR+PsqT8tmK8u9FTG
aR3nGymhDng2cxdznmXYzlUGCosiPZMY4+E7GQpanRxj2QwTqLI9K5AZwVpwuoPk
lvNHZwPxI7L/37AztoIIsuGX/Y3/lepI3i07MwCaV3YT0NiLNb+xrwWvP1gDkbEu
h4gOewBKmM/MuXCOs4eQtvltszi8BSyZYzL5kVxS+mJlIJz8+4f/IF0s6LBr0agV
p5Giu6v/Sr+x0ARn5d2ohz/bovp2Aa0BNDkpjPeb2y4dWmubLhp51pAfLMMhjSeO
mqHJTj2AcR8GhWu6FXlxjXXcOAKTVIg4uXLeSrj7yo5DVW1jdtGtWJ1auwRD19Yz
SkrdenUlSYSa8p/GzcN+mw0MXPJOgmh3KmmySaLaVMHOV0bsQUqSvIDYc671D3rM
MzMM9mjlwh34PzzRlrhJ9hUyEh9v9Fd67Cu6BhYFoJexJZ5nMcDdT5+xtpH0vsC0
fP0H5o562QGRJMJahy1W9SVQPd8WucFUv6UiIpcKuXxrCCQgKq6jup7Zanm9d92S
G18ipKUIh5zFwV38zVUt+KB487hsBE+T4VC0ckJ8ywfr7hJ7vsA2ECn/yb5849Af
sDvZ+3W9go/PRJ+HxhQY+Kunc0kq68FnsKM1zXHqrRwoD2g8+84efXEMqNKzJIrM
J/c5lLK5GOMmTepesBb0Lz3CQ/6/pHsaEKBRug3LOpjLExml7X1zLcSVnNCzU971
VX27bQfsbaHP6+i9MpyZt4AkY97znrAa2fyidmzbzbNR+JcJnySsTJtC6s806dqg
4lVrQIVbhtvvfmaAnUe8FFXc7nc8iiZotl3trzNmHiwlIGToEaQpf1Pll7sV+8rv
zcxmiU4y/3aS2EZWWOpPFPYu+DCSXP1CSyAR9eTU8oqSSPAvHpPUALEWYnlWbE6J
SMudZQfd36BtyObhxtw5nSAsjYIxvabkowjPQ++xL+OydCkBLcrwvb6oZy6HjTOv
C6zAWXkhKua4+/CepqlY9yKzJLAeQc44S3Xy4B3qZzFCuarb/T6MXQR7RZEt/egx
702hXgbw070Uo9C6no3jtnY3vlWo72tweugVy9Ityux6KRZNrXwGYzNbRTjbkYnl
c/yahVMQpE+PicCiaWGACiKLC8vUUdLjVDEYaDtqpdaVLg71FX10hr25qxwhd2D6
/PIO7WIopyWrZE42vuow6kPDne48mIqmnNentFVXMU+BT6zBP5PbVq+lPxa9tobH
P3Lqc+oIBB0BFNHUrO2S9H1qayoJtY2xP4URc1szRjmzS2KjRj9T+SRxF3tjKRBt
3B0Sgm9jD+vVLHl/EQTGoyHYod2rTxgXnQTJzEScbeutnArOmAPWYiY+y7FTTyXv
fk9W+mvAhkUGO5eiOuRZ9Tq6WzY0uN+SE2Fno8En0t0qQBOC5+r/mueYBWlHQksG
QQBdAifHhQKVE18lwykDC2UZGZNDn5yCTgzIdTI71MWn5nqo0d3i9EssOPECR/QG
oH4/1evVBa9NO3x/tnItqRiTtg33CpmAeIpNvFfi97yZ+svX5OCf4cEEhN+q4FR7
FnPQ5Zy5clYd/iB+OgOztU2u/oL4AUaz5w7idKhzx99S5BVUdS7CdzjOFCpWghEY
QTxJr4nRhwBIZ6ROcRw1sleeLnidHx077Bk0zPtfSMr1L+GLlUg3KZsMCeqqF+kp
hc5HbbpXd4lUoDSTMA2wKBmXZHEtYntX6UHFIB28c7BO15VGaXxfC+1KDp0qnmuP
U0Ofibm7ukoJ3V6IiiMkM0t4w1YwAahak/kSouxDPDAukgRxR1Rzs/JkaTJkY2ZF
6HlDajlN0DbSKzbrDG9THH5Hwkk59g31+L8+c7gOsXM30+JfZtw8xoCILp7Mn5qQ
L7edUHFIVOx9o77NLwmcxEldhQi2he9ZSgMwSRra1W+WAIVXhH2js+hUAK5cHMIZ
BPFzTIZaUqabW2wGYKV0Dl7pm6+XKSgWAIDdu+joqO5bTxpYY+69BmDO+QyEMGh7
7sDv7qcUp9czyAjnx1u6dWujQ2fOSoq+uFjx7eVMmD2tXPS82piBWQ2w2pnT2sTF
aHOOKXy85qPsP3YxUEDPsh4FZvX7IfhtDqSZ7x5RgYmF7t8at95XlDSNh79fM8xE
i8izfbvNTocxPwuCu1sDsnKY0apX1DuCqvhuhiPVkzlUhWODw6/athhn3cqOWX8A
8xHAJMyFEwi0rVHtKYafqbiYpeFdJgb7ifMhmTsVVa+A/p9nY5llMH9HawSNSb0i
bo9oYKr27ENyuwBHGqSv4F1A2EtZNcFNrl6XKvMg47+XTdLJrtJPbtSavcFEuo0K
wL2ca9AIn3iQ4J06tWTs3lwqQDWHm6StfCEe4Ap538eaK/G9aeDMGFB7POFGFP3p
1OwsDp7Ur5QHDpFXwckKbWdFPprxRAdS9kX/kNUr9aMH4WQAwXIuojFXBYz2NA5B
mz8Vo1O2LHvpP52+zd2riZwYhAPEd7bkhWy1GNIC8t7nLGCDhXCG4op7komS70cQ
bbh1rrvYqCwFLcbuhFvmT8sojbjKAJew7yCnIdMBvRwHw1+GUsJYJHiLlDZuEGB8
T0B95iMXQqIaKEyTZRY3OCCss1mk3koDf2VoCn4kjU8hGZkBnCc12uHjuN9sCZlD
UKnFJjFqcYloaEEP/9uaLtbBLsEWz+aBfwPrRWWVNgkggovDh53UJ5r6S6c1IoXQ
4A+uUKrv3UT+NAIV0LE3emb3C4YPWXpmGvdP4Nyk2fcWcQk8DGTFWsp5X2S0PqP6
nFc/aRhUvQB3QlxvXz9ajduQEfrNz5rKLscLVMka+lSGVgK+iT2KQxU4NNXjgLCE
KmQNGQleD20nl0u84/gnQHv7yt7B51mb7A5dM3YiWXVBjtxM9bvxNlAD2gT3tQDa
lbVcWqZ1oaY7F8IEqpPFfwrUtgmV7lrw9gRuQ6K2GkgXMuzycsmzE2nbTfzfBl2p
dOMpOx1X69sa9Ma3tWhbPWYifw3OAkG73gyJeeZ54/0J8A+XP1z5jqsKyYlA0SAy
wGllZmjo6kQ4f9wbEXwX3bI7Dw8xSz1FOTh+PdTKb1IhJ5hZbyGFjQXQKDq3VZZ0
93D5Oq9IOLsxoljosyQXOZWwwisl/oy7s0gcBJoxFEuIQflz2yAOJqAWuBGmRxQk
RTKBRzaJ0e0rBBV+LNiG862bTxy9XnVqU9d8y+qNifFpbzgE1RhdvmRTOAaWKgJi
6B+cedwREtMnVui3xZ6YzVRDPM0sTC3P01+rTHKep3EGY02wi2cjGpymRNHylFRz
WTW3Qk2nPsB4dbCVD0y5wGNDfkbypHogLsCrT7VskDoOk29m6dV22DLQ1LC+A/qW
UIWF+aCT5+ybQOk/fxRyr1ux4Ex6zxS5WEmH+K2GGjJQGgLsPTjxxLGXNdY1b7cP
CrMQ7lsFnhoqEMmlWZ/8dreJ7Ccux1FWf/DH3S0pn4wN/9+ZnBp6AqGfxcLjmGIJ
il5sS68WhDXYzIwk51zP9IcKvt0VPFZ4OFBODAvzQhAIj1S1NMeUVufDiDlJt8+w
3gw4VZmO7zZlLpwqDI/sXURFMTY+LpgKiW/k9yC8O/ncBP+0OZ9XnuOVziDtDFSx
46YwV6fiE1uf/NSayN99GeflD8PIDXyHAiGPajMDnAKUDiHGRX6J+H0K7moVP6OD
TCz+DyRZRkgdKv7aDk1F+i8COHsw4Qs60kmwQgwrs4UkaSmUOljG2K7UJqfCBKjG
4j86wuqzWQ2Wf8VfM5KVPrYErzULMQs2hbGhncdNS8GjQFOh9cwTb6w8+E4OQCJt
sD822YK5PiA+rPcoPOw/1gwppmIswWhv0jQCr5Bfp224VaMf06NTDWW3QgJfOS/C
VHt+1hLznUBiZXLTLxtLgxDYwuQ8NnPyofWLs0++mlAKK0SUNWv16ODy7clmrANS
lgCnSk+trXdCa/rlL85Ty/OC3kshLz1ASAz2cPbV814CKKT4d3QWxmRUenX1lN7s
K2zhFGXihFs5n/iDww19qNGcNJYMrW/6+HSe09oCaFHeI4K/ZeYOngiSujjZ1Hnu
OURivQjLp3PRQPbTRgjlZRJd4TVDd2+SMoTatOtoCM19zZAJY3AHXWMA3tTKWmNV
anCvbsggBHublu9/SqfKVicHISt0SS0W2tk0gaI5kQ9lO4cYH4Ff7YHhORnpN9WI
euQ649lbSGub3k/ALeLkBNqQSQRXHahzUr9xMtry0/yQTK0A9eORUz3T3GuPy7jh
ZvNkZZK35p4f19fxzdyWFXJcY8X8zcf1HjPavhMs7JkZDQmr6OiGpUHydIVnJFQn
UHYBoYawv4w0U6rce8sBuL2DszFOJPnJJhnGM79K7To5vD56zS1uD3UdketJyXnq
SG2OaeBlion5m8gLhiDVPHlBZwyDLl0djFadINgFmlIUM5MXzd/SiQkklSVBJA2/
Dy6+QytngAX6kT11Wusl+gWx114kCRwhnEkiQ2eflvicg7PEkTN6ZigwHijRsow0
oIXzaI3mxgBz6+TmDvYS6lCYgYUfBzIvJOyyDOcdJ9QI+dvtYEGRjBMHo3K5uimK
GXaIxA41HCIJbnOnFP0YnsOa4ImWrmuS5wxp2RSh2XdDGPhQj7kqRen48iPyt1C0
dZjGSsGtxCR2141Yim00vOHdoTMG/9llwqNgJtBq81XykUrN+LUnAm+6GfmNoh6m
YAI2qxQheyBK0nSHUqrC/wD5wbFBbDXbZyxjlpD8TTe0PFuWtOsidjd7kKdNgamN
5cEPQMto76nibFGOtVlZNaJxzKZdlMuB9kFVUlvVqQc8hz4uezuzJjEMYCkmkBxV
Ao74QygV6BJc8w00mPVVDoK39gc2dN6Tm4F12O2wwyTtrdwlha8DfJ8CWsRCiqr2
Hm6ypqAfP3w+FknfvWnORbhex27h5jLJI/OZWvHxw0xqQA9bl2LyvTkA7M4hdV85
CMIQnXRIYZYkYh27VQbv9568OQjqunsQdYAoQoZeW4iYKavIGZ4uoleArFOYUBcs
oNyjoHpXJ2sXV2D6/yjcTLXKfIU2J45SHmtJayL3x/yVeT311YjRWCIrTpZ5jhB/
1QxAIQzdFcufGfSX57IT1VFkPqAk0KEhxXySzhI0iD/WcQiQHI6OGCoVje5JqQNU
Y2prC8Dcd7eyiANKqvptUCTTMkk3uPHJnzUOAXAuZK/CW37bXjJm9+d0wGUi6cvh
TETBDOt6JRHz0mGw1mljYaXULouirjf0VW+oAjL0o3j4vjw2h1mOfTpNJl7E02jl
tL5m1Qa8bSzN+bRhay2EgOMX/Q8p/e3IaU0kwlyg8cH2qjcHd3NOu++O0LRur7/w
/GgiwcVYooiE43Ri2pa9HP3hfDEMs7Vg+ypXRheYo4e3zYagwOPj6Ign3UG6mlaj
4FkjLSmMKPAxJiZvckluRD2OlpXUzBxYRnOMXs6ciaoXN3sdzBBn37KZPskTw0B9
jgvQib8lkIxt77YsYmbAHKVwrPm1CU1bf6lpiIiHy7tIBMdVjFsgwuyFz091fVG2
SeWNR6jFwJMvlSUogkFk7QYM3rhMsvoVJl/E4bzjpBT06SVdTHKVoI0omy5frIZc
B1p1Fz6ayfFSNyo8mcHBK3R+BsRxWc3Gn/dxC8eeAgE5Lx7XcFo0WBatNhxpot5u
ZnD8M/J86HNgTOKx6fgiWrrGGJy3bkmWK9BO3uk4Z3MbMEBXv05xgz14C62k5JQG
ery3v6nKUtTb/1mGV1gdyC4nWmvOlCxq3S/cCcMj/g7I0kqNJX3aCQ2MqP6Vz+mm
X4Q2hHVejpoetTyMocYgPxtyagwGJTCYapMRDZf7916zDM7maQjovnajTJ+yl9k6
Ur+3b5iA0E2b51cAXGF4ny7V0n/bozt+OxAu4SDLqFvOX9TPEl/UgbHtowz9qyCr
f989zRimmvo9r+0swlbPkLZxIMjPtMXeHLeVkxRHHt6Cefa1s5ClPxupnZ5YCmw4
ozvDi5oWp2Fe2RWLEndHrisdSiVnPRrz7y86zt5k4Q5QE6Fy/ZEOaOUs4Uwj0f+0
RduY+2YBUMOGrK+vwROkyztShGRfqEukJMTFbRLF0Jf7nK7/4yPxMA0MtqemqRTa
r4qWbdvAsOUyDjrZ9PXwsWkp9KdrecUIeo73IksnFJolwfWHtMfUqhEAYr2P8tkJ
dmM+NkAg7B6aeqOoke43Zy0EjYVPv9JHWns5kIiryqw2Phzt1Fu9+zu52RC2h2ny
6R+ywdNg462Hu7z09r7OQ85Hbbd8a/G7UZYIyt7/Y4y0qMRRPFsF5nfbnci8BLuU
m+MQ4qtKEB9b7vz0Cf3BHXav0BGz7jk4y/1iVDzJeGURzQfgFH8A+GU1gx/rtoCS
ym+3ZHGHXoJ1FBNveWbblSdSzGFoXwJm2silniq3GLQ7Sty6zl6emLyFg0vBcqFV
OoIaVJ9EiBJ9GGH635ME3VaYakoAb2qkAaMa0LLqQK8YfySkCgCRHGTX9rpdxL4s
F51xIFEjjtpAl8W/VhJKc+debzur90aAePDlIbX/e/uXl4xJnCiO8abh1BbX5avU
sV63MFBGgMpjAeT+nrr0r63aonW4SI7+RT/ZQmDe8+FzVsKJveyTjE9QTP+eBCkI
3SB+w2V3yjjV/SZUMsF1SSFApAIC0JGJE1SnL9djIbLi1vPSsi/9cVd21LycGSjg
LWoWNtAGbAI92ku/SnepleWv9paeCItFjzS2zxKjWV1eBBLtaV3VGvKWt7IL56/2
bK7wDkxKET9SXycyoruLws3bk50lY7wsFWtImpkCK2lPJBmtnJzkrSzLytY8SdmP
fCBZvEnqezpY+gRmikxWbMyrm6LEUFwK+4rjOneeMPeRm112AAaZU30TESVcBFx8
mdN13yYvX1E+9gbFj1t9wHAJ5lW1alzVjGk7OllMUEq5WVpritCmCso7DUVGqBUS
oME22YwGQQh9GqSJ22Rri5JLQO5Eg+YmlhE+yMoOl6wg5LwNXYv/ovbpjTqo05sI
FtKRBpdvtF4EL2mKduWVjtdLSWOoU0TjdqmFQyO7iWEZ/Yhy7YLF7DBuW0B43A2b
U/ZGY4+1q7hCjCm+kHIOIxHwjEIb3IyVrOf/S88RpE19q4vgwp4VlOSJFjmFUwDf
IEMIElfc9U1uKchdM05nIMCdHcTHrg35sv01XaV+KNp9mxC2+i5lmpQKn0SpyHJk
WluEVpcsIS3Vr//4hZSM8ZnCwnc/u3d9tyQJEHAiwaXRN1J2dg48f+VC3M1tfhKp
TA2JRKwcy6mOMStMDljJ9ksG6OpTJSHtQkKWG/AxZecYm3fGjnIZnb6rubtwP4va
78Qo4FBWUEZAs9smYH4C4vZ8mcabfQl83V8ZuvDNYuksN9SBnUwMgv/l8P9mMvpJ
zIHWjGLzjLIw+Ykb+P7rDmTawHvHbHsErC1P3olDZQJUTHWQzEzDbb9I85AIfIhL
Q88sSiKzLLVxgAEZB4RdXiD2bFADYob5dWIJuMr0VTDXrYUbiU8y9UVX45ISYoL+
5KSC+h23AufWmmazhrEHVVMsFIIUGJkh+yS6+51rQJ2k2lPrMpfTL6CtEi5LWCT3
POAHjmbPBndmPZhohLdAPQic7Eepf1HIBT1YEgVkGxv+078A2c7a5OKcu3wGzmjY
/Q0azSRDzYJ1QdJuFJCRqqW2ScW6HXexMsYFDkeLRO156jnqVHFj7rK5HXKsptXd
m547xvqeAOjebsL7n9m0uiTDm/Pr9KAJuERDvPV7xlBCseS7ccMW6N5Ts4bt3CCz
7ki/W9XjihrxriRfQTATecQIYLDJUoR8IPs1rHqrvdnbvG9bkhIT3OJ+geemVdhu
RxzsVo3B0CQ5oVWsSWL6+WPdoYrm4qvT1FdDA6CgOEETueIjXKyc6Qvqsgq7aMQN
U/Tc2kTho1q6QSmN1J+1F2EDK9BUM6VVPigRMrAHTzEoIf/vNs/8GiLhosn/xOcL
G341Qwasbj0KoMU3TmRQuzseu57RHaJgosczz6ufMw0pNpGYoMazufDtd66octjF
w4EsbNsDU8qDHiAiiV0w8M9o2AO4a9WyCzBYzRC9gW7ui7wIRk6XhwwY0XyemLbc
hhiEYzT+DMVgEttyNcjxUc6q2AFbQzvixa+0TMKPorwkyl6CPE7aLR1ARpF3qsT0
64FpkMw9VzWEhT0kaNAKvQ==
`protect END_PROTECTED
