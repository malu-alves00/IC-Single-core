`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XmT5MfK+EFncV9HvOzlrygTX5pCUTJoE2IJXGN7cZXZAz8kNb4h1/Faar9NRzgTy
eH7bBBa2iljw9FcZpJgq7FdaFd9i2ELF2u2v8Zb+QHjeTshl2ALpLEgpkOXuMyRj
QMb1ULoPlMM0hIKyg14JZdjnkddLDqFpPXYkl2q/rNTs2sXnvdKleqw+TxJ4wBmI
fQGnlGKqr/b2fdnszthWfb8gAFkKYNOwgfoYbfBjCLLg5lNyVcZG40KzTQX3ox98
aLxQN7+ko3Dgp+BuDGUAICDTRKQe+VDmQTphy/3p2wcF3QdBcL5TkYHEbIFRFqZV
9TdEzt51CmcYd0J53CKwF5UCyqC2BPZfrOztCq8Unq8jeOMcZr0WGMduW00j+JLz
sQZrKPmYi+tCeInM71tPnIVknIF4Ap4IjotiUW66V/jpAGXYrVwXR/BOQsQrL7IF
aekDAq0lRCsMG6K5IeVaeIHFswnfaO0II+NkmW9vvMHo8AsnSwbkEl/IcUtAZ5pW
squNTuYPMO160lOxk0Tf1b0MzIEqROEPirTBBgBPNHdqWxF3VMUpckAmc1zUNg2v
wqZdcedLQSZvBIV06UpLF6AcwueDQgRbejhPLqKNvR12WxlCIh9ktFUcBhQW3Z9g
rr+iymYWAJ9MSTeJrSS69jlLIG1/ttdwntZ5SnwYEfUuhh/mklVs29B3prtGZ4VO
/iKtPJjcp9rCsOOnCTeagtl556TVntIw3/6OpVJvovp9MJjOs4+Ld0e/ap9JsQvQ
taI5czdV8Ru1f4tXl+EGzj5MHvHPune99A5lw4yEYZIMHofn4ChW6XjT5N5wbrNM
cOiwSE5YTvpRcBzCa9pRWVXbEx5xIHz/QX+Gv0AeFFSUpREhGMLNKYOqglkbAFXk
RmKfvGQ8vydpaOoBtb3dwPzqlg7G9kC8r9H3EANyLFsyizkh3DsDq3JajmpWz78N
EsUWqXHqDwNQ0olAhJWUhLwj8pgCMsOMrRMESR9lWsWk/klGwEw6QGD2DqptIaSE
kkZ5hweA0pDOe7BJSwpyakM0BZeza2/zJ5Qv+qwED+vqpq+9fBHSgopXzKlOa/ye
9S2JLFxNf+jFU+EbekPyZ5IPA6AVLbUvLiYN1OXe0nHcrGFmluP2u8tKgDyruVIA
3suHpLofKgNUjonDNoqvumJOQfy63gIvudZKSTUrWFHaXzkwuOjiwLxBQ5KMI4wq
1eWLtb09BJeKN2UV4f+tjePkTzHNw+7wgZraSbNy2YqiC5CGrWJ9IQKfm+1pAGkk
onVTKIbdxXkpnIrIfpOYdL/qgknxxM3yjcNDjV5U6MHSTiZiEBPfQ4UemezJKSOo
`protect END_PROTECTED
