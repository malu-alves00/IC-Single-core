`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xpVHX+MSEqFyCj3PW5Rjp/jkp8ePeIne5Cqvu7+httx2FEz/Yo1bv4qkotI1TQ3c
iq32yivn3SOH+/Vb58I4w9wxdkOoZsrr3WQyZtVB4JxbhW3bXlwDzPqL4Oyk9jhd
qqe/h9WxL5KTPrnOyZMaXq+wgPFrWo+KBnWykCTIHUdcYZNbO5qbILHHZN0pp69v
2lfrgpZOZrYu9S1wn8YS+AwpSHYELpSYqCytwvrUUUDsGXJnNvk/d/ZhYJwBDCz+
aYlkHYVG2KSDdk5EgQbxeCUPOzzHORoWWA0vMTHcEvL/v12jxeL9lPjhIeuHWuEd
UnZ/OJXZIwEOGExZcyelfS6jSMzmjTjRbe1x1fPeyostMBRJOB6r7R4rEtDb8V/w
pt/ldJ8e4rvDp9CVdrr+Zz68mZD2rmq/4xfK5G0bHntz28qcqJM3vrpO36npHzH2
W/iH7G8DX7n2iooqI+dI8q9zXzi6iYZJ84suS/yRXJUnTj2BuPj8FCKO275UOvZ6
ys+Q+H2r5/kuk6oferVxIrjrJKzKPYWRnnxZg6PXWy+yiNtW8mOVgNeLwnMV7R+u
TklwOic7x/JPaITxR4orG39mksFrzUVfbB4Qu6licOXMNO0+M4G5P6iHAj8TScti
Szo3DyqKD3M5mq9elaRtaXyz/MxxPNtfSVHWzv64Wt7ggHNmYLCB2ZUjwV/SM9Gh
WseekqAw/LqF17s8GIfKqRPwfyV2GfpjFXgdXMUOEuqlNsWtmqe0V6IWsRRYjAeJ
Lf155FOIUDDrZYy7pn/CwNskr1Yf4NbbUCEMch9Uq0CD6YJFoNWLtUKbNeyAAwZO
YJSWkwlJI1Ptr4pjoZDzKDBBKhaVm+XV57f0e2ZrHTC2EU/P0vNt7VVbGuxFZ4hq
CBetZpl9TI9Z9h2W+PNp+ZpSB+KTJf7HAtO4g8hy8qI8VAKjrpMpQdkiWtEHMPWX
v+sPU6FyqSIPxhb20Ulm60Wr5W49Rd2N2GNLOnP+iALDFtVZlB4m99DYuPtDimtJ
MO8B9rXH4KytE0awWubzDC6ppcWVSig0ao8F0jTK2Fm/9sQm7HBWLdjdQS/5+AxU
A9sO0EKsoTeNQ7dbRuT+fkTLOlm832xlBSwSQhhgg1ATqRoRaS98YR/tz6ABcZ72
tTZi8gQ+aIdAuJGuj+oy9XA8Lbo5xmPRHi3Gb2wVZ0VYCcRxG7bCbx7U0Zzpy40O
wqG2p28j9DjnT0sN0sNzsqpYPLEB7frgfqK83u03cjjjakJMmsKFLrd419SLe27w
lDbaqSl8FUnx+rwvZlPmNGjY5k/awD6rdCH0kJKgMNb8FGoGW/xF0ezjPpNdrZKf
7Ju9vQvqAAJ0n6Fq5FVG6r2T9K0S/nmNBmSlaeUHUG8+pGKmGH9Eet1JnrVIw6Po
ocYQceGtB7AtWZPAp25IsEUZV1ASpD2Pvl+wzEbLZzimMZuYE1hSy9R8e09THwaM
n5HDEucH6CLY1mFASuSFPuwuQcx2AxzNvGvLM6giW24mY5omxYNGjgmSfJwcQrpB
lW+HZUVQh2xVFQ61pOs8lOtga/AdDeN4+UtKtTzr0+JOjSmK4r26iYcDpBvTxFK/
bNZStqMFIvqBYQI+uYeOJTvCzyXeD3sAYG3tUGF9Rf9+hQkNJHgSdHb08xwbhTmc
Kap9xo0cwm5DZ3m0fTBPLRbByIPDNPWEygC6M0iqzQcbqG3KU4JdLsfiPpEiyGwT
MCoXLGMvHITaEWOGjBjX907pCwDwYVVZAS++8bq0Wxk6kXeew0la/wofJY1BDgE/
qSna0YTh9AuHTFcJwRDV0foyev6jml+95Uq1qrQBEqv8qzAqnXWEWUjuegRvPi8i
8NSOLnHiUe1JKp6e/Am7jQ==
`protect END_PROTECTED
