`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UOW/Jq2bIscjV5gkUN+52kmxUm5drWrwPYarAlKMRf3n3mEOWHx+qZHgxgZiaHsc
ptb/3QFizcCnQNx1l1MtygVM805oDY31jU4tVvWF72UqlU75tedExGxbtKOhybdp
tZNYMobM1yFy7t4GAbrp2GaPJYKp/kegcjF/3zDfPG1wAfhvqSFBsqTOeI/oRxNU
RgJ8U0M5+IKPYbQoJ+kYHh/EX9ZJ5zuQBo2SyDy68GjUyZjMdqOhjSrbWax0QPlw
xAAMYAYZH59NP7Y9hbllQxw+NNr1sBmouNX8JXMEekBwLS80NiKzfYEu2afW/GWn
Pm/0PNS9SEkydr9Usxm4hppTOnFzsJT8PyRBerHgtbOHy2XcvK6DaJPG753bqIir
GfxAkyb95kIIQjt/U7OAFOmZW9TvvpQEa6suuXfY/yTH9ONFmis78tZPef64nWtG
ugwm1NxrlOMvLyYGaC9NtDSghqmQckflGBAU6ueMgrPR38S2dXine/geQtjh834r
XE1X+LKUdKG61N+NceIxPB7YHDRYskAwqRx5LH+b7L4iGle0i0nK0JdzgC3Aa7kL
sDNLfMiXg53OSrEhNQQZ1aMO3iksww4AV4n/phA7qVaa3i1TuJhF6Quy6rIejcuq
anFpnF65dmSrtRGJIyK00a6CWLQ5aX+BbTyO9bokqHS0f0zi4Ab9OvjF0cQCQsLj
5wOVJQtphLBtiJDYg4uQpJp8vByNqvafDGfR1CfzoYJ2p7ApA4WTMpmlZ84sUfzE
OHslZblFo5SNw377T6Ahv1ud7EIHAMLSexhxPIGyqVMFZjTgt+zfwcrzEE+lczCj
HHvIwAp83IYvU/ixItTLoWWHZ9gf9subVQhHO0V4WmdXk4SoYy5eWXrNzTTAqKUF
RPD04oijqKkNt8+/iZcZklrKO9WP/vOfQSKUW+hkN+DUliR3gD49h/Q4SJXGXBgn
TtsTcGMhcC4AXY1VR5O9fDGMP/TkFmLRUM7vyldqjFJO0nTyxZyzLPkJJEP6bzWc
DnywMJBOfDLccksc2/8LlHoMbJGBa9u+RQMUyDKgwqlWH7EpmpKL9qyHMQ4G4Bl7
/Y2qI29rppJ0Q4BHozq+8HYMjfam0RS0BPclbsNeLzoxeMvOSJ8Wn9Ug4FCmMjMA
9Bkeg/xIyctBPZg8z72wpw19xxpFWePV7de3gNG84LWI4HDY2TqgC+sHfq5MHtMf
uncZcd9mYw2jzZ6/t6Xgl4jQiSATfRuvId85nJaHjBsaxYXshOye144k3CPdtxSE
xkhYrch2nDhXHjiMscpvrqkjI1+aCOq39Q5rk047ZW0uMjGSqZICNN5v7GFwDVyN
IdCly9heqkW4Sr8RfH23xN+3Sd5ntD3ojJ7x1zW7cjjGu6qG0L1mhysiuLrvZHdK
SY5RMKOtn0U+p0EYdyBVRetOy1gGGXv2oLYlkuZPHD8PEJ29zMUcZ9YFPCY7FsLm
jjTfH4/MVRbFrSdZnxIMgps1wWGUT1abg+KmZudCrHofdPm4twvgfDueZRO/6lq2
HqslRARUCl/G97zCtPXVqpIXGqQ9FQE0HVUY6mX5TMf/6frnqLLBIxbea6el62cR
hIJM/UH6X9xG6h8JFeBQAoDjFM0OeUuMwbV8YMZOrWxAikcA8dn3iO6qgIWEMx75
vh3TGtooNy2ilt0QNQfOCTtPlICpOMBlG/NJyuAiJlDZB8sMS0I7Y44SQiusqKrp
epYwFuSivKf+VdP+yC5DT1mwm4FAaH7oeoWti+7aj1A0C1NeenGT4iPmDhlt5PvZ
J19Oh81L5AM1g/FSTP6caznL7O/nYb5DXV1oZ/Y4NLocMQbn0qpHvtYFaWBnOUS7
Puu9aHiv7P9d3L1NuUEHcyED5lkbplqn1keu4HdmrCEWexKkOdvv/+Lc9hzfjrjf
JTPOSD178cQQ981Ri+purkfTm6ZYQHYZiPntnIsWX/qllEQyfykWfwJ3LSpP8X8L
sqm06AmHHDJTtEkAiITdw0oLRmNvpkU+E32xRwlneucVuUvD4JAqRF33I422untC
T8a73MZKpWXopogQWha1ObPUUiNRMaumaa4Uwfz5m58dPIaqOwGCESlv8PHpywo8
`protect END_PROTECTED
