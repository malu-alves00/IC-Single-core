`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RRjNkFCQsLxmvwOox42Bt81hJ1NTl7pBk4OcFK1TtneUo/oAgFxChQsmxefrAU76
Aynxpf8yF4QnqlCK/4SLueKT5R5TWtiSsoVOYlw6dJ0O/u81Ek3td2nQN2mFPlzR
nFpFMOuqSMTH78JrJxK6DK8re3e0dIlxnjvNplRW1BHnW5d7yYNhV8BHRSTKBezU
URkbTf0tui+S3ioOkXEUhYLq0uOXAvQT+Z6K2Jcz9y+BdtJuOUGFQCM7kVDHo66f
FLmZ6T8dfoBhhrPHZBWAVi12P6jssI+tKU0BgnW3GrXg2kJn8UXENoR4/WAKNRwV
z86korS27UYyBiS1zGAiL3uLnlcoNvrzmGeibPwY8k7+2Yl5DItvljDIXx1tcMra
3YGxXTN+eE4EWPs98MtC2+ll/hmDn8Q+Nz+TNcq7nYZD8ZNooGyI/mB0zmuNA/n5
kbTBs0CezGuoNmWA9mm+4O7ElD8Pl2hlTBPGQ/rbQ3gd2KJMxd8bLa07++t8X2MP
anDYXiZb+HcRB5aHJ1xHJWOvXzrRXoks6DRfQG7x+X8TJ2wJ70QJOPeUrR8Jl175
3+gvR53WEhs+BxSiYk3eRZUoL7WW66PC1xynWXkheDmmMHMGrtJJmj4JJHkNgBH0
Y7Iie8Qoqr9R9esezfbMlE/mV2JPVJ1BtwYQDJnr0rg32HqQi0Q89rprHzGdnWKM
HggCejizq8u93+wNhbcOBMbwBTezmFyNicTlckGOWGFj9VoVdEdygNimZ6/DbXKI
jbi1iw2DQjSwUPvoqQMRmy3Sah1yKJo+FPtWpmtySnvYznqEjpeD0T1AtLtkJ6lP
6qv1KNEGmpBZ6o8NYAJlAtqWe6t7ObdPhlTMrryaTNxX9hqVSPzLXC3YjMstgj9q
ISjNJEo4Eni5gMUUhHOV2srsiZKN12r4AJ33tpxC9L8moUi64uuF3tDFu0kt06JE
+h97xLNcfEKpGVtMaaChPw==
`protect END_PROTECTED
