`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fG9HpaHwppX76RPVULE97J4kibezlFw32cAMOu4kmr8c4hJRguBGx0kA4Uae+Jar
/tCI3wDTdKEDzJno1l36qPITCXpdCEv2gLMqtN2PRjKIKen6+8kcit371sLd4gZ8
gXqrENmodH1bZfr3T+QS5Hp9aOO5wErr1jvhS4MnzFUyBDIuMymJ+UoNlMf565Dm
gwfWc3gOT4pj7gsyWQ46hiBb7Rof6UfVEKndN/xjyinGZH1P/mTYg9PuuTro8eTl
6GQMhzbbIQXQwA7IX3RqXTI5DRr1wk6BIO8YlqIsNfbprdCnKKyduKsO4cUYRoWJ
+olIdWNMwA2fs9tVScIwP8mYudnzLqDzCH7c3PP9dj+MHM8Llp0WVniFIELEJW77
zry6/HvG87JxYbNgKUOUjasOahbVJdClh6tYhECFIDxaijzi5cvxuG2aoKdFFzHa
chunfOuSRgiL9I2zqKd5/Zpw6CYz0jw/kBguk8gQhaebcWWKqO4Eojs+9vIQsJP2
`protect END_PROTECTED
