`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RSSvwyQHlNcmR8PreF/x8tO4aTK24A/fB1QCHXa6L8i2lCWCbCE6zcN4ACx8d3nc
7wbqlxTWIroFrpizwWbq51VOwCqknXm8O1LAZXhnSam32cSxD8QH+RLPjflB98nd
KcSlQH5WYhvPguPtehgNITOpoI7ISAOenFzonZRkvkKb+FPm8PGALFTjKcDPG1FO
D2mVdyep642tmoaYo+C9OLPDWfvLBwIHJEqKo5pIpMvrfe7aoWY8ORDvhkUIr2FK
rXHz08qpz0EpVjFqlazhcB93t4aT+ZCYweKttdm7+50wYCpvnfGr0kRwt1WVNufS
NA1hnBt/5PxQXMLppNhCPJfTbCxLaTusXo1jw2w0jc7JpDJxV2YzhEcmi65g/aRV
QgpwYN/n3EynRp99opGma+j22QyKtBoJEMXSxYLmBBCljd7JC3TRik/437kmppGf
AYx0AsgeN0Bacn+Vy0AW1HTRDiGeAB3MkKYjlPZ7ii4goypjtP+9rQ2UoV+FmzCz
Wb0lxe/RePZE7/zRJEzjF3AERiaPQxUIfZ9N6uCfajtBQ5rlt/KBPe1jsjWoKRUo
+2vnycl7kHshIxAU/5xWxBACOQxOhzNgZBxdEBQLahu94JrovaktlRTly0NGZKjw
ePYoH7qUc0tQYVkca2XHIkjX4eRyMFBnfWDNe8H1BTmysyvIHIH+oq8s6sLd/v9B
eKgDVm88pnjtlfSJquhVMNABLAYK6kjynkr5KhTCtDM8/IT/dWlTtCbG7ND32uv4
9BHq6zzHGXPjEvvm1x4VcLdH3j4gHAAcp5np37CE7rCBVWxFBA8tuOMTVP7t54Ei
XvjcfOI1WdHDy+M6mP1QX/eDXRT6zjyABaIaOFhNZvt2jPMoWfYRweNnaRHNLyEB
erCGyV2TLq9Goazk9IY00izBnGgwLGe52jlicw5GDaFrIFdc/secO4qIX9HkDPSD
NZWNeLG88vt2EE0ttNDwkGMd06QLab5VL7QBwq69TpOKKaGmTdpmS8Tqp07889Y1
cRKiqDIY7WRQq7VuTLNtAdA/MF6XVgF9ZLr414zNS6ZAC1Mqtjy8N8eXWA5Esk1W
hAqja0dQHgAwiCJ8MP7DEe8oakmln/eb6IMf/7zy6aeX73OdBG0GM9LMKkGf8RBY
+TCGzY26LXMN0iGstEO1xDvRAfcSO78/XZ73kf9ZmjA4xyJwDMqXVuBleNpNVgMT
6R/ThkkM5aDvK9jkiFR7Z3Wu9tPadi+UiVblzpkWFPTlFGCrTobHhz+IgRI7k0A5
8evypVau94WmXOjVtXNYeJNZfovieyPdYSYExumO1G2MJz4hmHmS1y1L4agaCJDt
aIOxkhH+2WXsa0meqikb9CJBWKXHA24KW7XGq23hbhK1zQhwdqwa0I/MdGc/FM6H
XorWe9Y8VV+xCsP7fQKWJd5PRMmXECj65SCnCl61eLZiSwAo7nNOZ70wXP1H0Wfh
6nCy4RaRbGRdxNa2xsyBHlZ8gcDJ9Ay0tD6SkReyOJMVovm3qM5q7MPAEAbiHqwa
HIx9NlxZfgiLXc7PoAx7B9m3EIM40y/OQQ1kw5Z908w3OQdpgC9MQBD3KFx/nclJ
YarQD6jsiVPmomJMXelG2JluEAH0m+sL8KkOdjWig8Upq/B+nNCQalGTiK7SuIQe
THfCchCufoGhmUiD3eFB60/lrGlbFKhwFf9P7AXrkAXAH+YBUWa2Qtohq8mjceIp
AFfdYYsxE3XmSrFEp2JSvIMwFuncxjscSuc4+TczvZQ=
`protect END_PROTECTED
