`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0F9yXZanmU5FcWli3R2Y4MrRJpqf6Y7uThRLfUM6vCbFZ41R34UfGEn9yzezvApk
D0Co6Qk4Fpk4yOw4SPGEoixgyQckY/PP+ksgtbXdjIixP+WuiyR9hM7Pbw1fiNPj
z72w/OXvzwqYVZHbfMfn/4Wrv41oI+xoTyZODvVOKLdzFf2sPyQx5f53y4pozKs3
JRtEa8kgxLP6OPL+cRRDj7Lrl7iiHGsNYqomy4kwmF7pdrt9gKi37Lsl4Yv7a4Bs
7hcGB8P7IgMONyZAXupOyuiHLAVdJuvRXLo5hswtNO5co0j6p1Kp37k2EnUep0jR
hDelGkAOb3H5Qf5dVjSgLy4Ln544sTvQLWq9W2BqRhT1YoP1Dg4I+xuijE5B+QKA
vJr2JRGiFVSdZAoZGpZ1XSWRpNYd2lKjyin5YKbgTa12+osXuPcrRh01W6VcjrpU
nrQ396xtypgi4pIFPr7GCLiyai5zHf0UKcQkW0Aac37LC5bLyjUI6Z49irhmL+E2
5yEyB7wD67nYE6+KhfkPEDYeba2AXnv8T3gP3obK1PAPL9S+8fePTv6y/dlkhbP2
riON86uCHc18wjbi6LtbGx9NYY5UK0U/8MlPGX5ZkP0X16kV7lE9TupQR19re9P/
rmfSu21KUvAzxZYmF512kdKfEX4S2AVZc4Bt1CJpa5RBGWkTd0cegkmGB2nDUx0Q
ohKOHxzm9tkehbJmh84Wf8hykiMjUafraT57ZPwVR2cYS5jsiBytWVBkSugOdH5g
inuwkMqqUYtEhi8rnC81IPm+PO20Mc6V5nQp6o0nUqltAJWs3MNNDNUIXNV5JHAU
LAwUsI9fKbkT2ZNE2UxLN/Vx+aiNXItz+8+JFOTEGiQ2RuBPukacejNy4MDHGt8n
hzqqyekub0ZEEGn/kqOf7A+eyDd8BOldfny/hjFGEIjpoi3O5fV9r4TsknrmVZLu
LhP7mHnvnzgQ0ahtA8TWt2e3PCftIHlG+/NykQ96dJkVS7Ix4vlciOuVwA5YMkNQ
TPbt9LmzhILzyvf9mtjq3NxObOE63fKhXquwSYGWigqA8lKvSOFnDWM0+oZYhcJX
9KlkwyQHsV/ACMOiZFL5IQHrPce5cu89BpjP5F7XHsEXLT4kki5ZjKGwZ291OYCg
XOGfm/dH9y/7UJIgQNhxh1lrKZIVsSkQIc0x75mpuIx1oVtOfUHy0pHE7alE92Y5
NL3vJOfmVVxFFyuT1VN641AlgnEjWkvYlBDrGRcfXBaew1yWDyrvcIlHg/1c2zyM
PppQH3w94T/AYk1OJamqqD8ltlaS+e4g41KY2dbj39xclh4PF8ItsTJcDFwchcyV
7qk64H04z2APamRvTKsG7AHlfkmLcCsUiG6AwaIsruHEBOD0ij4hIPzObw96wg9A
2n4xqSjEMjAe41b1d8FwjeQQLhBl28BuLrjh9ftughVos84PbLUKBHMwszA+nXXS
UPYNKhAhWDIHtlaH4SDW9UOG4tl1WDJIb3aLp8mUWaDMhk1GUJfLThqWAK/oJllP
ktfQ+SLeX0YEXxNRHpa/EEhYM9ulvASoGZUxm6zMGky8f5EGlY+GcYMHNpCziNn1
OOA10B9YfYmvsnYpam7Fz+p1aVJwflYSP7nDGtJaz+vzmyJ9zbhC7rm80LwFJqVh
HSIFnFG+GqUAh0xAeCoKjOIVxyONphYSHUSc/sQRaW/ffv+VKuKcH0l9IX7sfWY6
g+UTeOXL7s+EQJPArqoVzjhAFPBJnYgUlXmLy51WWt/44AFXn6OMk7axLh7quKch
G9PRb5eZ3vfCbwZn/IwRnh2VGPaOlnEh3JsiEP0O7lUjx0w/OME8Ot5QRlskOqR+
47GqlAcfPMP+J/iEJ7D6Oz6apI9CwRhUpx+/WanNUbC1nNAYXO6Ad7vnNr2BL+Z0
JxODmoahOFszECE7hBHrMR6mmolNRDsRyIRIKKclkVOa9uEhLiYgaYJBRrjexMwF
JHVW4KTBJiu1GBUlBiaj30/C3YORePhlzNf6v6IGEZHgFM/1CqSCFtwZ+LqAzyCm
H703+3cleEw6IpVNKb4/QpyR4YVdz0FQ8FwHuaX7yrhhMIGlVSocm17J+MZ0BI4B
XoELFC+kr3WVHartB9yCeXv1fLIy10XemsfoB5YNU6ZC3WI2mXlnbtxRQlPgd1b+
8ETKI9Yx5hBTtK/AtObeVauIltgaNYVbkdmHzF2uc9ogf57pC3ftK9CDZdWSCNTC
WiwnWHMnFTa4H0xh/ry9zpJZ6C7ceMvfMKiC1TjhN52I6dq9Gi+UnbLUNLKStCKs
xTLh47h0SznPr8sVeLFJaoUtc+kvQVsAD8TGpeQ/zwEpNxGAkHlCgEWfJz5rO+dS
VhnP4WkNDrgRd6sth2Z8Wj3UPh0cklc8gsCXSUguQvjo6tdbA3rEPHiT3Hp/kiZe
K2lCAzsjWICnixpFgiMbsBxKizHRescUsBV0/ZiebVQjKW7ZiB1SKB8XKnmEX7df
B5ggntefCTIVF/iOySCWbC9ouvVQQU0mkVV3SnNVzFK3Lv8XObQ3q5ZbusYAYwwM
TSb4YYptKi9RiqzDRqjfiy1zos+WEvyTtOL1jOFuFC3IhKL/cFKI+JyMopXsV6D5
vo4IpcY//pUzOW4OqWRz3lT0kv9u/too+AtbWfcCgA4l/lH5s0ZAUn6XldvLfq6Z
Qx6Fr75QAmzhIkHIg19jiid1ukUIny94E+0vSF1+7kHv3y4NLVZqPmsYvQb1iT5r
jQt+yHUY3WEwqmnX5WolDLMOF5Aw0a50+ODd8QqJc9vsnmZZ6IzkOykmUoclE1ww
sRBfv5K1Herjr28CvTdihjiwIyZIop23PTkxL2wubIQ2/iJ1yh4m/LVrQ1U+jZ8+
gEYVgB9TEt7G8YjIbEqKMiXTRzJjdBuyw4LVsKpdwcEfH1F0Ypr71FZCX1DjndkI
YiP6hVT5p2wsclONZKBi8u6L3kqmH+P0Ws9foxl8/KmtywF6DJVQNbW0fAUpeq7v
Xzp91jsuQyBgz6FO1cJQPhS+CsxAA4zxIr38xDtm43omj8hKcmMW633HKpLpyTgg
UYMKuKRlgCmBVI69Hep6OVUQHHxkFWMJwCNsr1Hphza7Tl8RRmWXvYVtim1H6xkh
rDEQxmj0G267N5ggPg9uh3u47rc98jTpdxf/w8lqCvUd90UvCg/lnyzyCmPksQ0V
KQEGUYIHItkXw+GTRAjZ0EYcItdakytjdF4enwYHo5+zkYQJfKkZXSN5XpMHBG1k
jnP28OpfmHcPgH/hA8f/AvobUx1DO1hdEj8sT3ayB6mJX5grDNvJPULaqreHlgpf
pbU/LblTS5s9U4oF4NPA3H2bZ08Iow5eMpBvMbSTT89qWwcq4irhE3i1/WHhU0zx
cxunvPTPYBnQ21bhJaHQlWj3dz09OA3H1w+gCv+5tzECw85/0Xz9mlLvsRzbnMrY
85bdVlbSjGYEDf0DQ9izCTFaQ1HdxaAJLeshEv3gGLIW+Nr7BSNTt2BF/uQXbn6X
TQR9S+3g+SEUV8S60vbiftaX8amFYVMpCcEKID5YQ+2NDB29++SxdESmW0bQ7E1W
nS8BFQRrt44rdIpY/mH9mqxsfhOBM/YjJWVBQRiB1C+W/580T8NK73pAO1AjT5ly
`protect END_PROTECTED
