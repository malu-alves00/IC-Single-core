`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bsUXJmGmp6qeBmx00QZ4yXCjf4P1MsIlcdSWlQ9Un0esZ929N9nrYtfvALiPq5Qz
/6S6OTGafhRZywGNJbDE4PWfTHiwbFdqXQo2KvC5n/g44vNBNaaraN8nDBzJ9PpU
o3UCnsp/ou14JsbndDkJ/Dw5PiaWtRa8aJdM+QsSW0mpNnbhYnPNt6vE0sSJzNPI
sGQCyH1t7k+TYVKcyHJMt8MvHhkDI0eVjOYKSaD7H9IZthVnYtHperTCqkvwv659
Pzi0Coeb1WEyQs76gJ33YSHa2DZwIKVA0ndBFuCDVtaQUVBE6T+GX2FagzqhBK1f
6H7KhdSFR7BBh3P5ovjnTa4in1x6vVX5LKthBa7aFISrSbWmc8ria/yJC0WKkIQd
NqU84lgoAwNczk6lCNhUSaFElu5gEq8K2MW0h4cLTZhyCXb+SrChHUU1R0RbKpJ9
R/oNMMzOIcjIinHRqbK9eOUB4S3KN7im72CM/0VYsGudMZxmFq7wea6V7bOYMBrn
IneS91z/ibPCkpVd9VhvBbBAWB2uE6R3guUJMYeoIQqxelKZ2+b3nmiqWQnKPIhm
qwPG6XlSTpeLJpjbv57j12OAhQn8ckTzpf1KfU3RAftlmPQTcuibm33LhcCLVM8J
I1tOaW8H2cuHqwXCbDa64xSQbuKJa+HspVcHuK8YKLleoIVirZQmm/vKJlHdhB6O
8Zipzh4NEqT86ObBEAbAG+f4oV735jq9wqgYwM/FTEpbk/QTHYT6OI4YE1k/68mq
AFoTFwfH6lnr5rlpaxpmNQSxqDvoZxZVfvUQIm3lwmikS/w9wvvJ7N5AP+FcaSV/
hbKZJcTrME45X4GYsLUyAE0QGQszpejWRrOpNqEO4NKd9e3qI6bC8UlzipgsSypI
BAyJt19iFC2fP7lg8K2nI6phoz8bwsLZSJViE/TmoPkUWrjpUpdqJWC+7H51IZjR
`protect END_PROTECTED
