`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jQXwEoNdzEfUVcQ9c1WXTeeH8A3AcnoquhAHtK41xafYUo8s3SdzqBa6vvPF3rlJ
U/C9dzfeSZj6jaWd0HaLETwMFv2Ir5UpE8UUoF0e/JB0miEUrEmV16qeHKTqPPAr
UO/Myl7Eu3R6atr/jBBp9mSfAd+IdQ7djd59nCGcGzAxfQA2UcfqCQuxWwJfAXsy
2zCyK2yOYs5uK7dBaKykeGs0cc4Xp5MiTY//7PXgSfuyXa/nvXlv9FJ3DCqyHq/t
t0jkuOlsaH5GHdn2XZBWL1TR9frCkkmfZlwoMlibanzqtg1eiyBM/Rc9IL8r0dAB
Y0i7M5xINjUgWE0W0rC1kAHJFnjL/VROz/LwN4u/WHDKcYaP9jSCSMpwA4JAiNMn
xm2PN7a/VTqUcSw5weqvyBjRv/jzQ5EDJq/0vdf99jqRFq2xLxBaUECXtARjZMQr
pUonRh7AEw3oOwa6k+x+33zFJa/xzJkIO2MQEjQzzA/W2fCCe9k71qaYzAOvxLTI
k4UoAJhIycxqDsJkFDGwCl0xbEQ7IHMmKdbSBpTxLbBPiF7jv4fagpSVlINZrSWn
4hJqdoFL//+3LFPcIh1krrcB/bx5Gkr03c1wa+V1ej6NpEZRAw0DRwuMuP6LnkKZ
XByJM6pscq7j2rvCNLIpar2w+7c5Cb4tZbQSCZzHrVfVoWWsUnuq8Qtqy6tT5e5/
116XYbci5oRcVK/9hHL5I1Kdf0AsbOzNu8Uo+JLov5iquVpafa8cFiLxMm0buVjV
6iH44Dwf//lQEIYO/JSwQQ==
`protect END_PROTECTED
