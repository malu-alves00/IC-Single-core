`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eUl+8FM3dMrEtlc/iiS7Dk7Kg9CMNx7YZWcMeDGL0hlrdrlQ9Zbjf7bTdMRkhuIC
Fzrf9IaUZ7ZIVMIw9wRUV/uZxrHEAhUlVzbV025Bi+f2l+Wy6GjHZxIssZnHARrU
9kvjiLcf+Z1rR/0MR8Vd8QCXkucuNDhT2/0gvhvJMFEdxyg6HFv+D3xuON7TFIOD
ruF+Q+Aiq496upVu1PS6aag0wWyPWQqgMxC8AFIRXyiGHtAObVzSyWloL/0YYRZp
ot8Ed06kz7AYkfpDAIfNkmSSJondM5HI9e9+T0jNr/c7QqeZ1wQC1l2155R1719b
8mCH2weBW2JKUqHLOuoF085ugeSqBFLhyZRtspdMtYO0M2pbYrzWDIXwVhUrnjjo
FlsSYfJuxC7IDE1jX4UU2sV53UphF9Mh2ygKo6C2Q80d8rEkbySZP02K5c+Wclyr
yCpxHWQbqs8+dGzHKJqQmTG6pFwAVjpzITv61bgaDGU7ut0F1LutK4aCI9pVOzyD
Mmqes8nL/drDKE1EzsoVBM76MYHQHcbVhrvmbSiB5zANjwO5KyDk7w/JqzCZ5efn
DZvV9E+EX8GE9+P92nN0C7uLGa6bJkl6W3t6rhGwdAubDGW0QQyoVqN22TXUeceI
XV/5DAAJGaVjdU0B6zIMq1LN1lhedJwRWy93goK0QRp7xvbTagedeGVkPkLzKuKn
QrKpxDGzUIWJcj4+vTnf+/IqwsAq+f/neU+gMZIZDsp/wWZI1apOdcIcpM4iYyxd
6JpKFVk3C6n+66sn3iSLJaVpuRV7SpfF3Fu7M2jKOVPCP9cHEGsFjviRI/ahXHYP
K2sAYRZE4/a4HdqOuPVVmmFPwoQ+af18cs4XAj69gaEWMslaGWsxi1IWVEwFuYYq
SGgPRHgJiGdBERNv9qTWhx7jh9rgBcXSRribz9NP4HNUDxo80OXOxGKvJ+bRJm0O
9cBKHeFCzrDwImIsXtNCMxyrjKWmD9sKQH7YYgHx0Ja/wKNd6wZL58xAnoSH+sn0
MqjoCYsZpoUlJlbTfJly/OY45OhnvwJaa5VBKiu4i2gJnH276Ftd1us2sxu+ebgh
nMMddDcjuot97WdPbvHcz9zQLDYPdU4f8v64YIPR7u7TbOgs59uxNAqIM/pvwBwO
U3CpPNzcQrt8w9F8a7GnrsDbUXtaysKT1oiJqx6C9I9Q72GPvWpG4hOsy8aXL69c
QexGop7HN/y33Ba7RWcsBOGeACyDTr6+YT3AZjmbt0qUTZVGSLsbgmKjlWb2dweN
FuhJQS12x+X6voePLhylnfxgwyUhQ1jUovuW/8TL13rYIFImWVWVUHuune3E9kTJ
1ipY37ED3AWmOZug+qCoH1U93hdojada0Jkn5GbhFFLVnGNByb1t1+ArKcDCRE8K
StuoGW5UdBucmSJmCqi8yj+cQdfCzqoxdSl4OeSncg9U7F5Qh+YxvkhMkUjASZ3W
Qtk6viT7BpgQrOzkWBasZo5bh3zmjYMR4+fqUIiZXQzTB8s8dTZzpum9/z9speck
GmUTwVK0y2Zp9XSEENc2MAeQ9c06ZuO/nLs9vFennI/tATIL0sUT/ROLL1SFT5pm
w/NM+qPUXD6nP+MgAHGeXYCVN7zILOsuS7cRiOtpbt5NixLDEr56Qs/qbnhLe17S
DMPebCjxgmosNElGKFtGSngbXaFUgvbvy/gDDJlxhWg9TbR7Rgk46BxCMkhU6oxQ
87VcUh9mkiM3Jnwy2crnQzL5gNlDJ0ZvcXJsmmjzk6o++KqRG2ip8yO5frOV2hqP
aI8XX30J73MpOHTS5Bi7QzKjqyuZnhiCq/86hHk3Wl8rwJ2p7zxIPJkKEHI0cxv7
59QbMCrNYWISC+HsZiTp14eo8d7EMclkFHGLfNNGWRb033GU7IbKD6JiMztmApEJ
afln6YGRHGW00s9/Fc4s0IkvmkmTCGDdSaqqlJHrmW6yrnA620sciyw5E1Se/O4f
m1VPAiVGjfW5QuKfD+I3GvBK+mZYbLov7KB4XNdE/P1roGBN8zt35NO4+79xlomQ
C4RueWuAvm6ra8BNEgrhSa9WygBgPBEf3QETikn+Vi+2Nf8uZjLFlnI6w2wo2/x7
hq4KfRdzk+qAp7Mg1zLXUj+ULISqUyxvnM7drf5ET/tROwhGPJ2ArJJ7tGL7UTwU
xDC2/nmeKZp5XTpi6MMFqmjL5M8bj4hzI+pHau8QUTRnWn0TD7zw8dw0XwR+hzZD
R5tojUE9aTcbmDKx29G0sSBJNVAPzQtK5c6kopjnSmGBKeW4J2xoaStAo3H929AW
DrJwrfxisjQ5YdzDkWyU9b8D9QIVCp/M/wU5WUori+Ha0ey57I7h4tAV7wrhLI83
oF6OeObpvOnRtzbgadwsqCgdr/hPYbqofp8+Y9JsMdFP4qFkGr5aXU1sIi7bYcIu
+YRLBFlFQweV/V5WKvOnPp1MTnIKRCfNqZSlH5D0evZWRlmPaiEKI1T27XB5sG/b
8Rt96qgA5BXdtHkXZbAR3VqjhjzhlFXTtQhMSqj2uYCb2UFfViKWB/45lEdgHfwp
oCoOVzzkXGLVEN5ELX6IAcsiK/y4S3kCw3vdXOwIAdqEYZLGjqGtcZ2AMdxiI6Ko
Lcf+8t5jeJgg8rXnAZv8O1NN8eOAADnm6kmeocgbq88b9iiskfRE/OfUcoT3zWed
mW1rupGOZLZSRnpVel9DqxrVTlJPnm/zpnAzcsO98VTvCqsJq1qmMmAwFgf8rN/e
UuaxeCcU9E7nPZDVvlopQYGuwiWO35BW4K9Et9d59RTDB+SR5i77it3gPcIlKjCR
XuQ42XoYBHqp8dsIok9HniYbwrpvSnU1s3VCO14umMHhMUAgr39UtB++Prmj2YT5
Ny6w/M2zyeld+46Ipywj6Rxaf8hcYsquKK8SqKVFwdi0E0U1b3UfJdgThsiMKNJb
UxiaQ3YpvlTPemQQahGck3sQFr6i23LtsQhHmtcCHnmDc5Vhdajv3EcbFpwKbUdV
fzxZAN5dUceq2zyuShdc3DkTh0FauMz4ANf6RS1eF/QyJ81atxTzthT1RMFFRhQu
tKSHdnBBABAIHzOlusTSaOA3NdLrwPJRnoVxwjqS23ENVgZ+ffDp8Pgz8wBIyW0W
GhPsE8X+rnwU9tdmskomn6d37YlS7TXR5TexrqIxEj/E+mJZdwG+YFnQeC1Rp2qp
knaDaQBi/x37MQULnW0Lu4D53HZdrWsmpyi7hUk1YfIqbzID7k3g3vZ7LNIjBJg3
XoIkj9JfaNi5HTbknrPaho80FH9HObe5oLBo4GqMlLNCXamDQBLXGjUbx+xY+Ko9
MTMamqb3N/PAWfPTQm6phpytL0OtPlBkuQhzkm+sF/R/h2/LKHOJiwEEXPscsWsZ
5oXCIZKDHAtM/ciW4Ggs7Cx94eprXtmaet6sWCQ7hMVXvSJg20LrdVGxg12Sa0Cx
DLy2Zk8PSTlWkNNO/V33AN/R4myUiij88otI4HRSnB3j+B9EDGiLT583N60GyGOW
u/GVQzW+gsHMaLECjaQsSXvUDVo3/xNOBp46nfLJC2tNmXal5GjEwo3K2RDjcZ6k
PcCLhJ22dWsx8luzpS9g4O1X4UmUlk9OzaG/4i36OvMFFu3d7ShLX4Vpc99SEMIf
lmZges9GftqVKE2wkAXAN20Xr4B7JEwcTeefJffdg9b7UiUy08Fd9a9mvEP0wM+G
9FL7td63uGip0vw6OG/3uF42id4AtDTqvZtVb9ZKbXSCEFRwU01jj1/tRiGsu8Ha
hXxnNUnA21FkOlSxAkXBncIJi4POcudmECEVtlSZf68wd0XEBVaBLELuaKfXfAm6
5iC0fTt/RbwCzZAv98k6k91RFFRDKw5ImaRR/16Ly4TRNk2YbDoaeu0fUf9iBkaC
NzA8Cw2ds/4dYyhWtTlkht5wU09KBtQacZXWV0fDVfcnHgPLnO18xO4biYagF8FH
rP22e7vZQ98Lo7DPtzIcq1zgB0G0k57kxufkUMUKoW1aXu5zVdA8LlUuzqwqAyZ1
CnCUSeMjfyGCO6/FQv6gyTZVWs1AYlgCwsdOfpE2ZP2Cdk6aBvZhYuHdh1RbFsrw
X+Ep9wA6+uGtlEmdWx20Dr5iquvd+ZWMM9qaj7FcTZsYFz5kc0MaT7tlWTaNnE68
VH/L5eHovK8yC0IMsaUI22qDYF1ZiMlRFbbvKKFJWUn0a1NHrMBsiRaQhJeruNLy
XMRdDdpS8FcNIFn15xjIzpTSINJ5QRQ3z/xhNiwZUafx3JDCqMqVg9FWc5yiPUCW
QIPqbWUvew74HgFWQzTosDmqNKiKfe9Eisz+0imlHCiEMEqo8OE3mbNYCxcd8ci6
+BWdVRdjydHw2Cdu0YHM0Eps8HXYHnDkXSPqVIkwFXYhq5u/MCWpiHN6rcFV8Cn8
srCSdVauzDeUsoaS/vnX0rgHNddzvCZbnrpXZOH/Vd1IBM7luI7tMmy7BTqS9Sb2
Owcm/4w1GvgR6bFd7lI3/JTDBNbK5bxgrQO/6ACpaAwUG/6VjcqdMV/f0Cs1F2XZ
ErxxknQD+T/E1/trnu2s8N8wKB/h3dDP/raxeOmiOstdQT68C/oDl2q5exwMX7ZF
TREUCEBNSkJHQMSqqeim8SCAVr2SwLJBeOrPq1iq/WqL5k7MPTcHCyhVXhRKqEbJ
/Gikgroj0lc7yUhnHrHre6RpzXt64gYDNHnmU+6netvcnp8s6P2HTqYL7qdeIvJ8
wQOR0ocus+Z8RAKyDB5thNXU3/60qxyKn7XexWxSEOxD+Qc4NHLCqfxk5E0eIb2W
4y6IqSkLfFdGJQYwxkb2orvMDuszXnivd1rD3HAukrdUxx3KRClLe+5hNUJxn+ni
y2EStH2mI97nVQ6XvS5b/ikH3qSif11Pzut2SiSLHUa2xqULQAkx8Tba6JrVdplZ
4T8nktFt/RJEaqrAXmN96SD9359o6jPlWPDzwmfoozU/hpP2nUgincU8JecLoiri
J5dpjmdedRUieTwmPFeZYHqisJnxm4MX0+Up49YmSj2pr9ktzwgZaRlMbQ0IYR0w
Dmbt3G9nfLd5Dwbge8o7CwzzG2eeCbTUMn6p4b/ppvPmg3qZAdmiznPiwAowprA7
51o84bTukIcsKtxueGWQHoU+cftGgcAloxggF7dZ9gfDByiwguAVVlC/j3udqe/F
IW/1JSVnsOYRQbWCD/5K6F9JhDsue9FuBohPjXAUCncl0Bkz8jjhnMXS5cWpwDkN
VvC2NaJQJejwCqmqEM5p0vQ3Q0L+rp4BKsq2VuW/Ul26f7TsV8X436RgsbaYq+ZS
8Wb7izSyYEe7QutWcP4sKBwtFzcxBaJkckfK7V1tPeIAkwp8fSSZOA8+OGBDkMZr
7neJhx9F905Li3WARh6jdfI9YRhLcxpSJNXRU0fL7LVbBj/YMRmGx1lulN2q2UOI
iFxt7qTalvoL3o+TFsABImUv4jHw2CdGVyHU+4D2vX2xH8G1I898xFy35cPB+1mO
BiH8hmj6ptE4j71CzhT51VEfjUwoCbIR6OTD5Bxag7mNoJnO54YMTAVCDMV+jdcg
y7YHFk1maknDZ3m6b4TuyzK6AnI/pzm3WT9j/tVj/nzY+1leXA49Lg803jd5Zh0/
Ji5FvdqhUEFdMqZT1uoqlwZsQjmHAVDeQaw08R6ooGe3Z5yy/wDne6lYK73OVc3J
UMTBk9j0MWdKKzt7jBIwqS5ciAlsZS+sZVFwu4qNX+8t4U3B5ZJ/gwv2dtXfIghy
m13PvtONd6sDXiWKFkMfk9UG3adXH0jmPuD6gT9cNLCe3y/RwRzN/4+a3qVsnn0c
Ae8Co+mo5PncMX+4+VFrWnY3t+zVVibVCnRdDOmpeF/yz+7mMz5ytPg0r05e4cFC
F29YuaP3l4Xxgic2RYJBdO11vc3q4/8Hid1ZoPnHmfZmBXC70ZmZtjwayHFnAES5
zO3gstoOzf/v/eS2JA7ZCp2iqYTXO8ebvSnEbgi6uO6k5wd/FAZDKCnPnINNOGVe
ODhScFcB20MezSODj5+sFhD17lb8GBSDOpaqNa9O89XLoJ0saFdxTUnIGG2aMUlU
MV33uzCDFhm6KK20SXtsLeRWKNM3kw7V57+fzpa/hZi9R+nGZAk6WcTNnpdRXOzI
UJoDomSVQbNE2Vso+fiGJRSgpzC/BX5cqvZy+W6YA0ZIEm8h1WqDHSjdokhWU32N
/rFsX89sOh7di5vujcQnGXYt3eRRyhWU/vpE58AZV46uqmD4FIfgjlyGD6/eX+fS
Enj3EtQfh80hNQr3al+2KOfdx6j/s4czPko9x5a0J8V3UaRuGd2SWBHzePPr5BV0
m0f9kV7BvkgsGMKRgpErISGV7Zi2rUTqo121FZ08qhsr3uIDtL0rFhkrX/a5tlg8
Ofb+GRSf2bmhbrEyUfeFsd8oqN5Git4XW0W0LTnPRZAjobLE4XBIvJ//8AQvjsWY
Hx+l8W+Dvyb3EGFWQ/wVxeTwwef70CmnSF7UNlq2EqAQ9ZLkkra0nR8LKiYmnJl6
KDKovPbvl+i2L3xrTEVkRTI0Vlv1/XYmPjSmMSG90vU2xUdCqkynSqq5NmI0Ep4k
6/W3yzElUsaVbQZ1zCd82EUexTcvEI3cyHIu2YdcbXsjVsoqqAQhQ8QYyDBIualQ
ffyHQGrWRi5KjERHsEcM5rEN7bgKLbg1dePtBVtG8oYIhwTcKEBWc+LZA/U3PIwt
e584ktdZTAeXqdIM/qRNezsPQxnZ5OMoql2M2IM9L6djeun4yx6Pfg4aVR+5H8Z7
TulPWq0vIVOmPWCJKlE9XdzoolX9YDm/mhMr4FwvgydEgAz/a7eNeRIH/pEuWTc4
so38t2bl3lLY0COV8Rend0B1Pf/vTS0EprG7pjIL5mUqQ6tQl5UexFUyp8Rmc93V
UdSyNKDptxPy5zRCoV09rz/ykyJB/whATa4Y6Qr4QqiyMFQqGxK+z/rj1X2M/pvn
txA0C2VKoVSzhgZrcQ5Ao7Qe9KysBLpjy83kig12bCRm7ZiJ6W3Wew7hJLogptSN
YP6F8rXFq4LRaYWNCLo0KFQA/tktDBWTwKAoK8M2fg40h6VNU8G2QJDD7IzGg0Cr
P/urqrxAC3vM1gvZ0AKsVRhHLs0M/Vio/IRdMIKdaTjG2nimvKDlqTlJqE8NBPDP
3vE1Qq44Pukhs95TaZBw9GNphrKTJeZJpCZH5qJnjGACxPHyjvQEj4JcGmSOBWyO
ISRKBROvIIpWJF1jCo2F9jppsAtE6avRt9um1LMXnU2IIsLcXIpxBCMgtnggU/1S
fqjLbZCVjcu9IPZu586RBELwW3OXqlxObF9mUlzKYmhmHk8WNJ1lakshGGV+kPGq
JSuY4V0BoT00jxFGT3Rb6L6ps/2o1R7KSFgStKGrwAVLQsZVqEy7ipjThKSPjBQR
may+zElJEWmUcbX5+wcdcIwmDVNeMMJIKS3ekAXt71Wup7IPngKlVSWhKCI30PFK
Ee8fmn0CVzgVrqwh9/ZYGpk/xZR3nhyZiS7wys40ajDbOFZ0AaP8BSeht3c+x74h
gQVSijSdPgmzwEQ+0JJNae1kGzO9prBuDRJdJYj2cN+PHJB7E9IT/B7bD788Djle
gT6bCqPqGaXUNBNWsV6CE3YsfdZn8OMUlgZJjnSYh0/9HgX4EA2mrY5SPAfUNvqG
KEdJHQsriCwK4dtGvLadq2XMPjkKX2AmucRRuApqCTXnIp/YOdHPkOaFKGXyJHpb
ph/W0mh7Hi7vIt4wrloW2lIFIMxUjKLHXlcXvwPIAyGyYCXnJeuVTnVNkUgySBlM
Slg70/jrk/ef/SIO33XmHJ9fAgFbgK1NKmJMoUL+p9WXuyfkXRGz04tsZZuzEiI/
6bO+p4NIgEN/ER2PEknbBtFgFbs+5vGuL/d8+BCPVZD+CSWOMYahMyj9qw4q4jyv
Zm0P6ZHpAKODLdx6hZc/BoVz29ePyI7LFzNlCHO1DQRN+Ss3meupiVU9gMR+1fkO
tcEFWpsVTiwe/y+2W3XhN+FPf05+sspmq6M+60khMG1boszJGcPPFdEIBj9mKZ2I
Nci/Hs4pbs4Q4XhzqDCGQ860rMv4Q4y8prb6PRh6r9BKUwrRXYWRRkNXwVIl9MF5
XPGSd1djSyDhJ/KZT3LsvItKg+DwYqCF5B2bWPHpEVhiGskIU1ABbxsiegtiiMdR
SCzW7LxP/w6aXlc7OM77eyk6pDFaxgJZ2juCqYfE/utxitBLR4vhqHDKZ8ZOQzbc
VqTTU0tGLHbmU+q0lvtHIQlkk4JGUvaaWd3xNELcSc5wxxVN903plq7QAv0fqwHV
VmrE9QCEFUKiUKpSakr5vxM9Zp4VTn5QLs4ZNNGHL7NxqZkeD6Uf+Dq2OnsMsS8r
hBB0VA/LahEc6s790w39SV6D59k6CNNJ7HawMsPFajXpijmQ3vOe3/On9py4fOux
LSmfhh7D7Bha4W/B6NS7CkKi3TnWiCFpoozLIoatzmHrOQDrk0t0TlHy32Es1WcV
wIkzy9uYxw97oljgs8XNlaJkvrFcHPz+NOzwIHRjy9zdI7C0k20lfZqM6JA2/RIx
BVjdDfZyie7fHYzDaCg6chV5BPm1CXAahXqV3i3bbQsL5Zka+oVylbk4O46rJa9I
fAtRtk9erC5VoCRSh65/IxOH7wQZSyAmjkqscw+B2i3o0iTT1xjgQage2q55mUtn
SUKTZuhyxblVjGNcRemNMGOtxsdonZX0YDR0AEZqMF3BogaWtaBYwoD7Orf5/n/m
LGHMsz/2bSt27SQbqLWOofylfHoLuSQzGLEYsuODeoXbc0aJQkjdy3Y0Qm2i5sPO
0F2r86IcLdag5SOR5ZH2sTbkiVVRk3jfncWaQfRCjLH3o28yLI1dcx3MQBf4qYqS
hUC60buy2ABqeD5tEpeIJ/dtB4pRoHk2UaXwSdaF76NL+fDkJDyOd8TqCYTJDMiK
YCSkrooqojJmofleSc3aO0Aeh+Y+MBO6Yl+xN4X2s+WUpYyZWSNJvsyGr/dCZuPd
fjUNb7mNxD6Dwmi9DXQ0xw==
`protect END_PROTECTED
