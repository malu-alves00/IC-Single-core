`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bMshA6QpBS2RlR/EwV+mJ3G5Mkj7+ZqJQ04FXiHtlb7a/EeEJ7l4jzPJBa1iu8jU
tDfo9px0iwBY9ahXCtWQjpNBYqGKWCVHzO/aLUlq2wEhit/tXV5I/pJ9qUVmHbrw
KInEzDjTYiOfzdONLnIHffIEMmGLTU7zSQJcvvfGttn7cPdtf/uAmxqG4F2PZ+Qd
GN22w2b7Fk7KCMLOvkhmBwqL3jX9leKIe1nR5mUV7RUo8Rxhk5UQifKSvOcuTOq+
NIqdAi8GLto6t53x4sMoHV+UgmIAPCVxk+ekxzMhBUCd/74KyhCP67GHvYqMZ/st
z001JViwr7ZxSoPDAO/p2tBtNqaH7P68FrgclV1Z0fKY/CENUYFBqQ6p2kH+q2bV
0QeS/qaZOPP+Mtbv6zSnx/rWC9GhH/X9bzgocSaDup0SrGgXgSVujvjQJtvHJEXN
JLcpH0OEcJqtHZtfRzeq1J3q50pl/PbLZ077URS3JhmCVRZgCR+cA1LUugj+Khng
GL6RkE7JgO8E5X5oN8P6JtPA7sLvU+UAOZuO8qt1pmpmV+TvolOAJN3L1QmhD013
l+3Ol6cybk0btGeLpcg1CEL7jZbS0LRn2W5HRCQWg4k4MYt3FAI/avT+W+ck47q4
nsXibO3gnkLSpUGsYbIv4UBSwhjw4yFPWNkgIh5RpcewkmlzNQ51501Odj5lwXqz
yh29F5JIpPejqEZ9i1guR1fK9sWsJP+iXpkeNeeCANArz3STfGFg30kVNgTlDogV
RWhZqQDg2nJ/H+REYMlgdzPTzWP9apKXB/Fcic5cWH4lg6NXXV9TSlgQyWPEW6pU
iy56OiZCVXx/bnAtlNDoWFV4ikyYwALiwaRwKzNyCzF3o5Zz+WRyQtJNt2mXeHOM
Hdd5R0PcIXOtOctPj2Y+mPUnEyiNI+W+yyo4+qcL4i2zKaqPH1eA/K0M875T7zv9
`protect END_PROTECTED
