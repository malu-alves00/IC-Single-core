`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xQwMiO5990j7A42e8bUWwGlEOlRkYchTKK7bYVob0lkWjSEsua2pt1Vqjau4l+Bg
F1WmDrXC2k7z0+87b5WPFW+7T7fn2eNYQ+1SMvvovuUEfqnxxnn6dGsEAUtxhKQY
Jf6TpJMRr6IYJjPY/FE+wrWb1MZ8Bpu5GBOVe2VAgnCe/YXzhvPGu5bcqbU82syV
LhM+5EcnnUuBZ8trOeD4YV2x0IiGcQcSesAbUzPpqIcxAA1DiWXI9/FO2czK2peI
Fq0hTl3F/MnqgYEK3LoNm+y+7ch03DPfw5kF+ii6EZVWU26pHnqcU4pd/Xb2fYJg
HJnZUPgQ7Jx4pooZQ2jbsJAuzEJDsFcbvBAOtVXxqw71n1HOgSpF4AhAubxnylu1
WCUkPhrWB9FXoAfG3449p4fST0tD/wfxXU2hFpu/IoRkDangVZeAYbthndm+uXH1
HRpmquMHmypgnwMns2+LKpJ6tA3QaCTp2ul+1nKyl037TaeWrlprv0xbEd/A/9VN
Aa/KcIflWAaG9BWGjMuP+GyOlRHD6DIM/zE2X2Sj/sXgc/7hxsVQR8/RYbwJ7nXe
jB22b3rkMp+iobvU72KCjU7d5hYP+71+/csSJuoqnUaewdZ2F/C4RjrU3nXrkQjr
aBKMBxYfCnbpSfRUwmMNRDKrIoBtxFci26vnAJjQIsdxcXvfSdhMrLoEVVduFFFx
syeVY6eQEXkwGivoqPfSsWKMSDB7tYRTgRxORzdgVVzNHnNISSX42rFxTQxbaKMw
8NAkbfQdUL9kJ3BUmaIiQmv0QMLMY/H1Y3fCDZBTMehVBFMWuuH6T7G4jxs0G7X8
R9/9WLehL3ksGii0NwX/Hocu04egSy5mSVlOaIf21BZWleT9kVqteH95Yhf0kd+O
0S/+i+fapBVmiIABcA5Yb+RXCfs8MDlyyBN+nUHaBpYNzgpnwX1bFV8fkDiOkHOI
Hapq0YO5Z5BwFl7z0Ajc0UxAH5voHzzlrhYtoBGmJloLvn38WvEKMNo3awg0dx7i
s/yLWdy+wZrqSQdhhewq6jxScKn1pK0mhcvQCsxvfc+TpwBkTzEUOOeo0bsaPMi1
YL8umuYrq7QTxDmACG2NPg==
`protect END_PROTECTED
