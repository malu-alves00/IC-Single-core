`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uIPzz/oKUl4Q1vPqumh4FCy9LnRxUUOrkoLGFJlr6aM1WATb7m0TQLpEhR8P9Rra
U0Fr7kVM9JEeY1ecuhP/HdJA2hDdsvGe7zHRlgbMz8vnkXwcqb1FCyrzutnPZMu/
9yTixsUtib8lpvEsW2+ljOntDbMgYlNUmMghQNd+fOJmWxjm5W2bxfiA42ZmxfOG
dx2jR2zCYfsSC6WzjT6QlvGgApS5yAIYxexaMN/ljrJqLFJtFQ0+qWK4Wv9caZsy
XL7meXoq0TgxsQRkYo20O4V3GAA8bWcDaqKT32KwpGxVSv+0eFcOrwLcB7wpue48
V3O4EDLAtZWPy1RBzXjs2pEz+wp0skNMplXGwozeVhnIUeeFPkGC05iXlGGbDv/W
6pakFPXywbB6tzRn6vb1yr8HA0crLeaKQj6I4kHctWf1Eav0KjdT7yQu7z3optWk
ueoWivL0EmehFTjP3S71hwZKXSxo1BynRAOzfUhENM2FQB5QxZ0tqGn9DWM5xyI9
80E5om3P7rgdp0ad1BT2RTSa+etS/zCBJHjToWXdwYUlVCKi16ezRSwk+yX8e4ml
YEAfXX8Jz20QeoazdKFZbgqG+pFNZrod/KqWk9quhL60o210y3lZCSSzNSBePXYQ
VWc6rTSq9eoLD9GckSHWzywTq56dj0WML0YSxiE3QD3kbzCzIPEByRUtAHoCSahT
vDMtGGCZcai2DajmuYz4hiavVYGq138WTifEFi3CjEyJBvbP7kPyt5rocEwjhQFH
F9nfaAHYQ9m/MYZP/RW37+k7TGoenuRP9m0EQ/RqIdfDCM3nT5PaBKF4pqBRYpvf
Bav+eNoziiTdzsfZhYAxJQvAUnhJrW8KDny0cCSy+Kv/KtPLatU4S+ckqEA3prh8
6c2Uc/KJFM8Jf1c810BsFYYvvuwHwAkAzg7cvKrZY+tcrYYHcP9EzmnEvEEfjCbO
oAVlj9QfrRa/nRuPtYlDkx7Eir9AtiE/wGUkKGScfxtZgZKe7Z3jcaEiA3HvVHid
/KyJav4EEBysJZpclPcjJK0IiBN8dbBWMF1J7VffBXh34wGp/ezY9/5oN3hadAKZ
Kqwrwc8r4qDjRpbRw7pVWLFJ7zZGLSAgYKrvcXzDiTWMcoofEbGL8p8m7VerT+B5
0kYW/zoipf1U0jaWgL1LJFxTvl+G0OXDpMQDDMg2fvH4i46z3euU0oPOjL65q7Ay
u+UV4bY/y74N4Kh2uJAW6CENTmn7QtK5XmLByf9b+MzDrGnt8d+sC9iswIadVwU/
AfssE3bYwk/q8CufNKvFZQT/08EccBAB1z2+2MM0oaxLPqE1Yzz5l/qbs2Y7IQCo
aSwp+X7q5z7pTMg7FLiOkz/Gpnr+p6YGtSezWrLL/2qxY6xO1Q9USrw88SddHWmy
8Hxgysq+2fBRw990nP+3vgrHISPwLkYZxoMcQH1Vg760GFfTwtiVHz+pxr5Pl2x8
s6g0P0R537ye1C/TB2XbdPFthGeHXyzyY5naWkHuU+S8mf8WLVauPCpdFieVlXpL
FlJ/2ztB8fu9PNn9C4Mqb0Wt29fRkQrpCjBrc1Ikz4slj6OI/ENe0d6YvbVf3BqA
iKzdvNS4ET6BDfSPZ9s7JdbyNPka9VT2m3rM7TlBpTNP5JcjjV/VNfCJkx+YxMa4
aO4viBKvig9/djA3WsHwc1hMMOmm/HFIvk/kLpFsPX2Bqpnp/ktdjh5mTz2TeeYm
iGXZ66c4pMd4X0xRID3G1GbKY0NvpZsLwUY+nilrWYHI5S5JqUiHFUfT2apmJq3U
QOSXXHbHD+8TaC/GnhIqPVPNpjZIZ2nB9Rq9YVhrgNJvpu5722sAcLy2IGniPkhy
QGFWNWD2acjL5CgWF2ID8Ydv0EoemBljh+GVbeBaany3XWrjVysaDZWxEIui1Sev
I3dHP3neNd8cD+Ye0Bx7pXNn8NRZpjy6DVC27xc1m9Rj+0Gsn53dg4pP/alSJr+M
dZarw2sM23YdbQZTGTKyGukX20tpcJ2/ZTW2dsC6d4peqVpZKNFEpp+fPG6z21XK
hRZRRbNyBhj1CWFeJy0YkhJGtqbIgPcgjztXORBbtAs1/jgH9n+oclQPgB5wpWAl
Cx5YrVcYXoO5ZNthQHfYkUBMA2Jbyk43/NXiS8un7RfHncYW4K3ZGzR3Rl+S/nCU
Po252pzgapGDsBcFNlG8YH3+Nmib888PVi5S5WQa8ZmbdXlFWGrOzWkOYVECxHhh
lXMMMV+Jq9eq8pH0592eRXsiIQPyk6o+w4VG0CNhuUMHgqLKr7ZR8u+67rcV95GT
hg/fSxkc3Yb9pJpebPc4pdkcmot/qpzRxNhyrAr4iMFPZUKJZhuh/4ILyaeiqips
BoeGeUno3HEX8M+k4BehjpIAARcsaOVyFRRVHgkUgYJ7xlVVw5uogxvWQ0seFUMv
p8ufZCtgD84jkOy0DllPVoRURE1EhNdLydgN4rvCmA2LWUWL2DfPBmaBYEHNYtkD
RufuEYL34P0TfDOQq3STv6oL9ZzLxm8L3fYerJw+HXyKKPDg4z9zSY/NdKA1iuGn
PTBlRUcK7Yf/qiTXVHnNVsZWvq6XABd6eL+Fe0FzeWZw0KaWjybcDBVNYdF2oxYz
TA+T5u5/BrGDpQMLnDm/4A==
`protect END_PROTECTED
