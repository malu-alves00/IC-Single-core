`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QRmJQCRnJDsIwy4aeYceBaDofqhm7BlLjVxv8lrm/TZt8A+HA0Xtb9ArJqhauy5Z
f2io95ts5kEiwRnljjN5q3fwuhYttrIRM0+jqtSlWzECcCFrW5j1SR9gzdflYJip
4yx4f+MBOv9a6tsSSGidOUr9LvblP/5Goavuu692pNPd+W+zxSirs2kfvN5STUKH
nWQyTq002Oenr17kMDkCGJZyWfOoylTNzdzhk+3Aib1TEIdEBPMJAAhKtHUpwQBK
U634a9VsTvdQIocxwGU0yO8KJMHtbBKzC2dumS0A3fsnMnpooOUjQmq7QcCI124W
e6rOzzshASng5DsyMpvTsK6nTevWAnieR4oLIoV+Zj9MTlHIkYOITioiX8qt2Uqm
CSuwkzWIhA4uGd6LwOKwhqrs5Sdkn/QJSH6Iv1epauhnxzcB44dzHAMzb9nLeOpp
Ji2TrTWvIjVTlMLRbDvxgqAD4oHMrlfJE5cY3A3WgUNzkIKabicV0tTBl4Oj55q+
`protect END_PROTECTED
