`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cb26ZQubp7tXcnfb0mDNPC00Y9wf3dGNzlhptERXK5qx9n7vP+zXyc74N5+0lC7t
I5ZtSYkYZH+3LSajP1IK+JfX83hhe4ZUE1C1ZbrpwVAn/Gb2bp/VutjZp0TMYF3e
NmzqjdgTzOvGyjNAxgR/FXwiLyCnQJ0hQF/5sU/pWdUY8UzESW/LIjC/0FcT33yj
U7Rzvy902lGZJPoZ5QmavmTGMYgFLPfhiyZl44JEK8xZ/Ba/lV/BRi+YSEZqdbNc
R0k//XKCna/hIW35FfN6jtYTKPO1xruaheC9ADqbics2scIGEBmGqzm5p8ysA7WY
oLH8+RaZpXFROvqP86QI0D+aSLjT2vLcctSvI+yXl7F8M5oTN7jtxW2JljfX0ppk
2RvgN7Zw3mhH/1tdNlDMb5cRm9h1HKMXy+Te88Pvwnx9PG+Keb1PEHC298xRDu2z
wk3kfEmajoLCEcUIFHDmVMQgX+IuydHhV+v/bSNaHZpBfxpPanBREnQztO4u52r/
xdp5kUIDOknlPIW6WldQmCFjU+s69qZ1qgaOdXD23cf7NfiTn4wytt8P/Iff4Xm3
hxWFSg8ucq2jFlX4JdsBkKe8KPhtny4QSlDNz5NmzIISrYNBKBUX/HpptyHOupZD
C4zK3lQUir0s+9jmVhLEu6PjHwW69HE2lE5RB6GiCjEn1aKv7yUlcAcWFaYSPimR
oxY9o60d5s4r1+YKRw6kU4cpdtFhVQUwAwDUKTWwQhN5prGnXTifIgtI4S16hDeM
QoUw6rj1fbS8U2vv5XNmTOCZljgC+fKQJ0nXRlwhYI/Difz9ltIZ/hgZbd3P94AJ
5OzjZtXyAHHLlDurW+/XGPL6KqEc7iC9SmHtOoi75UDIi5HCQLB/WUKlr7CCOnp0
+BBaaVAno+6gp/kh2XzjcxD4Ykl574Z24t60HqXhWlSWGqLETo8MycK8DlRF/OiE
qiMgcAC87f/YmMVp7zXmK3a5dUXX5jxasRxqlSjtSTGGa1VjtjQ/0QLaWuLQkhiQ
GRaU/3cLTSL43vDT1GItQeFvBEc0/u3awfz0kAwseKztrdtZHVT9yZRRHyP9w+l4
7nF5jaUv3ZmSfLm+dm1Y4+K+mqqhekVVshsy5q8dxQrRL1zi5y7Bj/lvJnK6xJ3C
ASIxJyWI0kjHZWVseFyE+w==
`protect END_PROTECTED
