`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QZeRSgRpq67pOd/ch1uakI2Nglzjlq2P47LqqcbF76vV3odvfpFj4rZ8KVUtNBOS
p313EJMCjpit0LtnsnMM7kqXRlNURluLi8lcuXj5NgyWs6DBB7kd0um92EDJw2Ze
1AGj8HugVhDiNaPAdvnmgkwiPn1cM1oP96Y4tLUqZsmFjx87DO6ijbZnsDPuaXTk
HdiMbgj4sEN9a9kK4XzcCOxqXiWbvgoZVKAtTgIhctScfqIcxJAY2DWLdaLMyoI8
Zoj7uYMlSWbJ6RUxUT3cJz8nLgNu1Y7EMbXfB9DkfRQY/4a8efB85nqZVeCh+eHS
5l7cpYIu0B98kSFGL6H4vtGMga3iOfV8myAgT41X9Z1OVK0Iw6+Q1OWYCLJmv8v/
CoKJ8XP6Sz9utW+AZw28ZmmIEsc6hyRj9hkDx4JjQxNdfSLsk/I5UNMZzLMpxCjV
spAgPT0ZkSQh2xVJELCawKvq7fRRE74lmfwMgdwoX8wiRcE49lNaHPse+DYgG6TV
0Fxh6f1kGJQk/hIukuL7u4dIbD3G0s7QQxXQXG+Og9CTFLew2ZvUBbUWy5TxgRDK
q3mxoImKNu398lTsWz5iLUMViCQsVeCHLECZBRldvTN9nVoN/G9S9oPRYFJua08e
qzIbb+9dpte2lBfxyhJNR8z7Y6x+wbPU47DH5oh7SDB9zrZh9eU295PE5VT8XA+X
akhp6kYfrq1Zqvieo/6kbzOGX8+88F+W92+E9V3tXngNcSDfmX4xM+TXm2amIHhX
tunAYnG1mIPW9MvjxGKQgupIsVhGw7RxNKxeBmrCCfaTILqY54wcXatd0NKtgN2a
OmONyinB3dM6QsHv+HSC2mHE3QgUAakHjT9sjFNAKsGTGdTLlOyvzizTEM52tTQs
wsIB5TWAm9la46bfDXvoxByJiux3vVepKgG8icDV7K9506r7ailwB8DvgY0ROeYw
GJSbMyOYbc1qmqERvyNVXc19KMg5wIzlwhUpg0/7XKv2F0GBckxSeM0Waf2205dh
AvmvY/CwX0/i92JtbpauNvd+9ypFMFc1gsjnNpm8WT8vuRpN2woF6wJRHF8pdFKA
`protect END_PROTECTED
