`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cXzQi/T6fzx6+6X5DXvEdrBT5Nrs7lOzERUne98c5qnXURwGsNQMmilGdh6r+54P
ydxWEWZKq+Nfbp7nTB8/s22nWty1ELnDHW+8Qlrop9kveW8XJo6oCJ0O4hJpS3il
/IZkapaopJGUk+Er+kDX3QaiGxvmZI4ZBfgDQxk4NON6KdAOynfkhct85tFEI1RS
Xl+YoAxn9fzCgoFoPQ+IE28nxikKyA09PhJ7NdbvwVkzqRqYDVSpxDgenki2TMcq
yfTueRENhNU/ar/oUt/+3KZS0me/B0px3Ashg1f3o4UIC9gfUe9E/O738DDbihsK
6L2kN71x1LxXDDjj72mlUSNqXga6mLlxl5sJhWvPDI/Y4uOSIcfhMDE0yUf3k2iZ
Ye2xPoF2iQlm89WfOt6xmvRj19wci6VygppM6kfBitxLAj5A9Hl3PdKKgVIcfqsc
Xfj7dOznWaZznIhBhQGEzp0qdgS13+IWtJnUyXgmIqn64FWh6z2ErJR9/QQMdLh/
0eDV7QUsIbKW1A5je4rfVvf63+FrIxiLoBxEF5IvCwP1QUJdi/bpKz4fhDCHPU+L
KE1IOFIHoo3V6HHYQjritEOGAg1VMQZsa1zeXoSKjEQie6HJsz/iWg4mTbVjt6FH
WTHrOugmZ6vnFOTdKUJH0d2Ucj5K8ILMddlb2G6l6G8ytgy3w4M8bbhlohScLHx5
XgNM9cXspGKRd4diwt3RXSWjpQ8Q9LbJMFY04ZZ1F5QSgwiJMLPkBbtlfj11Zy2R
nDpLFD/H9ok98sYSBSYwp62O6DY6EWu9FQpBpuqSYf9SzflnHxngJStjOEsVHioz
h8HL1EBMTtqdsLqmOVj542lmEeXKFOuuimftF1SDkxYHK8ZtQ/SV2JmO17GNb+fo
6L5hgGI6Mk8kCKBy0RRXvN/5HBMEuqYB8+t7ljotFTkP9HhfQmzqLsdBGCKbNm6K
VjZlj+DUitTgW0KF4i1z2gaODlRioXAIA9BR/M7o6QlPfjFeFmeP+HWIkQ7hudz2
fcXw9ZukyC71hrT45dVfc0KhfFf1fvjqLC8WY/Xl/IOTDObDNR81S1XgQ5eDaIXh
vFUYnh+zgK+PRZnM2PEGSo9H2e9vRdrkXqEUCmZV1Ud2CdSZnTFolL7m4QYitYkd
/3VP7XqqqmEZ+DdGpPfJS5itQJm56vU12qpR0IzM/8953GgFk0Kx8BnxIjoLVbAH
LqyGwnjaoJTIJ0O4M1K+rw==
`protect END_PROTECTED
