`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cW4ghSUuh9ss1MF+Jm9FZuZeFPPldA+P01jHOH1gLePvv7DIbZGK7f4D+d3O24bl
+GbPUHWD0SOfEJeBAEcBC7cjXgM6wfZ8e7/OiDqVSLPU8zDAWcTrEQl2G6QuOSmD
QEhU8A09yHGAJRpmR2m0xdBTe5yKcuZBijCjjcg/KaJx56UuXyqTqsck8pdWcAaU
e7iN2I7BSKtCvjVoFkdecrGOSoJn5fNys7K4GDSX57xFU190nshY9x7ZgV25uEZ9
gYjsSJHvbZsoT4HhEwdPUilTvbChez5oSerhh6Kj/3FvicXEbANwL4zenqlrqTOK
Y8N2Wh6J7yakAgt5DHLDM+k2WefRx/GVYAfiYTQVEAUzJH3aQics8l3qkqn31Ipz
uXqo/8sg0UkIZE5iJPjxUXnE5F3NvmUQ7Iya1Lm8U1qdhzJXTk1AYJLVeG0fVv5i
HSw76Ay9W4KsMgl+ikm5D2CqBjpm00EBUfR3X9gy3uHLrh2VkQVp+9PYd7s8eOQ3
4RE43Yt1CUGdGZ/sck/RZdnALx2syEk0E1XsDGiWlo0E88/5X38w4i1bdWGpsj9T
aOBE/rYtJlQP7qsjkXEut0Rt4sK+ixuD1pnmES6+yB2Fv10gXnMqyLKq9px4cnoU
FCxycHpGAYnnRwbEJEVO7u0sR0jSqEW8xDZY4OlK6Plc6vINMalpIh92vdh3lysC
RsS43PqpUjRUDf48u89r2QN1mRonPIMeOB/KFfC0hora7KZZwSF4sCMSUbhiimE2
DaYyPtOljg2KJhL4HxWWUBqmW9YLfaMY3PH/hVeJAA4tJoehM2quaD5gAmo5bqaK
wccIJ7DY0sdQ9/RFQCtFeEePJNdHciBgBO8fhv42DYBrNXUAjkDavi8dLXnjHku0
0GC2Mo57U6zEjFXpujJcvvxAH3tHsOPLpNtoCrf/TcB1bfxTtrbPmWLw8M/DuDSO
ILeznqSuxe4B0rcf0ZNmwZtew88jtgmvLE/5rBhjsWn0/UrOSAs3k5kgVnywN9vb
n/6Z8Zmalrdy8bx6b2fy8qDttJYHIjvcPZcsSfGEf7+mZuMwezsgbojWej0U05NT
Q5aEa4rYWMAYjCz//N+iDeZAl2bQmUFk2isU1uUWgSx8HAzBvi+rLEd9PDeWzKkF
CJBug+dO2njLCa1X62GGpZTWw4V9EuBh7X5WVNe6OsyY+YlnP7r/NSWMUF882p01
qdEl9380gVuflYf+vkWOiq0lCIM2IRXlvNwm7XR2m+uOHiZj637pIUoZMkfBTQUc
NvzoGGDAxJwBUCXjVBtB3q4vgrx1WQgjswBRhIcyFOv/AlrLiFaSXB64jQRPu8iK
5eCVbmsomKcQJgtNkYykeoHNkHq9jEsiqld6zjrNFvRJclSw14lCBlB/tAF8Ga/j
yEJTrJD8Wxung+TiiNVR2TpMb7DKLG8Sjqhgeao3MKK+PiwqZyYkrQA4ZtCDrUzI
bdsPelXLlUzeRx1Vn8PJ1gNhTI6syZs8cVnzJWswrO1NVChdA1pH8+AWwcHY2l7M
BMlWePSZ+AbMper9OIzcs1pbYe1peJ85WL22ismJVKZIPrZuH3xOMnizXgeZI34D
09bYQC8yBOV3ZN1ZItvqg7eHkmxm8G+GoIUHyfdhvSZ0IwV64kmWl12p9e2gDI56
fBo5Os1tANEiKHmTHzrD2huv9xZCL+He55fYEvHWaZpoqK+HOG6OaOY6UJvjCkcH
QpIJGEiJbRPMTcmEJjeTRb2U6HGciDrvkHmodTuQ/0wQgeBG+WbZnd0Q40s7wEwG
HFPy/ohqFJF2ZA+Vj09vYHkP6eoGjjm750aJNSzCxYATdvj+Neopz5USJ9Ztroiu
5lmeXSl0A30eRIH0/IjNP4Lw6YAovB3hqneqrvMOj1vnVaCnzQ7eAPn5OD+JVmio
CaEUaaL44NlI5nFQcJnLOuaTvnP/bHdBur+LxR1LfpKxFzr9sKu/voQ9u/olVGcp
FN6Q/t+yfUCGG8C/e5qFp6AOmRMgw9W11iktaOqI4jfsl/aJQTPhW3jxg76I+/eE
GbhOm6du2AzvXkBU20S1Im2W5MQnYyO6rQl4KaLOI3/xCuXiKD1S7SsViW6fJfvH
43Orfthm2VD3FLQvQecuv/yX1EGbS3Rg6m5J9OePmBjVi2fLnB8GTIIug+VBMqL4
D7ZTt8eGc2m9obxP8EQhCZKhx7HjkcVib7eoxFMwWVBG9CJkfQNvoIJNBhwfgqiA
06yyyWsim8O7FJp97uMildzLVA7IlpL7Dlb8z/0BXMF78cy9hhTSavMmsuIMtzgP
I9rKbrsJzj8dy26DQs1DutwYPVhz+EPGpAMkIDe0i57nwhKvvvuOrrXvVpTCdBx2
0FKHTtbDaGgHakdvH730MFBGvHZ/SxMnChBF500npzp/uesVrcSLQ0ksilU3Gby8
vDyTMTcs/afYPYLt1elClDxBlyl4GNilPIm368/euexqdi8yihy8XeOrZDmVQT/D
YXmrvQIgONVDi366HttF8pcZq75qLq3FxJoVffAE5w8=
`protect END_PROTECTED
