`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
W4yrDHLZ9HtfQ+EEvBDfobjhD/QVacaxmSHbyvqYqle2SRwa2AYoNpKDzr3VLP+O
1994OoCT/d4RDnYeyMIg3safmTitz1bx6V8/IXX2/Nc6E7l5NzZnN3llYF5MzNSP
Pc/N1LX85hkt00syCbmNNQc5iw/2ud2Yvb1MpVqai717qZnyj4oGof9hoU2qP8aG
UsLyUk9dB0xLfFMnXqBASJ1iZHF9l3YUNi/tIrm9KmgEK3naysWoEGet/Ll7/WO1
5Ikek96tAUb53HO/EqzGGASbA768RCMZfnXce1PPcmO7C32Iu0AY0JoCwHVkPqIU
XJWvJi3+KvZ3/NnUWjsfM9mmGxQACeksn0yvwEra9xUtk9cSs8TQFa02/9bnt9Uv
/o+0Dpec/9tHGHyMMfiigKuyVfpyvsW3P4KS5VuDPTyf910LytqzxhQdWUaebTl+
kD/hl3S9hmxGCiDUMVllck3s5KfgagpAOzBTytT5UPWUZ2yT/7kYxN+h/HLGrEZj
olfU2zI4GQN5E6uT2yI5cZu/EaleiD2H1P1+AmwCJGtWuWohU+qMBO7wES3HCGdN
iKd2ajwpE9S6/VaqMlel1TsoAQFonnos/LgZg5qEZomfCG4JEtrX2RBcbr1SuQav
4exVSsTixwN6smMQ16aJ/Gq4Ot12kbuttJuV5JNvCLbbERo1jO7kRQ2VfuP7TS4i
qmdzovaLvGV/AmINXr4CbLi469Cd2DNgiE+y29aahS3fwuw/Ak1hM5Qzk0YXidZZ
MGAbruGt7/LdXEr2t1de5ZnpVUdIEsIjHwtF0Z9lmGWlvy7n+LYBy9OQKkaPH1N9
H+XbD4f4qXza9uLWLBVoMc1AWOlfjXSgvyx1bCm8uPHd+0bayRpmr/J4SlhkXeDu
6Seu0m66CF4UQh5mtmfI/4jIpKHVJ0WUNndyIHv1jyGu4ujLCno/EuiGlysEvAHh
FI8/fG2vibz6BDdyhkaxAApv6ZtkDZAw975olWqNzo8pbfyKRi4B17ttZW3ijlNr
qjXqD9HZjAg+5eKkF/DDk/MhBL54MBPnY5LOE8X58pSzcRvl21u0ay+8cgId0vmI
31klIqJsRAleBHiWcsUec5uzzljmRfoYfT2JOD/w2MjqgDTN4/z0iJVmGNjKK1SZ
7PBZ8hwsvVztnqQz/t/YoQ5LILL7Ju6qU5rDAHAb3wBkWdoVk/ziLaKlhfosC7VK
BsJMWPwjy7HEP3hR64vBYOO1br6dhCaT9fhvC070Gxmf++yHw03lzdLo+Zim4CF4
bZ+jFK5v0jlQH49cRTcRLpmiw6xlxRpxplgdUXr17KYbEBXZ8t9JxZ0Tu78Ey0l4
SFf/ilC3KIDfoyQMoyCKV7zzuEm9N0qjDEnXSgOaCtkrJwLSdD9mW78nCIQ2ft9t
rBC3kczrQZHaQin9ZnN+/fHNfR4mm6aDOhzy5sSawSJZ9D5p27y1ZA2lxUeYgDWt
MJMFyIQHAB5suXP2pXch0/3uUq/h2P23NysQddiECwQWEsq+yyeMXmPfFzzapnIF
`protect END_PROTECTED
