`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ryPqednKSuotuiGtitWvAPeHDxppcsyA2iIdPh2ErjeNXL4ltwUiWcAA3g4aFVQ6
OHMB6vE0u84R9njoYd2L/RVA/fm+SdIZ3NYRmkiP0++Xs5VODpraa2YQDlAaIuCr
bTD1wMDdOcvs3tcc4w1zMQZtiv9m8LDV/s+5wbxgI2dn6zRYl7n01ujczrNMEYJn
lKwVe4po4OREeTtSkwTqZs0pDznEBLURc6prsNl32dVO2ZzkAI33b3NNrbvM+sau
CcwsXgdJV5ahuL3QKVhew+95lp8t5jaqyeRnj7Aq3B10Gz2bcvyv6W6I7vPJlZoZ
031jBGFAjZQRFpv3QPLvcKwioFo6dUKaPf8lRJ52VQ344PDk7GHcs2LxK4keCP6h
sqQ1X7lDY2vr5hZdFQVCHKrlGCaskrgdhPs4Ewr8Y4NHrh45G3iKjmDv1oZRoLOs
0jFGBAKfeFcrTkNgzmOcTX/Z+9dF1T6QeKMf0oo9I6jpqneRMmJhz+GkbQMvORDQ
rp+PpgZwH5CYjiM79fSln2ez0sAVbQNYCixlbe/zhq/1dQottYBs4juJpHQN/JF1
uyLtOewTQdVm6SNF92XBvYXBI423O1Rh++wig0RURaJTR1Bzyqpct61Zsi+hj6GP
ax7nq2jVz8iG8C4X9fhj8CejhuNHnyuATZB1EN1eEND2Nsw+SChgwHrmB2tRdUZM
XZ9mmFchI1gJQnIowLY0xRhgjfFwl++1i9DAANOD4xt8eddS62bE/Bm5gALMMSme
M6DzjyTYzZnOg7Zva0czTiIDWbzjoU+QJIznRQwHpNXh2VC2uaFerw3xZCuoKr8E
2RuNfGqrPQLVg+Q+MIOM5J2gYWpfxVx5Y+aE7xiEn/Jrik2qwn5qUiVj9ifUOqbr
Ds+s2bkCp2uk2cPIt/a3un65T/StRKmsABGfsqrgtXZ2g3Ga6nV9tqU1WYIcJI+n
zajyqfOkDbNjaMf+cB+rHvlTe+sJz/tmGLhX/Hru1r5ushYLn4BlyM+Lw2ZPsA02
3OmPvoKHJjT4oPGAvZlLJolIUFjozL6IM+L5kS52FFvvuNEcq+oAa4ZJJ9TVz99Y
Z3vgqBSMuponNWr4JR185kmq6xjF4ndI2BCttCNXSnwX/OL13epdMkx5E9cxWQOw
774hrupEQeurOZYc7AWLyUv71UM64+TB+jL58AuLpSW3/uC/xwYm16IVw6yIVhdd
cZUicVnzZeBqzwyA1G9S1YG+eX4blBSeBF/x+6dUUCjaEuMOuRnfXwBFxjFofXNm
mTbnNr4wso33mKTSvvrKE1YmYvNeY2GUXDR84oeqGm5dTnwjMO56ej1vcNBYdcuH
qDALjZ9A2QSbMLX6pM/z1PVYOEPrXzPKrCkUxw937C4Y25r1SPN55T9DtFUpFvYv
DzfIh0HH8jyaK0nesx7kGJ4yxz/BvABNC5bX+59uD5Wka0TG/E1IASGEMfOTgMTW
tFHBufETnII0r/lNWnare+FAthYYN+/uPgOTautBrHem66UXgMYmyDQHZuy4xc7X
Mx/KIVMhaUhuV3s0DKfbPCh9M4j3+Cceo6a9DgkFAVn0gsdyQ7M2Uu47aG1F3TIk
KUZAqabwk1NnCrliKpOi7N/CKKLlsUkVrR6lIJNbCJHjD0+gt4toiEYU1kH7zLRG
Jz7yxhrtBRly8PDJW23jHhVhRsFTt40MbzWg9WI9y5KBkuNckg74K+GeAdZxKxlx
JGCDErh//Az0hzzYGvM3zD9NB4CaRfkwagWHHYVMY6ZtD8RhrMJgSczBfBbDuR/4
dbIYePwYIVUmQZgaKP77xLiEPLJ4PYKYTdsiwQgtyruPzC/zkI1qjfG156jZidO7
J8eVvJjNJnrKSn1HCfPqPBXhNFS3xBlgIsmHVxG6c7N2C5YxQAwyL//vP+WLwvSv
yeMzgWJPI1iIUi96CPuGS3ycyCr2aQofYAzTIZ/0E/I0NSI3ZR+7luCPOLLuvn1r
vkmp3GzP63uvUBxuHVXXV1OCltyCMPisF0Y0caXjrLRXn5HDG0QyRsq5XUBzz9g5
sfHHqdzrUFaTwtS2b5Z0ibj8MHy8SkHhijgs7OJ0g3tcxNLV7CxShb6R5lcMnHpH
ciU0JTObHanDVLrfxXC+1UL1x7YmkqcYRjnXZGje/EnsxE6AT9b6veYt6MxsaZUv
WeZaFdnvRHUtdcA959ER0WU15cmhO5UKFLXyWtcwSowVpkXAxKEfoTtV6i2Tjc0T
6sZMNEV9QG8g2JIyzvjFT+WB4eJDyELTLCnZTXezrGVoY/4XqGBDb/2w724T8w85
XFLvrn39R1I0eDSQ0VNZ1cK4MxnmcSAjGB3Ls7Y1v5OXqPyLfJzPoJ70QG6YkvXA
/RpMmQFsf/RuA0BUJyTP4rpV9MFo7GMtMgfm4/J0ZbCokc6R4wQEY9AT7t/7wult
qpCkzfAs+CmytNXIKmMnSzMhvAqrHcxF/8UezKj/+d5S0XQlVAjUAf9MR7Xdcp6N
OQqzy2RVnNhtmAbUMhjl38fEbHIbB6tczMzUZ+vPLr2t3TfIHIICD/CTbiCh4hiu
FWo/Ny0JYc+s30TK4vfc0O3W0A/yPoQOLcO+7Jyu3XfyKuydJB9qfb/ebMU2FsNv
+Jb1q1j4pUfAoKaC2z6P4eyINKQggam7aiMvwLJBqTN56bZqLHithItF5iP22QEn
qUpk0/ZIkIAuC9MYKXgP9SyR5f7kkuhzMgLwCEiA1Ynd95HHEEZgy6TVI/z5bIe5
fH+7AH/MSGC8WtpDOAatE7TuLrGZYgfwqJSlo4mpIWNuNv4IepJfvIKCCqcj0Shg
pMVw0l5ELYuPfGo307URWKl2bDBZ2Cf7P9KP1v730MruD6x3+YPJiYrBz85Rsc40
3N/Swmp+CrcGLmrQOM4GYiXbVoIThhZHp8EkaSidq5U9aQrtqqiK99n7YUpLhz2X
pP/ViWfL1yzNo5lX1WlgiO7qUEQ1w6sl9/T9AOnszk6BBRxLiVX/q0mxp5jmRuhC
4bLxlQtqBNEPawjBJrvqKqLAbjPv2wMWasvZTYirtZTTi4O3Yp1eKbLavMVsweD5
yEiTAWmbTJX5/6/4wpiuIM75XZzHFNQpgJkFHaMe1KUBqyfXFbZEqDwmLfdNDP9D
pM1iO24MbAEauwa7NEw9qqq7/1JYH19jtbzf3xto5ZTZ9n1u39os7ymXibZk9qlH
sreBEeedfvydNWE8Dy2Kh375ABTaxqvxVex8y1LbfbgHFxrl6dLodn1oDaX1B9kV
yfgaKXE8X83MQh/Y3dpwYNnLKu6krhaaKbp9nY4SbNG7rdk/etqZ9G8lV3kdZZwx
qrLm80jBDVS/7fdrm+bQpElc1YhbzRxhRAWWOaEmD5CAy0XbsbSQVdLbb6Vz+Kef
plQ1N+cHBr0EVogXPyIvcz4QRV610xbwaeCHcxlxojnrjdT14UGtFCZHP9BqgeBF
ZGjO42UTXK05+XbecWlZ/hzBgnutVAWL2I44175dz2JmRyF3WTMAPUPRXa9ytB5z
P+6h4V7I0wNUNYZgHUyByZhYQPI4YObx6VJsLLEKRld1iMmFYTrTqYOsxigW1HPb
QVmPKCDqZliwF6z+rO7bw5BxkKvse5nKpi7/9NRETHgxslxeiV8YNgrdJ8fYBdiz
TnLx8lVSy1zbzXUcvvOyL9RMLflc+hZ9TFZsGh5ov8f/tIp7GfpM7/3idXMy0SUE
0TAZgSuQ1Sl9Ah3lBSuNl76/mKZxNCKRC47rtppqyhyUlVsq3mpdfdcGzTySdmH7
AXu2ZoZe1EjH9pAKirLEtiT+ED31bAVweNe4WIyvnvjn6x4UIMdTkTqklX0z3P1a
YE41WCiExOMp4LyDXlV0O4ucDVFW3mYAm9iVKRBjujFwEPzNPUYCrwTneCbqvgSG
8f3MbueCKZBIfrThM5pOIHnfaUb+J8/2IUwpxw0l/g7u+D1vtMj42PAZ4U+NQyQc
7g7V6Bls3CBjIKDyyCwTslB1lbqZfuiQNv+105kcVkrL0Bd8W/jHUU0jR9xNML8w
fHGIy5SdMtKki9P5BnmkLO8M1LiQ02dO4/kvHUBdXmbOAewSYSTWZ+irm5lo2Nxq
1OHRc+3jc8NBBjpCJl920EOKgoDCmVAHTzBOe8FnexWqEj0bfzkK52/HEsWDfwzA
1AecBa6aXW6VitMd2fL2QHO0lCMxoGX5NUGcKnd3Jw+gBxQaFRvn4CsEkeqcADO+
Z0kHb1utbw/sYzKE/sz0jtbidQnaYO04NKexBYpKL3SaVw5pybrm/hGv1cWLb8MJ
gtu6c4DNVzz0CT2BOGjW3zIo41Z3cdsWpGAnVsV2JmelK02j27J2IpbKArQuj/Rh
jXyY2u9Pe5Y5uCVFOkdq2FMA0t/kUhMYY6b/MbUY7Y+5xYNYFNNkYk3QkNz4TH0g
xLIIHUUNf17AeqeF7+Mabbvm7zFfVFfH05zlyzXhjQ/Cg/w7Es9DeztmfnckvUqH
L4ACBEOkQkDOCU6/mLh/S9c0JWeC1iaYaQYFprOiXz/cTY5YLuoPW8IHNmHVdGNi
sEfv4iyBFviWhRzOup69Y3VUW9pxFNApE9TItu4rEKzCSWSdm2fc4be0bRqbQ9VQ
lGA/XZzsIopnEkF2L7U2CW/Fgf7hkeJeR9jLZiJ8aiuOG6A/14wYL6mhzKP4vULk
MHH0K4D9f022cPGf3w3q4vsPBgBS75xsJYi/k378UI7+Q9z0XAc2/kaojnMrsu32
/1lMTw2H3h/AglyH3/Amf0muoXNreaWxuD4uLMp2HIjz83cY60SvjCeHqf2FwDDY
7muU346DX2k+MDgbLRtdhFNNpNal959SWBFHC9qFd2X1N5z+wae7OVdKN5edxcwP
9N1l6VeeH+OMg4ru1NwmFkymH/KyDjfKikdDtI3XPErBjVc8iZzSWUeCAKNZfjWN
nTMxpfgbkQ8o0DNEvl38K9t2BvKZYqGAzvHL77YWdcABKEM3kJtOJh7BX7dNGpQw
hwiaVoxJWTGS2yZMiebh9GPVp9x172zwgAtJ80KkEGryTsDYaVz/yHivDyHndZ0L
ftVNYvyybK2hw6at50DhHc902JbvsYqQZcqBM7yUfV06iVMvDfJkfTvnMZIFRvK1
toDRNyEr5T6FwHYWwMzwPzWFJ0ZZrkmkzc4M1RAdg4FXzfNy6av+gTwcB3TBb+6r
RqhNgKVz834pMmRHz4VwCOe3cterGCzMh9fQGC+D1a2xSeYgp8Rv0otaS4cNfa5S
0YtNX2JLYPo/vE3jq3Me6J0FoNW1Z132seq6K+Mrl+GG+pjz/bQ5TRTiGakc+N98
Q4DjLF8FulniBsWSenNpuIZmg/CBBuOkMlaticAgI9QIilhWOS6UYJeh6nVA2PwJ
lbqiGzAOFzMGfb5WumAkiC8aIijNvf9bw3+L12ZhtQsAVVXTX5nVyoH2qMQk/vsw
0XmI8boOB6473qXzJ7LZHij/0xYN/Air/UdBWQVxdV0LANgZyR+hQfBN2apivOom
VtWFaVRkputRD/4iRVDaFmm2sWbYHl28CSKqKObbK6r6kAM7P7Dr7l8EbmzHUxTi
Qw60g1ftOMKL7ezIrcvbxZlM+o2cxJLPQO9gJEWhycb4u1OipmHQJzo3yKvHG3Z2
CGFTHUa5VWlytBfgVViar6OgpLVMdJMNmcmKGcQmmyUDtdSP001ido/0VVxv4KMY
i2e0UWBbb2p9EDLuO4mQFelMf+z23mtuY3S84rVjhCptRzJOzwd44kJitYDHeFAy
plTOfiXeTuBmUQ/mo5TvIaZR7vkBCLBOnA7Xs4teQgpR3V1fvtsyZOgx4xnlT2Ix
qCdptdJls185RqIItSF0xHibDm+ya638C04iNdsMHvNmaw+faepg0leykyksQ4T/
gvtQkI+V3zw5mVbXC6tpwML2L/HS/N/4r7l6ivpN9/gGaSOtFqrwRXUBrXmRJe6i
aERhwfxuXFOj3YDLFPTjZb7nkJZrhvrZ7ucWdrfztgALmUJP6OozNRNtoCtpth3X
OS4LbbBm+ZEvx7kseGyOdc3t/O/dgpJrosXqAC4sWaugvjYtPfgvreU+6XFVJ6RV
fvZpX4Bq/SX29PhddET8h8+VgkdZ5lGzJ/ethQsy89NYbAqcLv3ht70gJlnr8Kp1
cMLuUNkZtqPTEGBsHtP0Mwe4xTTfhvYH5ZaXHezqHcmnAtEP6iCKtMBemkYIOAaJ
jyFRd/9AcWzP93hlT1ewRIqbgjeYxS39aCMbBSVNPDpN7FgX8aaKtNf+OaEyBz7w
dwL5NndcxHtbSGY05RPN+trbIWYNtJHu3ruJ665VHAzGC0bAYdofBEjo1eKt3zEn
sGEtpL14W1koEQv+KbMlZewLpZt56L2kqRKvu/pPEwNLLYALljlBggoKPl2+1NOV
+vriYgVLvyjRXVWbUKODo+wUOwC3Pmq5wznimfR2MlELmlPYgA/1nPUPYlkunwbQ
tjEyLXbZZTq0FHoNMYcbPFoHEaxmqAYsZICOqeacFJV9LASptH73n6syTH3upztq
3Qns7aU0xxdHhRErFDzzmAOsqN7+DjJEXjU/q0n50wICVOwpg63+DmKOkDAW8/MP
MGTxB3FWRV1/iZN0N2e1jsgfPDHj5vGTh4IqiP9mwhmOEdface+sKYQn3W9JIPA+
5+b26byFHp4Rp4iXhglMsczt7J8u2guSZdbgkJBiwtRNXJA9Q+YWUF4rTKOqH+Ks
EbXqTBxjYB5p8nh//JGnNkIUcqk95mRKJVFbYmgV2P94lZ1p3Ue1j7GiUPDlFvQY
W/93+Ft4LNMbGIzDlK2ix0VrwYwQ4fGBNYgyqz+4XsjKbOjDDd2x85FFDC5ggVL3
a3NClAPXxAgUsb8XVA7GSkL3GaaSGphgqX+8zkdShlfzFMPEF4HtL1qZmfxpwjaw
lDNoo0cAwWZT/9wpvstemj5wauLAHzZD2WDPKicAm9r4pA2mHwV7CadjSTCjC+aJ
w3bN4EeCP8Fm86cmR4DOjYoNLT65VBAh4s8RiV9h423zNjipyvnbhmRhA1IKVsIx
w53eyyofX4Db4MC1WcUWKz+n5l7tltxNAWNzMneYjcmyk3djJcvNE2Lxh2LDESCr
L/hX3efjD3LcVMCW/rxQdBrXVGjkR/5cArMmeIRRiZXv1VvcJ5Dn9hwDKq7mZfJX
4arrlc+BMu7DY/RNlgxDHZs+GIavsizUpNnDqa+M+92jDOpYYmMxpPCSXTtLyjfy
0qi97xrDluYbE6CulQMVQyVxyjmiqcvdI6U5Se+Eohrl5lL8jUnzEQ+RUKAhbiAn
CbNkZHiWOMZVt5b2NcM89uyUarQDBvRnI1KM25sRZGq4CtD6jOESnd8/pogs5Lqu
PfJmZ40dWdhhqUAZ/om0hq6PU2e20OL9QeVvR/RFHqWOhGzYTHT/YN7B8sUbWTcn
UrDvxi8LfOfDv3kh5douqb0K5+bVS5APHC7LMC+K9TmLXm7rgRUGtJjtMcmNCs39
kS8MAJaj1nzXW7/zjrJ/XpoznyIfDoXa+YT+qrO69B8cKVPAMW9MltPplwuKGQqN
HYJwlCRWh3d+5wmcULllav3kSSjHuN1+dANDkDirQjHl3j+5KWiI1AZTfqOaEsj7
XC6VVwVxdiBsC2KPMdayIB+KKOb48BxRWMcJqrzuZTG2CyyrUfqGOTSJjCjupnnR
AZIU2aBtSUxM66Mwjenb71aWSgbA4BG1wTYX7FoONacasuUP4RsIia6DGdLnYgb4
o+G42is8qdpH4gdLyuTCMwcYeu4PWVlASC/rmLB3qOe/jo44+fB0FZvLMTKxvrah
IvjSAjO2mM5T6EvGOy1FYH7LMmZrMdgp6tEOIaQHmgLPYIsi31+gti4/FeJjlGtI
SiTofls02/sNBX3PXK8a6U4XgMRLi+2MSSSOTHdBWNihohpsmdyBAqB1j+ynHuK1
/j9aD+YTUyhF7TPwGV5zewI1AkmRJek4R8MEguF6ZYmb2kHKCJ8+85KuAQTPEm5T
5C904rsjvRFpCDbxPuNRGZI1HvqJM3XAZt5lg2skCxaekwkDOauVmFdpDgJ1foht
y+2cRyuORGyW89+wsA3OAylM1b+WZdbu9C0z+iHqJ6PUXHT0p869+/hoIC00ISFO
i3+TYKHMLN3GD5mhPOaT5IrFndj9y0n3Sd6mO9FAF9wfRbxryBS4hX0zptuOKc/t
DMkHhwIhmY/5b4sPzil5DxCyDnRcQzITFrkM2+r7KfmKW4rLHql2OOATqWxUJRRa
OJorrKHYqewYvrWgOrDRWkp6fqI8V9vdGdx222Pp8PEOSXDUHbkDlbmhZ8bJPDGs
b+n2tROc4cQ/goSNUx+KCwNUiZYeKxroe+tF/ib6+Ik0tqXYnAqls7S+CY2uPekI
NPdVTs6Q0gL2T7zpGHcFbVhwGNryPeGxOPT//ooJEiOfHAQ1jy/Rpb7Er31k7YOK
353MmwjnVs/T29r/nSeYvn138vvP0qrRBo0ps/64ZUbHTghjMROoGscAC3z8Doww
Krpam/Ux+gKHCVpbw298rhiv2ey7jXvSUBvK+M+nn4QHKoKdqVcnw6+FmGZJecsR
an3dRMQXCU/l0pHeDCRIvDwR8mo/2Yk+FkiRHjTKJVDfQyiu6rUS9wZSCFGIo2zs
zpbjIP/rregaYnpq8m5Ddh1JM10vqUhnqKHRzN5XKpSbn59X8b7bWq0AMYkOZ72G
/ELMVB8CAlQ0K1tqspgDe+HBgi61t7h2RAvVm9FxZdO5VyrOasWmuAb811kmRuQk
Pz1YvWmx6wLQ2A3pPqpKCk57KhvOnyVIIBvozA/H2iuckqzrbsny3d0O79TiXlnS
UVfNGIPGOLRQhhH4ibp6mhVsi/5CGZJPyYt47EjBH/uPIYbKotZVH4hC/eXYWnP5
JIsSil5r3PuhqdglWXuCXIkcUn7nVV0Iq5GbiCtuLS3kQ0+Oo6NNan2ZY9VozUNb
zipcMmDAVAnWs9FWX0D07j+XFLijZS88zaLunCbxKaAgzPRrSFr7PFGIlH0QIHa5
XFPM2/3n8hfRNmxWUWXCwLBYnPTq7R6sB9XyyfBtDrFRgjfUCPP8s1leqMshVUVJ
+oPxYfOY6CGdaYvS6/ZKg879SRuVwZbVMjts02U6i3qKSSidgg3EypEARsCk8udY
A5MDKEhqqyS38m5cb/YyhIqE7Q6z1lLDFPGXOt54A99dvhFQ6Ryh7IZNHSdO+nha
aUn6oKDd9gC03iE2hhBoCROYza3xTRF5yji5Xz6P3ihVOYAAEMuyGtTzZy6LW2pC
u+pooPfNrKQKMTcVpWJtypwn//m7Q3mH0xgLpXMxH4H0KumydZnsX1fxzyTgtgzU
g4ItEteaZ8fD9+F3+tuk9MDMGzIfDqXgIz45jrQIML/AcPtzoPgkxeEAHmCq6G8j
07RseNx58ISBVdPSAWdsimdSTZJ82dtHtER7egfpyoKLTjJYvuy1Xj+Ppa7n0YQ7
HcjWpobhKWxHTasD2bPfLHxU2+xFDAbxQNNJR+lFDCpEoDQUCyG7+X5WOy25JICs
3sLp7OVmAnPB2nm5yZdVvGyORXGHz3EpPKQqmNYkpZvZojp1HJ/NOyHeSml+JH87
3E1PK08V6TqDkg9jtle4bL5si7+j7t53cpCQ/D9m2Gvvdu8iStfwJeIrW+UyvzJD
fVklQLGr3VdTSPu+61QwI2WSPoz4Q33+yMuEsmzaqPyHiKdjCKVP58SyPKZ0Mxip
yhu2TX+avmE1mQX3ehL3e4qdvagOeBLkWGRWxt8T9cs8tIYdTapO617KZyZgNXov
P0OoGlTtG+NRM8gZGkH1npgg5jmtFGtyrXcxqi0yvsI2iVZRO2JyTTN+UiVzK/fP
qLvG55JgOJ89mghl9XMHcb5HgLNcpN1Ride5uOd2YoU7qDt9BL5q5QlibMaTLt9f
04mgytZ6b3MyBR0gk86cHvkXaW+NlXkLWYU/EvBrMF32Ysba3IsiDEuw2Xsn6VDy
kBcsFcYP/TCqGff0AQUQrSHpl8P8t46Nd3Rsgk3BTE0L+fDwUn90J66T9Rc8IQHB
O3Qquw6fPd62+L/kgWAhEI4Pk9D2HQA0//aAxh0CV30EkUZ0vUhYQkV+w8/dl/Vg
BNl1PY69tr2wPhVRnq0oXKoaiEaD+mWtETk1ptbcg4wcsnrvEpgxysQW9DHufWK+
CVe577MuZCn+675iU+5oS9WWVxoAo/zPKxd8lkn8mzv481Y75itZEfkkhxvjM+4W
cBeZM9oHN5zjO+I58Ud8GpsaZjKAKgufL1UMb+WcaQ0HSiKOKtldN/XvOsokLk/i
m6kpOp+zChSgCmsCqykptu2dV27d2FW1/Cb1S18C6HIzIV8+G5MLAL4lL3rkE5rQ
Df98m5Nfg36Lnpyfe8B4HMNNoMWAF7yh6/KEdIUCg2OP7yt+06b4ZkJ6g4h4jgLp
SH6Wk8NKr66MEb/gwR833aQiwEZ854BP6unNU3UXpIKvpN7T/Q5wOWazgOkSPBuz
08xwulhWdgKxJAb2xNRZPNPxrzVbXzyS81IjH2npOyv0/Mj7CzT7EGICOojEEs5R
synaEPMg9V14gI8Oug307PkyI87FJUDeKuzFbyKorp+Y6YtKs/CEeCDazL2ueFLw
iYmK1V5RXWmmTzdyE0gCtjnj6Nrf5uGZj8uy9fJUkfu0lYzF9KwpHes17A3nTUVL
mtu67omaoOB9tRA5R2FDQompFJiFQvBqr0tD7g3pWQi+FJ1lPq4MRutftdmQXHDQ
PGxFlRjMPdVNrJ2FiMUOGgpAaT2epq136GlLwQhVcIInzIyPbFSulCum0zw6Z1ip
R8NnvT0PK5aQGFRQ5EDK39NKMF9ORNqhfK6l16aNjY2p8KBPmHCyfpLH183/nuBj
nL1lVl0djTDcLOQeZKKLfl8APnQpr1VdcZprfOFkANxo49MI/9sVSZ+kLlYnbQVr
N0DeEi0K8NAGd2dfwhg/ZG8/OwBsLiRHhQS2Tgx6RoOfwZpu1mUBbg/2X588A6oO
KTTfsnQv7ysBVg9mH+HGQFXO1+QdEk2yXqno6Ur5enp0wQgyR1LhG1d1nsceWRaI
fs4U1aEMjJa47T45P36DLXHEPatXoghnv647aqUcRcwSvpF+tdq+A8znUmJw9vpm
k9wbuSPII9P6zO4XSOsY9LLkY+7ebqkR4S9FXi3+KK5OpYxYFpgbzBnUyBlaUt1Y
BmShY2Mn9Ni2vfI1onqzFs8rPPT73dcEe7neKPcu75lMoe51V3Zc+nhNUaBRbB3G
WtRLDl6Ezxh2ZzCuWpKq0CnzuIgNNG0bjTNKY/c3MPNWySsC8S8Lc3zp6elEam6E
9yW31XA0vRpSNattN6nz9kG/vhpXtpQHJcV/YIMAjNY+TV8r5IMtuAro5FD2HjPb
rPCGaewAL+x0DJlg8coHYasAudAsj13vlLqeSkjTA2eFE1oR9s0C6nb1ycEGeiUy
ovKPTJUA0d+u0fs2t4jVzROiv7UbqVGDdFMeKPjkOFklT3Hq4S/wXgEXrxWE4+gy
jCaZ0VvxIU08OC2UkhuTwhvw79JuBSW8aywEs3aTgFA5bB7ubQjeniVbkD9QTsS3
fTJyMSWgBHTXMbVLK3HzHn4z1bdJM2lmAwszIuPJtSozbNxY0JlgmkzEYn662Xuv
V9IJOb2dFRS7Y1ioC8CeprO3uM9E4vFV3c1rbXOEDKb3r0tKsCBR/sLdsxDkRf21
z7gq8IL7ARgH+W+WcoMyM7IcNIuD4XoaPC3q75b/D1PsvwZF+DRa/oYJkzCyZYwt
jKgKofVG++FWru6AQUxnLQkFl8fAxKHVbwsLHyUuExeyKasSVKdFF+WcfBrM68co
hJwYxd9NTcorVYwRqWvocV9NB3PUnue8rk4ne+DcFZlAQJRcoLDSkCr8jY6KmiIm
DxRy69OvsbuaIpKzc6KD2qgVUHV/DX/X6ma7KRR5AxIw3nfl6Adcv8tAEnNKfCFQ
BdcsxmyxdQ/ZWRTzhaCd+zi/GAtKH6MU6WAYASr1mG74CQzRjJ5ZSqklTBbaUkkq
8LV20gnp4oIPYJkS7h8SFhtWEZqQpKDp6bHimz9f942v+BHv1kOfRk2MzxXrb4sh
WsofvNYpWMhc10mVzNmC1JR7NWysAOMZ9KSkwqGSTvgjbPSpg0oYXtySiq+bctcB
fPsrUjv6Z05QPoGO2F2qmaC7u2xjPWtWH2ymKQVLyuDC6K29gy/kGv3BlEauy3tH
UPnJStCZWWTCPHe9mSuDB1IMYqpqm+DnR79vnQnt1qmhT8NXxV65qQnOcwhwy96f
LeyksQvH0zTr/PIkPOJ8Dh/4N5wZlceb2Pj4aeX9B81JE+IR8SOX1pfX5ahCyi3O
ob1inzwk7qOOSYsB7YRJecCpHI7aPYZ4wetT0Rrb71s1j3w8EPqoWAe7SckXNgSj
40SgEloRRIrg6LW4e1OzJfsNRL6vn/wl+z7Q8LFkffJmZutPWWr6WorWqZPv9sI3
DCOS2TPoWkpYJwbfKtbvsJBS/WnfZDpYbilQBYYJGKhvrF+TjxABpSCxlq58m890
2eindSYBWHtpMBGHKM8XRwkrdHbyon5cQYuLZnO+FSspYPzN8/43AW9an59j8m8l
S2YhfeaFPykEw1pH5/AsgNl4AYS/gaFoA6dFHI7Uf/L3fLYuSn9l/GEYGCfmWDLk
6n/5XYP4ASYqh032NpK1xIE0T4YxTfSgAm25SjkLlThbWjDSAwVFeBydVsYPIZN+
3Oct3AU8vK2uAFa3iR5e6Dpj+T8y9AtffDmB/9MT6cpzF6VqQTPZgM0kXVybeSrp
gbumKrdbvznOsA5u/1rsy2rwD1PutsLfpP/Tx5BObrfrJojO4vIDofHTG6QP1pGh
/1LY3y//AgzgtUW6aO7le2chGBc/5sDFSLFEAGd4cepuYa3yMiZFOzUN+AycxyJI
g9TrwYeHBKN2q/0c2/5nKU9iWiAi1kRcg5lPQ6swj7Mt/ZBeDLoDzUk9j6GmFs1x
qDxBW+SOWaKMZmo0U8K9u9u+vE4A+uFe0uSENHmlCXxdW+Dj+CHS+Ss3UI3fFFDu
VD93i8MIEWeiMG11vnAivnQzhs317cxiVCvzNg24AnMlh9QE4zbwbbxZiezpKY7Y
sUwEE/lMKZHt3OHiaJsSUJW51wO6/Fb6aJORFy3SNpfcL6LoiN/I6yhzIX+8NM2x
PFfPq9opUnlKivDs7Jbd5sDE9K4LQBt3O6pANXwYJgWAGMOB2ULVNrs52sV3VTFl
H44zmJ/eWqqcbFXewTYimCyyoK25yirrkxgGaVJZ9WgOWSU6vSE3UVsDn0HFC0LQ
w6KpM/JZuGDSsObwxyzxSPsBTxrWcVNS5YYQHDGONFXzbEeEhcguYS63+jfs2i0N
NrBrGnBU6s75g0ErQGvXp3Zmhxx/+j1oLyq2a8sxqc3RPZFF3Z62NaPBihvWEqPI
7O7KrYB5V9F095FB1qbLam2/7Z5Fr1eYqeWFUQ/x+o52bdbX23y89kwH2Rq6J4L6
aeK035kgi/5wcgsfdtMBV3q2koW4sC098rxBEgrLs5JgvFtfpVaiEkuG8BxGDF9F
3WYi0Qpe8Pbfa2uwvZXJfrEDbLhs1rYqfaOatASGBQqSgt66x1pGEsFvTHfW+JLQ
Ou103sYOK8YiY4AQPMR5SiCTbGsqWlI0e3eIJDLQm4THXyoaztF0k06hpxrH8Bbf
7E4MmArrBPM6naUjK2k5RvGBjGuKswwmV4yxW550jj3jqSRStEa7wxgH2KQGKN0n
UyPXyNibWtHIRpW541GPpn94g7/ITR/gw1KHHaVUEsluozDmZkU9uuECFSHEyD4a
O2oQ1ikoMesAw/1T3CuEN2pP5HEmhLreKqc6Dww1CfxLAbPrF5qDLyaTRX6T1T3L
1o6aIbJN+hbVTf5yxpP1n1AeGbd6YbFq+Pq6nG/SFSsf1sxuaxeX123xE9dO/2jD
RQU+u9rO4IIx9qpsokkiTBgitIBf2i24XkBgMAG8l3CDun/rZzP7DbgHMZVjprgH
hzJdUdRmoEtsFQHlAuIlLj9S+w7tFaIASeSJlPRi77/AWSl4SB7PqDQRoaRp4vtr
XODl6pRL9DT2KmfIV+jM5sbcjg9l4ldyMKyRWxBUTUZyMOquhVrUShhICvZGXSKZ
wBEyTyEL+G2jxU3+2XfR9DAnAC82x/T+xFaUdPlT7kl26YBXC7hDTc2PW+bdK2cR
Aa5B/Q8keBrq4qhiwmDMsRqfXzHw1/1cFOU6hWXKntLXG3rmMCWPwyOiFM9JyaCH
4sFL98RS1pJwRvn6drTPWFICYhctrsooR03+64sHbpuMlUjIIwKrRM4VSWoEg6eA
meoTHKwrNhecMTVQIb41qiAMI1IQ/ljbCv+xFgEDIjpOCmH3zVtnnCtr2L55rTZ/
SikowB67x6EReVsZ5S7TWfblnYPXt2YEIFkkKT/iu8/OkUBAoDJ3QSxdLg42ddiN
Mk2cu1NuJuovHcBrtkSPBXkhyRNLlA9cxErR1UA1mteZFYXnSZk9q5SNAKLgJgRz
YkAnQFvWHJiXQVQ3Arzo1vCC0uE6WOgVUSRrkbLPOGYAcoLhiZhWrQWna6ZDf7on
DOm/kYiOrSYIyQnL46pdEQbZNJsFiwO7jf2XYhm5mBWmMnKlSIsoSO4aMnQWbJfs
OC8rToXPYmmA49HgLI98JBnJD4hw3Fre3VKAeOo17lJPFZOPfK1fCQiUHcEsm1xv
biBMMa/YPQ0zArC6zHj6iMVnlq+M/7LnrQrVZd/C3U1JY9SWFkae4+Nz0UZuBIU0
3W1BJ8Yx2kMjt8StsKNLlZqJT+QJh/shtME07GBKDnB3T5M8FBKTrEMzIokJr9UZ
mL3OeQCL3HtsywUCIDTRzr+nP0rvsnNKC/7m6apD/f1DP2lM0+ED/r8+BaTajOqJ
VqdYK65czcKYzL6aQH4qEctPM0j0F7rM429wUd0oGcc3x6R7mCrj2Rl//NL6CgK7
W4CKi62c3Kyz5W9Yix90a6M5GWZZv2tGk6er6J7ugkUrdBwCosPda2ToZzc9aBQ3
tE6O/Naxqudnr0EuJ4ehgPUc1iLh//Ay69uRkTtOtvn6HUGcd0+hz60oSidOkh4s
zSgLxEk4OeFpGGAQDZzCHYqpiNQvJPbjccOv6D3QA+8L6ZF1gCSU0jTn+5bW3UU0
b2x1/Y+WgfEBGOJu8AAFPudZGlu4peSZccpCI0kjPBl8XBiPjwqVMqgaYMJ6vTgO
ytX3ScMXSPoZJb3ZNavRQdKMItfYjL+lPI2yCx9UkthHbbLws473KosUhH3YyVE5
FoAKxtJmQBPB0C3+zEGkWHKKt1U9CzJTfMFTh6BE2doOKC4G9WgICPcebk5bOs1l
QB+h0CRAF5Y8phdVIughmiIMBMBDcPQ22x98FzpP7Qv17O7yxM3qmhxbN7YK0XEb
vP051a2gWQIw5fYDsrsJc9RHebomSr2vt+vCXtoAH2TOonK7kYpDFYDJb1MOUStt
3HnyHch0a8Dd+vFlg+NKhaz773CUWOSWpIktDfaYYU/OOMgl+iRiaXaj6cKRXxkY
WQ8JEajw6q0VZdzD1cpcNAxi9dWWlnkrWSPhWE+ggSFXNg8HdkvrI+5BY/6BSot7
G1i+aj5K7AalHDa+1kY4s7BWE2B2mebervZJ+BXkJ9RBjjPbTkDQymS2cxyBxBLf
Q2WV7fllm9y9vhut2wmk9DYdn7OkIBvlPUYv6Q+B5DA7AGYQluKvePT/Dka4fvve
+nfSBOaiSQ554EHWu5xksyvABYUPs+PuBf4fApV0W2bW52dwSV/4AwwlrwO1DsAw
6HpvdQYFzztnGvT82bluMRKza1dRVvSKjXW0ipoGIq9XSKDGbXIS/LA5qcVeyX5/
wc4ttAmMUINedqdSX6+6ZolJS4GP2rfblyW3UgTYEX6hoMX8+yIP/OBVvfFt54uc
Qz2oXdOiKX8TYAkCM+SWRt/tHs0PACqCXfz2TCSSUQvVDnIgF408Nj6yh4iEz7qh
IX8d+JoJerYF8P/R8vyWWdz4SB4ViwPW1Kk3yhqKOGLOZ/9NpgW1XEfVCvX5Gomd
TzG/k4RM1gMmRijPeoTKjTFjbVseM0ArJ5gKKdpXNcObewd0Lc/8I0LFpgHWyhaO
unag2YmN13Y+s+XtG/U+DLEBl9brFoYCwjeAHADP1/aLZBX617MTLvCYM52xDkow
Qw4CgfCodIfm1twpRD8VepK/j1p7ujfl73vR9h2P+LX3xbkkGOpMFWDw70nAyvT9
93qZbT4c3zZShgnJfa4f1Wny/Sao28e2MDKqrat4GO+4GqITbPuUaCyRR9MFk+IO
T0hK9UGD9f8y5iJciun+vrAKfHEj4WlOHrI547NGgOkzSnMWOJCOm1RPWBeUCVLU
9Z2DH3KsZZi3+IACSurwckSORoxFXR2PyA4CGlKH59S6D7NwjyhU19Tjridfcgjk
P5klrvrZD+Dr7wFA2f37c6ajqaq1GiLEqcMacO2qNdSYI/JE9pM1pCloFtUjeB8r
2NraNrLuaIUY2aQHxk4R2Cqr/m7t8MjyWoRlc57gFFsOYydvv0go9iCX8F5vvB51
pTLxGA6ZOBi2AtlJUtxC5YTn+Y/PSuXY8E7YfVIREx/uFuJHVobwmxaL3GLguK16
SicmswOQig91MfOrL+nil/kDDPMk7olQpcilyy+v3dx1wDWvGArF6soZbg0LV6iZ
e+JWy1Cksj3BcKUllXLqXurzRjOaTbp5c2akvTaHQMMK1f+VYpKgYmOL8peQxjrk
zHMFRZoIYHbMiY8zuq7fLkRMtruOMQVZpFlkFWekOknGuHFQ7vSTVne+b85dYhcZ
Dc4hX12DyQZxjteNDPoOtSgzbc4VzIm4K5FOE04hJxqfZncdMEx7FsJJLzTlQtsv
Vh63vgGimHXDvBoVJ/XNipuuM4ZOerhfNoQs8v5jC5clfNvVET8vfWB7dAt+kiWm
H4yrid6v31wFGXigKgiZuQXgCL/tzmt3DQ01EdpaehbB5iqXfsJxXzE4UsqbI3y/
9eRY2yt59p7bFLBehJk53vFCHx46jDv7ub/QhsohbzlUZ6NZdQCxYCdWX11dZSLq
IAvRrn9FIB6IJHAUm9uXKq8DQRI7sUetuAnDMOrlH3wfKxw18OSv+rFTnT8o+WwV
7Pd/fZOvcN2EYjHoZmJgHlH9MHjP6x705d6RRtzHACzvcRO7bx9HbEt2kPoWDVNl
/AjmnABuCcQy8ewQQWq4JOTPefZeoC0OkIABrE+e0TxpwuhPdMR7OmJIKcZhkZC1
YAF0j9cTOIwSUFmUpIHk4MKQqF0xtWVXwZqM97qB8AdjrVVCw25EuTmCd6PruUv1
/yeIc+WYpd5Ld2TMb/eJb57dBi1JgyrQAvEAz3qGcQY0U/Pd8Zts4pJAGKyBXRj7
4PLwPAkRpTWBRUjF4XudMyWTiuq3PPmCT03k4sks0fJP+Kz38PKfPrbSWJSqc9/Y
rXH7tSANfKRrHlpAzIwdHXbWzfdc3rx7V/PZZiiHNNy7bteNBOEC0dGVzfiPEO5c
UlH9j7lUiYVcdCHhN/pS1yzMwfl4VQXYtc4xjfNlEy4+Nb1YE4VIdaLqsOd9TKa0
kNjSx9sOIOpHoR9fc2lm2e2wDjhXT9TZpJS6BSmO0rGqHS+gsEtIWmLHmBK02YxB
23XqDDbFJfJ/SSUGAOxWRg157Zi+3OnyiDnJHmDWH0eDHpx7WVKiGJjm4f2VRrYk
a8MMFafLEHIiju3bYsqpBpE6mN0pzlnbwKcrCzt1ixTZrkcg+f/SXq9l1KCCmCyQ
jkgQOIXk63neQ/QqzX+dYVUnwoz2oJalLXH5F6pP4m0RQR+Wo885Kn05yG3joSmG
U+JEEy4bxDv7nRLEeln6EWcgLOejANKJvhESW+MpQ3sEKxYFhzBJA9ztfrxaZtLk
qC7MoWTNvOzV5DKk1rhUSZLAE2iSB9xmhJNcngK6hzolqV7KDY0PsdwtvnV23XaO
jR19lu7Cdc7r0H/EA+GVkvZa5Dl39ZQvA8yH/daxs2VprZyM67598EwjbCLpXFgz
F2W6o7l+9pxS5//Rbq2YP+AtxeYq0ET3KHo66l77lRtUgl6eLb85KGnmgFjr6/0I
J0qAeriHdHDKdnK5khEag+wqI3BMa2sGEk4YhjysROVzkGkPuUGuc9CHM1/VIdnV
Fw70p1ggp6v1z/gJgrKRdCVzomvY2aE1LfrsbznWrjvJC033XH85bKfVuQrmI8C6
Kmsuf+KqtKXriAFjKvkcOgVwlwNU8p4F5sTpYNbtpKmLVpqpsHFH2DzLSyyMIqZI
rd8bwZR9E15JhfSf1wKqKDiIDL/0Z4cct2lrRwgaZHH3oTGnKnCOVDU9R3ZM0fsc
NdZ7lS3wpZQhk3SxCLWuC1BiNNn0WeKj9jldh+UUiFBkN5jFFKv98D/JbnL7C8gY
FS+4qyvnXzFB1Ph7rwXoYMuXcCf+M6F7Wrboh1vz8FOAOrwuOW0Iy05CvyMORO46
c4ezR6Avbxz2HWmFSWObw09k63mP+T9CkX1Fka3KEmwRvIe99pqYX8e+Z0dV6iWC
4VpPDEGof16CtFrPIKZASHcxfo1lYkWwR7A+gv3yUU9eQXXFh9EoId1i3XPmOlsX
9102WKtgnHJKnLZT44kyFfayFg83LWnMBoLHxfWrlhaeKch9yERrbk+EMc2Wb1co
B4Uq0BZgBbuVj5Wzi0LcjI+TPpO5749eDk2k5KPzR+QjevRKl8FOKuKFWctHNqhn
ndGkAeheHPJhAXII/7oHuFrFuhL352NgLgLz7h0ldEi5sJt5NMuc5s+HMSXZQW9j
vq+7e/eJ0mSJNraLOTujbaQEFTmf7tmDUmJ5XHuafXJiNajqSIkhaKM3Z1TpalJ7
l5paVR5RMTJxaJIyUEdwoZ0KeFUoR9UsylAJCnwS3kjFmN5rMZ/9Qdgm6WHQrlpE
8vcDP81QjCzTZJ+EqcLERTUlqL9ZXmxW7Imok5VTOwLu5wCTaOVY3Yhrj2ZgTWhs
6OWq4VV2xZ1LDxfsZWdomddjrX/rppCzMBj6ChsuxXJXIiNVqL58sLW7LC2IduOD
2mHBy+bBRA2tDHi5btCFTqF8UdyC88l+PWct18RifM7wELvOpzWJNnZIcO+ZL5oh
QQaEMI5CsA/rRNCAHCCxY+d9014ameHk9RK4Eld9e7gMhO2bNP8mLTGXw5ZbRkwO
O3JcG85W9N17SBcF6EhGSgt8LKYPmUxfi22H+xjwmB2MWJCmeoiTwqli+ZLW/K3Y
4IG3bPwalPVMwPuyo4hvdyxMvl4OAzayZp6EstxDXpdZlxYSTWh1qYDIEa8KAS1l
TPHGqa+7CnizzKd9RNrT/TDqtWbM01OC8i3+onrQAkGNaS48izrQZTf/Dos7ySnR
dkSuJQgAsXlmTR4uIRC3BcfBClVADOLGRnuRrXh2/PYOpAXaNmSh75lKzrlkyf+h
21i29PopLDMn+0f4HkPDNBjwrExQXDW8YQ1kj/9ZS2YfRp8Zy0CXbPfB+aXiq7FN
9xYtguIcDvZ9mVN6qrpNSmVEDAe1NVYHU4mMWBKURdV4h0P6uzluVusBPQW6DmUy
SgUJpI8D9ghFJVntnPedfY8zH2iGE1IAiPacNkTk2HAhvX37pswuEgztpdhml1L7
0KPQzNJ82siKSb9Lq7untBw0NCBzPOKzSIKbq+EdX32drnG767997zk/LWs1zt7K
oJE6BtFsG86W3TQW9JqhEX8Ble/uq9lKkhrAc7tQ4fLX1KNn7B1zStLB24AFtXfc
ifcW29eCLDiHFq0j6HN4Kc4VaOYBHBa6sBBvtLjUO+7j5TOYbxdhg16mt9IYDivI
mRwCi+MOr0OT/p+f/du3zw==
`protect END_PROTECTED
