`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hwnMsuyd2INN757E03Xj5C9P1936EExq8tMqVeXZcwpUt8t7oursd+qliA2V70iB
hFSmrU/sD+JntTwT/si/EwFpAHKSnE3EU0gnGKAU18cG+OT1giYtj/JgmwYw1QVC
/XZAo9lvN1gg4N/9s7KdgWQV5KMhBxoSnP7LDoKf/e0Vqq+ooE66recJYFVCx9/Y
G0+WoL0HSEt1mzQtrMKomd/QbmcKHFVAl3tLx/WZeDTikAMdcwRdkVpOg4WDTtDJ
hKnsp++9c9KQipjYWma2HJsK9ddnPYMfi8zcXRoxNCA8MQEWFF2iNk5dmUI4aFiF
nqiL4wpHOmt5iima/xOm1E3cE5aafv9SHVVVCecZni+Hcrt5M0fICrtMuyn95BXf
AQeqipEpVotdzt0Sv/ATjvuqi5MeTQOIbBsXcN7RjWGajZH3mMI4qWRGYpVtYlYa
nBY12uydDeYKi4qZFkkpc3t5iHn+ve1e3IYfZ+gf9a5/NTTfoQRjj3tP7iH5sGEh
HqDz2ciCsrzlSRokdv9e0xSQWFh6iG355THrtwMGHaL1jBjZRCngED3amNTluKQ6
rAbReP1uA0cETVBOIRv/p52aQvLNzmSb9HBUurirOAyLU6Dbud6oEHCXc4Qq5bzz
4yxEFuxwq5Kj/M8dNV/s3+3Op3vwenoxdXV2iM/jyp5ryl2cuFw6ObiuEL9AuTjR
QZC24mtIWtfCPkaZP7PGT/3xEBXQ/B7OP0Ecf8v1avPCAPhgJdD7CgxENvUCWPWJ
JoRBJ3PXloIWVM8e+Y3rCiC/rmxtvzerQXWbX2iUDMWcuDIVfQHpFzywbBKstR2B
aa64GDKQ38VlAImk7AS8SXZVF9ymPnIWWDrJVpFW+NvqL0GK8fLFXMAubNh7VUTE
hiDkZvXmzhBAevKx5MMiFGBUOktU5e72cGkVKdhTPI8YYQw3EsoEirRnqi3YDrzU
ZglbUBTXjuxaPeR5uPtpFQDdgVmCJ/FBFSzl2hn/LPv0KDOVO9M5pKa2vMcrLHNa
ipMkUpu8wGhBN62wqCeTeVjAe3MrQxmbVKkrYSfjl02n4CX19dP6SWVttx00khY8
DSQfy7KzYlrfKTuZya4K4xe2kkc63+GY/lRw5hGz9wcg8iUHdGdTJAfFZDopAUqI
KbpsRvKR4KZAk1bGYYBdZ+WEoY4RdE0zwHN17abnPSdOfiVwiOpAHVqWgkFJQeUo
r9b1Jc8LOWmB47TBulxs5pi/438qXHdqaUa7HD5e/iWvCfL0aLRDvdk3/usYEMdc
20L9NT5+t8XTy6r9PVjLse8/BJF+29SXz6BVhcvCbvgkpHaU4spXUdgNSjnrnc1J
Hb0u6PRJ5ZpHUK7w1S34AR7BZ5bosXREKpm4DAZ7sSfzwyWzgfiYYBSLKkbaDo8s
Tou/5S0PLaM5nZk1mONJL43yl7QAHIpbfVhFMCfCEZ51bQhulYP3EhpzRov6F2CJ
bFS7mo6aP8jUx3/7bN572A3D+Vut4iwkaEg3Cz9lc+lhSuBH0Oq93pDPyt6vEiij
50IhC9aZEyJV6ozUbnJoJI28NKHEK/ZVyAmFhETQXQVDhTydSV+IhygI+diKKDMe
5t06GssLwteMXt9EI16iGt2nCAE3QTlUrR25tcr9425DBGn0Tjf19u7OUFn+8bui
HvabgpBySIeukatm7pGOTWG0WI42tvnqlhz3LdzkEzwWgu+c2AyQY2574T0Axmi4
n1d5AOM4e3GG8+eFpCMyFU87qwJXRIMNI/G0twVaZOPnGlUFT0UFK9qMaRM353lt
lZHnxXJSM0C0OiJBIvxBWFP2zQXbEbfzQM+p+pu1JWxzn2Om8MFiH4T91dgCakd9
jLQSk8sRLkGycx1CFKChMQwS3iPn8QlCnc1C4FSLfXRX7ym54/wMjqkOLfL8Oeav
nkTkVxEC4wXlXUl7VZoswqbCVZfNWyLxrr+m6zVRtiaFHoY7MX0Tk0PTzwykZuYK
kT1jR9XNRkPl6hds4hLBBTwQyw7qrK/SQ2qwhe+0mEhsvZdALzVQz11WksRP85pO
gRrYzGHA7Np9i9YRs4cu1YMlfEEWBVcl30L8oPT3RrbjF5cTaLABGk1IHgi/MKhu
EV2L0pGmdeoItCzAHA9iLm2tU2ifudAKCSYA10Cf0mkRlEpfq/y9w/uDELqap349
3BZ7JdM+qxgOv7B75OgFihEtdlAh1Fw8E9QCOKDkxe0TMDlpIhksod1LodCj9KY4
bLfvmna43tTu4mZFBTcxWlwLZR40Nw5hygiK+cjnjgq1/XsHBELwA1PfBriACrWx
IbUMIU4cOi6tEA8i4Kytat0eWZzuP/l9LZJ8/RikBEEBzPeB9+cqF3Zyq9lvKtd0
YuEhbNa1tsNj6WUMUj/DHEJrS1j3n4sZw0CfWxMlphxtsTIV5+t7qW5UVFjPo/1B
ytJfzSEpuio/RNM/SoZerJT71+MMRTNC/sydtqL6FBLMk7AhwV5iPWwAhnSqrjIh
arElfXwhsjklNZ1vKF24/bWG7NnR8HOSxb6Bk3kLOCJ/kJUBA9+jIWsEZK2Z63vI
/LxCk6EZcrxh2BZrpPhho34FW7LAZ1hdFZ6iSXWhEutLbnnGC+kpwUN5iGYdxon0
Cn2OdoPaYrES1KsIzHZphhW6kDbx+xJcEiM7u7zvTORnAZJx6K3XncoP5Kzg0i0f
HhMMUT/Lrwr+oNHmc4RLv2/CxWwUXWOzQowP8gCrJqT3O+tEpc8sT7zKC5uhbpRl
eJvl6E6YLUXAcuDa0JKF+16PxoU+xI1tj04xPI9NwuP7bozWC8/J+Uhp/DGl8GZH
mjEbY9UXO/QpIH8sq1QJkPZaMLQJYwlWuucQbRvLsUx3QgiPBKlPgancNJXzG3DY
GmxlgyrpttZHrg7swlC+rjh0XBzzXtzKibvaqsP8pivsCHekyhqKZf9fqKN90Lu8
pGXVUJxrkmjgpfEfT9RBbR0z8LjOSFZPi331f08DHua3C/cnJVJf5M/dDg0QjHc0
u7OFOjynmKpD0sZxa76fxg2t048RZIQU5jvn5Njaw97tZUhflIJ7+gXNQkWg4dcY
IXAAf1+sEO2nqjlcJ+Y206lUd5ynz4iZoQAAvM+mtCjts1/Ub4/CZp2FDPsqoyPI
MhXtdx/xs1KwBCyl5smLl7SnegTNyuJz3kxKbgbDGQQIDkmmk2qQjqBeLJsM4KZo
o/nt81KnRCgCNmKfgSQqO9sEySfkT/oSOkL5ZSdpLmI8/JjCfPHmuTTuGSfK1xNd
8y5exzJdXti17ArlrSkzmSCJJYifQmcowqvjMUW0fR1ytj+7NKE9vsOXQb6LM7yF
44z0dfAOSncsyiYhPeLadkmaSPeHpHBWx5D315HMT3Yul4NY7dwoogZ8gb4MsKlp
ONDPylCiACD7RRNAlGdnrWj+yh9ffmcr4+2Tmhj0Mb44CrGt0FVcII3Qjqc+MkTO
G1KcRDSyqyzqSRE83ixjMRDqDHfIZCVFjrx6VKUF2RNcexU0CqW8NGDJD2/0prDs
gzG1vo+HwUreieLZSFH4AvZmksNJ+JYKvTbf5yWHU9s2p7sJcY/vj3tLw1JpgYUt
YXU0XumnWx+40Px5litM0v8pmFyYWIeXrt8VuZJ/8M6Loeb1AQRz4hNlJGy0cpnD
bKcpvNtpBeXE1PancmtwyXjkY3b64sVf5p6q0lQJntCZYml44A0HWOraP90BPSI9
aBlfSL6UNz/yePXgHEeZk+OX1BCqKZ3QxQMgALr1vhT/DUHEBL2eOqwqzEpam86D
m+Wl3mFTOSAuXvZwJdK9jXKiTHMCuqI0xezO3jGryY8p/TEmagG7Tml0zSvscoeR
IS4kCFoj6vHIGI2GJ+o5syMDGTihjkhcKvzfLPH8zjm/BeEcRMfjma4IYkTWaMea
6AjlUsJ93ObXxPFZqUWUNAsCSsB/xpGgwCmzBXyMmhizTz3jprR20LiY8CklgeN3
3qgXxjv2QlEQfTXDs3Kyzqvgno6PtUh6wCiQUCBXL/oRme2dpZ3Pem6ZBbcK/iJ5
SIUeboX8RWFpwg4xrnx19BGt/eOnD1WffKR3RM2gajV0SY9TQlLS+YpMY9XI4ynW
Cl0T92JarejfhQO44A4hPHxfN8iuMgBDUHqQ1lwy9HEKDsqAIyh7OjWGVlqeKx0/
gfU14K+TEZ2Zw/JSlXogkTXMJib9c3sJrvEKuETnw+6bEKdDKpF9WfvrCav8N/sf
snxKjbp2HqPcy+0fvrsvKiRTeHwIF6m8/civOgPizuz+64Hbqt+De9yq3YACazRg
V59Y3QVYTb1KLXLxhPiVLOGyWgUYdyZXV1j2lAwi7hdLxWnG5+aa1IhD4b9uhwFo
MlkuRsfR6qoUOqEnwrxoFs5QSGewY8pRMDI+fsE8fd6URXiEN4hcRF5j5xdjIsMa
Ilien6OQa6x3p1hfXLRw250Il1OkkI6NjBjvRZBQ/fzvEi+wFnVM+IAFIAZrhBDL
+A3gDgZd3abVq7WFVw2NtkfgAkwq6bx9A1a/2jwcLfoO5t29VvUPJjQSF0fHii4y
R0XV8XvjfZmpvPmBp2sDFZYq2ZH9ZqS1ZcRZ9u8yLd4SouWZGt5DbO2H7+QZEH8W
atC5QeVaay4ecDZx6dJzu50a3PUC+HBCoLGZVOdxH7FAZVxFgKyYA0TI0QNZtUi5
CQ4aMKTHYHoVXvKIrQgt75bX26zshNO6CNwKjWOlasDqptzN5ZzzflwJZa87TrkS
thK+3nzUs98y+qsjGrPLRH43EnsL+3bhqPqsAZRiQ3xs8cMDXbkwldWDnpTdGKop
uO4Gss3bWeT+NsN7/+JUKg3UIy5DntW2aCSkSIBC3ZD8T4RguTzcBn7nMVwsy8N2
eoqCtvpwQv9mDCdh8zI0Vm4/ZCVB4hNu6ORhCREmuYjdf3OtHdR+t3Tr61Q3Mh14
C+n+K5i8LQWaUlBBraVmRnlfK6lL+ldMZjQsrWx+2EadZo3K5PnLrR4jICWnbhLr
H+9bwTdcqYuXrAkEW5WhjK/1Ynqg84MQcBJTv2maAIQNqhS/psk081fX7HUkZa/X
yyV9zt7ZVKG/HrR9dRbp9uz9z3vVI+FZb/B0rgNHiH5uUdElk79pmkZYaI9Uk0BB
EE6qqkmBUpPZF4SYwUdlFPui7cg5dumumPHmS1j12awiCUgMo2Nf2m2GhH1v7bT8
ozg+otKXg+KAeJ0LowrgnFSfKUXDFt6D8q/Z4PDNk1I+LHvATOS0MYIuFmPRzmIG
DnahuF4Bgrpf9yqsE+lJIPXUf/ds8b9uIWwDKSVgRM3Cx9At0YYvU12QN6CL4yaH
/chCNMIIlxjxJMYxjp8M0sOtEIEl1sl7sDhodVV3PcN5m9DtNs9RpvqsAJijn8SM
lB0FtXCbkjkSbnLN/MKgSns+n21sj5ZqeS8rrBQgmwemIrY8tEMCuJAVTJK2hp4P
tg0sjC21fLGbM7SdzF9ybYq5BkrOQ9Genfl82IIMT7cioxB4H9yua6CFEPRICqw9
p2n93o+q4jcRm8k9Ub2sRqBVCzTYL6JIx74H1v0FQD/ZPeZWQeKoZqE4WVq9ft5K
+gsovnU/mCoVFPZhhWylb9xzDq7aqG2peRABoxRQNqnkXTNSFvRWrnsrGNwLbCz5
02h93W/aqDRt6v2WenSb5WsWQatVxPsbWaPMQWcGZH4nMdHLo7R6L6FOxV7oYXaS
Kj73ZkKbiDRSFc7b7KwtUKljRZ5PP2rMH3btfKLEtBEDXgTiwLKNHcp+tmFgCuJA
QqUIKY+aEi5x1+1ogci5PcUt30/CMYDdtzVqmUaheORFSUF2YDi7cLefb/B3mcA5
OHvZRkECLP0BkypMXctvHu/c6w+yMOpebQoqiY7/UauMAV5zYhA435vGNFQeNKPx
SWvuiiCOWSIfhpmiJMI7QwaYU53j4O2bsFkN2j4TEj/zthF1q0iM76ZXR1YtpREc
impM/lWmo8yJYM/7Hy5dFx2yqoSRt0GvfjDPfgo3T5RUZqm/X7YMr+VglgQr1KIw
NpI68R8D6PcNzNCW9YhndtY2995LJuRcBaS7utLVO+EgTO0oaOnMyYBBQ+oNwrVL
z/UXxQh1Y2Hhq10f30xdvW3c/eDTYi3SprtSpzyDw4cb7EF3II9eT0Y4F/eQ5/Td
eE54B8WVf0v+TcB8c14p0upmeppa0RFF76288ghxkllt1dFI6luro9ZyTxL7//w2
DtsXShGRi+zK7XBskfPPCw1V4auNbZ10h0gpG6wLmT+s63l/rtxFpb02ebzves0h
C008i9DRqUjgnlv3A3QXtrVRnidoseuFtZ1JMjvbV+z4+VAD+ybl2LaNh1/Y9K1B
CZZZ2Mq2TOYPzqlfdNSyeOoCUFpMAyG7Vw+kbwDEsG+fQV7I402ApArbumAyfnOx
01hVNBocSy8uHShNCVmxrfYYHBt4N/xF9gwOwwG2JXQq5Ww1NdB5yemcBHuSnkef
LCX2QQKm0t7sbWKM64LU+DRyBN7X/TTCwauZsU8mJcErXqyhqs27UM3GYmQEyEWL
Bb8OELz9b/SkYRBRkLCmKxieJFSJWHAlGw2446M9dBCnYqOwP49sdZJtdmhGK7Lr
Tw9hYgU8xyqeoKHLxVv6UcMl3GQL4NETg+eOKGz0fxiBDS+VE9bvG2GOw8G9pIwS
0Vpf92Tjqp+iqfYwnibi130UsJhN0qKxTowqJ4eJ4yO2C5eZjiXi8We2KGG78XHJ
uXKezANsdcMZ4khQJWVy9b3ZDr7JJdl9uUARZcxR640/oRJymQDQ1H8PPxje/XoY
NLxcymqsnD7fSO36/IKQLMzA+7g/Jd+HcGzDP0Fk8KDk2UDROz27saczbHTaq1xx
7z2I9JEO8FtSsrrb/P/+hR/ib/zvKj0T2Hjf+2zaaSDNUtLYh0MYPCgYY+2ASOmT
kdW1g9/O58ouGc+0i3tPOlPwGrqhbpDUEygaB8uK06W7MnpJYuEWpkQ+4CdslzBg
3QMckKeCAMdLTqe/PNzW0MEb0MDSaIM1++u3uAzLUIf+YjDkcx+phB7qFvTCuqQi
p42MY1EzwhL4L0wVnOY0zmV2b0mQlIS0h91kj/KStJQFW9IO6qNrC+5ikWQh44U3
w28UW65DvYNM9SUmWdGFR4nnaxz2MgGGNk9IrExKiZrBelJb1FIiZJBdIattDeeL
QCpK4l/7NZB/pfBoN6asT9lJdxFoNCuRGmsGH8V7rXrP3SOvmm89/rJdF24Zxev6
XcaFdduzNbUuE0BoNeos/yA3qeOBWSzVkBYB1q43KW/uGxQIf78T0P0Y1Yc2Jg92
y5NgecWBcij+RhKW8UDrKIeCoL7lFHscPs+8rF3FalsBd3Z7Inxcj4xBiiA8QbzG
2h/p1bfN/Ta+48DdmfBDoECn6LVOV/X3q0mc5HsWp5prOgjPd94CElyzZQjEo7pu
M/w9P2pq+4Xpz4sIuXhib0So7tp2U2yb61oYprACz7ULqPR87uDc3Y96XLINuBga
JCzEmf4/IMKjfOpUMyyF5RNb8DatWndSE5O1QXkaCXtuVKLFPibfBQRB5tPn+wsC
wAP7D0HUPE6R8BOwHtjLs/jcjItfAMz0UA8Y/t0eddi+gP0mWbMizyxxJ1+nUWYc
OuR91lR4ZF75WWLcRpC3FAHqGm2y8hA34Ioxx2EIctttQWlVPP7A/fwR+eT3Y1Jy
SY1QcgDT/+F1qXqiWSaS0uXkhXKhIccgG2R1aspq9uL/fHCVwA2e51Ni4wbX/HJD
iYCJbjdZv7J5PmJslAAOMozOjsXPY4uvAlEecrClCnhmtckJV1o8tDmPcIHdvB3H
5nyqLEWhMhihNy9U4QcgZnEYFgcqhIR2y94R3o1WJJ7LVA6tI7xGEcShT6devy4r
UQtzqEnczPiUJ9xiWaiHp+PPEgZ3RX6ixMMsK6JeYZ5QEF7+xrYbhTsrN0f4vtWE
3gQjnW9INgDJbVgTpmE9nPiDqK7XFrGLxtmEfaGBsZfoJs3hHy3pN45H1ld4i88d
kaPUFFN7t5lymNV9EOtzZR6Xwl1XMyoFAYPOZlXJKS9owmjdmwAGrzIWTp5i8jCi
AlBFATjPh5t2EnzuBwraRR5XCusLQBPl6vmjH4ka5F4dqdqLPWnqkzBBXHBhNsCr
lNUQSRpCgtN3wBAFYHipa1Hfd4LkPxQ/CAAkb6tJTs6AEpX13pWZbFAfEcocBcqy
MsDO7N95Xu/hXW1JfWHBkpEv4aSoUA4n/Rb6x5JDSZw3/bmJqUiTg8WQbFyLwZBU
JInp+/o3d2wi8e8tx173sDRJLb1bNVEHdpcOyaoaK1K8DY7XD1GCdpxPa7FVDwYf
wuiQfo6gDDL13AJj+pAkCTIEqpX9wyOmnGw+pxG4KeKoYsUnDRWd/HmaWwHJn45+
1q2Z1c8kxCWoaMrxjE9vceSGfEWzNlUwbXv1BvVDel7QH2WcsvESnM0uBIKw0UnV
ViOyqiX/6lUWShFsg7hLhikGy3QORySx+GAyscCAy+MWV8ni9iIE37Z5pdDvJeKW
pDhumk4FHLuaiglaBo8GUfNgKjTog551DmesgrwIa9QBsWA+mU/x9Glq5aBvRKpC
aw7TFQFUdw6Kg+sA/0NmF6SNl5WHpZudi+cu5m7oaHzeBVe2Cnbwt3ID+jflfZHt
JKtgMdZKIzzBGVvjfwR4SdumTNxQWqAj3YTwBbZzkh9wqrc3FUreznelZkgkIf97
feccKCId0Ie0sBy42Kj1qgvMOWO5BRB5CqzUU4ZebEFq3/2fV5F8swX7ZVKmopgr
mt7w002tG3pGNFJgmBH4xjlKI3sT1nWJmvgUOTPmQoN0TOJiHSmKqr0PlaG7buKP
qn9i+FwcnuGAbJ9VwjxqacF1yKGPB51O8zOaBqTDJ/KpkvpRlyHys4JUFW5gBv/L
B4a4LtAuZXw0DRgFbso2EciY1nG1S59FCOkuSlPaERiyrJQH4G5A4ieJacvfEi8F
ZFAc2TqcbQWSL75CLYYvmvKWKd4ahI0c11Bn5Jy57pGwxx8D7worcK9MvEfQVrYP
vnP/B0jc6vYNM8fgwRWsY2WIEqzQhCwla8j7naTu+95qo35axh/ztrNCE42XUAIr
9JCWyQ4pEaFP/coXr14+ux+4MZAp/4ST3gKrXdQ+nMvGUjV7zzNNtAM1OHhpCeAD
IL2pOQ19RUn9nLDCvzBC+fJQ4nR7Gv9r6flH8vPN68oYNp5ZX+fUWHxVGvmt6J+L
ETFFKun0nHNOI22BCmi9I4J2gFJ/Mhl7JDUVI4fPTCJgTEcazTtogI9+UHbgrm49
KoK4+xUBwvjWxqkz0Z9JOtUpKnd3JTn2pZLja3UpF7gzylQFDbrFhzxIGfGFLOWw
YLph5Df8nmApqfJFxb0pKMn9NjIXvXXhRh9Y6acW+N/vn2Cj+McjYrYnxFUAr1bl
wcVOpLU0PigJ/fUkYAqD3hWdMN45z8MqAmGhmhpWab+Bcreu9gbTZDwjon7YYklw
lKSIAluMu9SnWif8aAZqGpoQbXocJ9N9K041irPLlzs5fxJGcW8YZwKkUwxGMIgc
ngg++DQZU4UPq2aJ+io2XxGVvuQWLAj4tNDrUCjMQAW8lKp1lmRzFMVQVa86G//h
Uw4OxTY5qAWQ8LQReVJhazb84L0Geuwyj0d9ILDsUrclUaTCIf0v5hLcibGTLMg8
KS7NTzbFF1Q0okDDujhm4cDAjKrZtd2t589xtF40SXiaW9RqMX24OOiDGpWCy4ac
ti76jF6f2oPRJhx4XLU9Xn+IeX2Mky5LIT4Oa6KJbGXJFdnPBT3+9jEqdXd540Ie
8FWs/nTFtcPkmUpgnoWNmjzIjd+82RPZN9NPQR2eBEL2RfuRHCqhL1rpAmSiOMSt
XLe6k9OVUA9ETAyQyE2liFTAfAqKfsOztDmn5qcSDgEQHgrAcm3lbRqupCxE/1cV
BV1CQyGyOYwZx8bhoLOmFUv3xfF8PyYQEyvH16zuiap4KybPhkmXFhSVKHvxqh05
nnP15uDRH+kS8qZdTuh40cmHAFHm1Lo5PO8Tn6h6NDnLijryqO49tcZCkGDPQuNI
2UD2yPz3PgnHfj9c19iyw94IlDq2NrNojccUGZWNIpRysKztqSbOLPiZ0AnAZDVx
IJb7A+aHqJV38g66sY9zXKx7RGgtIvukw51szREZ1z08G5c31Ps9uv5nRAsuy3ug
JwvCHjjb+v24LkMURkRNOQqaUpVg+lDi7vi7lI2cmjESkorrMIG52MpplKRPeEiE
O5e0bgpVMMEGf/PCygH+04Ujcg2ihaXBX1nr8rMtIAvNlwhwobgKQnrEULn68S5V
OhLRAUI/RzJJdDODnQq41dEsQrZGJ4faX+KU6734hcd+jWsPK6UA8wm99skXIhzY
16tOUaeLtVYofnzZ4cTIK9Jwy+7OCnJvm+NUDlGrnWRMhqXhh4Vm29W6Y221BWFZ
/OLrHcSlczQODNfBaX/jPKhggtsvwERDzCisid6WuxqoeAkLfEAucI1knBot6p3X
zpKnTf8WGP/rBaajIjq9k/WXGoExSYOO7x+DLLl+uMQcJkHimxzjv82TioDKdn8B
2m5FazwGeJw1moKIN6LzwOghPT1Jedf0QNadW21MB6B6RHqWbLTO8oRnhSozDIxL
cp5djlX6O5/U7lEeBcN5NVb52ZAszOFjTMt9QyUytFRufODhhzjjc7Onm66nZr5m
mp8O2pocp0j0gmHicpi9g/0VGhqept+wHRIzL2hCDZM37h1wGGnw38rhGZOgobCJ
SytjbtcO1gVUKcf/pG2IGJUR4vRWeZaloMUn7k/I/kmKtUvk/DV4nEVMIvyq/OxC
93sXwsVqADYNbUTn0E1z3ZFoUYX3urv0j7w4sy36xEzIaJekTvDJVT3tJFY5TqQB
pkl9sewOKJ0YITdjXhD0y4DcJDvMzpCeIeMnvbZGe503fhIQ8Q5f3Sn88UVTv7Vc
SdDmighBV9/b3ri7otRQk+Oxw1Hg6ZkWqZuwt/ylHUN7sFHJRjCT+S5K8+tyO147
YXyD5LZI2c94JdZsmFdwIWx9tfVvge8DR9sTm4BQGdM7f+5BoTf5Sz2GtalXRbZk
ryxLY/tuwWVMgIM/r8Zsv5/ZO3u44vCJXYss3SUOBMWto+OH8rxPHhs2NVTvrUkG
c7ANk6SYmeh/khGAp12JKqOfDQoxDlB1iTzyJg34FS0YbqoPIVbB6bhJHQ09/ntl
mJ6yHd7DvXKPIQSA1dyzmO6pQYmE+eUroxaNvEW80P+WaXTxV+aHKDL3Rie1Rhf0
MmtH/KiV2xlRSMbzlHWw8FlNYQnbVkjQ5F6gKTA6sfbix9K7smnZJ6Vm0HGr24d6
5wC7IF2DL5wfOWnhu+VAoWbYoDP5yvvDUPgNqhvQ2ejwackBihLIMR5sK67w+Ibo
yON++kOCeURFTunmd0AYEpp1E8zw9cCz+da5M3dFHvZV27IBsHLtF+8VFC//pY8/
z71fi4rK8L9qQfsb2Oe/5ieVU4hCtPZ8/mL0sBz6rUbVInqnv9R+iApl4AkqqNS1
rOwOs6VtCcpC9IoEfI36WyJZnS6BathNoXISCgXwEwm3vrI2LJYJ6/xzyyvoOlU1
/R6fohXI0b7ZAYOf5e0Sg3gA+NCFuZWPgs+D+7JbXjcMfain32D+z1qlUbsnwtSp
VAGWE9E7aY1veOmNyIsjen0Djp+MVvYStAPQxUjk3FqOJiVIVllwz9G28eFcheNa
F7FzyqyVebq9G4tTVe/NORKce2Dmt9bP+yQxzBLCwiG+r2OZ7VSidOrjeyj0ATOh
tw2lKvy0lsrX/KQJzq3VgnwWJ2NQCWZEKjkBTJms3hFDrjJFzVR/j6lp2Rm3D6fM
A7mIsP7RurwOG6ik78eF4gTXEi+0OHcj3FEfPsTP3Pq5zB8s9MClk5VeBXl0pgXv
z7X0BGwNIJ/GSEdjUnpYgvAZ1UjKXaXzxyKiWqc3gdxwCV/Za6h3C/lkSD6hZQz2
TsIK95DAhBDpAglVHp4sMv+hstPT7QGKyuLA93E+nZbM8Lw5UpH5G5VlPslUmpPD
HygfV2QpvthL6yv1W/pQFL5Df68G9v4+4sK48Ccmu/2FODv4PH7dDv0edMG7cqBG
M4leWeM1dWE/tdQK6432pLS1zdiDfMxr1VV2cVXKOINt6+yzmlpon3ZGTcfOdgHq
GyWXR9r5sixODYwWrygr7PUt+DWqL71re2MMqLj5+JzjAiFpFRAHubNeqN7fPw5O
GS351zl9HMKg/gLc9I5rF17LWbbgxVY2FDBvbSgB9oVC5cop07dEYH3YgGXsag1H
Eay1keRiWYvgfBSnxSlI0Hz3IlcwdU5oUjjB1OxUXSHAclGfxUug58mTvlht3Hmz
mehc7dhd/9pUUNHcVm4AkKHM+k7f7kUcNx5ATia753hV10s6MXiUgrqB6+T09bF0
xbuan1Mc8moEY+ZkA1OELslW1SqElWljvv0nHegRtRVAXrR5PBDeGPWMT+g9bb26
qg4gRzQrn8uV/zU6cBGCscVyN+Wt7f7Ahqkq/zJGsZMtL5G2PiQK9jBa18aXD805
ICczA4LlD6TMxw+K72T5tgXQ5Mm4u4zMiKG1CIyW81NBOkxZOFs+8AZf0t80D0fe
4CEUIaufHB3X4xtE4WYC+3gQ7RutrQb5K7rpUz2zYx/vuud9AJ3WOfyaLrTHqD/L
XGB6To3MMEx9eOeKwNMDeZVCPjwbAW1zEmDi0F9UkHnkQ43/Ew452pcLS98ZFApQ
20Sc4pfoQUGeJXc+s+4axF5K4RLtxPO32YfFhU+KFItOodK6zEVPgbJM0ZZ6rftf
ucVz6G4NXZ+L4tGkrO+ZI/xlMtBFdHiWUY58RDfnD/Wj98U13jiRMnohi2X7p+8I
UKSMQfiynnTv6WFeQ68K8WjuKVA6e6TVlNnCtNKLHxd033Ia2pbg5GvEyXnRgWyg
X137INgDE9LulbmOAPNir1mjSdHwsKgpxlxZxOrfIN1GBKsYvgZYDLflzIyL4r0F
Ja1qlsi6LzRF+rPoqgTijsCK9tdE6oSlHN+9uNkpgkMzswgMng7MBCAjmv6e2Oln
j9zR9dmjsLZI+iX3lIKZW+T5uSW/IZViNyStcArvfEWp1wsFhLzBQQs1Y1EqU1ia
UC7rhLYTPZSKRWbP7P2pSWdFbyHVDRadk/8PpK5N10Ey3Xj70fbwubTfpUWaYpgs
JTsHTh+4QqX7bYPt+TM77OS9wBFYugRXF74cq6PD75DVdy9C3nayXQQGXBBSYQ3I
Z6k5g2Qh1Ab431fi9MynzIOfj5jpyTuxIzZpY5nGgazKSKtDa8xLmzFcKJH9rMas
Vqh3oUx1T7eKh4hQnb7EZ5XqRO8l9A+SxebnsdYJJLaWHp1oh7bYLiGH3NzPl3S8
k6fMRGHb2pE3voJ/0EzR6GDzR3ndBCOiLwjlmQy5IKxUTz2lfeFRd6bcO1RTmkGJ
VXvu+rv1AdIOMOJwOAxLEclgYJkdUvlF9othuxvdl2EGcWPaPpSgHQozs7EZSTtu
/DEUndYT7qyyTDUV3At7zpS6zy2YTPzPCEjOhvoB1UsyF68khBHCaei31gF4YNcU
tw6RmUfb6JmnOCeSNVYYtedh+7Fz+Bj0GZJsKAUZ8YIeBx9MV9e1nw5+6CNSNqP3
uBHetd7wK2d3v/en1W0tWdY201a2zGWmn15fk8ReXYR1tmmklUVt7LqE9h9rrCaw
wSF7lI7hqOYr6VBW7GJ8tb9a94QZI5k6C41y5TK/c3b/4F1BFjjdc3qi7hSskeaV
VjPuBw83WxITcO9sNx276m53fQ7GEdoK1q2Gb51m2B1RNvpNUm1iZ+t+GhBnbAhM
FbZ8mz3Cfv7IGQC3Sw5rD3+E+gi69RtE9uDTWwG242AHO2yysezWMkd5srWm9X4T
fxmvQAfFfk6xHZOXkokt8vI4iVJJTNzRw8Gj5Rp0txV3UtyToBUVH/3+M7kzT5wc
SLEHFeficTms5BbQYNorM2UO9DtFeXzYWuOs1TsE15I53z6v+AeT4P245iKT5dzk
U7/Ave77J2aea3dpZKsuj/dTTi7ehjH5UdNBxY6jMO5iwTpXvcz7tvzUgyD9zb7P
z+uzOIyRqqZTsp6zx1RRqNkZIbIiW4/OArRqmaJHrZCguVoggE2z8MyXNw6x/37d
EfsykAYRxFV8+r1lhByqZIcS5F0Jrs/CI7o7wbLtNSbLLlCd2WdPRAG66lde8XH0
XgRiLaVydxISpmoI/QkPL90zSlIz7iAn3t7xbgGBPpLJKbGPvScN/AkVN4nQnN2G
z4Sz6RAww6l/trnk7pVS2cgKo1rwzITbN2T1f2V+nRiZjqpAgcj+vF9tlptMoLwe
Bc7r//J9HCQtX1ArYFwMjLDjvewi6Zo6HN3Ai6ARXwxWSo1YnxSWZzRjqCvCG+dk
0AgQ+T5O6DAAHxSsuI7PjFz3PoGiASrIcAyeWCT9S68CQW1h2SQl9unfDzreSf9W
KQzlaB1ENsCgqSbyR7wPLGfX3Q38Ah0FhjrCxw4qmX2WNbeWD38NO6EycZgdHRZS
M/fPy/gsoM5c/ea749lHXaEuemwChABE68n8v18W8GxRxzJRGRxfbiSKcfLaghTZ
e6WF4d2VzQ/PSby22AGK730k1riPreBjGgVuOeFSCEfH7p7EG9jUA5n4BtHDIxlQ
mn6bz1tTEfFCN+Bi5S9R8o7vMf/hdO28gA76xBWhcW6XMeYxDJFIm/1+I7zsVPHo
MpmyZ1+cqjpEEw5IjXaFq2YEwbxO3i+jw3ai5JLC4S3cjRk8F8wMSYWnc315s2H9
pxXjbIByCk7BYikDaESz06UD8THFjrB4mm5hjsz/97K1er1uG4EP8acVfvxYuW8N
GTc9Z7/puetcUzFKIbHy1Km8qE8gsp2Okvu+kqgLcrKDtMesXUgUm5zjmVRThSS5
J6BtEDzdgIop3O/RaEYWku/AoX7N35HDu9JvW+NXuAzMWsWlu8liJ/851N2ZZN7d
rCzWeO7gOJJsFnk59WFEaBwVle5DrLvvCfDzgx1u2Qu4kFf/0G3UK7JmDrHVhxTB
aRslvNXi281H893kl3hW0nSgc0eqaK1PIC8WoLpTr8HAaBg3Lhq+qD6CCnXb+L+R
HAg9agslVeZDyQAamg9hwwxt4jG7atROsoXiv13rtKXmiig5lP1Gq9vaeUCEPezg
UHltKOUBdH35GbgkBNOyzXqBhkzwlRCemJtSvuS5lWmSJ229Wz6pvQQ2QUHEF7p/
Lhte9MCsm1tZCkPt/KdJvHUrUzZXnW1H4sGSev5Tna65Qo2X3CZMi1p+mrSlLUJP
5A7zoTmPEDrRIM4y5whvkuRG1uoaMMj42W01LZAva192yft7uPRK2sKqGOeNFS98
IlJqrVcEUhjHyaFxzowbj1cmdni2xeA5M3BhtsNB/yOoYXb6QW2G4lEFfiU91rb9
iHfF8tG88x2Dhp55GvufOFFYG4SCgAetA+D8k0Hb4dXx2DfiSq6Myz6S3MbOIdrw
HaooKxslmlC5fY0lD61A/7w+1wI5UzaktZWTcG8UgKfmdlOOuTe9QS0cyXtUq5SG
tW4n6Q+O4UBM1buR8mBULw/zDF9JlKv4MbbW0PDnpfMLjtbpOx8ryv/ktFJhVJde
w55bJsecDKJlsumvqNZiGT/xkEWlYkyV16vaPme1mFOI8kGO7YVFBS+SO70qaTnT
JIgHIky3Ey1JAPo1P50f57hSdx1kxQCn+/SFBfYoJGQUXyz+UjGIddsg1zm9p52M
Qw7OjCVbWSSA5lCXRuI9inTWmoO3WpPRH6yRxPHrNKR9Yc4D8K92RP6g2ockR4lA
k4DqWvIzPzOVwxY/jLDBtScxK4b4JZS6kr37/3aWCeCpeySCIp5q95n0yn3yUEEK
iI0lKl2e7G5E64GvYG3t7D6ITBW57y5O7PBUWXD2yWz0In+kJA652Gu1+twxTJZl
ptcc9fP8JYDKhnlPNxCoTOaelgkR1KyZf0YTCGnHkL7CAtjxiF8rCvw7Ofgfn+YJ
mZFCTrzmaEG12YNRjLOgoQA78o1M50Qp/G5gbXS3YSr3yT80um8MzWqkFFcVPE3D
MBlN0zmBDIUkkd4dU3g05MCwBvAmcpdmZ/wVL9N+Lp/53TKAJBsbGg9yfl6Z2or7
2Rsa1OwL/zWZyZNPadbLjUAijrfAZDlw1Lg3w8AhcENA7nMbz0HpBXJLeoBWIkYu
TiB0vqfNC0FKLCck2JoXrFfrrWCfJLlNZrzNJAu9vuDHwNPtiTt7tZE7hsDGG1t8
wHW8XvIzSmXp5YwYSFm7oMactrIBCzrh2UqzkTZJGmlw9wj9ttTT7iM7dWmj57Q6
aLbTprLX6BeiGenikeu6cDzl6rZsWSbR7cwgbLK9qgoWBIYeIZVhPlkei5EYARdv
wxt74MAXtdCuUddwR5NVn3BXYA6T7X4S+U1AeWPoWdeiYsMp0Oy1DOwBVKl2TZjs
c2VBCFZ7xyFzfKvdGkM840f5qYnDpX6X0HUyuPbXoSRphvUwlGJL1J3n3MnEPhbc
zTZRbutKmKIWdrHn3Zl226Je7pW1ongrbk2JiaSs7US6cRwIIGeu2szdM5zJEhRx
sdPg/eLRcx78Lzcck3n9LLECSKyBbcenZbptl7xYTBIXfWyj3XzeqGaTwmH+voKs
vja073sRM0xEkvzQ83RajKqeIV2mHL0Pm4slBW33onMNLRLoYTCAvxYMczKn+Xo4
e6UJ/RGuhBzqPuAFis28HjdkSR6wF91HhsldVjFyi67I0KnAnSvBZVGoUd97Y7ZV
QL9s5dlcsxmSBiehjbGWYygI3Wl66W2lMSRk3xklzNbwOT0eqt0Z7qtOYRL3+t61
9fjVJ/bEti7j2uRBQs9DylXYIJQMN8AoAlgBserqlMQA/RatMI/5h3FoRy5qORoS
xJlSSH27UvmMMEDtq6jOGv5AK6l/xCYO34eNDxflS5gMBxmncAq6ecJ1qdKZjXBA
Hdt+usEQIZuKvIG6Imq458cnv4t852EJlIVgUdgDhE5IrHcN69rk78CbF2iX6Gar
XD3NNFD9RasD5KnosH+5FipbPPSwD+JPFoZKhCtU+yhZKAfzuVjrq1tZR1y2XFgx
EjWsIeD1ZOflNLN3d+vOlXfShLhWOKNUbFbxS1zMDS90nsOvmZo11R8fmR2h2IC5
B2hW8dWndQY44A3TjYDl3pKb0P+18euO5AC0K3MabmaZ+O66sNKNWg3VEdP1K32C
9qFc3pXjEwjn5+p0PcAjDbr8goetBmedi8Rq7ZccDXyotfL4HwfKyedY+u7OYrze
ncv1jkr6445sn74QyqsHbVfGkLHcpSmb2UlDT0wg3yma3dszNCZ7ktvvTC25DWbl
3BFyauy5wc3RJW9vhT+qR2mwxs0d/rw0FeRu/CpNTx4b9jXNdHPW5A5XyhY27suv
OC+2Lu/vpoEglFbAN369O5J9261ZRlP38SbXAOCx59GRAaC9O65LaQ085zEb2Mlj
HikDdixKBVtU8slP6StL15joqgdWpUhj5MXqSj/ju6zXNwwpRJ7EQKM2JXSnHAHJ
+T/3m8qLmovsdLoieIq3iRAjd+EIdkv/BN0Ahp1Y3CjCBZ1kSZitx+dzQZTyclEa
5tBB9TnfQPES8Mo1r4NT3usjIMP6SjG4/czU9zL7RXXmJAP1jIjUFifkeC+Sc3KN
t8q8GyW8vD38wbtm+/ZDuGDpr/hfOZJwUIpYf2BX7M3yhYdrquKeQo1VqrwOxbsV
5eM6e8gis5BUU3M309uuMi2GNY4UB/tTZ+G/8D7FKEkrybYnY+4LAtvqtvS1ZO2o
IciL3cPLEyqGe9wfrVEPTUgeXYC/LyZQ6c8kERGu2JHlv1G+wi0RiLQFAyig4hQr
P7dfhoprrPskbS91ovJ+Dc1W6bZP6I148mnFSwEl4yvNTSRjIIVG2hAzSoIaiDFi
EON5R6BhTa7VRlNaBiMT+yVI0Y6qMCELGBSM32JnGvArQnYEUGaP0fmVfG/usxe1
7IWcPgV7s30AXUnWx5oovPcktv8dY5GIh/RB5+fdDgP5upUqc5qOfVZci35pyATK
KqaX2nIzpKk/OF39v4QqQOQ8KjCTC4GbYdTLm6lwdqyUhDEXYCNDHey9oarnulT7
vHQeyK5+giVtcAT0dR0KiTBAwsHm9keX3APMastKTSb+gOpvl+AGn/JLplARimVU
+tDrV9312ilMD96K/bf5Z5h9ZIgDQxzn32PFtKiAQPRDbATp5PtqTMYXWgzGVu+o
6Or7v5NOwfIV5OT2lg8DJCvdRmqQDtFtYt4vYNIeXr3xoyEI3tmacq1lz0wdZYMx
tgWpeBYg11ZMr1fdmR/m4RF3njbxM7nLKa2K1lGkD4W+FZFGw1ynlfS/A56A8zOi
11GWcLwLesyJ0XeoLkxGAhdL93DWlFGuBeS7G2Hv59KVnQyZKjmO8vAniip54W0K
xMj9i2X2s+Hh0EzzLYbQ3SojBd4fv6zcWucnxeTfvbLs9bMEU/oaypnEMa3Yddpi
2NaaepF1Y0w0uOiDRaczHrKka1+ICgovOk6SBkBw3ehO6SCfR2PQTcQ51m+rz3n5
fnvribHH536jlJKwemu6xl7hxIyy51WQJuExd+2AfPpCyLYHKHyAZ3HWmFfX6PYO
TBwCT7ZBEoghiNGbR13F5SYHpW5S1cIT9iZl03oVVpTOxSmUCymdx0gResAFdVB3
5rpQ9KD90R0zrKK4y+uaNWBzdVZJqjY2zP3d6sild2viPkg5OVV5C3+iHbz3Ka1A
fc9USfmwNlHqWEY5zplRO/rwPoMrKolcAW/SLDXYOlZrvdUorlSBJpjIFbV6Pjxd
FWGb1M53U/Z702Y7+Sy//4BXTSfdAqntTaNhWthRoPjADktcbNMRo7rWM6cZX/ue
RGng33motQ2vA9nwL/y1+POFDqp3UKdJPL19e2bdtFbDma04zkoyWULp0B+ykHSx
PZ3LbiCmoKoYQXaF+FJg48mWqVFFkugQArq3CXbZ6ICg6rI2YRcxg7Y59mLOWqot
pjl9Wcbo5AsOFcYPvWAjGte0rpv3N80mxf/G4jdetUDXU/9ZHNXM5xskz64lRK4t
7d9xfjUbkc5J9IiFGGTgdaYd3ZK7q9TuFZvzByhxuyXpeKPe95mEHTKFoECk2iRM
QEuTCtD5wiWgtM4xSS+6TFk6TUsQLUQLCIvfAPKq+dil/QZ3fA55i4swc+AFj/tN
v2zVb0efM/B9aIIBBExKM1N1AgeEBvfCC8iD1sowcWPqcEHhy3lvXvBVdGBtXhro
u/16EFnYQ32EpemZeTdqLjCeU9AFdey/4BAlIT1momBqlh/mWmECaadpg+/olg3U
iJBn6gOtgUIFHvjQDTmlgJUm41iok7Aw9Z6LgvlwGb+yKIUjEgShzQfyFqC1PE9z
AqPQea1NQU1zHemDQAmIjnVaNxVB7lXaKHEOtmfzMLlnK+Pso0fhRxqxsL6fUS5G
SQb0+hgAAlmdJnJtfMMWqQ7j+XChNHxPFuDvjVGmy7PE4Nbhblj726SG4hhfXCcj
TMZRiuG584teEyi7OSVpIT35zE7U8WAxDEIDA4KFvDzfMMSnL3Dsw10M1q3MVS7c
u58sPSAdDyXQXDVi5mXDWG+L0m+vOr06KcA7Fc3ucXKKcclPsedcRFeVt1hLrmeg
8zTaylRLYRcr8eg65Wzwp19UDLW5GVfglqo1VcJL7qB4EKS14bY6v8a948ltpc/+
Tmji+dEtca2dTtDQ4B5qSufO80Y9e878IEZaRxsQhvMl4v0THRST2i379kVnYS7I
QFBXMrfJeIt9JA3IynFSO890lieGFXZL54xYgjPJhWmYM6IWefuabBjr/kWEF3yD
bgCdNkekn66jF78gAAKYAyNcxhSuGg90B9tp256UiOCzxfXAPixl4p7KZ9aoYoae
sa+qpwNa0ot6MhJ6AxDVp7Q6vxN8IsIiV3TWsbc364TBHZ7AxRM94w8pMbIspAEE
Bi2P7BTjeG9DnfxU6LHLsqhW3ipoO3L/2ny3uMEfVfooxSsdFPFh59AElW4g2Z7g
ZfDbV2eIzIa7ESCnExnOCioywj3Dhl9L5ppXZVhBMkgLmZiGEFn95h72JUTe3/EW
4aSUMTQsDV/aSPzV39GgbTVAmCH54Vg2vcLKuuTcpdkkiUbuTIlLuipzH3FLITQX
woL+LOOlgqFnp9lhdeseEgJi+qNIHHuieRIYg4n7wkgGRYngwb7zdsRXZfDwOykA
OkQhu+jhOzOroCd2SZs7kuQpgZZb3nreVt+/fufcvqCpKdLkGa1TTqBIOVYa2oId
214WxzneApwAWn/FgFqviHmgCWcM9g7Cn9h4YENR43h5s36wdnXKPB0wZDC4a7xc
2UiSAjwdBL8W2XkctySHIWW/fLpvebNCn2TkcMbEwdjaQKbKc8Cep+3/dVzqBh1l
wEWpPah/h4afZMnFM9LT36pBbMmb+LTKXlEnNcAyBlAP6W5x92hGBT3xUFqwNXSe
9+WmxBKUAUoU6T5tqLVw24qa2ot27nb7nZQRmPA/hhMYrO7jtR42Dr/KDu6GfoKb
COjyVRcu1uyZKL9skPksPPqmPsItwiNlVPC4imq9pK35TlNW74gdHI2NkkU5Bmbr
4Hl+G3hnHlYFNM5bAL9IO/TGkSBC9IKnulexhhjpotOJAY8TAHc6LP8yCXynsg+R
Ss1Tn53KbEsaemeHTmeG2J6drQXk/CRwOjWCY1QDoZn88e1+AY9zASBSMiFCulX4
Fj8Rg+pvLcG39RB6rwZLyZw6rgfJToER1XKoUMOnq+ZtHTP7oXE3Cye+JynCpa88
RZhBS37S7LDcaXPCTyjAc61DA4t5l8e9uLYg/7GJuge/FpX04GLMiD5WVy03AbhH
TefbWCP1/Uk6SYzKDW9D5CDa4TpRW29r124m1+EOFw9z5HVwyOIQ7i9l6+2//Xg/
+5W0Co4S1SJXm71uKv2qtZXhbKqD2Y/oJfIaUZv7fxWdoXS5m8KMncqx3wsD3nSg
4/w3xj+ojKlcErePlu2DweIyZ9h11OyV8vc3Zq9TOz7/NESYJ/3h8AEdxV/aY5kf
X0nXmwDLAniEd9SjqUGdznp90toLA8MBaIsp/iy/76/jqCMErMjvuDXkTlr6DhVu
CFbDTD1eJzDi3kANY6bqdxLH4FSsluM27FVlf/C6eTo3ilCgF4ELuJtG5GPbdTzR
7MQfuCZ+TNcJpDOa3ASdv3YxsRsh5B8T0OXhiDHM63Z64SHCZC5aGoRivt7MDAUi
1OtJIIAYOiF2jAeX6rD8BGy4rXzS3KarCxQJr8QpEX2RV9h0CcCkobmpEtriUYWM
APa7JIYy29iUl34T2WMu+95ssV/BVnglABj8tp+S3QeHIobOqWp3kGCDG9lXDAnA
k1EyQRR1HIZPpmIKkEceEGvRPbJSToZZ2rxawSt2u3lHhGhFKk2kol4HnqcEJOzj
EPb58BOJXeMZ3NdoT74idQAVAVjiVj2+knJleg/Wu74YcgHaxJW6CvxS1/0eN6XG
pmbZNvn42NxKMwzrEHh+ZHcYe33/6GxN6eccm+0mc4ZwryoFSeyavY8HoFlrFK+a
ilv/4yMnnsqeRRy+rWqKDAfdiQdijIC/kgOGZG+LUMFZenyCmCgATmihBbh19ZV6
j+lz7pCYph6zYqVW5kkp0NL5NDnURjh32gh09ukHb286ZWWefWM/67tEi8uvgGfG
Hgf/EO0BOKi0IQXPdIQPAdlPcLZLpcQ49i9ePKRr01lbE+j3wyebyhO3NOL9KDP5
3VchK2I4eVykOrp12wLvscgvFCsGkHKOkO4087kr4IRnYd283V58NVZVvS6P9NdB
MlYC7kKuVDC4zyBgWfFql+RsOZqUp8QPwkG3baOG8YAnIUpOdrZEJKYCFXJVrsSA
Z8IW3B9hbbEYkvURdUKVmfIvU0IVVKllTTivnzOEFLQvg4IFGJX3ZQrPO3mInYZw
nP3Hbup2Ca00rgVj4FCLZtr1YNxrbUog4AtwtMinJS6WWbrVWNbNhb61shdZRoys
YU7Lu20QcTvUN1GmxZG/whpBTwUXBDXozL4VwgW5ZItTBBq8pQCXpHxTmEfYG/e5
g9ZbqQXtgaZttNRvYH5OHbTloNXDAYM+XVyGEprOngcxosJccUk7eO+ArVw4tBDV
+ge2Ktk/DzD82rJiXsqD+s2OP6qJPX2mpf4JwwUOusr4Q93U55HanU4QtMUrF2GJ
a8XWXPgjRYv/OVd/kLeME6Bx38LqKa/DQbpLhSbjZAv69UsBt1FlfwUgKz26zPRO
B+1213FDadU2YsrfF96WmtcRWozfFxgDbS0g1h+e3/ijpqe4eC1kBN5/VWUNKTau
5VEfdE30zL4Nqm7YaK2ts4Ghto3P40TKm7Y6ZbuKgsCfEAVshxFlEhGwy56y+O7o
yJD37qpxMXIb5yl36/De1u1Uz3SlsdOrJ7sL35iQAbunuU7Xlqht3ipx46thPscy
mkhJ6ON91viMSmtCEyZBvpaa+w3f1OnHfF81aa0V/lXF0MgggkY61pCQelIFvgtH
IiBFuuvAsZCB8muBAa6yCE9WQtQcto0yF39tZDQWKREcYyxQaHmspPRw1vg06kTz
qdQpOyY6rhHwWNuqTt3JNI10rHc3TTe9krIfawUAMhMiItA9GOIfJhrb2cY606z7
lLOqYVM6y/qwp2I6uHHlE6R20/icj0DRq8jaI13BfiNgh26O5LMU7dKPViHryayS
PFE4Pe5cqrVOe8LNdxkXSmnIhLBCicm6WuljZL3gOQ2U8g+RMnJVNwWpvz3U334V
gU6mpP4ez7p9p+sfRU0zOJptJhSMSibDZzkXgS+V3n7S5Q/sCviCQ0CxOMbqCK6i
2JmDVs2L+uCEm6gpdcUR9wEY/Ovp+KuOpO+vqROxrjXcLju//qQJqutjafBdWdIJ
FjZoSrH/6B8TRqoDYO6VkrDwUIE16ulKuGl2dm6Qj66tg6QwdnQ+KMZPa+HMgh98
zyCvMdmns2eW1q72OUhtuPId7RmW4niyPMvY67VtDGTBVji8V6qjPb5NftFWpX1U
4k2uI305oda2batWBGaM638gxQ7rruhveFvIv0Wm56C54fMHgSLkpb3nh6tDMbhm
ze4fNy/BgUvYrL/8XsOOBItOXPs+LukZKdhlApdZkc27o1hMC1MRRc7s01i+EcNJ
nwDhMq12XIBYA9SbL4P9li0M1grGtMgmBW0RxyZE6n756Ldpwcw2k2QWtbQxX/xO
THRu/QiEliHsSrO0wh2EdYcNwVTZdB6Ei7yLKTZ7zbuCnH2E8r+HsNZwtGLSWyPw
3FL0M1Xpn7IV39hJH++7syLiimozDzWvFfAOZpFxUXxicVLuxXZK/AjYBsWmyac/
Z0I6LrRWv6rGAd/QMSFD1787PVa9fBxe8Hd3Y+hOjyWW+vPn02EWW9DoqlguV08P
pr5P5ZXPOiGjSsD9gjRq4dhZghaKxAb4nFY+L90dU039Pr7kOpwD159xCn3C3c1d
bgxKYRsR87Ccco2L9gBGFyW1z4b6yAhxXgE6d7Oc7uz3EgX+eaV7dyN4CQ+fWcq8
/BmzDAgpZ4zsbFDwJhgPqN6j25HkcG4/5kITDxGwNrK5Ro/ua8vW198P7InrKNkz
xHLYXfAYmrXMl/K3dnRzDQQAuhFE3sWmDa8zd7imkWI7kjGJhr6l/KrOPaYPxGQ3
oNY8k3ue29hHfOavdeD4PVIDrVCxDVQOyujHPfh8yTLx3vYuv2mlNWUy2BuP32WY
pbIc6ckv3iOuvy2YcXn+QPLwks5/tIZhAGct8EdhKDBNe+mgVw6zTXtSInt9yQ4v
VV/GsmLkKN+ghUqoemP+x7atdsp84c6bQ7514LT4rFeI8BOtOStdq2vJWoN9EKl0
cteftzSR0rrnu90PUgqrMoqm32UPQK6I4ggefArifFNVnLIxbSkxqSG2xVSa3Cth
XsjQ5EB2aqASbUuKkXGegyOkDN+jlj4g/9ugVxzec2Je2uscKZ/XW+K0W4RlCKUR
MZXUNvGdZUSBiXh0r/wHh/g3hi2EMN9q4WfG0X4jRDCvINqbUjkjrRj8d1pJvOza
J1qZ6q81A+AwSUlE6UiB9O2aQEQAzya8zwaOHi83IXXginuWLtFAjyZgrYAo0MQh
jMcnJglBTkEGqrVRHUcG2o2EWEuI/cf0pVNixFDHQrVJthB2dgziA2oNGD+b1KVz
j7vx0ve1vs2x2XqFf8i1Ldn13RYnkTWnnBwrScYD6xlAN5XgdVjJ3j1JkHLuvrfT
tMbqDWS8ZU+b/1rh4WUnzlCJ83W4kmDgDJuL/WvToOMEnzAmfBfIdkY+q5yID5as
E3XTbKjh8hcRT37jBHqx62OmwrOwI8P1oVcmE3CzzGNQshkckS8j2WoCY0Aq5Fgo
B6aJsgX3BnfJTfZtZI6DW7+tgJWVnidikcx7+TIfT1lFKEXkM23umi5ZQ+L2UZDb
szpBdsB9nnbSOjZS9/5+H9twevSysLEq7MBKy7hKtBoJvBG5rLSCjLNp+ffw1g9j
fvjllPa8TrpgW9qngtskwLXSEJMg7K4is5nem6CI2qr1HbUtVjxW6z5o0TxijQ/I
ARzq6cujqRYqTAQeIf6IFBq27yhblaj0UoIljhdhS0tbRENp/KkSI8GxWh2VJ0Xz
gFQOSmRpjMdfoO16lcitlD3R5XmaEf/RKpNdEtqc4WIcyRh3AothBSKQD8lELIug
11tmcSHChAb6VMTTHc65UrEL7nLTOaRNll/dTpyD+wfoTnl4PeNy/pTY1Dp61LXb
U2TXqCy/pviup5OGkdRgA/5/tDHBRWBgzuIK0XXYkzWiqWPYtKOl2LJpOU14LlSA
YraNzuURNFamEC2R1dMjU6rZU+zMdIQMc4aR5rdW9I/Fb2Hw+2g9UAXbGJqZudZX
XaJslEpm77dDDsKwuqfLITUvF+8kxP0OfukXIt74yvVyDcdORfAHRmQAf+vKvQnq
kw/ii6RmreIGxrKTrF6Rakq6F50xGHNPMiEYti3GWWAV9zsTIBuTWX5fmjfDdpzu
fI/kvSf2F2kZNDx6X+N0yZPDteh953uhgJ9kTP8gbeI+COcOL4NwpQlXqig+tl4k
S/+5ZgI0TUdgrhzpI7HCBmpJ3CGfWmlI12GGBkXIFq9lH2VZuvUJ0bbxZnh4RToy
hc1AQeE79D8/i4rWrHIC2Ob/5U/wTyjKhwsUDIKnVTN2tEsVFpFCFZeWCevYfIV+
GrUu0L9Awb/FuVkSGQAr/vBjv2pUNQmQCxaBVdVyyThutYQfFqZ3WzOAAYbkUaGT
/2DQFQjJAcx4aZqsqEjknUYNUG1foSGUuU/xRsr6m0IWGjNy33nAI8HSEX31x61C
zzg5B6F1JUhLbywZTBQXnCvoNjZVRo/Ai2zOQiWuB9lddA9gWYGqsIw0wCSBiose
bK2VDPtqDYft3NslkqnTWQ/noGE0YKOr0U4a1KpQsWyWev4O8JhWGoU9PNSNhubF
y2jHn5thdFwzu6sb0NULHF3kekXcy0D1zeX1PEdShtV/NAWzI/4mvF66A8pgm2mq
qO0qFXjtmiNFlLZNyVvgwD4Pg+dx8+/dqlLX9xshPTD3UZrkvJN3IQ37hvwKHZx4
GsICQ/A9Zts3eYPi0/saa7DNqAiFu1S5/fdv7OIea+RH5p4fnhcaJwzwNVb7TfTo
6KrhonD87hGLRdVhDxhmXy+nntJw31Dd+GdCw38YbF9vHWCAlkaj6QI93DLtFLRl
U9fkazUFzt7GfPTvjLzwN57/c55eEuiBhEzdS0VRFw6KTfIMi5UfrPNNkhpUB5fg
aihKNkgf8cU+QSlvcIWm3rlkbFuK4l9GkdKkMJ9OdpOyZsR6aP0VpZ6aWOqlydiA
zqMlHN+u6HRyr7gLWVTXp4M/6G8UKsg0RASURFFanh+xZNu7Q9JDrdApuowXXbv5
jH8XCjHokA9qaU8VLenjMOSAS0tDo7C8NJo0KvfuMNeGcrLBLcK+PbSFnDHrfH6Y
WrboHqgYNPO2rGST7MY29tdB24VqLw9PPLJ+ay3xwpqDE6Llk79I2RECQqAd/Tqf
OrtvXuNkLmMwOMvx9iB9Mg5bVRUtBuwrUzOB969Yn2hrUCwUtjNnz05Abq3RJ8rS
6noBYj653OGkKu4s6EN129UICC3HY8BtjrsBLUFj5V2zqamy10knla0W4PMRgLQS
AgVSWr/70EJCi4fCxGJUdLgmLjwA7454mkroyo9S6BXYCdK7iNN6Iu7WGq/Bpnbe
r8B6g+Xoywvz328OXaE5buSS3DFfh8xWn8oZ5SO+IX12ZqYwcuAOqB5Fu+8iJKg/
m6o5JsKjr7t4kf/2MsjHYUrz2Q9UaZXxCMdBLDUnwE4j0cbI/AKOX2MExMYgjuyg
OqQjgus/NgmlX8cfek3g4bmwL2wGEOi/dN7YGM+K0KkWDgyu+/VGO4zjUFxAPmCI
FpeA8/fkrfj1lu3IoTS0ridHV2bWLUmh53t8gBNAS6TGFMQdeKN9HxHcwhif5CiY
T6+CmksmkfE5LfoEd3SVnMDM5zKa8jzefkvQ1OJlDxyluUmVrC2HeumnkCvDJmG8
aa11iaX2k54/HJqYMbFxnTSPK9MxuwO/Gv6pXwTrbVjJgobdkkiPIWKx+LvD85ui
i98XSVVeThSf/oe791QfPprzBVAYKYV6r2P+BxRgCzlVqOryITSc5piiD2YqIRZE
zQB5sbp6Nju9jdejwTj0y54p517rDrs0GSAQLgzowf4Mabkwb/TS7oICBY6zw7eM
W45v4auBZFpfxp6fNsc2rPky6c5a09bKyOTfaFuDDTVDT4JNWAuqsftToMsSOGfG
QlMQYa6EMBIBOa6FHoB9VQ+uEmYqF5kipqufpYtMFroJOMbbZcYb/TJgCYlYwvPa
b+FQPNhsFVwear95PeGfbK7+BXCwFAxLpgJ255mIkFYVK+PeYxfnECqSZUGEqgiy
cOjH9hNKeT65Y/KS7TvhKBSWwFQk6uIu7DPA/gfZv7Qdf9Vc//xPQnIjFssB9C8a
YajNZ01BqAAaKP/Pq/zMeCQdPmPN00/olxTvzdyRxhJ6/39pj0xW/5Xwl8otuEbq
6CWWMOIQcWikmeQbBnIm6/TNNz8DJeC40EpYB8z5ldJ+2LP+bjq0sekIHloG1ytI
DaI/ArKgeYg/dA1qdw+BZw9N7KAhBgwiUmEMsGWj2kwyjA121EeQTs4Mz4JXNu+V
IbLZzXtOM8tPdjbcIyDP03MawRfOFoxiTFWLUog9G0J9Z3n9N2gG1j7Ov8QzTagW
7J2nirP9EkUUsPp1YxtJwm5S1h2VAltJny2XR9tbRqVIpl6ajPI7MAFmsxqcb6DH
X5YwvPtjTf7zRcyjvrqlNXdY4gPdD1QzB6ZpDUrPpIlVlSflW6p7lDolhBM/3pxT
hHwge7PTPdnwDLrouRnrVXRt5tuNYQXQsygaZwYqiJfW69mbMBIB0/On4J2AzyBt
ajEUFA7KYTuc4bwatQPXPDCcX6jXeyj1lVXkn7EN6TQG5MDPtzcmKlYkM8VG/Hdg
0DQH9HKuWHTHvSjxY+oM3/mIN4fWLLuThfLeLo6TYvg9cV091IqpwDRuvRlSY9+9
fAFdRdVvY0jY3SELCmNp2HL4ioOCc7KTXrMKMOH1XEpdbX7IPloNUPslTBx9u5xX
Qd5TZDMASqq4JRk/be0/qf9cYK9l5uWUdTDGCzl+ZCdEWM9K/vuGxAlHJolBuAMP
Jteb3YDCZD44aUBwGjJJhwfrAimJh5r2yvEc5TI8AcXI+ZIs2u+hW5IJ8d0Xu6Gi
HxPu+wNfoYFaRVX/NSeIvs3PrV7neZPyUSeXnEndDq+ASecmkwsHUTZpvhHpiW6g
EjecLN7fkjrkmdABOjReCe88jMfIg74Eo07lztYilayJszWthwcRlEPrmEw7n18u
r9jueRO/CglMVTYHUay2cCUb+ycB2fdb0tX0oWe0A61fx7CBvwibKuzz3GWtJEUA
uaeObUqzhuNyLrhseQIk2vlgQeYLR4t+LCRniwByfHoyPU6KnPxCmrsVM9XQNPiP
xsYvzyRzh1NZFUQA7w5y41soIQWv6hgJcQBgquY6wrOWvHHu68jaJoH8tHVIR7+i
XrLOAnhPc62xExzyrVH+FhQ4BF9dH+d+sb9jxWhJYqxRH0ov5t1vZabMmVd+cQx/
er9CGXeDeOSLa1Zgb/XZIeEtKv2ErdHxTfj8CFH9JdSrxZLqOSLHhGz/PHuEHFTR
ODNvIxW7HqrXhbC6tFp7x0QND2dvaMe5dkDCUfeKRKZivyDpGtqDoCM5ROO+8f3g
fgv5xenmiFdmTC26Pt1iDe5/YcKGH7LIMTmQWrXuzTYE2f1xq/4ZSF9uHdqwB2I2
s7npgixuEWAfS090Y/4HtXfuftA1NncbMhLwauZjCaCoAcI/TzYtUD1gBfucDXKP
DjsACqn7akN5tbRE8GeEmpO1s1QUWxVhDSM3pvj++7BKRg2LmexS+tM0Q81hQHqC
uyRxsnU9JGCLrygWQLaly5ESg0ACt7Vgxs7BSP/rx6+Cn/Damxylh1oNKzGSwsq8
z/wPa9XOapQVrGSbTt8y3y3VQvYb7SSgZ76o17BB6p+fV7m6PfaZOQVP7q7GcAwb
Q/dQ0eShD6DO52vXIWhIjzliX8QpWnJUPSd4O/7Fm/rW0zZulCQ6XpfcnruxVOqk
x9vXCQGErdmjwH+Zuj7e0eQdYuIMnPUNuJ0dwugqrWiWkudINJblAWrFWPLi4Kf0
lUU2aW4PcS6/zA23Sj81hVMax1zT+buoSR0JQzBD93ZuC4L17MrxNy8hsThQwCVW
`protect END_PROTECTED
