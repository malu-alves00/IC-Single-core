`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YALyaoOR/LkVQ3vS9CoEB1UpjbcVJHnhlfMEDkL8tg9ePH+kLB05zjGvm6Q53VEg
GD85sJOQLsNT84viL3GBT8Ra9Cz+63C3QQOtuM4UA9PQLogkMO6SeM+e7SUcc2YV
5fBjuF/SARqI/ujsllNrHNUWHGkeYgkMWwPHa1lr3+zV2w0WgkkRoFRim+xR8SEu
gf36xdje9Lh/muMQ6DJKC99JoWFWHlIJ+AHqX0Wfh1G/XRbQfPRb3b+jSxvK8tFU
svPz7HK+nWc8/i60EuhsPUbz8AY/BAJe1mf2ck0rS2L2THfpOlwB6avstSvQhPds
kKg+C5IUfTkck7TWrRM7zAdd0njvYztmmiaoGpkdaJzG65mE7f3C2PSbA9At+z79
3AMb4ku81dpGTrnKK2I0QEnR9bv2d0b/S2VGGH6aGpSQ5JdNWV9w2aNncsKdKF8f
/sSvPpyXOBx8OvrjU6sUirFP58vjJJr69JQVaPh+PDFOC8/caF1wVYo205mVtQLJ
4wa+0SGmDkENJh0rnd3G0Y1oUpS3/95X30JqNuNhxd8uXy59tDnZ/2cpJ21cSv4Y
aQ9qTak53/LB0kaF2n+ZtAiicua9XEi5xKXxRGJKvBRnacTn7hFiVW5/+JTFxFWr
mDUY/sQzDpZIjIedGk0GjfysvCCWAB1XMX6k2PPSYsJxYvdacq9dUrPqZoCAZc7f
4kTICnTDvOnPhMtnU2Ud9Ye/rXZejmolNkMr/OPLNI67kvixCxX9g3SC/ngdxcl8
/Nkyoy6GCra9R+drboM3k/Kt8rWIXHC3p2oE4nuVxsdTSm4zDgMFr12yohlNEd8r
mR1aqJsGBG7s6KzRQDZUrBGzhyTupIdK+KOHuF0XDWX3B+OSUsYYv3MvgFMBkOJO
kePqcZBcv0H5heFhflMWPE68Q2O7MZecuIQ1O8vY+axHYYh32G48wDVN60/IKA4S
S/vi6C/c5mqUhn4lL/BFAqneS6qpQGk2PjjSvCgIC+ulLH1z+sFX96e1TG6Z+nTO
lrftnIp4+8dbAp09YItTRvYu0ewDfaxsi9hqUkBecRJylH8FDVRauKBSDWdRILgD
SpAFI+ruZx5AhSZiKNjgu1sqJeMUnD6wvQzyTq1vEnvYuGLsxP3q6x+g2CC1PlKN
thVOZWyaMMsbwghF7VSZVn2kahgPysLTfL0EkzPeWSYaFef7oSBOCD1BZXlaIyv3
Qk0wcKi1n9flwqP4ETIEaiCJOGbyNHc6yPWOkPeMP5emAZOIjNc3HKLjWDOUbj0W
4lD+ahgFrLZqdTbTfXTPhiGjOhB1LMotZTGWzIa/QTiCIjRRwHK170gWw+Y9qmih
tVJWu/NrPt6E1ID3+rQGjRUBRws2wH/176rIrBWv/C6cQowLpeitPMQUg7/pkMgM
P3VHXye0KH69oZMAcmngYiKQrXUD43DyGvYuZkVWnh7wp2Rh/dchVEP0B/Oc057R
JQFfgAtw34ZfeseCTFjsTPg8NYnP34Ayg+tNOc77Jbh4zJD+3/JNY9gP/OjndPWI
gCkLlESTewlPYtxgL1AppyRMRE6fsS2qF4PJALu5w8hr17Q32373ySfkFqbX4D83
tO6ptRS1XLjUNLWnrLV9t64l/3Q9Du5AV6M2rB3Yn3XRuElqNUIaUhI6lCgubSsx
TpZ/k2FI9Vk6Q+UzYt1i0+wWyirvgYs0dBDkW2tYSGml1TKOnHMu1AO1MxJR4bfV
SyLm7NK9Bt9UhqQ/azquqU/cd0sH0DMRkx+n9jDiMz+Xdq7i3NkkcTipfKnuR/gi
ZSwjL6e8ohdYr/jjD84v5GLzq6uHVSxt0a1hhBWBWgO4+YeWnPql05Ru5F5kIrNH
rWr9Py9VJKdBxe5A3LpgrwRvYwafBVbyy0Uixwb5oYVe8KIeirqtE5n4EcXCmTZv
D/sZjIH/fxRYP3uFSpOn1rSX8dK+K3tF+jsLea1BQkWZLDs1ZAd/9kzC0sjLZyPw
H5Gjnz1p3NLENQvripIQUkYgXmTxXyQroLcTxhxgrDulSZp3aQiSKycxuJWakIdn
geu5RAeWO5cCv201y3EbUyBiKGSMvFHD2435M0YtrGX5dTdQ4Rcc1kNWXUvmjAIv
1MsIKRYumdEo2imN/HqeGAfXuoIExDsooPwT9TxPpjWizqN0v2ZgLFnqIehH0qiG
24ZdnjuDvnU+fH+Ip8AH62zOoBJ2VwsZ/c2DpMamlgf/7hRq1WxReFWIXlHdr0ee
Jwdw48NGGZ//8sT2iGA78QUFTWrHqlGZWZKNqbRz13v5uidgyp/f3JVRpltTqKNz
sDhywrTiNWeS1hVia4xlO6zNdNNTe/Zs7A9kIWdjD4iG+hY/kLUE9yTb9nhYCgBR
rgPV1eZlvufU5fvAy+Y2HA/bH3zo/k1hsHkKfbtOlEFQOq32KVGH+NGXAL4xruX7
zLKNlMbLJ+4iR0SamgxxD5bc8tpDvDpyj+ETL35ZrcqM1B+LeJsj3N0Lq60Sewmp
enzasfQingH4WV7eWQIFnBZJSIQWPkpIW581zrKa3fZ6hanCFPkSUcT4MNPIDQxY
zB5Z/Ua6FDDr+tu5ezGlnNlq/DoFRmuS3Y9XdQGa8gVHPChTCHAjF1O7oLIFkEDd
XatpppoWGfI6Kwcv9jkFKDUXSFnKfr/HbpikToI1rW1PJIt/Uuyocg5seiHsuQDB
H5YHdVsq/p9XOOydUBdqZPqCoEXT00Qwl95jfXBr28fvMwIPvxBNS1+YvuPF68Z/
DuD6/GL6zk1+DtkoloA+eVwjIr13Lur29i+xKFe0cDB0gYtqPa1RqXBDj5fatIP4
erUoR1faqrP4fAyNwmZMDYXwgNXde4Ql0SqNumIcucVwpsMZ6gC4wUxwN1SIOMLF
fYuxGijaRvdwRcf1YuTNTy4tHc80pl3qzuNxaW30OZEtx+kRtJs9ucpk9fmXjWs9
RC8uWt6hAYAs/WYbeace5Pq/N54YbZdoGtZJJk/N0sSM/5jf4GvLG4JC91pMxuMV
OX0weKmgXRdi+SBGaNxowb06TE8UwNXCagHweK9hMt7ycYy2Qu/ox8rYDIuY1f6n
3dYOxGcfq2rGbDIn09qg7Qh/a4bDqEMi9fTtUvzXHxy7/cxxtTs7Cj1Xiesihj5z
/PlHf3r75s2LThrQ2lLPuxN6uttmGT4KItzOOwTPjjWE0hmZHsGU6eglhwlYxsta
+6isxIQ0B+1IPdQ9szY92Bb7qXSIVMmR9U5TuGS1AdaLV+heNmgzfvDrRsyZgjNS
3wX4+2vJSJWhM6nLQ3xCVlpBf8BEluNBQL/GIjQ6Nt0ERFhVN6/X5lIbVA5SCAU6
zXxdKh3eVufciVgVQbbQtby+aa24OX1Sf576OgdyrOyyZigU6RrLZyeKbw1pOqwA
CmejZD2v337hNuJyp9amAVVCG7iOMBZMUx6ARGkBWkGtJSzh4Sf/XWw12olFcQ/k
+9/ym/a/6OOeaGKv2cjmBtB3yYwgxhLDC8qp48Zx/UHJWvD+IbRCvTpfCBKMRQT9
7vV9u9eHBzylps6tUanBFWvdpNFyYCymxJrihdWs/0qsj5sogUVh/5NyvC5zOazl
haIO+maVAmVyGcu2ybXhknh1HWj9O+Du+GvFTQCJ6mY=
`protect END_PROTECTED
