`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
17dYNuVXMnaeVcvjkpbDByKVZ5miV93OIWM+pq+F86nLymd69nbqct/gPaSybRo8
lPuzvy1++jcLITafleA/bJePIapovxKJTJaXVisqcRZX7CBm9KqpsCkylNByzsCO
6MU+bj2fiXL2ilZ//azK7H6rJScBXOmN3hSNXbElEitDpaOzcG2aBJDM7rBUgsW6
oOewyUCOsp35i8n6OU/4bpeh3rc/pg8/mrs5mIkfbFmWWzDSjpfcw/fKnAr5uwnZ
uAnGxswadlyOQng4ka/z/INcuQ3BtAcXnblvPCxY0pN/W/Gty7eIu+ElYx7tOY0S
BFLe8HllTxMvitVhXMBerrw9/i22XLvJ4lwPyWxXQbIgaLyp460VtQ3wnh+ryhmO
DL9eL9spHDGlGkObl5X6bHz7MP5/5nqT0I0U1Eo5VRS/gOazqmUDByEvH/jpaFBm
P1f+Wxd1ZJ8PaCV9I7g8PwjwbStnoTCsaQprVKXT5tSI4OXsT1m9juB8vAosTP6L
R4jRSP6PR0otBRXbHngHqAE/1f2oe1eKvnpfYe8vXfbDGoBI3TFVzKqMToiixoqH
BTNVbxpo04op/gqay/Kz1/9RQb3IfJWVrTvEaUFi+AEFiEWXk+AdXHz4PqMFKp69
s2eCD0yEkW1rMVKSefVhxvBSHvLs12uQhOEAuAqLGX4Yuq311WTdHkT2mo9wO2qe
wPWS4GWbenYH3AE/j1wNN4J0FXTci8uSRs2EBJsBKoKbNCEdbALDl/pqIWeoRdRk
CRQEMl98Q0/Idk9RTjAKbMb1MheV5E8Kv4oScQJphiiuP2soqwd+KsBEXuJ1u+jn
Vj03T08mFq13aHCcWY0WvMvAa4HN6P8IvlPoe9opU4W3XqCqXAYYIeaQaqRJbvz0
rFGbq6gAzwiynz0uYfk272XLigklzrNJpia5UA6xn0FiCNxTYctV4/NYcM7v9M8a
3e0hBtDR1SKOo+YRXegh1go+Tm0Bt1RsWhQlM/hx9TrFe2+OIdnX0iQ68N6ON+m3
nI/u4QqobYpDBP4rsKouzsjPv6j4EMAQWQJlzpza2kmTgH+tVmOENoosqPqMWnd6
K7oRPV90Rv3mMTxlBH3uUV/r/HI1LBPRzUKRdX3g0sa8gezBcl5fXOjF9pHBDfXu
IuTg1v6QT1tNCCybn8udgNayv3QrSLcvjoMzdCPjq98PaaTpCrG3srRXxvptdORS
wluO46Ho71ROvJ2wncrG+WxVLpPv282DZhycvZDfRLPiD6mTWhZwL0HIucj8nzhS
PRTYdiVEuP1+ol79sfBC/hWfOpa0GXbBrMWo2FCE1BAB7pEOH4Qkab+R5lp/A2ws
eo+ekZEOQQ6rd2FSZM4SyQlPnVIfjkVe/3ol0Zs2LG6MvARna6FTL1wtxYjIaWcn
7wHefm95sesjMSSvNiuxMtHtjBZQEQbHDONHwcf3jr+82kZeSlRPMZAoLUxZ2f6q
zgfUUrxkhFZpfngEtTa/p3jOhbCkJte4Sok4CwZqftsNeIv2Lyzi+uObG5flMxnu
VqWglOb9PxBJzRjuGWfeIYy2B8Yearya1PUikUPHBLArXZghlvp51dBgYc1++AKw
XYH0HLutRRVtWyIkaRh+RnLR9eptclI6+19l6lbBaZDIco0gFzxvznC2iUtO+Lk2
FZN+or06DTCKm9rv8NMTjXztoPN3fNmOojNO+b1QJv3zfJcJNdT13bLP5Is4q1Q+
/rY6D+caNXXKX53ALEdgIcqnfO1OmzbEhMeGC/55yrU2K8CMZcTZr+d7mwuLwYok
fI8+7sQqB4+mHqvQQcSbYsUO2t/ewzlT9DWoKihR/ZMs8j+g73ULJgA4Jyk8LIqa
46MkiRqxfp4pgmy9dJmSDX1jpK3nW6mrn4qf7E/Tc0qkQSl85COI+Uakw/WlEuXr
fFDqqKa0OzKTjSwUENJOpDGS9rsolMqZrP8ZrILfsiaigqdOm6pacOIsSFkP+5Cu
lUYZLG674BLZ2d6TBLgzkzK2Jl+LZlwBfTo7MKmOpNROCv4+AKS9YlcxU3kjNhg9
SUuctG93eieA9KAzWdcCYhA5JHlWlMaLb14KvmHd8jsJbZyPosFlk6gbFYEhAMj1
jO9t4bqMd7+0YIWi9G9pUvhvYS//+Plrcg5BjRpEaoXrYefBsmKMmhHyyvXRhBCQ
BFA5+holeMm/NZ1owBbvnuEsnuM8R0Esg09mkw7PiKTp0S6VQK30Cjyaxt8tQiBD
LFgkvPgf0Av2e10VD5Gp9Eb0RUhg3UlmSB+NHDu1eAuHJnLWQzjLrNNGdjF/vuHu
wAGqWnmyo7YJ4kYciNnrxJvR93uzRV7GLBccWhwDywsCBxzU2GIYSxPT/ggKwmZi
KFt1KkGSxXLziscnfyG3Q0i9/t9i47Msf4hoH20wejxVaqst8gU8rtsoEyYnaosi
NssuF14527oJ1RhhJHOgguMonF7uvJ3OtiGpzChzzoXxM7/V7PeaZrg7VEo0VYf/
3jJLkMaG/n9E+QhFVHclkBi3YxgsXLR5OvDMfGk+GYNgFK4S+dxyG3e9Zd8HU4SV
p7CsCL4+zoTpQwOEEHPOznk8glfQeBTe0Ye8ycZewLVKrxgMNYa4D41X8kz+5JsL
P19M14eoOf3Yfbt+heKHp0A/fO796GbHYUfOJRRASVErMW+8i7YCdaI+GyJVQsJH
dod2OeDbDpZRT+hjjZ9GzJgt7/nrcVeUIpB4ON6fLJmgzsi7mNBAqAb8d1c9F6Mf
/LzN+SbH2VfPFfyjUYTdvgNmVI+51lTVRpQsAKCdZETYovZ6dTC2ZfN8gfvp8Nz9
hmMbSe7I2yPdoxT3vf/89wEgQK/YDoY9850XyWRba9KmMHsAaWQhf3ptpkOTCmMz
IUtgQIbI1CLXwv3avA6UKz5+5KmPm2vre0edsxJsngwsscSw7JiUJRXa224qNMXC
RcsxBp+tJTeGntbEoK2cG7kbrXVKj9hO086iIL9JsamMFS/sM1Jep2x6svhhlLTd
bnqppATmoakHPRVYN5pAz5lLAOarTYdnP0j7JeaCZywOztHy+bpDjGt8IsqU8O6D
jImUEOcBALu7BFicUQ7Kqzgq38SmnZy4+eUgSNia7gNdXP/Lk9lla7XsG3Z0yG9f
Y98vvSsVU0kD6Y3PHoySIYlB40vmQvo7iVQtOFKBzG97kYen3301MzUapfEothXD
gJ5nIjHFj6wx/KvEiGukQUFH9nv0tY4mDqhGyrcoYUEH3FAzunGnIeWp3lI/N2gi
s7A9Y93KlolUvWbRdzY5YRQ5PQTp25utjLYryUhxIJ38NOTzEaVUPKqoQau3nK+O
7uBDRS+RLmEuJDx6M68harodhBYfDxWMoRLLRtOLS6lFBJneh8ibx+M0dgv57mud
estI4/JwpAi2fvngYSha4Tp+pDXor2BMZEOqE7N9avYHf5Ednge+2n38EWjWqCLZ
yy5NjSO0767FxDZ7qYBO3tS/6tZ0oG34tMNOu50OQ5A=
`protect END_PROTECTED
