`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DyEmVRKGiKIGQjdYgV/Sfgz5e2mnD50IB+EMImA7WCBgCtawFFwl0QohRgzS/VG9
s/XeXBSUBc1AMmitHnaFFVPDzvF0T8uEjIi+ZodKFPnj6m5Rpqbz6k4awi7D58Ne
XqXfs8PZKt5itNZjLEhWe4VHSsnoqIeW4h0CuJxOQJnoIwwKQ59QounlAJMg9OpI
XGcCuk4mN6x1/w43t/LuC/SjeOFOMfiMC6OblbdGiBjTwnMK+8pE/rApgqtSx+uP
3/D/UGWuDkyQF+cOHNnryLmlI0t8T+EhfqTG7qbnvQVEP4NTTMApwbnJz5wndQSQ
tZ+9RHcYmz9LG04g/1Ji0htw7etjBJN2Ic/hDVVrvufrWdLCSoj0Hg3OIBd8lpxC
kHBaUtkw4gXWneCQVJaEq9OvovTLWMPTXP1WNCPE52y2OPrn49JEMoAzz8zehylm
/XaptKk9ookcME7vpRZx/KoOmzJ91roy8xI7JiWE8im+9JNQrLrHATSpVTaRVd8k
78YbCen31mSncj+FQMYuWQE5wm/bzrL1FY9iQ9inFR3ImtggEtr7x2/Nx3fNWQGH
aSkTTuyG4FzWJcUxJiK5KyTflKaYqZl5eAaiaW2+s/W2ELUlxVYtLllYENBiQ2Op
930AzmWjSFGyKWLcQGvAdMO/ZaHWGfIKgdPCI4K9rRRGedLO+W5rKyvNaYAzs/Ie
fPwiR2vKqGeKtXWgTJYoojhHKbdRYB6Rgegi7GmjnE9BxLVRj/wulKaOq0nd2h1h
8olNTtuL1StBR18df5ZK3KjaqtV9o0djkck7XYGEN9qLlgc8TlBJcjiVLAAh68N/
+7d+oJhz4B3Q+FfefjCPCBUSZcZ5Jbmr3gKoZiQjySFmziRNm/eX2AgxmI0wc4Ld
sTb7jlXzxIrBQAJXwUGAl/dncimoI4ic+o4kObyebAp5LQV0VTNIGA43TZNF4MA3
6PKcfqEcSSM7HH5Wj1Ho+Rh8KJT81wuMrarHrRuE0TAo2+tg/qLqIkwet2N2PY5A
9DM02VhIitxKl/hhuh1Xlyd4Gc9HJ8F6W7OJ3PLoBPnp8H+uAK4GLWMTtIdd1RKO
LguP7kaEyZ74kCcPQnkrx0mIPkCc4iOeoLwcSEYHMHPl+5xBpyAgra6g4em0y6xp
C875gKvHENfSPqTpxEuUi7HjhYu18GAXrkgGUnjrpbXHpadJBflegEEofkZcb7GB
nIflx+3JYKuuFWwuWpPjbtcgyQEHqkO5l1/21oyKQKBWpnCrKW0ktn0o6bNtWo6z
jBiJn6tIGbyMFVNOMMTsC6qjMw2j8dqqKv2+Xy1vHRKyO+7CbFuFv5ouJTKrHiMF
S1vIzSlPvAdClt6wPhbN9Wzk/dGVvRvGa5CXS4C6DoVQd7xACbgnICg1jYlIViqJ
CVzJv7GHdQ6FMfwRZuklsRGS8NHvS/TcyY82bBVGGZe6zdnuZkfHW9RanoPXa90w
BXY5i1VLG8ZcA7g9vmteKtK8un5OjTePiWGPSABgDiKI1R+5AEdAirT/JqnLzeDJ
r24y/o403txSrpl9r0ietjtihdEBRJAcTT84Gax3JVCw+/sKLUHwTtCfHdLEdMbd
Mrd3iBFOJvll22q3xZ0lHaKfiX9fC5rr/2+fHoNNtocg9ZJNHLMoejIvzPH+plPf
ajU+A5pf8ymzVKhbY9ub0IG4rs/pi1eqDdgTjUG66vJGRcLHc1/yLZfxXR1IW33N
hM8Hv5/EbbmDAtWSc1Y2Wup4yEI4QR3/BRLo4SWWDhlisnQZsSMilWtOMosAGPHe
C6PwMgLJUboDmnftHXeHO/9UOYVIU+KWxNFJXbKKSq1wzYJfsxLKdFWbgWXC2VxA
T66EgLjSb+AlKESkQrHNW891MeLocMseQkKJxHi3G+tshOXQN1c8kVoUW7Da1rqz
SLQedqVcaUJrliBpM6diXheSjZeIMdMlfY1JeqiL8VtbK7BJM6h4K0fyNIpd4yw8
z48SHEYS92P2hpvSu3mbB5dtS9OTEPBxS3BmtmlYkIfHYJKVloX8KFRpyH8jOQqS
uPa+0+irCs1N261ppE8wrTQCFZCrMs1dqkiyy7rp5T9T/YqDreuFAXLDvlt4zG0E
J9vUHns5yt70T2RNL9qi0bHdiT1TNvMWA6+sAkX0ZCI5Ln3OS2Swei4unh35yhd6
TxQAgfUv1fC2V8iKyLQw2ajY6KK4djDpb4/LnygCsiuy4Te2oIu1wZEukogINV/2
ToJjVtZqRiKJC3MM4ezH5UpWk5rW2X+iyyFvgAwoTaZD+lMfnzj4Auflcn44zmZu
K3PxoL9rg2kfQgIAss7HTQesQTYn/xGoGXoqvz+/+Z0S3l8HorutSIp+ZixWiHSW
z4deocArggzhTAqyA1qmkbGQAJ6Z+Rf8+tNaCbXEca4K+RzCB3wt6KDgE+uXadEO
uSmo98BEQcMBz9c35PN/5tMjyIcj+TcEdM6yXyxMhG1zsmZeCz1Okacuf3e6j52L
LIln82wKjIwj2TWTp7dvx3OGbmwz6M2LKPCghL3/runDc/K1NXM97wzWQvDHgTrI
yhNtVOj7Vn/3cknQkIesmGJJFk6xrqrTBJzr7DYflyyTFf8kjzwNyBAYKazBtqRK
Qtv6xE6BfspHdqvgGxQP0vEZ91crW59UzSsR79iM//bjYz4j60/csaqygUovyJXm
kf+VUHQqB6Ip9/tqO74FMzpdL2OrLwsx9kfvTa0m33g+ZAR7DmbKtRvCxSxcHWHg
1zI3josCwHGA3fHqcK2Fsf2cMv6NoWUsjSTbfFncmuimXaB+/ck5hTXf2ZwWZQ2c
GdCyorza+Uo3td8pt2ftkVxygESaOtVO3bzWSUjfnLI37o1h1PJ4BUDMqboauSWW
sL/8I2YeIyunAe7AIYJCIm8QAjsUoObl2SFq9S5175TSn09x9TFIBm7NlPKIolh/
JpwONIFclIm6ERuYdkDapnu9w3VEXaJRV7W+N6qNgvkF8UQLkaRLwAYW9Jaco60q
pWYsewkyJpsxQQ1H5bNr1+JjxybInUI2PczdpGOrms9gwHi9q3VAnDZzSFYlV4FD
hAPJExh84oE8SwdAle0XCjc0JjwQAuPl4Ot7LaeoAjzHJkGRrwYlzz1zTqhWa6oG
UrybbEWGuim26R31eAjS7mpMHxUiSH7A5wYi/4bNSkM6WW0NYUUo8p4xPv6B/V4v
rpXs55xNDAbbevmy3jAPpM2zPnp5ag83kkgfjbuBvpESq33eNfuuvGJXFTIYsNQd
jqW/jQvWuTlDzayVomKXAQkjH2IQLgyhu/52Fih2rvZ5bGuJHwGr/d8qOCNAQufY
OMIT//20YfsjvHsC8KssYUvC2emDvwuN2LW1z2lziFB5HQulOHS23ggMDm68I+9g
9XkoVj7f5zvlsrjbmy4m7DZkCcAtQSGcT+W/NhUf7Tx345uDro25OXlvZJp11BiF
szYezBpbIQYkBgeHZjDU4sy9zIh/oc7ecx8WV8+itlfA3Gtb6btqUOiJenl5LFPC
/QTTv5LCkvIzNaVYZ/G9hJDY+D6MjoxiYneT4ZjUa8qnzrHY1MaACGJdHoNxJEfU
HFA9K5P+0hGzBQzaJlSnhLPQO83njYbd+nAAXVfyDfHTy7Kt3dulL/6Grxko86Qg
iC0CdaL78Vylj8OaJi1m/9IkOt0FOKyKqW90Tm6KeoiZ3utlnSnpqpXJjbYzwdVT
lizztvdPzRC3ijS1YRaMOTF/ZpeECsluFrb5f7uyDD09iifcob/RSen3bYXl42ml
jLJyB52raPMWHZWaY0hhSS18V1AHkBPHDqJQkvfWwkieSL6QT2v7djm5UX6xZC6a
i0Ff2kBi5yeZTpqnUykh1Nw+yuq3ro7hgukpziltE0FwFgR5hdiD4/huZDgrO800
MsnPvb9ahaMu/+9v0PNFrX/PFzowt/H1S8Chp8dEQFXHqvNf3vdkJ8hZ20LP2z3B
NBx3yvyXvmcZ+VcABnlIv7U1YNaL9EDT9qITVRTOLs/gVUkraUYI6vUB47opeUD5
GboZ5CXtDoBU9cwmhQ6Qp534UPMZoUv2dxVFScUGA8ETabj/RmeX5WwY6QU8E+92
Cv+nIoRm4yzZtGkKYKH/TevmxnAsfRvrkdebacP9Pp1UyjjmbcHhKt75DmNj5n3m
1t1he6PSojTMlMNW/+UO2ocPMuant3dWy/lzcQQR0SzDh2kihohXq8SeFJWjHCyh
omOnAXtzEcUS0tsDK7C3oupZEdDE0TF/kOx7feiU0QWb8lU3rATdzxaBz4LhjOx1
xbuuAfipk0NqmaoGqcsT8Z65RKesKZBfMdk/ZJIOdaKk0zR4Cnb12wkRHT4YWfz+
gc8V4yVNc2B8IYgXe6LWHSYPe0v10Uon9HNXEKtS6rR0xlRAZAzhwSns/GxQQfW+
UqW6hPEks7GbaV0Ezd8hVT/AlG98zzCqLTansCNyvRj8EBQ/tJk80ZB5Mo6yjNYs
1lJbPyXJhfDi+GOuUXyLHAMshunAG0JiAmmSKnyLKuD0WvQJe3/ZrMZGiHKl0Kfg
KazKnLVqkoEnyX0WzlIPmL8//ASres5c7P9V4khomwTYdPQCtD62Cpdy9BC6getD
xdhVhGHSL0GlFsFDAts5azGmtbJ3ckB0PCShYuYJ39rGxpBPPj4JLodiHWs+nl0q
vBDoQ+KeCPRfzvL1sX7ezA53gnBRAVHwKnA4SG3VHTjrZOz4Zg2/2uVvG5yTd/Hg
sR9ctEnfwSNa71sckQuteXdP+2Km1FkCECVUDwbK0dwQXT/M0EwfoijYVaBlk3kc
qelT9hB8Sp/lhrhMYIGJjESfrZEH76jwAl/GteplTq11ojjLs11wdy+gwwSX2pL8
YOcTws87Ie7PuNbKi4HbfIidFA76UCg9Q/VrVO5AT77+P9zZvd82LphjXIaVSTK0
bfh4uqkyDN/TTwTc8mp6ZLrgPuOD+yh0t3RBoPjSDGZXH4hDuaSjrtO4OhMMMJ2W
AWhdgbN+R/q20TLQQW3EHG1I6u9+wsqCtxVQ2pAew4FSQMHIJHt1EGJbPcExbkId
S1QUiE3L68131B6MF8EwnOTlynPbBi+y/bdLTrsB9yFa/SEQqb7JID6Heryj4jcq
Rfhqs+DWgdumzvyZHDvSVc/Ov4qk0T6/2oPhF/u2ONfon96P7S90wke+xxWSA4b2
zafBvtFK3+6iFfMFEMQeBSgvQIVZoiceft+cSi0j4kNbFZELrvcIvQMOkyE6xDVB
CXQNy13ohZfIO2obVTM/B0eEBKbGB5fu5qEpI8TlWouV/D6+q9+wywL4OeX3Qe+R
KP9K8j14gLK0cfSmZLeihbZ7/nMEU1lJw0cDJFcYOmcxVVSOUAKJgfCGGesiaCYN
fkvo3UR4igB71apPE9jfUzcYe6K8f8purWMPuVdlp1Ql5RqonavcBXbhn98rqtWP
s4YEXylbRvg2L5Cj4wrCL/rYgkm/QhYBkPX2wrR7w77Mrwni+hod6mYvSlpCYx4R
RFLLEACkwQLENkDv6XnmbLacnWpVN98IgR7rie1N5KSZI2xohg1hi/lfKmrZcOqo
pAxK8nH/vBhyEuqLBhoIDyhWAcHaGGA7ft6PIsRo2wbtA/erNL74/TCPOelvM2l+
BPe2HIw+bZOC37wvJaMc02EoumOFE9/QkNxdzUHtrppdpJNPbK/ktn+zGXss08Us
xzxNDjpvlZGhpLdcUqFjtBUUc0J71PLTv1c0JyGjLf3VJNykBENvwmRmxucDl5q1
+2dIWRevM7o1JJAeY4CeDCxbrSoAqAxbXgLI2GZAqrRwuBPXyRcg59xSym1WeOBJ
7SZf0hW/T7qhI4HDtZQiinM00hH58lP6z+EhS1nQzLJhRKposJH+RtS8hvqqUjMo
lxNl/AnXTlXZKzfAeyQo+BGjwI8xAD06rwndJGPvd2bUg5ajlm50ZoTHQwW+/2Cz
ivQ6IFtROvVEH8c75aaJGvdNoI3QycKXzvGx2ypYzTXcZJaSLcVrysoSDMVeAJa8
cKyPGH7wAreOtAO4LHGbdRYGvzj/EzWwfMzxwvro0JG0C7nwsFF1t0twQJYw/Unk
n5PZchrZXouJWRy7fgNrqigtrRdKuc5kNFn+2gVYeniE/RT5JrsSyyoDYG+mxVt4
vWbrxB6N5okaJ8nktntKd6qQuNYIsjDWHUsmYJ80MAzpNTKg+sGtj4TdLqr0SLvQ
C6nzj6QRac2C9Xcoxx2ZiGjvdXYdS//jNBRAE1er6YQWmHzlJD865UTC8eVIQBRA
P+XLLIx7fbDXO/aDXRrkTSIEdM4QcCxBKk4A34mp4btw/LjKIAfZS6CCOLL+Hb3B
DKP0Dea3FJRigJkucF4xkpa+3Pvlzp6fg4sDFo0HiRGzl/fDyk5w/i1Ft+6aL70M
UDOqbDqZqMojl9QvaBVfTXYPRsaYZz+0kM1Q/OIIyaN/xTLgoi5Jwd0g/0m+RiRo
ECW1SDO6bB0K7y2msgfPDlnOIPD//ZiZRYpy5xapTdDrCj0cW+nkU2rnhFkGAH8F
M5yLaGMkQaBPckyTtnS2jcQc+hZjtj8bi9hmSADBjGVtUPgi8li8SVPLpwd1/JTR
5qHfWFhRIWUVCvAR+XdjCyf7kQfE+lzeo7JBIEIQJuPK9h+TaE109L5sj8RXe2oN
uQD5y3qwr0sH6Zf/KywSWilavVUR785O4MLa9MfMAx9qFXK/4n6T5HHNrCAv7s4s
/ufl8DI7okxztZCrKfg1IlH1U0HfvEAf903HrNCnKiIv9D3TEhHdSaH1VNEnsR5E
K7Ctp2dX9Eay5NQLjjXDeC0nPCRQpT4JzzM86gCj4OHxoCVQmIDz3G3GvSFHmMGv
uPxVPdYsW9k0Mh/49iiCazjbXKar/zrqNRrja5/cxETJPPkI5NgwYidoCNKk32ax
je+CJixFouhLzw5Cl3GypgiTR84d4/vJke4arQkx87P8aSGm6xndQk3TiOxL2wuf
WqKIZsViXMlwmYPa97pGmtmViajAgIjL15gpX0uHkfFf64CoyomD7QRIUet2xBif
hQ82OsLyujrZLLAxoSUQueP9fcKsCjZmet1W4JGd9L5sdNgTqVV5oIk7g7ae8CgO
/ExFQyzB6OutZX0f6HHHyki5pSkVWfM6Q5iKlCbedxEDiaVXW4JDp1fP8iJ4cYMC
LyxJ3uSAReEgJJZuYe6RUkFp/c05CmLIOx8+jCtnPSDaBYlFaO6xwCDJOa9ZppxC
n+JVNmYk7/GE3owqUqQHLidCLGsVpXjRIR/Bx2rklHutA3vXxdadmPDJkqm+MjsP
yIsIOOMVO9jcA9GQX7VCOUBJdEkUDEQROERIWCslRLgu5s0LlSAOo5aoY1KyNbKz
o+E1i/dM3mitDCEyDRbcw/erY0cGXpdHr+MGkbK5B3Lp0NWTb6NEg5jyjetiS2XS
yR6Sd4POMastu8nasZP7zNLr619W5Hqvw5C+O2v2pY3mUMsHTn8/u/vs7jwUI4tK
dnUQjcBU9M6yzi/I5u0ucjc1aUP/Kq11WBgSt0ler+ojRHEkEttGdDghr4XcHMI4
obIbggUf3IirZxqkZvWOgQhu0V5heS0Oqk0lWkCyO3SzfggDPan9N8grxh+gARMH
1VUtYLd29n6Uc1nILxYj+f9CUSNM7/7exgz6NWL9MCmvk6Bu/SUlT/6d1jOZlBrz
xuxIydAKZfzSP8AKgW8X/2fl64+fcweKLeFwQ8NqyuxgnP7ZE2z1xr4UaJ1fhodQ
fSCBzFvBxyk1MvSK6Gsu46bVI/bxJSgSJcgoVfhWZ8SxKhsJ6tZau14brW+LDx4/
l4j8dVY1oFrixQ3cbFSjBIONVmWlQQX55yHyJ3TCRppi78YX7AYv+3/JDyZY+cPn
6HPkhedevhvgzjfxghmnCKeLgHTD66HHG5RS+29YGSvFUoPccxWueVumSnBqrX4M
yul9nFpeFbxcvcjSwiXfc2eKLbEsatV/XMQajkRwFJ3pAtcL+GkacUGRV0TvRib3
tvOT3BY6CThfM9noY2XWlBNvfDq6nYoNxuWezt320ZwBO3T4GLCQpssojhvU4pZ9
JucjJDCVzGVD6gZvHMzGeZ02LDVP9sJp0F6ed+6guDrhSvuV1WqCP35S4esM7X17
8UG1k8dQ0QfQl1vkQNczL8EELdDfhBagYboVFxOBJbljtZkvdzLxx+0/xhejVLyd
fP0Qv9mHON5ixQk5DO+R+QNJQaq35KbroOv53ZTzywMLmD66aCojUKdgF+ehYKGf
VfSOHZBQtYy5r9CVY7y20RwkJITei+s76Yuw1EmtGmbZ2HKXPEJWAloVXn78V0U5
WCfk8arSU6thc231rYf7a0hR+eD9Ii8JyMwabuU1RVLndc9iEr1Uc7YXMc7zJnR+
xdgtIQIUbBdIOGLkLH4n/wV/J4dA/l1pqCbIe63zHhU93p7UdpoZgkN/1Ig/KOja
YvICoYk9u1uysi5AeWccSTrXSeEXGIAf6HZ199yISITIlhJaCwmgS535BKxAgR1b
TqzkkpAWCyRmgQ90a1Jp0BX95qNxi2LRz+I8OTtwdXjgxLgUeF2z/xxf7B55vfXw
hL+FGOIFtnOGJjy0eHuy3NSMJbwSRXnozs6JW/HRR4sCRevqPeRFsF+m34Dde2wr
m1agUJk+qAsLVDCHeliyuqTCSK7pPx7BV+Z7824ZIP0x7VnLqZaH+DJhQb4DMm+J
TywVFgoscPWOqGhsr1o8u0Rf/RyTTJqHbtjHw0ey+nsBplMxcYCzttSixOsC/NvB
b6W2ocxq8nb15ArotAaktAFJgV2142kZBv+KnTsT8Cma8UJQwQw8Itf0TD1WNutj
apidhwZcmMLyBoCfuwgSed6hJboqkLO585vrnbqrs24xLTcfZxqHkxMNJRVVP5nk
0AOtzlmbTtYtOKMzUVBvgrbIS+kiCiKro5frDa6+EzHi5wQeWxLWk7t3azqWnaJ0
ZSflNlIhM33QS/1iug4yRQ5YgAgu46A9eDLjmG8lJGiFdbxHN2vkaRsRUhCnJf0P
tCBPqdGxNnvsg81Q7zi7WV+41yw41a1qVPQDp/eJh6qLol7X14azTcpunBa48+bX
J1tniUq3p5HzmPs3L2PqlhVBKW2XiBhHj/0x8jl3PbuASPIlmxEkazXg6zeeNoOh
Vzh4oatG9/JOODTA8UOWmq0JuaFNXIBkH1BhCOyq8RV2aYz7VPBFZxmHquMD0S9Q
dQeQKwvc/9Xyc/K6SUaOgXdccj9HyZoTnu/SyZcApovUlihUpuEA3T+MvlU4EecN
EDVF4vad/y5oXhCbsnopC5VbRsgLpttteUkoRDlDcoh26O8oM+VhUXJjqxfxr3Cf
bBi3PaOh6xVnqbnUvgQ0eMqUI4byPKnQRvPYhgRku99D2pkIATGn8m8RtBxtP8uy
lb1rFD2eyKpdcmD+gFSgr7mQZo3+DpZvfMHXIgog/Lb3kZImDGg7btN1dduPI5Ol
VVo2E7kTaB++UKbemqJ9r7aFEKhddq+EJbffiNcWVDSLQLK4friJxsWMP/t/3GmC
A8/H1s9JgAX9DfeN1UIPuaUIWwhbS0KSuL5bHUi3nLXO/iW1HaxAldUsRa3DDpQ3
B58pdC8jwmpriO+D+djFUi4mEo369aU1lQrzgXlbE6TMMDn77uJt6fOPD4uiu7Ub
5HaCLZAMcojdI72exe7bm7gxfkH0DwirW+QY8Ui1aSHDabrepOEU8nJ+zSAkfUSF
qssk9VdBkLS3KklCv0kfaIdXGIf1s8FtlC1zok73rl+33f+z1gto2ljg9Z0ZqQQ5
onKEPvsn85cgmcTqzPfcXDE3ya9X6xJukDH5BOiE6M2gsisZPDuK4ggXPGub9SqZ
XfdTa7s76kyPy2KaVkPui4UVd7RsZ1wZ/avxLOEWld2KQAC0Y/mEO6Lsuc5f+BEo
LoIH1UBDCyaKrpp6Sf41BlOAdf1YI8k/Y5gf9ulcahv5HR4E06VrAYNZKkgepZiv
pYNnzbjN5/VGN77zsYNYlQvqsvCIRmgHfWh+wzNwoOYityWGp6+ZBxzU/N5okKzv
GT1iJO31TzaHJ+Qkvb5eiNLNtRzRBeL3tSgVkTmoAHwrttQpGdrjlNN8n9GxIaRr
PxOaEVSiH+gm+83pKDjJUV7r5MVSSHTGCmKlVQqN6rdgqnXBmw9st+7BIh+E+LsP
pAKYNMFtqa4tzu65mjgv9EdG4hSYYteeqJSL9SFjS3s8E821zKG3VxSch3lb+iaj
N8czS5DkWgi+8xVhoWSxAm0MC1x9W1vgZdqGz+T0FgC+jks9Zgv127q6YGXacTr9
mr4hc49Alsq8WcbBnAmUV2G4iLPlU/IvVDmtsrC9aIgQN7ro1NcXjGlzp6oRNBgP
X005lRjtfYRHn/UiGlL0cEt71Sac8BUp24nI1P8H/4EZm1RQ8J2chFuN6XWul8vF
FuvQevDa7t8T0OvyvYbBkVLtDDhstVWxo2fElyGEQ/6IzDD/1MPz/eVOjVX89v3q
GCCtIoS+wdq+NsVtayXaXQ==
`protect END_PROTECTED
