`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oASJRbMYO0bt/3lek1kh+lBJS9D1grDjNZ4+ybAcieiaucN60sV6ZpunCr1U8512
uUcpvRquXnMCrdl3Yq/yocyAcFWY9NcaIxeTUHgho0m3bwdkxWjEBhrua0pGuiDD
lusdtw0N/eWhKNCGOLrAYkYjgZeFpIFsH8hNY7JkE5FdPG2bGJpikbQH5cJ3u7T8
Swip5bAPWidTEyw8jTN9/9df/oEvkIgvfwYoYj1XjZ8bo9NGsZa6ad08+w96I3XW
pUA0yOolwc9nqLMJMNGfbZXwF0NomXRKhe8QaGYpr0UuR5QEzxhPpbNW1CPVF9Dd
osL6p4H6/vDUmqHP9Hct98mnMP7Sz7mD1iqj891gCzCK+/qKte+gnpE0ncZEdwOj
5poft5HzVnr9Y3vrrnTK2HiNwOM5HEA/7dCt0k8lnkvLyq3mOAYTNIlIMN54boSp
VWh2RwL/c5bGQ7lUe3uQ/qxc4503hlFLLDkSlzDM+1psCU/7+GeAI6biuISU8o7V
b9Eezt7ZAru6t82NB9KjYHrW09Kh+scq8F1wq6HMMI297zyCqrzVoiipPyHZgQIq
hKCqNLq6wREgd+apNwg6WxhBhliM70nwpGrClc6SCk48YtG2hOxdVYRcGxtWLyQL
qo5n4jkopzOKHXGsIfSIUZND0qKwx2Ctx+WO0eArDj8ZsYfbdK6Lflw22gs6NVkF
qaZBu0m3fjvNQP2PfoDlc7F6d5DOVY/Sweeemskz94+FZctC3uG3zBzb0c9nwtny
CxkiFaO7E9Z/IQkB7QoR7wJjzmEg5tuXjuJ/I4Mz7DfT0kO2QmSuazmhJSvK4byx
fv/EtGfD0gLRBRl5wPWhpqPL3qO8u+uhg82yamimF+U3cUae3Mm/vKMuMCFB6QTl
u6snT6f55rp+l0sGE7Zb7VDjE/4tP2B10YUEe7Jq1NxhrC2mxGDa9zeivabNOylD
1KSuQJc5sIshLHZf+JvBng3uI5Bx8Qktjy57WuYTc7D4FOa7cki5oXzHLalOTDcT
b6M4iDMhQ1L/WRv60M05QbIRk3rSXCKvtkjuQGffJhPmI1/+61jSPdGa2a6rLUOH
/LGzTC/yIWEsbeRKjd+yXh38GuRPVeYDx5FgQyRlKnQGEpxazhJgkkVAk7e4AuGf
3Cp/FvjRTfH8ZBKSjg0Hz4mCiX6TdE0D9nCJUiE1D2jYggbxLpB3vDlO4jcFFDfK
OlPtOPZrUE/iIInZj0x6dNPA5dOsi0WSKZVdOGmesKo4uM1NpFYTlYpYs3Fxf6gB
jQ6+Srh7leIqIGk9CSjXMUBICnklNdgHuRF0VXcGuKSSDKqDv6EdIwMeI/nrB8Td
6dkpATD4LsFllOGx7uBkru/hvhxt98qGMd8CI3EjxobcSKGT1ivU95kY0BMZhbju
xKQNXCOrPBhBi+xENkBOjKHyQWkdUXOZHroFl0DrOlsaWrSeSgFbhhMNinnSy3Ba
+KLzTqCAFzarwJwKKWNeTtzOatPZWQABhRHAITdVmlJ/nmjRpiPeWLPUymcyLFZl
Ppzpbq5tXGy9QVDh5w0OnEjlXWl4Grc5Evnn2J1PnB0YNZBgZCfDwV601ffoZIM+
bWHQ1maE8fsJmWqqU8uUrjCN3OftkjeBasWFwxHvfM29RHJoUVPderlxlsGIs2Dz
nQXrbLvvnB43Q8EgDqoDx2fuRDKew/9E3KYOAfeeqRo0lI8ASIa2uGk5/bcNpHSW
EwLHFTND6xo9SrgJC7BYpSNwWv0yD+OezMcru982btZqGRiTO44wU1RchxvCFhVi
ypIqLNtuwZNJ1KeUkVDgtxGuE1mVCRxcspcSMNvg+0H6Ydl16ZJFfnuU/JmfieT5
yG1olUm+JuZyRXKoSevQGifY7UkxTRiRQl8taCkmcq7xCjmH53Ex87/uanee0eQp
tSTBDEaEC5LGHBp5vUqdml7Z1C2TP7BkEl43XhS497ej/ycipYbYBIUZh/L2XdAg
v9iWkwFJZMKunjWqTDbqPrddLEy5sUAweMPTwSH4H7BtI/JZTHdJ5gLIiZn4CjY3
CtFlsKfJa6NCxjFCCTmqycVjE2XrGBG5avuAq19vbCaKnqQJMhwbzwGAj43n3V9X
6bJOb6MMtEx8iKNXtBD260mIUOeEe4au66iCRhvRLIM4fNK2kqnBwOz4rwNZ/xQw
93pdIXe5WBPQDYYQfrheNDIgh1MMc9Gy1j08wOxjih0AXftD44tDEhA1EhyGtEQ5
9kydqev0haUjY77Vc0HnQp7IOdAPtsYhRjNv+uKJIlcIW/p60J5L/EoB1XQF+Boi
2j333qYAXoTKg6ybEzlXKC+Hv/aMma8uFf0KUM5H0C6mqXvoQ3z+XPSd3lg46Fi0
urwoF6sdAAMMIIGCDs2xCCW8TVfUYVdaE0Fl0X9rN9vJjwW1llqMayGf3x1vEq++
Yao3t/pXfIy6aU35NAt+WtCeSsLfu6CKI3YZB6C3RKjGAuaf9whdSX5UnEocoV4k
zv0YYXvfthScEWvsGwaGB5AaV8ZbZ7u/kL/VfpYjkvVfrAO7PGiYAishvCmIT5OH
jgUUscNza+T6fcg8rFPKTNDjCdp4uoBUXP03ngZnuGiP+06bIym+QU5iKQWcINHm
HeOxjlHYX5x6xXYo4LFrnCxSBC4DRttyXhmC6J4SLa75Lmln9f5KRHuHHpM6G6K5
GjblGOKszA1Z17UdMzjF3CbT87KDl4/ZeionpUAxGFt3flrO/HMw5KjgJvcxWIHg
+HcfA5FZ+aNZuZd+nqg6+nRtYPwvj3QBlf1F3nOoHTmGxe6h91AJnl4xqIeN3n3T
3DvZV3cgnXczpmc1Jt/WJZj/cyEW7s9XxmqH5RJ7i2V4nO+0vwbcS0xCCE+//6Eq
6HoZp5Ic+I3NinvC+dzKLI8iuj5rY6MkgfRbjuoJFEvH413dvuOMkBVo6tK0qCBv
WZJcgNAKoTzS9+BuqRxfQWlPkKDbz7EyA+gMsSuUun6gEvoH6Jmp4hjoqyCekJI9
qPHLi4snR6coOuc6p7IWpjalmlzwELuIwX3va2RifD5eRF7sTS34i+n6U50+PWo5
BoIiWR7odtk9DfFQmZpDgDhPHHAPqXTdrpooGQpcmdlTeLLlszPJ9jx738uy4k5W
SoyrbJjanwnNhRfCKNevR+Y11mkYgL1p6UlvoHK622Yx2wGauMT14Tgw0M/FZadr
DFwrAZZzreCBU2RytOASgnKCIRK3zWJolpVNty4eiZTdBzRyMhBcPEoC1Qr05mic
B5+o3MMP2Heo0yNVilGr4I9iMNwXuY+xmxoU9OXUu3ajhwgGOEGx+KTy9kHwpGL9
7T2BerUMv4rX04m2h/j8tPEN3iQqGp5C+rlxCeuOFrskQqLpn+5uWTnYVjSB4p8A
oUcjMgDk94kBZGTlyTPj7lV9wJrT9tW8zMb/97bzZ7EMC60zYETBcriMrL1H2t8V
iM4JwF/+clH7hbtnadOo4ZR4ywVD29rK6r5/eUMSVs8Dwnn4Vux5H9NEIrmj96ot
p1Cibif3ZM9FJsNxtzL1vsZPqQrtxBJ1EIS0rzO0fLoOuoVv4M1G8kCRzY7WzhEq
2QRwhrt0RnplvStJVsbu8Toa42+OjRb27nKqjaZDH3SI0I8H9ua5M87pNKdsvfKg
5NnqR20clqASWqCtPnQUNc//LO81hvczBmskg2P+cYvlAYD9KLrIAYSNwrC+MQhd
FoxIA1IaF8HVARaUs4EtTltXSpEZnYXPDNQWVwae+19CgcUST6kWRk0EMLATU0On
9BulcoQudh8NrM0VSZX7OArjRoo/PnE+Rm1rcx6chabbUkybl7ECE2EXIvfePp6e
q/05yN+thVlCMtJMw7Qu+eP7qzcNO2XF8M10puLSPVdnu4aC9+i1zxwUxElTFJZ2
g9L3fRGUKc61EQJCDyxiFE1zanq2GLocdr2mWr53IX0rjnTQCzSYeQS8g5ycgZX9
y6A9h8lZT4emZeiXjCnbf6U6cgqUmTWkCS81X7pjeYytumRHxiMY256aHnJB4vRr
7CPR3Sd7GuFeb/BCmGMwoZo0Qo7HQyByFxtYthgchIfrtjXgVUQeyC8s6pAlEvBI
udbJu9p5tTIP+cyNyBqoQFeWAfRCy8y3Gf7EWsvCB7PcmxQbXrPDPSl2mb3tMTLB
LkCYwSdyRg6Sc3zwDvNk2aDIN8QK82Ne550gOmglJaiNeJHmUF/Df8CSYCM1qfxk
unNurPU3RlyHv8gBlW2oKg/dRXd0vUxtDDdxtUx6CExH5MPXop7nU7/6cQ3Uk/se
Cerm55gVK0XSYmnd5aTrsMXmPY59WKpvLFvHDj21bmVQjpk8J65aM7B5uIdbZb6+
tSPTRoGX6oGnxSZm01XF7G0pOOpObu47x5f4o+ISS7FHiPjgdWGdVS2njkiwKB3L
7rI0MWpA5tp+g8yAXBIluVKBdJNZPWfwz1MEKYO0ZWDCkRG1TxQSD2rtusrWEhi+
cRzOr6FlVWzTIu0isCYGccxfPIxphOlFN2erRahmQI+qPv4N103rDAxfYqJPh4TG
ERdeU5PIz8k+SVKxbcefbYklH0zK2JGW7E3HWyzxCpCpfF+Oe5HYhPKAen0dYPC4
PksLLs8FDicQcpkrM8Zd1nT/qWCrm+FEfWABCg+OoIng5RyIYjXfAtZ63bRslT17
7YVZswYAgdG4jS7VFL/hEk/9z8VvCEjJEh9XzRfviRVUCdD+wmhMHfHhEnZ2O62Z
JiEppoG0/OXYhdg9Vi+Mz0OXr3o9wWW6E6RjXU5/VGl8jWl9SgQfvbCzluoDFzEe
RDm3Pj3k0jvjRyBeLOyzUWqe6rO026LBYed/WK0Y55zFMEr5HWD/Xz/aWoXPY2Us
RcqfEe5mewULy9ziw7aq25mSzVRYesGVhd0R47p2bqZdlRjOacTXFb6qlKGmSJPo
rDOIbwPAeFAyhD0UGSF/oDbZ2KOX8VFDyzO7L/tK1z/HX0z89w17kWcq4oW3YJlI
b5s58y+W5IAXAKpqIzZGHIFPhqpVSFYxGU6CE9kADrfegMyrMVzgRD+51+AaQ1sf
2PVFF5svizNV0RwGF+gKZHGN6dFKIC0UzFIyEGJXbcEnzizfZFSxUV0srZ4tfSe6
KpwM/15Qnpoua6bI0dlPVBAdMXOtGTFiiYLIjTu7z814SqXI+YqZVsM72P9m6Dac
aEEiu5uu1G8ZFFbG16Klyi3kU3hD1PW8hrNiuARd9t04V+zsoe+P44kxrASKKHwm
Ac2gX/x++zP13tclHYdKeaeRvImTV2AbyPoPaAWVw32FhL8oVwhgwPycfy4PpAfh
QWIfJrtDcjnKHCXvzEJer3H0C95jHkV33zMJ/phRuMQ2vFRGMilGJbLHDG1HRsjj
6CWZNLyDH6gt+0xJt0CnX044x1dgLI9+1Yi8tlGzTL/8wMOBQ94e3xqxjLxjY1Xt
apSHhmgugh4XO7fcDTp4ylUyP1jmR8oJ16dTSwIXzuPx1PhQZV/+9g4TBuJAMBZM
WQaoIJgYTm2A9WmQfBDX81zRA8Fec3hnej0IS8y54XBbscDvjVG1CZnDgiIQEV3d
S1iWv2Kgce4UIn4a0EKMXQuY5zHK9AMFtl7n8rdNPXvL1gaEL9In0JaPGzN49J+2
S6bQUMTaPLum4e+89EAP8uEBg2NVOZfvMAf043WF2s0UiXgMD5EedHPSOmk8pAfX
9H/acoqpMQJ6zgWVfRQ9hDwrnMf1bffp6D/AE6IJAIXGF90RJuUQ6vANnbhaJdAL
XoEajxeZjJBxqaN+NCBnL0g/4vXgWsfBFYvct515Z8NIsRu1C7mjGSunhnCVWl1O
CWDEmfZVixdPZfY7oQRQwBXrFP/nAgqyAIQfDnHTKb3i0gSUOVgwLCDrKmax5TOg
RfAqDl9bpaeLKKlgRsEGwjqgRv68eIGNutcnQx/Y/CqYh/pdFDU7xB0d/K5/kT9d
ULCOMfoZsq1HsHab7+fiFW/vJHs7qyksOzIxNB82bcHSLhomUFLvNXwOC7Q3G53I
WI+//XKZG6Du0wYxSnOd94BfG0ymrgwlRxWUUOexr2BkW6yxjH4AAcNLj5jZkAp8
TbziCrCgWK4jVSG2aUuSHUo2saEpgxmLiQBjAraUUs6SV4XQX/6s/qBCh6UnKuRR
VxYcZbHWsxSIZ4iTsjqEhl6M7T0tK3ZAiUwoFlsvga89i7pHfJ7bcZCb6/zJmjeD
2Qq0iLXMvOT8qcPZNz0dQGmJluh6wWyR2ppE8sNfNcJYGts4octrh7F7DilUqr2O
lX1dMLw0Uh/d9p5pgH84zjTFisjBXhIIKjsh3AqIVHEvQ4V1zC2TtiIrD/dk4re1
DWIdtNKFzhGD57+0Y0ze7TBWnPSYwyU2r0cPf8xvkwZxDsJaAnUnijg7QMEKZVVH
S3rpVabZcGIU+H5h2XjcKBAI591/R24k4PjNDaMKDld38KjaJ5Ve6d7sEEc85QVg
CYwZ4FNWS1oZmVt2Hweq5lnrSzRhD7MlaKtWOciRAmvJz3icmCLiOwB4LFmjp0ku
8tFu433DmEaOqrjkWTRakgs6AQwjcHVajupWqeH+mix7+mEcHNt2SZ0dEIbf7YLm
YigF5Me6WdReGfKiZpIYHgdJzgx/+7z926+s1UzyH2rBIvMuUz8DArXqplw4k/K+
M7eft4rBjOkDYFsiBmz8Lv9IeYlEHQBOStQufpCt9/jnROgSu/QjrAGyeU0gz+W4
rQ7NsPnx8zTsm9s08zKYqHPbC5eBNMi2a++pF2FvOk9Szd57iQYJ1RERqaex63f0
09iNMb715QgsP7Pc0ozJsn/RQxBFCutY0YZtdADqhC3sX8LToDCKEdZ8+XXv9tgY
rPx+9iKUGVdTQx99Wyfz3Ii08XaXfhpvBLVpHGEEuGTNwEUXNS9iAFy+TzoJOtI1
KQ68bVJP6f6+hcPDv/XHKHC/boO4FEKqMMSGqLbOm359QP+u2A615CfT4/PwdgpP
1apbR07uGkcqDjKNKum3bO+sYFouzGGu0/yLHQ86S9UXRkOd0foYfqap3FFXUcVe
5tdIo322lZ5Zc1m34kf3jPI556DQNyJVHuknZImqthJehoJ8L5w/Qek1w5w4vGDm
YzwZUjvrrJh18TPZ/ayIBfgew8eZlQhlB9XsnZQaFpWGCUZOa/BR95CqgpIcacOa
tXcSTzu5Xvy0jxohwdKcxvLykoI/8wuj2JvZLtONs4zs5mP8JWnOADbDk0Nl3Q7K
NTyptUtBTl1TaU0IUltPv8XP2Mfvzi2xKo7DHBsDwLHsaR/v4SbFaSyKlzUTKlDq
n1BHO+ETycW2vIWw1HK7VwxxRUS5m3eucEWRWusJZ5qYhcAIJ+J0zHtDrpUQuRsA
YETyDrOwRcDr4mtrLVZBJJWxrXV0IxkDYuCEF/3BgZDMvZAOEVevj69x/HXjG8fN
JpkaO/4hzRrVaiLjqdTGJFn6qVErWh3Zg3hxF5LuX9saNKauZH84p/0B7nOZjp1H
jR34nA0RlP+YwC50sNmHs9K8n7/BzvHtK7ZZ1+n51mxxPsHlCd/6g4IAcsw+z9NU
W/tTRQhuZrS/e66JvZrIDZBrpcpHpELChkTNGrk13ABMqSwSMobya0v7s7MbSeT+
wmijzv1/19Kqbduvw0DD6hxN4/GYsg1vhOIpKTr4FTokmjyVW6gukyPjy0nb3AYS
49NmI/AgKvWJ9b8n/ScnmjurpjDjTOLpakVXyc+hVMLcl3aaNf6ySfbCL5q8YD4o
pVWeFud6rfyn6PvTplvlxZGCOdD/sDv8IKVuTx25THTFpvkZzCFbSRoubCpiFIkV
qW8BUIsneu0YrBia2lYv0CiAxJfSfZiPHM4OWJhFYi9+p39i2LkeHg5rzjt/C5lt
b83sp0Un/1Eu63jnJZa4gGnJwv940iIOmNZF55Rs1Ii7VdGxVltczilTo2886vN4
6EwiiutvxTkqxpmU+X3ZcmI3EIvWF2h+DwyENNFmlRcw2gSmlbgb1XGGerLmyH8H
kqclfg47YRN2NBmy4rE9GpODGizIu3Arm5BvXysNG6MB7GIHAYtm03Tq1W4qNs0M
gXa/ex/bD8PY4kqr8TwibB2gXtMscJJhn/BOovgmOJQ8VnqLLK5LSzt2IdIK/Bi2
b1co5gwuqPXwsJqzAech4JLLfZG7UeZd4QVQr5aU02StfdHywT7WUCrNZLfhno+4
SN7xinjDq9DUSM54AnwW3CbCmDOxU/i/VBgK8TMRHv/4t2JgpIk/qx8K3O0cDqxC
bUrVaApluyYnrHiTnFBLPqegcw2ayBFq+BOzInVuBHDjWmoI/B47q8vuVsCFKSHD
uaUFrpAH+iztp9Sfrqlny5HQTk2qlGs6TYkFTVkVOMap7g523Zs6Pb4y8orFXHt8
AXlLPtlIvUQ4/zLNrFkiNSqjYVrFMAvngsUx93Pw8ieA+m0OLZAr3kAxjQjOHdJZ
oibGcI8XFQAe2zuJviBDu5aOfEL+NuCtbs12KsTHr0gpon04qeX4MV/zCmwqWatT
DpfwHXZTd4NeE5na7ZCfNoz5o9dokZdgcdS+EoChux0plK6PN3jXaCAv6z7B0fr1
VSU9h7dLZF7hPBcOlAp31vsb0AbL0BjsaTA2N83G/1FthR61cJYHL6dQXnkUZnMQ
nDXgrmwAKNGRMV025OlaLFJIHZZkP31n4D7WHCA5dDtNdWagzjNxZVMUouj/bE4f
Ih3fKKDpnx0oTcv8rJKugJI9I9W3lLceaPyowFz4pQOZFT3YHUyGMeReVFCdhkDs
zmwudvCU83K6WTFx1iv6sYUZdL6TnJzMMlKPiqCJ4k/9JJYf9wob1Dq9NpRMfJDK
G7m+yAVjdflj1DRa9NxEmGJmV3FEwaMSAE4zuhqDWYp61YhD0ki1CyImEQ1lolbH
zj1rM0h6k5OkMSn45rbTYJuncI1a/hmcpYegpuL9fzjGD1LYRaNpL0fGaxW70UvA
waBTrfIxhOCLJiOPUzvM06Uo8qP6X7/mu7jzp58/+jypD4Wa1TPP1d/o0VCwUnIr
6x/wvLGSL0Qr1J8XId0bpxxCQaIIXxaHafxm22rriU2Tp8CokrFjvZVJqTMSucip
CHPYKfZuyUVGSq7Qnh4wsoDBQ4ojMAqzll03bNg+VwLuphvCMx+f8xiNm5+ULOGG
T6l++EO7QtaPAyT8nP/P0URMYMEphZgeF6bTHkfzULokus3GrT6VkdA9QzdqM/h8
u7CQ/tgi1dWprL77Ly1kQdOut5sXvlZ6xa1sl1V0gXKI73YCm7T8kRLI4VziL+g7
mtOXWuDLND5QItX4ei+hC21tdt0lcpRzAmQKFFOrk1NtTnpOcTXkwyvzG1bOkTOz
1n66HFZ1vYF6U/zjxM4moS4kQf26HPvt0Li6KvI9N75vj6/5G6o0+UPc7NF8e+W7
ZgW2UHzOZD/sj1hOocNcGVl9R56AhhzVY/y2MdknaAQeDLdbrbiSLWOLtXvJXJVQ
hG7LUZcQKLE1P//lqZgWTcfJEoSPqVMUcxq8WlXiYnDax3kJnnh/oeFTRXNT5PvT
YbQQdYy+J9S/KH8bGQczCawoBBo8REuTBN6EMLf6qIyOlqjIfcynWZxooSNDGswp
1xbvj4qe8Ug0F4GoDS3g52hrDy81w0ny/AHkChL2hJ3Q3PTW2YrfRR9vLqMGcEDM
abzCbmcBu5of9rwCc60hAuHG98oZsMXFOUqBpe840nM61zc/2D+MIXlErCUSn+HE
CN5OKm9sTrc9jIA7A55IlVDdYyCS/TvE0QVgmshEsW+p2D01I8VgFBFfQledtdds
R72JdTMbHEaHeij8YrfAYERSC+UIYXkrTr8W9hFquM9oS6ApCB8nNflzzBq6niLw
f8QVoP5C/Pj3HTomuaavMDp6kDkze1iZb+/rQJJEMYMGc6OFcVvY/VJNyxKDehS4
xiywbPSrsrBbODUUzpVQC0osq+um08REQ8/Ld3NiQost9Kra3SzSwUTbptvw1f2U
iaMSfpBFJIrfqO9kMj0lTj21Q2DE8eP9OZ0rtJiGdE4sS46OfmiLO2tm0VX9p70W
iHACcGVocgy27ReI8BaSyJqyy6U9oPAE9jXi0m1gTBYLp6mrdZ4/HDlQiTXa6hFP
5HsOB3SipffFCasewbmwSpoOVwFwj22tSq3EzWSgRNKqpW/KAvFREqwRP+ThGEU2
9Wnngr3oIQ6qSq/I+3sTwwtjUSFkSjYX6iSu2LV4/zwwacJvsiS4juBLbBdKFzT6
NojutYwseimw/TaPLS26WdQEmuiwpJg66dvxsLNOHlBCeBksZusEIGNtR0wc4l7F
S6u/MOtq3FWQMwti+/Pn+66GJJvFKRIHWvJKaM7nu/9kCn/JsKLnULLEUVj/7zvv
E5OaG8ibftGuvicaLfKcuFmTsCEba3Fi2lALYJFv4o5+bGBcOkI6YIipxZrZex1X
0m0SKGUlaLKX7wZaB7kAbki3A+h7U94rzqdE6S1dpgy6TQ1CpL/q7t5kQyK9V15Z
FAwIohmXUmkG4xMU3plTXHJJeSNzHPEIam2CLsOxFIvtLeoiFWm0o9NyvxKy0WAw
+1Pmds6xW4cLgaluFP3/6DVh6s7qe1NhPw6lkeMBl7PgCw2m0fn4uvOaxCx2RVy6
mzVStVjMhS3Qzlpuwq3KlVzhhzwqVKyGuX5i9w8Xvulvi6cQVQYFDXV3xyt9gVQc
YltuuaLbBqbnxpIU7RKjXYr2kjdNn432FVjvJMHlMEsT1v56ncKHisQ9YbPGK4yi
ziQslc4WHeMPMc2VPA6FZBwVC3cLqCvkBw3u2c9FeITYOyPiIjk5wjf107+XrrVg
FYcWxAEypiE5cBq4XPRGwT7gFr3kDeStiv/iwS1bYu1W1UXNk/vzCTosku16esf+
dyRhPOxEAhNsiP5OB1dv0pEkvBf/h+AxiqJntLDVSnKzxYYxSaKtCXshpVYHw7si
S6z1/FMhiiBxDsY3Aq/+sX46ga10Xth0AIom8vfT16jOL0DMhHyUy7rnQkMTEQ+y
MV9mGbkQJeMwpGO4YR6mTt/NbzQVbNoIYWPFoFADmN7GOx3FEM2D7UTukkyNqfkC
w2Tm3A/ZbutMEDOF2jesy40s1mJ59puC50+M9eaMEIsJDPoOklAWw1YL6kmiBMqf
yL+r1gjFLwbEPdk3AbvpIWM0EG1/+gqpeQLs9PKe6nRhnJtK91eOZcXO+sV3Lqb5
sVxIQSDzyn7bW3vKOaCuD6MI+CkDAZZgqhEVe6t0zq3ueCRAD0oNHVZDOqBDv4Tc
jAo4Eo2wa/hwMqqZSS4D03/WzDCpyaELnBNR6kUsdLP521alJP+g382h3akgmI2t
/SmYjDSASyLbyCdYJL8LJvJWbjjbJkY/n/pUbhvDGtDX2m/YQToZDpF1xe4wmtYk
7XjWlW4uVA/pgjahygF4YhK2KlFw2wvM0RdJHBBFkRoeF17sGsS/MriorcAuzH6G
kBOypWSc/DjESyJX5mqduKtIhFzQqkYHHcpQh96U3F39sZa/6tImKjXMzQQIyHLA
8uoCwYWYWd2IFM7RrOZ/O5VWpRz+g/PDqruGMvlHedoQ2eLxfsqqsHoEmo52c2YH
M/YKSBr8zEZhn87Cijlr8sbM9wHI1ucHFlKGgB8ymamY4ZwWDR/kxYGH792BQTIB
hZn2K0xqY981KSfk0fN+b6L4ld5ASA+7+ZWp3PZqRAPvgHdQkMQioKV9W5EQumUk
hodhaIaxEP0d1X4jfc64uxo1TBLquDhNrB/DLR/a8Xd59shpPg+Ubfwnum5WDrPN
tyR394CXi35CRdrLB7vTXB5CNuEz0aev9sMQHTfb5dcfFL1CvaDsQ/W1uBTbAuC8
+/dGqRqAylfy7LpK7hd6E19IvXjVR691t40kCrxCNLWuvM4EsqsOnOAbxej81sxl
DmuqwJOH/qQU76cc2z58GE2lu/ZC+Jz4auL7jYTAWLVHmFrsr7/XCJuM5ZU6S0DX
U381rmH/KN5pAd43DOpKyM5HxIw8xduWuDwKBRzON7Jw1Zk4WfABCEUFe+87A/T7
3yuCKPmn6zcpiEd9+iHsIYvZRvXq10vPuvWTqCSDJMhOd6j3uhshTqyKfCPx8ava
6iXxker7b7Uq50iCMfyJs8z7NRknjT174A49oul9WY8UuptHnm8o8vr1xdU0/HbE
x31BaXby/8pdExK+h3bhuffLtgGHXiBgxp7nWW7nu6h84SfiuA43juvzNpRcXNkX
soGFAqwBSsAt8zdJYJgTYy+1wI+kqqEmhfHknYmrHgyYsLyGahG7Ukqa8MOLwdBH
0o2bHCxxAhSj1HzFgxdoIuF+H5eexX5tSPz9oiCkJsR6ENwOTEDSoO8/0mbROvRh
y4EdHHh4e+GgTf9KMyHWeimDLU8S8FBhC2xpiCF5iZ4Qrt/bZNkyNQMdxTS56lTN
YTDhSQ50o2IxVteIjlZ+T309+6X/FCiblwydtLBA3YxYRNyPCnf9efWQbjV/34cd
qwvLHrImQqo0Mkx+7ltPYMdm5hIKpLthVslbEE8gNQmODTul6NKhHdcJpCec1HlT
vE5/zhXdIysnO08n2NTLY/PrjuKf2CMWPZIcxwaBqBkdF0NsyHms4LG2+uXKRTXu
InsQ6uDV+YeHljnGyVmi2rS/jEVLgqvPuZeKELdivZ1AOE/mVbYrHtsSHJRc7HuC
KzACeoLrdzdDqSVL2ffdYz1nTk9iyenkTUnww1ufwkJrGlMEMuFw49dVAEg68ojt
DdbHZsFUhPcSQhnsamXkAP2WBfXNTUHQU9/ACU97vNlpgT96D0tycdgrLx60u9rU
oLD0DJXSwOH5ZRAGfLF9tF02XQ1ymylujSuCKy/3i64IIH2i5sdDRIpdV7U9ddjt
LCEJG7ZP7BD9BunlHLcWJTHaICFp302gYY5svnk80RaYLwfeL1MGdCu+MjXAd/1N
Mgt9/UrLnx2ydtCnu2cXXZDF68V68X/T08YsER8MVpD15gvFIlVM2lWBiyL3B87j
rE2Ab2WMq+1OtUIJvBaGBGBEsq9BARF3BIojS/kYXZkIPsHiscF03TLQQK/gt52n
U1H/S0mN9YkNPRfsfUb+f8LTToMNb4AU9l/ipqu0OrkW4UlbqAIJ06qcB40OeMNK
oYudYzVh8+EfUHKg6TTfNSH0+LDmpZgMEw3OJ5BqBK2Tu5hr5JspULhX9cZkvACF
PUzs2xKDPA3sbsypzDx12MNcShex+j8XDuJA6A5I7qjTp6OtcjLjnbzqXzGcEcc2
WIXoumldcC0sEfO1eLhdCb0+xZIc0xmWYJbET7sPTlPKUGmWSObTyGGXdfq5AzUd
9Vfxxk+45Ft1hoxuwlW7fXucbIGHSmpt8ZnF0YCvkwLlzYaNY5Ih5BiAZyvoaciX
V9DZZVgFC7YZDZlP1pQBknYXOxVQ2GpqoMw/KfYj9Ua8YAbrGSncOj2DiiKdQrM8
Zrint6GMIhKeNx3M5PSTgqiQLnqLdhhJc6C6VbsGJQHsZmdQEGa1yyA57K+LpZNY
GGlfZkyLxKH0ikY/KyhJOGrSdgJIPpfon5/cve4CbSqJkJ6z4Q4FD8a1AZe30RLh
CE8AIQHt0zkEyy/Lwg7Dp4rgKe6AmAdSoDnp5WwsVK9rC2XXHsefe0/5Gls5xekI
E2xbAmus/LD6iJx6sv0cFGnTpCXSHVEs3607dTzVJqGSAJ7eC2AKc+p3GzwUPu8F
SPGvQrWuHmu71wdxw6MGsSvV/QKSqdsZzCGFMpnY6QShl9ZAvlJFbqh/XfmgEDJo
VI2zjdtibMoQDkuDMHxfyzsOc8IMuz8y/jet3hzT2uwUT49wuvnLzDoq3/NkfXuF
cwbso2dgVgmqmCcJIWxOqQ/P/y14cWz3J3IF1U9NEcW9XRtKLJsy1pbLrnPNtdA7
L5PVmVRbqePa/jyK2p5sfmxlbpPjFhCwCq/kNexUxW7G98+vhmKBgRRbudKdYkYq
8BG80g9/kVZp8UTnfxecx+l7ZcWdLuE7cdZAjbOVl5gEc3HrpCExwMTxNEdmvbjE
uB+6XyOEqR9Xyh1g9gdUTUsSa6N2MtMqqkABf7ewklQSdQq5tpROo2PApKG2ywg7
stH49iABKTDJRnEikJoriUOtUVpuVpLeGmPIGxw2WDWjyJb3Bej7Wx5EXb6PpR4e
xD/EnS2J0J/ZFDHvh4LA8gkW1EYJo4amnFuovzZR9sCv6DpjkW72IZ0pM9l4MxGW
HDpsKQ9jztXixOUcA1SJsKHeNtCuVmUSMFrr0pYA0UL14Yq9hbzcAyvwV9zQ//ja
rDL1d5qtdkYInu7j2vA5cbiFc5KyfKHorTogqWezDo6D3vMYvxy/tYgs1ap1C5cv
CMQHMooD3kArQOzLmX6KWOf/gng8xLPt7n3aajEVhBfYJr3yGfx7xLQ6SS4lNz1y
yVctifjZndCTRRqUIBi8hT2Hahgf/qOwODe/awPWO/vWovDU0B38mgqsRv4SIwrg
y15iKa15/eflJsxx7Xl+Ss6DjO3b9P6jpsOIZriDDoUKPaDIh9jAYrzbpWP3uiLO
nDlWwO+xWwHJACkjtrPLslGAZP8ZcF9CCT3NrZEXc7G+jux3gKIqKSfMs47KRTS/
2QrmiWxGeiARaZPEQNSMd2N1p7JVc1MVPm4ibhYoV+Oabqiz00wUYsQ5JuIX3806
pYnEzzfZsxJvCZZfeWFHXmGNMqoJjfvIFamo4yP0cvXxJm35U8Kf5P5CyK/O1Urg
fJRheqhkYOG1MF6bb8Xi4uwCQFhX0IyaNhA0kOLAoVWPNYdaESz0Tj+wPc/GO8uq
ZnE5CKkCV7E/ELyakeQ7eAl0XD65ccS3NQIykPq3it5M9UJagpsUASfKPExuoGzv
YtKzX0Nn5UlnFRlE10LLL7vPzFq+fLmpYoQir6Jr+oR8I7RFdsja+nzEZPYeGNUQ
ZnVT976U6lLDRZMyndIaBhZFqnOVtpVkSwvVt51SJRUlyg4WL1B4DwS9wqVwc1qI
EDS1B2a4tMyCqgWy1XU5DdUsJW1DskDQuSzz0JPZeP2BMGAd8ou5Gih8CHvzmd9U
AWD+LKyDup7j4LoDhHYNtBAEOVUmmAvAKHUeVrAMSGE0AAeYJ3mKkjeFo8MO2kfN
Lc1vWXK/du0ZVgoFRjRZVWqGGn38UQiZ5bp6Rj/qY5BGlJ1HqV8AamemcsvhOymV
5bJ75yv0dYAh6B+aNI9HAS6hmI0DxR+F5fo3454A7I0lkyocjuRaFAPWXj534I9W
Ii8bncFl7QtFNh1YPdNC0HEvjA8poaWF2uvH56m8kzP/frPan5b370JwdS8C9J3g
5gbXv9BO8JR0Q+ZpB0gH6tl5fmmPfas9dn0s7uiaObx+vupyh68LodRN08toPUDu
RL/M4esZByB0//K+uuk9uUOF2m0rW1w0jTHJIGPX3Oj1Iu7Juy6++ZPR/smR1wLm
oQa0gJqx4LhAy8PayKmBAh7v/BkjxzHq6NtjZBqZuYYBJ63xUmGU2pKTkqf0uU7g
dJ5J1OPfc7Eip1kvmfgkQ5XCCVjV92RdYWc5eStMZGpN+V3wl9dq5tNZ/cP9dte+
OBA8MEJ4WfUyjbT/qQysikJrSadykaVaPafqpzRgXXAF1iQCnCYFs16VW2fHrcbs
LUXE7vsjW2u8ao25tZKyEW71xrbnmB/bMcmZ8nHxxQSdmamnIjC8J0D0GSBMguVE
/FpvhEdh36ImS79zV2kSig/nuDvvrN/XOJkV7U+eU8Xh5ZpbGWFzeskA9wRC7rZy
Mwx2WO+O32IaSmWQY6y50wawx60iLieS92VHlNH/Ba7tvE6PVu0NHbrza8ofcXtP
h2SAwyef/MjNW3lG2BtTieswtEkpSK5KEwtWbMhU8sF7AIAz9FJRfDySEu5+259r
Khq9Yi4QVFzB5M5kcbZJM+N9UVdynl0Fiq3+L7GYBopDIvm4VfZKHapIPGLcVIdT
C69T55UvGcL8qr4DhinWn/zifkG2PeS7miG+NRDd+DFC5Yodlt7hbYqWui6ePLN7
DSjNH+KwmnxD8Kwz0cYMXwWgX/OA9/c8oc+WMBSrWIKFoivE9zlbMVfwGi1JDrer
RxmTitq1fHGm5fHb/x395CcUHKqAjRLRl8fKpsRmDKkScvsUdmDh25triF8JwBy4
Y7PVf7k9CXXgxI77W9kiQpAKXP/H6fYBrYulJQYYuWkJRf+5A/jYOE/BMh1hTodH
Gd1iZID831dzJxnb/Vfz2MA5UtRd2FqKnBalhhDCt7JYqFP9SRh6s8jNdiZJuXqU
DZ9ezjBQUk7C4u+KddLPQc+JLaN9ZQvX6Fo5ZNkNMcQN40MElWlp4D5reQIqY88n
sp7vLDMKTxIbWoRxVGQocf+6WDsj9j02kMPRLxl5UR+1c3OFnpkgVCSWDHfVSoc2
7gQtdhHRvankulP1Du2cduvFv+FUEDj1U8YXQPYJ90zztsnXAwqzM4O8ht41ltVf
gqt3iNblSwrYivDVOWzd3wFr7Gy1Y8rlLCZ9VpzY5cSk8mrdwTHebidCgFSojkZK
IbaR2/56hlRzwYPI6vGgIQiKLzgeZHhzwsP3PVju63SDPztXbGSgU1bTc1+jkRHx
PMftiBuHv/O7XYMlw2pSaq7AwX0HLy032PpTeLExVJwEV01/+kTUe8jjhxBQBtDL
l5wOPu/Kg3//7GjH09ApCQ9QKq3HG9/V0BEoSMOCpajsSbGoEuCGZHW3r9+dvlZG
vVRR8DNtBFr+i70Cf+GrnuMD92wILLi3x1kR4fEVWg7FpwKx8CJfDk02qPtk7p3N
8t3QttjLXyrc/cKQiSLfft8/rypywaIhW+1pEpQNzdjNHDLvf11VM8fLGg6RqLJK
DW5XwU2AySr8axV4mASy+lVgJXN+YmLU2Dfui6lDy9nuC61KabAGX7M+sy2zDQi0
J/iSZcpYnpxI9aO3ohfkWtpwJLaaydB8Qj/E1njb/RziiiidTlcLNsEpeEj67S1N
O/nt4ebJDe/oVaisX+D8EY/qiNQ04zt8EgFVQjryEDzVgTPCDb8t7p8UUdEQ0K4G
zTmbKrOxg0XNxkRacaJYR4y8y9mpACeakocN4n4U5o7muOhPBM8ahe3DfWlNRX7R
5AG+8u7hTnkj36x4dvLdBM8ypT40vXLYFwvd707BlP+7p0gn/mLJm0q87tdK27w0
3uu8A8SpttOfZ9OJ7MVI3k30naYlfjbq0vdYFGnsk1fjtyQP/3ihVTm89GOUXNJi
BB6dTJnFDHxJuImRKprFWfAWwnPQYccCxUMEGzq4CHas2uIpAUUDzZFSzXQAGqBn
9UDzJRn8kmRQjOSGelsSxrIQlbF9nCn64ep/CpNm/QtkeLqZjuJ42ETvdv5ahaE+
eoeTYzLAfNUEIBR3ql19iqeIymnVnswq7eSQx8odon0sGIEtBk6NLeTrx9uL+Qrc
rXkIUjo7q2L6OPEcE6PlYZ83bSbNqMMvIBCSgtPX1sH+Fb9Agoy90lVGaUeXfcyl
62entqsHPOb0Tek9YFv2K8nYeCKZI4V127NPSfuoQ0XLGbk6FwziK3LwDyKUyInU
YqhXZa2IrzD4MO5bHiNcm6gyOEGDNVdYDgFb4mjpOxOPR8WzQ0fheBFXsoRuGHbs
brMu+O+EEP5VlVDCNFdya/wRUgu4SMthrnKQL99RcwQB7Zm34QQX73ysXP7dJPcr
mOHep+K2xq6qO7Qd9a4T3EYp9geqD2s8lhPLtme9tpsWR0EL7wwbnnWYnDSUI6iC
qt/oOZ/eIBvzOzO+MzBNWdOEppxvFaiL8dCj4dRt+2exPXjmsFsOct2oPD3ee+VA
tir+zmwGl8/Pg8nlANEznCrlcM1LITeXywZyKGdpk+pSen1YC8hbiNWhRZybTF1X
KawxN+NOhMG7FIesNU1OFzrQ2HUYRpKdczJ1qPytzXDmtMn1nXtyFjR7sL37Iew9
i+JIVLvVdjnTIvGiw5StHTFqguhla1W14meF6yZvREKgDrQAZlFxVrh4VdYYhhqs
W4ohlD27vSlzapV2byup463DAcQZbs9b9ketUny+pJTBpOcVWyEYyLZwNbo7r4r5
vQ+opq/E++1HtHDW2yqFhLCKNV38ZHaFqqmSargEoNv0wSNoZXmxngHoaYVzUwag
vjPBBgF1FuPNsm1S/YKw/0NjpLif50CQMAqZn4yBZBl4luf3H3ujBbGW6n1fRTjW
RzgFeKJ1dwo6rbdkEcKqBCBAVhaOrio4oJNBbab5kX6XB/QUC01hzbAX4AnbRrys
p6S3NIpuL+Xt79IHMv3hAZ0DatYTUhBvP5ujfjr4ycMSX5FuJE4lXj3xuoC6jVgX
BVZu0SV8zNPC0ZHxmlzIcyml3jhLqz8SKgtQms9L11OrU0tYN2bPYfnCr7HZh5un
uwThLaKu4WgSOkGnctI51m34LvHeAVidluTS0LLJVgZVbzqgLh1+t9G5ZFMo3oSJ
h0TzafCjPJGd7MeDe1/5ayn39J0yxMK3YatYyu48SDzutFW0A40IqJuFJtbP0K4i
oS6xotUBVBWnTFOvoqWMtChPnU/xvGtaOiSNzjxgiFC2t7kORWND9yYtA4V6slMK
x91hBFYaU7UoDbRcHO2O8RZ+rJE5Q4UE+BKy6G066PvaD+kqQU1ipQVNITJ9KYHp
dRsE5sMM9MKM4ZFzWTsXZfSujerZv3OB2VxufkkFEfrhEc98Z81DRVWMUaW4rzTX
xJsGVRCFCRAIl0YqzOPQP3MkKwcQf6nEmWac6Yqmb7gMX2ixw48xx0fcxz9AvBwU
blgW2+ELNV55YfavQQ4ym7uXYOofxl26mtKGe08SdyBRJSj5uofm4eWkc9IIO2vJ
ffnG4ZpvRbkvKMVzMBwYh3jy8DjJG9RwXr52OttvLV7AzcRRg3nC0ioAZzptxR8Z
Zta9asGCCH/5W4o6BOxMFSbEahHP79QQXog70Uz+CoKEHEZ+iRdJWKOIWRvRe3aV
HMQN5p2R0pHme8LjRyX+JEOEW7VqPVPrVb6ICjm6Gf/Cc5bqR1bp4QxM9s37Mfij
MhX7l7czRMftE6Qt5Ufj0l102RyTnhfSIPe/du/7j3MyUgDaWE14xzJAr5s0WSvk
NfgKdhMp5oqDKDrsgIRjMHiRtS1B/5pfd5bqNAg2Tx24GmnyBTquchp0STejfp8b
1rFn6yhFct1qtJsgUhuf3ZLlz11DGKcuwVyN5TSJsSxM8Az2eI/w+6/yLWMBbxxl
399UN2VcstEdkxQC3QAmIhPF13Yuo5ScvsDQ5q6z7iNCOHyVT14p2wn5xEZDCUke
A8+YVER0TXNjqdkSSFyY+3ZDE9JDKQ7ZQxAGaoKShz4kvevcBxzdNOSeVG+ELLKs
0buddH7OCxgSKYZSEvnMsG7+8KPZFobdvj5Ox58bVUxOKJtYDGGYer3DyztZQAiI
gbjKJ/HxVTq73AqEKGim2zBBWsuGv/ervPNCxS38GRJQpjyOalsxJ3e9ZhP9lYR+
uuI0h68fS5GEixEsfE7GJ4edIPnRLsP5VBheQgR8bvYDVbQeNapZB+Jvm1ipAQta
VFOvFcq9QrHIxzpMQ5IXpldPnPz8WqnhU4Pjipp/ezKlMICNuPvLpO1PQwXiPHhe
`protect END_PROTECTED
