`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bMfofgj7AuGGiZfTMYvJdQSAR+NxKixxTa1eCg2nJbLCIFNNtFlxlZ7D3YWvoGCZ
xzWSEDcrcKzYpSGb2yWiqww0pka0dvAnj3bAR1Y0CXGqE2atMto7nNgEkw4umnx+
UEn56XDTwdUmwhigwUKPhl2tcZ1DjwDBbPNtqarto1epiFw3a2zjLAcImOc+2BNj
1vvu4+4mafiyBgv5O898KZfP42CjGhxU5f3hL3hIGvqXghXipKv2VIvdvCY9/Uxc
fEwyQoymAFpQkb7HVErTvW/tTNuP9GCEg4uMwZFSWgvPM61J7mAwqaVA3AURM9Ad
5xi2yc0/87C/ger59Mila3jozDcfnW6DrZaDYDJAn5bK/grp2nIm4oJbt5mdtwIb
0GfSK2ZqLzKj/Xhc4OFTQwthl76yO0f4pTiG+kupMchYcLCKJGZwIXUUaoUkacdF
0TyWSgvAz7TQmyXTwk4HH2KQbrWs33wjTme7qQ354i0EuP95l+wla6lNuS+R83dQ
WgbQBU8e5DYAdXrOi9VHGAbWriiS0VBR5b/mWZyIzEWo5gqV+uf9YJDFNr9bTzzJ
zjCzppNF6GoJT50/JTnfbmOZQo6DzObaNZ5TV3+rVps0sJqTjQa1cJ7rJmRdGMH7
A7Lhp0Jp/rcuHSES9dSwQ0sivPWUjlbW2rtAh/Bp3deMFCIy9pwU/dCj0PccfO7E
`protect END_PROTECTED
