`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OEGn6AK2nbSQHFIKHPLv0UYD85CtM3biXDOMdXgX02mXeb5D2UOwdl77QO0Zxtfl
2IWy66zjlmEl64IsOEMDBNkgaBqSawCTxINdeE0VcVMENQnDrpaNJFioRcabStXi
MaDhLdWgotuO4xACi/FuxY6GifWQ6ZXvxGCaCqcvx5h3Jx/K0DGPK7Mxt9ask19x
zpL232PLMsVVPRf5V6Ks0xIXDrnWiddwT+LGI86pBpoAfU3/kIjez+L6e71fd+YX
E+PMQVFHc8tuxKxHbX3k9JWSBp4ZjYvFrXltH31Cgn4RR9Hs3CKiYu7cOCFeXXbP
5fHqVLY1cUyuyyml7oQq9lp1BnsBpPE6nzxaioVCeNrvvbzkI8dF4nXGTd89LA3w
YrHwkawAsrXl1hUwUVQcQev2Bi8L6gMQtLIrqHvugwM2Et4IzWfKacpT5Kml18Vn
O7o1Q0yhOTtK0EdZgFlSUTxT4+/cG6LdwG72YeAx1BuoWlkM6BACc6U0BR0P8PyI
XEuX6J3yCtAdgtnJ0pSJsLY1Hpe0aqhoJjQlsa8AeHYEWxi3NoHSSo0AZAYEjsBr
KuJeYBDI83fFOpcmL+6nRnpd+kEtipmNYsCoK1Az+Q1+G2YnT+fLkYTp+/sefIjC
Pq4UCT0ieDurlzVqB6Ga/VxYkjzEre+X+hbvOnR8LzqsapAUr1kZk3xbxafKJAwR
Q43FC5z09vllUvk2bYdKB9xLms8ppGdW26R+5fXm56te4AV+aV3dYmC6Xn0E/tN5
N2+wOziVNPRb6roycQwRVNsjb+Y6mptBv9G/V1ms54IEh0O1z26ii7mRx2l7eebJ
lCA6R/jxJQCqLsAV/ZkFWjZ5lwiUz3a8C/fspsbtrnrOD/BOk0YBEodyokpmS2ck
N42gX6WVvu6SEoqjkCASF0Bbxc3+lPvwGIVp6hic5euFYc2jwO0MX/uJu/Te2a4w
KeMjWw2jay9CeofR5hmzis8oMpaREaLnxPiJrzCrGHUk6jIl5JPpwo3U+Bs4Mc86
2pSNl7gdB9HR3B0vOtfBDUPmW80qqBRP5PM4FvHOypASLWp7lFNQN1BP2TEhFhud
+FIEJX79jLzTHoExHTKgOSbFDNMdJk4FXHddfwOQFgCTBtWCLADt5RCHKIKSfIni
+IgUnA24lR5EPKUlFhqbdtEXxHryqEce9oIfTOmBnOBAQXLf6UGp9Y8JzxGWaNMd
Fm8liFfOk6ZpMH6KeumjuP4S0bD6w6E+3s5qB6jMVBgqYbji1bFwXK+cYzKa5iy5
FXOo+QN5gusjOMSLxPWepD+U72VgOxn8pW0cVt57N1k9fQej2faFy9HavCurZD+c
dv5oA/uIqVVnhNxbKeo+jvOCrmxP0YWyAIhFrnIdrnRMq1cm96+BAF6ugf3fdADC
VR+ofp0TsHFsgKIYNU/7F/euJRgunT3PfMuXzFDWcSVgyvV6HOd92MHu9flSKPQZ
v8AtQK942aMpHTxzCAt0KMQA/pWb4siP4urCv0Z4rNjBMjPaUAJC9w+qHsZ9ke4B
iaKn81JWJATXK/2OuC0NoqsBA/BNt+aOVGwsGLRe/7FLwvNrphadiAG3RvE4kMfd
0NiDshvNG7c4i9yYvVgRITL8uvqyNpTVOg9wsq2K602vW0IZQE394/P0oearSwma
rw523DWSow0RRI0CfwoVw2yhXPrFJUIVZhFwQZvTwywK5RLEW+gSWVFHUS5bUbir
EnGhe76SaFABhzHH502gNeDWGIognz7+I8lPiyKgu08t4C8OWPYUGOZC4WrSVLRt
UMAAAPpa98RsZz8OLKlCIjyeA5JZnp388dPxlXAGzrtEzubqubRMe/+x0PPdx7OW
6pFuU/F70Mg7fFjWNtHRodOn2mWhrXHzD/FupNslK41pxf6sZJafyALatm6/EIDv
wTr/0VXhHaksIxHNM78PVMijruSzRjdJrrULfJmwAngTz8GNNkqvsvsgk4ZcPY/y
hHn3Uxtv1Ks5lrKFehoC/Os2Aj/1uMDdFrmxKWBFAtHMpXcH05kOrnGK5reIRaMs
lX/d05p9KAN+VkoS3g4aQZHfdxoLJwCArYT3pu/Zoy8wOLY0N0SP/F0pCZ+RhTd8
N3RYProWtqahlL1+y+1e7neeE07ORWzAjGHMRKOjTpfNoUi/boZ1gSbXSOkXq7Sl
CfbnE3acWYsqYvxbho/pESFOgjXA/9j3nz05jP1vXJ6/+IItc53Y+iRuHzaejUeX
DpvUwnCVFrbcIS7yS3i230r/HFwrRjCcXTv8XLLGMxCceo3s4koNoeOqGbTjcLha
IoqdBFIiDmFP9/BeMPNhoNOy8cBB7CwMNhEsizu1vfb1DT+LOQ88z8NwCCjJstYW
sT9ED2IPMoafNdgYwZfk9+M493VaCQGXeZ10uUhnzNI4zu6h5NcIo85Wh0YNsfh1
UePKHPF+OSnRvIikxA8suFkw3pNWDZ8Xq/x7nx4TxbEkEAPwMsbAZa4vZHEdXVOn
mO/qumeOQT8YaUr/cS/5Ii8XETz6/UHWnqV7WjWpcUrUFYvlnxyHFPWwf+gfXCgn
z2Jq+GWglNxWBeBly3fFUrTtrSj7ipfbvm8OY4cL64o3DqfAitv3KSXqveE1xZTQ
Cu+pDRzzxk1CU4MahQJiOUi0PGvW3Crzt2v/KDGQEtel8nzQaol4ZChs3zXFZJ1O
kKPJOVagzz/8K/NZUuc7u3sVhtypGhk1uLMoO1VtsjpSPb3NS+RtkaFIufQYEsAB
KCYUZZrkUOaEktW2HFpLnjrQsUHQ1wJjPsq3aXEv1rvgW2hNZRq7CmJ0ni1UMMYQ
N+JlLNM+CLtQhQKHWDOsTzJFW1lyawsV+H6EakJWVQcrLgvk2RPHGAcPUlDMvjOO
LsEhKc8lYlKTpiVXeA/fC6pzLQLsf86NiOhckyXh0F2sWdWeVdniUxc2dcDziMEr
YKiha2nCJ/h1XH1T1DmJeVD1aQYHRopWhBXOaMGf3Z8f5xclUO5LnDVm+YEoOzyQ
G58GEpbJtZH2bV5OcZ/TFGasowRc21oZSecHBh4UMCPSnOYGFB7YQKiTcbMhbqZm
VfSc56f+H2ATL0qG6/1xScImqDB9inMVuRKCNWwuwauur5xxT0qxU9R4/IVsCD5U
Wsco3qpjldxyEy6VueKVF4YSxQpMivC91GwS9IKY/1jtDM0kyRWP5zUxeU0yJFUB
MxHgnVq0y+4d6m+wLGdM4ymZn2BiNSjgeGEM3hvHC1+WP1t8jjdGlQE0UosH6Fpi
iEpRPGdb7amgYbet+6VnMlongS1r01UmB4EXyHyZogdmGHRPSqhxedn32JtbnVfx
T16VvTX9bKlATzYQTiTKKUGB2IitW9sW7ZqIKPBP9fdyNU2hyF4fliULtTxEaRF8
G/JI76kM9YV1IJ86abLLMhGq4zzg0X1WyA2G3sxVSIkX4/IKEguqL82scj9fEt/k
Sn/6DA6AFi4Rz0DfXzlxEwz4bkbvYH9UJD4UPaAVV4S6Sfp+ZRrPcx28Y1l+Zewd
nKMFuspg2SKML91UsGJoLG+NdmoFCPS4lUrZbi4Ex2Qn4ij137P0WYvTZ8i6IBGL
kgcGp+7LfTKLi+5bv+QSNkMk1nG2R202vWKC+U329t38VUrVp8DKdelhEcj2+VfM
K4yopeqf/k+rRCqNZuCRac6rjzS3wbuFAxg81rJDqTCF6/O/aUleTkXA1Fbq/e3H
gKUgxzHMIIYHAgJSwhC421oVVwGUX1oZpjWuJlwPTh829SnqR6jLJWJ+zQGKWOV9
qKnBAIR5NzFdjc9vxLPWlkLI1v3QUXXm8lfoA+0lAuMhVB+XmrggoIkzR0mStp4H
5ry8gMQJpvagxjknE9jctmN6SD6+FZD2x0BjOKRtIgwjsygfRe8HMAjAC8Jw2P43
1NsNF1272rVCW3NjRTyLfM2t5xY+nYUMIybgSUfme6uIGSeQlBW0lXC3Yma+s7ni
xfv4mViH6iY8qP4AuV1p1Sljun8e9hKQFaXz23mf/k/oTw1SKGv8A6/etzEGoKhO
IWi5Taiwnf4tGOu/EhOnS/a2f6ZJnoVJG6+NzBflZOFjAiz6zA4Hy7hEF8JQJ1K1
psP9NUSXOElsrBtsGGvqJ5ImCmB8zbN8ZtLlAiXpMEP0VpnedDLa+7YgEi4/UIm5
Aq1B5CleMESwSAkCxSg701eVpKnVmnsGwBsNI9TBLpWRYyPuQlxamf+sFkjVVI3D
VViObZo8W0fR4CvTEXRg1i8Y2j0PU8QQhrwM0aMBWzVW4t4XVLX1ljKIoGXKxdRe
Hgg8+nxHNhn2PDcmiepFmKba5GRW8gj8RDNcC4jg6sdNDai9DxOzcyicvTWVGv3q
SwGdngFQWrEp7D6bi72qwya2mXdQO+n1d8PChBOps1Ueq/VPHv2wcnX1+jiQnMOo
oSOKEtWruJ3sl9G0PZiT8k4dVJG9bIasIjweMAk2Faj1V4hWGjGhPo4ipUEA8/Cu
rRsLW+UeVGTTqJrEDhkv1/0uhANC5Zq7MX+RODyh+3CYKyPLsYQxjVq1L6kTj4tZ
1XDNrKsRrEkABMezsqoRtYpPeTA1SFLN28qiy1P/7Yq45Ti9CUJfQd57Jk0b928Q
NgFY1U6uVTbtmi3jmMx/0a4hOPE+RzaHizWdDmBCsbFrd1V6gEMpAhIOjyPtTP9w
To4lLJ8eBAShiN6tw2qERRtXMYOVimJfggmWStAQMpVZ1132XdKUdWKTEA/6Ml1t
MqYTfBdRPUXQIzL9GSx2W/WSh4J4YfDU9zNq27CdPzhn8aWzRh4IoTgwN2nXfTJc
X/qAfp+AbgwVORTwPCFX5f92JcXiS4udr5k43cXNlDKeO1B6c4/j4/mHQrt7auyW
naqVZfvAujYwsaXw0axX/p+5KX8MiGbmJFOLBQrV5T67o5mI8Vt7bISa9EoOI+g/
u/yTjuJO9+Xg44h9JDjXmRc7yDhmP0IlnQ8zZrdrguojtf/n99Fd+nPDTK+woOT1
ZiZFNvHUS+j3SC0hMjv4E4wiii0Pspzxj4gCfhzR+W4odnGNReQnhVYna/EM4vEU
35bi3YqrEcZnYNoOe1coZ+phV5u9tY72eODKJbAsDwMxZCPFw3BJnbjo/3UgTcHU
mEyUHiDqRLTqj2RDCkz6xg56dFwejFGCmoxG9mFvvPS35JFYXMQ6Fa65atJPD7Ny
+ShsK8SDr69dWtz0S/BGWqHFOMyV2BjELQfRoVXTgOLtCjvUy2PY1yxeOviPZY/q
er9/QOZ8YR6FWbRhktuUAlcK4LAcLrH4puel1VyIW/C+tXTjKfgjv6k4a/OratLW
ay4sS1Np0Rw+/QJzwmscNggBDWRdDzKJxYnOQCgrcmBj2B2XP9v5z/KHCjzve6Vt
1hpQ4Agp2Hz6T+FevaZCzhCDJA5yMSAqo5HqolWfzFEaY5wFjBKN5JVOW+1cq338
m9aA8o37Z/UiueQ635zcNQ6uaJWWUgnlnEInTIp+0Z4m1Qk+B5bnlcTTDg30+9Dp
dpxX3Wrj21mVxsRielCNh+avlkThyMLVdBSU3phQ3Bc6hM05MPp/49J3IFIB1Iqt
u5GBb74SuwPr6NhoRUm5fQUiOfIN6+ySTPA+Ac+k9zGJdHfVvNbGBYYqqWZfcgZ9
0HuLke5LVZONnxHyAtJdvDCllG59fykD2MFPt2JycO7vH2NhvBmY1IMDwHkjJiaP
UyTKackJdWtZox1ut3EFxhouLSIrXTlEm0s6O6TPpWOawneoMrMSEwWb7bR/LvXR
J+lBd+yUIILt+4Ex+I8jNMLwWpzs+IBVDrzZVDzXoGukxnv+r2LFNq496Q/KCPPE
dk3wiSD1DXfAC8EXEkJIujQtJRFbGHjZ9Si+AAE20/CJ9yKLBnLZRRfusyUPLS7p
7QewOXrlgKrKoUNUNREORiBsKFFMA4QwbLL8fD7WV7MIn7ibjB6lF2qg/B0uMe8v
0APVZJY5BRAdlM3BpJiNd9lv8x03L44gA46r1I3L7P0Trh/sQDJDNM4tai6/Yd0A
B5v57npps7tDxvAfO2SULq/UYr2brUnkLY+AxfB0kjQze3LIqDoiiWFuFzAcg66o
mHUcNwXnRV72iFn45SxD9X6TC7D5kiMQ1YzJwkXVr0ga2/WmF/DCEVIxp2dnDyOO
wV1q1+yINUMKd6LwuIQb58cVztStBcfcIsBy6dGVamLAdFHVA7CafHxJZzFyvZ3Y
jMu7bPJiIouuZhrizaU9i71LxLIBWTP63Dp3dk4t9dkWbOqCfKo/Z9+EF/qGM+az
u/7IpMI91fR3OOvlso83KT29KoaQUidzhFh5xmmsCNE4rbMa2f6qTBuFCpGz12W3
8QnV8EjpAuJAaXJxFVGINBje/2Xt/hPfuHUhEmMSy3DXtJ0N4F+8rI88F6NfCYAF
WFPY7xBx3z9sueWzTS8Erh7JfcIXzt+o33HPvsECg473QLE9H3OLIXeA4aO5oJDW
kDROv6+IjDXi5SrNsXcqy4ZS9wdPBZKapYqHFmZosx/QFQRcwGB1GkUxS4xuTDuN
YScoBgQxsqcZq6fbyG0MxRnAc71myta+/K3hxBXrmK9j9cp1QKPe16+oCER61Lne
jPhqhJtKgVQVzeWs5MJaJLrwWK8YVEPJArPMC3vIwwg21xCuQlZAOI0nquB9NWMr
kspwIitSrFEyjU0NqSOFUl1th4CavTmZ2QgRErngETBQvHDz5W+n8Tw9h5CnQw+7
+HR0RsVa4R3vDx3+xDt7xj0U1ODpCk2bVjOO0G8Mrrlemb9TpRQF1W2IMcnh93Ue
fM/v72vfbferyg1aP3SS+xyG4lVHUAybS85bviaywN2LR91XG4nZSdvyWZ8AfPF4
7DmbU5lpHCdWiNyhZJdMeMZYeg9ZgGDIlC+8/MtdJpSHQvd6bsP0ByMx8mp2JLI+
68qCKTlroThkNuhlBECvneuFilYuaf/3491UiMUdCgIu2eDRqWursbeuFlt0hZjz
67jpg5PeTPQeh7lQ5E+kRTSlFvkGhUH6k1xOK06btyPgBlAMlsjPF3j0+HuHqQ/i
rv3E5DSdoo0IrwhaN7UcxX+odQnTTSdMmO9kgE1dokPU8aFTt13W9N8VnGWIDnHE
pM0gppuFt+Wl704PxMhhMrLKOVE9/TnCpmYoSn5aLMXDHdvAHA+w6UlKKvu+BuxA
JRkp890XWrjVld0dKva32QaXGbaXKzCkedY0Q5KGkIfkBwWuvkjFBjhsiXN7UtS0
hZbnPzC4o7bHJHqPH9LpLgV3A4+ToaY/pq5U3sC4O8CppjhiKae90BO2UYcoXNrC
VUdc2l7NdZftX+n2rdIBZeTf88L0B3s7d40hMV0pdr+BuLggvCVbZFugBKTCq7no
+6cpR7o/dF5UgVpKIn+C6f2GBjab1k4brnaBUNnvgba5oT+GLKunXRUep6ipFxHq
ZZcadz9PH/N00ZvHDBA1yKe1iHD04pEQfOBZmRmS2HpEflh+cVDTZpaiKAoesRpi
xooimtUJmpukkN1FZm1+1VgPiVj+LXmabUfEoMd+uZv6xYNpFAu0GFFBvBqLOFgK
eBYBell5/W4Ukq95p4cVFxmaTWwlJfbOP9WT6cgxIItRA7AI8RPabzSFijgPkhUZ
cjM5gaeMek70I66KFuQGYrqAkeab39YQ2CCuqOxqWCENuIOMr52AkvFBhe0aWTAv
3gIcYVNAVrBCOCFKf8Z3jvpwoKEzyxBpYW1vAQFHka8nM+h8/lNutLs8TshGp1Sq
q/ft9Oum3PHqIVGBqQZP9I8N+oJLXKxtqM/+ZOqOyZ+df9YNTFwwEta1ksGWI8Dm
cznCIjyQp+xh9ab785meiwi4MH0CINZTvLp6VTjFc1AWkdIKQd3kz72Xxqw3XPLj
b8nO+90uRSl08owShPHPjJ6zuePRDo7uPXIKwQI2EJ1LeVPsVF7zJLWTNeAN1PHS
u44unfVUG2tE8sHd/HimYwEqDF6v0KaE/8Ur5QmObVIzKswdfPgE6dps1Lr7p3yW
XZN6KRfHb4Qf07Ux9J+Rp15w+jx1Ex8xAw85BXDrjMSX5hhGcLpKKVfySs6Y0eGL
6uOVZGdMl1Wwhu9WX7HH4mnlWpUQAuMFbsBo3AmXo9NbqGqTqZvGWAkeTh6KLW8K
RqIHj1Txcf2siQHB9ijp0reuNmpAW+QCIU5Ej0oVAcxcGvP/jTiXiTl+7cEjkDp6
MOW2EaCacxF63Y7L2dVlvIcvizepdBQXY5DNwa8t/k2hpqYOHKpOeLZgVGJdWYmn
S/4k0jcoxgZar2IXwm9YIDqQYvze5CGcW1RXnTPLpmS4IHiRXWj021DM3AHT/Z2y
XNshDm6jw2BD6zfZuAp55hBVfdvn6F1K5kJ4J5i99OcFHb0bPY7fVrm6IK67g3a1
9xFIdzWuSAPtHYhyus7GJ3fulK17VX0+6hhLU8xBZSFfFyPbd+00evZQqMyRTjZz
EypxbWzaIlsEiGgSKZpcg+x9ardhlqpLxqwif8Cq08FkOm992thqRf1BjGkKIHp+
3QwAAw2N9zWwELWY27CjgZBNupygckyLTl3sWnKgJgBlcZXo1uza9DjxFWZTO/yM
uq5FGPigQ8aUC+MA4vi+eKko/Pf0VNifiZX8iw8Rd+rYxds0GzbRmcq88GbXCAEI
NgTQxxFcL1RspXKYYhpQ8fwQLDBgR1P+8EfDSQ5qRXBFwvzg10vQyTq6HdKfc+JA
20GkDCPpLYuMYD+AV2Bg4TVTPApnp9oYxUpMj6cOxt2FmW1M4VcJfU1IlKL+wZJw
wpQKzYE8FhPsLj7lcuHOqeGR43tHP4kN18oytgln8f9aTe5Xt4J8ZBFRUuo7ipQq
4vWgyGdNjhF+RLv4kv0OeUizsU89LFQebHmurLNq36msE0CdakO8I3vgA/Th5psE
8O4mWd1KjQ4QpTjIWdPGZLAJ/6VkwLSsM1Pl6iA7rYeryrV1/Xw4xLg/9ByfM1V7
aj8tJqsdHHpVP++Yx8cqiRbx61uiaIaRguLKc6t1qwdxQo2oHE9yOLzT22ktSgkL
yJFOvlmUDKywiHSP5xkJX1hSI4Zgl8uRp5bV8zynDxOnSfPlUCkVGV3yfUSreLS1
YxmCqYxZxrwd9YO23JGlr2goEa0cXcnzvrf4PnBztEYNVsM8v+ttrhjTmrvgQzxl
cnTK6d0XMEFFjYuJiH22w2T/wUDWBs351+4A34C+jNGLUlQrfT04GxNTigBREZSP
PWZYW3FAYBZvpvrTN+oBeqQyKtD+F7bSLx1RZZ6llkXQvBfPdBngD2vlEMY59HIY
xL9tOuTfa+bMimZoeIwGH8pmW6tuP5faP93Tw5FAWQg9Y+UBtr2x2Rp48xP3oihQ
MSX3RbKsbLFYO/OXHnUGO24ciSF5eyRiYyeeqHiVuycfwZ6Vzy5kpi5NmGJNFF60
X4tGz5LhUYZXhF3ac3ZKxBfL/RGE1jPBgSoM/zfiaX7zs//lIbv3qWeRyd+OD1nn
Lpyym/o+sD1fNpal3ltjSVhOsthiAiAjVymhg11vwO6TZ7FDVmiwyi1gBCqgnz7F
//aZkC2RU6JDgDKDq9xvtotWzPt3R7o3YVIoNFF+LScDMbDuUu8BCx5bCXJFPbXR
bnZ+KCz3Nq4PuvKlYm8cZsQTXiPf+62nGWmbYfazPyrL+97fTJE6lj9Om1C7MNAQ
nglTZIbeN0lUgwM4YtHMMOl73+gnSuy8yruQ4MnuvqhtMg+9MritzTFkav+j7mF7
eLALHqOxp73DSBz3fHaMl4PF/s2+DU7LgCi14j6WEpOygtTpz9+lzi/YQWIE9Hrv
C59s1NrVu72Y0VGKfyUeLyxcR6POG0ZevkENInGnQEouajR+cXRWB5Yr+9mKto9B
1H/lISWpUaCsS+18Qw4ibS1iNwg2xWLE3VOfoLbFhX7B3XQiDPGo+U+7rC4Hn9sp
h4fVOnDVOWxa71h35jjl/ClX3RWwe/BKRwl3v0ffSVKrBT4FfW48be88W3hCADKA
4mQsYNAvsHXvwPgKt5HWhyIajO0cypuC2eST3plfWaXw3ZqB+A5kLORvUChbuqIY
0Ulu3mRYEIcc7vh33VeJ2yvPQM59a7wqrfGU1hR7GGIyr48Sil2a5oGpeVWBIXwx
cdhZDWl1ugF7HWLFDOya53qd3B2aiC0ycsclReMHLaJGUWiZYkr70nsXHlqQUjhi
VovoM2mtKSiVVgdffUknBzDTqVgykuBw0Fv4f4wXGtlYkmIYwixzldemGLZfLGsW
6qCWSYRH26RtQ89umzTDI+mJb4q3G3WnOH4ZbpLPNGVmgthbd7lq/lxBtDoEqfmW
Rh4yXcH1ifld7Gp4o3l782k5tuGqGH53DA32qFi1ryQCdJjIIKFwpaA9piKdyi1V
p7eQfQZMGauIauFqeeIGOrD4ti+D7QIhiQ6iBuBNC4qD9tGuvOLpa39h2VdxmbfN
sZ/V6c4jYEI5Ifycc6q14hPgcnKGk46aqtczEyzTpnaixoD61GDt4Bj2KI0bK2AX
5TdAN+OK6lwfovACSvbA5axaqUvSoEkgC2EMmssxsKExS+Un/UkAdN2KDspjp7g5
cD+R3+SPJh+rleRD5zl7GVR5/QwNR9yWS3+XhntWrR/Qdn5YXqCmnxulbyQSQwcK
uI3VzlNfEevy68igxOjrF4J7R9TlqQ/UiMzL+vQWtqa3N1oJXdMBNMOi112HjDww
Q+ap9aSqO/ZEyLrmoFa3NxIdWBOL0xu71s3uX1H6pLSXp3bgm7RwQbJ2mPTfpJqU
sznQ24c0lP8z+n7vFcLq8hB4EMH5psN0pCEjM3H/z7cSGBJSVxdbENK3NK3+sz2r
rCj/SBZsCHGAQo9scrZSW2UZ1Eiq5xQKK/FXmteh9ViNozwIa8Uo6i/k+HwQHKS4
`protect END_PROTECTED
