`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GVySyGa6FnFstlMSe0A4c5s9PVmAD/W4/emmoC/BpabQ40JqIK0XQAgoIImC38ex
7tJI9gcl52IjCfuDNduAcOhzoq34uVW8p3vqTmJQQ+hfqtAxxvr+i4pVAqn1WNaf
ywrb4mOJuf5v1FYklJMJpBl3vrEh+aqncVKI9G88O5+mrYWuOf4W0v6LhP9CmUjc
0orlMGH7+E1iG+MKm7Llj+Hgp6B37EdZJGQRWoNrcESML3EoE9R/++ShDFBZdf3D
qg3cXASC5oElWJZbRJ+f9518TnI5RqrpOfNuDw0dDgVPV042GkY6nDm7qKKnFruF
PkOzImelXSKxgiiIGdYIuTbK9cxCFvKhDYL6aDTsrLgSnCKVcC7RCkknwueEi9mf
KNe7tIh8MvzXE/pnE/MmfK8JJJH6KQkRIy+N0Wu8w1YpXWt1oZETLadXco0BoHCG
sQtGAO0131b6BGDBLvp2k0slvy14MV8aqXE7uu83S9LckF0PLYEEtemA3760hP10
ymgRovpo8Q5BHPy3AAiXru55uF9uRfn+I6DDNXXwW7XriTdE5GJ5JNQxrHQAgXVr
QlA4OxVe6lnhrsNDMqE52zUn/x3w9xAEM5vPOwiC+ySbMrKkBe4vdX3mU/6pRinq
F0nM59fZjH92o6swBHNSVrPS6tTU2mGXf38B/0coY9lGLliU0rEZB9vU5I46a84q
2JeS5h8W/+d/R+Ngie8T2NUXr7O/8iI8N2VZF4scYN55aKoKDqCwRN9tmVWkNAHH
FBd7WgNdb/YTbuWT67xsiCfknUsg0dbLe/JrhuUA8TvpkUZgzDLmINbUx7FWOt8h
Dti01VAjkR8qkQzwoRCznBXJ36cx+gAVgONpUl8HPImpIMRswbp1o9lEyH637BLp
/ZuraRQY2S2vj2RcmGJodPmEht6YZKmumoxRq1aZ027gHPJTIHCQk7lGzHQ2rXWt
xlJlGNEU02WGLRZK9T9Q57j1ZSe9f2K1JZJJt0EeCRk4NxTOPja1LL4lU0yS9ahv
eWxQJOpn/Q0U/TD3P2wghnvX/T6F7SVli7SkAKouU+YoZbPzP+2q9M8LwsqNkuEi
DXYiMa9DfNKgfTmUgRWkxm4hl5n/CqiPDIFbYdWvKz7+3GQI+KXzFPF715nQNwww
k8gkfzvdq624VINpX0EC86aKtw9fwy9jv9u/yrF87EAShNJ5AlROY2/NGKIRmEfV
3LdkvcJlxzMufA9vEFDTTHUffBEbS/hxqn1d2itIf81RLoZatI+GIbz2rlY+g1/n
LbZE+Cuhy4hbiKivIdh83IKwWYx9IUMxjlngp7TeIPm+G3N/KfhySoHzMPj3CsPo
OvEnNqxTA4REQE5eQ56YpgfcHMnzxPN+xaaxokbWZfHZurEiGGQnL5frPbcJ6XaF
HZykQ3iCn5uN3cU7Miaj8Q==
`protect END_PROTECTED
