`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FwFuoOTDGcLBXoxI4sla9WMKHmSiTn6yKsMWOE66oefqkpitLLH1TKk9xXb6oHHF
fiw4tRe1wdXurIqOf4kYQbf1dTt6/jmVIituqVBi+pHkOu4ItVzLt21BOnCBdVpS
fuEp0wRB1lAsmQhT5uj5NYbIL3OUmqILXi4b+3qfXGBMoEThX/9pDQ6VfTX7PNHE
FDb369rNQZtY+8rf5q9rLKxqVY+xr+HALK6eo/zeiWNvK3I155hZq3oZa6ygje7V
MKXk9uV97ZeVOsGxt08Rmw/5reA+I8a1vzp/z70hflRFhgGiUsks4knBDkRS7sFq
7NBa3PPOEinhPwKrE2ikr2U2isEAEr65O5zsLt2S9646ReLCFCVxt3imi9/kgIZC
7GaZAWSXlExnW+VSTA7dksTPsTT3bq94cZsZoBKqD/7paln+g9wfaipOMG5iPT+R
OmZ1tZaOXjUlyTiAOxLvxneZ/FLTo7QTjyygfyJNwecWSLQePInnlrgCpdopOJXg
3KWfD+A300TwgSlttIrN14Jp5loRm9n52G/eWHesPzhrsoRcORG10/cqIp0tStAt
gygphJTB7A6aycDw9wkIco4h96p8c0T2RGS4RAXr7wsyzDm1ecZLLuY0GbYzUvPX
vs3xl2A9zV65NtHMLcfWFmap8JegM+eSKUKxQ/AvUXR86/AO30eOluqqyIEFwiqh
5TLj259KtaMx5HZjRXIoGowYLu5/dzitpPrHc1MwN9wpl6z6PrLp+OWUTRO/Oj+s
/RSGagwlcoxS3iu1hRSYW/EGcSVRReYarUQiS36JyBahWQNVQM/p5Mf/826zCDBO
zzrstMRKZuspGejT7b8krPO1kIMfbqVFY5Era9qOd3yyyTV8u46al/G1ioZ4lPu0
hgOa5MqHm0qfH2D9Fvq/cplDFrfzPTiuntEBbbZaFAQ39ZnTSrD/USF1filKWdon
uvXmcF0JgJXq1YA+H/zvSnGiNcnJnrVGPOpRo1lwPVKKZapdgLe3ytwHJNpljsBj
fhmNA3kap52f/NRa/rff7CbSboTAh95w9/ZqB9gCLkGzsIjpNYWUOXKat/3OCjIc
pvXxx6cGSFrxY/S2X/JxM3lLxeZ3EdTeBk4N3Z1/gZ/Mqowbd8MWtw8jHeIi/6EA
dfI9+BjfC+e9IUZVe9tiSJEFzN+A2u2utSdd1jlLVrPNG49uU/eQ96Nk6svMhOyg
Nzmd5jAbGMtFsVlhsKWcXumhc0adjK5aL2S47fWeleNk/WgbcivyOHllNA4SiH8S
zv1k2LdKW27wk720zCFNK8Z5o+daD8rcAWFLRE30ynlZkoRqyCIgEydk7Jf8ZkCu
CMBX5t1MLy86BYJPqHm4MoFFKp8tiwbGTkkF26jpJap71SZokdvfY+k06i8NKrbn
ZZd8p/rp5ar+CY+MAxRD9uYWXaOzcEF5wnygXgG38GAw2YrqveNHIW+OcAeJwo/r
DHBCDYW+jvpMMkY8kZIH447WsQVZbIcr/PcNPBLvPHd4XB6KT8BuZgqUElbVWet9
8zhmlQE3skrcEVE+bcOZ6Kg5WLl1XSaHK1y0br/fvd29szK0VG8q0AYeITkl/NYl
qJ+3t4amJ1JO2pM3c7Uf5+4IEqe7NyjR+SKTDwMuiOFitgzJFCTaWRYLeOL/q0mq
zTpGCaT9qM3jtkraJyWDRosx/5cSkx5wMb0ZAw/zAj/envi1JGvNrCVQg85FQQ/B
K3f10dgWRxLnx4+8kgkJaFpUrH8LGH3y2h/cp4Xic3rF81f58zUeOnjNUHLrjACz
y129YRSHvzSwmCNSQqbYjYpBKIVoCdWeMGEY8UcOiQY4SfNTA6JrNbRktUdPK9Pw
BsYueXuOfKxBoCkHT3VWlmfv93CtznY+2XeNdoPvbT659CphSI+bZNMFU219J1WJ
j1KBuUg5QV3t9TwLSIY2p0THhvIloz9E2D4Ygv04HxIxcb8kuihXGy0cymO5MvSz
KQ46apg5Cj7fyx1iUEK6QZQvcNCVqYc8sIx+uOL1bw9qJgwtWJ2+CqcIlarn5Tec
jwGOAUgPUVJnFiqAfQYjN4PwaL2o1VrmBKV6fxitakjY6UW3TR3VAAA0+cU+QJR2
eF3+TvIsNMHBfF19ZEbSbVJzqxSalMjPRo9ZG0t5S6oCNZF2OsbmE9p8yjFe5cGd
ip9rNWPfIHJtKqzAH9Rjy9yeXZyYvCKwWLToY9gboEm1X/2Y3k4mp3f5WfgYYXxg
lmdlIlgmZniI/XE7nnRNhuqR6B8dffTuucmpXUcaVG6ZZHS1eM1xVupk1xis+2pQ
PdJJS31O+XmUCvmp5AB/H+14ARuKW6FF9KqwugRkYpznyvZoUdDZWdJVPRqPQx1W
nZ9N/kWi7KKUxVXtSImMTlOPAS7/XNMi3Dd4OEtuN+Ng0bT+tBQM3iKF4EVV9B7P
tEQF/NhJiZuY/PdmXcMz5w==
`protect END_PROTECTED
