`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JTQ6J+3VZjshLtcR/DwPAkiz8Dnjjk8z7vtkC30ByrEO/gjER6EWcnMybbnKBoP+
Sx+H6TWwTJlpqZgTFvYpRrVgQE4fFA4+dfvWZ8P22ndXJb0SlZs8fCORmYJUso/d
Mj/CaPB3Ggraywh9OOXz3GcqvUGG2RSsACmhi12L4j4VQmQsg/QYhf/94OYc1Bxg
2UO+cmfGj7CijchysSRrec+xADXI2pBMWbOJdJK7lSAAI2MxNj5bOnPIwf2ui2+6
PQ+9EuGp1bFcWoWWFBlpiOhWAlIxiskm9LEXRwVW1f9CxOWsTqDaLqxWriU95vFp
yHf8F2I4cB6YdDyKnfJd4wwiPmstg0Ubr/Wfm/m0twi7y+AqbpGH+7JgaYOnBlfr
iF9I1iIkR0c5laV6NFKyfw3ax/6k8/iKaqUHHA3GPaQMcC4r4dA7Uoj1fQGnwMh6
sFv9hH/UXpS/GDHkzlYw2QqqojsuyRAXoHtM3vd+doU=
`protect END_PROTECTED
