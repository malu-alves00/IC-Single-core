`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8MuX8F+2IJ+Rv4Un3GZjhOpp7eE0+KnTbGKnEGiCbwyspI1pWYP4JJ4CLMyL/n3Y
NauN88XQDrsqi6lZ4uXZlAWbDL4Xh2vOgHb2QkNxcWoNRDEypaVNx/3QCOheAWJE
YCzfnaoi35F6QWsjqMpF9XaOBHPNG+ipG1oRb/jsSk3VQCCjzTVQvG5g/zcBJpSr
PAcanaHpIe42zSFWItUn4C1FtQ3sMgDCZMIyAeTZRj56WRb5FI8RozQbRqujyGqg
AL5rKBFrpu/sFaK4roxcLrHf9emfEs7hk6xPL26v+s2809HGef9Y+G5DSU00uPvT
CZGBUnUjYLT1uHHSqHIR3QqHcSObMjiWlSJK6zjsxpnuOKqPErKua8V5i8O2SE+X
m3s91lqeabwp5TKQVFfPIlu0ONmCvVQ5KmfIayEkeUwbtYJ+Yuowc4Acpp2rBch5
1CRv/+PW7Box/Fa/txNsNZ6bPTmDbJlyjRt8WXlV2qUbokm1UdkplsQ3I4wOQAoZ
iE0OpwrIh+8sGX+V4S75WvF6auOaKJt8gXykzVIeL4TVeo6m8cqDb/AwRLx3KjXa
N0Ns9DBMIohvvkjqjNzAF8Q/Yxk33UEpm0PdIrBJf6rRL/Ptn/xMXOYNl82ATEcS
3duhe15ltOnRuBFVR4WQ0XXADv9U56NMpZgdv0pvf7FTfR614AFSKLykewK7PKiJ
xXXPVJ7x3F+JhE4rxTH2wiQkBi+EJ5FIfMtSyF0lAsnYHE3mn3caQDD7Vvb5OHDX
kfO+UfhYVP3AnnPmiTmthOwozWuyeWPlbiuNoZg7go1fBg95GkOyDO18CbWPL9sH
0AN5Ajmg+AmNKQvAww9a0jzqtxHTsgNEYyd3/HUY4KYxVjpn1Jj1TdgmTyd9ap62
5TfAiy0FwlFOgw0HY+bxO9rgPi1faOXGy8ZX17+CpQZMvZeJt/UqX0lLIJP/kZGM
4o/WHQAH4FEYpksnOkGUIF7qpgwjXnubIZIBqoKTuqOYTJPK2hRkNlonALCuqa0/
S513SuTrXGfQjhPWxUEsIoWduKbzwCpyZLWK6KT6GSLFWRrZF/HvDFT78FCCPbf+
Ykley1/9EDymx5D2GHPXvd0p1yRbLkxZxXvu0E4gId+yUlWgE/MPQxHowc34LBf3
ChzghaQbqgDeDtL9ZDxfoOFdSCWVXweyq4SNA4j9CPg9ICEa+8Bdx8rsBtsjL3Ax
VQ0I3kAUCZkQiWpTN350ai4wMNqNKHrcblPZvQ8nzyiVDOdeDZ3gdOeewbboHDmY
BSwm8Zhd4tRj7Eu1qef4hi6LciIcsrHnVDDgZTNzxg8U0df/pASKPMeh++r4wtfE
aGlg4VVlWOOYtrdDhXLykI+x7Y/Fdngv4ZmPbqLmis3RUu9oUPxPUuKjvIwhzHq8
kMaM0mwMFOyuTbk45HThnvtaSsEm6asIOhItvRmIaEnr8ECwJIoaDrlK+t/tQdC9
UbkmwgSCkN7oLQ55jj7noIdZeqWpAcDaCNnGfQ8gsQCS7zHbBzpttndTIw8KbPKg
B7Xw8L/51wlIRkU+pWROyWJFZNQ9nzFCk+w3Di5e60HK9iQ7smfBkqm/2lQfkeRA
lQWXWxfLfk+s8Z8++mki3XvMHBlY4GWeLdraq1oldnHFJYY3clgtjf9hStMYaO7q
YDMGeHp5uSsNtDqVkLc7snamj865Mlw/04OdOXtg0Rv/as8672Goag50dtcT5sEK
tLSHcA6W02MtkshSUVywp/eV5tNQN8KAiRjOTct8vrzoLSMCqs7Hldwwsq9SDyq3
b5KKAPG4Z41ZmjRY1gSk6g==
`protect END_PROTECTED
