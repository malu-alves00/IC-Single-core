`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oGY37wKGUVoUDwPpD8wQtmve0/7SKrGMgATOxgP0pJiBzsiN6XB6jWbUzurUdRBS
ohC1GYGv5WQ5ptHzOmrVosc5rBXfKb5/kpHURhEJ8v9HELNUqjcLGazJK3rHLnVD
tExILvybxb6TIqR4uSNwCoPHFBVSzC1vfvj/tNZuHd68Dqzgy0oqu9wH48XZjlzd
pky8LGtlEjwkW7LkxrmIqxewxr1L1IlGe3qNFkg+75x0+JAqYlVbdGF7AmbRCHIf
/8Zr8YFEQ9iEbcBba5YzArKsBYTKBIIkKGR5hC3tRJvj4rKlGPbYKJQJm4vQkNBp
yCbh4BO4Hi9qsnMvstKRhuhAx1ywVtXKwOQpHRNVNvpguni4lQyqF9RiB1s6DYGT
DyTknfiOrKUL4eJqPEyHxo2nab3wIjWi9oVTVLcHri/Sf+Ypqsk1PSUPUIMbhVKn
WySXkA1DqTzVX7Ugfv8NIHCLO7pCslnYhNO3EPrk6PjPeUImiQki+N6gov7MJROZ
lTb9ilBvp7NRj+sRNglKX6fjpZAE8/Ys+5nwb/we4INBTKH3wB7BiVZHKvH3SgdM
Dcu2HygvECLjCeTe/jPhDktkMQ2a6S065Ynu8HiZeS2oNLRcRyB3h1cqLZjDLuRy
kWDeo73coo5eLTKs9w9QJcdxwo9EpR9Msj4avCqGtdXKMk7a87MzRBR8VdnHjNL/
G/yuSjfQ6JZ/RBzMFAIpPGbvINi+bka6wzwmKc6uO8d/L6/6qkXMLsBAFYEpMJVe
t/QKyPQNwWw0R+vPkdhKeW5+riFT1mWd7rlgXNEYqM9Oy2q37AOAspcC+1K0fzG/
okanwutEpAYMmL+jEXh6OzMyQZ5HasmHolYiDXFbNFuUeFMaJvMN7c9g1pE2Uarj
iMwe2BLmXxPpAPtYk0ICKyGFfmsXSUAq5kQrZMH1bXhYd7nTxnS/lbrzR7iDsQgJ
HMQUOacdW0aQKrv92Uy4s2sjp55tamsnqlguZYVgYfSsjd1fbeQ3/kwITA/zM7Wq
ECX9M0ffIAwKZy17ifvZwvg8Nb56lb7K0Cj8peWYw9Js+qa3jknCGQTxIbbUXJpf
rxt6rp8xkPSer5W6o92MXlNyZgFv/3NbgUQAMGOuMMKm6jexO5YJ1fPhql9hhV+E
Rle3YUZXtq6Tq8c4zde6JLSEuOHdFNotKkegzhgF8EKB0x3/1XsNnBecxSyB5mHW
O8oip6YeabsIn+x6FBt3jncPY3ajNjwZjVVI54PZG3gL+kKADNO1XiSno9xqsp2Q
hdgfELvibVuWwn/mcNZkZ4JAeO9FBTgPBJKszI8MFfboWLf+lmNeA4XoKuIUjqCv
Ysz5rQBng8en0YGQxLh5zbtY351B7ou1z7VFFyvM5nLVrw7OQknlrsoJnENgatGD
QNyTq23Y07wHNd4ijSjwZDGcyEq5rnfxdcR44uuE7xWwOslidakBoSWeqzetrRGT
GWnDsNMMhc6vLWXxrNJoztVvhKvWZxF2uVFB4D67BaIZdfyOIApYTXjUZR12mlml
7s0U3GDe9x8s2nu9eJ8ax2k4hJduDn16v8adti3yFzUocPEdtek3vaRZSKaDcTyK
oL7yKCbam3ytnYcrfW4rcnVntvVaZgK4+Pl74BYSWZ4q3rJVcmYVh/ZVyvN1M/Ra
Jgvp7YJvOIJ94rn89H4l/Mpx5P6W020CmZ3in7JY15kXE/8YbxD1HUSaouz/FCGv
BM09QmZIy3RcUpznQlAvUgavUMIU6T2AzlnphXNLaEGc4uk0cViU6SoV7sIyK+r9
SEu6bqvR8INQPHfVdlw/UJFY9iEK6HBB6zEWt1d9c+DVeVaw+smn+UBJk9RahVAf
HxcCyiApqH0BOpRcBEG+zH+5DSWopHfLYSczFNvZP+YJ6YVmpiVyCH2zWeaHZBLq
pO0yXKxgieCdwx3BDkRIyf6de80DKtqhRnmGUY+HewtfmweFAvZanLB7J+wC+Fvz
v8ON+uXZkuNSYBJ+yBz1x25I1+KlAI0wycwTE6DFDtersjXXQlHiCVUFSQk5zEU0
CxBZUm4XIDGoZso0cIyUgsTqVeT+5JD28Qeqe2KgBNw3klEFOQTsaLahe3Oz+gui
l4r+HRiWe4TS+z7HDCnjnmvR7A1SUBEEjCpr+krWFBIYYrDs/zAiHSAn+DXp2TLY
+btgTMDq8T1mVq1rmp1ibeehdUpvvb3Md2Z0x+gUrbUaM2dyHSAE2o/beNAx0JoP
W4+N82jJ9EsYAXiOE+pkU6bwswA41NA8f8GMgpcMlAedwRoEGxjNAVag399KT8PT
vR9tu7DCziosFOAW6NPyEfR94+3hW4shzpnxB8N2e5gdwwDejrUkebkdFgaR5c8/
SayBbjrIM5070uFFvZUH50gigULrqt7pj5Uq2CV7wBeu6YRO2Ow4mtYKsKHpcS/K
KbLb7bBdWLN1L/bj9dTOeUAvGpzY6MzZ8a7eV/yWoDtia/psQyaFQtd47ld4PcbL
Ad1qqplFhx+r4PGkEU7KupcGiaAR2bdRuy97xONxffJmhjgZyJSS5BhstcSRGSu6
FEP8s1FFik7wCRkjys/U5+J96gmeJKu4/ixoFoC4ZKBQquTGAf1/rgG1cfOCpJW7
vPoybsaPZNhxDEMM+uKis8+jCDoDPhg0+2krmcGxIj7reavHbuKI5YsTYNMI7GSa
tX7lmRHTr7kj3rv876sb5Ksgyf1yhbGItA6DpQXB32nh5T/Itu8zj6NtAc/hWq4i
bVKM87IOdTYK1eCr12mncMRMezFw1Dn0MgL3iZbi0EYJyde6PjKViIjMYbRzRJgE
qduK389GnYt8KjUcxiGLz0pvXR7EIzwNXltJtQanURyRrG/HpKe/Q4PGb2KO408S
BpQ73TpGfupPtYfKcmEKF7w2M2UHAQp0BmZS0gY/KUzoViDOvT++KVVHm6TYCfqp
a77XhtveUXTODn+Om+5T7CKrDEbibP/iUD9lCz0fRPzGPt9psXY96XHGcO4fQD3i
Vnx5DCAYnHdw40OBeRTA9TDZVf3IWRQu0CLGxfvaNBbuePZlusmL2mK9kbGIBW6k
/rS29DGpz3uYPNXID+8Z7HABV2HGyyBd4neqG/24iDAj+NbmJqfmbN3iUrPflVtk
xZSvxYGfHAviGhYl/65LYjwK0xTPs8P6CH2UD9yYb4CFVN1enX6VrKfjfpcH/T7+
rHLME3n0OT2tCMqGymNoDxuhFzrnHjXH4sJbwfBi8NxbGtxsuZf4QYrUMK0DO+7C
BR/5kWU3sOQJz9eJAmXZs+SDLPzkw2fjKq/6t7MJsxaXLzTPnUJ0ZudTGqkOmNdl
tXIJJrk9mvUccyjN9dphH5W/cfKEDGYSTw2Qg4Cs0D9tp7wzL8cLqmGDcmTYSro8
SQns/nRJHJmwqgFXsr6YZsJqSZBY/5mHeuW8QxQM/xEMJBNf1Op4dpQDH3WivSTL
c2CgPW+fFVy0yeEgSMx1lqMqw/n/Jebm0xn4PSg4pKz8NkxiSDQbB95JbGUqEFRB
gQMli3hYD3I2XP1KYOUSAQGTe0drdNDPXhLdONb/pMkCkYwru1PerQOfQ0s+Nexi
tCRWm/rc8fL1RZx9V3Vwq19sCmUW7Boq6UGZO0t4tt+G0kDA/YOtB3iWOKAD9j3p
JRD9+Q/4UG4qrPyKl27C00EbEbnrp1ONE3uQSqqUvrZgqsqe9NycoSdS27U9zET9
r0mD6IuYCw9AbDWtt+5sCrUT5+Pj38nHzQTz/Uej7UPPZ1j3SeO9VP90j/zmTD5z
wYFwrqLuxn8ippEZNIX8z0IWbtaRxHAV6harv/rGXWLtEgCwh99S6WAW4dQLs6Hn
1b7c8Zj/S1IGPbiKGasmd9aEDFyCSU7x+VqR2dixr6V6DvAT79v+JStHrZuPUPu3
dF6GAZcFiKBdxIG4tWSuFxiZWYS616W2T14L1I+m4SCEpydcNjNdaKxGhu635J61
UR6TPq1j6lYu7egN+wHyxxJoVooVZ6p9KlrmtbPJASqkoymfI2ZJFlRMJjboerhY
2YW7jAcU4iPCmfoznDxxIQ==
`protect END_PROTECTED
