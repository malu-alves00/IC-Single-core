`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5HW6yzeHNCQFjqL8NTAz/APe7dlDIXibOfT4RFzSWenInqY52qFKpVpze08rejdZ
cdTVdai+di/e58naiyb5E/wpWzcaVyQJS92tJtuXGnBzB+fdFAqiyuxJ2VLo7WDX
5pfI0b4mloo7EdASGsCWWZV63J7Bb77izIPNcIz5EuA+V+ZZxldOMcjDfPzxmNJQ
RobkQcV7ALVYtG1S32XSRdrQ0corhgZluD28w5vaoRjJU4I+rukgi4WOjEfjDc+Q
WbWkgthdY4Rs9dHyRgI2v6hbFr9xQI/Z/R3GlqDT/eqScUxfFuOt79aFERsDqPhq
qmz4VUJ1hHl3nmcxHw2SgOmiZK4lmbrc2/S94YILArQkgKkV75wNZKKYr8qg2zDj
gYTXvV+w5LKKWzznd5PfG/wBMHoT6Ry0/ZvcXizP7pLa1WMjR2QqprnfXJAAWcl/
TleXuvNtMiT6SF3pURh+QbSrdX3qOJLPjwbMJM/D7NDcH9NUjEtMfG6eFyEDw40J
pl/4YxTWX/1CMY+SXiXlVDoSBu8EAh3nEY7AxJe3CYdlgkoYHFfI0i3r7YbyjMlq
xA+xmvbetP2E4FhwUHxsoB16XguyhySAWnfHyaZKzW3N0CQ5Zsd1w8eKcGuf27bu
lXks3OtiCTzBxCP+gpBn57hTgkgO4p4H6ORokYjV+t/VnrEMA5dbNrhm3pNs8i2n
OeoKMNoSoXQYjYwqeMpIyS7eFyqa7gC7ocS0qv/Qq8SAbkiE9C0wB2jxA/EOXerg
As3YBh3JNw4zumjyxl6151jt80PhjTgwdy6CgbQn9X8M88DYZ4x0Vw2yjB9fMLML
RYp16Sh9vEb7ancmCt4tgXaUfhQMRyaGzwskSOR6eexphC9srtNJ7BYz/prsIQcY
rVkqJpJkUmIEr+NtBkJMAlcLFtDh1Na24MhHvlhMycN4vouyViK8y+kCsPyLG9T7
WMPJlhSkThnZNWqBsZGXTfgnbO8QkawTvXNPuA2sFNeU4Uye6CgY+7UoocApuI2Q
BmVfahmGUUYklNqlUWk2KDRlrBPB5ok+3L1JSn2En8JgmaCtEnu9N2fcgB6TUpvu
d+FH4z0391tTqp+fEYBNWAfydtfAOexof/Z0HHN5LsbAVMphm5GXBKXGtTBlOc/q
5kvY5/sN9iPs4YAwKLxunKPWRTlzx4jdScrnwUvrMGzI2WfPeZHNpHGcMfoYRux+
BlVN9kc2cD0S/uZc2rNAVlpqIXROrfcqa40IVdxqz6oEqy1W+tNLtiqijnDgEkXi
Cx28aPbkIkmDbbOWhA4JTGAYUvddZ5fqV3ZPRjg1hOrfpZW+fx0InSS8ewfvzz44
Qn9SIMoNKwL6Le7ysmq234UePp2K7F9YHOSj3SVzWKM0iZF+qn1VJKyCDSkdnzHX
/PxA83eLs0MlxZZk1lfj3NIkNp9thO09r6GGOuXsTnwYNrkfALHeeidan7XKvWVO
hIATu27hikD5OtiGdqilbL+zWCa4z4v6+7C7J35+J3Gkye2EKwKpcWLDLmaDYyig
RpWYH0bAGquoRXCmliIJL1YBt8pVBNTn+n2XPGUBk2ZGvw4sbkBn24czPGB+7yOb
m9OC8e/PR/9KevDmSYfG6gu5jvZooItqsqb7XWzdwtGnw9vk+sPyUByqyafdCZB2
P/t1aIL/v92z4q17sN9ntMl6MXbVDSsA6XDCnhwrGhLLQCGBpIf70q9WnDRejhk5
adBisrwceYwip6Lo8Iq2twqzmhwdVCNYhxAWeUrIVzTC3k1zn70Q+y/5gtcGKjnO
VSX5tUCEQzoZZv7padmi4MGDHYZk8EtqGLZzDw4ncLTLD+csIoDVek7HAuIuvmQQ
796gTNudKrZA5FgiDlwyuyyeMXqRVm4gmv4Ay/6QobUkh0qOQXLx6khw8n7r5cW+
1VQE8Bhou2XagliQEFui1fOwer2koc74uAt8EYRQhKRhJKLqhxiJEkrKNAb4WF9Y
3eHw8M/lXxXcY/8zPvi23NUV6qLkCvfFWTGyP85m+Tl82ucVMLDVkUuAmPbwbtJp
ntnDvsza3LhQtVjT4skFVv73TiZVGqAoFz1BOm/VL8DjeJhQFqfs5l02NiZsvO6S
YnManBWbfNKr1q/fWSuckuRRHsmXvrQOuZbeajoMz/pGu473gjIkBzzRXIxMbUCb
9Rn4sBRUP0ZP8gKWzMGh1S+nZzzO+Iy+8peHdmtqp1BAGtUsRs3FRAnrVJfMCuhH
2lNJjpp1mAEImbzZB7NlYhqjxxJfK838oK1SE8/pSJPvQZyIEM6P3xXePO2whe6y
UEyz4cFe+vJE7vcG3KRAOd5vLYDMGIJgY+9pDMxcTm7t00RKVGlgH7V+kcj2tUpM
+gIznjoLiUzsjxryWjC/f6Gcxarg8MOC6VKlOMAP1gMb2kaFBf9U7C1EkxiF5LZm
AXdlL08N0oKpyRXrdHPeE6g8mFdG6QpdEmi5R8zDRKmVnLc+3H9Uu5Axkx2WrCod
kCBrx9vNiB2Y4NRCbAkQkdiSzjY7VbZZNpWSo8fE3U0mfm4+MCsW3ZppWq+eGW1I
Rp51lU5aIrW0Jt3FDRa/RQPD3/JnhQpFfDH7hP7YRcYc1SN8DkrpUC2M6OMovTMX
OiKk4z1hUqwq38idAcnK6/qisky2HVKKH+HJpTNpLnrdcUVp/W8eMoSUuoK+L1qb
jqxLh0r6FNn6DphJTA7G+L2z9IWbf0eZhNE0Wwf1ie3MbPiL99BnESrZ3dZFaXHl
KdFTndOxGW6UM84gFbW/as/V47e/N6vkOFLWMFbi2kNedEjuXn3JJVmgLKUXD3YR
zBaBveuFuWTxEw9/rtPwgOVYVfESl640+Qhnbuu+6nRetagOfbkBXaKW1rDbBKo7
auwoWol5eOCJZ9x3UqcEVMMYq5RspknEVF+B9+Nh0MjLu0QRH/NXo3d5+XkKYhPj
D7vgIhtir5sbW+FEFuit5Q==
`protect END_PROTECTED
