`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EfWlHsc7UNrOTonO6nkEcj0rTrPdrMwBFVNzlD/0CvXFHuHN5Rs55sePjtz0ym7W
8qxdq1KBFanbveAHSZ1b4q/ZriK6EvbpK1z/SpwTJ5l4zuQhc85JE6WkNsa8JyeU
HEowTGhf83AJi48Kei8vgZoUJXaDquKynmHOHYOLtoQKX9rayF4lvv/SHfWS3iva
U85WdBlWjxmIEn81A8AP17jp/ERzuh4ujnl+UqBmzHBOTyFoMYfwvcqVo4lupYpC
lOUv8l118Ia1J0jxrJCvJsjsHANo0EUS0AafxZ/gEhbOpGyW5clJrpfo1ewqMLdT
DYbHYopzVwxVXelOI7KwkWFfdzkj8IFdC9Cbe6lK2riYRld4tBI+2Lus0E/3s2IT
XcpjXlDvyTbcOyeHrsZf6dHKKf+oiybu7eAToE7tV54w1EABp0G4FUt7c0rskJ1t
T/Dky3VYk7eiYZ/MGbbPTX2AVCLw5ovBMHzYxOxNrDGKAJ5Tg0py9xopNvCvFKBv
fD1jh4rJ9xvfHlTy8ehSy7ie2yXKNGfwl/9iwUj6Zj3Uul9WjTfoYnzCx9cbCPN4
X/qYunv7XzgMQf20+vGhvR3eQFAS1MQ8EwoFeHYT6XLmeYEfnHCalub5vjwEqlgl
bomvXcSFeUT5sQgZF4HP+ByA7pUmVhe1EmuGVWFFfYkofmYEkAR1sQIBQ2Qck/8E
PS0K/pzsxrt/X3tHf0jhn1hdDnYv1aZNP90uPSuFJiGVrmCZYk/pmsEOSEQisV9s
iVDQ6wVKpUxJurscyorYT5YwA8WrDUHdc6IDw1e9xzXT/b3oFdQhdHHx9khgB4Mg
j48ZFq305wr9PbvrvpEFsmUjPxEUirL659KBvItu4FPkRZXKkEbd4wSjbumwD7wt
fe+72NzVkstkvLFsLnZbdGuKfGGciwIWTCzVsZUHb+c++2qNPoqZSkn6zWObxZI4
sThdT61u76q6djM9GR6LMwxxq13ReAnh5k8kWVx9xYGTBFVZHGC6jM/QeGTlsAri
amwLtb9C5q6OH5XxALreCHE2UgftBksmwvLGymJ1zK+ZkxAWvZfboWOOQM4tCi7s
ePJOITkkaxB4Zf8/5msIqk+XszGb/XfiKlvuKUu1AMPmyiuuI9KfJ6x8JYdeUVnq
EHgBHX9PZFbEVCBud40n+1885EPBVFoRHRn9CQboEzJMkJlN+NjYXmJ5KcjhAq5k
90jaUeZi2+Mpk2lb863E/l41A2O0ZIZT19Y11xN8j7w1boip73QE1ABpH35gQ6qy
euSH1zoFvsZvyIVQy2rCCj0H0y5H1qG0q7TKZrpi0H7hvZ8ewAtW148I2LLJNclN
S0TpHc9Alq+Iagbr0R/BnwepiYPK9VzrhZ8rfR9WC2Y=
`protect END_PROTECTED
