`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8wpDv0hd3fRWyWJ/IdfbkuZ5ZjA6VqwM0w56G8PMi7B3lvumsQBlL/TiCFKoOGeq
SiHMaJyAKXGYxfiEd2fPC+SBo5vAKJBRz848O3pA6q9TxzQG0Qf3rYet6GmRacaP
1KrPyhxzx/hOUAtXWm0hYUF2/G04O8z8I+kxIGvQpioAbUO1lMEaCa/sgJgqKzqr
qgPpbmFhnTJ+UiFi4JkL6XSQ7arElGbdpcIM0K6xvAncTLhFyvggCkRO7vgqS+cA
q/nhM9GO6vc0BYFWEek00vm6mqN2xLW/TnoGjPqk+6Gj8OfASctL91EqsVnzrqAM
iZ24dhBaD9NCKH/IDVDsUyBUMnWaOCxYbYGVqHY994XuN4u5Ax4eD9mX2sirrR9Q
IeV7CnD3XbkWfVy++ZoS099hDv5JZ5F6jwZuQyhi1sTyUX1mDoVIzXjgfOincv3k
OJbrmA4le82kaxj0E0cMkvTuOBP8f1eNGdwS8u4Eo22+WtpMo686I5/x2RQgaLMg
xoy8dJKS26JZq2RnAQKNTwZ4plD9uye3ApMmFIdgAEQRx1iUHtWl85vmxEvreVse
JVaF7OWFir1na7rWMSiZU4BDxHeZPMFpAYRclqhI+1VVSo252L+85R5INOnTbHmM
WVm2YJe+KI5nqjIuBolN/Qu+Br+BAsJRA+1zeCwrFd5mA/PAlpVFHDL98fZ1VKSN
GlWNNV2G4+CFj3r+F2+d2PmF1J/a/vNwl3DS8rtnnO6lQpA7I8WJw38iHxQ3demI
4GuujWq3mjFHlodJeWNt0X6X2p/NZpYJN4yawswvyNp2eaO/2ShX/6FVB9p0DvGy
o4UkCoifVyTU44TgcbGDyXXQWHDLHHnqdykGg4JruA8SSsHOuhbfIrIg/UgxIcbV
P/JvWmjS2PNdwDi6DfjMtAGqRE09tUfdGlpGxu08VyjpEmkH0LKqUcJyJDFSBWS8
VtLcMDOWPMnHSaLyFOOwGeeNi9JwW2lO2mac6DjyBvFWK2lv2p/ZkdIzBFr3MkiS
Wzn9+JQUaizizR9hEc1Pwx6PeOwBI1EQJVmzWmrEIFY5881R3SDCuEaT+7Z3Me7H
wCoy0LxJ+xa/voKYxa9b/Sq2rZ/ZRdQBhI7mRLUKU8AwkakqHKAjsf+NQP9GKAeX
mjRkt4PsjBRaFnp2gSrxnjGkutVglhKjZqVvaYBMA0qt+OUWMRTz51a7su0GKjEO
AVp7lkTdVXimfeoYgCoU2hvbtM9Uo2xXfEuKmBfyAa3Knj67M/V/DAVljx8pj/Gp
ee57s307epjNnCXYvvO4PFOEvzTA9MTSfR3m/GhLMH94Mo/Zbup/mNbwJZjQ9Zil
/ms08kSOKhWI2/GMEKNbWi6xqhI3MBuO5Clv+eKizNKv/sm9JDKZ8kGgNQr31iGm
GXM2Zh11aEnXP6zXWBbvA9C1HYh0gbGK6aeU2v6b8OdxU+vwpeU4tKRKq2yvUZi7
tLanMMH6blUoKdaaI0+Narg2pEFYoV5Q5aZ8YZKjXKO8ORUni8Vn0GZ4/kzvxl1z
dvBrAlq97mAKFs1A+WtZ1u6CN5VW2AmUGy/lPpfv6hpl9k3ZYyOKrOP+QaNkF8F4
FXT5KosC1MEdzrk/Slnm9oPPYh+oUxLojHLKRuJZwy1RpzE1rkFIHUtQLTOGtsWJ
WOdhFMrPxgSqjNpgOvUzI6NoaC5XY330dpAeWv9kOcyQbzO3duGb4g889HumACBI
XFgPDu+OdTO+XCsjMM8VrjBHvUdmus/rb8GyFdDbSIMDdc5gPEETWN0QY2VSPuzJ
usYJe33BO7UAhEoUt5hsEMfWrCG2zBPhqGfH0yrc9KkQchXNrZySNQwmMzdLUDXE
AGfjyQ4IS8kEM6LOKuKk/Txw9fK7RWGBYvL88jAKYn3dOMfSRy1qGeCOA2qbW/83
7+hmucr5zDX2rkhWAilt/DUbquFibxL55dMCuNm9BzWWJtQcqjCGtMXUX7oFveGj
K1ch+p0CVP1bDkkITbxsX7RVwMCi26XJwtrqyI5zCeF4WMofziNeZNhPdAzMwjQb
r+gW7PbreyAM3kk+2trs4AYDr3To4yV49yXBDSPJhqwOJjecXIsKkvN5jrLB3qzo
BjhBjg8wg5E2H9dAiNlt4h83qnaIdUXCf1SHcIvGuTfzCk0U8QmgBWJsdSCv4B76
Ru8SUDOs1GrCPkIhPECzB2k8hluZ7VglLY+JtU9L/EukBE9vrbAHVvcB96K49/y9
d2NaVWC2hgn2HZ6gEA5Xm3MLYDEIkOD8AejjQ73MscfKwYyax4xU69GiKe+KjdPB
0Ou4QHecFGa2JThL3Ex4o3A2GuTT/pCsoI5aQQQkrRFkg6oNaeMlAG0wyjUnarcS
s36nP0tYhrozrNtu02VeQqGKQTKO/2ijdPoPTOTFlIYMjJhKsXqHEbdWbjGU3Wlx
CNuk/KCJ0Qh7+HixX4wNFe7Od+iU+2YAbuHDe9/en6f0xMD0dCsmq5Sq/b4Hj065
FVK5/NMOaA+WNYolVnVdrK5+b1DP89lvc9Uko1TgGUDPy4jM3FzRkcowPigf17ay
CN29oqkhNBS4TsMncqbE89+uBb5I7eKI2yFT9LG1+G/18LUiVcnBoP4B0UbM9mc1
iVb2ofRz8TIjwzZ23Uy/2PinqjXiZ3YznEGNESDaQ6ctl0XQhE3tJS8xsKJe7pjS
p7ClHk1IrD+gkGZaJuv7K7Z61PCbl4rTiyuDwDhMpHOx0zllmfYb4BWbYqRN3vLd
3neAXEyjQn2+jAOq1/tx8OUVU7jvg9XTeLVPZUvYQM9XAC2EWnFtsj4zHv/IrRzA
hpuVoIYRN8FjAyDocDES45aGeA+g/H9lfqpu9MSXeNrApsUBt004mEtSv/rOftCG
TaNLu4ka/sl2d1QZub+lg2uJ4NoHoY0Eu6oAqoaalozS2QMpl/iUVZjIkAToNmkW
PzB6kE8f/TDjxpOIqb7MjqD8+nQDIdj/is6xQgY9mF7W9gJz4WclFBqUEPK2r1yG
6I7kqWmk90k8iH5Jt9fIlrt9l4h2QRv/sMGX34QIIhqroWOzE74hfaMXcP9noUZo
Id9/gd0wZfNNk4F7bpU1y3pSETur1t671P6XAkSGvB+Paypacp1FIBs42aY+XnXV
WUPRHVMTe2QiZJEKXHV8TbZSyuIkrP2AuyEWAFgQ+APLw2IDIPZlgJw8yGjr83De
7pnXO1ZB62Z6rFKLmS95ZeJGG9yeSuljHpfeAYaWAfbO7w0tKYAJc4pBV4DwhOnH
FL+MnMT925dLJU2ze92wueIIQh43gV2+SvBg13T1juMXv2Ueboj9fsEPeAjah0Pt
xdKR3I795s8j5FbPx6kA2voNDI7JloQ5W1d10aJWRs+mXyWOo999V++zqAOyy+O+
JCRqyTQvCDtfvFC4+51+kB/EQRWhjbmxLMlkZnE6BuTMffztMxPsDmprAg9s9VLh
bXsqvf03ly50QcIeT8gpsAV7C45znmEzLxS+HsB7GqtKi4jPF+X4DV1LD+zeuZ/r
wFNQOiYf/XUVYpOCLbnSeQw6nUBTlaqGljGDGGNXXT4karBdDLgabq3/avnj+eV/
ktcwqBSBnsLh1EOhWu1oE3Ica9xZqweNNDaVIAObf/9tGaCt7rzcfUSNq3F/dIl9
kFr6nAFS1MfNt2qSkuQoIqOuZECSgb58MzuH57a/W/dDY9TOaNGtoV3gg8L008YQ
kmA1OLXUV1rFnrgOt+QOk10wqsuy1J59kCCWDP07eHA/Q4xozU+NIZHEClSQe0bG
HGhMmoR+/XLg69tqq64tVRpCJ5EjhD2f+uHfz66XDu+Vv7AnNc+z5bcwoBeQX6fd
CvcCM0w494Tt6W/6UAYwwH0SbXG1YNnaMWM4aGkWTksEOpXaA7xdOiygzCO1Ohzi
4jczrtRhbbYB9L92O4Z1ubwrI8qQsuRP+0ow1ZSVfYOh1PupLFC7rfwbRWh9sCXd
oNFCn1joLhXjGr4UwBGbuDfe8DgzQtKO1SpHhDrrLO9tewcXPeikQkGZWO/mXBPT
sDoOEhPMOWmYx+j0QCyRKcCf4E8NsrEABMm4uhdMT3c6KD/OPD3IgZhtkwMdznb4
fw0R8b/jkcaLEDFDTLWeAE1A4Twm5IZGBuw2//JWFQ1vSVTLcEmCf5VtAaaZ/fiV
Sw4cxPxSkmtFtOdnTBrx84Qy/kUJu3CTJCERJ4gge6dFF+y/k50lNWghDej7Mcdn
fx5eZHpqkCzoQhAwOAC0Rk2sW/kPwZhtc0CXNI731GHCtfBnbD8fVMyYVjWzX82J
eCxAN38uqZGk8tv7z7TRv5z0Ql/MC0dAkRoW5pyiR4Kuj7sxN978ToEJ8DjsXZW2
6s6ch5jzTw43m1yC0kALjvH5Bn4MwPPx+r4J0YvUhVsySK1DK7+vhkdc3M1xGVjs
FyUcu2DVfWcKOpHOcH8jRdv/0pVJrqxK8nA/6nIoLM80xfQL8DfDOeS8kLx//8HK
BHe43iLoowk49RTFUn9GgRQ97jW4zxjdZQQO0KeCYEq7bfib6gi2H3oK6fayB4Pr
xW0KQqodhdy97wJnmIuMm/t8wUwywPUb4n0sqWh8KcohKNCdDtABH86vVU/v7vLi
svlLMDh+Ex9W3PChV2jagoGi1sF/zoPuGOvSjoqii9Y92I+Vr+8c6IOWDZmSyGjS
fXG9PNTwZoxBmwR51qawWjtpA5P9RF8kaM1elFB+fKF+mj5Kp7ddiqa5iseOwsqy
5NEx/n1OHs5XLZoiGnUN9apTVRZyj/2ymr5XKrfy1bE7lUb8lCqjk4waua4XEok2
Jz5kB8ef4ocNSybDwh0zP/PvQYMZArdfbIFHE6IACEub17ZogLgQh5QegBjgIM/u
vUAdStPyfUEZN4xOkTSkWVNK4K6W3iew55Srm9KLaPkkVGp6InIXe5MZQMTpiBM/
vHl97rD+2+YS07XYIXGFCnLrYi4ODonlpYT1Gna+rwdGs6I4/trkJVlwzKY8ahrW
whs8VfGgrT+i4qXSdZvIv03Hq0hT7Y4KFKlZ6Ly1t7kPDfU7vwy4PDPXyHBfnhlr
RFaNkAcgthjtJfcez64dfAiodF/iiCqyCrN/LSf6GG1VBhz5FY5WTlksQa1jT60p
M+HR/HeRrbeFTzWoeLEAit3yk6mEKLnxJrA27fOidUWQoBdcWumAuDQVKPI/w1GZ
YDjRwOfq3fbfbJuDSMVW7GG+IZGKY/4HgUnDhnrY3h0skbF5+0ZWh5+Hx9aO/q/P
+ayyALnYoWkFHf4ocErRRdtHuQpWb++QcxxhPGCOnXf6iRVlLzPGOigxZ/FIviXP
rQIOLoXMPvto9aC4E0KcPFsJTN6lNMyuYa1r//dB+qYXLUKsNioWc32R0ahx14+P
ZKGu5bzkxiPys9lNU3FSNFg9b5dFuVLx2NXAWTOumKAC9Ib2j6piA8Sv8twoVN24
rdv5qB5MzPjgW1YWtjMv3AjyT8AKbwnvDxCJzwyLVuumRRipFiO62k29XdmIRgwv
udR5siT1Eg2Bt/GAa00GWM5yI7R+v0/WcZqpxU+Kca/A3iibWDQWW8DS9aWKRwis
vCQ2JqJSke7c7NR+R2JH2Q6ZnIhXZQnNv0x52bdL/vvv34CcGBZWwji6xP+zL6CB
4RgsjHJCFCFb7MapjG1rKSom06CYtcARNl9Zqv2Rj23SjeB8ygdKBlddcGkqQJbG
f4TK4Eg7ejxMnpXlRtD+lCQrKqYz/+vIxx4XD60WrAX0qHDMmrl2b03IouRUu01t
9vjePZgT757WV4Kger+UOH8Z0DseV1Zi2h1AwHwPIHA498IYp/wnujqP/nSWhwOD
V511XqjMWoS4sh/maaWh8nCAWTsmy+Kh2sKEVPIAUyKjVXBTLSFxBZiN0RXVr44f
A6uBO+axMcmsA9uiKpN9CfWLkkQUR56Gf0ihKppE2gN6mgbFWvrUvd9/PqorfNsE
XIi2J0vI7AXOsbdQdv+p/CWC+1ySfHLZlmDJb1yRvrIYhZ19As6lN4299080ExV4
C0dnR7GqPkbrpTOuBB2m97p43KIszGkHQXvPkjkwMKPBOTggK6i72HrsIqjra/pM
jSOTxxmzdmVlCO5LcKHxv4MuGgZuVvarRk4qiNW/NoovTj++z2xohhEgvY7xDNy7
+pCW6o+ezDquwu+e6L7VTNZhoNAVhwAuNotARLV2ubLVUqx4n9Tr2N7nijq7j8ng
5jIUZFx/gsW2V1B9OVCM49ThJ4mAtIpSdufS5CTCMA13Kii4ZpUbmDt9I1DT31BP
n6ocm+EQdT3pYJ1xWbYcUsQ+s9FVZsAEJX89U0H/evG92UbwqAMVnpuhD+fvhmHY
k+SXuXO5goFSRoJE/vOPvRe9wd/1fYEyGBiB5GJ6Qj2ge49fSWRyKuiUT7h3bGE4
+RsVO2NPRjjHJHIpKqbaaNwV10PImHmDPWE9MExxtIx9k2kqzUVR4K/U4ouyrzWE
vmVhZmoDAoJKCdfFdQQJ8hQHjLOa6qfnHPr2ytWba4AtrXKd7NbaAqVS1ScqRIxQ
SyGdZE/JqvHN52rRyNoPQpFDt73zQ+rtEus2eqySmVKkNfbDbaj7M4ii4XQIO0Y1
1frNm3TCRzSyWQxKtghO/9y2ZvyHBx2wrywIyFKk4Zt7JWN/Pr/6jQBql8wd+fcS
B7k5IMpf/7/dFEIW9KbIf5sXuhYiGeHJXOHSUsoSIq2VHYK8TuBCMjipaUJedSYv
pA3EEamHLPDOPXUEwIct0Zj/Xo8KPsBl/7eE5yPArKTI1yiiYCcuXERbsZDHcBcj
19BUf70ZK7xOJr/sy0bLUSJyfoxk3fnKtw3j5iOguoyPzgV2O4lCk6Rr1majEI+x
/16YAIz4WT4JcLuKE74Vbo3taLia+JmW+NGzq06FgeoVmlhDNWIvAKYIV8Qlh3rd
H58NAsKtl5m+xQl2t0W7kKWrAkgPO2aTFFmV8w9yKrKikM9XEBmvD1Oj68INJeOQ
JYjmti2/MNmgOyZPFqHVZmFzcabNHaRcF2+jVUhj/d0ynMURaIJObzGVED9F9/r1
6qsVbk+fRLWPBZCjkYxRRR25oCroD2xB78ql90QxhCAofFBWKV10xbxvJ15wBSoI
PIhYTDZ2dUhUvv3bc65uPJckMj5uLVRRizuhoXQewMF4KtXHSLj2Mc2GLdxgh/00
Q4S2BF5vCqJkSAaO+RWflIrxBBdaipCZ8Or4hyF4LhRGT6El6upv1i5lTAVbTI8c
jFCSqCzFrqT3Vmqg3WM70JN10yNmTtFlVl5IIKboeKhGxguvkAfUY9QAyp7TD+Wt
GERO6ND86tXdKSLgLJF1LwH2Etsb6l/tFkWNrzWHeWIuie2rWTHeiwGaSmTogsNP
9TLsrhPKKSCLpRURZMxyjYz2cBZjcz3FUOtR/0/xhO+4dV/30g03aPevBQYq+EZr
jo1pqLZvJfcpwsgIaRO5IziOPmZQSb75cLiHGZ6t1Q69o2ETGQjXzXmC5m+hdalR
svZwfRFKzFU7XnBtLF71qtYgxXpkQpy9QhgQEjmeUKkK1hH/572cafJ8YtQYtJxa
X/URxjsYcClmSg0pU+eGp1O3GPl+eecCn7nSYZcM9tBzBiWZzm3bifO/kFLcSv+k
vNGytMdJH2h/swEi7DpL8htEpn6IPn0N9Za+RprtN2vh5ODoiWihEjMYtN8gLhQ2
7NcawbmLJVDZ1mEjeKyeC/2q/m+/TX2FObMmruoDAloK9osDooMK58yKyTUznw3T
6YKPhpKFWo5RLexFu3Qq8zfcUsohqtUPOUmQ0ZOwoRYyHz9Z28iz0VhCBR2qVgSU
NJTS24st0WMw0HX1vepsKTO3oLezCkgQ8UlJCPi179EMfzLMPHnTQGzmhT8hFV5t
MkO4DFXQBKn4agC+/U1BD4ugd1xeWmICKVz8RWab15Se4S5GrLf7NU9FMVMZ1CZF
nH4l2IFLoLgb9G7yxjk6KQtCy5iSqX39BtluKHveVixVwp3tzLexB75vOm2pJ7YQ
hFkaRfQfMmO2MYl0MNRWhKm3lmCO/RjspKg1lw8PjjyohHfGOR7x7wi5/2L2l091
3W+qKiGRGGn5u75/6CAhVBLQdfQWLfrXpnd+FAdz+jrhGObUcBVgwySM+3PEn0wI
7EXYNjwgUZ8rCVLe/265n+vMuccGawO3R19/NpMT1TTLwIx+TFKsjFqlv8CkmrZg
eiqqkQSBnGDmPp3JUSMIIM4ieoxe76TlasyR8JUzT3A4ynoxBJdqNINpezQAmAGQ
8J9fAF27k+btjFf9BP3L3kaGetbwS1LxCKgSRqjUa+BuL/57WSFS/PhikEE79Ns8
Sr2xM6yJyur4nQJCAuCffiDv9YOVC9gvgEzjx1ldYIT5TY49hIToIX3E1WagmTw8
XH7xG9zOyaUr0fZOk/hFM9M4iSE39n4qEmxi/Ew7GPp/KVDLTbgHgRhOQ7k17j7S
0mH6Pt5Ttz5NFhYwi+b8QicFgXut+kW/7uaKLJRcgRJa0fg2a7IFJWzTqsreikAz
UtDbnC3KoElgOB+VFGgEyRh/EpSjm47cZJUlUyXhhU0Ji6h2OYBDfmeUnhXPUcWn
P6OQ9V2NvLx7OctIISzvvoSRmMtGfnitINwdg843YG3VrES/S7TfRWfJmK44MrHq
POhzAPBu0Gry4Gm0M9+yFaPnbEC7hGEITz9Iar95X/2sg+I5sBifMr0ZYNi2ealP
5fiVq34tyaGfKWbP42kCYDsvbVlD7lAV/q7scB17GGGmw5GkZnvzNuZ+GVj2ZW5m
yI+sg126d5t9H7/eFh7teEVUmTYjItIVXpDDSjjY4S/wrq8Yfit1D/a/njJtmgWv
SUzN4WpKKvP1JQMHVZhRJIucZ79XlafyY8++vlyyQTneL76cA0dhlpHl9bRYpEvT
qX04mPO0fJcosA6erhdsKItNtDH90bNY/JFcmwcKFtPDL/xbEsHCyMHUjLPZGSTN
3dC39GARdz1L6g0tUBbvBYLimZ+DBzi6mUwlMkBAwDk/pLymb1fLT40cV8Ddds+3
F8/GEZR9hZzY2SIeSIZlMvqZVfwt2C0vAPiCF/VpYSsCiTeE8zdf726VUNJ2Aq/n
XwbN17FGyuhHuhPq9zOHCZu1FLQHx3Z6pojQas/Hhx9m/ooOKaKI45jYyoI5sGKp
5CgXgUGWYP8ZZoSq9Ds0lYb4SX+graSjHFy5CQbU3vxwiZEZmAs5KuIUypOoxDGJ
GjumY5MBQLUme2qBe8RMd0YjS11NCccZBkqyFt7pTi1kul/tii57lSwGaqvzgetq
NpfiIcBOiju8EHHV8GIC8zaw+e/R7LxXbuXjkevPkoJcTLSSuKbSqra1Y0Hh8aoe
ly9L6SRHPEX5q/vvhSqurBKnOqRYFlQ+k1IAXQ/GjbUhk4A4s9v+6tUG/TsT8A0i
1E9e+TI/uyjQ+7/pU7Dtrf5qMW2DCWFsGYtRvbCrgh8MUHML8J6s1dHiZyaGpRIt
6/DXMYfSSvsdQIsDhbf8s2TNX+d6vIYQXYnh3HenDYR7/uHkHfsYVLo4xiVRAsJr
D4r745vvoDNMaRZH+P0LRe62kqbGClJSdE1mwqsVakftpWR5LzjonjzZzZXbdKP/
uRdZpCXFshVkLsTV8zcM6OKQnRW2iuEZaprO/C3ODXr+OvKdwfoizJJwXkERnjxZ
ZB0MpE0YKPajkeXWswstzJmi0UHo7wG6nP5vsywokt22mjlY68jh0A6IvbhANTTQ
AWtmoDPVU0yAvZ5izpWzSGvGf6c+3+0T7IP8IjD7JXHgrUravRh5l3ZeMp8cJwRS
xiXlcu5CK/257KpVg9JN1DDDwYqf3veN7oUmHk3JXi2OoLS7AIcKbsdmnCqiyBZv
WUytzfXN46061WhF6NrCepsvsUt8pGKmzpb5Wxg2MIXQKLNLbyK87Ti/uVoCHj3r
m8T3AVipw4RM+QKUly8DCgh6+78W6sRkSkKaaWR1u0gZzKP/9cAzMQn1Thrn5Jeb
WC86MGiTmewsNL2gasbeg2s/2dXIg3m+XYl9GI+iZLU6rI1k3mzJRc7blVi2Wt0r
/48AAESbCy7WR86l+SuywUHvuMJaQrXU9ZviPrvPQo9RoS2bhTDrGHHYDHIGSkvx
HXsKPkXYQMqYuLXQJxXHJJEBc4w5K4N8CUIvvi1LLD2Dtxx0BByqpX6yu2IKS/Xr
93fik4/xjXRol+EDLUQBoaKEqKkq4UD2Jt6AvlQDxfNowNTyZ+DF2UWuFLusVfzj
JR98nA2VT42kOsBMyKi6H16k+MUdqjzdyioqtHnTt26kGIZlUYNwdMqG4qoIivFi
szrw3lf+nNsQV3ut56HUw5WeYD3a9Fn7x8wp9B/R6b0Y8L7b2I/yH/T1O/gEjfUl
aYPbTkOyxrN0AdcEl11dd13l/el6+IFCGamgXDOTFdjUJe1WqLhVqxPU5gChEAx3
bYVQQZhAXI071jug3INoFBRvvUHiQbUf2JlpzHIlUVksEe7qU55jlCSRBobMjA+R
NKueZD0kNJSo3VxkUXfTotgYPVNdj+Qu2QKcyicv8Y1Zpz4LpOt1WxsnFupYqPZO
DY9y1AELBw2+OaqDxtPlODWXpYmoif7txhqjy/5S+1idPQfTI/jpVj76ICe3x9jB
kXrAt2M+fl48xPuqWxxJKfre/K2AlAX8ijY5UxV1qbXuID+lnswAYLLrXH8s7+GX
af6xjC9oO9lMtyjnpszRVPWSdIP2oAK3tAaK5Cv1ER9P5tXqdM74ODiCUqVQeLTC
xdq7IiGWsY2GMIUl9So3f5QrpkiHuxCBKuz72NeneYlxEx1KY9JkirMwlXZI9RSR
51LxqDa6lH/2vgOKykR9QlyeY3IsBPUSXwQC1eoAy/899Od5j1QpjbQp8saGIWOR
a2wQ7lLv+AR0sdCZ2aUbRdaCdAjn8JStebfKUlO8M+k1dmsvpysE+R758WUddWFT
mwH83EyklKUYncmhVnw0MaMDSscGQKjx1467czNx/zLudFHF9H8wQkXXIz5m00WG
x17Ej+XxCgVJBqZ9C6HqVgGAUTQ1TF5xjs/pvp5Je4wfrA3+nEteYwgAI6tSeM22
ljmmoG8j5BR9U4N6qnqEbKP93LGpWzPROjXdQtKbChnioqvjQxJjgTsHB4bOdelr
loGQZNVrDyaM1IJ4YY7GAQM+NwJ8stIKEGjbUDEt8f2v9luqfjYpVwn/w2nka5/F
d+2FpaEBDK+rvv6syZ5qxddp1GSsyGK8i2sRA7PHF0jYwG7k3vhWZ5vLFoKonpLp
dMtT9vcCy8XOeWj5Ziibs3RUDN3MkDPOonMX4ZCtKYGoxNaM+3005eP74GTaCaQs
H2F+GqWM2dZLFdI4Ul8yNvkfzmPX1ZAtTGP8UX19qqWfIuoQBCqtBHv5dAxJfZws
hW45nv/hSbSZytBqLl/+Aobsm/YnH8m66XOmMHaLKXBUflEjki0gF9FWTiggHwgS
rGEbqtkpWGDckk+rJy7LeGcgpR2vAF8Uhd7WE6NP02+YZ668tBf+0NB27rTZ9eCV
Mk8UE3n52cNT/S242Zpz51cyvtSD+yNlYFPNu/h6QHZtSUaGpLbe6G6TOOT+B9UZ
MEJK4D0IDTD+xxvh+FJuYGuW4M2KSqF3dN4izk2Afl6B5qQAMIyqjnWVjDl4h/Rg
f1ieUYusdj9M0aAMC6K8H5Ww6zhIj5mEQTHQ7ZGhLN75GFUJwjoo1dayCdgIQNIV
krg669KXu5NMzWxLRJrv3URTv9HwHcaOUWpBup07vpws3yWhwQ/hj5ak2k0blX5o
Gp/Wkc3PuyhQ4XyBLLODbummkFpIEIvtTRuUcs5VM5lDjG0OAqbiZwe6Ip7ymwIN
QTekS1sWsBIIjtwRIZDtWfl7OZsp1ydQZkr+qKMx+vtDxLcLEg4BoL+f5qz+saLP
6PbZAG2eP9fLhzXrpZUVjjWou8nHFoY2Yat+W4YWucNG0AK/a6AT5hDTq6ivPokx
wxAFcHjikh3IayNH2SGgnyy7CV81vFaWPVH/9SWZs92XMLZRcJK+E7xaDvkEupBi
06sfqL7dB3R6IWEcTAv8XIxA2+RorEYVJI7vPkpuHWzFEAUMDXu3Ps5kLj856oyW
QOltDVlgurenuuctlDj5Q3KeKLTK+KDdgYkFcA8XqfyKa3hbDRn5WUl8G+2pHlii
ezts7RQq57ZI4C91drfj9aQHV8E8XNTRAl3spq4lOLuPVgaTqjtECTZIkSOO1ce1
nYTrAaKydNfMClSpuchvj/PGf8UfovokSKJeth2IKao5n4rjqccQVLy4C/H2eNdJ
y5p/rGIPKwvGgyrSmzb2F3ZfMxnVkhHXJNS2xsiGsrDEDOP8EaygUSm+djPas9Rj
oaRammE7P51tBTnMALUxaOtELAVbpOQwZ6HKOjRO3WNj5t7Bo+HVcOd0/3ngb+YD
OKDdRBKPARkIl26nBp6e/d/1uW6TeFxseQpsvsjBD5VK5ROaY3IkgPkvrjqdkgqy
efc9FDYaTXOjoNz7Fgp9h26GuzMRCtxRIC8RTXkrfTvIqegDeCdYMfaqFpaZ+1Nb
UMqD4Y07mwrZwJ5ZJGika6Frvom+NIEUPzHV+2WGBPmPcP0fHZMWajcAPd0A7Smh
tgOjZ9usIDwSUUeVEh/tialFyKtP8TqtagIfrjJ9Oq814SNO5lKqOoVgr88SfylT
ICuKw7tSJ+BEMTd6/pglQR7sGqwrlwJYiXafwmt/sWkGlA9kLuP4SBdsXFNHm83A
gL3SO6xk6lKJR/mItnXzE7Tpjy19q/lvyQFbEMZPgL6MRrWWQGh+4WrMP1kNQovN
0Z6LVL+8slrRIrX38XWuDKxv63QhxvwKgIginJCNMrfLr0GFc6fHMeE5N1Sh/B89
AQRaxOeV9pj11MWDrhCjjSRJ9J6LkqAeqe+GkIRB+bCRMbw3D0vPZXJsv2T0aqML
QGascXlNTEChFV3nOJ6QJ5RhLL2Kl50Z4C3/zZ0VZ8GJ4Y2XOOz0LtOnX/5VR2NV
Sndz712ue6YpU+XKbZrerj5lzZ7CQjxKK11kUCJjbGwSE7aXcCNU+oKQ1VdgHBug
MirOEUXkRnznn4T8NoCAI6LdhvLqvvEs2qFGzR7cIHfub+Bpy9yqzilH1Am7kSNU
WGacEV6m89WOuZdv6QJI/cojvtS4MtuQl6ZmGYmDAWUxgWLr4RySNDNimZLN+F7u
z1lRk6EoA2zXUnkDyzlXveBZDAZC3aSo+OimzG0Mpf2wkab0NMq5GdqLnv+s5S4a
Ip5PlbzhtaThU2sFHG7SJoOoE0fk8EvFQ6HtElWuVxcaFrImFYOMAUL0Q3HlHuR0
03YIG+U57KFsPDM9izpisSTGzMe9YNhCxtIOZUpjvFdu83MMlLoSC5c69WCkgzt1
O+0Ok4doAH+fuIZCekoQjvDc8gIwXqftavq7f9rw2HjFYCcokVNpqfmSuPY0vge4
J+kb/TGbvK2SUkSFvFQPuqNsHDwYE90HiC74/k579zgSaqynEVjep7ztKIscYkiz
W6si9L8v6mXl9YKZHAgN+KH9MojSLsjMRDAeML3PTW0T6zg1F2D6mweCM4Y0I51w
WLGrdO8lKsv4STHVq+6otNlALOKW86Wz0I0YQ1pJxXmJIMJfa2TyVHeW37BkO+RS
JFjBRP/xwL8M/3A+8mlVQRzTHl80EZb50JvQQ8It3b8a2/FPExLTYYaCnuy4bIBV
oB2+Bb6I0ZUKD6KMqG+wJEznD3fOf7CM/CT+TTrRtnV89HOQ/93FZKuovh6Ijuam
Thyy1aDpDlZS8f5EH6IQuf2eVt3ZaShp+7Zw9E98MwfjXT2RtHmhBbLKreRIrsDz
Q5egeyG7UxEYg+qjCyjOjkqE43cityliDud9mjI3e/0EmrZTidkxgKeyWyLlCbIz
5+bjNXUv+Wm1VFv+5hEV719+kekJSWP5F79lgsb8ft5Xang82nTGUG8fZd0ZNyOC
idiqeWc+20I0ycE8Fq3djA6+XI4COlXYwWuxeeL4MAF/g7RZAQN7gFrs36Z7MsUE
0WQbrwI35hY/rgAY00astUFqEC0kQg9ZXEYaLTAv7oFwZi2Y4ElOeoD4TDWELhqJ
1e+dk/EzfIJRTDilf3pBUAkW2ZlVS2Jzli1/WmOxRZQkCl+L9/dysfMqEtOxUOVN
nhpdQ3n4zivWDRsKAU2mehRc12NKGz5PqgOWZ3SsrdSL7EXOPGtObhS3/ENfotCt
lyU+x5wYNW7ftBTWldfKtFAbeH9PUDxukrunkCd1Y3KdSGXWOyXoddW6KaWC5+/x
bLrU2IlRjyzV4mHAWJUhTnPZsuJipEJDYIp6u4XU6iC9YTZK7UjSkzluJOCb7jaY
Zu/LxG5sS1B+EIZxWozPwHlLV0qKKAG31i6bcHaBY/Bpe5+mYyptjdvCOUXTuQ89
4LCN4gvQCZvMZDzjy0gmo9AKN2bkfFQXISIMLmZzgBiOA9EuH+k+IQHPqu60DGF6
q5DMqRYXVhYZktVTCtqfOH8mwYynJCf7CGtym/7xOkCwCezNGDgVM+z4sQemsupH
Q/cz7WuSLePPe7kamECtTalCFufQdPQ6Yfp4yQgofH+vgP5D9nYsUeDtVRTDQajn
gmvoOzUZwajz6B0dCJmhHdsw9qiO20yxsnFLOid00Z82FRRQhq/v2FjElswkHBur
DogtLFvGX+bATtjTPtjKsqYSHoMu3ZCYuCBJKvPe9Alu6TEst6h+HW9rSGLHbizG
aV7HlndSWMDAq8CHPeAxUbncIY+z3hpxipeRRWIW00NNI/6Y+E+emBxOLKlo/yQe
3uoaqRvIgXTZWPKkX1mxjmlvwWMqPvcvAW3PlF7jaJty3Ou6nF+WruGPQvFHZIEK
k8Mh6EM67CDga9G+W60leg==
`protect END_PROTECTED
