`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OQML67X/cJUsLw5sY9IVvWkAjjgNjrba+Sa4ZHItz84SO+1Csw1BA/v7//mrD9x9
W+fCrSEfyzk+kH489KYn4+OCyWybAOetcog0R0z78GfMNVXzO+OLmst8wR4pHshi
GSY8ku9J8Ck+llGYHZtDme4AJVcT6iHFakxtqfNDKL/GwNj8xZSaUf4hlNerSN61
oWb78A4MrrUKNfyvROiWf7IU2mwdbjfHMIqtW1QSf2lCPejAYKtjf6tj6RKeXFTN
F9itA+lTxh8KT+opR9QXfv4OIaLiVNa9y6q26c1dBhJCpv9T1iQAL7UFpVcl5sVM
wUFVzD1uRU7gbmRSfZbEuNuMreAG6wAMRKtm9uK8RWtdL1i5MQ61PV3IaOZ/OU+B
lB0/92z20uO2wWQil9qs9nteLHZ4fnpGRqr3fskFskJgysiTc+aGNhQpG/DQP2Hn
sm7CsTl6PovhmJ5zjza5pyukD0P7Fcm7bWKqFQ1mFvKHQpb4OCKMO5+CMAaRUYBh
YO7MJ/aB/Lqa9JI3MfPzh1+vcDbaO/rzyi0QGzS2OX2JNjurW2CKeWtuNmq2A5vC
P0+NhT3l7v3REcyFbRdMnretVSwAFBJgPaFvIqly3R4xw6SrA7VVTcYQbygfB9Ab
ClvCjPzlx5EksmsNqYRM0SU7G8C/KkuAZT2TKR4HSmdxrOQwnGg9cvFibhJH6IvG
RAHdKNuLT3j7iQaExDhorcHaAwhhuu5HtShKbn3uVuwy3jRvmR/2AL1oPEKpebXm
1m/TLQp21zn5AW/3sh/CXbA/me8JS1u7WMOGzGNkqS5SrNJsT5aVmKpa6/TCdv8I
TCSQix3yhci4Yhh8jkyap7Gm2/7c8z8hqCqkAvo1PX/sthTX2C3+LCvBmaTgL2PZ
ALjVETgFa4lE/zxtKq4nv0PDqjk1WV6RkkxZXT0dePdu4XkNp695Ddmv92UpgtAv
sKyGJ1GAv98yKAzywSV0XIyYbJVR/GhhLYUR9WC65/DaJ88J14I0wLS373WQdYN1
uP2yZAKSrRXWV5BhP2KRacMwjc2BvDwoPYPFI7oVoaR7Zrnas2bR3TVaZxoW0OKx
z1IxzJ5Zrg+ZDcDY0uoJvjCclRr0GaIOqFBxpkmsnzZE1BJcNZOmX07pWcdkyN5d
G/L00ALkxtWUTBVofKZ8Lc23DPjkj7yHXjuo0v1JvcGLDR7iidf9huDw0XRsmj5s
oh++9WSOx7kRDIYWyjRqnYSdt51N9cSwVNfEIuuKe8TVD//9Dg8BVnWU3NNUZuEK
+e8CKXsr0bY6ASV/PsGE8aHch53FK00EIE0YSDdohucw4kHoo+9n/dpQ8OC4VN1j
1gzrt5aYCChQa6WfhzywV6fFOQnYNQqr16Ow3KjhbWo8VeMK8YZBLIeXeYkCk8/T
mmyLFyLQ36rPtic2XjoNeZYXm+YvMf8jczVDyUou2biXpTgkQapbStfBM79Gg+jj
C3OG9Fi1Z6CR5aH3CMejlkZzxc/0LqKpn2G1vfrn03rTWjmM//zl8ouhaxIvmq5z
vebPN1CjO1IN5FD9+a/tGZMM2UXVevaB5zn1kCxeciCE4rlXcDVI76PaCqO4nqHN
SqPFnp6nI/x7vUoGQF1nUcy9/9+Orv2gE3oAyOuKMy4LiHmcmAI6Ingi3QHacoBL
Ao92mGPBP1cXuHjvQ4gQCMpNF/GCDJ1iWsbkLmj481E8mU7LlyrqT00ueh4SqPCI
7F5WaiW0X8j3DWjslf1Twk3Qs020bFYHfTdifwKXnzr/2xbfm9XU7oITV/UFzz2R
Nj9BS+RbeClE70kt87RvJZb+qpIzQVpc9m7sqLvOweC+1J4FltHHC2zcQFJogvlX
lO13HKrHRkhCuGXBspuefQrfx+huxD+8Ekm9ifbNKv23Jp3ZiPpD3o5KySrJVc2g
SKt3YxJojFgFR4J0w+GoReXfH6jIRJ6VGvW3IRXCa5rt9U6I5iJdqEqrVZkhQseG
lqIKfvBd9TL3SIs7JW/OqF5dSzSb6yqHZwrTdlavASZJrRIij8zR1lfv7B7HeeQz
/y3fCX9EU2k1XFkTkzSy7c5yAMsYej0pokap8XwyMVfQy1trSnZk2CSm8j8vxbiK
3/BQ1iVfy+7xftBfvXP2HlEwWW2ptW1H14jxgZ3z0uBAY/K2487kEEBGSJ1Hs57E
EEa64KetgVwGJ2DMmcLGNqMH/xnyZYF+VF5Zackxv3ogDHxui/N7tVr6jfTCO+hV
l2jJV+/z/ADbrkjUrNf1MaJSIIBMHxixjgF7gFfVEgoWZTezxXsRXaGwvC8WNNUF
8hrayoS6yVVQhYUFmJXp3A==
`protect END_PROTECTED
