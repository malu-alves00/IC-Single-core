`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IEF80sY+OBu5yKhtoCdEHyZtiH3zVSs8z/tbO+7cEQ6JnSTiIlRgDDcPQETHE5O8
SuagX+yku/PVHCvK7CoSdG5Wdrq/C71ge/JIhiPCEOTamhVb14BQhZMBNuVRdHNf
NBD4+ptnbvYj6nRkcYAOeYPLsZuotj7+Dosa135Ay1zx36udYxxmBlvlBco/Ka08
iAev36WEqK7jr6jMtPoS63TY+guOm9ko/J2Fpn6o0nA2PRivscmbCcc2QmchTQdf
TiwJ8O+faiGlJKU3F5SLuF04n8XmHDUvn6TsjuK9dzk+73YpBS4DzUWCfyRWbVxf
hP3Lxu+qU48pJ6tFaQQ2XXbad9+Gc2ZdKzUlkkMm0gxScwlbzFEI7L7vbzIridvD
GJxmb7JnJTS6c59wropQGgMIkQEjD354Begz58CE1D685Ir1p0V/GO4pC+s0fJiE
p8xeWpFBZUy0T0dBYnaKm0y1cIx/D0BCfPVoBidPKOMh0c1LRLabKwn9rfs5Ylmk
sE6u6eO1H8sH2tvQ7XhvqEO0SXLo+T1Muk7r7efJoYLWIIOU7ruyj/9TOAgPUnvA
e2sAx+oE1bUuiRgug+Y036X4tU9isAIF0rQy7v17LejmgbqihuT7G38MQrUoupyx
dKTshEBLDwdvsf+J1Ul+Cx4XAm7+IxktA68thqGIuc6sP9zRSugni8RPIdCOx+ma
mZYjs5TVmjxmz+jL9qK4EVvT8bG67OYq66LZTd+i45v5CUkx+1fzL7+0w7tRs8dM
sBt25o3XN7Yhi7j6EF6lTjiMmCJdDGWGDKoeA/BBO+tqk+higNtKXWxYmvGui6dY
uovVtIP7LQViA7K00TtvEGhPzZ1wAc9QtU5slR2uRe5i9EU2V+ceVi2u0mwhUT1l
xbhsddCSbiU6ZxdxbVjR1JAKuXIbNEyrStvWXjnRO95s224LnoWSVhuqbzsz2OVA
DtZ/ZZvMjHpNYMPV9Mb+KF05NRvzDWWXzRnHaP59HxtSInRIzvgKNtKPjBta1i0+
+DC2+xjVKNhhv1L/a7/hRh2VNQmN1toYvYSLrmLa2l+SWKik5EMk+HsGczhe200J
AIKM344zfJGsM8Qgzvn9uho5EH8nc+yy4foooTV18CmW385KkovJTSq83pldpYMU
OjmhWqFrkEJKhsFMDs+TbO1frhnygrGYXojHg2XRWZovWt563xVU33CcUFSxj5tU
td2gppNsLcBbqQL8wD57CoXZEOAA25rcsErGmTaZ2K/tIc7SxV2ax5F37NzItyRi
mrczE3qP24KIi9fbGelAK3vKhh2W8s1OeE3jYf/Ah1CMSTaf2cUb1Dacy8zlD9zL
usphnoNiQ2jp4QhfaBHERqLgpK1vPbJ1zs0GEiYl7ORErVsK1j8iGPlX/60tIetf
sgID02qflvzN182cTlHeubWY1s14fTVVn3c21Z9UzhtE4+pMy6W+xFn1V2Opkeek
epwWpSDjBUlkMRq2upq/VOgOL5FEs6NgDxZAqXtMMv6TbRccM6DQE5XCvDdc0EUs
o+KzBeUsQGeo0AIJL7gEz9qEhVmNmsBxyVBrqE59PO0tHnv3segvpcoLwDds2bna
1q1aQR8YIXtI9ZZGYAib7D+KpyzBaE24pBJDSGYbUnmGy8YTocnytO+3cBUDyVcH
SwbpGz0Xe/MxYL4u4ZqaQlC99zHOM1xA4DddlsNFcaD+xEUtg7GSpE9ugIB9I+PX
EDYootQSb7cRGivtUBST1PrG6CSqxJalmcGbMFC/ixR/Ago8jDd0pyy7Ny4VCfyY
rhKjhMb1gftpA8xoPptrswwS0dtW54O+hQbTNC3brMV0LgXq2wxOJC+xdDjyvphF
69d4v/FchkhX5gJK+4Jbr/cVWDf1TfuaXy8nfdvVF44tRRdEUWKFASdfTSH9k0W9
BYYkFczfAicP9kXBiSKKF3+h7jB7BIABYzW8Et/a40GXXjNmbGbn1rXLCohyeJ8P
OFzjupm1r2eAyXmhfAHeWYJG71FPsxog3bsFlvquY1rwnrnhZcBTOZCG56cRLtVG
7kNzXL0/82uPuMjj29Rv3pBCEGxyppkdPXnDhdJZEmQt6F98aaDbh444njweatZx
hLmSzNw4WmlJz78+YFTo4KmV9b9tJZ76xW6w3q2KS69omfKJQrl4R6U9iDevncOk
34nZDbmFqQUzNPV0jK0XwGNgSoWVgmDkbN7WBdFTp5bjX5MuEaH1hdvT2o0BTQK6
gLwZD2LnBpYsXOG06xq1NXDoCGzdxp9stkMhfYq4uYSUU9iMXY24JeT6g7FHTKHH
PJIvcZ9pd9XH34Xf/nOph8LhuVhoa04F6EXKOjP0qXCvg6QneZUMJe8MPX3mt4hG
B8/9lHeoNPAZoRMzheWTYiEfn0nDVtBoFUZfka6xDJ5z6ILO8F2R06cN2E/yu+7r
ltKrpNM+POUWXxG7TmaB+HtndDg3yzcmHs4VsTNYTHOZ4PEUKLjDygGTp0JjShp3
OCwrXlqFG29hQr9E5VwN7xZkZJ75vfiPbK31YW6xejcc9VraQODWgYKUUpxRlBFe
WFixYCV/MZRpJcBjOuQw5GvCEdOjUjZ7VfkY70o6LoB6pku/EcLkMDZ5tVIG50UE
lahefx/3dMTAMDd2EkHfZYClT9E/oK06b9qqQ7KywCBIvRlDQf1PxlVMUB+++6cj
xW+5Bm4zcJKbkq+PRNQjjenviKKGsb4SRj9MzelyDaNaTK7cSKqpfAp3AhtyYuL7
cMzK6vq+9MenD35caLGk7qIOlyaaV2slz9LSVpcelJ5gSblRj0dwtXnYnH83okcx
Exg9ts10Z+jURXqghqe4ZpP9MxIUQMdDMLNuJ4+sJ8XbvkYIRBJC/P2FjtyP/yds
BADbZwfhhLfwvmE+Hr62FeMOUttgX51ElhkkIx0y5Y+OtiQRvIaiFF4Zva1yp3p0
vZ3KC5swuE2cqQxLiUyv7Rcf5P+qa9gVoc57vtvob/OAbRvMgqwQnxeasCW3LBUT
TedJ1GgSOUwY/Hu8l8TmjwP0bwmBzbZ5//MCiJAtsZMTiUUCa8AMWLbyxVCEAr5s
YJqfdW+UhSAeelsnmuZ0diqVUQ1HRl/+i48fbMfbOUTU6BNSljHIZDho0BFrlSiE
naKqmjXNU2iP64voYNLycY8RkNwwz1x8Iu53NZbvkrnqvt++z9TH11C12jAiFZJt
G/cSVv+hYKkhsYs0G8I7ZvovfYJqhtHw+VUXWazpNPzgwaHNs/8BfPs/+Kf1o+Ud
eRGRYJ5Y3awZQWNAKQNjLgAsB/2/xIUnimzoMEUkfDR3BxaKn9cBiVJfL1ThAOe3
SNTg6Dv6qS74yt97b86Gc5WhlxDGCNeFaPtl9LP/hWNC75AMF9irdTPt3jWwdSRF
IOJHfjV4lUrc3/2ZndfoELMpZPvw0G7cl0H4LwP1k9BVCdGfcbbFgY8DuN6ZQlzL
R736tBfWnqQ1ODdJH/XTAkDtkKzxu6m8wlNWaznamuTR9d7aab+QYjmnzxZYmn3I
Hn9IZ8YedhZFSOHIKKTWj8i0TLGBaXJ8u4qkJzlkTIQ9d8JzVbevm8LecQHFNeIp
yFOjgI2rIHIUjWNdz+nh9cWFUyvYk39MwTCnUpzTMynjvQrxsFNPqxC1PKmNTR3j
tli9NJlrAr8byf7V7ku/M8z2f4zKk+UhU8Q1HosRm1D8yhs5KXes5tTmja3SYeog
oIvQtXjTa1enrumB3vuvtG5NDuPTHP30KQssebH8xcr2JCjD7AiFWkkBq/BxlUrc
15iX8jsYeIgCeH0817SBzHZ//N19x/ryqqojws1AVlAA41xJg2erwHuMxVsU9Lw+
MGyV6cl4bbTFM9vVUDVVb7npvshkHfyX3pQmK+iARiXYIXZ26ou1fEgTqVyY21M6
45FD9PHc7mRK1TBGQiBYuHfzluZa+KWiDeL9iVNwvmVEXzK0V4f8xekJj3qbw/f/
qmwpyLec8m6dPGohD+kxGWvE8RBgbEsrLWvvP0nI/e57exUvQpfcRZGRmFYHTSwi
G4LiOA6A12hnJZbNDKPad0vV1HFKJbFhOpZHgsc9KfKybCkzo5DTamPxVrvKCo2y
EDlkZoxgtVjeN72J1k6ZBZnM0B2Ijz5E8ES3QRs8zoq3j2h/1Bb0N6woonSuBqor
emWpu22LBtlwtK1D18N4qaCilzQnjNmM0zNwXoXRzKtKRAhayrUUzz2gBKisdBYu
c8T0q1Ek0YNsSx7d3ZBIRyWbOuwGJJJVkwaG/jbfcjTy6a7T5FdPPZbmNP7ZpbIh
6QJEBLU6F4bSDuQm0mADrNq7sjIscOUWJbfM0SUxijqw1hwqHzPQ+c7tNZLitgKf
u8jWmRvjmujXoc4UTXgLh29s4BJWKkRODrSuubjGJI/SQw/7J9Rrg/USI/B789Jo
FE80JnYYGD0+G3RHOosk0hBzn5NlGNLQ1YwjcMkJ1ndC8e85nvNDal74v2hL+k2J
je8G/IAulNyyP8YodEhhTnXGSgqTi4BrgGZVOkpxJlP+z4JLX3IpSvUF0S26vg/F
7CUXyWNBRxCAi6WlMYm6MSZEzxwITlssqYz14lLXl9z+xCxjZdHNktqTt6lr0TS0
hD6WGXuF5fRslbpl+iqjqaeyZZZ3b4BN+4ohzBoEXH3GuSc5+pKIaKlhusL/v59o
Gk26pFJ7qbzmiPZ4aG60b3lvB+NthEpMnbmqRXcGt6Y5Voqcxlnrxgkhu/N8q6Wy
8lecs0WNgGjMkiBytRkBBUev7xT69+KnGxgDzjPLkQBcJT/kS5gVfAR8rpkh/a+s
bV2sbFPwEhx2piTjgxuIxYfKvixYXPFe9Hm9nkRu34ZF9mVyyusBb31J1PMNTl19
crBfzAM1hZoJTGGDqLID5TDrjm41RnUB88PbgOsM+7zYY9EzBH5BOHjdgfPyIQXq
Iyb6QmwOmI7fIaPW6IMMQfbHnB2JTGGajp3me/MeoOyjA/y1nMviRX8dGVYl84cu
PqVOEaOOjrnERIMZqZk9rKBRVzRnaQ+XXkaQWfosx88DC9fmxKJ5or83ve/6SfEY
N2ZQngzBLOhBfC//K1te8V+qZIOWgxfC+cxrniTCzyHLIhybApLVdcC1kJeDKmnZ
F5yfSco5R+tb4MFXnmetr9S+oYNt3sPkbTZ9lTMDKnitIV1xwQDip17E/eXUihWA
KBxo4esLWIMk1jjy2wNRFDBG5KK182pgMp13h3J1cTrsPzAOKGFLr2UyUr+0UVkv
mum9ibnL6/l6QITrymdYsYNCeuQCheQm1KFxiZPzsewPI32cT8CZT3VVrdoIPGo9
5KbZ9jzLNQNxJktOVDWEsU0vIOCbFJTlrE9Qju5DJHETweT6S9Vdctm5slUmlxJJ
eQo6Tv7vEX6JRR8afrFigxAEow5uFkZV6AL4wD2RwU3TyfhpB/sNgeu6Cxiqkgdn
pHD5+PoyG/UZ4KUDfuuRkxK95RqEZgAhKeduyTrSjv+isGCejYPSCgmrvy5mQwIB
zQnhafjm7Yt9DjRrcrnMjFp9Drk78pFH7eXgNC+Jo1/18TZNUrMyG0waSASy3pvr
Tc6oTUzyTGdq5e8706E3Eqsa+Je5qRFAtzlA3Yq6RSBAQ6IMqeJbLy8qNff3fu5L
6qlgBFoYwfmM7tDiYxmMjWMi/YVpL4tP1VIL/U7JHEmMAYjbOubrJ/2V35wgooIO
aAmG2iQuRwJ6mSyIHkrAVJ+1d/6wtBMrtOQaXVxvz1l+j6kcixyDPWVFboX30KgO
4p3fHwWfX8yypoVzVc8NoGnR7pcCK4wypQwNwn5N8rCo32tioAReItYyGzt0PuSu
Ir5aUZxy2TawwqwR3PEhOtdeRkx9NuTrZ2slaqwIPWXjDUZKmmsVsoXzTNlcOMw5
8vbrpA6gbO5U6JfHWeXyL2vtJCho95vPAzTRxoc7S/ir5puQbJMdb+vhQ7bnbuMk
lsTLO4bywode9EgGo2IXru6kpOHp4YBsoD4/tuq5NYxiByOUehLCir+4+9CYJDIm
a5lFRbpfvJ51C6+xMbLsJXKyX7PEkbsSy/lpr4cXtWp9CQN8bT6NsBeXdoQPQnoo
7nfRpxJCDlF4nDukjgEefc+3zAvWMOFdJHWJr7irJXNvaCW301AO30ZRHNj5tQ12
ZPuQ/J2w9emmXeUYtUdJwQT3OpnivucZVz8U/sKDQIh/TmMw+kgoYCmbRUDs7DPT
efpjLbl3lCg8nMU/q13zYbuK+kURFuqCFerh1fKs7PtJ2Eff/muEpj9pXuIUL0KX
b+KprSd5FKkZXy1WKtvGZhrAkTaUjMfdzdO9eNHaH9mTpPm2ae7TMTYkY1cC7PtO
eunaMT8ZE/KrWfGAxZ8aTOgdV8ShNCrMneZVOKXRoaWLDRJGR4yk1jaKhsmNaYVL
wvJ/SGojSZ86EtXT2g60hWxF6wIGktl5PU4p8GXOTgWcOWffRutGVh4vSRXV0NKU
eMCqpO4JWd0Y9gw6P0DD3MKgtixKReoC3K5mMV0JuRI/7Q5zJpkB+7Ntt717kD1d
C07L8APIRkya7WGMXEk88osNJ5HlIseVLGXO/oMzjwV/ICkMuhe1+/hWTV7rC7zM
cONfH3wP1an0FoFzEl7JCE6NZLE2HwUoNkTrvtpIdylzh09esY1Wh+Sia23LxAKQ
xk/DQ9tqF8NezwDhi/N/nPA2TC9J00yZyN48eMzZZVg3+dn5/ebR4ekndDtZxpkW
fNgciTSSJ7vhqv1aiaRKhulspV/R9BXcs9/EVPPain0iNJQ4YO9y4YlmLznqk9AS
z6Zt/uckWV3t4wEmJRHC/mWm2KcseTCQj8FOKn/p21Qatndn88v4qIut440Lswrx
EqlJj7kAZfrHaiNFypzliUA2dmFHrrpKIVUM+YlJ4FosGqKis8dB9zMF65IJIsCv
tu07z2AZyayqNgLHQXMwMrzffh8gDVVkcW7rce3nKrbY6djwkT2VzsL+kB4fNWMx
dP2mphh/vLF2h/in/QVPLGEE/RukMwFw/oF0bHPKxsLYAxE6f5HhxHVLOEbjJnNm
8q8oCMrwmI0HkHXg7ANpNKy3HtRr5pUfuyStXFczY7PTsmgIvjLn5CBhSV4llY4A
GKlz7+HfJt8xu0D8HpYDf5DNsVuxDg2mqHhCZ86mWZdrLryoj2Ed/frECmr7WZCn
rsa1Ba1kee5YjLyH3HfvZY8fklK/WRWutC+ek8Ht7QJCZbz+9oxahEYaRnhnHgNk
m248R/+0Kmz1gpnXFHL6yuysJr7dvTvrrNb1UKi8d4cSWFOONmqCns0qlDQyty68
Q5OribiP/ALSrEDIbh0Xx6JeHWiR3hU8gY4ao8qp0p8k3ODZdetynI4QHOsJ/gv2
fimXgvPQ5ktVFJgIk2yrfAXeW+MJCczc2yjnBqLiLxaed3Zl6EXnXuqent2E/ujQ
A6Ovx74zREO+YN/Ner2knTyEk2SOQXV5RCcXeqLp5r/PMw3jTrMvEkA6ubJGRxV3
mADFto8sw3zgdsAMiCr7qICdfo9wxtxqPtfKY2rNpkzlODCq28YDJKPHe3Ch8UQG
5ejGQU2KNid7VW4w7uRQ4jQby3QgfZ/18NbGJ8+B8tuNF8cgvMiRAdbNBnlQ8FHY
OWsLh4i6lCQEws/35q8/892ZIkEf9dGDHjiwPfIhedLDGerXLvjPQ7CuqH5iOn0I
20KJRDzvOid6bVoclXvyurcml9oYYzMmuJs+ECIykkMiGtJgBtWgmsodONSR3XvH
Tp6z1R7j/yBsHk/kIW/l0pMq2v4voOTyiHVm3a8xLtaycmPnWDWnx2bVkpiHUQoZ
u2UNnktKhzs0A+mgEDFrZS06bWYImz/thoxGb0vDxt906MJzG34dgdMRrTaxxVsl
lnjy5e3aArDzvdsSiqRXG8GV/M2kLnRZ+zz273QrASF0oAjYoPTQ5UetHlsfU2oQ
RqgnEJKB22k/lu93lgnKjlt7b4F05Q9GVrRausFePnzvyesFIZ0V8IULt0K3B03u
SAVPKtYZY9HKh2u8YQ1SuL1tCEUVXSkVhL+VBxtN83xLOVkyr6tR4NzeTxZ7DqTh
S7nKt11shVRlp/PDQjDV9pEQEWwm7QWTK08mLNIejUe+ZASgXYZs6dCbJjmZmLrt
`protect END_PROTECTED
