`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
614iF/eXAh/Z0ddsz1S4FHPYsDpw9ef2bE7Oi31qWEmtMXG7tUg8tUt2cvQcFhLy
qOS8QHTDhvZgd/EbgqLKqUGg7NLZnYx0eFnM/qCrf67QOTMBaZtr+8taVcY+h8Mn
VT9/7lVTfjFXaE1qHa/nRhaAks/NeVE5DcNCHFF6GZuRdUGdT5bywKyrMm5ym5/g
xqzPBsOYlH7iq5uKyKF8sLUcH4narXM93Xhrop2bLbvV5OxNe5gLugor+U0XWMvf
Te4zE3do896K+QMCkcf7j8R9fqtuYn0nub2sog9E5i1mGyLfeH7segX7pVNfbKp4
j/gcj0Vs58qAk0qGgvzb3RALb+cJZKSSIfsQpAMNUZJu9vNi/4lN7PVzrau5BGr4
NcEe9gdTwGklfHqolH3F0Ch/WKNx7I5ffwp6Vjr4GqDu+0QSQhw3D98RskUPQnxz
kf/Zf4PcLpI8EFWOpLQrAFPCs4f12VjwdalZ5ta5bYxMKqDTkeHY/0F8IKbRhQ2d
otncELVofTk7wj05Wp7r5IlTM1bm6jB/x69u+w32Won/XunY27aE3bCXJntqwt6h
RjZZhOqFSLZJ898c7R8+KqNcTle0WCtMuRVbAjG57xS5gqGwKvIJO4r+f+tGvYz3
VlnGmY65AARSi5YCxBilw8Qe6GobdVWn9PWXQUguSNQqk3vgGoxivT7jdVPNDEAf
DMieKQGjrBuDRMjqlcxOtZ5HvKGdkOBa7N/bufbDrkENl85HsEAJA74QlDubK/Ue
F4UH0GkQHOrbbjdaZof4rmIuhhEaJSF+ZJJ62/lGwuBLCtsRVY825f45CV7cxu/b
/ztHlOHqZHBIN+/W7avP4agdWwx4J4/MdHvjGtphbLedquBFrxvYX24AKj/WhsBd
br+AEfpFUVuEdDwou92C85oGUT7YtMpJ9EOvUY8CL3UqGUoaWdEHJT38HSlVYdtQ
Vr8uBE6CSomR5ldmefbaRkygF1VVSUGSALwJT39Jou9u256LPojbYJnW6iPSds03
s+R2oORDrovjewuI6oq7kKKPyYSX6qUCF5DAttUBPMSnKIOFc8UvF4uZdV0WXzeq
mkNiHjtFGq8JuyZ9ACHRanxXSB/G7kvqQjU980WrTeMoKuHJGpCWQEp8wjtvdv3d
g25hDrlvDYq0Jmcfo77IInFQ6BDpinYGbIQSpV9AGlE1YYrnipBBYIYbxZKjwk0V
vRxnN7axPh6sarRpRuTG3Exy1Cq4VoGol9DArYpI9yMrV0Nsr8wie12biL/1mAPJ
r9vb+KoBQv0J2hWTEu+HucZzSSzpDjVD63D3tK5Pr1ifAmmKk0HDUqk/FN+lgx7v
rCondhaGAJlxdNAdZcuFijODbZycmsu4itRvvWjAqYmXA3QMN7AeInANsc9w3age
8BWodPVHsxpPiXwV957dUGrOI1ZkXALCmd+Db7unaWMCy1rU7Xaq6IxZ+fDA/bmA
x5r7KmrJYGGQeS1cT0X6BQ8+2CzXaoHJ0+JkNduinBO0/Ym+4uZilrk42pJXk0Lp
GcIGp6CoAWaE8pgP7amkmVsPhb1JHhkxu+fQ9QamO21sneMfcIbnrk8eqpa/PVXU
quSiTdbXPPTz3tkxc7NloGhFNfDkA1f6MKIcOMiFgZCcjZKSZW+/QaX7tRKwYBHP
66g9ZIPqEk5Mn92qWTzZ2ZfYROAEv5zgNe0hXWszoVWhbYhpTp7YGjk3mTPaXVCB
B82+yoXZx1j5B/Y7CrhEjfTipEdsZ86HiSujxUgbeJvfE6fw934M3e5aYZn5YOzL
r2j+4Q/Rj5I7kF3hsGyTm994c/tiRi2/hJb68M6S1GDaGZjEApgvb5U0qL3TeN2t
ksUHTccWcgc9/lMMn4sz3/mDZvFW3FLl045NF4ZUgvGrJGwK6M6EFb4y3tCCaxMN
j1gGNLkm96kT8e1Hz7l5W6MdxP3qIHpcbGKXPLGFZ9BzHmM3TST/ctxqSOcFstMc
NuJ24R+n96r2OxGap8q1LmRp3GyTAGwg6C2C5URSgBDgqttQqRo29ocSUgzHYAyz
FnnTwjOPczybPmm1XQWQuauyrQNtLplkyWBsMJN2k9qSCR+cFu40ZtvtGBjMEnsY
4IEBQ7MUmxdFwQ58vhYeBI+7ASSHdb2pfbQx107GrOmI3cFw7JCqlpGPxqZYpQ1q
Te61g2GuZRe21h4wV/dWVwULXMFRt0AKzCl5kH3TcfKBbWa0IUgJRGN4Z/ZtSDe8
WfvKmJNOalG2hQ/iaoKSzM+vilGc9ZT19YTK7PON410=
`protect END_PROTECTED
