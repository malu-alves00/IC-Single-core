`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ezoNxQIiJ14ngGwv9GY548KThvhEgMuGKNpHhfUFvGllI/MSquEiFBR4WIiJ4Q9H
zxvZFvZ3OmAb6qpm2wQYIMc0HQKl8bsv6bKzt+XK5czTfBVSipmVUGO9EXVcn3f9
QYzjGLPyHc4H0TIzViKJfXfABM5Y6/1jzHcubh4raSJABpUQZQtFHbQsrvnYeA6N
9C+qDe4tzC0IfUYmr0NmrkryX/oCFuH0UUHH59lmg9oHV8oSe47sU4heO5V6Uoa+
PLLhDqtm9b4rO3Vtkecds8MYyLAmIJ0FPyUHbEBH0hBXBNY33+DD6Nut7vKhNoDo
J4gpRounok4DfIQyEzB4VyVU2wodQfDLVKVoBpPxQvtk6tuhgWntYRZzVIA9/IHq
lLc42cM4rw9mATI0m4uKlDlojGPWWZs6fjYy4+DWVd0JV8s8q16vwM0cApSeTeHQ
JW60XTYQZywes8KgdLbHcXLtpn7AtHwtxtY0rIWGGpLhYFwOcw2PmrtMJgGNUHx8
ip3lK1pOP/XMYl4G4EWou9TCrVYvGUmFPI+d2wX2dKT4yRMh8keDFowMLhPCeufz
MtiMhDVQAOQVw8vXGx3J2gh+P+UCzSurh3yeKxNF9PcAYKmlgUpQRRrJ6v/Uw4GC
NuX4iRD2U+JpFeF2U5LHJFtM5f66W8cyy+jqueIMOXuUhpJ4HaY4AHrFcUN2YsNQ
u7CO8/VqXfFZ8uefuOfriVLcP826uWTyo5+nBrjFWAogFdefWHcnuuInSvowVRAH
mg/9gKvNxQ4a1+dcvI2gJcVLMjWgPSJIDymhQ2MBtZN/4VamzmjXAJBuyxgyl9LZ
uFY/SHvsRYW9tu2m4mSJgtllVVp2bJ+R8cNp6rsQW8JpZzBTXjhJ6RrmxCl12WRK
f3gDn+VjfNywx13l1N/DbWD+UWdEcND8gf/WYL3bWe+hDKL9Axf5N4CXzFgwTfb1
78K5Po9czcF3lFysFTwX9KZ52SLR08K+bQW5ZPKWHJFJahmceDqYWDYXKLMLRbn9
0vzCCqm36vyLO4RTatyzYLZmoOUsjouyvseTMILTzK0=
`protect END_PROTECTED
