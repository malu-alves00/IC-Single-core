`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uffK4c9ufEOXXHpKh+OHyC+fC1FV/yRYV8DxxO19aDOpc+euJcuI64OYgOAS7keH
2r1Fmhdn/pEqc7AG3GySNuOO4i+dqRtxlcwwtM3bTLp8Y+IfYtkfIsEnNZt0eV1a
Wxp9r867fHGkltvc3/0rweMadwYxm/PA/wpucqYr8OeSxfWNX2BS1uwmzTseuPjD
73QkSUEIGBAqAQ7m/srm6N2RoG9yVR0Py2grJXO3ORYzcUWp09npKDmKQsI3jygK
jgd7+bPZK5LakZObsvem0lSk0geXcqfacY/c/x4X5YH/WOxXpRTFsucZwQm7RPo3
xhAzoPQ+cLklbaN/FsQkKyTYyUF7wphjTvxSCeNiPfzsK2UxNDslz87sNEsdgu1R
jpoq+rb714GEN2pgYKEqmqFf2krC7zc0a/n/doahPaYZo7B46n4MGScCJNb/kjlp
Zf3IU57KEepBK25LAPsKSgWrh4koSQXx29cg+bFoSYnvauY1yUHDV6aLdQ66wHOu
DINP+Fmq2CssHnOkuNvnB60lW+xijH5bMBdLDrWc3gmYhkjV7ZNLp9lTkEc1STIb
HlEfYfRB2LBko3sAIGj/i38vljtEPf0hBcazRXxBDd79bd7ClNwvIjYL7kr2c6Vp
u4lA0pXD9dOSW29jMZeHaaFOviHEGqVb4f1FpD2XeDAYiEwgcVxWnrMGUlVi1z6n
twXkEhIjU5oPj9CX3KsqP2nYy+OF+dN/JfvDxucGGSm3ct/bkVA5N8mNONlkZ+Zc
eX/JPRQNiRbiuRO2BMBd1k9wTXTtnCpLhJjpX+dYzrYKi+mIBJsux96eCB3uj0qE
EXRLhGTpwXa2VlXkTIfB590UHqssVJY1NcCGrfbpU0j9HunT++7jplhYcZ8Tvi28
2a/AhiM/MItjdVQ7okPXf90KZ4hdKR/w6LNywwsOJUgCbo8btaU4Zt9M4jKA9SzM
YLq8yiOlw+OtNIs4duVkl/2ubcN26T4cRuvS167B/Q23Yk7K1MN+blUk6geoXbcR
k5ljHeoYNrgwAG7lnvbfevq4ZHEWM62a5mDs8KjKp6EJ9cH4j7r6K8/aO9LIU342
+mL1MbmKRpnfGaCZifzJYFrUCI+mk9D0T9dpj4qS/uq2ID7uJPAjOF/UnBltQWeB
5WiI/vIT2q2kwfC2IWWMcnqx4ooUBqdkMahJyol6XROew7HUqynYMWzIYT/KTdOp
1mmHxag/xProeClnRiBE4cRMs7Vq1nwqiNFvuDNQAPrcJUjizVrBmxHi6h3/mJNA
AdttPFu3z8iH0rPg2FEmcC79U0FxzRE6vRjNyDRn7oK9jkESM9PVGnNf8kYracNX
fpAPfJR7cE0I9UUkoy1OlVEYwsNqvJ1tmhJGWh1lFFvcabDPtp2QWmqvT+n15Gk3
VEIt/Vt94iAhAqzmoclsCbrC6O9XAE47P7y6OaZofiSsvTkIvOYieQVA1rPUEYv3
SNhj0/S7JERAL4vr7BMhnzVylXgx0pzLTp5NboP+s6Zsifb3SG1UFRM6jy6eHm6j
tVpqJ/pxXv/DFuovLCpIuhpoGEhCG/Uz8XvoX9SvNuGLcjUPBjItp+ZPT++3W5jG
TydlgYmpFlcOhvfRE+Yo2rMx3ajCOmGfaI4t/+a9MKU8baHvbi3TjPsCNSen5o4Z
nST/DNGo68ahHbcZsiXbyhNd/r33OXj/Az1MjC3nYTj191SMmzB+zv1ymZ89upWS
spRvU5QGnrHvQiJu4mKsyTQVNl9DMfuYl2qMYxkHKU9NLVT4gLVdDq5XmUsSbLJB
dEvymIGcwEyQEljCizH+lhERhnoj3Xs449gFBlu8rSHfx3kqukzUUz6g94wr/WOF
VJ0PoRT45vq37xiEB1JJEN6s7V0ugU2hnD/WN/XtPMASZwJmkrzciMDGxd1QxxiH
MXWZfN7IiQZaB38395JzWPt8o76GJOxHIJB+xnx35wz6vV574XlBEpJebc87KexE
61nqdKfqyD+SPvqxEdlPF4pf1G+zO5YirMbVefvyQuM=
`protect END_PROTECTED
