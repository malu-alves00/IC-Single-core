`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ztTEutHMvpF/DPc9hK864WIk3K/jNgRgpn5MJB8hfhSpZiI8wngTBlpYPzrV8K86
BYlNDJq3rlRp5SQ3bojFB63l1v03FCawe8aFuWd/p8wEKCtA0Es7hkkic/qRbHko
LX+arUhdk7HQvW5LBbRIelI0UvTRlMMRQVdsETxdI4IdGKX7op4O/vdU7UkxU+vH
zUXILvWQRRCQHq89lXGYRurolJHcByOtOR9gVOm9AW/2eXbkVTl9fQp+6dYwjmI5
wJPtqswaLmPEmajOjrzEMIPw3bBzgo1iNo1BR3N/XIAmQQBiO34otzSQ1i0N77mv
82phh9AHznRwHVHGKnXFXzBhux0/f7Z1WOyFulSazsoe1Kmb9pv9eHxvN97TZwep
yOsTmeA1Sxa9gB4s6jOvZevE405v6vWrdazZ+7KnydzQVtpMXUTK9iISxC8ROtye
c5N7Pt5XCn73nf2zdHFwOIMHAv5bEy56l/9sm6aGSrwSSfbxMV471sda2TnBMtI6
bhi3hxd6iY4ulXW+uI+tlGnN1uT7QM0K938CuC/7D2/Xv5BeJdYgw5TdeomCFMdY
4z3LV+d1UUB2xlT2HRA5Tj0U4XwJPfjPDNQMIxTICvxkj4JVQv0faxe3VNzXluvB
ZXlXUrsGn2Tesx9nBupctRAuigiEMU3y5D9YPf1gbi9npFVzVFnnmO4NFnPUi8RE
ZfU5D9HyOwdkk5hggihvA5BkM7yRlCX8IIEbDc6zKgbSpxF70CmiEQplGe7RRid9
4OHDMxITy85tGTOLbV3NuHYxtYmBESKVEuZip03GJIBYX+76lt8HRiP1WjZgtJsN
6vGSEjloojZy97Gzk8S71TVRyiBBdI4O4/8NA3KvnDiOVLAFdRBD6BKJOklzBFcY
ILEOEAy7Zig7v0riTpx3Gd+9hLCbv4WJJddUaGANChhubtas59YEjDo0T0l/xoxI
EtAHUXqGL/sllYgNDDhdkAm4EKEWf2A0hGm03hiYLwUuqpwWp11sk55PnhQ7bSwz
Z//wD6r2Yi+jaDOjkpgtNY45arMsbiSuAHxSFIpafGVAWjjF+fjIh8BUhNhLWD4z
NtAECWstEOwhmyJ8kA+l+nxqQfLMV7FRcdLhPZv/3NaAd5zeAbab+w7sgeJ7DNOd
7Me6xe4x1VyAiI8EjGybxnJUemRKx3JSatM1qcaI7eYYel2OXjzikTw6vEB4Q3Do
kg+Wvc5gcn7IjNgJEfqqiU1tj+lk+QbrXOI+B2hCIa2bIB3S1MP9fKHroVzn/46z
n8PK5qwcVs++0C/vkV1QAdX0UFBy8EtMg4t5JdldI8oHP06L4iNc6YebGamTqRZi
tNrujrXtL1KtpxQDKE7748atb8tjVbI5PHVkyqCe2YAKxBfCzEDg0mO1MD1CYTxF
yFr7ZmxIvMguMjGA7W4PqzN9VGuFJfqs3/k1K1NZE3dDQtjww7RkiQi99wq8dQFp
wYf/Lhz8KOqIE115R3MB0yYzV2UmmAvKS/0PWdDdu5GHNKW/rtNF8dbngzpaqO6D
OzgpJxjRPIwXaX5qT7yG8ZYbIhXIFDcBh7YecIu8UKSxDGGLiCSKXbdLPlOmmqlV
6Zb8n5L2oSFWZMuderZQyMtMgY3+blbuwfQcY0CE5+HIONH+MExdCLWr885utHhI
oADed9auMuvA10SiLMSzbpU0FfEwyzZJI0n4WPDi2p2GcKkhcyDJ+2FHtJSetjGo
LuUKIWXCb6aBfBKgzsHpO2gZYuJ6Uwq90bAzSZPUJqdRe5eSfqWSErW9H0AZl0OZ
nPrGOmotoCxCbobNNKkREKMifM9vrN+z3ri60YNRwTMRgNDg89drQ3knFBmtTgR8
4tENmmym6Gt6GtWLeVgzoER7NE0P001hLM7chTfUowoS68yc2RFh4xA4JBDHtL63
g5xFzzlJgFb4PdvsNKGfTTCQ260NvpG2K/6pSepWcdLCrJwHENa7jHzn8NPg0P3k
Ub8n8BecsNBY2WrS0ipCBxiA6d2JS7YFWRomdtpnnbPleuMsFgvbtlqBaXCvzW7m
eoMe82gagoAjdZeDKgF3iNmDcWcTq6e+ZTWaW8wPLroWqAkDH2JmaB2jGNCl0w1Z
zOnUzcSgEXHCuwZWUn0o577LiSit99TlYWsK7YgLbvdpKyEolZx8F7ev74fFveIC
aHhpxNTbwbniBHYh7VIXBQjci82hLdMreFxAbPPRQ3dvv2NaVyRy8PwAuwQUssFB
VVSyJVtAHSznTuNZkrDK/ZYoYe63Peb/G6AXQodB/WNeoEVvriLSvnBveaAt7qHb
WojN1M1lcduf1vGUETz/1PCBkMeh7s3uU1K7F0diQgzNk7ddpfOBAbTcvR30WiMZ
u4DPcXPC/TA9DRI41uZX1kFRxo6H90ZJChSUZw9ImdbF+lnDpOMt2KE1MQcrHl4S
`protect END_PROTECTED
