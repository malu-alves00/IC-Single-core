`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xNpfRFxMDGfJbz97TDslVby3WpFByBokpy00evhbycHwguLeuZeMBal2jdigB43B
LnfWeP+y9rwpt58w8oYJ0uqzJSBbaT9kaNWNh4jcnTqUhMHOiThGd6EtEdGysz5V
yEGUk0vw7A7oIH94Dcjay4FbnDMT83bF2OSXRSLpyCwxJ+sApy4fMwFkiWzGlgfq
hZAWWcpRWwdmTMfpHl3V5zoPEKklT9cdINf1ufUG4nvLxRHnzsECglV79qn3+4/a
qdLhza9Iz+U8N+v4MTP5aVfAFFocZvuqtU1M+MeMpK35h317en+mnzunCVryr7vA
0DGeHRQsxyRpExKrLlk6zVPEryvWMWbVo7bCbR8QZKBOS/ohm3SDAoBbLYN2Gz9r
B7uKqmYTbYPmizOVsFYPnWDjL1n3MApJmovdI1LrZI2md0Ym3x6SN0iy85nNUDJ+
aymj0bi9Mr9RixeevOgot0mDmqjmnspX0TmotfLvo8e64j8VgJbs/QTxSLDDr0rz
ouHvsYdhLXfHDUhPlaf8ADt0Icg8ywHk3FKr8fT6LtW7yyJ0Exe6Zu9SX+JZ1IxH
gFKGtoIC2C8UdWBI9R78diQhTquhpmu2YnpKkKyEnO7EKXgSAd5zKYOcGSt0T3IH
RRFd4dDkb+pnsca7aw8sqbJsqZf5q+rDesulDxDO+Z3my/OxqQRF42/1qesqBPM3
JfSKARdPiCOJG2byeRFD05X+A6QLbnfdaw25NB/45vashSGpfrWTtigWQw2EzJjf
+gOkTJV1Y/pcS0nMFNkOQhnvmJqRbNtpC65pxu7U4vty27E2darJdDJlyPBKosCv
CypfCyUgOIVIR7OPJfWZP9EeI8zzFofaFrdSXOG9ieVdZGGASHqvXVaF982lp3Po
Ig44YresCpVSiyuMV81r3MYsn5L7MFU4eFjwYaRQJAEfHye6yCxkIBN/A+83m6DM
GajulMKA9iiRVwyitJUBqbc3Cpd69u4JRSvYVgmRhEAhBV4O6j8wp1ETwGqIt/oE
jEO32jyIU0i6kyckW87GpiPzzFn+XUIADsaHw218WjvAk7TQkQ+mrrD9WfO/vXd/
kbUnnpSo0znKcP/l6BuapQqWztWx2iug6oIjkpKLX7F40FF73Q2pUJMaMkicgp7u
m6KQcs6adwx5ZsSuc6ZZapcXfwEScI/+Mk69sRH0mddx0Xb6lNyDS4CNcbIwEtTI
V1AkvW7cCkYretFbIg3JGO/vgveH4VftvYBkh1grOqEYVkIDgsWxz+deeecRrI9e
1ZhGcDWCgiTPsPR6Se6KIAiIOb2BRUsVpw6LQUs8kPPxRoTBH2iXkBAaHw9xLvGn
v7hgo2iTAUW8ZhoKXyz+6jqVCETGUSsoedjgpmXdYlTQVaI+10+hEt12+3YIAAnr
LagcdbfZE757zR6FVs1d0iuJis2B9bt6x3oWDeXa6j0nlGZKYLSWK3wQUIygTLty
iR3PFzYao0BxBtYYSbs3aMd/dHZYlNGQbtIuKKHeoTM/u7IKUS+GfmhpBnLD3NNs
/N1u8uqZskrogWgl4JTP+tc/UnYvN2Ladjl6djWIjGOL/TfCKDGMb2I36BWBpb2V
UsB4jxq8OkLAybrQ6mtEePQ74o87W2VN7DISr+sH+cGfZ+K1vgxEYlilyp59hXLt
288JC8KJk30fVILI6mYSP3emTmMtuSMkOI+4p8aqGk0TKV6nA44j9etBpJqA40/4
+BZAStEzEEVVO5NU5qdkSxvXO10L2ZhaMkISqgfl9U8bX6M5srqnN/8fL0dSMhhF
owLY/Tfs+lx6KoPfu3PGstiVqgsmvHvP8d/vTlzvb6DC4jyjuLtZC9RP/k4CTqEE
sdAver4gjW2Pn/KQk20KteJSXk7dAW0yQDoB0/3kEiwl+jdBHSh38+tcBVrlpxcs
P6ecGj0LnbDMCof7gjBRGI1ADnrgQcEdL/Co6XNqlqbJoiQdERlVdHvy0vOXJyLL
raq1pZfXBiYgtROgPIl+k96GVw93ouV/sMynSWLqjMjDXvffRi1cekKI5MmjgM4f
fb2wo7rROGfVKacJ/BQnYzWChbtNp8ah4N4JkI3YWrvrFiuCJ7P0FwrZ5HKuIT3q
hDO5Ul1GpWCT55b611DY9Poay4G+NAz/xikbbQOT+17OBNzerwJz8ds7bFUz8msu
l3k/f66hnN3XPbT0VYQ+rcZXMhptAmNKYTGUFeXTZvK5QBffqTdp1uA6XstuYCrN
iYMU9CnXI390GFVkZ25Vb5maOH93g1d5WL8gftesXD7TJqpaW/XxDtYStpCgP+c6
sblCD8nFhdFlhy7KHpcWBHO5srJdMRg/inQ+wPPTqBV4YFuEgAk8y3W34rirw9GY
V/etx+cKUX0uNBhZUlwZY3BUX7hQ6xPKKGwHk57gjxCV+LCyMvZZZQg4WfWC5Xu1
gaT80UStb1HfKhwBfBsUPuAYjSe15GF99JTRsMf1NPGVtMPdL/09R32oJiPmKgFH
LXBrm+Wlr0JqfjmPgnkVxegvVb6QfSlXCumP+2MSm06HryUXRKWXk5X6kax3QnRf
prtNPaTiSv6YBUHVIGHPfldOwZ4txmiz0zG5quTmMe/SAxc3LKo4lTetcfQupMq3
39D6+aM6u7PRBLrLe+NG5AyXMInzFhj8hZlh8Zl5BPr1ZMjw7T5sBNJZZVYtmiBC
tywhdynAAh/YWdU+Fagm5qMaFf3030T07trXrbQ2cqySd/GctHoOs2mAAucHj5Gf
+q+OS9gqvLgsZRl9us10hsY5gch8ic8FiFf05cGj0mUwaPLL9I4NYMfD3YTO/L1o
TUd61KkUJCypUR9/YfFqenuk+OCTjyjrkOSSJ1JC4RIofSeO5u26z6n3u/kwyJee
j2JB/+9g8t1W7nCy9G1PTR0Vt0LPxR6z2S1t+ceUdKP1UcUXO+zfqvqmwUm3Qcgd
IYA6XQILq4OrHNOVvWiuNuztH4l5LIHI6JJIBdZxMX0RUXcr0iz97Kz+MO1iWdyj
Qmp0MGOKmtu/LmYZ8/fTGX8pa6qBtdRXTMhaayUJXE4xXhU1lXH20/u122hrNNR4
sqUvc/XJbqRGvdTx9gPl7AqHzd0wh2khGIi4UtyoMFmTNcM6NsnrEL7gP3946pNl
lHA/QVSHIqOwA9RLbBlRdkgJeJwVXMwhMolB+yPCtqQ2EA0A9eVhlSIfayZABy+q
gRr4NRiCajvSF7ZHX/30foGeUoBUZ7j7DV08HEqTeUaNwFnFX7Lfk6I+6G6jHXhK
gYnKr2awLJpHZFnL7oYA2UxiIAr/W5DuVfnYA494H4OohA3BJYJN1HiPdUZS++5k
xjoagSjcVo4TxGPvpC5gAbMJd7g/M9zBz5KYZ2A1J6xbiPrDDDd1SycepbG0TuI+
MU7AxFQPkeeLiveyEWLJwmEtHQOqzq2TlqGQDrxL4u6t+Lp6/PuPkDSBkw/iiZeB
D3r5HuTniGC/PW9qhT0aq/NXArWImq7opz6YmvX15fVv+TP0Xkr/PN/SC1wUtznC
sNyB4U3nAOcjLGmZdsLKmssN4kFFj0//noStHiX/xpjQoziAFSmNgI82Tg38s7l7
eqbpxyA5cVp0Vk3ivoGyJuxrFkx5GIkAQiE/PgMH0RdrFfqSh5KKnlfqYCb12axK
t4zaKLdXyFFXdOqI+w4pEWmEKqb+B4MGs57NSQYU6mfVCEDTTTJBObJRpcGCr5Tv
w74cSHMd/WUS0pEMWfTeI87Esbf7xIRDnoxwOAygVLap5oVKsKcJmZ6RFLAeJBCp
MrG7CPWTbP2k7KbxwWDGJ1AZAPG12+O3AsMBMqZ1Ltfuj4iI3ow1VQYkRgJ+6mMd
mjcHcJTgHX/SJpLQ9ItpAKGjFJXuqZf//cLNIt+656n537GsLYl6jfUC8b99wrcL
VKiA+8xt0J4ibSUdW2XHSO5UU9qNtCmK1b2QxSRb7qmPzrmM6e3Aq2DRUTgZRoul
zwlb9kmF6BRykFyHq/qrvpAM915s7pqrya0P3ReMrrADewIKJS2WR6kF8GbDOGsS
vIbA7UwxS1ztBEpIYjQxGn3LGF6noSEVBODVm6NAv/QgTdGHehp3i9pR+gDJZIOU
tIexIM8AIPZ8MJ54NFHrsF5oZOAE1ZG0AU+XwXoCys1wbMPPSWxr9cMsXJfQ/59o
TxiFEXNdGxueu9hjMfuXl/tyWBoeed4J1yBYM9JhCcj1V97eNjBTClk/DPsXRtp6
fdvMCD8NQ5CtBnt1CnNQRQeZa48eDcmFt7IWve0126BENnKjny3ZqwyPI47J7hQR
8fFBtVCxwvx99nLJZ4J5efTDKjfkgG1/zIgNxbbbCatXQTKFcPJJiRiXkwLLE3kB
YVDLR84sErACU2TdMNv0pFbl6pkctcy6ALgvpOYx4TQPBECWDWzsemHKXzHqC4A5
/DcEuBGcMkKPVxJ3CMhP0Hv+rShV6aiHosA04I1rn3ixZppDps0NMsbg4StgBleI
amyarmvpIeW040NBjE62SnCnwjJkeXetkWX4aZ4zl2PN4SNy0b96lImscozipO2x
/h0wgOxhKqQOEcWML0Wv1W1DnsKLuzlQmT0vCncIXmw0GaaSLY24Hzl7kMcpRpiq
EnUU4i6oldipu4BxzfA2J0tI3GhrV4WgOFsjw+aNmSAnoOBeU4YCEJV3U3hO/WVH
eOg4ic+m1VXEOWk/TKeIR50roIY8AHW9751/UG9XyMIjIL17wDbdb/ghWyvuGbge
Yqh8PdmBsbwYp7vIzQeniJgGl3pl3dKnYzO/tNHNhHucPBPnmTCe/mV+/sQ8PCnl
EsXr06oCUqyuwfjfxDo3c6UbwDJjMqersXcx8sd2mQVWxQSCt2t9May+R7MIx1XQ
ZqAcQarO8OFDVWyIM+f5K5IIHgEAfu+ZxMWwIeYsUV0Vogkr9dqqjKd89HKJmTCJ
nhHKEh2u7yPJ+dUeFbwSICMt6Vw7fPBYr0PA4RubOK+FCRSqfYk0WY/q3XctzMIl
n2st5Ac+v3aMdl41oS8pnEfLy9mxsm+He/rRLQecW5QahNsm2Pzgm8Ddd9oPzSgx
Ab1WP5BLPK7T08tlmn3MAeDdSOquIiJ0+YKtS7NvOqC3jR47ZKDhjaWt9O99Z2+t
+XS/zvlh1Il3L2GThwDyfU52D6IgIsio7DDQ7WelADA/4D/7LRePnJSytgs2cpCj
tHPiNcAAnj2IFcfC+KUcw7fgoAGPtr8OqCR/BxNc9sQEcgIr/QBteasj139omIcW
efpEKnU+IcSXsgidZRUhleMDttYDOkzWN9wjLURx1C9jDre9f+5PBqc9jfEmOW0m
EFq/6BNrkDx8M8eNmqQrh0g928oPAMfZKsZ0jUXalbEG3czPrg20DUi+7Nfa/fkV
iaw5vr0mZdAlvlyC7uDsVUziY6HtiastQar2YEZp+feYl/OISTCjP/sR8q9RER/r
1YVABSFVz78vxrM9+oVKlE3JEk7qW/lKg5dCvy/KRE87zSEEphbc77miFYWXwx9W
zORdq8HMqk5h8Vpmv3jNlpWpnz3D0hRmnjG28WUSvDo8FutUpiOGq9iF1nPZrzqh
clbsrRKMSmCqdGWcFCkOIDrk0mN6yAYDdsHp5iwkUz0DWReAe0sG2J1wBuoLSNGn
vddBlmk8aoYBV4DKRxom+iPathVt7nRYMCEjlobGnJ8RtKPGnLJmx3WnG8cFd0wQ
Rl+pH8deOGcgiE6uHXF+yYJsexEOx96D4pyBbTJWcR+HbfSnhRNO0IRT5KT4pHd+
tjtf7EFmemlFuiWXf7v1Pqk3dOlBpqj0qNazbwg/W5qdGn07yswxcaaDZbDJ7SWj
eDWayOIVYofY843gnfyYlmFIZi5GHemZaWjtIdiNybbk3gsRFmnDBXU+dfkU8Y0H
/ptsDvUm3AeSYxNR0LBHlR5Gb/9+FynUKVhd/tjn2yG0FXM40uNR7voJObgDfBT8
necRz/o2+3qfKut8pP8ZFah4hTQq2Cv7XcX9Iq+1slzNmd7gyteKSg8JGHU37TT/
ViQiy6AQ2jy0exGHwtUDIT7Y8wxk++lPZbxyRrA0Jhr8/0lc+zvYLQtDUtry31/B
+zWnJExAXVlCF4MoZ4QL4hrMMfjIdEhMFV8EgiraTVZTZYvc/DbsTDV1ZrATWmDy
7KSBCDQE5PZlfq1FlzP83NebkbIA/mCBqUUEtUO3/sWj+30OQeOCo2qlfBxfLhNw
k634IfxmCKpx93iaUeseyafSfSy+05AmKtTBy2NkyG6JLmeqR8zqIIUoss9OfqqV
RfIoevHQhyjTXpqsKz1K5jwX+ZCfywJP0DUQS+I7i5oCY+uVkElE+64aBqXJ1sNz
aCWlSW8SxCiSK5hiRDDdYFFYuYpCZ9Sr/fg+hKStF/BHgkd5C7J4CNMGqosaAuhQ
RkwQIX0Hnl1GA8a9muPaMdwQA65pboftQNBjygY9n/8xIwvxQntnkvBrYoA5HvuV
66kaUj768lJTEF4OY1BE53+BWaxnfwLq4Lpb2f2m7bprc8/jgWTaR1tk8g+m0VBl
2NpyE1FjxDczGQM7M1R8z95/zPMlVAYGkpT/Pqa9BLeBomMCr7raPe69lXXW0caa
i1C+W96KTeRYw41BHolnbd4kK+kCUFLYMUll8HSdQpLPLkSTIJdfXxNgBBtuXcGR
pFnw/pmdWBB2ktuTmBQriBLl1agkPly3buy9OIBJ1x2lWuxzC+OusPnG0uoO7NNP
19C5qXAj3DY/zqpyJf9+ygVJ9rOh/E53180dF+183ggkd3en8QP13upiYIKdHTBG
O7OaWc4xMznTej6w92T+oD2BK6H4FIh93CF916+HmqDizYyi9QTS56LRGxJ8KzWT
Cqnb/6URQ1rrBbtX8dGIBkh0uNoKBCbQbTGEI39B5ibyPl+xnZ4aXMaHFvKYz6P4
RUwG5WBNbpvyHGln8o89qnzYK+O5RMugxwI2B4xyjRW3fjEc8aeBt9YhaR7eQFx7
gNKP7mzz4QQDjeeGOwCRJbK2QyO20FScvpABgellaUjtkOyFwkgUCua89q+Rqb/J
oofl7V0OyRgpdmYBCVGBdSmmQmBKHXwj+xVXNIgfMTi9CCZP//0ict5G8J639XrZ
h8kKqXT2NfNDQ+n7+BBMmiU9cOueptrLBSr0h4ukzu3UtOB32uVIOKf3DrMBEUkt
fNlH1J1dGg7Qw8xqvRo70IdgiqyhiJvpgeI3mqE6ym1KWaeDgmnXNlhEKi2oYMaG
okYutAG7H846EfNk+CvFa1HaAOKeyva8K3Getscmy8XrwoL490/QfSxFcdL+uWfr
m/NYv0qgwBHsMAkXYBuL/VC9XypbjJjp42ZNMVQBpoYNjLrT7eYz8OsAULTIHo1X
3xq01ifWGTBhvh7Z83Yw/u+diCPIi5EvahU1Dk2Ge/G6E3xlxXHT1eEfA3ZdMWAs
po9LPH6DbyfG33MjoIQb/qyaiQTFoFrTqfDazsKucUGJtGfkvtbVFOuq1NHbcjvb
o3YwJwVxZEFQD/F/ji4mYGgJmsAtuR6P3BnWE05zUVDIN3blDmxhXypUlz/OLQ0H
JrU2DMqlav9p2fxeDzdtvb+vSnHtuVg2WUF1TuYVoA/i3Iuxp6LsZMc7iNfHQIOs
/2hANF7Z9M8PddohjU96XfMRZbBgTArr8SRJfbIhE2r7rhFm4/Q+/8FvohvJMd7O
NsOtGBI+CrbRd68c37KtXd4ZgjXVo1RSt6WZeFb8qtVw9iYNX2vNHUHdDcwAQ12b
Wa80z9zeWhENQYP8nS7/RwAJKgufKWPR5e4zE9mYzKs=
`protect END_PROTECTED
