`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zXQ0mRIWS9xqxhjzIUe3RkgGXe+H9tDamEWoVDT3MYEcQqmkbXO9WP1YCUAxp2fb
cqXsz3lwTJDC+Fsc9+rJoOiXsmREfxIz01jspUAhWXHyv42LejIbVrgLTWdmaKXb
4nd2dE4boradrmYbwoQJl993fIYjnM/wxcoK1+vzSYNQIFVLs431j33zjqmtzo50
arHnvZJbygc48zWrsw/H5kqFQdJw0hve2+SBNNk8ZcXBmBQ1Ij/5DdJxqIPoLwSu
AA9ffAzeUg2Oxrx+ia6VutPKdMVIIJWrJ27AZ4V+TPV4XR0AszniHD7OPuUXpR5a
XDLCP8HsMZUVWiHvibkecZ4wLHYJEbFJXuzsPMBGLHTByo32zeJ1ynlyjlMw0TKS
ZHH9WMzFPcJpeY5YUSVr+VTR8WMFNTw1J602zeKJC/FvKMLHc101ZBylUoJUl27X
C5qVW6GBhfSF+ul0OhMwBCtykLY6mQJQLJ9sjJ0xUIQ2U4g2KBDf/1aic3bjjEVh
M+AsVrU3/KSzBPaP7DjjDDEjINigzGFnjUUZWTPEkow44+1C4DucmCJNgQgxA+fW
El9ANn45NmrGBfvxGKYPWngxq/VzI0ePRyYgTgjsqgvbXvZIyyGv6qHs6wkY0hIq
UQLx7etXUovQnaFyWcXIB6aD4wnkad6W74f+NSkFNumuAo0ji0PHnmGuZCXZZ0Tk
9rHeCgJBEofxKebDKa1wRyCLYEeZL18VA5uPFQB6J0nksP2l8YfYAK0Qlh9Ue+X4
bkjrSw7GtkHipYWx/PoJqvGmRP6OYw7kc38VyrwoTkF/PH708RyvOW0kBFhCngsP
v0B+pN5f8JnXNInoAZlqEADsVDIYglUaP1b2A/4ULXiAd+EyGCalnc6TN0nd5FcC
ZqNlWqSFgCApBk9K9CqHapZ7IlnFhhUa0IxZQK2Qb05wFLvP5RvtdCdRXVy2Y4mV
2kBXHMWJOga2lbSqCbFfoVUGHCs7fB0675qVa8jvk3tjQ/YRNZS2WJa6+Zwzg/u1
+0GEn6LDdSoiUzTXwvE1vveUDC662kWFK4EqajL+q+Kbej45Q5RyvPWQibqG52JN
nWNrO8WwX1ThM6cQWa3YEPEpqDNrQb9P9H+gZsAjj9MzOVAHS6oQSrD6VNn41Nm+
eQ3oBI04a+cbkGbiLQpudbq91Rs4AwJoagFYvt1//sxd0AVKLm7PkuUMOk31Goi6
wr853QRZ2t6iw4SWcrBqxWdnUyuh/RfNqRnZ1XMMBOF2JJbAlq+4h0qbOj3mupm4
XqVgLcdNT4/zYmjsNcKePuJhyF7uX2UaoiS3MUG/EaHHkdwJLxZCFnCwsnTQFIg/
jd1ctSXAp7l+YpZgPJWnejkPhdz3TI9lHEKBU+Noh/LcJB7bLzu95XaGEp6qlcUW
/hrcg2bvYLcApUPxk7Abdjym8uWuNCTQ7tg0xQT9/Yg9A/+jBR6x76Otc/97h4CO
VbYZxGcbfbqIzQ1iEHZVEiNGHmEaLRsYnJVhEbesZG8l3tc7dlkePoDJOD6/FsvQ
fU2hNihk60ubxcUhMDWgzk0c7R9QjRBqGE/i0iM6TbSrMZ4x9NZtJamAwXDkUULV
1/eI4P21MjKbSpVsIHXbNZQveGxP1nXJdZu/fbov/hpTcqYTbCI1E1cv7Fa3/jEj
Ldk1mUSU3te3lNn1QzTX42vLaWiaWwWIfhwZt3jfcvaWCKuQZwdaq1MXSz+QBF/T
K2UsrFYhxsnD5k6tGkiehLuQ6n7SisOnv8U2tJufADYBVaCB9Vx0kPTgTtszQEyW
2vuFuSld6RZCXU55gfO6oS6RMfsN3rZfu4MDIk8h7hq5dcTRFWolVgW47ghLt/Sa
yZLlytIgg066PIOiHuJcjFdFdp4NWWQ/KtYqOvTb+TfGd6XnT6khX+/QIsQzb3Ak
Ya2ep2VtOYzIpwzF5Dab7wuWE49WKGZ07qJjPouPmVnBOaL9Qj0A3SMzpSbYxaWO
7fNjMmGXPpLMNaCZb0bibXCkKqxIrODsOmQ5fBvAeU9imSfcJA+xQLkumqbR0XdT
iOjVc21cCebfocAxwJtMGxKxcc8flu2lPhI0bhAYxwvw9fWfvH4TIAARV0A9JVka
NN/KqLzKwCk4rBgsgdsmJbAT3xZK6X+2cIHG82R3OkJuF2+L3LRxF4EzgKk3NVx0
OT6za+fPAy4fDw5aN4yhSW1R4pjNrXfqKE+ojrfZmP7mtTJ5/60ABDVxfQ/c3Ik6
lzVAf5xgJd6zCFvt5DzniOZiThQG8SPy+3nZQgODYAd7dSxSLE6vxGBY7v3fVsUO
b5XkItScJsmslrgggFzZ0dRvNgn4VZZzrM0Q4pa00r7EP/xXzLoYLEQQEGA8RvOi
VZUDgGIRu9TrfYlmvhHEhJLPUV0S0JAvgYZoZhgIO4JgaDmjOMI5eqc7ykoOmfGj
`protect END_PROTECTED
