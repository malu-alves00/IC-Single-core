`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XqyhdIPTTdC+gz0dFHZCDdhDJp2dq8vWj/7Pr8rvMTPzhnFVJ4abBjLe74hIvCob
11vAi6cYTVSvcJB6C5cXOFnTwyl6KlfmXr9D2KzgMhv6LGy+Yqq42mLP47VBDZxc
So1h8xzqjQFvuQuxaWfTgI9N8IRPrqT1z467NlSn12gdrtem6C+cYK38zwpQXBQF
MUw+t7HhRaqHXfRqy9Lo5rpmDUryqRSw0rm1pXVR1CGVHanit/SCITbYs+VdOI0q
az/lOdkHAO9MhvC9B9TZpEEoJUN8Cd8JpXxg5XVn2jECeBz84EeA/ELk8DV4EG78
jE0KyUHaz5ZzKQjcBkOYV+8vsQ0HZfz6wab1MczPlln+XCrled5r4r26cG/JsM3S
dt4EW/MXM886spY5B8/0XpH7pMReucHxsrwBMYdkCCYtVu9/gJQ+oiPiRjUhUDUU
+Q+SjZFlgiu2iqPxGQuq4VWgjMQHA1EQg4DWGedA8d0=
`protect END_PROTECTED
