`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AW+PEcQrnOga91l9m97q/U0XGhg6PeiX4D6N9BJHM+YOKVVkithKOXiaUvenpoV9
y6pv+oue5B9m1P5KU8qrjNevYW4ejSE4WXae9awNUKmUUFq6ztJAG7gnJSuQGW+3
XM87OPNjxcnxWL6LQ/Q9pQyiGS3DoJfMQZceky/KiixTfbLY3c7hVTeWhvffXa30
Ot6Qpv3k0OujiylRpovM9uo4GiemQ0lWlF8mz21BxuRtQLkbdgcWvg79e1JOR755
qCUS7w87cZnO510n3J6pZw+D2eOf98j3tQ+WZHBXyYQYx7vgvusfJSQQpzC7oy9Q
JPinqTOucr8pH4ANs4HpC0BK8hrHtZ+IYqzwD8BGru81s/L7bhWm2jzfTUIFk+8z
qub/P2IZaDOLKhP2675HtiKShUdypFo4JWYJwaAugNUIprhutftU9Ff7E3mkxe+E
FJgXepWoVRbGRD/R1WBInEHXW3IkPDaIjdAC5aalQ+pLBgHgh8jZ31BzoxXWf4BO
k6gsYqrtEtSpGtpqeSkYSPAIKIwKU2ZYGweYN8vNxL46a8yLtqDiMkNTMjkdEHQx
HvPM/bGblVNtMhfJFlZSiKTVgj77zlVFcpnSZN+DgM6CslqZ1DU6OnhR5wXk0KHA
Plhbn8ZeyWyWHZpznnamUIzoEF8xx1BaySSBwj3xj+6XAH9uOkvteS2Iwd6Bi4xB
1Pv47T+3XypP6DyMnvAmh0v2s5ie1KgJaXiwmnMYrqWUgXQvnrsCpM6Zb+9XPvY9
6QotNTZk9hZHmD530AT59b/TmY5c9TRRRcQc0ietMC2n8/9b+lof6UDD4CJF1Ffc
egXNiH2Bl89tr6R4c2SSqRqAQaxMsqlea5kvqThQBiiABmEmtiQuF6vRyDh3T7vt
QD+vQA5uCU+zw+nZg4LUs22hatzF3jMC+SWIxERzWEBn36LKmzj4jlJyniKurJe0
rsgDahLJoBLnCBO2RgvmoAK9EgmeI0FGKM1UNG9EqPzXGniIMSQ175X/hsDaOJZn
tkOlLB6SD6dFjEADxjdNiQcIcTexr7zAzxcFpdAgrOA=
`protect END_PROTECTED
