`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BKD9Fycx2zX/TiDJ34FXOrTqFnSBD7/W+fu2kBGYot0xrVZ8wEEeVrpO30t/JoaC
nuaH+KbmYCOpRTlRm55Iph+YaF8m1bQqKUbOOIQa/HlceHLK8Uc00++cEVivfD3q
1iB+/+IchCButCs5zTv7uXq6o2D/7ZT7rWJiOdhOL7lE9dYX34V7vglK5VweiC3e
Kz54V1S319R/NVLpOqJ+2+gPlFP83VvwYn+Hl+7bp08rgrb+8oxUiReHead6HjMM
eW6pF+TkuMROLPp/CYxj5HrREuqwYVSuDFOqhFwrIO263u54c6C6aT+njemYf1Wz
GuMmcasgMQ8OGQvGDn3RblJJ1meMH8BcFxXEJ57owT7VLqaVX6w0fraw7ENHMD/J
wtkB3IR4Rw9V+icVzRjCwbLLxFB4Qc48sPJkHLlqsU72pOm4G54cLeX4DTNlXYLR
FLDY0q1p7nY1t4LReMsHuJ75FAJSbbqTp9TOlH2p+zJKyg9oucX3OYgTtGyCiX9/
yhQg1YmDQ7MJcYHvP2nTBKZKNnUqWk7OpPyxrgTFTRhcRF1aqSlWOSKwqjsDocKo
7V5Pt01akZvC8UKBzygfauCC4ik23k/KsDtWT4RHQKCnrWx6Kz3OcZQQKuy2dRaZ
/174pcDX/2HFFhDlzet6fBTxS/ikm27jDCC43Aqhw+WOVw07eKNLsMZawZFYU4fb
SoqvoBhDHbnWLroN4zBSBmN7VCMNr+AA231GfSXigbN3iR8xNoQKC8KQNsBHEt1v
L59vVV3199NfvXKNidnRWgHa8uXe1vQcQndep7VpBwlAiBL/yYaIyLP+hHzjt+3M
`protect END_PROTECTED
