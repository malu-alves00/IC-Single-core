`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Idsl5xA9VvCvie8corLbeWGRRRzVskQ2nvy92zannJH/OZrLsYuy9DFNRy72JOOs
hagooI9ugWx9BtTXHSP1FpDIHNST3vBt6jdShp/sE1YZCvBg2x+HAe0GfY1u0IM0
A/0wi3ThQ1D2CTf66Erggs4mXRZc7iRgHROaWbzLN7Ebc0kglaq8t5LGMnclp+XD
wsylKHa3E1KJ2FiqNKKIwqhelYWYEUFHXmZaBNrvvzqKlyhiv3n+EBkRxZ9tb9mw
7RsM8K2W+zxZM+RkQyBnUSRuubuup58/X0hiA2HLEbk6B/axh+Efnsldvut8kRMi
WH09FxDI0yZRSK3Atppu1nz0NEQ8jlODGOZZLm/yzneCwaQ3JAUhOMRpDsSfiDO2
u6XYa2LAAuO9pc7UM643Fr5rJi+I5JBs/RTYlYnQH5SLc8jb/jC0V+LRvP8EQArL
/zZQQdm4QtplX8T84pLDmlqCaIAa7yLcv4bEYPVbuDaHGZiRcNalwbFazE+5Mb05
ExmY4HTrzKEmNUdi9geX7000EJg4Cf4oZ2XhP10GPSsmtXN9kX4YuTjrZtOpYcFG
rpFWltsFOfp8F0t3Pf3dtIgzCloO/JG3eN4J8U8b2mJYFlk6dAKbm2TzI/7e2owv
sqSvTB8mzX6OXLiqH+VDTdYYo9vck2ji59w6P6LuvY35ViZByH/1IFYLMP0QL+rU
6/dgLCJVkq2EN6y9fK471/0d2gt1TkY4RmOuJbTACbAmrs1b3GHb9T4YzGEPr6QE
Kdif+mBK+LjJrDmptAD+hKfncrqXFreaOIqySylzJ9BNcR7HxBIliwc7yoqS82Wt
`protect END_PROTECTED
