`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
f8NKJVan8thAROaCYknV0AoM4M2tXT82kmj3jXYLi649eXvR5oyGz9HLNxJaGNhd
v5oBKuLwFCb08u0VIumIBjC2tDJ3uP9H/csRDe1QOlP+BIT2wpVOFL8p7inEutxj
X7DRdGNKenqKnIVczRywYuemlsho63+s8U3+8a3MBxanQvx8g3HElt+6LuBqn9Yn
QFH8TuBpTjxA1WP7AIzzcaoFMgp+5G2fMQq9ewD7j7Uy3+2NLxCkdRKxW2Cuotg4
+Y6pQVbKjnRkYaeKB0mdYWdiWeYXT3VRbCiIi4KX940SUcBAn5rHWcKj7RqZ+QDq
7uQxxvEfRdtWvaCcr5dWa5jdGuYlDFGpx2YfQd43h+8M2lZQn58r+WmAktquBFE/
jL4i6GKn7B+ahHaiJOBLUnso9lWmOJQM76Nymne0GxXaqaDYazW6do0pnSwvhTI+
V/O1PjUqO90czj7RuVG2lSokNcSpWXPro7CPWbSMQTdg8BhKwLISe2e3+n2Qbkq7
hnGmauyE3MuDQOEOHqHqcoZLb8tQ2ql7JRUkgWno4VTfATsOlTRr4iPG2QpPqXgE
Vie8kCJgntDwWpQ+pniUdJFnDthT625Uh+qN+CmnIYal4Wegtxcuq/7YtiKQ3aFd
62XoaodWAWaGK9fF/glMxjhPjVD9JknqaZZTfTZd/FhGvlCjR71XVQg5dZwWQye6
DU6krolL5yBRy73mGUQa+xR8mqqH5OpoMCiPukz9HU16C8Ot6xAjHbDuRv1gPjuQ
UK0dTLh+oxjTVlfuUO5H+cVRTys2Y3/tbnR8rm7LSPWITOCthFIXTp8e/gjlTG5D
zEET0vNCiFhxvAhF2gaQlSmqURoNJrmyktsGj014EQroY2FTr/kDCPB5iJDtWfp3
N41mAfKaSkvdiogvPTEj8DXhsTnKO9yXJrgXyIsTskSYzPkQKhqG8Zjgg90xNHro
7yubFlUATbeG2vLnBM9Nnb2GG0rLxwc/FLLcRenmqpTUfneEkpqWrVnMpcyKJDaW
DzRtPHVS/2vnVhRP5GIwfuPuI1+fhBZPlfUA+j09RzxPKwpLl0EpE9PG01Of8JzM
b2nuaG3PbBNAlRHzx5A75z/nkGZcYyo+G1zoyjYCMJwcwz7xOz5d33sRhD6oGEoF
8HLycO8Drpv3rkT1willfjrtb/Slu5k2Uc9vW/D0b72U8U8dm6yUOobQsM9l+JY4
ruyhbIybkCGaV7DIURPbX8PCMGDaPYsV38T8jUoaHYjQHPhOJ2F5+th/nCXnc8kp
9Qn0DN+mMPaVJmLp5BtGS0QSushOPsyuL00jcTWvARyaffOSW5rbrj3SKcZbtjz8
UNGBclOt/PfjsHlPBFw37OpePv4qgrCxsxbXe3ZF4QvD3XWyArwtVvb9FEFrklqC
CTDZZMMMVfzK+M8sDEAzow6cXKkRW/1prDph2NJcbbmyAQQIFM+Z39F0vYFRkNud
eH89FA/jm6z6ATqZPvbKoHpEbEZLHAwgZzmDFs+JjHhSkqKvZKY+Ry1TCj+zCYNv
2ZVD/eX62SqXDWsctOy7TtMBfkQPkrulx3BNMi+eZF/qrLIHTh6xKZrHd+v1KiJP
TEp/YbiAJ+k+vMi+1cvjqWXHL9ak4DUjWHg3j3/obtwMG1vcru6158i+fI1pFB63
vm3GybkLtfsmfzmPC813xMS2XASeCQ+ad0k3mOpsU8DANFNrevtIZ0yQ27/G+rtA
DqnpamMmEU4YpG+brAmBhA==
`protect END_PROTECTED
