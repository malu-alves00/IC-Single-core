`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EHXndQ1T0b9RSxfS1O5Zgm/9LXnR2cz905/i/dTckb1pY94r95lX75mlY/HRd4Ur
vpWRiD56eTxiljX6WxI7IEsJ+7W34aW0ofJVXlvBrK9+BwtxWj5SHxDsXGljESPf
IINpbaS2yRyOp51Sgpohr2KQImCmiHozgAoNl6hm7AFAOPzK/rQWdP8sy6+MufoN
6IcPbeqbYGCHfbQYbfWi1pHW41BwCNT4eW5qD8J28LTzJxGT/R/vv7X4WcEDzT1g
3o2Ooff8qnKxUrQynnyxLnKcD3Qlptjtv5wu/kRsFNKG7c4vWceSu2u7qIq0H4nu
g9ZIR+nZSw61EIvizU/HepeDuSPhV9Rn5kxv6zyrR+kIP7YICGNq3glMc2sF3x7O
vuT+lru6LNPIgkPIerB98Zb6E3TtwQnhXpf4frZczG49PaE2D75ZTV0MA4mUqsO+
fbcQnHKk42pUmH6iZwXqSz5qcRNcMlZfRmExANvdxGt8uukX2RS+nE04/Vmg9iDq
QdonOzq/eNZkewpP999zKML/8gbhBVAvyUPVMxlCbUp9gr6nODfXbAvuLxv/IHIb
GMB0/0roF2T1Fvo3eno00jwyaehx3Q6xnzfgIKItNBpgo7OBCLZgpE49/KQcUBFS
`protect END_PROTECTED
