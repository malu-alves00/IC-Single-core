`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0wisH81wbueXzbXWtxYFMTtROGYOnyKpl2ZYx0zgGwlJ4/EDySMjGXaYwi6GQ3r3
whXlTVTZV1/F+FSIdqvyWnkBIkl1VhurXSKFDcD5/AHeF6JHWcEAgbdRhZPSu8LI
HGBeDLCFkr1CL9nWXp0zN3nbWmgW3OPZEOFkkEosHz7KB9YMtONyI3ei4IWsBgx7
w7eHlp0lMAy/V9VEFkyLI7pxVezvR/uGF2EiKKajTzT1i7HAiwV807fM/EqduOML
Sluotcur1NuAjpOykxYQG3XswaRptiZ/DeSpOT9PQjMTHkceuMzD1dx8eeJwvWBg
1IWzwYdXo4J0huL1Y/JlGRMhA+XeX7NdQAIGcpjXltLl+anxBt4ZzNjs3GdMOa8S
GVF8PDfr4dWpcidjqyG3bf3QEdyKoh6IF29VDCah7Rm2YkZ7d1KvrC6LWmPYwKIZ
8cZgZtvPZpxXO4mtuTY1Ylv6WY0S+t43EFccJjAVacoOC4uyTSE16OgAisbQo/zL
roazuFqVMpbxrGhtQWz4Q1nOSmnO04tQteXcqSSPGs+JHUseCRV+8Z0+pZeWWqMv
bAliQMKWsoZeImi+4HJpC948No3Dob0pxU4WLLr2v8Z9t+K/S42yTkYL6NEGQ8u8
QhSUslUFP+pPm7VAz2pm/xBtyM8Bpk32dxmrOwBx0k3k23gv5qwXxrHuXbuHyeQs
I05BW9Jq4/h6UreLfW1SG6DCWA3uHIDeKdPAfHljYf0K7LeUhuuLOTq2ZucSg7a8
maxMBA8tJ3+9iOcpjBUceA==
`protect END_PROTECTED
