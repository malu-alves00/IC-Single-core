`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nEXr05qfvMxZg9StwhVLa3uZ/DLYcNF2eaWtBRA9y/A4QN96FHKwSfo3IPbZvk5i
p/aO/fvMr+acPB+EYBMYRB9qCNNgRadSrZeKBDqPJDQEMT52X5J44HKIwuNe/M6R
BQ9iSmDmVwI7voAX6zK5ayNanrvaJnwz6lNs+dl6R9viLJp0m0Z11vPzMPjUfb2X
e4neTEomi/8nplKzxBeh7p6FSO8Gy580khrd5CtecJNQ+ODV/kT45yNYCLOZzEqr
Ba17VOLUKCjwf6JqiujJKPJoeXbOK3po6qDy4zahgWVzqnWIm2KoWJV1y3AY3esf
Mz7tH2UsMJ2mw9Lq3RdduhJP0az1MZt09XAM4z86ew9uxR/7HAsutIPuDR2RGca+
1U3zqn5KRIseKILisfgG0driav1xLQrj+TkmKv89/tW8v33tUU/iwTbGkX8RyEtw
p44zQTN0zUU3zyhHLJcUOvN0OYskFAglZBL69Pt/9qeF4mVufMHVPJk+ka1NOAgf
u4eKm2N0Y4nxoE6X9txeP8S6d0dAjS2mr0PNCVWsL/cji4j62O7V+WcwPVrKkRLs
/X1Q+q4T2qz9y/9iOvDcmqUe/Shx1/VoafbfNWjut+RpntO0/5UgSJvQe9HCoODt
7khDczh0VSWxo93UdwiqssFwYbD4fCOjXwSU1VArY58O6ayZiea81NHNZOmSeYuk
ofJSwmIGsItOj3Y/wSfgE9vfFDka3sTfa2NGO4NbkkE7O+HRmJtEKkqg7bkuHIB6
RGpv2/2+YS2KNm1pq/lIwdNMeKIeUef0rGJI0In0rJ7ixbnuzrOVVZm2Ywb/1iI/
bYj38DIe8Vprg4T4z1QVVw/xYpx8MjbAoLCnV5My3nVXV33NrO0tMFqaNOTulaRO
ocpl1leht4Du7qB7U/DX7PIowrrGzTy0nsxwP9lMcb6k5cLvrmXVZDgHIzymE9qw
/82P1OS+rZgXWZAqLPnYn8dOlqmQLAJs24s8hKuRd7jRHN4mrJhgtZ3qfRogLXEj
RRYfMexbgcCFSPN85M7sXmc743k4mq28tuCNw/0HhLlFLQsEtSKk0Gl/5tVm21dg
b91K95f/u+7o6ICT9lxShJqOsS3twYQ59xdYWGd/IHQgviN0tsJoexkE3AxleB5L
jRi7Q5oEy+jDsR3nsXOIeM0UkK2fcIbsQH86c4FqcK0EwOf4ebuAmenvBqk36srr
bvICn1Wuziv57gD8pMs7kPGxGoPJXuA6atjBJ1/hm91Jc78HUXlForwHj95ANnnz
qQ/tz/Sj1/ugQpfCxq6HoZJ5BepYPY4aVJE5X6wEbDAmhYGsTVD6WAqXPtxB4J25
jbLFk4Sl0bz4IDIlMc9evc7KamDqaktxebeAn6O2YOmJYc0wKkWlTtiE73uYUkXs
QeAkGCZ35LogHjrn4A7T7jE7zCfQFudurUn/2t6+3+vlktmy1+4o7BHzXXzgk5Xl
Nd6ltKk7hLAg14KqmGflATvts2KrLdK2wuIIYAi1b/P4XaA00AHXxVtuQiAjZZ/B
mR3dAojEbPDDONc6gS5mQbNuw/rRmaou/AAdCLf96MwPz1KO5NODfHcsRKcdXnu6
UvBXZbHBQJBQcLfDGjDW6X6bnAb2DS6sZfvAxTZ8wFmFlB8PNB0ZKw6MSQFF/I7A
h2dmxVIbR3fbNZ5JcJ/OB4lG6lsVK/KF5yg2B7a6/eCPRf/IEUm59x9DGrqfEP7j
CjETQfEVbHMhNreInT40DgbJUHU0kPcFMJrWlGqrxf2r4++XXojxj8s7BQUC8jv/
0P5CIk7zsgsnj7kGdLNqFquV4saTnYoSi072YX6MhpHIU85Y8V85wHzbVZB8XNmw
0UrGYaBSPdsIXbHL5DHo8V57fXwc/wkeSEa2nkcLWlF/wRIeFOhpdO5Nhdd/MDaf
8Sdf3UvBAkTMO5OK8lNN/HEPk8lb7DpBoF7LjGU1MkXooous9slzSxdgcWjceyWD
uJ7ddqtbscj4RHHdzxhAC0oDE1UqYdeRym/FPyLatNEwYYlr9TePz3FG7gYvAOF0
Ph9B46w/eWfR8SjaHUDiPSnsump5U+r9Tt+YZgxnWiJWT1UWsGrz0OZj2EHrh98Z
mRrfxN1f7PMQtsnavrlmQ2Ou1yKjGI5QCnDP2J7gpjOSqPhaPtpSSHce6tklWv2W
gsK/slknB/QAmPnIVQ2W8CrtHv09a0n5GBjREPTPMrJXlABAkApsjlwB+rDRCanT
ftoqi6QvEbPv4PTl0421XJx/ObosPg2tq9la1INJ6XyZFrNvm47mBPIlVRh0LVJp
dieT8buDejjrbnzK8KWWfRc3+ifzScBLXG2HT7AmiSDgVuYPhenVt4/hAGvMo1Sw
0Vr7ROtvE+4KkejK68u0WZ3S+5xg26UJUJuOWiViEUbADD4nP4Fl/0i8uM2x15Mt
jzPR984lHxUtdYaymVEirUSiXR8OsMUa9IpbwfISZrpEjx/rXBrilufffn9xRrkc
EF41fRCgQg8xMpqWsYj27/rkSVlb5q01fwxREjjZPKv/ffgBRpMKi/YQRHBEPnOt
UMypCAFADcNjLUT9aGsZ4zFCbgUhPE8g0fTMllwQZzy7q1UtteqAxHHGtJRTXnqm
VU6DMAAEV8cOxwnudKZUaxau0dmbkNp0pRhyPFYZfav5BQSQGaQs/H/z9WxJU9R4
LFUdaamNqnJdF7WmXPGcwvpcHrpybgxcCB4tiKJgWV8N59qEt2KT3sXBqrAjBDTa
d1GPkohVZ7jNRfvsxnxlvD2vDHrDppN9F9M7bcwo+EKqM2TF+EA05nPo2mxMgcR6
ylOe4nhRamOskEcwEzNk6v4lHzhBtQg9xemPKJ/Rq9ENyYoRXrp4oeAYQaoM8LWP
GBLKbv/pQC1zYBADdQzKWNpjVSJDSdUEG2elB9YmGAi9VaxL1OwMNh48J9Vfsppy
UTxd/mIF2LrS3wHDdgZLqYLYXcjZApuz4TrRfeG3KdFgA6WpkUZ9/iucMpGKD1xZ
v9lcR/SOUjdptKIyJVnvfcH2c6nlbLfJi6Cdddqd4Ygz5ZMUoSwPuJ8Jz6E+HAb3
camuXvgsjguN+FAkF6GOUyIBdPpSX+ZV3FF2Iey8eoxizb4FujPBg6AyyDBKpoHi
SmaNuRcTXOUV6d9lx0OfDKEIAqAyCJAK3BbLHa8mmJoOp22due5QSyg54Dc/hzAF
OCLUeAaa5FKJF+UsPSnUWkTDSXBV2kOH19/17z9Wh/hZo98DzijGJq0vdl7qGgoW
N+JPaoFTxkai/ANO3kGAWOhvOMZltCx3BZIIjWyy9J7ZQ33F/Mez9JoHpRiJpMZr
hrHpPi+5zjiOugbS+lQboymOL/Hno/3P+L3S7JJ/Sb7dOgbl6zkZuPxqgioL1kvt
RKjczrjPCICJbhR2cwBoEkLgb0mUdkMvgoPWDIoaPZ3GrXWtuUbbK3j0x1piKPL0
wkIxc0mc/sgTqD8fS3BS8uqPpHFwY7SDhxxu1wctKQ8768T0eY0OARc6Lmg9TFbm
or74/ZRd8eDRRssyRUcAUPs2UOS3JAn+BoxUs1cQe5PtA7cvQ1b59aI5VkOJgIan
JEoH8cUnpivuzXaDX31Y7GVdhaQEHuTS3KJdcCnANkYwv3XjZnKJe9kdfbKKgRsO
ClDDZ2qG3zDTgiA3gpXOp1+H+pnbcgMTttTHG5OSZbY9vHIcR1spslyOwIzQA/8b
LMinGvzB/dmCe5v0yGCo209USXH3uqoQi8hqjn1kCS6pBOQInbzsgeIfxc3XdSM8
BT3s/EkmPG6ABiD9kYxDPQi1xeiEJJS5tapXPyU/SN+Y/m/JIguRlmquuU5KLL/o
4Vhin8is0j8S5PIM14QcOrrTtbN/dKNob1c03fxr4RyhQQ9+ONNQqoKXPIERKtDp
+ZOassb/MNKJVRJ+Sfy/JhrY7dm5DcPXAN9G6/hHI0i6WyIfSeDwl55aJF+NAsRx
multixf+aEayDWRoFN7kpVWrXfL+MPX/bSjKJAMWY4YGrfTDAF7b/OhY0qukKhoR
fo6/sVUV7oDKCiHl4OrbT0adiIxhP1oJRyjHGeha84YaDZkhhuxohJmDn/AMY0A0
+P2lptlhf2yjQomNtCa6o6Ej1rVg3i+mPaYkH8ybCnzvW762jb4gpboxpIalHaLn
9K7KQ3QSB1bdrrH1ODEub5ClgOqxplTU7Xp/FCG2zl5jNBS7CjjDSWoDj7y4Wnr3
YE28UcVH8GPDs7GuY9v65BdfGhSbWIUGJH87QGlihlFkOso42hqglJ6xC64rtdW4
ZTtVk7pn/DL0QdeVHpmP7YZPX3S1eXRR1QxKb2CyEdlLNPcnFUOjthtGmKH5mZhk
69rqi61jySuSZODttWVwTFw9TibveIlGkh/RyYVZbiyB4Bdmy/NY7SYvtEYBKJAx
ZoWg1KYu037XXPYHiu1NCaQ5ybFhk2BxicfZa4C2m4JZV5yI3uTf1ns/tvz8b9Ms
lwAX7F3MkAZ9kP04fPs2TKCAj/f/XUnO3dIJSTw5b/6TANSUY3eUjKQdWYGZ5nAK
6aU8HYWLNpcNJUnbyLgKpgMyG5krEULPXmJoNRJk8QdAj3bvUyDO7yBLyqnTwqye
7Csh8OmA+2Jdj5JJaO3JaqRGjs/bNQiHA/M33zjYsctTbvC21e72zUQlmmLTKQcu
opficr2ftMe4rHlDuy9/Yg/qnH44RnnzLDkVUgR/RV3KGbmY1uMHEak8NMgfdvH7
mWGRKnWUxdk4DhUsQaMpN5eJMkdb1qOnl8352HDh7OFvs2oBoZVvuD038ZBc5LzB
JJ6OGFhDYHtBNaUd7slFRhqiJKF6Y57XxuiLdtaXtlBshdaicpYLAA8HAXvzFUyI
D1MBJZ5VMs1Jafo5Hqf+Iek46mfkk6NiYAD4GlkrcHBT4P7WPuTLiMEOUSi4z3zh
f31WkB9ITSHxPGojVb0f8jZb81FhofdocJ0R0mQNGJgRnMgK2Z+GA90QhSgSEyUx
MdtpDSMu7aN6nXkw3KFUqBbrcrK7JQV33Nu+bib2mS/nRMcMlPWVGrC6dOuyyl+s
Vg9w1SXUZzwnFdB0WW9PXoz1rHSUeYlHdBGVzmkZcXLjX+SWMDaCJfYf93Lyf0VL
WsNkI9vg2YkM6LsA2me/FT74duVcoVGJloC4TVIe6ATgcNwhN+XHrkFQC7XcuYwG
/qwNu9r8neV6DCVhFk1zkF4ADKjFM7Tj2mioaic0HDYTsQ1xHsQUL1LbPN0d57vP
S4jZNBJeS6oHkzoj7EecVR8UTiHz7VzSkHNG/tXrrlYy7mMkB+8AT+F+KajZYXZN
VjUhdcHspplTR2kjKwSobGaItpL77W4hJ/3eoaBnYJiQmEGD27M7ZIFtyIVRSP1S
z/rROzWYe9Ea4/0BIN0DWvQDhcy168Ptolq6QMTW2d9Fx5ap+KYX7p0jMXM4cAIU
z+XYeHiK/CE+7m3iWanJ7mC3AT6SAOMuY7QyS5g05JbsSz4aQKKTVB1SSYslX4E1
GIz7lhsUOFfqQOI7sFo+DvBxwY6F/Wc36HYvtA4wiBV/SgsXrEj91CsoHnrpluji
C2ny5hZgupvehpaj8zHmBiWjiCg0tpmkhH7DdMaPaWB9lFeqOUfsO6+LUzQRAQJU
gZJXg9NzBJF4B1sXr3O0lsbr6LqqdJjjTToBBJOdr5e3bEqw7pJdPG3okYUwOVdd
nyQ5Fyck/cUFAL7Z62sD042XYcdMSafv6PWB0AIAzT2RoDjTspy1+GrGvt8rO6Ap
+NmrQnRF1JfZ+l21R24ZdW6iZS8dMKYY922ed4UoXspXp8IkIg3kawkN88SitvOj
igcuUUabhXhD1yhn2XCbTD0KtXV202Wwv0ZVXCnAzvp0UUfUAXB46WrP1IeOkJYM
Dax0GuDusNHdsOP7l7tvqJ3E9U/6LOa8GGk3ScKcEHDIyyy5J2WYz/e0IUSNXJUE
m9axXrz7pDcKUzqv+JEuN+Itse+Vqpx4Fn7UuCd0LSf22d6b0PyYpFtT8wtRgyKL
l45bSdrQAzPaWMmieZY6CHNW/bssOgMVa7NV+dxNMbCyX8FvNdYdujAE8lezDN6d
lfUqx0B+0LEpTSbjmIXLY0EUPbcWmU2kytnKJmsvDrc1MHyX1ufNrp7uzPzHLV7K
KVztULooN4gvJmPdnLJcWT7ZcAdojYJABN/R+hjGPZPcSsXCPKxiEiDCF70zD9SR
iO9Y45OiBwdfig291nPywf/3eP5/JLQeTSNFPTokp5GDbVYrmnxVEaD7ZT4EPTVg
ymc7KAwK2ZtMPmSnaa0v9VSRoEsncmCbPB1Ij872jPA0WqUTDhOdVmvrp7Ae49XJ
ExtO3SFvYMOiFg56K9XWi8HIjHhAvO4CytWZB3mYc1vPC8c3k5qL03QYsp1KFpMk
ZNUQLYPiN2A0Ps6vw+VKVFefXbg6q9BZeRMciLowjaUj1ItWi7P9iRouKkgUvX6e
UvZkcw5gVCp1c5sUJZ9bIL3FL1AabFeREhUoig//nJqJa4aceUmH8V/pJiCj5wKh
yOsLjP3Vqsflh7vHgRvNWsz/vK1OgXnlWeke11iZMsX6XjH9DZQeahErCg5pKgDz
THp8xWOqNo2Q8V+EsSAGFktdInWtcsEFsoCxjhYZ/MKM8qwKL6wkGcGcE0fNEBHZ
lTCyL+YPLMCf4TkZeuUGsXRpBJJ2yfpMVCrWM5BdPEWdkaC9j3Oep6MimVJp9xIy
qzkqjSGIHof/zrfpVduOkG/R8NqiK4r0dzj7BIYIsQ5R0FVsjPGV8X/NWjxRqcfr
QQ8/dg+4b5v2I1j+7T0i1urO9OCZa7IhnYt2QLo/FILg+UBILa9Mx/7h/m3ay9kj
QUaBLIJuw+Zs8MZLwhzIkFnzHRbo0y+vH4JRUYAHWWpjG3AZmhMY67qPg9KYSOut
nmn54Zy9fAOpP7Wm3Ebp00l1KEk0cCxOdUhZ/n+k/iG7dUhGedeCIOL1xkQ/R+Cw
G6oxu3DK8pmWftkPMc9L8YVXIX54xOKaH6qvzCK+49zDWJ6THf93ru6I9XJaGxc5
c9LWAe9hO2G64s8Ca/clasy+BaSD0TeS8MJBHQ9HuIzo/roolR4npgt4ZadoUyLt
ExP2TRVyWsXpspNquxo3D1qU1BN9EVmePtQHqMlhnL/wbsKlUg4l0HWvHEzbx/uB
QrH7kD+0DYRubwdtAZ2V/5T9YMFiAuq29VCZr9ASvyvm2tNfde7iIcxUD8dmpC1X
f5Dsg/zBYgPju3R+1wH7EuAjGW3z0s94ZYRWbIbILZa9X3z7QSpPxZxA0eWtFPj8
ed30R+O6ey+JeQ3tFudiSfw/oCbeO0k10MCpSRFAf543YhlkY2STB/7zWGldVJzC
JaZN7f25idNXZEIffy3PDVL4u9MMtIAXvk4xGh/Xma+OjaOS6eKmv1rix0vfJbHF
PBtu2AoHyp2ykJb/cEmBjjfZ+Cs9W3Hz6vypnbNgtNy+YLy1z9AEJVbm7qcIHQf3
sLAPEPNYFqHZ9k2nUAAVuo9DZGhAwO9gONeVwrLkdVyA3z+Oq+E+OTE3DzFD/xiP
cTP0mFRnDDdWR052Ywms2984859A9nxgm3KFNknwsCoFUDAOitdXmQ3q2kT+Ijoe
2Tz/4wxkkbeCOVAFZOUZJF2ygJu6l19O19lkcXtcKAuC7cHHXEgJITSL0+zkEbIo
qaGGocEqbXYNt1zOMzddM12l6k17ebatXvqqeaG6BFMeSx43AkUdsLh/Pv/VQpjz
ODXq3YrbXGtVXnWsPIVXm2Pc5OMa6qJLxZmRrh0dnbOwl+p5LMT/iKC48/GfFaO5
DW2Mv6k8EQDY5lEA6bSZQ4RGy90TqA6C2GXVmEFGOJ5CJi/MDZmZqGfu6/AOUr34
CMQKGDwFSGzBvUBvTc37vMX+ic/Srk71QBcOorI1gTgCHa0tVyWmebL5kvUcDgeS
sioPTch7nnFSrdSSwR8YMv/sEfhwQGW8mZq54WdN7YXyMw8fPlHPCILrCWgu6pRc
HPuqu6nyiwgftkNXfmVFXIXu5oQ8vcA19AleplDpVW2R7wdkTrvVrgR4aLPPvGIl
9w3kEmTADTbrMiQJpguL8oDdKoJUKUG4ripDW1/bM+2p6REt+NuGif+Z2XcbtTCH
hEta4jbbgc7SxS5UMcD9+nljgmRB2MCUVcjU0VV6WEo=
`protect END_PROTECTED
