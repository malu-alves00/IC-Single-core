`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CJQ3GW9iK/3T7PfJPlbdLrl8/1cU9N+QgA1jeAWH3DLIxwL7IN1rtlpUEF0ISEaa
mxZ+EzCDRQE6p38sN7J3402xjNWlPlJXM92GGCtoWz6TX2hrnrvUUcMfijJKzTOH
9hutpm2XUwY0qYsjt/VVo6NXFkc7Lr1hLPNg2Q3AwZciUTluL7Y19HbGfrTR9OUR
gf1NYvJ90VPob2FAtgkBaqG4jxS3Usf0EMM/sCt62I0Wfvw4lsP5vv5ELAJi6izy
sBXORkyKb/7OXBDEjcyLhd5rcW8KOkehxH5Iq/1Vj6gQgOH7uWn4h/V5vg8TNfgX
hXzsdWTDjNMRBBj6u/pZPd5QrobkHEkW5TpQOXXzpvHGQd8Hs6X/TzfJJt3PTJlv
p0yBEzHh49L9x2XvWSY/NkqHW4cGnuNOhGj9uluRFaM=
`protect END_PROTECTED
