`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Q9VCH23rZEepxVsUreIfatR0TbGVuNlOeoxP36UD0+wMaIwnEInOkn1L7OBV5Qo6
+dLqcTbnkyw4LZLGiXEHPh2P+OyaRlRVs62BuBzIQdPTsuCcefpYcuUIcNGQD7sd
gfj/Jb/uEKrMF34rNo3zA08vera0enUoyMzdJMWYdbXiKWISnVnQzqamuRYLdH+f
zQMnKL8cT3fGX4yiYq/yvjyNm5YohoRt8fvFjy17WuVWymBdor3k0fB5byap9AVw
V3njadcguM9xEbDpT9yFaQor1q3IgbAg0yJBiA6hQygOZe2NhgEpxdTP9EYL2qTn
oHMFIGiXa+dUHHt2iZz1flEx9jaBTDNWmVodtR0MN86vH/+I1AjfvOIKPeOIkyxz
nOX+4Xl+QxjWdnAbBh8PPvp5NS5xuakLceT9Nmwdr+mjFrLv++xxMwHupd8Nb3LP
eA++RSmiKzYFyYsjS+WhUVylwcq1PY9BvcA3GllkpfnJ7Y5yaBEufo1ZHpoTfkDN
BmcbeFO5yKzsNuGxER0wH4/MV9lns6jH2aXWo5Nf4P/VmU75uqQhP02k+xOodlgS
mp1395BvG4VzWqlRt8wsY+paOXc5rEErtdfyYOuadMhnTGyjxnhNU1l6KdrH4xqK
/X8a9+2obtt6jouNJO9s2VeekD6PGKJwhUyKNYnNGH8pCC8gcl15Y+HbJQ5TIbwM
uYkZeqZWkajURzU69nxYY8eBuOWknF5SFWyYwLB93mtJ3OOMkE0Zl3XYFtT3KGBY
QC7EEPWXTidDZU5GsgouCJUEFv9GRVZt9PpVG/bVib6DmqLLhrAEjiLGarxJbViK
XanERToPa+PCE+3PVxMtBzmiBavfzZztK23I+IzGbw1zXcyRiDzQ0aQoRWpoGO5D
zAGWr6gQ4jl/oZCMc8bFdXO8HsmKHVAWh4lQkFbOX7xUJr8Ow0qqXpHhGxaC4p3V
7K1M3V5N2iIfcvZVVsHFRgAqEgtGWpCX3X8VODmB8DopXve92O/TTt39DVsUwLUX
Aqk59RxS6n8N4EwEZOtEtUTPa8iumkP3Cq11BrT867Wp3cwN1tuyuJkNpNyfgfLo
CiMKaw0Nn+9zHZAR297Zj49jcZXms/sxqyIyKTOJgQBPaWjTd1KG7vsppxRmVvDI
8eS6yZy91nfqzJAYpBcr+an98fFVsh+R4o7pXInlpReL+XxZszmaX+1GWBSncM3D
zb0pUhC+oQDW/LxPoCqaDGElvOj82WfUQ/VTN1QBzQ/93vOm6Xr9wfJulCUOji6P
g/uxe74QR+6IKhX7Lk3aJp/eOk8/A3EOXVypbaidJCLQvQ4SHr0s1e7YHwQK9NuV
S4ydCWdsI/TmYKGLP8K54TY0XX8XsAvCGwH2pmFM2RJ2fUizqd2gDlhEJ5Icf8EA
eP4nEmQe967yMllu3uxQ5XMx6Uc/KgI/ygxnwO1ywQi6i2XfJTGScpGjtihGTuVb
4Tw83d19DCxAygBgGHMawo2lj4nmJkXD/kMW/NnV9GahOOl5BXwqmQ1tHoWXhXP9
3nP52rdtDbQTClYr+Uh5F4u1yMJhuNfKa8LkBSFZf3S6tM6g/9hzuh2ZxZ6SQpUh
VarvgCIE2L2r/UGqNfqOlTSE11f1Ss/fLlAVtZ6zO0gXXAsBL29fxi/CKwQlvpqf
IWYcRuc6J+rWsaRSjKB97WQwKzI8lMRKP1Rjz6hFGV/YOFQZ/Akmo4lubUjkbXGJ
YcDeCG15j2lPPBu/anhizFXGJsE+UOufu/CcFHpqPPU/hglfJwyU+mWmonNCgMAM
e1+8kLuJULHwsYdokmRfsAMB3IhOgxZWdWwzqpPfpmmPDFFdQsSPKZE1lwdBqsis
jK9tVhMamd6G1lbWBjU85zu+Pl1r81oqlJxtQSAJ9qcLGdp9g1LC0zlphY9I4Bc5
E7/vI1zlfJyA23H7vMr1xYdbQJ/7qg964hwY0PfkSUUAiF/c0UsJ6/gQ3hZr4wCR
bZ+uY6zcRHau1e99h0bmfA==
`protect END_PROTECTED
