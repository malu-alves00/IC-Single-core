`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sGHQMVPf9hsxKZzLvZolcNXM84xEoNRJuL+whlFTcw86ckGih9SyfmulyWd4V1s5
wZBA2ugYnnjhIdlZpXYAEsBAsOKHIFxatuPI/hiHYD4/TcgfwNBKhypjr+tmYyq8
NbivK3Ahcf1V4BievCySIMgFOmXNZU7tfLlf3I5/OPaOIzJuMHaUS/WJy+sJS7wI
8kecf5rHBj+4b9Qrezj55MoZfRxTEexH5J/CSH6wQCChb51ZwviQrB6+jZZ7EO8i
aueHuOFJjIcWkuDgecAzIR3vu6UBzq0f8spMfAEj2zzWXa4YcuOjWm3Aslo7dFo4
yZALfPJQIcZfg+eXkzbK9xeHHeGpIWIA5hdjjkWoWSDjKBbw0YwMe+BJedBPD7xO
GeP9/Lc56nL5Jo/9xUjP6LOBdEXYBzvluDatytrJiY++K4A9aLvYGGQqyolJ20fn
ovKZrjyTdXvp+EU0eav5Zk36I17dTRNVhy8iR9ziWticPP0aJA1/FRmcTUgAZKw2
MYugVL/R3slA/1v8mLY/ysX3InoOlmPg+X9cq4JLOcT6WFi5IYG2nWrnuYN3HDB4
bXoxKOdhoqWNoRacLvPpo4L8EglqDjBjuqw2hJ9zNZY9VAC9rOReGK0NUIWXHVGK
RkDNdRcZLZC6JUmB3x2lyZgPjMPB/7+gDgKG8KF1xHERd+d30+sRzZxdEedhYBvC
lmIgJwmRoSNkJsT6vHjlPuzp22+zoHEtydiPF71/kvnAQJkA07PDmOuSEi62Yep9
QN1PieGRHtpB5tMku4lSmRBpX9/ftaTt5KBqFRpcL/fqiSVlxSMsKR/06AGYj5FL
8bHJAkJWUy2XvzfEiqKGEwS7ySmHRgIkJuoh10afU3s0SCPB0X0y5/F8XchQK6/0
FaQjVwQswOlH/Km1yY5dzmDH5kPTNTqLHaWter80V7ySKjTHpRdWlKKK25eiYA8A
GUdLS+WD3ZBRuh4UB7KDmR++vPV/9/mG2+fLoX+EKZB0VVCnzsPn9gk7pFiqWZxX
wNxiIr9JxtjBRFKv2Uyjb72hPcJYVmB4ejR03sGjuxsn3WgclWe78o4f+6r0VGpx
uwNIdkim6beF7gIV1IRAv6y8Dxc+JxZq1Lmjl8a4rl7f+RVfbeAINzXKeMC/BBeM
Zcj4ofRoqBYSZSB4dT7PQY/Dy5/sHyhaHFu4vPGXJRDvoYRUTnjHeBP+BHvu2bxZ
UEtZCGFo2ie9cTX8q5/eZWYxESjQ5EKV+CAoLnzdnhm+/u3DgQf/KUER88y1GBh+
8FXrfBmTxtiIxrL0FTf0F+C0sqZuFSWB0X4aWEVNIPrdx6hpurFyWoD5go6TBwmY
/YT+PgvJOG+1th4rRaHuI5G2hwF5/5gSDUnlOhH+RGfZvjlMHY+DR7HBp1rL/4Rn
DuRY8HnAh62ZnVykqdY5qlzaqG62YV+TdnMBTHPRIXQXHXQq1b8NC32aoMqj8l0V
p+7pRcwmeHSc4h/xR5wgxakTxGlLio0yG2jvudFwuSxxNDieX4frsKPDoM4Y42VE
OZez1Y6WJVqqzgXRp6AzxD8nOhQ4WLHElR555dmxCScAg6qQT9MZBkFp9L6Nzqqm
BFiU1onNKtlNBhNdilUg9OAjmDrncgp6xYGhQ5xM6A2iUHTxnOwBcQnamcBPMcAG
IGZlKMWizdUz2pJcK47jPg8U1qQdctUSeuHUrO8TjhZNqoYla/6R23cij5b/b/BU
LNvQN88bpcSIhJiva3k0gbX0v8UYV+cigAmE352bC734l8+bRSxdBa+w4j4SJEze
DZ/nXae9pTnbLDzwIVFDjCKuoylMyW706/SxAggP/G5dAG327AJEkCsKhtsEDwZu
1UQTovfnzj8GdBNU3vXMghimlCIB3MgqOBd8mqLczbderbQRam0J88Z4zizalGXK
wDOs1NvZo33CakHbr2fIZYT5kvWHViNdBXS4ronYg4u201yCS2KKUenMFT78MarK
c4lUFZWu506APx5wELH4ulH7cLshMojrGs2wFpK4guhF0AwSaN/SWUD+HX0TtZu7
XEOMz8oqtbk9741qJGt7qkUxDv1hnwRSL3c0TcSJo/tlj/PIc1w+5/lFOKNnXgbQ
EuyOckphJ4iYraVBpjImnKsDJG5x6Eo+qe0FZu5KtNLx5o/AJkJNSOkYadRSju5+
yKU3gJV2N2xD68JpxoLq8hYZvkjmPUYjZYjBCPnyR6HDbdGvUTiUc0Wr0HvNFQdE
bL9D1Nd6qC63Nnm5rdYZwj/tbXwTA0c5IRhhXhNeFxl//ARkAvReLIoxYmnvz/ij
agQiuk1G8zrTnNvQrKYJlsy4LIMV5NuYC4sAeiBtvP0DUgwoq6mN746eGxSH0IYK
hhGbtG6hP6dcJ+cYJz+ndyOBU7C+LocwRxPKFPK47TNPDY0RuTCi+q+Vv3AxLAFy
6shDEMSfPEPZpxSw4ifrg7KZrlKRQRhjvA5EOzOCzrqcRYL5Z6lgZ5PIqqdgiB9j
/nxEuKNU+zBkBdPTg0jOCDeWuLutiIYypvv0FUtuSulDn+csdj5bu32jnBjb1Q40
1/Kt8ML7Hdx5wuEdq3rX2mQ7SgIkVcOYQqebwNdL2etakGR01jFKH5oLcqb3x1C/
pWUW4fKF9ZJ6yCwj0qtHkrqQ4q+LcdrqjV/Sybb575aj3jayKSNMgLNriwZD4YJ1
ulXfaPcQvdabSxN+TtZWNUGSEvVHpa9x+BQJlPawXlQOmESWORAVICtoTsUkG6mJ
9nwo94fzyxcOr95/wqivqFNrJcFq0wtfbP3uGIxZIbx9rnE3hPqshTde9rWCT5b5
2UjPJIbA06fpwBUodalQRWue6xrBNOC/vuWCxSCEGB26+zXjr/OPeiX7HJuAAZuN
FBhfFRvyzzvG7fQXZBJhcbD0YCGXTuvM0GjYKs/9Fs6KnrNQx5afsd2orRwEMXb8
4bfhQ/80zSP3a6+1OTGsWC/zled5yQBGPVa5/GqM2+6PWr6Oftl2LUuRoKFgciSh
y9+bm1OC4QPkhMUAw9nbc7cM4bcWeld75Hb8Qvl9Ov1IwztazM2a6SCjXktn2Zhb
m2z6uljgE+vud9D0YpOiotDL2nl6tiKxyqULXYVKbEjMhxBw7EQvHBcXbQHBBssd
TpQk9tPlPzW4ADj1w1am+Kb1O4lAimg/j2oip37Z3imh7U0sH8X4at90/Hq2IACA
LTiyadlqdtK/1wfeq7zgkH2gNX+LCA3IzdouC476MU5SWLlOtXBKeIIa4Bktgxi0
Q9zIXV7OQKHTzpLwYNPj8WJaqLeE78XNNwgo70sZzPSZKGaHIujUIG5iBcN3CBkt
Yfzo+P8Wawi/zx5bhdFCl7WDVSjP2Z1EWL7yyrtwikCPFXP+fTdL0YxVNknxQ3ts
xifPbJCDzWk2a83AfJSrOGOoDHEkvZ9RBL/Y0wilxLzp/iwgBFjfTxEh4qhKTKKV
5Iu47vgkyw6hINv7pm4cqF5TUVOsRRo2SLLuROXdWHOJbZ8H2lEw1W0BP3vBCz37
+ceJ/0yumbyVYZ6kcpodcQQBU9DyfaE0LqR2wzN4oX14+i/eZWpx8dy2w/fZgQ/O
tfqoCVy+X9aLHu1hTPBee18Vrxl7EacooVIEQO3H4tbr3r6vBP+bHkgWTqjfb6eO
4UElac80CLTafsKmQTOtJtin1rUIxyvLZp+kP8HX0nvpvoqvztW5PuNTDA6QAXlU
OeHMyvroWdBOyLqoQDCAcxx6oJaOVZsHr5BH3RPNHQTnob9IEgC4hMo02ZP1xdXv
5so4ohH/Af/TWlSQUkCFLIoWy/Y9oAo+w4ZxWRvY7hxPmxrhU95dWoXIaRXFDHX7
ycMc7e0JcuFVI68XaGs8sORO9V08XDZfjwDwIB7gWB/3/pbHPgo3IXN0fFbUsOKu
OlrWt7Rdz+2eI402za8RMighrFi4CNuUYbQc/R5kSVp2bL8s/uUNq5UPDgw45H4F
V7W2mj29+mtI4+f2S2VA6WZhM92WQIl9vkSpym8c7fhFQkGDXah2hQY97oG3CbgB
3nj/pGanXhtzLwp2ogwn+adDvQEQC/8ceIsb3cdCykW9jLo3pjsU4kudgtMBVWgn
iMTybqBlY1UGKI2KwdWxMHWIygdzEgr9cI8rAMkkDAN0tIrVTIzlkjZzp7KxzU4k
ORc/s3xAiZ91gL3C5kxOltlMHv+3+EjFicoHpCvJf21SGWSbY3LEccoyUIgEwDKB
DwAYtKs52PkMf+KUZ56z2tViXaXRCMSpEm+4hQ4Qye3Il1DaEnWVJfsh32GKkYws
K22Cb5QvpWPwS0KD25/X7STcMKFcmQmDa69B3QmkAG4sYa+qW63Qy6VEZmp+jVJ8
jrSFEwJD/ex8k4tZsfmTP7vY8RQ8Cy07/bpn/j8xpxvPDURawMwrJWwXnJRS6uZ/
WrH123oM9M5lUQii6Q2w35fNlba3ZH17rkMCHQ3tZaDYGd9PaqjIuq6hKH5Svn7e
CUvE4amXVhIIgIAK++dGZB2DquYMvAsXogltl5z4MPYDoSDWZE9FBxF8j67itCAw
orWbODX0yE3y5E9Dzuwnj4/ka7P+OmDCqK8802/I60xt9bKcI9/jNz3tQDESAPr9
Mg421FFklBlCoESBOCc8Zt2kEt1t6sXY86YaaXPUiImyM6BIBrzlFXDNGqL5+bek
IesB1FzYJMzhXe57ndc2xbqYApaCswXCR+Lr8gTlOlhL7vW3KRSwZ8MQrCxrgCAg
jlUbAv2ZayCD0tub4LgXZZxuB0oCCSLLy+C51tIjC+cZcwrEB/wRUbkPMMO1WgAJ
tid0/v+0epioRw18uUBEheJlKOR30OIe74hDt6kzTBqSM5SZR8WGrNJhLYO5Ue/p
jHyitMOG2aun53cYYfI1xKcDF+MsgI1nVVVane/iHuJIeblTvGMRNX3CCoGe2njq
mr5hYx6rEigKpnpKdZIYRB0yWisaTG5ECaBORUiveSmkzFwX4TWnuIOif/RscZuA
/BoYHJ6BdcWogCLqVPDWmcpg1bS9NMrXx4rSyS/OQnPIUduyznHHCa5ULbv1cKeq
4/J9GatkYv8yri7RojBzv7WgCV9SpsNP/B4+eutZ3p6BOJ777zS/tWr0TR1n1zBp
VwgGJdWDc6SGmFK2YqmyF01D5zd1qBrV69+YJA1eagmyx5ZmOSHN1QHjVgvJ5YCF
lQmjWuC+PdNZmZNSLKBTwfps46SXVpVcWIpHlN5tnF6bZ2ZWAXiU6IdnLBNFqRCu
lqeWeB5LDyCGCiIpzqnK4tLVduY8XAZrKPFa0f5rJAo5MZtETMju92un4MHTIiZE
QT3G9h6NR0DW/6IpVqMCQmgIo725vZijMYFP2a2m6GWbNZxhRQtsQ5bbRjvf28WF
a1m6Q8ir2vySMoGTb3gvln+dt+TIu/p+bk0taaQubcpioCJORU8AOk0vGt8jBb62
6DidbpZdLo4AAF1OdVk9gbF5V1/J+nSb/KPjwyM8NGDV/l5q/HoegYaxGCKs/zj3
y7+GJ8owBEkC4dDf1PGjdQWg1pHMURGddRCbPywkQNAIfmn17H2drjwumGDYAx/I
5mp24zlryeN2/P1ptKQXL1CZXjRXq4k+903sIploRc4Og+ww646Z8oWtjfe9C5vC
eJagZjodNbJMvClkGNF0LFyUVpo1jPqfHXgK91NccZjqGTS8d5Pw1RslufWlCi3U
aUj0zkHD7bVEI6Gkpuz7KYTCgVDDHx9AdeTe5MZh5Cjup4/zK1DOxEj62KNCNs79
NHdwfg/Gb4Xsmkr9k0dh6DuYJ7q/zH+Rwqb/wKAvgLiYpS4Sd2u9y+zIkV3wD8B9
8WesW7aRuiv058b00QJANxh55yMxDZz6s5SCigv81fSuVoF0m9IW8/K79CdBaAzo
gpFmKlbyFUScW3bgE0t7tgODmS4zfkOBLRlGMY0rk5FS402PEk6X4oNYWEa3fUAF
GZR/reFsFARCY7FwMo5C0MDk9qHdrudCspvU/mBBaudMj7HY9fuUThvZnTqxoc4G
v5LCTqAwuhOCIG1OMhk7Oyxl2/HlmbkX7Rq3ICDYmNTPf+vtHvSeyoslanA3myzA
77Y8S1O5PcpU11OM5NcwgOquTR9owkWGFHc1aAueavUTNtpYJNH25hT4rkeDlwp7
6iBbm3i73NOYTlB6f8booQw0hZu1ztdgFAS5Z5U/r8XYu1abN6/P2T3fPiahIziF
jjubFuE67Uq5ZA4p57x8NJcS7hpxmr7mqTuF/G3VXyq6JwAQLmXVLkae3gzcLGGh
JiXy7jojFK7m3NVx0YUBqGao2MmJbVYDCwMdjIk+yNWuvjK+INvsLcT8votH6xZr
FbuFeCZQQwYQ2fSY0L9ZAd2Q+gwpCLQqFl7dq9MrK6m4QWgFXBHR9cwO+ABhsbyg
PLctHkIGp7OfW4IaTJdBqTwwpkl3/6KyB12bGEcTuQ+j1ry2Z2nLIGXSbLa4jTTF
QpLofwAJETHHptyFfoJmrGGVeLEM8h8yObJo4aFloWN1rBg/MoKcYloISZzS2l2A
zJJ9/mvQY5Cc8o9atXQ9CI8O4QXcWXjQ0gLA6xeAAVurpbo5xFhA86HTF3hfYP83
rIK8NiJX0uXdQnftEiuukXYS02LEqT27d3XHFj2x4cLiq7Cznm8eT7nQiPlSKBJq
yG7Cv45IAQLjGpSMbL/pWCbU96Ovilv2XAwKdID1fRZvS8j6wwitH/LUd5wbwKO0
tqKnSCaYikxEVRXTTIWLU1HtZV4/CWc24nCvEcayZc8ae3UuBROL22xCOe4xJI7z
kXEE/GUKI5yhfIopvRvvKtEFPnO3/IrmmvLEd6Y3aH+w68UlSlI+P3hvKM6YK/l9
In1MCZGL5QfBTuXOlFJW8i/rEniKceKzeq+VUm+QZRI6BRutICowHAbk6//XDMVy
rz9/uc00ldU8eN49rV5pEIzRcDoqg9kLiRDBhgUCNs4EzSQ6ruwsH5lV4JJTOUXe
LRdwFAccTLChPBRoIywgBfy0aHw0rjOZt7Etg3E/lhu6MVFsP3NXNlNviHqUZIAe
9TcLb99krRX/vZmrHYVi18eb1CJ/RqxDGrysrKBf1WqvLDRxBG1qG46VudG5M2Rw
Gd/Cqyj7XvkVOmAS3IBX3nHg9lKiZIRfPlPr/Wh6guY/hcB6/vmQupC97VJ/xy70
zC5FckZbCcwkNZTc6a1idfJkS0oFQX+4KYMrnM3amOLxjdpMRtuO8DQBTffUvBhC
VyEzirVXTkLdNohBMa34+mOl4dDYdUJ/X67ofj5yAXhMbr23XaCFhtr++NUOfAr8
MF8EEow84Uck3jF5vq7hmBiSSM+jbQFPz9Tqd5G5p6gc1ORKy5dLLkYWlyS1yRRC
3h2+64etFV4NQeoMn5v6Irx9CCQ0zhqYAe/h7rHIzmD71AwTqiUUXLLdyTFmiHwI
8AwObWjpvfi3R1bLf2w4U9oNwnem/M2awgjLDQbF80wZ3WWGjcIgNWRaJp+TLUbr
FJ+06ov/xsr34l4+r51fng2HSdzMi/XqgeA5n7j2jeAjDdu7gUxUff/kv8GMgIHh
sXDgGq0RxHondX3SXk5hbBfrfqvAgqOwzzuNf9iBsij+CcOYXJfB/xB89hpappKE
lfKuHAXjHccjgd90Eusm4oTRvoRU7M3enpvV+lLY8HO+/uzwu0/kzLp+bqL8Boj/
vWkC4bmFtuTmcQ7beU/aUWLxUQU30tc2hm4A9xHkUmgbBLDN5yBF1JHBBmtwziBK
e6N5tUwJ8i0vO3mfs3DnJ2d2yFIb97n4q3GzBdVCVodXzNXu3uhMX8yrBtALnwMu
TsuhvQg9T0lhz2b63BGMqoph9GmoP4/6HqPytUZNPL66+MPcLbiSPtkdP9n6K4kG
lj1IxXnEfwC5PGtza/EfbgmqDCaRQ64z3HfUpCGT/64ux/z9aLL5PlFUucg3eYro
R+zEbH2jRuP81ANMoVRmMigRABa29c3LuXFjG4L+joYRB6gdETOrXLLJkZXGbT8p
DW5OdmkGuxuaLzyjSfx/XTpMBq0CJmU62OHfbqLA5IgeQiN4TWis/iRkwF4sxyro
YsAPoib6KC/LTdFtaUMaFkbNh1OpI7H8OWemRve+/tlZRKuKzxSqQN0AojHTMy81
vZqEnGEY5XUv/WnMg563mcD847gHyc+P/J+ie63Nk3PeKbOzl+fjqlr/eOo1jmK2
Uc2VowLr4CA5PG0ZjlmqMu96DA+Ntd+FSlcNKlO4jp5znWEiAc+BEYvdudrfAnoN
EfJGXsM2eY5llKHsvhAk+Vpg50iKpWyHUTp6ilYGyQpgucRaymLZx42+RqNZAqvV
YE27ck5uW8u4UKvqOHc2Aq3/sYwkj5q5mQVYF6FJzAYX7Gr2IuFk8oINSdFHvBth
m80g+lyEodsr6IQI+vp2tm0Vl52Tk4heZe+aA5JJ8EdFSF7HB0xWPg4OB305tvH2
rDlla8jaAWSrTr3vjVv1sY/u+voLgufORvgk8d+xPtmWih2FEDunJjNrcf60TRB8
rp5ZbhVnIPRrioqEkHCgKgb8W/4K0Q66BwDnX9dBW3DQKTwHcnFHpsIz5XBGj0G4
+jKRY+OJn9MpwvDdms6vfn2AO02YRbHcIpZQLZA/olDGU8Kn9fwOtg5HLukZP/ym
PK5TszVfKwlqY+C9b0QHROelF66jFm1no/8reqLz0gvYJJal8QXpyccOTeADz8CY
Q1okUOUSJG45AibdgFE8qe2Y6CQ6FsY5qreJu5isCpGVcMB7gZNMIoZvQ51eRlna
U5ittTh4coXT9FkpuyoROx3DDt8OJArbAsZM5uxLp4dq1X3LTTYAIbYp0YfcMg11
U8Ra7kszhnKP2BhRUKqhgIhfcE6+EaXKig3215mV7ZDk1BjvAZbJtAlptLQRTlZ1
dAZNJa6nAvde3CuZ+5RubV51mmyvdRRVC3U9JxkLDR/9rZeUbHBla6QjUMqzzjz2
5H6wJQhVCrQaeIa0G9C7LaxZ/J9aPYGYSrpcj63WiXLi3ajNKmzbHvsea0f/V/H9
ApfHNdgeeYFUvPC54C5eH8c6GdNTpYNOfLmyF8WEzTPdGTe3iCJoQE/uVAl4bZKL
2FJl+7gk1ZM8Mtjf/VVFoJB/hYJHtDqWptAQkMyr3Q4mq14A35oDD5GJfA8O0gMi
VHdhDdA7JVEsoRoJVH1M1zN+RD5J0IiSbYb0gF77tM8oFZv/JaZbJpoSiV1c4u50
cj0EAmyAIGSwIC981cQomO0Ugr2g5bjYo48MxU+veha5WbxDxCo2nDCkVy63/Lpr
NnyxW1p/4vbfW46+EYeiVG185OlNtZfmqQDf5tlqKvvVtTW5kVNgmjxrD83lrIKv
1t0412EPv7u63MrmWYH9V0jDQ9Ty9kyq+wQkju0+4B2yPmo2eDzjSBcjA71SeA/0
10vgWw6hsZhYvD1DyBjI5QaYOo/828Lr3/9o7f3OepjsmgsDaNPGPkEhqNbvApS0
VaLpTtYLSGjNxxf3/vxRreJQXZ0M3siuhnfkAZi3tZsYU3V94sBVRovdjI/LeZrJ
1o3N8IdU0HYh9x1mUi5pmqdqAhw0Z+wSZkKRhwk+eMVziYIprbCr/xQNhpU0QCU/
EdPs5H6XIJprdDqITGx6EzOcXZfYyGSmvql5V+B4Y3VjHp2t0rmbv7YgJPIdbFri
+V+GqoeTav2Mf8BgBH067LFPjyPzurTFlTBXem7li0JuI9udODMQy54UrPbT682Z
yPb5G0j01hJXVRkaap1BLGp9Bns5eZSY5l6GM0dMScc80ZEWqyOaXwyv5asphpV5
lsnTwn1xk9uqIZjcKgzgAqrR1q9yfGNG0OEc0fExylnOb0g6LQbF0Gg8OT5D+ljS
lVKl+dlymQo8t4xyR3Njd7hM8bv/tBen6dgPceyejGC2Von7aRePIBnyVyHPELFg
F0w/54grpn3WDt6l0S/jX9sT0lqylK5Ajj8ymLp6ItHLy1EduSPyUKebrMMWRPu8
8/hBJUnI8FjS3xhCzr5dM40oBPXL7hobSi89WoEHfbk3AxO4F/zvrEramNI09uYK
06goKa+2qUoLcdm4BEL3IeOkNv1KfVFVkYgBv9U0KAxC9KEKccad2bP07NZdxGKB
rUOTjtUOWzQzg0ykQ1bV/LawgDbWqzkzdyqm4Pj1UGJCbbeoe1ZsqzHayY6W4xjX
V5Tgey6Qx+sQrhyQLv6Bgs3AlLoGtboaI0j9scCt1D7tDpizF1KyxdLuI4HS4fc4
2CHjMem2T9WN/TNsA9YZggW/Qk2i06k/z0yPNulsIx2+FAwfNiO7QovSE+leBNeM
XhHh2uNLmiNKN4CwTXg2cxyg09uOYJI7B19tb/V1Aeyk2Wj6ZgJzmVcUzT+jVv+d
EERF/Fb2rvYUf/xuUUZa2+XA8qywy8ilImF8pZ48lZuLgNJcxcGluf/YXSykmj91
LD822ed2EnGksz9CCaRxa/lrcweGbJFXjdxGmKKoiLubcTS6rMBj5iYrc/D/8dPW
cn8QkjHAG9r2Za5g1z4cViDA3w6h2xbtBbTdsxjJ6LQjsS5/MmVM4A3MIe6Xnr9w
NAaPXM27fN4bF9/HRxuPQBVFQPZEcEREaT44EH1PjqqF2DVTlgAFE+j8pe3CtXrE
8mtOGM4OuU48tvbUzHPA2MBAPNV+akG4Vd5+4W8fhMYeK3/Vo6Dpt3ugayHHukIR
CE8GcWnUP+3iCeQpvEr+mRgROc4vzvVP3qq4jiAPhHqoc8dJjGarZcRXxmR6c/Em
cjYIEuEThjffWbRXuPkbN5ROagE5YvWZuW+sIMp0h8x29qKhWNXOpMF7GNaw3t8n
VAUUGwbtiCG8LZP0NlZhQ9ubghRNDovQrVx2v6SxIYmqERhaEbUhpYujQDNivBLL
GAGG3NCfF5doYwSDGknOXV9usrWJVdsf8QvkTuGyvq//TfJtxzRKKXXhPdRZWVhO
C+xFyVk7Ak4eA8D15Zc4BAegiK5nbjN9qpDaAjg+LDMCzkfcZXannNqjhKbhBGCG
VBkcp3KrcaSFZZnoYVcJw2A354xLJ/nz2stR25WNAjHMd8AH9mEwg+7v7YhJZi2u
xtUBuFfPrwcmRfHc7A6AmYNuVAtGdbfEsiObVksNZ4pNOYe8kYAjr2GE2lmmH0Bm
6mAc+5IHFaeZskpRF0QomthLBStee/CTjwf+I1G17x3CCSdBSVsTTn9VuoPL6Yw3
l6ISpMJAFoRrvH6+tXwSIcjTxHe6s6+KLRGROTSljTkd2xVN/geRcnQzwX+NBBSy
bEGwj8ssXNL71wN19UkwyxfuxQWlcc1OvS+VQj2s4oZysH9XbZ2b857laC/3/XkC
NPKAQPlO0w0wkHzBG+P4HXIYITkCfeBoxoypdcdcPTbrOtqyRx2/k9Hviu/3EqW3
dLzvQGlNoFF2jFYpVkN11K7svjxjV31Da9H4BpvPyBsn3REOMS+KgvP7wenKxgLc
/eAllS+nCwdpBdf+EHcCMX/NuKon/ld0TMA7Rpzu+31Z7DS0t7r5At0/dty9cA/k
S06MgzxBD3svQDYOs/pNzHmtbh/5a4fORAFNLM+lo+9OYwXy4bmRCB4EYnzrMEdy
yv+KGpfJGfZD56t2gYbtkwnkrxxt6JmvRWYpM8RFyCyTnIGgGIBz10KAsYVhE8pc
0gXjl9OtxFov/RMywfBF1/FgpK5l6y67Wz+6QmTC7PLepBlsGBHTS67aaSFUiSSQ
b7cWL/CI40/Rr8SfBZnhpGxJx9jvv066NzlUUki8IIS4AEzq4fJbEqaAdyYzU2dt
fTKZUkrJA6LptOrznlapHMxtEYFc8h5HzCdKYbnsGzSLctS9ATegZ+1fKbaOfnWq
J0nZQ5rVan5OYLTVCn63amEeomvbUT2Xrp8q8h+CT9/espgRkJxq0R1e7jfPLiP/
/L4eBVp2oTnjtam7CQxG+/SDIDqLc9S9GWqLx1pTAN84D3kZvPVvDoXmua2/gHFx
0MS6rTKaTX9OXk8h21xNQYn+OJ1qYGGzTM5DeoArITK5fnjvJQhlI2KZqwK2CQUK
8N3XpeBM5YIM7P08I1kwKSpEtf3sWA9knS6E89T6enUpV+rBUtn/L3GtC/Ex5BLz
8OR6TPVkrPCsWpSt/e8nAPRQi9lLb2dGksF6w4V2Avey8T2NpdgbqLoBu7Gornh5
YOnwF3CavO3FZ2TTgvjwMuWmMAXzgx/nSOiT3gkyC7Sqb+6wXLUP3Rh1BUDfcRJP
sAsfQL7pnVVvHYw/uXFxmZdyD3xliUkDPL8MF1q5sYXIVuQk+NjzYwGadm6o+JgG
mMcXRHxnrpZBSbAtSRn5vR20X+atRfyatno7J9MXSwD+Jymms8o0h+nYLp7Y9ZRa
ol8VrS1S22cwAjAhlOo1tx+ciDvMK3BthdNc1NiLEypTX372I6ANWDg9q1pg0nyY
6QwWXu47Bul3ceiFI8EzwzDOH8exnko3HOp3fdJIUqWaBdQjmgvq0a1KiHrRVYB8
ClEIh2mvqBzGH4Ncl68e6lEClEuifva/5A+yzLKbVAEdyYTMUqIrCFguTWm93YJc
wdBHUL9vHOZzBw45tFWfkun2mb2oqyLzobxmQQQK2b+gcpfmhQl99XVeksBY20EB
BExjrZOq86E6YckXZ1wOe5rgoLmsjDL4usjK1nmUci88RsQaEipYWsSRSuN3N61X
FNYRUQruEkGO5D4Y4J6iID3jg3a3RH6XsTh+Sxy2sCu/jq7GM42uMcC0qpEYd/Ne
7zfej/6/66O87sTDf7kuNil4vHpf9tXJoN+1OaRskX85QhHAMJbap9xi5L3/S16R
nNQFvYdIyCRP+R9TV5JxOqXCsOBcke7roN7LZwZ/UXH5ZmN8m0qrczYOHBIjs2+R
cxae7sXssLDRdQewjGrkDvLMAr7FuZuNcfM9SR6CjD2cjTN8kRZLKCrndCavuY24
N2c+ZQj72d38vXb93Ng3QJOlHP75G2SaS/4YiNMaxJMy+U1lN22aXPtKqAVSAX0O
fN3FjfIFLIseWyUzoJNqzTB2PNm4GrITaNiFOHwWh40gCfzbocM2sh0nxL8D4odC
We3qqvIT47jKS+rkGmsrAj8pYOffKiJxNr6uHY4p/uEEwARWOlKPSgJO/8VkGHVR
PZq2Bib/1vEOE5blOQW3stiwO24GV4c5es7BXVFBLwjigeZVgrlAo2a9dXlISBzM
n85KZ4kxik+HIK5zV1dUhr+Iw9YJWc/8cBt9TovL4nkPtcXdkg/Cd0L4k90amvuO
Cub0Tax80JxybEVoFMCPuHO0RFRHleQCwZkzRnvoYHFeivuTjwISa4ayw9ALVVRz
HqMRGumFt1PdMKcE92bkciGYkMrTBSArqRIgthTv5h5IxfccZWXAbvyf42oWHtQJ
/EzsGITgsYHzO0xV11VypYIE387PCK2zjP4L9hy5vijl6TUBzMXdsYSCm75a2H5W
c6PMJ7yruvVX+oBgfnydEGLkUEGMlCvETHGZZQGcf7EKUf9IdeSbBsl4jlzQ92pc
3TegrjqU9gc7N0pnKmYT9TsEuYrH5ZjoMqAcpceD6dYcNV8gm+1oUyrE3VhvQEUF
NO6JpOpOXXlW/PiQ3HWGUgFRzY5+JuQU2EoZ/SOJb3Ey776L9EM89BzGgN7MrP1j
pOn3hvqz0PMWRy7/YUb4IYL/0Mekyh4yADc6kHMp0Hxy7z7Evds2FnjWD4wNgtwr
3YgzzOzKL6K6YNZwLYbPYyeGBESS+kBO/piRaQbrrChM8gnU1B3gzT2T2hNjRMJu
pALc2+l2K0XqvLy4GbMwsPp1RXZBwh1729iRZqQMMJA=
`protect END_PROTECTED
