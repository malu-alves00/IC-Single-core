`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
msbqSECdzG4GFPgR1EwKbtbOIaq1fCkFQUeKUYK6KO09b47SyUqAKVYfKPNA8K5I
VTf4a6livEbn55Xem8/8pcuWDs3sZ/h/fTxyenppatdDodj+lFb2iBM2PYOFbEfr
1ZLQYh7gA/Pp3g+yhM6gUCj2MtSX7OVLyrL6WnDhEH94ruy5PLfKKHcx1ZZIzotH
LT0c7GCUN35g/ImSWUaR8cyEE4yaHNpMht/ew270tmjd61JCOBjh3iG6axPVPKoM
2sTIBX1ICzJ2EkzA4rLF9vcxk3UHFG8z1biz57OD6uAJBh8AwKBJ/Q18/I+l05oQ
ys1rh6KG2h2Q0dJRP7Pw9+YV4i9PVCtmksC68wrZsrvp9pa37rVl/Tw7ddpmqe5n
4IXSgG0Nv5v28j13sPLvy2+iswZ7lV4fXbxAx5XdINn5IpM89yrr6WBvwLRGeF1I
LTH/bp1Ae8qyMAGGsmeHLBU8cuNvxT0VdLe9aw+/PhtMWq/xmN+nWwUznGOqmiNA
IvLNc5pstMg4S9d1tZozgrH5qaxH2zYWYDoEJqL48hSgyjpEVpJtXXZ656DEGnN/
b30e0//JyeUeQ9oW0kzCsStkauYTdqHZxFLEHSoqQrn5DvidBmFxSB5pnTZYgtp8
OpRXVlmo4wxJ0n+JxJ7X1a6RxjMixIJGGVxljj2k5vpH3DAnudmab8Vzk3O1Bbqf
Cn3JI2pqda8Bhh7bxXaC7zPp57BQfwswSIadrxFtqJ4X7x8Ohm6uqjfXVxu5g40/
fKuNbg26nENvRdqSdh7AXr+od/DpVgGzpCoi2X9wP+jGvGDgu9rS93Sd7gphwpuK
iUFYqi+DlsrrbCMHnXNYm9B7pNYPszW9jS7667ETL4cfnU8OMpIXvNmgqi+EcfVL
7I2KABi5Eyc3KFoBveGHasbEmVj0OlMbmP/N1d9GymJ2aRQdNaXwIqoLP4BczyrV
skBaT0tPP+CfoRLRY+8XT1bOlGgkx9SPDOjxFCDBL0HItadJDBRi0066JiTrrzYq
EkcCjFvUnt4dGbDMSYvkX/RCFGhbhRlAS6ujRiPj4DE3TeLIhbmXbvIG39dn3I/A
wBZ1LNiez1UGCi7fOaeKyDyWIg0pk4GLekFldB5sC52O9WRpH9ciIppr9agb9T5D
NFqT+1Lsc7t9uCgkgG2522WQpoqmZ+nYQHNF1yl+XypBHROLOLanEo12sghpWHWM
q/FiiWzdi1xqUymZfQzvpfvC5E7NpHQBKduk0+C9A/+4Wl3MOsG1dDPUfu9Smv7f
X91Sw+VCNnDjHu1T7DQER1xUmW2dufLtafQQRqXPPnADxn1NhMWqcNjE0OK0Ud5c
InpbPm55q4eBn9C2tGJUBSktKJaM1gWYLd0yrkMVaYWfwACr+xKQCHGuizJ/0/TN
4k9zAywkKKp/SA40+nnoYWKwlSfC6/YuKB07FLCAMRkK2IW4sQ/PYB/MHvwA/lXC
mKt1rJPh9rGl7vp/+7D4i+hBnVt9rRJVhxd3xQBPkDOryNvvtD491VfdeU7GmwI8
mvtRrybqL2mDX3bCLMDSiS9sKyPSoxfyrfM/lA29lKf5QlLAeetaBWW74oqH9xSn
cmmoix4/IeFSaJ5zc9PWlvih79sUBkX+MtqwGmh+y2JCnr7siY0PZvq6uL9FXfSj
RX8K/2jZrn3HpFSRzAgJ6lZivA9jH9Uh9VpTFhuk/jFqef9h2vQcIxroF+ABE5MV
kmeNtNRrGzzl9pfy0qGSjWfpYXbNZsFs51grYWxbEXMsoIA4tK45PVOqDA9rfvDU
XPaPOwdLS7ea8QH6aLlq9F6o/rgexdBXZQMYdaoqr5QEUTacXmwx+hZ3UfbA5Maj
CyxpNE8kUZC5EnuqDE7m9rBIz6CrmLoUybdeysasNi871luZiimwrTX9b2U2UDDx
kC8icxx3uTNFgI+OYieXN335R2T653AAm3ZLeCG0By7A3hcla5aqw0XMR+byBEVN
5UBW6gARG1mk7MFj+rcuVhahOJVGEtRj5v7vs6NTYNwjujg83QDnJrqRs8F/wgQ1
Vq5AmXrZSPW8a4K573cW1YkgTQxxM3WFRQSg3WntwZV9OHb8kajLpXKDE6rW0bEI
QQyDpkBu2p6iffPNeTT8ApsXJTFcuyOmFTa4hY/5+MkhBvxmXr618Fwi0E4O/kS9
Q2vSZvoA7a1Cp+lYEtaIyg2vY/6VzIGni9We13RuZomxazLgKrQzCz5hVTae847O
sZ5b1fmcxOtjalK3/6G4J2T8O0fKJNc8YB50LJcg7UGBjpDTkhnyQ1wGASLgFA3u
JIR11rX9SaT4CJ4Md4EgiANcfPOgu7EIiY3Pvn25IJWIBBbuTFYAdjOAgF5R55Bi
OTNcAxksPqfUVI+KGXWuehLt1eCsAr1elIArjh9F51X4L6Y7imToLFLPhbVSyHuU
KP1lrNjvNn2NS+cuvCMVmFbiXNkzCSvuDTThGlXuC8X9L3PtQWhW33/hgauyhGtW
6XjXRV7t6GHKc+FDaXUBg3bteQmq5ulxnSqxmfpYAXQZ4x20NKBSZ/afTe8RRDXQ
hX110EhiadgUsYkL+fpQqXSFhxyakzYPyRaYuQXkgrF4fw8FlZJvr6m5w7l842Z+
S3qNbD8PSr1EV+jRjJty+1jOANuU6jQZshK3VdEYCTvhutIMJaYcDBx1NxyTDI3D
0UtmnsWC091ZpyAwYDY/bAVIYvSJ/8v3IpYGReuCjMNprrcCXNMqllE44OcGuips
`protect END_PROTECTED
