`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TqAsW6+FdMWHY8KxGaZnuliVjmoiJuIeMxVbY6p/yVQ1uscyHD2/Cgs2MNj1uYQX
GNtXjEpuJr54Q4QXOuhouuEmSlkzekdp+WN3mVDkNMU5do7lWg4bihjFxt0H+6U5
gjSiKPApcdDur0tQ3Irc87CW6dZ0y2xR7P7e7hjaB1ONjmb+n5JLzCdriTab5zda
F5ueFZ+rsh4LRgADFnV+KEJzm0ltR+QDU5jE1IaKAJatS4SNUkBSBY3+Kkm55w0u
K1lfFn6/GIcEj75Zb769yp/wASlbVhHHEMfkSDLwHWv5VpLyfCJVcCd4bzED3yD3
jJUKMKvsMofAHgz11QAGbITZxyNsGhL59iEHLQ08Wcp0Z2Q2Gp/6dWlcjo3bgCoU
k3iDTAdNYHGLFgPlNuVRQFEpR+pUo8wbB26BO+JlRAoyyJfqRvstZpxqcinyR0R0
NBGDSrFFSrSDiCEpIRjXS1epstsixQehgMJp1ypGPKsF0rbt7jtMmiHG+evJ54OY
/nwP3KclGu3wJBPjtQlPaF55/E2bhtOMCRZvaE1dZh76DuLiCOjW59BxBo5QdBsR
Pkid4Th/ggs8yr5Vq7H+tcGXP/peYSO+ObquGIO4L2spXP3Hz/VXPqiYD0QI8Nh2
WGyjhCzbjdVHEDo5N0JEZFV2IJuQigc2+sm1AUbPKEo93EEDJK7ztHz4bBy79mrm
UI5YECxLNlYr119LZKVcRv2dtZ3W2lQUA9VIkq1SxqkRCo1tbhfhLUoc5E64O3Ri
Q7r5WgCp8Q5yBVLnuVN2RKBg1mF/OXwLOOscDTbDpYu39zybexagpZl2tu3dB5AK
dcMPpBjEq/r3HdO9ULVPdcRALabwxmxFjJgO8RMpZqV16uNV4Yk9MlSWhirM8SpN
PG7tCMZFSv6zdhlCnBpu53ExPr4ARa6KnzVtQtK23T091tMk/yi1fas1KSrE61fa
2FB3VJe4zchY+WfD8ElNHRNkVwluMGnskV2+5+OeH/XEIM4v8ZwYEPVmSGygPmNi
xSa3XqxKTLghN2b+/VORNrxF4kgjDEq5f7Uu/lqBdhzOrarGAQE8MJzg/kZ25QQT
x31iAP8n/y+AkO8+CDHWi0y2J0HkMIzXRsmZ02MAHEbbiKmDvuPyPj9JjoteAbCC
nGd010JVfMgCTifPqp+FUCKfzSCMIi1hUJrsIydUw9BaZeLURpknG7J7BHshUBSg
AlvGJdB5Merhvbs6SrGG1St+rd8PDA/GBC/E88JxeHyzW+4qhKXunqLEFN6t/ziJ
DuT2SwAxM3zBGUKIR8Knp18vp0+hDlkbksoheZy3CFyOBoj/KYxleir9A63/haBq
npuOWPJdHmWvaxdioruX7JCMzX2GpTdtKWrWYxh01PTjV/SJ1QnVOQ8cUwhQwjGd
zzGz12icHBGIlSIIwjGeH8SczMKujQ+qnyzq9oB0/7UQfRpWvKCGpRm44qo2cI0X
TkQGbHnRpIP1Pdhb/lMX5XVt8VsBn6R78a8bOB8tuJTdtwiB4rLBQuniuG15Xamo
DU3yz5rwwQ3RPKwoc/1Qtb5+T/Y1YWIqRAyIMXMbk1Rvno4KiwqmtTaI/7qXWwhF
UN/Ruf6ea/VbbcsRfZPWTNZGs2Z5UpjR+0fydanzrNYf9TrFPglrS36eEi7UMwFY
q5bMaJHXsFmjF5y3f4dGFeqedxIXDT3jaM+y8AoNIdbh6Faoo6zPWdHw7j45zxLl
wvuTBKAiIR2UI3hdPZVOy564L0ns+uqHSg6NzR3K3FDGeNAAePylOQBSX67TPbo+
JJWdrohG7uJfgRLgOYBnQw4Ba+cmSy8NGg4ithlZObKWFmUD3ECJrzvkcn1kB+2S
6uZ4yP3DLjs9etpWpAnsqC6NfIRODo5k14K29CXOhHwChatMYlFeHrVu4lFp0PzE
s91lILyRit/fF/j2O4UhGGhPLCh5w1ld3BovTYUFP6C34l7wal8XuXMO4lzK4IPE
rRwaLOpccu1DmO2aSettRBv0cu8zyeyKHakP8stg7UdkD4+4tZHO6KQoac0VVxQt
UfLr322IFMR/XplC3S/DCOTS77Nt0dBDxP9bTHOBvzkyKlq2Xxi63E9eTsRawdjB
T7/aRm7ZCxajT3X6pB821ZRJE/z1wgKbhBUKz7V8P7IpKnmW3aY5Dc0AV4YJEn6J
HDyPz5jz5HRVASAM8Tj0+tofdTicDZ/Ub72LuT0YcaiGJu2fcJSEYcYh174c77Ib
xDHypEYwCxSBUQkk5N5U0doaaVV7/k3ncBtUkU/fz1FGdwAWUdFBAMa9s/kRbWzf
v1bI2Olz6XzR1krI0AzdQFwkH0CDJ/tuvLc+g4C+4gg/MXHuxoXlSMRuR7qFO1Ky
Soxqp46FxxxiipznaPW3+7hDioOxyZBS1gC0ofJz5AsJtqN00UY37yLasZps7v2O
H2jd+paKCIva1UT2avEnyWc3KfzE7T13nIaQm2s5idqWs2w2UMv+1WbRe3QHobrk
WoEOf1R5iFDKttMbtFjS1RenfdkAJ7r3setF48PrjiJa3sJdnwYXnNdiRA56ayQe
ihzL1dEBdzOYWnrEQ6vV0Rk/BDtb1S5mrebfcdPGlcWnq1Tiy9d4TSeMKDyp0mTW
JpOE2vZgdkBp5SW/OLFKXJ3v4dPyGONeGwoveOM7ehLsKg7UJNCJsNkl5fbJIIhQ
/mbwdIm3GqojmFYC76XxYtW1Lhr+fzOboYQp8UghY4btipbi9RkBUv0JCfbsw/X0
BlldkpY86o2iNyJM+mT+DuR5UB6SJcPIBwDoK2aGX2vNu9c6mShr50bbf/yQTQTc
IeG3zK/nSDeDnZsSpyFjsaMOv+2lDGwzVvkqZuhk/m+n0VsVWf82imXmkB4h6Nb2
mKHBUqro+uDKhB+wkVoRpyvi2UoKz9bQF0f8gau0znomtV0OMI+6JxxXfDb590q+
fzesZuFDboTAgLT94nQSbjdNXeB8qA5GcxcRklPy/7sPPiH0ZHfnYMYqrFjDH8eI
EO5NtwqV8I7JdTszzNP0PBjjUIb42/wjHEIoyDOGTKd8epv/dh5CoBCR9/uc3e3F
xtxHJVu7IQ+nZKUZAL52YLt70UK90pXubiEvgkqvajIRpz5omLBlkfcSDEsvOdWl
/JEX3Js0PiugyUWSKa28BHJzT2yUd/QrgDkRqp/F2D6VRJ7Z3vIgp5xmQoGqwQ9X
x1Jgb0+E8rrlspOMhOnAeEO2Q2u0tFVVMYEfKsTK6d5jsO9GPrNQ73OKj+kdrjRV
CBT18CpAwi8usjRUgWrunXXpfSdeKaktZTnndIWgqd6lxulNudhNXASM8g3qe9Vd
0476lR8gmqqZvjBXYhLq2uwRgJjTlQHUUEEhvGVwXklMchY99sTEKFkFVrYNRypL
VBiu9ncbMEu8t8czwG7gOWuRE5ZEb/yBTOA7I1iGvLMfTno2sFQ/aGXReSLNq4zO
uedv6cfqDsrZ31wTH38n7iLk/gID8xjAYRG4uGfUZLJZfDgBWEf25Zjc29OpwDki
m+X3JGq8ytz/3jHqMVsPnSMME8+7ZlDxVg3nEPGs5qDapsAD3LypakIbkNsYYzpL
QCtNstLYL+QTEMfIGuFUbxI0pmeIT2lHcfOZp2FljjhloGFRGO3miPQ4LQ5/D6eW
nPPyfFQCuCQh+53J/205rDsZVWIgy02oOYgPXFuCG2Qdf60sP3pikbg+l9HxLG+C
lMaHtMKi5AN06jwqg3Vk3ApwAsVpwd6LLHlHskIMA1UrcJpmHhqZowzLaz5uP38z
hyDCJqfhifrg7EhmXV1o4zjp4fZVN8AJCPeXACctWsgRRp5hNJFMh4QTuDAEsh3T
WeH0ODbOV67hJ7dngmouob/1JjOI7IgyRYOcwpilVXww4dnxKARWyE/6UUFrnaoT
7ECiIcmNp3B19oBSl9M2S21eTRXV8EuvokokUeK0LWm8qehtMwYQYnWNNb6a6NSB
b2Z1xwHc8fH4KI1TiOVuubR05v/FDdcnr0xhaqqUDckZUuOrYWgSS1eSs71e17TN
GkkHyPnRGPp3AHz7vEwsSYprPxkd2TIMJn+dNig2EYAnkjYPlrbfwPm3LrtVabID
emC0Hi+ruS/rmikUpDGtCDHOUd7q+3zT6dc4Tx0PTKttjl8tAmVLqlbW3QvJiuH0
81xgU8heDtbzfEHlu9KbFAXz1P9MDQO1ma5IbmCguNMHhEb3JAUlkkCs2bG6jb9n
v2kZS9XTJxwbZrBf72q+tQ==
`protect END_PROTECTED
