`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jnrpfrcz+XvrWJj2cEis+ziUBtA6vMnMLaToEHr2kIG21A0CpxfpIuJ5TWv4tm4U
xMRdrH3AdVvOjCtJl2Ejb7jgX55SpjQSVFiZuiCxBizyqeVuQ2xA62Q4yrpIKO2N
X9gZ/ZnzhMtreRjIqPwT+M1f1BVBl72B+sehmDnAoWD+QM36OfVyrofbudX5rc63
KXARfsEHZwb1nuTqrf7eW3EprKhtV4OrXckvPnzgQi7mB1qIFU1F+2JEN0ZU8qKW
U2CH/5jekUq4gALF1ottGxsg/UXC7b/NFTh5AqC2oT5Zs9zUyOwd2ZcSNy9Iz5PA
YtljLYW+mlmPrktMKVm8aM5wCnsj1VP+Fx5SuitUVsTkxDL2S9RYkPM9AG933nPN
2eXAD6ksnarY2vpvEtLbIBsTxOlyL1+WcLC7Tk0CcZyrkVGeoMQz4WLdhrWjRwpu
fsE6ChAIIdPR6fgST79SVNwfOuUeLu7aHvNaq3a/lDyn1doR4AMQErMoxHKi2WGE
z9eduXWN7Lje8bIicbsG8TAVsI85v1XdAG7e9cgN0u88udvktQXQw9fBbJ06Sjmm
ezLqOc00jjp/McM3+0qe3OU311fkubw4Dt4lFuf3k10+mJcFQlawdDzuH9xtbA65
b3rrHHYpUDEpfyGoBImSQeUJ3umxlEQpGlNZcS1Lbu1yRohBqzJsjH6LDtANzmy4
AGGRfA59ao5wchxiTvW1ddI0FTLGv2cCrSI1vq6jFMoXi+HmZ1xyyqVfLs26M9DN
/asyKMIce2hcvDjXE0DKsKGBH47A8WOl3orkpxfUxFYbM0tgt9Uh67BS6MmFSWpn
cMXXcd0ITetVIHZt48dSy3riXvgrgK1TSrgP+7D25aTxjXjq2d1AldagQSmvzace
VIjgSRux2PVq1TbXvczYNhSB6ocIRL2vXZvCQdiJEapuZuzVNi0cjBB7AiL0T4Ac
PT/EfIaoF9FbZ97qgjDT4oSRvW6BI1qTpC8oNflo3M53sRvK25z2do+PeDm+2vzU
W7cOdgL2ER7wlIAwItSLrLa6gphHFd7yCrpogOYWvQQJnybIx5sNEGLpQu7BeZww
5znfUaOvRmhxnxVdQ2D2zUyQpT+AVRsU7I6wPFpY2cY2U234V+8UnxZspQ6bXayp
mSnXD28qP8R36elWJ3pmKtk5eLxlGyR+jNb2H/KZb8DG85VYTPsglJY39xA9oz+c
t3ol7Xbtwv3tjToIQjcq7Rt5qAVLH89G4l0hhUAa+BJnng7SW8Kv9TAgOYIQAKH5
C1wijAL24jCgm8FhZsYis9Q2cVqN3UlGpT9Xe6kdukZILs7FaAKD6UrZgsNcLErE
wFQKUWTq7ln/G7pZfpN57hr8zo5/aEJW/5S95bLfF9rQiyYN9//dn1FefDq62m8A
L+KPkbqg1vWMUSVvXrcgTr1uPID+D6JLszKB6u35wBH58Qqcl12XkWd4LkrUYic7
5BKpe7F5+9t4N7UrRx02rrRxConBJIHRnvBWkvUpeL9VK6FSFVm3Kyu2FwFk0/BI
x+LYrbwYR9t5wzzp9pHOzKhJqS4rC7dLYPd5PAEtwVKTI6fQXwruivVHU6DJNnfK
U5MCRa9tU7y3JkUhA7QVf5nfvXwNDves2567yOqUfqMvgSJ9/wPLv6Qs1xYrJXTY
tbOTul4cMOHPqXydVS+mB2p0JtnJFVGXO5NUZklm+x0SRyDKb1gym3dDL1r4jJJ9
NphBOneZVWYAZvCBb9/8CAMCYz35kXm21HcIdvEg1hyF8kE9Zaokswxa0xRHBzkO
4G4QiAtXWIk2ow74AXM5Jg72ZXdu5fal0yIyggOtPEcgaR2uZVptRUR8uhTz/sfc
FxRJrlkjAYdBkjhDlZX5U9Bfbk3kpwkOtf+nHEC+98CP1lOhhHT4iSDp8z1KDihC
bXNFWGOwufpXXf1YrptRMf19hMX2+/Snig7GTSZVpTB2CRPfCxxfCwqfu+rxeoul
tBl1YQdbOQR8CC75+vTHC+Cu3T2ZKbDal0YvNRpTlTjyL/xMEikV/XQKHIOnVal8
D4ELmwrDvJXVXLj/PRV16V71IIU3le3dNxU0I+3pt0JyoqHWtYLelqs/5QpKGx7+
RsQRj8+sv+yUf48PBTWoNgzAXyk047ZtOIqlOWf6WJ5r7SXcjCwppctohFtE1zvN
bsJjkyEdRCLiIamjsoGmnmdH+6qz/o1f7m68lMq4p/jh+6Cg4BjAA+B7D6G22wpB
VYMmQj7zioWpfJIRypOfcskwtydD2exR7/5zwG7BphTnbEux89V+Bw4TnTntS1IN
X5E/4doBU/O1LFUpVZVs1Y5w3mkcg+N4BwwY63i7YelTiwnmYDkysSnyI7eK6QOv
EGgw2O3YbzsfB5KErWh9jjlJ6sxiEtB2C+EaQvFk8Y29ChZ89WjR9PbuhXF715/v
luNo9Q44wwCp1JwZtFPNn/+cajQ9cBWej5XgArMIJQlcMrqHy7pxF6KU3ewWKFeU
SoclYFsrcNWTFwyUfGkUcS1D981Yq45vNKFYna+59ojN7vXXrEbX8IvefUvnABgc
gnYpofyxuCOQRcPAd9WpjFQwMEBXOVy8nKwLCMSOwiS/u3rw9Dr5V2x/QB38RmNb
wb3KTgzGSejBQ4y6ag7GaFrixZrtIeFYZJwXJPG30oyolHiuhdkQhqnnbxTz/0lR
G4pObiBHGzhfILnRFr/uIVoNdsCC8ejw61cOa61+idxBqujiBP3rUvshT4/amhsG
hJnvpX5GQgE+pNxv1PLk9SSmx/fF3/ldpK997zSxxNbbyN0r9g5MAd6PNm9QgmOm
Rw1CHwA9mSxv4OA1qwFGu3DjMcw2Pg7ITbbHROgbceO2yje2J6yFHUvx+VFb4jMD
s7IXoueZwnCjCVJNhA51Fa2Ban6FzVlAq4H7DbYy3XfJk9mY30jj4wjYSmQSiz6E
DFfDBdMQo5u0+7X/PVp46YtbcRFlV94r6VKIQUqzbIuSNnEsYFcOLWYqSk40xStl
NmsV01YrVqClVwFNGNn+Uz7yM7u9+DQKe+H3a7RPbmy+ob3+taR+hONG6giTPa83
UEiO3gX/pLVQMFaEgI2WJk1s8NusJFMo82E2C05lgwOsD/M97NvmwJfDHr/VQqF/
Pb+P8dFIaNddvAtdj6DkufVRnYsWV0d1y3e/13nhmBAvHGcE/VC1WE3enUB/PCTc
Z3XNo72JBn/0Ui5Me7yjHr+BQEzh+UeUCdXXKN5viti7NHJONcRmjuiBmiJstSH8
x/5Y+MJ3IARdgqJ13rhRucEiKXAdO2Vikdl+JBrA9zpk8yBGpY5N7VPlmFt3z/v4
kHMMo1r9+vBPq7w7NakHVILjQ1ENzWawrGnORsdWCUTwCWWbm+S+asNM/z5um1fL
`protect END_PROTECTED
