`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hm+t2dCTysI3a8bCMBXyyL9ouOZ+e54scGoW5gZhQEEaRpuC5oJOpQVovakVL1gc
+GwcTYJUZhr4hjUnu6lysBsKuP88SRaNsTHTjvjTTIe0wJGxV5mpcOeGtyheT/TQ
aLNcSfAxg3Y9p4GSovAHnD+qVrPx0JIuY9fP8kkEhj/R6PxS6Ar8dBgwMWOYUnhM
a2oeR/vdUDmnkl4PXnmZPQ3BeJ79cBk9jfadB0L0KaHkhKGIaZ6kFNNjMXFEqrN6
Tt/BU20PizM/ZNOM+hAR8pjssTk9oPbxZi/YDaCKRGwQHfNCyXmJlj7qGIW6mz/c
m+X13J20DXokYSgaSB7D7/OlZXQGrw1kl+5eUQMdoIOauebKeRn7YJCwpWc4Kq4Q
twvKMD2CNG930W/RctC9wS+eZt4nNIQwVLEOtf7TgkSYoHQJArKc6tBNHvYOO3Kv
cwzuZYJ0+1sm5WJIughO3leTkmcx4u+GRbA1wT6hUcJwv0pC/Mwr5ZbLKgIdzgay
LM0IUTdl28pZkI561kq4RNYFnIB1WR+dnNX/NNB7B5zCSN9/C3A4ngIuMIe0YxDv
VKofk48usrO4ZVMpBspk8sXWhCTkp3G00U8mo9XbIG+8NYksuCNFd4WIl59ZWgKv
7gNK3fPXaPuc9PUYdE2oWe3XYHL0iir5OLabZL0103+vsV3IGZ1dooO1LH+/KaKX
PXoOdTj8IMOhLTzVSxicF6chmH8+gGJRAsqanap69vLVZuTncLsWyEvFxKCV9n73
QmSFK7Y2uuGSZG2i78iGKJmGkYxlhPKwlIh0sFupmd0KPS9pt3kOfzJXyE94QLzx
FC6W9pQxaGbemYr7XfWwICdh1oQPBnmTz5IIwqj30SbEtUQseSBtR9A0aMk2SSrx
OOBehYOULeZ/+gTR0v7wgSpbZCL2kk/wc4fLKoAYUvcnmsnlUNds8vsHsCCgeZ4V
A78T58RkqUingS6G47MgLknsMV+Kg48d78luhE3xXNvOTnPl0moe43ecaCCEPmZm
W4tM/i77nKjGVV6UQAHI3I+0+dBXWxZvevd3MDvMoaqyZs/AShk+k4vmAiiSAgph
7EM42hWCdrDaC+K5GWpeh5z2LQcEfnRTbwuEey35HWyzS9JfoSiPTorTVoNDlhoa
NdEn9FyOnxVEnoSyS+ELelTVAPcdRrnmq9LmQnF9eK/ifwzrGy7Omx689YRqbs0S
eCt1cUCdGfkbx9KoK7NZ+vTA+C2lXPdABe9NWe4WgVDmGVpL/m+w/dlr+C/aguLk
fHRtgBmT4DE+USpaOTJ8QIjTuHo1K8Lyd72LqfpZW2twA36ZmuLyW6UQxlnvBORp
ymB4N8qRnBVnHJhBg7ORfgL5VKpsDZYdmEJs5U70k5OZeZYKsDpHtTR0Xc0NT9KJ
nXGqWAFNyF01q4Wnyn2JBKsW+SaPvRiQHliaM9PftOYQtKNQniH0CepNGoVV0KO0
63AKcFeIVldWb0U7UyhkT+ntSZyj8qzyXTG3snOdFRsa4hJWfFNNB882Z2tPwErH
zIVd0k8u7z2udw+Q5Gi47yDf1yefQIArJ+liOrytDonYZGLtqmZX5NBtVc20QOo0
/ZdPkWX7Kw2zR0er5Gumx/z8dSPe10w5XvEnec5q0MM6XwWVB2xWSoTR8OYgdw+M
MMSPf4UgjILit36r86wDpxCrAZAdIz1smWlXw+XX1VfGIrKyZ7Q+HyqWvgrgnEwd
ns7naAUuI0/bd8pQ5p7Ubzw+aRV/IXAXHDv/xq31SHhsEYP8gcVz18QxRKU9tsfr
mQzpMfNxgllbasBy7bK7JohC7spldMYF10SuglmRTsXOCeWzbRPwDrw8ImOS5PzR
BKQW8VvoI807sa/S4ZaX2phpin+du0fjpFcUgrnZ0o5735ZRCMlTopL4Hlyiao94
0WHCMeP9iUnumBBSgi68BDOmznr7aiB0YPZkCc3Dv+9M5JitJ/axkNq7gqEvEMfd
4D2jl1JqLbw6doH5qI/0+Llo9UY5XHXs+LWJR+TDgeK6PuEisCN2RHIVczy9woZ6
MxzUMmfRVLQSV2ClfAjypLR+qEUfEhZMfyWUfY38xl1GyI03N+Pb6TE/56kwftzz
5MyUShLpA57dx8KlljfktFBaShrCkyaM95HC7Fara4QMMkI/cbJSBMavBE3v/wmb
8gHfJYpKyvp22wy0vEmg0gdLLqAdzxzazsDZ/k54uiUAORO2EUDp90Y5lLr9kWsv
ed5oKkFk0GgHZTd1KkepZz0RVH5Aljn34/i1Qjdh1qjuQNfVoy8KdPX5Pc7IJHu/
0ck7s7+ot4Inxq0X6+P27RTAbngS4U+5k5ugQe+Mbl4pTPxeG0oe7tkG/+LwW+Ur
IO+AZIcXNtnrd6ZVHr+O15TnopyqZw+Eah6w9E6YAamEpnrnXfMg7M8xla8DysrP
`protect END_PROTECTED
