`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5v8HyC+/U3kShPkEOnehgR8Ns8cLIpdJMoVVKfYIB7iccONQ6KK6XxEOHttuw5LM
49NmMLf3r3j0alOXpBBFEsq0lINWSWSY2HkxvYuMn19OGHNgozDBmX0AnHjNxa0u
ZhRXxYBlSkY1Nv5LO0Rc9GSd1Gsh3VvRgwM/D2OQO0qCSYXUY17qcMGRk68IrSRt
cW7PXMa+UWHPX6fFGsOBKB8JwS7Kw6cz8wYAsfV2mOjWwVcDKM3PjHJ7bRVhQvFC
96S0wlfPC+dt105q0IgecbJ3q0jzAgOEQ0Vnc4S89XE/jwNvz/0cb4tQU2MK4PMl
1jWv+fbkkszb5uyxwIhbT3YuzTYPlI1/EDmxmIu9QSBv76+ETo0uhKfUcudYtM6j
odl6jGhhJ5WLhPHBif8DSj+8sczlOHBIvaZ2XXhCsWLaEpN5IJDGJFwx+QAI8zu8
pjL5yqoV2NPzQeWUAr/e8CvsrADSPWuJ42eVzkSbGeU5c2+gOwzV8RhBIoNkmF+N
EAXBoWhkFRzka4IQd5XhM9giCjx0quwIpefX3gNXUjKUc+FGEbCz3y2SPid8LLab
B9+KqdqF0fgW0GomQOzvZq/QTNGkxjPA5RgUKUpQ2YYegEtRlRo7zz8HPAU7vPTc
Exxddb049qRtk/hFYIzlN8jkOiBjM8kJSQwgu2lOq1Mm6y4If+XjB9A/0LMBtgrE
KDzulYYo9CqqIVSBVIg+13awqDRNwhcZqjFyv9S8ao3o5TcjPNnJfdOlRfHyIKD8
53t5TJFO6Ckl8Hw0vj8b1yuwmIKQwGAFN4NV0fdLnl6JhAB9NhfG0aHAUH4bTmMj
eSSfbiBmnEV3BmADTStsg9V8+mEflz1TWAlskviDByh4/KngOAALXHBRKJWX4GqZ
ShPr7+cyj9k9fbs4KLF0RQHdW28j4k9hxuW6QicbSJ3qOii7YYtPeEFL6f3fR+XZ
`protect END_PROTECTED
