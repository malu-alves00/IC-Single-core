`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3IJlwME5ZJQ63ISU2VPlSd4c8fijU8prZlydZxPnRXdo8323IOPIfexvyqa231pC
Z+4sktS6FRDgAFuHeXKkrO2aRzmjpVKCvjqX274XNbsH2jWm32JBAjbptxdtdSSp
BF9NG0UbZ/sz7k6ZqLhoPPSUhXRHMCS1Va4FJ1s61dbFu3E4uLlIs+JosR4yQIPZ
Rk8S3BXs2fSFCWj/YXtMTFzel2b2PTX2kvvptQIbcIpYatGkJjYH2DqYsMdWaJ1z
GwSawVd7DWVcofLOwv4cDdSIZ/6YFTOqpncHDInMrO01fYaEICoAMLXCE9NV9UGi
NND0B8xw+4vC89GrfFX9bGSXo3m5drXlHNqFWaQhdhl00ZO7+vTk9Ozqe0lFAiCf
lhHfL1egebB0ROlADoHIwNKOCwMWA/xhnIkR3whw7ZKWNKG10s1yqyS6h7CpUpYI
loKkTBscx2vsolLkP5Huml839imgO5qHajEYFUkbbmfx+UHmi6QaG3nyMjoTkbgG
pODw+IZKfADBPBqnZuNeB7FXypnpkhKzB9Gccr1XPaGCjIFuInzTDEXz9JDOaWwY
lpUlu7vlb2ZoyD/RjjJR+fawoYwuaFBipVxM0vbeyt20l7GAvNarfrqmXv6rV5IF
bNQt3kOr2KIQwJUn5/SMo+BRoz5QI8n0vatZvNYB8XatsHYUvIWzVMSHTt4+CFOw
kQtcWT2P2LAXcHGemq8OkO7iZne4LAVZQGh/k905J4elNduJFYbwKzLWa2sZl6QD
1tMSbGfKiOerzMSG4vflojlgPJWVOjjmyzZw88znHuCSZIdRG3g1ZHtShGHwrikq
Za/bPNLzawyhYapsTi4AiYg+SxuwZaS7JddM8ZfkNP5r8K5aJ1Ubc9aU++cQ/qjm
X2Z6bVvwgOufFa6trt0/NNethXidTpL3zUEC0treRer3goRcnX9kH0Mf2aOQ1uYp
nGM7mlrqtX3h8JDMWMdARCThDYFF72sZiavuQ4YHq39ApH6zMcita7knpKC06O+I
3CDdOelrvya943b4OGSaiGZ16g2RTHUJqBf1h802xDwUdExDYVjyvvKkbv4ZIImm
mbRmhV9M/t0qod5taMtS5hJSy2vb0nYSs6dc7LjNiFFby18GwTelfToD6V9N3SaE
N/KsXU3MYEhapg4WSq41rjOVsNzipcVlMa7wfZdglMk3JWoBosha2foZvEcMHo5P
`protect END_PROTECTED
