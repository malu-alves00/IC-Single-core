`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FsKNgtbw6Fh3Pes1Yzya489GsTUmgihR/8f7q+TQ63ZlQ9D5beUXlhiedUC+VXB8
iOulSHedRIT5NG8Hf93hpEKoYB9Ntld9oItuRejRgQZLp9PRqaQ8n3iCD2/IYcLe
JOo6hoVNAQazrZpZTgc+gZKwTohsMGxpn1n1/aHx7zFiAvcitbfz7m6jdF63xm78
Z3Q8fxRMapODJroXeNHgrGTGYo6PYrpl7cdIoBFHzhFcsCwPaVsCptP36qWjQS1u
RTvlZMPMuL9gtZMYrwaQeMia01pYfYQX+Gvs+BbfsuIXDS88QMCETKZ4F5tCm+0N
fwvHXGuKNWaFnP4NyfT1d8xPHweviZwRsrntZJxado1RyoAEnsw5QdS9h9pkhOLP
Rew3AW0NK33wkr05QJoIbwD1/03Mq6k+K20TxqJeBVk/AptI1co5W61ahfSbZdKz
wwVWSFBvVSA8T2D+f4IJT2pD3ViPZWrjPpzqMEMwkuilj63GHdry8DXWVnFCM4cq
sS+5xSfJFPXsSaZEcOR8wmxvd40hSQLWekqMJMKg9TMdMvg2yxvxq8xp0xWM4qmj
OdOAMa6zr6xpkAIiTQP2q2hEHpShCAgcqiy8UwDSqsAD2RjEP2A87kz8NSy7HnKs
rh/ymoRxW9IMh82nHLJDZS/NOZ7WttmdSU7CZHXx7dm2TzlYI+mD3JmDMknxxa4t
CopRTvTz8QPpHsOiDyR/ysJu3auCAIuhZNcl2MGUlutkBLdSI4utZ9ZS0S2UjF/6
9aUdYE5BlgKRrslWQfBIcoznx+slVnz+dIS1rkTPVcrbAa1iWr1JDGHIcUXjObPa
hKxVNCz/Zf46u1W+tPRa4bpMPsX0IfopCjIgLiYRJHhDWzZVq2YwwVfjonaOnkac
ZcB5fnM6tfBM4/s/Fu3+zEsTPVjUR6hpul2ZRUeGXmAR6SyUDtPwMM/V3lZPo488
QwL4N5l5Da/2De9UUmNV0PZgFQ0ymQOMILPYcBEG03PF1KhvRrP8pp9H5qykLK+T
+YqD+yRbtbt+wr9ngtsSmJxFr11B2wvnfAi9iJVPAadhoDaacvDBk2KDnswRjsvc
KnU0IM5NXYgFK8CWML6PXB03iu7KSVRWYYEWEo+dHoPjlfcOjCveefzTjaljMi2E
H89mUafn/bQN+ehN3H/VtDFP9Ag7TD/CX0/xS1oVz7Ia+ngV9YFODK6c+ls2ivzC
Zgs87Rp0NuqbAGYsF6eVaPSe4oZumAgC/mNI3D3ht7SjBfVZijK72dMRFwAq8qy6
N4mY/xr3wHSCD8PyJrG5yckJiceRb7VDe/TT1BXhswB6wc6/errtwQOz7It3RoQK
TvzYYqjCQqKLZnsj6FFTatkeOmy0RaVMPA7rou4AAkcX4biEsOkxdPaMN01CHqBu
vfkOU7JbsbDmygJxATR1wFP96Mo4mkkcJYVILglQPlHoJNjv2M9O9ua+MLtDfaIV
uqDOSE9pRgWLQ54hu0NG6/IDMVg/0TqGX6RLGJYoIDrVaLzh/yNU8gRAC44E5OOG
+n7mlIVw9oTzWsUSn5Z0e/A66Id7K8n7pfLsdxIBuzk6akkNmaAN/PQZdYPycY12
Hf9ak3fi/SeK6gqIaOMjp82tfjhOov29PrqrnN4f8UXl+7wjKn6UaT5REN2yJ1uc
x9vO5LzTggrcuei9SAVXiZ4TSRTktbgKvxtDkWktQejt7IopaJ3KMf+QwrBixmOB
QvF268lXCoqi8ilx6R6fGDVWXFW2OLj5Q0L7044+illvjf01/4C+q0KDCRjECDYK
XIh7liuxRft91u11PCyN5P81Iu188ihmEo3IrmCu80FPO0Q5KpX2ycPEaGkPRk6r
qh6djRGUXs3IzIgkK/dTvZ6osCJHiMJ21YhOVFghk4bE0K+/elkT27z4slipr1Em
sIfblVMYFupM1qakzoHQm089DEvF5Pj5+XupFf1y18PcPfvvyggfSWLDff6SlyeY
d+40/TXUhb3yrUkoWnrfBbQhVMglSR0ZYLi5Fv1lYBjKwhjyluSZxkXvBB/X4Nly
u8Em4m0eBw4UXoFwmJUj/yUsNizO72KetWgG8Z25W97mCG7XcKBzmYfXSfe8CZcy
OdCqM5Mcs2RdfJ9sBKjhULhQcOoidIDqKrt2vk1qqZVJDW72yRZbh939sM+1wUJl
0ezetSaAU731gJWVWf7YJXCL9dwsPsoUbPT5OS+OgQl22DKN9e2LHtfmbpxNj/Id
Ao3viM1jfOt0ooFwY7ldyh1kZfmh/G2w9se5HzplTMFns8ut5Gsy1obKZPOQsnMO
L4TmAm79xwK3BdG71E1HIRQzBbWowrRWth8QyBtZ8e7kb7i8lpAf0pKDAagiLLpn
OxLrGUq4yWgoHoj/l1rzoT7IqyoWZKZZ0i5eEOBqVlv3djtLFigFu2V25z94aDA3
8E3by1F4Hkvfv799w2clarU8QjZJJ0pVDphEs5iYaScz70UX7i84/iv98v/V2cZq
PsSVmofjewcfNyl4AEMmaJzWBfsgrkIMWAtwocG/7WKdPxddQce4vDZjVoZsY8Vi
+J1+1PhRqwx2xRF1X4CBnL6cCGGEPfaI93ePZcz6z9RgNCVyEyF/amW4kWyIXSBq
5F6n1kfZgeTY5hGeghuTihffXMCXmcgeKweOnnvACBmylFp5eam/mJFwv56OuT4b
wlIY/KMyvXUmCDD3/A0BlAqYWEbhGgSESqNLEl6NWQ0OyUQUN3zcEl/7bg8qdAf0
IyTiD3PQcoUHzcu2jlaNJ6yWtepwxGGED4zBcoPE+z6sjDTKM+UM9Li4DvzqkfNk
`protect END_PROTECTED
