`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YI5v8zznWIbBPo4bhnvVbwQK6E332JAfx9XmEolzucE/KNcOOf2b5+eeL2WTRKZ4
8u8xNl/Wm5QDAE7mUQ3xibmqEICnvz0xTL+4LglcF+iJpk5tNvYkb6OWYP/ALY4/
tq5IqV59hIDirP2p5r9jhGRVJh7TPPUSXFpkX/wLgfukgCJ0oYWRfm09NxNGWeQa
ObgRva5OHCK7ISL2yC2o5BMKmKKdTll+pXfcQb+dOOM+IKOULmKFb9+BAiJ1oqfC
nnLgcHyj85BYze8OVaRWm11OzDgIPTA+LnTBzlr8JGvsm6V8m6p4Ql/dzs4qjB0F
F3cbi0jz8tHC1r/rtIP7jrnr4E7AgJ2ksqoM/RGv6CzxE7dSqc69ug98L4y406Vc
r8Y3BGX5QEgfEc6c0QTaWXOTbSyIqgpNWxvAlzl+bGHODqqxPbDAtBNg218ue3pG
BTlvgLX8mMMyiBSgoJowbxgGqdrSMzsP1HVYRL2GXbplV+YKowdrUTo3jrD9esDY
XGVvv+2DNSrAX3eQf9pjl9/8L2lvXFmuQHrkKVLiB+RUXJ7kOncZoo1QSSfs+1OM
HMi9cFHm5WKpfMwKsZaFQsJWjTsMhb007fgDJOK8nYhbRpuO3VEuLyRd2ltV/Xf2
lBfrmMGLg5T+78jFVvFOnakU2er38FJGeMBvEcawajIOIErxdAUiRZ9lONZMS6g5
tR8cEWU0qeGbMqmcIzqjOh75duDou41haqzmy+CVTIyGpz1RVNQxSkS6P0Wcf8Oz
Kl4/Opq6165NsDefvi2YVOUPZvVqrIIehcIL+8jY0evWYfGo3xbKEH/2h4hSq6rO
tIzW45AfR+VsSvsj1a7f50ZCZvVvA3KJ1P2qUPXl0dUz5izLsjigBJEpDHzH+gFQ
ytr50aUNNUeP5gosisXGUkRSD3Shdr02XNddZ8N3IpjXn6qUjHaJ7mPlyA96ApPB
71AMkE/nkaWdBoVd8oOPJUDSauRnF5nGeya6hoCLfAhSC67j75d9UVr+PgxJKsei
BajMVfq3VE1ua0x67DsVIYvYMj5W8jMqUVlYiPy5EZsXk0GGcZGWZjOCHPu/1AJe
t1Xlo5U4ZqZkG6ZgdqJO65wh2AshA3EL6UjU32MgYOxJZIlY7PVNxgQOMfkN4sY5
bsjQkOVVO78KhJeMp2Ib4USJH+IWl7/XfA8RGsI7bETPDMk0nbHhNBQcyf4zh/ez
FSXz6igL+xyQ+lb0D7dcoi5iD7vuun+r5d8OA+O1MxcMpT681cQIPYXnuUAvDnER
whtgmEzMADKBAzqQy8758MSK3g7HQigSD9JEvHOs++2kk7pmJ9z/38w3hK6ghxFC
mNBjy8bc5w/Y8DnkVgdb7/yW3H0nO0W3tJ4+AZ3n9JwLY887PnqY0KA7OjYRPtIY
ujmAAAVfyTjEJd68yV9ScDTD7foyB9GhJf+RqH9hoWCzXqzE66GLyP/TIsiVypmH
G4aeDYsPbeiuY6UYuuLOYrfsH2SDS0DKe0Y8gF2bXwoWralpb4So3rs0hjLCYP6c
UBgo5Ga7Rj50k7iBsPk7G7VeEROwjF9bGVe+ErGd2kOS6rpNAzF05HauRGVsAxD5
z5ItwQV0HWwfwTi01zWR4vqSWWjI/TFlsd55hXl1ouBeT3xwCAZJKvP2mo1fX5S7
VH9+yDlMYALic0q0Sk15rSyNShgZgTVhRMRyIrH5v8zQWSNGvgxKThiDiyXS/CcJ
z/SM5EuTUJbDOFyLezXZd7hdSwWrSIRmm9YZaPzX559YxDqAmsKBCIbFlBaQ26M+
vueWrSC7+20YutazttcCj/J6dUdYAYmcmASxzzHFJbU5n2q0umXchiUWHLKHb7P2
wQLSTqBve0+K/5BglqakC+Ihzy5T3O6yOjyU5HtTd4SaBJzY+xhGPvb04BLp4zJA
zjTPaTAiW+lXh1qhaN967MRsFjvN1lejrZ8WchUipn/ETW4fGqoRv541wXTEP9AD
N8BLjoCaCJVIPSOzhpM+tJzpRnx4E4dvhMq9k7hIdOtfzTjxB+kAQYlrG3e4wY6B
Xs6xxpEXKU68FewJuAgoMVVMzOlzpOKXOHL9riw8wqEcVCVENaN4pWjiDAd+ONoM
RWVhAUB4+OT/fCXO88WS1HeMvDldDR9o9tZXZKAL0/WSwJjqTF+E/i5WUzvKXpdp
MpQJVzfGrW6BoMJFQyeZZM3waCf8p7aoaRHSQznwcttVv1LHa2YtQLNmTcGho4Mr
nsBtptwyTLBX7GjCYIFyzgeD2nalntOd/bIpIFjHHKM=
`protect END_PROTECTED
