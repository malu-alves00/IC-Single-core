`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Xq9PkUEW7Ozijax0btzPhpUgI6aDQePp7Qb9sdbE0uhP0+bYujW3fJeW0+GDpvdk
itTF9RC1cPaz/fPsmsJq8YlsrqEVj+eRnyZGSZTFedHMqSPK3MAiZPF7A+oHzJ6H
XZeLSl2Kcv6f1JMeGOH2F+9/ibEgDahu/HHPHSPbzXsRYTrB9h4Nufxe8zdz6VN+
8k7lDaFK7QMQxt0joh2UH9ldo/fBmW+sVOaLo/F/7cLYaN5UZjxAFHPlSHNLTTeG
x+O0iFLA6oyz+/V/dzaUVT3eqxHSP73Shlv1L/DyM3e+DeXFirafG5NpGmcryiwB
oyB8UgoinJa1KVyvGcKwbEGDs/pC7RITgSGTAoSuCkzp9FF153sAWOGQv6P22Z5H
oM1WKpi5eNNaXlYmJ3hM14wEsw58j3P0j5Q4VClY3QxAI/aVY5YnlUf7e6GcRUYD
ck3NdR+hbYcdh81XiIHN/+mfr2FBp0kMdgUrPZrb8gTwHKMDcF+mHbaWNWufz1CR
ahfptAJctayiP2lZiwnRTo2ta9vJAUi4XSQ3zxbHpUOmC45r5YRbTD0YbgtTvDzq
5IDIWRNDWQrrTeE66u4apTIsp9O+DP+aYdSm1w+SnHPClkSYrEoeEalMc5RbPZeL
73njkOSMNL85TjsglTZdlMt0imyGbmmmIot6pdU3IQi7q/X8UFsMEpTJoay6VUas
fVJS/YiV/M6ewKXhmHwryvdji+dfwvfn/aDWPrc3OX+lc3Sd9tiCcSNC/y1s6XIH
oeyHYq2zjV4hYgZTXGhgxlPA+bYIAQCNPEfPrihpIx+xZt6IymFbqHzRfj+YGSyH
YKu8zfpY9ODSorhc694VdBasdels8Yhk0Q+90inPdh7vwbuuLTIg8UXuw9nHuE07
rjxlANjd1Hp7LSHvR34DJnVlamUmUz2WoDGOydsSz1Xq28H10QXHrTesFiZutuie
HMudARl8SxxiIRHcnZNsalVBWQimlW8AmnCBtz7QCTE4vWP9zcophAQrXvXqhvPQ
+3Y1pU0iriYut/sqY2C/RDJg2a2Ag8ERXAsNAopQ7lvH1UpQOJreXycbawj6Xx0T
u3BIrocP5m1cAJ75dcix0XDvO/cDvewfEh4DUY0GyaWvd+YsA9+p6JMhIMhvKi1s
TsC+fsu0GV9qBRTI0sZQodfy5y/gpNBEvbkJARDJgZOvUIO70HA2n18E2oSKUZ/o
2BIDwDzdnG64KNXSCL0RavFZlZicq/x5/+QT6mud7ehFFI+cs53XNvKgGahP3O2t
9NshPQ/1Fs+/PmTcLynei2MQHGJ6khLZLsJNNTFKmg9XMjdz/Ev66Lp0qEfF0L8z
5QsAx5ZfssjKoYUgnv4HGPDzIe84qfAc2kjSKx1euieIpKoYFC2wfRbK6WO7PJy/
BBqlib70KXtV266H0MkShGQM7lb0H0wGxUnd6vD16kYFfMPKFQNl2XFacIO/K7zW
2O+B4nEKdqk2g7lpPOY18L88dkVxcmcT+YyDLVYH8cpHbwj0gg2OKmSK8ClKbpix
Z47iWpyn1+dcUlRgJP4vBOZq8QkNYZDXVsO/yaFbl6uaCHiYPblt8hBJ5vhp8uz0
chPY/jPVh0wnQo4qcp5VG7NuTYWCVPYj8Wn9C3GHQ7HoiIkIRIuJUd3utCzxy8RD
lRCjT4YF035a2vLM0k5L1uKHBOW3gqdoVtD26ZipqXExDwQpQqsbOBxI3cfRYsjD
Vso6AH8b45i+GoCOrqVzK3+OF9M1Zkbg9k33sgLP2f4NkvjotgZM9FzPJrQOsfYc
S0ZkcYxrAxkYjcBwIoAyEwvDd5Shh65Df1DYGwLkK0D2Ut6dtZkBtJJVdZmc6vNn
1C473lrufBtI53e6/K/nmLnT+PG4hORkDryulyaCF8/O8tjn3xpeNSHqCNTbDD/9
uWi5fULMDdmv0r3i0L2oksVtHmLwlNbFdTEJC8QXX2QTIqFPzi1s5wwx0CC5n8GJ
TZ40BzTOuUwZYqK1XjX5i53rTSLXnvbMe05IFc3SAr5+6y6vznAHBIIsMx8icM0E
Opi4GRSVq5HPFEdzTXvyuk1aZkjqliimH6rfcndD0pFrECn69mQJ77Dvgl715z32
O3nXOr0rweesXl4EjNBKfbaCDG4UDQ/LkfB1qLjLfL9iVg2UahVVwkxIIX+kiJQx
MbqKGSxiRtLiHoGUKMyJUoXjVruN87RqEFcDpGf19shFtrNN7CLMij1+fwFtSLuc
omERni9a8CnwwIwE/5niRhLeA8xaT0HQmUMKjJfpTIsF6WFkH6tNpHAvy9g8xvVs
Pl5xCOl7wKVzegzJdGkrbFi+ZFJ/QiZaekb9ocvCJORNTwM5U0RvpL037bPYjhYH
W6HRoZK7SaH8yxklbSXM9xaySud9EvNNNqWWAvgBlKWodTSk9WtWi8bPtvF9KZhM
cYPXbycOpDqb+o1K17Ta/ABvmPEvozPLYqSxCjpPyYMIS0WvDDTBiNmhp/dFJ5qY
/FXhsYT5FMn93rRwHaMAPwpYo5iT06leOlaFEwawN4jFAi/EUlq6Ywut+b47YgEd
wRM0r4ym3G6kQh5Rm7TZg6yP29hsDLA8HGnLWMAmazOpRGafP8rMmYh/oGY18e9V
C2aIImKXi1sxgNEV1rgIoP4PGuXnXPTxTVUZfZruHzvf3VXEEAY1dHdh22caggGb
mGofeRkE1duEy+W4KXpwrljGaFJNyoBkZCWJudHo/eJIS7CgIRv/Fk6hB5OnNlRk
pFCNvcn79yWQ+zC2FucNb7MADZ938y7sxG8zm0ipHG832EP1OQRccK9Ra+a+5Ztj
nskC64OLg8D8j79jWlMOIYKHl7yNZC3bb4EFocnLsGMpj7YAv3BG7HL0OvT3QZw3
MZQ4dgtbqJb3dU2UuEpoapGPkDxT0TIZz3fppR1nBBxLa2WkRU1WZfM7Zvjbl51y
1sOZtzc+8e2V0CieDj+jTrSffPgfVQLENCoiECSUMLxvxrxgurVnTBvoiKWOXjQ+
IjMzJLLiZKwC6AoM8IgF9JEKOkRAeGl8d/9amTAD1kL9my1s8sW82rpkYspr4s/k
H/fyUt53E7O0woUjBa4DMNh7YF3966ps07TgGSImJGAvlzciY0MG2tlXUvPIelXR
NyCVnNSgxKLFF6w0ovYCqtmpmzD6y+i32u4O8HhbR8iHFloiR2oc9yY9qE+VbUh8
J2vj+/yhTLyrspJo9zdbGOxJeGqBLGBnbZv99M33A/8v5aCaowk274qdSvueHqY2
mYsCJW6L2APy+hzx42CTuHnogVrlv983Tj2n7x5fSsmNpzA9wvgh6v9hlmTS4VgI
P0xdZPXWP311hDUIv3F2PuET5U1E2eSx0bVo+nDtlnVmbyVDd7IXvpCOg72O/s2m
5yWFa+xJSvSc2Lq/NCd9qtJdnptgl7uH31x5gm3vCmZf2imphzOhilRDoUV/aoZR
/C0tGYaiQFsR4naFkaM2pccYtI6nL0v0zIZdrKp24r+kPW3M79xR+TOhfW5rZ0NM
vT5+zFDeAViDsAMKMsFDFA0VBHOmiWX7PbdcmEEWoTTZ8mw0I4prdV9yoKMMa1no
wrDBYPHKvEMR2cU2Gs383Q8gh8e5A5KmbiycClQHCCWA3HKN8Rf8JnGhK0CFrzkB
B2KAmRqTtRGwmnIVMq09B3MSE7wBIPStiLPyJ1h8eIvUsbMG3O6bZsC24J54l8Fz
ib1lalP0vjBXQtc4JGhaLlJ79K7AYefdQWaLK0840Z0Iuqm1hPdqjBx8FQx/jUN4
9qo7Omhwz0ZyzvmtW3a2KO1oGqk3iHttHqdmri0orIHhzsMpEkjlaNYSEtFfcNl+
rhZkOMehWZqYJDB5tiYVKlndTWPleSIHqwJ2i+ErwUdLW7K/dqN/EIuQzKvYG7r/
TiU9uuKgi/UxsTBIX9cATsMQL6HR9Y9kWYmbu47RsbWBNpOzHYUug5k8DaH7uXF+
m9SqWIfol35bLgCn/f54NLd6k6BjH7Y4Bi0SANpx+wUUMB/yrvBFU4EUPxmXwnUh
bJatZFyu2LQpzwYwADbl5pfFEqiH1As3feuBAlLksG/7OBV4s3aKsPzD0qjCAlm1
LKAacI0kZzqvCGnRkbdEWaf4ET46ls2rhcj8D6Y91oDlnBP0fv8UVQwdUFv/OG0i
Q92uM2TN7oFQ/86W7vX27mltbr8qxsOAvXth0w1h9Wav+3CVC3MNdEJ+sbZyqJJD
9vxnJot5olDoilJSZE23cNrScRYc4chXrnuH9TvUB72tQHVwtfKOjSIEMkPbon1U
/67oXd96YaVBtxrd8Pbi7s78f/S2PthlyJD61XD9P8TetqyX7e6w+sH592WgRhXp
hy03e/Oerbwuu8qnhMKc7L1GXcCXcSqp4yrGdM9Ura3dl2iDYr5ZZ4L84419T2P3
aeDylqQkoVmOZcbL4+a3xaUyzLiPuo2Y118Gt7WstVFZcEIL62DEIY58NvoUrDDy
dp4TRdCHm5J162BxOJHuc2dTCNSCy+uhulwp0v9EDsVahszBGCrMnm0m0BDu9Fns
10hEV+c8Z2PJmoncSonk6e4ef4lgf5W/IrapTAYWUBSKrX5ZTqjoyGfc7EH33rlc
0QOUWPTDgyn+aDWyzI+mXhvWBg3DD8elxvAvGUTcs4Pzko8E5kUFwYzADs2B4mPl
PFvHv4rPXbN71jSdNUUJHqvUw+6ihHZfmMQyYFdjFQ05iuLizWGsqRClHL+0bOjS
A5Fd3AnTqbIwQJWoCMUZpvZAbR7Skq4W6TuCBBJLroMtFOck/9jc1fxsoAjhzNaG
50ss5tNPEimp6qbGy0nPOrx9es1ZHwrLsY5/wikf4Ibiejs1X9vjqWoll5Kun69L
ebssqS/LN6iri0nwTWyukAlFl4/8X9AfKPzK386R8WzbE4SKq5j8iTSkN9P172EG
LSqcs1LcUWamUzztBubj2uBkIKjipSOh8KEmSrDZQQ2wH3GG0wsFTHQSQHwHTyj1
/yScnWLu88r0Gfa25Tt5BxTmrOwuKdCRsXGuXZAvQDpd7YkFYFbpux8h+8JVZ1lw
CQwdu6P4oNKeIBHB65ernikdJ93kCUtj0Xb+lrlIFdETde/zVKuLYujYL3swkwAM
ncpn9XxJTrOZE4Q6E3m/Vod4/Sqw7wMBysnmBGZBoVCxn03OAG7BRTY3dVUDyVKd
iwsp3+5snmmXwif5Ls7W9ZT7ZpniHNdk8+jSt3+Dcc/IIauP4DP5iNNGqxGVGio0
EXFycj5U61YxGE99n5GK0LoUWf1Fx2ZimYaDUKuGtrK6EeI2/ztKGYi12oYV9oVY
X1ISqc2jCh80rnries2/0kJgUGerPczeSTEJrJerPlg9sy0SFfSdlHQJc8vAUVId
3JJ8E8HdtGrp1PvopoivqwfylVBYgaigQoLrQNnF6J62EWuzIk0vYBO8Ty60tI/v
7RAKxdI4ja6+hN4tH6FwrNaQ/0OJJ++NAX3gtYg/IQMZU/8aUEsWuwEQahzSq/Gz
+ffBWzTvgZR2maQS7m+qXm0wMi7o2JYrOi9ZX8sF39CoOz2+8wKBDhK13U5afZQF
2Vl+qOt8NLutaDGwfpSw2erps3ozdFiKKrZoX8YocCtbvpg+be8O4oTlACjeCika
uFm92mNjzQOtluROyjTg3DDS0F3uVnPozEt/sR0BzZKU+qP5JILUXrzW5S9iMtl/
7/pZGiffaYxMvi2GRzv6Ti5j8A3bzGCSe7yEaIe0+6sVB8uRqcHVE90sCSiSfYbe
5LzAFxvPG9MOJtzDOnVveeBwKUnXkwscoSrMbCb7SeuM1z95rbV+NDPxQtVayP9t
LIz3EOTdF3vjYHJPCfwCSDBHak1U4AllrnxAyLzo1pXixV9W3ZYPJVqsX5fQ59Gc
OkC6HCC/70ObO2i0nVNZGd3giWmVm7v/fDR1GBDZlbUszxw56DQtX6KM1mfXALVQ
QYxRTDSxXTLkkT9S4BtiGO5iuFCw5MyECeCujGgmuNvFB9QL/wHBy3LMWae31wgL
Al5M9+zAMZupWN5mwRh4acHd5tpehmajKQuTrjlUR7Rj+/GG0gF9sMYSnf8dXuMs
KD1HyBrDIjefRkFSQWZA3TjGhYOqz6Xn7iu7cVlFfWtjXZ05QOJOEEESdecydxQp
oDT7OnGMgG+F/QEvxpW0PtkMrICMLi23gz1HTjlFTCxApq74tlxN/dzpD9+5yzo+
X3ZlztorhxOYoPM6ae/4zipaxgnWhvJtwFJy0Q+ZiqckfIy2rJPRUtdScSzfVIfa
wamceNs5EMERw9qefgK7HeolDrl6mYRh76kJcuUgWBQwAjCCzE0DrqUPAscLOQ5A
y2u0/Y4pP02MY6M/pWt3X3aVLmJWTvd8IvNmTzgs/mqos2eNa2idHRNC1XxGXK3y
W5A8PUiC+sp77D8X80lGsoWQUnw78rQ//bsQeTOvCrTKVd5RCASNBXIIfihXxozo
177rZj8kmcSbUo5BDbt+I+rSwOvfQZm3+Olp6owrAfzqfI11XgxYmc6URDR1Bvqy
NCTmsMEu9QhwYVjVL0JtzGNtiHHkeMJRySmrMXQENazFNVmThBPXtQCbqBOAGdDA
6dDJCaZE0jYlgYw1CzkSOuQnS/BKvCcN3V7s1+A+RTrjA2OGPKNXEDZCORTOwv0e
nBADy8hPVTQ/2Z6FTpu5uTsBpkCPUAE74G6PfIkY4WtnWY2FOkVKisbchQhExgxJ
1k39atAjOa+mErcjn8GPqtYGYZeo8oOjXJfJE+PdTQ7lFsyQm/p80RrlMWCc4vAN
OJvtBmbqJMxrjksujClUkJfG7h7EpRH8JaZZ8TrXvGVCzMECMpHXoQ9LM2RVhTwQ
6K6Sh3rvedWVO7gkKDKUktRMGG++wg3yrR6OipfSwnGDRyHOgxxCGQSZTv0uDYqC
TOVvPLXCqYfAqhudK233SaNjD31d1owQuST6ml0U/vcRS9UHfGt78mfNaemgF67C
gwgfHBDYaCg7qK+8pyA2mev2qWWV4aWHJL+LOf2Fh2/PjurklCnG3SN9BWPtM9wv
32LDdPU2LTWsL6MM9J3/2cSnv+ccX2zt9+NBatFFvP+OSTXusGjDCqrRL355PqQs
7eANTqxpArO6B3ddYHsEAsu/39jfDX+tF0CWKwnEIcOEbXwhqaq66eDDJzh4QaS1
HVtPJwReC8XRxXLm/O/yq/lQ6VxopHVJMSfejm3scwZCd0Nql9kqe6+QXPO+X3ff
GIdjbDFpK408DB/nlEqk/C8HGNVo7HE+OChhVxx0Mz6sEEVFa9umLUGbFyduFp5s
ZmKUwuFFFPl5V4FDRULaWW2HX5G5quubhtx2GzCUFRHCp2WNfIoKmXQ1fzM31eV6
TpWiecEhQFlsRoNURKhz5RBSwLoMc2EyTfYu/pog1IxltQiJYip4oQEXnEsOLJ2x
7GH5r+OUMu0dh1bkssqzTXo7t+4PsqnK7Z0xdQafxp+QZi23W53Vmf4owy8QlEu5
yVito6AGDGETC7CyY+VVZEbFvNkGpfpe6CELru5kX+Xs/nNFB2LdciNOQVeyxDQW
IzYAIUqnIK0aSeAl7QQvKSi/GHb9XLBJ7t3p3hubJaKnBALxY7wC3keGoZRE0DUB
rspO61RP35Zf7IJQNDxyadzYZ5zvU/BLzMg42dhvnrpkgdqPl8e4SfYqCWC+3Tkk
4Ami5tG3KrQ3tyVQGf47V+OAixgG8ahIoLGFdpJ6DbhVI0t7h3DDiZp4NwxCfeJI
3T0ksioMisv7WXBjIO5BMIC8znd1ou4RY4SNUqR5YqqvVpoffsYhxhyewLT+PVAi
1mhyU2fAXppwWA+Ji2G7xV4JiHN2nEXyXg5io+BIWZm9sRBEdnmZ20NHrw6IwZlE
YiCtzWcIY/SZ3kMraiwB9qAMIJYsYZyHMEkem9stVb+6nf852H69yaDbn+iyva4u
IT5GEov/ZbggQ2PzxdR5P+vjfSUNnvgLFU2LpyRl/QVmUu6q43cM1LZ0LrteY6l3
y7IMXzge767WF8xrPAi/oM37Mge22oANLVZKsW6rO7YB23083M4XF9Tx/RsM4YwF
cfTKew1cu0E5UTTmKgIpO9YoIWDM8n9lb5aYrTSNXGaSYWMXjHWenddX+EQ2Bn21
eariGX1wJEFuo2Ai95FX473AxghI3C4weaIPiPMtR+CtJuHYP3fIt+hz18lr82Vq
qM8RP9J+7+LPWVXUMxlnRdZpwY8nZv4fmnz3n2Tr8FJBnH0yF0DnywYXht7BPo+e
5leWalO8QfA6C/ZVkTX9Rd5APWQKv3iewZzcSyCh5SmIoDPFE0YrfDCJDJcyaNHP
BBkvorDfBzoV7Rbc9iczdL9NjTR9g2N/Cf6iZuqnLgJ1Gp3+YJmcCG95xjzkbmT7
nriQPcUC5BMuRzZL3Ktsx5KPXf48vGzJcHWzgJny+MQcodjJ0LMUNVPO4Ml9RryO
TnYoC0rNZHBe9TxxPesjmWW4YinEKoHl6S9kjL64d2qEvNK0+jSZjcqrZoSaPsQL
1HA4SAJoHE8GRhKlTDqAsBOkztFlQc0ifjwAbcHoLK9gIVzyZVlcooQyUFiDHrS0
JTi2n1wiAdY0J7YuvsBTeX6XdqezfhD5Jo3cxrXX8wyhCp91gQZh7bvKfmjVqXuy
b8tTLbgHZ+hikUVrIe5EAUy7QVGSS8JvAyev1q/lmqwcIssuQVrPQeRcsclBNqO3
cvDQ+xEPay078GGRsXbpTKPT8+Aq8wihP47CeRZ/YM6sDLspGANbNznJU45NZHvG
vhQrWXaRGtBnV7a6vYD/ySm0b4IL9+L7jLtenphQ35EnoYvVkGT4XwtYwpHvOSLd
dUG8p6zvhUfiukjwKJvnaG8iO+TEMDpW92UDUB9AEVa8Eu+RlDVdRQH+y/iWflHT
MbdL12S4jIDl+5DEtWJEdNWtBTctd0nr+JEpqzMJeHO7ziIN6bWK3ked09rvWvjL
O6EYRW72z92/FVnFkjmlwvfvbjmCZsuMWB/As8/5WBxQlN8m9GLYH6oRjOsioJDS
67vMiepmSa/XxdktSX+mDEzPG4JlgGSwIGKwNvYXlyPCYbEC09fQ100TeKOiAEgL
aUwwDFlcF8ABLQBUMpCUBpEqG+ALE+/yRZDeUREvsHvF5ISNXyiiT1UzEjmKAHHd
4dmLtdmhezBywB7MQ+vbJBMsRHXZGgLUwqopChgagRyv3GZlDZU3b76fGZY2rRbx
VKSRyytkSwp0msuznGykOXhNeoBxCCVPWFgSIklhMyaiNtHHSug3vKPgTo+hW3Ov
SvcWDut8N3dLxM+/Ckvc+L51k7nf1013xiUrgqCYqRO4Ezm3uryt9Q4WG/VgQ7ZD
+WmmhJuczCDsOUxVtyM69hczoyi9s2/D2LSY3fVuywt2wgCN0d4UYXn52gdcO+uI
U9Jmm6s2+kB/Gd8haFehuWMJZ5yk4SVVf978gnbBRxb8gB6vQsYrC4t7RMCLOC+y
R4+DMOTWdS+zzbgF1Lft2y5BXU+Pq9Y9+rooZk4aZG/2gaQE1lqDnvdrinL/Drj2
iB0t9Tdq5kmvft0nnp0BjhJqol4dGREc3+nCC3jmq+TRLO9taM93BqzpsuUO7rgI
0viC/YTvEbdcdIBrFI/n7yQmpboq30yJQPc9Sn74U88Rh1V3Ks+mu3Kg2xAjisuk
5wzWuDrN8L+XZjb7Py5Y6piiXWgnSI8OhPtuRNJi78iN+Bw10YSlfqG3rtlCZd7E
RGNunvbTKfywcXbkICMEg82rkgf17tvaHM2P9M0w0fJOFDIKDuFMZ2uMtWmSWxpP
yEjaYs2CNVjm1+P+S479pxxlA5dabPm4Cd6bYOEKg8GYVMJVYcg2tHEzZpFWqkuN
LKDLM59MYiN3zOoqjNmpjpXh6dE29Hj5RauqN7i2a+k96H3RGW2je1mlP9j5Q71w
wMEz4L6Evq21/XdrTt9FKcJLX8ebuXHj5vYDuyGWQinxA96Z6asjt4/RpmIYFqBS
yHbNpxyYdO54W1ZZvQIID7k1lb4fkcpzm20qOhixKrpg/a0KZ6lRYMYHmTcV4pN1
KF7lLUHXIAvk+jqxEoGWs3UkgEFTEHYQMHaaihqFryququAefW55dpqySqDyt2pa
EVRQ+buqQFQUTYZ1ZcE1NOPTa81FTfVAQST8rjb1MZNFpMhz1RfTHK/JcFq+wzYZ
v1ISaP1EvBmuSQzWh3qRuXx4B9y+9xeLaxx590p3EyxYDnAPXF7pbw0lQBT7qVGI
hMyOG0aYVE1cB5NyN642Zm9pgTLbdANgTWaHyXwElVjgbBIK8nTUkAfvgRXagLr9
NeeuOIXTPEKaJJeveThO8hfrEQMwm7TE0JcpIS7OOOCnA1lOawCLoXCQHxC4sBEN
qn6MUOG0ZfW1AsgSIzfgJU5kA3nToUSDu65boj1muQhdmGqtmQtnHqNnue4MzJfz
lcokZr6aYEBW8D2G10l/HIeKvkinqgTBfXo1OIKEe2EUdqewHX8DKkAEZaGFOycd
6damhOqEk3ebr/0GDtYIcB/jafZv9kOWggOasxd4OVye6zaxt1xs9KD28j/0OFwk
rMQMAN/un+DOY9Krp3soJVz3lwDS6VZzQ9D+NrG8mtu+A0E3yVU4QzwLjOqZ7HvB
z+ipaI9uPCKVZGl86uupFSR+2BFoTw7dDJN+2B5imNsaUGI1eQDoS1SPfnTLRLb5
0pBY5a62K3i9g03JTy+IyUNOQzoO3dMep0lXgUDp5hQM7s3YZL5iOkjavoVXYeFO
KjrsIqNh46iEPFwFus/I3IZKYhJFKsyD+zCX5F/htRZ+btmzqr0t+q1ND8z/lMNH
WDLV+lVSi2rTQfndq5FdUJase+Cu/aG/0N97X/14Dw6SKMbP8gq9a+TDf7vDAJc9
Mqkht4/i0KD7bfUCZsvYWXQzkRM0efI26J1jqBtYu7yA/03IgNfB70X/q4p7cXGN
MjXXv3z/BBkn41xP+6OT794ZS1V2GuGAfrpeQuyiLbmT2+N0Udo1VMH3bIdK43/n
whvTzpZWbb1IkvW5FaDlTV5SVGaYDcQk7RG1QFMv3+CggTo0DR6E82gk6x/I60/L
Vc3cipZCTTJTds4H+B5HdGym9/Ahe+QxwRLIJ9NnlRUdc4+bgnJ3DQQ2fd/dUKfo
XIf5/ULR/9nkupaAx47gEeiRztL0mT/5ooOm4RJ7ckMiTxi6LQl7NUbGklDTNv1F
wApsBgqZ/v+VpMLr7cpEwH+DZCyXdlu6gAmqynoL5umgwLoenH7YwTIApA3epxv9
SAEqEH0arlZRkUJKMpuBRwDITbe6i1qUAF7fcqgBAfK2wzFpkx0JmOBnhmX9OW77
uKpULAif6XaGiC/W/de2j0AvkWJGq6m5cCQk3jLQPszwF6a2fwGidAKfKkuhdbnN
VrBrO6bC8rcJrNSEF0MsB7QS4/ysxSEX3jfZVFkFu9yTzdCLTq0TqHEROS7YIn0G
3kXrO/7x1TpGOL4KZPTNQquclv/QnE4WDKqGTHHmO2utnzvmBgpZSKXLzLvPnks7
HaJioxeAJsk7df8zVb10dHxUvu+eOtEv42SZH12OyjCeZkuwR0Q5VqZ42f3ysHa8
vrvVLBAgLtjKbcCArX83dTb9o/hgdsgdt0vCNDTjybFXzlCc8HA4pwsNTlExJPGJ
YLtSKaOElRKKn6TEicxxEA9DufLFiySw9fB0Af3+Mvz2hnBGAHghg65Y4TA2Xv/z
iTy2Ey8/TO3DcKPUMis2fbZt2TfRd5aLo0YdYE0XYVI59VlBHw3O8yxMgM8aPXqL
xupBZ0BylivIG5/XE7cArHSGN6O+Pje69Gq96dX/RvoumjBXrZkvuJJzv0WD3pML
QmTRWRr7V0pSxqXYAfj0/7N1oNVZVw6ZpKS7x0Q9UKLmM28ksc7io0ID4+bCa8lI
NqI0WbQ4lyKxMbZuO/PuelvGxYIGB792dUPnhJzZa+rGBYxLO9zxoNxi00txZ0Tg
e6IBtYEn62x+JZ3vZ6eCnczFLweCWS8XbKsv610GtdP1Vbdssj8oFzvx9tzdaOLr
fJyJDcq21ShKMjEB8w4cKeKm7PXZhU6iislD7duWTkQjjgm9cKA3cGs9iYhF3wxI
YhVoGizDjFuE45xtKXJ1ksXqxLuHqG8qXPlh7z19iEoFnG74k0YXSXj3NSVszXMS
3ZOKxwFQA4nNMeKbDroM/wHDAp11gARCwyoY6pwzJP3J7ew3UD7EX6lgX21wX2tJ
d8lmYd/sbe571SU551HHMjlvh+Zm0r5LOjqRPL9gUPWgPG2mnuHbgF4yglKzBdVt
k1tmo0JbTDtFzAcJeZQTobc7mFWKI47TsWfHujvBgr2CTn5l8WUzvYejetUZKaA2
LlXt1yDkeLaYVE7RNVyIrxjSzQArU36+ujeztDXLwZluujaN2c7QCyxqPrVjCG1/
EuW3FGy34LMi31TKh0Q3emLdr9Nw3rmpyRUlnkIQFn90WaqACb7C+hDLoIfijCIU
BT6dt6vA38f5A87coC34hndk8PEMwxt6wn0t+6pQXJTeXzbbqZ4r/xMew52ROCk7
xoVT9BiqObJfvJnCATbEkcms9LrediP8meAxXpFmH34Fc4XqTQdrHbLYApSQNFuK
SFarF42YOrTuW1VJ/aDS0flb6yFM++C4xhz7YYcal65xT1asZfePUZx2frXHh5ZN
TtfVqg61qLwLe2P4Y4kMP/LYEsuRdIgwT/vp0Q9JZK5YMBG17aFS2YBd4BzC8ZBb
oRjkg3/tOsrDEztUO3CoKtVVimKyGLtYF9xZnD2z81LwsepHMseajbd2vOgkO3x0
C1m1b3jKhL5PgsEXkvtPDhhTaTD1jbr8Qrge9UBv+GVKq5AZKSuMJ23Eglsykmvv
x0WG9MOyPdXW4cpBmkjH+d3uP9V0Q+XzP7/jkov/+R/DAymoUqt+7/lwnpQ68tzQ
sv59rhT+iDKMStfrUciBUIiWjfDi+27yZLNCYNErt31dpLqHqhOjMOHf5j9IaIql
5XyuAC7VCY0v7Nk8CIzd8eSyCONoNCjo40sQGF8P9mPcvcIAGqTW9JKnDx7ZZ4HO
KktniK4YvtEAGPm0lk5rm38qyDCbfnU0xmDNP1kl6Ly5X7ZpQVlD8dYcw45h7pgT
6Tp4NUQWZHNsbm5TDYgftjc9RAqiLNJKqddBQshp8QJa6MEc1ZrTGmM7R9KJmuGc
7MCQdtplWEgRQowxxRU/ESfIOG96WM+4u8+yshtRknyhDfrN8pBp+VH3o19gqM9M
eGP3dCyX+4fjQETStD7vyjWSNXdAfrVkODexHxCpQiJcd2l5GG2sWS6xZT9uh6+L
hXi6r797O0SOJ8Lj4a8MIJNIBGeek0m82l3e7imDnpXEf+Up6o0EPQ2aHnEhfeuT
Zt9dZYgBuXmowyx0tknFCc2npULqZ/HVmgmWb6MvAzGj6/3LBY9B9bYCyA7hlpgH
Zx6jNbD7nAgkPDA1fVFUVjHVQ6mhCR2ZxXRLuIEdkLI8DiIq7+rkrqc1/dYsmL64
VVjBABAEelfGDvm6eU5Mu7pDw8Esuv/LJK95OOtCCxt3bZffsmualX3gF40tF0yP
myXdyt/2fkdta04t3BI5CD7yu4ZIOiUqo0wKHHTAkkiXUTDycaQp18fYwYf/Mb0W
tlp1U9tFlsV+8q8EYVWaAg1HdaKiornHkLr5D6cU4tC5RSNCuUnUadav2gYazuYE
hmaWF6amSoG/rOUsyn5m1OOU02+ikAEJRfouRmPCTyI8LRnKlctctozj125HxJtC
xPLCwtOs/I+CT6wfIkrvcE5ZH3QW9bmTu+nZmwIfMyJDmGiEvQiPnZKjBM1e+RJ4
HfvgG5QUihKHfbUlQRPS333k8pzbpGMbe5q7/ZWOCt8mxnHBsknhrcbQ9epMZklZ
0xBPYqDacjUGRtDzXFnXL5Is/XxKD5LvTK5eY2OOU4fm7wLTaZ6Lmd2GTz5px2On
0LyfNpp1qST4XYPo7CM7k57caqukmwJeSLV9A8mpnBcNXuz62gLwKV0zvF/GZiWR
QrLrX6AT+K035NLST4hFVnrDJuwUel8vmt/EY6IXNco1/bLNzlg1nIF5jyolIaJt
RHRJHcBc9o17kPkNeSAEVc8qC5ApqCYpz+iAt1zU9VirkDHLIyaWlXxQlEQK/HL8
czWPr53K/V6f7X9AFOucyNue+WU4+hdfO6XJOZmDWFled3CJyRXVIH26x99KztdK
GAGThgsHsUIpq5A2xIqqxEh3oW9QTnRwTVxVYeKAfhBgRa9KQCQbPZpJeDrzNRd4
J37xIcfwwxiI7IUNvDoF7/ms/v1MmGM2NFFuHzgjGgWE6W9WGj7dq0+i7yqXZDe9
H8zzHHOWfaNp9d5ptwEhJZT2/83or4lbTLQpXrzvvkQuQAtjlZeg4eO9062TYEs3
MQUiSb9khL4CA61i9iOKTvjLifVTqawK8V3ERiYwqXieSD2I/TjzchhrEWlFUvqT
JdrhRSdyb/wCbALf+iXqrsbBr7at4fcWqkiKHPMrID4FW+oNQO5kkYn7MsxQJsX9
yDlHtK7j+DV6yX2esupJun1wAXFhSG3UWRXd77TB+f3AI8+oR04NdMlLNxkNaVBa
qYNLxw1M4JJ6lvNoKVSzH0g9ZK1IIAJ+yzuqIFWJXZMdSFq6X0dtnhS0nRoOKTNj
u0ixLPk3mXAD/kHBGIeTWXf3Julj4nOz0kxpQnFZsmbVM5hmebvW3+gkHVpOsQ06
eSMxRjPzMZH86DZZT0UTK+4AV1XUpCGC94LhlG/vzSTVE9BCaw+QtXT39+sGx0d3
DbWXVjyo13lUt4s7AUvkRCEn/PZ8MffvjpGVWZZQz2Op3GvHNEL/ryf4VP/ml/Sd
QncWziQNJSYC99inwyrdOBLVjQxmBUtct5+3dYXdHp9zwYrHo+I+qKjVBhryyAqW
FF/Xt31sf6U9BDhXqpSRQPpZRuT60Z8f9s5nY5PnTO8UowAhQNZcYgZm37bF3PkC
nMFPplKgmlAJvseStEgEXISPI3WoJt9z1bu531hFYJosLShwesOcWAnzJWi9dQ2U
QT9ib8pK/I1GRAtW44BjhYK3x5xdqQEE3fb31e5q1JkSAMI0gTj3/Z+81Xe5D+d0
z8PkxpbD1S6mQ4GCfG/fdX4Ujbtig6wWKwUVVWe8H1TeU0pIyGwIfTK82zg7KFra
OUw0jSlsdR+/WK7Ng7FGZ9672tVI6OsAPvpm0BI4jybhWdl8UreKcZZDpwkBigg2
cskcJYjYKvX/zCXzpGWpHz81eCx7+x6JqPFyZY5d9FjnU1tD6gZWWx46jT2KR2p4
JL5Q33coJUY1iP0F3bIrbTxq5HA6vljSARlcBlanLe2yfaMKe7FhcHxZB//X87od
LWlfo1CnFoMvm2/BXb7S3zzY3F3i2ALLeRWWLK+9+FUnRfVVzb2HuhE9MhDMk9kJ
CxsecEe1jTer+UMM6+RulfYCtqx16FAusGtANNN3U7EWH8jRtwMaBqjYWjl90l8G
I1AUObAFg58x9xmlU1kFfqlyfmJeagYqrm5UPhH9ty4ARwtvjlOZYT8QDnsc2L8J
H410fOx7tK+JjwcXWyWAbh6lcMi/Pt5v33st9w5Qoqavk7B4xcvPvt3sgNxp1lHm
JkBpIcIIOOwDsC8MbbBLBdPX06XGDls2OjC7/Ghoe4yzvZgyYyTGRQyKVIa741Ja
Sz82kQsy6JuI4Qs2y95tn6yrJcwFTgz8299BrBdCkIOF3bjXsDsh6F4Tn8bcNinj
N9x//ItmxL2xAWsAnpA4nlVm8cdqUOYHj+krwVtnaJcvStVbzbsWNku2zSrqeC/h
/eyj2Soynfj4VGlz3+PVNHruS1tAsgrxVzC/cNHifUDTYa8IB9LuavBVKSKH/RPW
xm5E5SJnu1Jo8SRzIdevUVhn3XjTdPSfrazW6Y98rw5cgj4pbU4FSKkhtO049rle
M7FqSGj53zoIF1jBVOl6nqfrGreJLKVc0zjrkqnAr+l7169So/PdC1u2h/mP71Pn
vroraFoXv2jj4zR8Kwqpq9RBe1GWOyVoKjU9QBBZWJ/eVf9JbFGOGLKX4fF7wkZD
LrGHu7/nhiA94QfP/ukYQTV1E2Dv0Tpg2bxGGaahwlo0SpvrnQVBb5eVISfQ3owN
ZeGpx+t8vINyJ1eOf0klfmfNr6xpoJMQ71jA0q1N4PFzRN6KOqWGiaiNP22MwY2x
FJpa9hECiPdfORxOOp1z9jLfiJq2rvk2YjcYZRrBWA8WsZTNihWpL/s8x+Z54Aa7
nG0vdleay1ws+W7t2hxCNhmcznBWshxYA8fPLViKjgV5wiaJsCj7EFCowL/8e67Z
ObGcEe0+7+Lq2QIF3Wb5Pf0DtkZueNLQ1ep6WJ3z9qo3kRhUn9fbuPcSYD/ErqJo
EqYGw39Y2o+UBrck+xK2ueoMbswoAAHm/afShB4juZ/fBiHBvqoh1JLcxMqB9/+s
hv4PxgVnLV2uqj51O4+dWcUNeX5OgzOXV9zgM2yCm89YUDMM/tMLL8MqFbfQnGE3
brKPoyawa0QhSq5GewmXOfhyiQ4TRQdpbHxUvYN8RML4ERRbVQlmVPr8H6jIiRJH
TmBCtEcyxcDw6F+FaH6iwoJNzTOTzkJp5dCup0Rlx5zdkA6lXID3AgvyMlbo7NgD
7Zyk1mKlGFt+VLfdTkwhg/7HAoulBe5uBEPkEcdH1DacMywk2w/CfeMnmpX0vtlC
Hr6NJ2PRVUP5tg5XknbnSsfH9hexrKllJZXSWRfZ++2vGa+yYj8CaZZ6WyoNvN2j
x/VKFHzViSHLE3rtMBNUtD9K0vHUWUVEOROUZtlZGzq/t4YnCwALNek/GoYcuLVE
4bbTGt6aJ8J68fKtJOz4ehQ5meayZA9d00/eYEDfeMJQyJ24WyJgBlSGxzax1yoL
RxnMKtg8HS5FucLAxZVAuW/MWfR8yHwbn0biNBX8aG7Lz+N24fk08+qwTnnN0RrR
I1v0u8N5LuDWWIx56qd5lDa+7g3SFIwnR2sBtavXLGOe1g4cNEyv9bdN9hqTjjs+
na1MbVmUYSudwboPQyJvXA/wT0dAKXnrpxzeAfNOS++O6y5T1E3KqyeviLEn5h6z
iC5tRNEWbfH7aD6MvDtDSorSGGM13z9gPF10tHCu1F3p1w72NkLTKQ0X+fo0CQGA
elhT5hJMK8nuqDMGyxHjWknu+Jc/sIH5xO2dm4C4xZYLxJGZTwk1DFKfW9TqQL0E
iCL3e2VQm8H1ni+ZXj8piHzPGqToQOcDzd8hj3qdEg6uYBniltGpZHddSuVn0qay
t0dmbS+RHuItN0921sH85a9XBU7gVF2Y+/fHTA0+mOTwTE3jWp1mSocAbmm7CCJF
GZlRU8E0vkXUsTvJzBwoZvkeyM9EaxM8OyTA8LWIUOvx/c/F/aBpZV1qbmSpp6D3
dY4GkmJLJmYYpTn73IzjE5Jd/+PyWz77hA4hAhTAbKA3LB2fkdmOD7/6++kRwkXw
HKDy9U9Z1VNZlGYF/MiPfC/v67V8TqFpd1vTtLYDOZsAf4AZ3WbP1enjNA4cC+xq
AM0+hX2lXTdQpfEH8EFERfqS/CyobxQv7nzKj48xhRMrbkkvTGB1lCyTEfIGq5X8
8XA6wSyFeL6Tlx8dgC/mx4BM2sjMq1EElYgGUv61tamGWweDH6poXF6Izo4/vjC1
YbU5Dj3nthNsCrJmI5sR0CZX3WvPToVTrhOi7VjA70+357+HyPIvzNQi1YzeOEkg
xqDyuW5NuQ7JPCGWOQ5BwRSy4rYJsKV6NZBR7uCX4hn1+HlDrc77Q7s5rp35jPBs
eO6g7SmMKZBR2Hyb7Wn8P/9LA9G/prmFrcwswVdUQ2DxmyIplZi1DPQvgyP5bsWc
QzurBnt9UdgYVvZt1/tyOIxdWZyxosQGgu2gyPPMJG0MA4Kso16T4WesYP9eim7M
mQPyn0CHj8Sp4nnC/GCARp13xlZ7nxGAI/Iw5ShFtoc11b3ps77Hglg/d7RqwHtq
TOalPsV/oTcVw5mXJRciPhVyEvD/ykiL0AiVYQ6jnjO8zInMPp623hriFFntqqZf
QvhNiqpvBbbiCKvPOKSJxpGgJ6Yh2ZiFmu/74zWzjShvqfvA6ymGZj1GuZDgFPxW
dj7lXakGRiHVVwed0BzQZCTesYUh2OlcNpCRmcuuPY10Wr/k8Qwn/dbaZuzSOADl
OZQ1gTr9z9Up50/0HbAETjvoPk+W6MCP+T52QJeVeeRPVz37sHVHiqza9MAcCU/s
vFjLNduUbM0mV6lKaa2GAeMd/uq1gJ2nK2QsCNLsgukYXT3EUvqJkGq2pCrDOa86
HhodgwP9/bZ6DWixKTiq9sNBy7ht8OOD3KftvFzI99GJYynNlLzcPatPgelmxZ34
2UlQEo8Rgcgj489HAwjirNPX4FiDL/mlz1j2BRr7FOM0FVK7tdWtYZqaG6yaM0Zw
zJZAkKbWWtSJNZQ7nMhpHiNKS/zk7VPiHl5KubxxnG86W2Bvoj3TPNbhVoDzpKEH
bYabLUWwJpOOW3EyA1gLEng2UhNCUsDoGnDaenJW7xr/Ob1eZxxh9E5ZFWUFiHwl
9r5rdcp5UkrLGLwx7spwQJB0u4vlzV5zvjmkXOcUAMLb7iIXeW4EVm9TmwyxDjw/
whKTfn+5JNRo+rbJOb9yNY41kQ1Y/Lte41naQkpNx5HXb8N1EfatZz4HBsnJ3jc4
mQ/4akbWzUWmKwirsAo6osxk1tjU6GQ0lJJ/EfWE2QpNb1XWZ6LHqJQEMWm3Xgkz
GoZ851jq1n/Bscy6RV+W0v8jHGTX1dz0/2lBDksmqz97pdVtCuefoZiWpUFU1s71
bGuRRiDcIM6HEfB4U1qEyFe1Plow41AlN14mg5HkXV+tdtC5EBJpHY3DX7G2XyJy
0oKT2d4v9Ec9RMGRkAC0XSf4S7imfqi4QgQG02QUhiUSnzS5ay3NHSuuk2/Bsas8
7CCgJ2DsP/Agzq5TFu6JDxQXPCGJVvWh97gw0ziDR5g89fwYIoxY8JkW8tfHlkzi
Bh6gZdJwgsiwJr4GDR/omfxM/n1XaBdFipq6hiula30IxpwqLH56uUmbYYFX8Uwk
OLo87dQ7lrZu/ID0COUp2YxTOcrpoFEVtKua5jPySlc9Ai5ghmRTSqlsWuPhvkWm
ivAcYYINFBire2ZkGenbBFSDAkPH2JPaoEE923zqVLeDsbFIlH2oFIwkNv7oHdZc
HPdHJe5FVfvlkrfN+t4rRyF3iuVeIRsKbwlW6u3XU6UTFEhQQrxh9ehz3/tJc52e
5QG4W1gBhuz3q2Z31J5ab4g4QS+PMrQAhbGvT6sdttMOy4U4VN+cUquux9OBlQ5S
OYcice4d8ANosHWS0zHib4siqrN4zcdzT0HyI1xSlDP75UIoaUccdKuf7fix54qs
Y7w8rotCfiYg6oGi4M/X786GyCpJYeS/UqerEaerRWaexWPSxmgcfkxrbnpbWc0r
CvJP7501X/99wgozPUHpuaQzomkY5cAX1478mnjmdPwsgtCHouWh2O8F1M4afb6t
p6FntOAmKdw8WuUtUH4WpA65vP/ORnsCOgZ1cJO4iwQh3H7gov84fFfQEqeaCuvQ
b7iHzOSUdo0z04/88FVU0Fx2YVkyQAeEh6eHiXIP0/r/EKW+54QjZ2G+o7ewLY1b
CO7aC9zhObFt1BXwNnu8n6RFYppGBGY9slJzVInifilVx0kVlJ47eVy9nsxbj0YP
gyMeZ11K0eLXAChh4BZ5mV0f5brsAEhlwrmeZ8Hl4th14oyV2lNJPVU/VdAB//NY
D8eGmkY5CbqA51rqD+CWLF2R02Qc7DQdqO3vB+zA2YGDwrXjeKo6xvVO9NGNTna7
4gMDW0D8kI27CLWDyefVdTA0VGWnZ+7b+glk7LA3u6lhSy7C6RWuOz3qjE/qJN3c
YjaQvgMIY99kASJGNZuTlhmst4yfUm01R+tmZ5cpr6iygwxD/OvNZa5r3JSt5lnc
3dgxLRzJC1x6J7WtXyv7mmit09IO80yxofQzYmyqT9uWDmFhCPbvOfLcM/iDM46G
kI2/0qJJattVAhoyPidYk4dIayaH6vCTLEisGjIPxyAyCYXOQNzrtNWMaSqD4R9c
gkJNfTxj8P3gIIk1s3FfCx0snasnd3VCXc03kDkGhwY/sm4Ekl61hM+ZScc+Sr8E
ZwfOJctpvErGKfDvmBWmsTZs852keojBv8D3m4zbtPtRZzvNqQ75o3CMzfCZwlgy
V5vVmadc5EnJOq8eDgtoJ+OHCrlB8pJ+z67lMqwyYcTMyZq97gM3aH0jfQJX5eoE
9/PAp27T+Q0ToqiiHpmBnWOZfkWEVK1AhKTQG+G/bFuzkjUQ2e6u+bNgGoi1BJwl
UstCqAKI/ohtk2vd3kS0AgrnUkF0h1jNJtQci38DRZIenf6VfB9++CEb9myw5JIK
Ly4MrJp1zxCgqfaMWXlHTsddpoQKGW63xqvMkAG1dMpJ5vIRbZ6SCRklXfWEpKrW
uBB+CqobJZZf0VBkZvZAEz2JB8gV+zzHIh7b4hDYg59mRCvT3HIQc0Zc/H9yAg29
ZC3QBIF1a1u+BtyqMsHOPHMQPPIyn2oT2RUsWxdKpSQrWIpHl3i3pqFdOT83k5Gi
p1yQf1pPFAVj8fTMMYs+584X0CibwnwRBHCPmjaz7D1Mx6r3e9SpwmbW0bO6k6rS
Py3J20QhoI6JTvZxdT42o5lJJNZqDsaj/tz2xnSXw7qvphB/hgJbZsBzWTHTd5Sr
huR95ATWULsK66z6V2WWGCZgco9HZ8zexN7s0LeyXzZ+NzCLsI4KK0uXGzSb9Q1Q
H5je0cuKEXBuUygV6KGP/uS4btpegpdRH1n77WuFzF38XfbQzvgNYGGkn4vcca8d
smva4yb9UvlBCD2HxYF3b+jIq/Gpqmvk2YZtaiDzFwkJlnX+a5XCZ1/mOxa8FnUe
msyN/8NBs0fYXPnhqqPpK8pin2mq3apnOWKYzGGBWsCOiiQxHT/IX3p0VYNQxJ2I
o0sxBkLL3qnvlri2ZsteNazzXaZfjnTjFxMAFygvEa5wrodshwPdCyUWruKf3xI1
eRn0hvQ9H6Xpc6lkRRmDlLVyLAugT6Okder47RITUMLFrqlZL+v1XMVQWGHtVkFN
cmyT82bNRueyynmi/12S4bnVhI40X9BQuA/+NIT2Ck5YnrwiMK3WMyC2m7D3Plnf
JxbkGwiwmUkVOdsvBYE2K3zqc23QsYlcF0X1PGvlvfVmTHh8oYAcb3FoZbBtp9m2
k6S9MLWdF6PyHaQ+fvt9Scqrir/tstWwd7sIveM6KLyQ3teLhHi+lY4reXn34jDK
ik5AdNVBuMHp67dIL4gZ2GBf9P9UF5P06A8giSDMMkM7OV2cBoB3HQVKvMYp7/PM
X87Cs2FwN3NbKYCgdCfxHbbxKx3ZxsZznmop2LTVPEl9r/NlzBbPyW9konva4bcS
c9anCZvk2MII7O036Yzk5yrThH/VU37naTCOADzwJrofIOp/gXnsOzjMaq7pkn65
WIliFQtazVAVaBL0kNfTnrY5FX0k0UvD/9EV2mYYPKs+rRrl83CgMD/8cGpF5spq
MnOMkQfCHw6CvCIop3Wi3w+scuH/nhLbTSS4nrB71it6nhFgbY26ezIcBragYjig
U2SQ3iPdNzDntu/GYahb6JjtWHXjiiUkmQu+wJcuHVgLoQPyZQqZ4C/FlrMTaWSh
T86oA8ap7CZEz3flVlIrVonCIdr69V8QHReBGnZ5znHcQ3fUgt/9M2fL/UDelqaS
gEM8OXRBBrLl3l9E+XwFPo0ETA6Kl4/Mz6ZWTawrUUn5NtlqoIqOW84MHzC4aIT+
PHTEc563ZU3kJmjAzV9o3w4zntV5tDbfI+9HGYHihuwQD7UuhCWhh3hF/YsR6Pza
MRfRp3qxuR8m7+DRYPklzt5Cw+sAp89PLYAy7bVJ6BEJFzOJ5gVI/3Tzpkv1c8P0
t3XAybLW9IZxEOHi0GbD/7UMkDNHe6rQvMC+IGmr+/cmhep19UDRisR4LeCKSqLz
lLfXK4EFQeHElLYP/x5nKBFeYj+UP3o4SOzGX+fEiHs6G/G2dN+uaMcuIib2ri82
/d+9wREgU5qLVdoo06HvRaZD3LwrlElA5Qlc2TGSpFrPzZVhkomktbyYpmWCaGKX
E6VGW4TtQQVFZwF1NAnZER7YW2nNMgXclPM+zNotxIBIeQlWnxPshKgUHNAWf60i
coVhBiPcvjEg4aL3vXxTM/kotJ+43jB6huvP9ECClx18BC0haU6CSonTf0FcO9bb
HvQUFpFTUO/kRXwbJK2Y7BNaUKn1KOixfZAYa/2Ncjeb7zNFGnEK1gkVb5/suKqE
BtsqFg3NotJopFMpcwtRzQRqw6gXTGsoPPf1tka5hDJHM8C6X/K3nwa092ULKKmV
bSGsRuknkCsDjOgONYuBQjxWRawhVnCDzaJ+nsaLxZXPMgopZOyrzgbssWxhK+eW
+GzP7OqTr+cqtSAHFWlEfFV8lUvGQazvkS83R0G/aKdOVtlmLOIHjgaZOLcj15lx
RSgKSsj14lds5Yml1wk+hzW5zBGZ5RbaysSbO4G/E1p0+SaI9rONKB2JDg9jR5gW
QXpCH27zC92EgrXMLoNDmY+V1r4PhFOtzEmWnq7TL8jCesSRbc1LSEIew2ZW7UEF
cTH35j596Enj2GusRxsScWe9xL6pW2A5WAQWuUKNUvJbnBMaZmNx2Y3TL4HdXdLb
K0W8JybFR60UGCi8woyxaudr3LwKeWdYxUBb35Cu5DWs5faikq1+7lwi/mUSUoY3
oey6csu5LQ3/cscWlXTvEOsRtf1kfhdfohM2YNKOFJFZMv9g7xv63GlJX8z/vIzm
iKBA3OZo7564CS/bNeYS/0A632ALRQDkW9qLc4bgCXAFPTVinbyDFuUVU7XQTxDX
JMsMMV8tMiUXnjcU7/oMNH77PLKqp+2eJ9x6LZ5Lu2MK7jhRIa/yf+Hl6yz9M0Ru
Hj3DnUt/iuJ3nj68XDnaPCrcV7aGWpB8XUnG7p7D6di2FhcPtV9Lcgl4MSao3z6U
XuLwkhaVLpAKzs2xVfesuJLK36aZgdrAPk1f592oSI22e49yx45XeZdM8UYe4agf
v87WAfNuY0rU/7E8XdFPdeMSj2T/phIE8Udr+8+ykMVj5iQujkjYTphp9l3CZn+8
9vsW/CQ7u3f61W0J8yLmp7e/u1yBjGgdEdge8Jw8A9fTMCkOywf6eZmhibXxHBWC
WO9U97Jt5D4H/zUmXLmsrMaUgSq46D8ENh8S10pAEgPowehU424gA8aCAebtlHb7
IRoNJr7gRFm9H0FkHaNKfu7yAuNkzSMKebI/IJ/duPCIRuq22MdAsDWp/7al02zY
fkqljKfdxUC+K750iq5aqkzfoJrtxFeUb859cM7MLEQmrHP/AuxT4oyA4Fuy2A+O
Dqg04dtGnnFW0vKGcHIcNQcsb+f3KsEIEldV1fEhsY2OaCGOqJWT0ovNZvaWXuoU
bCdD6aUTgKoPE93vBnufBzYYbcOK6u49X5E9j15ZOeL8GYhbm37d3jVaCkWLTnKf
lRfZ6MzjvF6H8Q+iTTlTIg7vNp7bLXLBdnR0/m6u82VZP2I1cJ6Sl2RihIWqbPjK
d1ocolM/rq3lvrDWjYQhTIHurbPApZ1X41OcSNbNDJHKS6LbzIm6s+QCNB0l2+2Y
i1MBUIHLYeQ52oHxlfv7Nk1tRoT1aeUg5ujh508a2i6+volGao/4StG2hIO8657O
0gilwtsALuwcXrIrIcND4S9L6IdsDSjIrdNYr+vyXPEz9Tesx/TaE+fYMiFypaRT
UeNZJmpjpVsqRkER71oFoTcaierjqCqxSKLLRBQS4if4nKN/3E3yS0WWrpx+6PWY
RIizoqQJuy4dQ192JCMM9ZSyHPY0SCXEhr9zbJ0bbLArFHGuHU0ewChUJtYfCd0F
mTgpBjXOGmtXqShAiwnP8jtEVRcAhwsX+PeSYmo50CdsYMpHx2kt2Nliv4hVN0xd
ZsJpBPduCJNnaNYXziWDMynGJZIzw/LqgYE4rM60yik3iqivQurSlBI1yyB/O161
2lkt8fedKEXKrJvUJ0A/80A6KeZALGdDP4Cgfwgjh60qZMTU4tXASfBm0vWLcMmu
DfwRo5MINOAbSBRKLNvJGXS4p097YJm4LFyhca4tzom6RS4tjmOhXbH5Qm9+8XLP
ejKNw5BWiMtXEZQhrSCr1RlNxR6JaMbdPymLV/UFjITUIScy/olvpDv51LaBH2Os
Kpk3HvehzKpbZCduQM5OhVP+/cCrGfahE+vQ/96ikw696tS4Cjuvd/8PTPAG5vHy
ZkqcXrGeozbYY0e8FLjvmjN2IF8vfyu4FQL9/Mf355/aqUMy9XuNYoZLXxm6I/4h
Dd5swcTSEoS1Jz6nMglTo3eqXq71NpWsATD+5nfCFfbBChNscneKAyE5wPws3tEL
9PD5mqkd5PIg+frzoNnSNoemh+GRHiYCDdjEcsqpVavxIk8+EzClBN/j43y1o1Tw
s4HsE79t2q4QSj1OkZq5GqjRq2CCnqrNIxDgvkiZz09QDGDgAYqXc7v29jRMjKjC
0N2Y7FjimDZICwPq6HGC67XJMS2Klux4Qjq8f3zm64HFgVC1R3tYyQBM1XOhUNr7
XhsUeIBRFWremU1HNHFrVBqvsl9jdhE/uE38symG2lNpko/cst0oOc6Cj8d9U64C
pIYXv+KVZnxxh1KlWssQ+GMb7tVLqcsSlgJVVQwCdSu7NrKslK3+57iMJsKXk3yp
CGaKy8fVRhLT4ff9w3lwMmSSPhz4ticLX3M/LRm8l6lgqSbgNYUIkzEdv5nVh7jT
O561pXCiF+j/REdXEBRKDee76ZUEdo4vHFUhDUVGO/Xc9dJkTeds4ZyZLi5DdmnJ
NPxjLQXCXynkcPeDolVvQLxUhFIq3KkgDhBlH27y/PDUs3+zsvYsliaTUPmQzxfp
TacG7Kvr1v2zs43V8KaKh1lrjDhUCzRCLvChLKvmCslOKqHYsX5Ogec1SA41X0p7
CPTJlR3ZvEKhmuxvs7BcsF1q2y2msNcRJodTgWGLnUrtffQSglVMOgQ7fDQphsQ8
9Z8dKRl9R5439hTN/VLB85ttlYgphsSVHr4LAiHwRNDGgDkh3YWRGQ8R1buR0c35
dI5b5cXQCIcg52Z9nEDd3yjbMg7pYJGqMqSzKBHZA+tj445x+GSv3snRrmn/cS8c
f9CaC/PsBpBmJ4Hw3AQBTPr+Lxe2Ol8f29+e9SyCEKG3FEI1iFPY4VOH41YQRZSs
3pG7yZEoYV7V9l1XzDo9U9Qyzp95xnFvqxw5mScOeYQr4tNifsLnNFJQuCj4HAiz
1FcGKVnGdjEL6utjyX6CRW5eCc/WSTu1CwWuFWVxubYgqwMzNVSQkEH/BGgZq13j
3xLMT5Bo9EqBbmRuLqXQJ+qxee5j+A8aJokwq35+2mlNqgQ5o1xHqbwAH+qqHF+o
RPEk1Oj3ZhRqwzU0BM2KqLKEPMAcEjcU+YJmd3ylgNJhG35+KXCrh+/pjbzuGHfw
/WmicTNIlUCZo5VRZhgz1KxdHV6kladBSibyCK5nu4RnJGIiesOpRKzReNAWJ4tK
2BPnPiK/O1AAahlVGIjnoP8UtaMY8cjgE3WPqglYcjI1BqREm34CvzzAfwRKvbwD
gYmWJ39OkfpFFkvP/cyW++T5rfc1VJwM7T46qAWsoMuhBorMLH4QNFDv8Iy3hELN
8PbhoPs41w9heb7nCMo3bG8PggiDxrJ1/XxwnrqPIqtZ5x6ONsIQ9ykeE8xh+xyE
Jc/lDWl6VBZ6jRsnqTPflfUs6JGhyA/fYfgeglGPrMaLx+tSD2tn6VItsd50yw5n
ugdee+QR1VlIlhrQJOwXjprnHUSFdx01eyu0kAeOIWzt2J1mkjdTazJ1BWeGkgyd
/xz6ap0fkiXcmuPwWSp/8SxtxtMU7fq7xH4D5oZG5HywqcLV31uzJ2qw5IlzwQ1B
S60ZVwI2u67yvqdSBdYqksWo1rvx35iXHdtfiwWOEWjJfcnNoaYY018J/o6ABik2
RCblbNdqw9RlMxgSXyT+7Ra3irmzKqMnEWAeKxDq9IM/2O2HS8y8Giu/YJQg87gI
V+eV9lEzDl0K5C/DpSBIOxoYLnO8gAYQ5vw5eXscMQ0I8mMvj4q1xymPYuaLsRTs
X8Na4X7ZYQATQ8erxdC6FlDEQheDvRMUN9EnqA8kQtFlg91udxMdw+oMwRsSF6Lb
6nf/ypMs75OUsFaTRrcdq/s1UtHJKPOE4weicoF5wTNRLUOnn0nQxQqZT2FGQYCT
akdOV/kJ/1MAPAICPke8wM1uRCz6W0W62IutYv2+bje08vBQCp10Dl6Ef6oN6SEC
0kTlowafUbex95GkzMB/mB34sUsghQ4R5EF4lBF8vVtRmnz+DXNL6ySi5o+ILViT
2FiIU+Qwy5CqFkk4ZfmR7uxxTu19fS+L8Si9wAKQ92a0AGGj9XMlYW74cLVNblUi
EUgt+IQId4PwKiWAzZSrZi0WgQgUdMoYmvqGQ2RCRt4kLvuOcXL3I9yI+u8HdCw8
5JA1i4GlJlVtr09THLbiaMGKFybYUK1xBLNPYJ181881MGZcEqw6Znu4d6GyK7M3
9ICfaLN35Hc8X81prcM0OZp21NPnv8AgeStYopQqfakaS9BnQpStS5GO3IC0/+/2
+ObSzO26t1Mo7yvQR49vU12sqWun4k7n2swrsF4A97YC0cAkBvO8dbVRZC/sYPYE
brD5Ur9EjVof6ub0bZezw4HwxPkpYKUV/DZ0BmJTOZp3nX0oVWXeJNxMh0TAoO15
jS9su33i2rpvtH/IFm7D+wbPkg2XNW/keZ+KP0g/PyKQIrNKx3NRyIHbQMNDDAsD
sNElghzuLVjXm4O/gdMQg5eL36+zGjfbjJniJxtQMI+/Lc+okc8Av0yZ8rvC80Sf
6k1HhkQOmtPByJEKg3dpdxlPI6wePKHGIzzW7J17a3FtHvlZg0PB/3M0aTv9T0Cs
eUFNgssGztm9N9mQyZ6zswPEb4rgyCFZttSC4KPgktjLWcoz8QU0Wn/2SddvJoNB
EtuGM7VMTKDc2u4DTCbtJu0lvAsJYTASGRoIPoxrypREr/cnlBtwbL23aPRn3YZX
8k3vN/l4E69eknFb0wkfiN0+jB1dq3cU4ZCpEhaQNGMdWVvVE9djc6VKp+I/sK9K
Aatj+KVGyumiD1rcCwu0zG5wru19QWQgpyXAgFUsUlojP49VyQjRjKzWOMFpejVX
FNxbN6eAJErBGOuZP1dvaEhBHkF80wEtYZgz0DnQ4ShA7EAxShVdldKDuGy3Kl4R
XwzfAgTGGrIWClXYlg9drjSIALHYwQqaFWsTiZ7+YAnGcaxaUu/CjoVg7cL26KMY
kFxtd0QTNCK3O7By10Bw9fjWHaMTf4wN+z/xT29xMQjijUMwh61+qBgEnSSMCANr
UIu3l7FlDM5G37608uJd4kU+60Xb0wv7GlmsDrZSO3crNOoLMuITiQavIg4Z+Om3
omoY2spvpiTFt4s5GG3ebP8X1GtidAL323P/mnojb77Y885FI5bSF2p6HGr28Lt8
xqHrcXyoAX4NFb9S+Qp0iXlPjf4xyUlp6Exkmk4N+Ua/74yfCeTCJvMfdNK5GbVJ
CDFeT/aq7Hs3ktcjFrmWFP3HEcqtkHNj87QE83gK/y6WQ1sxiPUlsBVAy+plJVOc
IQ3JJd+ZwET6rFdn3UdOHx4jkQBTviLFEZEqOyzWQtAy2H0zSh8PsbwlnXlC/qt2
mwdtwIbfyrqUv//NqC/kelIJnLMI+znfsmuxL8XrL0KxTdPMLG+qVTdcnNygrhFV
sg0+1PDZiMwGmBQVT+E/48Jt3uapU9GEyEBOgW3Eo9HkGPkxho39snqj+zu6u3WX
zt4qz7e77LzEr41sDvbJ2qKjAcLg9d3sM7XnLieeLgF6GeIzcsVJiIH7KjpHzCZd
BvSzXb2NtGl5wdZ0PQPvdWrxt/UwVmE7wGmBeQD//cjVexCPZjSA1B8bwnmdedyU
dGue5SF4ix9RQOgvEITZGkh1xbv9EQDSNnLee7GhLZq+viUuLokhqLo0ub7N3RU/
mZ1FgNaHbOm1LIILYcr5iQCUyvFAAgN5ny/P+v8FbPyXJ//JSpDJfxNu+LhzLbQX
Nsb/0oyrVGXFowi4/pXOwK6ys3lXZU0p+KdOuv8ZYPw0aXMSzxzqkTTqA0vKUZx+
irCi8Mx3RzDC8JQr63fRSqS09g/QJdtjtPxJj5GKEVOxlu4VeQizxvzbh6eDM7go
V5iqO8iOwnxGZz82+ipGOFBStFdw8yCtP1XRVVdJAAh96IwW8HNip8tC+Xedf0JB
h1Sv7o0O3KL/qhAWRvgpJgXYpXRnG4f4z9sc3UDEvnmyHUtXT39iiQA/shXUp7yN
tyzYP+Z1Ao6qqTIp6WVFFRWhEUNSYleX0ckXuMxbvOHJRIDMaULZM1hUpYT0tSKq
Pe4rAWwZSSVwvcJxbJPn6KtO+JwUPsM6WCqnTmU6Y194phttAwYwzUmsdoWT8dtj
8F8Pm0SAliNfcwFR5ti4igF+3ud6Nhxv1SkrEi8L8Tr6QOQJyB3OiQEHZsRyu2Jq
dc6pqWR/z4DlGMPNHsYyIUrUxImnVZYFWRDz6BtJRWiFVxr0qRzk7Lwy63zRurMe
X6kY8DlfZQmeDYtpLmI3N3wxfNTDTF2+3qITDKuBhIm7MZStuRVXhFQCH8cwPfMV
yRxXgGWk9NonMlBETWxgVuLK2OmNm8uxf12L2qcS42wmAWaNvRMfsjl3SIV1vfiW
9YW2zKl8+ULMjqJ1jDiZ1PTshzHvO/aPTfyp2T52aowWD41HtMhz0NClCfIBACnt
4ZJGse0REi70RM+xp1J/Jr20RQ2VujQbSoOj02E1oc1cI7fuNl21nbEjtiKqi8Dv
KP6o5VaenTZm3qywb639Xl/hHmMSZXPo1neeQ96WLaYE9PY2tSmlGgMLGZzR0jXm
7gbKUCuhz6+faG00ZuLK83R/vm9E0O2e5va2qkUpOI6jP5rmdG/AAU7JJi0WysKR
FsxFo8AxhQ/38yPlGTSIHFacJcLmZL6MNFP5sCn6vmqhtEW602pLIYuS9TEeRTyJ
sDpNG6lqZswwpErnSQJfuOHSclxKgeIQYfhQ1C8Zrtzu0WEvdiR25VhxThpx01Z7
2n0gj2c1ld4ZPPCaUJfAtx5p51ug852z5EocznKExNsHJxZe/RVJcbJA06Y26eAQ
f8KKVCU8HSJ/22FcVVgSORS3BRXt3hyXVX/VD6h7bKdEUJzEgBb0rCERy5ffy39+
YRIV7ArTbOdxUdh529qE7MZF2haJ2ae/hrEZ2iNp6Ju16Nv1KgdABA07FmC7AHEX
II0z0B+sse1NQog8cliy2AT7fUvBbL43rXm8heL62eUdzC6/d3wLaSvxgfQmnG2M
svLMq08dFPine6FhvKf895tVvnwXVAAnyN9O4j8aNoHj18loA/BHGztSgJK2RoXC
ptsU3in8D4gZIooabsjlFsZEkfAJLCFXdGt3TdAp9xZ50axrTGz9hgSqyzqJHfyy
WV4s1zM3BVaKRdYoV9he1swZHr92mUZdOeWIzH9KM7/gPJq0M0KNpHyyETil13mg
Z9+m90jVyL1jAzaOfH37vuDImYT09b2QwM4jKIt/bUYAe8ZyQzsBaC4mbCobi1Vd
ZsDjV4VNsUYHR2pTGbDaQmJP1HNr/EEMfNyIzkIStUiu5RbssggkaIgW+eB3h7/j
h+lh+EfrqTY3R8Ve/5sy+sZsVJ5lJkKUhJFwRyPjY+hYI45gj5pphwZdu2EdJ8s6
58aJZ5hO95YD3mUP4Angy2T7BkCfX/qtFQ4uUlzsTQme2DwKKOPzZ7uPh2zWFqJ/
Yl2cFF1h8V7STSA5U46nIokKMVuVsXiFDk9HoueftaCnKr1OWqCO5LVmRPdivaqH
eiE5T5rAztZp5/7UwtXjDvfCu/eEI1Kiel5Tj9GwCskHm8Bx9MKfXPnwIdNgNJqP
tbMr4rltyEcTbAAX45TdBj/py1kghkeDuBHSAR61F/e6YNpm2vwWLfNS8FpYtoR8
NxSe8jdmeYmj3WYJvVbcoyNcIenjlAdxmIlEmGmKp1Y+KA3mIYcnmFhdelA+9Noq
6YEwMgw2NT/6cOE9HclTbCHGvmMTIMF5PDn1QGEoXWVxiRtuQl98R8ida1bzZ6WT
3CIQ4m/HsO6wXF5sOcXK18qFdeDQfT0PIPhEQhRPNR9ejAz68YTVhPM65GHd/Ykd
a0uDXgAbi56fnaxMRUC+okFfCt8r7oAZwFwGsbL3raxGuUYHOhJlgIxoB+hSwHCH
VRPP+q6678h5XJO/Q4v33SocZnOVMcXUtXpL+BIjJsHAAVZ/Y4GUJQULNx9beosl
G9EbJkOQwreHF9FlNJjScKLDSA5DU0Q9CepaSEJZiGHVLMq5rnkW5wMFMzXwNDqK
Fe1YBjiVGbekXKjBxXTwXWR16iIxg/OW86Vf6joPXi5Sxf3i9ZJDlr4YVFLezwdr
3ou3IP0d0a7SGPeEvz2Nakv/zwaMBIvbRrRnfm548G5mC1BMfs4EDtx9eFQXnKRe
n52vk7LszWl7173ZdfHye30D4rvemkellM94HD3QhU0UpDRuiiySGozlOa7tgNFD
6NZ8P+MSCmLeO6km+GRiprTcDnOEWOTaBgUQZAZy1w4+FYbDdKpQcWSmBnDgDzWi
QfZVz+Ovrx9MPUmCJbNIPlbIeUMFN6j/mnBzvz5HbzuzTdxzlDhBTBLl7fhmZ6Mb
3LIK8sBtc5tpXlQh/3AvV8/x1Q3HFKK2fMOWVFwQQr6k8bf4k7Q3+aOEI+rpTaNj
0r8jrtNy8Y43LdGS8SEhf71Oeb3MEhC7E/hOFCCXk94ZZNolZUBGgFa6ALLQkKHk
KAYGd6uYTE5ZWdCBOTp98xU/hmC/vglzpf8D8kTf4fcRd3q39q5Bf9S+kFExZ3Kp
7NHevFv8+OE+erB/N9oVEF5tDR48zgOCwxkgn4vzh3IHJHQAKCvaNtfrLBNpAYhw
n2J3xpCwIUUXXrsH5t4owBZt2jfm2YBrSBlUIG8MahS0tCGhUGWxrrCaY8+eey+X
gv22czyQ+0D6JTzUEdiLCIWnV2dULZmP18RvsW1TdNwcL+sFmWPMrYOjIRfP5CGF
12myz6QX65lf5S47KdtKgzWKLz5Py+YcY3j+JnR+1HoQLorvckVqxEiz97Xu6TV4
4MQgD784AMIOQoKd0yUTNY0PpTlkmcJfNRcXnOtKIEehdEcbrXvqDLkatMgMj7HC
7kim3MBvBLrcaZtFjW33jXJlq2UbAAqMRdnXiJ1L0bdC4enWqAxU0q5i4QXtuqvU
e2UsxgcZsUbFb/kTO9dRYm7oD3m2UG6op3gg5l3+Uj6gYLmShAbHj0i9XTAXi5jQ
TDAu7bcyhukkrZn7xpOsh10d5zUqg7i6JjpMZmsc2VvUs1VIgIrGsDXrT/xBBI3H
GYccbBfMsothkp5f/RTG0A7B8Rr63yngj2qtqSledjMrlOGoeJVlzqKQcUnRS1ZL
O7cZmGZk1+MwDtLiGhHT6vQSd9C3Bf6VI0Kd+hLKMKmC27O1K1UJ0SdKqYfHtbIH
zVag6JEiJVGH/JKMJGf/IM+1T0k8opooFnUlEP9JQcR0MMCym0497NrlJEkmYnre
2pN2B9/2dCTj0pltGK5OfeuugRULn7rvYUL8Sr+oFqDY88BRaGGLtXIJkzNjEP9b
6yb9362zF+8DPIhWJ3qKJQN0dOW5NrZrGjqnJZ0behrsJE7Thp+vYfjSdfsnWZvQ
FUTUMVTu8O46TdtBvR3qJ9wkv5bLyH4Yqlb0Dj2XSjnhMzLRXMfR751SYNQDqloG
9tSbMLpHPLAGS+mGzcNPPDFBeLzplCL9XSJ2uUPPtTPkTU2p/2uxN08tKqazcK/s
AkS6hlFuVNOYGCQeUlZbibpoeJMDN3YlbRVQc5swep8NoDC71vqGGdhc5yv3AHmY
SQ++46+k7xzzEZFOJgYRfx86ULScOcMEtPsGbEK0Ls8rserNeH23AEOwOfnJyGVC
5csbuBO7jB/RLm+aLelM3lPS+hbHERh2gAFfLxJC1LN7pFfMkJbtq7FwDG5fchRP
63fHHzEszTuIBMISn4qwRU467G71knvbLY436KGSqB6zGibf3iOnFhYn/QfzntFa
XByHuU6hgyjXNen+8ZrznjyTnl9zZ4oVjudk9G13yx4=
`protect END_PROTECTED
