`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XX0nG8kVz59DbpGvVPIlOqx4O7M9poGPPCSH1qgkMHWC3FbaoCjq2EKGlsiOIrpc
Rf/1MZa3+VP68nOTEGrWYlko+0NrIEovge5Hp6UBkn64j6G1dTJGfQP8AYVnHrus
64bLm6kb5avHgVrw1sM/E6+G/Svqs2BMWfwYU5c6X2kx52jgPY/3MTROpIE82EiI
6poExCSU/fTS0rXXLelBYHA9ORpMeknbXE/lldZzHGIS1fSpfbXaV+KwCHUaoxAl
3/q6zmzvUEj7oy8RRMI8ePYfrGakcROU6vZrFh6hh18ESRduyrD2sqsEorCTwu2H
KFww98iHra2HcwKWosfJumS5NQonMuG2IPK9EY6cXrg=
`protect END_PROTECTED
