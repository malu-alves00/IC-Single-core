`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hkoLZg5wQYUs8MPlmBJgaA8Yl92OaBA9CCBpy+a3w+enkinfu0eIa+lZIMGWsUf5
XfC7CZmp8BrPaVnguSjHDP/o8vw6m6QnvB93VjMA5Q8VEcUjvGP2WDMRQ5Qc/4x5
11FBi/JQldIXGIJCRZHaFvf8g24PEL5b897QAOjQkE25xvUIZuMXgO47gX4LLZmU
zVxfadEzOZfNgl9boouMUyiYzweQq8B5h2hM7okrkb4Oj+rVtoIYX0bwol8kDjx3
I4q401uEozQkkTmsOlQLtE+0kGqosg5Qv4KDBTgVlB92kJ9unIt3phBbLPLfbZSc
2Z3GSHr2nTwQF47wPkLh2+kQY46VakFx4ZV+PjoRMD3bOuPMQ/F6u4dFXkNpWiPb
XrZtqbOrruC3AO96TUxdlK5B7e2Y8Py5Qd+UZjA0JGRuXBJ9ar9wqs++OMXj1oiB
/7DgOoKbnO0H1w4WC7ZYCpDVzoSPvFGcbHQ4BA4VokoRLfly3D2MQqEzMpuMQ6Up
xFyfBDI8NgEPH4TuJeSUAQA2S+DJweSH88kLbwkfWIFl10KpYPBx1Ky8AcTMrE80
/f23ZWcrM43X4FuXuRcGcIHQU3YqaVa8cWK93+v3lF7wDLj1r7MM97XmNd2Ds+7d
OryNd3orMQDWa2r6op8HuFVX5lWbd39Q4USisgrCVLmvEaerUdDhsyAXlHffBn2O
yK52UFUiFbpQLRzOAtO5Uo0gctYGCaK/VVfqVeR/A3AHPyGmkb8bHgyhq36twwu0
nkctO3S25ncvfrtjZocgtr79U0XqhaatXfISkKIzixJB81/TC2POFPZ2jq2Dmkdg
/k/r4ufF2NkZ3KJGQnEG+w==
`protect END_PROTECTED
