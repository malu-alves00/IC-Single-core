`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+YgjiJZEv5xkUs/y4eZrHLcePahkyNB2Pl4wuUW46IBmtMWjH9uM3PHCgbis1h1F
SY9DZfct31xekVBiQqALSs4EnOaVsnkUxM1GUw5iH9UoFFPs1uK3x88IIE/bI7jU
ETShF11GA5pJMVU+ml11GmHuJaU7QS8E6XnrIs4e4VoAupBYSy3Lzg/NNDdFCvke
AErwfhcsOUtM7S1QT5ZPnSmjEYfaBnAK3C0tes6VpKMcI2pq/Ty3RF5aCgbfRc6+
t8a2NtAY2k4axWv7cG4Yvfl5QiCGrFkEdzkFnn3JyGToa2Zg0uIvLNAnhadILrIp
ssFkOArxQP9eCOF4n9KN4Pd4AbWf5Z+LM6AZYCWYDZByEepHapvuSPANJ+mFFM34
cMK/Mv3wkg9TUgYtipmSNR0zhaqQqB1NJQFQ3TAI3kzOw30zyl9cTbEzYABk9GOb
kwyp2OIf0aaIo+9ggRS1ypyhupp09ku1YqBc69IsowjI3VqqRBGg37NEUEMeIFHl
KunJlLKNDkxZgg3IjNsO09eiqc49ZB8ly8TcTaAK1PTkzbWNTp8pVCsF9eflaR0x
Ob8lYotKGYuIULgfk+TPnS6Lb0g56ni3l4oWKl0b3N+XjMCj0IT7b9+/XjFyl5EX
VNs/k1OOYfIbznyWkTPGi7x2n62mWG+kSGzqtE/632SevLX0LJumqVn82X3Yw8G3
08C+7f2Mf5LWWcEnO5A5Gh9jwVM88Y0E7+eox6+ZTMwmWlYC7ZSAv8rJur9N316L
t3g1z9FfSiiUUF0rZd1HEP/UxwhiXOQaVCzGcARLfvmnX1OEsmbf2h7wwWvDlHbi
wwIAE804TcYHn3l6mfvhgMOAu6omIeX88rT8rxDQsTqcMr39azz8j7PgCM6WCb74
qh6H7ftUu8VpikMhnoHQJwFf5hDtORZupb2L0ZA2cNeO9EDPqu1RtGUHmUB7WFaj
1Gu8FCrN3h8pE1uFCeSi4AGUtXP2exiWpi8Y40DmEKif/LGarYpM8aBusf/oVsVp
kxEzNbdDhKKGc7HatP73ztadD+EECFmjoOBRAatm+fNAgDVK8p1hy24pcdpZvFZj
l1HSAX1lEi1kNYQIvTvFEMSbUG7U7v0QF2TQ8ni3WRv1vlLTiQ2G+uqGVaD193o1
6jMrk2P2DNwh+JOpGUEeXlaJM9TJUTlgzGcZrKgLbFYOLN8t00sZ7VhonpkX+FTh
CRKhR5FvvJrM43Yih1aULXK901tOvXOfmYLI8K1F5BXje4vg5mfIdlWk9nfjtslL
gEy9MXi++owkY80tHMQ4u9M8+XoXfRBl0FIlUhrqzEEwJJxPwgy3UXcyT6gEm8JJ
mxBILzzPngztab7Tk7hrnAl6RJqqLIYGz/kc8CPWcoc3aM3j/864g9NKtSBEi3o9
PrfKdiJaUXUYOqeIZRXMUTT59ZqboVAUFaL9LeVJwNI7yffsDWub0haiYSHwS5Ix
KkGhgmhFqEVY0ys0BK3aLLUjyF6Rwt+/uDPGLvJDeh94cxHn6hb46WVwVm844nJU
lFmcAYqD5C60QyyXzD4HO206cIkm+wj1HhIs0h3yN72iWtBoxiUCxc3X3x7kzG6w
h6ZCSnvbZ4e/aZIOGJ489YLdZfPBTPLe44lDN3DSTOqXEMq+ITsSDZdyn9ySNd57
eIQUYm5676XbTR2T9LMqHhg1+c7HlTOcFjVSIEdbqMeFbm1qETq70HIVVhY6UbMV
Lm350TCGUOwaoGmcFr2swJJa1FIwaWjUMmunM98HJprs6bj/MTK95n7ukTyYYteN
FH/HTMeT+pGecS3rBZEzEGurBR7Ode53Ld/T4ASdHxwGHu72ZnuO69Jftigv+f1Y
pyBUf2wD+fd4vZqp34k15zZhlO8slye19cstfcszufopVBRJVrHpzai7yc8zaZos
QVN9anJFlRUJAP4o2j2zk3qHVH9z5m9aAw9wIvCfZ42ecLajlJqZ+fs7jpRffOwI
w2FpWvb+vF0ScbAqPoMQwpzeIsGrscKCMnN9A1fBJ1Y77DAzCA0Ord6gnGl2/Fjd
C0Qa1xBFkSR6P2LqKgH5eI+c/QWnbMc+T42V9LtnQaZjN9XoSipAOiaCTU+wPcm6
VT0zap1vPuSb38Uakd+GQ6gTzNrRnxNV8euiBpR7vrRxQWO3RKIv1FIxObBE/m3T
WLtg023HlYxrkSZpQQHMd+W2sMyPtF1vEjO1EqcPHQzXR7mO4Gi2XtlnLMdO3VXV
vjYgQw6LHg7mX7yoQ9woyZAzJ1NBicGv51wp9QjKevBOKGAPKQJtz/hgVa0RKR9e
BhmlfCvvtPWY4gfE5y9u+yfmKxpX0FkeboV39zxwX12X2bEL11x/e8CqADlU61G7
uMsqO8kAbFNT9zYuYVj/wGyz/NKftq3PCaIRLVO7vs/mtkT3mEuOuH0lxLRFJOwZ
UZRvvtAUsgOmn2IkzZk37BIS6DceZbISOc3wax6UJFmZijzmJibWkgHbrGZjanGH
mOLXXx+mBsVcPp81+XhqBD5uAmxa72tQEiki/1/W7bpHFt6mTKVrtohRYOfbZaa+
SNv7fK2t+LQOe1TBI3aSQ1lT3cwvo+SeyVE4IsxdGlS6t5I1WCaSQOhDMYb+EYKc
vnYWW4Q5qSYvdImOmQ9ePKN28TzxNhNuhg+uImmTCH4zjKcM0EfzOlNLllBoddUV
UtdtVjWl7OGO/hKxFL8Ws17vIkQClqHe4FW6A6R21NwADiBGYYeF4+E7HTbo+trm
mi4GKtQ3eg9aa/nmGYvNR1s+sN824Ul9t3TTXxmwXXmUF/aDMn+LsPXimcdB/146
GVspDRcj6/cAC/WenNgFs/t04gF2O9zZvXB/Fw1V2R4UFMdAguODsPO/q1AnIGz9
uXkTa73855y4NTwKByIXm9Ey0hiQZnvQm6ZHN//NFgMlGHNngf3qmI1EC82Yv8/9
oj/9QtXgkp4g7KkuG0RwSrnHV3U88/YMc5GA63ujoOg/TicNcQcQLLh/eUctIwOn
EL5D7Z16JoCvf6uLMDGECFG3cjjdNpRXc6DGu7TJ8yUPFVglgld9Gx3O9TMDwi2J
xOFgbRsV+hY+Y++NOsEAnwPGUc6BR1S5nez5vEQCIIQLtgay8NQDC3GRh5bEreQx
M3idaTBZriI76F040y1jtjxy5yIsThxoHDLsWAepsxtbUE55sVOdgaQZJAFlUdkL
YJpgnGrgt00cEGb/tvPZD9Qbhc3M7IHCYMiKh9ikjCU/r6rVKAF7p9IfjSnQXC2f
cynU4IrbbzLh6VQuBfYlyqfZth86YPQYbXWQQEKKHm8zxHEYGfsI7vlPFup/6iLj
TfTGw50xoSTBKVc2EGz+hLOCYEADDhyF/DVOBcbvu8HHfxBli5i+kqpicS0iukJf
I5kqFLIL2QHNpFj/LF5tYYvVWM1NekO504MANd9Y2XQtY0fkD9OfCKFThehH/fgO
vgeaIinjWixRTKlJ3zqa7Ax4GfTTBuV1TkMhdqr8NjGfmGqUGtgnICijz1CiKRoI
Kbb95P0074k5zYEDYJSFQ4IgeT/VPzir8tlu7t+u3x/Tf90aHcpknkcG07xxYRCV
qIJORtFCd03UADtZzKGkJy/ooEqovH8RCOomxZCkJLCyXWGOK5PoeSiGlkRRaw02
DO093RNxRh+skx+K/McP+oGdGXWfQRo3ZJXeifWi//tQ1o3Fg46BzRx+xpNGML7x
7E3G/ouSjwwQX4NQLP9Zbec1Iua8IJaYpmf02w20pii4NKUP3Lh+jAFeAnA4eZje
vCoX7wRN6OUSz2Ht8XehfFplQNvBMYFDH3uqweWKbiV9NIdaNvp7RIhyh8UY50me
QT+z63NSWv5U5BYDSXStVRdBoYkfTkSRhRLkvy94ZDfkZ5UE0pliUOSYu5CnVvIX
9IFVTXPUYc8AbwD1xevGJcKkuyA5GpBc6ATS8aeEaH06e+K+q3EJ8ZiTMKoqBKqh
KaR7zYONDsf6An21gQJwK1gkdLqI+CCm60Vw9CqiNnH+fVs4AaIuPVXQTSFWt0Ow
dluEQr5IXkKdXRB5g3Tg3g/95qfb1VMvU5/ceAyJKZuq5S5+cVswyFeihhrlfSKn
juqdl7eRE4DGzFTDgFNi5jeL48qnE4PDv51U5A1+7o+DCho7vcEO/d0DT58u6EVo
68yZnjXF519GoR5hW3L/yIrgLRBhVH2b+IgenShGSQcKCPmaiXkAAteJN9zKJhhz
fotBXKCtAR+2U7yLD8xlptFfLhHHKPKOwAM/S/OA5XIfUFT8rcOs/grjcD7OSz4u
NZEV/trU/k8U8nYtBkRX0rvArmgLKuhrkZvZUll9TxEru2N8GpJt8PaRDB8vA46w
YqIyPv0c8RreU/m9ANGMZObua6p2IMpxfvBh1xq/tv8PZSbFTmPAMXNiFKzWcaha
d8sSwkDUGfbJyj8HNPe2xfiCSMUUDhOjHBKPL+R/fa+TcH/uXaKsiX/hrNnuhQ42
y1TZrfgBOoWH1atv/zFcwWbSMsbLtuMChEC7PsDH183aqT67KqvkjapLvKwG1Wi0
DL2okcBIr0Ga+stW5fgB1Nhu5DA/3CxRlCGAXGurphyr6CgaPQwdYjZHnwFpc4KG
Sq8oJkKCf+1xzl5XHeNJ2H/P1OKKWt3ODeYrkFwKL7F8FVEiUwj9us7Aad72eCp2
PQzqi10Ij8eRyDpq/KHv/u8zhJPZ0s6Gh4sXOvgJe2Je+pbLGRbtIa2c1mCEUXIT
0AIP8+xWBmvOPeRcF8eQqN0H/vhtjMEHaNBf9K1i5XcAtocxFEkwJq6mJqPmkkEZ
tSq7UOQgfVRViqTCvr5/rl7le4i3XhbgZCUfqPNNVGCWH6e58RgwRz/Gd24wdBLk
dl476KrTbyn+TE00kzxWJlDeuNViRoGRp2fVnzfbX6U/vQ0CMXznUhcGLXWjDAg+
iGXYUkQDnmO1MoJPhRTTmm2g/BSxnz/rU270tKZk14IH1/WWEU/sDpan9vTQ6VqL
pG/dZmLgNA8B/0vMT0LVcQzRJLL2Hs7DwQ9A3L9qP/4nKVAGVIlrfhJLP8hQG4p3
woVwTmID9QHA2TxldKT0Cq4Oj8FK+lsrjDtiE4coemLS0E+EztvuCU9QGgZKTqAV
53kWH7vFEHILz8NRsQr3RD3J43+JMDD7yx1ESltn3v0dJw29wsE4Ooj0ySplA/1A
4nk/NhF2QOFFRwirmzuZAE0+yDX/iqBhMNfaPDI68uDRypyo4JO/S+IKqTzsjTFH
rZoMkecS0Mc41QcmPZ4w1b4BVhgcDb6ybeOr1/jQ7UADKHX/4nJkP1ftncMd4iIP
ftwOD0VJtuyVbBsstfTzhxXL2eivE394Zu+bSzCRSWrQ/CAHViPEjZbxq7QMVBxq
36bu6WndxAE7VMymL41PpdwO6LOmyePktFcYW+XN6XVysr4lCiy2t79KvS8DQv48
bPf5c67B9zCLl3Rku82QOf4Bb9PcaE+migMUiD7sE3GtvELcGZuQoBuYxjGA7PdB
3jnJ/QLkBofrLZ53WG8WUKJOm2wjYNGSxeBlHp3k8AWs0Z/nPSoC/dPs2Kv/bYSL
sduDapOJ0K4FmfFsY7sKsi80JnUBEOh30KzUP+6QbxOql34PGpeiCQ5gED0lOjw/
xqwd/R76lr2jmnp/2sl3yyIesVNKI1DN35bkk2NZJRb5vfQLEKWEp38neitLKEZ/
1TRSxg2+a7zNTeOdBztzpZqY6DHULeucz4Q7P0KklsiwB9YP39gMyBfmcJEwr5XJ
pRjMf0UojAb/c8HgtB6TlFUF9y6rFZKA1yQsFuf94y1A+zPrTxfLeQMTDvKi4/L0
iObpITHLZF7GhCX1GzSuOQWRSBXviiNAyUyIqO1lZg58LzwbnT4wTyTfSsziDF38
aN20vbq63HPac018CUgS6LioGYRn678qNElT8QYkJ7FT1dDdEyGKdlLC3BYtFVcL
gTUfYsJaEMTF3pcHhULduzPQHv6lquXmtEu99NtuNgH/v0gOc11usbxAtdXj/5DY
9QUsfkbS2JXTYDToKG9AsJa93wWUQwqVUlraCa7Wp7izmvHStMMDZyU3C6zUg8aO
Vy264yvohG+EY1QUUvcNtvq7R6VgLvR+5KftW6+LRsydi2Lczz8oaf3gfhFKYfsQ
yn96ANQpkDv/+XQJ7QzwoZy+LUSTZMvMRB7rNJ9KsXfGGdB7W41NfDvQC8VcqWm4
aG1K2+NtpPjlN+pjfvB23kcy4RPzzOBic8Gfchk49wN7G59Qm7vMEhHpzvN/EF0e
j6emQn0czQsAILyQxNo2cr0Ssmj2SMbyBq5AEH6R7FvSXk5sHvzyA/gcsxhBBcoc
Uu1zmDWCi3+9nLQHvVUIxmvvdskLqzGIbwQOPJszjym3d/7CVfWpfm73Qh59t4uy
jWG8QNKkmgeISTs24LC5gw6O5G3YQtCm8FgrPheYcmlyQ6vcOW5CXVQYuyNfqGVr
Yek9mKXfrEA+y6CGzVqGqOgEgm+koiXflClsF/1cceWEhZqLvxwmkBWpcL3u9Pvz
msaE7Z2lKelMVt+LV+FPGHnjxvhBw+tA2R01mwTWstaZCXBuzHM1QAdx6/UCNqkI
k+Zc7n3T0d96qCyzgb0k4cDrVsEXUjgo/OqlnXuTiyylEuwzYskPZJ4lEULC2vcH
bYptQnBz2B2cmyrvvdML6A+evMI4w4wx1aBARX6vl1gYASlvcVnKyiriAT82ozw1
WJO/V3P9ccE2UK8/JCRyQKwadhRd0QivIh4n0AG4iILey4oyEHNIeGrzieFGyOKf
4YcJuCQ24KIcgdn0j+2pS8uPIoYD3zkRWzK1nKKm+IRMy6AdkMtBpPf6kO+A4T5J
hlNIqIFf8Q5h2Sp/KcPsaIEQCmDR5L4shcXFmtvuz2g1nJKFuOjPLW5wqV85HbA3
LoJpKCVBN205fVqjf5jsrhj97ROPv3lx79LDBu4Rh+mVZepiv9kPnSgsVcAIjGNT
nXuBwawdJJDMN+veXeavLWJAnugLwU2YYR8mF8Q0aaC6hwtSNXHUzhZ1vJCzAiW+
faehYRUjbd573cP3ZPc+num34mMb9PTEW4Z9xEYBgGzvxgcloiDXxoUGSfPynghx
hRf17n3bKE8S0VTSOaD7gjbmo8jDW5eI0bNqesMsujC5bwL0lU5Bcsua0z+wDuII
R4Y+DLQ7TXer7qbDup2MKcvKTrT3B3NyslMcp2VkI1DfgfHmjUnvgkJ3SLbezzIs
l6dnT4KTrTKti5SbXduH4yCwKPb/zyilGzDDPBpAUhyWmFw2BywConw/C17I/pMD
gayOoOfQse/rVFGC4tTU8VIBztxbdtU/5m5beaWnWdwKrGE/V0biaFTGLmzgoD0z
SS5yRaeEskcMhTlhvsveu5gHJOMheJKpAnfZstC3CjJVQQXoZmGdz+ya7OmoLpRn
rJXXqS6vDeZVUpoWmptb5/bqEQZFEuTU/e6OtIzte6TmJnsMP1BLjSWxZGv8RXIH
aQ9zsibqtgLGpp0XJDMHmuaCPwcQ/Q1TVQLSTNVevRye8D2DbkK1bAXYewJmTlis
CLV1SwMa92SZCHm+nggO+kPAcs/oEpP+Vnf04rR+i0P4/w/rhAAVu+PASPWClWGa
mpDphwFaqbocMLT9bzDs/HGXWsMzXCxFtpIU2OQpHgYCn1A5dxflNtME09ZtO0yX
R2MsH+wRwOQDOH7QAc/+tn6fNBqP7QfTDqVz0gN2+3hYOrWFr4lA6K4Cp79teZtU
YPD4Qdhc+plA9BWiMwRnO4Ax24wdoz23NutjEhNNQaiQhi5ksZQvqD2wqemmlp8u
P4M6aCLaFtbmW6kGIkapS/Xr7knD3JhJ1QtAxirgJpXLcFfX6Cy/1sORJaFvlRQi
5KDukvYeCgW2mdoqQtIGihwipXeEhh5OP0pe1ZgY3/84byXCcSdHK3qQTDlLGnF3
nAaEZn8+18yvHuJvxzx8D+5NWDv1sfQJ794MvmRLuDOujzEkd7LDrouZEeDBxrDC
9AGLQ1DUmZKRprGsLpMpNOCNyLxspBkVF13jKTTrt3D9xAHOhKUxbzEHSdlNzz3W
2jsLIdI6zY4dZslH7J6C7muQez3RerA6A7ZSL0v6FGDXHBVGbhN3Q+yd/88OFnFL
8vJp7InhF4IszoH9+kqH1irknK+gnkYbcXo2p+8IoqBR/9WNI09i3nwh3qteD4fW
40sDSmUReRL81RkqlTmWtg4XHH9sqLZVB8R+yv6kq34Lr4IrLUKVEjqPe7v2O1id
ZtT/gwtVfxPWtbGM+d6/79nkzuw5t4cI13V7Yg26n/73gD52tVieUK584SXgIhOh
0jBJXshoJgzy+82QTO5s0pXHtIkbqG0gRbi3079KRjVXRW/FZKQKiiSoPfrjmxZ9
QI/GyztXfi6/LHoKbXMkTCoWz+kIlNGqJ5fgUhF819cebm4Bh/EzS2EEqcfrzOA5
eWXjash+IU2iRE1025PQVwjfXRftMsyjLn6C2HDUI41fyqFCNJxSE/GqQZC56xzA
WuoN9fORcLxK9ga78K1/6q3c/bhWxZwnQQVRNITWNefv8ehnWF6Z9u6x7kIUk34L
25PDN3JAR9wn+S4NGXKaRL3qjBDCPfO9MCFSxFnjBoPvISqZX4TW88P1XM9+DxqN
1bZuDWQzOFtkVi28S+w3L9ziwKFSjQy6PpFphicW89X5pPu0GjzQxIwg+2cRnKCp
6jgA4goUjmQWyajFdIUlHlmY+cuqdhVHmTUsPcQyiUDGjPPgCL6TiFYzEF3/uwbj
WHgGRkUY2TjYZJqR4W/6OH0MNSUdQ2R03z937nrnCwsXGc6NuOt8yxtdHzk+jm5X
dFI+aZc6wJUIDgyC4rhcPsrPwl7EngoEGkJMx7tSZk55Oyux2DGnZZtVhQnB/mxD
Ua/feBOyZP76r8o7YyU9jRh3QOzfH4QfiVSPvUZ3BsG3k00VhK9XB4I/3+Io7VYJ
wKK1emR4kHbWOY33Z1sroAUE9swBnQkCpYXw42iEmxdTuYDPTokV6rdNddUTMQlw
z7wO0MhmQFQtGswM9YFFZO8jC3soLI3GRdyhzbFYOCF+eZ44blKWQwNueQcKAL9I
Pb39XCRyf67sciX+biEDapwD+CjxQq9x40wmZ3ReFU2zxoKkda2IUB22rTrozPgb
4Ya0z0Kiyls3ClBC0BFNYBK60zaJVN460zSZzaMDotYzFgEQA8u11Sw7QPBVH73t
l24Hw9asBF3X+lIH51fgmbX7EnUxPAyX9KkoY1nvlbTmOZrQDzfWplAxcdbaBqIx
HFDJ8Z5Rk6bTLeIMTUXmVymoxvlo4qxf6ykazuRNiPnbpF57EpAaJoJK3rKtMstP
DmCNxKpLafzujB1OFQT38lFsYv4o7CHTL3UcuzeTpRpQWro8+HOl+oElS+OTWXUZ
mkHmU/pwYUSxqwivb4vSNvsDTAfg4nFVowkZ2KMoEuhOPn2Gs1BE6d0W65fAupyD
d6oR8IEQYU2qmcexyfXS+vg+Fg1c4ccLeIDAeCkyi+Gkg7xogOGsbfNLJ8mDoVtU
xZhcPiPW/9MLLn/udjqcJnCs/zECZF1Ihc2Ef0sEn7H3unuhWFMy24j3bQcGN4so
nxmOl2X5Jb0tnm9jviVXvMKku0CrDtSXLWgrSZfDiUrdQG0xVreeH+2ym7uzdyMB
B9LIT0mf5I8qGdePvYjwuVPg2nVQ9aRg7sNcF4y384VDpUT9YVwtBAp26cUA+CHc
IRBw/+smqEH+C/BYt3tplecwjB9NrlI3OEZvmt83nO2ssBdqCM8df1L8n1uSGg8F
rvmdFAK1swQFnkgOSAhto1meUnD1hFbCogoBeBivzM1goTCMuTDaAqA5B6+KiWpd
XrSyAepAzLYrEPKBWvBIWnd9hEr6xnznnnedwEnewXarBk/KKeE0fYsC2FttnxSP
CZNRMnJEbw+Gnjv4gPnrsTfewdRZ6u6i/JLNicMmWDpVBRLNh+cblKZJOEtbyV+r
tP1atwjsuIqTV+Wd9pmwlzCdYoZUuDpCtQBG2NK1q3myh+xur77eKKnHrIj9jtzA
NrAqF6SfvMiqp6F4XXbl/cHkcjG9SxefrDY4Lz7KZGBvdQVwPA0LS/VgOPxuxqzU
JSDTVjMayOCOcO0nYEgBjQ0/SoJMfLzMhWmftjrvptsvg4/DtavuvTO5EUxh4jDd
VlQpl8WHrIT+YWtqSZYdaUec34HipzQnoAgfe/6Uc2dqvPuhSJiEdhr63QSZeGte
lY3cmw6diBpZw8ZtvkJ+4WANNrsMmtNSi5ivMoiN5YQYdikyCJZQN57r6CXvIlye
hLc7k/criaTifqNFrnVqzmdXSzzm7ZGRnZCgp/lKYMLazyeXedLTrYZR/WUVpMUk
B3m0jri9xFYgMrT0OCf0iEQx6jfQWhiXtFTWIACiXAP8eCw/Xr+KlZKhbXRG7NER
St/ATQWu3esfmV3VBtsTtSpyynQqcfDOM8AmgFBgKJ2+Eb1DnZZr2cGAw/PWRKFr
UVbyuHJ7bbYfdwiyl4884TILNju6d/BA1G3twXuq8g40L+RuaJ58dluELKCuZx2/
fnM3DNF9ahO7GGL0EPoLQVJnEXvcSmkybAl0LyuZFq8sTM3niBt9eIpq/SWvsxxs
edEWKQOA7sutU+FKUoGqmK58IzZxj9pr607+A9vNybdPelVh5E+O2KnOsPZFwv+V
rQ4wiHZGcUWfzpvaz11ylMBmZAjJ9n2km6CAKP1R5uupp9P1jVW3uCWA2a7yish2
cfYdQSeB92qgI4AWIY7yhkUqOQt2omGkMsOVbViF1rK2Miq1HfMnbc2DtRYY2LGV
JsNLXvp2sogINbnDd/UOIFn1XFtozq6BdHnvpaxQsLC+1jfzxIyI4wm5HAe94b/P
`protect END_PROTECTED
