`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
67VqAytLA9DHCWV+gzBo/eKniDMStjH2FSO1WRaegedG7qY90NtJ1leOIEuvRkE+
qgdQ0GMj/q0bUWf5NAyHQhU1wOuQzHaARwV5X7qlaXEpB5VErYyOaipZEhQYPZDp
ShJXQFGB8I1KoI/hAshvfEktyMi6GgSzPAp2R9GIE8yiqNVNS4BEBDn12uN2I9gl
TOJvK7jEr4t3HNSrRO7+ka1elulM9xXab8Z5EPXt295spvw4ddPf+sjmqtCWl5XS
Xc8tKKn0J5RdObtpYHohV0cPCwcypXs/yiAAKJ8r7V4F9/EYV1XvHuqdx3+QaHB6
jr33YLZvdOoSFRoitToLfmbOPDK0DnNXrCD3cmUrfumgKZuVmLgSnN98kLSpImQX
cDZmg9nZ/owWJwruAS3m+XlQ1dfyFlBBMSpmmQ3dmL5XqluNC42yGH12M9V8c3En
P2BL2neHu3nwL3OzU5on2w==
`protect END_PROTECTED
