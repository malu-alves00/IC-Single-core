`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Jxxz/3crMk5rOAGucWmqqNZfIwqZJqvIpI+bruBOTLeit/IyJHAP2CHqUYkX0GZj
y85X//6oPBhTL2m7icLfGN4xOSwmytnTlFODm5yveWhwdI3hY53+J/Ct4nC1COaV
xTgbocdcGipyZxmPMU0jLxpIH3De55WlhnAGP4XK4f7rOuyGFPDisFn37nHPFN1m
DutxzS4CX694/ppiMGXWUEcTGtBP+dOdfkHDjfZIXu0rO/LhhMzw894UeDGZS9nF
pu5Ppnx2TdUd9Ooo0xR3UCDf1LIVCLNDsEzghLSXh30+Pp6aNzHEhQSuk+amVwor
swqTXy8kyOTX4LwwLjNnEKe5Mm5e6eB3X5+T2ERS2WonvjxwjOGOWk6BI5QLRZbu
B9Y1DfO6LF0m9mPicKwoBHQ3MdqJDu4ydoriarxF7Kj2IehiTWrMmWr7zgNC2BUZ
qDEL9DqHm/XP5xhLvOufqsmd3NybJHHsfgrDVHAY//5oY9O8bwgGrv82zVb6x0P7
KzXaGwRvVGsOrFJ/j/KqE8oF9HCZxz7HCcvx0q0v6Xgjw93TwhaasPv/O+vRcJrg
LmSj7FfEYAOoKvsyFDsgWvvojifvnqNp0/mnn4KEb2nXo51gA7w2vGLZhPgH5WlH
tCiY0feaMWLr9GDo39QznSUv9e5Jo0o/7RBOJvbw+KW9PSrxINMkSL9g17fzZlxe
SxmfWZ2+oD/3tgavnfYalChMZAW0PDKt8VdgnACWG4kraf9HnCLnUUExJ4bz1vMq
4ZiLqLW7my1Kf24E0D3u1T0rUeH0749QT8eWI5GQL78Mq+/FpjcECWzLE6kmxD9v
r/aafbdBy/0VNrcD9vvCU9GOi1kWD1ldW0QGlHIr2tjBHk8tvaGQoQH9ddZnceUb
VEN5NvujfJQAKOCTh8RDF61qjQsSlMO32W2EaIlX87aRVmrtYUZRLKHKKtlNgTaL
zv6wCsKUEWQv+QjSPwXszEjEF9aIrgYLesLve+YWoUjOVIAOUHPvPSAfitSfzlI0
`protect END_PROTECTED
