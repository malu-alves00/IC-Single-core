`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aI7n2DvHppwvvm39Go60qnTA9lDTk3+aqog/pLnqkBUQ+D4T8RYe9nJRnSWfp/eS
gTQrwKyK1KPOjnXALgPyZ27bY0vu1Y/fSJo6+pWZSkLE4lu/zhC8YUIkEmOHOhHq
sVrSGHZZU2s1sVyIDnXqHatRvjwOumbGonXlyZ3FV/hJMEGe9tFivulu2WMK6BE3
sSShOJsZn8MeCdiZ8khkFZUqDKclsM9mospiUDBxpEhpJHjNSE8jAAZeT2Mm2TQk
xjzHru5vSQnKW3kUXs/vz1ZUN29yi6zyfwm3xW+Ad857fWdYJM5HH1LtpZ1R7joV
fDEgL7xBi31WYWdVDuNXAA==
`protect END_PROTECTED
