`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8lRHMMXgv4SUaaXvMmuD9XLjRlzoK273xi6QwqvswCqI589GlMnnZiO7URh+YrBU
wzf67HmXrtBtCahAhMyIIv3/Y9DB7tbszYRBHysHZb30qEb54NDnyLcznrFJP7cU
WoZWP7k5xXi0KLRV18M934gzUGhBFhsSiLoAlwbVLyBcCfO71L2YFzxkZokGHJRw
VdqxK8PLupd1Q37KqEuwRk5iF+lwE6z1M0cQa5U+TFT+3ddym6NwZAuugRVv1wSp
Msczjz/N4NKQEqjb1nUot6JyUEFT68Mz2Mj/zWKR+D8zAZ6FPlWtKccm9VtORdG6
9/Q/5HgDA7Vcvs4UnqJIGXtwoWbsHC8H2C06T6i7397VV96XFnz6CrwMILONcEjK
Icp39T+q/2VkCzNJwC68ZjXffpF4HufeFFvc6HaDla4oFaSM54hyDVi6ID16ErMA
yK4VZfVUYD8X7PHcqk7Gkv5Y351mmN/YZFUy9VwG5MMuvzHPyDSguLnJY48dHVMp
s6Ba/lls787NfW+p0kAF8T3zDDMPZvdZuVZj1Uc/sCuoasBoKBO9yvAsEeJl3igt
U13kX5Sr3ZFNJCTx3u80n/GKqTcS4UFEIf1lJDQtPKafLtP67fiYB0AGnOW5Yr6Y
hvf9QYgvLWp/EDHRD6Mkq0LPLrnC7V78veBgTq8fgjhg76DjWLBUQsiCn/zcCsBy
Y1xjoaBI983f7z7GTW/gT1RUieZAVPTyEujkZ9I8Q2ynXoTr/fIGRIgAiIs2Nga4
FjjW9kSSI/Ejb16iP3P+jYvdTLQzfATdsxn6lAmUgnRP7MO1ahDkFrjZ9tt6WrA4
fAJw839FquBImnTAVYdyKb5L6hSixNQR1Ab7yMS/izRKfA/6Zn3xGMiti9PKcRx3
UTnrGTR7qXcUNYlj8nZ2/3rEHNvVbHt9G9qy7v9gmp2I3M4EXEKeszZjxsTiYb3R
P4TH9i0ehaZ/DghjjtPOsL7XCRpLJ+F4wl5gZBxr8WlABoMPA1b1l/I1Tp2/5cFW
lAX9WNQ0U1zrXe4p9Ieey7cDvzs/Z3p1M0R1P0ALNeHktsfSwgSvh+zilAs5c21/
lMcG6kwTaTia81Zpbeb7jABNNolMqFGq3DcfWRGJeOeFMSQ2QqraB6PKCyNkKKU+
wxjg88vRZr/UI5w7ucUn/c0Cgve4lxjhWB/NSk3t/DtAUj32LTveN43gUxUI8r0C
dq90bzIf8c3mLBiJoA4r8TiUQ1PBYe94qh88B+MNk7P2NPM+yHh92VQsJSSOGd6S
rM1oYc/tohIzG3uMwa5TzTpIPrOsBOQtQqFO/QnzZFygoQNlxgskrX0JRqD4Dxjy
bwzt5qw2PPfa/0AEkDqDp6NExfY4ORKaX5LIbSel9NlVfVBrJG9TDOidk1grrAzr
Co8S5J+8yH8/qt5hE3CXVQO3yJCUS8jsTzwzDvLj5RA9ahvq7oXAE8D9iRi4CG/W
mFMZLJHcsM8Nu+w3KsU8ZmFWpWQwIn7NUQ/TUiTztNGBGvbVzsWP9tbosFLa24Kf
KRz+ctgBCl3CJc1NnWI+c2m/OElmz08S9iAxjJiwo2qiM17CV07SM/zQ9Q0xR7uO
qsvRbCh1luCSJRBaT6nAT3HT/e4aXzsV24Lr9TIValL3nWedNPh2zyY1S7WGCP4K
8ayl6VQEaGizo5MrXOwlSHMfIGzd8M/V8iwOrZYGXO8OOop7ogLuOfxotX0PJ2Ug
G/GCSQXXHw4SXgxbvGX+/VCHxN8fB2MWsdpit1MvduKRQwmDT2/vjY52rMt/vdwK
GCfi1RYTv3txQm0xw3+YVM4ngIFKgBU0hJIK9Z5TmE34BaYYiOgV10y5CnEjjScs
+cnlzsm9+lTEHRHIZccOVfpKo3G/dS68g3FJO0Ii/ij99E3nKTQd/PcT8eoAcDSK
8059SgIZMYnKWZRQWBMVFS5I25+S8/eDSWCKZDha878gl7D4GZ5utbje3C7Pklfq
PdQecCWYKDRX7KcHtucMfqzK+jG8yq7oQmczEqejt36zTyTnwuRukg9sShz4jIJi
sHjsHYcMCQaALDJTzxJgvld6dl7A5Ji99f0YtEPUd7mylsA4hz3hTyJeybfy/ldN
/2P5w+n7DhoduU2/f5gEeu+4DOjoeNkGhbzw36Acr7w2P9HHv2zxRJtUsStmaxVh
3SEj0R9T/H9vSRhnC04ZbKypDE/GG9OOofiYyEju03+kImaLBcdx454mcUVmO11Y
Dize7UDhf1AxdQ5Dso6soUOFW93h5AHkUOjqSbx7z6KHOJCNGhvEYTF5o1+whdwf
3JZy+YGNHGIt7sqERf1vnSxGJFUo1/IV+7vylKKZTmNobIWyKf7F1T4bS5bW2rkF
QunsRHfIzk9g7dt2djPAOJrdYc0GG0fTeSiL4R0ZiVou5j+uvXxEuRqmdYaJamjT
l8aQfsUtaq+rKOWfzKft1dtuhYDaNUOvKEQLaVyz2w0rXGsRWkgYjuhSbvIiuYIk
sg3lrbOr0X82H0hIkBwWnLsfWlNjTNaWM7ORc608tUYqRzr1kD+Xkedlj2uYgh6c
VO+frA3BuE0kMO1FO2TPW6thMgzjspUPJON9k1H2sxsXGTOx87agJMcJLtysKRAZ
iRYVIxEq+QX6vzu1tb35kkb2c1qvyKvPU9muDV5VorxoLhW5qPhbjcGywmbJRpHe
sNEtc6dAZm/naXLv6AN+8gkIm6dupv1PGKT/IBPI8Xto6nfJHwxz5fqhcauaL4gl
qrgi/Qqw9mziFlGeazZK9P0N4uDypI4pIEZtud4Iy61k628DAPzt77YhR9SEoOdR
lXzfbhbBYump6614HDZyZKu7gTb1aFwhlPckM9D2vpkGERDRh2ZNxnLLZAWpMs6x
TyyX3ny7BHgZDN5kbWhzrg0jxeuu+Fct9ezHdjsjyH2hsXXtAfjhggC9GEIhiOzE
ZqHgcQu3L972c6xtY8uJ6k6rbeoLuSJNg2WqmMhEvVQDMe2zmNBEs4iuPqwmgJoE
sGdAUCU7Q3ZX/4CIcIEP3q9HSyRIJ3UiYPtdUFnyqgMmyDcBAUd3TQB5bSTjs+iG
NcWkTIU1wwJZGxGeNKB6PZJ/nqh1q981kT2dtSecC5Ql8aZZCYLvvyC2ERaveko2
VtJ/AhAKd0Q+3+IOlxvrM+aM+OUpYEEaevHr+BY/WRkJDLhdZw/UXppKFWVHsfk5
g2297cGHIm5n6oE7bHur/P2fjeFNwNFBoILn63/HWXxF+jw9uVUPCXQWJwDKSqvD
Bqa8vbh236GyLQp/S9+caS7aYW1k4SDPQGk50lSVLn9KFyoo/vvWhyVS7L8t+QZ0
hWlEb4M1Le7//m2BPwhPavo7+bBIv3Ntmufr9kUTlKO57xkS72VvUDdI5NVfZ+nJ
mmPuDV+ebVTcDMcwy1BvuXWeqtfyW3MezqmiRTOOnehNYFiSUrc9f1x+HTLctOtp
h4Ils0SMRn8CbGmmXUxo4VMzbB0wZdcVaqzSziipiTfGGgBDvWomCdqfgIcsWKmB
Uj2TmAVZTl9tdHuZ3OczhS7QxKMED2/LgcURlGKC4V0tV1bvBF6snRlMnLQjpeEM
82BWbRchnMk40f+Jqs6KLfM/Mgn1OQQ4LCoRl5Pc0nXTlcQaOGFpaUlZIwJYagfs
Ac4O84/0KJOrGCvRTNRMMc+Z+YmGcsb6nCVSorUSuvrc4sdBz+CPPuJuQ0RbzmPL
36MwXRsibh+zWglro7PMHMYUcmd2KeXtxERzaCWcdJnpgubD5/SvgMKB7UoM+2sg
LS4yl/cqWiTZzMeMaEuSSH0dX5wmyDICOkRYk6SPnLH7DsPDIHQZw8n1b1d3o3gr
DeTU8ajxYXEDkKzQ7woSBf1XFLKdaaukL+QdfpLZrI4vQYQSSA+t2tEAa+TMwlP4
yU5UdpQAHiC4qPCN7kdP7FyVZoarEn400dcD/V69pCotCubR/OW/DbqVZHf1GKJe
obH4vUdEAP6027tSuuzO4Xi5ZgHkgQ9xc2VckGOc2E21pts6cBwV4q/XLvYwFew0
0gqGofo/94x8UKQMkAPLWLJJzkI+6doqD8Pk6K+x94uLKWnguRTnA4JrlDyF7jNP
98zh0YEw2S4EBsHqqEgLLLdlWd/jdvDwV80qXRS0zD01ojaZPYfXzznAirH2VuMj
cGMyqmCMEmclJJEzVeWADs6sv8N0s86R95fwmO/QDFYBcv7yiz6WffplPTKktyV8
eD+drX0oBGyHKKD1M0ZTHrHb4rgQUdka4kFuDTdwpGRg9lkJzAosIekVu0sqe1nt
gHlLiwW1U9fOUq7RapWIqiJK2VDZJ6wCx7gCThaZZh+m/qL7QfqVKWnZH6dKeJid
U18/uEB4HSdsw9GZyiR14yGqofQGj0j7awmlAXm8Z+cysjRghy757IXpXjmXa1vQ
GBjRHzmmmEKwt3kb0vWvliIfUMf4mv4q3maONf2poDAnlw5JqaO7xkNdx5gJaf+6
`protect END_PROTECTED
