`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
F6+zbZW7k81FIRI9bpW949cWxq0LgyfrkqMptb7X1Qqgq1O5zdxo1s953njSs555
iwLf+IpHA5+9mUHhcBLcd3COe13xM2rxjyrJxbuCbiunNa62nVMrImRprA7GjSji
U8i8yPVAQ/yXp/P+NLdPbkLEPkM87aqBRWh+h6MA3+PF08qJ2szDabx+95nTFg8W
O91GAFXkbe1U3pQU1FPAcEpShq4eqUEo5ZvrnFVoQ8KI8DR9NGpddVX6ogujmBTr
9eLmICCjPF9KM8dPtmSrr+BjtQ73EkH76il/QhMDeqdkKnQ+zO+t1zcV4XgFHZNr
mHaqM0lJNPDaGHsJEt3eBJzUoWznDB0YBZPdy8m1G1u30QX+NeBQaoKek7FNAITE
m6g9p2+HPmKkJHuKBb49xVZEE7MSVJDyOi+NRyn4CGamrkgmgENaLdHzrXYytFk9
EwUCVDCdQH+mprYyPo55ubNhJ5xM1bVC2hHToNHg4lXceUcAAhrIG+5sc85Lmd1P
tpImVWLDum0eHSC18rfKoqxMVdSKqaF+O+o1mgEIeU/48IJobhi49kaYgVSuLxYD
aUwLVveNooRCb/8Ttw364kC+ndOIymrBG/ENuHNxdLym+JumW41+pXfaHO0E5641
z7mQ0Lfnbw6+CBtalvgQd+MMk/xTiWpzP2fBTaZP0iAirZbyuzqf0+DMDbmtc+7S
A1oXB3rqedRsoQUtWyZ3C13zR0a5KuqC2Zvq28p/3kiJrW7pZbKtjnOsNFAXevlT
559sG9s58kg9VtrPZ+uC1O1TSPPWUI045R05IsmRp/JpFtrKHw2SItV66SmvuB5/
a5IxqGg8uwbvhg3MykdHpjugk/oeq1Ovfc4n1XMYTHCxzqtvzpgJGgdceqzWuieN
rMiXv7EExjJzvFB5zkyz3O/W3mTgaLZFFm2ftTtDJ4m0fUXLXT7h+292IPCaUj7i
LwAAllbLLfk7TkyBoe40pb0OMx4uHR4ySDPVs65elPS0o+XuWcI1drjgT8jBD71M
yoLUeOI82Y+h2761BF1Mq4FHSibVjq0b6Av4ghc3oIFY05PfNl3b2AvGxRTpt3TD
UT3y9uz+cWC8jL1bKApUCpfe4sVyOppv45EgDySRwhwEfLNmYA0M04VT/P5TNWq6
0YeFYPPA2H/V0TwKpjz40o0/3FAgzeydGwYZoQtgQo7mjscBnKmwCLrg26Ahaybi
iT2FYgIyx7WtJT2Ddt+5w/PRQmr2qy4mm7tkS8d/brHTkNyVUK9PkOPHzFeFs2bQ
RlvQkvDGJvx2fmI9uvv7uldMDPVKF878S30id9o9ifkytGkX1BnZgvxo3j5aZo3l
9EMdQaZcLcu6pO1fY2InBJJAQ9DKFcAbP5/YPC7Bj/EPXAIGhHdygHnJmrvotZa9
nE+dhRCWQDVqtuaqqlDUEZ2dho8RN9v6qkbx9+PyoCPTG0M8U8frmPA3HPfVx2MW
2aQIqKwzxbeuEGfg4S1Ais78E88lHAf2bIXLNjR3xkY3LOyGB3ObgLZeA8xM6uyu
HU84vl5DlxQWBSmS7UyNuOfyEqBOiHH4QrHcdbjQzPbck7mWdGWyBPijlmAEra7s
f2WL92RsvV8DOOrnCho5pbefLtYAxhGNagoXXELXg3mGvQsY1SN58pZXn1chQ4SX
MEVtvwR9NPWvy9CXOSK7zeeModHhnWbOXfPMwY+Znl9AILDiunWCdN4LCKlFy6ZM
WGWoGcb+J+v+zPWsiKQjUSq+zTE+tJJsSWO1XZEGk1+YBxfWsfn5kFcWi9qouWlC
gq0Fx1br5EKEb6PuQm4Taa7+QDnCYJSlnrCRf+2FWWsE25rRO56vHrzUVJc4xnxX
g8mph7hbdb+dqagVDk9azjOZDi9bzodS4PDECiH6V87Z1QJ5iXdfCy1YyxMh97WJ
ajp/rcJ1XIfpwBFNww9VZvwhVsmytZUuhyXx4kx466INTXkQyav2hTzhMGKAnbwo
EM6M3y78iAnTvHKNsbA3XDR+DFvo9X3MwR0Jm/0C/kQhEaGuW/qW4ZLHjePVUJ1g
WekiWmHeKlRHxIESJ9KyuumGp2UffUWrS/aB46gJxdfM/lTfuujhLYfXQvmUCXN7
Cj5wsxdoY+sDjr1eKQTcpIirX1mYgUJs2njDQFHpydjlV4SwPxqtbLX/VMyOAqkB
Q89w5UsP0ScN5ExJjPHEKdQ1+BLVUxaHiIz6fYY4XglmxS0KeUEO5PCUaHwHaFmY
x/rzveitkMSbt9TYBcXWRw02xN7xbsqfS8S96NZNo6CbT1pqjsFMXL/qRZScUJsa
GHgkQ5Y1K6MUd4MsQOwd8T35WBX67HSs0TOAfSfvPT6uy2aTm9H18wbHujKy7t+0
WejAv9iwmaeFRv0I01S8k6WuOLALHOlUT+StbUnRtT4adQv170CYzn3zhUxs8cBG
72kQQyMTFCLrRzxYwAj7h2DS2nlPXfCyJm8FX6CSRGF7fKpcbhcweCYlNOVn5W60
Qalro9uxvXvUQikU10R0LFFwu1KWqLhjwXFa2ezxXX41ji7ZtpdZ+tXi78BxGi0d
3ecm0yhF1rB/Dckbwo5hYqFkcSeoRlbalC/lmNr75LC5pgnUBNu/mi3RlCoBGiNs
PIWOuKAWeJRR73pX5d6ohwNi9MFxybpJKbCbYcoABpwht6DNv1uvZZu2erJAI5gu
iz6E7RZW46++aYzxx18pkBrauuoQFCt9/hBRIltcbC4OfZMSGWXMZC5or3eyLd4U
9WZ7yGG25gCcGTjN0CSfqh57lpKQU1gpfOB5qWOjV8Crd02/WxeFxczCGXnQo23T
XBxYBGxbUAZbpvVc+FhCEv51brIidfE3otO45SX87uvM4Y9Ya+b9AJj627cCd2nA
d1AGBOU19ZUakT6XXj6uHSGR80LIcmlCr4Et43kcBIraOEL4OIX//XGfph3ZTMpx
IJkoG7R1YyMxUkgWBoV4DktzUMPl5vN6BMaogy17L4kXRJYeO4mLyDrW9Dj7H4Yg
+neWJUUBZh9bglNTyaqT4qyysumXnWY+aSRSbmGtexKUxbw9VovNHFNuzAXeV0Ib
o12NpWnOAOyBuEZyL/6RS8mNcTls7jwHDyGRsUqKQkQE30dU9nQl2J5JI0yUIL50
465wQ5LLWv77LR5I/hh3vtMKGnaON+oMs2JlTCMAqs1ULMnTY4DxBIheYFhQHdHf
Se0alSMF2ryublT6fWUsAx1EcUmQZuTdTx6INXwAJtTQMNVSlrcBmqTRXdqwmy2D
VqhFNgHaaGzjmep9dbMj4g==
`protect END_PROTECTED
