`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+9aqk/4FmMgLvNbKVhhOiBus+YvfcX+cn4pPKJTMc3wBhY43ER3KntM3IZyo+pMl
zpfXDfpWjfqT12B5xWfi8TpCS0tCf5Y5wuHK+ii8UI3hYKIYY3/miqY41JnrN/v6
6IbmoGbq65IKeKOX6GEvxqi/R6JcW/uN7zqXxneq3NUcMkDd/Sf0pkA1qUWdl6lI
ZMwJHV/cbGPES0Qzs53EwS5PgNbBXERXg3B2B2r+ZZZ8XuLCO53hoee6H4xTTkCX
/GD8tFrt7MWD1cfX3VJ6be0mmdWikdtzQOfrUoCBabKxJndsYtC7VhkxidKIuBgT
jQDCc52W/CIGU1gNI+ZOpHIv4Nq+DfZ/ySGUTuFH3Zfdy9AEVgZPiEZgf0uy1wJL
a9D3J4SHBDW3Ni0pyk+zsmNfzlaRWmLgEUimtu9TlIcFE0y7cSKl7eyStPyo9Jlt
cYqC4KHQr1iqvDocnOKTPycQHBf8Vrb314F7pszmpsdVbrRDCNg5tuvniiGFfY7a
/0lTFuW7IIy8F/KGak4zANUnutj8cM8wWMABfs6EjDoyLF2XkCfWaWkp84jZQvSi
UxeRfp7BOCjlYjwAlTdOI3ty901+hVnDXkk+Rur7U+hmjBF8NyUjH5jhuVOW0cSa
aGZ+jQ3asGTPXOR5WOI6dJbj2n3Ipi5NnxixgYrvmProEEMtznII47coQvBwArIL
OOZlYFOOJV0GGuGANv2vOcBXBuEL0WnMapGbaDBukbi4SP+K4EeaitWOySXDqD2i
rMUz9CK+kO/Fm7Qjqbr9Voq4TeMSY2l43PT5ekk184K0kKmqAnVrZ/Fjou8IT9G3
YVEsFyRSxzY6gHdtmY2B3L5/GWNb4qtJ+cRHiKegtOgj2CA3Ohekw22pcguSFuYn
EKcddOZhgCjWxINig5W/mNX2bblHXn0PDWoHHLOQOb4=
`protect END_PROTECTED
