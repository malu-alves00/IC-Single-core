`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
F0eBeRCSRcJrNbFqxhgqcZ+9BfxmmYbVdRhs3wTspK/izaPxDpL2dBVHV+UVTwnt
hE37vjc5pPWtPUrtpYsUu5QYSO4psdE5RjgudZ/b7dHAUohPc2K+4mg1XhiydOMI
hb3sgo4RZNKXqmqxh3/fYaRzluQT/XXMi8maXUUClx9zoXDLddHxqm2OEprn/Jg6
z5c23sz0lxjcqtiv0ocZvgxm0HRj9235PNVAmieVCj/sNSI6gVHnrL3Af/8Y8qmw
brjFBdy20dlhieiMWAk9xAMdjjI38Atx02yX7mSXWH4PEYwCqyDPb0LP7mFLqWWK
vAOz9wHo1IN2ruSOHkE4vJV/J0ed4/q4nC5atQt5ecSS+u06Y9rhB6Vq6pvCiuuT
Qwpeomy/lOge2AKJLogzkAkGmx9hbyBjQlNdxcO0nqUyZYhkaeAIbWi14cTvOcBw
w7PRM9t2svwxcBJrNOrUP5mwjud9+7uxgHLGuOLQO2YMQQmACOrHOVMYNzFFbvKc
hewz7RttylljGlHFJcUyMK4vehyDCLdWKSkTHCuAwrTcnbRyTGOewN2X3aNcId9k
rkw2eqaeCJzBtg5pgAhPtJt2aFjSQbZ6BxqJZP2QUjzsSYfRDgsrk4jDR7NvdWRD
+az5Ztt+p/err27gx14WhUnaYG1Q3/kcm/rqIcRrMhY5+MP+vhI9WFBcfp0zDybm
IW8xQoSU1T46lG4xjB7BgZrQsHroJahDLXNuP8Ue5BN2Fbx6Y2bL9vxsbeU3DNJz
TocNm9O7Yb+6opHdgjW04aKteCVuc418zV0h85aO/48Tw8m9XbpKmuxhmYLdiwQT
ILn92CG2qFKecNb31f6qyQzitzejL2jFanR0nKMQPrGs1J1XTPVS9Y3HZHaTBQI7
0IDJJoB1rXwneG1jukSfjciDl0u1FRtzpHa5q6dksmxVKmsauaKtaDoXIWD/DMCB
L5HLNQHVFvfSm98nI4Kb76WleAglTbsA2Pe1y+TonWgfPla9gUI6uxr40FIXWisW
dRFcwlNpGU2omudGERNZ58/YQOq3rM4k9st0kjtmM1lpU/McVij/gSRJQi0yHtUa
Jpj149qOLsLLShl46VDQh7HbRCnxVpA8UpIgeAuC4UX6u2LtNcbSwUVkjfsjF5Dp
7cTU8/Eq4g3YQScjIMfcBxIx6qQ/4bXexTiXZJGiwatxKBCIIMhtoMY1bMu1hf8O
uWQIK2vOWsk4eUNiQwNFPqiIj0w8m83yjAozKGtl8uMmeOrvW94lCDyo/U+LZFGu
fr5B94AVYnFwY6/5lLih+PyCeOerf4r/FpH6oBW1bCqozDY4g+9Im2NQBuN8uuPU
lacqMC1Pn70ltBGfhXoLu2z6LvNfFbX0+bqC/5Es+E/VHc0HbF9P5g1gS09XaxBR
TC1vIHKhNCiP9wrdKOsPgoeezBVIvfOZlSNi8tqdgDK8D5wy2B50RWPk8WP2NIhI
ELob9hfvipBYTjjPHjPwva3F36XUtx139/TCsp6InrZwzw31WfIUM1PoLh3nczW1
HyKwnTwoqxYgbM7cURmUROhC98YHtokhMSTWz5ntXgziSW0++lpYAMaT4qZDaScO
l3oHdccnyk5QYd/q4tASbTs0jK9kGLohLi6dTK4USubqXjjivJuQcuKgK6+T1xHC
`protect END_PROTECTED
