`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pcXwG2DfXqCQA8bLMMzeQTD/MPrBUA2cR/BFgGa8G1eEFNbgQk88TvkEkCGdYn+I
8TbeyaKTZM7Ph8keyL6H6dny1yVbi7vPOMPZuAaFfm+llIYFpT6G+D/yuPNQ2oA0
w5j1zQy2JL3/z4feh5zt/b+EbC+iGdnlYXpJ7/Fgt5Ki/UzNmNcoY9q/1pQTdS5r
yAGFd7V82LyU/ewkPmshA15rPLiexOlB6jyfkxvx1IKhbtVWBG1V8RSM0hpKtUzb
Jpa2Gu4+0qTkMolO0MAU+vUbm0OQkBUolFEWaAoh2Fh/gbDk/pRceOZvxRo8Qz2o
9DYKWE7shtZ4p7PgI+pfhms1B5Q0iNW25uTglc77eSWpP3CjO5c2wlTEZLO6pBB4
HmuVMCueODD4Dyg1QJnC9aTyAvxRt2Ini9HLjgdIeQQE2HCc3L6jGDWuLHxv+HQA
NKBq9lBvknR9n/IKFAcLRDteuQfz4F1PyY5MvwBstflzSAfWYpw94y+cfI/jXvht
59RmJbPtLnPsDTeGdP82qwrkfQCmD37/p8bFMS2webESuXLaigEE3d8ILtwPlm7C
9QqZ9kCokrsx7Hx75VLYAuX/nFQknE04eG+qSWHvuEACRy9McaUSG8fLf3+iSIiW
eY/4sbJ0sGZTq05DMF2F2P8iXxRv/bRmC2bU8ySLtYgA7T95kfVclTIGXJTaieBC
0Yo1Y6CciKcbYfg2z8VVqWHxwCDKVVwb3NegXjbkG+2Zbu2ftfx1OvnJ3/sytk1X
ex+lnnNchF7D8ewtPDHZSr3CjlmPh9Q2+wJdgn8zN2tm5GfiLTuSZDqRjsqrxmSl
Kj8AwWQFyZz+fytMZsQSoxL8VJzCzg1c4h4zhshAVQfSBO/KZcl7o6krtNY7kK+s
nV628IT3vW/plAGqnXywMdgIpCPWCcYBgYIT7/mZgZMNRaioOHqzLyTvqgbB+evV
7YALfzxZj0uMTpqnBZRF3k2RFeKb6lnFhIGPz+A0nXLsJsfBXCDakb862uJ2SFS3
1JHc0daNY+7AhYghKGpeGJ8yfq0/ri2N2WeU7k6dy01LopqfCKz1NWrgoiE8v4PC
WcMyUcHgrdvLLWG/ovDt4NklSVldK68N5rE6BOCnaCdL4L8H5rUJJm6IL8ml31VL
w0hmsoMtdV0H1K1ZMY14mTCbjG3rUxSmVnOynzMVufUf+ci+n2YaHkLStQghuNUt
7XVv63I2XNJ9zobbn9WpUduGtVPT3mfrUl7KDdKfvh4XYqNr1iNKmA06WXC2ZDS+
q/lhLyeJ35SNsANGtB5Z/cRc1v5MZ6h0RDf60Vqc2mjktsGeWr12hYjvPsLD4eJM
+2B4vCmjILrN0yS0ANL782HaU2Fr7bbJl8s2Z6+u1CVLuF5HsXRszWhTI93GOhLu
1B2xXqQjwxSALP2C6Nfhqv3gm2JUS/jhVXmYD4Jv+v+1UZAU/3a3oqC8fqm2eZso
CpHUNK9dBgsXjMHoyJBJxJsM0gd3VBnhavcORflcrcASzdRRE9vftklu1p7XqeV9
Xr+jXnLH8Pp9m2PvFM5Spmi1c4xKuNuIazm8TFmKouqXOk54fUSScjqmv10+O/km
0xdqDfCgcrmuPBfZlP/oJS7JrLCDeZw+nC+ysGD6FJ/GRvQ93Ec3WxeOU4RLpX2n
Anh76/8B6SUXjAljGFfeuasQe6rW8fLweDaXSs8m0Tc4enGmTT9SGKBELaxgxwxy
WNrYAKHiXTIC9IvKsxjT76qNmC2D6145/Wwfyc4+m7oJuwidfkUSLdq1ZfV6Y9q6
/cWCszrffWFcR5Gd7pRecXV3uHfA8wLvR/QkUpRoPPc2aTnPLKFtSIZJruIrAvBT
P6NbSCuZxZCD0DVu46Sp3kLFGjKATe4l6MP9dOIVmfMmbjHt3u+bwTfGNMCoryLm
+ZyKBzj1xTaC2TThw1QZflqcVuX7wHVtryWZpJI6SrmbRCVPbUWd0cV+SByYYkHz
yrH5x2k4ozwtnJJJFEZ0Vr+1GbjtqKEu1Q7rt5dGMYSvyRaebU/7+M7jnW/NI1rb
SMzED8L91JDim2Yr+1MquEXxV2XUFTsbPShFlkyTa2doJUuTY9KeMuvJPhyUeQuH
J8mljXkQyuWDNqaxf50v5QMVdQYhe6GJau1NRWHu1CRVzaz+f333kOBZk0irGv0E
WEja12jWCAwVLxcdd8kTZO2sqefAQbhvsCwU4ZWVCGjAJQEiq1fdnuLFiep+W6lT
/6S3wLHBciOyWMBvZjLnwIffpUySmMeN152T3ykRWqhd5u7O6OEtFJ6isw2ssIO9
sqnpbDCubyoXoRyx+0R+2md+4Quo7gldOKoT1AC9WY3o8COI81l6+UFnZh475O/3
/gO9qaGot5NWiSCuxzo+0SVz0WwdugY+tz42MpXBFPjVRZ0gBrlI7CiEIcZ43ZRa
Z4C+YO80UpJ01EW4vwFxkyxi/mZ1QmepmV8OG2VIO42+mIc4KylWRIXhLxNiMeVl
6aFhGW0H/+kQSjdcD4V0aSIrLXboMbhhIfGJz0VMwYK0dIcsyE2e3GCbTO2kxrD5
7LWfSlkNxyh2PcfYpUlRDwGdf9EMcKrR7wL2le6bL8WRaiPTjVI/bOvNVCZNhmiK
Up6XkbrKbdj8Cx/8CnGbUKzLc3bQOCDnsbyQpgd7Yl83HwwI1KyKjtlfHHmRBi2W
lhwY17LiVUdGS0IZ8613AHqaJTcFZeNha4BXQGmimHHMZlnEhT+Ovl0F27rfIpIY
uu8C8zKBC7SuXUnAaB5h4/uU0CwSBC9+ULp/JFZERnRmAgUCTjw0t+oOuH+Hau8B
or6TjlGWCIwtOpV7KvxzRQio5vsd1s8lK/lCbKWNAUq2Nfejj5RqCkI+Bd9d6qxQ
qJogDb+dAdyHg5qkGLyALXJshXh/Qkv+dTjhnKmoIMOIRreeFbHm+D9R+niK827f
H+exBLnPtu2PMmMSKrai3fGGRzCJZsCGTjbH6iYP8w+INZyuPs/Y071PS3UIoAOR
93Dvvfjt3w1ktoqtX8wbDAcryPQzEDtjqBfsvguhOYq0Er59Vm56y2TeSkVMy0q+
v4N6AbjQLp6NjlsmKnjB0YuktN5eQgP1uWSBWkDu8iTPhFBVxX/WBJO6GRNEfl0x
n/i9Cmqbf6+b/o83WHOWMnUCHTHvM4XwtIq8zc64s3M17aib4vPmDQ/AlivbkNT7
a8KB3cSHvRLV6MqtMUTxQlHOiCQMXHBoN/FNSqaUbBJYUoxJ0XafXDCkQvAv+8px
xJoHW1O/HEAegZB5KtQJ3yUKWA5RK6A1eClJHZz3nQEEZJrypiqsqilarObhVyhY
a9P77ig65kW7TLzbwC0yKmmNI8uzDB4TJums/Sc94oNL+FBylDd8Sn+HMRcV8ac5
oHYN0svQMxcZo5Ap3TJxNxO7luNOXQWELFVRdQTgYG9deNra7rc36kFmYZNcmbYX
+u8+ZFaPbeX4brUvuD5/aI7ZePjQiMSPo6s0zzLDpN9/SnAkB4sAxUUa5zkkIipC
gSfZoW1b0YC2CapP3E+Ezya9XmmfGgQt1d2jc5POk5TRTTqB08jsWRanDw8xSwtI
fzE2J/AoouH0w66lRhGXxUmKQeKmx8HpYi4zIPaoe/9oCMmaoAlN1IGFkIYc5eFQ
zW5CS5hjEd2Qs8K29vSF1Z3BHPvoEGZj2qo789xyi6VoEk5G9bDkjNKFMLJHoQNN
5YHO0eXb9yGJcM5oaRJVRyGY7ijaC05sEbRdS/4P4RXo1tM0ARhWtq6Y1u6WL/ab
od+ltrxXCMUoMjW6QP1w0/gaINweIlxDkG0U6agYPjUfMz/wZVlLgsc2Lpiv/Bkd
kJGmyI858YuTEkJCQtY+gjzTBbZUZLZ6qif23fEEs2jpCMSUJFPTa/eOsuRAqbGG
ME4JMD8F+3OedxdgEj6WvFVyaYaHZa6jmdIk+5cFMtrD3eZZmrIQYeTVehMqFYPR
zeno9aRmeZzhMvxwQnr8cm6ZaLBQUlfRdw9qngrCBYVRItz7rTD5Vf6PhhDIHU5S
fTsITu1lkn0rX0msKE3BsFByaS0m8LSRo1MYZZUpFWlfZVL16/EwEvckAEipnzYo
sRQcHoWe2PZfNm1ThdO6+597Z/9WnZfAX4AWeWhx7/3ZTt5NZdHZD9NOpPZnwIsb
82BnEvkfgOgm40eMiIfaZmbaxh7IEX5OcWk7vqpBGxHzb2t12JSFbxQYkcwFwJ5y
19g78YOG2s9Mu33g5RQTqP/GeEqz4dyiOj5TQXyt2083lV+TcE2USs+5wA2Tfuuw
AndzLwg4L4sVczneN9tl9MnSsK+lDmhsGqXzd36SeGFHYSpua6F8goKkSYXaZXXu
12gAt1l7dSKcJX2+nfd/8/JHUVK4PcT8X1qVNvs9DbQU9U8bkcWUMIwLLsRqW+4Z
1RCh1zglB47RezLS4u3tlfEF7F1wmgMBa42FbF+uDlIGqSHZ5nGYLxIoRmplVP0O
Rmeqfa1bmeHcywYBeMG2rd+ewdcdQdkx/OiDcV9QPbp/nFoDIiPJvQWBQXWg5ifY
cG0gKwfTGbY4LAW6s806FSO7mSE8MIwUcuZp4rvDekOgwPVs8rKVrtz8FtGApwlt
3an/A13glRF/sB4lSjQMNYNq7gNaEHTHfwuE5Xs31abwgrGVhuHFcBEJUTgcZ8p3
AbPwBQM6ax7elOiXIUl8BTKnrSGTwZfzDAsa9KkTYVPEjVpXXwXXHd1VRt22NE+e
Wm4sQIOhvolLcA+93uzwRHrYiUS81ZTdZfUBUq2CRR59Qhja+0HNO8AbtGFIqp2x
soHrOY7KEMmrNF0hYd/JbkjNxCrJbdD8tXt4qrwSQKArvPZ7+39Er+u+XuQoVqzo
xEjeFz5kCFcSmvqJL1PdBvO93DU6/++PsUNBzg4Fo3/mJfoA1gr/S7l6cqIUYeZt
`protect END_PROTECTED
