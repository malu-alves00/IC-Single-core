`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
49ujFcnCb2i4AHKH/KW5UDkn2BAbQsYaHoggK+ZRXG8A4z3YGDWYleMyRSINrq+N
s0N+5sbSLMhbnY59H2fjEnV1eXBg36QDSoCW+ilVXU4AXd9fe/0W+f3ebjYuI1Xx
Q/he5b5LvrfW3HWnxMPb+cxm3ThRD1GvaRSKk4fPqJ5oelVlXfklYJtyFHdSRYHp
gJZzryzkz1VG4tDKYG+Q2vaPVZ7b+GLnxHk1kG/iVj7L92Jn7D8s3yjoLichQroR
qBTC1EgP2pYHYeo0OE7s9JCuhQuUKv30DI8eJWDgJ/3zwJb5ng9LvrGsbfKQrQbl
NUuAwHHgnNvPEftNJEZr6gwHGIlSTth+ljxEEnr9OwLWTdZ20dSOhojJe/YnX/3C
QhYzqGTBl2sxGf0XA+2BDvRdZ3zLRa1GnKDLsxeNwnP7ubI3mnnEhBgd+DmUsswM
JahlRUeLG5JImFvrbYYEOY+KeZICzR9rcFk/9DMCXJsxg8wW0zI4o7yjWl9sHiV/
WlA5xIno3LtYwJaFcsF65AXSQ966mXPSMowd35U3BIJfjzRvdXSV8r/fi64qZB63
6cX1Nzi/aGdOZCjwlJC3QqkEUyBFEQw+kUpijxycoPOuSPCcgK1+VkXsYbkNkrhP
/6IIi/bEu/g9wj6s90lxO1zUjlLq7nCOXBdmBaYgACjtxH7gY0R6LHuwEQHSpVR2
BFB0fPyTORF/9QbdfCa1hASNMhPPsLi0AsBxIRtvLtmrd0RL5Z4ljECiUAHvvuH0
TKrLK0A3kKXaHD8Ml+6AIZHpMhhWT+oE1++QsInxQF0N+hr8DD9WXcbIHxCDSg7e
6ogYFpAXLWTa0pcjMtFyfjCu8t0t9GzoZ9AQZVPXPhAFXfZG5I1+l204gkTupDTQ
o22K/9NshD3hACty698fnNpzeWqWoWZWllE/kE47lUMbz9TIuOPvMx0d67BNQ07Q
0A4MBl3rbKHmO0nGJutSu8SVUXhFykAxnkJkDMIt0XSIw/Ryv+SudFSUci2Xywvc
sgXuhHvybhobBLlnSFHaTpEdxV3xKkMgbJcgzOYE7774vK/ockR3Ks2JFPouWFdJ
Skq6c9Zs/q3L65llQUOJC3PwHg7Vcu4pQYmnREvgDLvyijjgrBvNs8i1M3h0iKpx
xXjIgPegEZu7hiDN7QS+0InLpqUOXGtWLZHVp1fQWBTt74sJEDKgpRvAAT8kOJn1
MfBNidqKlhb9QPwrTjZomF80YV2YgViv1B/QAuC2I4erUtLxcbYSLCJUVrXWQHa3
7GoSMOLisY02xS2u8WF1oa1RYq8I4+8ArqkEPj4y93+37P+YhJ8M94tX8+4sDX6G
QOfTpnYnq2TdOypAdE7+1z1b/RCU2B/g2yJHhOttHz7BUXvKCrvCI+BNynES6XBa
mlS7x5MKv4Zvof6Aa//0AdF3AZd0MsE6afUzqxvRmpCoPZ3jK3WfzSD3gfRebSVG
Za16KqxJjWlOXu64f3DaiOupdeV3XKFeu/z+1+xmeFEnocPat7qGs6T2KMTrdjsP
6xrySL8400pYRrygS7w/T/SbL4un/6ZnCBttjSX9HjR+Fr+1smasbLgOcdjhQyvy
Qie38xhIOFd/tDTSP+GZloFirYqn2zkeazYvuRdZGT36I70ScycKW5CGvTKrcO57
r+RZyjF0cesVr/OHJLkCrKfpG8oRSY1H7g+NTGfZY3vdMFyMir8oT2BjUFi4PDrr
rCF6HcGHjMHGr2kx5hedMRTMDUGJwNRaKUO3yoUgr6NO0j4bkrv8fSg8vwvoPeBA
OCON52U9/R+rnrQlBqGEBLfPhP4QxfrmB+1il3bzRMfxeN5Nhl1q/L325TVrhUbi
fttM4O0pEsOOQsTHI95hLhxuzJx0zJMTQ+O8vIbGh0tNCOdD6yRsEaEw0Li3u11F
nlHpX1v3GiFicN8X1wlKZf9KWZFnUrib0sm19iwkDK6ZrZ8LN3UY7nruj0hDeuzl
l6cqQDriGijGsIQHyTtJtNUi5QINAZC3pGBSe545O8Th1d38BjKAFudSrhT1f94X
BcEsJYAtq8fl0qsw3kDeSejMMzfs+7Rzw58D6ZIARUvWOpzYwhKK1e2hnRZmPLwi
CUaVmPgwOxuPINvuucr71sLeQVfTMzHZ54A4poROfWHsoE3ZH3JpAC6ItJngm4Co
/3ZRcpTJR+8pLLE9TGnn+GjDOTNmh0tGrY2E/YkB8pW96BNq/AUPoQ6bPOOK3J0R
O6zrrNs14VQOwDm37Mm74sT/WV5KdR2yfLoD6AzVYfgg7K+6IEi2KBHUMam/zRLt
dbazZFNtm6pdljNKTEiM9TkxpT5LEu4Vtq6ObqngHDT3J7KlANZEl4lqLFkIsbWj
vAAiHngCPV45RLgOGHk1wjYs9rAYul98yVvbRnPcEXnrVkk4ppp2+33dm1QCmVRF
HlhATiUohvNocJdKaydi3wCi2BPRPeKgOSVBQ6oxTlY0QupF/oFllIsqz0rk1KG3
jEQQyOVnpwC6sjCjp8Dk+SIIoddtTs05+lWSuQfZam7rWX2OcUY9pFZh0mhiHpZ3
9i23o8Iirzf5d40fBx4m5KnH5fcXvEB0N3IgS7eiFjJbuBRCCmRQ1LRrSw5VgCWR
bliwEMsP0Ad1BX5sSPN58TGb5TjdI/0fzhYXtO6byLbUXHBL11o5QO8pzsmHDIqX
ubgPWFVDfq5Rqo1aZpfuAxPEtmraXzkGvnUn7TVJILgWiPAks2l7h+NsC9tXko5j
vTdEJqk8H8WDW390ezl5G10FV87wCt7ClhQ9OcGzLXG2XmmHS43d2TMfQ0yqTjso
ZtBN3yEp2DTGZPEKjDxaYevZbaGAHxtgkXOZUs+SYI/NwzMo6sEHXABOPIK6hVJP
UQtP4ROfEOyQxY/U+7z76o4woQwldbXY6ogfSixo+jmAjb1S/ODFhfSlpV5w2Sr0
KPonUcSOjYN1J6oVFcXBN3HMDlFJn6+/RUGqiBo/QHetdZPSliFFxARlCwky6TSB
duBjjiPx7/zsRF6DwS801Gcrme7L+8C8P4ldmxtZqwm5Ql2CEp0cPPPBpKaiw4j+
e823MldgFi2UHRhFJxEa5wqv42q7BlNlT6wUJznuCHLkXaiS7gLch65gLCyO9Tic
FxqiQNzfCoprTZp4VRWQsrfEiMiOdQWMKkxUPASiXs4jsKK+TW7ncfQkFIkeNuzW
BYvJxGpUsAmseXRgZny9sxNhtIzIe6XjDQAsP2ulqET1SKL01ACe/OjzTV2uP3M/
0Ha+RkrFiPS11g5TYNhVPC9lOdcRX51X6e8oCg1g4dSIoq5YGG9fbxfIEQszLXUG
pPqPnefHhq9fu49HIEL3c7CORo9kWa6roBYYF9miPfMxUoq6djd6cTcRSg9BdYsQ
JZPWbvQeQ2x8dUSsF/EojBkOVjAdYMxsFS1CJrrgSqHPY5d85MsCqnQXGKuwPQbT
dZofHz0zrY6rkEseux+FpN0FTDyQl+odvCQMS7GjyKDHUxqB9gljwLwBfl7AhgCP
sQi0XzIBd5V+sjw8MNDhkLJvNOGNikOWCdsYrrAc0EmlrkEIg/8MqTb++DU4utBe
Rs9ohSyg88QTe3gfBrAyv7oyp59VFhLtNFT1dDE7s8sotr3m05+B7E7+LwEnGV5q
C741g/Zz4SsDhpAZtKSaQozM8hSayzoc7onnpoHBHl0dIUZvIdec0S2KW8cnPbyB
7X9kWen53u/aebkyMMqQHBaxYx8vs2mr+zkG3mZQ7/nNps6bOmqNLuQ8iBAWg4fe
hUnLhvURqsKax7R1op55MWyXjaxWOubextrtRrJnEsqNobSVHOIFu/QKnLSEwZDj
ZRE307WL9scFsNiD8G01jn6PDDoK2cJizK04TDdcssqaAIIQqqcmqrkKo35SJBCK
O02x9gF0Uv9dcMQ+HS/vk6z2UmyVKs2gg/tj19vOPqalweytnj+FM9/RPMIBdhbv
ScrBnsobP4PgQ5OrzBbobmYdBocvaxWR6OsUpjvZHXGTzA4tDGPrUBboHhOEs0qt
c7zCVWVHj8r54N/rnrwyqb88z9HOBL4UQ4PRtK2lLBsosxmi0lJQm7RL/xs/MKez
9mih4NwwQdDI5L1i8Qk4/pcSSuZcGyfIYK1nfr05+xMVyNgCViXhTkOKpBjgdtVe
QX9OkkOszaeGnmZm6PRupNbG/JPEdqMlk+YB3i342pRhaMP7Q29hp+19i1HA3lc+
qfQMVyYIUhmi5UlboZYZN4iTBrCiQvE6p6b59qQy1zZg5mdfJkr8gcmguObqEHAI
kgZKDMnJ2rAg0DMaEAaEk3W/nfQBAmCM8rVGItbLyt6Kfv8MuH+Vx0xG0lQHurJV
BL1XOWNrLARHd9dOY3a+dTgkp2HDHd9TPCDE/L2goK0iDqvBOCtbs3iZchghiB/4
7UqTbdTC4Xz676NG2vZTfexgGyBplkNAAu8H0OXXqQrzaVO3ZMNAkHebecorKoih
EGiezpL48FFflTpNCyoc42yNdRpZUMlMdSp+YIAbO/90e5E4e+OW1VydSCNdnJAo
qVRqijh1pPQIWtJBNOKThl2i6TeduM1xzWsAkD2tt+lW052S7GRfA9x3FcFBOzSE
Apiwu9PPcyYFO6Wb6R+zNxJZMHoKomdNzy84z78dBvqDV1Fjkm2genJNV+1P5mDJ
6xy9kkH33N+YKIZ0v442l0b4mlyeqt5zu6gX7xEfHz2pqdGGzfFCspfTPaQGih2B
JV3jw53hzIRpdBhJZHzUJUFiilZULwdozRipaDgVutIzmRlWC9wuQyag3fwb7tBK
T7p3RG2nW2pE9HDnYNejHmH0xljf7wEL23J4lHny8CWR354o2dsjTQ3EZkjKy4H6
NOY/lGInXvxyqXhe2sxWlP9kVl42Mpu8ktlbYQXSRbt3V/cP9ez0yvX9eP/dMxep
g89qPk6wu7oSpEvxiPyLFBUI3vAPSUzpez84F1bgyhWwjvQRVZlo6j0znVP6ftgH
A9gxEI+GrcjbvjvtmobFe2j3fh4LcBhb53dMZkg0WgxocuTbvryxd9PIXDWo1n2b
F5xnG/OXItF+174Z7tFKDylBxf6LK1fTHj/LOISpBNYuciTRaY+Gg0S1Il1Z3KN0
bFy4ogR9GndqQgA+TfYN7ptFCInTAV6rKdO2ngb8/KMVdYgDcagUg02Q9CspcYtg
tyMouVAe1pdprZubKtw5oUpJizTIlcj8xnV92e/k3s0MtMTITZNDsLg0FIFN6+R9
oVFDec+XF/3Ih06/6/YggyZhnGvb/K57FfuGz1Z7IL4c/0RetqHCPIOUeXJDxeM/
0zkdg4OMX2PH27vO5cDpvoYYgBYuiON1Ki9NkOXw+TyE4seaQVMqjgzkqQ5TRB+c
8p2woYDPcigsPx8BuNNspY6NUs4YNVqdI4Foq13ZD82AlIl79MzuuElp43aqJCqr
wwiTGwpAPr/VEHy7O1hIvE9GbcYNKxj8YazQaE6dN2k5fdX+Jfxp2lcO/q+dlynj
CdXIqr5QPoWk1HTEU+zXpR9e4QZcDB9PQfCUKAg9MRCj71V88PqdbGUQ/peZLCPD
ZbvP6qnYsaJlxIkCWhEoNKfAHWHF+JIKFq//uvl0unSbkRhra12axBkx3YdnWin5
UAfnc7l2XY966Y+Cxf21HUOZPvQ78+UfrEybWRb9c+cjLKqFwWyyudDzhv9T+rNY
l6gEIYJ39y2Jyz/k2hwUwdeE4jTmeGxZHVcWQfYGBmVrFw7L3lSZH24qyiEq44Tk
kwopC4p81esAbDCHtVGYVIcbxlNDCFQdJkQHjSgmMy9ltKwLGsdN2abrBR/hKNzF
gx9Sf2fyqKYheoqhFSZ4bXYssExHFrZ0BoonUgevPgmx3ZhgT3govxj5KVDjMB1o
sH7B+33slWI6DL9UKmmcs1R0tDejITS/cQ8HvwqGp86lZLZ++gPotgCUCo+fHiPy
3PXrpjb1iTGB28OCwI65UCiukEE37qi3JrVOBNPdJkOsNHEabrp04vHr3+Kb4tsA
AFn3RvsQDgE41ir79w6LCTb2no+K7e95wR6PZLk0cDWGf2lxk780o0KonpX5FOHZ
pdD88sPeuxlwb+yhcSc2okTvY6InTHi1BwOx6Zln2+2nCFfSXSHRXMAQCkBsqEiT
IM2ko8E5Tg+8kiRz59BFLEpGHq7IComt5ImYSzS402td3PnSUkM13gCMLXPp5nA0
7OH4lqVfidZQQ14cuwA6o17F5dM/TMhiZBEWHc4hvfC5l+synSuAWOFqeZNzAjvS
f5/yy6QdYTH1St63f6VmpaAnk0VsPqA0TVq/nWhm8GmQ18LK492UVI4Q7KS48k69
kg5luLMgaaihm99R80edoK10qXLU9dn46/8qt6OwyyzYL1Kp53IcNBMPezHVweVQ
vG7gFf0D37Rd8PYrVYOx0TwN66U5V4HNxQZU5Xg53p0gj5YxTARtiEIEA2ckFNWM
TmvLMmwMS02wzB0BpUOAgJ13FAZOwU/M2NgJjkdS2plDa/Imd1v+aefMiMDenBWi
665dNbiEa53Eny4AJugDtQQj+VL+Gpr69FlRyY8kksj5/FSyb2mt+mgeEx1F9Z4G
P6LthlZlPuyDl/pqlrTBcyjHFzO6rkCm8m790jk2HLBqp3OGTVFvu9Bn1CK3DLrU
0jtrA5xEvhNBnTkd3mz3Ce+ZkdD9h4Gw62q5UraMK2ZVVzNiXmbpIYooa5h4BX78
oZhqHJm5gAfdFAYOh7i/lgg9rBPbM4o5ZmPbGEelUaDzTZDKXVfn7GDmffMfDUMJ
uxb1onx785cn2w057Whb5YzLkRMySHSsHc33kfYlz53tMM+unO6qvWfN9Ue6LfRA
XPwvNn2ywQLYemV22doAgz30/HCbFBvcWpBiwKBo74kmPvlkb8hDUFCN/8G4kszQ
XK34U1HuLTV+ypcz8hZVcrLGcu2toK7qx6gxtZFqK+ARGI3ZWGGK/kxCSG15ynVe
SiTGp74D+wro/zuPAA8Xk4P1ZnARQT7bCsM4rq8yazIRzkgiF+yUPoH736X94xRH
xpJ4pkd29sV5/nnArwJWqM9u/KGZ5tmq2aIKx3+Ob8LKfRVtBAF/wMr6A24EaJD6
Os5S8WoV9SdNhTl4lL2TkXBviMwuMACZCXhC04hS6KQi9V9VtgKfdCvobo56Y80J
tB3vgn7rgwcC4ul1MQNXO0PBDJKGDaFLP3JWNYsmlHSKz0Q2mNhOK3v3bOQZkgIj
Gen6ZPOgd4XSCLvWowrmyy/w5IploH2ZR9BYinBpNJ+BsYF8L5m4MqtvyKNbYYYu
zEmODc33JZaQ9VKvRgPhXiF00hTacN5jJDMJ0GYC4jqrz3/vTQccGLuoIa/8qYWK
JjtRole01gpP3sqaulrIfOXEstCsHpW6ybXB6kAC1gKmyQmpQUTuIUBFjGBx/H65
IMaiFJdQcePZ0ldGeb7sEeYar77Vdc9dfSXe6f0BvsVDOiMwWvXLUq2bvW3fVYZn
8w/p6ACvBYb7f/WWJzRNcREpjJ5ffvqouX+MpmiNUSJDdx5OVhgFKMIBvVaXFBlB
YikboKYsob0KtFCTO3SG6csqyfoSHzl1gXDtwfrkPe2x4Bw1M2ApiueEdA9ilh7t
kuCfHpzF8nrx9Y9SGNdmfdTvCmVO4T7w0WXP3o4FiosrjBU+NVseS1P5fggC1bZo
qLNT2njHH8tRezV+GYvh6fB4Q289RJtyjXhYS447gt0suVOdojL3ehC+XvasmPYm
NqgQmW4bNZmdYkpbtuF8T1tdN0gVj6Mccca7tUbyo0tFh2gobCpqKI6rVaS6nSpI
1b6tOufmpfKazSEBnB2yWJCgQ8ecJtHH58ZkRuDo/oTpdDDDZywGDWLxAK21CGwi
3Sy/PJvtK+Bt5mDznvgSdB8GZAygigw5eEFHb3mVHeSudLQMcyzzjQuqGcIceGBv
85xbFbMiU73J+arMmuazPQkudr6rlB8cqltv0Ckar1VJB8rXRVEyWrbPn871UVp7
9/G5jJKGZ5bX/8vjvasylxlcTXvbWDv6GQpS4jcJPEenW8UGKfOEPs8DcL2Ppg2e
9aR+It4/wiutPdOdqz0faZ/6RwgvxmNVTqP3yINoVTHjVNQjK5Dey9tzKof44jg/
D4FKnR1X0o7ssWfg+l2QwEJFgumL2YdhbkL0GM4S9t+IiDAmpaaJaV3MkyhTK8hg
4azYDgs9jrvo42lzD/q3SXCjmtoIg0tZGJxtP0r43rWcZpw+AJf/bav4RpfFI1CZ
0Rqh9dknPDRZqcxujuD1WAoabuExSDGWg4JDYmzclC5i7SaxhfcuujVLGM6cyYxW
+7LqLM8pFi+WlH4qC3AfRggu+S1Rs4k+hLwCX1pUYXTK86nBPPFSQuccZfwSIIJH
36gdM2goSBjBujMRxBSnDVNfd55E4Z/uJPrDJG2qDhxgQJ7MTD6akLgMvP23oTrl
iPxTE5CNClny4qbXW+W+QQ4Ujkig37/bGFKopGKXzMdr1tbtr5eMK/YnWBisu7E2
RrSHvRMNgSFKGpfGxoMH6hUsgSDez/VpGOT007fE18WEqON4Rx6Bn/BGpjHECm1R
bcVycmykzAuJ69LtYd41DTUppLc/4n1LBbh275kSSDiDxUtc+qLTer70fOrUWbvD
vztVDjWoPOHhyciYxkYH4rN13iE2WqsdswVdwywLQsg1xpRAYKARV4HTwZg8ygvv
FjNYVbqnt8D3y+b0o3eb8QI0FNuRqV7kQDgucaaL/1EmRrll3VFJbf2QklamzR7E
C1+wbviXlhqdXJ/NjGD0u7B94fE1XerxDNxBEreU9L26rV40TvYHJjfFdc4XHJCS
LKmeifNzBnjlwmUreuk9ZemQm+3XC9O5quheYoQ4riTKBqTjV4FFQpf2KtZtvFAE
0EzZTEstV4yQlbVe6E0reuO7wb2ftR59j1W6OhWmjnMxQgI23A9tGPJUViSgDD83
mj0OLhAd/pmtz2C/sC5wTqGDFaMo+yUv944+M12MNZoP+v+fKthU68CFo29Z0pld
ej1FHiW9eeRcMdhytjp0+R4Y3yCskv/cc4BFSjmDNDNOjvKcn6HVgj0zUNulFxuN
8KTa3K+J3atEEsFdWLzDZoIBnyLDjpEsifq+eHkZdm7XO5VATbv/jZeNYkvF4w2S
1pKJyUdys7vFbMZDPqiIwGA3NyikzicS/fXNrPYy7AWpTeQZlQoF+C5gJRG8fyn/
3L8PGFjVpXPAYwsp1vRRgUB6kVfwxSLHbsxmwahMULcJdPkWuH9tzohqcYeTXWLk
Ious24gbbFl09X3X4ju0maecsGwOPy/wfYEuKmcrhM3AltldjiT8yNC78QGYwFyU
tu06fvlB3BIQgfpMMJfJRqiI+3y8VaDv7a64+w47eNWD21UIzA0sQRpqwPdumzA7
aneTeseZStQTy1m8l0uN+Jo8jdiPuogvB/mrNXLHXgV0HEgftTuhLjl4tKQmhfNK
CrxGEgYbalWq+bHerbQal+aMgHstvsJ/AF48BsnnXTdPfzY/CY1t6igkERsyhmNR
/cuuiXXpWBMjdfn9nT79Q4SA0LMlpXyy+w/4BfkYhThg/3N8byTwHmrJJiFCEM3Q
o0PFA1RU8N+OjxA7JMcjtyvKj984/QHa6wdH++HcbxWKcD3TOi+L/r+2gyScKaTX
GffjsW6pVJyFlOLxcIOJyI4qn2RwgLfiRDhahTqLCs4OFwe+Q1DDQvZ65Jqrp7f4
WjdZs+oA6yBKcpAjUazHhPrFEFq2nLw26nTgzfkbkMDiolGOFxbzxR05A1JNI2i2
DXORE1z82X7TkIuppT8bKMOU+Hy7Bz165pzSo+IBD3zN+ew8YTuPyiWewrAZolum
4u7cHMT7ERYJEsxDot8uRIETKIiJZ1mfkSUnR8y/8vXWPJJ1+9pmMnwPn4LLJC99
J2YkWB8M+0TEsGgqVNwlZR9+dYIucp7Wkpzu/ZlvZLue39Fy8gISSjZxSCNOFQHD
u/R9e4aNqxEAfOtrP1y/5crj46WE1rKCir27+yAQFPtHFO5Kcr7EaW6sSx9N5GSA
FSw77q17GoNHHfz7ytmbX7OBX3Jk8QanrWED4dwtXwej/u64U0DptMN69oL2hcdw
8o/fJn6P7s9XxEpfxY8NftR1rzbOahAchdEc+t8InvvZMswPNlf40qBirWA1yic2
UO6qHrwqzLklh1N5F2oAqZR3SaSeNuG4F/anEO3daCNeQNBhH91C4xOVtugc2dIr
jyK4ksAzePyME4VKm/0j51pKC7CaWXU7ZLve6J7DMgCku/odtdpw/J6SlmB+EM2D
fcjJ+glFW2xM0qMyB2BhYSMrEMunvv/jgoKOnrfyfHsQ8EPjEhibovJSqs5cInns
HCybJM7vyDJSP1S/rHQ3mqD/xNxcEApeIEamaIgPdK1zloHVWVRdeztKoAISLjM6
GEjIyY2GbNdkoJY+NfoLRnBB3VTe2xzQQEqsC0OkPWErJN96nYgC2UMBKG/g9mSu
RDnvd73kHDZHv+tUTUrVLESDLbeRr5vS99yf6O9ZKloCBUl6PNFbXlwzZfZe8sI9
ly/eSS3+qMEIl7Pf4fQTvN0N4ILvQhnW6DeBi30/z5W+zBkfniZlDnOMWgwSGs3T
ZOsOrkLdD/fazgK2OMf20aOg5v26bjmqxNM1R8XbLjlWCa6xrRLOoGqg4AYotVmw
ZsBbeAEjUs9Pg8EyIjMEXczYNc8Bwl9deZFYic4fpztMCIwwYBOEBs3lvTwaNqHT
ZLOXNwiZ8+/0tk6SAFY3PZebm17oFXBdMa0iGka0Ay0eunxN9LB5djxhxuvoAvSY
df4nAS/B9dQwNn/+0nbPPsnBlaAJv1rnPntyJhUyEboUHpi3dd00OHWKsUlyCGCn
zXGaEssX3tJMqEBtval5/GYRrtOr+iIpTDl2/+r1VKIE5NYFdWasVYUU9gFkJJQj
enB7Amaa7eQenFV9x0WStE8Ia1OucIiWYxQWTjWpojyBF7pQ3h7iMbbOPI9jGkTR
N2jNdloGuYeSLAQyg6gJktcREA1gRXTYU31CBtKRLhL77LKlghHw6qt0DIPhlHYJ
WDPu59YQpMjAS/Bic7jSMAQmzfEZBWiuw6Ig8cONNKTCHCxBLd8NqP+5W2zBDLFr
PqQ0GsyQaIB/cCIdWuiHtaQmPJnWuCFjoBg+ttlMyRqxXUcwjjpmpy6Co5gejr2V
1Xv9WoK7YO4a3D+aAh3H8oU59WGRS/iT9PgTiEO79xn0Cs0kW/xtfQqhMMsfGsYV
fSTiuJBAxwk149U6qw6ZeVgWIkv6bWYl7UrCZbkrj8eqRH6YCTiMPwGgLs3brIdK
cFxVRevN42dYa7SKNZto2C+Mq2B6S/d04XDq4nLWqkf5GFCSVnPg73DGfQDNjbfv
P9UBt4KuF7OdS8cyL1POpHsvhNJO8LU7zELi5jbvi9Zftavag/53610JeudkLNka
Mni8TT8DepUhV46ZWiELa9HiKSOCNmh6de3Hz6B1INEk2GF66sgOMK+VHz2rflgZ
FucN82A9RtbJqNOHUBKIzQMzq5PpGj/VcfGE1+PHoSQKy9yRyATNQmPcWUiXNMoP
8DD2C3GV/8Etbur4rlmYEA2XhrmyOO+s3Cgoxbet9bIH833LOYLOI4zNhiYfUo4N
aC5YUiPT8RougHIaAzJkzXCCtehmxmrr0sNIrEfI6Kvf/LSjL4XVhHuSliXIJxiA
5U1FOnyrz03mMFJfa+EXRXrjljYqtbby0bkMXpojCUihD0t0+qS0aA0yqkzqy6W/
iWfcAVTCb52/N46oMl+kKwtfHBx4x/V0acKr6COpr+F+HZbfk1OpODdxOG9wrbhp
ZmmImzQ+/9Grzdt7nF+NmNPLqBfrdf1x/3IPCb2epq4z7i4CsUO1d/lzqOc5KRvW
ZpQj5weNwYkyzHBw4QjSbAx9Lm+pLooZj0/xCJurkvSbttQFA40rh/A2Gov1BZWq
VERqaHvpQGrloAVzLTQpBebLh7K/z1Ns6i/kWp+hRzt4mKxUFAOI+h+1HRGm3mHF
coVYqiylrNmeHsdD0LNOv2JuoOOsdmZBzuJfmw/i4Eit/i62SIRObWo9LT7PZRr9
pXPiw1pRyMDiXvydtO7Swdf7JT1KxP1qtutSayuaVPdsSZoRZ4AnKda663ZcKqDI
xjDL46cbDGaPGOoJ+VS7OH0Dqc0hNpcJuHarZ06l8kwcTnTi3/Z05SiywD7hwCnJ
d5/G+4JiXtOYDQrG9mm7d4ZJ/fy8iWXLqSQVadvsMOrCX/4txcVl5W/nl93UvCFr
ztW4z5XiK0XLf95oR2TuRynC/kR6Md8We9EgC1dhY/rHWEeNBxWtYeMjvxCFJCoe
5DmZcHIWhkevSElf7TsgBlMCG9uBjZSA9YWee5Pjbeq/bzv7jY3yL5O0pn4KOF7D
NDMpL4oxElMyBwf+rOzaaR1mEdBE/JLu81vw7HEJJXyBU3y5V8fgqJzK/q75KJ1t
fMse9o8/r1T0VmGsxM14jWww3j0FVkljDcKxguOHHvuHrZQ6khGaJ+1AtHmj8tzV
p4ApNsL22/drk5o3sTn2aI1wk8n4Yxg1H0P7W6kMHYO0DTKqxYCn/HLL92NCfF16
hP+x5YTN64CRd48fcIbVzTTxHVxZou/S/2zjk+ZrIwFqIRiKenvTWy7wQPnsnecS
Q9HdrhMRuYqBQtih+hFuLcXdX3C2VFP5hqUO2aUBWDMSjf76SYyd7YTZYcb8dyWl
rKKnL2acqDfrBb32v1tIPlHUjtO+qqv9atfMuxUHVf9slog5rMKSAkTJsSvXCPed
QA0IGthH4FGg2+026q2epa9quBTGG2mfVTqvpnI/KKd+iIqY5zlVmgSwZcqqGVce
zZbHMwpFQGrzIQbc4JtSMgtsURnf/4Dcy7sFvIY/t0zYrK0XX/rZoPaz+azulD3I
xTQeLu8+RxE1pA0gsWcPDsiPiViH32uZcMV8GjcpITSx/RE9rZfUuIgjBbDdkVYf
1HEZLWeeMZ0xoyEzUSuZfTUUK6thvSdOkOfVgzbfp38WrWmVNVSaS0qNIml1PR6i
ZhzUxUM3557mppOHwQjnUO7u98tPcu7k7muQh+LjTWsMfRnu4X66tKTi1NQj19Fg
FSvpv36AVUltNId2TENS3llYUnCHlV0Ty1W9ykUI+EPH9UFy1buImcnGimUjNF6C
GnLPx5trbz3eT6b13YV3vi7uzQUOND3XmP6SkZUET7rOnux2kjVZfPepzJxB3wbM
zDYgTOG2Vt+fRPcW2oQVifn8vwuFja5muMOURayrppysu+sJmcY8I/B0Aj0apJIa
Pn6xTIipQuIfJMhzxus0atTU/mHFgX4KtKSkvIR+StrM2Y22wpjvsjjMjVnYUl15
LM45SKg6liruv2zanQdXKf1BVY9sPSq9uX9v1ntjpUFg5kNOmJ96BZJJ1Lxg+z2J
b9MUHgN43AyC51r1KxsBWk4Oo2mKfRiUobpf/kcuqx8MmOCH6UiWZnFkUVRvGcYH
6rJisjds+E6MAgVCPQYHW3ZIY9UTouU5A+Pla6pKjlIYwcOSSeNgSup+Tw6abIMb
3AgLK6rjEdxO+uwmv9un7ibwHHHWrfRab9qWvn5e7YR7XMoE11Clcssgc1j5uRpr
RBf32/zVZ9qYvOms5N4kMXcoDX3YrjNqWvFPb8ktZSLhbf1UZBuEckbEKkjNBKAg
bOMwKcVGfJ0PyGMOyTFh5RMsajIS8v7MP3VqjYbwLTHT7qvUPuQ56dPSQf07/d2v
d+H28vkPeKfn9aAR58GscsH99vSPwtGG7vInpEQvberc8i2e+Wa9VN/DNF1hmAY2
N0bYTPwV+smRUbeiNrVpcOd0Vew1HKk9JdXv+DG1hc8uthHO1VknoxbPEtvKnqdE
uyWFot+MXv+UHNWoIyOg2HmHk4j4zJeqOhV6/2WreXQwtH8kqmnyI9UxLKlvp8JP
V6Mo/dfOork8UceT3KOF2uSfC1ZS73QTj9yBv4//S3GoF61/XcZ9QYlFr7q6OTn8
PazjfMg+iX3s0BoenkoGsVgW8+xo8m8qqQZSYvU7eDgNt8jmM/K61U5MPFOhgjzd
5LLgDC0MyR+nMp9EFb6CtsqiF/8bTM1s15DO7C6zEX78ci5qKlW9c3R0wFoz0Zc1
PQTLxwmCoUEVW1NVGDf88OC0zWuOPN67W1gLB5+fdBvoU+laj2BsYFe3wNvXJ4mH
eCiVekMUp6YHYYTLyW1B5Zi4vGKZeTPIjBzSt0lf1wKJu5b11uJd8bvQKLKqhkuX
PjBrEZthgZXfvk8y+e56I33HOmkm0vZJd5EK3gdF/3scBX8NHXl34nBWJKrGk5kA
FmxE2ths9rkkCAGa8PuGva+0bXetPOKKolEwpDzH2Pcfz3Jsbkfno2drXThJWrIk
02bRcaen7UHrEf0go3pKKMIXhVQCWDWGhM2hgmqs23qwJ6tIbHhlCUtTG0DOyyNz
Gi56FtpSjE8UCp7Xxehv6sAmZn7crXDZ4POnwixZMF4jUcZYppuo4I93EPq0WB/q
PP4wNnIZcX6c8exUtxqqpJ4CAsFJ/b+nwUrBBYfEyi9twUaKKxY9YqLFae+aWyQj
nHvlOA/8HS1NrWqYc8NVU2cflm3ExXVujRb+fTtQ6r03tb2ouZNXm/a2jLMfmLUk
oQQhStMtinFUKCzLglk/GIP2GMqx7ejs2jyBI8TXCd+8daMmSB7FbSgWEtCOBDlM
QSI8Nzje/4PpuRTYrf2F4VfLt79g7kutlBSR7zRZNC93azrNtRwL4ROz5VMFsmjI
IJCnTLCHT+53oXZn6oD8JA==
`protect END_PROTECTED
