`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3MD6Fxs8hqN5O1EmSHzPNMNVs+gCJ069Kp7U42G91fwKxSEEZu+CH94aLD+aR/Is
WVfdin5y45HwzodyLKQ/k6NXQtYYI59aTV/QW9rDid43WtwXKRo4VSNkd0K9xsJC
rLn57fUvr/FR41zpOg/h5z6ZkT3e2E2oUJjSZuTWfIcGGGDamwOpTsezKREzrkF1
d28rPE8Ds7dyxWf0VXMC2d0KGMN+50zqc2JXysauecw38K8eYHFGzmwLacxCBR05
8Xa83KE0cHue7AajdqraW3w1MGPAhTrPOB+UdBoc1O6pGIntQiCoTGM5B0xiEoxk
vadsNF5wvNYyR95WJr5z+3i0/pg3lDTTI7ps7m+pXtPXDDyznKHKBDyutosoNv+z
BRaOGZgs3cqejJHkkOk8CL+INMqB/gYw4gN85yCeDGWGD61So80gkGz0Lly8OJJS
C/k+ipZLb9ZX4U3hWU4+hwH+vlpFG4jXMyWD6mGLzIpkWn+X5WtZ6qWcoQpzw5st
lcWhX6mANoVC5KNWpXvlZ7VSHdEuAHQMg2uaDxvfbqRE23Yv2xMbpWMwK2QDjEaz
guQheAGHGH0yHhXVG7ougqCnHz4+CWTEH7FQiNv79/NSjzYGKyz3pAd57VcKcEpU
pUO9AvvD4ApFrhUznOEP78ecsy/DJyHRHZxgvTsjZX85SXet5abVtwBYYAg2NQLd
+oS3lmJosFvwVUSTyDJX9P5ZcxwLeCSF+Uk2s3eZE9ie+CxNDc1cgRr6nPz6bmkR
CyDg5X+9C4Vtd/kP3yL+ATH8tOKQKGSV9T7W821N5EvWAPtFViB0dGNF406k1os9
9k0FEZygsvjArxckJYe2CTF/zZWARV2XHuj2RFKyewdlmILmUWa52N75rBUhr9dP
RfohB0nLcijXVxeaMOy3Wz6Y35uoinLsJMz4JKDdUTdCKKl2NamQFoyZMCow8Q0b
DmDBFguXo9jbMHO4r9H6sZMJVaCn95IJnywwkTeidmqpV0ahNqpfLbC4pZ0+RgxG
k2L0kAN5JsVYm2Y1cGidD3mmq9vaW9oHZSHp9hqGG0QAKNvora37sfoAvcCYn6DB
dVsEA9bShNDFxS+DWQDa3rEyYZxPooGQVqpqO9VEF8XA02uOCEJfVUTWZ4LWeXy2
0bj5oeY6w0Yz50CU6dfxJseAAGc1KdXpUlLpq0CVTBcGMreQz5+caCeA9sdDJxjB
/z8vUyhzrlxlcl7T7QS1ddBJj3bXuZDNK0har7PwINHe7GYXdAj3XSOwyh8zsEUK
oOrQMiL8xYkWTy5oFFptZ0XmQjdBG/7lRzXP/ZyvtDOBEpi4sLjyQp/0iwGMEp7u
14oikl3rNM8A8zqqTkZtFZf3d6VAy/Shm/ndtRZspclvLnpOnqHeJt1NC8T/3JrT
T3OKXwo57lTCSJn/yDdYRpzbZiKSuk2zBI3A3Q02r0UaAq4W0h5GLUi+/ZuX6O5l
xZYoT8I5uBadqmCbqC80WqYYWstcNGk/flC06Qp3nj0/aQbjxgh9zAg9xrglvCIQ
Q+HrYzxtEBfiEAQFQSq9vOXV7Tvr0F5oYQJu1BsEJvyIAX+fTKtccPFfbv0iq/86
8SxvM+znBCLVdjHcri19tkMUNE7ZOqF5OYd+JmU5xa3BcnspWrSK1odCjXBw4hjv
N3A3KG+Ltol8Fw9qJJz5qOLA9On9G8jToMIo287PdSRxu2h6zkODDhjy5E6Gw1N+
kA0NZfykG222gwl0M6pfTm58mjM5pE87SU0A8+V/O/pbEOsN5lLtdzqvfky+pA47
xe4TBLANIMHuijaq3rc3qfrlR+mpA2TnYCt0R2JKw0I6p7A1RsY0FKdjHLVgpu2d
eLGZVnf3h41s2I3MGE3Ma22sL1wkNXOZppc8kOoX/7hoFFGamVey2AuqGK7zEM+T
du8jfFmKH37tdYtSPpzD9sX3P4y5gzoTQGo+onEXFkiJUTfnWFS3qYdAIjREFSfR
WD7lLzMvj6Q0TthNIMBn23xrsaAZWOfWBEey+SoBJQJQd7stcsODnbHEZt5hqDv1
f89aeFpgUxQ5A9QOL6MMW55OBlhkmwT1P+6NVQOo4NFF+6i/OweG5hhW6w0UAIGH
W/cj3Ptk/eTGiLCOgCeQixnc+ZS6W2q6zNsa6mCyczueBUiwW+ZzQZO06+itAI/d
`protect END_PROTECTED
