`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
D+m8IbbwgMYAH0MYz6CfdU3fPUTj82mBxGT70IdnUIu8mcu5+HLWRq1SCIYQUKsg
zTVmhnmjR9gqMAThYtFPzfCUGNGPOXiXqPZekeLtfn3AcrMwAfkbsQ/diXHccRoH
XfZ095A2CKekxkhTQHvmVvueGHSSdBN+6DqYXseDVeklYIK8CLqbH/1/iWSq1tmN
9q5ptJo4NE288lDmIMjMVwqswZqkVFjJIZbPZJ4VDGW340Y5nX7jr3K+fPMgva1A
ZZy61vZGcrJKMISkb5Z9nRf5pLDHvNoxilXhEcaGR9T3rNZfMr+DLhB/9WA52IiO
zDWpiYkDvxCnoTTMDJ0btzYgoI6vfKyOQkku12uJdPV/9E8R6dNAVSzM9dQUl6vo
1PBcG+bCgm7S10F62vgJ3CGyFrlml2y5x57iZ/qbalxwV43v3aqQWm0likZJRIgR
oSUv0+KJaN8baty9R9tmGwgc60cwqd+UbncOyhZz/pV+BPABc51mSwJAtq0y5sCJ
p+8hCt3iYlBVGh0gPRz7/WAD6IFf0vR+Cx9csrHoBZm9hI8u/2VXQpgZ6dpjQ4Mw
XbrNfXaK0t1yr4GUHJcXXBipQdS1tBBg1TgUfQu0F7H42cBjrVVZYrMhE66Bn3yt
ETlhNVG6FDf7C46x4kwGXGe1t86DdPG6h2SDbEGReSQuTP1NwtxLKF2pzvEmxziN
ymyg5sTOMHVANJfybzgHGuHEquZYqMmNDzYb1RhT6O54h8f3JimAFTAQmpaa6nrS
HnXc9B3xXAn4EvJQLQcrfgwMpBjhRSWvRXprZgmR0uXq0VJpf6eATQypzK770IeY
2k6v5wpVxWCDJDHphnLAkb0KxCuJ6G01/64VS3Ti1+THyAtW91w+URRtjq6mCGKv
tTvtxvqzFQv9X3g/5XRFJ84UAA61xrFMaZejgnrcQt27ox+7J+Roe8fggWLCxN8A
CXfvj6o1S3aOIJihux0un6Y5NZFhbsZOyhfur1TuZAb7dO+W9jSp6HqEKpUOQw9+
nW83BbNB3Cw7swHSLcKkKQjctG8cIFq/s7a+Cwpe6pWOpB/x2kwTlw9YRbGX2R2B
2dLWDLlI26mvZm717oS+KinQH8kY/TDPhooNU/SXhbtm0gQPOqZWyoEwPakRwZTP
yNOYAPKupA4jKpbOM+kXLOXccKdoaN9tEOC7HvrzvA/f1kXtzke6eSWEpQMaEsk4
bYjg7MvIvnVwFp63hNpoWsj0c1QCiwskWTeQshdQ6pG/EpxsAUplUFmHXK3TDOvA
MIokLo9url+xfqHXJ68fez1VLEgCKmzIJ//kHYeyP39DN+kCkl1JKO/KLeOJDrLs
nzbwd6emTLIkqs9ALaPPbm5VYkG24SAqhiT4lu7srUMKj6/fbl8eriu9mgcHjuhk
5ypH6ApFutHHnmeAj4vq+8smANaxLaJKeU26qEt3fzqb+R5td7du8I1Dv/dCKJrV
gIzgGD64dtUcCYzKdTZ0wQF9Ycw+aTkQJUmBVCAXjwwZULJ2XB0F+jrcZg3nRmDb
sZdkldu3DLj5TTsRwxFTpjOM8rCiVUopMVrJv39S6HfLDvCFeqrkbMvW/whBgJve
5mAZ6pGN1h0i4uZl4KuJkjMsA7DyyeQyXaFrrc9L54i0DAS+XFuMmZ4hD52cqdtB
CtaqsIoybRPAoHs1cNVciaQXp6v1fXp/9SgsnGnokeQ5fS3+QRRBEAC354Lylykh
f1qDHpqyZGTFK3OhMKvSvKizRg6WEgjSKo1eI6m59SWTYC0GMPkXKTVMHi1OSh1j
yMmrEVG6VRl047uC6hItiEKwVmb635kr0/hV4WlfEZBzefX9sq9JFJyoV2dQvC8Z
/XE1Zg8b6r5ya3a6Kp1QZjAciwLhBHi51OIddM8bWgozTmGCIeEYTDBj3MufYwGm
cLf0Esq22JnWnAfHECmA+0BTUGQlBehx9m/Ht9zvKlH9shBMVo7PpjjlUB/cCrgk
NIKuN3AtlsDCYyICHzYkx9Z6MmHfGfSupOHU87DLTgnKgFfUseBtz/XVn+IMmaEu
o/c6Jisnsg9BmWPvDyzhPfE321qu48UOdnKRCZpAn9Z60/1yTDIkqOrEpGV/X91T
sa+nwX/M/KnoyyN3WgxY88hZp7jCEEJS4SwSgaG3/7IJpx92yZ8eVWGShjbWWt/Q
fic69sVpYlX1nvowlOns593sUmUJa8LOFXcVSlWLh9ZOmD06lmUGMJO1e88ESF31
qqqMMODekjs8N4w4AGF60DLyYndPymtrUGHesDxiTJtfbmXbDcGzh5hSGi349aum
O9ye/HxXNgwcR4tJpYMMU/XPTRLG8dgX9BPJiiEs7sy/MIRD3PPbeCOYMMR1Z8aU
Dxm9qGB6Me4/PQb5OYcQLGSe0Qvw2QAEGNpvNEUy2pm/gZzCmngN23cE560/dIAC
CCS1FxabpgcCOB8Zn+P63nzbsGbMPbBZTWMgn+5G9ps=
`protect END_PROTECTED
