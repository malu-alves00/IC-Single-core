`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VnlpryJzuDuM0J/9iTtxkB9Bl6qzLqWWCr48fWf1lCkH2865yXHHqahtw5L+mDSr
14nSZ6c0aqPdXDSSCBXXPxzWYoPtLBDPTkMpjKrkx0Lg1uTYNMwkhxD0PaBarcYV
OwW1XHAhnUS86RHmpTDiURokQy6ZOevwe+jiQ3gZR/GfIwN+v/9s1nKsLpYRHK9a
YFN79FKEPRtOGsgfroM8bwClANyuRmSr0WOTXQT7sqwL8yvfuVUQBFqhD8Xr1XvT
2QqYc/8FGXY55c8TWaL3szWtuV9/1cHZBtIDHk09E4KqN8aDQawxe3pzX1V8rsEd
Y2YDTNfpQa5MJ3lze6AtlTaxIk1PjGrXbhohitTAE9evu0CZ0rpVuNB2lTQWif4g
JvmF3h9zOvq8uQIZSGcR0dWbvP9pgxvoYEj6xSpF4xQ6xynR1j4DMGGF1WCW4qTb
18pvLLanrvfBERE2OpJbNZUpzE6qADY4vcaaKMy9X7RsznJQMyy/0dZ4/xYMaPyW
HcZ/O1Xp/GMAWXNFoS2cu2Jort5Z+JkCG5CTp7+oLOxF0XCbqLVP5I1bylV2FIsZ
`protect END_PROTECTED
