`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nbpCrF1UzDYs8OPZ0d3ifgZZfVbQ40OQ60om2esGwdeaQl+o4MLTu//ZuOUt0xHa
5zCfNtGQTW/i+6p2FFuwgN4dcALziIy4FiPe8U/0MhIkUKmb4iZgFF1fgmPTx9Ko
wJCoJMOi7twtqsN7DIo/CqRa0+3SNNRc1fWbZ7WqRUkyxyIucREpbCtqkm0S8NMD
SPWKsfe4QVgh4sPyN5nHHvxq+mZQwdmApJnDDeWwTPiP+E3tRFTYRTbIJCpbbx7s
ykWSNP2EtAHVtRG7pu0uNshXWB9W/WZv8/KcgdJP6Y07I2jXFvbULaExhnJlR+Dx
6DuLHIbOKPZT5nM/3xEeebq76JMfzV+GfhW5ZDTAQ2yVfMIYCtla38SKFXHhfZa3
9joa7nmNExSdgmLVrzkyiFIpLK648vyFoPPi+r2vQrl5hmyGFS5C9N72X+pk+PBP
jLzVGn/xlxX9SwcsaFgS98xav1bdnxURBA2cs5jN1/u8yE/Mt0DI3uN67KIxUc/C
EKzj4ge6Me1TymANP4dIPIb03XwERSS0Sx4Z3yvuK9sSxkzE7ToLF3McAPCxhdyl
7tA1k+C1Ju91qXvISINWqgcUL47D0Ei9X8c4HKgwch5TwOOgWK8Px1ObuRuJdxbN
UYDVEW7FAamZpcfhxpKkJZYzvjW5jsDTS+X6C4vNtKg/K/i3/vmqjGBfyqTonWNb
o5TQjy17DxfS0pWluxOiSG7pEuJMA9UovExgC5Nh9Q32dSelYwH9D7BgQySMLjp8
53MneryGKTGUzwuZ3FCAWAzpWAETJ3w6ORq9uhioPBiDvVEkosf4MBDLaA3JC/iP
WAwaTq/++S2C11bsy6q8SOCCxuK9eoYNW6PXN+uFMW8Ai4tuRbXWxBh/lVNyttf2
cUFZ747L1l/7vLa27aqfEEjR/zBwX5eRTqCBfKM291R2lRU0SM5fjs0H/+ReSJCq
W3Z8LZOQ6asSyO3EisQBHqPhCm0kTKjQ2vLvShzarJdvXCR9IFXa4jde2P/MD9MU
Fc8fJ6EUU43UK+BvL4egsEyKSmMcyP7UfqeZMu17Osdejs3G9WlPqx68Ic/dhn7J
EtpF99B2PCVGDHW3VWrGm+XJ52AYfbHIKU1jasu21SkYgy6Oee6aAQFV/Taf5Znv
cP5/gxBDccfPcYKZ03FfLtUkEJ1qQ9utrIbopgpVZv2ekpgE3Zw6vyyY2i50GiR0
Vu4KpmO9xQ9T29jzORiigjs7Lq5hvGhFaOXSnQWkcRmSk9cTJV/DsEClc7MYvG0S
OGCZVL3qbFk4NU9+E6n5l6KgHtXGyZusAIPEdJk+JJn1Zb8oe+hdX6d4SJdAqwCz
M9zNT3/sr8hUbHdfJ/JV4u57iQJsLzj82op9MtedfwN06JtmnPShoPqTZLa5zqXs
gHN0yUVMBxnDZT/3kcdW/BFXeWzzc+6g4LmX1S91gWc=
`protect END_PROTECTED
