`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XWUfsF6TIraDVWZ+z73ZF36WbzrnOnV1RAml9z5RzofAiFzHlM4fiPykVWlZ+qnI
ba8u202lNumz7oUyoLiJyFFZIPsJywly1JfHaPIESdSPJk6dvro7UsqahGnmKshn
D3S3Ilyrh3znVHXyIEpMOYaYcM7yNlcY2yO5sfGLu/++1Gh/7Fjkw3OplpSXKOPY
i1OGl4PXXhbOZ4HaaafNCWt7ZDYFHRppLzu125a558YpjFMgAeXc+nBOIREsyUIu
5p4iNON6OJgsbWxEKogQIGYLltC3yFYPTcZOMoVNEmqnSeoTU1fNYXUdyRi6jax9
ILQySOv7tE+l/kFTli4mIwRYiHHokJoF6mrie+ySaINLEnOYz5ALGr5pWvMuMtfP
V+sTc8Pg7FmfS8/fllJc5xgod4rZiiA9PyMaWcXZ6JxtN9YNhV5VDz+v9EYbDTHP
zsBTM96yjmMISuHQsYrNI+eUzEyC+9lpOVVBiFRwaAE=
`protect END_PROTECTED
