`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Rn8EaOE99sH96yf3dbzKovAdRkd6NbH+0xuduJH7VtRLmfRWgBWWoxBua7LDKkd5
e5kMwhfImI36/Q1sp+yV5+RPY2W5qu1xzZ3HPQOnyBewByu77JpWQAbMuCm9w5Dx
wX9LTiSlTmaMR5WRK+5XdKndV105Y30LYe3iNVRHzJvMiLzkc2SrYpKacGEACBAj
ugVO+hRJoYp0EoNADwK0VqvMenC9OuyISqo0B8kGJXfqhFibiEYVlykHIAHFRswE
zZ7PCEwKBvu9OxmeDOwUCPHBVUKAKjaOgCSrSd01TEJV7Zw2sWmheLAkLDIwfCvf
jrydcwKmr7ADUdcW0B+BkkhZQBv1AhB8/GHUsLyFz1jAItbj1q7zylVw0Szjb9rU
wzm/XwNXXUsYFLfah4+qm5PcAdAR13V68jAN9Wc8HmaENYp0OsCoOnFw+8lGXCjo
2z+W7ow+W9yv8Mkrcnficy0rsnlaJbWmXuCfZs/GYVH2CGD/zn9CoSbhDXYJcGze
QkKoWZQRtxlvak+J/qN/4d0SVJTYLrbEg/AIT6CNpps+hrty0jQW0F57jDxSOR18
fCccMMApVZn8yjuevviI+vemyJSOWu973t4E7RcT3qDmCsM5gfOjfeVmRVIHJg5j
YbwfsymiExlU5rMkmsYwxGHHxNC1P2ij0ZAoAGFmJU38OXAkENs/TbBBQ85017iA
bNs8Rqup1spxLAj74sk9ZxlCFi2DVFe1kWGBaEjE7qtxFJn/VES8q1fB/duqxEzC
4I7UgfKCBYu5b0TCh7aa7PGZRql8vwPEPpM/p7HAPRtjd/EOJsU6JmImZv9ihrOE
0PUelsS64gJ+6PItmSpofKWyus1dGbxYO+hns9xUPM39A4EFCqqhTxQ+kjqXZ7BG
8t3LTQw5VgOZ4atq8z54qjCOXX7UPCtA4rd5Sy+GOlxw8po6WNAOVfTg21bzwhiQ
EcYNohHLvBTPD6wfYUE/oHVPkmhsYaWdOtYYGTWEYT9dcaLWI1a3LFZfheG+UcFf
rCE7d69XAIrrntMEq3xX+u0EN/h9AU3+LSP0C98om7D7cz+X3tDghKH66Lbrpw7V
xQN3U+vNoMEvM+LF2OLQwQ==
`protect END_PROTECTED
