`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
j2bSttA3pvngkijoLtdqseiYNeLLhQJd6MsthES73haYT+LPSaJfVKIER+1FsZnT
Zr+jJziO78UDn5X5vKkMUoNVpXVwvyM3WLZ2Unhx7TEdSdjBGi5CW8qEQF53lhFd
PfVr7+O84TJlZVHx67UZQa59yvITyceAt6TogSKVPHXkqgxLAs/QLOFRNqHLtO59
wZm2LpDfP1M8Aj26TtOd9jJftJ4Sdd0IdGPbOHkoDCkvZyqjdS2oNtxoXUIJkuQZ
mGCTeRTAW+ORbN+81n9ZrYBbgr5aGWRL3PelW2UpfIK0eJS2p5oDVaZ/Wq1mnQ+j
S1f9UKHA6EmFc2elG30Dpiung0s98wEFHshi2DreSTuLJfQp8K7klNM0xG14Mb/J
vsHfkL91NEFhticMzWZgi9oTJ5JPF8gYmjKoyfv1a6EpwueYcZs7YAPQ3gu5meIG
+mVBQwIyK9ObDZznMQVz5xMqrVNolR+zXECJi7NuC3DatXxdh3XlAY8suEYH4ZKG
FmdYM0pmf7pA0bysuR8VWi+LDQgAGAtd3i14UE9c+tMfgjHPnReajyk+0q3D8c0r
MaXrbhtUefoMZnXDOOACOHUPvdrbaf+s2PSQ5cD1EWPsbz8qBKbkOk0qEkcLa4Mp
s5YMaFbYsEd39rkc7zolK34alcH8MWowIa+Qm8ueT6UE1gGFaS/7+q6C1/Wz36QR
LkVSAalBhA6uDsa3rpN4XahRmM32psEPSyOrIG23so/Lec+Th9o902M5Zc3EsFba
bPIVmFMULjU7+kHf5pcI7NCSjlVnpBqQek4TPdkWaezfUB7nMCm0Q0g2dE/idjXo
`protect END_PROTECTED
