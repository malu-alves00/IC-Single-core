`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XrdWBCb7YTk9v+pNawq4rLSVOfH0f2NVpBenI1Uqdl7paLyhxSZjCwF+48bM3Wfl
MOlRTyPiAel5g0D5JyJdkxtbEwCt3122ClapfpO14WrjIa48kLNG67DcMPlnT9PU
pJsbVY1j2woc+6n04ffAPYag9gFOxa3K9PU4RdKANQDuwxrfQ5jRKw+544rxMG14
KZQ005BZsoXVoJ8o7atb6z5vqTK6AxRrErVCH8Pv2iH5pyv6YfzB8owmSpa2wPyk
ggAKJtWDfajQLC8KFwSWV2sIsUsctlW9TJqwxoPKs2ZGS5MNAAhqf6tVDVvsGUxh
LnIIZOT7Ta+9FUgE/uIHJ1Akbemxr9E7uye4Gh6jSTQ0xsWacdR+ZMDR4lcngT2q
FT6F1PzjZeAadk851EGu/TIMl+VvE9D9FSLwBXjOEmGM57fjjH6T00KYu56j5eIx
/H+fAaQ02eDxXpRuW6iQY23y23qcuZBFtO6wP13xeoRjeTuThOJvunJZvmL7eJKT
lndeMlNy5a4Vuz+RCNx/34gLuFFYB3zK4j0Pqa9U+2UVFXuSTsp0jRrm8FQ6TXdV
R7bdjG5FdoOfqj7fAlqEqefwN7h7td1SkZcveSXIhxFJaBFVY6/efiNHqB21HQXN
GX1yqR7r/GkEcd9AjBfyLuqQvzQ/TurkAY1UHbkJvtEVu4A3WzTD/irFzdRSGaN3
8MTflXBa18hzRUf1v9aEma3qOftWdxywIcsIrIKyz5fyoLPyA0eCP9zm9dYeL/2C
+GVTbLuuAGE/oihPq0L2CAtS5dA6+vHr/Zsn3HxdztpxsgWRsAznXw+3nMBtflwq
SL3bo+9a2EHZKKwuqrMPAVAO7I5Bywe5YxejBubG9zQp4lD4+VqItioV2gMgxIet
j97y/WOs+XX3rEFI1Rfg0c/UttOI7Jea5/5f/jo/TkLx2As9Gz/XYK79hs6whfVH
o8XS8/+w3VcquPXNut1mlktGkY7AMlZu7fOK/SQrtu88cpFF98XnTpwuBEWz1of3
HisVaULGEe1kMHMVhfnWS/+90Dpt5k4uEnf7ZBqx85lzMH4ViVYvIemNhNr6eikN
s5AFzFDJAwUW0xlpE3iV/4j+uhhxTC7ajq/YTqXYwxP/H4JB7Ce8B+apOrRDFOAq
8xl62NmzP6r8YZJ75tfJCJSZWtHkt7BDdYTpjj86hiuqM4GtwxHSEOmIFZUAMx9i
N+3KCs6FHHeZ1un7LD/RbaI6QEFAHjU3XUdOKdzUsdzA2NfknwSLThulJ6A+BqRl
ytsEIcWTbcPuNmGw0ee8hU2xRMC/YT7nrkORBU/R5+iJb5Hy0zUtvSWmarIqa7b/
SDwna0qTel4mz4CfLMeTvASD9M6j0YxUwB8y+hhMrBqsFRyCBNCUGerm0noADh6d
y+nUiVQQOotDqKMDcdrlXgwtrkTljsZdDxxGGNaZA6vXqDU2gIf2qfs1SXo759a4
gNkwDkZc7qFl5z4jw5XV0CdLpUbT8xe/1nzf/YtCHUcFMLVgulLeNoDSKNvetzCV
FGLY9CMZuAPbz43lV0Hld/R4chUDW7Uq0xw7drHMTld12kUQdQAD1vkIn86euRsO
0MjvqSWkSuxqWtZMVTXZCiULJL1AFicS7PGCr+LBeKj6i6MVt/ZzTjL8qRqvFNxu
gQKMqk3DYHJkMZW1LCgiTGgFdsdcqb6MvFN3ONjJO+GyVRkwDpDOCUPIU91VlUEl
xX7cVBaIVzfTa8G8xbeZ4WDrDk4EvRgL+9AXh8dOnU28JiADPoc1U5p6YzMnUDe1
HuaFoFK4WAeAhR3O66uCGyGn67gUZmhv1zL7k+XHsFRD8pOPvsMheBF8eDOTPIfF
00Z5Tea0SZOmR6HoB4fOIdu6nyke4ezdA6uIAz4LKgV7xIZ6VGI3TWbSdNmj4Tvd
Ok6n/46hAdBR25emShndvKb6vHZD/ZWdA2m63QtufEpdtkxd+Y7GFgdP4MPtxy1K
rvyLJMb8trw1BqnErtU7QyXNg9HSQAXolH8tM7BB06Y6rLipS69OZTRt0j7q7zwP
LCm//+ko1mOYtRov9Vz7JwmbiCoewwNMJsgw8y5ZtdpKQXuVGd6FbndNWSIX3hdS
XQN4JKGYalyT/uvv8wl1pA4Wg4e11NBra9svPdZtCNsznxRmrwLa6RUwyI8kn+cC
G+awRTYUAZfDB8cSfvZ0JPWzEIPL1dXxKAA63S+5oeFSOfFRIGLXOeQ22xWJp5Qk
OEehdlx5UFZAWHfjw4fIH9SDj7dJ7wEhMqETiBo8AFU6AT+B48ePeTZXZd9ogoqq
jJkCpYsUqYajZI989k3Bgt8lav/Ogr5P5VQhrnkHpW368YScRXJf0Z9dviYnrtjp
f8VPmGyyYdhENFiAW4bJBfiqfDlkO1EfmEaAvh7w8OjCb2Lv9CGl1fFuJ6+2vHZk
fIeGLm7EBO9hAkAnovZcRH5Hcu+AiH5DXCJvqqXIJZFyFEkrgNFhHCzazCV7fpTA
7AQt4ACKTR2zUzrh8T8Lf6A1TjFH/NS9LHnq6Jdc0VyNmXvtkzLzYNw+JdWARJ/f
03X41GdG7tlKKE2aR+W9DGNPsvLPOTHRORR1R6a3biBOopHBNhpVLCPB2d0leoP5
UYetGkqt6+VAoIQjMQKc2vC/QhU85KM9+5N2UhMM2ZugZokiDLUSxKNG/OzqjA1e
CqOo8Y1NSh3NpcYSIlkiOE+LEsZemfpFkrUUfeJ3zf5AhQqc8PPkwVQ/4Qt2P6Fl
O99QBlJGYPhdu6F8ZP9PUCC29GmnRfOJaqrTT3O476hrVIgMszArO13xoj4cAS8d
5ZUjZodjOsvWWLmk5MRfToSpxQ6TyxAENW36B0ds4FvV5jv98DqrZJEaq46JW80V
d8Pw9hjd9qi4ZHfN2QFpD89HWLqo2wkKTwmlqYB+Mgo1gbUjh9GD8N1+7cPJg09y
fJeXLwAQ9lUl8WE0i7Rk84FzGCxw4giCs6Tuvl7R45o7KdroaM8YSbYgT6YW6qww
ftVy5zYbwnV30LE8WubArapcwK/tqnJ8T7wCBxYoTZL73p1kdCBYYR+Ss7u5/nIs
2Xy2AkCR+yvc5L8bTHWbT/5LKi95WdiejOoenUd/JoKZf7utgDSMgJnt42bGHbDi
4GiGHHIyZW2i5NwbSx85ozbtQeD5oyKNANG+w0hEdD51wFTgrg56ycy9v+bwXNvS
ruHlEcNuaxWGw1sudvXmp0MXpK+E5McXqrhL6c+PEwZlTQ9xkjBQ3Cu3tYcleeDx
/e0KYboqfbLHLS8JHeT57l23Vvz8pSgEYZJxH3t90TggeEBIJEpeYCp7+df0d0QX
zxL0GyFu6K0SDbCgobJlUXkgztIPFSmeDngsKDPax74GXrkCsa4t/nkC69M51wue
/DzQU5qALD7/v/r2z4drA5xYi1FGIWwZyF22phvldmI1ULd3KoGdPUYesJ1PRiWo
s7f46KZab8UKomKykvXElFU1+ukRACt9qC34f744gj+C6zozsEiT3tcsnx998ulG
5MqF90mjsM5Sv4la1cb6IRtzM121VIpYjkY0BJsWXzgprw/U5uUsooNFtY+lGpcz
yl0I/QX+Q1SJqKtOyUv2LBQZjbDNVu5e9m3msTLut/YcsYCSvnwbcnHhuWiRveWD
BKLoyXN9zFd18juPS/9VGMUKlksr9niTaa65DTFgdIe3wlt50NNrXGNoPzW9Zj5v
qGfs63E1hqCZ/BzpwtnlIsd89S6QwrUSIHbSFR8VNISnVLaOOybIytoeJHDogNgo
uDy6JMuONfh3j7+Kk9gufJtIGREnO2Z+pMmpiFda2uMIyMUApreRUxyNsv03ScwD
CUrEcxfo1hJ8DqWezz86u7lupKxWzZDRbPNi2usWMsMvmWOqtP39Z5xRyYcDPSzU
W2E4urcwQo3XIUWWv1mJZuUgWRDXB5FU5EN+/c9ip7y37PBY2Uqf09VJUJN9W7Un
dQ2zdOmUFPF52mk9izTDeIKcw25iIXwNHqIblFSXF4LtGZ515+VFtgKU7FJdFla/
3IVwis30RxFwykV/IeSHJohyHg6nS8sB6K+K9JckhNOrJMG65nNckgb8WJWEv9rh
apv+eLVa7wEJDEdeFf6GsSIkwOlj8/pH2c/xt9G/uitB3omRaUSyPB3pYrJdUvpN
DDfNvtoe4dXt7dmBWgPDlBoidpB3W6XxSM5FKTjAmpaIh8GBqhov6QL3TDHxPXyH
ERKcIeNDDHMqnMNt5XIt2i4nKZgo0RdFzDfAGb3QeeZT4UNkC7rIUrf+FpaTZ2H+
OBkueyDWvXV8PHNIC9wExjN8E+ThXt9WXQGn3laXY2Zq59aHLi4y7Bbnq9pw5mab
iWe32wPPmRimxey0g2ynJNy8JodrxfytDJcUlJ+ST0T/mpw3Fv/18EFw20/vwYgI
AmVZYr/w6uuAu8jK9KPYrD1n2oaTzTgz61XlupeT5aGUfdHMfJd9UDI9G0oeYny8
O51vpbz1MapmVPEPomburkCJISiDn44EdDm+WtS5TtSTgWeASf1qxa9IdT0ElJQl
CU90ZiL9rF14M1bhAlx//kAFPTPuusqf52dy4Ml5Ln/WqQLH11JQu+fCJLXjwQ28
01pifNdLorPwOVIVQTUzNA==
`protect END_PROTECTED
