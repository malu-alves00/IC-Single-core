`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
44geH23LoYbTsyiin6KTGLnSObxjJo/UvLFk6jEjPZzUOz/pF/cS2CtJMcTsQKkb
Q3csy+74CzABhUrixs6fkZvmG+UgKKhX/Jl7g2yk+6ZngLnwAv0ygV2Ba9w0GJzv
lhL1B9DZfJBYFqq1ZjA+7O0psQPIzkhL8bPoA8xONF0Gys1Ov8FsXT/iSppyVzWc
zMD3S9a1fFFXO1tBTyrcT2Fq2aYOBmz6v7Ekn5Xq4sVgRoVHYUOoQGUGR2akKlNv
dUSLxtCd2Ne1j3Y1yKjB/fD1AY0RnhY8RKebkOtPqEh+yF/mqQLd4LWmjU4N6EGK
DNYO7V37z2XluyBt/xRLNiHhH/6Tz2nO77wUTLKbE4Qa3XSMS8yTWSWPhTAcx8fa
MGtJh9nkl4xSgwQuNdXp/zHkx7cqviWtMyVVeXc2GlsInPRF4i9JGJX4rpw+TXPq
QdhD5eyVdBO8lVvzxx/I2BigmwYDpt5PGDVdCCVVwTqUyei1tNfek2StpeHZYizU
7sRMVvAXmIan4cjqZ4mctVUlDIYJpN0HHTr8OVfc2zHLD/HU6WbfhOWsMVNKvf+V
ygfBU2z1sDyMGnbFlxnVVYazg4FkBVK/x81obUQGCcHRFR9G98BosF+LbhSCmv1U
0GVdDkgyR1uuAmLQudkgfNiNkkLzHlPzBCsvDnArbzrS9AuS1TYDmz/WvugEawOT
5w6WIo79qifkcU2ZqleNEtJyIeB7+vF3Ucca8PECgQxcRPzV5OsnQ0xUt3jP1gPZ
7TJb+OZn/BV9ju+NUtSNp5atsOM0vTHMN958ohWTZ2V6NY/Eb12DvgU+dlOtoFr3
BvsL8YqWDQIknF1qYZtcnw==
`protect END_PROTECTED
