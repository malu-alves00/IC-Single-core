`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3BOh4fL7mY4Gv0ezoRG1Inwsteu59t9g6kl7bFW2iQta2BWWxtLYqJGqVMECAXrn
Xje/N7pU0FWwjnoKcVXU+lNToR9opmplQhVtM5kOSU/LQvliEdvI3Ycjnxi1sVGU
pvQMIFvTA8ydK1GrbXB/uEIApNa/abUldU4UcbPefUPu969xOttl9TFmo5u/NixV
NB/46Vp8DF7uvzvEFbkr7ZPyBCZRmgTtqge5AFjQ0EbuCIvsLfonupslltTF0O8+
AEHK56xlk0C6ipWtkSLhLzGDpC8JL9+ukryZ6qCCEtJjeOP0FZxybFeOEjxZfMgu
QtMN4VgfTAKD7ZATrrYaE/0pkU8Ql5o345SlfrdK5kpElsOvvrQ+J0Y/WU25S70K
xsVwbUduJZxYHHa2SnG+yShpL5R4mv21vsShOuZggl1hGjY2t6Aeka/dvIUVlxS2
XfbnnSAq8cjwzWvrNpoELXU9ZN8m3kbr4BwJulDY/FA=
`protect END_PROTECTED
