`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dBOHSVpNziWZMqZkOcDNABiA90Cj4G8WpMZ4QrCCHTVS5vENWOeA0ki6JGPnWuEB
YJMTuNzAkcz5Q2X0/vL/I2C+WThGG/DqIGZOKbKrwsTj+IaOlBbCcpXw8iILxBjj
nQny2GtRKn73Q0Jr8TvYtw9PlslDPKgkSZjxXq8bxS5v/SwSIu+d83tM0Np3iJtF
Fxl3d++VUc9H1Fz/8L23MAjbI8N+ocA4N2LEFpGD5eUEW/ZssM24L5coy1oFtvGy
g1a+Rpfxwg8ryHgTBD5d3ywDvniN3trgP71ZEvlA9iH7l531UOb7yPZL7uaC55ev
yomty6HRqNZPzuIp9jPaR8U0/x1CQjkxfWqyMBaCszoOtnKjZUzebLN8IFA+qHCp
cp15XiD8XalK1OtEE80PXWelQO9CaNmylFUaaes95T4lJ7reXDrdBSsClhB2WhZw
7gHnSt5rAbhd8eudw2bFp0bS6d1CQNBECTi76arR7d63k5/zHNCGsYC52G1cWoVz
Fweey0rvOM5X62BaFM+fAwhRjvaDIZHGN7Nf722Zdu8sZBGxqmmlV/F8f5+gzETx
DcHn2i1QoXNtb8TMZVBUo52/GFCf0ZJSsd6tFu2+8PRlBIgAK4lmfqNc2LW/AvVW
8RplMvpoPky11X0bZyCutjtyPbMo5vtswSGP3oQtWII1rUOplPoVIt8LOSWZMb/u
QBtrIU9wO6ROg9VIn08yb+EEX0mEDPAtjLpRdhnx6i0uO8cXtDyzNmPup0KQjs9t
MBm/iIoj00Ur3GBWqmuXkC4OqFPACBhbEnVf1yaizkew0Owu1sBLoNzAbz1er/hV
loFzbAvJPPta+yposACWGp/LXvAvOav2OZA4OlKzXdGfT5+fJ7+Oy0qBPqeO4F3o
IcdQ/cWKWLwS7ccKGVpHHAUXNZv+NH3WmKgCrD+Gqfyyq4NKQuM/muxlgJBZORiv
`protect END_PROTECTED
