`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3bCTezcCnQnOLlyzMRBQHW+EJWHq93w0Grmnjrbyklnf0YNKW5kHCxco0bEhRfyK
uDuNntdzECfZaEkiX8QTWBcIon3QSgbctH2p6V8TFCSByl1qyxAiD6kxWNaTfxMu
QMPH3C0IUfjK+iLj4MK/1NuVSEUGCX6QRXfqVO5RhCPf60DuaQ4zSJyuEJPidzrS
8wmNtzsB+/AEiv8pwS77i5OSLf40rxLmVwWiJiMimtihQnDIDJfRqXOsqqvQOQsM
qFe1Q8ZHQHnjoW+x42ooQ5NwSUdr1jEt2GA5eDRBUx0gVUFRJyoUxECVqEhSIDXW
4rfhW2qs7uTx6M0vMNlrWe9qysyOOT6C2dAbOM5TwBSgOfc3E/3U6QWRjxA4AaT2
PdJ2byPbOLJERBIwRI620Gp56Fjz0IcW2+uFnVMBz+cmo7iRR6e0/dHhnEtZ9xPJ
UbJ67TTJ7KbiRLCJqt2PEeephfnQrZGQrSXd9M/1/z8stUTfFzPH8GrXaBp7TQdD
/8O1Zo21fJQ4s1gdRDgq2Z56H7oRPmdN22BvlOLW3OaKS6VwveX6li9yDMXGw/My
4Mkh8j6WuiRWauDlK4lPDaeMpRzgduaod30C2PVMHqHbz/IiE3CObttbjsAjovyP
HAXkA31WQ1y6nuxugVnjUGFAp7wxEBlMpMjPQFDbgxb9d+XhnEz65Dtu+oQ3aiS+
+df0tO21JaVoSzMkGczZ8uLNkUXNaTYraNbXhWBodqg9DCcLLVsv9crNZ1YLqcc2
EB5SHJd/pkFnyZF2krZRfYB3duYYpu5YrFm/q0+1/z/3+4rUC2nokYsfEZDyfR4Q
B96aoCFNjPLcZipHBvNnatuLWaUUI/dDAC2Nvs6lJCcPQiqisvgctubyMuN3MXBs
R44f2efecg8d8c2XqHbIr63neACJMkFlmb7jHmEhCjx9RI64TppVQ0YP86TvonJh
cKyFhr5hH34p3E3YE5iKO+rRxdJCkXZ6WEo4PfsLK+GCfuq68BntVjdK2KRZ9oAx
yxoONtC040EpPLEHSsUEPmQSftRRCbksiczVcW8Z2oTqahnFxTmzZDaUGqHhmAYi
05CTnSmX/hE5HxQQpSjpUfwCOm1sOYSClldoZZTPzFTW/1JSrpgM3ORKKCMBjX2p
zDFUarshhuzYdrcF5tDbNjZMm/dNOi+bV86iUOQDDH2IJlF7knu98chDZud4iWmz
vbe92byZ1L1JAqmd5gvy4cCcMTy2zrnzO1U0b0DPh5YzYsyfA1mm5MtmzimXM2W3
/y1smzRqBfaeePkwOywmR7IpyGMUw0bJFQkzGUAhaA49x+dlZRHv52IKp2OCGv0q
DaJwT/j6KIs9LzLk0p0tmivrYTaWe9xeJcc2yCCyhH0MV8XlKKUzinqMP1XG1ZiM
5t8t4A1WFHp+TgbRKJ+EGcWCeW9pS19kEr5AHoS9dGiZSc+K0tStpeVieprAp4oQ
aaN95n5MBsfdOzYUKXux6h1N+YSVj4vSLyTd2zeIpLedObl1DjQG1VVcq9F8dgaK
k1liFTqf5tBNoN6Y1vnYX1bbed6uxDMgI3nrVIAqGBkWZjIHDmoAtIVbMCON7P9B
WcVeg+rknRTNFVQaqb967FF6KPJfGESKPz2clv1vtsuYCpOFvdWzX+dbrEzviMt8
0wrgae5jKX458KOytIC19cCPjOVHyle3Sl8QKFXK0DRQroHvykU8kM8JerRX+IfC
Sd7Ej9FECaEebSVRYCxLgYwFHTM9Y3dA/j9R9SK3o2bySXRsJZnJ656u7HxHWbKg
c4kjBAa3FpCOtCCIWT1syyhuVJKVBLB+RoJUUdLfFTIfJpuZSsMaQ+rFtjg2TUep
8jULmrwSwUS3pKJiDjpHVx0payYXRoywDonhLt4CI6jiaLTzm39G1kxoLXnAIyb2
rD53QDBvch+XV7bUHRT/+iXRAgI/wrIWk1R6Ar5/VDn5ESFTV4KFLtmIaJpdv1+O
wt8b3K9E3HHjABeTAdrYewI1GNHp5d8D6ubhIRYHvs5sn2a4lxmKUBaqk8MgLrHa
RUbR4JKbtx0uz/EuHKnzhibldgRFyZetOHIy8a/nxHCiYdCZHURJfGRCYNrszU6K
zn1Tq33mdqsH/DH1A4Es3hbI+X9nvsvAbSXYaLnVVS7HjJgGCXcOksfSjkLaHk3j
w+Ats+b7xt177UOS/r4FQhgKSpaBDbVUtIEQExLfR6HWd6iHUzppZP6iJK7TQw2g
99dBQS112GtpFohrDktIenguKMD+1FZIP2L73QBAG8V5at7JPIz4pbape46hFO21
YZB9JO5cLJtioqlZ3L3k+ilIFN6urvqyDnJxp2aR9aCSsmLDQCuuletl+wbDF9I9
tHNo801eWsXKWIQ9xBjBUjzytL1R+vQrmyTvUP0ZNWk=
`protect END_PROTECTED
