`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bYOQiACy9FyNa3IjSnSwJRgkQKpymQ3ZBv6EDP4mcrTyFnbD4VmciZIIcpuD6Jxj
W/nRJWaFrXCBxu3TDndynjfws7YVj4CSjaArewb08cvACKMyu35smRy1qAaelMMY
viZqn2NEMswtfQGPID5DD5skE0+75JFo/Bu4HDiW+FM0/7S96gf/fRTPELSQXMSa
qgyus6HaTB+e5+YTXq5aitpkzkj76gVARSiRPmqkSXE4kWPkRmXfCO9uFa0lfW5e
t44YgoplovM4y76J981yXJn4o41auUUFjIkOv7FzE8Uh23qxaptHleeDqsPqjKqx
j9mjrbqcYQvor9+Ppgs4xD0YHSQ2oNeS1Se0m5bfjHzixnjC/2e0kH9Xs+8Ohvtm
XlWvmX1xdrvHRa7q7jSOu8sIhZL1tqHHi6TCbUCfiv00VnsPGqtX5XtBXxzC8tZu
6I5rK4c3e5Ds7vw0p2E3CMcmUMFdgfvEzBczJi5f0BltSuHygryazRBVgz0HvLsL
N3S3RpXxjcN6LbhNOIaImH2nN4luTSMo7Gs53F0UDRywqh62lceLoL5gqOTQ5E0L
GiFThtu5LalCdnCrkyv38skhD2hB4Ml/6ZpMciQaYWWnrHx5rQgNem9B7CQeVF66
lsHaU4iKyfMy4uhNOrR3PQ==
`protect END_PROTECTED
