`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DLDnzMCJ71U6gaArfNuSPjnGZIr/+YKrsrUEKUUSAn8unK5rj3FN9SyPj8lemv1l
eApkbh1e10z8TkJwVTi9Pf92ionC3dBDdAtyFdPNrhx/Gb37r4jnlQp8COsD2GAt
iguMujmWcGas37duSoeN0RhImUhrwf+urkH0+5G+zqTqbETxZdZtMsVAlHnoYc5i
NZEIcrw/Hb1EAzfJa1b7tkjmZzMkr+HGp+X5APkWhwcxG/8sc84J+x7MaixWu6EU
GUOq3Gzx5i6PJl2IyWpo/bqGZ8FxGQytFXV7S9xocoflUD9c1jJgDNSShLK0+DfU
jeEuXQlVqDBBnDMRuuUXyszeLzAFyQS2lnjf/GXDn7tdmEhmq0Y1oyp18Gwt1Q2N
as3eLwTavqOZ7YmwqPJa8vFPbxHsfE49qDmgcG79HM57ZXBDj1JZg7In4HmBPOBp
dWx5OrHK84qqLN0S9uNmNlDu3xp8fTvl92pttButJ/7cGN46arEJ1Kz93low+lWg
z/ArJHeuIln6TdaX1ffz1umE8xdmKIELskiWt+ZBY+jARcLiPpvBYB2WV3vKaTmB
UBL8/bqTGohz0D5vhzJzOmMbCt2KafDVAXSO8eGwlUcdHCsudnXcbkNKkQOUPvSz
QxfkcpR2ueUIlja9ozB609jeoX5ttTazbNAM1N5T6R9TO2TGfai0f9qufDBVwE2E
MTz/cymhrnF0TIP+0XCioT3r7b731vGrEUL0fReBIEExZL40hRE+bmLqnQd+Dha+
6//P98IZgoN0WfdvkyklhJlwQmRyDvU78HzeVhioh5mhQfXUtoOBsaLUXHyCNQIj
Do7OwNEZvyLggiLLiRwILr8HhVKp8tTzlNM4QMRv56UMcDc+J1Sp0YG0GeUynw/1
5LgPYViB5fGqTqjiSfJNXifeWJRiYqY6rgemGU6j/IemjJxuG/Re9zQRpxeJypHN
+STfSZeCZuB2cmGY3+WszKEKxmuUw6tkHcWMReQgno15E5XHp0/MiaIiN4eoKquJ
A6RwRsAL8On+AnS8OP6FgcGgC2wpnmL5GF7FmIiKvCPrUMoC2838pUrdk0j1fVWH
N9EE0tZZXo32CmznXM25ZTaMmsqgBKAnO1agutI13SFIBcJA7lqM7Us4Dx/k6YrB
db6aHW5X1/HqY7pIuCsBkZLUcIPfsq/xwJFpSpnIT6ADpvaFul8b2cIfFqoRXPtJ
b78C9l7b3nrOBBPfLTTbWltRqvC+uk1ZdZVar7CZkySY/hSsYEHrkY/59DL896S1
vJcy5+c2GeQUF4r/n8ju7IU6P6FmI7DBkamELaQ+vqK/oYIQUMj8RPZT89yOwX5+
dSzYh71M3RuBfEJRRPQ9ntyAlRzMkuhb37yIF3vhXqL7RtiJXcp3nya5KsJUOONb
ler1r7yz/UhMRJtPS7inNrxUuaIJodc9uoDLvGC+KfHu3iyFYrRV/SzKkDdD8mx5
3IwVW7zCyHVFg9tXwXKxR0dnDQ2y885D78cvOGvOj9uSa/NLJ12arWYkEgfoItjL
5EJUv9e3j/RAtPdUQIm5QnI9SezHxYZoGNgdbRPLWiVzbJIbWgb7DcM8EIkFX4ad
r/7L28QRIHeu0dE+ALYw+YQ1at2Kz2GH4HCG2UOry1Pth0rIrdvPbxpwWptzcjxC
vomTpNAGhx7pRLvjqv2SfgD5NHiiWnFAgJeH58afIJ8jIA3LU897704hR9+vMkmT
E/msAVBt1GK+EJlkkkHrZeFpjDK9lWe8R9lwN9EggtistcXMcHGWbuh/fUy0ixLt
zVpVDhYLQV6XGPU3wX25noBPNvAe5Y0oWkOur6wUS8ggMfXM3gsj2afMS1My3hlb
UvloC6PUlT6VdKSA3Pnys5xFkbe+acW754UaWCniuBClv1cKIQ8jFGjZ3Jbc/bRE
U16G2omr3dbtcyd2z9vCW0Sb0APcP0ldlBNAcIBkAJUpwW/89ml+4xGmViWO5hWm
4YWVEcjriIxP+9l+WXKIU8PMs8ngQb5U1xFCOVbU9gACtoTxRLFVOWztD/o1JJ9n
0clTBtvDA/AdI2CpQgzq58DPdZ8T4jstrKoOcOgroKYazFhyojy4ymZiMyYAleRe
ahd7Zq9w1fP/GzDknpvrS8qXhOJunYWZDtrFF8pWSzc5ONB5/aTKqimgSSffY5lB
WX1XmW+nFUV2IY07VNRX8gpR9c7QoGoV20+/WfxgTxXhCm+YrhZVZ4L3um2jSTHZ
UpeRbrxu+2gNvTtGW4tmp/WI7jA6ErPF8jIURBV6S0uqkVqqWHOjWFVZP0D2EtId
LKc5jM58dcFhde3AozKRBt287XWQkqreFahGrMJDvYDuhPnqsIh2KBWQ1uYsiWdU
31IXz8c/yAuLVU7XPdX9gQ0X0qc4e5Sj1xR0iKyN35ugefRoNfhb0JkLbvBoJQx5
K5buZw3gFgTEjyuxYia4pwYhsM+TFs3XKNaWUgFUhnutdji/ieF0irjlFZhdxehP
i1oAQ6EYyGG/11c1irPaph7/HF4jWvV2sIz06+QuKVjR6xLJGKuZTeBlGXb8HrT0
QEd4X2jbqghsbPYt6wi6VTjucMFGtSvnmDAgR0FT1IxhpIr21+Srsa3ZF2/eLPBg
FqaIY2z0soI+BqKVegNe6yNE+PnfwX0b1B1w9tqVzAd/gqEPYMxMpVs57JQ+x1+9
FK/IDeKA0uSgJasJYQn9pO7yFsMi6w6K88tB4xHD5PnbTwU1arlbwBFWfZne3+1W
lt38fxWpaLdTtieOaGNjxGKIeyayBM0LMuBB5Ro7LlELt3z5Mrx4q5l0pmuSQgbB
EjEeD01MTuwF4HwCXupB0fuLvrYoDt9A2sSR1oK9zWXycaXY8ouiloiBsuDkKshJ
QYkcyfO5CIVLRGYzGOZH5G1cdZdeJsbJnSt8zKHXhKLS1lMROYpoahg7gDdpk+Tb
FUUyxucyh/wGYZeF5zuMB8Mbg9HndnOGGqG7E1SgoyH3xyPGqALk15EeWgUHV5Js
jyeomnEGPQePrGdLWVSC5nZfn3Fr2eVndiRdvSp0+8cCX/YGI2XoprzNqKx8uutR
cQS1cCzN1v5+wCp/Gz1LEmhHvkajC4SFClahbQqMAA3TZH/p8bA0WQcpHUnku0u2
N+TxgF1a/6FxTLqc745yhQeC5zWWt8AcCXXS8VkwJ9HCnJDy1d+wWENUZ7t/yC84
wemcIM75S2h4PRQLSWrmZtD9VFdDgZhyBC5khrS4oIsWETqDX7+Qv2UkwuLB9fJ/
OY0MONqZTyLagtnhxM6yA7fLBFb7zB7fR40xQOOJpMewonq06EZc8NEwaUVLRt0x
Md6UPEkbrvZpGObvPdjsx2DPyjgP+hQttYtH8iVi9qGXFATTEju1sTIdk4L7DKQk
NkLNllqf/Ol48O66pk6LPHOYcpOMef2P72KsFdkimXM2yt0aPotRGXPXpRYRAEiO
0raQJWPk5vaw7/cKWVmNv7qI50Xkz9AOfasbn0Q9/mfaSl7UxqVsFjjL3B+fuc+x
K2t7IJlDsh/Ntmx1wZhZT3cVNnh5fXRctSarUnOXqTnL8DmlDCbyIUGNsuKcaZbB
PZaXoy5dE7FcowlrsWOIGO3VHQeH1CkxyNWAgPYDkx5k9pnuy9EjZFg3Ru4OiBWS
jjzvnoknRqvNZAK0AqAnyHn07DdB+a/Jd+lckdRLlF6RHOcRxM8FktVfC7t0RflR
jATEOidHyqbIV1A2p6E2Srf+wMVzzLEny8j98mB9u3BHdxwl+enINTrGJ0cUN/zC
eAP3YSeu/BX73f4q73MkEq0Vrn4pe+uUoVC+sqgbRXUXGbhNU/1jax591KpdjbLB
+ySy9h9v/eT5HOrzJ8Gt2PSHSl1viOBnBc2BxeH3HAMBpBsdGiuxm0wbnpgp4VNt
H9dygOnyA9aUhC2Kh7yBI151n1NRKH5t9/jnJ5NckvtSAidtKz5Gi3HOFixST/DD
+Z6ZtmlqMb4EGcq7cAJXKb8+JY3hwXRT+Eoa/lA4WYU9G+oekgdSpwPnUoBYdQnR
G2GPByH6KS5TT2whqqFzBJuX3CfPB5mBDmalloRxH7FxI15Is25eRuDfDbXui8Oj
8RIHpgnJWFoC/0Hpjd9uxtUYnF8DW2+/mDV6MtbKFP1lO4gZkuZzmyoL2t872ksh
Y6Rlqzo0/1p7YMEHtL8J0cbm6Chrl00k6EMEqPY+6hc/ssUfB7I5uRNrbFEnoJ8T
XSQK7SB1DI9Ege/od5oKRfyNRt7LKFWJIY8WVCyTNJUGm9VNHZSF8EXv7/kyhgTM
gYRC454K4VxAYvSmjTF+fS3k9Ngt7QpyLqyRlzcWCI3rN6EtfRA1NzC6MCNY/Ahh
pmVhSzudVlnYVG002yOrhMVBOXTt+loz08ZRwJs10Hzt8wD1rq/jlPV0S+BGEhaf
Y+zP/uE/V1PN8pgXp7Z0Yx47aIUXiPkRVLR4lLWc4ZTWStyGhLgjOtsTcuokqKMU
d6wBWeJYlCy+ENNChYJ1eUyaPBWyhfLrRI3rnYzjGCUWECprB0CZYLvdU5MiV4tM
0H46rXVmr/LZPOS6f5U864zqx6GgbyzHgtwpZSJZsVnEDOVgt3qBDHZqmOq7LJXj
W5vT+9DQJ0vAxCGAtV7HaIFrhWaIU1PNFK3BJE2+2JEruCq9bLN0fK/RLJ1Sf5T+
UYXDx536ICRluUJwQktJzkJvOlwmTwPMvRiuGiQjeYA=
`protect END_PROTECTED
