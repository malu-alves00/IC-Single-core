`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
o2pyn9R5fhooqNwfX1nczcr8WC5T299ozs8pFFXBJi3qjZKhqKCxn8f22uN/rQcx
xJ0zby5VnkBKHaTruUJgWet+3PhHh8AwN71HfdYNch22o6u1UcEq0iUQrrVgCHWP
UAFrgW4ec9nZz9buM58AqAtlvlxHvlDAI6TcfBxsiR80kQ+L/wQDyjOHQr4mzwUJ
0g2YUE+CmNDljBCA1TaheVecSeUJh3k8o0aWsyvjQn+/A5r/rxC2ensP8LO5vJ5f
ChUR6/vdkV9kGoPTG8xQ5IJuhoVrMVIrp1NWPl+NqMZuTqY4SSWV7sEahVAz+XcY
bn0BcVFP2BTA/c0QPsoRWuDJEpXsKtuPt9MJTzL3yYMwCUksZltIQ+VEzRfvwk7O
g12iiKzyWvqOplqfQXpwqD++nTX+s+Tq6NQ3hqel2KNUv4MLyJHJWZBca83fe3SC
urWNe4ZsBvFX+7BJRrBlHQ5KR7wWGFndffO9WKhLecgHfGDTMg6M42XvRv2ae4Sk
7waeUTZAJaB74mUpeN8LKuH2tPKFsQLBR6N+Sj8ZS/AT2UhmwIQYXVCkbNWKprA0
w03HsUII46M/HCJKMtMg1uSeXakMhMmIk+EimrkWFEVli9Sr2l//17+h6AGyz47L
`protect END_PROTECTED
