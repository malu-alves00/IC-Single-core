`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RmEnmyHXmEbBM3zS9/2FvAdImCbS6TA/CGTktvkjLsbNczvCxfZP9QR3Y+/fLCwS
9gTTbo/4dwZJpTfrRHoRnEaZA5DasW/KDfLJfxgNZ4BwJJzfXvhym7Tx4A3Jb6/S
4+Z6szqFhD+R6GWG9BgXvrjPVJAheXEOefkUFxFKAFwN4NAena34qaAaMtz5rHZd
tIkA2Qaj+BINl4x8/ljjaep/pCmE6WlGocxJPaoVejBtBk58u+lnpJ2TWYjSYPOW
d4ynJFgSKKJ1cHlZG6MOSR575vUhfPrThGgxNpOR98utVqHwI3DCSMJt/O5O3wS5
WWtBoLaufdJcqc3S5z3hLRrMcjz2iC04G/Y+7pEmVvjjEj0EfhZri2wL8Kq3iOPx
fiKjRUvkcJufJCyLXpIEPwmYgpilLtC7G/OZjNFfzdiyqTQttYQRWi8zJG6QtdsP
EzRLD/vkmH5joBiHAAtEYOk4Et0unayQfEno8y3pcQIOyOnfJHsIKj9racUOs9dB
B14wwT+VkplocTCwR7QZ/Qu2Nw2QeogE16hywnphjOyK3TvVGbTtFRGoix2nV81x
gsXmkWbZ5hf3nNERb6sMBT+bHJlBIqMfUoCD5RNSI5wzBBVMnW0ybMEk/ZGeUuBL
oR+uYvR7f7uJb8CBbPXQKb+xciERnbeiwp7pfm/dqU6Q5mSszund/zgaSMu78wBz
JOHQhBudWKY7F15vvHYqLqiurYFn1na9w1H7WyggYTVC1dsHWJJ89SBMvaAsz3WI
RQ9aRgWE12EJJW5yFeEker6jJDjcoxXuUmh2cO8wr1yvnrBB71rQAuC9r7ZjeX6+
tpyrIX1TAJU0VxMjHpGTURtitjrxZ/3ZXNFJyJxy9E56dUsJFKsgRCbUztKhHB96
T9mltA0w2t95RpUkLcx6FCpx5iYx/+2JsI1CJ0Xdzxg5dyOeutsLNfXlKc3RVmtm
GRN7wcn5E0Dc467Gf4/GfSZ0ePc3x95Rh30D+gY8IrueBIxczXv4TCzInGTjfVM+
WBWoTXjzrPN/tOpmSd7WVFDP1ieii9FRv4EIfsAMoAwIymjtI8YG+Widjrsk94V7
kHinWDq2weffQYe6tIHfm27taiWe99DbRT4JG5q750UjZUYP0OCUjkMm5k55Orvb
bq68f0V1FYOi0PGJRgze+oyCKVktrabe5urObXx63tHprubVBdaq5WBbhDgilolW
WupMq5f2HsAzFg4NkjJ0jOPZVtLu9d637eVt1CNkD/7VQwyvBp2SFHoI+mtee8PJ
zh/O/snkZp3noLWIybZjXmOCVnC5PObtRivxy98xxjkciBBrO9evsmei+NM8nsKF
ZkmiCfICfifk6DhRJat5JNRJvebPoYeo2MwhtafSl2L07/WsZ9rOER3iDtdU/Gb8
RG2s8BWpB5CNf/yOgRgGepNJcLamV8MgIOhNQQFFUrYJ7tFhC6XS6K6ZKdKRbpNe
ihg8n+o2EgaAopScr0XuqTljgKBNnYYdkNN0O5o2dsiq7eiXfsAp8BbzVo6LK7we
VeyFGhW7I2kQNyB5NHwHfCsgB42xtaGzkfWR+ZIG0MuXKYKVuYaCHanwdYv5ljZm
3Dp0ZX95c59gfdrD9E3Eb4HWRL7QoZq3E79VjhaYbPZischlTmPk1XjQGgCZ5ZFr
0qQhZ4fQN5Urhw1WB1pqvH4gRQWdqcmB4K3K/mMVdxGWdG+xEmmvMHnqXDmYzHl0
MMzy8f0A0ivbiQrchhqKC8TVB/BFgebN08iyDAl7eEG72S6xUttP+qWsKqyEu1R8
2HG9uZ1Fi0N+DOJYnZ0kSqvASbw37oWceMIWwRJaNIhF8CWui3G32DQN5COf8Yi5
YiwVxj253kMjsWWLgviR1nzdwh0tKDu28ibWR0uNi1Kk5DiqyFvAwl8PiyvLuQqR
x9vmsJGM0fJLCx9g1gXDCewcuSBA7vkBhdLJOwT/FWEoR9OBQ/cs36L3b8oP0XWi
dbx7yZ3P9ZySH7Np5C+FQwBQiFxRkZmQlf545gUsTiuTf/exuclv8US6yDDB9YFY
id3701ysNp3tfkDLQNQbTbvSACiOXIbDtBN44tryuzTLPEOZpzQC+eqyI8ehqPkW
/C0ELGPlqs7QvK7xVSksFzxNE/lCEBj9e6nn2BiltbU1bs3X4Phszbkm3kWxDySu
2XbWzX2CwHFkfp2IenfytmPfe1f7ePDeGx3bK2RmMH7OgCwDV0EbrUuEGZlmZ+hK
pYSRW/vMDEoNs0Eryacv4gEkVp+G/fIGiCqNmluURxsVk7Nw3TfRxexfeHnLtvdK
KuOSNXHvGLfioXtLB+SpeetN4wj+oPdE8kNJ4zaGlEneS5xoxDW4hPyNs41ASO+C
Uqr96/SJ58xU0RTG+QDDBHonUtHQEOntc8sYz4qt7h8kpHUfhHTVQ4+4krcKb+0a
rasv6J+bm/g/a69cAW1/0RCFgxjMbcqRyJwfXSdL6ZkA4MRxnQ9nWZ1heUwVWBKi
xtUcMZ1+OpCTMH2dcZ9kBvKopRH4xLJaFjyzttnXc7PdhJ4bl249B7ymjE1nP7eH
YZfFtfvlhuMhov3OIDRcTnMHGS0R2fb+1m71V4x8g9c56jx7K/YoclH3D7VYwmdX
Qkyefmu5D/oN1TqXnazZubPId41rzMoKTNfg9lBwpO6kysvyCMZ8QLcQfhDYZogh
wnvXrJZpYP6V+SRF8AGrouliNv7KqjxkzBDkYrZnCtzYTY3NSFVeHEk8Abnk6t8s
W7ipKKWg2QqMGUBf2/rFPH4CR90lxzwiFo3ImzMrfsZgBSNDRwkMmDNWUxWMosRJ
wQAw8ElmA1rJ72RIjqDephmy/aDa0wzCAsMVlmRkcdrCzXtyitIcvgsxtovL/xSW
GuLqsq+PWLtciQ4jV2VarezfU9ZMzj7IrITqTxBtMe9Qqyr8JUa4XpsgP0hUsAzX
7tFuVRmWxoPKpTef+MYbq1dK3phCfz/D/uX1Rf510grFWKJ/DnRiJvWdup/AVt2R
nSO6iHyeQIOyNxa941f5wiLPTMEEy4NMC7zEw6U1fHYeOssBIG+3TTSXYK8fFiw9
4n3qnh+48bYvMo1Rg0fuYTTTLmyG4KoD7bxm0e19kaSiKQGDh9hX3IjtdHElKTIP
Da1IP6qQaHz84/INcI1QOtnuPadvDkmiDjtvXGwdM0ElLmVnONn7ZDPQ3cvnXvSE
rhKPjLkNJ43bSiIAEfRVtRU+f69EgE+v9bhio+0v25Anoby3lCNs0NP/HXlYXxH+
vvognd9gJRBGjhFaFnFzBC+7Zy1FM4GrThWl9n0lpkBNlOJcPk6hC2uWQvMmYtu3
xXZArMKzfYhrQ3Bvkb5+2dAxKTekCHpErmaQtezaTODRHS648Xcvn35RHGPsUXsn
1gnoxFtl5YRJkEiWlojYY5rUbkJr6KowWZLeffMzPGiI7/mxzUAoaj8HtiS+wp4s
C6tWb+USO8uiGWOIw5cFL4XTGRV5jvVhUXwErNsluIc0j24WeGbOH4geBXiIuKmB
+7MjlK19kUP7DQvcg6TD6Ysjh2VSgafFD2RtZfze8WaOvFrusuF78UUjp1/r+XQd
zicAkwWzGUsNgG2EdifPC0ZQDFo5RIM+6wH51ZzTOHmjx40ezFt3KC+ippwlOpFw
rkvIyeaN1Sq7ajVS8T5qjwDlY9dWyQ+QmOmqnrx4INfD3svbnCok+2ZWQX1CpMg8
pjCv00YN5lKZceoaQiK9658iCKXg9PtvjTcVRo4zl66zN1q/LwdGT8eQNgy6Kl5l
m+f4AhqioSIJMOVtSImtbmo9NTXUHW1JEjQhimOBooQv2hnyKSeI9D8L7oBxySj3
lWsnNudu1RkA9nbQePALRV16OlF2JwrgCUp+cyK5wM5CIlkKu5yL6HkSi68Cpea3
z3UFL1aFOSCwOmhrUn9UzDD+eOGPN7Xb6IkcTiAuNNHnHSva7Vr9rxpupiLsGt2k
FHqWN11mwm5NaM7N44RTwxBIwMt8wG2L9JnJnKTLujgROl4q3H9bJqXSiDfRfLlT
Quyh/lACX1hcKcs2FxFgK++8FC5hxt/jjPUIi9sudTOBgGeXNiZA9IEtKqwSK+Ti
cPCaXJSS3kgS9t/ieh9D85QlnyKDWwHeujR6OSwMOqkmpgx5yxZ4YsZlFkJKAyk8
wHHjV9Cmusmf9lp3TXNKalDJ+Hic1NgB8YK3XKmghNmr0tr4Fg4bFWoImNV90p/1
HFfOBFvS3n5O32Md4LhGSYTg8+rOmNHrRpKXbQD/FOqedwry5CQs5zCSiYL2HbT5
FLyLHZ0SWwydAA0F4TQ+02aiJdrO2lYP5Tj05o4thgLhVNW9NdFWCvxGBD93JLJX
GQwzKwgG5M7uHOj8SKiAENSLseNphZ70THWqSXu5+mPS7nih2iFvMt7cf0KiYSvL
BY11a9TwhN3rTiDlwnXZU02fNvP1lTCXllw0Dv4FBCkj0bwkOpFu6kEmN4HwTvkB
KHdC17CPrCPScDE0qWAa/3HV9HU7OU4qMKVeF/HNnmz3Mq3Gif4+Ch3XGsPJ5q+x
1CdMJqAnu4Qufo0KC/ezAo85tCTJfX3R5foBpx4UoBXETTDDSnTg0hNsB77ERsst
i7fbI713CutqGoi1PZcr19o1pnPc+1gsy0U+aCYl5djvLjYuh9qsUDUa27HXDAZ0
gKMjX7hIcm7laGFTFxR8kzhQeD4nsc78qyLz6hRdZGJsz/fV4ZeSvp406KEQbsTo
+5wmr/Avf+byLzjVQZrm0YDVTrIohviYiAosJVZtk3MsuFme3qfsNJihaUxvI98M
MlXbIPuD01PAr6uBx5p5MRoDD4Tj0VUUw//wpY91LvbpKl/XI/VFS9DM6x8j5I/r
IwvO9XkCcSgbaSPC7iKppA/I43YejAlA9fhJFQe1cqvvcuK+uAqWaLDv0XAqne6T
LV4mlhRfi5JjIvFsf4ZmyXGaBBn7KUIp1Rv1q6+S5f7AlZc38ezAmluj8mULl1UB
ZLZmYGtAs+APb7Gahkjyf0bQlwEpcKnX1iGLUruFKgorv8Ice6rf87Z7pKCUn6bh
Lm1Q0iItIx3Y9vK86Y1OxcWJ4tw6MnZeHTsiJG9WMUUBz5VjUAWD8en5Yibcro0I
sOeKacAcmgGFiNSWg5K+kH/16jKH9ZfPLLAN/BNkHEcy61CVl48qQeJyjcNK3Sc0
OylpIi96syLjxjAMm3t1JRrFXHn/bqt/77KAIxjLTpLO/y9UHLVA9rwrgnrmznGl
8HhArnlEo9SCKx5T3f54MWLNhlrKT1lOdn6NLtjJRXLKB72JYo7ucJ5n1MCZVQhe
goKpIP/7Q2OBTRPR5D6bNkX7XUu6uspIOCHCoFOJRvOSKa3w40B/rcu7pZB7WuVV
iAl+F9Kmsrw0n1AJE3KV8v0SUZsxbKmnyAQUMrUAs+S5KdnkvLxqPHNUWUE5DVka
Ciixw/mgDKsXC3OT99nd+ClyLS4ztv299V2lVGWEpKD1JnXzsWYjPQQMTUuOcZqU
D2ox+e5b6cKN9o6X1nKzz0q7fZXB48MQKSwOce3sxDwi+jyE6UgkXjA488DgATE1
nN8INsOm5+uqRMCZOneK53bEriAy94Sj4OWczUWmZie3stkeNsJsFdn0lPIJkoRy
H/djXTg8pXY9o/QaoCRAxe3sdqjXShEp/Olu4k/+g+hniIjmNUO+gmM5SQ/iLtn2
h4zkr+KRCJocWdevWijXZ2JF5FCFHVXtG0CZDTqyDTJLM9DcLed4I9wtbDDiEQNZ
KlP4G2U7PiniS/1zmIDabsOFfSurYZ+PuPA1qGOjzSKsU2pXeSYQKlKtKOE7Jdov
mLWeLvBuvGOMm7tRjBc3Dnn5w8ZRQQrciZ3YXylZ2NkEd/16oRFt5kWIW/zarhFZ
gRU5vi4V6lUFxLuB/GX92Gj4+WBcuTw05bSmyficeaYnJn2NoOR22hwY/92BQ3u1
LIuarv/3+1vFk5jStANooia5l05tORnSLXquWB4TK24+qpIcCLIxzYJjNItMl+PS
97B/5jAbrCXxMe6FWtZnogUK7OZodbOEOPli8zUxvdV7cxuInVpqnVYU0hfPBeD3
6zXjLmKclHTfa6G36LcdS7rIlhg0KydWVuWCCZpM3SDZUuWdjRPnE16YgP35Np9w
qc4TeK4KEhCx9mCmduoedbsY4av3UFN0QNAZ0qKipCtqTDZv8KRB0JeUPQi97Iel
HeB4s3AsmgB8rQBCucLWQi2FQSG3qLBfeK6GCKW27/nMI5t9Tt2b1gkm+AZC54tg
O+J2o8/zOQ4Kjo3KZeWzM6My5MRpK5R5Va9wlHvpVE46taXfkAKqMIK1qXeBSJhA
hVpWl5IXy5gfg9rCkn2IjWPgEHnlTUUzKIUA3Lvczv4yH8+1Sav9orUPao+8PbZw
/cmZVh0DlutvJDfLTKQzS1ggTO+mUUyZlCXoS6edU3uMKeKRHv0BCFEF4/Ddb5Jk
QmXoNPoFuQzNdEk64j3QEz1FmWt21w15hTedhQyn235tYDNMFokS4jEOTjWbgMii
61glFGrb6uNT7SVfVrC/j893/BcPuYNpqLgsThsNIbgyXV/h2/rXcxC+un0ovN7r
S2zkJTrYrOk3he/1eaNA4B50Pb+7x8ENHz+9dc8xDMHHnLpNNzSP/tyrm5DVHWOb
RFLzq6EcCTgtL4Rpmg9/fb/dVIs1zQ9wxelD8Ko92ARCzsak1jyJDXKUXP7xR9A3
FWyuQYtVduG37GCjIsyB7wUbZfvnxbdWWXOFOiW7qw9e/qUSZtoLU3t9ClhkrApm
6ji5mYRw5nCfngEiajNzmsAiaWfwFUswgXA+txfveCr1yYjCpMu8SzBk1NPUTVSB
FriO01Z2bZv3RHg19fCPEaquIJnk/seBGZEn8nNTHLZsSrgGRtoD5h97dZgNAS/3
/FRznWcdnh7ulmJQd3dcxG/4HmL0YVIx3mLg371QqXIQ+0ufXXdGZ3mTr8vY0jej
u1kyaAcsQwpRuY98KppLqcL3yhXYHevUqT9PG0TaccMBoESMGG5ckSaesffrKbN2
uIdew/CpaYht1A5L02EU9S78lv/qF5ppct6Ge/f9HBSfAWz4C49Rb5AR/Qw63CKG
TRUP1Roh2cL/ayZRuVctbyScaJFbyn77QMsYyriz1tAN0fqccPLkgmGgWc2Tc9lu
YLRBlmYHINcmGAH0t0Wj7Wwe7+CJnyDYhEZcHDdOVkxNcYTcyTi+iD6XbdVJnLz6
G+q8S2iLzEn+wWd6buZSnpHTXPgl2fBkrw6lcJoXQSWyniM1XnFmJuCHE91vMqij
Pbzv76CaVmoje3SgoZZwkoE6ODgS6MQORrvgElSy/biLCtE9288EsDgDVnW4lBAk
ioDBYhqS53Baufg6AwzWaFTXZhW34ip8YuSfT1p6Zj+LQjq40TqC9bwejYbBt4XJ
fMCeqa4NUUMJvu6+Mq2clN0cIXKnLxa3xsTiOieKsa5g9t9kuAxqvy51rz4EGqIq
c30zG9KT5q/wPkWTpfjx0IIp98n8dJ0pDR+vwDzLtjha0Y3MPpyjD4I/kCvBOfFf
fS9iqyODWsr2Db4QCkqyEo2FKwCbi8Qg/g+q0xNeQhoYvuxUaNPGPx3V6ViBtpU7
St3TXOtZLJJ3Zrnqg2qLSZ0TVlLlabMKtC4PT2GaMEHZi/5Hv2vCt1RMkwcq4bCR
0BiBN0vqDufuL7Kw/GNkk+OCKdinPBVn+D1/Wyb8gE0y10peFtXU6pRPEovFhHaI
EjTFD15rNlyt0mCZ+fHgekZuaJQcXGgp6x2oaa4YI1J2S0N3M2pQzjV1YfzCMZQT
d+0d7gNRrD686eHz6dRfdivnXwXUHqCA+fs8rrd7TFf+ynp0Wf1KJ9DECfyY+eiH
idmOIPnllpvpNtR/Tn4/ATarJSALwS0wInVguk3tg9g88Ns7cpyur4vXkpuXVlSm
tAPe/8Q04N55DluP26G0G5mzOvcyzoPeM1RjF/B3hFh3CQ66XN32K+l1hxfhg0+N
XEnFqgATld1aT/UrVy37yvWyRvethgrRKSsWhdZPu657mikFdex9lEjcRqT1gqda
nUuJ0LxPNbs9o3wXA8eIIOvdW708tRq/atzQc0xyx9aKWJW9BFbwpzur6IcP+WqQ
vKsAUrd8eY9FYXm3ZCjWcssya+7gcXWs6tBTDyh5RbE7VgFLgMiWpqb6BgtpBwcH
flQxNjLvWNxUpjtgV6b5n5V/ib3wwwVbJtI17s/V1HBug8OJIgJ6PxdY3sP3wdYt
Z/wlSAbY3UZ5vfnCiTXY75OEKiY4GSpd36RIvoB662dF/erjrWA1T3ZwqWnIntS9
rzbk+6j4K4VBYUzjmAPpUsk2Hr8SgTDpkwLX1mi2kPQz8vPKQdIHoPaX5h5SEEIl
VKzkwc7K6SQHAKT9cLmW0qUfyuvPCWu4+Ibw0itaAW+mK//Cez3TJbxAtNU+VWc3
pBHI1tch6CiXk58NjeTomnAnqDac3K7VXe1euNQDjs4n3ZtsYoHwQnG7kwizGxXt
pZ+eDhui0TqFcXViiV5XxNMNMOUfAr3tKFB+YDwEXVl9D3dZMOppiX1NybQpJblK
Fs/en3tohrD5s/6fN4/s+17A9cxnfchCzkc38y6qoWCmQYj3OxX+pOTcg4Xk/9Zh
f6VsmhWAH4RgnsvGo1p/24bZ0zB/9arABc+LrNu9E1YyLL6v5QNTcETcKrzqa9iE
GR+oRn1gqHFzkKifxWr5niGFFUiDspVBwyxZKcOSHopHnOmDtsDj9a2zt14Jy3xB
A7HyQwGeJs8fMGO8oda7UAqfbTuwkthckf/jBCwlvsMeOODhVPZtiOUs2o5SlhSm
NEdKB9wrLN0yeihZZDppcUbg8bny6yOBNMZHgdCZrXh5Z8S+u/e+/f5ONIbZHCHV
hL/I2EeudefPMk5ki+xIyBgU+a5AdAiHpGBLX56touxjHoc0egOuzU/Uurk8guki
A4KZFMDoAEn1Q1D1PbpB9mYsSnEEJfXWEr6eUGmujuf8V9gmdsM6pw1FzG5jQsVO
ep6QY7RzA/ivWVI955ZiKc65JfZCQ8xU2nKHU9S7DluCXtxbU7HFytYZWZSQNDHb
7qgzHG8D7kcBAnZvP/HRihVVpn+ZDX/2b9338SSG4F8Yvt2z89tXmt9colJlbv7x
C1eSzVuOIq7rq2v+KIEQ2XXONrpryw9Ngzew2+EzmVRc2kXSOSD1GrXOTwWQfxb9
KQc59iRviqAaYRAtPfZ+O4QPjNZVRqd3bcIzlRcE8wlCjwdsgFYGLuA5bMdHjqVo
WGKtt08zayCip9pm90bQxVwX1Ya+wWfgTBPQLWAQ901vnbp+NliQwNRDM5K7I2zp
qfL/Vf/7SMUvjXY6kZUjOda9w9g1KkAMpMELu404SjCQzB0xD5iFv7ryvUbqWdvs
n0SsCfmAPZQXddm5AjqeWuwX4KXTo3IG3oRgDdAQUXz6h8VuVF6deC0im4/nEdI0
3d5WjW4Y0CLxUIl+Bm3E1ednS2QG/WKm7t3F+LIKaYM2JG86rhn+oDdiHoGnPk3W
JcyaQeDGeGU1kPiNeGk4O1FCD8qdQnN64hSJrC1RMUQik+oyZqfAkjEtY8czSnqS
1twYUvA267ywVyOVyl/FZUVeDsqd5/i7ISQ4QY4lfJgToO0FyV8BS+oAxsifrgdo
RgC537RFPX2NZEtwGURTblkerMdVj1M3jA7Ypk4Rvn7VgBMhd1D7lwKiCLgy+Nr2
hfPiDpwc0Il60jrGk+9HPkw0qUfIl1GmE/HUS2JoOL0pTjRpe48J0pXbpyhdID8V
E3K/fGAuUBQiHgMXHxJYi9YugTsvfqjsyS376Bk2xfcdx5PE4GngED2ReXJMICcu
O13tf16+RX2Sw7WWqiEFURS2U4Rv6ZNoihnmVF1sQwqmcmkLWN7i+IToTfJtNu+N
1nQCltjtYUnsaVasnCWNHqHlrQbLFGiZQDQ+gCB8G2VC9f0s9p2Fsho6YRzg8//x
T+HM4X9HjA8gE9ZEZa0u2LpUA5/9coKE59kk8p0H8M2Uz1uEOMcXtjkcWZXxHu5u
aR/OK/50Cic6ZNI4p8UpRp2L8Qjn1kaYCCUTWbGYreVb2X6QoCTjn6Kro4WdVGGQ
1XDwGvWOd/Wr/GiXSWFafwrTY1qlUZustSY3tjC5IOsVjRLP54eO4o8rMZI3wGYY
kXf7pPV3ti2OHMQuCzmKQh+4SyEsl+dT2YC8LM+CdhY1x/nUjPM2m5PLI8KPh/vM
oHWVYD85HbtseoRkaW0XPauTXEY1Zy5WVb6KLEjNPaS+uEy2ZOHINBBCDb8KNdWI
/DNhJQP/ev6umPlDxXOd7rLMrKgE2fK5nFexRAgMbalkGt7XsAkFmGPMhsmkj3v+
m4RmxXuhdiBYQYR9xbqX7hAA/cMcudODL5feFQjxCBwKkeKJzu8foF/nAS80cUw9
1rfsITMSLQiQtvPHDhK5N4k3I91qjpenFN1mCOtGsNccv9dUO6VDpeuAQ5LUwzgr
QnerugcQby62VKU6h8UdkEYkEEPy0DBzsSD9gfUu2TmiB27XzEWPHRXduBJtBf05
dHLWFxHW7Rl1vaJiob5kOpHgjiN5AK05cwH8UZxGwmb5ytCz40fRsTqLHBxS0UZ9
GkRHdF2wZHR1HSFnIiJT+1r+rXt+BsxmMh/vQNMV3sfgx1XGnCmVTveb9q4irIOI
n9g8lDN4Q5mF6vFbRXEWXkrVBqK4yWExLDkFvuGsORX+4y4kOMi01Dg17OkfhZxq
Kbg4HbQJAJJBMWefF5Zzelb1+U3vrgATl62HjHXuq0iydaZdvFenoZhDsroO8g00
chmC4CkVkeHXXz/P5f45+DTLTKhIFt9Yi52KGqPqr/za+XEB4MVSJ9lzClHAr5bg
c2v8T/Kw8/7N6t//rnA6mpPsJGftaXIWNNDu6bl7uoDz7gZRcWwnd6El8IW282KB
KWGRbTMYfAVEIoIwK1lzX7pH8c7S+fSUytgCDPdqFqZL930UrAplU/MKidzRJ8K8
LH4s3tW7ptli5Am5B47IySloDZN57yWRuzjGcYzPeWXf7/jCCnXseyAmloLnh6q/
byGpteuhzNQwFMMD4auHBzHH/g6l3TYfa7zb7JdAPmwEodtv+537BMNF991sPDBF
dVmg+0doSkxHS6YB/9XIgML+ow8n1bhUmpuoZENNDQdTKWLo7mvRmSXp0Nl04SWl
EqAFpv9eW/1z44aHoy96P9qK5zXuCO+gRSVeQyuYi4MU89UIUXZGksaqtHxhAuLR
3X6LxGmcR07zojbGu59ZOg0QLbpjjWQUFljhv8FwvyLwlvLe+UGsy1JSkPGC5wgP
BJFrMT+/7+QTgMMtu3mtRu669HsBNHsHvJKdfUB9Q8AFcU4oVBYD2pMeCw6CBqI2
VbGGxL/zVfu6VlID6Bsu82r/zH11g/59dDDBe/Uwhs5qdZG+MlnemTn8e+TTFA7N
dl95TYP6qZnHXOX4EuXm1sN2r3bLGQzteuxy96NntkfAAnFheh7FZvPbiTiwYygS
dNk6C3YDVtT4g/0qgZ2USs2QrKhA4OrbYjDyqHpLZ1annj4EG6zk/DYGmyk9Fl/k
mfuKNkcf1z8GqtM7rgtfmH5miIKoUGDHMu/wuHyOauCOzaucVa6KSa+8cyEEv3pX
VL+3tyeg0BiuQ5HnVeZATLDSxLgAMcj5dPQuoAu2My5GIhZp2QYizCsme7/UJwdP
I/3f7myOP+Q1iBn2LzDKC/ZdOKViNtm0EOpIC+dKFPbeeAp1Y9mZJHbl3pf5AfVD
L0l6k6sGwwaKGDw9OoqPE6WZBM/yhJvbiYmvFGcpBr8SpnI+kfI7mThhW+wU5hld
Q0+xLfH4iJ9X93UGdTZURR2IogFwuAMh3e0d+c5lVvOilINVo6QLllfLix5lae9X
fcQWxNPjH6EHBZXoBtDe3+fGgNrZx86gIcOcgg8W3sgWP281Ak5WomgU4NS+pcP1
PTviwI3Lk1X5CdHY1N6pVENASICNi5m47kXOBxBuXOJ2+p1++3OowwJjFaV3k+SJ
PuvMIHR9MMefWgCbL4Y4Dqw4uuBefBn4Ih2jSC0hr5IVUhMyqALk0wF/r3xJf8+s
uTHSARg8cZztjBT2/F38cvrjG9UAKyoedjfe2AknTuuQDJ2ENkapSN+QFpugf5rb
x1NUHcGqnskbZQNhb5niATP8upEM3fcQBSIJDiDzUvtG1GH/nPnXsIugcDURhDUV
nNfhnZAGXcI242b7mL2FKr32Kbkz2ZBIT5Sjihlv1VasW3xvAwq6ZJvA819/+M5L
3It7Ue9YuR11qPoInv8957eQSvP+vYJ7JskitU1IQZxnv8jb9zc4/jCL/t4ZKL5B
p6vGd0DaID9W56cRvHf0qZMZ7ZuSbHg5sr5mUzmEDLLkON+nbPsBS7k2auMxwtGr
Ht1gEU+acbkiw430hc6jGVXphU9AAFaiaAC+Qjgv8YZmnXPY4rN4Zoxj6LFClGvZ
KPIuYrR2AvsIHnMo6RAPq3WpYVJ4EKuNPazi+Xa/P4WBCqzuYRenFybdDMdaTMtq
//qq1bXcabHlArBiv3awdns0pgjTRDX6RBJ/Y+gJhunkHraJoiSr5FEkUjl5qFWZ
YSwi3hzmWYs4NcvFKOBCrYDpSR2N5K0fJfNDy+Cc4l2gE6G2IP/8Yp45bOGawIz8
vYi9xugT15JtK0RT2MAGNL8RSkQw5jds12VR6UfJtPh62IY1i+KchF+CO6fWKWon
JlepAkr9gRiqWfPfy0H/g83QRJU5ZOwv8smC/TYvguebVHjlG5YNQnJbIDiuvMsC
N/Ew0hRfAwRyrSzj3rQvcviqG8zx7G76SUAH2Qumt5lWv7IQRz+A1eU8x7jSvMZK
nhRZc+qmH4vtu2hCLkDu0cUytyGIIhvCFg5P/uKrF8xEZ88FTp09QaykJtW6tJqk
i7c01Am8WrM45gFQsnTZ4ETbCqcc/lfHWJi1sSc/8UsIhGNfYo+3y/CC4PzNw88S
9r7ZI+UUTvjMxqsQ3Kt7E2OJnfkLfZUC4+9XP4M3zVzxymZoV0Dwyh67aBiewouH
eXlxrUul3ugKggoK/AYTF9tKsVAMfUeVdjZkmT0YKf7L9W/MaxZX8G+RomKcYw5A
dRj5h+OcZp7wfyCOT/LPDa1FtfvLHQJh2R5Tz9Lt2npG5ydcHJfB4rBQ9GEaYS7V
tyV+RhnA0eA+PijwVULNW7t6YDdLvqApsm23KYqls9bw+iHKZSp8tadZgIeEzXvw
mSXQJptCADwvjIPS9DF3mYofORylXCot/UUKHRkfpEdSFrAyvNB34QvdRDESE4Lr
iDnj43943ne0p+p7zMwYQp/TcldIK65wkoY9aDHRv+V1BtnD0QobNDM+DnGH3c74
04oxAvfeHh4whyabfpy1Eoywa5yIejb0AmD8zeVS4LO47s5jWfnXXtCxsFLOhKVA
e5+7Bv2AtzXpBG59h+t6miMl5A3zH+VRPJBW0Lgd6K3mjFiZWPl/DbL3ud+sNOKV
KsifQ0R/WArVLs+XTiPKYnTac2TAK+axve6A/QTTvz4hXFIOJYxclYSKZMTY0/GP
wIehQCNXQoN3IP7Qg26veREqY5HqfNRKfU04847piCCO0LxsE/5405yJ+JFna96f
byhsiwpu4wIy4rScvr3TG9IrqATH4Kj8tLajysisWlxTAvFk/qiJowqdXHO2F5bm
AT3DiKCxgAc9KZPbxlcQlt9kGe5wDuYkhmC6xZPi84zA0f24C85uuivDdj7feOKb
mufMhdrXawP4J+Es3Kuwkv0YU0iI4PsHlDRX6VQZRRwBbrQ4jg6/0PwieEghqIgr
fMFkN0VkWw/Xlehu3zNdxlqt1hM/4Xs+0IBAaTsFYD1Ckb4MhW098rRHr83hPpTq
hZqC2xRe5xSAiQLLwyjbBF3tUgKlRi8b+7301cdpVNgdbgNbBEhW7MDfo/URLxpI
zvaDb0iBuPi1Flk0+cKpymJAsUcsZBJcbDe7bHHQI5huidGX9oyjY9ZMMN3C/ZqQ
CnJHGvx1myQ3NdyZ88OUeQkT6AvyLJgj7wgZooD04pF+fOkzxw+QBsTV0h9k8CtN
iKUGhM58AlDyIHByEFYwsxXqBAC/BrY5JfExBE6RJJtY1n7chEDy8NL4M/s6qRge
tVBg4qSY8G3hp6BM1mQ9rXdGiA/iaQtymMTtvMy6bDOOF9T5LKfedzhgzoAYfoJK
lPsPBZ9g0zDPSvAuDGpujyjX06T0WkuKPXYSA5eZE7Wa7yMD6r2IOO73RQEPfZm4
jqWfyDbP6+NenpeTH3s5MOPn+GoW0QQG8bhMHfuG0C1zms7+jl+W4t4+G0vzgPH+
P/Bz1x8mLeLB8+GSSWEs7zfz2c2QEXpu7iY6aaI71PXBsheSRfTXDkf/f2T+PArv
M9GJN7bVsmIKMZPL8fTxX7CjCXVXLF2HdCmqHezPyMzhzcpHUMV3EmvopMkiyLjn
wenVWesHFYcy5ZzEYi5P51W/eFxyiEhu61jHT8PkfzmNBN6pLZDZqm7Ca9sb2QX/
SDbu8SiAoTNl99xWyd3QOaQ5yUNg+6Vpbc+dpzmjcT/kkBDqhYkOXHgf6BKz7rr3
E545A7L5P4TmTU9RAyQPbl75NX9dJew1PnND3nsJjxBP5ox5ICES42IAaEZRs3u4
a+N6tpjEZWGuI0MdSnlM8TpXPhegqlRPEWd5y53gAdZmOr1G7dPk78sY5f7hb9GE
wujQPCxyNClairsSkAy3fY/pv0f7lsqDs8TjNLKoy6amU67Abb/wFgcqSMLbMQ4G
i7BjAeUse0Wkg6unBXPnM/ifuBVlBleN+7uolAgpYUYTgSRLlPSulLgAWwuzNa1l
s2MIWrlB22al2AM59vFaEuj1I/iYhYymbwRZ+kTNeITUYF7aw4zddmkalz7EVguH
Um0r0EBWvRYGleYtMpvqEyWL9UgV+W6gpoyx6xm9c6FJYNFTJKY0mVc33n7qBVhc
2+mXHdt6Q8ytclJeXYfCntTrjGARXbBWE62FSzxvpCVLbhkta6aaLa5mNA0dRpHN
xCrBJhjAcMM+p37nLlL9SY1jEwrLkmtnv+kWlfM1AA3F4Xhszn92kvGdDz4zEKwa
GhDLie3p/j5x7rQeqelb8Z/Y58qBQiXnaJ1eTKvF+Ayi/OmLSddncXGcXJP9M/hw
vL/d1c8kn+Spl43iYsb1qTUXucrQdNBsFqO3hEFVHXL+bWnljsQ9VzwBMWbHJ0xG
hPUQ7XmJLyGgk1/NIDvDKkrJLi9ccI1YI2eFuScJ1pmxi126uHH/0YtFNZJT03hX
bTTNOSjJp3On5UvYLpKpNcJN0jyTcLoHBeegKNEwNGR4dP4d5+864CbgCuMOe7Ue
m/MWTcPrrGGTCpfecIxhew/L8C6JzXdqIyOHXSY1AKdlWSIV5NxFGNAovxeCwbCO
X3I/Vg25QibU23pks+fgsL+oMmENegwh1rQNz63UWTwciVtmfbvmUfeg0FmfYLa+
N7iM6allfs6v3trFywoQRbMCZgvFoVegTNsw3pUwHojlUNk0NJDSyCtRgNLqZRhc
zGBUfW71g81iQLhXrfWIOMBYHMmqj7ktgRJ72CWJ9nEiLFB18u9csISfErBm1zz5
C6eCsAGgB60JVLLS3vpyNDicB9lButebnbVeiXehstNjHutAqeK7Bsk+SzG/pvrG
gMgEzYRsEQ9eBV5dIo4+xmKg+GNSVrjVxHzNPfGv1/nHC39DvE/tXDIPMJKTJOKY
EKWNrqsKK8Xw2K4YcNsl/FjijTDWSsy/6eI9c164x53R1FfSA9F6P6DkFsrD3TpE
xA+PqIGjhbu73Imulp+BbPU+mX+x8sYmhWpt855cjm8S7fEcqwZNYOVD3icd89ev
nPaetC+nk2LNP50rim5UwYqlPwKzobxKHm8ep5kL3S8crCE8d8/Jn0YEPgCGFTUr
UILqOXvAMAlult1WpMefAfPp44zT/RAbCZFw6IztSutFaJHmZV8et9LFLCCZP8Is
F3kbe8gZgq4jfaOB8FpqnAjcz6LY2ZTUT2T3N5FMpnZWwD4BmwF0vEcdLxSL+gMy
YEK5gZcYFwxSSI1diyg/yNAy4AKLpmX1Ly8aNs1sQ9paNE0o13U1uIEv0im/3biI
PsMBmfeS6syBqCrApUS0iQFThYipgo6dJRfF7ISwfdeFCKg4AdXZDPwoiQanOqzT
oweeN+wgSY5bNYZqoYJwI1g3I+UUVsuhgk7RaY/TXAKug888f6Shr7hsaFalsmtr
cY05Q5Tnl+MBsLUKG1AYeHvJs7ixGch4GyvwhJuckx08OaV5h61xD9mVYmethCcy
f4BCO3NUxy3X3RDbmyN6ulXNy+bFwBVs3MZt6aaBeT+p/9NaIn25VHboWqNlNrM8
kBZvfDM3ILR+we6Mk5hk5dwVzHqul90a2nXi5KltnPXjhlQbpwfNJVSpjDJRJXr/
zrUvMGiW33rkx6ZU2Gt8sRGR5nVSEIE4KweZ1L060gg/BTrckkEkJCsxkmDOYaq7
jtauUFr/n1gOAb4PElull04kFdm4KAk2nsZN5RIperOGRhXIXpDmpCs0HWZmPyQO
E1vqvSu7mUxA6o2R8S9yHET3UUFMYrlFdpc9OPQSXnJSp/qsZ0mKP1803jkWwWa+
FEJigydCuPbKrVktpeR0nvu3nI+tqmuW1KDMsbY1/cB43xvjmjcgUd/HiRn7m+Pg
itvGJfbicnflqrhS0bqgcsU2ITd+UIQYUB+4DzqZp4iFvq6vDnIaLhvXbjEmC4jO
YyXfr4l/mNLcN5kc4VIXrHS5SE+kkVTj42pr3Wm1LFva+Pr2iVBMzVlSWQeB3nVt
QuFiMhopYUIwYDoPO5SNAEV+UHT18HvWCMZdON7LzUDIK+TOqBrda9GL+DLj7o3N
GhjMOllA9eL9Ag45RrN+FJzIa1jKu1kvN0i4uzoJ4fMQkDVfyPRKBcgE61plfq+9
qxQ3xdmiimTQ2lUVqSPSNimFx4XW3YzY/K0nbMWy4qojAndXbM2oH5GEN1Uo9bbL
fnVdJqtRROVDH4ko3+b6KxhUC3SRmaDbYRBK/cMU97UmxQImfTzl059cLjJL9jbn
L+a4SHE5YwCMEopDeHS2eOpdJmEdjmggaqFPMNWfuYhcgBMLOSEwesw2oa1/56Rf
BSNoK5KtW96+B7wgWL5egLlJMexwBRSf91WgLxRUjy3doDL5LpMk5mmbmkNWECgQ
JU4X+nMUpV/TzM3XIzzR2Tm8VN6UvRIpU+JSAyTFjc/Z0B82YD4ydjET01lTJ6YS
PiiA8IMOtmWSsuzl2HmkRyxBf29SBguiIgDwM9cPzL/knPtJCvKpjgMD7JbHpEXA
6Ao+SINdCFvNp8f+CrngQt9Y4FO5IxcOdLn6ajapag/ZAsjtDWEunNec77tlqjpI
B7xsa1IYIOrkogHTHNy0uvORXDEGlLhjiDbIP5G++3gNgFP+3rQifnt0PMFXbokf
JKhZkWm8SJYP9y+RHYg6p4R/LpQhK8OYJXRE2RCqhKXoRDS9uBqci29MK+Aqww83
kdDf3inM75+sHiCkNxy2Vpzr38H7WjG/JQgHYGZPR385sDrSP7U9HR+ddiqeX6tU
P/5swOEu2mLwCuCMQJse3XsVrv5Fjh5cYXi3gR2O8mheArdezQVIwg471VyqJPrw
vpCfI0JcyDABoVCtxFITUGr3801pq6Xmuk8NxAV5BxcLDlVpZBFUa6mQHDUaoUJc
oHK82QL6ChzyJMOzz7H353SpKkNG8KuvmyYkDLlDtjrR+LPPhuQamyhfgO5G8MXE
LAwGIDE3PX1cQl15+EM/V1fVkCnt9YdsGwgWOJbuXQ5JL/TllTURfaIH2+wDDFBo
w1TEgABoM8ejILufQs7AB2/fvYGYQJTizR6sWaVnANRWhfRczdNUsvo1tD6yLipq
yHoen4jqi92nBL2DZNeTDgXosZRkIN8AvPY5YFw+3EDFPyR08VMSuEFR4yiZeoJc
hvRNCvaSC0sgaXxx0RkM/U77ZZCfO7BxvmyXUwhkgMzFkiNge2DNPOV1M+mHk+ro
h7cyHKHBkJkKsurbw/ChBCw8uRcEw0ak0Qv57xMVeckamM/z1tlrKdtZ/5+NtQy4
iJQTcUj7gWmjHvWERNYe/qMY5Ys0f9KXHMSub/CUIiyLgSYip1XXeXHOms2RPpNh
kFWzmctonhJeFvc05FqY8OHo90eTat4AEowqx0CRZxf6ht2YyusXdDceWzoPBGHx
n4ia3m1uBEBo0spsqd9PtZfrc/YGoVbWUBAlqPDVi8dQAm42qSwGfg+AV1HSppWo
Z3RXJz6vmngbfNHphd1CS1WNbCW62xMul6jCPTuI49Vh7ftXmm/tPKvWA12q9Zct
3lqqk/bpRl9LtKSPhLV/a4whtxevLbEzKXYXwv4v6GMZc4aXjyq/zootiPHUrGmc
FcVsCkhe+insBdWTDoYsRHdU7nzhMb9S8KdN8ajxzenwY82HwYKUAD4NkNufsDWS
iwPYJ4DJtaP3zZG/mWn7PgCzT2sHpxeC2o3Dw+a+gfKOviy8wMl5x6KU4omejiMH
jCoyQk70wkyAQqYw8nNUzUQm9Zc68LACYMV82BKemhtBqvZVX0p/OVSqcnf+HbjI
LLaudORe9/Nd+uRT5hT8e0t1O+CBjyMmb3+XoxLwyj/9sPSzvC7V2OcuAO34NiXo
dbvVUnD69e3BXpUys48/MXr7YQnKrIf/h/9uRgaFNKD5wSFE31Cj7JsDjT6MOITe
aJj6yMF43S+W6xW6ckOjVRwm+Xr3utDl2J24l6VZTmVFTF1i4wgmsoF+y6eH03nR
A+3t1F7ww+s+bO9/Depb+VxjDvKLpe437jDVBdEUBTv30cl2Kpnk7J/MbmvCsc1k
vX02NKv2H2p2l/1GMBJWBuR6XlHT/ajThvNnIVT8bzMczwTpQnhprzbrcbMTL0jF
xF0j1lBGG6cKAjSJpEe81N57a+zMnxXzC6LMcnsasQZXi5LMoGxntppVgB+x10d0
5BgQz2LiaBgJn6BRqMn7JOZuHm9voiSkSTZqx8GZAxQRHjuw2YC/8J2bDVonaJan
I4ooWnm6KUMEqg6wKUvat9abjROEXpKSslNJMkAjBdPpvXoXCylPaoz5uczYMaNS
dc3odrWSmclCTv24oULyYMB9h604g93/qNM7cT1BQ8rLr/WWE5fs850FcBw3dBCe
HmKgg8StWNZ0EZymtLRI4Zw+tkFZqXLMmi3IQVn8IStUiyYXfuDsvvZBuK3BqOmv
oSYnPTUtM73G9N2bmLfIkbk1sRuBAY6B94wrlscFVI6ng/OYowy9uywUZoK3awTH
93H8OUb/V15S5cbeTvj2RFAymvOHE6mMa7TWdVqXxiTbFKcWL60IgVHAVfu2QCrG
XpMdXMuLXFApAL6Nc76ms3gCqc1Y+sPGXJHk5FDQEwgATIxnkLtSFu7wvd4cZ+3U
j0Ky0fTdhucFGgC+8AnPEpRdyipLY0kUBBbslUpFlVabgc06jbfSG1B28LUxiEpo
wCSbIO3F69xbXSaet3RAyMfN+rtRUUpkknDqQRl6VIpBfCXJIMJRcetLa1Bdw9K2
rfdYRSonr7nKbL393cOMPLlGRre/7Kbmsf8ZK/O1/wpDm+IzX4So88D9Ub7G0nS2
w9VJLaQXI2pQaAKfQQ2P7sf8j0rzq6akMXlHRj8IjB9QgmvkyInh8NgZZSILfaN1
E6WdltyaUckd1KCnwci3jW730199P7MLETACOiSqlw7DQvNoVZ5jF1DmqKT+xGUB
kJtnVifsMznoMvuwNjlEVMxLmGRh1Alk+zcuyQXmzprJQrbfyx56bNFgNrGi18Y0
KIhRKgKgekefG+SvLNMSXz7PCOMRq958A9zKltZBaRLrvg6vg44hIYSviuQLVT8h
BQCvBeagUqladMiAHloXG3ZEWtOKQOPgKfpOQgymJoCjDa5IPMR73jzu1UR5Pkqc
qhAvMUoOJJCm0gC/g0ZpzFOjmAxhhMMz+IcheIs886DkOFq4bV8HVlRGd0UTL6+9
AM4DpjEyIfe4QAdmI5eL2RtGRe3WFYtjgH4z7A8q6QW94++ppwMt3GUIzKj5S9JC
ci+0OFOdBok/lw3BCaOHrsfPrd7BPueB77GCRpGqNDuvO/NwK1Ofvv8Q5LU/+gaM
niqEF+fy4+sOhMMzbl9Xc5QqhB9v7JYfvWiqZI9+ItL1M8AyGhCdZ0JdH2IpIs1g
03pV8E1BXHLs4p7MJa8c/hAGcbg0XRNob/YyUfpNuAGpJkhDyWZCh/JbSdLryX5g
1FkeSVE+Ggw+IrPd+/wm+pa01Zx5feKGEykOSuIRcjYrUNGjslU+TA0LsxPPxCA3
NcPrPZZMVWaC+gKr+B1Zwg/kvkMIPZKcrUGVWVevHABsCwAxNA/Gr1QBNkOHEi6E
Rpb6/Q08Rl7csHZZlJa99zlJMaDK9KiATsWRcPKMFutrAX4gorfjwBM9HwuEX18P
5kk46gg7qqyZQ47yDTpd6OECQEinBiMiid7xNvZJNV3tnR+8sOa5rkObXW5s8FNb
QRArvibiRdG8T3XIW1Jv+4P6aPhMs/T+ZcAyylQMAE5y7RdRezzKDkOj+J+mD7Fe
vDyLSColaGVZfNbaJiChya7GT+eoIDv6loDg/rXWZ7RgEscPxFFzkclky4C7GauP
bRTi1fnju6Adp+LDcOZHJbeN5Huzkpkk5bJXWhzR+GLsQ3FsNh6M40QBAdoEgSFI
i49nSPy/ckAcceiVxurrUg6SoFh7m5AqUDnWgZ55X9Nt3x7JwB9YFccTsriz+iJG
OVCKimBsePGD0+HLajcgqU9NQhhMdgzsk4fSIZUdv9w0Ra9LYdFGIbPfiBODvlKZ
wJkBtox0yxiZd/faMl3dfFZRbPOsYbSej6KhTbxow76zYXPDr3eJ1b1+YqXeIV9t
gVD1GPkJh7sbjDJRFX13dVkSbDG3DH+hQ9Hr3/T24QefwZB/pYi85HSKWibUpyCX
8dDG87XR9GKEd+3KxayiMEpFICObq1+piw/5tjz5OVcjWg90ln48UnKGc/2JlQBY
hnxu5GutpOzVZJs4Po9Rs//+zPgL650YTzMnVxE4Ii6V7daNvhwx5Tf0obF08NHm
RGIkGTI1O7wXrTl0errI58uPbCdxIVn7ZUbAvDjREQsEmk/HxHecCZdKev/xIJq0
uE2r5sLZzOvaLhuQk3g708RgOda2lP8qt51KCvMRK3HO8LBHcSXOA5S4AkrYEhea
vHNT0eATf/eQo8ODPjGR+GrR9568sn+qfK41ptA85dvbu+d6er4WQ4oLOV7B3GC3
Gc1eCTF6+vRQWt4fOFuwAIfH2h7payjAKMCKCialpHwFWq63tac5t/S8LnQMB8B3
FmLz8MTGwtmkd6jjXuOak7eY9HFPBoawF9qo1JwoUYwRnwZ9HXIJBIzSFBNibpL6
lLpecFVvveQ+zyH6q3wsfKctZMsQvXEp7xG9sXeWpUiXcbuPHhuzo+QYz6PxzP1X
darkJBdCUaFd3Qm3nJz9rkdVAp6j/rF1WkwrR4RdVlnyn9AX5OuYJjNMc9t7q2I5
OA45n7CcIZSIAKeLPLNLAelXG+CgYgssBg6yA/1uzklEk28XfqysnxpyCeOfRVYM
FrX4neYpyVCNYo86fzobar7ArSaVQzrc+SVoDBYpBXHmnTTJGa+Zb86p/x+fvhdJ
fIJ22UheWUn/Wtf8++GaLDK96kKrnBkBahYYq4E50tKjuJfPB6vlvOMzPE9IM6jU
14jRD9RUcPDjE2UmGZzmKFlbPJY5e5IHxWBIlpsI3r3ufbd+ElMdze+tyal1daQ6
OXXpodolMn2a25V/+ZiWPVUDUCO8vwNDezDE+xcB9IltrpGdUeSYfoqWiJcpP3XG
XU5AfuV3FrReh81LL5YhuiKBfFKxLLYlvRoCpX0qG3aSkWeCnyjEY6PlxV6qG55e
4WyJsYjf3rsD6ALKAiuNdWES5hjKCDe6hipGzdgzh1Da5nYAQjVy+fcQhjEFni7k
MRawEtDGAMut5d6dpVSeMobwfvEL2Wesd9XnkI0GsRh3vtS3lPobYxbOgYYuIgZl
XG/cIAYwiYr01RNCCZLSrBLu386HvWn/RLiBQQNdp5PNSBhl5uL34+YbxUnn+CKC
Fr37uY8kWfU13cMP8gCZriZ0zoxh0NAzCzqARuu0T1XlLhtHPWXAL3+lT7wcWizK
4585DaT9qhDLwwoFpmnBUkBKqgmKx8NtisLTUlXgswLRJwlpPAkYGZ5+3CkkVxR+
dH7ZXdR2QcTtfFyUzZtqk0ws3mMKeli3VR0/iMRw+B221l0fFTV6syNmUfWE6o2X
ywuC9iHqfElX4wtH85Ht/K/Vg+egZb1phdVXXI8mA84cyZgxxvZxo5a+a20/izhQ
TwpUQZtbKpPgiRHwHKZJeHh06uNhm8KJaPfnEySeCFGToD92BCzAyFlxhIAy0s9W
SCuDO2oKCtUgiXZZmPQDVsuhjvAXfVFs1r0k7Fjn+qrQSZzLClLGO8EpuHjYCfM8
yphjvWvHocVuDT9K9wcaNrCJAZAzmddfqeNHQMQ9re8C0dzyetgj2LDI3m/28E7H
kXS5bmwnufbgxJKaKgVHEKfWHSR1Dg0Z7hk2sFH8ll09kCQkB+z+lNp+t57Klu2U
hueFc64buthGP1Gdh0ROW45inpad7UGh+ntOh//M+L4qoBntti3G0p+JPxbeghze
5+s2QedRdtt4QugIRN7EydpLco5sP3bH6IKg7w7LT1O/Saktk2/msCwd6p2bhgdl
HqVD7THckYh4fvkgV0ZGmbiD+zElbJTKO5AV0pFTQkHKNynU0UkRKh8xPChYav75
rp1A+Y0UMLjgj3Cb89dIDEFHElHKpP6MzDDysiApqh2SDlESO6yiSgNWb0rxGFzr
jePaRjlZHHresIYM6u7y07v4YCK0gIIbG50ZxR7y2OMdN9uWMkFCmttfEyOFB59D
ImY3Q9pdLZCGyLK1m1XUVxiOZSAYznpdwBXpDKe2RVBA8aEvPsQG8JY9fdew8bkZ
mhX0B05x3EwdOus6MciT99zJBJ3k9Nj2NBP2FuPmbPahNrwuYyMaNAg+G919eNHL
KplMr+TCgNVtsMCFZi4W8f9zIQrtEF3IGdDP0Iq3MO0fwEQ80AsRfG4hHNEHJsUk
JQrUXibipbHrPrr/9v2oEaHSUEUQNQ7lWAPyvEHv1soLeELjPtqlYieJst6FOusc
5RdlitLF180D9EeH8eheS4n6pMckvchiWpqsnLiI7AcWx1Paf80MATwxDkivcSeJ
JT3LUl7ax4ZSLKL3/IiJR/tl3oFG8JNnjXuKxYEQTBxZ4gUmhCO+4O1UsU+LuYZo
drFcwTbLjLe9dup2zm0lUNDFqlcRuetFitpIDXIUmOWJinz8s1dMndlYM/SS5stp
JiFqFB87y0QX7ykUwotpE7G0M0DemdkJaTClDDd+FdbD+O0Ualczkar0FOCAItvu
nks/Iyp0Cd7SOCMKGbezvLvDX43YbLXVJwC4QfVNCzWUQJBRWOR8dW+o6lCA8igz
IdwzBBfMLfySnQLPIrrAEJHZ6ctRrL9h2dK7CAQXuO8UJEsPdHN4/B0L8qosks6C
/vtk12D7FccsoRfYh+VEB2F91i5Tp3xHa2bqtaxzRnrHPf28Sy9Ga7J7PNPQXd70
HCOJcahYr7R60ZwxRoS1yt0ki+Vq293x3HMGwG9jau1arfQzd68eQIriXZe3mBlI
GYSpXLawRnX2SucFshde+iRnwnLvu3pD6CmEUIpHQIL9Xa7vLM8kWjoMQ6xOwy8e
t/5H+p/SinyYseNtb9mL+qqqIjIL9KulERdOTuPo/IXdXF2zu7hZMt86OMiBo4pM
FlRF/LVrp0uAAH6gEWIhE7fN22ioTpq1oqExPq99oKRv9uJwnJnDaTgx3v22DcfF
gHvDerBr7+1RXSHO9Gh0CS5UDTXgPtJ/J6S3E4lkEJnhFLFnqWDXz+xCce+WfIDz
NxP9/WhSJtrPbIPatTjGAxJK20i5MlHs0u7j5Gca0ewRApVxf6GJwAN6bmx1xW/i
OUFoMEWEQmN0iDeaOCFGqWqPSPtd/TZBKqiNSDveRhG0tFEMWbylEzEiYMS9Cj+i
25tVwHQmNcIvXTEcSBDMtR8afeqDIZZ8lCa6zJuqjpn/wgk0TSNT+rwn75oE4geR
vPU7pXOkKYAPOx3RkIhN3zVI5oqVr0xgtxfPeHxl7cf4SnTbfP8K917Awit7R6pS
Gba180NkJSDhkFuqFGjdfwSV86HlJwxKvVYF9Y5ZHWbvll5Tpa5TTYe5nBMOM6X6
Pf93HH5q0Fps1Ig41UrX5C9ok03bmrXmGJ9BNrR15soQcbrSAVnPLapTd9PrbRK9
pMxbaKso80gAs5XLl3Hchn6cfvsRAxC6Cf8RKr5KYOGXGlsEwjbfEwVzZH0l4xO5
/Q8LsCq3RhpMUccr01t3n4DwDHfO1RzDagoExMb4aL9OPCSp2vxoZ/bmIFZOLXLB
kAp0nfmGsOvnSCQUzEvblhDFnjFUU9XeE/BQPCQl82D67Z8/35Is3ChLNLxN3a8G
78EzmSmXc0PW4IKjk6jWn58mbytB9PSKBjcxzJwIsfYNL0VSCw5vH1pDwM4ytkk+
+dZNu/QuSCMXJG3Oaw63UqLAh71IICWw1ZjK6bJiuiGE4tjgCUUOdxOnzjLF5AZJ
AonWeEYEjU0wnnaog3JbB0g4Av6mb+in62cfTfJAbNIxDBR7GIKJAKb0lmvnmYCf
gyEIJO3mpSuBIiJKz0cy81Qd/nUS3YBEz9TBBNcaZrwxWrbEl9/X1bGpdsN1SKkY
Z7XqkwAlHylCZ+yZEuJYC0PMd4Z5ImmLjFMcxQjS90FIiVHrNgdpIuJnnbjG6SuV
zTX7uzlZwCaV970VGLPx5RC5WdZgEHG4Iv7Hmu+0CuLjkZbC/kvjljemeRaEZ4lw
U0uLI29ffm+n9mJ0DoqA3+3bRWNh3Qn6sSgpJcUFd2/w66oJmdTk5ex7h1JCypzW
Y0G/o8c7ETWFQ6jT9yiM/Y/8QnMoTvHYjBvoXNLtj5lqr1jdNlpp6K26KRyQFVOC
2/toYtOyeagpEP8Dv18AQU/1YmVwktvAy767O3Sa99xgqxIAKBv3CwAdxfumg2HC
5BxCW84vSa62+c2p7Dul1tk0nETw10SuOW4RrjHJumN/UOo+3bl91FlsjOv+DnVJ
cF2I5bHt1lKjzuGDlKLzCUmTcFU7PZCyVzrjoFFW+AsvCYqbP36UHZaAKUBc7tu3
jWOgwg744HLKodnp3q6/14+gym4a/Lrp7502QLJVHnwbrwXGUc6Z/m8B4fsptiLu
7sYnwPni+RgExTeVNbn5C6LgEqeRAiCPqNYcIRUwKUuWKwhfTKx0rdVOVtc05+3T
482BiwAzXr4qfT9+tM64e2pnxYzrWvlyEO3lbhKL64PKEdUc8hz8+4gaC6KNkyGl
CTMmQWHcIJA9tis+HcpOKf82tiVYZk48S+QsNEahwYAxsfH2TdksS6TkGqLIIRjV
kNEy2SxtPT9nVmbi5bWAw8Jo4+yx46SW6oa7u/1UBwCXkorIVXdGt60HBvWQ7lX2
LiuEJfxC+3TDMCbMDywfu9S9alD2YmOlBwFD9FzsLmwasXoEtlU5MotI4d6ar4R2
JtkraDC3TTdjgFLpwbURaYMUs+sl98MAs8Yj4CBbWTLVRZ7ARmVJ18R5YXg8vopp
RonEFFfCSOONMuNA9/2hYceWrqu7PxPTwQ+AAr8uSGDvfLKll/xzvN7jgR1a/CND
MhsRUu9qqqYVXWZRsm6s1JcOUDxIjXRWxyGHs6VXrJJ/0hxh1ZYJGTJeS00Np/Cy
aX4Ao4GxO1lpg+FIgfaQ/OcQFHGB8cp3VxrlZFhoy0IyCXscUF2nInJrYn6xdgfm
7By1Xz8DNrxhrb8AjuMxK3lvsFPPNtH5Z732MII9rVoP1MUiQPPH2U8i8EYio4tk
FXIuvp51fm+Of/Kj7fXn2AqEEe4U6yVLqhwVvmZ2Y3ibFIsS+fDSy6qVipWepPWO
F53dnrNhCu/hybWphDv9nGT84P3ii9LM4RyBqeRtBRpCeZlDmo7JirrHN1MYmowb
FY6gAvHwlNyXLQJFCCDPmu7mbU3uHnKt+hwrkldwlEFxy/BVhn8opUd2wpuWyCSo
+/PyuSkUijoJpe+onryrwDkhI0lr/6y0G7+HE40OFGztPuyirVsxdfXVfTjqEcrW
hhfJC7jtSEBXech+bLEAeSzFLAmwD5W9nNPN1smZIepHfKbz920I/dBFxS4SuB/Q
ZAfk7IsRgd7bEhidhpmHPNQajjWlPoxiYq6Yp0Z9YS57pgGWdTAFbPbS2gFmRQhX
yHwwcjTFVc3eggeUC/2NXQKANIDlY7KGcT+8RZP0Kk1LL/uSX1eeSXEImD9VG2EL
SmiB9fRpPErNBe2S3n1xHf6ZRPVHyCjBdOafobxeOrrCBr9qYAWDpLcEYPPgFVGc
QfHsXCSLgqMkZeHk/rlOPS9PixpZFZIb4sQ5gqMRPUIk9kjw9noiurQ3zV2mpuUQ
34AS9KztsD5LPAxe6e3TDFZ6oRnURY/dL6x32tCw+lJidNOMyFlzd0A1KFLSXeXE
hLNv9PwLPq9gUU2VVXTYsNFejhRyj7KXPBTF1v0yKexYc92uJRzMjdpHbJBq5cGh
4SDLHEClDnbP6AGP6vNT0WsuU8VnUw6eyekLITtRu2OOb61jsVVznS8jy0n/791p
rHvXxSH94i/lLfUPeqlxOA1SYJy9GbSLbyhd82Mt7BDqFlfo2ReQRi/bgdQgOSoq
j2aTWthRDxdCwhVMNxeOSnerXnQsCnfpIZpYtGCe/otpndO3WxUigBQ3Wf9OITj0
c1YRurqM3l4KrUeGsnTJcoKAbckoy27fD95gWE13UeR4GjRVEphT47i1fJ99tkAl
/o1Bk/4THbjIoj+G/HI74BUEIuB8f/GnHyzro/1M6aQ30joZI28f+HGRu5AXb1d7
Hru0v59IpVZ4FAIZILgDItdOZDDdufOZy68dcvlQA0DLC8WAcI+tzDcrWzetvHQf
uhmGQvEXqfRG7Jhmlx/mQDgt/ugc5KNsWOFDDOWMfI7BMf7xuRaqB8MS6PJBvkOZ
Wo60GM1MqJx6EKPXs84UrQq7sQtq9DWrk9Izr3XIxxp8TJmvsdRqWKl81Btp4Jno
HKYmbLrX8h1HJnZsGcygUGfGM0zIQ6k73kUZ96WwlnCPkqc3ssyMlyU/b/kOBp0j
5y10ikOJJ+DN0dUZUwap0OX+FPk9gUcsWYUNa+OpgfrT8NLwUKvBlNHd50X3IGEY
Dqt9YyMo1Cxv8WsBmnbyMaG/qyVuYR9HSw23nUc8ZZuqvGQYZT+UIYRkEAm+3Svt
NC/W6zM8d2oSN6z2qNRRJoQ6VlMgs7h9HelmPygEIDBfNNYbsRsDOSG4dkyfGDHz
J1R2cDzPKiSFyB4y5tCqVDpgWREDoDkl27wE2hg1lUg0ehrUvykBjEn88H3du5U8
6XQ7fmB1NeZ2mFDDEjWByQuC7VEjg3+m22ukOaK/8M71nVWJbB4N+Z1o7RV8PUyz
kPQ62ZyMnOgGx4ordPoUQYS261LLZCAe13IXS0UurKetJUItEn+Rji8Sq9TspHg/
g/awdNLfhIr7LrawwsNx5oZj9xUucLgWK1L2io+562QsyzRzF97bEfusCCr1r5G8
oOW59PiGGEg2oaAbBRhk1Az6naZiCWX3iK09Wu1sBMa4w4f3u6tb/UbCQVU18hVE
nmgx3COc+N296E83x/XqTmEpCndj/udG/qtdMwSEM5XLI6i5kPyAI/pi3jVpZEHs
nbuhFa1wamHjdKyCfzX4IOlY66/0qqv1DXOAYAjbHORZPM2jSD8Dr6SSCIaPZLZ9
OLd/CtjIZVUOtzpQr96DgubKsG+I1LEbZN2qs4KsHligsW+ogPHa2ZILgELU2ng8
j31kdFSgorkrJh5mw9AY67r1VZFvInrJ+mzs1j4mbNGsZtmnRcWj7QViM/qXHW1w
g8wcqe3WLYRast1q3yaHqGkzWc3OoKFDPVm9NL5Uphzn6sNJKGyNSl/bTyf7eHAN
JZ13d48QjSy4foiZcvVeMfm2hoROQ3cEymOdiZlgquO6Df8ewyGduF99SmrO2Qny
a5qkobxeJX6be44mRV+Gay84i14CeK+SAu9X68eGvic8qOY0s3B7XxIUmsHCeX79
ac0qyZs2faMyBcEAkjwpE3GBeu+wL3yuuw4tkOlUNt3N5/pscNmwb6xTPypfMY3w
f1z/4n7ms0UyJGPEuN5hGl4BOS4myKpfnLOiQ+70mY3M37czHJ7Xyjo9ovlDa4+O
akCOPevOkRVhcihvcnCfspR8xYcC4oyr9XGvUOLIr9zk0wYn3sJFtbMWAy1RmTI0
cSBJhBGVlDnrWks1Iou+vEc51+iH3TpbYpYqwF/pBuW7kIZLoj0HyxBsV2LtQMB5
JQrrafGf2MqWCPjPiEw0irSkfW1CdWRZwdwaIHzN8KxvjCJeiBuMRs7jGPCRpI7j
bKHTU0fhQFt+nZ7+i2nfhl+2OVtPnfUPAiH2oNiw/Fs7lCxzjnazqN6m/jJ4G14B
wacd4XPb9REOyIaIQ00mVJPZdoy6GolV/pOIwPSmjmOTqirdA1v16fryVAF6VSFm
BO0gEHo4Rq6NOLfdaoF2Q2IFO3vVHDCFYef2STBrpve9SkcTQZIkVdo3j1DfgZ0x
+aBCTTZo29Xp8/spE55rLKmcfFA4hvzX9uz4C1sHuJrxugPk3gJDH6vCDXovdWkl
MFpXSYYS4QN13kzs2Fb6qvpYQsM0r1gHTgbblUtf/A/R6iavusKAfZ10XOENG1wn
ftDhjSECGhZGvLDUXhJsgoJ4o/fBupPdNYq9Ntz4zolEdcbV6dHvZ8SdjU3ssv5P
7eknIYi2KOeb83oHA3iJirXeKMN9n1i8bwusX0C4D11peNyVak9ze3FTOP6tIgKN
ocO4G0VuxaKWn/YuAMFUHanWmDRAjI1DP1OmyzVOXdXQBcfIRE71Q+9PtiyZIQTw
eCsRo10KSM2uUCSG+TkpftLBc9h0+b+P92ZS4VrORhpYphRR8O/PIVS2oiqAQa/f
n181QKtdPmLRNfVinN0x1gLWS1Mhs1ylUVLdEuD+xPAkJ/M9oyA/A8nDIOI6I5sc
bAdEsTZh5rpxcG/bzA1hSY3xbMqn8ao+4NNmPE0KA+lFZ5U8r36AzMqG0LGeWdIs
blv1RMp+aUJxd3WPiZH8jJ7fOku0+Yds2sXUvEvBne8PQ7lN6URcLhMnhzQN8Xxq
bCdkF8KkBhzeBUJblnFJ5A1wLVfpH3IMfDecc8VD4+m8OHb7Ns7USEWdidCv0Fs5
idqrj7gfAJMzuH+6TPdrbnNrPTXqqsRcbxcWDnl1/uJY1unKXyVmoB5VrAwImkQD
qI5hSnzVJKb28Mc0spLSg0Sv6fwhGG7PbyaE8GxeBY89/FAMrlMWnTaz3yiZsjHS
ZO72AWQ6xDpBuqHPKZs5XvvmssxSbjKPfVaXacPynKNmtlLmx9VVASDv53oxker3
2gMmFUdsaAgcVSVI3Fhd43d9uP4SfVRgZuxYgPJFOwXzrwXqGaoBq+Hsk2ii9JR6
no7dz8yxnXejq1xnGGjcGlOU4YNQahjBpRoZ5HOgpwWrr4EUqaHOdEfoMkXXAEjh
xjgdiDA+X+7ovIdqiO54aV/rifYAFvXMJt3+mbwqtUfdcYqN/o3HUVMR0NKc/Ew6
9jC+OnMOCD4i2CdA9zmnbsYIXjlmkprUv0xitpgIvaz9RqKiGOzhUQEmxzooBuuP
Qqi5valsZqX31RMd96ti4zMlTFDG03pw5T3sWdndcSeAwjiInVHUPwAMeS/BDZ/R
ODiTNsMiM52nuaPn3O1beBFXHXMI2G4PBK2ayyDFWtzfzb1UJNKXlVYIF6acf3Ca
wzw9LXn9En+yolpBNAOiy0LmvDcpvtzIG9BUBVY1BtCGT/M7JMrHs6xmhO/tdOc5
G2cWqRPt0HWj6B1S5X6oE1I7sMC4D3h+6fRhS7PS9t/wxfv3ah4n1nF7sIkBhWnX
ELMX2SgwmKsWzDT8Y51C9Naw7TMjgMKd816U0URTlNQSCcf6RCwHa8SKn2PG84MK
0t4o1HlGspdFJyT+b4bPwIT+255Q8nj2kriCACp16tUwTxgyTbj+Ojhol1Peizvy
seHggnoERgTpHMX8NFGXC8IZmOa8alzEbsj9yGNIjwuhVzjoXTfhpNuBmJiZCaNU
Btbwp6jasy+4EAs7zbTGxQUfr/7N7LaDP6BWPEbmDONKcD/uGGJthUNiC0aGjVek
DhC6Wz0Y5KwCv1Uo6sBIbZeRoEuDqHcwMQSqLb+Lnuqzg8MI3Ws9flBM5Mp8x/yb
blgAXJNf0ogW2Wru34D+4ivEGYmoFtBtafLUCzVJzVWeVrAacZKT48w8pEG8rCGu
dqXqi3kdbPFPiq8o6R4GXQkQlAGPYQSD4leJE+Xzg2YXzQivcKUYDCZRJTgKr/Sg
iCqUWX2tJp/jfQ6+FBHe1KXjGn4sROIdeipuy1lYXgQkzHuslOp/bqTamL7/dxvk
7LBN+PQxf1akqsevi/U/FNsR0Nz9ai+/O69OEAk9U3ulgf76CJyKhFo53GEamqsG
HAJXB6h9Iwl6wnA+Ha+RkaTx4YCJgSDZSQjiBwyFLkYTJnz3stmdKYgQSWDs+ytL
yd1QN1xYTzXJP7lJcoEWjCTxlXMYCkTv0FLr0UDm6c4j9/OGNIR6y5hG6Aq360yy
vgX0kQxEJ7ljMy1+P48z/UkdLpytoBls33pEk+2rHsUzkYtZQ+I1A4H3v7UsgnBT
bmi7Q+qT1UtAoBtjgAHssqT8S7ftDiYaVQ65QvzZbzpZ7lfUXXEi8URrElnu5NLp
Om/GNSZWjSzlawW7iVF+liKet0M6G0V7h2rhlnSacQTBZRLMqOs2UTyh+ZoYKINC
v26/fTw7oHwjmOiEOmqLuBJOL2JLRFFcxQ4V2RyarwRmLBFDYZCuBoQ4qF+RDi68
PA//wp73g0jEz1zawwXlDHmqAe3WHQTYgYKHyEG+4Inr4V6II5sH8jrKkrHIXDhU
vSVmfArnBhon09MOWgjtrJWz1zXtjl0H2DXzYO6a62iAf5cz/0r1JM40XGIb/ULY
w/QV+FNkU6G3XNM6XwarcRnyPELROoOOWarm8HL33bzhcD7bJjNs/SckASDZEtsP
2S5iIyvQ4HpLmSE7dQm1TSIgYbV/FRu5VIMXhRENvXdYbEUH5L1fqsvHK6j5qRDi
HPrf0mXiCzHN/Ulb9fU1Bl5aDsEEKXWuI6ikNERp8tzqz0GISCed3SSJMP9BALSe
r6ogKjCzhnCajy2Uzs5YntnZZ359lD9IRSdeWtiaPz9b8tsflE/pRgISNmnh583l
WDgyr4OK7yTvifH4Gz637NZE2qF9OIq94SuCdbJUOpUHAcx90Fi3IGmAH+nDrlRu
YU+Mw60Cb6fT5tRcUXCPaLN7NL+zd8OW7t+V83+19blj1I+1uXb2gVOeBxQdmaUo
imJfyWxoh5TNNnZJjhOvIwNEtmjgtSn2bB8CL9K64aNj7RV5dv3bFakZC5m6KpCF
IG3XYKuOtysdumsgbuQCy7RIExDGFmaZiqWKTML+bsn+RSp/iTv5nbLNaA3VYtwz
oR7C5vwN1y12aaK/DPHH2i5M26ha6zGj5vHheG6NxpdXfHwy0xhuaZ+U5vcl5GMC
M4jMmvRQNHO65+9pxj8ncWFHN5SNP7rNW9nfCLyQc6GijXzYQQDcjq4YZSTl/lSz
vyWQMMJAtf7gxREHFGhjFpllJOBlKwxv30QczhgJiXp6TLuyTUgBhpq0+aR36aQp
HVyB0jHOzj1sT+nG8lrreWlaiJTKvGc8I5kkiLiy7luUCWicKILtQ8dgg3hkb+4L
gU4DwToucMcPQSoHQPFILCako+1SHuk0gKtxz1OxmAJlMVNZzwmB06ybjs1AEtJ+
GdD8XYq3fg1C8F2zgc+NU6AJcXCue70Ufdad/jf2XRpSpQq45pdsVeKBufzhrazw
Ds6TW3wWdo0Qefngtcm73VZuPGmRi9LzeqqXiTY0uNf2Z4HA7bIPu+Z4GwO13y+F
SmWZuNFGGwvBw1mMHIhHQ/61YcxtaziuIZHqUDWov29QZ5KO7MntnZ+4vQmU2h9A
GF/TpW1UHKEBKizFB85A6Ty1EQTLMwOViU9ZybYsjFNiqEs5WDEkzo9ehPxh7Dcc
KzmOAsFzXTIRfnA2Lzya94gx7o1JnafiR4ISbVkPCQWpQkckaDbvCCrw3/fGYvPE
feVvH44VLZQwpwgEO11ygCEVcNeEqDeEGdo017s2Vy2aSlVdOgSqofSSYLy3OoHq
JERORwwM1Ea72nuyXHeluWmkH2QYSf47LTBOjrc0cgf7cLztXbmzW53UbtdYe2RS
mbuw5TsXf++G+5IzPI7rxbHJtSUM3HXfivlOsHEOupBRNfO0/D3yYMuIWtk+2F/+
Y/rEgUMXpKVxT5BmMyL2ezinhRcbPJN12zog9DHJfEEIUnMt1xA0A6l8rvPQIS7c
hnVOc1pVu5QU+ASrWb2Ty2FPZ3Iflwd7uUEeYvtHUdKT5q/SyfRBgX1EpPfn8FJn
ltSg7t4Cd7QOwrhLW0lW7rLsd7k0utqrzdUTGW9y0dSHd/E5Al0k4YiCDIKRFZPk
jot6q/NDnhkpNxULyFgWW40+S6SwSxfh8g11zo93MlsofkNIKJdA2v9vm66HIsSz
9x8yOh7aOfW2KkVo51coNuyEcsSWjA1g8CuZB/kPBG0md9kpq6iFiClhC60YCV9V
83J++N1suDQXuT+1qOkrwLRgaKCtH+OrlY4XFrjj+9Fvf+oWDCSa6OCDyXNdJlSH
03LvMBztrEgjY/AVeUafQ8+UUlN8Toc/xyW8HTm5FeYknXv16lLAtTTs/PRY+zsU
wkgnI7Vba4GCKl6co3CpUFwbuQlXFqmTumBZSdeyn3NiY7Zw135KQRSOuKScMgbk
CNRe2HQxbLS9STnDUTEdiQfMom6cza9GWj9/yHk8EMNdfWyMzemP4FzHVgVWsHqV
riwiN1rZwgrD7C5HgyjlQ+DYgHafoGQigE65CHYNTbfnyqr6xPSyl2j2nTL7g1lm
YzIXTdEtHSXO9TEb54F8bgLdAen9RZcKhOqLbgiBNnOffb7Iv6WJKYGCwHMm6T3G
T67WqfQ/Lh1yQm0VNI1Ly/mAMXh1sWwgn0nauvnwMVbMPS5xaHJA3LieO1kUR8c+
tti5U84PU4bm8OUoU2S9w2um/eRFHAf+JXvRzXSsl0nUrFuo8DXFiVy+q4AVIDMw
ordy+Rg4k5J32C5cbL/Vt2lt1e0lwhXY1Dr5VX1/5g3uaNQeUm11rwfYVNw+SZ31
8E5FUOyDGU1giBz+T56E6Hnr7SnqrU75rEPaHQXr+eqjXITZKvf7+zl/4d6lFKT0
3hWhJxrYOUMU3MZGYN+KR4dKvpjAKRhnnvhJSGOzmWkyHz4v0GLnxR4NZrIeS9Nd
l57Um9SuNMTod3kharQBHu51H3qba3kbFZOdjrQa2up8eAvG5/9dm5Be+NTm37dH
HmxQ+buTjvnxhaaj77J0sY35Kr3lc3t12hu0AsF1YdzrWqywZSy3Rt03Cx/00eUX
kwcbhrwzD1BJybKQgxGxOhRufnfIjN94FvBvIfqyqLEya+gCC2/dintVQehowa87
RIE+1mSzVeRPFv4A/YqmrKpuZFygZjYQDTnA0r58xvNTTWKq88q1oA05U2KUclvg
KvejdEJ7Q8y+PcWvTFkNoI8KtrrjzgnWNBOoXCcnRMYAJPIEXJQuw+03kqMwkHSI
ITS9IMtNe3WYLB6BJnH02v5zf3//288o6GoWovle1rzlQLr2iWu8ed3xPnL4FLHa
KKiHaWE4nuviyTdJPGPp4bXeEK/WgYmn4mrFgX/KcUz1QuxX9L7cJd5rT1iRz2Kc
eswxiikqVvlmoOc1DSRdyssTLI3eARjIY9DMLyHDyfpVuYYeLV6naOQlsxSgibJX
ge5SycO66zv2/RU/wCinHialmqy1cnSTwDoU72k6B6yqujqvxnR8AmtYsPK0L8i9
xucMKxGxpO4XA4WhTtJzJcTYXbDQ8U9ywkl0lFxUb+DZ8k0YxxHRFTF4fBkfX6dt
QOQ9GyuwMMQD6ijcpBR2vuAtU+pq3/FIcsZDjwuHTVb6Y5LkviP4sFhnjk7Xlvr6
2P7lMpTL+RaSpwQfFAhi84fZFQFZzuC58vOR2o4mo461YQQ+QBBdXnFhOSazmLLN
8gYMRCcANYpYVA3RyhBwy/atsUdttbdOfajZIXDo4KDhkNivIvl56fJnuLQceX2i
Nuaa8jF+AH7L3XH3vU2U8wAA7lIrEjRfsP12mI9YZ5/MukweynLGyHbznQOaY/wI
HBpd3oBnTgpPk4lRAv9JifMEWxmVNEZdNZegIGhLP4Sw0LDbE/TdraTjCOvpjJtj
O9DJsu5DTpf5AD3Iszxx7BkcLNU3qtk0kn+Pa35maBwSGjGbHEjQTwT2I8QlfGim
rwfdgMnqkcjrhmEQOt50DO4ernIKeEJQ3V6slAFziMpCzVnWU8bIbwewyX/Vg90Q
8EnPIP0o2wy6OSPx0A7Pjrp373JUbuO9bQnVUQixeUA3Bny3RzuDJuHsA6eJhq69
by/gQrHzYiyn48kodKmn0YmufvbgeDlEPAHCV4E/6JS70JQGyCx6qpjrGPmiUa5Y
Be8tXvwtBbP8BULCjoGfnTmt9xEDQa0jMAHb6wLaxs9WmvrqKofDae1+9lwxpbl7
Qzod+W5rzEXYZq4XFf3YHfUQ9AodhfMiQ7BCqO9Ivclt32R62olTAnu4UTX13YTz
S8D9Uyaw7mwUZgak/6AnMdlR3Rp3fRvmDxbqVcyPMdUfGEGvzjS0vRjf/DUoJad6
GIZEdUeVRcDL862bGcY7X/80tveaFLkfuuAsB++hnuzITkgGX3D0/enKxGGe9Pzn
zuzK7rtB2uCeVCff/HfkmCCDC7CJcfdeRgIVc2Pn5/qqHwWfCAr0ekY9WDKrsd1Y
Xr/oAJo8Qb3foS+WHat3z4lo6W6Sbgqv1GUS9DXE71kAiinypsiur2JbCivm5V0r
CldajzXQ088XHGLGPX1nRM3WkTG8ITNwax0K0T6F0V/6pXtkJ9CWVmhakGjUTcAQ
jkBxu5QBefv2yQtw775KB0fSkTdbeYYJ8QYSblMysoo+CSR2gGepHNsbMHooeLLe
2HVD1yG5cuI60CEMQxHVFvHU4qpdsvzUcaV2SHH8Eve2RDxvaXaouUWR4gdqOqoU
bFJ7detk3V2wLIB+QlusgQC5clSoBj8L+4CFYA0Yl54lMn/ixU4rodoZW5vKe9v8
Q9tufm2hWQvTUaPhgROAQUeB2YNevptacBnvwFL3FTmE89oH9uGL+YAKlK4m/ODr
9f3Z5WWjgkuDeyEnnFNesMeH/1/+nuyvMDcnHvqHWZUk8Kp05hGAmnCnGs8Gk/SI
ms9vAdGQXhZwjkhhru42Wy9rjMres6py/oFqltqdnk3uk1JSB2cMvEUCQ1EDhbD1
Hjk1h7+bGgLtOVBTLhnCHla5xtV4FVuF9rR075tZtUwomB+8Bh5Kzi9sC3OSNCkP
Ak6p57ltZ//Pk2mtQdOB5RwaN0lblwXBOSEH6bpHYJEd0vmyX7cTIHrtJ61Ont7t
78xMK2va7EralVZl3eH/EYQ2ChknsbBtiuBePEnxJmWbAGJXw0pKSitVyQcFQc2N
wlj9Hn4I4nkjF2NG/07Ovg1l6hF2wY+OopdWAVAAmajdGq/J38Xiqk5LzbCon//U
FSD8weU2xeV+q4RW3N9XFfqLCR4h26URVOvQHFe/GwO++Srad0+md5g+72t1/GC1
wW2339CGch4bWmgIGdi+vqswoMJByoFxT0Tpsbj9NLEc0lkHjlrld9fHgL05gZmC
ZmYSW6ctOjNUh4I9F3G0LFAL1LsmRf0F4QiuHZMy4JF0+OouWRO1YU1eqZdAY+g8
+jOfVNloFBWA4/cLfZ8FBziIpLsZ+ECRGrCTDPPuuc4tk9e/vHN+hf/qWEWBz+i4
9O4dp64FIOdyZOdJcDPwU1CPj8y5EIO4ytPNRSgiY5uzUlOVoDsCe7hhkdzAyQJL
wUoTaLcfTQvxnOT3XePJW+ppvDnE7Qn4moYZ3PUecY6B7HR0hwbXFsoYxYVNahFn
NpAtH/DNLuvPpPcJYZoyWRcO2SgIPd6d+odw37J1i10T9hhIpOn0MX3ca1Jc8WQp
fciV9Fu1Jn6TVSS+5xH8r2IeJTg3rcr5xyx/2iddwLKuo1xXm1VLnUbj0pC8RyzU
A6ZQnzSiuvM8DzFu5hJBpdNO+7AYC8swuoCVo6QKQ3FcVOCiEBsdxyUm4OK63Pu6
y/uyZMC9ar9Cl8SRnkLH9aJ7E8agvqx+n8zAOET8PdhE6nI/d0okS048r0xRJ04t
OH1QXcwbIC+xXzE48aRUViucBMaZ8Ph7fDAKaf84mCZfpWv47fJUmf8QsGoqUTNc
sRmMdGaMOogRj50b7xTXSa0mneow8jh+zyV8v3ktOUraXMCkCAXS9KdQtzo9oDVc
L4YT50okrXsrmUS0aDp15hMUHoeZ32bTblwsPpOfNQUDiVnrdZO6p46HPLdWTXtD
9J+RRW3Y1aBAxbZPgdqzzTl7JkotD8E1zfM7wcTOLNC1Ydt9Ueza33D3oFm00ynp
dAFJ72u1uJEVMrxLfHENRe066WUkiwk8XEswhOjmPGC1VJFIj0aXEejAp7LUKQGz
zs+ebfEAfqNg7wGC+8V0BapBPFeM3/xYKOVQib1azHbxlJl4JPuBD8CaE2XKFeLg
qgpheIF9StLtqefJgnJn3TuC4FN2I5hbYz8YB8IFonmR5x3cFSZ3QABcRxVjv+HN
VhasAnzv33nH8r0WKSK3XKH6bFBDCD0ibwq7VLIZhf0HBAMQn//X1xMqMpva+yES
kHsOAjPtQFnPNUgId+C5ZmotnVBW9F4UGO7DcHq3eosOR7O0Hr3BgKzp0BlvPmZy
PrcOMqJtFsYsMMT7l8nHW3eAuRlsSqyOBDrPuiSy1AODTou7R7gNkBKwmMhWBNrB
Yd9ATTIkyDhwvWffzln4PvxL73yP6DSvdYwQUh4teS/k6b+1mhRaulP7CLUGra/P
/wg3pX+uzE1Wm4hThoUGya5liwgBz0IkEoDoBTNiMzQtbK6crY/MYtZ6k/teAeVE
G5n2fgegS9dmI7tTTisRd/gGEaQw6BUib80nBfMpuDoP8fqM8WAC1UHkawmu3vZL
VX8u9JCkAuNfRJxfOR+7hwXMflL+uOvrx4uMlblzTT29ZfL+a4LVCJKuchlVUH6z
/JDxaxEwgo0ZJl6e9ZF8PmcIXZwLPSOshi4N3ErWhth8Jrm9ebI547evjp4pJUtK
SelZgAHH6W3n2ahHopoXIdZM0eiZ9967r91cph2hCfUcAPanp5fbzrHU/K6VDDFx
sIOs5/L/ZnDKr0NZ3CwgYjxXoUYAhReZvH5FXb2Mp6iQ2Pl7s6tuOFMXYl9fHcSa
bc+uH0yNZUh5cdKq87s1GfCEll9pjnk+MwXZGYKL6/DNd4DYCJLo5RALeRClZAwk
qhTQOqCK49+QtYczuUT/C5gQbNv0BzfkiybDpPBT6NNLmSxdg5MlslyM3kKFJX3A
Fj+XENG22wq3oyKJ8/KoE0f/j6VIOnQEWAf69ruBLNz77JsLz3/CiALGQzCJZId2
KGuQcCanlXKPotyj0Cs8aTxUMnpsmazPFPbiXJqZMsHjLbN/2+e+GUPaNCL9oywB
N/udSGfK6hsFNl17gOMRhhkvgsrA9ST8GsZ9MOeO5O8iRlIBwf5q997LARfVXZib
3CuEc5npuokkg9y3jxa6rslWSj4c/BC1JcXNCbzZWgr7GwaugQEz6oE4vTnR29P7
l5BVemw2p7XqtkaFwdZn8tP1yKfO1M4wcnJN5C2rm1WAfzqj9SkmjundV+8ugoSl
bmsAB0RXGM1OtPPuxC2zjlyEuhENePypiShCoEKJPFW8SOi6/fHcAmqgRGlkBYmz
LFSf7CPlozVJlC6W8sXG4NrdDYUiSmp7gntA3dsp3FuXK+d4AVj6ub5OUEjeCGIp
dHMrgqfEiLFLKed4rkUfauPosCh4NoSSM9zPNX2wWczMNM5IQWAmBg1hdTDwqMlG
416OHYI7uupxLjwVcQXJeunnNnnvSkLnurqE+Sy+QnajNpY1C3Q3Q7vNlmcpjJUn
UqAjJFYUzo8eVlccflbqKHlpo2MrRt2An036dqK6TQ4xXpYqcCxpUGWRim4MFHaT
jFPgv1l4Nr+iBI05a9oj3VZM3E7m+xv0cPF8i+yqEUixPhb+jZRlDqJTKlBrFeRo
URxH013U2ZdfBNtrySTD7TzPcjI9RVLaIfQMoCBglOZSiqaZELTp8u/AIBa6TGFB
wR83/gHwZRDXyCjUANJXzZwVrTUEKLqWChpWSKCJLaQTWoqvO+fN9/7mHp26FT5v
8MBTfKcch2reZ/c6eIWFjdE7jNYfsFpVomD2SpHObSoDKD9lZeDoZihgWTgZSbUe
f73sn87/wQnYIJbyh8Z3Lyan9pSKwikdLRdL370PYwd1lxMYWv5mQ6HlWsduS2BJ
UKOCXrX2UOpXPG83SR2c4qJVURwS90jWFLdV1xEOdJQ89RCM6yQGr7n4T3mYmr2G
INYJKThXoraTATrJFelDeDsVS1svRzBgC9nDheCkKGji+ctpnZc5QAfygbn6wZFN
FYB1CmRpsBBGhF4SMIHtpoJAAtAWnRQZt1n7QJDGn7WHuMrTQX4raxrgguyUfsMy
C/2Yw9qlWGK/oSnMcSYy1F3E1c7D13MPKru/SpKjl+btfbcqc6BMBFj0FVUxPw8H
9+qpjG65WggB/9TiG711nk+ZDUdVLXr/g+1bWGygmxy/haoTaN+VYU3Br/aLSGLu
G0hClZiJSPOF6rKlxYzeTxqRQIQjMkiaz6qUPugo3l4loFFZQf9wdheuT+hVplux
MQZf/PDdixhz0smGxOeFphlNQibrC3/cdGN1IXDxk2yLd+5gVASY0QyRwTGVdlCR
tv4ybylMZDvwa4b4r4BGis/WlhndNWxDXDFA07wVJWEVn7o4vBT89+9sBZR5xcZL
9isNL0uNdR24FIoevPTnGVwo/z9869Rj4Ow2KZeap6tE/xm5BS4369Izh5TBNCKf
ywlLT/3xDysAx50yo47K4Rtn3CCfz8xQrDCR7ro/sN/Kc5p6Q+MNnMoJtkKeHgTQ
UH38f5ezJEst8Q4EBZnkQC6Y94nBXWKcaeIxO9JogeJ5n0fjBTGE/j7to9k6cqF6
+EHRfhhU2hifKBpnZZjNJvLPRVKAxbeFUXrD0b5itKP4ugrNLcbCAj4KH7cXghCI
rZPSSqBR90vW1+LlTAAO3TsvC+5PdpDfR5KNJj1pVt0u0fcrNjoRIkk45KwjL/91
lwbNBWdeZngaQZFnbnvSzNWZZchc3BfRP3MEe2myYF3/RxOSvCR+EfLmkcZjdzNQ
kghY8EPGFjsIxUtNHzStsB7EQ3jH+zKvRIWczEOcgy2U2jUwHhMxANJQmXtfQpcs
oQV5FIGqz0gwZ5+HBJyzxsYB916NnMfUEhLXVtiKF5wEAMJ7vm8MORwQtRO98+Ek
1abtwiO5roJkixUeA3xVQ1dTqW4SyW7/8MLfBragNgBdDHbAEK7Qn9uK+Rbqn5zT
2AP+QZUSOMrGqXPLsfXDc9g7x9WqacBV0HiJP7p0XhzrA+QUlRJ3UlTu0HqJgVog
YyQVwoYD7nHZIhPJZJXHKEwm9Te3VkXfqcAUVZX4KhPVJZl+IyTpBomZwe3k3tSr
LiXwKwG/4YfwOdkgd5VSVTV02Eo/yPB1XEX2/Swxuh201PDjtgRVilqU6Vdv/ixH
Efzip/XOXX2TCvWDY+7L5OmfOD+H7iRCcKtMvf8h0pZs3PreXn2RdAc7MzTs9PeJ
DoVAb/gocIEh2I20ighwIOfj/0VtVmLclLv0bng6n3HtgnQ/MEtXfnSo+q0vW2Ew
pERAy46N/EKeHrFwBXgER7jpOAZCDV8WM9bheBTsq6DzcbgEWrBEcPtMfwK0qLqj
IGrpSUxSfi8t5dELwbqGMnq30wNbCo72+UO+FKdR4qUm9H01hL1un/uU8CMH3Uac
y4cM4xThX7r9+UW7e+Q1V1jTgORSVjyJeU+QtaTvMzK36yJtS7W5NxfCszfLnC9/
tJpcMeav2anN3jEfCqekgGLYG4fCTPREgfzoonATODJQXzocKGEp703LquPHgf6j
YrGrnnVT92/KsW73PuMiNd2UNaKyssoEjbbZO+4gKhTW/yxebyoCt4RXj2fo97Ea
pjC56OQND0ye4t/GeXWH7RqbRhU184USKM+rN05ZylvfCPRAUCF92k5G6ZcqWGM+
Q+bwwUO42WyiHciG0ILLaYFft+hlWTA35V93oNMXLkUPR2tt7LLQHi2HkIpusHoS
ai+7H60pMwqxfGND8YRswlF8creDdc/zvwIpNnKxRHgieqwE6Oin1D//BYhVmat7
CWwVG2qhghGpW4gyFRfQD+mE722KIgyvZNcNljb+i9DxwwW9qd9cjdyINOVXZgtf
TqqTMn01qlbMRA53wwXTPDl0OVbiGrORJztX9FCdfj1JcInBO2BfMhG//H7YrrPz
QJAwFwTSQg5FGx48yVUkVYMarOf5grf9brzuwdkGinbubvU9Sbak1b8+XbmD0Chq
G9UK7HmXTN1bmjE2QDZASCJ34MZUmgQs0hfa7Vv1TCA+gf8HP4vP4XDI2oARnRdg
vUaY3E8lStEQpf1GvPvqWBUnbVLZUXwykpUSsy7LlTVhqVzmoifypkyf7O6TSFT0
rmssFUKf4r2F4xcOUOf9HxT37MCqOsh3A6YG3+Pmu/86kx364DrnFSqj26FwDXnu
vr6hWs1t3INdbLvip1jJ+RFwl+8ZWQOk2VrbHgs+VEolUHzwXi+zfXZR3oZN9XIS
C0NYCX7hjrbaZDsHv78MqdAjlJ2dZIVsqhMRSL1ctNcuRe5UcPMJMPMXNhfc70ui
ql879YI70ec/FfX2pToM+OD0LhDsbR6oHEdTI5wK1DpdSb+SYZOZQAic+BstRfyI
3AiqjKFbzZ1gSqmSqCPeJdgS+ZXnoAmAVcdguT/TTcypu07AcBILMMzKHsBoVJuN
7RRPG48GodJzwd3TiP8/l//cKITlwYaQDgoVpc7O0zn+baqMkl9EbbkA7PxHfxMz
cN3S5/zmXt42NdMnq/h5inD3/0DSYaZKc2JY5MFcfjWDBX5ZFiOfaG7kzcyw8+9y
/H+8y0ZPdGEek6ivVAAfRdxaOhq3+D9J7TZobrdvOp9nAxiX2ls1ULvxQZ0B8DZ6
zKkMk+KZ+cVhoRVFoXOIKPbS8yqyO9vYzZ5quhhhXjrhcLRC3psW7PSLvCNAJsB1
8+ZFB3GhI4Hq1mqttfFe03VMCwC3tHaizkHd8dpC2YkaE6d56vjpBKXGHVNE5niM
L7mSPhLvCD3Nl93B7BEo7oagYzdfbEhQt6Hc8acbV3Zpnf/5BtbPEXrTQx5D/2wu
FzoMbnWR2PR7THlWjGwYptQMtYMPJbxCVOrsxkDiIlRFat7y4zirnepGoVkceMHX
66QG7JXgQfMaLlNMEXlBhH+Y/69SDZzgBqWjVWIVRh7HHbQ+ZLPC88bOWJ9k2FQc
pjIB7ORGrEg20DVEYsAGB/KPOD0AG78YNsTJ+gBz/HHPvkoCsLBOvtBc27zAOnbL
LnS8iyTzhh/Jwqe/LmSTcrvd/3Q734rqH41ljeqcrh11G26I37K5X/wQUIqWKoC9
j+bl1OIQ0PaKuGPaqIpmydShCapyoGCJRICZvEEeu+0SAP6HlMWVHExrmKcWzii7
Wa6+DJloPBBtNHgWZ8CU0tJvKnYdIuVMAqYA40mpQgbBUBlt7PtquocYikbXoAd1
K3vEwGUzCCK5wh5/QD6T/sv0FX/sOKoLI9dh/SG1W7MOQj+zgaQ5TxXXYVf4FARM
4JiKZvSCVpmGdYBIUL/UscaoB+UFdZq8dM+0GjKHnaTzSiBZfXvNpZza2e9O5aH5
wbgEQvWi5KZoCgom00QtY5jtqhtJ8hQ6EcySmCMR5SdWgvl+yRNA8BLS9uY1WUaL
KtjE5r8jQrATmLoemVizu+pW0jpxTqBVAE2IanhFHMsaqL90XR9LEa+A2kS1GAgK
kA5/Evgz+h1KLxuFrcSRIWXvbHJta6OItghkghywifN6/5Rkme33IvCULisaco2w
1d+eC3VOX0B6ubK0yWyp6xVWI+k+3mAaRIjsDK7HPvP1wX3edasAtVfjybmYYTYl
g8N0SIATAqsnuyIaLnKa6luO6rHAXbIhCrGXwDEOVRm8TXnrDXfcFJQz8PeypNkH
RXwDclpa1Zkb/WODsfebKSApXm6D9AN/xOYyCmkly2mwjgUAuxuPqcFAx5J7U1iR
B9IsZcETIstY1O8YFpLCue1jp/7gwCQlgZlqHMQQba8aV6uwKh84fEaHVBuEV/Gr
wSLRwt3niimOhDFZMzKYtc1qedenPb+uLTv6+N1Kt9B5JCyJD536PkK3LSQBluwI
YfSNGuP78vLbMNeIWsmG8siW7wN2hVvZNG1fDHl1qVxcp987pyRL7IxmMmQovfkR
lYVv8PiNF+wpB1mJWSWZYZHkPSeNXdDZQAZLKbG5rU/GVqQQiZ6eRvRaGOk57yXL
v0lpZV1CNAyVxkL4gh37GYTgfGL12wT+o8uySr/WCf2iOApAhBFHXZxK2ls4uFCy
ujXPo2Iscc1LLhCT1F5oajCBcFYfR/+WaCVJ6LXCUlrXBWis8z0buHroB3mHuymH
hBa38OcaQiXRTMp5lWFI1QTgnfcBvbaP3ErLpov7qbSRymxc18KTYvthnf7tZTOG
GfhJfdbpo4qThCuGjY9c5dUPc5hXWZbQhVYIegJh/b3f9vUjCwlaN6YjLQBPttVC
9ONN/Pbk1RV95K9kA4Z17KuV298n4lx7toUNcwXgyeaDgNi5fg0nJUVT/U8YaSE/
l4nLAmw8NsHxgNLo9ajjLxI+Zosm0oZ4k1GZbVSXm7rMsec7baCFzgyj7nWkY9us
8P11GsL/G6Dnzdr1LuPj3oQT8Z3SyoRW7Tq71wPcoiaopbGAsLFqwHUg+ejbve5S
bDC6OyRlZFG6OjSdTCUTmfTrVOejvx+UXJcT5/pZB3j5HBbBEZZ5r3coze2HlZLs
vQtZaRWG70Ze3haRoYyHdZE95p8EgYl+60kvcj8OG2NMKMaO1jZUkDyKLS0Z6eL/
oDkye2OWxX5YA2lxZfP43loWNEs2jNk1NMh50YiyW7NvCw2uXSeE1uxo49lttPks
N4t+9vEv8s+bRNAxCsWmG3M7ujcK0WAfxg4QsAbRJ64ChukFsevEkAuKufEAyzZX
qL0JN9MvRCKM5xNeaIrXGiRb2d3L1lKakr28griTRRdY1KMXoO4bvPI9Akd3PesT
9Ir/ASSppkRZphICytVjWFkiYZtWfBmuzFfBr8gxnHB5+lAZBKFN3VJ7zzoZFVBc
sxNlO19k6mGOS83YaEBCE7uv4DgQpbAJKJlEf1MEHYk2XVCHG7QMH3PRNj6v0BPQ
o5whKkCaiApBHhWDA4rqvElPyfO8NcMkZbbPNUBJUS8cDdq5o4NGH7x+JRIjcutL
4LkJGBXlOLtJXrdk3I+LAdDvhAHUpSCXMAPLUHLoc5C1/nXhN3OiMCXN8scMugF2
JzoPz2gzx/WmutZpQMgOMG/oTLomcxf0Kn0QQr+fJehoom6yyIrJgczMSHSvTSqx
XGJbJybgbv5xkGdwmoJlPCjF68Ng0IKOBKBU37QBIp3ydZzNDIFQq6o8o6ldqSHt
DLJfwlVdfBEBTKxKBOdVvZqmdt6+YkbaMIkjwlCyfRj+PowSjHTAmsYvDpdQ7grj
CPPz11INigtmjqPhON4YftocLImHrXH7qSwOGaHJTSOWbpEuOtwSgg7wzgOkmqvi
heTTKPjscOYWk12IgPpWMcLAWRj1aUepRPKR2fARaa4Z8dSSPWNHiwktnpYSaW+r
CAnkag2vMq9jSOdlQIXhEpB3I/m6hp4BRmCNw42gB+z/rUwKG9veDkfL6z2nIaMX
AoLXoMcoJtJdd+z0+shZcvRpLA063y8g8bhAO4hCsZPS94fTJNlgtt1P6Z9+yIqB
/wYx/LtRVW/Q+5XZyauDd74k9vr93y6sCjMdvFjxBwPnjEhVKwU983mwFyNsMDJa
oF2H4bsjVrMt5kHtQHIAhOh08LYuKuRKlg/nC1dDBce/awZvIzhUV7L+GX4YEhtF
DGx1gH99DkyI5+ObopcqpeaY6LrCePNCLSg5YBxwqkP/Lr3BxDcJt5tZpp/UyOmm
KhQE/tsYT4RE4sWefUKkubY6k7Grx7j3ooC18jzbAVw/GpB1uHmbfnYO00IZURYW
bMJAEzwoDoB6Ol24Tb0U16bLhyesBgOjJ8AbdFXb37PXwAqnfZANEVI+KCuIEsnB
jYqDL/l6Ixt7MaaSNdE/oM5r1dWFHSDThFDH96ftv0npq0Cv7B0IGBlTS85IwsRI
0MFf8riMfNXbm68zWlWBzXvN+VCqpmyPcCdJLiAQEcKqs+hHeK11IoW76Nnas92e
pbCDbsablY3zleu6Nvu5bnn3nDOHpLsybRWJs+RsO9/Dq7Mp4+JPdo+ccRYUVblA
kS5obcqrdMhQSLAcGew/CEOoc2BZTNrV3NTHET2Or4BlLt0UwXAdkFv9pa4K2tcu
/QgNBNH+5co9WhPpMrTYFdPzYnlRO1svXwnDDnosYKAyodZ1v+DOJSVZ7obmolko
VhZwMj5KMZ+wYnvsioRTvHMX/Fl3E3BYcYXuKPWzLtaF+9uyp8EyzhXm+4qzzgoN
F2CwPG+lZ3weHvbZ1CV8KqgPNpt8ATomCo0J2vBN4XzTvOGLg9YGKyvZpEwrmTiF
Wjva3ttx9t4u0xGsZvGUolA/Byaz8WhLu6kusaa94+EYvP3gKnFv0OtV05NyX0fo
JxswnfaNNADLIWxoeLNF6ztVisAwQ9g1ykR8mSLJEuA74+FLnbO6zMNri5xBPV+D
mJwIHTZxLemNw27LGEPYL5HQbyFnn5huj/19lZjoiH8g5SdHuNtBUWbaCfn03pAa
PxHHgLoY3r1A/HtjUmbjXBfQybihqNK4j1ecoLgmdnf8oIzEikDV8UfAXJIukW+W
gpysbchgUaSwENIR0GgEUaUav0+DIVE1bG0AFePqWPcFPSp2oPy60YUQoAJeD4j1
NaJJuF4vLGj2opt+Bq6u9e0e4wYNImLsEArA2CNHEIj4zV4g3sIzL1b0UZ23Wgrm
9ttJKQ2OEk4d8dx1UC3mLXZvtRi3TnrZ2g6nkyFTSLYabaqDqdE6NlB8LzRNVqcL
CzgzhNkUKNtcqGBGXAEzOhFaur12BsZ256P0XmxmE1ZdegZ8edWWSmyJnNy6fxtI
BsFiK18fOL0a6lKTzlwYF32u3VPgrdNyBcuq6BMnib7BZ+ZgQhYAwAm4RhGqrYxu
FYUrLxS9S7SEcbfV5Ipt3HmEpTZamEE8VQ1mujM2jyOMqNwnOItdxYJesTQAcgA4
P0BIARlG9aUskLQTRyhY6vPxly1eIY7MlGEABA6622HJjgDLxkTs/EC9vp0P108Q
xi0fy/7pBVnk5A6gs2XNbvv743elET+qUGJ6fYEsjVAMJQxoPzkccc7843OO8F4n
WjG8Sed1KBJdkM9nxGFbbJv5zE0B0/jZ+OnPCC5WxQjPOkhQTYDblXJjWG853y5E
GIW88cV2c5AZiLRHklNi4ZhjvcD8hYIu1JZD7NwsN984oHGar9XuBT9TZ7gp69kF
wzF9ehIHFYflkSO5R0JTMQnuYYNOUmSrom1S0PypkH1LXtPzReHpsoOXIETalcWu
IsHE8P3BFXxV7IgaP3pZLUWT6/6n/lRhmZRY3GaobdPA1qqO1mlHZirPaNtt0Bkj
o0/8Tca7dQDLOVII0tNqT0BZQ+CzhoJqlFkIziZJ5TZOQdQlJeYcFGwNJHvFbu9n
OocomNBliE9zk9Yw97HM+b/bVgijr7+9tAp9fdGesPN0WZvytpJv3CurmXfikwk1
N/9T3yl8o/YM2XV35/z2Hom6l0sICWdlxASF0R/5HlIQaH83AxGUmlg33j5Bha0q
zWQT8jyCD5WryEHNL6gKKHSF5fT0B3ECNPV8oVylZc2i0xEEeM0GmmwWYCSiH3GX
e075iqri+6sQikhxDxj/nIJyqI6gVHGCX0j/VkkJB+0antDnVDR64B/cUrnQlJNa
Wvr1+vaSEXVjW20VHSBCy5zWH6lJJ4FpJf8NsxBzELPiePPA357wSdAIEBxegR1v
FbBmjtpj7pSJBARaTep/xPZ4rPM/TAILrGpu7ZNlsxoWX8sDlkieJl3xpxIjcLnk
2jc7W4eGGl14Skzco3yKJB+6FB2fzqJ/bO5kNH7Pt80r2OJRjg8tfEG6SQWxH/VE
mVo1G6ouKlfyxMZ7mFxB3aUZvsGpVhvOpcpQphy9+v403N4C+zicXLsOe2vj3pmB
UxfIdH1BazHVuJDtaXtp5NtNNboh7aS7k5wFu0s0RVjvEvd8ga/5e/VDPOYeuafR
cmove64ej8uTz1JBGxIXuBSy7m42RBXxv9K57RvqYNPFNeqHtVw6ne53NdwqAwT2
TpNjD7r83menJ2dv69hhHBzgURkS9HTedk6wIiDk8yI5a8vENUeQjm38eJzkIgV1
M+ZQXD3QimrLyAkTB1LX84+vQeaKao4EE22frlPr/3ciF3X6DE9tajrxtsqLyZX2
w0dSGEZ39Nmsmm73rz3dlWm0dWZKOjrvFlFJ1ILL4kg6rtksIpomfq0q12ekFYZW
mqNS2/q2unN7L63ssAy6w50mVYFeC5z1xgUY3vPeDG5FJIyEGcy1FLu//FIz+z0z
Mb7qUWxI2azYRZrfr7/LPiRC8fFo5fUuyZpKODdUAaPWGndZhDiSkDOIxK8McRW0
UGyrCHyhP3LueFIN4US3pHXvC+G7sE8i6V6j7Hq+K8M9U4mRFaBlLuloNQb+eR9F
5sxGmX/3hLaBj+p3SBtKSGpORn2I2s4AXzeAGMuI8i/xe/ko+2akl2+Z/0DZNxys
lVV1SeNrQp0oiuw50NBOzjsRicyXYavwsVEq8njlz/yJaaIlMb9aVMabikQUtLfa
b420NcRP8SsIrLbGsUgDcFCcBlmMJqIUvTGq15iPx3N6su6PXDA2Faof7l+BRfl1
5efEBozmpOQ27GA7cgQvr+Pu/QdCO0d9iq0LshSFDHXuPLwO4Jx1G6yxJn3dDaCQ
POaHpSj/UW7uuBlxEPcJE52hmtDkTZJep8qcluixGqBU1LPNgTCbGS8/xF2JL6uF
xVw63eWpMrba3HhsxMhTv2352I8GhZE2xtG5ODcvldCKSbWEK9xtFcAVlY79t46z
/wXj4fmjksDeit94SQPDviT3nBSyxroKa+jTmO4FvbppM1nKKwlo2Rjt8A5NLtPO
PrhjmxGq8EB4LYhx/+KIh7l7llps9ycdyIi0n2lm29pQ3c+ke41PvU6yibaslzI/
a3vUwUUbKjfuFdFkYFxTWKdyGc9cD/lLRmBEiaAOhn7EgW/P2QOFP/594YC+Jb2j
7ye4nImUZznJTXzGJ6j4jGpVW923uQvOCQ/WJDIO/UmJGTG+al1/sFuNeEi+ON5x
kqzzVtdTPkY4rXlaGj0eWJ7TUlTgPRe3ZdzmZ5xcJPbARAPdHVtswK3KYe2fB/JD
lMNhdfOS3CcIoV+JlXsLa/orQdq2oIAeqdGaOokX+UQMuhXbwxR/6cbYUFpVkT34
HpFW6CHDRcGxd2D4dgB1i5BPWNbdzX0+AvY0wtW5dsuo2hcfRARdzUvoWqfhkAFH
TPboFDgD6KSzL6z57MxoK579K4PdQlLswhXxuE+IdcI0ppFIlNKv/KDNVMTV1JDA
dEnOh/oOb3GlQpfzbddrWABNRTvfgTWPeqXNWohUphXmGuCz0T1L6WZrYqv27RCg
AjIhLTIcQMFeQalAtbFucloh6l2E1/Sh0aQ1VZIdhzfTvLUwTQXxK7ZM/jedCbGa
ErZz4vG2Np32UZtDHUefGqEbTh0DtSDCTfMTGfy3qY/BMhhtAm1GSEE8a7JWXyEX
4lk5qkGx7BTEUs/IPyAlFszBs8igclhAA4CDAYycC32YjixHyp3dlLJIMJ429ry7
siY2DgLbuGZ/EJToYpvt9gOlr+Eiq9hFc1OLa2EY1mhek4oe9XvGO5+TnqvshWQi
G+1AcMh2KAmsiVI5MgqBOXMxf7KoJBewrqtDcNO7WTth7c235PMmZLbylNwea545
FySPQrENW1IbSAaUFM7jGP6iXZaycUtEEdlgutnQ8oeOuDwmWV+r9VwgLeeabYPP
IysD9IcSSMpScFbGvkCioSa/ckgsq0Pdbe4K9XAfZzig+yMMuoa+2ElaiWiCgx61
pEv5beR5IMkxiCeYw1/yIkbaxBABIuUPV6dgE/pJ49Nw1zK4vJzO0auwn6kgfPmh
C9ENLCZTMkqRBZOK8v7mqSkVxQBFWjVrVSU5ROOkEbF/tn/oi+hONjOsrtbw2xf8
aoQS0Wp6rzgMtIjIO3nvIrf3qkdXZVnEAbzxNpcNHCFywN57U4/Mt5H/FPM2WfKy
9nurUPBWEihixZF1yJHNoBL55k5RV5Y8hqZZQFdb1qefAFLY3RBbgWe23qPu7LJ2
m758osehEjQRnQoj4Z02vioo/zgHwmHRCyVEYeXg43UQCwzQaKyZzCsgpqTSzn+W
WeHavbPHOYfDQvOBLm7G2rgFQEjk2parAQm98GNu+Nm+SuQ6s1Hr2Ys5xs4h9YAN
cLDBpkUr/9k21vWaZEZY73bgKwM+LEOlgA4qyrz9zLbulsdkb9+PmG5Luz7CbrI/
b1AnCHBHKRR31cuB5QwJp9i14rkH8jp772GRpT2zfE8mbUCkCv5TlQNuGSI5dS9Y
Xm0C9f9a9QiwvSRrtCOgnYCswgCBrGP48K7ZY231fo0Sq9pw/KE2yvmyluF/SS61
lf9Fg/NFt6GAc1vNpIu2fUuhKRPY3RGnnvLW0dl315vS5EM1MnFmOshzJ7OMDOlT
UGEX2OsWUQzx82vEhvTsYGbGFJ5HPAd7TMbDuSiceZdC3XUFMrUReRrfZJy6/r/s
Vl5CI5hCvl+2CTGgodFutpogstqEr9aGWLrQxjqeB9+JtQ5hd/Qcp48T/nxC9ARy
86DKzakyMSo8WbkR+JtoUs6I9wsaNj/TDtERHGKGlxP0mqkovQJwzvGKiVYAlO1E
CoB+52d+nWBdsNBBou8EmL3I2sL7JvMLsCnk1ozJ78QH9yP9MmZX5dGJATS+9Ly3
MzOwuvYua/lvfFlpZzkyHOYoifj6Hm2ubU/W5E557GHMLXO4ncpfS7+S2PHrgyb6
TaFugckpkgCImrncU8Wby+urbwPYYJKeaqTXYDTeLvEpknVdq2MpDC2F109hlFQT
SSy1v4AHBE7m7co3udMk9lNeVPw8WtwpVZ1pUfH8dl/mL0tMhrgPLf5/P05gIlt8
0ZbyIHE/k3V1kf3bwbFYDxYDx5xca3IQrojyUSynfZogTRqtFwskVYJ/N9qi+DXa
br+Lr8k0IIvSHYsUmKfGV16GBhWOmpqoXXlwi+z8payWmC6OkcQhaxtfUVXCf0oW
QplGQ4erY0DzJhlYLCxY+1R6w8qkyk0OnIG9ZnutHDYtsBjrf3L2kv7WI2akH2je
D+qrFVfy0Z4PGEt8yoyxxEtAAjMxhaUgc4V3ikbLAonl+eXw8PVfCRLi/SKQHIUl
e6D9dqunKuLFmsxn4AKBPBGaXXWsjNbpNgMrl3q7K2wYzhKHSefk64uss70rPgP+
nMqckPonex5tgb6Nlw1ePe5WB7ulI3UT33gM0P3bWi8O/aW4jYg3wuT4oMukSFXJ
bihslg6p5VlxFo4BlXmEcuMk7gtCfu5NMG87sBMWGaSzMhJfWbPzwfRbrqda/Q0P
5Js5Rvmbec20vRGj69TRknRB5s2l34oTzReIIzF4vdKcp8xPB0v9F+9Ou9RJJtgc
w838Ygik3IgjO7JUKEMV3eE0GGUB0UPdUEbfQQ4Cxjm2ZkKbCxu5FqlvgYD1Ph3E
ig8pscyycuscrHoIm+wFFkk6Jb0QItC9/jfjZWeIUSy0V55AWw7FIIK0wVRgOQrr
JqU3nCdccuIdW4CDVUz0mjcfAIr9m2y9sB9xXGLjYmLb4ZR0BF7gjTSmCS9eMER0
nCMASVGn9D5kFA2mYD7VBymZ6HV7CaE4eFBd1U2EtdulyM8QFevifYJBRJgHel+2
B456wrxyIDdsHOjFpWm+FeXCZ/spkEMfpFOHu3/IPoa9qyC6MYYU4bFIhDFqfe3J
81BTxzNAS95TG1YyY5m4xmoDRTY+SWjHxCvjVlVZ/iwC6wjJ1A3x2MFOX6zg3VUV
Ii0vfRZEfCT0BB5WPXOOeKnGSeVfo36meYvWNNx1VPrKh7tkREWvWziO4V5cr1/u
CYdTCnlVxuGmHxQFislxORJo6aqaeOAo09LoyDyVOBOjzHVnMPzCzrBaq949j1+z
aLUkVlybRGWlh7qZkrRy3lsTBy7VguJO8j+NUXLLNVa2/jUCaDFWSLY39OUww7jN
3UQDr9F3EiLWYpfYuXGwNK2bl+QdK9tzPjGHMFvRGIUDLwXwc7in3o+xYZQ1a4Vb
6pdkAAmedJqlD2B1uqQt315mfb0kQ7Y0NnaWNbI1Q+lmClzEMUvZdpyaJDIfN/rQ
QamEDi9VKlFH3hDd/CdeIhwK3Gxchg6m9MtDGWFEUkaBZ7yCzTqKi2Mb8gTV7nr5
2KJs9CxU/ajQRbLrU1EBrL9c4CXCpx19R84pqz8liFhedTbN1H7LOy9l+izmtON6
nd/iXoB9RNyKBQ3cReXiifX2LQPR9EdpIlQCiCh2r2K5xt0o7ZYEaBDi/wG+dIix
BDF1VrFD6lPnF1OsHCe+ZDlAw/wo/UmfBQeABAsq6PHhryrBfWJuWa9pwO720MNk
cD/L88lHYRNt8eNV6oNmGMAWnRN4pdVdVZy0K2mcaMUa01iWl5+tluUCVuu1oyTB
bNV02AGpatUEt1HwlFs9JKnoTBk5Q3XSaPnSgz5/dOHmpaTBskJZoORvwl2J1mJS
JSQU97euhS9tTfk+lmmbWJHBvdHWTshsoaNoxHfrfj/sOYpw1kmAG+8usyKwNtmM
RFUKZFdMlbfohMj875/ZY2z6NMxlAALYbrlpqGyazCDhXjuU7gaa3+ejtTqHjayD
ZEBCxNyBKP6pLW5+Mim6fFZbGqfOvHyEyOuGEds6jqONTXvd5vGY+UZBGp+AVHgD
gsyv3P7VADCeHjNlFfraapg5xRZHrY0YV6QTbV8tSTazSG3Rgj604e0WCooWOGm9
PFHBx9vvOIi1t6qn2YHqkz43R5VzQajx9n2IFFYiUpfbmWISE1dPkb/UZ6//o8NS
rRX+pJKlg5l2iiW6oiv9g/VGwE1hPWoq/RMcsq+soiJahnJt7NOK49ft6hE5t2LY
3sYaiVPcFmXz+4fqMLTwM+ZKoUHjOC/xOB7SwalJdTjx2TkoSUGm7Umc9iLSWS5R
nkFGHW5M+SEjAnks4qcen8oVdBuyTR3L2iVsmgcm0VUgQT09UEbMPQbrPuE8YgQb
lOn7/I9DxVkLLo/1QHBoMGuOWZj312FkD+RyVkQpRh7I0/nKmfDR1QzmuAsnEpdk
YOIXzt1WLawkF0xm2bbtPtBIZrCSK2Tjzr1g9cgUfpHbN+YHe8ZXSlS+XIcCASX4
XM9N0c7BnQv1nt/xUiVOEZEZqziFxUo/q4m83AZu1KYuJ3ZsZQK4sd8aKUTz7wqB
ynfQaC3iDmNXNyuvAaDPnURNFgjE/JwZ+1gT25HAQ840raPVC75GG/u/bh55rOf1
6tmtBA0ycHa1WAOnXQsqtc5SK5Y4fXXkM4wvQBkCYODaLcDDIkNtp+Vcd9ka8Nnb
OG4pLnutRI28zg9DtfJ2nboxwvFJRyCgIuVAmWXrpz1LGZvgm2unDl/XOmoXnyyv
hNkZIsBIt1qKYTmrSisTDlBfOg4d95ppJVKQPJ+DOe2agvSExXK5UhaB4MxIwyKD
CKaRl0kCMyPLhl4c/MeFZVMdwkY8TS2tIyeSr+i4TXLvawDT7cnOhMWtGrUT9gpP
3EIBoKiKas5ysOpHgwlq8TOJ39GjZOsrlllJIkSj6Cg9LrmeEYSQzbLKkv8cES6G
GHpsGpZZ3AP35GbLGOy4kYmioKEZRIWy3y76F9S0NI5MgqwaSiWMZGFYAGl3r2IL
A2wR9VEoENEhXlc8ZK4ldsarQqYhq651MlJltzSIgRt1+nsGQy1Tlpo9W9tmhC5a
axbeH/ZY8BtjJl0Fx1sxeoDa8wGDAAGQt1C/p2mw0c0M9PTYGNdoFzsJOguf0AIM
duv1odb8HAqXEm7rfig9WzXDiGxkTmVTq1Ffe7xtJhHtfhSyIrL0Cz+4EViLABfx
UDnKTkFA9kq3bGA5HV00dSfmJ0TBWoazAkZgWysy/SQcXCv130P8i6sRpxTeIUlz
eS79cTJ6hUu7t32gUkW1jSkH70TWfHEohYE7T+S+7bakVONT7kBRz/3+7KKFQXvc
Cc3JBnaYQGVC92I4mmxyp8Mboi5gnKWmEWuxJO56QYdXCZU+vc+Az0aa53iNI6rR
UGGMVulRvI2tYcajxPTwbpdcyfdh7uLZuT3cRw4OjvrsAzrq1Z3JdEVkMBThtVuL
Wwxy822qNk5DbfqAWmGI74AegRBw64/Htll17LF6lX8sj258+n/iJ6BF79/veHzM
hsKtNEIofAG1OG2mQrUv14g0kriz6ZH6f4gdtXpx5n53qlVhLtQ2YhIOR5VQwsUU
2r4aAxWh3t+5sXc8I+Z1LPYHFs5Q1opDRTVtHVWgK9sa4rIlhCubbfr3KTb7bVnQ
ojhhUpLOLNoMNORfBeqDW/CjMmc3LRIKxS42JyTrMSU1BC2XWM7pX3nt+M1UnuL9
d6qn0pryTBaVwgRU+a1oQVEnf5wgRS/Vw6TykbriRhjhus3njEj5uhMCJia1otrH
xGaJ+BQkTBkra3pSkspC6+OAGa1F5mlhUUd89n5j9pkqlidX2L3xH0seH+WcVxzj
rwOp9AuXUhLOv+3ZD3xm3/2zwTPdoAepDK063oF1fOCzbEpSukUxJhomdVbBVg7j
n4HbirKT6LHKpddS/q3kNgJxajwD8DyhNotufZOgt1lMghHYTjkDqhQWecRVEvB7
kn49tcyrbXmAYthtdWychkEUdPK4A4u2l/Rb8vveZs24suFZ4w6E/SkoxIA7piNg
DhuWj6RVU+PpVxvdWnQgKueoD/o4u5SJuZ9nOVaIR6VCK7uxUYRuu/YeUnk0r2Mu
uhlO73TILK9iOzWqlsXeXgiefHFZ6HEBV71CkD9QeDLiK80Wz0vHX5RzLvdPRx5y
daCBeVZSS2LBytChXANO75byiFdDfAXcQ00d2NS0DUFZBe9DYaR3RqirCe9WA6TS
PtEecQ9aqW45e4LKiPdxgH8RTujKP88vt4N/Kes8VEmENNSs6ysBXvQGBltumz7E
93lp4CKfFpZvos/R+FFYur/pGyp7qz823u4EGL+q47mCfJq7hUW2bPNegCRAnXu3
w8/Ea54X/H00VAbFpbk+qs8dnZToea20hvjgeqw/lBFYhvbmLalA3VjFcAeLan2T
YTrFYZn/HZFxOLA+UuyekemYkm8KmUieSXQvzXn/wIZ/959r3clN5qhKC+OvvZa2
W8u3PfVVGWBZlCFrbAxf9aQlh+OoyaHPdoSmoZEqVW0xSKlOtRZe6GITOr/dBXyf
UPrcMPAnu5DY0+hkcot1CRDy4moKz0UNeffLp2FIKppOWHNpqJkdvuxwvdsER3UH
nH5GHr3h4ocQufGmUpqo+bZsARkupp7CUeHctaQgQO/6RjWdCB7BhI1jid89cXAj
HzuoL5mtHQSaW4TMBpgelSmTFiLD7Y93F1Wx4Po3cbk+jhNtgqzWMLfTQMJc6qTG
v13x6Suj1kOU3FcSnUZ84fdrXa8afCsNiXZxMmNXmjsLQ3ftP7PKBamN1EvEn5oO
ZoVcGg5sF9v4/vT4r3vIPPsa3tWZ9GhmDYFMe3Dl39AfNxw3K1naGKMeQxhJGps+
XJUWzYm8DkvKVjMSSfpoCYvVYwDBaND9jLQI2YYQ7+s3bBGa2uEna1uU7JA1b8rL
KN+Qt7axv46TayOCMBqls0846s5zUTUxbnv3MntZRaUOCw0hBUA8OuiyyILW4ghG
0iAoqJruSSw2gSZbV5K4A2WzIxSBdV1WsznOua9YR1sQrV7b6W8CwHbfljDMmqXi
jYWGCIi+mHRJqK7/otRlzLKJ5YVLKudSLx1FRfTTdEBX2jpvmEU3N1x9oiUGlJ8K
bBEz9ZbLSkZcbCOJKq/GbYUAxWNmpwU2eLfTbdDektsQ4+fwoiiDHw2jXBUrrYtN
qiuHzjrXvvszhvRPBG8k9e+c1GTt5D5PEL9fZ8qu/XBiNgLCVlxpIqdCdws6sA5A
CpcGzGQzBxqYuvdoQyF/i3v6ZHDgI7LDc7mVpuH5gyiMaY813+YjKFopIlDVNkHG
H6cya8FXSrjH6iOK6Yfhm+/09BctgOTJZGm2w26yscmucPVn2kX2ZL3ofqsl3hsU
fBd18xXQQHLRCOTa9M4tczb4P0C0wHNoNQuIMMgvaYkWXlcF0siJ4ecVcJsIx6I7
aWG5zkMG8KwvEk7R5JUgM7dJBYnDj1lJqPAXJcRoC6Bj7KnfVHkRVSrGD0h0CEoR
jDMFbSye5AmX0G0nfba7vulrwCFGkYUr9fnzsP1QXPFNULadkQmdHX68LOdIcPuu
39smPDfxkoIi2IoaaJ/uT2Qv/eLVon74Huzo5XtpOlc+S0LXurYGiroBXJuNU1bK
GtGc+XfJ02o+APjir7HwkCiS/T4C2i1wJzGQzkqMF4y9rhfZfoBkG/NYPXX+Q3E5
3nNs79+q1bEtkaf8TtDAYu/b2VQ+jhR67wXZKhk2TRT9/ssx8xmw/NvRorLe7JH0
YVtfOLdT/ktkBPhgyhg7BbfABpQu46vhm8ju5EFeaSqFb/uKBmEs8u5PlNnaYMnu
R3T0F4XwG0/96ydTwbwohOjOwDV+lS1cqOe50uOIEF9vuLjiAah0CjGmZOZBgWca
mvdxP6zIsnD4y6EEpbLxHHGV7Xjw8XYVt+m4Mmhcl8h/JpC2ZKWTXrm8Lay9JiJB
9jvcn3JXPpabxdQYJUdVBv9akqxEI1ps69RZH58ZO5G2m+f/ZOOT/tLBkIvKe6bX
GEpPM2+CWIyoe5SDV85ynQtVb826dFlNI6cMevJbkLjLT3DNo5yQ5mvui0n5cupy
JEC8/Cn3E/4WQZ/w7ucJGgVF8u8hjX9+kRDe9StUfB1d5i4xwkhnlSvGYFUs9pgd
Mojdr18QqkfTc8jhSZfTLJwGKnNthoLG5oxs7duA6IWRnrFd0AKyKABUw3zGFTOY
HWwEZ4pBV+pAXt/2d/HY+171kMUdFpNnTXp/g7eQeU1gmQoka3USb/L110YwPp2p
pjZDGCm7jHPpP+ZwZi+1M6pUfYYAOzXK7EZY6aJJnF7bY6dPggWZxMksuOCDscFy
wTyU/JhW4o0i4ZlkVXYC1nTLIOYwbEAffEVF3N3ff8oE3SMF4ZjzhMSgPTZ92toT
rKl559Esb1FxytXv1W1Ew21x/kgcdaajkC/uWFZKiJP21TJmK1PK1KvzTC2oxWx1
lIkTpZ55oau917JwkGQPyPaBryN5hHhNsgjczHpBDHm8Tfw61bDVd+KyGbZyS2VW
7TfYt7hXt/DJW3Fmwcd/RQkR4WHJpAQmwkehl5L9Rc8Qi0ogkaLy0ikMe9jK4k6N
08Q5BoDYGzLlo5sFdZnQx2EnAwNYHWoryBmUfEPlyo6a+zqnSuBcKv/rQDm+LBIR
K2mjZPIEyJ9umrSk2NptvjzGwkVGszmnKA2iryvvimgQXUb1axZWidDJ8BFjK9pJ
o8lPYpIRfbBic2ugNRT9cJBiIwF+YcMjdzzWz/Su1Gglp2I2wNBjBIyNoeTIUDaA
AVynLNTp4KD0f33mba75dSszrWacYpHmcxZZFsr6Hy7tK09GN6CeP4OfCM3S5Beq
AROeAA5PYndTa/oEtAZl6l8Dei4BXQuNQWfasKrEexOOG05oFKprLRtO94Z52CCt
KpBfVONPFOVMZBWL6P7ZOC/1W0W2VsWmedp+MzfoRtNxMDJh9CeBjKXAner4RmY5
G58XOvME16kH49NUfIiKt9975A5s5XhpxAgQ/898F4a6FRYGzOEWQcaBgDz9d0zv
fQqXF+Kx7t3jAYSbGTIKHhnWD1ZA3HkulmbHV/vX2+C6d8S24WGdLWefXDa5KAnK
WfXIpOjo98OjM+WZGGOS0K0IGhm4Qq45M8qagG9cT6I7G3eMS0MlyaWrEEeKMfIB
quiSen433Cpwnw4a60nEq/I5rIjTZ5NJw9h7cae8xfBiPWf2pKHcD0AzfEvXP7P9
hVW47l51NEtWZSrNI/+D4s+QaEd0zlRV3iyCREN0SkY=
`protect END_PROTECTED
