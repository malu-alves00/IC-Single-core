`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yRdBk0Ahk5cUAANaAOJmBgH7RpF8EcGS8kICohEKsbRaqR4bReYZQB0Y3tau07/S
1S7YIJsTEHa5i+PVQiuchj3TFBWgUR381SVUyZv9eI8C52zsjlVwoO372bM7Z4Px
KgjXHLrfhE6Vw7xE6kGWLJZIYbcO1eOcUFriqOAPWwXFHz1uBbZvybUJ0qyv3mp9
TdRNhNBbvoJpryk4J0sRottu7199BWbbx8mZl7RF+knWfuHjJtUdqgCStxj6szGM
KL6dWnPSQueLTFwdMKGiYljbRBi6v3NEA6UP0RbtPZrhiirEpE8Lz+rRDPaBNBxJ
+Vyysm7c025m8QtihUw43mcleWWnftcJFm7s9U6eDo0bKIkFbCS05ujQw8qjbMig
5+g398RlZgaGK42faxlggsdNW+qas8SrQ19hNSV4c42q3/RcyCqLAasoPX165WmP
FShz5t0O/KauSZKrrDocpT+6PGptln75hveLUu4hOu6Y/k54nfFUQuUyZSpFWUR3
IASNKigneE5wrQnvflzoQS08CX4r1YDnMYPAhQFwc3fZGO+8285nQ8g9yxMnwhqp
3kZN/mZKGjvFHJLQ1H1Cu4wnN9A5ZtEWeHE7AYBgr6lGXIdqB7WXjQrITYHvrLU5
ilQeIsr579THdD1PyshMokORp4XuI8tA2BHK1NDNejUUYmb+XSlELPmoo/lA8Wb1
7pcNtZGYlsU3mtqNqZDjnfOvJt17OVp3NVkf9uVfoLxc11dhM3KB758pkBR2+Vqc
n5filLUjPvXNp5gwGx8qT/jdSSluGASLbm3hUDEzfJqzXf69XjBTYXt5WdUiDzCS
uqU+5ZVYOvbGhVgn/pOjHN5CRBruuQXmPZ3UPGMf3E2Gu5cJnJ1CY972X/Ifxkop
M5QRlRt54aXb2iNtls6yPDGFU1yNcqYex7HzJs7lxvoKo9/ZlTjRgQWH4ZxAV+N5
c8yYzTpldKU42aIrncYxJzQRdZdW1swzRpWHZ02zTZhh1RXqM+BTgLV9lvU5JQP0
m9/s5/1Bg+/r7Bw/KlWHNdZbjq8t7dTLRe3iqYae1WP+s/s02K1SrGzPUXdFozPF
dqf3W0xz/vKQdKo6seP2269orNjgfu6+5KB43KMU5qPBs3InbG2nt0/7BvMtPVfg
jjH1tbatf0gT2RuAElFIg1SndXr30fHU9XwY/lM2M/Q+qqg7kI9+Kb7mkCefghCv
rjb8VcrtXhvzVDBChB58mHS0WDs0gPAYqtdbzNrvAABvmeI5zvAsR6YkFM6kDYhg
CKWXjFlkpL9ttPvsOnzBTQwh2bJEE93g1x7I1wsgSFBpT+0WbKqL8vWiZjkPMmTl
EgIFxNz7ndqGaqjECrtHnIfmh5Pua831qKpYdKrZv6MWqLO/wi/x2LRCOXKsevF4
hjTJyqyRayVaHhYQ9TJFx9FpGAUUaE4R6xmNv4+o/iUr18zArNOax4AELGoKKEmI
iT5OUN5+/+eNeK6bdEAQXZKg6691JT8PHDRwSx1yq16XDAOh694+/ZLsJFPQrbX3
HilMU3Lee9ZMkemAVAicCsts41PSXccT1t170E1xtcHRIFdIc5QqTzFUzwd6FJD9
LSs3geVTHtpfXfOaRfiFxr0v8G1v+gEZLfPrfHw1JeKVG9vtSHoVidgOY1CVm6S9
F8swVLi5nwUOnlADPjZsYBOasve7UKBNmeSa4jCmXq3RDklIj6WiYPLCIbED2YEq
gMeJmyONtTpx5DysJx08882B92DIT6RBGM+2QiN8tHhuSJgEy/gyC2cAQrQqY0DN
JrwENAHjWcpGAg9FFi6ieXIFVIjfIMGX8Qk9e44yhC49HPGz9HK4REky1zIkWDai
kWPui8+ABHztqzSeCFYxOpHbofFYyYZ17I/rYiLV1lV/nA8qjmJYrD1Vv7wokQT3
BEt2saCOP7QRw5f4JD5PCF4WbSW2K9Lo/iLdT9icVNATioul6Gtzbws785OoC8jl
sKHZyuwG4sq0NEiV00U+Io2/f5Ihc4vr9td3a1kzHWUvdJBxLbYyJ0yBC2Rjo/y7
tARFeJUYxae48z/8XQ+KHv4ItpoldXaRPFWBvtPeV1lZXKj0mBF0n75NMSZH/9qf
Vvk1f5WXlDpuTucUkwTkLDFY3YobkH8RP5Ue8eE8TECqD2Lr6MRxcr/772pBCMQI
FupmmPplOfYTD/mQZFJmuujGg37WutvgpygD62E6y6K0cPPj1ly6NuZnLqZuxkl/
GOPAClSFp1Mubwcgxla/qE9VYIfhLKXQsINDb5QhM7/Ci0Z37celgqIOvRynUFdI
zcfGVltQXIRozMpVuMBFM81r5i+E/FRMNgUDJ+ZrW0L/BwxSFc5NYOn8vbfmo33d
MMYpxmxkx51qlEHlDdVD5urq08Ya8yesaolBOYgYi8eZM6SWoTL98Hv80JAiW+lo
/d62X0CNwu9z84UYyMu39JNzrI7RYzYl/mO+t3v7Vbq0J8hgoh7BdIfnjywfmi0D
VgnRXZOsickjA9tt19iExu1LdseyNPNI1iBbok4ZBhW4ue6LbAwAJOcZaPvMxih9
6Hi7Nwd/HPGKkFNeocWgdYIZeZ4G/y5nF/u6wIgVczU6eDR5tblILfp5ZERwEDZx
7Q0VhEA3vy9tsxQSjOG+hyBL4ZdgGMgDG1CDPRTGa65MX0Kznv4EGh34pi1omfHK
jK5x6YNzxSk3PrOuNDTZJg7AslEdQheYwbD6WnffYhGmyS9W65tin6+x5L/5Ht/l
eWUTbyws0PwmQC7f8/9LdqnoQY0dqf2SwTUvF4hWLt3/3yovPHF2B4zjN5l38un6
l9Zg75orjRwyRhuvqPt9vZESJpPBfUWIz0N7RyDtm5+tUkuTPL+t7KtMY20DwTU+
/EclsPDhJrm0Llw/VqDykl1NDgvSeDXCk5DMsb9AXisvmwmqxAkB9E+o3C5akyKk
w3RjPBzij8uFqYq/v8qT3KznMj7WB5mZowi9Ie9Cbi77TCP6WOlkpycQL/F9wxyd
VsVC3GkRwg9Zagek+ZyoCkcV2/4F/dejFlFb4liCSFDnY3o7fA6JBi7ItHFeodtt
0VdTVsPUqoopmpUksRdJXcRtIU9JjhyxghLX7g5TTmeo4ahBIJi4IkN5pDL5+EYR
aw/7/sV+gCJfObTYC/nLswiywzGbEKKY4UHjm1HR8EL1J1bo6XeUMPyfZcvV1kwg
8UrM/BPZg0XGhMp4uKezSwNBjcrpHTdajt4KcUgwxjgmMRk8VFRMXAyYNfrJxBUv
BUF2Cg12+tmfQ2Mwrjh91qSqJSL82n9CZduDEzIVMAHAIkv7EP1Ml9cppYMnf6sw
/I6GuUC5XtoQ2GJBWCZm2bt+vHoyZfIlih7UjeVRvzGr8Qrz0lrjEKumBpHeBP4/
No3G8RzwBfGueiiFH7YkJsFN0RSuDEw0OrhhCN6FHuAVNn+3YjlDWHKnZ5FmzmvR
eq1g/np16xlrh7dYJ2alZrdo6Y/C4GXUpVMEVX/4WqJlcb2Fs1MeBj+ub2jxzgEO
nG+oGPZyQgrrWe8wtPZdN7w9+zs18qTuFWBYupIdmmQ6L7G0g0A+MoXRzX85znEN
P7S+aHtHKpbvRcjXO7BLIJb35Ox3anPOcbNjOU9gSvkUylGgHqU0LgXOi6ahohLg
xLO8AO0tvRF6HU4xs31SPLZ7J7dmjqq9EL2moPSVsOCYJY2xhdRogVLEvwAhXycB
XJF6hSE4jXHB5fdIrvXHGDVPuPYEj2YuXKhEEvW1FZrjHmbnD4mb7OF25griScKp
2nbtIZ4RNEsMvRvf9irkKZRraeGlik7O7++pzn1+3WWvX/3NOClQ4XG0psUfgfc6
J7/jzqZrzc9bZ6c/cM9hi79lCOaMNy4fMa4luWV3cf9unOEYOuLlmdTktf5+kpAC
2wXVsrx1IwoYJzwvGMGIOYKAEQmQWz4VLt2AlIVgjgNJJ38geB+lT4Twb1+DlclB
f0fFV9WIG/wh1g/e1WIgVTHwwEJ7jR+3x9bL3BTBWLnYZCNqG7Fe5UaBVb1Xo8hI
a9CPkR7N8JWLKY4PaAEJc5PaIOTFx+uDkG3OO1Fpogwf4Rggwr9JE6T0ARUFXEEG
A3DZQDCevjIl/gI6/eRepzMxCQQ4iOfrRBjxFZLwG7L8O8/lMScjZc1CeSy/fRz2
z8OgYMBTq2y0kYzCkihqvcGQNa4Htu8RzslERk2KDi4Ib9RLae8LIs8cogKj3+d+
dFL6w51U0wwJxXe3MJr0b76hPWcAwSr6TofOIbU+tgZ9tK27bF9wgFLbbAn6Ld3G
zIIG3JxsQR4HZj+V4acqImp85ufv46EHrFD47u+pI+mfynLA8g4d/a0jwVQhieVm
sibD1201GOfTV+Jw+CO8kcLwSNUKtI2eGsmkAKqUbRabqoBbXAoWoggPzJ4NJvLV
C0GU94pe2AE9+wxnXL8qBuNLeSqA2qwvmDCPk46qLAAEqhsbR4AGoAK9lePBtbTL
31O/O00e/GD1EFYl1VBwPyrc7y+uc/r5tRbyhKspoqvdmBBOJ9QL2dnnmMUn+DON
Ns7c1vfo5ToMzU/Urzl+zCPksJVVb017kRVvfPdHFWtqS8IcaM3vOcM3fuRJBIOv
E9+IfEG8YHxARO3c0AdW2c41OgIuxineCpVWxIiAc4Iby5kmLIo3GbmxTdbru7qE
y/EKbNa9a0qFORzA+V8i+ml6KdvpqaqfNDZw8wz79Sbylps5zDzq1ZjDcDTUEAqH
WcBoE3SyP9tWmOzY2MNenz4V4HhVw/CKtNSohqdlob+98AyeE76niehaxq6uHqzH
6W7bDQOj5R6wRJaJatgHcVQZ5Oq0de93GWmHaim7IE7+KILmSe0y+o8k9aK2E9Ut
nPw4A9HdIMEADV2/0OiwM3orNRSY8YMFJ2mq+Z7LMLFd0S3snERODrjkh0B6vdZu
EaGNcRc5++pQ6+VhSyixQMCy99ntOmUqINMqCkYVU24lclBRbp6ls0zIkNUKlvmI
Nc5Rp9Cs7srJR2EM8/hJHWFl5NM8svQpvbpLCWHgd3SfcpOKE8hDW27/u9boZiFw
DtBD1oMnh7SQioSxp0I6AtYiXFokzbpKfexLGTg7j/CgTyuHClut81jUd7gZ0h43
VTTxn0DCyOyTVZ9I5pqGqPBXBpvqIkdxbtic19ZOVuMveKiWuOs7rTDMQgVIHpfy
pJOakmyYQsBm4VLNmu7zxkMSz7N8mtwl1NGOtLc7wSUD0MW/V5As67q9gvsHRhz9
TJRSYOCGtv4LQ00wUGbrVNmpw+mOoIxxtqZE2Y41G+Tu/ufl/o9yk4gZQEj1uUUw
svFtQ4QdMnVmDHWPOoK4Tdu/j2G5qbZaHcBOlTKVLPLpjo6ZT4Dd47jalcEqegRZ
tXPqmP/BOO6sur+qMh58lvKxMAxgu0p7JboXv6mb/92Ig+U+ZZ4CnHvTCp0cRRQx
xGj5x/WBSxrR+5TXBT+UHPTmLMSfSpihPxmBfd3DIF4LJX1DZ+fqnrr9+w0PgZoT
Sg2WriSgW4OZ/HCMFaiCFFXlBG96dGvwKcr5kZI/2+ItWrTfrSFpg2lXsM6QJegc
vt5dIpWpnpHKsQVQtNeRgMCzFy+Nvfb2H0qIJ6PkDUE47F67rgkH6p+dHq3F8Ty0
wOf7Jr44DhjG0+a8I/Ll8jHcvkR5YDebZMde08XWqB1duIlm1N8ZEJDi6V1Xc4Xe
jG+lXsypR48eByvZ2xHXQWAigXg2rXjfP1ZaRXly/PKXLau52O/iA6Rl5mbqKlR3
f1GjwQyM7n2cnqwvaQi6AqL/KQ9uoW2GLB3YYO8eng0wPWOYl5Ftdh0NMierSxNd
+Xjdyhx+NEoxlOfLvhyW5kmSzoVqHkCRr8OkRXTFI/E+5vRpBj+VtK00fjBD4O+5
H3+i7NUjPBnVcs1jWlxtXUyqndxSeop8bHy6fjSvRlUDSM2+nCPkCjihZlmaNomk
1hOqCMAC+Ha12+Vb4COq9DluqWMJdBSqVqNqhOrWkI7Cp5tGPCzZ2oaoGo7gITSc
58ueqaiSZiju7aXpaPnd+ulto9RVXZCPA4U2bOC3FdNf2UxfQbXW33/4AbtzuCHt
5/cWpxTIlGvxNlub5Q5Mp2YvFS4LpRzkhzznThEC3BcJoYQKlzDavCTxWUG+PGq1
CuACENA+bZpQYw8lfWZI9VxU2t9RlxCyE0zUrSEg0nhJIsijqVSk/1dZeZXn1dgc
J/Vfm7tHlWkPgCRXE+g9CQIg7lVkefP5EE7zuNm93eUrOmxB8A+LWINHi0MicsSa
D47xTig0bOciePDoCzOUky4QLHJ9e8JmyueV8IUAZ1U1x9Dr14mLNUmsegVi8lVC
Ce6H+c6edbVxRJw3ukFHlvMGiN+Rka4Rff1bltg+fIvr3hHZ1ByTcAG97HIsMAiS
yacdfp2vgdJUicYCH08KqE/pLfqjCYxCUglke8SdCpI0gwFu6Fo1HA8rqrrwB0s/
MD7TWIIIJEqeiJIBS7BzH48O9dHNltfRXmZzsUEusu/oeqhx82RvX/qcR2D6ARy1
b8JpMzG73kcjIika4UHJiIn+rfMpbaH+hWJ2jpqxR4vq/0wQxvmh8d+R1l5MXaye
cSKCP22Sk6/+QTSNi7SwlUWQO2ucMf5nucYaBycEpgcNHivs67At2hM1qNdmbxYC
ScwteYY0m37meivWp+aTpEEv/MpYfqTP/wB5S0XAEW5xL6yoL0OhdRDKP1uXlOme
yBe84Vo8CelJLC1enD5Q2qtp7Bp2Wl30x+2AgzaCLivCF5V1+v3eCuZJ26PCliIn
XAVcvlIZdI/hSnZ6fHVVTdWygRIrtumovOSCmn1CoacfftsXzyi/c7F8H7sAJUbZ
`protect END_PROTECTED
