`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MJocWArO5UDRh20C0xq6n9asxW0+Jp1neXSD8XSeElR62Hzvp3LGY7tJ5kEBav7H
ann5tfoqPZruZ64O5CfoeLXl/+CEwNA8oeZNwtjpwjgGOKLd/toUj6mp38fS0GlY
J0ZoX9scEhNw6BAvHxcaSUAKTnxmJVeJYPd3ysN70C4x3lDbkRX3qtnm0yT5ZF8W
NyYCnuAhCX1jo1+n1J3K9QCo3D9ia6iNbUGrV723iYp+js+bljYSB0gYLihm0vlM
gUsMSkOjdVIHAn3TOnI836lWg73Okpbu/x1pcw+YHJH0jJl4e/g0VyJW//c48t2G
dZLNIh0vjBEJnCnvs8dc2T+gOxw/Q90drcUyT56+p2QNyYrSPvKbcPSqNXpOrrc5
djbzc1/El8AInr6P4OtW7L7zzy+loNfyJ4ZJYUVa6iAxxXVODIH3IqDItYHVgs/k
a6jk/Ggj8iBsh7/MYCnji9lcFH2PcPBm6Th/q0Gf1UidtLLJI455EN7ijNEfLABn
HjHFj20x2y+TpAO3IuuLxUuhCIf7CVVqN/6D8JHDs5fulPBtyeSIFPYSD5Hl6cVJ
aSC7xPtL8T0E5NTPMfWmEszANmVIspoV4Jxbjexx7GpLcSlAiRPZFnNJ4orRR/0q
+4qtypSN1QOIWq4AxVtv+WHQUsDyr8E4I0Vl2q4qTSkQOb6MLaLKZAu/mD7bEdDa
1q93BmS+/0gikbG5ilmxdF+s53GybXvTxe/mfb2p8ecWc/9uT/zLrL/XoNvnT+gS
R+MTjxWD+thaWr82RGokn8MlVnXH33v/xbLvqZrBMh50/mRibZUXBiwndFk+dysB
csXM+aG7UOqkqa5cfZ1nDuQtu39XkCDewwxx5GGugjz+psQ4LzykJFk1i7dIH3sG
NPhHfFE7m4T7BFG5PAJ3y0DTCsOy4udxs0VjM6Y9kmWI3tFsSmhVWFmnUHmlLNQl
dY/T8OPb7yr03BVbCRSqyxdK22b5jyC2ibbRr0rbmzRKxq0vdkNEZhMpa/Nl8Ihi
VTnkv/4+PhNF63/Xs8YFv/6kWbzM4BNzLpLN8p5T5YawcYXEZ4r95aJpauk10hft
pbdnrM4B9P04+7OVCjA43m0ss6ycamXrtj+gIWFTMWRguPWu0vpFIvaYQ9FCs24i
kUfoA256Jhoq3I+i0dXLWYhPj4L+7uFyJbRppcaXw8iBEDRasQ2bA+9nnOj18VL1
ehN6jaEPckfFkQS77mA1TivSxOrRtCcuwXlytt2F7GzFV/aP61eUDnKasBi262+M
8g2RfX0aHREnAYCJ2vyK2gAYUh2S7m06n8yD6EACwCfw3KQRrYECJ1yNk9tFFhap
+gNaH/ksBVyWDoyY0HzMqLBjUXK1luLckFsaJlEtGvFeChqMdYCelW1hqvP5WUC7
JvOBv0n0yfLBjGnbH7Ky/qK5xNS3We3tQ49QhmGQsbsGzllk0zxzi3wre8b55sTP
6rqZv2MUmwV+6Fa0m0POMEDLsrmMe6L7JdPtyMZ2gyT7Dl2Hg7glpm623dwxEFfM
AMTQnPFNfyE+TCA6aZB45zkHvTCvIOWSrwcuCLzCxADDSRGXC1+gTUOjIONYrrM1
GJmrA9CA4o7XxyHHG2k+TtH6WCGJZWoXec1lQEcvRxWUeML8zNC0usPaz6/AVMQJ
yMfFlZqrWDkL2iz4By3LdKRPXxUH0YNM0E7Xu76cl+SKJWFCktqr8yrcyf1zMkOz
zJkHdThHAetotbjee1t63BhPJgvbc6qgB35M4T7zKQ3ZWOQUZ+ooJKu78J3trMnK
Cqkip61onmbWiITQdzzuP2Hs5LcYtLX4g3UJGORVavIiLMd3uIJRgq3zXO68g41J
k5lp4FlV1PRdUjUTVT1u+zZMiq5od+NUBdHJ6IjtOePmYg81eL5zXQdglWfYsQXL
CzUNOCuT0fV4E8EkiLjVjpaNBeDuiJUC3/E4eu5EFHqxI+AmaIyrCpfCGJOh4pCc
ZlUFBftJjc19QIgRwrdcW16qHJXlKL5Vb/vcG5qb3HFoXIHcGUZDXTbrKmhjWl2f
ETcSuujNf50V4x8SBXgBqgbvIk3fIQ8G4mRLmG3Icuu+3FiLG2YVR57B+OiXnlR2
2+Ixqpq/ueRZ6Mb2NmkB7EORyBmjdUevA0/yp0lJO8kI0QBTezTsErOXlfqiR+MJ
coIzthGMFt24/J8bHmbl0W8D5MlmSjdGlLQJzDoZEw8zLS5gQirYulRIIje27fDn
9EAlgOnrhFcXYVOG9ZurzR7v8C/eHeWbUzhEohdwe0Fnf7fLNQtpzMA4uLpBVxa1
Y9gP8UFwE7VjUauJLn22d/ae7/t4+7TkXYdlmRD57qTQuo+Q4743qSaiARP4HZOy
YFOAiQeRdYSZn4kCC8lCrLUCUqO24m1TIDFvOINkI+4CpY3m9T/3asD4ikAMygWP
DGxdlm8RlW3EDmf5KatQ8T0WyE2NmR4+Fz5G11SkyWyYsp2nATkaXBRc6znVE0tz
1v4GiBZGLO0Y8ooP8RLqce79BcJRBiO/dTDAKLHgXCkaeZL4DAz0EfGTvldiOZs/
3FPNNmfi+GcfbjKeSMo1fDrB/bSrzgyRpOIi56ZRD3JY5adktoFsszkGJOYkTCkC
XCQtP6w2NttfaSU4Wbv7jiBKxJ74bWfIym0Q3coWyViEsZmj/eX6hGl1/U14qVtZ
yqnrLIh1Fa6D2W9+nNeLSB+OnqXzQYMRizTsY+iDqg9f2xngJWtn8ASusPupjHaP
TMRmSvoyT71k4ibC7yEpbUj/dUpcduH+V0EC/3jeBa8GB63tSV5839cc7IWhLKsx
Otw0gM87tqc3cDazWxNH6RCMrxqWCDN6/RC0ae03rMjbjzNVdjsWWBzB5+BvsgRq
9Izlu6/hpmYepjon44sbzDoBH9HQxB/AO2pPx7WDTWwCp573szdEiIn63a563W2w
2idfgcq7j8aSk70S1/f9KAZwmBUvyA7UORFutGUer8PmNA3PRYxBoFhDNp5rb/oD
boZB4LxT5WQZlTbilwavARZKquc/bxNH/3JiaIrFrcfPV5vIQijQ1onqFONwIlo0
3b9KrRjpAMWvHxpsPwS9qZBrGgaT0cn7mbrUcztQPHG6QegBXjsbMm0x06y/XRGD
JVAgiXlIyRAsZorczk/BV30sR7SQ+4SZmNmdgsg5zodnyRYFiLcjAxruGjZkBuUZ
hPC9pXxQdNGdXhtq7/EMcreA1zjv7Ak0MyN6wKDi2G9Z8xOlfstGJ0wCUrsX8lql
bf5YpAkyEmbmX7dPewRjoQEDe3TlpkNvjyZp75b/8pKz/SaQJVa09XUozeJ2csYa
ZuQJI39xSeETlz/dZU2ld+Aqh4AnwZqYQf53BES0u+0Is4VZBteI2LI2KtB0cnmE
sA/eAvD335FWe/0Ngi283fmOrE1u+ScmuOlxCNqqpp5AP/RCWxXZyTDW9OzTemKC
flQMqhoy24evAY/61UpoDHIEZm7Amb0kXruDPW2ajdY0AkPEf82UOGqTTg/OIxmt
nfleuhnsWs3r1YR7k20Zb4s7DU+if3RS1IyRoBzyS7H1eMYGYS/pzTIkLDY7PoKE
/t0WnsLWy1p69/jKSbQ8kRu2oZepDUwcunQrhKhpeqeox8BdRNNnaVQQSfgPzaFz
2gKjAd/S4u5PyKwuoyjZo54Dk6UEXbGbF2MGC4MsG33YFN2ixkQC6L580/mViXwU
9jf9lkUk+6zR73AFcruR6+eIWfRrsEIcTWtjXDCaNOnYcnkwd+Qp1Q1eow6loZKT
LVgm48pNRPibx942z6Kzb+e92FARsmdn4QCFL+qF7jN+xO4kvGUnu30qQF2Zt1a+
1De71WYHzLmCJsIuTJFYsKzTtbca7PTTatwzj5cctUW9ccUkkMytRA73TaFWxoOj
6mMNI7aJbKZBqexq3x3/B/eEJyMDCR/5hk7RIo3fKXQgI/XFbTwFJxGLnh4ffZ1O
H/rtWG1pFUtLrvsv3wkK4JHF5XVgQ9JoyoqMVnzBgJcghVByeeuZHA7QgrHuyB6e
+sC2lLq2veXXRqBMSo7TQ8bsHItMepO0cQrPFtC/+b1s8ma97aWo4tkViMkz3Xoh
bZuEMqlwYykA1Q2TGWntfFtjA4ZJ/kJZRGoRt3lqufnd+JuV58t1Z0qgSIuvBR33
KiUX+DeEBPaMofQUoBpC4S3pXjIqSAsetxg7T7kFVIjqxG1ahgtZiRoWbKQ81ui7
APBzAxvICxxqW37KbOufZHQFCfRrYTe0+xlxN6hrNEPnPey77eUxSCRMb45TQTCY
3J1+m17iFnpqk8QA4n7aywxwl90ebuWKsk1mk1sXo02m9BDmTUxmhf42l0/80lAe
IoD7TuokI6h0e6MbXYDsb4EMFbWx95slwhVwS/zCS2Z/pmdYiXU1lJS0mSMg8fAT
Yh2t9aHlmBAlBCTrBuMZr5q1Bz8iQJmvrSkSPSERuEJyBbpcjW4B6zl5bm+GE45t
WfB7iC3g7HpCOmEm9kon7+pu9B9uht1Zc9/gL1RprQiAO0UGSAS9T993kqqv5+Te
pJ5Mm0CSqlkPpSM/EgqD2A==
`protect END_PROTECTED
