`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9arEb4dM2ucOgp1Ex/6cSxDshcqclNHZgJwhmxxBUurAcByR4r3GbxkyEIBMiNeP
aAQfSt/g5NXf+9ougYfqwxArQM47oyidqIgXmR+jUJzwFqupO/lHalhF2ft79GIr
zmjdl/BDRROuKIM2un73QsPFJY9BPJg6tEEVLOj+RsNc/DJ5oKR6WdTUHhpNhEE9
i40jJDPhV+7Mas5jeSMIyvSD/PpzIAEdhFTV1q5w4Z+nkVhXtOyj0vqtdK0luweJ
q5gO9uNoO7fMXJSOfcEC+RIwQ8bTHEKfCRG+5GiJG28Ba7eEv+k8Z8h4Ue01pbvE
vZexxysA4DYnZeyRbnQfP9nKiCU041pGkmCqsw9g+QWGUJdepIKmbrcelkktiCTy
`protect END_PROTECTED
