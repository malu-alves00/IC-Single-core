`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4zAsooLpzazJVadAzr3XQ7w+rvTlXvfzPq+b+K1X/alStDSGcyJcDfkJtw9br/Po
5paB0SV6bzN2X2rQUM3E5uNFAX4nqJx05Fb+gXtyu2JaS4pOTRRQdwTukkDiFP1K
OAwdCgBCvaVbBvyIba8f1UNc3Rg/FmxGGbxAzyjmfnZLlNUji1+q7eCRzk1sIIWk
9JOVON1pZAKOQHZ/umtJzSMClcrsD8Ukd9g9VdVQv5O9Ji1ki5L3cfmTEgDIOW00
iziTwWPe00sQEhhIkqeLLhInE6WYLTS8ZfeCxufu7rWHq+6IMLpn/v+aAfCCVBLv
4/9QVNbtALfc1036HBgqnh3OmFU8atxpzvRGJza/Dc6tbD+BVtQp5ZkvlAVIHvsp
BIIgTXhr7WasHpw7g40cDSXrnhbqEw3/ONxoBmtBcKs=
`protect END_PROTECTED
