`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RaJIkinvkav4P1klL+wr+QhDiH3DE6ZdynUyr7xdwes4gdeDMatKMSJqUlQGqWbZ
KVvuT7ZHVZz2zCOwtRZpbGCtOV8+ZRcLxU9bnxqc7GFailYHHrrHovPMzs0tS5Oi
fVSnXCgrpw8QEbK+aCUXGiX0YPq/joO2rw+GdXfmVq78bts/xUOKflAUCq+cF6Mu
N51Dtbjh+/kgasQni/GLqh8Ogli3yIfPx+uP9hrnLtjaFiyBASvLO6190ErK1IGC
A4Mo2c70i2vQnZnJUcoFVuNzK3MIQ4muiLb1/tWudrmJ5gFk7/qltWuW6FzXvtZ8
wl0hs5bhawx66TGMMejWd3PfYqjR1om51YGbmh+X9Tdv3dFEMo/iG4Q3Ub/+swtc
58K9p4Ha1O6kV/RxFRUFBIs8PvdJLnkW0swIjsHW9OVIy1w01C7BMj7IeEKSO3aC
0fiCldigPSdD07EzD9AVZBrc5xlmrrDADtT++oZ3buSLg0hB1zKYgUf2to+iRtCw
Btwd92ULZdQzzceDFSIbtDHcpiIp76O45Wh2YEEfV1vwtjEb7fTcg1lbRE9LqTFn
425L/fYgyihNeS5uEkLW0vF/Xcl3ltpGUnAxSLi4iFicBURyxrekuUsZsa1ShN6s
2lfsqFa9epDeEXQQDyJlu8Gg4i9KQSSkPHLyJSd8LKiI4blmLo5gEXDcs6AyaNky
JQmV1lFBXlLupqWJ9lTFkUWTj9DhTnu+4OJHKmFN1X6gQL78395XrD7PwElCNGGc
nmhaLx9ijEiMvuA3c0LUgAA4p7EOmp0p6j2/HdTAzIBLZeIcHUX65ftVJgfRxEBa
CJMVpczj6Hn99Zx/2f9fiT8QsdXDh/QpDWUAWX4qgjHk6spWKzn3ZElHN3SiHyy7
`protect END_PROTECTED
