`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
a4Sf5JZzxqTdvCTq6c4wgs2+qpAGE79SaUnGYWRZ9sqp5DgeOL/1T+IRAu6ZO8/3
Yk5fJwfEcb9sHrIGJPFMNFs7jFr/Q02zKDGNNK1IFkASPotrsxPow8ZQkkfi35rO
+uWHTeK7c+oshWFIvACpoHdkJ62yLqSBgGmhW/H1CartPu383+YxnHa3YHHvzVS5
78l9YAJQKWeoFZJRYUW9iHoDDp57b4iNX+KQMN41iudO5ZRvESSzUQcTnKqpVkAM
2M7/cRHxRBAf1jqe0yw7LubJIgZ/8BGCmWftYWGD+XrZaeBex9rZEmUFJAK65g+I
YP/ZZhTX3V8wnXkS1gHmjb9Wi/VS1V0k/h0GNEnkWY2xZMHL7lL/jTLYzkJpF/S2
kYWD6kYXkhSNOid4LKp9YhFkYroQdpOCAds76DPFgknynQLnPmRH3YVYQdUewrlg
Q0zkaOj45FMWSF02tiHwVbSYbd/YtwLsjSQFT9ZE/dYyubkR4npTR6uEHe7/vE51
IEA8kRqRyCCsRGnbBGyhZQ2CbvatIu/jzdcix9xMqs3xhKL8zANw0WWMbsc5SEyb
ShMSr+LjSF/rrBObqsej5Ncyj0jelQXjMfQZEWpSDcrfnpJXEMHbXTXqDrr+U5ky
2nWUtFQ4swdIX1HJU3xJ7MHLd4rmhhl2SDbIM6s4pWOLpdROQgNFQBUhALd/yO1J
XN8jbcrLp8N8SRJEI+920CwMnPXJXml4ulqWi3IzYEAMd3rdvYZU/McKw8/AwCPs
4MTgDtwV2aFRMQAih5siwpCYv4PDzt3qUz3phk6Wj3ERlqQt9qPJD4/3u2h8Zbk4
npL1YpsTNAczXHEAKwnVBn8rlf7lM97KRQvYPi74KEGxbpMU/tVUIW0317R2Ixvg
S7K9lffGZYjPX6Du5IrCl57ZGQwsfsCWZmDU8IUbRG1DHEVJSykShyjOJLlyuxs4
rofrMljgAdEOZLteE0JBZEDR+PPFyed9gOGPoqVVWysSYARAlQFfaviazkWGtYDj
MFubiQqfBQsO8eyl68kcAjwmgx+JVivD7CjF9g+1Os3pKcbEeWq2+xuzSxcc8LsS
Zj77gYcVibMPoyb0IDu2Om0qM9zeKeIqmXayRcH0LjQbHtZkRior2Wbv7ydw8hvc
VyEndIDxfy/jR121tcXXhNpz7oVQzVvpTKAmrhvD8fFcaOAnwrtjKQdmZdk9NDqi
jnFsG33htYSrdCZeLinx6qJ5mbYMh5KSMOhq7jFBEoOB/G+is8M9oov6O4GmdKbs
W3MEiggh++rSxtXkEkXzsfuysSKYPLkztXdrg31Q5ycCsDmSOomjbZtcciCUpmPY
hqpZf5rBFgnYnjRZ3lgYg7trR4xpZQdGsIIUd6FBG4l732DdP7qR9sxANgLAkRGZ
ubWVcyLmUnX8e0abDGgeYBAHMkAhgiIc9uAtHDQst5CLWcI7+lPcGE1tGpJvD7a6
vYMdLl+jquiqfNeGJHLaOLJoWy6l2zMW1fdTqQp4meQoaQSvrDAyUR6c3WVnsj42
zl50j7737D4c3QHxDjOBTQdiP0IDEWgP5zMs4PlzUaLjU0/W3IkTbrbg9egsybX2
raM9t9Qrhn2atsnrfAGCJCv3mYlsnhBwMFHdWyb9uwb+6bJeKyJa2SJX6QAFtuDm
ZbbrMJubfYPSLCSISwjGhTKCXC/4D8W5ler0qjDFQ7/SNqYZS/RURa8t8aHJBwor
/am4bVfk4SZcelxAWqa3M4D2EL1MyVgKi6ofDxbusTWQAlhcnW2onEAMwnv6X7Ik
+5/g7Cc1jM691XLpWTqN1lgC1v27DNILYlWjInjKDp+KP/0v7c6gIOA4+a2nj93R
RzXkK0z/F8Yq6DEcYwVQ3H3GLXAVRxGaicIoNrT3fjHVeQ94UoSRnQeMojfsat52
ura44+5yRqLcjW6mVpuLefAzGs4V6lhK2+OBk6DCUtkSlN2FzZcdWSLzfVSRbZNI
QFIC2ipD8ma5V0BID916fgCWT+CQm6AzU3h9lXqVKRmXc7U6WC0VFqV+RZqV6u4O
tbD2bRY2Y0s1bMFgQqhDl20B5qVXI3Zfak4c5z3h3BkDlJwjwyDBN2FasaBblaMo
6XKPyU8Rs/XsHSS04mEyLTzh/DV/ji20s+Q7QL5W3pBeBNonVdQ6KjtjBEfk+ga9
Q13SFqpChfyP1PrE5H+ll3DMPYcFleiH14EqTD1GHm6/zI9z9uNSQ4onoz+X9ZAw
dsVv9jlECmiPFmV6kLGqQcstRz7K+FeRy9pYZErCaXHl5Rd4sgNoU1M4dpQmmPXP
8vRlwRu8oyWs7DGVChKEpVQN9padSk46p1Drtpja5yrX4NF3DXL7TE8DyDXK84ud
T4CA73IXE+1D4NyfStZ90S4uiP7UFfOzfmvkinP8RiIa3siZu/EHNmd+BDH4AKGu
9xaQ8JhqFzOtAZmPMuwM0MBZEHGa54JM+NSL/URDmThIrG6HWJinPqS9EKF1ITRk
U7zUsBan9+jETHVspnMg6G9UCBiycHOWlSHTpUXsiO4DqrkhV9OnGra7ShNYuTow
D4EzYpLRHzsK1WuUERtMNaph+S4b+kHqDZae7dY2b3ahc+AjM/Gq/hWFWs5ADHgS
CCaDotM8IWgkADUAgdiU/zRADn8A6KR4hp2FILvZw/Sapf41q9mHeFGFJ0tJ//qL
4Ll8pVFkpcVimx634Q9FoE67qz5Riz0y4DZljikwXMxQ3cMB+/7ZTvWSlv+iEkrb
pmT+dAikcopXkaTiGsAD4MiKjRsQ1ytWA5JXqGcfa+sITyHWTnG07B3+pMGfhKuB
uRuosaCGSCeM1F95JlWe3g694hyxv8K2Ie1gowsHPhGwTDh8yAIp26GCI/lH4Ats
TWcaAI/yybGxJ8ncZlUuAQgggXPVNI00ndHnyvfF+HlFOnB91vASQmHmwBX93LI+
Js0rcVfl+KEenLpi6aQSTjFHIhovNazIyvdzUzKIz1bIV+g85iCrqvVeB8S8r8/i
D7GTt5UtVmdOW8ljlFkClXmYuoqyHJ+DyAn0tMLc+Vbx9/DAL9YKbQcB7vOuwTez
Qpz5Jar3uybmVsm01FsO7vBxdSwNUHAwIL2mQx42NSxIwRTPmfeLwncAJYXxM5Zm
x+Db9haQlmZBXxz7Yxm5y8vzmFqDIXx+rmmBb3xjZ6S97jKBqUGPu7piAtiTmqTt
EYKP/N6q5OwMt2Pv5yoGnZnK0Htolh31eq23TahDVODFZn6KqQROGcE4f5QKRTAq
+LlPcBZevdF4lPnUnZ0WauZke0+HFagP4zvVGIP5NZlB5IEmmBLoeFOMxuudmgDO
h0vJyl+dq2a9PxSbhlu+C5/SVLqJTFPxlgca4yoNptdcvx6yQU46Rg6bY12IIHOV
gNkpzlFwDebCW1bXICdlVsW+suOslhDsDGjBTFWH3EokA4HbQA6p3PGvfJqb1mic
24jGHrM2LOgYeiW8ryMybjN2/hNmIKglUR6L/LQvg62VRXv2Qrxb0/x8ttHupMhO
1BaMkjCxeQBuTKsIBZ98XyhiOC9kS+qX/e982a6lc/WE9wRzu9hgcCyHQy7gy3Bc
5+kXy2NQdVhaFcDSxFXDl5A4MWjtkYUCpgIC68gbfCNPkq5sCzOsZaK0RwJ0LhIM
Q5aFn+swsM8ZG8ksytmtAbDtuE5+VJXEczHVpTeNJVTyHkOKDNkTQua2HUsv8wsC
SqeWz6UPE8QikF5ogeIndleRA5uDcj6je/Rxjx+C8ijSolYpANXJAMbGscmziH18
xs9nUE3PHbu8+XxJa3oHuE36FQGBWJkZvDX8rjC5l3oENbWYt3waLzqb3aPosNeg
LMo5YJLK8TSiuc0wEAYkB5QqKrKJVOnVghejpRWo+wWfZ5Pz3Gvs+3mJxnqUKPGa
P7iiKNwjCwAyrZ3iTIbVWyUoTmZdwOM0LvXqaqRyA7WQ5QpOEKrVPZvVNvnrw+qf
6VdriTp7YQxBytkYLorkVJOmJYgx/C6QQySZj2RNtwKYRdA4z2LeCgCy+Mo2+TAD
bbzkmQ62/6G2uuUOWiEqfrt6zzkMJb/EZswRJyiUCMlK1jsScq1IbLuvRRsF6suQ
78hH1ZX2n+MV0jvDTK835fbCeQJVuJy3AWbHf7NxmdGaeg9RPpHYa9jhjzaz/PtT
gwyLISFTtSZ9lhYewjXIe8CQw2kpEfeetmBXCf8xPwoju1zko83jSP2AdtimebjV
9t9nPB1ZV3RXdgntTSCzYRwAJSUCb2/bvhVIWZ96w5EamEGsJYqTlgznLdcPo3hh
LpTjTmEEqwsvcwoGNE5uFT7aOEidsBQqR/vOU3QIyGAnovCYByvw8Ept+9jK5hrd
n882k6O3dSRT/qHBCgqYwBxLtv4Wi5JujUTtbYR2ZeGgiSilaA/ZzXaTkSQHpLjr
8nDe1CFhtssZUgQBdb+sdweDYZtjy1lU+b+glzI47Zm/kgTp6Wvge0UhD7spk36q
tEYPmKN9B0a8epWBiwKEbfxfibPktFTDpQovfYCMtXfFUWEvv0pMf6OVV6XUiYJN
MC+DoTTCaMHV2iNavIszSLXnKHOW1eyTh7QrrFJcOt7hQr7iaXxxKjonIUABrRNf
emEu8yTLz2FhJwOYRUFAKzwwYAoO1ePhWPaE2AS+RtabiACX2lY0CDE/5XZHUUvt
7fWCMCF12BwDkWIP281SmZCUylgLaQq1u03OU4YAbMhdh//F+8ciO36bP2n+rzYu
058v8wfYtFvoCJ+tu7UejvvLBiH+qeGbv/WQTqAE7fSorIJxYEOYqF1uZ6Qvl4zd
y9/ArY9G23u4jFrSske3ep503SD4Rr1PIbZd5szlmW8BEcDDrXIBV6x2NRbVrP9m
N3CxGMU4Mj2U2HeCvqyUEOjONp0iJiTqhR/ikh2hbodvCVc3pTASzrimLabtMLcc
yFeIZV21w/QjR7nRVfduWWug6/MzaMpGc8r5O+htlgTUy32AmVzKut8OGBp/vvYB
WheRz1G5mpSwU2kiFNbPJzwdo87qPMbM1YYD7rkTwxVc4fnw1BlN4KlQ8yCXO4nI
RLwKN00YEYXDotQd9O74Wm59bSIZWaJ4mWGBgw+y6iXP6IlS2rTNsLn3+3pReI/0
aDUC5TKusM7Q8+DWS45FKefNlFIPrdqwyDBmlwGRYW4XHyvCkRZ1q1uaBHOp0qOf
XXVbwy2+TvYhAY50ri0d7zFGZiQ0PXw5V9bSI6xrIujLJuugSzoEy2VbOGqjSnmH
fFv3QxKqYmzD4NXQOGPkDUR0xCccwTBDnAUpUCAjK6HFbWQLvS91CoqUc09M3RWz
CIQpmGtyHEfydYcbOoKaiNZsDz9Acd/0PgvNByq8XuNXrIH8peZpp0xfhiQanWGz
cfz4/S7YcsJlPtJQTLcrL/Are4oeKtA4M2ZaacsbmucpUS0Q85RfZzD3oMygxVLG
37HJMhAnrKcujlTR87bGoVGUqHUnzzy3x+5eYNCpF1a4ft+eeaFubdvWddd7fW/K
DWUQZQaeDG7fosFcnZcMJGOITvnKAlSC5p8u1HkuaQEBmYZyrmG0O+Mkd49EefGG
Y6H4qZvL1B3LkGEscdFC7QZb+T7CVOPk3ryOR6qd+7Ws81nhF8dhMIlj3E3gfnEZ
46tmjlFz8P6/3D3TmVjRfCICyMb09JfNr0Rj1QgiUKbcgvbgiB20GwGWqFcNy6cx
57Us7Y0hCJadhGaGGki3PCqLuEe2s805ZLdICi0KXp5mQ/XZaZa+yxwcxb3y2WFT
N7t/KUDhxqhirAj1lo6ZSZDhWVDx3N5htklTehlU70tQj6/7vnc2o0leh0C6G/pM
Vxo/E979OnYSzdRRDoybSuflZX+3Y7g37y8B9V9LHhhv4wt4SwsSxhmFc4BZY2/u
yCIDr39HCxSzOxXq18w5jdSku/2ZBVmVOs8lwDGNVIzekqlt/2BovXYS48ZtK/jb
rELhSWp52U0ANf+1wTFJUsdQsESWAV+vUCFAqbOWg9njKfsqlvfHqU/HoU9wyqJi
f+CWEgtssd5dEhY1VcIPX7FHIcBkpdFD0snTzz8eBaGoG67+Tsm47QF/fhxwWzrQ
PmjkA/EI6uzOMpvo0jEI/dbezodAKrjXnoVpmRudYZFr2yPzK/U0c6rgU7YtXPtN
jfkRCvOfwtwsL3ykR9cnFXdwwRCGA6YPCLXG+FWHRZdKtBLxm9vVurCyJf7MX9j1
eq5KEoypMzW7yujoF/RNGvhcAgC9vcg3n2iQA3dSFEVb2m2PNWfd653G9k2jD8Kb
isixHiu1tx8xX9Yo/ndhF7pZGMDG2WbBGBNZvcPjymVpQhao9yAxPaw6yDWtKLSK
EZL3aDOXjQ607rCbvINourMuqdih7BuQVor+4AMffNtqjnEbVlTfZoCcU86dB0Km
JcpqVE6XjBCsYm2KACEZo8Kxb3q/ua0wUj4yFoiZUaer5o31+7RfBvqi/iIIHY6C
ZsjTnDpPtnefYrimqku2XrV8vPhpbTUpz2j5tmibrdwIXmBnj9KLKgIQrzCEJnD5
W3V96msYGrBUZXwB4lzoZT0E9wu3jhVcP6qlJ++TktxR7bmbKGHRAvi/COegMqb9
M54PRqPSmiuuMfFeHC10DX4jnPh8rRp/kg1wG8ona0B222/LSgEGOVN1RbLjSOP8
mhKIA+tJwYhkkCHUaqGOqpjwfInn9Rh6d4ayMewTQ+v3KKZx44IPoZhYWeQfxxyQ
bKRwrlpRF3X0exujBVEKQMeyJ/KoTQKxBdPqXvb7aoFSQHMNRZt8RNzVk/R+3BsH
nrUhzOXLCkaVFsUZRbw0QH0a9D7BbTzrkPpLklHo6lqe1EQ4vjljTt/O1wJWRiYy
LGmyWlLimq384HpG8rR1LRI/7cFei0vjWU/oImqe64eWQPFMTymT9aYOLJXNf/Xh
5IBBUQovoWSfNnv4IJZdVytm98tXC3FW4wFvlKPcOAPL+rrReZhP16YDHsC1QqE7
UVotFVu8sao2IbP0yEhaXwYfu0g4R4xFJyZ9oi3NXBz5y8OaHrozOVx8HgoAcK0B
NaO3GbuG48yoG/s0qqPvobyaTVX2onNSzBqexCgXxfeYuDwn5DoMW7uOOYU4wb++
M2x0vuas2NQeWxG6C1clSrTF+HTtlO5jLeJzB6SOlRecth9u1BVSimLHzCTeHMoK
kqXxCuIJ9o2AMmrdX/oHjvrC4MpMxH9xeQgRPpN/zYMeS5SWEjRfUFx3PwwX1YW2
t+xaXhXargtFwqgUYq3/kiNTDxBcpL2yepn00QhOQK7Z6W8C8RxOQaUnFQpRzI83
2HRle7qHeWXdLlvw7GtR5xDZbhxMxnk/jwG8lK/TLFrWDkVlnW8WtWyNQbzQj/YE
Uprd80Zwj2Z3MEP+Z5u6Q+g1uhryQRGTKoAiYQtclH9UNR1XTBsH679uCEoI/zBb
ReFBJW1gmxvB0jnQGkieKY1mTM+kWlvyHHWGZBBs/qBEm4I6yIXFF+K58MqthpWl
w/wwHHXVhUh/A51NmvM6s4xHPW64BAI0KwTKL4N6bMJDmIl99rFWogQLsae9Rq7g
+30DcHHTvxZf0Kyi0ux06J2fBlddTS+3S5UJGSR41dsCQH9cFAO10soePmZtORMX
zAMqdjhFMAeJGyn3Nnw21fXnLwug4mc72IqgVfvOMYQ4F6a8pdHhCoj1rOoVVOxY
oXWdHVQyTDZlNIHR73ZdWJEHW/7G9yrxRZy51emY9H5chablVt8ZBBD9S3OSRjSG
MzfhCuRLBj8KUVLXodwxAJzUxwnYNpmI7rwKpTRwgF8BuYS1S9QPkOjXM4Auwmsf
TRKxgZHOs+sI0TyJHOAy7PM5xeZjp5txVTFxOX/bihK1b94JobGgMTTFPDD2FMr6
6kxLQqFiSQrGpCUspvp+PVyz15ndmUxBSr+094HYT4DMm57mvzZfTyWaGymMt3zn
di8paei+il7hF+YxL+DF0+usRRCyiPDe3ab6OOB6vHfvdEKPYCjbJc+pMLpmHQeo
bwFY2xH03RW7AsdJrpMDHvMtqSlkPfYNhK7i246NMhKgofHK7YVM0cfJ8USy37ux
mBRZKZB/QKduZjD7FIlMcFvbw7J7rTUwdUkKAe0Zc5R9d4J+0t8jaX+2iGuZYw5N
AL8fp1h/jsO41HUZGw2oFBtfN1s4pmLw9Od3OTDJx/qE0ln0HdBkYD/6T0AmBpP6
nmKWPQ1NrRIjmcfJdScTYgXiubNoieQirn1PwuSJCOf8yWWNqNGVEOFX51dGZYsq
R9xdys8dgWaslJfXXhjsR8QbMhjoldEyBkW85se/KrZLYji3Aca0uBS0N8anIO77
XDQNV0azDAKbvCZvVJCGdYVFZ9WAIA7o9HZoOzDhtK0YLl18CDeqR13mE/u8GeP+
fmFJoMG8IyIAYRliwRQOx8ZViJMfJW0500b9+NL1G22UD04kBlOL3cH5mWIJTluw
+T04/wDuPtMCaNTCdRd7/WuQ8H9A+wNWUS/S/nJ0GmdUkhGKtSx6E6DDQEkbSVnb
BfefoJycbe2Gk1c5twsE10z+iLfV6MG+rh6nL8txPxKagkono02gQBNqnPsM6idK
xFVRS+AykiUXpsKbnM2iIgT32cBfnU0+vISkJGLpefDcOW1ZTNiO8bgR7Z4Tz+L5
i35b+vI2h60a/t7XXekGayU7HZ2vCfYj2uyMxZOkyX9mqck8VY/Vv9k+0wGCzyEw
0GEk5YVK6idSPOpdjKRKPPHR98bgffSVeCC3NC7ozVivWoM0jNcfdOADta2ynjWh
KxvUsFeZylCdwfZQyPP7ATtvsJp+X2DuWqdFsZ28eUbdkgrTBeLeKm/rkrJbOPDT
MKLs+SqkhQqNpR3ah/VGwSg/Ykj5bx2XdzvHl1FNEixQ0d03xAPu5XN+oepD1G1y
RlpB6XYJMhZUgvv49o+LGhhmwOKGvCj23KAUtuYFZCekn/X6XoRWAOHW8JkXgZ4m
LPGj6fRoCAdHPcYDeWYXXUKi6+9eIueiBJyNnGMDBCYjKgDqrOM+IPx+oSkEz3Yi
sfemygZ/lI1V7RXkntb96txkDb2igyv7dPFll/SJvlnYkrwEpeB8OA0M52CsfXr0
pS6lIumF6aNTi/KV8+l/A5QG2ETnmdh69vHSKxg7BvSPYekAnONX0k8B88PjX3rm
uZkRtvHcf+iPtTBy3Ie0fnPxpzyZ5h73WUx0h1+yVBgG6uYBi+Mimj/yAiCJ8G3u
jbyhUDApnFNX2RJ4vDRi62UOFynmd2rj9StbVWQO/VX6HiALwd3Y4rZZz8KTtAi4
X9N1HvYeXkUdDBZhmjCgnt3MMKssrPEZReZmpFCPl5Dv5Er+qwbUD7wG+6uuoUtb
gnnnNlt/C3oZWJvNvmxI2KZ8BouFjbjsQn10BWvyFuKi1r+uq/JVFRxmHz6kx52j
+WlUFBOWDIEPvhCkpkPTCMhJwocMgi3OQebdUojlwwqHQvuoiW6ZqUOcT0E7E2KL
v14TaHpz3FIoUUmleatBlOpZfJzM9aW0R3rlIKjBO+Fe0vAThMUuYAW1PwOizT6T
XIJiReYSuKJruETFkfxlR5u5lo4mLRmfO+Rtgd58PNTYk6FrQLO7zYvVof+e7abN
pEobiqN6emlFB1Gc06YKFEbxVIilr+xxjiVddGN/gIs0phccGYwedkma8WkalrmM
nDf2MGNqrBxARZVc2+JRE6dU7Quf4JmWQblTPMByaWyPhdjXCOW/kncMlO3ufKcw
krWqFA9lkqgBR2sMHxa9wRCookPsEMeKHRcOI91iRHrKQbCUstWpd6WisCVUH0yR
8jy5Okeabn+89IwUFvF0E2dTxX3fxAlfBl7vY1yhr5IRxaW1Ill0/pb50aM49UtT
RslBFkz6CSSO0WcuibAN82aDZp7kWL7kow+14vEBBg6fPJYBEq7ieQsXFXmygtEE
KOzAerRTgtmiIWy/062jr+WWlcrbqdgJ7mqPBX5j5g1T5GTneGhvLmS9fWy8oIRm
JFq1aQZCIcM7dJwVw+BJlgtpLkz78/Gt9/ArmpfT9FDB9QA1/2uOixQJpDl/FRS1
Ya4PqYkzTRy2G+ZZ0pfrOc5l1su9Ru9yzD8RhqpuXuzDcLPhjel7Lu0YlyBVRs9L
iNr7IMiphGkL70PKmoBZ/iJmdwPaoZJqGCOJiV+rgd+WYfdqXc++BAx4jNEnpUdj
/5JLyLiakK3pHTD87w4PqkL0o24mCsVtV4uM/PTVciQFD1cFgBYdmUkfudxIyWvu
EOqoDst2zrYjyBou0sJAeoWPXry7BVkAqGfwGJB6y/vGdJe4clM3J3OFw0r8lGGX
qsPDz+Qy2xXZqN1qjJDiPsWaE5Be182pKosUQHqixwUVerc7F96qWUOI6mLYTqLE
QcPDtZvhlZN8+6Qw05PhoJdyBYelCDM21R/09UmAF4WMr80tKx/NYdJrZyaUNKs7
X9bejAU+EMtA0t4n/RySkZBQ3I5AnzmV2qrNS4f5ZNmNLlEhq6Hgz0NNHIxgZ8Bj
ybPUzqwnbU8LXFfdzGGmMJvkeKz5h3zFToKfN8MtaEJuqncFkmnoEgluguqt0sF+
2Csci1JA0MZphB2QIfsMiFclTWsnfuJSsEADx6zfqZa8LyFdS0zWgCNgPGBXA77W
HQ6H+oB+IQ1mCcb/gu5WeCewUJOX3oENRuIVjw99nPFn6E9KsFE2ILHb9A6+9aG8
svzZxFN9qqtnx2tGG8WTkHNuAdlkvqwj/JlXlCdI/dyVs35ZHH1yg6FLESVp5BCd
4SIG5bpoWiqO11bQBlmxE761osWRuSxk3mR8kFcU7iCCzBkDCgkq1Ectt9RPAzxH
Y48f1cTqhEwJIxzA3CRcql4uSR34UO8cH3ReMxCg0mcYhfcU26e/KL76F+KuK6zg
/1PuY1zIBAg5foPj6lS2n0xshdS2d257BUC/NmJhzB5WhFf9WiL9Hn8LoNqYv9X+
zWs8boj+LNzROUlDqXLEjJYi72VHjqvEnqPaDXj7Cj20n/sgPzDtGefnbB1gp7df
uXx8wK5nn2n21JfBkN/g8+0z/t/sZzEtyerxGvNy4CFbbOcL/gaI/QVbaDsIutir
O2ND9AW5z8KOAfQg7kknzI2eGceUrnHf80AS5XMBqU/ELH/KL6rRNUhsHx92HU45
MTbzSPy7Sq47Kt7vbfXGCixCA+US9lN2LnqOCeszjCKJkNX8NmHoxTo9kB3w01Si
x1xxHkCoxYjFLAPqYOzw1FWT3V4RpFFHh/l0S2faxGx7YM3g0PHrD5VIPKBJl/H2
doChUIDHKaXBHjCGOwC8Uu+8m1YwveKcDFnZQ+cd93+gvLosUKlls79GZfgP01Rj
bTBKhwjvr209HmbIDKHfxstLblMxVgH7U0+8JVP20KwSjxOrrbCI5oSBGmHJezme
4zm8pqWzE3y/6j+rTVXAt8w0JhEoA+T7Z3y9OCn/o91dczbdUMM78Bw4ZEbBKFKl
dihRDdWiPGBD3/lFdPl3PGqh+yiIPwbbRtUDdVljAfJJbCzkubu4qqTx75g+sEY0
gGkGaJNhhuFSzTyIyY/0RDkmEy5iDIk/12vCJjyYUdox7Ij3wzriJJT75Vr2YOP7
pvgvsckg6QHefikWT0bRqsoDf464OnWUERpWDc+bdsQDmZB1AwRQn1KwSpKtlm5Z
hpKz0AxbB55KvtQw/Cw1ujzB/FS8sZy0c84OQaf+owc+JeZidGCKqWZG47GFpDxM
ZUptOJ00exoatavjewUpIsanpu797XzQaaqiRVhaTXYe4wnN7vz9ejSEwcDK+0su
1eXSgegdrFx9H0W1eISdZ2PHhA6PhadOtUqAMbx55F3IWQKxt14rx/EOxaxEyxeN
e9PMt/cOMuIgLe7BDDvG86CSajy6TC0G4mdTP2x76HGOo7OL53pMF0TIyuJdvoUU
2Cp5lU15WuloMcwCobzFihFH31ovQ8PSa3UzYcxXv9bq8JM/7JOiDR/eNLWwpyGI
nI6bJYjh8sGXfY5irCaQR2c0xGBUWbvmoKc0ZB/yDo2Q7Broias+uezbs7oOac+X
zOfRNV3O58sFVKdiGrBK2BzvkBxsZd6UGOHQ8PefrQVXT4QcVhyqxQz3eKdL3B0z
mbLI0Eepc0NsuuU4RCwbR/lvKazw/rWCvmnq/fCbllZMuuxQhFVoHTFn1Px8CWBO
zristF2vI+Y5a+k5Sdjft1RLF80fihPZ7P2hWWgB+OeDTisPWg6qB5/ix21eOIGQ
b6WJz8HwfNtIBsC3JbruEiJ+ExtzmNPZx41LiZeeX3i5V+5W3Ac0tABtX5EIMTBm
i2c/uHEmsoDSEX5mwp0SW5E5zwCYssne0tv2+u8XmiNR+9tAF+8dudPtlnGEKL3K
35O/nVF2DC75JZFLwT11mnkCSTyZvqFRQDK3dnmtou4s/2Jf+yF5MQ+1HMwywHkN
wHv+fAmJjeuzx+N/22kSIdqT0pABPD1N58JUW1J+amSn5LANfeTKgEWGnIVX5DZw
`protect END_PROTECTED
