`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jHpU+yxiK0lTfTNzOunHd1yTSGuCoM77dRysXObgMkcZSe4xTF/7RYPNEISIySk/
JLOKYVi70EK6hkXhQO/ssQHbNr9gUVmCPgyzPxmeNQiNqtuzCSgNZiJuSo7fjaKJ
klU1k6sPqXENZgYeOpfeCp+Wj/HAfeDjpVvIb/FfPs0AhEnc+XeGxuiOsRRzKSQj
p8kNnxbiSR1APmT8ohbdvOAUJqNE89aaBGuTUYyO593BxgjJztzy8mTJzHVTv6WA
/XpTD7up1AxNqXLO3y/1DNWJvcAgC8IckJYf16NZ2/nAGdINcAdabwlo5p33MeoB
s7paZ64DI4QVx1+ceAs7W/cjkWI/WVu2dEwsVieBsqDV4MA1elkaOJz7k1e237CM
I98MAfGk6/Ob/efwW602DoKE/VBbbWY9+6Rc6hpB8jq76L9qqoIybwemENoflKZR
kRSOFV3g/FVHDKp4r3lanOz5b0iYv5uyMhQPDCyxF/xZAqvExB5on3op/69iNaOe
hKzqtNSsAF9kHyAhbXRpIGVu7ba2h83V3XjPNuUnI36f/f4p+0DlQYB42puBJuwE
6z7e8LC/D/vQrcFjrHXGYH9BVHR2UY+V1Sh6OvTTxSXoEcdVwQEkFgFP5u7mg26i
59WZms9pyo2zjLUhM9qp3KMfbgPu6iQ/ZL4+plBFUyOhYprLaqIkJi+GxnY/V10/
O0Fr1gcUSyeQWHr3HE6Yt4pOCyoZ6Nh8ogIEqcSkxQms2y2V/K4hrPu3Y8WUyc9H
yFlmtiX+i4NpeFAy5i3+huNdW4Npq0pNTs7zS3+8rNXvAsmdOeMv7UO6w/ahqwiL
gAYfPwvubGbawb70kHPojHpMkDS8p55LFNW8yQCvzfIMj8Z0VJnW5z3tlKx3WqvF
xTPC/GbO4SMmnfTKccskw5gTdpkEFBqubPRiKUHxec6yKlxMgSkPLAu+wu8ykHJz
/8UhefAkZ/87jp5479jg1TlpVYI4+r0ksvHG41dDdF0kpLGvbN9gVaO/osSCxfS9
nd9GiL/iYEayua55stRyIdQVr+0x51qWsYqiNQN0T0CumkmRmQFnsonpAAmVpJbn
7dc4j8mhDMkxWnM/b+WrjMIL1cEKe3bEb+rHSBCB4mT6Q7C85iCpGGCN1jhk9DkA
mSFEEeKz5EyCWaWgr8POn6aGwdUN0gaYBpDrxc7IRI1FSFFSNn+Uouj5DrXns4YQ
uzn7rbAnFLkSs/WaTBLYiHNdRzRPU0LgUug7oQsU4i6H4ZSRJhH4SIx2JgEkN6un
A+V3oyIz7g4K69LHLKbLo+mTkfysBcsdZiK5a6Ht8Aq+utBQkFS8BZdA9BtysgJH
Hy+6VD3Pi1YH6iS3yDnps0Lxde11nau78mP1+BMx9jxcc5y7MRFpQtegWXSsvuuL
MjpmsBbK6GxJpQX6aMeny6nATToiiMva9ZcESziacq8h1Pc+sDAOmFByQv70D3cD
TM8qAp8Yf6qjrRyc0xvvu49SdZudreLuewg7+UU8Z53NmGjD9I6REO6piy2UB/Fs
iRN0FfXvUyUuHpggJVYEh9tnnYzO+qRvUem3vJb3Y0V43L3mOzlxMjuXPeODWUKS
scEsvdcFhySUGgg1MbTedCeuoY2Q7k1Fbn/jUsNf4jWNjHSGneI5MvlMKm7q/MAX
OkYB1bLXQGbQbQyrzMKxfIoD/gwm+yQUzy4GjdcrXdJYDTTMsKDuYbheVkp8qBhV
GCbWojRvHehyot7y3gF8/dzyOG3SSRKlkuMLiCsYdtM1d+fWg4U6WYTU73+XYeuW
OykNtE7dbdOdKKdWaLt8Af1JOke6mlVEf6C7DJvtJlFUqy22L+edKJ1PJH2on99B
p+PWudPHBoYh6kgqjhUoS0Mqitsci6UrGtU/JKA19lhisMa2Quk5F8kcNihpDaTL
t7hQ8ToXAi+wXTeblrdXBy6wKaNLo866B6JwaU4c3H89RbhYDWP0538prXKlTIK8
00BFgihKV8mP9/dAJvcvvDV3npEum550oEzMLor9ZK8KpQc8tWv8vkinZZas2cC9
rviiy9U5z+rz6Z+qalNXFlX9d68nAW7eVwvNjwQ49VuK1VdkQOji0UiX1ymiR9c3
dedGtOoqtVjzy1EQMNiFrohmiaxB37e9gFtMzinGXoPlE2W25pEAB1V6uFTZJDOj
WJQ1zKihIxHSjr0qL8ZGiglCRfOyWeKB7HpOHaASZ45dpKqQciL0HhaC0ZK6StoB
B2fTmkHekVXnnQgkMSJMMf2rQ84Q/+2bGsODT9K8vS+RTV3Wq5oa2ixKh/ZIQjO4
lZDzpAOpn40058FADNCqcr9BdRIYMyBvBj1JnRPLHoSn93FY2fyzNl1LC1ciRJRD
bCY4+TXveoo27PUr41yslYU90S6xRFu/p0psanSwMSW4/tOpmgPdxcQYElopb2fR
VvZFxI8S6uN3rC2gyHwfXC04MyniVUJk7NEp48qeQnTBRFvaDjnLVkE0ZJKp4DnG
V/ADOWyokNxnmY/iJbF8669okfu/yOXz9Y05d0Tw5+UvHr3S/u2C1sl+u3Q0J3Bm
PTCyTr3/SQkAoxTxT8UAi7/DkQiNPWyVJwtqsWzvCxoq574yd+V5PN3h2FKMvjRn
oz0E1nRLkksRQQWPSFwIl7ksSZ/gb4WimpJoYEQmNz/8B2sRG4IVWButNE1yVPet
/2cJlc0xfdV1jSasy/NdTwuXemz168UxWnpDbBqkLaHFittmduT6nVKQvsUd9ja2
OoVEsxziY1o0cn/Vqt3aqDUPsD0Km9QrEULqCGWAEZthoW+3hV6egSyulXcXPX7c
9oZhdqLqNRm+sGzmwrc1LAsxZTn9uOqK6v0fo4XrYcF/hV7EteiAH/Dput6oEoy6
ze51COeOLyznQQrj/Hhazm1xhV8kwM2EggsIGCEpv5Um5s4Mo/shvrOYy4GhY6dz
YABYOLSf88cKCUNdP9RAhMLllp3lJZjd6wwwdx2xBKAwhE/Jbr5qjMje9ptdP51K
XSYlV5EjJmql+NwycrKOThZJVW+trhvvH/zDtgXmjz1crZtcPTMjtutoa2A3zReB
KVRQBVboE8KF/LGORcGf30n5ujKgHYYPPST8iWOeGYrR8lqry1r+/3QP0/eU+qeI
oE022mQ4ksyWm52qX37UMm8sSM8GzVWH8N71fp/PhFVL0gEkejLqoXeuhNAkt2q9
0hCvPCdk8WgKzTM+K7k4QipeFmNeXZ6h3MXaRp9Ym0UoyfhjIuogxY6KeFvWzYAW
dAwADKB6VVDbHTZlYg9WcQKqUglWEedXEORphH9rQzswHjZC9YXL5AZidWpS8WtB
FJRtrYVsA2niPTXokIvJKn4e5g21GhuPSHDqpF28BIewGNB+amGYvpikUigAC/He
a5yS0C5qokgXpURccsRgyP7BYUGD+ePUrHMjrj0/WXbrE5dWhfmrTc3CRKBFidnL
oeigN/vI/zO8m1TZ8GKeewMP6fysopdQ85BZq0D5AxEJesOdVEbw7EsT/PI1E+2Q
VVG0WqK6bKMaAdTQTT6nvS2tjBINXqdLWEft6otSlg6H1sdPs7s5CV9i4VfcTdGq
Mj55moWK4cdSVZcw7e5zeN99t8s+JyDRSEByEOpuT/Pm9FZA0aapo69g+h4pPvDY
MzaxukRRkLKQMcyc30H6Camm/HRwQ85uXcRAo8Gp2LGQn2/+hW8eZgD/yrH1zX7C
SU3X9UZkWK9vu+TUv2GJ/hs/WRJjQEDATfa3u+CYzsCK5HB2d0R2xRZfle/xUjM0
q2ZCNwJ4N3RQkpLXKXJuOWz9rBEiQvSIcOS7HhkKahPwfPSpeXgH3j1v2i3h06sg
YO9EBlyO9XGP751jqKowgo6+87c6klJMp964qeViKxcGQ7HqCXcw63Mh69MY/gc9
Kn4dfIjwV6EXe1lx0hTlYqUmV34vJbpCedJj34xAaB+6jfEFizT1ch5PXn7CSRSN
JPy0g8v+/b0838Ecw9y9g1sfkQzx7TDEGbGewBzul4hoLJ+6bZWrNsZBO30bx88h
hMWiqiOT32d++x6NVncRPO6DQsmNYOit7Gq4VuyW+SymdW+rNIFafhpUOo0wmZcB
hhzWDZbhqbT75YWLTBgpdsnhqzREFjnZvgWcopyCt6+TKoNXcuDNILLsHXWprlw9
BprCuPJvDGxo3h5LTm6qPvhLldu8YGsL2RZJ0m7cTta3q74yAo+G/k1oluLw9Z4k
vmjO7G5JUwto1QE5ndW56xJErWLnjM+Oj/5ibfO+5H+F5kk7ha2zTD192k52OUyR
CswltCl9394cn4YXhanDIJcmMuRUQTMqt6Cpaw+s8zajckqEOhamk0CP1q3kUVQd
u4dMIo0jJXTnDqSgniwmI4QHfZTBxj0dIsRur2qkdjp1qeUFnlJLos4E9uw4igiP
pRuQrs6EPmtGQA2JA+IkQn3AqoIWEzoKfTjfEiiK28DqkcQrV/t9lGsMHRmeMPlc
twQCTkXZm4kirrZ92CcxqtC1t02S06Uw/LAo2TjBNZHHb5EgC+AFBmV23EB++oDp
1T2fmHx6+4dznYvJYOlp0aGTcXUpuPORpT1Mq4UhHG2VlErTtF+2BTwlkDqlwpiu
2nkkWjvtZ/kbWaI0m5keVz4oOBPrkrHTWO9Scdbxc39I2v9vMa/N8hTzeZT5W3fS
bn/iBMTBCtuIOpMvFdtvJPqkpCOUKiEA8DfMxLleEV+nyiICDuFlIwV4pO2CSQfw
UuneNnQTPjRlZ45Q6TTvBvCE4x5WHY3utXP1zZRw10nfRejCNMXnCpKAfIYFjJUK
FixgwOhCcw2F6+3XaGtn4ccV8Payp30cUdPboYUD1trp+Z4B3HZ3Bn34I45RcSsF
Nvb9ccslPvbH8xtTa9ulMVQmFNlQ6Y97yvDnEp0nPMqZoCmEND4Ry+ujMZajTxA1
QcYCdDRSklyRKa8Ot4Jn932rcfJpSJvcZJyoTT9gLFIDdF3P8LyN+G2aLSJm/w7O
CVB97Jlu3uRMF2ILnjdQgnZ9gSaTS6Fp9ANnhRwxX4rOm/ybOpQauinYKilngYwV
DWF8zmw4cJ8zPA+iSytjPIP3EBe69PXNxdRTF3yEgPRlGFYdQdV1m9yOz6vq5U5K
WFJ++x0z0rE86VNw5xi+hm8yuvqG+zrRoGNNNqnMlXLqCffUTyatLZjfix38PH0H
yt817B0sRenBRl1n3q95/oRgxTAs5JKsW5y7WPi0VwQGWdXVESEJXwPFqwP7q7Ss
MqHcFWHJU40+ivGtiJhxa7ESxieYG+f0zAexhU3X5PS1M8xcizqBwzeJ3foTO7W9
YTcc8AdEWMoongWTlEwGqQSKwWFei8D9Af8sOpvqmMKcbBIH+lGrnIQHh94gKP3H
nr0Z7LwedYowCy1kUoi70rnpgJuYUBnFkLr3RlQfF96sDv8lCzl8P75xPiEgghMh
lM9WQaJZqgTtucGET4EIgiGRyiwLIOInU8r1ODE5s0GbWdSt/OLh419w2+Hreh02
FUPev7tecyBO/qwYDQsKycbhFwmfTBCOMJxLpKsnmnh7gKHTbaIXwACcipjBi8me
EQQAH4l5y4k3V2HEexbJgZRDz7oNU7sUCawG3RqQzSaylQISM8GntkFWkEq6/Bg4
8Dpu/ZNqfhm3xhoI1MQshs9KHGLJb373Vfid9WdZT7D/VjbU4iMKEAnuoiTem855
KCUvKPEHkhH+999GDLhMGep57zKzuIpDKT0fGwxxNu5W5PVzhZk0SFD0RbAR/FFf
adHcaVNiVHCla1Y1QGTn1hJhhUWy0uCqhBwqxEzg4ORNTF5FUGu4yNqEIRB+rfce
cMoYN8illWNoeYejwHbj6NQVVIBwaOkvaJezPS+TTaVonUtIPvIgAMdxp7PhX5H/
oQfQq0xW94sMRie1L5x9hfn3nzjz/AS27yVrRq1vDQiweExkLJApqy/tRE9W4l7/
FXIkKPwv0A2yNTN+vdLwJhq7iwK5VOc+D4SFiAoH8gTZ6fM5FQfgLLtTueadYhPA
`protect END_PROTECTED
