`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bzuSQQsRCFJv7DZ9wPg5OKUDyVrwXe9NfBuUBGzmHIFDBLKkai6KE4tj8zOJCT2J
+klfRjdq1mG1bN3YkHKXXZ48i0aAgDBDKk/TAotze6LGNwjoF6PtXBMtyBJkSXxp
jTFFIM3JNSNRcNryX9/0CB3BE2fSkERLCqRWhTtmMuHbpNZD2MXorSJQHPlbKp0+
LRrqqYGB7w4NulbvJuj+9y9vzn0+quwxZ3cgYBC/KuxXcPq3wNC8LOkCEmKOE0Ln
Pb4BTgwOf5QYV4WWJ8C6dk852IbyK5AbZ6dzTR4Ol+js3KFvRyaVl8IRfpPLHxpi
DrzMcbRBu0LZ+dj2scn7qDLfCdGyX0276GPtEWqUcpb9UMip2UgCtNubevrkxE3G
2LqnutRrPVCuNF8Lz2MbqPgbrHrMKYZz3/7P2wPqRE0+NGK9o/w7yB5AnJPa+STj
EvyyQEWKo2uf9slabTObZEGCuPXbH+FiTJ+CrnzZiFeZhidHTr4YUhJiSc7iYmJ+
oRsN48nJIWKgzkU46a55pM+KIgLCWb87LvqGfIve7Es8Dh5G6BWfH+frAzmjpQn7
29IEebc5HjbfnX1fuyNNxF4rrCVcQt8lTRL7VBhJX/5Y4jGGcGFqvXYWsC0WSrxd
A32+y6XKRiRVa4DyvywkVe8h9j21JkjxIwCc1QMvAHB+Huy/yKsKKS/xB0OOjvdy
vrQi2nxp/X4X7AOmlAiyfmGgaXaA3fWFiPRYN8mLN1z7I6/aoeip67WMhoNKnp/f
djiE+wPfwKuby5QqiPx6fbDHr5nTbEuTHAiHqJxAANeCW/SGRFVcshBKsCz63Tc2
WKtWxwFLBg67AC7v+R8kSjmINCLb+/PETT3Prw5CJVFcY0AoaDAE1AytmweclCk1
Bl2bCS0QTydG1JJ/GAjJQhsEXsaHLAc7RRJCz4HH7rA8SiWv4gbaYllT4k7fmVnF
mhcI7Rwu8Zmjg4/f5ecXH00Apm7rWGbexq8SuKwo3jEM1LshPeDDfI+wKs7g7T1L
v2aE8qGBSwPoQQwgREwU4fGTkmGSJsbLPLiQYmH+y71xXrxYYkZzF4wzNf8W2Csk
6korDrCzy760PhaSo+8dNJdjzxXrDgVp51g+bpTviuD2k61+scsnnJdrjwSd6p6E
I6ZaJUK4PpCBr1fn0Q/p/jVGLGT9s+Jb/x1F94tOX7IBL9lu8HqfmluvEyAUQ6iA
P2CZlpdK8UyR4JX4RJ+fknDghkeAEZN/Vf8nvTr5V00=
`protect END_PROTECTED
