`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WNAK2CvYQ1VlpdWebqOmXmz8CpEPK1QQnvKKlzvYrfhOG0S96zXu5Iv9WYBwkq7h
JMtzmO1/661vziYuw9+X8sbN/bHUbGCn9hhL/gk6sZ7d104EVnS4+v85uyAkJ8QC
PUZ6BX+bvF0RErziXTWrT/5ndgSuYkL4ruQE/Cu4u7KgOhuvBKkoDIGrHDSNpfi/
tKPoXcG2rCQcCq/4MILlY/kZSxc+aVihPoXyZmStqtIPr7l8eIRmizVpGokDGiEW
zyd6hx18/cI3llr7W4f4ByQXyyASkSlbm16E4EEb+gnc+/MYWgzzSAGX1U2JBwA0
2I+ChFor3eSfriwcO0nSw4YFRakA5OM5N8bo1bcwErHIKQwazACtGGbbnlHeYLCP
sMlUZzZo8/YiQpLbrY11Pv1FjsyZj2i3PPQY6j3Dd1zclt87jJVYYak5tJW5UmWr
Ky1xDGlhsAKhglDei4hSaMrtUUutqteG3TNuOxB9DMOzf2VLwNKuxH5zoxPAfGUe
ay68SLdfcww4HIFwlm/qxurB+NE0fDgJnG/L6dQwBLrdZmJxEzGgDBnSmjohjS2O
kYf2UIfn/ec3oDaYo5E8R2ZOqq6XjxGbyWzlRJudHSMF/lGSCLO2w6J+liCaZW71
1oX8QSYf5UF8dA12tgzV1dVe2QjUaec89hfEk84Pn3Aj9qJ6pYEQotSU1kyPKa5z
2L0IiA3ufIdcaVzZ0Rtu47Yg2/msL5VCtbZfnkBqymTbo+77NXTzxb5L5ryJPIne
2Z2fbsTtVzDH1ZYGFrb0Ofg3VvE+9oPIXGZdE1B0WlesAbw5AZxSieb05Ots17zI
qlTA+3BaMd7AmJtyCDygLkJIr9wjStTRxg+lbN3arQtDFH3j6eXhfkxf03MgucJt
xc1J3qMqJzKuYu/VCxSU+ID1f1FplrL/EWLqGm05MDZ5yL8X6DAe799nQk3jc3b3
kPPHWUoiFzthQ7CHc34JsTtuv2NFVw2YlVaqeIYiEpOrz5NaJ7zKG/rahxbIvF5O
F4Y9PrZqj1gydY7Tb1vARzZmDeNqNK02FvtMCup6vnzC9eBQTFBo8m+FTizQ3Cci
j19lRKSknTHD4a9QR0tnGcf0tidSsHoDqiEydBjOkQAe3lODphFp1WJtL3cdgjfy
jLZ7uiKAXz5/V99i7aPtNOrgmhpjAeSEHJznYlazuspOdsI9u9og99tBH2cgpe+a
TC9UcujLe9FaiveKSGGbXmfNVgfUqSGLWiAtxP+4aVi2ppUk6Z18/4v6zQMjDR0j
E0BRZbTQE9jsTDWLn9J5E1pX4IonhnmJm7KB526OwqcHPouZXYUCuJHM5kdIM3zw
1HLsxSsHlKWUm2d/8qZhedOYxdN5wLDU6bs30sFHt8WFCHkgEIWa/8+os4NrLSRr
cdTVevm+Sypyp+i1DKJIg505l7N2cTLow2+aM3xJo/cT6qZ05d6fUvajE8Yc+p0w
jwk+RuxAIoY5bpZFzLcRwpPJ1yb6ZEmxse9Rt5MuSaRbi4kmm0f6W1K4qdfmBd6K
JXJcAcPLrUCOCL3WY+OrMoul7bmGRymvM0oILTWI/OGo9Ck+VuTLeVFYj0mSuoIn
0IS1qa4Tri7ndB4YnRtKfSYdL2ISnZnFz3PJy9bT0V0MCcq2OqSZOVJb94mlj5lg
IOrwsawzcWSVl+FqWH8BlaAMLcynQtU+isB1y3gxx/9nSW6iFWWMygV4MAj09wNv
OeDSdDllWVuUnVpT08avQkSgwA0pLtIGDsIC9E7jlgHAKPTxlMjTOJceI1Ns0Hnf
Cr4o2N/ZU6pVymKdw1GjaQ8CO2U7RoA8LBDOgsdWtQJiBJBkkxpzNZzM5jKRtRPG
xOzCLiWFmBsaICQMktgleMr+yqV3bbAoXvjchAes+xlkPlWGVK9YhzcLSNiM+MLa
fWzcrRQdlksfA2+cKB7yYt6QiNNi8XWJINfmM3TsjvExGmfGUMARQHYF7Lhry2Ag
/D7/w0t1SFDLBuIt2GcPgHe7xz5N4b+VHsPB157f+yHpZ0WUmIIlNcw1YowJRr2v
PWravStQueJap3B3c1hA1NO+dnv5Z6+DVhXmk2yJVdiInjkZXi3o0J2trK+97+WM
gvpwT2cNGoVfFdZO6YZXT82JtlrjqSNcdLL0sA1bAkQvxI10yjBDqy6V/f6rD1Ch
thkEmp5Re829FyGADribBTP+IzvF+0PyZyAVrAbLbvmRSQKBJKptEBvQwhhG2o86
kov3nJHJHsEtKkbVNDfJ5KImOruQVgg+ZcUpqAQ9Tc2c0ay4U03KgLy/KwRXnsGm
ZD5mQSuplcIQ2L1WItTRzcl5IXHBHW/kzfROqS3XOPTxNDkJQNETalFr4tuAusCo
9JkBCgViGK+QFCexE00BG319gp78tcvmvHBUpPVCdNkC64KySSVl4+WlbphSznsk
ymLEzugIwbuxQJKBV96Ka1Y25Nw/a5+jN+24MXlpewv7j/I/yEA3Og/m8nWrb/7m
LWAQGNCNWVW06QbszezDG0mK68EvrnAie5+MPiKhp5Pr9wOuKB5PPIvNNbrfefZG
/Xx5eMbQdzPkHcfca8hmmgwLdV98/DTQPT76Qul1w7RH0DYYQ1YVy58uwsKI6Zwa
yoBS4kHjZAaJK8xPsAAFJYvLujJzOOzzveJwzZZ5maO6LQsuZyLFXNMFh2mn1gKJ
lsThdlIpErwV7MeckksZGziMja1bMl4jz6J+WwzRgZunMGcS/FQ2LgIB3v7paNPK
Hzb0+Ax8SbqsmE/eIs36WpCEjFrxVY7LDEJQ9TBAf0k6bWAhrc2LUH37fIDzTcAS
Ree/5RTLuD/2QNvrnrHYxGbe391UPGC+5RiGydhNi2BNzW8zotKBcs84lUtm7aZz
QE/XRDPMS9vPgW/HP4kthoU90znmMcdcKI7Xjv4fGoK8NDPPhbvHL2OptudUCWLX
itwX0205BC0l1IMns1z7w9xFHjIKKt7eyYkmRORtib6K4lP9pu+FpXRyiIA3NxFr
8ofLCCSTJyUmT9MSOyRYKSR9L0RApLPhVu494YP1CiNsZ8cD87Ay/vq898v+I1JD
xuiJLfDQ97SVGSCPkA2vnLaBTEC3F8VDb0ix9aJVLp6b5m4cooTtXiOWkyPvusct
PtTdhfulmO8mrGbpXqHMgF+8G0wlq+ZqPHLLd3wAYt8f3tNYFKIcAGSCBtOt4WgU
JahHzlKMZ7jbmhE7FrLwqnBc8/3HSrrd0QwHyBfjKPNe0Sm5OhcaPr0NytNBZwVw
6s8kAzA08OPnDgI8ed6WFAaaU+7fGNWSfbjJDGrQ6GLnRUebzaKTj0QRZhgpMCTP
oKowF9R0tQMosWs1fPLhqy51HUGNU/YkTuEDDByVALWjwm78lAgRfLqn9n4HbDd1
lo8gDcnD9QcYAUkkZFS8ExuBOt4ByEb1qi1d1KX1ZAGBOVomX0jZSkdGLp+ah/XY
RFJKoc3GS28cRuZ8IzWtADssxAXr0U5sO3xljEcIMO9UBHajx95sYp0CoXMpSO+e
hLzXw3zu7gdjYVQhxFt7Ce9gHD1C5QonhkDNBiQTuZXCryHt93YXj30it5ahELgL
HkhlUXGyESkV92t4UrP9gIfHHrlr5/9A2yBm1ywwRwUzRSBv7Iscj+Z09DXdX5Ew
Ej3/sPuUJHsHYR5CfqT+X8lPDigLrLvrk+H2HtVx1TJq+o3jx6wRtP5zlF6/yw7F
YBUlF2KfPrYH40QLT8STOm3Ff6UWVNdRdxBDFCjtEOISlkV0ICCpdQY1tvSSvroV
Wp8TRzQFxAP2BhL8nty6pGQS5WasDWX9EgYawzeDfyLaHceCPDV2MVPr2Nu6fi5+
+gCaReCaJc4I313pjhj87BkzrB6IN9sTX6SI8PmYzy3wKNWjtqdPLgrzAJ1HYY7m
rSSgG2DbHreA/TdFD/AIPtHgN1QMjVFg9rBq9ZC583kWZ7ANzgMILVElLbOq5jeK
XYcazz1mLczS1fpfxgnT52rDfDtj7NHfb7ghntkRLz8wy0EdCwXD9XMaSMxVXiwD
TSrYnZ/LIv77LffrPVLbeqzWXzTrsCYD0qCMtA6dmQgDUcEGCbT7wQe7QP1x8plg
Jh1OC44AC+SYZvjLnkWc8HPb2ol4Bukb3t+LBldZKjvivxzAxpJvsKVi6FJzV4H+
2L01EnG3JhV8w4gFqjRpwWY9PjDuU56Q4rgjAFtop+DmVsjVeBD5xRHUVBYOu2P7
5eqhgl7Iq3TT6+MpI/82WBioGITCwF3hbfYDx3KzGuLEq5SuTXPpEqq7ly17eufe
rn+VL+QL6ZRLFM72sRNg8i/PtZlwjNUkAPv52lIcFKQUHTKlXnB1w8aAWgGW5XH7
ZWhGCkuzeAbdJCHRc66EP38V5xQlH3q/+MtXT6CSxkw7j4Mu36oh2/03CkRMlSO9
UX7+LsxOqbHkgfxEoU3lVHKIOX7fm6C1M3JQ/u9PFtafCnjNgEMKNO1qhDj0rLPs
tHCMOemkfen03Drnx6PIzMZHFAgJ+24cbx9XHrYK/J3Lj+VBiaqB2+sLweWns5sa
GngXYIgaGaQpgFXRwkPWWccCFk1z3evelYxIA6rFQGWbyjSITQvsn603G3iVJcMd
KtHD56yYSPIutpKt0forcMOAdD2J9mFM5NaWL8YzjgHaaJMkTgGoPDj48LZBFQ6c
xd+MdxgosdOyEmHYqtdGvOmkEmn0IRziu9G0DYJ0cWaQUHCpmBh+93wRB39QHWfF
J8416mQbrK231QSesjidneqaOesYUkBb54t1p1BVDrjWEVB6mkEbRsHYx9GIot5+
hzERcfB4yVyi5uyKKI3ZxFe5vjw8urB1YFbgzJ6dd5Ed8VucX1+340GlCp9HWOnD
a7rCdvX4MhMxtRacdeErcRgOhmKCqM9Ke8fXKkSNusyfPDWOmhFv7OPrgD5v5nyd
JNHpeN0gOygIzUtMcnKp715mzjCR7nuLMSw11upSDM1Sui/YAEVmVSqI6opidRoE
4uHlO7ouQ0bZuBRDgMoY/CqbU2S+bgk+mwbag36GdW0c7/eicZmk0wdezTA2F4vI
mVGqCN1s55R8Vqmm4aybtz+6VXG02Ciy2f3TlN4zii5ZWTG91pG/tlxnMXCpL4mr
Mc1a9HfXUBfHn+y6OUM3qU8wer9b1irUh/uY1bDwE8H/FuZepkzRn97NPQUrspqx
9J8BzpMVkeTTNwTL3YYIkKZyjV4/xyA//DehldvoKxmlysYHDvTQvu67a6gFDNkJ
8LCjh7qYslguPH/Rv0bTiZqqoAteHS/3gTw74QDYPhHIU8n5nrTtkB+wJeWh0hh/
lmhkpVQMaX7yBiWve400ITgR2Gn0V5ZsQvqZDkykFXccIZV5eZ6pP02uXywctYuW
luLgQasPjMyPqyBZkEkdj3UUTb3BfLMAJnYT+g+mFLLMQfNHW10EMUtQL5YDS7NA
RPS/JGe5pitRh7sjSUYe9PGrzVhonRrxEpANhfN8dQm3HR96BURKk1acc6lVzh81
wksM6cavC1w0RvH42344dCp1M28WEOrZ9chJDVgdTINSykT+5Axpa4Tk+nLPwqrc
uBEPf18+52X7j3xBjNEXL1c0JlW1zskLIWtKO7g+7smu3KW3lpJe9BfeoU2T/0jV
drehnyHtm9NlfUaNipLTmPAoGBO5dhSo0QXSN1+dMqxuJa1yJqip4tUWii23o6pj
qhhLlBM8KHcpGQiJiIWTIXw6MAWg0yRFMUsu2qy0OajMjOAg0yblA8Uvx5NhIxa8
ouNtbrc5rfNTenDiYOz1HreMxaC8hQA4u25H9ve7ng1jbV1ntoZCNUTpqDhlZyXR
nccQPNSDbibwZedEif6VR82IBZLy5fgMDYSc+JamcqwCn7/OuIJguNLlWeNK3fti
TV1ar/No2SQ/Z6ASVdZv/KyB1fxHwrnG+4sxhVjcAuiTIPGLjTutmzVgbNptyZ+C
3OaRRTXJAlHloUIEiXdkjqB1GJQJlj1Rq8PCmpt5mK6BbZ/EaMtdvn2w1a7VyUz9
dE5Hmf2iO6R8rwznC9as6f37EyK9HIMHSWeV5074/108UYCo0/Ubif3CbkGgFVig
synM2KoMBNNvigYZeBsIZcKB84t1yvDFl/YHdD+kWwH9oziMwNW6j+8K/LZNmX/c
39L/hPIjY+BSd/8xMCl7ExUa/UUPxCtd+kptbSlYHOORGdnONTdrFnuC6spctQi/
ivPX3oDzPcweIyxd5DCk60L/Td66u4fKKFWD8yTOuj3puXoElZeL/Vbzvt/PQpil
s38PiiTLHo0ynxHrJLHOmoEL4kSCSb1D0S6ofqTnp4VP9PllrL3Bb0jiCduDtVs5
lCnC7yLafWVwZBwhn7L1lvkLHyc1Lv0X3vPbwV1qVM7UlfWXCU3CqLRtNzji7qg0
s4cO3GvlkxFC9uPiznAQP+nMsjqFGsL7WgXW8X7QjjxBcOTa5hSWO3jePhelUBPi
rPKNg9pgW/a/bYpKw2ePeJz25XRQ4bDAEwK/dVbKiZV4/1aquxUGaSxFafFaWbY5
bPz1Cym7OtWQ29ieW8Jdu4eEBhlw+/W8PYHIJTVsdDKKLZjlcBJvHf4LyOEESOGb
4nAMCKW2N5qoF/QZULsQP1EDq5HkyWq8s5n4+PDW+XcIaITGFMcVvfN5zzQBR3wA
hOm1ahM2/BKeHI1WsieLIRY+XSY/+wj4DzNDDxcNAs0eQic1UxCt8/V9euNCt6Vc
scASGWV5HR62n19gs+YrUhdPTfl1JnhdynGYTvuofPlC/bx4u/eVUnnhFSVNlviZ
OWjZOog+IfyeKL/QMgDgZp+F8LBA68UqFSJ6OBWQQL6PDPtG6lWpLhbWei+KCEDW
p9kf1yiHl1N06xO7Be+mANhJgvbAK7KUskbwftQt/rvaaA/Kmti8UL+2mYTM6KEX
00aee80Eh1gJ4ClgUESEA2z0tZggVhM+SoCG3eeTyvPfFVyUwZGmO4kSNJNEmN7Y
KsIOVZWE0EJ9BJRO0WBBheeZCuL3KoAb3lPkAxNZ7OC7qBpywT0kEqJHKwUnyy8H
lkykasgMlwGmiLzJndI1Cis5g9vpoffnI65LGPpo/4tVkPlVSV37Dt6Maz8V1H7k
grGvRGhFKFK4INAQRPJNCh/tJzeUcwO8v18irBpBVVRcFivC370KsQ6z5WNqTcYT
7LUGIYsAqjHiG8b2DbWbyOVVvqm0esckvLDChZ1I2ANXnTYNu9hy0e4Nye2/HNmN
qSNsjYjweXTP7lNrTDBIC4X6maS46JNn2KrxkxDJazh27QNJsf5/5Gfm6xqfi10s
+SFF95Fjfb79oudTD+h3VKW7A1I8fMuYAgnf7/2Dka0OCXncSIw3Apk8a9urwpUt
seewm0So92VXuiMZaLrL/vhw3fPbP3Bhg7P1znEySeLt7VjRf0aY5Wq80auM/f1N
nojEJTTkwwOWj+Xd8wOkUSsjheXq89gR2wt0B6b4jhYKNpV2tEWLrkmHp1K5qmGa
JHiABWIU0rP7mnJ+k7wejfSYxgU96HDAJg3/6Zm4/voDEP/1k2ucoCiB36obBUJJ
TScHimgYkiv25G9/28MlWBazSGPaz4ItLGKtBCF9Le9QgASR9RP3cl8vKJ229YzA
blf5Q/mBx5EaOUhmTHRWrry+YD/awM2G21toG90M162eC+K4kBQxijGEEx/8bWu7
VLgnf2ewEQEefisrVLSvSBENrhe8N/v73+psHiKXVVaWfcC2cMd9/EfK/ZtZH0Us
JEoSuJniIx+6xqR6AqEeskxausvQh9auM7ZOPMwqQsuN/wje8S4MXD23MfxGfkC+
EaDts6uFcfaBspC15bSRREPUWaFYoZyPVUIo1lw32RUmgKi4uyGGgq33l/mPm8mW
OAtQTaZQomfJDXH2fAgtKWmOgmVrFvAzua2P2/iNsPUV4q8n4cTUiXHXYCzn05GB
U7Aid652flc5wkWo+jt5qmB/j8HFlHugcALAnpFy/IH1ZJ6sv7CsKQy3yZaP+hWx
jeoP3pSBUa7Oz3XdMGriKq55/naqx1zVIjGKIowwgP8/3lqJabSu+SA8ymbKZbfF
1YQkRgmYhKng1lHleeB/0l0Dzsv2Rx04AQDe03LGjUgZo/HLCasYV1N2Aqgbs+qI
1Inu5JEc93uNR2qzTaEDY0L295pV7SlM5+JM/8V97QJkACyty6JHrWQ16dM/HExW
w18nRfQvCe3Y17t+fNexOyEpacXdoJRtHZcE0mAPij4gCKqFD91i1v31fD4oeJUg
V02O8IPfYsasMuwG1fsAAP1Y7fuiiGvkSnA0xyb/D3iAz9/LY8i/TqdS8hYZkNxt
yTvJ6LnFX8/B5DYGjhC+enOpBs9wzdhf151H1cP8haOSQqCeNxVizYMsHHfGsaxS
aO4VQc8qcZD7MfN6V+Z8AYwYy7sd+752mFRANKV2BPVwTxSWSwa1Cvn8qOPtMgt5
L6wzJ7d+YDoXK2MQSB5oAS7C0mVFqYudlNd2nWteWF6L/cJdNIwNFIaLAU25A7nU
sdG408MgeVNEHKCLeXM+z0qjlLTbRmwowMQvCiD6ht27X6FTigiKQEqZNLDHKsNT
vbsmXL7voXp4rJv6ofq2X86R3Q3xath1kdMw+cLPLiduFkB72Z7Dl3lWqL/x0+Ac
6LD0Itn6YBrClnxuxLB4PVGt72LmgKjlJNmUZkIB/CoMB5UiSrCfDkrwvah3Ov5B
AY3qK0kvkXUhjcov1bTsh/C5qvBXWO40cJEkm3uYcxPVhPB6//oBJ8kCs0tBELZf
trcQoieIyKIH1y4Iv9NTBgKvTiFKVthVrGhxCydLG/M+wHvapQOfSUaUtyDAQysi
z3IW/E2qWPaB7NSMpAtLpQ+cR0nP10DoVA2Zr6/qt3su2yzxhEuu0qecJOkVP6gS
SZiqXt4JWdhTXrZtrfW3pf+LFfNq0c+gzsVrj1lfqW4E4c9BsJsrZt3vEHM0g0XM
BrY6gazsyH8qPJhUseSUb2LxacjD+UQaIDOxzo3jJGlZ3xCKpUB5Y/xiGolScAzm
SKlzthBxIBEginDFNc1gIEorvcFkXZO1f27UR6t7AbXIkmgTFO/jffXZy16wLYNC
wNo5YNnazZ8yK71laCmsuqEZPGsUPI/6sMlkjt+jJR/QtRExJue7gddYzaZ0NeOt
nSlLjTdFrL6PskqfHjcPB6teuhWwHiclZCxD8kjGlX1Rg/zwuenUFacYUtl8v/Rx
CB/dDms71BxMZ8e3A49I0NimSoPKMXxchRc7lvC2R+3QVTnNl/7gQYkVDcER3Egq
8maieOTcPqD9Xu82iVX+d6fUDyn0/Wr82W7S+2MKb9mMKJk5aZmJdxIZA+KyXv4y
Bw14M6vvjaoqf2l1WeZXgGII+2phLtMUUYjHzhyF3ghKRQLiXUJ6yTl+QothxLlZ
a84u/5gkBPEHuXQ2zCdHV+BPVN4cXs0PxPjovmpv+ViY5DX+5uSTXdQHiGz6xXad
3jTGT3MpkH+bdUrNmUXvr4jX28P7hQ092N3tqii4qMfB3VQNx0jagkLBscSiSyqw
G69foLoH1sZFsZiTJi+RIIOn0W7rJzLjMZzr5jlmnW8Jwf2BrZuisPCZD9mv10r8
4SISWBSfCYFjaJNCOkBGw9LN3O1ol8Fsz1/Vv9QCwx3WoYBE9cKTGqv7JmCy3LVm
E+oTxGFj58GZE46h78/Ar3c6L7qcg6ajkQdFhALjZykKQn5zu3KgTrRyS7/pfHvn
HiR6VvDQOog9UKjzhsWndwP3qFlH6mYeNOM0JYRDM2+Zto5Xa8VBL+VMaEp2nCPL
P6CBRDf7bMWLiAkTZwqMDjcrIe0nDSFpdsH/xMZjYItitavucTK4e9ClOO17b9N4
stzPu+Ep7j8DMqgwKvoXArHEOL6M2O4KryAo0dBCzDYmnHR68mDRfO3F0xEfSfAU
iyO4l0EGDpKp3o9Ee3guggAmc2GMc81bkay59HupP2UP81JWQJ15NUSueQAK/19b
2vtxbRm8rDgeOIyUH9Zj0aoXTdkQ/Q9Mh/wLjwuqnLiLCkd4EN6xDNYuxxdtcbr5
1EXamjMTTQP9zirylzgkmpygprnCQmhQ0h7YKIT+viP9PeqtdSX/oa4MOU6Rv2Iy
mLZcKF1YMqOwswhHboZtrpfed8QKKBwFoqL4/xaNkmN068YjOFopV7tF1Jv1tH4T
XrFS5ElEmkUSt6NbltnDWIwAmOpWbGk8Kqh0Jue7nccl+REOjoLPB6yRsXWGs71A
dSG/e90ldYs+pKYOcmgPBZZweBwbyiOMTypcZDX+w5V0rsu/IpTAFwW4nuKjz837
Uq54qXUfImFQv0QxyU01yztQ4yP67x033+qRq8He0OBRFnnG9ONJt/hWHK3LLaKY
KSU9oqpyJK3tTmF7UFLXFe6U/xZgHh7umLsWpyegWPxXImxWeNg7XF2E+KaoInWZ
mvstxw2JN7aQEedb3ASD7aOvpWuR3ird7D3LicaGLnS/9VxP/23mmMnYbnpAJ2qS
TOkD6lGGDZV0Vvp3M5L8CJbVjqcGkt/zAPi7q57vr719ejTGDk3fG8yi3FZne2al
YBqZHQFIuRMoVx+G7dZtsT2LNKP33K64JNAzSjScY84mnVVVbm0cRbrtN09Ah6lE
yUqyDDZrkSt1kr4fmZ90IiXe29n27ASDFVf5sDN1lfRFlx0lGNHaDwIUwuff5CVy
KZBSCTiWX8owX+GJ3dKmb/wYiGumLvAwXOMzjKkeIJudnZjGdrZLqq9/cJaM+lb9
n+efujGHSaoSJ/bTGQmKUwTSoH63D5Db3sklCvizjGZhLGM2GALodCyEEXlqPye8
tGDMiSSIq5dAcoTdwtSQHQLnMT92GPrjo+rSlNvmSytno+sDO7BDVIot8gmBipiZ
j+96e3b2F92vFcthahvm6deDxu8hSt0NZJATbgci7bYZdA/tetTPiNfez3DOuunb
q3mVz3yCr6EOo/CHKYXvpYGZ6Ropxf+xc7U+Q+lVNhp8ZLOxW8N2zDMr9381r/Ep
C7rc0WGVO3QSWl+2g/Nu/0ThiniykTivrfkz9GUNNfpxsP3Gkldn8EgRxNisvBOF
oyIAkMDjVOwI6JNnlQ0KW9TVSSakv8/lH+znEyTV7WPYIwLiEACcElzg/aH+eTDT
xKjDN3obioTytjGYbxHdcoa7RGl0DfOgs6D40D73OsW3nHg8xvPP4RfBXVGmXXjb
dY6lD7MoYqYclzhYXYJIOjZOXPnXS8lrnBdzT5/AIeQVwqVHAm41MQQ4CIgGMeVN
mYfaJj14Le3p2OhnW85cBgQYy3LfJc864vKb0gWngajZuDK1FYnct4m2A0OY9da2
awR2NqkZfMBoBayc6o7dGEkv+Ea6sIcCMlI3j/EzPDae+hVKvKLf7XDKV5nHkS4a
eAVCRoPeO6wVPkFekFdNypA42oJEs2abuMSrTbuCPQj3YOwqTm1UTNj5L+XUG0MY
t8LJx3xqNQiLgQQMZUr+dVDiqYE2F05+KoFV8Bzc+DeFO0DZw1l0aVbIctYpzkGo
oQt3x/PP7Xs14Wn/89DyTW/Ey3pSb1rKetGkEsoFitCQAh6iapsFYegrMlRiuHCF
UnzqQI8DpQUCh2dizqEokbX8G4cnSpN9DKEsN0++Hs0rfxgRMwlJlGY0kBdxAcR9
l9ixEDrKGZx8u5GslJBNDc0qfhE8WkJcWyYBwaug4umEKlJ9L5b43YfpiRDWg+oA
Q0ctND49rJatwcXfCus28RtnHh+Fs+5xoGfegV/J4LIJZc6c+L1c29TSfQd0FK0Q
UgGavKxvyuj8LO/XlII0iS4Iez+9X4kV4Ols/S0s6oaJfiBvD8cC60mw+EggdCEs
PgPaxBeu8vx4qmXyxaPE+ODsLBnG2YManPI4SLkpBDfNv/91NpUVBuZxESAfPRYZ
S0K+wI1g6FSMigLv+A9ZUBk0HEm9RdNCWFYJrV4gHneEYdxeUG/x8hZoXGjhWUYI
lMCgo3n6UoriZgY6Cbe1GNISLYV81FtIsMU4MFJciKU4AbbR88lsw+sxQG0TDPw8
Z4gdJfzQfofTV9rYXOwSK8oYXI+qED2K3Fm2qeglhFYfRzMFaINMIgEmCdoY221X
WSILIgfiWzQOWCx+ynlfSQbU449G/Gz76I3bpBaBm5WWypJq4aFqYjMhgisfT5RR
LhPnEIMhkuAM6OBjylLu7mZHSG/Md+HRHodxdPHcjPdFXO4d4d5aQ2v2dtjLbAAR
73hZ+W1+DOjC5ooIzDd87IU5SikxOWu4z/Pp+wo2hjP+IZ8SJ3Ug1EQUwLvl7qf0
pHkhJQzZXXktY79PpsL1Vd/CoKUsbhZKkg3OO7q7VgvBSwIeW3p737YzA2ZkXbKw
pHMJP0Fo+om7DIGH9D+PXCUMfShHFFnC6nxPo5rmwtvM2gKnaUsuHn32VJrr5xQM
Nj5W1x4WQWvDSAx4Q0SeOhVrhxfBBlLHCeOEESb1LY2xtvUvX/7DLAtB3tSl7gl0
vsY5LHLpnxGLQwrOsLpY52t/buANBYvI0kS63ErpxZUniV+HhQn/Dgeix1jMZari
FLOW4RSOd+no20Yx+GGzXBw0qRQuKq8ttNMaiBFNzE833ED9uiNtva7JNRy9NwKi
YM1FTmxE6XhmrkFIJ+l0VhwLDHOlg3Vk6iJF6fW0eSUlClVPpGcg9FUw5imCYyIY
xZLqkqRkB0VAKgDLlcLo+fsumYySRNv6g/YP5j+c1fpn3lRhMtARTAHFJ+a9hwOd
6T0Odjw428r8tsGjeZB2tnCHbv+F1epl93R0EcwmJwlPW0w4+3wAWQ4cXkDhtIJl
KBq3lIqBs3GvB2rvxLXCVhA4FnebBfQAvjXnRWT7xgSPvvdlxmStj90D0aisfQm8
lbYQVYkaWGN5dHwphib3HGUJTY550uM0aP0ngDkc2kW1PO/OzN+jg1OYCgGs3QYa
QA0kII1aFo2q7C5TG2R8UyV6+P8iqZN/3exVyePORrDrDVtE23yR6xEWdOJgxBYC
TcjDcmA3i7x0ii19qWY1naZe/6rmBuX4Ua4eQt0RCsUNXkPRTXhRDCm3lEpvXsTF
TPSxMYC/CnwJVS+ju1lCVOpuf+LKx6Kmoc9PzODFMzz+XkJ9fSr9BpSKr6kfEmdR
3e3mFvLIQZmWrYmdCvZHKrphsK0UqGX3O81l10+hV/iUKkVVVYm6v9jtRnVlebc6
RLjGIK/E7qzoP91wssbJrfDejXY6Hhqc7Ic2I3SPg4B3xvLWzvmrHu6hy/ppKuz5
DLwnUBSfg7OK1EXf+TLeJYCLs130eiA7rtzOKbnFeuI=
`protect END_PROTECTED
