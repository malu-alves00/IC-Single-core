`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BrnxXQUWRKN5wtBDCPORwi44TlPD4cU6GJWwpyYQDTJ4kDzd1keiGYbzOyntBIMz
/15buIp2WH27xTm7OrH2Z86RDSkK22sOhag29ETMUUe99OZLXoYncIETYcoKhiaT
pHkPgKl71f+HYITSHXveX5ZqTX5+MMcHWJ0cYpwHby23mT9WjyUw8EDCFoUnFi1y
6/vn2WEXCeeUg43T9kaLos1qnW7oZPFaUyOGR/rs7h5OMN3BSmkboroCgWalYiVW
wtNSRlaKOBD7T7H7YqFfOi66jFfEjyzOg4/PrqJgcAG6rbkpQBbAMNzVkTrrIl2H
JKmuVpi5qpKuSUMJrp0DIRmj3V6HobczKpDai8uGmp4lbcdZzItts1e4VmKieGjO
7Vl9jq5Z/jkEM7ljcqUN/SDX4wqsyvAQJMO8qKUj3V87/NT5QOz3HtaCrrhpkEd2
rXDHYnEdwM1Z24UHHJwa0XrUJJs5696MQouu8DlC0seQyY9Wt6dA3IgCGJAJUpIR
XSBbcuTSqEJSiWbM02R4ASVy8njLPSFvphYNpXclDcDJ85mN8TXGe5QIxqw7SY5a
/CNxNznDwMz9rzpha/0kbPwFBoUGkLDjjy1IMcF5+cYn9YPyBzB/SFSxtSgdAoL2
`protect END_PROTECTED
