`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
d8+XpQxd5lvXx6aVmtYhFIjOwZgFtqX93DGKb0AQ0t3vDjxke4RLC80wBUBlvnjB
mfhAjpnKZYzGe6RmeCCcbmNzKrhE4aVnFa9BRZUCwJ8RS2u8od4m1Hb7Vcz7yYU0
wsGrazvfn6HdeV/XEcQsdcAjcwGjN4wgBaoZwYvz65XgkRFKpiQMxTz2uStdVz6P
ABEfbQEmE9fUKfWQYMAWOCxVzs2Zcia9qG0apZcP8j7gDh6p7cOG0IvLPi4itRju
7+GTE4gKdxMeLjdJN2go+m1I1gKdtl+RvrvI28GBBeJacozaBpKe+RPkTsVEBaly
KQBqE2/BUCp00VDAYp5d4JN3h0ANaByup0q0igxSDdKDmzc55gxrQ9Ikdd+UKCrw
wZ1fDn2QmzCcdISc+lWO9HjvKrFjZWiYBrSxHtLc4Pij19BAn6ntqtWQ7BFuk+G3
ippfx8B8mSc5JBfgDPp0zFKdMfddJrngZ6/GAiPNziIerbZWhogougG78pj9w+NL
C1N4hclKkGBN5vfoorpN5aDdYcFHG2pq3ESAmlCDGpzmeHKf6UjenR9tEs/AZxIe
wt3c63gubbVQdBhffC74RQhr6zwZYIhS1puFH5H8E555Mgf2p0tFCk7u5QuN1JS8
K0lOjFhmVlCYNHL1NBcHfix8gECZzj5ZpG/DIPei8FRraY8XGYH6kRjI59PNM82U
A/nJaidyeUPKQZn4jVKlR6iHJNKDfdOpPPD6VTAegUejrGuv8rlpzkf0D229rMLA
RnHQGOIgOZN5orjkaQQrkmmrc2IMK2qXF2X1SDtDqwZIO7mZTL0TFV7OjPjGqMNB
8dUWyg9byfZ524431GA0Mn+fO2LiapuXUtSpCanocSZbxo7s1O2KnnTQrf1FO9K3
fC+hS96FAYeKhZ3iR4aVq2jiJXbMrdjtY6ClW6Pl/alg2PqCrpwCAXauVO1aE+xL
4VRMJEBmjdOYN78b92zkY4quIPfw17EOI78wPZckK3GQiFi60Nszsg0DzzlFF1OS
tDX4IhIm9KDrk2gudyR7kztvW5p/HV2/XY9jvOohqGVhSUfZap/a/oR/V8L08KNd
JmqO6tQ2DP/SxjjfjFwwC5NkG7Sy6fOYpPmJjXr011zfvzBxEnH6BP6qjkTTUUCu
DMOpAmQIV0sjpHRCh+MQjA==
`protect END_PROTECTED
