`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
D2OsjW+Gy/wyK5VKtWUl4NMwI0e25dEOY7vqV0jOfig2eq5RPHXV6u8ymB7cd/6M
QRjpg0MkoHcoOPpqO6o8CKNzGXasQN1/MLuUmYb9JxeILnAqEaZ0i3C+XFLAV0a0
Wr9K8nhic824eLTcNP9fBWjqaqXA4bIv9M13cL/gH7JRRMle0Xg+oHiJVx/KK6ba
HjZifIW5icN8wnKI98hFTG2HQ4rziVgw1tPfuX45KbAwQDxhTSM/QX7WF3lz91v/
Y3EsVd4B66jGDtpbwiBzOMgdWHbXJAO2tlEH2twcWtK+OvJoNZNmhuvwwhPXKoPL
YW17Z+03alFhzPnmhrDiZdhQE9L5MP0pOu0oBuocI8ZEm7nrRTBjQTw72tmj9c+b
KeoHmJU75oVfCOOpqLCv0OIjzStM4DL0sYiF5YcQOFufHN40wsj5nIeD9zj5QRxz
SK0ixAVDou2RAGke859wfHR9Pnvf9ocyu2qEvINk4oPsZJdEkHXpdJwswqGmA/En
aj4yZ8+fkfue7/U4WegyPOTiX3+NkeZrdAVWIhqLQ04/dUxfoC1kmfiXAFeaVwPn
fo4lyY9MnHTVZTDtv0030fw4l3ZTZUUku+OgUX2B0kPA3CfOKlijk8AMlLxU15yy
g9+lhxQg/+5AD5aJy3L76+rGdsjcpM4nJT45J6kNBj66QIK7aLMrjFzQ6mDvqf9Z
MGDl5UjHrPIkRDjMDWTDdxycLXQIIo5BSMir5wLymJDGgV9ik+MB/+WkowrclCxK
4AH/TgZlkgDjFINZpkP/P+jfkMaee7RHIHJ4xbtwjBk+JXzQJ0bp3RmnerKgESBZ
+vDDonKBtYzhn50vjMCZQggkkUNhVl5cnxf3lUYEaAQJKQeE7iUjg+XJ+pnNUpfk
0WqoFpnFNjfc9XpGhazml38PTloelOYyVMbsynBdIr5AUiqUCj52+iURbROGHdj7
CHbCM1/Nu/cGEiz+CfwBvoAFNXG9oiCny64n0AYp3ydhaijnW2I04+XFAQwvpBv9
q5Xdlu0ZtaeXKgk6uiCZltI4WQI6whfeS7kmYgiCfoXUMtb5YF44VPbjYcCnFe0s
oXP7vtz6/HVhIfmKlm70nHdgWrvjm0J1tDRIBqiz1t9NuwpQFWHOcF1ITa614e2k
8aA/MwEq5HK8kwtXMc0tcwt0yKF1P5xLgzzmAdGUWz9WMmn4jPLrXDgJGjtm5Nwh
YuECOkQX1wtkC9ylA8D82saKjUZlZDfEKpyBhNGRPjDdztwpqRdFXeKk9Lc/5Hei
SAjATU9bhzNBK4asdudmzlXfPUnS1e3eoEyQ+9rflHHC3TWPPvGUMivghXLn4JoH
pGBorslp2n5qLkzVjYDnOXZ3xF2HG3Oxjd9ZNuW7D+oN49tZ0lLvaNia8qkAOp6u
MMvd8FDy830LmXiTUT/sNS7F/Ti/KWE/ZuorQ2FbjVjbWRIiC5NImuTB4+QYy9V3
p4zndVJFb0Vv7hZSNTALK9L4r7UnkgR6textwdzNAtxxH/+MCJq+HLqgkNAeicJN
ZJotvXFG/9hSuKgNQgAgsiqzdRVXLn56gjrJm/rdxuaq+/jsHYogb9bhMGAxzLXh
/WYc6StPGbApDHC5UHLK3ofZCl/+3AdvF3Vsg5JWHQvVrcOj9j0Zs0ni5ZxsKo1F
CnS2Q70xrCuAeLAlpwUpz6/FJAJh0TnWTCeouy3gVwzEQIev4Ir+HyQDFGZB0ZsW
y1XmSbK86KsWHHWBzDOAIXQ/jre21kJ3YEYzFcOomFZthpbi/QCV8o+STA/o2Xl1
bRSnfH8aW2/83b8CbKsRkbhxtlcVPTSQHSOdakk6aOGGkz+xoi+gWctpUnWYbCw7
TUZpYE5lxARczETmr35xhUT9kU3izVo6JJLp1T6kbj2RvBeUYf+kx7a3gWR31u04
OGWny2TqIKsZltTL/xBLQzqbJ/A1uQw8JDT1wYS4/6YGe3QOL2blh2nUpmwlRNDe
Dy5XoDrsN6z5NT4Q3q0h4ZaeO2Ostac7tk5n7Z82JoNbxcSXTKmUEEkQgDm4Lmtj
hXOdOFqIL1enW5AkAEe2JDUeYTXaXTC/97pP4nLUrrNggk90rZidyiKX2b0mA8fe
4jmmsqINx5lcHewyir813JDs7jH1v76/lmS1aTDHKNBpTqVONthMAMVdepsyfo3B
KFi98ETjI8ZF/s0i6+4N3SOfdUAIMfD7fIOPAFsBwtAjFj8oSALMYcqaRGtrlsDE
BhMg/Pf2uvf67zOEyVFQb4vXfDMgK5F8pHWxFJeGnhQuxxcm14f7PXG9yj45vSFf
8IVOSOuPteJDgBL+b9mqOAcF2prh3kUeZwUqobYaHKB7GjAykSA+BRMt1/gh/GxN
ZKvj4PlONoNUNBpP49lb08LK70AQicK+XKk/HRRptHE5Xfdfh780kJBFhlq+wYAF
swxrl1+oOu1OsBTrF0Ee6jut2vs5iZmZrZF008Fg9bhTR1N0vGpSxSKvFva7xDd7
YefdfT+ZHSQ86Va5qj/Iv0Y0dpBvhRqf7SrFOOY99hINXutGXQHdz2bEkb9l3G2o
0Pv761YmyARLwplCTmy6yG5xwcaBDQmYUPnl8i85+OLqDsnmPMl5aTlMnAfBCNJF
4wZcPcdxKAMyQ7FDy6prtA==
`protect END_PROTECTED
