`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
b4rpWbSRSnXxyJFBMnON2Q4Mh9GZaC6tILByYREILmr1RFKnz4cn325drGnTptGg
WGfE97520h+dUiq1KMu6j7EEyxFBvG08m7YnDcR7ptbW8S7d40DUIp0OQ7lTq6Qg
dsafdRU1QsGSf0KT3IhH3P9PlaIbF0ZNZks1sk2Wdxidigd5bqzV2zRIdy94oAC7
hb+MiNAHDKvS/oZZkxdLRSW2t/WJ/kdQcJJ/r+9W4Mg+/droqpIpFo9iButB9M4k
J0SwTqm2I4I8rwBawqF+PoCVCNgfu9LpqzF6QUQOJqnCUlyq8pkzWT5/IldGc9j0
TRJHtoucimd06LcrDW7gP+FNRwcaLalfXUEbm3nCd028Q1wsE3UKDO8PVVgkALXH
f9PVijmenpvzMBOAFMs5x52hRA+mLSRdqNmYKUKekrP46b/lIAnLFJA5I/7cQLyB
`protect END_PROTECTED
