`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IGI8KePpH+uMFbyn5mR5ZAlppEjMdpS8J09B4BMZf52eBNHl7PkTXMtII+ltSeu0
RtKWBOcXs79CPv9XFGgGhyfqe3TAs+ocF6FzoqzECnNwe1EiB737+pQ4tU3tY6qL
duYJ1Fk1QrQdN2wlftKFO3IPAc3xQN7aSdQ+cYDSfnnpl2vk50IleyAMPUcxBXfL
MGoML1XYu+Iph1/jvuCLUtE644103D6/xSNrz2q/dJuMf96YTiISw47XTBGDKPwN
DZiUqFeakmZ3lZOPOiCkBc4bjXY6R+JlMGokWF+fQtEUmE5V+FFZ7APjMdi08gvX
mqmVoeMKaqJWiHp1CHvPHQqmUUEZ/+WqSBnYNdqqnqm7DD0H+VEUpmr+yMgZ7LDk
QV/YUUZh49iXsaSil9JdS/fEFHnPe+LJGDCb6mRPuSCbK1yGR/9EmJNbjHTPj4aZ
7LTY7jlxhgcaIVtuaqHx1DGeyh3wYZfcEW85UFseLYTy8Vft+v7kSE04lhbwWjgM
9gf0hJYG0SYFsHQnTu5JeajuB3ZF8JdWLWFURC8DYrNpjr8vYxoRHgUqNrU4uTmN
/3SfLbyqalRwKl2T6jCwMyEQ0s8GCEZr+DErZNbQk06Kxu7qZZXvsc7Zo+G/v7ME
N+/sgP/lgH7ly4E1mY0S18CrBOqWlfpi9bRA/443kdc9zpOn8DN0gG6QE7wrsmtR
a3mm0RmWG95lWcIWRGFJ2pYkMvkQdS3vWfQhhvUxBRYP9ma0KCY7PiHtGKAZzkcp
XhH9qooqk8KB9B+1xgvlbDHN901np4JiC3RUA2lQXK/W/h228dSdJbLEMpYvecfx
wpn2UkYF6CFqfu818MCykMJLj+sv2WsVSMlQ62D6XCF4KrHP4A/OFqWmnHoYyVrJ
48qyoe8EFMWOIpsOAUt95n9wxmHhNZAmkbyYYVBlYGm9jLspvWBtfcuyO96tV0v/
NcPF2S8YEhIdwv0FGmf2tZSgz2VCHHFMyrPOW1MIPsH8kwocyWFUhhsDyNMYzuEl
sAFMpVgi0JTRf05PMzwPmZTZWC/rTW5FFwJyyFnJ8zkB1MYAuTpB+lxSmpnYuRoo
`protect END_PROTECTED
