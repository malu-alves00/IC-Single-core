`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
e3otykdVbHI/QTblUcqNa05lEx5ZTBkytlapIZQVNaYErTZZbifTj1LeJdPMwoLU
x0NZHFh6XTTEZ0UWfVEK9t2wSjzLWGXx22TNwfEhwmprhOD1is0+qLm1k8tgpHyw
D5nwyNhUKg1T2FwSkD4Fa8JU+4S6lIuzmbBXoOdRek2gbWx6erO+5hrT9k7TY9h0
eYeQFo/ClhwAQZUsUCr1s7sQWkyzDHYEYQcsrATwbNzUxFYIjvSEq2kGPq8LMYr+
R0DsGQ22ew39+TJmVwL8E5rP1h3SeXuns/CNwlCvXKHaTMNFrWOga1SSjP4gKCYu
AVQAoH2Uod14fIkg0/fgmuRAQNnazaQZzS2Kfrc08jX3JvSURiNW221D2AcuDsGY
+uw6xLEDGTdGGLqCZKO6WhDLrjeguj8Jf4WQR4+Hob/siH8N211amFaXiYAWjPox
n4k04cpIWQnIm/9dJbCr89z+CgSlHtAOSzEHgZ5Jsg3UBIUHW7lJ1kN4xoCwQVtU
N4A3/DkrvW3x59fGKckFqOJpnuR9Tkvjt4K5CYMiVU7jj4JWIQz/pr/sRp7VFOZO
gtynBCqfGM1YXG0X6CZj0NoMPkIEbe7ShW7CCw22W15wg3joNMlHaMDfdEVGhZqo
4g9fkVf79PSBaFQq4JTLciCb2NjwE/Ztz3TWCtEJgero7AQg0VeYLtpDdaGPw+e5
EmiR+FL+j0cTXX873qI7nfpQSBaqwbTiTRwtnd0YPFo9EPou4uJkDpKOqV+acLxq
ra1wd1F5TZKDsKJxPQ0ULYqq7Syrg9V6m6GRr0KBWrLgmLMYLx9o5Tsq+R+mdzhv
DC2kzhzM9Evc/RgmPyYmHekecqflICtpm7q5TvGSbBfOE8OEU4LJ8plPKDpFRoDj
12cqKGzJWW8ePixZSgc4MLOpu09zJST1MoBz2k7nPvl0d2ZBj4httm3wo42qCrbH
0PRQOB65YVKYfEwR9a3t5Zswfl9n5bZJLLYZakRgPh/lh1l/aneNoDeQbDKhxoHa
4OJsTjV+llc19uI6BoQmrhBRZrnYBYACr1XmDF8JG+NthqagPG+jmuURVib8MfAK
Ok9toUnG1ZuuHDwhEiTTr4G5MBBla7ad4kbEL2IJaP5PuIbDgnK8Ct9xd2gDdj8A
KGwZldUIDBJxNM1L2Z2qQJzGtv1E96OvEbYZVqErpxYTKtyQMTaPgJQOXz8JTWYP
tOstmbN8zGylc2pLXupETc5E6PbZn3g8J14r9CreHYxqh2XNR4uwGF2f677nB++z
aqE8iiUTQLZXNq1hgBPvGgiO3L38a3CcQZx3f/bq5N4ZX7sZqbgV3MRSng1dhDpg
YshstFdglqOdaXE5URHdvWBAQRioGsPF1vHdp7Duo3Qp7mOu5LU5qmssNz9idLwo
9sQVEOx1eTjRTiBOqilnmJDTRc/8vWnW/WPvCu5KzcvIfzche7s0IGN6EoAaYlW3
vYepU2XHyQbuWJvvJ54FbXA+SkOBdp7OSIHF9kumVR53iVXkfjnRdidm//Yl09fQ
t7T1iW8mfZ4YyCbxnW5KMvUujBBCON6MZN54VJfFNWjCGDkU2UqG7Oc5WhAFYMKo
qqY9qBudKE4pao/0oKpUEbdWu/98CUkjln9J0LyaNrSsV913aEw4pzjBdcpNl0A1
p+3o6hZfXrElX4qFZo670e+8NVzkUBgnCiBYbUoiNgGhbH/FfOIGFPJbQLL3CDav
ivm3/WRp/9W9qTggnhvA929lrbxHvaRWDzhmBRUwKXD+gASJn2D8KcNMzIWbfTGy
volvVc6NTYkP1PABWCqgBv4cdcbjfhTcO5wPxu7rmcX4Cyg7jQ06VaQ/4j0PdeNU
SoxzRYhvcTknKwXIJohYcnzyHwhSteIrxsBGSxja5nl+6QmIC3OioS/vpVI86kpg
M5rFOOOo/QnBgX6ctd3EHlrboJnOfRvrnqYzJIU3uBNY8nJpizsidCXSxAsZS2Wl
/XegHkNESMf1lLkz/S0wwfpMayTKOF1NEmMk1iT9okoxlmy8OcvpNuWxjoHixpv3
uAnTlGY1rVHb4J8Fjf+IDyihhWMSnmDgPlKaK2INYXGDRTOO8TT52rzKrQvNeq40
lhagnhch2wBLvfbR8wevTsigwjwhPf3Fi356MD8rpEowec3sCa3uccE+kq8mapoI
EpIC3yeLiBDN4ptqhrO1m6A1GPQPTumGbK98N96g+ulhYjzBDv2mO+JvKSac8VEA
iYJ/p2ElbIV+Ht4ymwhBPDiXG7Ay3DGjRy+s8nxLRXLRFQkdbveaP7LAN9p30yFG
j76HTX6cvQwuet5R8GtwjpYJDSjExPvUnnjGQY1F3pvkj/PwCPT0AcpH1709MMb5
CHUk/7Fq5bryzN1/UXT7kLKgNkqio5izZVtvOb/+n5iJOnvsuDmtj3H5HXe6Ilzn
+P8GxnpNag16TIHXqh19j24B0NFi4hMbftU+XmSVU0cadboaaET0LNbexugKEFq2
Et8zY82BnAlso802j3qxGhuq8hNpZ2tWPe/iieIMAqmRmAr3SSAnBecuU17VwfXk
RHEx7p0WySUGMWnYEXwvMguNQXcyNl9has+jCyRa4F1x5+LR7FfHvwX4xquL8pSy
t1lutV+QAaCyKtC9bjlwEe9FbXNwBacNP9MBCZQsHVWwvO2F/rly+7Vn2KSTDFlX
AVQBV9ihdgob3Gpc1+39AbGA0qEcgqOsziqUzK9ZabN0NgboprZQjndKqE8xz0wR
J5i2y8+Dz9D07xQ9WyTt46vfhmEWJZ2cKk9ZLd837Xi787qKRQ/jsQxMnSLI6g6t
Jmr3QEwr0uOv9/AqQbYZNE6WVc3WjcxG0Cg+gTQfUcNB/RUM2b5pgYl4AgTZMKSM
cRdgn59Tki4OI0E4f72opBVurcOC16yw5uUtRUkmbueE/rACmEU6YPBFvcx28yw6
8/W3ElQYyTYVCLKuDXRL3lBy376YpAJG28NQnjURm8rAWKxrkCp6Evp9XDVszJVm
KRAzGSS+1sOkXgAcEoxKt1eeXbu0FeAjOVzEWSKkDVTN1UDswARkv3qD60l/9rQ0
Ggvw4Nwql4zPpHyQHmR+Md+TrdFFpKm/1y4F7TQiFi3W/Tj2xTVsXrHoZXNDYXJ4
IV4rIoJgLSvN0arzribersSFXvqcPtxJnpML4fDPTKIlYntrbJg0gz8SCXOnxsrL
w/d3LAA7vwovt21Ee0RjeL7t0EfrzE8i/5rBmt4oDPFogidTy39HyfYsIwIyfzRC
vyEjWzoBNVTGlwnrGUTdQHahbhNH3mBd4aF8LVwS0F1OmtIjeRzfIc6QiYUsCslw
AtOQ7ZOxOHH1YlOe5146mcfxm+Z8GNQpChZjOYkbhVOV5/7xvdy89McUpZ/hYUwn
4bLm+KU577K/J4niFoSRRTzyXW4c5iAv1mooR+8QFgDqVyTA5Djwi8WQl6nAD4jr
Y3YnO38DuxoUlduZTP0+QlYMOpu/7H1wP15eHyde214+iDbHK6JKwJU/dOUE/BOS
ODhFi/gvgy95LcXijW1iSUDn1+P4Q2en6nJWzZewv+u96rf0G7nhSYAkPZWkTgBm
bR/Aqd5v3sUTCbx2XUX9Vkp15rUewNf99FnG/Cw8iM0Sic8eubzhVg2SLvlhNQ8U
dGp3S/mInWxMDkyUjTa0mwXLZwsjYeIPjBvCBljaZeyjTVBTg5lYGwB4xX30j8JL
WxxaJCV3IsP/EXUcwUGpKRMsoGemN3tuZ36MSiTIaELnYw77DfDQ0w+ZMJgYQ2bX
GMxlOlIPMqhhLebgVZpxrkwvebQTR1SiMbbPLGluT8TXgwk9R10bAQNqL6tuqwrR
v23pavDRCcLiz9zSaOLin/aaOg/E7dC607H6qW0FZRjdB1ZQhifgsH2H4Dzqcwbh
PwjvVQXbTfghq25lyQ7GJnsuCUsfGspGpFvQ9L+yRgUAvmALk6rgVJ70IWLPROl3
/FbzBID2Ho3KGciI7MJCwaA1zwfYczSC68ndwZDA4FALzQ77cSsXbmWVIPYdVncf
AQyp8fj8tmLOu1m8NzbXfUsmBJm/ZeqEvrWBq/9Q7ELKz/99UYk+2oxCz4836v8k
oUZNRerJCJ2hpC2eedxOYlyBdyhtQIvJMAHoUUvff7vbO6ke2SHvnz+p7UPeJfPP
PobjN3czkRicUdPmhlfVmCycWHuWe88Mi56s4XFqCdiy4tiYeXIR5qyHs2fxMw1T
gPuhp6tmMocios4QF537P6SBLvvn/E1iHLCneWUL8JgcW6bM+qg1tow/v4bQkMPr
W0/aDLhdxEvyUjEIviJbRAzB17+6QhJjWzyBsFP3N/w2rfg3PNNMk2Z9oJPnjHXg
pPLDQ33WVnNnKRUZ2HeSiz4E3WIi1UMxrL8DTIKn9/pr/CNsdVMJkW3XXfB8Lx7c
hNJOtdLEL6V7hU94LoVKIKAt4b3LVdoF9rnrlkQa86+C7L3nJBu1HAtvqus4Dj5L
AWoUU8Pq44B110ItdwBWEVEthBgckz398en2weyr4aBZIOuvxzMx9W3AAeeDsolD
JY0D9FG2RGudPCUuwntdn74FPEIR06m3YRzwwene/GOSWqXB84aT55zvcdwltPbz
wwJhpDzGMYQ+Qrfb2IQukhUNIzyxibZ7oCXnApwuXRFFRdIaHMPcHE8io6To87te
qCG49qEwiS6a606Kg6I9t6SRl2ya2ASSKpi9nWLeGko=
`protect END_PROTECTED
