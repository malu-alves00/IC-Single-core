`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vBXjnw9rmJO66s76yHMNCblxWVKcvDDwcKfDSkWN4J31ba2UErZ8+zhnDixFNiJM
lE1WTZOA7/zXZtcPlQxaf/yY4Xw4J1JeVnOKn29hxLGkAPowjRNo91US3DXOVER8
crBiMaAfpnXEcK9iFyXByrhIHEpmofvg4FLe6jWbnAiVWF54QXSL6zUGK3mcpA/E
vMqhNBbjkVL+3IQfFySFfyASEHrJh73gFLGZnwCYlGcfkx+v/3GxM09Z2i06QEJV
aCpp1sCZ/FZS/w3K8vvPkEHRN3g+HcqhGDVjgy0LZmD7wBybmxfo/xqISbvmNfOQ
Jfx5VWEMogcFZsahCikmWyxmtBHK0hONkH3P6LNiVjM6vmbKc9WY1dBt8ZY4pjJI
mfOEjael5l5CImaMA5h3zhTVixIJ6TtM4k1lDI1RNPE9G/PmUIk3llgmnZBmUXfd
2OI3mM2Mg3ZjSqwpbkuNr1h9NrdpQI/dGDo6rQ//B9WD7xnYdNfC7HzVut1YUHb2
wW3P2H5PtS0z1h/giEYJEkXB6EJbZu4JGOPJFQJV8/QN67J9LTjVBTGP7CaDGFN1
Kvj8Q3QeoxZDysSXNKetF8oT+MMYRHjkhzvBRSh2/BTQHp+Aq1nXeInxlwllwtH7
/XjwfNste5BoQGcB5z3CaWkbgnzxGkkjlARfnulYjW6YR3zltnMTmP28AMXqlXKU
Nh9oQcu+HdvXY1MkJcyInFAOVfWIX9BktWuoQgq3CVdDX/AQsrQexNoMGGUmZuhC
4EbE9xRuLYaCtADK6QmMXTQ9bAcGhpHVWvqsBBthbbBpMdsPRbA0tMsAlSPMY/yG
nxO3jBFsYFr4kQlvS7V1LrHJ5dH6MRqZpgeJBJbrQzxU/gnzitU6pG+VHy7VqtDc
ZfjzdrnrOpwbTAAy58F1+AveJ6xtDADM/CuWnGqb+BsJxQTGb9PFLoL8rmRF040T
/H1eRT0osUDP0YDhtHYdeMtb3xRZXrqCGD+T+6+gCJeAGEQ5dJ48wtDRrplD/CFG
sAxEQ5Dme77+TBtxW7oyVExRXs8vr9a+n3EnZcSYnXy1hauDz14hNLx8dfCWmZM7
7maa2v+tBa1jkWo9iGMZuUHwTSdEw7g2/EcXN+yArsTwQ3e2GDiSkF/4V+KYZ6cc
AFoaWJ+WsvkKe1XNab+ic5Vts01vBXhJFLqEZ7wveWM5XsicvMdCWX1xP5JhIXyo
JVHYcLOg3ehtU28QUx+2Jq7PGO5WgjOKm1i11aM+eX06oU+jVsbLfPJ2exlzriBM
YdLd019YDYfGS7qBH/GacPFm6pPn7PDBz2Lh/6wgia2Q8kMbuwZnV6hY7uSsIJSb
r3f9GD53amBxQgsIEwjyTBARtwXfi4VcrLwzUuj3NJukFvUzCgs1TIVPMEXNgZtM
VTeeZzijKIph3+UKtnc/CHYDdAgmxPLNzF/r+t9+P+iTKcmgiUD1g4Lc0KTcGTnL
k8fSy9qiujouMbQxCcWrwH1hOdWDxcta+kt8UfM5L6nmm2fqkA5cTuWXCOQ9cXjV
+Cg7WO2lATyQrMX0nNmujszTDz24f+jI0xYWKg3siPDq2xHrke/L/YV5wltngdVD
Qrc+LZE1vGioGyfyEdxQM3SXF7SKtEWa8Kqd3xqQ2JCKARGas7YW9xGz+KSJ62dz
cyTAGIr4wmkTprcpn7UlJM04N/FL3ZSt78aofOAo/kF48xNQJ/eRS+JbkRGcaPWv
uUyUgR/AXiddSWctxDEar19l7fGFn5HBob3r5N6BoJ5e/1ud/MYpK+7iE9tL6ff+
Kbs/DPz5UupR2CifUQ5aw4/EhyZvxCXfYRyP1/ahGpozDzib+02WwW10BTMVvf+t
+9mqqfpz/YXtxluYsrIWokRGqijaheP/99x6k9HDxgO5Kt3GewBDzKK4cohP7AqL
YhIlH+5ST7yg03MmvDZOfcMcx/AXRuv0O+k2aBaNUmuuIcfX/vBnz3+TPKeskJ9Q
z81XSTyPBO5JWhhmWdAlhu3G7pbSdONWYXt5OVXMCJ70ZM/EXGOXpPPxrpoRsIo1
yuvw+xegXBH6pCODQtZLARGgR1jZQgCGuM5+qS0iV0h5+M7Ngz7XzH8liTyifVWH
tmPc+VWdBYJX4p19KJB4LVMsm/b3rhQJnW2aiWWt5patZBZa2rdKnTH4UUraGSTM
txVJ1eRQiOKGsYsV2k3UDnkCDL1zrqYDB5w/8AroS6OPU7MkLsm8MF96avoBXdYl
Xd4ZO8K0vhVsoHgtFfhzfnn9XT8EE7OJj8mc0zyANJH/Zpdm5vOFqK8UvD1T94Uv
7H30iByAYh9fVgRDh/d7kmdK//7MsqfSTCgplzICiLBd5mXFpcbIYx+itg1R9TgB
Ypd+dRm2MqDAbSnENS41N0m0WnTIvVxPoBFojrLMunciym8Rml+dw0TQOZU8sF5q
zxmwhu4ADql2Qg+iQ9igzg==
`protect END_PROTECTED
