`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/VWk9X4aZbXu/jTUJTsuY/KbPcu6G5L8h7Xv5yU5hePXWxdW05RqU/NmUd2+0DXq
uadALe81pl0UfEGBuokxUpknR6AQd41qOHyArYZdibJ5fT3ELrCNJD2pBgTm57EY
v25EJ53j6CjHgwI0yOJhMcE5FFB9m8ucJRF8jG8OXKkD9Q3xBiwOJ0M1lxxmpovd
ZPqvBBmaO5iWdenb/wItAF+1nkmV7ubgdWVlfD/w4JqkLeclpCzUoU14+5l6yRQs
3w+HzCEUgQXi6NTxw+8a4364DjKm4I2arrydUBhW3QjsmwAWQZFJCjYMhJcqmgZH
BiQPA8jzeGXalqUkWzhGWopxksjVMxh2NqBalurGuX7ebJ+xrHru6glpg7SrzIMt
E+WJp3rJrO9Zm5hvs7y5Fzgcz8GMfsZtS/Ge4KJUFagsW5EXAaefoCrUsGGeENQ3
nrAQmv8Sip0vkhRJ4eLllzrssaakyty4Fxe9XDq4aSaSMsdwlmI8kk3z7K5ixi1M
dyyyFuwvL9DbopbULQFEjFgT4scocN1V/XU1ttxxXBlxcimqPMpPcMuPDN6QKmds
B7vlweOFD6khehnM73RYeN263GaVSvlq//m3QCMZcnhrnjrhddVEDw+jNxneL88E
UdlpbY3rPMtHFPopUnR8ABJthRLASGP+ynU4HTjVT7ZrZzssyvoUFS55A7zXIquR
hWGsQD8wiw307kgRLuexx+gKM6/j1LbJk+VKzbP4xJiDhY5tcB/ibJDXt7bC2Dy1
RU7WJGM4xLPa4mbnEwhgGG+cdaxhSErJHKVCjxGjLFENJy2X+Mc5GUSshQ9HkQDP
p7RvCiG+3atSutQfC3tXGKirKIwvzgZMvRYWwwLeXJ3kHQFZBfqjcQtUQcdCQffU
F9gDBmWWL9EaxooEUQ8NBef8W/9+vie7Gh1HsWQjJGNwIUN5z8w3quTtnbuApmed
xc7IHLmgM5jxrguxY6MdalowVfTJfTCYbnTdh1yz4G3fDvXnBDDoqzbvpakg5G4d
1VNyhuU4pFm2pEplUXhdoHqsdjYWhTF/dbKIFVW/SB2F8cT/US3B3E5InUvp0qnX
sQ8xfXTyR/D6ebQajX3H5d0d8pPU9eh1oZQDjaELNUCEofjeivpAbMxN7I2DpGJ4
Ys6PRnIknG3hrp1yQCCtSYI5glSkndxoOaSdFkdx9H9hKBGfA6qMIJiD0WF5jPit
NnzuYw5Mb7xMKyJNNHjvgAJ/X+6l6evMgHpLBE6wCIzDQKPMn0VuXXHuwxUJUuYo
yxBreYZk066059oybwz+A2LEGooy2GjdLYGxgQdaMjT24EDi/2k+/pXnE0iPkc/L
Z2337rnQ/hhj24s/7aX3CYSIGJLikEhcn+Qhe+0CT2itOSPdCUzYKlu4qvJ85Oz1
OW5zBivskJ0OKTZBQPnKBeBHQXJkYJDW6aBym9s1HI/e3FvmGGuCiKhDZibvE1Lx
FZ+mzziDvBAiY/c971SHtDq6gbWGsenG3vriWKVYpUdkBWRYYMChcjM18nd8bFEc
Awmmh3I3ARKHs38fLDTvw7ImNTFG7W5Omo6wAAzzdNYA7XaFwiVhM4ktM8kjYpeJ
Pw5vnvgvJ5NFE4yH81MZ7DusCuixwqkJZ923kjjwbasy0ftLTX91t78cxXOjmKxZ
oDmvbaZjkukVBr2qQxB7u5NJCdMmc8rSOv5WWtPv83/Yk4THy6uI8Bd564NJpDKE
2YiT+tOPxKpYH6QaYGwlY96QSsS8M5B/80O6ud5QHWyhWzIKearVvuUhpjub6TqS
yc3tssAycmrNeLTy4uGz+4e8paq7MbUboiQkOZ+obtJ6SPt19BIgiYvT7tf0ZHce
YOH3gumKsuvXmL+5/rXmWKpb8J7J7x9HuVtyosMZmlu2uZ7iwB88oL2QibZXiVu/
1z3h6JE14JU6aBaUJ6l/IjsjrncUTroBwGM0L6JxV1rhqhiCMowGOkd0El5dimTn
BRghOIQCixykbZTkk+Eer9JqHshkRFd4LVP6WhNDXTCtLRBF1CDC9yqIBtrPIaVA
XSHYKMQ86aoA8eLetOmgGSFP9h3GiycI76gIRx6NScfPoOTTirQPbIgLJ1zQoz5X
yH/RQVsm1jysc5w7EYHhNYRHEN1u/s1XlL1h/kaQMMq3Vrrcn/r0PG8VJFE84tnG
JKHPNWaIrB7XBqmtA7o/BHDRgm0QfmZPaNyQCXpmx+pbzxs5mUtMLQFFPh8CQ5Cz
fLETENxo59qRcOsnF7o/AhzvhINdLd2K6RUCTe5FIvVzm5KWV4jn8eyvYf+gCC0P
ckJytswkWfxnzsrMdXKjRynltm/nPrABHxnv/sqTELG2oTkOY8JgkszLcfCqS+72
IseQiRtvna4sdZ35f8JrcS/O6o0dRd5Sz9IJPktRWw49lqbmfJuN6WyWqtKTTRJf
XTT2qdNiC8VxoNmSHN7tQ25HX/X6KyUXwoxgeq+MokrHGBEXw21blcThLyoA8qEj
x+75zqI/L0ruxI6K+/0rdPy4FQoWFFatYgdjfGI0Vy17bh6bOIu8r1nEUoSKmVh6
4Llhu7gQG3uWBQOPRIk3IV45oU8tFUeqAIcqxUS+R18EtcpgD2jnKjdw36UQknRU
twG58gbj3WeQKretKqUg44c3h4lZ3IT4zJzG42gW+nBRJyWjiUIeJRKFHgDhgH8A
dBb/pnpuUNbTa59hzXF52jHRF6E/mWd2CZXsVFDWIOm0eof0O3cdluBRdmgcSt16
WmKh1P48hlUBFGsJyf3/OgfKfkZnnLZurAVibY11fjE7C1cN3rab0cLGtoTPZ0d9
UyAMK47iAsjf83MxjirvKkmQVguNQuewBtdtLMD3kW4zxBEDvFf5N81hsqfEi5h/
81XTfhluoNjDzXW47V+wC9vyRixx5a1lxiTmeigHqApGLQ1zpRZxw6IGgHiTZofN
pqhrF7sURqu29Cw9YCh3AuqtRkCV1Rs2QlyXywaprSx4YE80ewN8dQydV8Wn8rfn
ttyMuatcA9y6WvQ/vBjd20GXhfxoF7OiMWFUnEUscczfm127UcNVPHT/to0zb6tJ
u30eO11moWaCKwZ78AvOMBP4G8e40FLz49Ks7pJ9OLppPI72fZxYD40+vaukAwcg
faoJL6Ja5sQ5UlMyGCegjh+hVJOePjkINsQIJ+nHoJ9iMb4POAXMPU3LKLbXG88C
JOD4HUt6/BmlTEc4jhIyzSnIV9L+ikGVAHipDAq67a7ngnhuGvnCpgzQHbbsD8Za
aWkayUL+fJtBvZrWCMiP1YbpXEw1KTKqREeFGlHPRBlHy2EKT7hPef+mWnA3wbZ3
9dzQCTbDPqbNoVRenA+t1KuciK758+ED7mpv2rJrzAjh8cFdwH9J2pkQe8O8e2HI
HHUaoEFFkPG0OiXWctIrLCsvL4fTbIJ+Xv9paLYdDlyXMnQDH6n8uXyr0eDvOqTa
2kCRoehGdYHfNekKgnChYo4OyZPqkpVg20/gyp8rD4Alb/GUdWRsHhJMyS3DKcH6
o3GOGepPRQXWrYZsmRmKjcn1wpkweqH03KmVSbnBXpNtO/mS8cn42u/CcZFV2M0M
asHAtX5fQnOnEgHPSEA7v3zmxvZqhSGECf18AQEznQ56ttlBISu6A2Aq3yxM4mvM
PYyMDP3cAAkkqI0Y5SdLAgPKjJF3qqPikyh5gY9bLXOS2H2Vr5fPZnggi0Nio+T6
qNuxGqZPdqZiuj7ib5/4nM1aU6svRpwuEy2mE4ZGDm0rpWK+Fa3x7u/XeMs5AcfD
P9lHGeQKn3uTd400ZOxf57WX3H98LZrcQ6sEhGplm2WKfUliGh+hMN1vZcvB05hu
zynNmop0hbna2l/XsQYUk7fa0S5njLfmF7Pxl7I341MkerW3LsgtsyRYLGAvd78T
+euspKbQmF76zWV0PgLoTw5lEdpFarS1BNuCXMXsPa7CD/fraMtSu7iASIR0gMc4
2Add083yKcmH2UzDk7+I+B7D+ZPaNtQ8MwbLrL2TlGZOvOpykTZ3Oyip40ni1yFu
vUbd/8MIEQjUnuuXQprSf1iG/U0wo9tiNG7HHlLUqtvYs656v0yGxRRhx5pfn2hH
I/f9384ULD3EUopZ1QKrKRLq2Qry0y/YfPywltNAksbedLhc/o23L0POAsTZdM4N
7/DxVCcQx0wUcT8etxAqipOGXIZ70JrU/ET9jcIO6KFOmYgpLe5ZoSCqAXYywMJh
DfoJwunzuFa0EpFH9DssdXitKBChFFq51vC47Pib3IcLhx1rz3yiYaaTyB0RG9v8
ZEXiAwfk+3k6DCDuTKNPV4hU0cDUVAxy0X/JGpCaumMepu+LAIvBqCf8Dha6aGWa
tBYcLi9+ET9X6u9SNsxSX1jZ5d6A0QRZ1p88LdSlFncbVS/TkmgL/v/oVY5+TXki
MY73IrtOuVrwmdegQBIuEEdeqJCtshz6kvLeIzWylGfSPiP7PBFPpr0AjFY6WMW0
SsaQyl67MEIHidq27NeZhqBCFbfXdllrd7bapUDTjQkdAp0CylUpcLcxRXdwk84t
pyAT/C2hbzRJ4TwdgTAgsRltMt6l1K0gJeyNmGVv25SEOf1ZSDM18UszrEloO6bb
QEMwoz9PIqYfN7i4Hgo5IFsjkT2LbtbM9huzTKCePqQ8A0fkEqBZiCPK2EN99bQO
YcAOz9Nzp89zHEQ1vNgXjVqUYnadcjPGs6duFp7/Jr7FQR/Jb2tCNE43yxDqT8jd
F8MGFBpzPrefWNR3lL58I0T/VBRGc6uuOK+Cg/Ayx4DQUzy7VObdVcjOqc2+UqaP
wn5yjDvJQlUNNiTV+YvefbvQkdt+NxH23z8ygkeHtemNQLcvZFSeyjTFU1e5m72h
aGeB+bKfViHjVcLHawVcjHE/d/u8M+tAkeMeLvovFGF6R3kHzRjykTPUkQ6qTrkn
15pUvN8QRNfD9/wIa4/sxwHF/UZrA1UEdvG85HmvX8zvra1Hp8ykT91RBeFSLvix
eMxluvDMfDTRLcdRdsx50ZkR9VBMe94IDuuUYT9JY62GGU0usovb+BTTnvUEKQHv
jbLi+S8SlV/ufk2l9IUat6TdfIcr2+9Lt+fGrWOfW3p4uSfszqHwdjRb1iPy4dje
eeRUZ/rqvzxJ8EL7ZtnptQW7SmO2NIafs+P6UeWc4eOGdhk7h7V6S2TxkDhWwJ3q
I/RwdaGzWIQSd8V9x/Kv5uUcHbi9odJVLrGJETGaLQd9efhT8njr1hPM5ho3bzcE
hESNqDknHd3An4YqUee8TParSxHPMNCR6f776EyylvBXDjo0+th/t8pd7KB3pu3F
hs66HSQ+xLYTXMEtnCl6+In/kUFL6k/QLlan8aUK2mx+8ARSEJsljzJ57r4zPnUn
ATlgU9o/RNdZgpdSeUbTu52pZMlafNAM0FchQeBGyH2IgfSi6NZ6HXHx43GM4yXZ
aGBzfkK0arRstxdnYjztccgUm9mk8JPmIBNkIUOgdTojUZp7FYht72LWjA6HHtL0
efe6JEYMw0VCOcPFuxbU1wIdvNDQ5yP69WQgw6xcJm4EJ6PeiphAbQ/pSJS7Xizw
FNGzc9AaQmbCERJLD16S4ozIYe+VR3a+Ox6qLLZBZaftLk8czp4SG7yRGi+OvuIA
OxvEU7JLEuDzTjQd9fkDN/Z0zEcHDUizHp7/GSxKESQJExWBXPSFKGx1dxkXPgNB
LYJ6QsXC+dQca0OknUYIX6B3MA/dQuCmSGCt3xMcwYZbT3D40nJ9VHULAIRDTCs7
TsmkLYEOFRI7XbzohkzVE4+sPDWs8xtyu80a6RQJRAYvM5mW0YM3ctytVx09UVAf
QZZBg3RGTfD9vauRRDnONHTse9ypoAJQk2RxkGDo+idDfzMeCPG4nGqTdUtkA45s
TPN9hj6Q2XZqvBBSaAH/hrtIqo8SI4ZNZ06xZIh4piCX5X2iU8X54B8Fiif8/2IB
Cc4jKzy82m9s0AzZIq5OzYXBH0ttpZ5sUlw8XlIjQ0L7X7lLPJoNlyqpoCgOeeiV
GB+7m+jUHOt1gFE1Ii0vJKib1H6TE7dmY/Labe2TCt2+9BVbNhy3w9H2XefQVAxH
vugSFORptQPFJOQ/nTzM65FWYwHxIRvRyPkWg1xl+xZ8AWBB2/MJsGKLJ+qzKGtU
RrOPxrQb0uYj36OBYMzOp2F2pZez53Sxu6Cpk75NMqguZjWn8EhdTFCOAm8CzqQj
+30LGylMCVMCwBTatlSG9eieaXJuMrzSe79adv2YFRI8/k4voXRtxpE2XC1FyPDX
QuC5cvCspPYtBkO+O0SmK4hTVmbXQ0ejw/7qVvtu6RiZ/LXhCe0Op+8k5gUesdWk
nQuln3wxfQbLsRJIBoLLEic2GOA01LfWgptQ9sKMRD/aVuW5Mk1NE2zz/hLn5gEl
o5eoB+2x5ZWNzyY2utVkvEUSIadTd6BqtUZ5xy2Ydar+wAGWvcQQltGD6WdIXrDy
t4ZVaBgCv65LJyekEotbJP1GYFVVVwRqPQUsc+FTneGNAJoH+mKwNyLnwn4C+FhC
vgGuDrk/y/2/+/ZOaz0fi5ZealEnvgXjN5vpf5T312s4uffKTaZfDZX3rVUZ59xi
pKFD3zs4G00Toz36KqB/nFXwfU8VNDsbxVNTw4GjoBwnXpq/l9vA8bxJ09xIllSL
BUkM7dxA2USeIwvRbHdAHrvgjvGknvolItA+BHAX75UeQk9OPpQAP3X0aED6D/DA
AkkdJcRksNydznPlIcoi7cXwCEsqgoGg/BGmjGNRFx6ZmP717G40BcUXJEimCyCY
WkF5qb7KS6wftJ0fTbDXeRgFqrIMlQq9QY+/XTjbSp/DxQgT4win5NMDvXcpVOsY
a1BaFGm7MQ31dsY747nbjBw3GSG7IcXjvwiwCKymGZkXA/tExW4tf9BufNeHJXzF
i61x3Ig56soGThcRhZ7bMJlWTdhEYMGbOPaMcPKKbV0Ysz3nzKBk/jP7VIkoWcuK
h44Df0HN31uGmPgSzp9+rZ6dEQYGmOKShxdbLxSGtLDF7XnnFiPnD5ZmhCqHKGnQ
LA1m4qpqTOcrbdud7hCetW+8dMUbKdj+RmQWnB8XPzoYKj0hVNH49OOuZ59IM3va
xgAuj2Mccg9vIWTZpC1W1OTzOP26YM6wx4lzVZxlEPVwYeRywKazN/Wk/rUH5BcB
LK9pxyatkkp2hTRkvjWyL3dL27wDIRGGu/Ywsl5WgvF/jZBI/c58nwBl0KjtsV26
MOdHhM/Q7vwqSPjR9JmY/y8wFkE8yUlqbPYv6nkpBtu+Ti0AqgvhSO28Ev+ULaLu
mTbbnpKcjMqVB27WIK10dfPaVApUPmpMj/sDExPQB68VK3/5nGqTSnjJ9mfKcjRE
B0Ly3iPhDt8XQiUE/WbpUDCJMDo4oVCG6jl/hQySFETb0r79NWKPdY6cX1JSCTxW
z+RWI0imMcKVG5ccqW3b3jyF9uSTqnRt3vPpdfP8pnJcvQBy5w5kxU+88I8VEqVM
ksT1szXkoVVSe8pIlyDovOvx9XzKMN3LrBH3vmpJJW3EqgGGHAXg+lFs9wKy8rRu
AXIQkX2MrvLBIOwcxz9WGGp7GrvxVe5gFPEbx0OofpcXWi44bMGIGpgrsOSxH8Uk
9dPlsrnenS3GrjS2+VwjvcnH8pQK/Uo8852xBmlHeRf2YAuPdveUydqLn8OnywTY
zxOywoycwj+aFwkbDz5CZsrLMuOygkLd6M3KJT56SPp+Bezc4usKSOv+Pn/LygNk
LkEVKmikaLnvYBNrhnA26zoo/lDIp705QuhqrDzVFYr5FDSP0PkRxVUbsVGv3p7j
tzT5RBY6ThFtSO8+SFdz9jJrsg8ySzmkgoRAtk3w9I3VJjfo5pD7PryhQq3CYoXP
GIFmXvdBVo+a57iGHF9urzcWn8whT5DSrYkYEw2bubohvUZcuiTuvrlTIC7pjZiz
yUFhj8dTAgcVJPn8Nlh4Dm84g9XU31RO6h4DZAk93vWVuvW9HrQ8Z2j6HZ3rg7jB
MwsDuzk2Ypn+hRt2UCYnm54SC35CXZbi64ydLxOxsbjvZXKmje+RvSmmqNyleUR7
wE9EoqVv5Q05dCmtTTHy4dfHw8VpzdtHadAJ+LCZXUs7rD3WIn0s3W6s6BgLa1Ki
5AZ9Y9ffDawxggBvzx5QiFJcoiMyXlPYxRCtzFQdp/yT84RGeEZGbDt+QxqXyARq
S46SnURYVK1quRCsZSxZxNGwRx3qCB6PqpFCuuOzd2KmLqcL5uN+N9Y+mpfySgZ5
3d+RjksnXzsf0wgUrEN2n9YzdLdWIjWK//Qmwq7Q5zeoKTafyafnxQnatsv1ctFw
B7F1UuukTlV42QgxxWU5uFXW2BwocupvL1s4Hhdhm7n/OL31Vj7/BwTMPnS6Bjo9
m7qac+chFIzYcprxRluoqGzdNsiW2h4SRJM9LwQ2bBjFN2gobx21C96e9BMrTL+V
h3EBCuWW5RSXYRrrHTQ3r27IK8wR2bYNE2ljaAH7YVzoUZQmSbs1gJVb9pCM+BIw
Xs3zBdqch8jhkBH6/n4xCpzecKl4tdgBtnW+/mH54zYzt9yFqaLYoIcaTea6+OtU
uPsG/ncq8e4DotYTRaThfM/ATT2NLUgxDfFGOpcDaGiks49EaSJ+PmG5h3yO+9Gc
YJC+JYvvkGEAAMlCrEuHGhX9kWkWa8p1dYbiHRy4Z4FLe3fsCpqPwjYUrpr5lhCG
aM79lgQVT+V8R4isQzj6koznJRrmb0x78vDvCIKKCnfWVOoeo3Ahwbzww+VmIDhr
bX411hnoFzLA8zys2iuwrDjoMxcvcMOqp1XSvQc1CuXQ4r5H9TIdhYdK0345Cj9E
P68YxC3bz0tD+A6dnhCfagNxLjlBGo9qdMxds19FaDbp6ehVxMKO97xbbV6WPBZx
AjmzsUMh6zImgd/kIIwG2LJofKS7h4coIk4ATQtvKoBh8H62kjNLMXBGF5t/l7W5
RK+u6A7uyEZNCRV7+BLXvBy0N3r+WVqLkoYHVu63IQc4tr5qVycOkG2svEOV9/Ip
4mQ3Ewgccerx5M0vd0TvHU3iMhsLb1Pku1ORG23mIpxIeWCcFF6QjWjOYOI0BeCM
+3Rls81G5whVTjyH/YdRGPUDisgBLZcKdbthMspGyatVo0WnLU/tpwbTZFQDpsWg
PrlbLn28ngaLGWPxUG0bTMzEDmnxKqhSctOP40niO1lfGXm4UToErYNDWep+6/5S
Bs+mcTU34zZyjUfsPJw79RrMBFbpyiv5E3FwvSZ2q8me+WOCzuR+S2tu7BNB5K1U
D6+W/HOY3qEpE0C0GzXNdcjR8CKgczPGgf2JTxvzb+At4K98Ae+rp/ICMj3ue7ru
r4zPnauPgJ/2OYoUZkHE905MgNk2CFDd3MQOSFaEldZDOmfRxlE2AfUF/E/uVfVb
2MV7CTA9E6TOYbEk0VyH9Ax2pToEoLT7mSCyPprOVWK4Ko7QXAG1zioOPbNi4EK1
GQ/rJcw0BNmVd99g2BX7oMeg9EFk1Wzj1aYrp+dPtevNjvuym8ol6keZWLfvhZ8d
jF/jQ2k9TTP8uOAiJ4gCb6xfgr6YMiqWWjwjnbo6iM7TVVJ4h2cnW7KxCqheDkpO
L3MxIrms1TYNUFbM3K2iZSt/duoa0dtnFyxRvJ6Z3c3xksfwlvDjp/Z7nYMT0Cnt
PiVVM/68UT8wyzeVVAZ77JSNlpCWatREvcCghVRvSUZNVZfukKCykKe/tHQrl/qM
TzLDfcfEJYaZTDks4uAkiDbQk3VmWzNdHGZC0tpVF2ogm/oNZcmWz4LGFBM2UFZa
GZ77tJtvfBUy78F39yaHCWhwgy+8vbO9PKnZuZpWAYE=
`protect END_PROTECTED
