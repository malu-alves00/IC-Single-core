`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hOUPQCIW5+YMOw2aNnDmCTeGYW17COcrgGWiAvGIRUsQKG3Nx7ZlSgcuse+uob+v
z0Qf+igqKKx8eAuJNcD82MYDWRRLM8xfRnRuudkfa4beRP8IVwa/HLFsk90z60mm
1TsMI9HbgVDqwzgxwRb4+doKUH31UqrRBjJbQAAEj+mkgIdYIx2xcL/kAzrqzUTW
Mr98TEZv4a3WI94llamuY+XAi3jHt/N5HaSms9uTHz8PGY55RQuAjI5drOvt5qo7
HyXOs9IcNUCf1x737oM5cmtU5vprQnSaWYpIfV2ul+WmzcBMDIUfjwhjx2AHVohj
c8EwJj46SjUCAGfhxXK9llhlwr4u2TzzHb1OkRninKj7Z+W4p7FEGMMZHmoRPNK3
wyBy5dHNz4I2xx6WUqbe2g6WegizZVgg7T83FrNKH1+cHIrXplJBz00SfAzvklxR
pxAnRds4Sjs/IS8sjYZ/aRN6u4VI4GI+oRLyqQVP57fRFnrzH2KvJUNNXfzxhoJm
QbtqP+kjRp+rklJanPKQN1Cv6hRagqhgK3QiDlErQFRm6qeww8QVIOqY20377rMI
8L3yPz1HZpEhjvbBhxL+ulzvikWZZWd0yV1tIQ7isCSmBkbRXVGhUQMcLzLMRLGM
Xh17pf/RES01OuImibRh8rAdj8zF56GoKTGwrhhv4qn/W+3+NYg83zjC3sSpdAm8
goaACWXP6sLPB+AN6i5ffDKIV1gAC4gAcqvoqZviniAU8G+mBxMJlZc/QhVU3al/
WKPITul1QyIyRiLYHazCczChwBrh60zOpe2KAr8ghJwQrC/KZPSNPO3B+BomJY5l
V0nowZ7yHNjDkzruhBRCIKtVrO0AnjkDFyPXbJwXniPY27Hb7HOZ/BIFgOSnO4sW
Tg+7znVBTG622PmMKufujiSES44IJ63kC96B+9g8oXj8KG1fb/6KgMfwzVAGexdA
bWg9qiSP29XP8WCrMKQRZp0xB3QnguGIm9E0I7ZuYRiMgCbebYYM9CAxjS9jEEhj
IPMZq5lDdWKBzE3l4QtlR1liiQiD8UF1mru4GtEUYMmjQrMRrHkR/yuLPgaLc/Dj
9ilbYG862ZUSvhZvB2pJ84ECazsKla2dmcfSSbe02rEQMkDFKG8JbbwmjWHm3UiY
G3ARYjJenHJK3xK6w2WUyq5DAloBqlKkiZP2B2wnZbJxeVzoLgdfpP8skYpxIEF1
rGNWio7zetZFONPR0uvaVyAz4gVe8w0y/j2/2HBG4rYD52YEln1ptuZtvhAVd8SG
jzmu5tRB5yNpVrq1n1SrbpYB6+pCH8OGqDhb2gyFEpR933ApL93h+l9rS5XIgzUL
SWuE4i/ON/iEuEjEMLcXH7z8dS71rjQFs9Y3FT4EWl7LEsySDYFnkY0MkCgTvP5V
HfMHbqSzKB0f3IqD6OlFdUOOM6yJL+7Tn0KV022u89AwmOiUYNRolVTZdiQ3iKBD
hm4LrFqO0a17AO87ChluP+452pH5BZPtXcgs8k7PuOFO7LMzJDQSgGdcPt9RsM+8
Shf+Jn1sPe+Ec20eQ1e+IcxfjcRj/u8K2Tdr+Z7pb5XzSS+z9bsnosBMnQEIXnyE
wS2T2IBiollw044U+VQJUg==
`protect END_PROTECTED
