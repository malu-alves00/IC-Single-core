`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zcgfTw5jQ6kS7pRlu152reC61MsImixbEHV3vFCgRdIJXtsvNRBbQE9zvn3eRD38
wP4pnbbTLuyPae4WOgFTfpil46UURaLcgUUweHzP1zM3UetET4V7zIE8D2rt1iF0
UBRezDtgrAkJiqrL58/h3EDqEISuArVFG5X1eAIroGNnzrCPK1J/+i3TTxG1LTYo
DnDcvEGLT5Hz/B/11GIeH/KFBfLlmJdCi8jtfotZViWPpW4hLy6fvftebe3qqF0d
Q1rC2VXa/V1loUXCdof/7+2rAVaBFbc/6XmnnCMaIdbTKoB1SlOTZ/jdSCwYR854
4zrah8XKEHyC+n8e02ZMwvjrw+iV5F6CqJPv1uEpVHorS5Wb8xIMH5U3srPiIM61
r5+WKik5TyVi1DLOzXrfxwND6AxbIc6EwsU7y9szC404OCLRGisAiUFrVk2F3i6I
ssVDi59cvIgfSNK+zDBOmhUQsSTDb4gCViMvvWbwMh5TRyW6/IToA7JWDiQc23tI
EzntBfEcgqphlTO4Kqkofx7+hR0+Na7YKuy07vDk7bJPFqjuDa+XyPTSnCKNnvsl
TN5d1cINyWxxU10B7MCUBI+fT7g73v2J39NlplXle0QYwyUtRuJdD41WTyMT/kyM
aernO87a/uYg8ExFfUIbVNS8xbQcI+acWJ6N4zY8Twx5EV4xXx6Lhw7F+F4AbRBy
PvKwsBTIetnWwpV0e+vjNoUciZuxb0Yus0mV0u79ZbSLxT+Pa7ugmlhG96yW1Fy/
5w27Lsdd7w9aeCdcM+WJA+xZlTk4uQGR8Wyr8ti8zgWFYtostK9e5qLkZyCS4F+V
tMW4OqT8RFqn+yd1REQsqOPhYjaVayq4Hi0BnoPPtMn2TNsCpTfItxTvhRRoadIC
FbKF8/wN3tvTK3eY5rnSvRMtvb0TAF+Glweq+kHPALa0nTLxgxCXHkj9Rv0Tbecs
JJyCBAABC3EPC26rbu4XmdJIM5mW4To+hKDObITJHePOarMT9lrB4sEI5pdT0ylR
tsTdYWtVMyi2/mD0GD1/B3ju81fUqX3qOR7kQV6Q9QdjTe+mYH4E0nfRIef3lOha
ED52jXT4okN3fExpO1/VaJVB/JpQk5afUwjVt6w6QD1d9TT7IWOXxHxr/ZFelaYD
34CbXhesEy/daINmMr/05G6wr96S4EUXzHU7d8StVocD/zY5kuZUcJOpaZLWteAL
`protect END_PROTECTED
