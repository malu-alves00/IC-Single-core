`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Xvu2vges2uk8JIBoFiNiddz+rhsm7DuGxlHQefsdjSM42I3TvgU0Ft7gaEbK8A2S
LR5K6JKyxHrkeW1xQjpwtsNwGUmQ01EQOkDKlWuR47YY8+lKtgIiq1TksZoVzyPo
5yvwOVOOv4KtpBzAVaJWdwR9JG0Of15wdrB5fp5b7y1jovJxBTFXXYDyt9Vb6EPu
f14wkgxbU4+6DiMDoxZCMv8hkiJjmkQMPjt6zA+mVHOif6ila8tX67kTB9ArHM4X
Ij29hrAI9Rsk4Mny2lDOiN4qCpjYAgXbRhQzuypaRdu9h72fspngDn9GBnD6h07m
ImFMKEs97QRTGH+jgFOY9jIAIy5UPnXPsjVAhlein2E/fvGMG+opXbfESrUoR9Zn
wA47heyvNOmEorIbIZEusroo5nLHuVmqaDOMyYaumdXihTqTKz+ByIvShxRvVFJ0
AsPxRv0S+TYU2BH4YoDrtpJVQVqFx2+mQsnExz6dseHAqu5NCOFCkJH+5x06UABc
6/8hVDu+udABndX8c+9xyRRBi6BZNTbFZc38rQanqpj6C1y0JpomBsz4MJEd0YXN
ct7VQighIBix+dohDikEZ2zSCfEw9tX4JAL2RJGJ/HyNMdtF5W/Ih5rX1EHoOWpe
0C2yarUNUQ3uxhL3YN3LuV27lPUEqWq+cGqOL4558Cfsn98gRbEOm8t2Mm3BAI0e
UY/jOJF06w5JNofWJSsJtJVExddU2FbfQnF8SsmTpWQeXeswNDo+JGvlA20WnMe0
MYf4NHfmtMskvDU2iFHso7EUUnD9f7UHllY2Bl0QuCP6X9YoqRbCu0fmn0YcT4+V
whrgsM8kYsW+Rljha90DZKQ56yXyX7aDTYl8PhIjpGyZ/vwVZWveM/ur6fPGW0f/
T1oI/uNfKC53li2f3py/hZUmetgnMRmtlKHc/xn0MJHmmd2AyxKQlHIPhqVBermk
jOHiMWvbGNBNkHHpbBuEG1ifeus7RlG/GQkYS5/AEpZT7Bf710LTMOXjHbeZ650V
15s1Mh/GFIdldi3m8CR2edHrfCONzpH6xpZIW1bso7WDNkt6h7xUU1KyCBkc8HHc
krlcw+RVHiZ5g8oHQQD4PQnli1vmEm/ViQAqchllUcrsbrB8S8t9YHdUuFcG4eNk
X/swEJ2cCLNFx63HkaRIPaqGedIjr0AwuAqY48KIrcQfUve57cf/Uwdf6dOH+8LZ
d8cjkfgN0m0kmNgrMDR81lndKGsCk6FE3BilCEYBL4fg4Aof7m8nV7wAdWpeUv70
om3lTS001GCF0u67YQizsn8HRRlF6Bykpq50BYY+z2aCtHOzYd5V87OpIxFUBW4/
DAyRxiDF9tqKFu/4uZIdD+Ikfq4kT88QcyzVRw6vqf882VafermWSfeKGqCvJHZT
845K0DF2Fh4dxxG4z720qnulU97lCl7N4bitCI1OnIjJ3AAUz550gEZUcp0aRZNj
IewkgGMjF0m9YJZdT3Ab5aNOo41byakCD4aifJS3Cxn4+4XPoG2zzk1w0NIQPqU4
QkXX/xV+gfbY/zyXk2jyFKO383Lin7pXBaeQGivUKNAiLx2hwdyjEP3FMoMs2y0F
iorR339cNLFYdvjRFCFIWCsatqo9xvPOjHc6Vv+Y29l3xR4AJ/8cfj7obSakDR+M
82doFz9t3Rpo0AaW3cKFOL9vywrPGIkVCNalEBBOCNbnsmOUlIqaq+BODsg/MMeG
G6TrRDFYUsP5kmMOa3sOlpE6+qe42SaCbj7iyOINLE92ugIhfZ7dmDfu6ElaBg87
Z5jTrZ0UYybmabaFf86A6ZrEb8D36icEGvLAOJc9qnwYcXrmZEIGhmyiz++lWB0u
3hla5qpURE64NtJEo/EgMCo0RR7jhVoKHwLWWwXgjTeW9fBPbq/kEHNJc1S+vaAE
2azMwNYUbC9n69k5uPPrlJSbGGYHmlSDDEoo7Z0aM4dEM+p6SFKsKjNqfjVElAkZ
9E4sU5m9bikn74iiW7meOgEOoN5PydRFGWYDdahtaZuPgXBzUgLwPNpbvpN32iF0
4kbqBkJm4miSKD1aZvc3AGKg24deykXQsXiAzWr92DFQLPpW7XSVm37i/CepxsUP
E3RIEEk1+qFBo2ytDh0tlcOSdzUjc+dLhUKxDjFfGBKhSNEPx+ThFlSaNCvIpTyd
iXyuUzdkKqDEZOVzdj5DXp78h/XwaSK4QRSyOPBjEOmHj7IdaLcfQKODsuTZ0hcu
Y9kNHuDigmrQ226UHgS69829Owk+cOvcKsOLRRAtoFhtRB//c6KpSBpcp/LmsegL
cvjtuX6IQtanl2/ySu86s/gQkQ4Ua+ztc5lAN0WwRX7H5Nmn95TgYWBHgakKHa2a
DjQRu3KaUVTbMiAozx5ZrSsMQDC2n/dAE6h7scg2n7JaT8UHSk2fnQorSPrKdxBQ
lut1ue905JbgjWifcaIf5yAKXf6MQ3MUQFX89YMrUV/MkMrKYK0PuEmIi+U5vFdE
Lmnf5OXw9X1WeRwV1X3544FSXk7tfSVdj6HPP84bVXGZ6xh7L0024tQgEApq0Cr7
NThxPaHlKBviQxAaNh9tXXsKMGIMsRSakyhEGqIJniQR5KZJ7L1nOvu6qm81Zoro
xag8dGWfRS6iCzCwud5wRsDOvP+unnNe/jlnBFXrxzgPWuD89tn14OiB8ZC71Ysw
TTXNc5EBk+5Fi2eju7ZnA066kdtT9tNHxp06ckwvbi0u7iLGgjwBHSBWxMiDNpfe
L3cb3rgalUV4aGxi6LhtbwpB8xnnxvRfduESn6z2zrNk+xuKAUGpekYKKT7JPMzs
zOw2w/QjQKu8KQH60qvmGjaRpPVeZriF79HpUrMuD/8uAgKHfkssZybadkj/75xF
F9IYMX/L7SpGIbB8SEEGaOw1U2dvhKu8plYhIeQsChAqXcgq5hoSr8Bry5ng8COR
jSsONFJNsL1VaxX4stJwKk1kIlYEyIVxRPIbeY2V0nza+ifTQ0R3jtY5ejCmcugA
PrNQ++LPnD/BvT9y4kQ0lmkakhLVQ1nLo2R7RB8bBCE=
`protect END_PROTECTED
