`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2eMoUi9yWHj6pGoTWgfgJZC82LHlkAiFwkwTHpcB+hwJmtbxty27Wm7ntjI2gsJK
oCftSKT+ijHcHAZofECMg+aTk2/l5S8iFyMOutxWcGK8Q8392EZDPgrLg/0ASX4X
phYGgwD90+G3abo/z9MFtqyaV7mmZgfDG0Ka8PEx7S4q1TJidnlhbLaECY3b4Abx
QaVIPAnhUuzTzOCAgddunwX8XQAAjm2Jh/iXy+RwjLeeu1KQfvEVMwSBbGbfvrzO
ae6i2S7zQjgZr6b1iDnv82SvEfl/1L0fT0r6m+c5yNyx7EXHnXJAbI8FwFehfn10
hfbidp7jAohWUv/XGD8KZzN0P/8+lCUUwM/MjAC8jV7pvQFJt/ZehxFW47XGS7y9
nf2i2ivakbU5YVRU++JjqO8PZ041q/icLyfgzJHGJ1/jHFchEVn522Qsl8+sx5QG
fKPyVQthBMegv1pCV1MI8g1rTS+8C1FZK2ecZXn6QvVuWojAet4p3bIxQkKGrCmV
2vPEVsymJyaQ3AFQPKbQ2WJN4gim4A8uJ8lDR4bbHRKj8rBOIvG+kpTPol1BYLBy
9+MiQvk8KqEwC2pWndRC4crT2GlPpXJmMYevAqBmxTXuy6dzF5vUvEGS6mgw0e4l
9wijSmqtTnX0k0E7PQ3WM4lB75ANKtcbct7yrmenbFptTcsV3Ok1Vns0KP7hqW7z
YxYvbtpFRYn4wN/azzJgUKOmqPbsWr1ElBPh5y8aF8gjo7CGEO61TvyeioAmH+34
tL+hE8n+MXsftVrS82yg29ELw7y5cFPyBihghiafGNF+vql4Q4BrWAtMxKeP6kFG
HQlItyFEvB8T1xx27+HJzGTzxLqNbEllFMbTqvYCJIx7HTuUmKKqsie49FpnHuHm
hBaSud3cnp5Z2WClmLsL7LtgTD0hy2LN4zOwiARgLQTPByp2P2zbLOhkWi8YH79y
ZYk96KFsaYRuraopJHBODt072J11zx7LC1etwKEgWBuxuyptcRK+maGpkAegvTQ+
GHQVPY7HoTtdQMVMtahghUAof+5k/96qZgI4caGttscInQuDjT+L2nr90RnXarnY
2KlfIaEL77mnkNef/7ffXzo+XNeHxUaim0Ym1XOvy0eZgST66+gSEhwSG0slEWEz
vQry9rJqGJm50EhUlm/+jK9EWRRtZm/N88Jy3auyshskvK5xEqkxZoe3zmsSww6L
W+zGaUQm3Wkptoofy+cUM4bw8pV9LlGFpoAx4A9ZqfUY2UzltbK5Mkdp6HX62SrP
XnefDC0HBPUygZrQNhYba7IIMhg6TYRfQALYIESCMkVeND5sINKkOR881wjhx/uZ
8/aJ86UJd94OA3eoZPHVT7AFs5ojSW6AoZuhPgquDSbop8tV5pzoO7yUlmeZk1r/
2grMPZL6fvt3gfNh/CDoIWCMPMjxOsb1UBf1udQzdgc4qe7LZYMk9c7y0whXoCzj
9MDYd7Ng07qe/a4rYg9csZcgL2AHXNS7QhLUpCwXJdbeaSb7WAqzbpRGBBG3LXBU
CJqb++H+m22jIoffIi6ytnAty6mghyDJMHOtexO6PNcWuUtEQx9zP8lMdwp7s8hs
ICB3lzIBkjINNd9Z8f9K/zZMC5C5d7pKTv79doq7FI61/7C72IYYrrY+RxVV8APE
jk7QEdkqjlcva1zMfeSnfmNc8X5IAQ06t0bIIKXJXC3bjsK24H5grTGIlKyYx7ZH
cJxGbJP/Uqq7lGYAsPIn4MEi5NZE7SLS9bi+zkTBSAckXvvjsUB1h86s98sjE8th
IJXxH/iK2q3c6j215GStxFW+2jY+frEAL47gZuzmnPdu/ezo4gzvyOhao5mOadyq
Z/BmP/+n3X9ARjgLJPrWYR2Wu0lgBmaAjFZvw0vKciCQhcjuhZf7c3SezBLKo7Ib
tuhpzO1RiatH6/JekIEWlk16VoGONaYUKnQWCO8IRxsaRaIdTSIrZLnXyReefd7P
yIawzRJlIAZE1fV9uKMrhBdVGJrx1jsXBriX1JKf4A4yog68NMphbFoxklM5qTln
+1Spmn0iAKDo3Y+Yd/3TlRTeyGxiggsn63hKC2SWGUUEACjO08ikDKlU6SoFTjCT
ETQNs5hzNb0qFklg+vyxUKCoRM1KxGQdp/Va2zz9wHrYfAwdU0Fd/QEu3f1Dq6ih
CzeIT8oC5CsUiFv2x8SDSatV7tKzbsKFWyUrtdOp3mJHUFPmibFU2S2OUDS334Bl
zMhoOgZYsk4FzlUX9cL0anXw31Y73va+5T2jnbbxXbTYx9+c7bqirrt1ysW8n2l8
Us3dbDpFhgCo793Kpo2XRmHb3TF7pwqTf6MQqtMvTgzffhNoFDcvN3Lnc6RBpVwe
2kSpFiPPKkkmkgv9rnKDKywl573+UOmeW/EK587761ZFb91gAgmZegh8sYntoN5v
nz/TxjJ7ytiBHfePxPJtDB13qrrSggNxV2ZtZSQmOVioFiVtoW5nIzOW1rVvOLKt
tigUhj0U2SxbxlLm+k4RjWzhugaeW289G2F+8FaPeaITZeyrIYV9qRAPdQdLuTFM
FbgLBYS0EggpukrjfMS+pZ82X1UeCCLyqCCRE38/JUT9gZON56V1jtsLM7J3Y417
ThTrotQnBbdqNtY7FykxluCrt+z2YuA8lBXSFEXyEnT88S+j4MoPVRb3TNejaeUf
E1+4mhUSbEO6lxCYNku6ccliZLK4qmuTjG4UNv4rA9/5OG2AhjgRkwTrFX926Xtw
NF0EK/15tfrZmPicsGFs32LsGhPb1eNjj+BuuQ9ssyuIKujRfYY+trXkx7b4ZTHU
5OAsZs6TojkkSiMBm0pZa1efEAyBjptWVOwCKfIEN5o6ldVD3VXnGnHXGDuz9ucs
Kdi3eAaQihaERY3L4/iGSHMkzvtIGxNl33/96CCCr03HU5e48ZtK6wfx64wjw1Lo
Kw+OquC1Ehe8uhfa9xdjhyLkm1GbxvWhj+laJdDcZl9g8nuKS4aPqrk2xUYxKfdv
hBQ3F0C28w6NphsmDT9so0jb/MyCZwwCRFcdSaPMcl5Y8Py9kKv2xxroIx5GOPEx
FIM6Qb7KTaGfmfGoK4YntRz2fl52qDI3XnxGgTm8IpssE9h9cN78U7sWQuFXjFFX
5BAUKvZUgL7gH7GBXpfYLRnvAWR4WiCQ2QrjdcfqlEzhpurjPGK3o/lkWcM/+N+x
VSyTY3KibwsqL8O+p6BGbMqN8AyZfcWOJdsKu21fL7FvsS+RuOPt0Jp5tr+58M6y
QqJcBGPhWB6+zxGwF7CFxBjceJDwPXTEBOofLG9Z/bLestjXNzQgqdn0EpjXZv9v
s41Bc0SqJ3PNfMHG6X58x4aMwdH7PhqNG0CcAc8pBJ0j8G1fXXGU+ke3QGWvGq96
b4XLQGanTPzfW+qaFby28mPRyiouP3hiTZ2jCRUsNMt1SNx45ziLeBYRRUnDLnyI
iJLXFZ+HdpRt7tBH0sARvcONLEI722MZfsaoizdV9nQHx7v7Y++r0txcJedwEm2t
zeldQjNB8ZAuJmxqAXkNQCWQH2zuIOCEiPSBBOlHniBGWQm+6mXGfXHzrpMhfxRn
rjoh2Z4yRAQ+hJzrG54qxjDK7fgk1JLkaLeHpbEZwIvZUl5lIxri1b+q6xu9kDaP
TFAcdQrnR8inaO6vLzpkIU28zDWzlGg9j+ADeo8YsBb9BT1+bnJO30VW5ASxucdL
Nm5aWvgisaIVXEL3p/NOTsoGvfoeb5TjzJuMwPD3SLW3RebIDOzxV4lA33AkSJ/L
RynX0o68O5/PW1PrOnS1J87PM3HmQXdwUQ6JWXQuuzkJHPQh39JWRWxKi4OmrQ9V
Gn9Q+g53afKrww+4bc8I5weMPmZGSC/pcl2R9i1KQ8D6Iokq2KnTmmm8OLCtOe5c
tsvvTT6PYhSazEzPwEjuBYQyVEkD+FhJo2MnCqPTtgH9MDBckHoUUpoCVA9s1ZRu
E18ExNIpKwBO5rHTBwRd7XKUFo0+L2a7iYblODiIR8T1UG7xabNbgu/nzPq0GIYx
2DJNexPwV5ey52LgjdsFZoWCIk1Z57MY3lc6PTfvpkVbL+ICk3tX2JWnV3kV1j/r
sBn/RRvpLcg0MgtEvCTv9cGgjcMI03xg8jBzZgPhHXc7DVeD1oT3OWd3z5LR8fxt
M9TFOn/SQFYqEvTlbUt4ps+ayVAkpvzS9S1pHPJ1yeWgaajx1kRAbEq0Nfn9TOaa
BoplrMBF4EEEuRrsESowrwouJGhLbk0agFsvAVnXjmdITXqKLSpjSZ599BItSzFE
2W8FKc8ynwK6D5DOVcu0T01UEsnm6JCiSjx5ExQKAZUqWtCHUQrmpoXOXeW8iUcY
43bm9qIjzKHb2AawmLaFKJG3hL0kb9BkWumqLJ6ZzsTrCMWdMHpbaN0O3HZv979d
UQyaxZrdsyc1+6h7x0ShO/SmFROSo23UAYNVmv4TYhIRYnSK+KUZD7MYZ53QY3bQ
7PaEwXFw7BUI/HU5c9JfM/WP5TzWXcCQ1N20agPe5r/icF2lhdOp4znA+8YQRJ0q
ekWJ8rhTpDmZv5VZqXxMYup+hVjFAzECPAH4gJ0+D/Ea3voJ6a6Dxvj1RylkOk6k
vQ1eIm1mk7Qa45KpL7ItF2VG+Nm2XElV0tRumBfxJFrQp9DTnWukbA5RCOs7mgf/
0fmPFNNH8uE7olme2kzHcOmhjRZTa+3JRmbCLnk29k81NLdgeNsge+qw+SVNpLko
6cggUhnPn4ya3UDhMxGreaOZtNQlFtm39ZFik+KS8MBN10fXfoi38JRPbOTQOz+6
QJIJrq9Uy8j+zFypSMSJtiZTbll/oXZRo+Lo7V/bO1CiyDKDyPfR7v98tleHPJeu
SEJT3CnsDhU7KhBMKkjNzZQz7f2p9RAPaD7WV+YPoD/mC7dSa9Wcbq7iaXfce9zY
TIwbS/4n9s7gJHf0sISio7hrq2ruHJpR8B8MhlIRDSbVnxTd9MV98Vk6s2ec56mL
Y0ZX9yGx+tj+4UQ03RR0V+KB1e79R93K3R80TN+qL9SsMfYUzQs3Nbb48rHNpSNT
lgIh4w1B9VWnXECWpCgR2Mp0+/YDwdES/B9nmuSygTiOzpfEltaRX3fRret+P91k
86pFiVAAU7zI8a6El3/kAV987rbVpvNFQzf0Nl2F3uhb1farRGZNTSHCC52861E8
aENeDsGp5zicgbz6NcoDNiecVqrgohhWlHUqW9DzFRBdEmxiOTIbzTNrO1PPS8NE
XAH5Anf+7AL7gughAw8TzvQw0xzKeIiXJjBNTMiNVGrHrameTwNwD3gEN0QM8nfk
EbHf6Sumqx1z5Ieq5rC2tRaoL7zFpCf8jOOtooUenGBxTX3+8/yfMBHjgWVZiPpg
kaM+5bFhVCIb2tu31dXC2vJ8HhdXxvlBqMaPwLDnCB59vgwF5Ab7fyGdzSEs3gb6
laKLc+hqQ9efdYy4elS/76MAOUuBzjVAEoCV3YoGBR4+9PovWuZyh7Qc8eZTHAHS
i8OUn9CHbrFCeinTrpAb61aTbFZL9FbwYUL/tr4T08sHxp2YbuaOlkj3L55w1zVz
vUn2mknwxG8Enbf+DCUvhKq6Vlj8q7ZRPRJ6lC1I4nd+WkOqQzZsIbYcn+9MxIf2
3DJaJL8NJKYZbhJAsLdZKAznrUaL0gjBVHMYgYuIh4fIMwslzD+XtQ6tbsFD7NFv
TPpZ5vZ5AaB+vQ8KXuMWJ9DMgtHHgQcMmtoAJEJKPcQKiV8xliCvzksSHDFEVULx
L4PXTnC8BdNxHjZ7Hquw0K2kK8BAsA0Y4QjWLclXGQBPo74H/EIUXjVIFDe0oFo/
rmV1TSM7prhM6KFaEfGB+Na60uervuAr0LM4BDzNYr4b/1akVcV6garfzL3tCOO5
fRKF5Gzx7BlDmrL1cR4JPm8otV3YoREZnvQsIt/ApJl6vZBNl6I72FzkfGijKLlW
P0tcCmchSWiPRrUeSdzKzY228lPj5e00tiFtyTjly1nEepxoeK0UpEDNw6dQHQ7z
Csw21oJlrMXrkWK6QQXeG4oxysn+n7VKYVvA0RfT7ec1LZTWn6PDu+cO5ZOSezd8
cIdmmiCuYvxUq6SVQGnEHSRg7YnF4vWf8y4EkpmTwvxTS+gVFo+VAi0QGULFEjVX
uXrRxL83QI68WfC97nm5f7z+qowNaNZ2khfVgsLRV/4NyYvGC5Vvxfem3rWOwXYO
wbjuMy0Ik+VjxTswlFdQ5/W8GE2gr+dO7LvDGLWXemE3/YRM8V3MMbgSAHwBA7Ij
e2I7JSDgJAKfNXzouenO0D3P2aqLYbguesVMAywV4kcMQNGBzlNNoLw7HPZkKGaI
hR1B06fyVMPjnUv+jmk6WPZnI2QJX0CGiVyQYzTygNGhmyTK3WL+0fclPuxmBA6x
nIeslh7WEqxpc8YKW1E86sfSMLglXwlrDGMy126XZoWw6Q23skwlJYamEaJVn1sY
5ZV/bYi0w9gQ/PpPzm4pU3INa1NYARUFbtvU7TVGY0TEmNP0epAXTxsdrbja5l6+
TzCYTDVMbT4HukW6cQUB3izDwIw98HioVxiswX8qtPzokdWO05jeHKQNwpCOjr30
UsRYuC3ZgBvCySk1uFCxz8PV2BKJt6vagZ2almMvbttbj9YLd65qkonQ9M2QG4+F
I7HfKYEndViLf4qtU0WbOo7/iQKaRBeZ32SGn//N4Dqw1actYebhiPGK/0Oo8NuD
+9eY/4AzMEXzl2rHq51EBjkfSMWLStp0oZQwQBVh7qGTbOYhfr2ZF48jtpfAMauV
JO95mK+ah7bGuqwBPkVw1vuRiVLiAj/vKxHbdWBkd25VY9BqX6W5DHEMCLUBnIxB
BYjZXJNGJkEJzRhSuhNhbngNNDcv1zTUt89vdlkuXVra0CdIBZjesq1BB5wOIFx2
OHgiyuDI6qyD5OZIrWiN06THd0NwokHhneRGf8WbcCI+eBX1kECOI8cKiSdRNh2b
fUcljVe1f+9Bm86YLqzb+WRn7QrOV1m5Y3CzQ/gWRtRHkvHVBop0J8CLfUHsIKvN
gM4D7WAkuhaOd8EPZtJgn8oTRfJ+rLFoIVyUfhp6cuBdoHh9tdOntZq4F7rqLTbK
eZv9rPlcW8fcsmjA0PFjKF5cOS1BE4Y294Gjle6bNgaKkdpU4i2IzI9v8fJwOhm7
Q1VAQu5yneYZi+zI6ISjYOV23CgtVZpRykwcELArUu5ynstDMTSuKY7rClgCL7rE
QJlLL9kNTD47L96csJQHqQgtHxblK14H6KR+1MAjbYiRWr0UiC4nVYiuT+snhwJz
AQ70Mncl6rXww2e3F+AtRv3NNn6aovpHrD3jp/9sFCYwHzuANV1CTf5BNQla3Kk/
9ggNzlOwcBhkvM5by/0cGickpiK8gMjNS/s3synEorsLP0JX4gq7/d6HoRoB87Iv
LIaOefaN3Ubm4nxcZ/X7B46IxMoVwJU+77BuSTf/JHGrObFAh74l3w+GrzGOQt4O
kYQQ5nYjvW3AANr3h4b6Fl0g+6qi2HraibX9QP1U48bLsmqzUnWj5B2cU6wjULzo
N6dNWkhd9WfsFE4HY5EY7PnL0dTjeAnFW8fR6muzd5kMk77/mEUnJwMVtaMAW8kp
Prs0LndsxwMTGHhf0MnDQAZCdow2oqkm5jO2m7V7lKH7sWvMA8CkS5CWx95W0Ogl
Ndw4zIQDsiV0T25pTAHMTXpw+4x3yeAqEMTHXU0nd0DXZZMEPP1ShgFMpJYvUo3y
A5H1DQ5zHiqovywr28gD/aV7SBRfxq3RbrNHtl7+blKi3740p6MoTqqe6rCq8elz
BVCiUgJpqHMuQevUmmrxClENx/1papwCiJWXQDSD1vN3HxkxdA83uZrMcouOTkE2
wyPIhxTNx2b99ux9uCtPQdIPPiZNnoOcQD8hwlux9HOl16wXhuhxr0H+GMVF+5Rb
MdBgNydS5+oVct+ureKC4Y0R6goVN0se8SNqLK/8i5UtI3gYbkxSWCLfM+gQq+56
4X4oxXJsHdMSfPf6N/90EckpbkT74ZhkTubupMUd2HC4MhEG9qY9VkkxBAfHSdPK
rpLaUFdsm0k2EC7stYdkczvVBUDpZ4mWO090UTMKuZDyu1WW6Q78uRLHJVM1WDYa
3on5O0aoaeKrDywDkhZy/nOUiy3dysou/2HnpTs1OwAI/hPK81snltO6uWkTULmo
0E5lZaUvOMi1l2YSPznrtxj2cnawwl+Zj2IfRPBEoaH44VV1DIioyJHhO5L/CITH
MVh5ADe1iSWo2NU9GzsLFQ08vzvXMqbUb+JvCO6alpVib1H3y2aPqWktPsd/zaN/
h8DJSdAnAJSLzGx4UZXpB3WWUVqtsnB9ZbLKfaqApa0eVCnjpF1CUwlUSC8hl0YL
HTPBu8VfwHK4awFNRNuoO4YXaC8dZ8VWxqwFX/rgB5UZOkECF8LI2mXJlt2dvALk
OivvI3aEs0PTXvdwio+coUr8AQ4GBUraqE2XVmPf4kAOzhmWttmtmfs+qtMYy+xv
ytdKVrjLTkQK9fDWCgrnEarMYZdUWCw4MZHAqjpVKD1kKdE6c0jk/jfhe1Bn0WjT
gL8UUzk+19qPrWp9Glfi9fx3tX7mBmXUTsl7fojOmm75oEj1Rkq5Bhu9PepLZiJn
cP4rE+rIvSp4RQI/DTIW3RT0Z+DAYEm4kY3oLlZ18FNb3BRDiWN0Tr3lU50AXZsD
JUePLUuFpJdCMeQR12xvKIp6EaXPgzMeBwjNxo9Dtdo7CWLui+8ZA0iNp5RkJha0
1lpg+bKjC8uC5aBvyJyiZzcP+yUais0PepCgttoLg+wDZelUswHgcym0SJXKLGAu
x7vGHm4N9IYcDG4lqZa9MwTd/BFB6l86JP+hioqKNHIrodywJTKYGTGUbsSHK2hF
QJ5yBssffB7oNYW1MafdkdTduYjipnaWAOXcu3sKonP2PLUXsSOboM1/gpKZRRPh
7fqLKYm1l04yNKMARATzoRjZLg44w2tNqvMxfWJYsXEQrCf/MwvRwWurQ5bTMPgT
xOzOQaWgLgX19lFCtsbpTPqB+szOgUVrGMEpczVHNW/u2JynstnpAP4F4oBi+K0B
Q8iGFrNwoqnGJf4Ir3+Fm3H582wxyzWcKpKftJ1AOCwp1PAXPUP9jqEEv7Ls2blw
SZ/ayg+H6SxUAxr/PgEmLhe2nipf8zP9Y8zkxJmrm+J3tpN1/Ov+YcKKSx49cNX2
cxlbAwKBdjpeTbV+H3+kJv/9vu005MpEoYGiwZ9yn3R4h2yvhAOfPzSlamlQnOpx
3ZyrXo/ruCvPmsD92Pw7MC8vRK48MXu8k4odD7cm/eDmzCZSGDVDXCJgM22WU+41
wLtYOXlQ6N7zz+XrSSzUzu2fWAG3JDcJb4oYiSp3i4OXoDjC8M5lbSlPEm5vMc/v
mXbrjUwgtBeucaQt5XyFf+psiCV710UgI5HoUobe4mok65oQjwmRfxJ1YJcx4D1r
IaUcrdM9BvrrXLIR+gVmdSxsHtN9rCDjpiNxhqoltGsNebckR0HWt63dxhsQ9CC+
luaLzuTeSH7/eJOGGXpDYkOoM8PDcla7GuBCIoYWH8R7zsQBzZnToGpT4Sl1/2sz
gq3ExM9BXATd4ubsFA6FXrE9u371SfbkJyrBhw9GwItRQfGvZn0sH9hC1c11Pf21
Z2uXKM43zjr+EYq4l9sSpV6zXw6ZjLnkat0mmd+Efa2D1NZdwJTzOMRpdQmFw1ej
0Evw4k7LLWPtnAP2il3lrYbqMbBBozAGnGkO0f5oMiHg/V9W6zyJU5S8jarXtTXr
m+ejyYkyyszZdkyQLskbgqu87YQILmT8vdrcCMgmKx2P18BG9466bUUO4VXYt3dr
LIQx2zBxbeoX+kkOECvBI8l+0X6gYwBAfIy/pn9mfZE1Fdf/rrAw+U4jaC2+bEDi
4Byne2r1GecKBjCNiWJPn1azeAm+9V1MJNovvKEgavAZX76mItuh/OyeFKmvgDoN
8Qu8AcAbFh561WrRm5Ks+dRJQuBYJkm3xd0FZ6Q0woi95l7l4qR2dSvB+kLdBhAT
NRQXV7njcXzBZbTKO29qXFAH4YJJLVI3ZKCtysv03E9RVcDlEOwlJs5ZWaYGcnME
8NAoGxldOlqPlqy4kFd3FvO5MnYV217J96uq7tYjIlO3ts1W27cq1iFA18sE5Yaq
2TJ49+ONr3ITtqLjsVx2p4lK29CDbCFldjgwjAF/IqHE8wenL5zXJnJNexFuLiNE
fzQOyPrgakcrhkz3t4Xswaw3T4gDEA03TceR4KBiTgbSsEk98CvWeFiz21B+KD5u
nUPgaRdfqpsvvB8SWa8YCK51UQK+HVJYlHVaUkm6YJ2IfTQsJJGRaqEMZXlnQfol
PcwQeIEMUiEmaVHE5meeZRRPKg41Z98QXxDWqh+gEAEPO+zabvu4goHbqwOfyjvQ
aAE8zIbk2iJ2roOvbEA+ublspG15+5vOJtpbgzzZV0eA9WCvaVaOUlBAKILRTtsT
KDtZhagSPoVlqf3iVxzxlPgQpnrnG7t77oArPrQNVPO0OVgYAMynTx/UnOa1U4oC
wUtQFtvD6zingjylYe/ND9F4xS/Fht4vJhRY9WsJHrT7g69A20yyqt4qmehWEV7X
V3dv+3hI8TO8HphqmG1KhcnmJOOWQtEBx8aheqxr/23TRw6aqg6241sufnLTVai+
I8SvNcLqbXuRRnI1RZVNjzew2HIJaKLW4BqQYVnC5m8sM8xH8daWGbgbcW/R41Lt
noxueyscSqklphHRJHTJT4ajnE9SeSOEDos1oiGdSWWRNLUI2lw0MyeZI72nbe+Z
q4aLcygNR5nr2QqMRBR//TiDmyZBbD3eDPr+hHsrKhnL9D1SCkozFn0wnbXQzjbI
xUNGBh0pmQ9uCkwvUnxl38wjuqEVojjDaSiOMM2ojGaDzHaTeVjHRS4iRwkiLkz2
z1oaY6CyCFQrdC45ZdcCnWWTruwFFEuRMM+Qj5ql5BvW4Un7QAbM5zI62S4koPjg
qBWuhZQI3mwchCKQDHgUdu2/m4w1L5gA7/ugLPuptULFy+6DlFsOCVSTcpkBQZt2
uRFr0wAh7ikn+bCo7SLK+gO/UosY3taCxWt++P6wqDenxyCvysNtOPnhYkKct1gK
0q1siGiZoKoRrl7CDbqfE5+F29CfELHkV9GuX4ciwK7MiF0m2xW7Z61ydKXBV0k+
2r1dP677wSZdwGhQ4o0psbEYheEXvDIcEuTxdSeAMCDerllQOSby7toNr2cTAUKo
5bLOougspz/q4U5pCJY9Li9mHbeALqUILAdkktOKJTT/falth9TPQfMKqzHMQbDG
38qbDiPv6FLco8AMlHTUqTNfDPr9lmUTBHc6g+L07Wvh2H5a5zBjwRx3QexDI6jg
YY4vtgF2JfKhvSOXyHGZQLcO5e0AsBgaZoDGHXlK4TNX63cPOT2DKX4JFlB5uxJ+
vGC1BgECTJNEDLz72yl9LEXbPlzPPBLmvdEZKqobNixPa9nU+eqEPjaMXhJgJx8O
xx1RMpJozyYfAtDq0fnMmu42WrFZpdqRfGbBotb4nsS4Xktw6svxC+j7Z3NX11Bs
rp+RtNKLvaUjVC2xaMWhV1nHnpEBI7BerzYbQ9xQD3Cy2dtD8wcVTnsBTvQI6n+9
JiPopfqLjmcrANxAGSMl+LTKNIPcQmEPC3/TXNivfoAnWfb/0FILfApGsvqiBjto
V4qoOVpwqMG6D80a5tfBbNKD/IycAKB3SJ24PacmHWEvBysFlNUbmHEtSr1mIZ+2
Xi282RHDDCxskbUY+iQLquzB9p8xY2C6CEel3tzshrxLiivePm7NNdeEhXPLEyJu
GN+T8wp9XMAjET6xS/5o7X8oQ5GOrZBLSnLIRD9S74vvXxEj466CUMCkAPSqlBuT
9pxjF85u98vhNB0K6vK1R0+nMk9yg7wPRC/KNkgwASyszDhHOUUSw/xSVHPr77R6
JzaRGDtq2btn1aLmYJX2toK8FonafNeJHkA3qKWY+D95WHt3ZVV4ElAmrWNOXrcA
8dG0pdEG7E+RWzCIBQiYgo/lc5aQ3kK14MBkoa116SxGgKgbT3dImKHB3S5r8/N4
FiddOjvmxV74XZxRfT7qWItaaUlVJp4JH65zk+gV8Oh4myHWqmrr+2gf4O8g8k91
R2TFUIs26CBehGekZJQUukglxI1niUo3BP97zEXQucK1HPfncBQ+TjqeS8CdYkZz
2gL83oU/DWc3fg5b8KYTSttLxs3WM8VeATP0kZui8Z8iwuIcuBW6BDxTZPFVsw9a
qMdpmxXGZ6l5wVsHdgfmb0EoLiD1YCUCv3IvMUOVwr20PFwhsKUtSRQW/bGXZgql
b1izUwsHOG/OBz9KYIdd4VQG+VqGN1lJpN8N2Ot/s+qh6cDTKO14unFJSmLVCPr2
DOZcdn7ltv/pW7Nq7cVnux6cuP7TvxexqQXZKjaX80/XWs4XouD9JCpG6YOX5K0V
G/Co+9OQ6H3kfHqmq1P2tkZsBegXzvk0szh0JPmgbF/DFVqoUajvSC0ZGNvIckcl
U/q2NCB5g5ncHaBTAeBILn/PkVFxZnpS90wB/z9VOi5nHe0thSNoX5kD1faCK5FQ
9kujTlGFIMz9LwL2ca/C4/wVydK1RYc6R9/2Dm41lXxk3NbqCYfWkaqSfLUzc4OM
sSMjUQfP8qUDh/QKN0rTDsAZik+9RXj7L5WLeNINaTT8WXcVFxyvkjrjsfnDWVZt
Mp2bwG5OlLczPt/hB4G1TLGd9+kHXFmoBBh7XdTJS+1Tjx4mkHkPw1ZZOK6aKlj1
Oy6soXAAA/y0DIutXr8Bpm+kg96TJtNlwcPa+k86g+GddguQg38NKE0nmSBviavO
VI0R4uZor3ri2PmxHl+popzih1SxespqFdL6IL/bvU0Lo6mH7IQu5olqj4VIslG0
cmCiiiQS8Sd4qGLwi1RUl79wLJJJmLpU3i3vwEG4+WMQq1sw8IyA0D7piyzz0Exo
zFI60u++hkY+e7YZRdauC9a8b/lb26uJYXv+Sl+2EREoEA5ftPPEgyC+b2FlSmA0
Cj5l3ou+rG2J0IkACMOc1TG8l/1AhHFPn11F4c6iDRWVygMr9F1kO77OeW6PLJ1d
BKT0ZPig70fyDtlGbTS87b/xiJa+OhWRgcKYiRy9kWNZ8h3yCEzCEk5jySmhbehn
pXoy+Jh0OQcOOh8VrWS3m1SzysmHF6DKRMRhH/u1YNNwkU7T8DJ9lhb0y5zr1dDq
crbhu4Cb7VezVWmmVSDcYLD4Gb1zVkEQitYSrIVdA2o9Xc5Ao/6v3IKWovr1RAGm
9LJNYleuGIs/fa1RNfloQAAWUxDVgmbl7U57+Oe0DlcH1IhzwsJ7CyUU3rw1lhP5
M00a4HNuioFYY0b9DoZN5TxBcfw14IFdKM2AASax5F2QRX+03igeNVGRWKEhl2In
b/YjZ+XPvWfZIJZvO6d2JGnbYn3f29lTeBMl5PmqHgCkoxWZoevZza1fdc9Q7ED2
VY544QEB4k8FxU59PtL1nlwa0GAkDkim6EPa7+chQI8RqLSy5BuCtryX4LnY35Lh
ywQ9jf75zZyQ4WWs8kpDShkQurZFzp87TmVrpxQeQx4v3u6/j+wsSb3mf8qLW06W
tFny6m+RfVk+549Va4WPB7HiIRkzY5NrgxxIkMDb/eNfMWrUz0HYTZykVxp46bL0
j2izNRVBG+OKrTsbtGtkruhRB2SrWy89HM+qlXWn/bVuk3AarVgJk1W0GBX4mLco
lud8zhXV+NdCXT8ldUeoGMQMKyoL6xhDtvShVDpC8XQq4rWuQDh4XX48K92Y1orN
9AjUtmrGdJJCM2DivicG9YHI/vPIUgxnRv+SZuqBXIoARYlCdATR4N7mUZmwSOM6
YpyqbDIXum3aewEdEh2FaMtbJPHcjkE9TXbnD1E37lEAqvUlr6WRB6QgR2Ho0LXO
X9XCMRlVxcKf+OiFBX0WJ7EKqFJnq99RI6DWVrs/MabfhphfGV+wvrLCv/SMBX6O
0Et+srOkWagor3Jmd6ILtkPPWRQ/TmY2pZWATax/PKScbcgdcacTHWEJZh0gy8hv
RuR0hA7VtHI0ze4qoUx25egoN6bnwg118Xagpq7xKyGBtwcCY1o0szCumeFEm18B
dKxp2hGev/4Vi0MlYjkAqll4yxoUmFi91MfC/CIPKKb8Tsy+ZM4KjbtPhhaNyQz/
itq8lTR5hv6ZtoGpoH5rsZS16Tjkk9OK/fw027fR3/utoF4Tw4m6C9D3oACvXjDV
2JOJEfD6OYDEv9YGrcwu5Lpai8Z0hfDC3BDcEapmJSfw2L/c5E0S/6OroPlM7+fm
NAgT8oyCYgjyC1EJfUST5FlFRFo8TNsF5QENdjZJ/maqarBacRhXDnMuw5NVLdlg
BCq4sn/zwTU7MWj89OmqDKHwWOYN2lzBwtsTQngy0DF5/THayQBZmmECnwNYDpNt
oJUPsQl+j2OKzpvB2RFGcSPcSU4ll0p1G8R7Dd96cQts92InvseAT2YnFm+cwOQQ
nmG/pquvAGL72FJgAIW3/esSDIm2SDZ0EIWUE5uVhUdzjju37ornzJzbpqKjfEcn
lGsAmMM8YqS9RcfBOLxnGDnZSxsFXHN0fRNmE7BsYGv/gVV31H0tpxN0Pr5qocUC
PPUG3558ZKX3H6Kv/65FXz8ajc6lVC0X8N2y+tQDhFYpazpL4K0RzjxFrJt+sSWq
8U+w/vndy8ABHebl1Ktsz0w6ISQ5tzl8JWJlitvLJneR9jb5FxPfBXIDNPLu/tYy
8J22GYWtVLwBawAdIJVW5XweXTHyZ6x3tE3r8cM37RBy2lK11Z9SbXVJH3h1v7D5
s/n04HscofO8Oqa/6WXxK0eDCkth7+0OaIgwjtkmFWpkTroMCM12QBIRC2em6C9G
KBgQgTAkCXY7KLHv6h8Sx3bNJ8qTKI/KCm2Q4p14rMv6zhybhYOyH0Do8osZKiI+
0LQASEk7so5gGs2mng3Zhit80w7j8IgPb973DkqEDKHTRLOYFXLJcVYz2xoaOUCa
+7koRirELltCTGkz0+59yu80stecyyH5Hb8ktURCTpwH6yWZm79dndrEFVJZ1aI9
Eeneezz9G+IUy5b8gDSDJo5lrZRJBEL+0t2/4SOITtk0n7zwypcKfmSl2fB8ovZX
pm7sKruy0yEsoyUp2B7MdpeM1fvqT2gUezZMho0EK+QwnNLJfEEoGm2KCkly9RWJ
Tu5eCf2Bqnjxd9lWLWRz/aXG3AASXOqGEdWeWQ7QCI0L7klD8hGgjt6v8JmgH/+M
w0CiBIllPTot6k89/uKLiYqodwfurYq2i8JdcS8nPh4DvPsMSPQajW7HoXb1ygq4
QXY6kcyEgro5YUY238VAm1IAcISH7Isp0GHr/9041i60snv29JeSERh3j3Idzk5j
mOOuJuEbKz35WTzL92od9AuXck4xiTYHbiKJFyB46zIDUMk3pVwefxf7q+EfkKj8
75SiqsaalAWvNEWYHchBEw2WlKhCSbAXC7D1S2Cnr3YZ3CTF5BWlx8jISZ9YBnY4
de4/C4DUMy4YL2hDEorxjw1S/Wzwt9L2H06s5hdjCSw01pPl+oElHh4mVRL4GEwW
EZSH3coLVtRG07hWYJx8bSjpB9QS1Rvicykjaob90CE8s8mw8vN2KpwNNfJaLmiH
Lxu/OMw5jag+eNBPn/2OzPLi0Gyw5CkUm75j0oXJi04IQhz58l/sv2mDs2dNMllB
+hkFCH3LkFuXdbbdQYDY5lz6cnbu5EJ9/sUCGoeP1H7XsMsmxBH3xDlihp+O+/kX
4wu2HwsuxRe+2c5PusVWkNQHPd5kGAwGhZ8Lp9NQE49GJRNVs7ahLZ2FrjOFpmmG
p8CAviiaD6+PnYM9ei0Rt6IraJQdFEQcsoHZTWQMHowcUIM/m+KwfEVd/T+Qw52/
AB8kpZoZhYuSpEkqlyY1SFnj1BU49u/PIlfdcNI/MYuyLB+jytG+rpv0yklVpn8M
6vlRrj1DqDgedKea+Q5O2NUfY8VJdn7sLHdo9BCNE8RQgSTZGhc4bLOQ81Byum/z
NvepYjjnCKLU/SISJ/UG+XQUS/gViFNI20nfo4PypnO5X2wfGu5FgupEfgwciENM
a9yO6kNE+LByGHk/FZaT8bXyGF5/lYILzVLQjGLISdLXobd875BXTHif+/wR9/Hk
xodIV/KNtKd0taXRxfNYgJbhvFTPmNKmnNezlHw17UIOllD2HTUENdQL+D4NjKkb
3dZ6P8HAk1ZmSFnSRsqK3rofZhDw2LhMm7eYuJCcJjjDE/r49OmfM40pVuQ9NlXC
ebDNj29/73fN+vIwF+Hem58bwgZb3ZGJD3yxW3WGNR50sNASzb9k8qnmHYcUgJ3M
HkkDzWTOxNAPWH8NtniyPlbiPg5hqOoWPIM9FehapcD3nLwgS9KGVDbPNlBSLX6n
cRNLvwPyVVp9ltv88GUSp/5IHIhL2B6G+YU9ST9PaahHKnHy1uBqGbH7DgGxMrNI
smfG27a6VsB5AwPKB0Db5tH70+gVr/HUDASx1iz0w3BAq+wkTh+caITB/LMyLehJ
cYDXAvPPtdz5zAFe8Lcwc0lWDMdaMNBSbotPX5d4y5ipYa4AJB5Vumn1bhUhzBDr
18pv41a0swBcDzFsFyKTlJFb6liycFDxDp6uHyG3FsJ8I/SWyuM6uhibpblekP7/
une9nIP5iRtY2hdxKv9YzCWdNcnnYJKh/heYq+i25yvfNSHuJxNp7Bmh1Kcx8wMX
AemKdzRHVxF9bBfwifwPedvqW8clg345SIoTgfaQv1mLRgIe1hlFeRlQZoVRl9lr
0ja71CBHvPC98mNpBv8+0QrX6I3OhTGqoSaNjIxZJ8BwIKrJQ/DJj8n/KuN+9WnK
J5eik0OYhXco0negYM4oJzdq1C/OxqouyubLgxaEKvzekHkXDXkenissk3eiyz6x
5zlrnhx3xSc5Bv8yyg3d8step/24GBMAlsdGTBEJHFqp3x40TnUwMJpRfRJcMB/j
0ToXK3KFzglJjhWL2aPlUiobUJXYjA/0DmtQiR0hOjoCnAXl6WE6J/Hjat5wF4+M
hAaeVKGDy/xJir3jkE6RsH3iAmEosxibcMwLr37zfPph6oB3j0iikVOU7R/XuLwk
nxgfk239sEmdwDY/gWPOrv6GuSDwaujpM2hdXBw+KPpZMwtWmg05dF7S8OxVAA7K
iU3pfIiqOinFODtidqYR+b9Nfj3wjfmLVbJFaL13WUxgJD3N8yJjbsEIxJqtx85j
cGLTWqTSTnmhEJW6UMmjkjDwTBH3FmNVvKyrkBZ/5qNzrkhdKLCxlgwkAUktc0QX
1HoL/d/s1DovljouMAXgQq3+Lp/b6nr1mSL5WEhXmjdgj1rVRMqt4HEj1f9rkK76
WVcan+oudwB3sll1ZoPkZfTAUQekE5Wdo5Ixolwr5SKcMuOrX1FMHPbI6Cv2UPW3
JKx+0NP1zw95rLoITt9uyHXNXRWm7lXKw4Ia/7+aIdJm6U8TSl3dY2m7ZlX/g6sR
zQ+3JzpDDuHvFsu40GOoQMzJzP/lwlONCpMQCnzQ4eraRSmS2M12EJZZ4grfbApm
vfmCQoyTpDpTKm+sEPo3fxTLB1C91J7YVnGv4ADq5HYPwLYUnKdo8HXrRu5QZCOJ
oKTWnrGVbdQyaLys2OnifRzRanY1Q10ouerP4rQGZxRnbtuPd5rBj5Vf+R6GE9aB
kKIOkxslrxEZUB303JiZWgL8GjRiuFF9qNHPQKhEAtup3ICJc8EPq30aae5cLMRS
vOL8I8lCgqlLOm/19BTRbO/AzJmsTyGSb87hkqU0JUqQohb3bmtrGhDiY2M/f/+B
7H0YMdkOz03ArJOMA+CD+E+31J9HIxWTMcmY5FDXVsjRmnBBqXeAICAtInrD2XBr
4Jn9mOYLppkMQX1yAeyhZqI52Z+7S11VKm9F3eYRO3p4jOxk8PlJcl6d+19/DqXw
ijFUZQMSuZHb90kB7e4vOGzdgbemhiWS4xgTTOA9uNbx/vhxIy6iwXhWFLuXbcD9
pbsbRHgNLxzzrV9JC3fXv5WP3EE6c/1ZcEYYzKb/HVdv35elvJ8ypHkEqUfIPb+x
tLIj6wILcgIGHFT4gyC8BpLkSEcNmbR3jr7AWZpb1F5vj9iTwqBVVPetG4jAQsNK
vureLOV39Zs+UuW55YUUMOdBkFNHqhmNouxa2hEZs73W1euRJjFM8kd5PdkJd/cd
VjhJ6HA37I5tHFqlTNdpMDtPSt1Phqzu3gAXZ0JCGhO9RNGtars9nZaMqv/CZ9/K
x6KZCLW+e+e8w6G0aN0rop/WUDIP/7V+W/8NpcY7udUA9QJ/JVAZwoCM4vh634J9
UcFsttUFDtVv/SP1wLbgDRo9A5R0Wrwbi8t46ymYQOc0++yieIIhYIY3HMS/DjW4
4QaX6fGTkRl15PTx2iZsF4tkwbNPoBw+2O1HdqwT6fszhov7syyHg7B267IUqLAt
xv4l8AajjHhCnlWX1PqXRvbbQKU+QbixCZlMFZyjevHxjmjA33DRcJLYMNhX1+fe
8wQs3gMNS4dWfqUgW/zE+8BAdjf4UVdVAkGjLshCP0hCodMbA53/ylL4BLDGt46i
nxp8ODwA/Khy3bdoXbqP3teXMTAWlQTwOHd5SISrwkU15eySFC/BtelT+ojHtkgE
cra004jV0F88zrqHXM3XHoN2API/fP++zqTmLkrSBsgQEyIRTIiScH2MWRMOXJdf
y8Ij+kruLrGiq1qcgucuV9XhL0xBHKolYDPr9OQmkm4a7WhV9EEuUvLWG9HrzDgZ
1EIvSHBcuqN4qkz1WgAfQE/x85sfcET9yfr8NqvtzJqPuNedtMbH8CWE4n8z5Vz5
K3MkHMaWrT9PV+3V1rxy/nf72NZIQddtZLAtqGzCiRepfxbvYDUy5Wew+GA7y1KH
sBwI3wyBNzazYEpgCqrdy3/54AhLGT8IGhhgoAb4MUz3RASQBsz9qsJ+nNVVOCTR
6dRsswtLEjZGRPuO95LkAFbG+U3QQzFaT32Gs0v6+8SKRT5i5tuIZOg9KivpwIHN
aLbcWBPWEulY29BG1pVQByIS+2UD1XG5rlXy1wfGexIDO09KMUNK90E8ZA/JbOdE
2Jr1z7pVGWOR0Zi/qLmktPCJLg9YXpSGx/3os/HBy5jhgNFue9vmTkHWsxQC3788
6eeLdKxEk7rZadtU/kNg0Dk+fRvNj9KhFgtM6gqg8Pke38tSeHqzomd4wEGr5h31
8Ekln+pGPv46UTEWvSt46Nvkfb4Qyb66T6TYnTogbSGkBMDgUv2gmgLHmQ/OKr7M
Umi4/SUMec9cJAVd/N6D4CHTkQnQ18ujC1JrmkOED9MQf9QlPHKDwBXMPTin/nIH
rvz21LO4SRV0SlIMA3rAVaSbcuNOyxdcuVm8EVZcQUM/XIOCaCVCZSyxp9j4+ShY
asYeXzBsG5Po5HhmRTNKFIJdoQN4j2kXVDn1OuYpBm2SradPBaStIfvVOOIdvtVu
c7RtY+p867yCmXO1/vWKuMB/aCFEizQwLJDSOmRciHDuhSuCxk9apKPKP318VJEJ
wfzYMoZnAAOgaoPPePwap6SHIhIlAu0d5RR8T30lRmuTKgtCjZg9+N8tfOTFxf33
G0+8eF3OBEBi2WLQNwS4WgIkRTGmxkR7LWD5bRwr0xih6Bp/Gigl8GFECmN8jxtE
xxAbe9+GoZs7f23wKqouk/UZEctmR8P3Wnve9LbJA+9igDEst7fdQSzvKnR+bTSO
250xoRDGHArU5aqkllW5qr/LhWC5jV+oa6/z0hSklUsCA8VObDjCs8jDQN8j07jJ
Jlev/clupE9EMhhFc3EYcXkLsrsN6m3SkLcS9DjVITAZjKMb+I76uHkhzMMGt3Oo
dsSJWVuHi9YbV/SUx6tfG07FS+xpni9OhQ8ihCN4jKUh1Zb5EEZd9az19gomUaNF
Sey4a96ZaSm1jLm+N6Uy2UTv2HSdOeOLpxnMZnFxn6aoCIXsAziavxxo/MeKHMah
i4ezkdhf4AxXTIRl9B/ixnpBKAR5aof9nGKH/ddBXVwfSTlpJlbtsEhIqaof9mfp
L1KEKHaL5UCVOt9QPOyrleI6kE+4Bw5y2PrXLVjrbL3XtF8d9Gbslt9xBzUnmIBe
PNy0nnCN7Ep4aep4jC8x0+ycLwl0pMdtn1eMHknDXlonWRuxCAP7qQk+ZsmHIZm/
/jZm1IOztXrohvlc/wHnrenp7KwCnrR8q7XvPuN0rced4BCSr/8xkOlUs0DdVYE0
yKKyRq0FQ/ZQCYJHqs1+gATnLqbMyRFYaOCbzKreLjHiCQW26M9X8e0zWJsfaaSl
xGh0G6PlDsuXY9j+awkPfv7hLdKn2tPPKJ5tywAp/sFUXCtZ5bfS5+uauOTqfhLv
rnirQgMjAJRZ0Suk4SPcq6LExuqViqg4dycMljNi+6nVzeYIa0mG0Z9zCP+dbaPK
RE83xFrrKjP/Y1tLPHuLZp+hw/OJNcOWBu0wUM2wEcQw8PQNpQAScIR6fQu1YrF9
dRPC28NeypRRGeACcCDEX2pYmLlxpaYQmMLDmNqMKR/EmG3z0v4KcogHEklQAz3r
9l5E80falRNvKOhAv0wmgMaZOb+7Qiv0MEz62RLhBLsakLNxHW1SSauy8hIBAKV6
E2bYldgTjW501fAXLk+4Tmq4zyLii6qRPQGr423vs037Ll/VDjYNQdlB4GBJda8E
2O5z98p0IEYNpQtNLCnRFAJDpZHgr2f2a8NnLqTxdDGw2MEhHPcQLDPFhPM/xx2/
OFTr7tUk9JlCrnc84UVcTZnRnax3gov0HIDZkIM4YifOiIqQrWKM/XK7D4N48Cj/
0FXLL5vYCWHsuYls6d6ZyH0dIyJy5wh9zY/r3IqwWMk5x5xcCY/A2Xs7C11ncXky
LfTvUbfic9kmy25gTWeiEXughiAFtphwdxC1dX7JTEfJlexa4VF5HD0EciTpBjJA
9RmqXbrdX38DFy/BaNZAK2gymkVQCW8itpw2uTq7/LNjRJIfwlfhqZcDnv4uSKyx
EYnHJpC1/V19WioR05kH/h1IG+kIJwFNnq3s5UJfkrX8j2DPsTCMsg4yDvmOLwfz
MKg8qqjMS9ZWQWM1ln3RB6sEhaEA0RpMMqn3l9osQWb0qNVvhCOHjQ1816hzfA3a
yMNpPB7UEJNMzMUV+MoAJxhMQvxriw3ESwY8ZjmnBZCA78SDsUeN9naCKU96xM/i
j0Z6ddq0JUOdZ6xTke5y4y7BoR6XoVJJ2aCQOCevglBHT3u/+AKtGULgK93McZ/f
fIKqktZpGelsCor0xa2vYi4jxGlna9yAQCvjAAB/rRdj2p6luJ/5UiEMNVqazBXZ
99kSmfl7qte+vYORUm7XKyYVhWWk95iseJz5I+zrWp6vu1NUVFCT8FyXQT3nG8gh
Mr7d1pkDRRbOTIwbskpb0tY7lX+zT+UPPLlWQSuQG1QIDRADIUSPYVibiadkGIca
EIcm0ClW1MhGmbrmuqBJtZTus8TzEM7YEGd0az27j2DWeNtUt3La8hWgVcmx/H8f
MLZ3tsntPtyYuvYRb82GKYR18ztb3II3lYW0TqDMSYtQD7mKmDPOMCiBFiXM63xD
/zJqP5Yb4fIIEWPnDRX7US7PkDVW+mw3h2WBHkPXwoTtlaqHxsJmD3yPDy4jJTpx
Obl+brJ+UbfPttsLpYQBRzJIjtbjIt1E4E1j96nVf5wmfLL14wvQRsXYMrjcSN1j
X+x5XPj5LX7CtaTZZ9fR7SAhrjPzLdcrxLKYmCkjCnFn/1turkdLsZoRpVhSxwr7
19urynpprXAPEdwJx6LMCxCTrBtuYZWR8aH9qCicNItbCuJaULZbJc7d8T24JArX
B0VdNq3ujIYgt87Sq7wkXv7rhHnZipxJzTH0I+m421UTb+PkjXcYApn+LT1vTp10
UlLCRIZQ0KNItJ/F6b83Y89s3p1Khwaq32ppbmTmh2PlnXZ0rTbvCheojcIkdJg8
ed4MNLfaFJTOjm7Y2vYr7zV0h4W0W1PCFdlJ4viq8EcwlbWLzK+c06ZsOtTfq3q2
RhvfoQv9KzSYwGvsxi72EcXp3QfnkbwyIm659PCwLbCXTLyrJT4pKE5UNBy9uXnG
6L608SJL5T4fLssbk/V2U56uoKeOlFmEPzkjeUnytGIG+/+qlKtyA8hz21lWPB3Z
K9P5NEq619AiYWeL7r5djVxb58xZ1D12OdnXKBbRaZwt3+ogzF5e8BgzWeCsgNTE
nIOgH0qcIL3163qUcPVu78Mvj5HRDrRAFU0sQXgg4PYSd6ksT2qmdcSPDutSWZNL
7AhPHMbwsXkFJBhmVTH1pIny8dy1leLZtuGrqi1axUamhLVZ4Ra2uYhP6V4b9ZL1
Iv2Bh6EUTPm8Wyf3lh0V3Bo8tiK+EtTmKpxtfudihr4kfPiPZxytHHaa2Pvcw+JG
5yUV1vCTM3EUTUdra9ngPJdYCWF2lDC0g0zjsHpZ+AaZSh26zQ6Y7MF09dFsVo4t
9BvcPmQxAi5uDO1Lr/1iOC0bBM2B4DSMGsZafbi1sOmmf+vId70/l1sHhIRAnC/h
bLG39QwfajVLW/mDgwnnYB+apfIYDTrtR6SVHzqEMJaV7iXILTaWrhCepAK34OFZ
WeFaILNkGtjBkO5Xxdqrn7C4qqLFcltoMJcye6h6kniLWyc1LiBVq88XopRwM9rE
LUkHPkxMGUJKDzre8vbkWVy0i1e8qib02gseXuEe8gZPih2vAyTiwhAWWP8RVGXJ
LvFp8wNzF+oKoYyQx3BfkZ3ZcvdnwOvQ+dK5j/iGfaDk4p/GmkQLlnlm8a0Wt0I/
cKlnl/CDyCUfR1dshHaqBXJPEpmIKeN2FaS+R6gA4mbVyEMkqyuIfgzP+mdg6meL
/fcCsI04JUQ6D8cflwTAdx/UP3winBozSJ1GukHS/ihVIikV5W+0k5WlpncG6iRR
o1dG8C3VErtmdfKRTOFlSAKL+gYYZqel1kKskdSVEAMD5KCUo937zxCLNjBrc/B8
x9OvYRw05K1DR4iSA/emw6Juig+u3L6BhVBUMv+XBrLOIUbQ1PmrODVGUPHTmfBJ
DAGkAGmRHzHyS/o6lPbIIOt+CSKavvJc58C3Q3blTLpOJyRKYvPUm8HkBpciiat1
5QgOBor2MLw9w/5xEw2jhkYnMAqr+csNwgSjvkTLXmOgIPDBscGYvDxLCtYX39mj
Uqj1gfJkAPwUjWs5A7pZjTzkhNc9Q7YHLlcIMNC6ODfcgcdaybXhXaTUTR3MZxQx
lZF4UwMZckIDXLxU8QDBdqhmUBCFZ+1rp7VaDLVNIbyOiOitmqciPXGW49L0vFTt
Lg+rOSmsoQm/zhR2oQRyffq6v2PFHl5UOWH/v3nWRcey4KOgKwZNenClOudQQSUG
UPomuEu3RC3lFh6sKBuC0CMf/Gi6nT+kNoJwGhOcr2Xb/IHbcMbTrcSyhg3Awez/
PhWRg7tRjDgw0ziV34NPz6km/W9SVLDblDPQ7vAGPeM7SqXMV6XCcPm5BW0k5siN
VGyYQDT5MNb934Cg6MTaVXqHzsUqY3Hxl9yzxqDIzMglAB9zJpvhTQEQBbRqmxpK
8Wo0+4EXKvaUmj1qsPOa76xpspi3s2KaAPhsVKDfknnMQpKtCp0fIcUex1wB0RwG
CmZRDyujo9w160rRXlg4JGCfxFUa73zT6G3utdHN91DtBovECUNPVAwvFiCGR0SL
kzk0mVRuFGVnp8q4q4Ae60nJsouExl/Poz3jG7m53GITuAz0fD4JVIcI6J6ATCcd
KDAuRo3jyQwciis3O95rZkGhOSyCC1S0Pnf+sanM9iKpCE/JklDceKXg43QddKQe
EM6sf0yc7cPYND9NsaIBfSAmsAY520afdYVyltjmHt3pvYasoSbGc/Sd6KTnMgRv
sf6WzmEEOC6Tf8Kxp+nlrDOpL+9nT2ZPmvx1UXK3lykouICMbtXCDEGI3N0MEpCL
P42Ci+zJRIBbaEkTi1cNkKhgm+cyWd8ZN0JmxmVkEaq/FAdk2mDzYLuGwJ9xdC3h
oRf1NelorGSSiXY05h5tYiPilRqMOe5GJVEFwWBF9eEOKz4pGlL5xUSkcfeYHkzH
UUknJ04fV/psQlgZIE+z8Yik4PYaNLWb5wM4U5CCdET2zvAe13a98KvVTtb2ilZK
Wcjj7kVp4tvh7nMtN3seclEnl6yxZZFmtc+qb2Pj74HWzqPEcbRHte1BNRVrHIJd
b4jDI8mY1SyON4tlLVtTfj5zBXAUExQsPpyUsuZKnOxDJVco3pvIUTLSakg7vV9X
Cpya885K6DTiDNyNadWIIAWhS/IZaGMjKFmYI57TdWEK8HiISp9AMjnBuMheJwqm
oNNbhnP9xEMZrnA4FCVtz0HJbiIdnA4y9Poo5unZVYFPcj56S8ZFnWe7BqalLE8M
Sfslx5TBoyXaCQylu/1R6hKSTkl4NDq4qTgO/qwIhV/px2Wfwa+s+hzMoWWwYANM
w9197dDMf3WIpvyiuVghmPHKD4GtuqUPbODPgCk6T2sHzgQzNP+283T4qGN3/o+e
HL47E9tW4eeUQPfDQHShp4OAzYsE/vClk9MtEKQmvmAu6jUUjVZ2zq6rKk2+GPvH
+dw4J3y/myFB4zA0qWFLE1VbI7IHIKF4hfuQwM00pMIC6EJX9qALOLgqUk1QhKfu
b7Afz6X2oR9QTn+IsPrtAmqUPBbK5pOswoW30/VzdlM+y2hukmOrTnx9AHPjKnw/
g+VDCwTZMS7LeloMPP6x+wacrLFgDe+b+N0mpc6hWf5+IQZKJbjKdhDnTESGX5na
8S4qZXzw8qGgGgMumRETTsdwZpGH1LhZ/HZdOw+XEsGGVkXpKu2wC0pwKZATyY9B
MlCzbl2o/+o/0slVs1VhSGFgoJJROQWCjMaQ5v9OIsKeJvQlq6k4XzlCTH57H6BT
BAeM9bRbAo99GoSphyoeoj6CmE6x2ND7PWqNTUktV76eP4bR5+LhZhDSTNUfry9X
JY5WLaMXF8ZIYMuQHYw8ha3v01bNxke4sqiQkYgQgm/9PJjPOIcxOwfN084K+CG3
Tg40v0Vy3Sd6fH0KLCAzQ1FpI0tu4B4O00DcXxGzHJy3o12dDDM3mqGklnKdcoT5
5rEj/3F+CosZSb8JJZmVjYJmiW1wBbcY7kZVkbWdJPiQ+aEbgVsk1kJD8A/pvdsG
gzp7FzCcvXQycV9tTkYIFLIWT086HBOQMOOIPJDzRJ26hbWzpsnVqVq4Y+L3oMy5
CgWHwzupTLzzVH1tp5hufp6YtKjUlA4txS8glpiNoNlUOOeb+ph/wTowhV45+Anm
XTK3viiNjBxdmKT8nk4uEnIhl/wDPSro9DkB8o/rDSF4HVXjz9nj5q49V2yBxTxL
eIrA4QT6EqTmbSb/tlEKOWno3xHPGeiStmsdGdgnLXg2GH92fq433gE/NL6tTmjJ
2+l49TrOaKZij37XYrJGF/wxwX2DAL9G1Ergc95JAhrHPNa2goO2fJ2oCv3eIol1
H64kYVfgGno3ltOS19b1FWIe0+9o3G94QUk4lEDjSjyi+Pn3b5Q8g/D3AT/WZmPl
+pUXD1ZLVw1nUCSBkvHOvfdqfP6UpA/90fRymnK+S3u2gdWjFFlFcxUtrq60BR0x
AScSsBizMHoiybPBXrQnua/5ZLF1TA+9qut6V0Gc+pmVifVWjCQWuRRDheoE6ari
9AsQ9RDexyRaVZwP988jIXNi/5y8isaHBVF0H/jmkiYPWfdloIrMsUuoqai/VbAl
ao04T5/c8O3BITic8Wc3rqWSDPKPcp11LjDCCbVwsPidOCiDyKen7+emOtRw8ekm
crUM9oKuq85rm4aD7fGhl1NAzKhP+TgvinIVHBu0sfAIB5HdeHGrK3Mnxuf/AsGM
0YGVrfKbMcg8S8uzBSyfroecQNBirXeBR3+L/sr48j8hzX5nltIaTeoCXNF7u6Wl
CeX1ip9Mnw4hmdeH7CoOPtgwKDkuzLXT7NBuCCm5AtMuUpvmAKXKWA7TDJ8PhNH4
Vf2nAR99mJsHp6edqrYrj1Ck0PXfHWFRZF3+8/cmPjt7/69sdGMVDWgLs9qnd2Jb
pOGKORzt19ayBdNnYpk5paC7++sOOLsGsToVQkZVwBS8UD7F/yQlFtAtGEMwy7X+
RNXHEsTumKFRkPRXPr9CYFL2FmRd7hubyIKm0uD5pnyCOmkcVgGpjQ8M0SP08r2h
ODh9NsKk/J4d8a50I+DH+EiiA+3LVV0gsq1WdPGWVEuBLrB6v60Y+UMUU4eO13Bq
HkzWBzNqx29WbPq4I2M5s+oHYlAZmiKNQYLUPUGEjSK8zQdIOunHCuB8JjBEb9+q
F3Ll96KMA1ovejqRQLyBf5+W/iGDI0RyrSFK6cTg7sO6DfJ6Hkx1SIHuIKsTP8FB
f7T73xCMkCcxyo7PUw809lSJgPLBx97kCMKzfFAwyGeTrk0Icg//VLDoAo78849U
hzegMn2P/iWN/f8ULRrxFY/F4LAkBUNB+49emUFJvDAs4D+OB+hJt9k01tw/l09U
ilnV+Dk7VjiRksujs+hRoPE/4e1QLJ481nMk/bAl3oPUljVwcqq3N5Ykuj8d2OPO
HbsHeqnrJA8T0e7nid2AC6jeRklU+RchvrbYv7q4juD+dUYtG2TmVo5QG+QD55Tt
Nascwhk/4bgzBXxwN5JexBO+f5me2tMn2psX78HVqZNkCbNXfOy52pXUtiubBnGZ
dU7hqSlpFU5Jty7Ox+f2zOFONlAJnnF2KtMzoBqDaL7wM7u/KavMhuXFbACXjWMt
UvGIMatBlrm4VK01l2KsV6xTA5WkJ4m4KtSqh7IlJW9HyS+d9s56gaVw51lbZwM5
eebLUGLhtMXDG6Dy7Uu8eKMkBoBvQ3b25bEamWK/kiAkT3iUBOl3Gwl/JE1Wi71v
1TC40rz5ojdxQANRCZn5SU2baX32qzERGDYPevjWVgny+D0tq4FFLB8YQmMexXi6
mb9esi05Ppp5/Ab9q2VUTPnLIXmZIz+LlxN9u9HMed2Og7z9Z/0Y0LFbm7LGvrNH
o/NaxTYXzXPp0A4uwoNu0OCajJbbHJjXOGH5mmy//noJesOkM2QANg2U0JeYnGKC
B/P7uSXa2qZ1zrcGpjVr1ObDtekQ2cCCvfRmFvUoyEqkB4E5GNdO6KSXUrBj1BvB
zb2uCAJn9oaWMFjQ7imdwmWURQqBrMKyCJPK9ibh+GrAJ3yt3jGE8TD5TrzMekA0
QcZzwfqvJYOXchphXulziD9a10uRWtJzxFBpuFQEqfqArEQtu/zcQGa9B0vHRE6X
/862mk/eAZwMuN47eSP5P0mxPZz18PkjOO3PaJU2mbAxP5wnHfLIIOWGhzbefckZ
04NLfXxoe5U93uPit7gnnwHDfiMoUrOL3FuSk0MUl9lM7+NacQ1ltPQHsjt44u8Y
qh9tHZbJN6zjr+WOG7/mzXcKd3T6t6SaSUNVC1NiwgOsCWYeDf325FIlnQVAawlW
MUkirAkU6ggtWIazmVeqKJ/H/hQb0GO4Mj1RPXBnH3QCu4K8VFbkE6/G4R1/CNA2
L82lOzqdLZ2wUUYz8XFXsNV5LvyM/b+dNDtMyc2nCrdxC3+Mqtbi/B/O/CQ5H0Zy
jklXpxfefW+D9TQePWSlo3s49VRmLblpRNerAU/IJjmlGSTV5t5sHoMd0v1qhhJN
KYIorGNP9r9jDOjvNiHUEZkMSadLM5nDkyioRVyC9NEGHN6ku5T4w72dC42ho669
B7s78X39uo4qAxQh6RViSd967SCaogq5kHvpnHMXMoMsfhI98DewHQEx6urjWf6P
j7agYl1Lk9FGQArxaZzDFuE0LQCBQ+neAj3IkxTlrhluKaVbo9kJ1bwbgikYVbK6
chLZEhxeabiHht79Shmmf18vzJ8zNwHScT5+/JTFEErQy3NsyWxz4MoUbMv4MFb1
QmGox7u40+48LgkTgXPkMBNwMwBNaZMqPvXYpZRgcLFN/Hs7Utucw0zdnuPV8Yp5
OZ89lI2DAtbtb5QS+CqB5MmHlUsXQYklT+XChXr5NpLId02Zlyvb/K1H5cSPhiCq
Ja72Iw9OKFynI02HflQlZc+7s2yd9O4TfbkVFCcsg/10DK0a77nZ7CDp/QWoo6YN
i4AGBS8NH5P6uteY/omwpHXZgAEiHzeXMKcUx143tSRcKgmbmu23cpgIdm2q2eF2
9uolLczOVnloaVDer1xR92h2vOmZgspsG3zn0w/1jhDjvhlRkBPxHO8NuNXXgvG1
Zq1+UDajyo6sOW1eYuMmDJVjFlLZjx9HQvR9KFPBklkGuLjLoTpW85Xm7tL9MVu8
u+iITCJO5L7tkgJu0mjzB7BFa9CvxSZVhiVXF5e+B6iJinAaRYPMsBhZn5P0UBBo
rRXOrJ7WKnmgMYvWJFMIkJJ2grGWI3ik9t3PDOBmezYTtkzDH16qwmE2buLOefkC
cqau9XforVRENLBO4+GaMXgqo3XXUpVUQ5LAmw99dwrsII3rGZj40Be7JBMgCr4o
cILA92JHa2Pym9zoSfXQtnQkx8ua+jnGp9b2pxf4Rr44eSlPdFL7KI7yZZpZ/mQ7
20mSBglVBtReXemDorpGu1skM2dsFW4IMPVgaegnpE9BIzeZ7Wd2We2kxfrYAoIX
TkhwKTTnELdCubZFMR+qb4jJoKV462Rw6+ODbxX0QdLPHYSIfz0wummXWkg/L5Dp
u8E6YrHOJQCgCymXDfxceoOPS90DeMRgfStfynIsv7NFdC7LiSQaxB0UYVlvBnWn
j1O5iFiWd27sgb9qPDS3zP5MEC6KNofCOBZdvc+cGHeoDkLOC6q0Uci7GEOA05YJ
0EUT/3G13HMYbZnVU+YSFn+5N51T+VmqFnaqWxVCEqrbOrR7pgbv8midZ3hDTQFb
Pr/9K49QjRkkW3oUYSf6sqMWoaNY6PTr/rrR+NT3cGIpkZOpB5TzlyVF/SZ52wF+
qRDirb3BLZqBAN8Rztbx0WjCbszAUotQfN5cSaNflMFu1h4eplSB8Zvc8B92yw3M
7dbMDFgBrkO6N2Y8X/CzWITuLEnKa5fEGcHAu9ht+bwYSXsQS2OGw0whVp2jeLZj
AB9tFX5BP2iskxuSsDRG9mHXPEAXaHlJeiItcgbt0F3eRQUVk7cno/y4Wp20reoF
SnzqERDPSHiDnqGymNAkU/INRr0FkeTNjLtGJee9j+kHisd8F+HezYbQXxICDJjU
3RJofrJAAByYd0hsBRM9pJTOl+FmD47nYD/YFI+09ZfeusJOAWWbmAQiKZG+IEev
Vwav/0LjoGfZHjNKtYIeqKXY1ASvv165GOJDqh5izozOymu7+saMZbl+Uc5jlasM
AKxq7kc4bIN02BdJsNKFUaqeYPK4i8Ai29Gv2A8yDGKHuqwM6EUTOz2cmDlt84HF
I+xcj+hFzw/LvyDTXI7eNZN8NNiSKrEpbcCR2xVNkeLzEIyV5IERJSdjmIzjY9hI
hDn02Zw2biaRugX2oSyUPoC/J946n4rILq+W3VnZH3TbfobW723N4QJOL8l/OMKU
SqLs8u/3Oil+QFChrjSPbeOg17et+rF2d6cbTLDAmAzUkeGziK5AWpDk1NqEo2/s
SVXE13TIPwZkLZpM4en85yV52w/ii5MBQ5g9QhsKvzM8Wz2T/FXb2FrirP9yJlhY
Q8/VN5LOuPkfDU9CRdK/mfLzHxkh+Tez+l0xIrtg01BYYE+c0hnoOKtldCW3oVVw
77rqxYegLy8CzsLfQ00b5Y0T+Jpg/Khaqeg11Cu8x+dpDow0f97Musfc/JagjhCK
zgDgZHVXkbuHfAVdM2YI8PeLvHX7/FLSRjTEQAsjUoqHTuul78AA86dqNM15jK0b
/5dWUvfCk09yMqXLwfU0en+kqS2QbLc0CX9RC0mTc/rcjQkoyigfVd5UbHMYuWTi
BOO4pZSvgSe4Nzy6s3mMXw+nj0Wwv9TbHYPcmlNBYKozKSCrbvc06t+eqkWvLnqi
mEBcjGg7I1hCxAn1Ft02zn/F8E40ZnJroB63l0G00HAraBOpxor/hiNGUdVpvCg6
KxT0L/CR6TjOoha7MuyOpIUp9wECkI4zY0XfOSHn4ky2pXWISO5AoXUq+ijfqb6T
1pM3ABh+OS/yP2VOG0DzXMVmS4ITwo7CTtA5rElv9O80RXZzobL+T/PUb4TYhKPT
9jTeGh3K+ZHOBfNFRqlpjMoHaTf7RyaTuo4Vn5TXWaHXbQzqNSEgavcJgh9YEN7G
ku1/8qhY6f1wbNJdZ6bP+dxw1mUqynI8728MgVFIk8CG/fN3ilvzFqKcJ0ta1VIy
l4PUfZ8FFVb0paKAKe/oZe8e6jg7BZ3MubtuHYxZG1twQD4kR6mv7vKS6MPir7wh
mT8G2ZtBSkUPmmBTFoOPvfvAkyDvcQobtjaYpemyiRs9NjChCghkAGKjiUopRhMF
0XTR1+ijgAxht4fw9HqjNpRgKHbl9Gazy6rMYG9yMktO0jkix4H02H7g2XgSIk9e
GfFykP4V3V3nC9ad2dvHQQjeuKi/2fO04xYYOEjbfIcflFfcw/jMvbJykXog/wCC
v9sPwCXgIc0u811e+WcQhYDSFSbmi6aulozazniaSoEr3zdEnQUyUfYRMLvcJ12J
lZFTUsFxwBNMrNRHOuCZesP3rrr9Wif/li5a8o1eqCRtZULc2InHbSzNzH+bElBn
PFJmR9gI9HQxXE/Z//XkYeoukTRbSd+ZndFL7bKBnuxbupN2C71WomXwyeaZgHPz
AIZzs9lQx1cXzy1fqxKSMiFevLF9ImeqzU4GMX15V4rcN+7hBTSjGd0EswOW/5u8
Myl5zP2K6pBSZKsaL9enGF7jPIP6aLBbd/QFCcvGnDOGm7q9HYLMMXKFE2QtA7IA
ipGQ3SWmRhO2vIJsFyqZCv1kR/Ef5GnUHMS4bfr8VL9zUtOaL+BC5FiOBa2mfqVo
0zVEOq5jlK+2aWauZawjkJilB0zaw4RK1A/v3r/E301i69X/NA8ppVKqMXQ2ttsh
5t9A/c4baRRQbTtwwt5EwEErDbidRnOBLvi+ypFZOyIyQPFgIeLjcsyhEaqXdIra
6Tk6H0EaAsOVZeYAqVAZWOyxnAzVYlLz0pd789/Ycz1Xy7kmyunHdBGDVAyAcuQp
gKpTLCfHE+hmTc5BKFOhAMd9UZkz6hMv0t8vDoQ4hI+GMcBPrH4C2oKRL8ronu+P
m4NLETdbOMpFPYwhDNlhxLPFP3QeYtpcNOYjLKqAaM8VOmghmkEr3dL0XwS67tVt
15rXwY2LNmXEaWvTb/DHJS0QxDvgfhEJk7jxv3+HPDCtZVC9bXfhoiCYx86NzZB4
qt0OE9Vjwcpz1u76ZGe+UoLsXNuq8/O+xE6G6whDJUWsLGAyvg7NG4ZUDfY8HGxs
ZkVu9NDjsA30pS+qdjEnBzxOpA35XcHpkse1CX7A+BnosVDwcpg+eiDECdozG9bs
b9jmVpSo5SD6uBSbGDFWGHgu03i23vkLZym2KJqRqmSghHvluipgKM3O1TtvFS2D
nal2YEq6XAnqG0c2ZYe2NL9OTl+shSo3jjUf1spBYxo+CpDbWc50G3FpbU8M2Fc5
Zmyx9sEPrYJuNAkDULIOg3eSXwpQa0hlJwx/TQSbPUg+0kOSKIPbQ1kyf+lQ/D24
62mNzpf7eGwU+GlOdnsTgsR6fUV4uUfroD+AO4O9A6zGIoJCMn6KrYhg3WNHn7Dr
vdD7FHG1cJEH+kl2lP4lcQWkP9onjw+tkk106KxsU9+mJwZgZDl7G/Vt2oS+7HgF
Mq8uE0tJe6JXn2gW4qFb8vGB8LYGIML4j3be1TOZDJqspl70RJFqb1EMqkGO4Ey/
Mbbo0uxg842gWo5W0HzCDObkjYHqM5AzXsJQkeQJ/UfctpI/miV8fnciD9R4c4mN
BueOy1oQsQfGR+tKoxVXdfWg+9jXTlm0aJOoeXJXCp+/rbI6kwZ2gP6F1fgzeyol
9bD3hYFuhb0fAUmC9x3tSsg3tvEmoVqc3sO+9DG3LiyhvXU9fgWQ5xA2nvbFXHRN
JYzDhI8x8LTMdixA5LaYp9MMoJV0dkqra8VqVZMTkm9PF5LwU3hjFpppg7gSErPD
A2Sd2/1f/KWrIvUQ+QguqPPF+mH0laf5b0H8O5tBds9hN/QHsYs0uOQZdi2/gVZg
eijXXFa2M6w2TaKiffe5zcsLyQqMWbVO4+FLXPYz4ZgJTcedh5gzidyGk6hhrg0I
uUdtifM0UDwRtDQxLqCyXPrxdqRYSDZoXJObAgiLbWBwAOVyJFFo4+yu3LN64O3V
4H9scfKOWf0SEczm9HYxDaBfV91OqJ6WTOamCdiLSiahgpL0HGKawXZZ8qbJIzX2
sTlvJdEylItrDrhaCwQQl8AXxL/UADt0yy6rzeQeavGLGcMG18xxDlLdDyREPKqH
JBDIy+dZSEt95Ad5Qs0lMMQbaX6oA51p92DYWnfppX/y/jl1+fqG5AADghg+ltSQ
zy6zJUYTpWUp5RVCZfyeyM8MX3CslD47MIh9xlSmdF41ti7OTg2OiZ9fv+kX0nQD
OCpIO98+w2PnMKZ1QDK+rfoH9gA5LP9LUU6H7PMJHB6MAFeul+3u/Udyb5e5R1TY
Kb77quPYNQ9BPAn7E3sZ/1jU1IWY6fDVGHd7ttQM2InU5MgAaYSnyW77qgT7s0c6
Zp/2bO3hJ/CkFAmd6apfxKb/7F9YyQKmx9jg40PuV0TCkTvzkOGF+xcMmrUn16ue
byqnDzWAVmjS+uXRXDnm+RVGR/EA6M5K5HmeH4KcaXUfBflzKEnMxdTeoQ7zW4iE
iRqIrmLGREYN5YMNp2bj3IGhJUQWij6MCc4UawjP+UNlmn3ES3ZvDMnnUXmL5i1e
eYxFveUSF7MrGhUOMK8Uab0AnimGBhXqTz9HYeaO0299wTLizAX5yy4ClW6NEYEr
0LlwShtaux/gsI+nYECz3gjJ/D+ClvuIL++2+RpyuNNTrZJGZUh83qDlFZoekLkt
HyGMJRcP03zr9EWvN8/BpBMJHIta/R6Q805ZyKiwW9C6njZxNFPQ5VKkVJhzWv3l
VcjNfh2l9g+l4Pf7g/ip2Sk436m/mUTQwDDCV33C50O6cwxVFgB6WP1ou0uTCqWf
C6gVHcj/oSO7h3vkpW4qlpkgCn7oHNTV5MJ7MmV3c5xQFAmUe1wj84gCZX8+8gnv
iRiSXB2Wok6BQWMtYaaxV8rS5ktV3FsE9z/y/AxLjPeZ6S/L7W1uA8e1ZqhZpjQn
wGEkopgnZMQMoBONjZZ1UlHWZjoqCFwdmZ2uskk3phC4OPzEVxOD8s7XMKHfTuLD
D1qWCYCTDC22QttOmSkssKmFJ53Jm/QpacCbkwxepfqm409U+meXYQHAcUirVdy+
MupH/wgKG59cwUarC8ABzuofodqtJxrF9Ow/jaEzXeE9y4TWH4nIBe6I4NotoUpW
6VQP5+fsM0jq7oNKnXfFiuf+WqayH5PA7TV08BIdmSYNP4ZwB7HbVbqimTCZAzTB
6uMrc6O2mdhfcKg7CErRX0eTpWvKfN4Qxj0VyGcB7vpiyBhBHUHwYJz6ibFFiji+
u+tT3ny6ip718bDN9OLj88cPKt2SjPJwBd+TPH7o++gMHU/8hJ5b2dHdaNeQN8A8
kE1eWPl3QtfQjHjdTVcqS7Ml1ccu8IaAaS8wBGhzCRnLK2KCHFy/FKroJ0G+EsOh
WMwFENW7rD00BPB+wPvKBf6nDEqF2C9HJxh1/yxkSKMeKYTwwdiQwRL4PHtNZF8e
SBbUsVHGd3MFz5kNjdRaPc9oQTF7XtaDPX8yVxryyhXw5lmtfsUX8ZU7I3yLgVbI
6JReIXqInPEviWopwscggyw+jLh4u+RyNsiQPXR9UTfbxJTUboZMxJvlvcB7hQ9F
kUZ4urZ9ChjXlsNoRqiMV0ks6YhBLcOFzpyyPTOZg0S4TnSHZa/QAMhFg9MVyIhp
6WxpC/kWoVDeQsbE0JDwHEJqSvbWKl+8IHyEpzCACncXkriXS1aP+0Gr6UzOvred
ia4+n4/X0ZzsUl5fc5M4Rib6A167Sw9NhpWLoeyrQy1//MNoxJgsiVHVnP7+aPvg
5EssGPf0n0NYq6CVuYSB+66sACPSVKG7sw1bKE6aeNLifIwwWAIi5FAVZyNRfg+m
QsEi/SGgueOXjTM2UdEaDTBSW9bp6lutxYZrFGi48tQs91cu3FyNunSUgx8329ks
P0yJHOBFyWtdw3xEfguiXI60D8bBSgXUU/hq0pTu29YQA/g9w6tW9Vd9ep9ywzmQ
6hrwjnSGMpxiWKYvqRC3D4cVfcLBHa0hpTO3+AXsjUPILeX6VOBTXgLfYDmzY4eT
yx/vegRutGyMZyJ2vy1nPnnLyx04cQlj29E+BkddHV0B19XJfFx500k2zFiS9uhF
c/h6xzYx5NTvrZvy+uTaHb35Rgs0gx93h/tiV1gCug4Jh7SnMqo8ClunE1iytt1o
+txCeAhI+NobcFevWCTm2Xl0dqY1CMT1SryU811VHGJkBvLrjhAB/Dz4HD+rt535
HtURMGXa955em/lj733O0dyEvAidUEmFV6TzSDqkWGjs4WyfCgq1GzmzIp6yXOi0
1mNS5Wso5JzpaouBEcRLaefHeI2wPkzTua7bB2yZNYCLg/LkHw3/srbpOH6XEYzz
aJkqOPhcIkYSqPejosZ8LaUBYuQgkhhwc8iLEa2wsCmjFJ9xVqfyH4zkd92s4aOd
hsfUOKxjIVLfbOys2kV0W5LKUAluW+JjPD0qdCgy5pcIy/TiuAZdeDZu7jMr0i+a
eBKmN7i9oUAEmhlOJXrg3ADW33bUyYyG9SIxhkV+KRaDHUX1mqEE1se95SHlu1np
ThgyrhRHc+wLXpwjOWpSF/Q7/riM1NbNrCvz2bn7mCpDmD5RmN1Ftyf6z+51ql8t
HFxPHnWxcTkaAnFsJr1jUz8Jv99BMypVNcKIPACkVdW1UUx08DlLad+kdZiP4xYX
4PA/XQ4z+sMm88Loegq2QZpSDNN0GHnyKUjLEOa+SNIfp+zX6+kIgPYv6vxdP8kh
ZEkwuwXLq9NWVv635nK+ccQHuzIQObHJAcWofwnxA7DxBV81NjFBkj+mLH5cgwvb
Enzf7EXNt+znJSVTKiURGE8mzba0LbhwctXN+hLq+WPy+kAsuiNaPVx8raHYRGUg
gZiTvf1LFb9K1d+b/nebQZyJtPYKvF88dIuWrdlXlC2IZzRBDJYChzC6Uw5pXzHi
vRgsopmXXpXlj8SwPohtZc4gF+iJW8tYKalCTd4mNw15vPdagx7cDqrDBBgIbCW4
gsOlgwowxK9zJ5zgliL1c3GrcjQbzBtx6sfMnqpBZYKkkEdsPq1XG0GwSiaYx9Mc
d5NWoUwwNCkwuLpbn4/+WdftNjt6lSauhhbiGKTJ6sdaacqtXm+XLL3QaOnbMwsx
9zSB0IEyK5BgAtLyX5ZY4/Iez2BvvgHlP8Nt8Q5ODQNPJXUcYTuMiYpGCIQXWeKI
WCyT59/9bf6XOkGmWHPv4VOi7Crf+Jr2kmmZ2SRwb6GyahuIA0KQnaqEXsCmzd/H
FhFg3YnDe8n73+DaXFVS59pGLYoC4v3NH47FzHyAGbIJKnnNWTc++srJWYkzSNX1
FJv5KIF732rEV5IqTMyCarNemQd9pxIIxlnkrWTWkHNGM0iAsbskze1oyValxnlD
M/S9Jq/6/zBZWdpwP3aB1HKCEsdTQYtvgZq7s5RuK20orfRNqxE8OCUaBaQ2D4AG
o7UdTd1vKGmyczkxuQo0vy7Y45OVAyDwZOJKIgd64EQPaQc9rgGd3BiXeW94O9NP
bF/X6lcpnyVchU2w35z3AzWlq/y4En4Qtbn0nvv4WfqoiCSi2K9rH/xYO9a5y/ZQ
PmZNXL0cHzpYL7755jFCss0g3BZ1LDDy+PSl+StQNo4CESJwsPnF7v8ibBMiZV6O
HV4BWU2UycUVdMlm6z6i3vWal053CVLex7JJhOgwGc7GTadYxODFC6rGIIsM7voB
jOicEAgdjNxJPQgioa55cJZ9mxrMnmTjY3eg2rjQ9ZEYhJkmU3BR8JcVeIFnKPxi
oR8hz5SOikc99C48RdjONbiHHzL7kaTPu7Kpb7EF2PXEyF3A6ML96PTvNJBCV0OB
qwAMmXWTCuG1PF1AuvAkLVSwedKcQnmDnNTk9diktVdQ6pVYH+iL/A5Wt+QWH4lh
cNnizcjViBIY5otU2aLSaUxeuyHAuPojkNbS91y59trEMATbqCJaZkUzZnPLoN5Q
QdIhGl0OBAXEUtoEA8abbpXyFJnW+vbZIkr7SseOlUdW6AwFi2/HN+0DhrDvNQrY
CfJGHqd0YUSxYpME9rGjUXcoTaXbHdy7iMgtjLcZpwCvjvuk3aeXhAtE4gEic7mJ
JeW/9D+DsW7C5hYMm7cSD4ClButck3ybZPXI1WlsW43N03NNeow7FIxSzka7QeFx
lrGAllttQqu0eQSRXX1HrXZ+JkyVvVcDRETOSXhLZblmCf+iaKPAdXR5TpSrZ1d9
eZz35yyHlnKd4Foe2PQCQq+UB+MAiRdMuIPKDIlvJ+kWpHtgxgfjX6nqpiHR82LZ
uYg3IhIZpMDdseaBZpQnWTIN/iNRXaTXuxa2q19MjfI+DiTCNhZdL1WM/lAfml3g
SSDoKUrSs+rtqBguljkY0tcgjLci+Q8roV0s4HRPe9spp2WR9SRFNHRvEef+UqrK
AiHo4UniqO+Tq4H5Q/Qjur0/xMwvmUiZhzqrHGOFa1b9uLEst8isxJvMZ+5JJEl7
u3GtOTlXajPEG+hEhM0TGpWpjGuEXY1vrUpoPVH0A+6u7kSJKY2PcpemHgb0pq89
KBHh2FhnPN+D6DM05PFfyDk5GItHHjA4ABIRFNZfwY+XLmEMpwYNEtpVsdg6bgaE
FeF6xEOMfdkNMHV1nQuJMxGCRhRbBawyq9U+EzxZCFDqYZLSpgLHR8VOWutzRmCj
cWWfEl/kaV62+S21eEwsiauPa+ZVNCTEYGY91kNJUaxsJFeFK1DgAsXjwF+stz8S
l/tq64ZwJkRjK13HUixMdVkVVq6jv7+G5JVLy49mYbRRJLHEMvnwFxKCSqtVCmUj
75Y0AsyXRjL5Wg08cyUIYvFXCwn+sPNP2GtkClVlAZtJ4XQFPP049BboJlxvoNeV
h6stdx+z9DoTJM/W79XDrgaPbcixjHt1ZxAy5kXbra7P07nRBUqsYvvP4481imGV
h72Ztf0i1XuzENrHMIUNfVZlFirmJXd93/JXawPnVh/Y1ge1YKG1sw+pLB0o8XTq
OItfJNT9Zr3YwY7uSaaVaiP7/RxS6bYfG84ucI13MyvqxHTqPAeX8A8wid5QymiZ
RtR2Xp1BcuhnB0vys8SXv7lqOEnk/bWB93R8Q0xi053mG8N7uQzDIzl5JPfNb/RP
zPQHVSg7OBxRgsoRkCUTTWMOQXBq+aOGOkcQiLYwssqD4MZHNKkgzk+otJv8lkTy
HZH5GLqD6Naesm2fWrWYB/NGhX04iDyRXDlqoA8JvggcPRi0OFvpMZEkHWn+sim4
VxSqkVzCwkFgL+NSKvYQJA3FrvFiI4tlPjetgbAPI7dKczoIMXFQj78aN/jBbN+J
aePNx4iVMb3pgyng4FdvLvtUxv4pFdLmpQp+xPjjb9i1+LPl83N4vKj+Mvi4IjDo
sdC4hnsji01Wf2H48Xmp74dXhr15Ndkl5h3zDw1NVVt30lWvx6FHBHIvbH3//CEv
1ZOCV2i7hWlz4IuYtrzkESxd0P96dWOFESqknzm6Tli29/atsXWuYPvaWqgRm9sl
69QjpvN754SvEaWk24pZZW2prdbio4i57rowm6EqV8h10x35NH1tcDGqeLrVyCIY
wBBY866pkUdJVU884eGlKl6t7LiyIQzo6076eu7R5qSUOkfkcdv/SfnxBj0nKHM0
DtA14vtDWW87s1HF8TyZMw4/EQTFdZ3ZWH3vsy8dAzNy/3GNebsT20v5LUbF1T/q
GUQ90AnB3trzKk4r639/BXFmg/xWbO3VBEduC5ww1IkmByUk4plPRP9ke84FqteG
aKGU3fjLvKpIcZnTD532x0u+CD0ptXgevWr96RCct3JqCQR+rwF0G5GGnMFm0nOD
TPK071qMQ8EIlub6dOQ10353M0ARjTgaLIqTvOcAF+Ysr1n7pC0HNNRijYnmMZbi
iLV14iLJSYq6NkLHielWkOD2mT2spvVxv+BcpEy8K5z0tLPD6LtVzc6dUhX66fFa
iodo1hh4O6JNJTAtT2pbDV8rXJWrPiHSqDzaGfaHrFnZ6MOZUeFFJ2pfzNBsk53W
0xf6YnN2N3eW0AaWx8S/FpQou6JZLXo+MpElDeJiGWW9j4cjJ7YQm7kBak01g+Jz
2ZZ7OpNFnJKd1HUjjppFv04sToKrVD/qatpyBSrIEV6+2ObGcODj5AQsuXy1BVgr
32xjaQCUpah6fuMmYl6af2JQTt5r4WMLgS3mC4seLeAwc9e64O6J+ppEFliOq95l
ZJEkT3QB1ZN2J+Nc2eHBhoU12arcviKQhSnhajKZfaYuobpP5bMOP9lfxH0G8+DE
/YtK30jyGLuQ7p3N+asXVYUnZLSoNhQwbTjl7/ttuKEMpYB4RdVLA93RscgOH6qr
z2SALvgyejD3dy6D5ziYdeKWP5I4oE3O+ebAh9bivv/d1JfTlgR8BggmVrrbNL3C
cm1dxcLN2yXB6x6cLgkmcq/lCUmYyWUYVDOCOf9yofjnz92B+aFk1pgsPTHCKOs/
tpD174DXVFwAoyKOjaSPIVWFWLby3+ykp0W81aH5+wNHrgRHzZph5S96hdv3WFjx
q2Xw4IzDtDgdnTD/qp4PqpJm/pAxEEgMgs2HUGohUAZ/bb6CJ/yxsKP1K33TED8m
uRITi3BREINthHwxLR1snpt4F4Y+2FW510WmLEi03+1z/8J+xs1aeR8o/3vutQF8
uxPL7sdWrkM9JI2nf2087hX6fNDhB6p4ABp5qlSTIsVPsC4cWWrv1Y5DUh6qwuEb
PAPyHgy1T1BFcp0AhFO4wo1louB049dOTALcX7sxeLCeD65ipwDw9n4kayPkt6vd
c/efWVsarly0jVeX+d621kgeb5wX1yYcTTsgUKzDJYVjlgppoyPxE0yZgIu9S2MF
7f7egV2SLZFUANJgUnj1XQLa2ughinogMvhVxgWHsz9X0Ge0ym0mOcL/AEPI7bOI
cWwIasPH5DhZBmhpHOt+zRPrXCG8YMBE0oVJb8/6tvaOA/pmC2of1JRwh37TX/xr
UegF9S5lwflBq2LgBS49KKg9lWImUp5G5nQhW/yoU4NHht/IdFVhngKgtx9GvJ37
4cm5USCrM7p6aBdt5UcPSyqNiw11y1eKXIDerM6QWx534GEChw77aMVaXwhCKvdY
N3xz8lz0PE3MSyEKyjuU9wFbA1Arq+vdJobR4GhATfP0ywyG7k5YyO84Jxf2Nt/O
0yN7fspPF9iqVp0efkGbbrg1UV6zJCMOOf+DsaKIshQNRHEVTFnReBudNSZvFase
lrU93pN3gUHM6wYUoZyqu87UmGFlYnNwalKJJ2UwURtjLH+B4KraMZH7LTCPUEKs
L7bNHN7kpSFivJZme/QodUqb/ApyRfiiIRzoTG+jy1IuZ9DbLSQZ2jvsNBwQOHj+
vbCG8pg0684eOZ0NsTbw+NhNMDVBm5f8JpfRLgE/421zYO73qcqNk0ap5i+Q2vXQ
8eKNo11bcXSrsWAu6rpZnOJKoEyoKqf5CFKl8OXY3x/XG63S6Dto38UBWLj2RXue
dwQqKXDoaezbqbQCoNSi7ypNLSJLnK5SdlwrYo2ySkQU3rFIaBWB+FoGEHfYX5qD
hUzXZUpq6qXS10B3L6WgpWnFfdzM/8rcLfJFBOfIEcVH6dyHP8aSkzZMZuFrbf5l
2qX+tBfY83pIkvLXRO9TgwWzx6SqoDzu0nXJD5WSBX/JBtTaPEFeaFxx7uDkf8kE
RzLTR7AZZZ6yI16csZlNxlbolnV+4MSk5RmjaDvPvp8FVsHoptoTYQkS93BPR/wG
BnDC6FMpDytNT/y4yy3y3qqQeMcWMUXU9aL0bqQhGSi/do5H9zZUIbpADzjTo6Rm
kaOi7N0HUAM61ml2a2wJkPb/PQW+ZNNDESvrrHsrS4IR7XQjl6EkuiB/11oD6Q4Q
O1K3kQgD6RbcOlbqLvC9Jt5Frdul9pVTCaxJSJf+X9Crp6TWCsM6cUOG4L49ZTU1
slKeVj/QERd3IbaRNWfci/r7AWcvD9r/H7abOM8j96+2YjiAB0KJ0/iQudrP4t9Y
HgA2yi2hy1C3w2fAXERHwvYK2XeLdALLLvdTxlWxxrYHRrktCYjI0GA2I3vMST4Y
8x95Lo0gZ1QNbZXfZkV+E/pp3StISEURfA+rX46OAF916rmgNznnBUVrFNcsNhg6
2hQUN+RXoa8fD8CgZ4r33fqJE1AYjcJWFTrnwrEhNURWJU6PuOYqJLncjVTOFhxj
1gDNthMXskH/OKwaatCjqBQPVn+gN0mVvJEx03fvpMgpEz9T5dx7VEhRKBOfy0L6
xdeEXQXxMQNTTzI4/6yX6oQt9gt1HtJo/vk8y+xJoZaRNVfehPP8hSqsLe5yz2Rv
bNrMWa0JA4RmJBDVTM8d7aktwsyqqeXgIwIx7jPEFytsJ7leMshkIHbaVVweP0X5
TiBWu0trV4AZNQVum1CQoeRae/l+/WS1TFbDbz73t7sD18UYhCt0tOX+eHNrGUKe
Q4W371A1ciAEABaao+8eywpaDl86cCREaDBS6G0POLab8nZT7pOrA84Ac+oOdQR9
XLisAQ7sOqaL3H5bXv78mTE6bbFaSGMuqoJOJcJIObEafTYUk+1oqZugnFLdQ2pM
h5eZT17bjZFsGP48kL5kvzV3NBmppZJivkQQ6fp3AatQWZFP5ZP4NEGoioOlLuSQ
2c7DLwNiSCoxHPsr6jH+exC/8dVFiYr8nQOkzztsp/JDB39quI9w7BcsCIS3uD+i
NUjm3LHTjqqRvdYbCYIHOfRbn2i51P9uvdPb6CGbVNwhCCSeYlwpzvweFMX8H69o
FxqSO6BNM98V8XMNCf5Fgx19Y+Oq/kLL6M/+H60U8de5n8pguEyZHKrg3ZFpFMpL
KHjo05yrYw3AaN/kFQAvwgV4hUwTRnwkNib6QTwFJVr4olbbhQ+atoIXBe7iB0IP
5YmL4bhW9D9tqVl6EMsrxeBjg34OCywtphh4Tht1Fz3m5bye3h/pxava4fiBkmbR
DHdAYWv7kHHGzf9P284YkTzfuFYfUB3h8F2Nnntv4VMfnCI1xM6fsBZ/NobxVST2
DAXA7lV9olBfoctS1kA25o5We7vRIC+JlZ1fZUYQoGbBsgC4B5tDY7wKGzbkLArf
TAipqzf4jB2BAge2/U2PETzb59Zld9EKe5Nvcaha/Z2N70pmUmaYjIOTmz08ZS9c
tfSR3BmozL7c/2UrzREtRFKCLYfWbL/qf5bdW8KAV7G3xhKCVE2tmlz1y4QvyDn/
GeFhX5S4cdipcarVHrLFxOY0VPg9CyfMwfjg1I1BDfIBV61F/IH4sak52On6s9Pa
2zq+NxciVMobgVpVorUUA0Bfzz3Qd/7fH9QaUVWD7EZmUSmcJYsavQD63YKoBuWe
22Bag0Dy5kdrvY+6DWYd3h/uAUx45ISznK4s1F/svX7mVyR8T4VXbBA34EuQJtqX
553Nw562q1kcAVPPgujM3VvD9uHl6J6mVshprzus9+8aPgNzdUqRANNo5kBcz9aW
8o6f7/TG+1lVpcFQ3UZlyCgZzIuzYuG8W40NB6VF/AxkmH3KBG4NajcMfdwQx9n/
kexlS2HmeywnyPhMh0AGmmv4StCKadcIZ9HuW2RMG8MYCXQ089kvgowwVYAHCW2e
JXoLlMg8g4IfQRckB7Lu5KQH9ncIqSJkH2dK9khKNCzuzvRvUs23suITSPSpy7Se
exy4elxxQD4C+0XAoQdHqVxx+rna1xahv2DXjvDzAbqEcZMT57/HRzAidxYE40Se
aw2/esN7kru9eQCsCrYEXLqepvcdWsM0DgRTn0ZWju3xxPp0lJmVd5llvZtYXVZ+
h9+ermS4aC721MGwmgAcIoOfEjUAeU1hDfk7a0WstckJ5ui845Co5YH0dw47pXCl
PH5DwG6KeP8jgT45+T2jWOZdEaPGfuYH690299xNjL+yG56fCzi2EIzVhQF/gbaQ
xb9YmRcn3J5HLJpeJ6kfQ2K4p1S57Vid/KVZ3lEut9ZvidvdO7Di3X3cN2TkmO4F
Eq4IdK/pB6lwH25ZNRZjgayI3SJI/MrHkXUuHWKMxO5RRgVyWSuJpnZ+KgrShHCe
FjhqzqOPPbvJePHyyqwh/sYTE71OO/Z0G/XBgqqnfjcJ1gSTmsDX0Rh40gL83nif
1eLD96I5qJtyiyi8rxDCRqAyig2kzTZh8IQv7BLNUkzknZ+VpdNs0ae1UB9HLcgq
aOXApUMjj1FOuiLehi9OeDyrHaydLTtWzUYuhMHr6VapdOsJ6xnz6bpAqpJ+bSld
5OSnYexuoeel1I7JZnZjwM6+tzvF0paSByqt2q1Uikc0yaWtTRP8mAVEqmtGvIxA
emrzHG8AX60ux06qpUbFH1EXFgkF6adw0ySEKLnEnnphsMIq4iE9WVwez5qogZz/
ro2eIRIg0/biWD62XT5tIPJCXWB6biNTq32SVAR8REUP3iKW2Rf4Ms5/9J5GlMF0
eREEQxbGIdpaWUC5u+zmqbu6GdE54P+SVU/Jv8i391qj8cIOsOGdadm3PfXf9kvB
TJg5NOLvSzeYJJXjay3n/SwyA1V4solugs3ShKJL6Ty/pAItT6hSem/1G9XYACSa
g+8Lohyv+Sdy4h9cD4zkZpckzW4vVBBJGu+mg4vZyW2xy+l5yrDELQGdnhCbIIff
rFAYaMlStSXP/mDxxzt6ih9EGaxV2JcsfU4a34bdERzE5/W6ooh6ECYnM8PPyRCl
V2eigL5AW+LI84gHwdLpmYSz79H/GeSs3D5OPCIgv7aa9FJahVFocHc2jswUJjyH
X9Egd9YogOCwU/DOcTq+T3dcD2fWklzy7RPWGQGtFkaVkLe8IHl5YrpphN1yso5n
TF5mdQw7JhQW7uk3mKgCoVoImjt4iBQKB4P68EkIPl2QoXI7I+CehRqRELLHnMsB
oAE+1bMGC+LFXDa1w3KASEQwMmSSi6J/4FnjmK7S5KXQcRNW5uQ0m4XfKBRnMqEo
fA62qxLs1SoJMXOZUIWJXs610rp2bzNmGMqdpmOkst81QETOlmvQJEPd4Drg316d
DLb56UAxscS0i4cwD5otbZgqEU9BbmwsW4oKQWAfSk1J1JG6Jkmv44ZtRvRuCeza
k15r/cSLnpksRGUuQnSw6ycA9bVFkoaIJAw3WExXcvvgzTCjm4WLPbRRE7mYUsT5
oH1kj7WkBTZhKmbYb/4ea0tdXnyH6P9f2lMqvwuAOMbGNhZLRzcnbS5oOznB8xbb
s4OzogyluzapoNYyV/xMUbZdwItfgM0IYoGKLBMupAuOTp6qEn/E8NnnGOxYsKZb
aJ80ARfpN9dsHNHBTIo3n1KEyYUTt7mjF9ZBnZ8343DWCf/g5PAevbwzo/J3Sm70
Xsy1O2coSiM4lRsbtyYkIrdBT2T76Dt2a+WXf0KLxYzBjPbxa1kDZzaqPJo0WbQo
+ATfikQ7M5usb1Zpek/HuDcA2m66TDXbroYoIYRJHdi4TNnQ1RRkU95WeEF/Ar6M
KfiGS3cY1IYw7cyvo5aXvgPPmcU1S83V17WOmuQeLjPHraY2t2rZIw3SYE37QQ91
mCUepSIT14sOmtqTfSqoXcFDWSzuHZWfjFf4ADpsNJVln1s6i8OVz2aeO4y8ixll
P2LWEMTyzj8Hznh+6JylQxhT3/KmeJkvOPD7LE50UYQcrOpKUw+a+5hlqwcMp7Xu
kLlMciNht/gzldhf9C6qblo4Z8YYM5kbCpIGisl4l/8RQF8LtPThzdOkuMdXae5s
sSEhWFPOF/1sfa5+ETPOO19gH0aypamzD9PpYTrml7D8iUOc2uaekxDPK7CILYhu
lkkYSSCOxjLAleOWbBM4gqhONBdISiydnwAhEHs865X/HYqRk5/OUShFLgSDtP5M
E4g8LZAuzS2UsRNyv/DPb3TzLW9+AabxDXr9pNE+vzAI3J6q9TTfQ5z8fErBJjc2
Lm+kARs1kYEqQA4ZbuBSwz7S/rxiDA0ruTJ85+iHAM1GF9Tuo17O1A6rEQ3kgVOu
WgOU44WRwL8kAG+g56x18oKpBQOuBXUGbORihs7jGqSZGFgoX+0ulCAWBMxAkhe2
tmGeZGAV07fZrMCGUriyIfyTfPE/3rvFm+mi2FRKd4QNqO5dE+NDLK99Vp5i8mwm
vSRKPoeKqW7R/E9auP4yvDvfuOt7CV7q59GMHfbajTh0pzFLdMtZHb4hmW2BV5Kb
zdFR0JjZ4K83uXXy8NoUaP3iIkom9kqJIuASemQIxGrARlfc1tLayqTO8sZSA8W6
WErW8K7UgQpCV8qhHr+zWaq/qF9kVpi3Pcg/yOBsf2t+Ulewi5y3p43aX4jiFgPz
k0FvyT0Hu8chhLYj8Ps5AA670JgLycKbRKiNrIfTCLe4De0a9CR0zlLUEtjjnlRW
L8zw74OOq00volAcA5wYey32HkP/N5pAGgBSQuRgRVyDyfTsmyr6a0M5DgLFrsYP
6s3aur6KchOo5mtkvTBH2Mws/QQRoOiNGkD5WaJhwrlSn960oI4rxLuSj2TpPRu/
4R/l8pECxYLhtV/PmIjcJbyW6BZLJXN1E0aQcI8di8N4DsE0b6CfGmnzoiJxxTho
7pQ5dmtMsjOGa/3GICIqTx6OeHMjkeoMrIuhDghvpFFKLD7rfNudFVMcQe9LsH54
YAS5rV+7k4pT1GFE7oCHmHvltL0nZtFyXCy8xI34NCHG/Kcqaw3VLmPXVMETONL3
QsUfxU+kou04BTK6zvkr8yy444bLOqx/OHYtTIkGks9vsHOTyROhWopJHx9YPoLD
cTYJbSJytwYHlHO8GLGU7VU9y5xip/yRv12/8oFDgN5It1hd3cvqLqiYa3t1Reys
qHwRvkMy8R877g+1TTd2QsvuOZULEfuw2bPpRMUJAh24q+M722hysqd2GX81HK60
w7nPxBBJQ/KtLlE7hq0jY/Xlj3tur7FaI2rJLQqEArVeTT7/Wy2AtcqRR4rztd0x
I8XPH2nkGL7PQfqJgaguhcA/hXSr1kh34l64VCL5l4DPaq1j3oTgaSLhYIjwpNq8
3/p+r7RU+nQ+dkRuCUCn/ZnOWLteWjgeG9XMKus0AUOZ93QiBP4UZjCskdUgZZe6
1tll6boQqG4wE1FvNd6PE1NMYvtf/dt8rudUDCbJ0QMURCeblB2BMNDzvQsTjrAs
hC9RqOud2/QKNwYv97PpI+rpTysS6x47e/wfWBvpZYNfaoLziF/CuGXE+ig1bLpD
Wgy7x1jx1YVWPk6nxNv3oq/rORf2uZ06Cnr5jBa+91BaE9gz+rNQOj+lO0qT7Q98
7pu4XCcakPhHxfCz3juuQvbeQQahMKQ4dA+fBGDE8vsqU6LfngT/aNRgIvOdbMUY
UhT5GR8cPNWS35ZWpvS3/MFIrVRdcfyrvPMKZcoocRfpmAUmTC6HgR5jBAEU4LAn
6Z+FjtaC3ty4DCYCuZcHlHsQp8+Qcc7f9dIp8LbI6BYej4wfJfFGOAPSnUwXL5Aw
thP4l730EPd/a8UTbiK9mOZcW9djWp3aUn1Ac1sjiQ/iaF/MWsFHBCPwnk2iR8mb
0LDn9t5nThK027EoZV+K4iMuMHGk7XWQKT02RZ5WThT2702oiHEaOPYUdgvFG3fi
988ctBHyYkzKBdweoSOFiqm/vQ5H3/Afn0CDX9i+5qu9L3Xbn0j2laJ/WT+NWmoj
6y2l7BtovkMNNC0Y1j7qYvXA672WP42WEQClEjOMDQMnVIxSVt9o1qukX9woEJSo
pE/cTzj3qbakBWpHWE34c/tljjSondzUkXH8L7DLkhDwtGGeFF/ibiW7lyW3wqhQ
4S28HhhY87gFUpJ+hwAt9m1hQV1eXTm8Z/lW8OLNnhPJWjDsOdYVpprwuYuSoxut
gg/HTgHN07WMLWgjsoS+/PL4X8exccUmlpC6gO/Ca18ikWsZPdDKeD8fPsBCSiQ3
h9Jj4t3s0CIR8n6x1+zSxLW39EBK2jAHFaEctreJlwQdrg/Ns36MvWAVY4Vu1tct
q94T0GXMwBj+kdj6nQPtzYJa0W3qhu/pHsVkqaTJXVoZgXofcYH//QFwi28ZAjdy
UJR8ljV8S0YqrZERhuh1hbkGuPBeYC88WvMNdvZypew=
`protect END_PROTECTED
