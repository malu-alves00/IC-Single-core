`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/2AT0QZ16fCcO1ymFKplHzCAb9nt2nR1URG2a5B+/6WZ1mCpFK9fWnTn1uL4ze8g
BeTKmaX0kIHowHYnTlWNudrIN+gSRw+uJiLHyU63NQJqyotuLuUiDD8DAULNMX37
HMqVjbQZpIgjEBNVlEcWJu1MzN9FBkGUGvOxJ+c//+bsrTAW8YYASZS05lJ/six7
npKTiZeFlY/ADE5TCnRBOV82LIw0gBetrFnH0aJ1UsWvL9mSDlELZtvuIkg6vHFX
Kfe8b1ri3Y2h8DBAzx+Kc/Skgph9ScBVbvynTRSJ9I3W17mlbS9Qhkese/FuaRho
AvGglNSWq/aGW+ltLdrUVUaNfarEgV+hngobko6wZvC1nayIWv53lLjToTIK8Fyn
9bAQeECAkMvlLhPI8w6EJB8GkCMlpKZfld+9++DwIOju6TplvoBS4d2L9oKbdp30
7tizXdnOF+gGsTsLGURJFOtZCCvs2BaN5VLIK5809aBDoJQ2JfZEZ/eTYw0ti3Jp
vA0gSz8OgNx5DEwOb4RNnY5Eym9YP4pSgb1pWCF4/e9ZClXv5pWfGRNSk+5xUtGv
IvFOB7bXVkYdqJg+SdaY14EWz6NIjFgujkOoV85UnykHsJt1e6E9c+SUbwZ8sFGT
9Udi2N7pw7GsB4vLd4amxIo1fT6lafW09UyDKdTHoa61vBhJ3rnLV4zFthH98T5C
EYZqGyi2sgIJXQAkiT6Bu93qDrXfkWYe5YemporbSVHUN9gMJUCdgS625dxN6cf+
Qtl7EZCZi4BDEsbi4Ho+Je4w8c1pqb59UJQ2Wz0/jYYF8gdHecn7Y85INIEYELDL
N+HhunZXjIUo0vsR63s64Plo+QzCqX2xf/q3FtYUWFHI0v/zwZeZQN1UQxgglx5f
FHqER66pCdqvkbXepp1gfJlfmHufwTYY3NkjRvzgCJdZPjRICvqOxGTJjl1+P3Pc
qkwc1pzsLH4/45/M2QLeBxQRCCn46OSWKVRpYYYXjwsX6WDIroU0EcYjyP57E19o
67AEtDEI+BDz5wxqjrmT6Pc4WzmaT7LlBVI51GDs7fu1xyONKPMtwxGJVIY8qXvd
oUQETT0orEPGfq05p4bYYIyrGg8/AjGvgXJ59oYIKXgIbuMOjlfv9f16IofgVJi3
X6nM4pcKIF6K+ynzUhSMNg2FentvLigX3pjQZ+pPCQaKpHfiB9Ubk+vr5yBFQkxz
ZzRkO+CLpPhtcfDZtaMJ+VhUMNCJDCpUl3mTnLbQVJk8r7xOw0Bv729FYI+chXUw
Z4qt9/m5W0Qf3j/IpgK5jCxiDBou9rRZNCYOrF9iM3Pq9fYUQBa4iPZN14I4fnLf
ftqmFTyjFZOOSeNAhCVKwVvkWm9kIdMVP0OLscHzvrU7H2Hkau3/MGtOVW8C14/l
llINHLA255cdcDBW6pNLCUPJ3zAgWPCACJhELAndLBRlR5R1+uQ9GVOIAqVWxjbQ
ecHW12+yHIMV9205TXM+7PQQBaEg4oJ2+Wy58tKqjXTRk9tWInWHstUzZkAO7fBp
I02MwG3MKy15b+hgPpuiCIfHZgauTypSGrd3Ne8bzsq8ZdS2yv9VZjbsnnPSKYcR
xkKhLOC7/rUJg8BcNRSgvkD5qyS0Wpy0PsxpHwjI8p76/uOduGDwtn9rV0jbl5Eo
2bTs07GI4/SI8GffmTBAKYfIFQfybRdcaG5OiEHA+PFhNkowaItwMjKbPK4uOkKL
A+AzhMFutn/p9oKckBznKQn+cCYU4yWN4/jikAhD6SxANVigXLCRbhwavudTWjsC
98b/TU/WLsdOVT3V4ExgnBgbpKHtHkIIIhq3aTCTqEECuyIP1f3t9c2qTIwqA+lR
VIuS6EXRgYJzxFsowYWxZw==
`protect END_PROTECTED
