`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8/jcxDO0BTm80h72OQLBtablShqxlFEXnVYT2r6IEyA9HihhFcl9YPltMpB4GsGQ
z5vJyEkrFHaLuzH55rAO1Bz3nT56ItZIrq5x5/hFwapUVNvFy5fscejwy7YqyEEU
6jAjShpOZBF0IKNrSPt+dc6Baxn6xuXIgafBVaWOCXnh/5JmZ9/FABl6K52LErDx
6ACvDo/LK/ubOq1kvssQ9FEKaHbinWY5iT/dv1G6Sp7tP+3JWw8d5zOSi+stnMpd
O9/G4Z91+9tK96rBVQNNbn5PBkT2ax9f7uc6wMMSmIBKJhm4z2Ji4UG+h1eJ15gs
XOe6Ta7qJ4Xs78UpNSTkGPyQUCKbiiidK4FV2CDX+LO937sZ0/lVJA1c2cRKx2mm
m4HQTWt4tS8pSjTHEZkSzbSeIQb/qXasTFh81Wc+aQR6zPrCCVOZuS5o6lWTssgq
wyMfrOnsZ+m2RaKNvz0FiyXSj5RCWZzJejpuspn27TMR0eQ/HDUN1dgcRMNLouTi
iV1XBrdSI8T752CbTVg4SUjCOGGRFstzgLhiZ+CGCo0LTwA4d70UkNymZDMNZ3u4
0+k//ShcUc82P45E9e89kcrpn+Ihmk0nGQEeF48cb1zbW0QU+OiMkCyvoJ3ZMoaO
PgdYeOGcaR40Nwjz51VZeNCwlx7UBgawrmcpg0QwDIozqE/fD0OPe/7oomlh0Jgp
+ySEFuZyDeply7iYIo4/k+limGqgDEGyUFx2KGtLSKA4gWa8E0KclLlIAdT4fxmn
SSlFPFN+AenrgJxBjCQiFit1t59KtBik9Ix0+hShPY3sj7N500E8+nywYDx9bCpR
d/yzJoZu7YpE277oZrXf9g==
`protect END_PROTECTED
