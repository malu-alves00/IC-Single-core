`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jmcuQFDlLtJNooQyrXbELPKxuBwfCM0sP6T7TjHHtyDYz3hjpuDGZBkhFaBUsKiB
wYuIyLVX82aMic7MHvlfBo59dHGHvfSXA2RJwuazNb/jGIb+0Sy1FZd+G6wveSI0
o1UekRUHtMQsy9/XyeJMyKEuLaMlK6lfNOf21EzU9TQFAmdrht0nUu7NE5oRVsdl
`protect END_PROTECTED
