`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0uljubMzmdVlETPX60UlnCDm14WEYTeiSHmcwdIVoJwKZlcWx+h+f8x83FvsTw2y
yaP2G53KwavJAPijuHZe8IWjI57NfNvGpWZvdhC2ixpxaQ1WsSFyhm53GIksFR13
Q6SkkOye+qbIP8QgaNQg//LHie4a/6TmUOOJWwFE0Shwn8nNQli47Cv3C2VXcguN
6wLWN0N5H7WX21EMfaBlwwFdT1jSCpN+IDz0Kx4sCspz89jl3GdYjEODv4dBSNLs
lbe4G9mz5ShzLyAW1wW/tJ6jyYnwDzHXQEQRI7xvxno92CR4MIM8WAHeqsXWOKMq
/DuC+obw6JDx2mj5I9pu9Q23CXOGiArpWYzk8Nvmrpz/YNR4tiXkVnPpuNkPsy/w
XoHwiSyN7DEyBol3a2xyLU0KOSc7kmemrbPDQWmsul41+NzHvl5s08BWUHTFLHaL
IA/IVxD0kPSxV6Pn7fGvxFProE1xuPk2GoTd2hVytj/R8QmllU/vUIO0j2R+L/wu
mpaNvmiiJRkaNSRbzzwTPd3mW0N4moG/GtC6Qd54QZnYVU+LFFbzH4VmyMQYXeIw
jQVDqAYelaJHIF1ITj+G04IA5dVJnAb0JlzwTadsw+wqZgyoyMS2gKhqlL6uR3Ou
zzyb5pZEnoeyXA8N074/cFSVUEjRUyhaW/rW1CxzyLTvtCayDSHZbNIV24B+qlQk
PsdSz3bjwcLosCxgV99XGVrTTC3egtUB+LL6RDO/x+ikJ/aviMDjXDJwRlTghARP
rTlZN9aHMmmDXOUsG1EfxjVQeV/KXauinId5f3KyUrxaTSVfaYqRm5ZMZjwCNrtN
oriGSFY5MN2Hw+KTZlbd8pEsdAaRS8HAL5cnXSEy+CHKCIcSi+tmb3odr3fvRdEP
mnf7mtQP9cWht4c7hk3QSG3QoXlbo2wYF75VXcX5ClZ3TOmfcgPnIYpljjRnmOZj
7BzLMJl7Rsh6JnJJi4nozH88Y6zyrVqBRZBQ5A3DbvPxjdKZg0Y7pG9D2dd7Mmap
NlF279Lw4PaJ5YAL3mxDfVltvD1l4j2GyeDPEqQs2fc0wOb/Ogq3cSQ0zNA1bIZm
RxnX5gZdQz1NmVOb2m2NHqmA4NlFwJzr5NAgPreqRlpDRjkKrRATutiIXkgTuoZV
YyzHjYVWeWznj9lJ5Q+zkzFLfQ9kN1BBJ3C7Jqcjw7HJGFdfhqBu2UAlLmu/W5pf
zpauy1spkItQLH1U56nlvE6vX3rIWQUvH8bhoBu48E2T1Ll7tgwUiAFj5X4MQ9cl
J9tZAaAB9bpnNNwjAoOmdXGjYTzW1SNGL0qDcrHs+jMt/LQXryXjqEvT627lDE/D
IDdCECdvZfees7Cl2Ih2EAkNkK6kEYVd33Kk6DxULN9iXrbajH8FzTmZ3dWxONh2
GC0jEBUIMW2AqR9oyBP+y5Mj3FHaU0Gvgg/WHbkcVeyQFLAjtjf2cvPrjnw2bA9W
fqKMGl3pK/QOWR/zFl4G4KjQrV0ffvNI9kK0K+3rJyeTbywwIiiav780hhf+fNDw
Zyu878bliOxrdDW1W+GmDAojIyZCRZcoJjJ/vz2KrQ/X5pbDio/y4cwKqnHonU6k
p/fAb1o/K8WgDKe5tdsGcmzVsUXwB6hK19DpXqdCbfE+Yss7gE0zjKYfQMblccYs
epSCDp5qh+FwfJ905vvmT5/I1aQqIbRB+xgcbqAx46xnbzlba8wVoG7C7aMoF5GN
f8bN74AS9Z14eWJOldLMlxMmm+PfXn/jitZS8koS1Oqw5vi0cEM0t0UF8w4jSiMM
scXRkevs7H+ZK2CIC6MYi/s4/pLaaBH3Lm0ShVuZuYJCqV4GjTs9jFZxDNxZcg9T
t641lqSR1QQGPGTKeQxN6n7odq7+b2TTQVLUOv6Z1tNonrzKFp9Ccwo2RKjXDf8r
Ei1o6aoNE2fjySqTySCtYcnzKlF8brAtX9ZlyrMpmMHBw4m7XsJ31O2ar/grTzD+
lqrj9YqQI/u6IyZKZsLVT9LOSDH3uFVc71wln4DeEowd+FlfpKWJIAlRR6osoV+F
vHiBJcRv8lPKzm8B9klRHy89ptkStOrnpdJ/X6M5OFJJ0nvry5dlHcv6iurf1++Q
88FPvI7L3XHnFKDB/0wpkb13SLxSI1dpdfBw61x+xNIgg7ajBy5oFYHq7HyKc5GO
TsaBplHzym5Z7PYKQYxdqtXbI92Zqp+L47spVy5xTj2PvSxj5okAuR4Wm7vy1R4c
OUh6RpFsHPe//7n4/lsUVVlwFBVus01F4otMub4rwv+i7Cm0JR+1G5nAT6B0/uWp
odX9zCbPoq1YgKRpd0Mnm8jvm3mlwfFzUnQ12EUEpabrE+vXAByMMgGVNBGjQ2kG
6BdgFbrfCZGu0SKXJT0Y1tmnuk9KcbT+bgeXQ6iEJYHlPtJ1RXwxT1H3kpvYjrjF
M9m/jfU+zSAduGDmWdnQnAD+YYIFw1jAnDB3UBYloJp5wTcF43LjxXWHkx8DKd94
CRCR3nOZuaKvSbFar0Yae//0OctuOgEV1Rw2+5bM4b1Cef5TMx6QxW7hNV4t/0BP
/1rzsmYLV8HepBskQnwsUdYUtQ8Bg6vO4tCaMUa66615KgCDUYoQkIyldzQ8WaB3
hU8qs0+rly8ZDnrU6+CfIavZcsZ5G4n/E9bdz7n/EvkCBIjGSeV/kA9poS7DgoXR
r8r8HgnI7KpQjBLo90g28v/wPyRjbZqKCja+gBCQUYEh1IR0wsEQ9G5Abjopp7e5
sgDVk4Hgj9PyEqxfmPbJuVlnRY5AqgqL/Jw1LeosSe6qmk9TWHpYwjE+BQAQ2elf
mntNhETVBOljNOIkHfT7/LiYqnCLvsYpw6u8eYCSy1VUoyBzCr9Jot+pym4/wKwc
W/2CWjrR7GJ3hZG1xlH51bpFtzNXvTmx1RpY65abp1Z16NFsJBNquG0vTgJ2zOSw
gYQUDWK5fLXkG1ADPbatVZvO95t06GZP6xjgyHF3rso54u4KKbNVnYpGuIsVjPDV
qAMUL9AtShaiBUMwsS0vWK5TxNsQLGvG6SYPyqbvpjTmptztKd1iI+ijmRVzUoTX
/gXYxqUj2NDGTmBjXaKF7eoopNH5dCbxCrAFfM28u06MbkHYvqZF6I9f7GwGcW0q
Cyz4Irz4gIeaN2nXYF7kCNj+On3i6AzMsu3Vfb0slcEILDo1OEIde0Z0dKhLuVHY
mOvo8g2+KTp1a2/8i1X5Iw4NK4IPM2X1MBgxBcRAgZqV33D62GIlhl9Xd812ZI0G
29XXWSkpNRZPa5D4fIT7+6cJIhXffNqkTyogRadSZUZ2PU2ApFmkk2i/xjm/eziL
Ttibmspmdry05wO6Y2UgslFfatnQ3n8UAMLKZiE19BetI23mhLVuhtFsd+OMLOjy
iZ1zrGTS8WO//ndZnWEYCqnWJH8DLb1uF/pMvNeIuFEvQZ85Wz9hTZ1rOvk7z8Hh
JALJkUxumnG0NL2XZpUSII+LoGZXm7C6b/oqyMHyysizKHcvNywfNHfgiA3Q1QWn
pdKFJX14KP9ypwJrqOwI2giV6K29FfG6OmphH0bRF7kBNnjUcG3e/f7s5u+K04HT
o++OAmw8JAPvnG97iL++prPi4bSPuBY8S80rykyaxOl4rWKRZXwWpWc9MIGzOEX7
8KHQ0Rqba1QNGBZGe+cKQzUxEUegdzWoDqw1bmY10fd/DG8tlx0D8EQs0oI1F8fL
bVqP+K/GToAq4Mb2Yf3e/u7AYXuHQpZfGq8TOfszCijD/4lP5XsDXO7edEPs83xJ
PmPv+95AqNHzNMC7u19Y316wz6Ft+mq1QcG4oa4Wca1nosT+/24aPbyiCA5GkkVe
rEqBS0Y2TvRkiNVrHtH+HQRgpYAHojX4QB3zaU5xdOU9N6szYwFWKPW8VwPTtzc0
Xhr4+Iq03lsy1CMfeS/F2Mf1hYbmP7vehgqVAlMImeDKt1ZKAvyIVShKgb03//qt
asMsuLIoY5VRaaI4Vj6d0N5NtBhu2CeoZTyUwo01yF8mxH7QDRjGsiEr8w2zCcAi
7YIq0271NFcCjguChLhjvMA6ya0sP8l1YIZABxZH4sj6lJAFthyX4I2yv2WrNIDz
SV5sNjWKQZMiWLQZQxTfnNCr4NipQ6y8V30x4Pf7gmtp4iuJfwxZx/IGrPeRzAq+
PjiuOpbPPtIsYITW691maw3xgQ0G9SilYYAwXKVWi/ZXflag2c6tAO8CKUeURTuk
ArlwB5YLupkFLzmcPN9ZY/VwFFwSVTvBoMCxT1OyT1LuSqQSkGAXExPYHs6fwUGG
3SO9b6kk5kx9HCxQFpROmTXURKTXGH5fdx+7S9291O89bwpsUMSS46jwnBe+EwQH
/wi51qqiSANQ4yHef9NNy60WGpRhSdl8PQRYt3NgcIoeblYDsOr4u1sfvFzY9fgs
xcLjdN8yWVN3ttkKwyk0JR9Ah3DysT2k6uzaP7QUPYURPQH2rjbtgFTYP9oe0ctB
tR7TjQunbc7pioy+iZ6xyCcZGetkclYM54DMBuIxfVlvHCILbBvFArs8Dr2XTNyU
6PPBkGhyek4+CRiVaWXID/yRNk0W0Vwid8qtrEzphfyzg7X8ROdrLevyDFEQADkC
+ABB74RiuSPOnzho5y+bkuViI1UoHih/agk4jX5RGFpCqXrtxnmAhcKoS7XzYkMn
Hlm+JhX+Zofl2ZCPAImiRWVTfLon+z91GjdO2WZblpfvYyGbAbBfzBwN0FLjWpmm
rhrrcF6znQIbdrACeoROUJRzC2ywfX5T21vhL5KJk3PPfYZQvEV/6sYJHha5HzTn
8bch9afTf4577gudY5cGBHig6sIcGcaF6ykLP+ld50mQcprhb5UKLNsFsBTKcwNd
inMH09nT1XhzXmHL6F4ufEoHqUcwfwwi7dzSadQBLAQU/eUq3M68J8iZQUMypvxC
0FFjR0zJosMEf4on3F+t8aXzhPqsp5tGJH28mTwmqZ9GDAfw1N9Fm6gdxkvD68A2
BWz2mhW281zY3pJDPSZJ/MZgUJ3PXYnvBndc/zeOyx/kC/fuZqAkpwdpI1ICtDgS
03nIjNA4drz8Mjh4PE7Nk6LGIGgC8u5Ee3qckjE0FHa0PyUPoCFN6O6bf9xasEP9
912Dy1EO1UtT6AinLJm2e+8aBzA4WLg/Hccyc7efnS/8FM+DresHwaWcwlOlYE+S
kNtQ/ULu4oIO+IM9vEZJcRdxBYCZeJK+yaNI/gyPnXfMhMyMWqFATF75lzB/PpIT
DASDIfcm1f2H6TaS6yPkhO3tgfOZq/8SUV7LYTxTaNP2jr++4CuC73/LKQsu7hNm
SingPqzOT0vpRl94esbPitKZ/6cj1VJbJ5WxdMrrqV6Aqs8dsEdYw1WkmzjQs6bj
Z0pZZ5z9nE7LFuqMurilK/EUlHxwhxJKhwNXROQR0Da/k/N5saHJAYJdq5UKhaUs
jTCW7a+o92sDe9VhtcJ1+r0uo2Mv+BlIEbqaGJYRmJbHcko2xJWAFJk6/YJpLcsh
eNddCKor8wwW2KNsiwZbf6Mo8q+t3kTaI7U0yk2aY23g4AGPTalmRwjySDb+XLhx
F+ONXABQH2PdVAtSZN/EnhfK1m80Hcpf1DeS4Q1CMF+8d4SiF644K37ipOD8WXiS
Pmw1dTZpWKyzi2jCGaRtKNUSVit8FJFohZMAiWRgHJTWPBnpVaf60NR4gUwOlQAe
CW7KT6NsO8ENqaoJzgI4BMo1SMbGxJEFYoZ0i1jDxidtqkefPR/SWqYNdPmF/KVn
KAPltqv4LY/gdfQIQYnRkMVlXwvEPREWd163v/dtj14ExbNJoneSkyNvbBnnNzyt
ZaAL96znWCJjNYNCL/dtXuYnFpmq5Gvk1z2C3sqLZZ4FsrpRJe2dltjK9o/j4tWS
HOLho8S3etN8cQRPm8oBKW5zJCktz0kt3FM3i7A4DWVxOfY4T/YgsZ8zJYovrnfa
X3vuJNHm4zJrFcpCj8BBmL3BriJnYLLNlAqBrZITGyykCGOEIrE2mWal7jEXS0Tn
+/mmkOKbgr7ZNLkSJ4AzVcLMxVY+CnqVP69MVsaQVTyWirjGX1YLzGt+gizL54Fm
w7Mf2HtpLwmmXR5Jj/Nh6jwdcG5hho5bYiceqAozve/7PX24RxP8DJW/tGIgD8P3
fp0xwnlcNyded4Z8sEDamM7K6NE0Q06I8pEiX76V02SV22HwZ9tq0hkb2MXSk+8d
WITQTUKgaDAXO8MYnSaqAuDPuF9oCSnqNzAH+8PhELnOTrDGXfdH+QOPlQ7stL7H
K/zxVZcZ33bEkYquyZ4/KX7927Ddln7OETCk4J08eKFIQXYxEfr1VyDZ1ijQLuA4
wwjmZMH5IQ8Yp8H/8UVyHgw8jVuz4sQmGfa2tGO9p9Hfe+gsUMthulY0N03JmKds
JlN9L5EUMtoO/Rh2dX5xxrdtmWxeLmxL0O92lFqTI76Pe0Pog5F5QPjdvrXUQcvy
3Y2KrPV6483QYanuodleGLG/KVNS6VlaEhZ3fPjJYeHZYEQHuiGYy3kVknUEhRjY
94nrZlo5oRKWe1Ud53Fj7OJQJEeMuk2ZrzKx7YdCJtclL/PbkL9X3+Q3ekne44s8
d6zv/65gQ+1cF54kQswMRckS//a4hsp6r1wTI1jTDmV1JbPGVG3fotnW8sTpfZMN
n2tIv5c6QtXX5R0nbCtkQf4dFd5jajv5yhnd22iAMcxMawgPl7WmFlJARLUhmi52
eN0CAoReyOMbJMrNEmncbpoCHX01xNgsQK8tA0cw0MCd+z6VThncWQjD2gBVs9hc
DXff2pV+FqXTMgtvBY2xzMIlOVzMEMNsqYYnao8TqE4vZ+CnqNSfJxGtu8BED4BB
iQqc5r5aBGCg4Ek08gXRsOT72HoWLN1270jRZ0T2SEwI+NlsGcBxLvYXKQ2g46xO
Cd9/3UNte4SCrjkyZlkqMWVggVhACD32MnsvQRr3BmaoKKtkimIXgSW3CPuABgRw
2/6KFu3/IDEqAXe4sHXtD0XC5/pgOkf5dmIMZJAjre8LaXGiEDXeTjp/kS1ZDpGd
oJ/dJgKMsMJgQGOEqUnM//mc2deUHEUbRx/xCDAMRNHSOC6ctvqkdHWz/qscdS1m
FgJYFclc+OPKUjvrXCYgxo1eA9EQCq20FvaW7RUbuVQVDW40Uw/DWLAGXwkiFSBG
6j2pgfO2k4KFZrIeMUQmwqnacMZdZJBqzwfc9+pCQmI5ZH71ZaZZ30QkGT1gopGr
to2RAayIdNfb0G5P9rouVp8EpRK2px97mvDCCKKuZACK4CuW7iOneOucJs19F+TE
3iEe+R7i040K738HJqyQp93FGb1pLc5cWlB7K3anw1s4R/3/MPrpCAIn6kG2yU5V
6HqNRkpxnA5082zXrAm3wpR756F1sJfVALfnyIEvcHkqux8tKeF6vuY+MiktD2Db
/bDyMbrM7P+UF7+xtB/uRrasSZ7xxR0NXUwc4IreZ8LXiWU4R/a8XpNb7h6uqTRu
EAymPmmYAKfnURp6CkHRqFbM4ckWGGtbl3cT4np4oMz9juwbyPV3+mYN/4oevGkB
5eYVZdk8ShyMDqCUkp8MxhKiglMfmyth9to9hleWeplHCIOUXczaJNK05R1wYP1N
EzYqQdju4gpCxcQ+914hPeAayhwpYP+Hh75Y2qvsVtIFVxHFcEMIDzVdPb1UvK7c
NWx8M3K75CLIxuGI+lWJDVZ3/0SnjLZ9NzBIQJQK9priw2jxNdZeXlrw0S0jcWwL
bx6winfraXXNJifpuLMt09DSlY65I1tHV4aEwm5f9dlTowU84HjNZybodcKqxS0n
gJfOKfEBOIZZDrowGaSal8QT+sPDrFTxmrbo+bxYbgAiBik4qXpYy30cQBFD8QRy
zIzxTcidO7t4Q8UsvCV2eE9ueE/GIo+BOmPoXhJRyF9XW1+AekLw86EIVVfAP6pG
ccOVHUkXB5DhYyPjPmRryN96HA2A1+ijGoauQ7I8J+pwwCL1GgZDH0dyLSYnDyak
QXefZGt80KXemlDR7/k/Z68rTYqxy2eySPTk2qABrPzMVYZGszCeRuSrX2MZKRre
SkQTLFgJXg4c1XKA2nz6qgJErIgUQ02AqNEkuSMgPxhnIVwpK0u42d3jWV6d0R8j
2rk49zvr69p50my+uiyLAvwsRd4FkGsSrfTlSEXu7DhcRPVElZjnUY4/aDPEXich
M9fvP8ZKjOkf3hE/0yc1CvllDQrNsQKYyo0PzvMPXw+4AcrRIgOLBlL+NDZOCHWq
wMkDwhPpI5eoC2W0Oiz/pbF14HMWx3xCngiAe3yMzr0Tc54igM1xJbNWfY1BdStY
k5MqANmKrqdMcr00BsKvV8XHp8IDdE7c1ccicDsF9jyjipVkeVpaAZJKjG+UNfsT
GvjF3uS1lhnCmCv5iqaAl3FQFd2NJhyEKjT5EqF7EI+N0Z1jum3sLcluK5HsyL8l
cW36nAgtYH/efTWfep1s9FUagcXTwthi7xM0KJIUM9Oo5rp4vu9hV+A5buU7Nfl/
pB9FrGk6S976a4IKMtWyjZhj8SuwLh7GszjvF3xIZ99K3E1UKNrp51c036wSzhB8
BDNx0P0JouVtC/9bHJyypEWQA4p6sjqTADbJJfNxNVyjc6A+kgxibFYzSvuRi3RT
MbU4WJXwuJ3celnzokavPnb/dobBN9Bn6eI8jtDrvrIrxqLtTrX7l9ONWUI//igU
eMso+vGKfY0JWtP15gx/5XqZUXirBBhdqByh3kbJDHjSSTA5rWOKCxCLKds+NegL
Lr73tL3q797g1IdNpEaqH7XkV0XVY1Q88NdZwd/rxijTvjNRWEtJn4eTkuML37NM
OrctqSQn9ejaxohKg3/tGXO98cUteUjoD2mMDrK8HaAha0c67gbw6OxS364iwthK
VrlFseWdLCTZUGWl9xwZcs9US6Z5wbIxIoOLSpCAExaIfAJqc9oyuPaQLKA34axJ
4rvUgu+xZpx4WTV2Qw37gBawrh+uTXtMPz1aoOPEwnj7OPf43ljSOy0ecRC+Ruii
Fyn5CPpekfoB9C1hWqF13ScLclWE16qS4jUYkKL5zP1ieN+3KecqAuZF/e4VEaU6
eSoDUGrw9gQUiwiYCAUJqDcMasCM9TsMUwiWAT2vFEuQUDnIQw1+wSBfP+6X6qm0
Mhxjz4++RkGocCr50gZStoT0ZAd17KEho8WArYLuG0thJSmc7KUDmCDYt3wWx5pc
X663MsuyrMkpw34A8T/WS9KS2EG7B82k5WqDGjebkzsr/ZP+LlbXRYVXp8B4CV5N
HSzGus4mO//he6mcRQ7qCa8v1KvXCTHsfXjjffcAUU6QD1znz66TOJQAKf+Xt5XP
Wyzt5ozXd96lnfdLJ1k1Rtwhg1pH8iJYLm2ijYt4cpJzaNsU4d8qL/NkZJ22ojcE
6PT7/1HpGDGlh6vJawAaWrHbWxDZZhuuCNLe7MdVlaAdibJzhQ/snPay2gKfNrTs
0AJ49fhdlUpudRXa2598Co0FSrE7VpfSIg5QX5lyJuVAS3NIeZfgQMfavDW+dwzW
2XATRqE2DRuTptJqVPVpvptpMDQ/IVfalr1GMJVPjzWdcz2aWrBORCqKj0U4ax6v
/gmFyqEnIjEQY/a14oMG65y4J9cKCNq1SlEddeRGadObQAeUB84TdN6MHQtoWRP8
vI+w4sWVcqJN3WQNvaQIH2GyMAJLUOdG8159xCKnM2/vKo1WCLTYS+dMQK3VGWgB
u7vM6cJWPRUH/H74WhYsjAuL7Tl9Tak1BDXk0B1CRWZP8Spd2F0Mc5tDxGcljC92
KvvL9V3iIAMawGj3/QuKlkCeZdYulfzq3BF9yEP8dVj2FJDarLeYkle/ej7XIOSm
DMQ2J9MJJ9nalQoRU0OuF0SXstyfOSjMP3+OKWovsP02+NzvmDzj+ynDcmcbCj6W
diOqmtMAsPa04B52FJyFNW9CHjUGA6ZQHp6BmYQBSHWLlPtqlKt2xA78Bh4wZ7XS
HfPLC4CZkCP8VI5IkgXwWfviddVXvCqcxj3CfZsXcYMgl6v4gQo8lcjP5WSAB8Pd
AQt6uln/xoVMmbURGPYzJAZ0fwPDyffUvAWdaRIvkA8g8QMvvWzj2fK47oWPnrL3
ZU+p7cOLiwGwVZi6H/bH/v7PcJHwwqPGwyOY5pf2TuckwFSHIyWz6OCnNIPIuIyB
Yj3LPO4Up7XI2QfYoL+9LwzfLcVCNWXvaDaaCEE58NJIk34BW+7/KPGEBRhKXPqr
FfszDn5bNiAAbmKvNctTg6MWynaCS7T7WsUsifC/8Xy8SF5d6X839DiXq0yOKomU
bdHgWxHg7HAJXqj4QFdXWCUcd+cmPZyJsFmZ5fehRvDxyUgmA2XIxZEwSqiE5Ii5
PTArT49tYO+rrsqpLK8BQh5Xs90tV9Wk/96Z4959VoZGHRz3M4xmhJtSvPywu63r
cjIW6x5SAbSLdlpnGSatgMvEGVLKpJvUhi598zCFVfXkcKGGvlFAZJ2PofxdqUA1
xD20oa8SNutn89ZqNG6azrX2swk0iqWnjuoAY9xDixYvDrLQ2zoO/nVdo8SPrv2L
Wc0LbVrq98UVzoN0RWPqiV25SJqh1PgMXe2Yj2H5bMkhEjIHdcaHy8voAaTIMBgS
3k1Ao7dBnQv5tXvoG24eX2i8eRL7h7k+00m8j7r8541/cP0QB98He7/vsRDL+VuI
C0NecJV0zAtEciwlcDTMbZs5ux4jTuO6G22QR4zgpOHlguqmT5WtmeIogIXca9+8
gBTFBp0sA9MNwqn8iBBWNz8BRgqb65560pcL1fzzW414ldTkx6yBcCn0FG/71cTP
HbvARVEaBydVQGI8D+v7tUvYFk69eb00MMP7pI9r9M57BA5NbmttSTBRzghGyiha
dRPbYokb3Okd5txlU2AocuOp9yEb0O1tckCTw8C0tsIZ40Ak1ChZZ6Bq/hezldtu
tISvDBK+08Q5T9yMnae00FzBgA1SotzOtrTUycSJlbxiKe7kVdj4iQ2PKl1IOthN
sb2TUnm6Th1vVnXNLrlSJUl/c0P8q8a8rtJCx0AR+AjGZ55RL4kbcx6R5e4EXr55
VguCnxt8XdWQ1LYICYGAI64OsLW02ZQSWjDjyfip7Psr2fS0Ehjd5FjT4Bxd7gAx
Nv8XGGzBDjMScEskvVi7QtAkW+xmlUPZnPa/debF1Iez4vVZQ82cLSIXqdlNjW+Y
pWAd4uO/q6xuNCUSqVXcreZ/hHPN6iXYzCY3kA42XD+wkiqFYKprh7V3i2fde789
hRS9wRIsBOgGSstMbgQxeboMeeOi8hyIji1bu7r5pZaXXhF8ISKoG/IA/8Bq6uit
zBEBkIJNC5Rd4ILMXKZNW9Y8oR8ckLY56/DpDj+dyK9ucsv+IriFw8hC+nwmrZg+
wQOew4CSfGhbaBQMFLgRJm4AXiIfoy5syCPiG0hPK5NopVHdDvY4rh0BFjZXp3kR
qQK8nrbHf4jU5de7rC8U3eMQ6wvS2gM9cjgtF91tJxvb+z8vqfO7yqZGznXZgJz9
AT6MVd3O8UD3E5gX59pL+k/U3uNoGGIc6BjRB72OnVkFfGkcX6xZbq36Mfn9UEKZ
YfVqevG+CBwuaAhEt4vV/lQ9/fCx3BRAr90CGGRGLsZhq/PZjWPAmkEg8nfDEZ3Y
mwGvh1R+ROSnpLPPD8pX3YX5TpoFzrCGKVdPVlmRy1RynyPsh6W8MD3jmUQte9MP
o7YcL7ZbDrQjwOPyUQMWjVBre90vR/t+1zK2PX1zVQH2cS+eNpabKEbvpWYEetdw
bWDUVBy0a5tjdI876wL5V3UZaQ4Z+5Z5Z0WHWlqMSQB7Eir7iXFq+CzugMPdo89v
Chmlc6D3OKUiqd4bJk3EULTTPRD/b+9uUEoPNk9jfph1R+61ceIfeP4saROW/Bc8
ICQMoxW8y6+qaIMuW6EwQzMkR3/5eqKefCBmxEQEE5out1RTt8aemsxIDw6E2iip
u1GfdGJ+EQqVWqONkpc4pEtgrDBJxTUpiXjyPDujHOpbjQwbSqeYQUNYScPBNbwp
bwnDrTWunB5R8GKOAQaugtgnvPaYTZisLRlt02xlkJ9Z+8cIb3lsHxgJ1fT/+iar
vuiv2v5T0wx3aM7lgJTvNpXPj7cSAytFPameH70pK5iBzxB5LumqgSXaAQGvTLRJ
x7DpSOhb5gmRRBjMCeFpzdT51i+/rmN0oZun7sCq1TkIm2bOuOvPAsKpQF+3CDjA
3CrXJagWUoLe3Y/DoJsmzl7QiWwftkYnjGIMDmjruCr9TMwvcaNGgqtLuxydzL7N
b0kVQw09BUxP9bUYCMpPrVjdTHhKLhwdqqMA7/HGZGDHlZuHMk/Pf8ptdbWLR/Xz
2boLBnA/nlRXYGqTTfosIF+eY9BKXKkogIkRBCZp6cksR6HmMTa1CIM7aFRmtA4R
kJ56ca7ORCE73FbphPYeCrpoLi+CU33iosaw6g8iRV4+XYcxFzpHK5pFqgG4B6YT
LX0pIRn3vs7Lj+WCR2PpjvPZmboHPk3wmjlfru6Cs3JCF3t7r9IhryQ1BX9RAAtZ
cRxBNZuFeWlxJN67XuwoB5/mZ0F9bL+E8RgyS0fGP4dybagfcs+dlfPY5ZrSN2aX
TWqMSWPMW88R9znZpWESVuSSNkekbXNfM5RG2PqXJ7pe0zniR1WvfFJF8Y1uDk/M
HYex7NGJmM5mfHVbBGiuTwhmOWHaacJJmVEfMJnLZiiBpjLmzBECraLkbomc4Ne+
W8A6aRr+eHJ63LoBWDt6wu2Lp94Av6u1XzqZdEY/ZjAeCydEVO2OGfvPjSIpgFSv
YNvOlQmUnBvo4M1Agz3Vm3pjcEdoex3aiSZDLOtPugkgWQi/fRHsVjTqq5gx+IlI
1LEP012Nvoavu6LHEdTpPEdJWCcq2CUNkIuZb4vA4/WjUXD1n1fUVsczcKMcLQoA
s1jTjfBjZgHxoN8jgIFElDtqt8ILyA3mkgm8ZkVhdHdlRDLnVaWVARNnK2q+7E8D
kfAQSBthI+0rLRA1qQg7CUMc8C/w150yhbZBJ/jKoYFedciXdeO2jkY8RgF8aIKI
fP26oz4GYC5MwfPLHQimYXnmmWcSaek/wme/SiuHyEXFXv9+kwTMIdYzbG+0aY1Y
3S/ebLCdA4Go8z4tKuGZLriWt9FDjC0tmDEbUOHb2/Cq67vQxNhStB2y78XhgYjq
FZSR79ItEf7Ha4yNgFocR8KxqL8LBbwz93EzmPgAL4ERCiGbtwEOPygkEalqeAUs
jOR1XcggToQGqNfIk0xZMrTCL9NA2erd7t5A/8U3Dk9GpY6K716GJtnUD/aO8U4V
EpZRuipDWDWiBiZsnDCR2MUIc07DB+MTwtHjg44UROJAkQCocxKyIcNsjbFqmyO/
Ua/0sl6OOiEkPpIXGyS2gcRY+oLFTYcbcppEVUT7dof/Cf99cWn/GKECVc1L2gnz
Uz66KHL4RRxUtHh4TMzUwjzGhq+i7lfIJZTG92XGnpNtD+KDEQQ6240IkdAQVIhm
b8JP+MKM/dyEJ/VHYPmsLPmWQ41a8W8xvSoKFgIoRY4tiK/eji3IXhmWLJ0pnfa6
XTzMCxMYxIN11UwbxsSk9+T+8JRjEiN6U8jPKIGU7xj7JthA3KsZBT2wUjP8845U
OVZlGOYzSDzWu2atSecMBXZHYqjqMFOALlRs7wAR3t24Rk656MHpghGVbFeZpheV
TPrcYvhnjNPve4GyT+qi25xaqnOsPbyOdyFqW/uHDSE2rlb/GM3uNvJTDW2LkMjq
1jR81jG15uYVO3Rws8/A8KLlI57bD5IPNAMCpAyhY1y1dVqoODWsKnqXSKtYY/j2
OFq1bDq3YZpJTz6g/OwsrKwDgTe+mDJ4Z7Y80eJ7RiYolzuf+EWuMUe30HDLJgOF
9n5IRn7aMbY/UMllzjYYIAbFCekNL8fPu1k+ohK9GDEemMsMcgwxSXcQnGTVAH9M
7puhMvDp9zsj9g2QxraTXVIG+7uTcpp1gY5rsY8JVKd4uQ59Lsf6TeFi7WwHcgIz
avcp39G7w1gEkUnIih+HML2YUpexIRGzCfF44N8q9beRLw7tvFYOgNIMp7jGB5U3
Yo96P7bLDVn4Y1pccs9FYiUItTqOAWtJ2+FeUe+/VUXZnWiz3F7H0zj218BXF+Km
ZB4rgBK9qqtxs9xg8jP0rjb8C1Y+Dy8DvElNi+rsAerhv5yPi9GkfZselTfeA/3U
NYFGmG8mRAA/zhmphJYrZKL0zQWaKNX7dhM1O5ZD9xorzaZ1Obf2fE+E9PzqasZA
RsOmrbOl14mtPTim4I/nk7WH3ZUdomWq5IW1lJwJlJzp1TaEGlP1jGF0vhQP2WHJ
93biF+eGTocFszGSebTQ1HnEYPXOjBjTgtV9QlHf2r3buhqp6lxBXTsvrXuZTDZM
FX4dJY9QvWyd8asRHQ+1vTnptz/aI7DGtbx+YClo/N3yK7At5xce3QKcYaZ2XPxQ
0SOx7d9g0nTjnABuqOWF0l9nOyDBuocLmW2jy9Ab0zGo2JEZ0hDcBnYVUGpufQC4
t2wgW5UaN85vLezZua2TTNZCeUABRqU4ZBu1/GeiYZtnhYipW1XSgxyB8Ar2TIsL
jJ+wKXHOtLUONPZl2Ojkd/5qy0Pc7JM13nw1Fo3IuMJOcD/2vE9Tok9Jcg15uRJb
TyPylkHh+cdmicXOj8xezTXTiS05M2GAgJQjicGQ/XVKU1sAcsUPk1RSbxx+V0hq
KtYTaHGYQav44bgRVb1kI3Q5TIRrhpQ/RCqNGL9DWvoXu+LxJwXrK+mkf78o/ynB
Y2YMkcXj3AHccSWlLC5trQDWoPpOwefWWMforM/XG4u0ooNA6ZfKeC6jbpl/fKse
SBVtgIHjdUwp/hCictu+KiDP5Sc6KGVT8UQZoLasintGzdSrTZspyysEEP9Vrpmp
T5iiBm4H8bIi94q/o+Dz1JlMOPcH4iNjni+jhlxgE28dp5hXgaaSQzf7M4HmkFAG
cKR3Bw4IU7Xntvi8olohhxkxGDbVfUnWUyulpP9WGAYKHcaWtaAzxO2YQFN8o4TR
eQzlW4aEpQpa1HhWLF8wUf1BtbXKEDmGrZ5otxyYIwnW0MPtqe2qfO0ZJ875zxR8
d1pu4AdPeZE1+46GXKubD5HUvgpoLz9f8HjVNazLRm8W790i65PUaK+6BJHehX2Y
gecMhTWX8HXj/kXAqH7TdEhIuyVZiSlvpWC6nmqN4XXScBJTZ/V2fEU1wJOYlWIt
tBdCvoL+9c4LVMRc1O6oqy69M2uw9/N3eBnuTNNFWiJi12VGTlzYL6CLOl/y3p0d
+olGWEh/fu4MXQObo3CMmNwrcfLxpEv8s7Wb66b6T0M+2+FcyUNSOeWCI0HwvRqJ
tAw38C2JDRrBNQleHw8Co274BaYqRjsHy8A6CG5MgM31cQq2ooo6breUKe5yhszB
TBMTovx6ctyfdIPfHkGzLPfpKGuS92ozpv5EGZZ6dqLy5/GP0eOzSGClVMqDU+73
5fYyr1qkHHpVGst7tzp3Q4lB/uqZSsu2S5h80gSHXUY=
`protect END_PROTECTED
