`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MC2QADYvbwBdRxJkGFYF8qoZxrR27CPSHvy5xSiHaEAu2u0lVLHKoRs3jypwu+M8
O1jmqyHqe0mk6fLQXYlqw7cw1afqttwcw68Z0fO6qEqzmptbma5NJIqSe0g+0IMa
lq4Lu1uJvLSjCFjvIielPpwbSySes7EEHeDnz7c+Bf+bkWy1ypYntKmJWeBXL7BU
ptQsyitHVs4jCrUMPEblFrukt9rpwTgP2cN7Ns7LDG+aZ3E5aAPQ5xNdS1czjWqv
ASveZSFcSASzcWgxYv3xcPXLznZJkuiQyMvvFPYBA1EDtRTVkFVERyePbZM8XSFd
fQZ4eU2EbqmIY3Uqx+ze5Y8KX8JkzfBHO+Elx7YCKCgqCOBaUhMc8FB+ICMBCu2k
HF0gCaeulGNbT8iaf6DNg3OK+mWor2dmjVWZ/H25AZwqS838umxfYCUj9Ray3sPm
WUugQM5KaO7NRQcndI7Bzryg8iV2Cuqq4PsObxQ7OGD0Gi85hDIvrwqEN62ooYH3
Sl9tQxx89i5hvx9J2UnDGd+Q98YtrAXL7T1KtXExPKUPCCvspF1h6wLzihXOwNY0
ITVU8AENW2+M95kmyKSDM28fdfDvuoFSvEfWoecHIW6btMPpeCI59PzBGjRY1U+O
HZkfuYY6tc0vnFzx7VZNkGzORIl6uk2ZWtSrSL3kh66FaojiH333O7FTzMckfofF
4v5DRxyXD+pPs1+CV1qNpnYkRHLc4ZYf5edHnZoz3hVdy691sCYp+wGc1ZGdr9UM
nlll3qjmF+UwyRLxAEIeUGq/KM+M7IDFUBITx+DoRMR1p4H9VEmb7vdRFsV3ZtaX
ly9sxa+SFA8wbkLd/6T7U9L6yvEtQ0HzQLJtBGV64xmYzxlq0efvyjNMjzMMn1ml
VRUaOBxILwI/+fr6OsZvJzXwp+2ZCqq0eaTQ1qRWy6X4k4MawjbcGMeTFjXCO0b+
KPVVnEl/54FqkFZB7s4j+OObzslgPNV1pceCer01+fZlazRQL/ykXNSq8TfzH+a0
4dZ9Fd5tH66UlcxceEv+uCLF7zeeLH0l8OPDevUYdCbGXSLPpJnrL+Yku2P9YcIE
/j2h2x1ut3Gc2bZUErgEumN8HF/3GJxfq//F6bNSPWKuxbgElFkeVHgE69WMtUFp
7az6+s4j5AYkEJauFHNBf15XUUhfboS2QEcb3Lt4OBBslyC2V2kfLWGN+7KvOyCq
xY7CIRrSWvczkIpbq4UQzc5w82TJenecKA7YrFnOPspadsZEBf3WI97N00o9LjJr
gQgc9tF0+8ZZi2iLhUXurLqA6FBMJfJjsAQKZlDMkb/WkB/YDVtXPRFHpC0Ve+a0
RvXr97q5GH0uzHm2VhCyUvIpWQEUb2LPOOCHRmcM43txMaiBOjaiwlAhwB7WeOh5
FD9/jV9nuIZDhYVXn/CFAbFpMh7r6+GL6Hdtq8MJNF8CUhg/DqFOmzybxYc1ibsC
I/Y1Qeu0MKZkF9JG4cRrfw==
`protect END_PROTECTED
