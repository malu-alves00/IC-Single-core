`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TYRhpr/7EB1MdKHXTI4P2W0EVQUyM3pGx69n2TrNg/DW/KBSoJxzTGm5eGqSppcr
fKo+RV04zKLNxQyxc64DquPRXnu1mhj50OOqN+dMYbNoRow+Tw/Zb7wiYMltBNaz
XEnkes+F10e9v690mS+3/kbNLs28HX1n7ae9FoH+ZrdCVtsN6dn2Wt0nes8j14Ir
pxS8YIF0KsdPTMI+I4B6SiRTULDhhf8AXanNHsiffV72iKzC0loQvA1cZcNLKlOW
pUpJc+QWlthQHmQi73GbmWCkmMbvKnZGZPmnjtbeNunKwzPd8VepsaglQr9/W35P
EQNrRUVS/OP88hCs17LKEvxw3t/q22GOJiD8eV6/vpmgr5MyRcVX6PCyqM+uIrWL
xeeNQ+BZMJpbploIBKcObR+x4vFX2kEszWsDZN1b+TJhoFRUH75uhd7noeQZYiWD
GqrBiZyqjOOdRLQfOartf5wj0POPa5m6zuksfHg8koE=
`protect END_PROTECTED
