`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dwjMKHsKHfwKzhunLmxjXRV4voVn3F/k6NPtrF7p15vuAxxrSRUAYI7cP7di017v
TXVAG3z4DCGzFNdp9kRJahUVaFN4vwHb/Dm2QlScBxtqKToyA29hBQMzgi+r/XHs
DYun5ta8Ok17kv+bSadblI0apSEijjFsPUXdyq2sb+HtM634zgyV5Or2GNcu73Nu
S9ljfSjNTZq5v33Wc9yu5MV8HDx5eLLNnPVGfCXGRF5tGXv8YqtXflpOo+i9mr8t
U/u+zlzDyagirdEQYYgiY9MOzaaOd59NkXD5kErQOmK7QI4y9M5etayzBD+wBF4e
qUhHWCxrtqFe7b4566LfYjxWIni73DrjykPvH0ZnY6z4xvG38S/OPGk2634Hw5Xk
Ks3N0q5e4mPQV8ZHCvadhQeaogtAjCdqxaqtWjj19UUfpiPqVOooVF6R3p1Kqoxx
Np8nmYJkycQJX606ToUbJBVrGM4AVC38kZ6R76ATa6hsYjd7F29Doz8ykCUVcSJs
EUP92R4jiA/if75yJNB98ejm+tC/iPGphA79mIsODwBgNqeg9NES/ON9R9lFJ6Sp
nWQ1j1PYjQiycumpKNqOHV1FD1W9itrZ3bxl079agQOgGEBjX+f44sTaPHJRpL0T
aMKQOUTXnOc7eSCyeZmjX72Ij43cdzBdb8ySE396CQhNsc9Ol6VWPBH8BzuwLYjq
0AOregq69mnLAtB3WV4fKk/YaQT1C3qZBAyhdgktAQhRjc84hDb+tw86sqTGjCt9
S0iJRBrcxX/+333PT9YYJWiFL6RVgge7SgS4fHrztspHZ7p/O+sNVHguPJo0dNKL
+uq9gKIVB+4JjSEsCaBBrs8Cs5JvT9cUZI0UaJYQsC5dOFxObpAg5VPYn26kzliC
ncU1pHsw27dgCUxdDUIdb8SpULlFT4D69G1B6z4ude1p8gYC1AGtE2hjYEgu7piB
CBd5zzgWMgIeMMC61jIiR5Kg0t2d9+ABef0buvD92Tr8Y+ssORTmB2MiwbLx+MPN
gaMXtQcIWacVDz/oOIyFtSv8Or1QDxI0kfCGCDwgYhDfYNKsKcQSZ348Kx1MzGDJ
efsjOKaji23zNGkEsqbl5d7Cwvw5ogbitP7vqDaA326li7v9K2qB3XUQwwJ1N1PX
M3V4nFLV8GHB6XcYZ6CRbx9YD+srkyYwqbmS3lQRRCcdwg+MwMnrBCyhkHScL5lV
5yDaXNnEYlzkS5fK2TXhVwYyg1FsocqTxQ4n/snno1oK78SFqIZbHq3nTAbzql8X
D3zBD4vMxeYUiVEeHN+81siJ2kChFRdh1jLbC0Ypwqot8WwLIuyEB1VK+++4Onsw
0ditWebcLlWztfyCyDBQ4LWKXQM8ffGT8EDQw+9UumhNRDffRl7W7D2l54gk+pV9
xkl2QMyuByjuUMT+tFskD1S8aefZbadmRoBKhR7QHLOEYU8KKTzHLF8AiAStWcfu
yug4onluaqk/hyEXZbNFpRJS5QMQlljqVFyr7661J5Q4iQ4Snq+pSI+JrtJbSUAb
x82Ra1L5s16kb2t4E5fdpTZfP0cGJKsfR4O6llPAk/70HYYFh+MwtJJRDBOBUH0C
J9ML7QzkeWYRBEkLTPKV0X5D/LGHir23z7zCArXbrzEH4kBArbjvanuYh2Kwap/s
n7cOBjqw+BNJEfiZlu4ZVU0kRqHGXw2rscdRFInPfxXduXHB+BTS+AXfHriJ0Kvq
uPjQRZ8bC+KOa7Eu+tHBZAPqrcmJnb2mhLSVs7JK6t1jTGD/OuZhvGK4u2iADMeA
mbt3xzKkrTOaeoqYsOg75zg5tslZfmC9vGex3MNV/cxnX+5ZjjumU7CrQeLrfi9V
Sqbs8ttBgH1zbcNq0ksqCkxiW/sfwp/kVQuFpQfI6sNPUXKwceuhzglXTKhxphIA
zYwJrOgFEX3nRKTxpmWPy7GtxPbKZ2Gi4dLP7PtnzyIVFcuXKZfHxefERJW3cbN6
wxwYPzCujAnbpQo5q1e7C0hCj56KSlWS17EbmmsUOr5IURaebteAXiWuSKyG/zbR
SwAkq6aM/JUmmQnnAjJojO8g0eJVy6+HCzEjDvSu9IS1FIMosNTbQbZxNQFWfbCf
zn5Tpiq08c+SjTcPaB5jVO5TMvFcZKgki82pOakMpwWdb+ux9v8yIpbngOd7zkzk
+kg6ji0p/nw73tY+jigzPsIS5Uxh2UlrxzxnIq7hp/ZgB9YFCtx1C9QWNsfgObx6
0AXqbTI6fCP+jdU/Q/o9So6yLHx3dJ+utVAkEbAUTMWU35DRauXf0MVPbCYHXN9w
ycT3E9CExT7uPKYJzrhe2nM7GzaGAMeJ3puySaPl7CIAMSVOFN6TCYoAZ+wncbHL
jQIDuEIA9WBWwICOxv36xdV8YtQLJMTbmxAaN2w5Z2mtSiQ21Vhc2Ck5vmIME1Xw
AqP52JtN8Cy9UDwaJu+ZyGNADcp9wVaJ22xXXukfVSV0zDSJzNTVZnfSh1Hj7cZX
qgV1knnOKAnih7huNCDcMp0p4Xb0JPkzmvb7UsY8eNiS2N2Wfmr4P7kX+/s5B8Sl
RviI90yHHR6tBjdzBovf1J8TumlufvVkAwtk9HQyZB8FxfyfVQ0ogTseWSUnhax3
twTYysQyquZEeni287penYtAQ3ksnLrUQe9AnSYl7gQvm3uNAfukl2fPcmqcydgZ
k9739zgTh8dEf1HS5aBYLfOK+SfOWUbpRQwjfl/RkP5zaS8I2sypoVgLvh7Vu7S3
jicZeqG9o97LEPdUvGKeXuNsCzAsZIKKYv16H+sa+DHjUIfekochGtw2CWNjCliY
+gFpHcdWUQRXz39PRWxGA9fSbX/Vn94CPz9AJqVB1dEpUbqlijQF/7tCGM6KKSfW
7wQhz19MZC42rArjnW1/2MiFjr/L2Q6gBzfnTxK+QyhBukgy5Gpq4Sth2qH4FmK2
qy0yrEDRkhYEQYPPJh2535LKohPPz7foJO/tQUzi1+YS3YzZGP1HPIYFnKUbA3kc
uSoowzfJOygBPPUGzO753F4/+cwljp8ysVcVEOn9SEr5pCI8lh14hCukXPv1BEMl
BK8qL/fsAnzZAAY5DxGUnci4GS9QdXpXLoZ+VczelLFqS4xgVNzK4JWjZIx3WnPM
B+A3H9i8ZA3u6cv57YmgcjYdYIScJSXsdRZLUTy0r/QJkJIcWOJIf+M2gtOXKELX
8Fko0Dw3vc/tX5ZaqydsM68FEIW4ayQmHKItkhD6DJMjgwGCwZlTyayLsXtKbSAC
mVCFPgrC4f3BQOiW2pJ8sjcfJCUdJ/XmnzeyV/3T/q9ZqpX3Qxiqa4Dm5mEbNv5y
YAf+hJ/JWAVytFhIVwa2uucbsM5AieYW0JXJh9mpeqz9/6P6BBiJZI2iXpnR9VQy
sqNivx7kWxUlggNslEetDO/bJH1t0HBfC6ndY9S/nA7xLjxWEHC8rDm/nkOr6OPw
JGSMLBBHf2oWsS9NZlDvfFvyI9TbGuSzsjfHixayJ1gpQU9Gew5x1bRPv2tZTYxL
emrjPw0CujHUhz6hIJsXoMF2kvtlRhqbGFPhFYfB7XyYAir5QrV02BUJjLSTJmIM
/63PeRrdy5en3K+6dq+QRx2iD72r/4JgLPglirl8d5fwNBUTonYBKGjkKGvPNINp
CucwuTzXp/wSqy9DLpr/zQ0YJnv+zyN8P43FPDSo82f6LAu9zzfkO/Hd9ASbG5mD
dKE2ULvKBPqxB7zwFmrxazXXJVAtwnfLLqhp89C3QN2cofAj3NjsyGRnEz81KGYJ
UXPvxXI23twzLYJlxa448gIldCJLGd3Sl8NCai4/2nc6zyzPO/QQtzLCOTDyO14r
xYRjSfXEJKZo2GPMpsKpH6RYKaDTI6ReNis/i8Va098QxQqP1JBHZENZZCGHZNAS
/XGr7HyjQuKbD2kKgKeNi7Hsnpohd5IntLVGh68tYzalCLu0WFbJEFPM3pVgrvLG
kxozMPGegeeSj+fDhsV0MYAvfPO0wecbQ8t245200l1Bn2iBpEyv75WYqwtGO+8n
cWZHMLtN3q/siYcJgyswsp+YNG8EYhfpiPAqTXNOu2H+72IabqirBgbDuvSpZpsP
iBhqvOaotDf0F/K+ebiJFeaa5HHY51lCuSCKx9ZXg7WGHYQpgXSLlwFaBkGUghyD
TfLzHPTl9e0Z/jHTvFGfbO/pG4KWot84NnDNoLudo2tCCx6yKb99XNOVlFtJtHDS
P+nNqgq+uvqG5n7BKy4lJ+TH02+uc5B4jSbC4qIDJdSLr/3jooFCaLVbCxK/aRFu
6Rx45KwxA/b+ufSpu1XWp2D8mEQY7r8c3wrYEqSATIU6AwNQ9pAgdogb7PcHQyoW
JAWocQbwWGihWuoRclLzCl1xScvfrZUbpqkhg7H6AmV3NZQ9jZ76njy98XpdmB2K
toU+9Q0r1wILumE6aeGsQflWH0fIJx3kfKttsuBUtGRsm6B89Hh1hu4azFDgsdIb
z8Yk+1G9skhvNzHs1ESqnNDG66jbx5A39BUL0Oy1ee+jEElJZKYKF5F2J908/HiL
/UGXckUP+Es4LIqiZ9vDfocNKq2rPUk8W5DL6j+qOoZr+YcCniqSbZWLVyWLYg92
vCM+hyBTEwvdNcwPfv4Sc2qngQYCNXENqi/toFBQur/bV7fsyEiV4DwRdDTso3DV
Pk+XdrxneXlcN6IvVI0JyIgmXt7fHsu9Y16ys4jFK+Agm/0ajsrSaL4IvqddvxcF
uPmfTsvH7Kqvo1xyIEDsXOki9m/MlnigLRZlZmCatQ1Dkk4ttfd0R0oWg5FXtd/2
aOoXGHyX3dkNcTOlzSRvyDsYGH4hevESS71hB4eDzFFLQ/Gs1ujLlJrq2d66Xtm0
fPpKcHS+RiDIJwzTpLzQu37CRlvTPwfx0pNTXBXOP9gg1zKS9WNYPKax/F4c9Nbw
V7gH6glUkAHWtbyjz0f/G7MYAKLaz8eaevjv+qhTA7JNTp3SBjt9RLZH/kMeaTwu
BaIoUyJvifnTmUIky4goA6UVE5TiW9Sr/zA2x1aIxx4AtLjte0FkD1M5qMTSVeGV
5V5taPjTk9nXPM2S10RncsjwcoYjHgaHyNxxjoCS1Nxo0GAi1lOwhLPM5kWzuUsh
zX75tQw4KIxAgOIABVQCHvahU7bZMvR+Pt0EA5iOqsjvK7FpeQNdFfE96+DGwWCj
loLPV1q6GRw3kO8+tKPhD3vpRtyPk0Ee7IMiwibjY8gwT457zCZmDsxaRLu53FBT
YchELjZYjSUqbc45oiq6bG8xUT5154x2ZGBAwGswCXKM0pc99SWcLGNJ/QiN7Z6H
EsHYs2m4oxyb871Nk/HnLoQkk7f5TLoLHpk3gUI0E+fc4dR2mvBAlv1PYQkwK02e
nZE8L1ITyiCBmXkT4+WhvnW8KTtUHNA6F6oR2D0f5Fpa4iF3FlPG+di19yyHyCCM
/h/x/I+fbW+rFZ4RspgU/LaAH1RhFcyVNdvsCCZW4xhitTDAQnp6y2+Mkd4+KcU2
MJT6ZbPkccNbBiINTmJEsfJSDocTfPPjGb1BMIQmyms3i9K3CrH/IGaEr5EJsc+Q
IWOqDBz6727Opcm4jJXiwAhsdRUqUGQGWx2NMv21jlpLS63BJLI2ZWg6YMNZyVuu
t/ADGgULGFiYZh3wV89fk+noHqEopEJL2QBewyzEdxqQ4r/5UKJNT3Tqof0tdjTo
OmXbjW1Qpk4ZAJpMpVlDii52afiQ7tgwZP1UiUqMaUgnx/NVP+Kd8SQC5Zqf2BJp
FlC8EuqVU17kdBhH89i3bwFhEM48DSWNmROv80JL08nkGnDGg8KJ/lCPsVXnSbVx
uoBxXFVjHQOi4Hg3FRnvVIbTcY4EbgOJeqis+2vsBbG9tOX394FHShPPmy/BpvSy
evv0xbO0Px27QdlYuRI1qLcPeOzLMnUzGK+PSH8WzLzxvxL7ugFmyIjEWQGZQ+GL
QM2n0Qg4LQlrBlZt05avPHpZVAqQvD91XtoMS31HRixzP5x6DAejqEVOTKJ4tdio
YU+SOikboMEjGjNZaaxUd/AbZbvGhP1kFzUQJItdj2jzKyizkA6KuEh+3lSp1729
1hTJ9yiyKzkcsWICinSZa1iOgdP5OW4npgB9QdqNibSZosy+bI7ly9cRE5JL/Jlb
+/l4WKw8pn/SWgKek+qUlHY1zoh6gYR6/okCO90pLN5g6KC4YNTNHZVTy3U2iwqh
qp5IMAFl79/sQVsoGsH/3NMQc4rB+AK4/ppjEwDzxrvuu3Pb6XWDeFkMACkSGmpg
fqyuG3l7Q5C8KHfOUB7OqY81fQYO/CDXAx0qn+lVVc8uUNPIRBmjRM84r6bS8F5c
Ew/pDD19YBpsSBI47SSVPoVRzCqXo/p82xEarFoBwU3UAXkrna8R5C5jBjkdXCp6
qBRxZ7vEge9ziQ/RzVgjY/6PhEbDuS/VDPGz9MMgXxGh9YXJXkn4I6bofm5H/Kad
68t2BopRiihEw00wADt6ddBggZMY2+C07yuAgWmYpwGpytgqY4o90TTwH+BR0Zcq
A+1a49q/QsZ6YWSZb/J3xAmoB5YgoeN1ooupZh/xE775yILS6worjIzEhJE4O1/J
N8+MTTul6Gr0tOmFu36SV1hEz0z4rODrBT9f3uRdoY4IsZb5asuxCey/JHB5QsF4
4J01f7LEbfWBDobxfG2NAHHIqRzF6CBXBdk/j0VSZSY0A3uxXiSGMdBiwBzCKdbl
8VTMw3z82cwLh1pHpSH5eGceVzP58jkYlHtmWKijhHgAY9fDUp52kZdrddccwvCp
Qx/mG5+gCaaVEjDevPBz3qpwiA08NTPJsmu2+cGBl4G5KMHlQSxX4oBjDD7x1l0r
EPVMGbSeFHVHckD3tSb1IfOO9nO1X6rF8ydAPWMDF7ABVAOYoGIMzGq//OTsmGIm
plsiZtCDlLqO3oPEFdCoXB2amn8GAJV3E+B7dlm4af3IuoT8pOWQKQUTsUUVhqCR
+VNLcr3NQSe8qv19x52VQZI+EGn/TH8/RXvqv/9ivCEzzPB8bv2UtgYk6aBJIce2
Yp6MlzSVkr3PiKwTOE8OCwuc3cjmI4WfyDQUXXE/DTMDcVLJPt9CjT9ZGUcTxBXO
vlyU4N5vFOORr9hKL1EDSYkHiILnBHXHAnMVrggsoC7HH7wnKcwE6oj8iE8mW1/9
bk7CWvR5zc743nb++j/ZyNZN86x1u51KoqVN3rCTYbcdhopwGbQwq2gm91C+T6NA
B1Ga8UqHzwnX0T/pdplEP3UiNeF2hyBBZdh3GXaGNgKoE3Ka7lVzSBrZEibC835A
LR7inuzaspaLNgsDlBJ8Hvli3OEFste6vGioRCUaQRLRetjBnnNlHA13x32DQF85
M5ijHEi86N4krSTp4p3QSo9/c0z0rjTiu3Ng6WnqQa2BLmzUCjinCeoQpvQWjUFk
nkuXavw75In+m2Lit+5Q9U3u+nXzvAwRfa8Z1jVG3il6D/sPLlSDEFG4tZOyli+y
WDWJp5w9eNqbjyZN3ct/iQfyGDkGNlT6+wSksKoGvN6KUZFNufjCjWVJRbHe5fXf
7Bdzcg0mmMCJKrhggRMYK5VUKBkDsubikH2U1C5sBMEz+RDfqchLWUfEvoW71F9U
hX0hrg9DmqTM6GaDEIKMPJeF4vOpwYCNOsWrKE5XLUOwdd6dQjGD5ICDsghT+/DT
LqDlATKvCwgIAL3j6IFZUjv0QcxGL8EZGJchOLtmPtpboiEYW2EBV65ER6+QdJiH
n5873KfmSy5giS3GC/LUF+Cb5fPZGTWK+g0jmWcpagrXz3p94Fxu8Y728WD5LCsp
rONVM9JmsRKunGMqz+xdHODEopL6ibMFXFjlm8FIPY9R25ryeWJ9nJrweiEcu7vk
mxy6UkcLGg41bAs5nlFf802FOiz0a0jezNIVN8pCC/Nvphy8NAuP1V/fvFJyUoFS
k339sDiKRngutofuwaFsIv//+RzC0VRXndUqeWJ3BpweBro861kBOIMS+86A5XvR
9UZdd8n2Omty1jYr638x6asfnHSa8JiChQMv6Utr6hCN2BBBRdmIGsanCorls3eE
X+DX0t9Os8M3Sq7kafG3eZ7wz5VccUBSGM5EedHn/dlpRSOZsiuOgG5/d0ap3uLv
93gpahG3sBehBVOOBW6xNjEo4WqTEm99w748PJ6VsFOQyDoAQhO8xZx0Gu1bUIVs
PLZb03pKxIex+rtHolxQZ1E5DpWE5Ilxx3extF/truhDBqndRAnOXd0uLIv0daHP
ZpK6YwYx8ZeFCCY89+FtbqKYezd2h9Uy3JTnK8onbyo50iHdaGBgy3pRDrpndgqh
dNqtvxmI+EV6+0viZz1p0fQPWr0oxXju0mwwf3xJ8SVPegJ1/21YM7xhwdX+RvFF
DuAtnL+rNOV//jjulk6/wiBorHvNzkdeFbGoCPKBCh9435SlNqjzy/+t9Avy8+h3
GxnpibNG2XwAoSY7oCeCZsrVlZ9JB8DVcK0zRMS2SfbGyV17amYqzTG4kj9JqcnE
stCkyjFhRTf+etNkFnsdMCznIX0unwPT8IkzUhNDo6aSEQu0yFXhrwHZB4v6pm5T
09OJzTGC2FZ9IV6l9s4Drmp/NUFzunAKvCuQO5ZaUtQQcWHiMOZRO7PZUIecX5We
fAujMd2nMMUSJ/E78NUOc0Z3TG0Kb6C0P6qdqYlWgyPmp2ltatpl9C6bg1V4nKzL
26J/83MlyoGkF+Aj/6+SzUkqyCrh4Piybqfyz4V3I8JrYARY71k6ljePv1dFAghK
v2jJ+3nNUDKHJVeT1K77XcF/2G8m01Dww8/L3wfw8cNRmcbTDoRp0lvhlTszeIpJ
If8QaAd5xyjMAlym3uaGpP7Q8TChcaVi0r0Ql4PDaCwigBfhbNgZwqIKXjpZOf+E
ePf84wyC2UBe/nhv+QXOmMObZYeF8TPfCJ5/eSoxGYOArDEX5E2zEnZoBjleUPwP
hPvv325LY9KDIEBGMvTN4L0tQndvnaAnHJRCEP7EviBFQsfeqU68SA48Ij1FVYnx
hnryLNBXKZVBBuZboqzbJno7GgeOdi7Ua8OMRVhnUAQaiRbQJLWEMxe4oquhZBHy
tukFYGn3IAoQcGQyQ0S4Kw/OxZ7ilhwbBFCIuZuwgrbMeuFL6VLABYB0DZ8rpA2u
GJF9oAJ0RpvZ9pVyAE5msxOJFF75D53b2mQvsMe59m0Mu3gR+lMHNG4J1SXyFtVn
YJxwM2gD342uTKm1lhwvWS0KKTSbUZz2+gyt+oNPi2BmMVCj631CbhzDi7hG38cA
oFEKijVNw52tu36QZD3Y+7m+AaS8tL6Tf93gtvT+8vC9i6I8OaXSB1mmOkrS5vI+
XpoqFZTWzOQ/sBLPz3XKe/KW+BrJmdJHP7KTBLw+fdW+Y3qPB2ENkfbmck1mYlrB
IvwOypioA/PVdhsVeAOLauTz5BQQCwfZFf4em+QWcklQir8SKow2bh1sZwHX4zhx
RskkFuR6aUv7XQGhoI1Zr1J6RYb3Ev3mlifOtazhbocLU8ATlx1UqhOTyQqqnz5U
fAlWekeXsVAQHjYaHsoat99qLmhFjSNgie+DWCAfCs3RhBmiev2Nq9Ce921mMKoe
Svbj0Yy4sH51UG00/D5yb3raYIv8GyFcAqaEUQZzy32RBxT1iATzRtTR6ZJs+wMy
xEg3CYtx13XOyDsLEiwsyrz6UE8tWMnm1MobxlOUfYEt29htq4e5vT4YOFC83e2k
JYgchxU7su1YopQMYM6IyBd4xBRS5oDLkjEMsdWiLjZi2fjFcweGUh1bDle0cPKN
y8C0VYG4mjicSzHswqjwiB7cGPGOCmCiZFE0DotahFWZxBc/0UgAJADApva3sbLF
eaQUHFb0Rm7chj2B+5HiAxWpfehkU2bucQTFuhsaiw8y65wSNvMvs8mz/XHbr9+s
Q6yzNbilG1IqRCLNtEYd5+kw0vtbrv92YpQZQh727m0qUqQ/GX2b/g7KurJ2pZBo
i7UAX12UqYQIFZKmCR0uZzdF2Mi6G6himq1Rd5a7hrTTlO84Zgv6591oz/xmsu3u
hpSuWcs/ivRyXHrXqBoaAtEPh3j1IfBgjQ5QI0KS9GsEXisX9kIjTaGw9Ni8cU47
6BcpwTULE/7CiFTMV8CFtFg9lA5HUX0Q1pCaBwBDrWuTha2PtyOH3eIKdp+zKQRc
0pDFAfkHqvzz48AJ71SFgIbz/tqJIOm+MiGJ6avqN7USjGXUUNiVUWZsmJFkVidn
fD5fkIGUbcmVSy0HYugbNA2iyjh2LC6PjfnRTlr5nids17hpn1JfmgaPsMuzgWXW
+Z9A3+d19rQTpU0SwIFJKoFiraoybipdn/RuBPGvX+3NwDmm/BDaRsShnRrsHgi/
nFWJRtahUHlVuliz6o71pV/M0uZAXxIFf8Y57NQw6ainAylSbeDix8sjK6X48sGQ
8+qI4il+/S9QIXHLVqDzZCCdHFPoUaHUi2JGMYr9gMEEXbdU3goHryvp14FLyqPh
xGBI0VDMKI5uca+/jQ2GiNznrqaqYXLqEzmLRoLSShoYDdYuDsFoM7jhZt7RxKAm
i119xh7cI3iRB3XPGOWqUCD4GMYrJ2h3U+hWi3ZdrRL7lxCoocFJO/BJZ+qnQons
wlkiGfb7cT3rC4ZIIcjU8oZaPD/Rxy9GGJsF7ap9Sl7UcI+9KLXqwX6FPQVJpBAh
CXOBNeD0TAIBZrdn2x6OjquNnFZ4Y0sXVu5UjeWf8A0jf6wNLbPBUP1vXYdyP66Q
xxw7KCVMNSk0YIBhDKAsSQKQiKARqVVhFPwspJHMe2CCbPPVNJ92rccTLUEbAWOE
MfipFuh9MH645RH7gfr7WnkUhxrlmUX03yPYo+AhMrQqt87a5KGyM/bSC36MmYXp
4o3q0fwOYP9nMo2jXcFISCFFhxPDJzIs7RPrlt+6ObyvC+AepcTwUysYtxamFMpN
/qjADsihrJZQgFJK3JWmToOu3I/D0K19l/KJkJnkgH8ovXj2+C6xq6ztA8rMdMyx
xFM1auP1qfAzgA75E6mgjCAWXXZNTuOpeGWGjs/HOP7h8+66lVVoijjc0b/o87Bv
40X8uX0N1s2GQUkA/w94n9+JTJgQ8Tw9rOUSXuCbYytXQRLIQAh9m1vZF9GwX5dl
dtSlFgXf5+dp3q0ugjNfewp8Q9yN+dBSjI+vfCybvv1B+LIo0DhvgJS2VjsPo8Lg
el3ZQjhEVzL0wSsdRAC8u4EmPp0W9IxdUZGyZtqwfBKi+lsP1mjXl+uJ+xVaAyMg
M/2OOEHi4bJ86HaZHkuVPo+bbMpuikK92iyf6l4dLJvH361izazy89JNYIQu1Yng
RZ0bBEb80eMR9o5q5R0SeubrhdsK9jSQqzAf9ouY1GlsbcSvSVl5wzytySxzC+6Z
iZeJuSlFbo7g93AiUAQK1UM77tVF9mOe3ZGHHBWymJ3W6jAUDDUnZ/tQBZAYrBoF
r9cxrioFcmOHsHwB2zf9k1vsJh4veD2XUvgA2BgAN4UPvWHE9FaDv8mUntmf2pCJ
am1FvUsuchhdzZakwMeIc6PPRZ0wzBVRiJxnom5aVCoOOQyVah6HYedckVpLVgUQ
e7CJMWevBgRN3HntPthib+9bRgcPoRSaCk/eW5eolYL+s/RVDrhPUd+cxydt7Wah
jHRZXf3Ct2ZCAe39zbVJq966zbl41M9qVfsTRegyqBPFiG6+yDdGpaNIlarL93Zh
I49eunCR38OCnMIA6xRhwYZiZ5mvm6oOxlmibiHt6yH5sA1EdcHnfq/AGXEgYrCm
m17SHwjkzW2V5t1sFkxBRgwEVKThHwjN80+sNb3bjaq9Q6HfC5z+tegSRQSK1GPG
hNe00s+m/l8nvJd1oieKvVXsdLNVAs0kAS7ncj0bViGaQtze+g713WJwlZ26s9Kn
6GUWy4CaOtCrX49C5FTeKfnf0lJ2hV7kKmLODNJievlhL2XSzXSg1OQfIhMEUpwM
XefxtEaxK3nrRM60Dm5syoByi/MKCVLv019v1+uAq5/s0tYJLoP3fl5titeDTaUg
LV9nmkFdAe/cvM/3GYuNmh00om4l2ofKP5q0Y07MjKsJS7LbrfYcKGYIMDlFjSG+
nJb1Aq58jvv/WxBN5iD8jKXKtKhrl4DRZlwawhpyDIOk9/HIqTzItjxTCgiymXVC
PybQ1HVgFxbn1a4MtFOs+LAkFzlhlZoL4UnixY4/mEkJ1j1RXoaPSzupFslo33r8
SF5hOAHAcAg04TPRMcnDbdBJMxQxURrT+2p/1VJGQi2eOfDWJ8w/WJyFIFC7+1/S
o3T5YZo0QXmzpKGtH/sPH9sRqcbp0PDF1q2De/5sTDK39WrXYZmHfRI3Iq0Da/bB
Q96y4QJEWyP1ZsSH6AKuZ1ZNt3jWknXr4iez6aBTUSKEve5RqwN4xFjcjh5+ryDc
t5pJhluLcq3zIAFaI3EOF1PJPcE0uuddCwBJMyqnFyCI336SpgTXzUTd0w2uVuya
+102j2Hz5JQWXlL57Bg2ZeCShY7R11SIVCnCJmcLwuNk6oHlyLER2o7ISiHPlWVE
cvi5j3RkxVicYumvRBquYP8B9Ho6TEuOyXj8hrqPbz9/QE108W0oNqE6abdL2wDR
eDdAfqSbVo7iPDtPAmQenTWDG9vPeVcuS33iCkjgnFQg1Ltlvi5EoFJdOT3uURoO
Q9Rw/DJStQ7K7aCHoI7NIIYrkt6hj2BJasHb75vtA8FL4r7scHsRRWcF9d8i2EHN
5weLXvlTLKB+CBdwWwT0NqsVcIwZu6pmx21VGzY14+kNjtIaczVhuohCHG9P50gu
cWfhzcPZvDZnkUvuk43fMCH2AUIlqJk/EjLcDps8jLRJKatmcG1Ju9PPmOrb6rnW
xggTn4VEXQ2NM2hEQkPz5fvZvhbBqau1HI3JNwM9QpSvWpsVfeG0mgBG9SNxWxi2
YD1EnUJzmHHd/A8ixgwlvmDMKCUTz7VDmZBKBZ8hKPSsJU+oGgI3GSIHai/VTp66
IOWfLZmy9xBkbhIJ22DyJRgSF1xULeR9TSel4OXc/t510HJ5QH1UkdwQjowEdF7t
EG21ZliKLkL06rjVzUhjUJfpRPLucdcGIHvaSHfCHSOCTETDBC0fnKwsXDc6q014
YTG58E2lMOdURyyjecE0Bg69hS3oeFnOBBf2Bqw83Mg4h3fj2/zTn7ft/X8D8goG
cffSf3vLDrEQT5CJJMug1riFCh+bmz4RnBiZeSaZbaV+HjOjOgPunyXrXWTpfhdU
aKr71IAEih/ViAmg9NaWk9cF6rZf2w/kqIANFlfnrF3Pmbe6LM4yw7a2rhUxaN0B
UVFWU8qPhJnnrNfk+O0fa8gnv18evcq9rpZ6uXriK449w+NBjSk5PV1HbvYZ1bhB
7LMIoXaq8gsFDS8hYvmxTY3bJr8AbMs0Y8IjSj6EH22OfQye4cPZHrHoBVr5uBUa
Tam+pm6kI+nV1XUUh2AeeKxDqoLZTOaPJETZ6gL1IENtJSRn2ton9FDoqejUdYc3
Dl6KxjUMs1CrL5Kj/SnIWrFbVLNrCH+sjg2FOOuMV6+r7Wyw+1FAQMOJiXJHueEG
aHHPEyK+RV6y4Or+ro9oPCJoM5B9w3R3ppneZaIsSGWPj/3poOcIhheUcJKOOZcS
BGyYWt8YIfS75wAubp3VY6Lrb4ZcyZcG0wLTWfuKrpeygIYH2AqMuKp0MpI7P8ey
Ze80XKDLZAHm7ZedGxob0ZmDjzaOlF6XTaGPcdvgFMN5B8So5A0iVrskYNWz/Yr/
znUEBm3m2+h4NCsGA1QPXgNYk98lTfAl/2jCfulIcaCNmFJnXWvlBFZjeJ4HHY74
kIDIFviKY5H6XFOBfv5zG6dIrQFo+jPs+DsmX1MSWYgIHQofX1OlyAwApoVIJmBL
W0sTbDPibNPfEaXVlVt41Nq9wDmy9YifK1OTk5N4Pt6pKzRibnUKdpO3hs0i+hS/
aw68IwaYbxUGb9/XDYnsHmNRA5zBAm4LZVsdsG975UvgmM89zcIVbLe186mck6r+
+JBavjGwuLAQyKUTg9N6v1U7NqJwP1G4Xne5tOqGSBCnVZgS+xZYosEHjG4Yyvhy
XT1/MyrYhaCNisQTTrvbt9mNFEIRhKt5HgWSink3zH1KqBdzIASNwid5F+YPjWBf
RPHYb1XBrcztdCNV1IoODastJkSlEG338Txc4ahWqUDOXkhPi/JYGITsSlTlPK1+
KKuJGXSTLN1kCtj07qHSAR9ltqWSYDQSbF7rLpbzoFtNfGeNjZuZUWqY7zMfClbS
FX/kW+n/jCATe47VAbq59h/3ytWdfgqWICeFo3xGA+BOF83tGj9WxUQ4odgMlpd6
8eRZsojORU6QadkQ/WTw0KT76YPMVq0xHQX2blLPY35KjkJo04XmEVT9DqNXgyR+
we+U9YvVqzcXWEAjON3Z7z1KwzFecKoPZfkyYLAXSn+0b4cAzI2BC+E16AwyOIpt
Noyp6Zp0sjkpe7b3mtuhhHE7JpBN2myL9BgsimnRjsrSIm5sVhC4tMXU3QdV6vBo
DSv/rwhvYIae5Fqcue89C91d2Aq7JJx6PJXWDBnc5blOBJe2fqt2dZ7BPES9PIMw
rpvWn2A/9DvYQPO5Lza3wKbc8wQ96f9V22Di2R/E/GlERuQkjKue5ShXdx7ENUb+
Kw1ZzLQnCW9I1KBQZ7LUOfdYQmrxE8KjdetPOclmIZlCIOUCbxPZHX6yFSfKFITX
IIZWH4WqNhLdSKDd8kyt9Pb2rCAz8Kbqo+JZ+Gicqb0G+7moErZl6CktcyhaIbX1
OLSJmeoBlKMeGJOJgZ67dSxrMPw5ZTBjRH0CMXYKx8LdouTU0v6lQ7N2XRnYwFkK
nRh0QvHl+TM7FVdChumAxul0XZgxObuqQR3s/SKaNYpuMJA9clMpwOdt8LkrBA3H
vsOr4WAeDH0Qo6IQ6zAJty/aa3IEnXhng5JyXS8jVg0E4NJbki28FliSh6bvXGmu
FBHTiCxS6zFf4fm9H03acIolLtuGd2xOG3Xj7zdu1HWP0F29cyxAY6azqeapbAiv
GDHi5QaoVMYiKsdF+C42Nyb1YyzlO1ZfOwo9R2xAExR4Ix9jgClJxN4TC/7K290i
PKIMb4JHGQFah72562ihi/9p31giovgjojGeTZk/QllrJO/kl4zlkKAESZrpFyrq
PjHQPPQIsUAP85Vd8Yij/p9596kwM79zxvnMEF7A3TZuABkcCsKxQlAIJ521fq7A
2MF+SCPXnhmlDFlaHvgCFJCI34FBsFyFvb1wbdXjdUdrbBfgghwxBlx/L3+cUPWK
VScxUY56sPYlAC3AnlMUq9ZDFBmhoohdd/c64lujociE9DcXzALSqOYCYr2Q/f5B
VVWEK0F2CIKrRsKhxq6SUrzOrX0I4d+XwN/AxvecLzOTGfN/SEoRzChh4ebWwxoz
h1eeZUvC0aFXqinjNC5XssuW7CBWd9+ZJuah4Dmejlf0WqdTvetmHdO5tbj7lfh5
9e89vi1tAIALM3Yc6zsv6MVnhVbkkxsp6xYLf8HagB/7eCiWTXMeP7ZheOYDBY4a
7ol0khWIGeGYXKn9XyF1zKbi80VYOz0NZprY7DFyfl3LxSX+uPdr1U+wGtRjTTLf
gZ8p8tv4BrzH7s2FDcD/s9C/Xy1Tq78UM1lKVg01HrSm9AJpXBqV60QZnLviEtN2
AljidFcCrdhOVjLg7iyGaC5YxfpK6SR2Iifxzwy8CBrD/o8vyT26oscRU0VxZSUg
eQyx02KR7Cs110ng4HuunpJpjYQTPhScsUB/9iwtdDggoUVvDLASEa/j8QTxMNTS
LppBA8auBFusBmEFUqAc8OwJfVaUwwWPnRFGF8YhsPuqCRf23k+LsYiIDL285Lj4
u+QWH1nuA8EM6l57R/T6Q4I4VM58pdShn2UEzvEBe7tPSzpQg4OTvaDaxF+wZTvA
P25I6e6nLT30W8ax4DVJFkGlgMlOpjzUhbQnNxVxTyvLFHqAguvSFAGTmDOhc2qY
jAtdwQjVxHtSiVYmXwz5rW3svtKPmsmQGsr0M9cEf0jsjKBsOmClFZJ/zve+s5ma
VxlbQY5EnQEUWEok0Qmx7h9J2ccsV3EfrgZG9M1tLdymnjyDjCNn5h7qWDpgBQnh
WivJMEutSnAqwefG8lJEFG7XpZYtPzia7VycwZtkEyqImOM+qFYD+CYOOe8muQjM
8jE4qtsCJ7nW4gPUUeGHQjVor1rQFSdiRPyxDHWNu7q5FpFb5it/VOqT+9pLQ4Ab
jkbpTtj+/s8AlEJxhBVfu55Az+uWwDpP+5iULpJCHbfz93f0yw7u87LBlTwsqZ72
N6VoKuCNZEY4o/5OnnEMbJFBrvZLOlrpU5nEqNqoCS52KqEylSv7RNwD+M0kRHCe
AIeRTPqJNrw1AQStLQGcPLSzvSIoEZIydAaG8dy0PbK+sQhIsVvL8Pg6Oxyo0KMR
j7Yy3e8RKJyBzJlLjqQjNv/zmJ14HRCPh0JByFrYhPQ7KizoENUY/kgyaMg5QNEN
RYDGBFqm3DZOCDU0X9SZqz2shvB9Uwconyu1V2/X3lTkYZ1d+q+DdSnGXIFXDS+s
WVRWz2C3K6VQ+daxVZSSyy0036+esVfzGaC11i3lUnzA2pt0KE9Cy8jAcI6Oj8Uw
OBR4YP/XuWlOlMBn3tynQ7PEv8PItevlKl3XsoerbJZ5DYxk6S8V3rcB+9w9Jdu8
rkpGeNg1D4fMFHZQG1pJGUCA0ONxoFBPPFKhu7/DkP6huIf38kWsUgN13CV85ljA
bTrepizBvmDzzoVlmm5j2Dh+weCU2YLpFh5JvVtdkFVImWGd/l+E4GC714yLSc33
Kyz0sSicPbkExo2RQjq/JJRZpvGeLsDg/mWdRlHLySFp5/RO8utNdSnSYfCOu61K
gh3P7c451qytKQgrBi5mhkGAGR1kIUAJVGxp/gKzJnLH80UhMWeJCH7b96kTOUg5
AVeVjTwsNB+6+Fu5sXKAMh+vXganPjxGfwJpnsBhuM0PYcM+qQUybZmAOdI+JpkO
4mL8IKTiG2S1n0xyXt2B0ExUyWAhXa3F6BGTw9CrS08Ah3Uv12erI5ty0xkisLs+
wG/Cexs7DB/5VlGOpmliVAXXAYsMBg/W22h2jBwoJzrbc9+8bNjI9tB42SOOKR9O
ewYgppWZUE+GLZqRgiRJqMohyZYewj4Shw8VamP9r92eVexpJBfHLmX4af9EI/DF
PjVgs+zd/PFKMV9O9aa9WWof/me5svTtXp6hiLWgfTQ3rdkvUOaeF2RPtfrNQlf/
Ms+2pq+Bljgjhm5Nle7/a0XEyLTGHa6acPsy9eRqQI11xOp1QUB4k3cZiLDXkYa1
BqMxT6loGucgwIo4I2oeqgLbITyROi+yO//LpxuymIJeNWfcbVxBtAx4diNmLLLT
zqWIZk1vdMwUhXn6HBWVUE4YhBlbwU/prJeXlEt9VYf2AjiWR9MF9AwEQJiPQSqM
Vdb/JtwGFeLE0U0esf0LaqJuaZjrFIlBGZPtgBXLVY757ce5r5RJgoCTZNmHn2ah
uQfxlU8qPhkbB+BzzOnGYI+1ca44NDzjXajASSQJWfHxlgavRtZFMbQKSddN3U7r
3uHOhMX0O0idUZ6iwuRzIEixY+NWWDnk1hWJgGGuavYOemK6b2qu+CQbzE1RF/kR
WDgXeyFe7mzq3Vndx3fxjg6xv9M27eo/v+Ll8e0G5ge3EjNp/nhTp1Tmi5r1LUWT
YBblFiCXp9JczfsmneYOTFNDfPVsUvu7CJ/+LoeeVXIiOpAlKVjebimN+l5ZDiVG
ywZ3XrUm6AvyCJqfVQI61K/ge2/cSFAazU60MW3GUir7GUVk0QzLfIolNCjYjTyZ
Krqn8ALSFXom4lgQ2+kzYYTjbf6rAXRNFRKCwZjd8bSGIlSCtXTAYNmDv/vXaeNs
W1yEWB/OhgFOaDYiwS7bfdwSbA0hy/MEFj3rWn6cRpJLVorQ9oHYyRethNp4ENME
yThVbynw/LSpqp4/Dbw/MfUDFzQImhGjTngMPSNh97adYsjABcLefsuG1DSxzHaY
a3i1/Go5WhYOsvMag1cx++sPiGGmXW5DDG9KiJ0/GR/4SdtCJe6rXfE5YjIkaEmb
86Y6FBkIhfaJdtLXbEmvMlJQhiPIBKQnVGyezu68Waew3Jat10ldxrckjYawnkKp
Nn0JGizxjBhWpdHIRRb24JQkZtDPXvYdBoJ2ucpB/+9IM8iOY+px65iC9JkvK++1
/pnn/5Fn0vcYOI8ZT1vCU1VetYVC/49dpDbDHsdQdP2/2rSM/0KYcKc3rHzLJv+j
8UZ1u8077Pza1YCj7KCm9h08SbOqE8hbtCTfq9Qr/16Bu9UjqzV3mVr99eSke6bg
eJOej6wgQf9fzgjHC0Q9b9wvP7MeCljHII110Ea3J96eoXbCWzz6uXP/PYxgiWCs
/suzwpmTWkig/h0XqzOdd22SF8gaGMKTxzhZezgUL2hneJJMfj2dZUn9W0qwofgv
ShzfBoKNbjxrWIi0CvgX4AB42fcQ5z2AUL8WdYXpTCT0ylM1EM3NLccDK0lx95wR
mcsUtUS7ywVj1Eyh/myj/Wt65ASYQ8KUHUXnF0QRAYKAeRt666gTI413sL4pMdfI
RpDR1ss7Ggl1ObWHYthYx1rtHm1mTQUYxDXmhW+8ZsqaZZoEFIGjjRc8xE7dFDeB
0Ybe5107OO5kq7eJLccxq6YmAlFkLciK8PNN/f+D6CZYeHkM+/j/XtItO7UheaYD
4UyMyLxncQ2GP16o5rVN7NgqvJIIEZgXuzXc0lddU9xfisE8Eol5UT60EAb4d4wR
tePxFZ57mEAtGYHBcCrj5Uon1ivdXC2OsJ8d0J5FapK6AULo1zQzzVdCqpIg0hzd
1m2HBl8sCnoLnMXSf/o/nC6ybSfFMSNXbgL/xIKwZg5JEFMfZ0i4AkDhEArjV+Wv
rknqg7P8GAZygA7N0XL7xpGy3x0oc8Q5Z2g+HMTwBvsWC4zp+yi/MUjaYv9O1QH5
BFh35E3hMN8cJquqKv98kZlbvOvFLu5VzlkyUqPrmzbl0v+RM2RQepGSLg9ha/wC
fdppxavbnlXl5042Q5TWI+RZykOM++FWSubQ55nUAQAvBdNzS/e6H86HheyXjRov
ey2D/EIJ8u8V6cGgkiQj7yyZP8A6GsItMtooid2kzDu6BAXlt08zU8SsBbjsDRcg
FUxXuq2w4Bg82m25N2+D4inC2JFUeZ4wh/NML9RYyG16J+RMLE/mz/AVf1yFcH3M
PDChDl0iZnwUdcIDLdzUs5jyA8xdNfIPQdHGKPWkEs9Ti3XPB+aiT9ezOS6kwkXV
GNEDLJRoMWsVW+E9Y9K6inWKy/Fc2NxgTMsHHrp/jckaYZWpP0Ef2u1rzVSQzck0
PH95SEQmAMSNdjlclYxOsivBumJVhZ5iks5/1geWxo8CffC876kXp2/E3gaEjKwy
+aPA7n85FvQ1k7niUHpGd2rP8qi1vDHL93l8Y4Fn41cemKa0wcWZ8YwK04Rooh44
QvCwADNqKds/Lc7rvBGFJzvAE59naQVm+wGz6svHjF0puU91dmZz5ClWuBIfkemp
TizXCHo7578OC7uWRLC2inFbvRQ8g4T/GCkrPzzVsSZXMeBPSnunSqrivx5hwpmS
IjR7ffGWXo08oJxK556SV06FNHfNzsSvyk5kteDwzAHck3D26+6524NDJQChvbMH
2wd+eaX/qJ0jJMRWeiCHzsv8Fb64DSoGctRPY5YSEGf3LuqMwvADhTzajIpzuZbT
FRgqvuu3ltdMglc/9h2xoV9GPVBinjVRqXER0MjS9Xoi9gEKiWUdt7oLjywAtKEQ
h7QVz7o0Tv+XsHAuOrHOVR7T0kb3guZ0XENH94N2hcuZF1caoGF5tdCkoe8X5+q+
WeVnBvld9+v7lKhiLCJZbv1exRlDlkZMwhOPqcVskPqQyN/qrBv0Xozg2/U+RknT
NEJF6+Xbjslhptef2k+YuFo9Agkh2o/JDbE3RfSlcraRhAqZYB8eyV+9jREjpbyJ
f4GLF0PJqEEzZyX5Ae+QW5wIuSCurE9HTg7IBMQAlvgDw54wwNmB7KtqtEYXDPCv
BYGg2mRet+tffvtwIDuZVjRwTpCKgVmJFoRoE7GN5+dicfz9NR4zdfQN8vccMQyK
3r9btt0f54jGf3b080ZglPcwDAePunilS/VzgMmz1lh7F8wiUmT5g4F4DlrLRbYL
ThtCA2y+ut55vtdhtitQiEQ7J5qZ1DSuJipSaWR0WxfzV0F3LjBuTb7JBdND7yPB
wwqOsuiIgokd6ClXyu2Z86JrNhdRFW65fdVSb5t/yeHtZTFjquBZo7mC9iuCHb1M
P8pK7zuJd3PqakW9PgoDBHxdrkcPR6CSIs3h1y0UxxZ5S7K6xnnaS+61fmmEzHWw
x4SS8oNvUwDxAxgIyQNt6kEvhp49g1/+TTzLtW1zdWI/5/uRHPVjwtPTlI4KnS5e
VSQo+mqyurAnEazFZE2zEE2Ssr1ZQNiFsGreUTBFdeQdqXVlhdaZQOZJ5ainTLgv
ww953En194OdlFUZWzPYWocjPtzscvFDIfUfSyEu3nF8ac3t9vzARi4R2Liuzjp7
hQAqkgIyoA0E+9Dct8SJU6qarKH2z9tH5TAab5DsofM91MHIiAewDHFctskeHUg6
NM2PnsWrPQiBBXyEAUCfAOuwNU0whBrbNcXFzpx5LR1oNzFmgNAhKrIFmbH5dtLc
sbZwdBGAK6CfyJaF3fIWE0DxFjBI30Gt1MRNVmrKbHOYidESXMtIUB4/HVV7Tgp9
yr4Uy0F5SThyCFkfaoiZYEB26MxS3yMB/U71YkC7beNhM/zlPQ2WZIGbt1yeWi/Z
U1oLsDJAiFND6yz4rPby7LsGFoc1pJO8jrs1X3M0D7X2zEHGzbJtCKc8zl9tP3bR
vr9d05iJJ2LlQXb/Svyu7lofAeWH/32pRNqOZqElAkcxVFey1NVUMMJIckMZY801
I4yPRDc8f5ISAgoJXdum3D/fu89YPj79ZfZ2tC2qtzN8Nwj3hrwvzg/I9oWUJcLS
/zRS/QW7z7wJU9nxuHF9M+lB8GWvQmHYqPXbaAja/hlNSxsvpGxKGQ3yT0+foRoQ
nr4Ux3u2gZKPI/71SauFWFfCS5JVHjatnJg+yrD5Gl1H5cbsHU9x7QTbVWs+rTZN
Yy+iEHmqbPtLo5bwmO5nK80cqTyGoDBeQ9+P90AFsrulFaMRp5EhKMKXxT2iBeNE
aKiZV7jYVxIlMHMDh0ZGzhp9ZXUJxIIJYwWUVV2d436Ec/z1YUx44GGnRSPv6alO
W0VbohCTBA2W+gGwmtEIlp8AIJcKamJ/LEi7J4yncvTxxlXbLNuzS7JW7tz186cq
Gkib3Qtbh7lqfb1JrepCKOz+x7hMw60UPF2/nGjbU2lkpPA8m7Mf95CdduvsNhx6
5XrJHDQrUowP0FDfD2aOW+GLXnKC/nMXINkPsCtK4uSPOlY1uEaSnGtMKjWNk4NX
iETMeX5EUQxteSNnXSK39O8VDY2noc9VrH1z7cihijGhClKH4Ft7tb006wXjeHlG
tiFyalt+FKRx7AjP9SFazVyQiXGhokj3jeXn0elxdVrf6bR4mKB1XL3eQEmJO2LQ
SIVH0Dl7fqRVwt6uD6zErBGIjDPW6CA9v6X52+m6ifXCzpj4udnpZKPrVyvHfhQz
wgEBh+oobWQNfrXh25jpS9LBoNl2uPMD882Ez8KeamL6uKRB03vMEdyFwGDKf++n
NszzBge7EGeF8iJaY7nneA8xfdhxEpw9PGOGqEPYLpY/05bBT4OLcFtpdxacJ+nD
jwrqdoFg78Si1OlHwBonsNT8uEAgmoRz/YWdJb4hjuR1l+pyeUKHOUz2DOSjRlaG
gcWb569K28j2JSB4juCngYQOcKnl14hzUSd3WdadPZMJYRhs+x7sdgWiEJ1euuFR
pBNMAKReOOOJamBtouZQzWQFG1Nv0yBu3SCmlxRmzq1gQ+PJ2uf4l6t365zCBAQC
kPSxc+9bGZTRy4kj99OlOnpx3aMY1lsvmo27v7MP9yy/YAKIORQxwD4WGxSBHwL/
BCSYkCgftEQxVDO0lxgVDnmur49Tkj+rt+Psmd+cHhfkfjSs7WScDKTzE+R5D5Gk
16H7gGHmogKW1Um0hNVf6M/s54NqEthnn/tkFQGBzoO5MbUsNYOSXS7r4zDxxqxB
VqnhKidxpcd0SGWHWdmuBbeo3ONQYatevvpml5XyszLQc8UMSseq2lHh28wV4qCO
uGRMD3Ds+oM1yw9euWBGRbKKRqYV/vZIAzjRr/vdlUzbRLUts9Dhx2+SFTlQV3Bf
UUzw4dC6oQV0vyXDXnfoaJgDxtLr3UHtywl5DAVsOc3a4lP+WUui/y4e/brZMGn8
bkOdwvkYyRS9rKE8S4nZ+nFMbi0sTrdaXSzK92yV4S1JmSq7HotiRrN2ok2c0KyB
8k/ETmPZX2cf99DhmgJYDCVvLKc6qu/iE77tDFU+n7nQiPr+ZIRYPRwRUxDhEY8N
+Zwvt7XJa00D/PhyDqe+1vQdifcKyfqBlGqLqD3GfjddND8IjWuAv8+XebHQ+sxO
rrc8UbO19a5bGr2XNv05hpAxlUHAZIHcG044ktXuxVbFefUKKgBvSNQSKR3aaXt6
QOCZjm6a35YZ5BPyMBDacl74xtE2aQPYoEZURV62L4dsL+Ukh2S2CKjJU0UTqkLA
5MNyEL/HFUsXDccbSvWc/qzObfi5pdZbCuB241bikllEF8RvrbLp3NXpq8X2vop1
Vh2RfnTsmXr0wwl9ir/K/6/dmb4hBrULn80FgGb2nKakXpc0YiUVDOmnlSNRTZca
fD8iKs8oI58qmmzQOyFtWu5uEAbRwZzOcuTDD2rUTjaNj/fW9UzDKRrbjhNORasg
dnfbopnqlb8W6zss+juNMnN7QZqhCRsEaqZMK5oxehfqF06Oj6Qnwm+wQU2XZqdB
IjBVA0CXtQRlu/5Xo9N9ofnQRdXGIDVW+ispVIlaITPodu+ofGqU4N9s8775TG2Z
BqfjXMhsnvBhikSOnRdJmpAKjcWJBTk4CST2hu/0oFeSG5SV/A7xwi/VINZRoISl
3Qu5mZ8s5TBCTmjHTfQ8ZjTHA7nNtpoKXtaBDOEwH8kGYxnc/9D28Tf24+hEp8Rg
L5LuU/qHLFBWt61npB1ZJhfIc+PhKfqi8OdjpeEi2G5gqMRzya0xZcKi8vYa8D8G
qySddM+Igw5gdwzVe9Qdw19v68BihgfdXrr+HR6OvAwuTdQnVNqRPHFX7R0w/vGz
P4Rz5fZ6R2MKVWjD52R6vtrkIwoxKVPdIuziw0M8/iAms6Eqa8VPDenisfxxhPtf
Q8XCUaimz+9s9MbRxugTrBwbONbZKUIpjsYDjuvFOU1RVCWSFiUUweBW0hrB9I+i
TlqSnmDTkevs8OC/BKL0UYRuLNEe68ByzZg32Xb8Deb+ypLhoQq11HIwfMxrkFJ3
9hMc/a8LlRfU9KRNDEGLWqg5GcFxO91etgN6BDyjtCsNyH1ysEICIlEqWgfhM30D
aPND5I8D02qPq4MK8sivq/dVwERZDMTHPQGoa1lNdbTJnQn825xNjKkyyXcbjTxf
G+62JkumYJkVg1j2PEnYSgFK3N9+9ILTZSivJ7KNESh5mH4+pTcrpYzoiDdg8HGn
VDqXFEkcSXIRoNXTbyQYXJOVr4J+pzQIYejPgn5GDw9ppmBV4CdlhjH/r48LvUAM
NZMN5YCwMYKyzHxRBRejDEETUxFLeyFyVauKBZ/BzXgwH3n8KBiaNm0D37tJ/3jI
UBnE43rS7O91AnERb2iANdU1iXHLfdcgsYUHPyWlR7hApUgsVuPuIX9zuDJzpXZt
h3OX+penvQkCISrKftiP2f9Hz8kRZKylejf2kZksckKmOboBIymU5ydj9LPopNGr
S6bPtYuCtm/JJzVBmRxWUen161RNp82T/elW1IqnP246cxSfOAw7aiIH26NZZmAJ
lHT6mVkODkDDk28SdnjDmRwiJHpEn/TDHkRjaHzcEO9JaKnIIHHxoxtaRkUcrv4x
sdnhKlCOHeQzSeKMtwUBBhTMHsWMXN7cYZMasPdRc5R4cPXszIPfpgD+qD6LjM0V
9BEQ4yKu+0tXHm3NNdonE9sih2LEYuCVXnj0v+b+WpZ6Glmns8tcZlY6B433fL8i
doW1p2qEWqff7zPcGCi+uSh85jizrb6s5yIqUHGXA0iuuMvozAkR10M4pL9a9v7y
jjHVwJaF3Hh1QLXs5sh9ASbIJfxFMhGKxHfKaEJ2JFXg8L9Toh1XFDEAFVYSppuV
RQzJ7rs89YeEz2N9NZ5klW1GItYWdaqBBanmn3wZQTJ02r/+NcEcuiafQhtjFy7H
bHAESPvoYCXx+WYekWGi+XlmjovReA4qchPpifXYvmWYpVY/u6C2eFyFF5UIRs6e
YVaYYu7h2vCN4byr0DPlUWiltYiSEywdMReoLna7Z+/0JJy/qV3JNSqptAopgHxv
2emkRP/kw0877eotZ1h3tWNjCbm/CyTh/yB2qygFO2GpnsHNEi8ozIlpxd53+6kA
jRMOv+Ql81Gzo7M6A8XPSh3x6LXZv2o1aXkPh/9CnNRaskFzVHX3IjHlbkLAn7E6
x1iNsN5uysC8tcTQwRiffIPayfRhNFfG1l4Aduelq4cvxAp8trIKBx9/zH+pJOoJ
9XfONNuuWBGhcdBts4caTnc893U1Hp99ldFBcT+sWVMj2buQasR+E9RmkaHclkX0
AWeDIQMvNABGT3x3P/LcF0Li9ulscuW4+595/vLc7DfYSwQ4LDEteyAbKJKpbYZ5
u9wR0bjmEw4XZ/lzu7pIcWJf3peslS8VPxw/97GSLzXthFWxDjq4ZcjABSX2/Ess
WUUl0hGDgbIDNfNtlkR8Iiw+NDU1JngBpK5PGeemov7CB5Bn9gw8rO5Q9KJJdNJU
iqTEQn4/nunWv7l1WopzKw5j9JsSS88fRHHBAd9hagJXB0AADsyUWgyMtp2Qkmmd
PJRUvlesqv0OlHDw0mwnMMyPgdSyqWYLtNYb5ArC6WnLpjpFm8o8JhsfhbNQ8CGT
uJZX8U2+kObzhbYsHV6nCWj3BU9nxNFhes3TeHWajr5fSl7CnJZb1PdFt3I3qfcA
d5bIhE20GuHwtBNbbyxlLFsXAV9ZoMUYCxf+A7iiJ41NjXA8B8gD1begxMOXHLhb
VuHl897eKWd3Unm4gprDdCmiXukBuoX5Zi0HHb3C8QmFgEmccIIW3pL+iqEC4JEb
tzfxCxCZDCe0VPYNky0DOSfNVVdCBtYfZT1sGWrxJL0DtniSJLECMFCG3l+lsuxa
bNXOWHgd7J9prWblwedtCX0CZm6Halju52y6j0rwCyo80G2x5zf+hUTr5e69frv8
NJ0rbMk0lVCbkHXyMDRqwor30f1JggpJT4P+olV0cYM+y6dz6kqhYwVzeZl80PQM
3zSdi8NkrMYxRjUZEUx4hy3x86WiNFyXF3WHztV+qGYbafXbWTFgCmXQ1I8ZgWT7
VV+5s3vW2KxOSWe9YTTIzH+vQbVhDoHtraoXZfb+W9fCs9vdZL6I6S7rexaubLmj
rfEuMVR5lj36p/cTCEN85lyvRvQI785/+EYpvkupaG5oNiUYRk2591oUc+EvzYaC
M/3MuHb8L5VJc7LmkmfGqtD0CHu1BS4MbMURRti2oPSLLVHx442BrFyIGuBTiZHh
tZ9Eb2KOVeGJAdP4hLqslUN7iX6GqK8BKsqdXddIdIvQvMu/rWfQOhjJEA00y8q+
9pfBrpOiPQRXGiRaVSSs3Kut7tpMF0rrOIat9pKlyfFF5910OjU988yz8MUekUkb
kWCf0A4zTnPqZ8rDumnLatn5U0nHiFCr3WBKa5RirTL47zbsYT/ZA0ol4JIAC0vP
BsIwhk+VanXuNBg1xeQgnitpb01baiKgxjK1GGfoaYRbsULWG/TH+zhdg6Lupogd
PZbbudPi4g4Vnu5yZOZZBY8i31ZGlyseAzbmoBhZwDKgznDi/XxpG6Ae/5cTzM/U
MXC1oACtDl3GPdBFgXUBesw33nqqGGakDqZXYjlF09DDU8WY/U8cM3JKzZte/MU7
LGAxU+xtoThlAePAsOWFqaerpmUsSdiCy0xsLOq7s+8Uwfy2XPG5lQGc+33xjzXu
JwxRMRrxdJrJWrUXLsHmPJPrYWvHKetT0VZxqEpZFXkNjePuCc9ofA2EQKeIZAkk
Xh3qrpFDyRDgwaS8NnAtOIJfd1wGssXFjXklwHwxjgWIXkV6g2Vze4QgNBA0XZrj
z0Rr0DkmomAYmJvPoZJ5hwDmsEqzD4L/grUtt7mSbEsbplCkh6PSw8buloxKW5j/
9AK/8HWGGLugKikNAXnqWakziQZrO2BiklXPGhRuhMPFUyXtTM3qOTFsr/Axu19h
kMZRaHhiNQqiubr7pHR7EPoJU+ZWVEWyzLFNG7YDJWvfaITXtTtVaqnAXPHEi33t
UuhVOCFYGNbEPdt5GjFNkUhsOziaHfsdOZoCLERVcIkMluXphWnAbGr9QBs6lHwX
qQ+zyHDTl8fRDB7ol4FWoproUyUUyHdcE50wBkTSlOTcdn4iDyh8ldlH9/ozkH7z
eohW9XO0ssVJaku5GK6WVOJIc8DKuYCq8G3RgbPatCW9QSzUEtyyOvV/BRF1jIGg
Q/xpwsmusl4CSPKusZusdWKC121ZTTWZgGSl6y04pIz5a4fbQVGzOgQhRdDDMqQ0
7jRxY4ThUMDEpzqbDbMTYxSb4zpezBB73Up+qYdDM8F2G1eIAQtPFavnKksWn+eW
E3npD1UbaGSyMhHV79hnSCFKDJWYQdZOPLTQJP8Rjmevt2CgmacUEiPc5LVI5nk6
X05YH5UItABSp5JTV030yFA0bkhsuLnHRwUhwWlCnN0wNgXDoGpy6PwQFxVmcdRQ
2iJNby00PWNGZaKYxyEKeAMNtpEKihxh8a/TKMGVhKVWjzhNCk38McMbNILBxtCO
BWOgKMj1Oom0n0JCdi6q9o8LYLPytGf+fa/TtTBIBRZlV0AwwrgxT/tm/8gkkDaG
2ONmaDsPVuX0MeKYtZdJyBlgg/DZ4UJzry5YNyhNSSqSSjlqnHRjs/zRffJ4F4br
rqDEmBf2ySsxHLLJRc4ci6XxdJz+fPJcUnjm4wDkgPj7i6fEEhVBPllUOCbP0fR5
fNqW/Kq1hbho45kIhjtk7rv1tUHcIFnCN5RkbqsPidfTBy+mc/WblpO1rMS0UMCt
7Z/UDfDKs0m4YOMoYCmRAS40EP8LmadCIjrgCmM7qAlnJ2omjkbKWmLFvDMiwFYx
G/X+X+xgj2G+9fbFRNDdjgWsSt5dclyN7GA9F/o0BdxAi3lZo1xF/t7IXIRli6KP
WlJYk0urVD50jMV5yJwsema/jHoOkI2VIhFufsuJEYGZWSlXda68f0OQlNLl9LED
mV/BlidOt7Iu4U7vtwpFwmuXFIPjK2VnPN2MUR1TAv/jF//i6OIonYLYU/o0WaYA
oz7hwiNd27zyxYD1mJxEthYhp2W7UuWZjwJla0y6uGh6eBj0AjwReVSB7hWJi0ps
Dy5gL38OseMwCJ0oyJB2jbs8P8nEKYbdI0FL/3ru8SgZJp4AIbeGr99sDPsjbHAN
KzlGWHPF2ob3eyC55qiJq/jyf+Jzt+cDomNuDU5Ft1vQpklHLdGRjEuXWE9VryL/
7l9B+m9L0z22CG7TeX2K+/znrEmG+UfElP83rXVTrhz2Ab9xJLKAGHBjeJ3mBqHT
tpuf4aWVA5193WvwXYCzE/ofukrlf1Lre1xEIG7ZqXg3zxbU5dUbXdme9e7GnxPW
XNwCFmAomYY3oaSPVuVYLrotvUVo++vnahHsdj0JU2l8ELdhRirp1gJq41LcSdke
6jFzmLBqXeR6bbfz9G8kkmkLh+wKuYQV5wutGe8AsR/6l3arxF22toE3D7+8/ntR
DsPhx2MwHMpo/AXjPxv1zOKb06/nfoGu/wFNg2qxns6xq0+SL7Wd94xexwpKpOZd
ypNj2L6yvT1q7Gt8xHf9KZk1EvcQADTwSv23ikBYC/RtSII+5cHRF+N/+GxsgM7B
q/eUQal9dougaNqEo5bCfnBUguynyC8f8bJOabpuJMqcBU97uBQ8pOm8gjOKanFc
WtBWYQz+wDmTK/csixhZjhWCAKwFag9llCEdPHI5Tvdx6yEFy3CLDSBEtWvLBN3h
OBXGGE5RP1HalthoRjPUkUQ8QZDXVz8t/SQuBasBSsHJrqaquuWjij9i7XOXg2s7
2a+h8eykyLw5UfjCATsqp6JLskZesi0FYb65h1jWD5uCwbLaIy1PyskBO+Kbi7A6
cTxISjKngsng69Ovh9Q1y9j2jY4snNFrLnGiT1WWWACnKQGAQNfKGSBl33Tu5NGK
9mPFEvg+o4HfEKxAoVngDLvjxxueL6h0XTm6JqNzzJmurbHXGbDJsiBy1FPhm2qg
Pc5SE8EV9lOCd/CPUHTOMNjY8XknXdiR1AhhF6LF1so23tD703pW2uzZydC00APB
ODsPsAWWOqudIVOFqJ8cwahRWP1nN0YTVNgVCm5Wd0SSJorgEdS9T6SFdktdMMIO
yObSl9VpeA3nT3hFzQT7bWhpqAdA2rRNQIVx6ceMEOdV6d5hI8KS2v6HBLOnx0Q2
u7HpvyBst5zZ9r0n55BjP8h9fdvZlj1xrTWPruAjJ1Hs6LC70960yCvsmFGnqs1j
nHRF8cax/2cyiqcqSiP2ZD9n7HRlRqASEKWKSkcIhpe1IOOUiYyCUOCmnbhfRfQQ
oWKyR/bWxSORNnQeFEIzo7e98xvqCTUS3K6d8OENwmnQn3Hptc5tvirCwMgS2MXt
PISBFi9SUpNAvgsxCodeA2x5Ir3eMc867dYnW07ypt5va09gCanwmux+Xo+vD3An
22YtXBS3qWBYMq3TxKJmS+YYbnojUG5tdOtvtVZqbsqioh3OHaG4KrJkS3kdGtVw
VcQwJS4N4c2kq3dyGut1ou0nWc2wDIDnEdAz2/09Iohxgir7d5JrN4PPz907swyY
d1Ec6P8LT6arAqCh4xD3zDtoWbODabDOWH+hcISOleQ4IPM5IoTJ7ZOz9P3z+1aP
nDjWYZmE/OVxVUQ3Vz1Ub8XlyoHP72V5HGy1TLVSpZQQ6dO6DZ8QwMSldyey8pl4
GHlxaReFXKtHNEjscR+lhmiwwJ1LvoJBrgMPbx5A164kChPdU1Gv8ziWBulOHhzd
jRY+9CSsGH/rRMJczNhHBReE8vIk8UwXccvVlB9nHrQcRjg3j2Tj/WFfFzgSJg8e
IE6Lh2AXhebi24MXQQoaSGc3NaE4dfifR27A27PjUDTD9g/WI34/KO7iTCwpdXWu
TQ36kGu/BANlzxme9a0euagAIpzZZRFxwQRu7M54ha4kdipOtr6lUaYH87ckhsRx
ljjl8h/e9PLw73FL8JWAMeut5MHOYr7kLkq3Y3bdx9lIgBzD27YE2Fpip+ZOBu+d
UEy38SomMsrpWFLY0rICw+d65ZEzeCprM3SyCBZ+N8KDwbracA5vyysqhEXY13qz
YZIjTOa2dO0ZdnuP2iu2at6HiCxrfrS00G40pWb09gVWDClRlkb4Xpcxqc3SftrO
CuOX3rDrZKwXwTPzQ0PM4c3W2155wjz30CcOvoCj5T24Gwv+EFTZQ5sqhPCmhR+G
BvmH/Erlb8w+eXN0iLw1Rbb3esTBlceP/EtUY0lBxOfyyTEm7svBUdtY85VLAs4r
1mzKGAow9BYftTe4ebzI8cyiaEen98qNl4YFb1t6zmJi71dhpQOQaUZtXz4Zxd1f
eNZ+OQVjFnK4UM/mbwKwOtx0LTRaHWK65Ou4ynXfzGg+1iWd4zyaX7LitKL+rx37
j/nm06MQOAyQG3PvTSC8j5Vl2kAES4TveLROOMNHsVrowSgPm08KU4mpgZBeSjYx
Is0f/xnLPlztFvtf0QtT2kjSrXhoORfpYjXt1yQwWi89CAq6EVIZdFpkR1xjaY0Z
luEtp/fozuW+ROUqr9r5VnIXmsvGlriVIqgrBoGgKNhElFTA/6Caa8zJJghf/IYr
0mz2SqS3rQNx/ek+R0uFIVWFKJSjR3bvBVxNqLdJkL4r8uSrnghKDbwM4WG+VqnI
qqyCr4hWaXe08miOH6sGG5tAt348iHxhd05027P0kAGb8RvFd8/rOgN8BKN7ptcY
Non/cuCR6vpVxcjMzyfxwXTAFrOxDBuDG9YBmJJz2DOdaTqiG1aizcMgx8/Pxleu
KPKG4CoL5KvnxABl1GOgu1YatEuxFxvY7ZwXgxqWCA1V046DCaUrZqWfTZ5ZMY6M
06A3uiyJG5ckGaQzH9JrBRHSv+i/vAR7XqR0bcU0TVz0h7Ws7NVVlYYtOM7YHYgu
Ov2nTryy76CrpES0FQbycnLlBvcP/hpnN46g9BZoJOjT8RUmValaGot13vrd6zwY
blC+7palEHkyTY8tC9LX0Zx27mvPettMGax5MGeBc82x7+mFtr7/r+lyZ4jcAjI7
4DxAV7rMet4DczrgzKB/eI6NZIhaKVYkBLUbsHdtvkSB/o5YH+DfNk4v1btj+ycB
20MgGEsGQAnVhnPadnAzSQ3OXfqvYSVQgki/OT30ipwiCtEtvR/MBXdzzPhTZ0B/
iVbkr72/3Q9I/G95RRq0b4aJWKBLzXeNPN7JVUCc1lrFXmsSDtrJP9SJIxA2e2j0
oQPTjX9CBnbs9Iy2TFoirGrG2vMdjZgaxIRcOdWiodzpUrJkSTaLUpTtyKLX1Yex
AqjMuEvTRJ2EXKjMaU/QdxWhejO32E//gLDhy30rQqg8TOU9hFJuvsO29qRz0zZ9
n2G8PmHHRQnlZhpztpNSBYYk6Yim1gnUZ6D3WAdXJgh0m/fwpKcTC2PWhV5KmX2l
ttIeqjcOwdoHhTD3qA0L3s7bp0cZP9gJmaZuOPHz5M025T5S85MWsy9vapCL4zTX
rrEIXhf0PQ7kQzA0sSWYkMeewZ4ylCA61ENoAF4o4V1g5Kdjd2v0yxIb69zYEcEW
EMFsj45ZHwGtRjAy3kFXPB/NdkFUWXIEBIkOU5GXIqVs0/phc5Ep7WN3MxAEOh2J
liOv11Ais/OEgoP4+9e4xE/KV5bbTQXVjf02RMWmRxP+WIQU7AHvwFwBDjqwSd8G
MQhnw670wtDDFOBmACagSL54KYLQYvbxDkuXxovxjOsCaVo34ZDOtknqzbH+1bgr
f5QxeUw/FQrBIbJ2fmgBr7yGWCG1GyEB8fEnLYyK7JiUM1vgotqHObaqQCkQ0Q5X
Mscrd1dlw0T6bBVjT0cf/Um03IbHjNOemzVJ+TPqPtbY0A7EzxU9U3IbyffLG3Fl
rq9hkk9uxWLTukWYVPWj26R2VQZrsWR6EFv8FLznhoMMqJ83ryM/JlgZsw/gWPzB
iKAoLVd+bLa2P2CtM+tb9iYCTLtZFE/TUOw11ajszDh+drIXCg4CFybGAIzcdSTY
JNdyNMh+5jv1URCLV7GZBDTsIE3G16h0lO/fd2+ydxtP1/aQi4i5uSV3ihaaOz6W
2kNu3/3KQG9TZ9oaSM1Mn7KvPJN+KIxcoZLI02lmS+VsVg7+rimf/AtH1wdyMnlw
2rZ5RHG0TqYx69WfyPgmewHHwIIIXH19UIrXpFeBHmtI3zFXC2Ik6eBYDyF7WeVs
hXAfQAWDazko+UTiP+RkzKUPWWvXLbQoyHLAX5XkVrvgeMN8Wnw6YSOC4VT67JgR
uq105wQqutCzU8orfQGJCB+Ib0Q0gn3vz5sQRAAyUSn0i7HQ41Bsfl33YM3/JJKk
v7HvV45bEj4lFdfbpSFxf3FzFz6hW4hnhC5dOroUZbNNm0igfLIi8djxPXMl5ers
jc5xPGoXrMkXxnpqC1ILpdYQV9xrJVmAJqqwmxeS2TLswhpLwBPV8POCO6+pj6ON
MH85ZqsEt6e9p8j5npoF0SLbcB/j3N9BO3p7QS+jIXjwq3lElbNT1N1rwtleX/9d
kN5HQjWC7wosPsax9ovBLCiZix5B2j4Ez+9zEt6rSUvDKQg908Ws/6ZTTxMO9G+F
wwvR6Nn4xd+crvTfKQMCfyDHU5HaMcZsdp6Sr5cUmAVOMhLgPpRipGFWiAorZjjG
UPeJ/ILiXpizz9ll/mWRjbMdSw7OVHWNdmTNoCqlIMJT1FTQyIA4GXhVhsoNUREP
XLnMl6Wmczy9KkdPv5lvh8b+8NWNQjTYqQ1B7yBEXOKHB/jlAK1DTKx2rmtp4QK4
JBRyzIPN1PhLRK3R+8VA2KuScrr9ebMKlF2bI/mLjV/+CBt1Ju9Z9lCzkZgdAzcC
PFypyNNq2GcDEHghkGFe8EbSRv0Pg1k1VpTOGB9PMKs+ylucI34wQyyYPjc7/HRw
gAAkIutKOBaV8btl7tiNsusfaB2Xkl7aVqgJC8UPvWZVncZKHIe/wtU/XGbJ2Xwm
rK4QJ4P80+gHTXP73LeDSk48nZJiNe0ZaFRu7usJL7D0AyQIh+YzCD92p1avz5/6
/2t9L0neStEOhIW4Vmc4IBZ8nuKsFL8nkEaOavkRbXJJqMNoOM1UM1b4j3+BQOmN
0fCcxM2P2diFvIR74EZZHOrbxWSBa1hHrs/q4un4pItNrAiHpnm3YMcYqYMN4Hdb
nEdVRB/2jV7J5jdw5v6qYtefNJwMhyP7009BbthyvbqUN6asnZbN/fwHetD//noj
D1YsAkFBt/4F4HuYEaBl6VQIXApmxHumlc6UeI8b17JKgHeT9T+Q3HSPxjxCyot6
jyR0HmIavXhD99GXx5jz4Lk2zfd8UXUbsVKFVEHjfbhcz9Xfzmd+Bpl6WmYQYOx6
Z/3OrvRq180SabYtR0fEWDAxuTm2o6Z99HP5pg2H8tOzUaXSXJWnH+Z9paEbMDCl
X0G/ghMSbOQM5bEFPxFb+c7lJ+vymQXMYgX5EpAJytzctKDvWFOMcMhW8JKOC/EQ
pqq6iWFcPpQ+xH9XRA6CbO1zWSA4zmorEa2/gG0nz8PHo/OlRTMUgN5vYMqU3ca+
20ixREmE8IJZhkxn238Gvtzo6VXu4RpMhwb8yIWZrkuv+ctBl7eHaifvP2lbqEx5
9GNJr2aY+g43domh0hC7S2CmmOF4k13nXEx928vadckn1D3XL7HbaWCygmornKk9
NG3WxFjBODMs0bonUBeTOS9fsZ/9Ez1N/XIc7Os+WyP5moN3aUdCOjUvSEi/T5ov
0kyC8bG4tFrZ3DiJZxy4aIgxBClAxM9wk7z6v9EXmGsNH9gSF1YgijrTvx9bj9v8
Og0fSMG8IFiIbTq6p1Soon+D4ZNu4cZx3Y6gS9ylRETzVrVCAFhRrux/hHxGEa3Z
s9+mdQA1sUkP4bqvHJy8dObuIj1GGF04zwmz0UbtZSnd0ZUQCCP6yKRMFeh16E3V
GNClq7tyM5yU7TJL+4FRGe9G6YC6Rxh26wnWxtOfU/aJJ+fk65mIuhRCkGL9iU9c
TvcAr0Uv5+dvFdxiQmJ1as5DLqeOdtt7aladF/nIQ/rjOOSEul0S0pjItl1SVaRM
9EyQDuMYkcuztHH+ODHIDgEBt0s0uz6pm1/IONGrmEylwL/OTrD7/G+KoMcbftKk
VOlywtwVvqQ1DzcXx/6jA1O4tNCRRGdsvJPCmOQNcS+NkjtI7YhUnrlHsWuk7VMV
wZNJIowfyL002TM7x+g0xX9GCflh3CVbiT2UvIggFpGDgBA+nGV8cT/YiIRSLZ1d
y0A/jh3GvTYAYVw1xHs1zdBtD9Z8rByLl3LQ6OgDlETITfHy1RMbnmiPZm8tF04P
iZiwtG+g7X9LoMfcGEWjlH9zUqese8HM5u32oDmG/8R3wG9ZJK9+ooZjIVfY8AGF
Ohy7R17GoDxKiBL8XVl8Fwmy38A0qs9jq90Kd/A+2hLulknJEmzJJyQ7NBzcPdce
j9KRCzXvo28ubjzFRoeTwlv+LUVfMJsZQJhFNz0yZRr3Qp1CbMm0Av0S0Z9VHIff
4er6gXaDDZpeVzkHsiDg4twZ4Mwb7t62stfKRJPvTMFHtlkSoz+I5Fxmu9hQ+5y/
L9yLKTcZwp9UOFeAnec/TREviYa9olJYBqN7M4D+emrJTVbx6E7ywBgpDHF1g2ec
/mcjCSkFw/oO6BXJrcwjK0L4M0QnfB3pPdJQWP/nnhKEQpD1Fm+P5kiQxJlDvxp4
S9ES6Be+QOHWMcdlQDCe1m9dMVfv4Srunb800KavE5LMxivx65+rgwcUzQD7NDeD
gpUut5FSEIJcAjBeQ8LkQBVSTJxgmjoMhtRj7SNeSNOknJIcUAAxt/BUi5ThnRnH
2bb7zHvrSIjcL5GJVERu3xXG12htEoPMoYszTG1DGCiSGxDilYCLz6ZUz58GqeL4
IxJWZAQTHXS7H86BfWbJSXA+LOQkG46pwfZoUBSchXM42j1pP8K3BUC+WkiTdPYw
ywQUfsLj49FKSWBNKBlYXD32+lNshmAKeDknMJhbbc+Yx2z7uWQ8CW9VaBid334W
1FKTaK0mSWrtv+YGcJR1lgbpBalxWj/tGPHtCDN8ScyrZRAs5Je95g7nQMlBwqlp
a8J94NsGs/ztd7Bed/ixLe1/8pk5Pr7dy1lueEhFnEeUE6JUK7ip14ClNuE8+XDR
IguhcCpRIRoaAqH18r/v4aLcWoolXHme3zIiFs44fDRcT4T5LSSI5RvWQbp1mDWI
1p9/L/O+LRvqnX+cHB5pqbwqGXYFnmNdddjccy6GMMyh3TIeIsjleHd/2fDN9wdH
28FAnyPQrNb/OwXFT+emoKqzlHOSHPwVXxiA4MoNeoMjLZeh87hPGrkVRYVOlTDq
e7bFFs0+TMTqvFkB1/7O1Tifwh7xii2E8x2v9ce3GkGvupyrCPR0N2wc5gy6YIYf
Yr09e5m3iemLYSLA334y+1KO7sBNt5sZj9ii33ChygZ5JI75MPN+ZXY7D6aGRUd8
hek04oG7EVXL17M+AW7ZJY0rCBY7n4ML4JihmUQtCD6x0DTiPVHHkVz4pZ8v6Xsc
ZqMBTKGv41eP2+EQHa9CjK2BOusuURq5nBL5Kcz7ix3wpXZ7+DCatnxN67kzj/tZ
vX0ra4d/X1HcI+DAEWBQpfq2vBq+Nw4C+P0EByzI5iCvle1TYuO40oFyq9n05Gqt
yyob6+ZK80Y0mt7a0BKESSP1mSufH2abJkmZTADpF063nJ5Cymd3eP2T55EPDXyn
A2qQc4J5+V8b0xh58/4a9PsfF5Ea4chXQ84GWXBYzUIqCHVsbqoqjM7hzYS9ipB5
8AD9/4JGvpnJQMVbaxoyM0d/oAPc9ZAbGxruFE1MgmobfBJhKARAh/RR1OmM3KrY
y79CSyH/ER5Cvv5BAf5xgpX48zCuIF6MoIurQUm/nnCsKI3KEESfUXeHXuLhfc4A
Xw8Va+mP5UNLbTMzrlfFyXSwVTAB3vGxvW4FDES6thJ0CwYaY90h5+92+0EnBfnM
d4p63HkZQ3GRU0zai7DeIuBleaI4EnO/QzdhXNX28VA1HyG0p1L/K4gaMmpwZNpF
lRQWuzo4aCh1nWsKS2MpY0zXxYNelZ91n5ymLXwlibkF0odTaAZ57TYpJJDjsyCZ
WqdWHF2BdAbMOW8wYiNY4D7swS6J1d4kIbZiENQbf6La3r/WC0PyOPI4xsuJZSvm
x+jBGgowQ2NBeCC47gzDvTmYRp5O62W7jpH3LFzaVJeQx3vtg11udUI+NgRHSihN
gYe+oG5aB+tb/qFEOywU4sLXCDIp16TtDxqh0qcEXiiXPBkfBfBahqEKEo0F3iPT
zULvtA28WMvwjIW0qyfUgGQsBVjM1iA/0FJMKeHfIptluIxMcfHOTc0GomdAiXRT
t9DjCSe1xiTfUVq85xL/O2EhL78bwMTt9gQjHkvEbOC+emdkpBqbnkhy+xw93uFV
PkAT1MPsKg8Q9uVTB58PIGe2mjDbyrlXJYnEAp995+KmD1h1Q8UnWElbm+GSfWzg
6EFjvKTMgi/LDxl2N3wFrksCHZgNNfsacJIl4whtLRwB77Gt8+d9MXwZZaXyT7LH
xgTxH0UPvZaMmrl1VDJpsdPv+Tm2woBQpK52K4uW7TujLUbOB+pSR5A+XvTuNOoz
B9WRviIBx/Y7fmIjFuMDGw+uF4Mc3ZaAYV9DB8H1/k6YLiYOHlFL3VQf9Zys1Htw
zx4Dl5YEP6vjabYgm1/GCqDPbPl/w0ZVoErDBKnzQvDfoauz1CJ8rikDsjAuDAWu
C7Ym+10qZZxcrGsYVyb3MMdSUg+q4CaMVVUEBkqmYZcc18oZJnc6f9TfwM+XUuPa
O/NIR2qjbx1TbREDC0WRH9QjOCmFpxhGZuVrzIJ+Q9uqxDVKG4iPJH2OMUceYKoG
ghicTOpF3DAaez1OVwbq4lCqJkxspPTpkHNBDqNthEy6/T2zPcGrn+UcmpQ3+8NR
LvyIrCvqvk79PcGJkKNBVrbaDZe8En/bAwJowKBlpAuUmRoAi/NP9lMjmf6Htywj
a/JjZh0d5S4PUrrPnde+NefPNX+KEibe8W/PxoE60e5mqiodlwMyBYPd14oNVIVO
PYjg50dytsfj4z7jNUBTO+hit6aBYgE6Xuh4gPrXT9jl1n9RCWm6HgzaylVnzq3b
odtktTdB0p3MlCh9qoNgSkMQjod1meSHMdlNyfoSOzqLt6TThy2Sc9aSaEPrjVdz
bgDXi0RIwd3SNmR0TmKYzczclizR13I5SLFY3RMkZpC9NW4Er13nIyKwF6HaHy5o
BgxxFZ/W13aGsOjp73w+7ayFC9SixIQwUS3qaJdxzztI6h0B/gUXmwnldj0OmUKp
z9QGJtBuUkA8T8QKfSFy3hPvxN0VQxfZT/i04Q7FnC1WqqvYYpaNUkCGiaCG995/
vxTpQycNlSOXDXjHJbxdl9Cabk6z/40wvKnl04uqf/ATtC52zhnRkWqdzAizIQEd
lu74mh+mrCzDSryMFylz0Vpn+MdinpcaeVUSvAp5/GfGXPPZxsRDoAJjncDVk17U
efdxOwHjDhO8xysutUdWKnt0nx7UXo1JP/GaR3CCuLKfCaNoO23Cnp1hYxKAWQLy
6LZuGScJfe2DGbXI/yFlR3t7uzVuR1DLynFnhbbB0AzPhdLgj72K85VrToy/Etof
Jwd3RReDU5GXG0AXQDRRyQeXGr2ncr+tysE8uoNScXlAhOCaif5cq+vF267OeoXR
Y1ygqZNdrZt+/HBBbKazhQl8q+1haeJVvXRniq2BrYs9wOdj+01XPdZTRm+rThGd
PSx3Nf951942Xj36MrMuTadvJ2jO16wff0XulD/SpXpdvh3TLvgijkDvd1AoIbYW
/c+kK8LArkftr6TxYo3TgVm7HfJOvpGxgxIaR8gRrR+lj48Cg7NcHBLK995awM2D
UEwRni6uea4SblYVthrA/0K3VKuSbs1Ig/7Rai78SsKnlKo3+hVN/BgBFFqT2vPT
TJCGQmrO8YDo7K7vbO1JTYYpIsZ1gIMtTWhPziDgUMDunGb4zRT0w05uUPG4Tjob
kalrd1IkqjEbV+tifYPpWL+4B7AyPNG7XaW/D1kZvpGKwq7+JDa1xZoM4jSjrPXO
LQ/URZdEYuyXVbF++UJoDQRsGNgwrTjtjvn1HTzQ2zyypJ11M8XYVm0qWYFmJM5f
8nEJeSHuAScTRepQGl+0OLxOZzP5ZxcN+n/v8JDGWmfM53JuHFmo7krEVRii5s42
gE/o9L60vXtslKH4wqTn/3ihPgGp1l+La/CnUu3Ew0a8VdBFcgq78udbLxQSmtly
M4Zo/hKJkoKg3+IRLtwz2xjrxmQDwRkRMfQdfc+NsHv+FoBwq3AcLfq5H+LFxsDo
l8ujOUkA+0o8EQSIO5PUzF/sufODK/RzRJAuykhf9PvqI7giu4wME5ykDlHGZDLQ
AfttYLhHRJ+HwR9Cy+5Kauq8np0/IjcbBOvnBwcBtWQZwkX7xMzhjhe/1huUuVWO
mDE+yGSJkolnR0FII4fngT6jzkvvo/Y7Sr6UbTZc8CeI9AbtnTI+vOO7uKN0mffw
qPzPtu2ndNM7ekqkkqFf5ymp3Py3Lk14VTfsWBvsFAIfkeUF2Sfhq6hPgnClKsxv
4ORetK3EfD0r8EFqA8guG3auBR/a4ANbee2h4A51PjAbDidjcEdrrIbN4lKFU893
dHsisCFdmDcrYPjoMFWgvsTDpV2hfGguCrBlb7Ramf7P2odvjo62xhxl9bv3As0M
L4CJQxKtmr6x44GZOoHck8rwZxzfkfv42LwMVX9GBNwEwVJUQK1ydnlr4IJRAt0h
uK5Q3ummwBD+4O8Br96lyfZtZtX5DnwNJb766xGDpbiRHtlNI+n3vyEuzuQy4+3h
VWO1WBR6bjNUX6VlO9W6EWESllrg9pnSe8KphSQBI/+AiN/GSf55mSq/eOtcR7Oa
c0dvRPDMJePSdwQYeQrqk3DKl3GwBnxqN3Slni8k1dWoDViQ4dn9iQ3xPejafO6v
nADIbsjWFFYb+ZXsRyJvJpZt0iazsjUvKg4d3GcPL7AhnHDy4P/ecaS3sDH7Z1JR
1jXSgnylW7vnDrzjv06EibXyRTP/V7UjvXjmfGqNvGJzxtlTmZgK1axXV4gQq+QZ
qCGZZgTdnqLvOgUvuC8goL4jHNnLMPKzCT3g1q7zlGrZT5n4cCn609L5Kw1jPu82
2Q9xsCQ4jfFP24ICp6Me529kPHDvZSRW41R21ZQ1c2tt8BbvMTTD4wCK4vanHaJL
4HdIOoMvLnU+FalggMCw7Bx1ci32cjlkwWw0gO3EZSBaL8yL334hyMmI5EWmm9oD
ZBUJqzdTaPt+oTkNXL/R566rFwbwCCtzlNu8xcLGpdeNswC6i9DjgkP3S0x97T8e
Yzszge9m68bsaKqLDlQm4yPKdWNz7WrPwEhyc04AcRXi+mmqMdgaBs+Ie6pqsLHb
8HKsnILtJ5Qz8wCRxk5XwtLK5M6Kp9a5lIiR0mWfJUX35Cyvp+DkAb6Lx50gXe+p
fnggBoZIp+8Zkvhg2HGeJ94frJLHjgnhZ2aVxPVoXhJN1kbLR4SX7QdrcTz5wsvy
ZNTJWZyEqJY4i1EjYrJo1FqyF3faEZwn0nO5/7JHr5R7N14FupVLkxL6bc2RVvcs
asspBZlBiFossVtSAsZqzTvC81GAd1HH8Lo1NFbu0Cu6dIXAbqJWuWg+9p9TFgD/
9UCgogEfaUYisPbMLNayzY7Eblv1e5VB/kS+Ro5+ifsnxcXudZeMfpB7FabSN4s3
d28rvxgmwEIcPU6iRyIuIZ+kreO5+SKP3eVQa2gY7kPJ6XvzwAQdecQ/fsyHyTbP
E43eOvSZH89bSvINywqQcXa4ywr5YcrxA8rDbw/uOegSlc3ZAWwEFLyITiGwrulg
E7DHC8VNz5ndtFp4BkDR282nPiQMzLLFOJvOsIrC22ONpDMfsn66j2zJu/NkQpnq
rI8BrNqU7zHay8aMEMFhrQqnGiA/QGavip3LJfNtSjf3DgMljbYuBs2tYuU3Tn6p
RoG0Nte7yqRwW9/3nIjiHKm10K3mlX9PXZ4KP4pbPkCrLDMYOLWiN9vpNUipci1r
dNlDIovKlaO2Rb29X2wW6izPz/x1XQ+dzZzsRzVEIEMlSk7zbs29S7n2UYGT74J7
6qEATGMQPrI5pH3eupEFQbXRSH8i7oZ/eWrRC8hdZBr/vFmoIZh9FP3vhjt1lRQv
tIscjtlnCHjmn96AsTWe6L3ATY4S+VcVJ6q5+tKptMzgTuGtDnEtyy4Rzy2Fzsuz
61a2mWZdrdj8Gb3mMUWEU9nhPCdbHy89Tdyzz+TMH5p2R+qtcZua8HaPj2SkpoNd
KkgZag0oAw0VvEHWjl/stwGJ8w/aSO8Kji8xUZG6AUwGtSrYu2wFC36uIQmNDNyK
ea3VKX4pKt9dlpEw8ZWs8CWDVLs6JTAxzz/ewmVlHlGk273BtJ2Bt/hdn5h0ppDk
rds3GhyWIXSP7J4LknNpC6F92QweCv9HfVE2TYeUtn5PTa4+PszgSX/wv2/PuxEa
gBzt2Gc1PDzj2smfKV6hjU5Be8E27P7Glu66E4lfKKDfJw8KLH2Ly6qRNFnLB8KP
PXzTr83kzWBHbx5RY1RpS4lMJrD5MxLIcL3gvetrQsr+WaTmYmIR2zHQCKwDnjqR
sD1KS+O7KLdVKSUUB+SU/SLqR1y65zJa23ug4NpAr67N3rv5ukuoZUbeHvGWFpSl
MXB8vg+TV0Oih7mUX+YkAJobLNJH3xM0vF0E6G7ctPBkhIqQROU4Y6SFcgAfO00j
+93zqpB+j5XFUlj0zo4MOrfkGR6fJFh402Qai/bei99PoDzEdC3chSA0thQp357i
MDZ152X8ad4FEZpyPbTNhXZfkVZJuQnZQ5LOb0i7OtxKnkOLg3UlAvZXf2gPDHLx
Wy9D9r8HDDBa8wfv+vn+suEKjnR7q8JozKyzFtRD/Ri3qVAslHKoWY+WRq2+1Kir
nn2jRHCHCnsYmlRWXDYz2bE1flE5pB44BY3d9iJSfZ+3ApGR5XyJUMkqLPvKOV7f
yBGDWCzrqXP8tw6xB9L+CXWOkEejywNM5jRmzcgyWFHmrVhHvCnJ78a6+bTGNTHK
BGWSoWlZXBzt+XKcz8mYD7dED+XGmq28TgnFaNrHNCcGcd9c9nILJLRJ1NaHrSwG
7FmvNCi6CbSCuDc10h9uWARKWHm9NrwZyE8i4574OXAwOafZsDQ/hiyC8zOP8ZsM
ZlsDDX+peNrWTiwZmOAkYNRpU5o7DNnM5HFQ0GpEfNKCc6RUQ7Jlg9DdfvRf0lQb
4XZU8DCIyRgYNXTB+MkvqpMes5HujWLekOw7tOGBPC4znLu+M6FTp9HBsPvDlmMe
9aMJx0RjK8xSXI5qd2ktHKQF4zXTFlqJxITkDuSpnXJbOOChuWFgjEJk3OLaf1+s
hjQX9297KotwDirmch3txneYetPv6wAYJltVuXMLjZ+wn3y64lliFARrhTjqPk+p
iJYaR+BOLbi8qcC0DwXwtm6vf0F4BU5YyUs62/OKB/kX9SJfnjjV+WT8w8ChfYAf
tGN99f2tLW17IyVV9knoZpQ9sqmLYagosMRDSI5Ovx+ymXPy7sBv2jnyAcFX8irA
GbaKJw0JOxsI07PilZmHNLqYTUJzrGXLS/A2Tp3sVhvHfE41I2ouZo6AyIoUAGEz
+7om1lA8xlAlXKnHYWGFIOWvp/cpSObQ9mPpw9aNTru5k8jRXiQa1KRScX8pT0nJ
6l5Q6ZQv8lTL2i19EulM6vGL9JOLr1Z5O4GCKnlT7S+movT0SL5O4c5EGlybgXrD
b9x8HojeBb19d1N9Xy61pNj07iCcxwqVLskfFpozXEP61HvpO4PERQWrEnrsumSs
mGtYt5WrHmAOMLjuMohcy7wz3ioaIUll8ct3CpEtW6M9saYQYxSYQfJEVdBTND54
ruJ67VSFZzePAeryfjDMpb1LQWlv0zcv6FpaTg+dvSZZoyqBn37aqxmiMwezGx4k
N67RfII1NGtelOr7hKpht3nKWO/OgUkSGxXELh6By7x9RX2Oma9SDr6YrX+A0eiz
7aB6uFufe76Aan9BzeWO18JddDwtnQVuC1RPWy39jEjdfYzJEwy61P+sz0Tlc1OY
FtApDRLL2VteBZMItQmaibQyLeW53skPFJU93ag0pF1rSq/F2iveMi6mW58sIInA
vYlQphFp+ZtMsZ5Ig+d6vRruKIhe+94qTIBBy6xhyVOp4OznfllXHdUggCfczULP
KiK7uKHnkxM4g+MrW2ZqTfP5N8QkwgYPiuKsVCorTWKz/IZLxqU4KhygXnSOlTIY
64YTSbebGUIKJIRiJ1FtbiiXfrb8DVYbGEKBI+0+RRAIea3jmBd9ykKz2CYokXJ1
gjD6zYXyOZYopjZyHhsVq5vHZVFNEjGXnh299p8vSqoB9V5sNLHG7fUzivEyiTST
8dqyjQUnkwUHTa2LW2CVgtD9Dqgs/dew6uTll4dPI75I37UKBo86ilO/4JNudtN6
WUJZl0vKdSr2ibvZeUvcncNGBtqt9AciwM/Dac2rC+CktWy8xHQHL33xBDTMF+4R
7YYKR3l2dOPdB/RP0QYm4cYAQVukU/GFh0Npb/rOBU9uSnXO1fd4IT9dDFU2e0dX
OvUz8C0Xy2x5HW0hu9HVMr68rJ/uiQSXZPPPwL7LfVghCLzkYg2/7jBvAfS1c8It
Dz0g3MJ8MLSu3C1SmSuP5S3odg8Mp6tFx3crTlv3AxPYZNBBy+t9lCrgtFf2hwPG
OIiz7TOcmCdgJVoFB4NxmDYCYajuA1XSUASaDRteHknJy2hKff20faZEh5sRENjm
3o3GHl6D5sE82mn3Jdh+gtP+hCqy/Bcz3aaI+fZDAhIvCK1/DebcT975hOUM/g1W
Y8TFEWshTH61Cx224rMa+qLPUY1jvf+ergFtbdEGYPIbPx/X0WG9+b4AEor3Eitf
lHzTFj7c51zEV0IPjUBI9QNMsn2wgic/cxvWGLT5bMiCgbKyTp7SoA5jCuUY1hxn
PqCUulRhETxyPo3pScMAiMf9dRPVH7Sx3GVjAss4oG88EiuLPM8h/TZFGMPmgvq2
oLGPjJorUk/fDAPtfIUFblwap33rHABa8NplEUzclMVKasKLAzBeS1QrZpz5dshV
8U8/p0Zvp/BZy1z/yoSbhh+IB2od4MlCovTAPjVRTSNNsKxRjOi/RuE/I3W3ZjD0
wXpUo7SvJrFSZ5n5yPGs6Q8m7+h7Z+5BYhKqg9S2kNFnYQTgYON4IPVMIh99XpX0
R+7HRAr8V1cTbmXgMkg1Rx8+jNjWa9m0Lz1XDk3ml7u3kvThv7Vceg45G2PxXq71
s4nLiWMfiHVsOG5zFYMohyGGY5M8YKfC9CcvHYU9xL++SGBfRjcdNkw1M7KAHXUe
aVN6o3Dq0r+bNpsM+rR2k4gRtTIgkW60Nn12CN2rUXXQzwUtBebq4fxWYl9uNGr3
ORGAhpblYNA6o9K9VU+YM1flRdnYh9d1tiuklU6ESyZs+hQV2+8DtIx3cavEqN1e
wC+8gjS34mA5wR/dkDd0wY+SsFksTkVeGO4AhckcQr/G+V7Gwk8qMgeh8besYzPd
VBEg+o+TxUYb3Y8OfCqJUoLie7hp38kLG+8E7X/7cCa41WBDA/RLmztcD6jMKnj6
O0B3I6b6wXgnG/ORu4d/5N2cUYTVd1DfjclSLPuSxi3MSwqlTAgtPLwXP6r65sAo
NaSm+HR+QTsLKeNSrPz7RY5H5ZL5edF0NWzwf1Em6Hqbr79OXqESU/RlAUNeXmI8
Rd96vh9YLK+JdPPNZEP5YwoLZ3bGjkHMzwKFpibXJtPz/jBgvEqcHLLjaKlnGAHy
F6QjN0uIB8fABvCzXkHz9VZZqSnuLi9Tg5NVc+x33cJmTIvh/4EKjM8awtmRdToF
gu4nayDTilXPOvBe25XYTnAtWxr0NjoBE9qhsViRgxAIRaZbqllYyoyQaIwWQ5bk
XLJYwsGV2pPQY8ixAe7gA/OvdVscTPrB9croOz0uZU1vhR15b6+y6kzpk1kBxpPr
J7Dc66xculnh5B/n6R/58ehtrwc72NLspGlvS6dJZZjR/iLigcCoj0/ht/7mR7o8
s1n4xNVY1T2aXYUZWJw1+LXWTztGySa4Ht+ahCxJAa6hpSdlqiBQSRmmMuzU2yDh
dnMg2TPtu4teb++9xx+1vvYvjJZ85cp+wbNNRB3313pWoW+rQQVadlqy1v0BLgqQ
eC0d2ZzqdLIaAoC7V+d5X9eELXKEj8F4j1RbEzj/GU4XXV1GNrYRJNZn+0xN8vFV
XWkWhvgD0G7EGeKP5BQErbtqXDWdV6uZp/a1YwS5oGKa5eejUopAJ9ev67umT9BT
ivFZfsGrw20EguiZJYJ8GwJmWHIznXYj3vAMFv9GedKv+H41MSzh7WG8lI7ZsPWw
5zpOKZwiNPjCBrbi1O5Omrp6BJNC95WCGzROXJry+joQBWs84GhOvN5k8fOtNyx1
jDwGuc5WDXvL3e+DmcDCT4zXjg0p3XNA8yjMsgot1zUU4iKdYN+umZc+Odqy0rGu
H2CROw0Q2P7MN0Wdg0hIBDwXTvPazhbgvm3yqCO/+AnksjsvXnQIGdUjqnaLbs+X
D1JlsrBCdcChhmJtDli1PpuIwq500Q0sSuAdobMqwWcSL+5Nn2CeNQ9AnktCumob
gaQUdN8ehfm23w15hVuRh7F+jtPVzrXpQp/LwajC21cEvaObGmwnfEi8837jR3Rr
6bgRYvSatz64AOQsNKy+pRUPthV4YlXmBuLTSbZ4UhzGkNCyvlJOT2InadAypxj6
QXyIvzDHmwADbgTBOevuBG6k7FIWbJ/5T5dPDSKvruMSZkhg3tFY+MQbuh/MeVCs
wysYrVoneO2grcTbG8P6JHQ97Ybc5Btvk+ne8EGYubmqZK0QZMDSbSVMcuPvDhpd
iZ7aWmlrbcc4J+69lPZLdteLDHF0ilmhrm8+4HkSH6hRXe2+TUJhGA9OkJ0VNS1s
agldr/10vBonOoM/CwkK/koyNrwie035yIO7mNlaPfv4YMooc44zOehGQXdy16Ur
C89MTIDc3oClvKMfR0HiRnsslTXpWSjyQgsC/RCVpA+HxFT6yTmbvpBkNlWJGu4S
QVc+3byydsTn2j2+LuT/zPcKz6IwwxrzJpTkBrVtgs2LBNsUEytrZea6vT/UH88r
G5hAEbknqoSDaZ43iWUCKdrpStD/q1r9ZG1toJd2jdLnfxuZot51zvn7+HYNDy5k
OSJYHq/tOhiyCUV+XnLbXOMpGAT3ASmMaBwBQ9sr+KixoOhHUfZvSSPEGFTOSPfR
WIK/+A/3Wg9NoSz2miaUDM3JMHKrLSQ3tfqFi4ORLj6RlNGKSKIV+7+tH3f7TPTX
CnSz86kEuqxVZZcHnvLJ6osJVNGTyU2Le1sJYClk5S9Njhvp2T5DwqPA+/sSnBFu
CvKb62WYiXHltIZ7obCjgrD4gCDOnNQ8kiemPJcbfNVPM88LzuvgTkeNd0RzYyUJ
KTGbBoUeTpkCKkPbizGwEQ51vYDR7oWyHr0E+roaf/qgary44pvKNvD99haAjvO8
IvvmtG1tL43JiLaC3lpMIRn95O69vg5PPd+zc3BwD4/W6ZN7zsXCgVk1prr8Ms8v
wAgnONF7QqecWxhGVAGd6z6B5Jwrlgm81dMn7BObcWcSFO+nAbTdfdxQMSFwSGe4
B9GsnzifXcZTICZ/B5WRVwOv6hhG3N9VkqxJZ3sm0dQNFsolAwmcaEw2HMttQmG1
i5BN1vhRSbjowAfX+k39nC3L88xRCH4RnNi9+wMyGBDP4Dh0wJbbLosHd30NfIOw
Tyt3zYFrz/H6IC8gTrs8C83YNWKdaj7oUFncMymdna3hBpvpVXeqfeGnfglPxwmI
wBF+KuE9f/9fjFrgAJ1kSQovSMpCStwZwO8/6aacg2s6yo3s85N6jOao/A+bTJnG
BkFPUkG0/svwF/ZqwfmrkYUh9xqm4ZwURxNjc3KPpHtRiqJ6fh8PwGfCAqyKcWLV
lzdK2LOgg7KWJN1EVg96SzVIYCLDSPSMI/NBz/DTGiHbquk8o0gt0MLADddehVw5
6mOA1hN2w0zW9o0Xe/LYs4m9NVTEtDxvy3nU1WVjpoC8Kqv10ZWv7cwsuvLnO+T8
FQ0VGL1uYGq2/wAXD3GECir2rttxUie6hKccElZ3/U/UgnO1hUWPJxXzywDclUMZ
wPtEuF2aY8yNDpSQEzBBnZvSafGOuBtHoRR36TGKtbNoFGCz5YtUTXzyH6CFChfh
+BZ3U7WyuJDmB2R0FSwICvMoN0wrn33xjR+ziK+LJIa4UkEEM9dDmbWyDlXE5bhn
yTamovdq/iLUNG9MAVeDdscdgkWM3GkRiewPWQtUUCz54+5NXEPNSzWNzaXQfpkx
SfXhWWsbMgdhnTvKCw40vIYt3O9S0NTFJzKzK0lZb7PxgH+RQ67Xll9ATFovvVVE
Wf89iTMQr4uwBRvuP+MhWNrYRu6vyOA1JVlceVOVTWZJo2zBKuwrO8kLFGd482wl
j3kYSJrtLijUQuUp6bsgFjzJz1Tm0CRTigxZM2BMeFhuleYrPihK0KjK4UevOvLR
OcGHkQS8Bibt5HntdzhJYDBM/naADCfiQuawnucDcInbPOzKYz56DpJ4rUHW3rHo
plPwfniiDxRaPzYXorx2M8KkraYqoREMEfk8beIkhXHJ5ZwnnWGhhakFx4AwCi5m
xF/3KwjpfyQtqjt701Z3+Oo+a/Uwvfv3cznr/Kqjbl18Icf9Ngu7mE+XrkBaMXad
fwGmyzYQKq+syYREJ4yMhcMmG5tIZKP48rJqm9BAQI0EK+JmpvOAUlx1zduzo4RE
BkBdliBEJYcK4c6c8GAKedOlWClxk5ypu5f3crI+K/3Nbh7ckn24RntKzBrPu1I0
4+E0Iz50umvVlQybAbLPZm8tTIzt15CQtbFjT0Wa5a9pGVNmQNn+DgBs+2rU+hSC
mOoyY5cZa+wajngylzWK7t/7SwgcoIvBHfH96Q45Y1sbF320GmsEIElX8RYXuriY
ORe9U3ymW5+sZDfQqqBe6S895Z4RP9cX7pCuXzCJJEJTPuZxtuv6S2OYvZ7w+dvO
lvdTXYP2xeLyWPtZN+OlKXHUH15aNyArFq7Vf1oz5mIa1wP+mBI7JkViNflBDUOx
eNXIZgdWVw/3NYI/EIz5Eq+aN/zbspwJ7Vd/1OkRvB4M45mWUttwz12s2jow74WM
oaj96zuOGI1ic+px7N9QsDk6SUMjfs0Hs0wYSFkwmSOWKzdGBi8jvim4j/mcD2UI
JEzF3RA0O9bXldRNFOhRpWoKkT7aJC5mDJOraqdV0JzT6Ds8bkhgAMFN/wetIA0/
/XPgyMN9l1VexVe79EXz+fj/Szo/kKRmbNGUHuKTMgymAicIJoc/h8iOxVzg7WUs
hMVVRImqaPPRvdR1ktQA51wtkuw/pqZUMMVkv6CUSZpcfo+1tRk5S9YvJOOdPBbi
r1Ez9YVyMwLeNHUKjNk3kBaLMIijH/r0SogDoMiDBGeMr5se60MV5rk321/Je0z4
u7H4FlsTsxAw6kYVr78+8Ycpi7eCW4TyvtjYTwPmLW1AU479Ou8m1HW72Lfbx3uV
lgrQ7xHxooTMsx7bTMxqm9DdGGXlfWCiP6Ufej1cMM151CHGkFnLwuHcLPPL073X
kGbyHsQWj8IGstKMbGk40OuXqC/5EP4YPItolpKuORtKSd+b+OGWy2kQwtAgUlNj
QibGLjWwXGa4tfCtYeB7eRyofPcHiq3ANrn4RzvJkI6AtX9ndaqRROXxLjZBaUnV
V6bjLfBrbGryOR5fCFQfj0uRbe9rQ+ULmt1E4q8iIoTc3xD2YypYujspaiHqcp/L
4bJMTwxds2vj4H2R94vGI/akX4Dkeppb12FOD1gl5ptWEPfoxBwaafdi+Bg5nI1T
vnq1YhFkcLIpY7B/jfUIyajJa/SD3xjuYYzT5CvNpxfmPaNZngeBYpIoxYfXg7lW
j7pjdzK3YLcDkIjbBH4fUa6Dhnmci11z3Z7MQAN+UPO60usvzzHYkoPFwXZwPAHo
7qorz6ywFUMjRazkgf6D6TN8R0Mi9GNpeMtEHz9aj2zuOp+i7aiXrHbr+VJ8hw9e
NRiRtyveuQ3SdcYppQ9vrYhgLccaHGFK6IOqDDJtSh+16YVeNCqHT8zAPSwGvCfF
eP2hU9fmhXGSOxHQpsK0qBsQ+zKIzbUpOSeClbkMpmGicOJvzHs3ae+5+XJ7gkUS
5IzXXerlhTkCtCCFCfCCr1My/kNVxP9h7zsJjR1l3/2RXqL3asilRGDIqu2tKk0Q
tcgUcVpAgV9Wfo3bEC7M5g6+y3lX27YKTkVem3T3zM9rJDA8zMtdEmFnNaTs5+AX
2zIoldgnuJ6mmGcaMI5zxIhuBpCmmULjBF/eE2yqLghobVPcUfrc0nQJCBwm4C2/
yO4mD5zHVL7FmRjuZE4I1jBw7WAN6AwM0cIzfT+OPNXKkSx9K9Qk8uZkX+GPMvMU
AMlYK4yFFxQ0Ij7TjBAlE39zD8u+o2XePDKfqhtIyXZfry5FbSB9xXbxwa/8bSqk
P6FJF+wQ2GLgn8VjF1RYiBo3U//2yky/Zfu1uZeT/upfgNXeAkYgDBGOADKnm4Wm
wOuVHG+53yC7p3z+jtXn/6NYxDfPPL27RjtuVHWhZ4BmfO7YWOFUndpGTJmjy9XY
9etb8M7jX7ZmYtKwglWmX/H7PLQs8/3Dl1DQDIgPlBVCkU5dugHyPTTz99jgmaat
UhGdrq6pJ+/PByHdNsGHuiZ53xpsf0upA8TcecMbjjKyvH8bMILVY07l/wszqh7X
RJxN3eq3SyWcoC//DoSiLxYCAq03UDd2POqLMleHFLimclHR+bYhpJho4udKks43
L4/Ph+84W33QW6wj1hYad8x1JBHiWxUi2G+ZhiUMiZlo3gtmcfoP9DTYRKds0sHR
ag9AnPtxPgfqd1RO9r8pP1HqAH3EZMZx8p2595CkUUrKxOLzq1QdJTpVdTLRaABi
pKfcYsA8BoR5VocXFMB4/4HgeNMQzjZRQLsORQcJFnwsKsnvSWNYE/QDUP6CtldU
+GTVEtiYufEwvLp0i3g7JIUPCXJhTRlEhp2z7fKwiFjXbQLhFHu3i1w9lqfWr6Og
TmtK7XLUB8SjTGda0B2A9K6Ezj5TwoJbd8tSjBvNc2daxTTbWkoHInOBbsFCb2so
xjLr1up41kUcLiTYwnMaO6N4ZmLevBNznrVSjYnL1cILJa3lUiE6lpHPLhvuszzq
Iut/yyGuibgb8HC+JltNF/7Bq6/KQVkGKS4gElcWloB8y2xtvCRkwD1M2RLcmiHr
bV9WvE4hz52WJVAKvcMQh2redNPEfNhoeuWV0sWDCFGt4ZgHMOsKmm6KCOf3H3Ls
HYQ6BjdNVv3/8W8PYUzLs6WtGSMwhfBG4+w+PZHDM0Y6wPgmQwUQ7vB3/kLOCVZM
m60u6yvPd1opdjtPrEjZCfvFvikUDLpDyxxCmSOHRcruyJbr8cjeowCr/L49qeox
85QISCP2Cd77u6A9SWMUhw2hXbotyvA31Um8Gp9VLG+731w/ZJqlecvKwz6QqGG6
9NkCuoqLn2DNdfM0CZqTZBS5bNnPpSku9kfwsTGZbMxw3O3iIbg5J58Quxon7aNI
eZE9gZ+QbtVWYCR1BO461QMbXMkIP36QWES+fx70yw5ZnbD2SgPxRKJFlKGJTqVn
LYMKE9oQPTWCUdL/MjVRBUSXeAaOMyEHScJlSzdHuFpoDjlmf2a12FeUOZM42lgR
rQQh/u5OAlL+z585EbrSOgl7Aqyv1zQJxMtLlM9Uw+B4Qajdr5AIcANL2CDbRgSJ
zx9+6KHcG+jpjshIkp172QoM1lingzefQI5zw9rbWInbPpBNJ0lhWEFMd9azJ0xF
n1dPFcvK1lOodWqQKtzeTzL+KzJnFEKliT+tD4xfPer1nJd5MJAr5MbFeFDatpoY
OLVrzLLxgdd2lYQDSij7i7DEy5DDWpSXT4PZCtllqJOAj78SNJFLEweL/Xyg1X6o
Lta6B/SmTA4PkFys1QKD4Q4lXGNwbj5A0E8iN/tFgxYNhc0Hkrhfj8Ut8CkU2IMX
n9X2giyFE4hl4XebK5euBlXURQEda8TxgNdgO0ctbmn8lMOeFdxM8Yu+XfoT7+cv
OEurAf/H9G+Z6sUA9tL3PpsjS4I9lHtuJKgARL6ez9tQA8H/QdquAiRYkt/r6RqT
W5kRijbz1zV7vBMPk0eWAl/FBr0XdtaJPGyxSyPBu7gx9/82Uz1xJDa7sFQlmJyp
6v9K9XeAzTcwxi/t0zvnJMDd9TSAoQnsm9FiDpOK34bgHmu5G+ydQpvx7AUIOoQq
yKQZmJDD083jWeCqs4VFdUiCfx0Fz2Mnfm0s1bcPcg/3guRuC9Mgs1qYk+UnpdiD
KucLyNg08EMMNIP93X4qknPCVpr4oSqHFxVfTQ/eCLgzntDkSG5ot4Sb7+I1UAsB
NqapKRIO98Twe4WDyVvJpYgqN9Td8f46Dk97sLhTJ8tkf5rwtgqKhXYIDfSZg5Fv
QYgCQ37zdjKeLktLjLSy9TBGYJNUGfl6GHZJJlpK0gOF3EtQ9sehHUM6oMLcoixC
qG6w7zcoH33SI6/i4FMRPRke3hNrU7Bfo8Q8ItKDY0DJnH7fVCBh43aWnOnpfPPX
0XLcHKW6sHKCE4vMvQxXKlXcdW1CyiwJp+eTJaVfNI7aTUfpeE/6xjAEfzTRJ+kv
4Ssr5Ylgw8niR9mEIeW72ocy0doXgNJKyD3vCAZ1QNKbT979WecnMt1L2t5hkXRQ
sYEbTDfb4ReOTj4Eh2Rjsd6MP1YaC/fIUtPJY4zVOMdkRs+gUoSQzNpM3vS3oubY
IQ64OsramnpLDsmJ/Gmnaq9ZP5nbx6VKB8MaKSKXl+VWGX8leFPbD1d8EBhUbcR5
HkgtMRSBqOxpA5GFvB+gA+c0KEziPxIF1UDfUAYLz2X1No1UviR8KJNFfmFQGEGd
f1nX4C5LblVJORyh3/yGlPTWsdTLRWWsseoqxfHFPW4DAhKRofkQnxuPkWxY9Pr6
AY9qrCdkVX8ADIFHOLErUY6dMjTbcQPYufcv30qzR+Ru8ctmvUHUAIE0pdBxUw+8
mP2cJjF7tWfpZxTd7ydTyJKGFUTknddoQMMIgv90wtxc9P9RM2MGzyjhRWVs/Gzd
HgSaIxNYOx/zB1Gggs6buW/uQN2bB8TlBP5EjAcVH+O3onCLI/aawBBS6FwkXG1k
ijPVgkFVuhBI+2fy7iljMduMgDsAV2p0ZhJlLQo2SvgVZdT57a21C6Wmk+PtMNNA
hVtzDMcMh9huuOZ041PjxPBdjEia2eTkEM4rHbNZYOZWbPp71DIL7NQ8yaZ+TIDy
RNjKZU8k8Hbt/yJDGMO7++SoKayAPmfyeRBhiJWOOL6Tza0RGuEGfsTvUJ81ClPC
9yaV3XlEVyzx+cH+wLh9Gj2XYg4ZClkywGI/aYzPQioPUI+8DVkAeeXKbDTxK52g
2RuUOoG4NjB5g9j0iOduZylQ3KXQYEl94998oUK2AiZx7U3H1EqLtCNWaLlW4350
J3GdOvtTxm8n/qWj4CuS0oUKkHihTRGZJAAD6O18pQhhN/uUilRFUV5oBjowh8JB
rDCtB0RKMNPuFqTYtnRp+mRIe6b1HJ0H+JN6zREuVdpIyDN8lOKkGsJiPBs246zR
r52lStS65qi+jBChJuJIzpZkyp1wBKdFMaMV+K94MzLjouBR9HI7nbjUa7Rh9siy
D1D2+nbUyMA3oPSsgbZuq6SOjvPJBw2WR+N2CnAV9hw8b2wY2Fcq2itLsJvKWRVS
QmUevjSBnivj9pQ2kuPBiw4A59lvUatdar+9b6GdAAEJvYFAy5QE61z6v1o0Mr/6
mLs9H4FlFgxS2m1xDBZXPO5uWr6Y8tAOCdS81ivylBuU/Hmopt4O3WossuZEvgQR
Zyzib2jbhRolCDwpdb01n220QSM+jORZFwkW/iYbi08q6qhoyBQ2isllGKsB8+Ii
LfwH4ma2vI2p9JFtmscRHKfRlogXzvzXuXJsrW6tK03LTDf5tEZ6Fq+f2vwOwnCD
CvtJRZ8/eKTSsj7ie7ksTtdOpW68eHC4oLPJ9NL7BRWym5c7JHr1AYGpb1HZU8gB
86cazF6H7yWk0H8XGjTChFs6Y0YFg9b7SM74nemKUEfBfpr9fZKdGgqqinRObTuZ
L+lcPhTl7JgKJsGrBDSGmjKtK2m72JijJk3sKlSN07X+VTzatSBpNTCSsi8BO2g3
bpJN9Xr8aVioQ6ehOIeFOqggLQnpL5tJHMnC48+iLmBpBS8dOEd9+enKsvqAmjBh
nCp2ZFJfdU8BMNmEMfVR+x3kCrq0vaR0XmwnmzsDj3cyQ/DUyOp+oLQtwNO8EBvS
f1aU/N/DbLaTJb2fxd6MQpX0RuT+U6UOBL24/OIRdvu5gfhI28ExajuKo3Q8Easa
qjuXuGqcsXOMynPu5JsdDNx5v+bjQDhkdZsPWtIaIRyz0CQRvRxmjz6/MluOuC+D
domJ58B0BBQQr5TKDHDlWznzHF8EPxBAfTCo5HiegM6ZWZv3bPHwsCPcFUpsOHHM
7+Ceg2C9MMrttBvPUsd5+jKxp3y3czbeEyhXZyXrCIFDDQdkB3e3B3GnupdrmoQx
bP+LNOF7BqoVZOgJ7YbtfAOs/Yp5Sa6AaBg2KfUma7fmmNiFgQLmCZyMBH3mE5At
13OR4EfxWRHHom5O5WRtSWyMrYsBjH6SKI30r2hRRGvFMOCGahF9w7+HiKMpqU4+
2XOwL2Rcqb3cmkQhhwkx5z6ZAWteVtNtXgOFkF1G0F6h91WbnoOW2uq2pa8Dw8k7
DEJks4lQgkN8TGeO0pti8BexYmDouQsQZb8HoKw7Lq1XBtsp1l6Z7HgUo7AFmKOy
2gAQ/QIE9KhaU4f6dXKT0OrB2wLqeGQeeqnXn5kPmBB8bCmgk/F2mqqdcOt+rcKb
uTnPVAFYmVT8staWBVrxLW4JAtAFFZpcHNV2seX6FeJUgq9xdEJeDUOdWoKuO9Ff
QDEFPAglitL5WRzQDqi8pkcRugpTy/2QXn9Nf1ureGYYYzn0Qy5DR9d8PVNXPaP5
nBnJAK6z1V1qh5hZySg0UoJLeqxapHI5CoL/+/Lihy98xsAv0xQP/4CDfq+DMljn
1aP2FrbdLjVyTaNy3v6uXPfmypOronjgMu59WMroiyCf40VBwx+Gz1SKY/Wrm4u3
TQiqIh6zoUt3/zxot8PKahrPeQI7glhYiRdsoShxtxyH+8IEf4GPX0tDY2t9VU7k
L5Q5RQDzIL/6uU+jHqLXele/U28oxghLE8erHy1EA6XYmtfJYbRmoP5b6ahrYRxf
K2Laa2lsEVCgjsuw7XL/p5TQoKwLLBHxVa7WX5KENhMMWuluy3uMUwsUJ75pmEy0
1NSXOOve/tWbY8wQzidzknMmKmncDfVXo7z1J8T9bss9RR0Vr9/aLAKZedWEWEOW
T4paijFiaGxYezP8uBRvwP8uri32s9MM0sEMIntStZ1ONkdNwUbXIZYXgvi3Z5fw
COUzd+tQkVn+UrYHatOOJDg/GC3xB52UUHua023rmiSyqgYn44A4W1oMQ2/86FDF
C8P3TDMm7z6IYCbFaxEKRahG9lAl3PosnLfhZJRvi+lgHH6gdLo5oyDfN6U7yaWh
U1aLXltjJVSxPSR0QF7P24hdrJ/SumFyY8IzCQu8PbsOpNB+31uKH8hjUvX6VD25
Tywp2hNQmk+4mOiK5iL35DWjK0xXb8A9E//OxtZrIftPklNbAV+2sxX7p4sKuwAu
bsA7BN/Z0i7n8P6kZZCGwVOagnoXpDF0rHDrPHWIMeo1F/Qc8dUgOtZIE/JzyVE2
KEfC1CqF8ukl2BouxwBRTMPv5g0mx948knLx7zcIPXoYfdkX99f5oSWH4Gc0J0gz
FHzOrJbGpcagxPjUubELb38Mg1+6lDnxG4i+Pmgltsq/6awBFNejveg+u1/TBDRn
A1gyw4Ze68EJLNIX4yhxuW0Y+akHY0kJmRRwUduB+uJ4foUNxhyHppGfxgKTQ+lX
G1PEKr5mE26YYa3P3Kqc8RQwEbEncpzXerRyGc+3O1gygFVgZYDc4oSFSbeAOHli
uZG3hVRVvzfymkPswofC1CtRShlCaaCP9HFAariYL/GIjAUwQNK84nMlQYKSLP6u
eW9OjPfPTlHfx9Pl1IioJJOdV/gK8/vpLeMxBblJvshjxm6uSdN+QgqRzJrqOb+U
rUsOt5J6OP58s7pSzmS4iy3980QxFXz0HPM7JtvVqfrsRPh/Hkxksw6j9iU25Y2H
ExEFeqrJ0RFMvpL1Jyfq5uMw9nyI4KN5QzIx0KSJWeXOmb3Nt788ueBuQoanue3z
4hFFR4dEMq3Z3geGc3zcpqRNuNy+uXqckGfbCPxoECl2sh5yezWfvRnEXRq5+HeC
J4Ki4hEjVL0om3/m1SnRGbGylmvxzFgT4nI4OYBEH/CciWl2/nedyg6vkclWtpcV
oJlpSThVwci8G5heP+WjvkrX/aiBoo6HWhz7FFezJPheZ36/JUgGnIN4Ml8uNs2x
giDN1AJbCmVFuE31dwRj7U9e4Rfr5Evu9n9BcQplC2Tq6H7wrxUHv8w8YY68vadx
XoW4rhlCmUZPhr30NoyzD6qROXn05pN6aNIiHLeo+uaIQyvJAXBTJHxSTGryRvFD
5bju0ejKCanymM6G2Mx37hByOd4gLaDwJBszsk6MJ48VYa89W+iyZHJUH0Hgbgc/
DIUhYG+vnmUxWoTQ97gvSCsXTd2UKS6H9bYH0f7Xv/cI6fviTltf+/7u5FK9/Ug3
0K3air7bPA4i17vibYGgm8EoVfRCe/pD4roBKeuLwH8tM9NlDeT/QTNiBCRJ0SRX
BjrseNMd3lcp6SCMk8h9L83oMe9tMDN6JgzwyIFvyM6PBjmgS3F4ov1CrpA+je8K
hVUEWFM9/ZyAkEu621ghE518cQWt1qlXViQuhp7sZXS2CCRftuwVA46sekzXId5h
n+lzL/XioJhlQkVWhvMY5uR50VQsifb6zKjIgPbEQ5bTwfRgpQm6xBy00Xc1dKAS
ZdS59FXZhQF+Ne/wCfkprpOTaT4Q3ljDuxF4gtIk9fpfUV3+RyHoI+KlGxd2gYw3
lAhxkaOd4I9kZ0oow+AlTdUf6acZTyu7b257APXQA3+1JmZ2Rc8yMK+uUppo7Vt8
JpYgXegpNi+/92r07MXnxKKtnVqyjQDOFHlKLgBEH6pw3ocGSBJNXaWLZ7cZU0z2
OqJEFJdEwANs0Y5UUZGQOdPQQS6oorsoGOTJGT72kEVdhVv4uwqDVc8SnaF4Lw3t
AOFRz+xaYXaO9IFpEi1ZJNWxst/kF3mmj4roRAw5XzxTocIYls6sIVwGLdBf46LS
J/TssSv3tzJq5/AW8/6MFnxKZM120DsJMeUSCuR8OBjJW65TUIBNQfvmSDYB6N+P
8qi1FxI9ZFFQFPsCQ7i4y0UrmhHm59zbYbXI//EdVmm8Yj9fEOmI5hndDFbTDHk9
lRAASX+U1gXehLNyCTeS49ifXvWtER4d1LxyTrnbmGpj5jKvqWoxMy77caegSvf3
xdNjx6riLT9OgzRhEDjKpwwcoP+x50Rf+f5/UuerXcH32v4VRQOrEuCvg08pXTlN
J2yxxB/4/avggVlLAD6PsJ9v1Dh1YXJhR2F1Aa+H0PFIQdzjf3aRZBDMKJhBYrIn
nBtTsLGimSaHNuH1w/ZHNUhKzw787UCTxT+zIGB2wf7Pm62Bb/9EKps0Fcgpjh/D
YIPd2dA2NwUhlGMGu/AMahNTA5qyke3YsZeaC3uh/RUFuh6MZBteUKw/A+a3pL5h
tL0l2XRqjfVM31UZFM84S5sVPEv+KaviZoHpXijj/AT1UcGtAN7y+tvD9rUzdvct
njzDUKOn0Py95mVCfm5NVGm7ASVactZS9kmjSbBjvdsB49+/W+SHBmYKDuapB1y9
di5mj8elUY8nzIsXemGl4XvfYPvlyEuWSMwEIGsWR5M+Rgi7VldlCsh2tcK/0S0F
0QDB0E5mtFqD3wRRah/w0Zsl4wvsxL+f997u1e8h9BQb12BIt2eV+A5MpLr/1fA/
MtnWhjri6IgotRA8Os7MeejlYdCCQ2qvfDOLzYVQtX1yqQf8R/M7XiJZpK0dLUYN
3eW3xM8osxFcOT8nZh6uxrtDdmsnjPJXi468R2xzpGge3e2LMS2HNjwE4wULgD1p
/qCsEf8Tj9/Mj/pUQjsj2I2jNwnKcj2zPa86AOHRahPdHozKoV9Sz+x7Bc3BFcgh
o7QuYAQ9yrXeDSN7GP+7NirVAiOiebF8SoIuzrExPuvlzKvOJYc2aXJoorzcQ3XZ
jr1GtxTkwkkG+m5aZFcyUHQTwzRo/3CSP93K8shrxGAljqgxV5uftstoqfTXi1i8
prXu9gDtv2dAAktdW5jSkOjWFjdT1+cYvfSBcCiwvWrTDwedV42+74wchz0kDGz/
3i1DjJFZbF6KJ5/X3Ph/1Lc6ZdmOn8C1AtC/arIiJ+DQQEZPPdbRpMjx8i5kC8pU
kAfhlCLLDuLdNQJjEypxisTND9z3nwSZ/kd5Ftt1wgwc4OosLCtaNePPQWZkQTkF
He/0GP+vNNwEn/pUNm30n67JcjfnkwnjlrLP4SEp8/kATQO/R9CKbECvUp/fDxgE
Jk2q3JnXs0O6pdMWrA6MpghV43ThMvOlruWSeLIsLl6qc+r9TuNNn3fNA8Vu8SpM
aQoYPXap24Pz7ukTlKWEHrJ7Va8gl95+YNPXetH+508i8shyjMqXUWFCR1uHuT4Z
YIuKiqDK4da+gcH26IKqaZ5rbJWu4f1MQ0Sk1g51hXGHFe67C/O+haXb8fDxc+oz
rzi0vdd2ziXByt3EBX/DUpEJFtD/GxRWOqImrem7i4Xxk4hsSCH1pRhze1kQO9Hn
9CI3xdSfLPdkUsH6f4AAtply38ZFY/bq6aWC6f0rSEKq+vH/cqhUHJM9hzSODMfC
kfeCSXzS8YzvFuvrfsVvKkitYXD32IFOBPq8WwTkqErLORyR+Wd6nEmYceoiMtHA
CD1UF8eoBYEYly4O9j5VSRd8QeRSRQT8fIzXmwPAmqwNa4JDCHfyBsxXWitRUrdS
TwHqddaul0UDFWE9e3QXKFdM6YCwf7p9ICN1OZrQvOS/OY5i1U7Y464Tm+vhp+u4
SgDVRRHjMYlrHJkFalXwiyTWtuw3PO+tSHcNiWyCsd4Kw73520fasEsUXgYWKtYZ
g+gzynwzpOCyqudE0qhXDcfXYcDXAZEpox8NWGKLYWc0j5Ii9UtXlO3C7mDOIx47
Hd7Y7K9PneYZ184au8csSX002ACqZ2rUTFnUFYt9DjfAcsGEtZ7JzEwqqmcsLrVj
cy+hSqgwvSvX48UdXvQcbTEFAkjmbzHEJRwAPjvuHmfv7AEMGYiCDzoZ8yhd0zSE
mmn4ZWwAlN32zTk7Oy3LKo1Ume06rs0ktQS/JYrcdUfTjOiTMtmcRjfq9Ilyq3pF
GwQPl6fBJRSO5AysSeyK7ntBZwAKps1w6zerBY9+kJqNYXJkfkuvsQTTq+6gk2kk
QfoUNQvAO45fGm+iDRySUv0S0v4lb4/5AbFgqHpDzNvzJbE1kgLHsa3mrVPhvZKl
mz1o8zJ7fu5DLG4xDxy+oV93dyKRKZmimxAnsJgANFdG47EUN7u8KEY/HRVa8b7H
cYZ8L8cABz6PEhNeuZ2e9JyIzXwEi2jTpX28XIP+krCC1XUxP1x++NXnUoDIR5d7
bx/DN4k1FEJqXaPRwoGFfRh8TeFeATm5AODAvmOtFrvjplWWLdf3Xv2EMs/9QCSL
ZvHCerSZlkew+AkpC65iKMKshP5fnmcRTbwqtVkDUVx4loTSkqCaVLcmA8UoD2Ll
pFar0/qIZpbIeMSG39VSi5TQ87uJdVCRO9kyEgREDww3IY8DNpJ75UyzUFcbxuag
38dq3m45mZzV8ygJAVzvbvJ1Oh8jOJAhPMtdqEIpHHpml7yyCA6gRCl53ombxgKP
R+9nP0BHLKdHjRIYKfgNnvWrEcTmAzWWg8XvAJV1cEUyddDDDzKakjWdhgcWq84M
lDLRsKK9SF3cy0b6SNQS46nUf7/ySU+Pg7YeLu7o2FfzigBLLZSvb8mcjesIrxn2
d7iy9r2RHw7H4Frce4pvVc5sjDxs7130RagJSNYF+CHWFjYXS3qYvIxmWpvo+vBh
m39EmYhUAk3Kf6P0lRIXe2Y4HKSqbJhCP+ZXlqKoZuXWtwNaY8RXk0o0F0QPiWUV
i/FOGyC3fgqODca4n4c7CTMw+Lqr2Zx47JIunHdFKd6hWHlaRDWCbKJFvTzhMbEu
ar//1OIFNo2ziSvC5SyX2ledTTFfqC0BeKgDyPkCcfQoViOhRpFRAi7lTdofduPm
tlC6iNrpdT40Z71QzZKT4ZNM7aal8zXqW2hStEgUR2YCeSA0mjIglSogUGy2NVru
fI/uTln6fBPanO1rgj8G5PrHTCNCfifwFXXnHNpBPJ1/Um0eS5AI3Di/JWCWVM6y
9lgNya+AlNKDRWtic15Hz8DEnuHnv+5oQdqJ/hsDYpdjfsVMNLSQHtAZtkxOT06q
ioUwPjqmTCGjrOkuQRCVe0EgcdxlKkajqoJMDw1bGa+UFS9tJZdqzSdZLRvUqpk0
SnPopIcpZSIuWnFs0s1b1W9H/Z1SDVU9EHu5nMQVx2QEbUBYfi8RXcIACxW5/uSA
3q/4UId8ZSmo4kTktI5/ohmmpJbxadxGqSZvGml2WCpljdVwgCEakuECmsWTffr8
4Nl1F1B5lFgugwDlLydeJH7/EqO/qiJxHfwsumQq0RL/3LPFpV/ZJlEDwQ8gdDRQ
GmAZ0LYzy0LLrxVs2N92ECSyUC6XWB+jTk0YQmI0QqTvhtyNltSIVVPZoQE4oBPv
+rjXUCBhrGS4RPH8uDUviQEwBLDwQxUsCyqjqDAutjxLF8Q9Q3dX1FqGELEhDrfP
pI/oAIPtnYnU0T3EqAyjxfwL6dVvkCMFcbGaueBbe5iuAV57ZGRJBQwaWmoHGg5M
oRbaEPGRtNC5+AH7D6LjoZkG9KEYRf7VtvOmceOo84jGSNzWs+aNDVkVUJKaUk1X
X/OGaORQyCS9mL6kthG+s+lCgR7kRuuKcjY48rPpjkcbPk+7TKbR3B2oO2we96wP
kwyEfDf/2X5CNzYwpS1OeeGcc6tqIZWtIJa2SePpiGO760YsHoPRhfOtE5Oa4Rv3
eMHXnDGneG8zGPaz21M3GXFfgW/TevoqiJRIKRDiuJURGGsdMbLXQlG1DGJdjeOj
O6vsJzEq/sYwB9a0S3UxxpILWiOLOOgSZT4c8AaPr7AUv2Hz+AI1iLIRhrceOpH+
AXP2PJ3aZUHbROBn4EXbS6B9NOvv1xDkJcR2a3Wp222BT6sbzheU/hIxrCrV/TLd
1OtFhfYwr1GAxvGXrxIFRgbDZsXZu0gaVmp492hPlQbjLWV6UhSRMtJR3oqCmca7
3LySAQwEsQwMpn4r+aZOJDcVdRojWSBOZ+GMntPvWyakmABNBmPa7z1vy/S4gRJY
cxb+eSlIEx2xdz7DRV0G8cVODWp5Fui3VrL1avMX73pV/EOHeYNKCnuMYT8s0KWl
dWRi1IuVwBRh/ZnPNvWjHltWP3pv9eMPmHZiWypbrPoRM5KDvlk7EYm2zrXXW+iH
KPcamXW21TU/Z65xzVxb+2vV+yWs6HtLoIwCTPKktII7cUP3eY8lBrIjp5TSIcG6
V7CXw2KNQkql7KXSwFjYlIwKucZCq3sCE74SerfZgzDkaK9bvXh03+jC4DShMkU5
x7tJ00s/Kp4uSYRH/jkkue3GvRfi7qoR2CyUj2IDQMjKAY7vF5Ro+KdJyPcg3S0j
CqeSxysu89VJKuaVMbx0AjQIKstWcQUTHa+Kln+W/yqsZaFRWaXRg/way8DULral
vAaHI6DT9tJ54JZpW3VoMt/2deqqESIgugK8bwh9ikZRPGxIp4iQTRZ7TvHVByq7
Yz/rAZR9o7sBfqQ+mCQKPaSADr1FA9+xFBwgcdwmJg1ZsO4I0CaK8bCtH4SVVSwD
IGjOw9+reedRws13dPUut4m1KjopYCUzDOunjAW8dycuBa18G708jPSr3BQaU8EK
42XH0UQZcjpJq+MYbN0SoBpFDIKV0CueOTT6RHO7Gz31CLTEGM9BX81lJtc6AI96
HenpIU2+/vKgd/GItHKjy8c38hQ5CAhHBhDh+zkP1a2BbZFYeTCLu/6xuXHv1mS9
aJWK6juw3LrVRnAR1O8hsDgl7OVUqDIaCxsOVaJsU67v7ggIsRqSiVWziR5fQQGs
I7d3vogrOhp+B2bplP8GUxSj6/T2NZRALBVqZbxFc1NAnXr4kygWWk6OmEVawqfr
1nGoXKgkxvVkFSU5YlCoN243k673ku+8v5Uf2P4nLWu8FQ15Ikg9HuqXJoh0D8R0
Gg+l5BgTAQLfhrYJfJrNmdzKNzHNhMNp1JBSmBOA34/WywuhqAeIiUp33UJWeM2c
8pqgjCGZWf6xJX6uXCTL/vP8Ot8LnhQoWG+MIw6InCrQrkiC9r3NezIGAMrGlwX8
dFB+Vowcf08JKYkf1/FbmI5BZlKWuN4DhqpyTN/tfXZMaYf43F6n57VdHw1kkbRr
XtX4xv91FIZgWvj7mT5fcK9PnHrbvWgCx7hcN6RB9VTEkKoREQfZDvBHe3y630tU
NGsuBht7o4qlt6H8/Ma+pSN9fm+nfzPWxIGigHxu7bDYKlFkVkvM7B5fETlhnG1r
wDP4uAblt9ms+I/OULnXWwHGdS6fXVMHaptaNSFXw+AtiwGV9TW2BZ1mvWypsHeY
Onvn1pg7zIZrTbqLbKclnhEKb+xj4V8s0yHoE67WYsoQbs5xShms4SolkJFzHiI0
jp0iCdpiUqXcphRZJQnWmz+f9bTx9/aSHEJj1G5H/jJMmv52tFOa72lzwJRqfX8U
jwbbgJOjdZl6KtmQe9L4fcsxvFGUhVH7q/dQ2zq0bcK6ca6aAMIUn/ItC6A7dMNH
5JAeC758KOTedZJbS5pYGPRqGrVr0eOnmgvGQ9mDqanWwscrQXVKmf7/cNe2bq+C
lfFV6hYvg+9shRMFAbmeMFE96UM8+iOCea4qquFWdjWah8lGTFunBPTsuItbIm4g
779rk7kk15wTZk1tzWPx2ULNuTZNGHv7hPO8ewurrukySx4mgPCH8sCV2SQsgkCN
gmkIopCa6h3GmZVcygnsbJneRh9NiY//aGWMYw+SNxSVhCobsSF09fecJAvoncVn
4AmjX9COne2nxoVO3ZY/aBMD/9yGwYsMbaFGvsYgkJ2LV9s87fgpcB7ogZgUUqMy
8FFJDOX3m5uFjmYhKdIqI43X5Z1uCV36WG5qMe5R1TBAxX4Bu1V+524Zdhx2uznH
wMwaYuYkN9Xcwk+rMCMiN4YHdxCGrPbhssRBYCqPE04Cl7H8mJUjRSURg3T9Eac4
eGIy73Rju8/X2Hk7n1NHA+7HAbd+jkf+inGpY2mvlsaCrJvdwenPK+eCU+UfWnAC
Lud2rxQNeMrijRwNP0DqbscJ8VVWfmxBHhmknbQffp45SEBG2aAvtm2fJ171JdtE
Ru+dI2Zsf4t5kG36H+D5fOoXqZeIxRajhHuyccATelEs0WWBEhEB4mrwuDLWE2YV
4ldWwFD4OkxvnCO6BBhbwUj0V9R2F8p/DriUcZcmRdWYmbucZVUXOm/KizaxqbMB
oxKZVcngthp8nz2oHZSH3k2ru9Vtu9oAg4jxaJe7EJMmdgpSRNOoQyCB808aZZEg
wLHe1hOhIQSet1uVQaLYZvL1cNzlFl2+WZ+iSnvIn/iRAlB04mmQ+M8je8pFBZ7e
myyifWDc9vcjvWUaPrg8mdDIaZM0rjAb2J/al1rA/KAaJzIP2LBXmYFFK1qIvpwF
JthFXqP+aWER0HCn5FitIldkzakJgyJz5T5yXCCVtc1s4IJZPGwLY2dlIZp8oitx
+lMX+gT0CPQ6/2aSXOIPZhcPF14mpSTwXxA7vIpUvxs3p9rYStn8IYzF6Trl8mam
Rhu9H3r3w65oZtwGXn/XebjBTciZYYCIafvChE8lhHnPKPEFXINxA4uPTEsRb040
eGllnG6IJtu3xXhhyAd3jEdwzjPZOeC6VWUqOfcoY6J+YwfceeLTISI2Iof+A/H6
hPUyc4BdTiliisQdB2SIhQnQDY5xxJ3F9iZW0XJDo9q+zk+o5TPdTZZMlNgjDwik
Wa/lDSYy7moPAUtZUp0whttkgqwYS6wdgJew77WwuV/Y2JvCDMG4TLOYy7BQLLrw
uLMjAyShwP8aUJobSj8a8ozZ7lXAGMXHSzStmHgpHHFzukYobLtw9j+ft0RIQSvG
OMlhUM8i5ZT63xcPid6aQfz19vtgLl4fX0mRczTu7knUVMb/TUMqqob2oGdBXS+S
BsiJQHtP6k4Un8hIGTIN8lbUVEyw4wLraFQkXima/cP6YnmiMHAbq3UBDTv5/lrr
YbbkzhrqQ/u6Md2EU/bAijLHEElL/GTLSyMBbj53DZoxAxsoGl9gjZHTV4U9bR/e
DHvcJRHxHaoYiQ5dAkqq7YDHmjZcYCi9TVwqqew8l0FrDXMFfUwKkTpUWjeCQHZZ
z7pfg/pH5JQnsHZceZN7iwLpbZDevbVwAhxw5hYXlZ8URR5/NvK87+YiOjtbJmSY
vxX/T7hOz4seaaNCHpI7beiXaSEE/PTk37sBvlMY1zfXALbdsg8cV5PTXHmF5lI6
yDN3yjbCO/BjLltBSECQ7oJGqHG56FDAwveI6nZZOfq54ySOMluA37v/TLMGeWSL
nyHa4iZpkZpgfa4+vUBisVGJZiy4kZ2nirpnqOlbvRQLLpO45shGr0CmJFqJ8Y1M
D3J5Xj1xnf/n21dqEnRuNW3k9+ZicNtt95L6YG54iYUUXfUSfgIQj/y+E97LDlHT
cYuuXIJR8umN/nwUfzKc+Q2Or8s6/4JRn/yhzwnpzhLxXzzJENwSC2WoBxqy6Wbk
5LpCFH63A4BnehosO59fKXRjmv1i+2w3oFHJlhW/ZqucgFZiy34aV7ingNd9u+Yi
KfOuHDPIA8nSBOrLJ9YFQCI6/7wZqXTSIXLbXaojTy+D9fue0QkTE+43HCD2B5um
iBuHCMwxUktJZ7OA1Jj+MlhGfuo0Ed2MRveQdLbjATieWWH+wg/0234CD50hE9/b
Ez5wzDMsoDTIv1zpNWL1IA8pumZ7fLDhWkqSH3AbnGPCeGyODAQKlderjE9oD1x+
hzMXh+TZ6I3wH3zhzvmcITow9wxRe8sGheorbJun45ETywNyii8fj5IpAR2qrVgO
xp+dHYHaxKilyw0s//31+mGgR9l3I24sHPsXyDXQBvMyhy2/9gj1fa9SAfeGLHJA
EVVSe3D51ZAnooFzxL3VRKqa4SWGYbRSkJQ+yzS2b1UPnaskdHaValpJZkHAETKH
LutgqxBuOaW9uS+lPZAmhABRPWfCCMkwT7Ct04cppjZBuPVYniPebpGuf9Lx/1Ou
PwImo9XKTQScUxYK18yhNWBrk32jhhZB89bUxysN5M5+zzLEssyaJeSqMYFVY5eQ
hy9sCzri6wy6CNrMWlMWe6o3q3LRMyShaWKSZnIDqHg0BzOMf96EyXWWsWXuKs6u
hhpv4DG2VzHB2feuRTgBTNkXlsJpbPLZqzQKzYkAbmFX5GC/yWLlE6kcjIoD+WQh
feC8NRyZP9e2OUO/ze/zsHDt2Upoe3iaTqUXNvatPYhOs3Uud7bBtTJbPvRQIfHi
Gq5Si5WvjJClXektsrGmD0vHOpQtfsEikGre0zo5prL8rlTEI8opVZtQvwxjD360
CZBj/hpVMoL5+SHGSNP+580EdQqK87oi/qnfvRioFAl8OuFaKj4AEdEMvapdRXgU
Ly24zhwbuwgIOFsiFNKc7G7X0fsqecbfHluxUD9tQ04Z2FXboJ2RibqK/gMeG5lH
K3e1H+yc42CWeEULlaT/kdren4BlKtJQB3YvDvPDLAswZvIRWwdYCwavlift05gi
6htk4yVdKqfrqqyXnB9b804BxP+RBT6yzB3ENYVUNFpDU5yUSCgD8d7lM9vze0rK
Qe1bxVtNxuHYTPWb+O/86gvSQ0A8AD5/NDNHtg9fCGAT9h6l2/ufdzV4zFy44Lh3
Humb35+YbVbbDVR9YuHwOcyDTI14aainebLx95fs4x9O7Y4n3Rx3DfOODBj6/AS0
Y8EExtrWc+DZqpuDsOsOmlE6hsGLKgWfeKLcislA62Q73B+KIdLDlYAOkFsscth7
IH5Xf7yiuckRp5DXDavVrPWRG2hL20HNFCEEeaiqOBwnc56wPJ6P0jTXjluq6SWX
5QPe85/9dKjThD+WrMCZIUvWySloIWpA9IQ0WDolW/e9Nf4Dthf95eN8QeThauAc
yikNd2baKNcWZ7GopkOv1tNZJbVaj8qqff6MqpSzBdA0xTf7dAOHCw8iqQvqn5U6
AGN6799atdxxt9dOuGYMveptJ74nXaf09JS0D0PQ71s/xG4iHCs9d2uj/5zVxJUb
t04CY5DEBAlODOG3Kf/hqMGLzDg7nTwj5pVaTj8Qq9TOx4/VtIgilNoyrbJoLI23
Q8YqziU+/Hi1pK71n1be0uERvUrUk6jBvG+7gMRzzrKr4TgxpehCo6QEa96ZS8hi
pbHfk+7Nvu89TiqhQ6fe+zC6l6yMzYSln4lHBuWrzU2gvpyPqiUNk/qNsH7VBbpl
8A+tJ3K75rHBeBEg36dpw4/Vwzn56FJ1m4p16QqFyzJS+tOGM87FjfAg9jsgju4V
FNWrCGkUWzf4HQnf/T8d/V/IkQ6YMSsAFObEy9bTCiTxCYZBRKvsdbJiB1l+WSnv
tc0+9U3iUldqK5hRL405kCGC4Zslk2MtuGBE5pTTLZWG7+zkQbT42w4WoBwcj5gk
YtdIdUhXwUs2XUFkcQAw1GhJPILwYuD7MdqKl+Zm7qvWJAn4YjpKn/p+NIeB+7Ux
Fp3jhfFrAfF3/Fzt2JDvcWUgpDGbzOrhJ4xslUShOA+AkXIKA3WIwMkKk6iVcT6o
VKQ5xcZGJRuLiRsFo3Ek4a+Ppif+6f/FAVL3wh0PTjnGYSskfP2c0vkzR4E0f8y4
hAd4vv/kNYlKSjdBuuS7XATsPZMHpNS9TIdvbsmsVjuGmdq0rAGeo12uUvL7OOvr
sPzXh/s73qC0hRmqGuu3bMjQqSQlN34xXY9r7x8q1jN81CYjIrEd7gqLYp/9l8I/
1c55h3ZSks4tDfuWelLSNBH615J6IM6/XVkUPOjDfSHskqZN4y/oUgkg81WFbICt
eAm1ak+2E85D/yTFbtX548NOy1Os81HbtCRjKveI+NHdUhUWTHuUmiOP79doWXH2
UdES30AVFWvcNdj69AvIW45v/4AakbCJijkPS/1aFS4JBtnUppm+sFeGQRs3qXLB
JfHq3H0MZlh9X1qM9aJER3QDsTDoXysBzvJ53rBN4oLhNGOYvIcOM2D1E+kFatSk
f2xgZZgMzz7NA9zFtPgOx08bbItkhOPA+ks4RzUnuZq8KSHINZ8D3S0Llp1Me6j0
BG8Pd1gv21x54Pfza53bCWgaA+0H7IU+SK3xqgBhEAmgb7sUlcVc4PFCn2vMqLUF
oK8YDAK+p7E6d2BkWrtig+MatNJIemPzh8KYX2dYrwcGL2LjwG8UdbW2GW1v0SET
0qW+iCdP6l/nmxQHw6roiHsAHRq4lya46X3cqTcItoENKvTD64gELPUtatHrFve/
tQc0TW7cJgf+CNIM+UG+kHKrUOmw++HRz5LhraoviLqcs3iv+Qi1bcw2zyXY2aR8
1zPFjhWhs217kdahYpMNDiFIIAbibylvfkYMnEu05lKKROBdaElZlK+BELqaBJVH
Vkk6RimOtFBMUEYqSdPf82zhBJdZwXTkBCQVxs+dp+BbNYemY/mxweBCjh9gxZyN
7ai926Qc8IOSqGjDeI+m5J0eCm8QhgKVBj4xi7u+ZWkVnIhjCeaiqshl/HP2fBQ3
WtEHej/P6Oohfv65KDA54NsYtzTDNfzGwRCNUfoV7aL1RrpQSfvqNBkalADJj6uC
z0qO27fjySedSpARKAJ7RA4N7L5YyAFGtAh0X+bs4tAVBF1QoB0l76SmUPneK+82
Q5SZ7fGYuoiSREGmd5y7ZcQuJ2Kr6UZ9Yj9bUsKqSx/65GGzgj+mcQwMdNFcqyKU
8vs5tWGzXjhrPSrwz7Svr0cspgO0zIFZEGnuksSCmQKmY4uwN5fphvWqFhbHLMSL
KidyzTR1KDZ8dLiNKYFZRLF/Yw2nW3GFpWBoCcvQqX+w/AUDphmt5zpE4reJdoz6
kehEnFx+KSqN6FGEHxsqeG2KrZyDpB0Q2nsXoZA1419OFO/oiSG/TGkqmDYop70H
6AwB7qej0NCj99o0JCfiJJshgf4wNIRfQRUQRPeXnpTJjuoNjfeXK5PcfKf2kUEw
TFmsdQmhUGKepAldqzK/QAq53DHI26jxU2yjG8ktIoX7IcY1zd3z1F9hDf1UUtqn
UaGGAqGCIegYJoHHe7DvNiy93OXUwe0BP7KVPMHsAVaNS218fQcCVuK3M5o/rMzk
SqI2q2AEo3Jsx8uUJh8r6i/CK4OzwnDiVAjtAZ4cCJWez/5hkRFwZFzdYoFK+VYK
q5Yu8/1WZ+DVFtinjyVR4tAE7JvEPnonKAHpkIG/WI2nTEXE3gs7yHPKPEiTQBdb
0aIPG740PrpxJ3Ki327uE7kf9CT/kQcx+/cl9fYcjGZjO1nSPb8kDXFXIFMSODfN
2Bypfy97JvLzopZYTBDGpUmaAJPTcLE4080i/UeE060NCfEy4oOcpfk6e8T9Ijni
Hcj+WQZ+/THPNJAoA3V4WCfk/iud/1ssNTfeoyC64UaFAtCNWN0KwEDDJdw6/C8z
AuJA9HFwHe+i/oYbER9UTm5MANcGjaM7mlwuvnpMTZDoE4+BkW9wyXxUN3BL1rDa
AyavBnaEOREMrLYjmUUa+zOH2+ufyeAOg+dyESOiOCvupwrSXJ6hCoLKvgMdALaP
1qQd//4lzcicuTKaBzUmWCKNJFY7MORwWoW7Pi+M9alsBeZmmbrDPXRx2xtvIJbr
ybXw0yZGpOOZsqiUxOkgTsaMNa+0xactsbPeROrcOixs62c8yqOx1tPLDz4ABQr+
tElJ7co/y2ZcOIxM9wQgishBLSDtdOpv4vMyeHQS6EzG7QPZHp+h99gudt9Oy5Ig
ImuttrdLnvpnR50pxoUSOa2rDPxtlBPae3oZ+1eHrG6HFplF2QU0I5r40Bwvmjg7
+YZteAVFNPAd8z3htCBScMevjg140Ksw1pAV4anYdPN62wiSJfcM3OapHdiCEly8
ygZs648kOp1nfz0c/LRTmD527yVcGJqK87JkWS8jCqnxQuMwTTBqZQZ+PkiXHG3W
508P1RogLUdvk0sqjkGw++VbqWITOcXdCjl3bt7SwDSPZZeMw4szqhb5cwzJOEef
Uat+lAZhJ1CqwbNw3AjJk12MS481BLXpjGtkKNMzEMd20QhVuxoX17z+5NTDihkK
47QY81NDteStmxmL4T/W2bWXOBtqyqZImYnNL62nbhDtjt9qMyRvAZ2z45ACRLKo
SW/hfZWIUOWIZpiUJIMMXZyNeXNXm+lhOQsJRZrN6MxgBVknfIRL7iJroBNjUxU8
F9dckK6cWfeWGSIwgU+K2Wxsz+jiMu9Zn8LBY0j7wwvdzrstGG/loQWhsXfrnv4j
MaDOGjBN7koMPhKLcYFZfMQFiy9KCa+mpPZFuMn+IA2CJTt0hf4talOWDmKw+K5w
EMgGgPyuwuus+4fjCBMAHiajS2pnYALd32dnLJO73L3dy+HrBmsVpAIUKwzFYTYX
Ro4y5b1wDj4T7s0ek7Zyofpir/vjyYsQw2ksVWxhcoy9zzxcZIN+YnQ6KMawZAJg
vO0jmduT5yuIM5zhckdQOrg3b4YHgAADwOnELXmIaE6+vfdcyv1lw+40XpVYyqWs
VcPhQ9g8dBrTJTBrQ7pyhJfRltW0djLYCBFHGyR1HCNKNJFN2xuXthyVNsw1ZVfY
xOhthsWvPE9KhSIIeBXeG8qwS0+bssqo+xBv2TQntmcLCVYqxLghWgDeadOUI5Oo
xy32FlRVoW2yrEoApyvNB1F1xWvjU8Iu098A2+vEv8QGc9ZxYy5OboY6TubzzPTa
GHC5+VbAjfzuZwKo3SRp7nhnUBmWdoWGSiTXSmB1rjR0PhGBxKvXdjQPWXfcBf1t
HYfoRTWxWyb9Wz7x970wC7hM5ymLGgD0qvGBy9Kf4K0tfLJj+tgf5MCVKpqnE4Y1
gXp3Ot1wDudI8DwT2Nu35MM0JdfSl0EVwGuIACMJ3sqpPau7r0cy3Pv+grLSqKmO
5OrDPnG10S5ZzR6m8OdkbxJ9xvVn57JoDTrhGAX6Rytytwyr45qxzQpGswzIKwA+
k3cSLvUtWebppWue1rx2TOeVpXHRBFzb/hnhyGEU5ArkFOrqzhN46X/0Pi6XzXYF
rahHtOBluFqA9x727dlU5dcnVBdCNAGaodUlau7pGcB0bQi5vhXS4Kg2l3371Qyl
EYDYHTGDVw8vQHjXn2pmWw83zDnB4lP7XN8YOefqfXQmVAYMHQWv/6gnzoTRtbYx
GWVQbUOsBCMMDTbp7cnzACxObeKxniP+eJkybvraZxpv8QNOJeBilKWM7cYUzZwK
mAZcgnmUBBoSRq8WCgG66EhhNo92jk3AYuUfIL6hYxwKkUIRiKva0Fobh6i7gTCc
eXpkF7HJJXSlJt8jTV6YmmeoRX/2uZUZDY0L5mClrTkdPyk47uy4PmJpb+IltX17
SRC9Xq9w+sfgPt3ZTA7lMy1getjgZXOmgDB5NsUA/QHGINH1TEKD8sZBPCGvu0dR
8NxuOeoG0WX3vTQlPEch24cAjgwUQuvchNa8oADf1cWiQ+ChnCxZovlPgGw2mkXv
QW8CoiQgvXIy/AghZwlulyNXPMOu5e3Fne7TydGIf6VqNArNN4N2fp3OL+iQdp2b
XzHRDRMICwaLyKDqlyezU4azqKZIaCiEGHmOBlMlTukOtbxYBWQrqXZhlgOXYOrz
E/ZCcp7OVwSui61mJGL9t66/38rnHYQzeOB493hCAiGJXXVHyT8Wb+XB0rOXUK4p
ZzeO3ZcEdVkisvz2W+GXOrZbgkXfsi1+3ngp396/1sLil3qdvXUExi7m8fldjdVB
pJm24rU86AQF01bptIJx1woxrWUv+7v5OHibOUqs1PsolWgaruTULswWeSDxsDQh
1CF15MDuoToZSKy/LuCGBZdX3bp8lZj5SmYNiq3S21yUckzX5ZB53at0WZRUAh6k
AzyTPZS4C+2330i9DcrQ9CnyOWuPOl99+1hUW8gzCgAhiyZbbpG6Ao3eUKqt9fEL
L0WvFZ1lD5FlU1azJXzoIEQs4qu5OpP1x/T43MCI9Rj133b9eXEFI/fGZ6wZqxGm
jUXVpt/9gjVof6C9KH3xwM2yLTso+01r94DZHzcgyqnx6Wv6Bk++VJW3YuqDPWeV
66Cd2gtH5LGkMnkREUuNmiCfGIFH3rkbXV8+VYjO+Jy+0Ky8gsAuckMfYAie+KNq
gOV1Xn3FiUklrjanoyBSeQwT+nBfP+fknJnieYBQvTtcjJafWFS+p+QIV54a9P15
Dh0CqT3A3VCA/FsEtbSwEFwSDOua5BV7JStSi0wTqQPB902px6wO6Lg7s+SOe/i2
e133kCOroYhYaXNOl1u3rg/W4jedOI4wzRYSCbR3cNs1s9K7MJkXV2FE8dgRabKL
Gl0aBRWh2XSw/h86uDlfybPjKM6Y8eJq5SCbMgGvKGxBjCCe5nBhT/09hzRCcDtT
Lfl9I4fAIwqiINj8SroXz0vPruAQeGOE84vYTN1vIlVo8CuFJAUARc0oZzWg1Jch
JEwVDIBfr+/ln5dSwOYj7J/iITnbdGdlUvm/celO0jngooNPPSzRiLBUIixP3MBL
XSNRSMfLX+AJaPfIflI+zfmnc6ucz2wGAsKn/DywNPBXZckdxoYPNGztrV6aEyvx
lVzZwOuteeXxCNCrJT3Mil6z0AW7pCrgJgxtOBRl4wphAFF1dQgOm3D3M3zPmOJz
uyNzZYEvmeW2P2HLugl2CGrzYeR9MmV3pERPfuMU9Z5fFlI0JqXvxDLVsyhFIvrr
B/1YIxC2cDDoZtLQyDcTGxhoPD9ugsZUMPMi4b/xhpVuhhYhHP2oLE1/XPonFv9M
tKOb55eSRqZJZEou1weB9eyLKmkRQ7ZLndcnSA7z3bZ57fNzF32txg4KORc5Ppd8
HtmggY8PppqA43tus66aPbp76AGNSIaZFNfymc31EeE5s7G7ixHyah3jO/s7N8Ax
B6rj152GeVkNlicoPh27+9UJItoCEhlUMkLLq6f+p9MfIXemwq+Qa8Qpqi/JVaSD
3vQtGHmuQU33BssfLGm8dVIA1airTrX7io5fEm+MaeFpJMY3n2QWnMgl3S9Fe5J2
ugkRqLpRKYDrXK5u2vSRRTb/Z4UXsEklAwy9k8jiUqBKiQmteJZG8n8xVOGpVtFb
F2fQsM0m7B/1AW7crrn9dyO5vQMe8V5FfA1hjr3gRPDluoBOjdfy3SI7LEn/O7o2
a2Ge5/xdS7bBHVqYHrMfDPCOzKYBro5ggDbhyUtlqcwh1K0KioqySWUgDyWwwFgp
zXVuelC61CCPijH5ag/OzNDSi7sg0cpSV61ZFuGUAdky7/HkfwZ7c8JWP37WVhyo
DRKlfZ2WGzBo1i6z+Pv+PQuRwbygqwi/cZl5zG3RmD1xXeIdX3woJ76BK/l1EgEq
aFM0PTOwNAHzoEh4HiyoSY7zDdzkTNTbO5MQPrCa6PcSXfbf/FNh6ot7/NfDLN7X
ux6iLCyczKwuDeNsp9A75lvpFaWTTJ5xa+WTcMrvmjA5usEHho+MQGOgFAAfyvFm
Qvhmo8OlG/PEXBMXLM6VykJWrm4ymfwaeKJi0exOZfeHKfo1Nxs+lHhEOYFdjLa+
/bb3/QorypGMQjYFj3/Qzn6Duhp3zRoxMBfL56KunY5I/+dVnprdFe6Tx3NRumun
oS3UNGDDYYMtnYA3rXCYZ8avrR+lKvdjAyjuupVQ/L2U131Mn1DdbxaAiEyc7YTd
NaDEaBAf3Fs5iFvRSoteoYQJUiq48OS+FZPcv9U6wBW6fL7Y+T2t7K0WTe8ff1ls
PhkIpRX/itvRRWn15CbljTLDDb5Bb1BIZ1r22jcQG/AkMgMfR/qkemxKIl1eMot/
zhVMPEah+KYXCgE411Z3W4IKydXa5WVML9XMrhNJ1laezO/rY0Wm+UI3OWavTl94
llK0K41keePXswoTmErS1vaklXFs3ONlwzGIY1Xd7bBm1VK4hDMaHR9mtqJe0dhm
Tw6ghZ940Q6WgGmHzjsDi14VEidLgBRnsvOfu40Gl1gsfPf0sTG2rDMVrTgHjOPO
0pp8aF86JUYAipbjNzTdTuNsf+dhJBfDN753Sc3JnFzCvBIN4yTAJhZwAdzWTcJf
weUSYB3firhcyEjvLyKmxfM1exct/RJoZD2i7ixOirXKy7zFA7esw1FHbL7IqdPZ
EghhTFnudmlkKR3H5uPozF2/9LHgd7Nk6yPSdDpErGh8pSTfkcWU8fZ8ytvJpaQ9
cPYe2ucH4BbxuQu6/goOnIHhl3bdDnWtSSPivnBvbjxRqDK+2lZDlb5BRrFNdzAo
5aurVcPET+8ku+7G092NSJgVY3F+hACFdKXKUAVPSPDe2+Y0gwQc1sVVpu4VnXRQ
fPkkbL9JAQfIRgtXmsZIfenKOOw44QGKxTEXh5NjL3oZnthp9OMiSepVcdCg3fG0
4PA5d46+/Ho7cLxb2tplq05kE1lPYlg4TlyksE2Y2lUcyQWzXTx3Ys2FCPiLWZvo
WI7R7jDignoHdjV+EozkQ/mr/7s03aEqtFOqw8VSPVbIeEbshBDtyNX77L6vZ3yY
LrOtu9g20ZrS6LoMIbO0Jd/cQyl4/5NpCEsrHEG40VGyFGee/LWENh+6/uCGeR6I
h+c5tY/Yyq1/OQtIysaeuZA8RXAQU4N3gm3owbfp2zyriJdW5nKz/uwyD1ujT4vI
reP8U0kyHFttKxechDPTLRtooZiUhsNoOdfDpftGUHp5lEDDXjxOFb5as5HpwE4k
Vi5XdjEI/B2jJNQCXeCIMtyjtIiArgQECwMfjK1KTx9MFpLz0c0tu3iMiTU8jZwI
92Nmyh45Xnjd02m3fIOVrig/tUh0QrHvKIwV76r93CAQqxTZs5SFJ0fI9Vj96VVw
So6RT0+KmfZUdFgYCupipLNsMSdDI8yyASAKr7hQ9IpY0RyTbG/8+lURdZczUyCI
yjgTcwd4SZWNyy5Dka+BCd22IPQrWL6Ukl0qtnO0JzHckR2B2lRQAjC5J9xfpAJZ
qwWos6BPJzDXnkObm6X2l68GCjd1P/T0VfNqxT9UFOjG+EEtAkVedjMY8Mf2l4Aa
QQEhUWPEvhgHjQk0iYT6lUZJVdEEvwBnskK9pf0kElJoyhCslpw1L1kqY+kgqi9O
9TkB2PO7qIRpMNs3pKqXHZwRYxsyGttT33DpMKUDhKU2tgu2q5F9si76vVsM8FvU
2SbP49vTgwIPjiSXlamYOJ4oXFFa9vOQXw4IF24jReZHG0m7HHDQMATD/dh62CRo
biM45/jTJjgLLEewDG4WcdnWGs8o2F9NVCEalezCiO4CRCBy1dqD5Lo+zCdkkEq7
aojIL0o4rOGIFspJrvHGmiAb8/p7Hzm54TefS2uF6a236tjOrphzmiX3W3VmeHTX
sbORn91CgvSTHOXkdyexz3GidllCfc3DM2WIa43jlz/UMBGeWSUzjDX513DCg06f
/DthDwtlduufSs8NJuSVgO0pqJdCPueRtOC8xEqyyDgrHNX5qZ1DLHCp0oB0tqOn
V8MvC+EnCVvsw12ece3T+Y57wnEn5PQ02/RqUn1y6kU41dZi/f762s+eaQCsf8ju
815SNi6QxlVu4Qr5Xl7RRd+X09tKsTmov7bwmjPtN50a31OJEtNJvUqmYTaniID5
QINQ3oZ0PWc+/kG0lNE0lQv9yWf84+w2j2PSfCJUOplnw46s4oAAHgZlFgaCCD75
YAnYdi16v+lTUUGdWkBeQjUxCKAl4E6QTf9TQeFaThfM73wvOnmq9MTm2uPcQIVb
+ELFzTIxzRZrXkOqN1/jufNAyXh5vZqvbXYNA9X/a1galWIrsghxyyRE9O67J92O
9HVN1eOo5/AE4zANZJKjBx9LbR8GjQxmhw+EQtwrjL/aRkGZE7txCLxC/5H07t86
QONu3wEQkhUTUJ1Pf7IlM26vuNVmVPIfGUSfgFDmARIYoF8XNhW6uZM3DZFrrFfM
N20ZJSC6Ok9qVVqlQoZxYRlxYszSQsQnHlTRhYcxosFVmXM1bdcfwNgjQtvury0M
OXbssRRvDqHb7fuSipDcZsH2/smEx+R6lujn6nh0xQlAZ1E1tvmW8c06z4uKy5nZ
EwT9p4vDQ/cuRRUFfVob4NtYSnVD0pvY+VSgEaz2P3hxEnY6YTAFIPYsPn2RUf8q
EZDQRYtDJBr1EtlN8+J9EHJO6vavxiSMEtIgGCKnTDqkzdmScCfP7lYQ2RRHcdUv
/lNFJ5Beh9GQ6UQiw/zmeMITSL7fo+8OegRH5z3j2B4M1Jks4FKKhAEkylt/W5l3
0r9ljnHsYE5pMZtfyoBh5FWLNCLf8t9viTkdJU05ZXawsy2gYbtDj/Cf1vo1SP6P
oGLv+hovZdYgwe/VnX+ikfYxsl5AY0HTZz791nCAvafRTiDMYLARD1DawRrq6mws
Im4l7fxypZWzIUsIo1yJxOXUUasjjO3IzQzMvzvpCt5OPYlrjNIF2OECwblhJRYy
Q+CwbKoWUPHcfzkaAPoyDOGST3I8PwYlMKOX94L3T72Dx6pB7b/VTYAZ7bR9t8tF
Tsk9zB4wKqR6w0PCxUpk0TWx9LOYwvi7CEf5pYAigYcm3pcUtF4GchirfG9BEssQ
D6GoY5H+oj/LPHkB8nkKxdlji41kIfbA+Ay8qjFkunUmonO+cOwQbbh/0CmH4pgV
mCit3vqS/kkO0ww+l/DzS83Y7JUg01E8IWJK09Gm964Spu5dRTy/nv0cOrDZQX7z
zJaajy3ghvIItQe69u+DvNHDQSyHtIwf/g8K6KnhzfuhPg0ctuuebe6Ptph2dICP
vnMuym/sY0wx9XR4Vh4HVslJrDJzfxzPq1UUWydWFfN6/pxSLfNfX2TfoE8G7wTC
r5GN4JW22VzXX9gsKpDIO+VEl2lcFMOrmaTRw9VRqp3kb3C1RsivaO8mOFBALTnA
85Y16EW4NMv0VVwtJobAKSizrOgKct7HDFs/1/la35A3Iip73Xp1yjMK2TA+Zg2l
3Tny4SH6YGnv2ImxdoKTUtrOBNVnCedXz3mXij4ZT4kRc34kbkNF0+HwhegDsDwX
SRjnF3puCLFEWOdrCls1YsZ2w4Hu8z3+I2KlENJk9gJWbs6bfA5mnnd7csK8qDcX
afUsRcgUBYmx9YD/Bb+7mm+Vu0H+lGWzyUWrR6AxQA1sutaSDGojXjIQM7D6yDec
R7XIkfwqtAYTPyMjxhdfmphT4s652NjWE28H14vULcQ56H73NgC/puJY9c0D9Mo7
PmygcUCALh/spj0yBKIteHvCcoUlCPJ39DW0DvFJzvYBo3EAyKNl++dfT/VfG3+Q
LLlYz4QhsSX29qk5WL0n3Z5bSJd7pBUMC2R9X46jmAlUOp3mwy5BCIMQVFbDc6oQ
Sx0dnKc7W0oYRIJaO0dRLQED0cEibX0wiNHo5AhH9AoNuvBH1eHwZEXUgq3doZz0
ksNS+A5KevbXDgv8uGobueO1N52os0uIBtvHi0I7o1Isv5kZPiG68E52KZDWTZAH
SfwOXIBfmqPT0dVh+8WthcFgBra9vXxnUlcOgTWIDP7yC7pA4YX1ge+PpTQR0jb/
+z3GKcyO3FN8GiI83HgDQ8bho8O0iBCrxWaqHhGh1DYRaZYkeN3YgC5Ue3VuYh7d
6AQYMH4H2t0+zHoUbiPsqtlRLTz1zGk+pV7vxbKFCD4j2Fl6KJLsre92V3r20YfB
zoDzGW8zAGIoiO7NiTAPsh0FqVpwRtEnER9NuXU3xg6T+3lAv8nPphmhjh1gLg/2
0+5IGcwcjgU5ziOCwAjlcHwLcXvIfOp8qvvrfiGu78n+uIgmTXC0IRIDHO+EdlVQ
g9WXC0ap56sMOzanl1ZxIJx/FA/7vjO97TNAGs4hk7SRTrdxdEqLXzCu/AmGh08Y
PYXB445LYp0DB1ds4gQ60t78NzVJOqWzDWkB/NjGzHhAyA3+xRSXi59DquMjo7TH
2KfgP356ohkU0nh+S9+00dLV0gUxr2fBO7wzF/6WIhPVnrwAfRatX7OPsoRZt9CW
dghZDzUdoWY5jptXryWB/RQRQ09fqw2MB8x829WDyZtsqjOccBlZBUE6VvS7K2eH
tE2i9BcqtlKwVQEndFT0qOGTVeznNytjhQKbvlOasPKDkZGLpst9p1L5JMYlucvx
14YUGXI345HBHLZWwvYeAjTxXU8jBqkUpjbw7vE6n+CdZJUrEeFNZc+jmav2LBk2
P3aA1XkC4LhnwDPdAz/vSR03B2KKGam9pEo7RHThqmfK3zxLf8+yJnG9s7Wh9cBf
wClDimzTSGksIkqHfN3ycledpVU15SR20x1sP7KchU7Fp5QA8Qi2WpMD1U+xHLvC
Aaq86mC/6tyqbry93cAzvsXulETJxIXckCKX3HwMOkgYcFQfZIAj5YDO7xsGWi1f
h7LVo5b2GbdQbnq7Z4uQ/4UpudSdKNDjKyILHenOstsOHO7OM1DWDrbUwWsLuA4H
A0dWE5PLG24+EsSExCTGQvEYLrBNX7DlVbI1x0sfBY78wMp1L87Fws69LNX8KEHP
KLPQmvBmkzUzrcBafESwlj3gUqYMQou2FfYKHdhCuidSI1LEvmbDRxe6ZfSSiiBY
dYyffFL1ANaN2RNeZDb33Ok3B+kXx8dwuk3VHf6Jh5adCAMKR6Y4EeqZk7VkypCA
9q3W731WmO6VjC6oz695ZzLs4qK9RZQ53U2IxKDh+LWdnSacdRpy+hn2QDHckh87
eSIZCthhz9eGMhScs5VkuFj4j9tY6iLY0RDGzXubVLNZp4Y9U1qWf9WmFXVFSLl1
OMDFmzhMhaJdIsO4m41af1OS2qOk+TvPdmJSvaV33gsmmrFlyLMTU4KTk+U5nboT
O7L86ZcKoYpqnWtZbd/pufmGPUi0lu71F/cHqEUjj+SuptU9/5bskFIMX4oLzCSq
U46OitYlsCg2QRnqCONHWc3pJ2547FlSg+OZiMIUbHP+kvPG/K8Zcl8jhXfmsn+X
ymnELgdsqDV6GIlVtO0gx7XRuqWt2+aGmQ+UCrAbvD9/XxruTC7fjqFdH42G7Stk
oJqW+gdwClxHrfA9PF1uGnvELFklNfTeaafLQmqFbNWwwTKqxJ8CRtdP8m0+S+OE
kAAP3XKNS6cUziwqX3hbLpS83vy5x7NoqpLhE4gtw+AN81K41KW94J5R+JCChFvw
m3JmhtPgU7K8dNbo/0SW1cTlbia4RS52lODAMBcLscjuxk6CYNvp2GHbXrVyyG87
FPpUq7VvscTaeijqpDDfiT0rBFfW7X/PK/0niqIGRxwiARO+4Gu95H2dW7uNYBWn
PA5FrR7FKWoOdQaCZVYKi56+YHmhN65FR7jEITvVzEhy9vuvX2cewFMWenHMmTyT
HapLlkQNHJOgAjTzLPtHwcCYNoc42Al07KeCSXISACVLU1wVWFksV5v/3CI0Oo9c
PkmesfT+SVzoE/fHLZe7ztQko1M5IjEBQuerTylTzSbcwLqy4nTSUuDIarm2RIL3
fOic+becQnvxaZbPKgQwwUtXDLs1RJVGdqFH5QaxDmYcmrhonC7yVvX6xlPF2uck
ybGXJ5DOhu9Iy23d7oVjFH3SsDBSPWeaOAhV+mdNVFob4PGVfkncYNjxvjPbyhWs
GGq0SEj3Wa0xnpCrQ5hwj6F5ePKQZdQVUZYxRTkIYnfOYGdPsRwTg2c80l73gxwV
TXEfZB2xXApChNqqGN2rHJ0ehhSEy7c5SrekESoaW6r/p3UeTUX8UDLxmozArxF6
/2XMc7eEEEW2zvcVn3NrS6NUAjs8SmqHty52TpKfG3v/OXnxESNve1gAbC1fogO/
jTziM6ZAij34eUYO8B/RQfAwqH8IxkyIgP00SYRcBAJfykc5gAUmC/ChCLZ3crow
UaPGL5ocwyH+ILAJg8hC09yMKIqHjupYEg0Qn++vrIqHTuDhVTCmyY8RWXI6gJVN
88pH006FT3JkqWrzIdAJmjEM5MOsgdP2HyIox4T9UUQWYUdmRh0PThxoAzgtTxF3
oemvjfXwIuSjVkRWXuJMsojpnLSjtDDdcCupr9+1sNybdlhfPNgSPyNbzbWp3dvO
+7tXwaJs504grQngUueXBxl+VFChCBZ0+gEBRgxZlVdfwLc9eAVPeOMCtJQd/Uut
jvrG9D9x0hOj8GiCieh6H+tLb+TUIEu8QMUPOfyTYv2Rjg107lSOXrKnM//sF7Rn
8ftJZKXoVEBSR8AQ2t5LnnumAFaN7QyOV3O3LGxfvkd+e0dtKCM5eTgkF+FwaBRW
Mjn4iAUUsnnD8qt6tds7W1c134C+UgQFHJRVxf+Mh0GX4fwZTkgjA2qoZe4IaBx1
NumGmhCM8cY1QLG2ibNNzj83Sg6X5YbNnvdrifFE0jlYjRn/F0cJWcL8hxfAvBZY
/BzQ4waLCVcrdVH5aJcNlgIVBxtQiC/iKw5vfrsOhPDd9TaPCHtOxIU7s+0g1TXS
y11NNNo/EuQ8WyOx1xiB2IQ3IRGMNK+8NUNLvzfSVmp+2o/zvrvE7LRjvh2p/tLs
yIhc9tHMKw9NTGI57iGhMqtDL/dd0uQEm1qtKFhHkLQql95XQiE9fxB0H0u9Ft0e
b4racs1jbA+j2XShJ02BIb5zyrq4gQ2p3Fc/zi5F7sH/n5abWfFW/9rHerKwdk2v
kUe3mCfQgCSkiZ6Q3Bi1PwMuRE6V4WM+D5xvOjKretkpduoyeEQWrwM94rzWJU4Q
Z7P0oNfWOhk7xelXPAudCxe9XzjVjdFUtt1JWK2tkM1RiwmvEGpWnmn2dcx9i6Ax
chnhINoDgSyg7poy4wREDqggQBr/l8wl6bvMp0seNR2MpMRYQvbYLGoHGcBxJivT
cWFdwbLa/guPmk/S/Hbwp6XEhGObCqkH6jFpT6vYhAib/DWGWzaWePmG6CiA4HmM
gTKwvS9KehA/seIj9I8g5v5IcH5E/DjVjX7hKC5YyP5yEL6b2r6qIAfUZlk9dA4+
mwYvozZJQ3RviHZ98WIyiJpLbt0/kE9SLT5L2rnxrGKAoLQ+PTTjQ56NxmLAxf31
ENa0uWiXm5yFLtono8wIWBzrDaFZICAGH3eOTlE1V90PkTyeWstkJBiiZMBXltzK
e2ObEulkzeppl5TQJ44lBQBi9G7341vNk+m1oMeilPsUtQru4YkHhzFAPpu2C1I/
GC5cy3gpZcR+rHMlXPCz3JcS5omAR1nZxCJDsTwNJtxFg031QW5+YVux4jnFA97H
LCh822mutJKDaYhowMSK2Or3i6s6zrQqicDVzbHUjWMippFkVvBYlauz8xSV2rma
f5+tuSfuZiiSbtgkjoCUt/dtqPKpLtMw9DcwuJ/YqyzFl64z6xuE77vFmW3/MXOk
o+IAqJ5dBIHgbiBFlJfHHdpwZoZWFbv6Bg2IMNelDX6hc8rGo17sXV2xW8+GYsSi
RCI8q//31iujJKqIhFbLdxTMBio0OrjgLQmNL4JuJ4xlG0Vv8rPFgajSDlQEOHJM
bAcjH17QzpjLRi0U0s3YsLNs4D25owrm4WOhhN3P6Q6J44Z8leThE2Q9IintX/rd
v07sjk2cQD6sJYS6yAw7PShevD9/s3cLhhJmoHuI9TyFqY6DoMY/L7HWGHuyuLQo
1IvqOabKgp5Pzg8Yl0VMAXNr3XtnsgZ8+mx7XKqE/ftIAYux6FbVTBjDXWj3IYVY
Xz+Twf7ywVtegXMrPcGPAYV3pdraZ8qsHJgCTRP3YHqQCByroHoMFkbzYb29sB2w
UIx2rOq6TR/h60RhtYrwSKWZXsIWGT41qpEeLr8dCUzfNjweDZc1wC/jwhniS3EE
JUBVCUCR8Gzl8YaXI6AglVv4LJ0L0d5Wb1n32ALUKvdJxc+WYP7PS+9IF8s0lqKj
Ycl++ky/g0AGq6BU8oSwS55yZpnIjs/t6SUKN50F2lQtzf2HLnzHb0K4G4RAaL4Z
qEURmhzWp9zkuH2CQHrNcVbXHhusHLE92Siv8+kdS7qcxps8zdkzhUb9eSCgchtZ
DC3skNZZVkTeFcFZXgxnxdLKbEz9u4oGgmCgeYM8MYj/qB+MbJqiaqA5W1Xn+cdI
5+06hdqWVQc0zjYfXG+KxWtYPRV/9mr6B725GjhttVe/3eLTR396xa5vNvP33ym6
EzIxnCOtj/145fEN8CGrNx8VeM2N6bh1byVgVfocQAJfIiXjn+zMaPHCBuNf22Gi
4hB3JqwocFCJ+BSWBLOPI3eBFSlaTo1XB9ru81tYpWl87a+hbdx/184FdYCShtvU
BGOn+6Edr0a20LDd2XIbUGpbJTTFOk+A/jVeaUPx04Rt96f75ixxD43HIW7NhKGT
xwm1ryuqj254eI9YsZGzAzQAA8PVbCJuzZ3LIiC62o7lZnrIvTOXTM1CkZ8AJ2lQ
svpWoaHAE/QyiPL2uzNC1G6Im5u1z3DgvnJERznEqod3mX7UN6Lmlr8btdbtQNY9
mK07kqTryNF4yklW7h6fyErP0V4ynKygKa1QEr8FLNG3vrh9La9Mui0siQcECedo
ojgDFYv1lVWvtcXPZ1FPdOnFLjhaY8luXxp+N2yxCCpOwJErCNzcDPBcmI3SUEFx
0Lbb+y5t0eiaSD4NPSZ8mGclytxQhCGzqKWlZio8/xCiCS6n+tlfQrnuXsJdxRG2
lHN1SgLrl98Lp2Vl5N5R/53ieLl4ICaZCcfqgCC88imgAEbIdqA7k1qWDk9LJhV7
L9dsRL4DdUrNQb3NZfuPBBTKnKsNnU8Dfe64pF9Aqumd3AIIONVv5WmCcmIeafWu
Bi5lhkJjpSW+BV7k3F1bTegMyHnbYcMwQ6+NvRQ6LpuFv8xsm5G6Ht+BeHuuhTTc
MnJWljcNxPo+zKMLJmx5btaDgnXyn+zuuvRhPcPUdzudzwtrzo08ATHe6fjAV20y
Xx8kw3Mp6HOO2eHUCnghIyYwwluhFbItxpbu2XnmL1q552WIqinatC77bIPmHuFp
uMxjhlUQtm1Hyx50TsUQwNbGSFyo0hFI/5NaeyFhOAOE8jPs0/gXCGF6DQeSO49n
1xUtTRqD7CLZ7GO9fe2lA5rFxidmo4++zsJFN748bHDO7PwQ8i/Rtpdxla6zcN0N
HEb9ji9pzws7qviAhZzMHCGXfLRs2L0UDQYijVnX0bmU3SwNHvzruJuQwnX87B0G
xn85gP8DcLmcyBWCcTO7uphzn4CYOWvbr+oR4dxn83izL+/3ta+FgP107m8P34gL
MYyi8xHb24QE0D3JRYacqfAn4VNAGiEKAvj4r+MSzlOaN61FXqhRZEfneslfDNDf
9AaCEXCMFZdrcBbUNR3wM+XddYH/aOeHI5w4LhmmAYI99RsqCer0v3RFUEeh7PPE
YDH2/tNGFpnWD9ub/k/EeEECq6gpD+bJ3a2RBBxrkbH7i9v7j4Q04EpMu0Ikt4wk
p+UnA9txMw+2R3EwgK9ESO6PvaTiacTnpFTd501V6ZIWKIdHuOKZrrbwWIPIVM+v
DlhL/JoYuI7lMOEbYYWVcgqoGQ8J7m+U0IcMnLht9qLI2VBV2kT+AovzXJS1SQ6A
xmOCZYAf1/fvlTDLk7r2ftd4mLSBDeALyQ+eQgGihkNUbehAu4HpL4y2mQ4ICnvI
27Fvjpudk6/qtF2iq57ZbSDP257JeKkyRlYog/WnFNYaleQDIqbdCUmjXAaRndLT
gsxXu3S7ksQEh+ZgpuWFStty+FmZ647hA4ILRuPeAIeNAiczo+b+qgX6RZW0KBpd
FbLYGMOS/sLX+nbNwAYpS6mEOZh6+a4MHdLj3CAvHt6vod9m9Y/W8S4Mt419XiyM
/43/guH/UglW1Av2CljsxfTLhMfSPgLljph/LAImX1LQZ3/Y39McjB2LCkBGwBPp
+pqCQNVFawj5rGmXGpR6K493VTZL8O5Pj2JBdotZq4sgyWSePVs+tLbIKCGYChJH
zyXEk4sivFoazoBToyLp2TAtBYnNe9lWqCTxm7Hk5h/rTWA4pZt1evAH174iw4bS
cLRkqSyBcyWfZ8nL0BiTogqxkEdkzHqhXSaNzUJSVApbwAO0m3Qnye5d8fPFhAKY
RYp0OFHcfujBAzCdx8A+ZSMiRHM0RjHbRjkD9IA5w6bj54YjdW/9+pFUdbxAgaPk
DljFwR5hFGJmvsSB04MjEoukD3Cj+peOPw1ZAxjqEdS9ilb1eBeIX1GzL+HIaOC6
QyudCYPKdn2O0p/XxoJhjm2brVayGcC2bFUJdD9Hz529pPsCZZbbi7sUOSV0PP3F
ZxuaClHDw0bc3nFS9z2t287c2Ym2kFq2MwgBgQf7aiJ0aO7ykxScdkrxweHwuekA
TPKh8TnXbR5XBulqYuPis/7F8blCEhAkDOPaa7IO/H13olhmqLPhKfDKoPXWI2qL
jXstsUvJhFx6ukJEl/u+sT8JB3vDn6yLPMGEah6xKy/j9Skir960+tsI1jlYE9XN
4fvlAiZ1xpk04WP2VVEDlILmZC0b1FSquuw33tcSdBF7V8BvaVF8Ct3eFIobvj9n
hROLVC+MEpVi7VL+hhUuF6P8OPzVXkDha/KqJMLqKv3DePWcao0BsjFgWpaUp414
7TOeMq1TNryQx7Q0z8qtDMxzccGbETTal4Pt4YqAwLmbqjiVPPTiACoaVFyzyY2s
GRi8TRds8STE1IsPb1SJvSr0Aqlr9yPb68z5Or4yRhuJ8MGv1Co2uswD0G1oHTZ0
529snoiJcyc6Si5lkh5tFIk1SBxif3fob0nIrqyJW6gDnAbAPYkSiP+FX7VjJ2pz
goI5FK8Sq3WB6rdupT9fmYNNSSm+AxzgZLiJM0nNpnfTX7DT3YebGeK4lnvyCIlp
qJEJsvaNVaLT/ohE919ObckeOE2trsuv+YyDdqDn0mEpqlR3PtCElKuBgogGfIK+
QMwa90iPkezuRpuc7ZSq6RIYwg9Uc1CAi8viqW94tPHBwl9TsYXjbqk37gLjIhMN
dZEG//rXX8426Szt8NrzWfuw6/48QVbA/ZuShVdPM394xDS4JtsFoWpqlh3xrDiQ
9OgfFpeRUqmDUs0th0W7smUC6RtBdntY7zi52GqrLmiZHoGMffWjcr9/0hNHGLjK
QLdFXJtGFv6/ClC4oD6qgGLVtqn/HaHyxlUqziqNKMYUh/5l1ppTlt2QrzCEb3my
y7DAS1pEdeuYKLWvdkd0ouo3G0sSNodbvftePHNu126SJfnDykhE+IRI1N8O8DL4
iC1XaHy2i6bsqzJqpJxRl1KwHgyYLRxBTrBFshq99a5H6Ij/zdTv0op4yEmAHFLm
GWZckGVddgz09QabjkqOGxnklevRZAENQBpEQUYsCJxmywVEipo7bAgcZf2u+NYD
T1pRllXf5YZiEW40Vj0l2qu6jIQga6LTYA1ahRwZQ0LvQOgAjpvnaDhjALaWYEci
FA5k+R+NuVqwZWEZdQS2FbhfrTHElHr0lK8lYlfpkMyQ2H7pqIgAuyKKjri1nFRF
Q8asE8mMEhT2Tjxt6WpjP6IYgX9GYI84CT5tYiztZszJ+vCsz0tAmzW6UehOAWfT
waOYhc5XtlXcby026F69S2QZWPJaE3hhdI4HGOAv0kUvPEKThSOwT8dxCZpVZn91
8ZPHdlI0baUA1Y75zpciw4trk/CiVSDT5Gfp3eFTodaJGe6kR8NLf5E9SJKgXzub
BL//+DMVeo/J5q4Y3gVLvf7DbUhAHzzuteuUORvoBntAnu29v4fjFo2fDAst8VBX
Lh2sjtXovzfntVSio3wh9Ha4ccNfxf44dxX93KFpDDyDtlen9tAOsPkQ0mEc4vf3
z83e9WuxGBh3AkzYNhXdrsheGMjKaOoUAnTUjcZM+1Beuhzn8R03oeeP/tS+e+xP
yITUV9lsTVb4ZtTcI+tNN2ygAlCEgvaYavGhIFgbo7rYT6ngLHCtnW9fBecGFAd1
chMeWuVZMm+zfnHfbiqDAWuhMSo+41GzwZ4jxAFQF8I+iDMJkAhz4CGFV0OIsDSy
vHkUqIEqFO0yb7il1ZO6/bofaVUatdBm+kTNoQeGFi8ZQZCetR/8r+6pz3B0xE1g
jdZOav+Wkg3Ceh8RfXqdiewQXSTybA+U1D2toidbkLrpuVADc82Nrr/g/IqCd2ji
Rc+pnR7a0pCzfBUP1S6+5uixBn0BZpnilln9icm3WmuPQfrDeVavwNMtHXd0brn6
p0N09wtsHDL1/Al1Cg9gYRniuO7zwdPS1sFd7mC38BdUOL1MpQ7Dz9c/2NXnKHB/
1FDwNtrDqoRnASi5tSo8IAY7t9ZhZhp7dsBQCfrA+y8cCGGkMQjgbOLPsQU+93x8
fjpS/+pCJWGqNFaQGHxLDX0nS6hjAIXHKeMRoesH7lYqjDZT/2Z+0CF3npzTsiLE
413SK8+7uxOiYg1C08XgfTUttMLT4oMhMswxsxmmctMjjBbnm6d9mP+O78W07gDR
01jAtbspqYvsDH9BkHMNRwoS29RvrYF4+M03zwOtasPtuoIAsD9npdnvefXA3NRO
fuJSn0EXtWIt1ePvpJfYTWTPsf6DmnA3/B/L3et1ov9rb+AvTXuHpKKG9+B3vRS1
8UH0TBQgcjFFxO5nkEureNCDp3MEorFiGF42LCEZ+XMEzXdDfZ7uDS4T3EvaIEGp
FeWgvyJLTVD8IawX97Y/gGXxAVzCiFIX55AZV3XZrO54fCyqhPtIFDqxZAHsG6r/
fETD/Nzpj9Fb8nd53aOig3kwZ2Vvyk8pOH26RnfFT6hCz8x9DD5WdDGjZNnRmXZi
+kepkQIlwzmZJXn6ZMCkutdD3UkwOBZr4i7T8/lSG4QHrydI/ghqGOR8KNiLO+kj
PAog3oL9F77C+WGglFgZNFPz1VTDYD1oFkHp+XbSFbIT2um1CKeMnTRIWSw1gczL
F0u5F/leKGLFyd+Yv0hI9m+GCQD6DO1Uy3g6x/IrDYyJc9JpN9lK2SMgHHsM4Vp/
RsENVa3Ul5fw32Rkg8F++waFr0a+RF2ZCAzeLSN78hzO7hRlyJjXyXyIMz2zYz3c
8k41aKhq2E8W6V2XbWP/VkjlWo1tqn3KlGdlM7oZ1BgSHoDY30MpJnh7e9bG4g+L
oO9NsbNM9zmFkBAib3weVO1rds9NgI+rFp8XUuRvJhIeYWR4Q3aAZsNy2PkvCk6l
vL3wD32L/V30+FTmamr+nru3Sjir+9/lH4ejF+c2NpIXGDtXq/eqy0VMpqTEWHP6
9HyE01jWjOZAo2LitFH3BEwr23StOjd5qbi+30m9haxdvEbhjlXUfB9GnDzBAAY4
+wOkqlBwju+3Dgw6Ru10X4EHjduoiZgFQTnxyEwvcJ1vgNeEN4r6IuQ1diukq5ol
y5F5QslNXUnySJO7P9+kbB+p/vmrhmk5KdFmJgMF6cuPYEb5wFbgGYPK8GVZX15j
LY7zDr7ttUdn8TScxKrN68TPHSwvGEZz/DQ4Ak8/24fwVjQXzSa2VnhipQHRgNQQ
7kD7UhVevOU+WFUxWPNqjNp+x/aQzLyvOqWjj0P2QtDi4mepoIRx46PoI4OZznBz
k52YKSw87HycmZklsH0rWoT8HUhHbXaSJIZgMFhXNByQLZeb9OQq6In+QqT+O1yX
wOOGNN041nCfknLEq2vT+QEEzc4C8C5Z1jmP3BZHnK4qLqt2cgx84yPsdpqPYRrK
iBTvsSuhSfeNefCCiLNBld2RNfMMn7VZLqtvln+PgC56Oy3sSFUv1T2aESiLGV0h
HPhHzuNejysqK5EyTbKKeSyHssT5j1qtZQRmx1af0gKzkv4AbOh6L3R9f8XsiLtM
U6X9QbyxODE4aMhDtslDVRGDel3jUb0AvW9Sh6loHiW5DLYKXQXlqJ9OFMVq6p7a
D63/C58Q9asJbmnrDGFcSSnJdqVJ7hIO5iAlMWZf+jddjaP3Y0XOBKiPoGqqzCac
RxKKrgDlIr9N2EifL9hmGvrFDN94B2yoUsUGHzDju5fO8eKZAUql8J4zfAFE6JPz
YP1uWn/+tX+y/7eF8GLJi01mzkmPB0+JGTlr0KhASNBuLIxV5bkL81bjVWyrsJW0
OpZiTLhAd9GYIlplqgNcsghU0ZbYSEJ7EHhM47I4evsqWmAACQnq5o5DfLtbjxD/
eZ8GsLaO4B7xOdEs0xdGpHqEYBvrbRJTsVzoykUFWM9mAlj+rYGUPAP85ojKz+os
zxk5vMpvEAI35ENI1z9EzRgZtMG9iEOlI/fpm+LLGoazoJ2QcgewP+KpVtPL25ZW
4dBWN26CfZAMJJ0u/SxS8DM32BKDNnj2IqezieOak8CCP5byTfvicI8oQ/HbmyBR
k5wInMNDKtMLHMfOpA0D+l4gvet4Oq416aT89w4IUHBIc9RMqK/lu679GHCP+USh
ND4Up+6Fxq0OOAB/5iU6akRUOccr4w69F2oBOXEfmNLdAacGlt5fG/h2KzBO1WLE
W66vNmcRTKuWkWA5qN2iw1zIWMRPY6dI24VLTN/Onp22X0qAvywWVO7+SMc54kEh
UBNZPlkxyOMRE+6nFnuUbEVZFDun1qROPEcK11bjVQsA7QtZq54i/OalFC/80Q/r
zJzEQo+NBOyERjZl1bmC1t1Pn9C4/ZluHovnafOrM/SpzvdyiVwQFyW2EK+4F114
plB4N2sC+NSENhf6GwU9GRkl5eEnDDZeE+aHKced+dWzXvFi1TPJ/lWzBJYSaUmn
eQ1XNSWEHHbkBORHPUgAdGym4v9i3JHjftB0CuTYLoO7y3yBaZAodKbsT6zt8bb4
UwTUtL2D3aBySsUD+9euEAP0ja4xBnyXz9kG3xTL/1/tn39fOJibLDh6ABJrHCUz
rJcdZMep52/mf9aMchsTuuc4d3h4tumOLFfAlUBrJOgO0pat/XriHUdnQ9uHVrYb
39NTOJoP3bVpIMI6AUxfC++4IYMy8ir1uYCvCEqdbACuMGsLfBz3RD52uiUqbL8o
GlhXPwYO3/p/ke1V2zbxsjAW2p2NRn6Eb5fRhrDMu002DNu8Rhu5QHWsJajsLYzl
9GUX6qRdX4BDmVDRoVAfY32hIdjEaSSDhUMK/fRFfeZa4tJicfDNR4NLopJ2NwXP
Tl8/JOFEmofgK8Wu7PD7HzdB3umCedN3WEFPLjGlzxQJZrSMJ5Zm6a8lnuXFsWiM
1roWhnAhr8kDln18ptzq9Ki8oyXkv7uBGiYwNMcFGejAi/1cYsDth5Dj9ma8BCdq
9GRvND6Cz5jPjIYFO5+uXKdFYHsgwhPBayDelf/tFXU1O27zDS+cTTYSjbef/gHs
7BnCo2WEooUe11ecKUAoVIB5y5qbA0xuWdmpCBiIiRQxDvCqZWlMecC2VPy6oN9x
NRQ+jDDFPj0Ab7VBlWbBU5+VEJg8MfuzDHbcjfSmrvfIRaPjHqEUIorrzEeRB3Ol
tKJyPQ1Hgwft1ky12CchY9oOWyF3fr3PYhaqjyV/4v0KKC9fYmiEVRRtwBIsdbDb
WWupgBAujrf1Uv86Hb1/Ei0JwO3LlC3RFhrc4RA6b9Zi4Cp9F1KtOXQkoUo/SJcp
0yOmrwDsmdF8vS///8dtB7RRLuryIDSKV0lrBCq49V3lVLrb/zfU5YkY3nX+u+KR
0gV4PX3MFYkK6Rog8K2JqjksIctSsTT41XTAHnJBmFxP4Y1nyh91zZFUsiHEi1h+
RvNLgUF3W8Kcd4zTXKgm7q7I89JhS6qFhZB7ZPBj2Xe7MIxJvOV7WH78qoW/WAXM
y8qNPI6zDMpYCmpOLZHA4tmoMMDzVPlQPptwdmPFiAjXN3NEizXEOkK2qbPWq8ZQ
HYZP/qu5SRUcvGILHCoaPdtur4kKILA3lHXz0IB1SlT/LYf6C/F2RlCYDG/63k5o
zr1hYez9dCh0WA94pY0bjxMl4l5YaskP9zRNB0bw785EOiKk9JZSQTIEREskWoRh
VjuiUYcwXHMGc2h+C++l7SDkf4zId4T7MLcgDnWx8vCzVkCgjjOp+i1vv6Ujx2bu
ha1rh+tDEkHVuIBcEiw/YRc22ImrUmioN7afXcFMlDtWf0u2RioJtiK77ve1S8a3
D/lWSOYQQWXbtFUnCOXdwuGN+01rkMI6zXnkhdrRjGs7F5S3JZnDUGc35c48TfKj
yshAUpNdUi6FVFoAYfNnZ2ds/uui9PErHGxTrwSusW5euVa/IDixxq4Q4PFrL7Rm
4x9V8kqdAO+UsirHADNXDgBzS721gy+gfuqp669mlhXEOBXidJuqmS9VKxkIfPYt
smFLgBpo/LaJvkOs53EqKf0VH1J2Yx1edTwPHjuNkjwnnkqOGOSMuoCExTXhGJZL
cFs7jyb3gwuvzR8uefLr2Dn06r+vsFGGw2o+xu2u5FC5rhGwE6aT4yOPYwoz9VPi
Aqdjk0vhZoFHKc2Ge4SWMSJFCuXKhI6yjagtlFjfcsLcEEfDtmHYckwrOK1ett87
TNHOBAhXj4qEAINSrJTiKI9HglwxJrCJjXQxLROuN6XjnQuSPN0up13SrUxB0MmB
jGURPOi04Prs2safO1fQWTGOWy/7bVqWEiTB1mqVUuTNX+uM/W1xSgejW8xbZyYl
y3KPZ6YWT+z3r+AfsKfPZAjwA2JJ+Q4wBarkGEmScX89sO28QQzHQ0OlHqik/Mlv
sv+n99I5jVrRJiKva6c5FwkNWQY6WLwiVRMH5upKC4oeG33UvaXScyVXVNkJmiMy
0h7Whmm92QYIyROXcysmmNratA0G+yFjeBeAQMYiS5pg+kwQ7S6xyqXj+ak9omgp
hakbblSjiwwyKHgQ//FjL7mTekA+lqUVUhEneCYUJ1sr8y5LzkN/qDibvYUj2JrC
Ut0AD4vgq3jYBm3G870xd9a8xGD738PLnDY4FgkM38C/nx3Zbc8B/GjQ8hqZtweu
0vHNKVBYQpGnkl0Hf8FpcWrUFLzBpI6YKCBdovxPe8iT3y6c4635blZO8z7Fl6YO
tTq+RQxv5bpNWcmTWitDKazYC+YiwDjq8y4p+LRl7RrHte+gvBUuOj92lvWSjtkH
ddTw0rw8J1YJ/WF/vKZVWJce2w1xdNl4D5l7OnB8b4E5VE+WSaVf3SOhHOd7Mjnz
aZyhKm06Co7VTnaYgBhBsKTEfubedPVO9HSu/Mspntob+aoJLPPSve0STmAu2RSx
iP9oW+G+BLgrKYgZ8n5zDPp82kt5nO5p3tkV1pBFOHjeosk2E79pzFNMy9RoGj8k
l+cu6/Fj7y9QW6CZC/xsKkUP604Fmg7knGkDnUleFWcB23fOeSTLkEvto41DLMqK
NZVE96Dqpnr6tT8uA8Gak8UPae2G/y67S9AoxaON7VMsn7oSWx6C7dZz3mMAaYmd
FLZnAHRtd/j1W+tnT8m/GMtVs4hNX0M+gUEZ/Yf+XfTXjinCfSNbvlfuMUtdyX4l
UfcZtC+qqUYjq+zRaxszoGREb/YxIHbSY+rexXBidFvqgkB4PLOI0bVPQd3aIcEI
rz/mfTw17640ahtjCo59BZ3EsllzB97buESLjeTfU1nNypbIvM5IBOHvCaIQVkXB
LuM/05D7W8wqfZlc5aCQ795DRCEGig6z9NPTDVu3BQNgTN1pL+SR5zMSs2KhrK2w
VtJIuNKU6Z44jAYc9s7Xvwr6966i4TByOgZt+7n0JZlI4EkyPyPPvFHnC2gNs9p4
BwwinNKdONN2w+AiCu5xQVjDMfPcdA/6rzxuH+KCN8HP2JlUU3ZXpbtWRmuAxo4P
83pfDBXjc2UqKHly3YDmS87u5wYEfUN2oqF5uV01fhGIDIle7tPf5GSb7nxonCmO
tGpohjfnllfamIdZXXhjMcwckclrID0Cm3HDnKbtwRBSs1/XLv9fhkmElFi35dDK
aiLBFBef5v7G6iAuD87Brq+BqaZOLpJN2J1+p3Qxds+cpZXEwrZV8nhqmMOePixc
xB5XkaDN9L+VZbQqh1dKJnEnc+z47CVWRQxY55FbSPr5ZT70qjL0EhanqQqvWeb1
yG/0YgLuvDqrECZ1OE0FBKzPJBf/IDxHEJ2BKDpu8Kl9J6Cn53CsKPv0aWKmCn0S
3kkQIWxyhuwUHgXSyY+708LS0/EqGN5YZEEtzqI3t9SVnGoH3u076EvZ85Q6VQV2
z5hePOkYlyGpUFhPwXMzLKgDsaLMYWunPF1HQmWlWO0HgbBF2YU4zQCLIhgP3fIN
nU7MQSeqCGBK+0eYV+tCnR+ccmlpTMAbnfivj3CVKDNecxSGyvGHEiHp+LVvnbw3
ugh2SlMuXYKHRXIGq6tThs7d1S09285hPqfyftBK0mpbEVVJMqsRq+dpaA4JTnJV
GQ+/CIHG8HsVnCxXrUoPKyRSRtJzsMXNEafU2EITM6sL7AaJdGf3fIlwM4/Ul7gF
fZS7y2nw2hI6N0qKJqqHlUa8eQ2C/PepmB08z39N2HRtMLEqcHh03cvbgnXUVpTR
1CfJKKUqK7rLHRR7eMx4QCJopFFxI8e70Jd6dHPJo6+YZ2mN7VqTmuASAA6H2FXA
uOwGkesvSdjEKUDPTlwMFRfayaKbwr2d3Dxjc5rDgqz/swuqDD9kLpuNqCpD/HZJ
E6juIv/AtUPxEPXzmPGmiVEaNTs6hMaSHFULeO7OSiJxWXjm4C9NPoxkluw+1RE+
nGL/33LXoFqxkjLOgoun/zAHWBbixJgeG2QyqWRv22a9r2tswVat8jLIkVLZxG2E
kmNBPzoP0IkZK03lZr6GICYOah6ZfiSeXPmiEoON8ArA20bGh2neo5gcaZar1rBX
Isyr2DfZijwqV78hIEG/rPIN0NyRq8WVPlUAR2QgKcP7J+irjeoQojINOQPU6y6g
o4Wegvq8f5TWM1rTh2f0bSyi6nppVAa59WzXZmqG6pKBIX7ES2Kn0fKpA+gOgYvn
yGUrtbca9hmTltFk5mr7NblF0ClLDPDvYlnBtWJmyHi5taAEIm7dstUeFDmP4CL5
TQhHRzN9sjBITZdSaexU87ZCdGJSBAmMkocTjbmhJBi6HTeZWApcaEpZZHQvn1xl
QGXtmCNWu5+mIB3nJZmXXARpN/GkTQ4p2BbNlol7Xr7cvx6HUfRy4VpbTukhZui/
yKQmebxhS3Z+S6MEapcpduMB55egqdM9Du70Mfz5ks2wMiVczxbcJ8584CUtrvm9
rslhn4LFs1V6wEPI/0XsTGkEl5hsL91R1/Q+ibIC6nRH7OkA9I4phbtIi+8MvMir
0knVeRdFUfXyIdCWqR96uRLpveumfpNrh3YVPsnvlth7Uby6F4iNiN324v95HxDR
hqDPnwNp9NXUkuIiwNoDaqN5ARuf4U0+D7JSbRzFZb9dcKa7sMcwfcTIZMs01Anw
U/V9QTUTJOam+Nna/AbLUHNnbFkN8Uw3ypxQGA1bA7/+TNEA+y6YBfN50D5BSD+X
01w0rrDNga+m+qYPyQsa95gR0CpIfkz4SqQwBkBWT+vrCbhBwIJtx7PyzfxtnJsc
WiozG7r67v6THDkm4OZk/0dW+OxO4hxtaMvwcJBLiGgJc21xj2scTsXjUE+lHzdJ
XWvnRxV2yrGdSvTf+4yyfXKe/0vP+LAJinM6oh32hVMTyNU+Xiiwu3XSslXCDk8m
YH60ot+oY1l7+wRGL2Kvi5bMW7wXCBtNrT555KKSa0uNSQ8aDtgstIA7wtjDbKoJ
WBhuedqemzGt227imkySYeJX0BiE4WazSAFFki04lCKTi7KG/A6DMpB4ZAKHITZf
S1fXlogM/5poB2/JDeCYK3+Ch/S/JXJ69rlYiiqOJqYn4VgMclDm7kE3t9boX3Ei
EWQdJjZQUx68HZVWZRiBz09YhFOmMQNgIQ0+YAyuxFQy6452BjGRKzgP3U3C669J
10mUjpWc22GevSHboY4LQ90DGqj2H7RT9dmRlenzSuN7/luL+yjhXnzYGTVr9REm
DjWH1JwzrgrBdmX1TbiMkGAX4ukaPBDq3o2+GH3DwQLENv0L5YocODF8ooS5Nvdp
JywxxOmrgrenfcGX6I3rCfuqvPgwlDf+30bTRgsHBwm8tLQzxToCmEkel/C78JdE
sOfMn0rLtuo6/gtycmLdGxMtQ64e70BQZI6GS9M4LuUI7AYk6hIiUviK/jWArASo
krD5AqYOSsOwtP2U+t0GMAak8FCSgRXPLTJeBru1mP9/9MVsDqnyWvDAGMHmLG0R
YT/vKtAKnYFvEGTRzY3bfTDJblJAo3m5kO+OVRM8XHJKZoL130oAb+V6iQ4DkWqL
7cxrLsbbTES9Ubhckv6s1E6BOeOtrNT042w+MfuYq9Up++bDYPAqELYO4wk9wYrW
ZtufEZmbsUJPiKa2XwvzejqCCj1QtEJKAOhAVMtUXwRZXLSbzy1VG0BBdB55LWiI
+BaGbyHPaQM5sk096cR++hyMEwqotyP74SOEvk0sbIxrnghk0hv+tPrN8Wl2Yaad
HFZm8jXMVjEWhl3mYU61PjVVPkbsPIIfkTasvxbk1+6OGl86ApN+tclDqPAD8NgS
oOUOLGC7numHpKoJXQ4zvuDjWdCZyFNVgsyMMoxUvjECF7BhDBN+j+fH+MdZ+E3S
53XYnUD4FN75yDT1cv5UBlyYvVk2NwUMWyoVeytGH354l/JzBQX7WbnDWyXhRuZ+
t6GYtqVD8zBJ/Iqcg9oA1PDL18+OysE1DXWfENGoUaAXxJFRwPB3xdg6GJxzJJhY
Wtpix9WkdX44F3TCJWUwGfdDKrcvTReipxrJrUxoa9KQmBMybxa/fE9orDtS6SDX
ZDuYwFh2e/yHP2z8RU299ghFW41NUJ70PrtYqPXEOcI+8dE6l9RAuTZ6PxewBI1H
Go6AeBkZOJHFAjdP1qI+7S1BbzZrn6SIUdDUrsL9q7yBH0K55i17TaQGccOBwOtm
6auQhrhJnbmGhP/2we8KCaz2rWFwh5ZbkxVmyYUeHtZkUY1zbJH9n/2rLZGBIuZw
dOLBDX3+cSLlyrg4pcUgbSp2TnTjZP6qK2Wxr0rCS+rjTRpLTEZIxqsYOG/P/PBk
CbGatqprjZpk9fJB0tduQlUcDgdWcJgHKMiDykyKSNFNjZ6BRPw4GKMIy/ZygJx9
MQxaJp1wf09jM3uod9oVVv36UIWAVETSSC4YZuihDvLoBKheVUJrkJ8HK66LXGF2
UkJ4zKamRqfJ3+CpSo8y7Xb+g6SqvgPc4CIzrENNevDMem66vWHBaBH2KyWneddr
RGz4D0CWZ64dMV+zGsqTRFMlMnML2CDgMhyQ8sLNetqlmdZwVhC4uoXirnUJcjCF
Q3h6wneNdsSH14D5+xpvgiuUPdP0Qa6pVWJK4a4btY24zuGQl6bmEYzZtuxAiShm
wOYLXvOo7tylJHXdzm5rscxFH/o0IeqJ5rd1fKzZhtpfgOGS+h2pbbZTB3z8oQCL
vtlwj5tgM0Sh5+VWiWHPPsohVWoTr6vDv5QdnRXHMEDP3FNwmyQfpn8vBW5D2a+d
SUF5XW9Uw9SmP9wC+ZhoDaKzFVWQH4miZhhODIl21YpFfeZdR9mw8IWDdnTrs4nq
b08TqGgqbf41o5QuOTfm5Q/aphd+Po83FHDTEMtOgeRM7OGXXFoNjQVdaAPBVqVA
v/0I5Opyol/4DcBgAWXxS0WLvpcDDVdz/DeFVLvwBkwXdjRv1dlojENMM0Yxlngt
xXQdVfkEZnm5XEFRz3j7grnjlBfCwa+7UPZkP6ovAxWXQjczDfZ6Z/Ouh3e665b3
Tx14bhyZvPH8Ppr7Fd5bLIhLa8aQHn047Wue7yYlKANyiPr89qWuQ0YrMSoH5jia
k1/UX5sD8e0sWT2/CcD0KyXn/5xJ+YWXIguKAlbnh2bfKAoVXrKljSqnSxFv7HA5
11RdLBO/fVvhI8Fg3fiRGMmgIKoAIS6KLG8H4k357rlndVGHIDzbxKPEigW2s1jw
vAsk2Qv2bwA2OoDuNyTi+cl4hyPATE4jd6txcho1DmO3cgRrDpUr/sx8nEF1P5Vs
rmO3qMCRhH4oHIJoTpEaghIkz2KKDh5/+pKkTSA4qPkwORLnfAPaGiB/ySCFH8BA
8DHpTl+AkqPTc0dXSaMru1FIWhRIAq1Wu4u9YIjfMBOKTDqGMVojGJaFG6PZx4xL
Hn8Fwmv9p8qGaOjFTZl2EBjlC/XB2YlCFfv2auCxYV2e/t4nTMsN+GN0OCgPhwUp
v/EifTKSabWx2BdCHWPil5Rxv6tQVTZJyKusz+yTq99S+1dKf8I37SDFthtiESCs
YDWeekhnQg4byujw9bsmBpxbR5D1lJq0fC4399mM1ax1eROEDAGmk4DTUUBZyeBE
e51O14yEh923ojL+aEbDY9to/Nqxamnd+JssEA+dG7paAhUKPlNkeNhYWSoCHgrk
zuNl3QSpgQKvL/q8TwjMcQ4u5z2tlr+wgGsGrLmoL3dIRFpq0iv+6rlyTtyMRcVL
zXceKwz1rcMJBl9wWHdXogBh0EVZjmmq6T3Ax62BFDS6kuFCcUfjesrH5SOjzHi6
HXxhD8a0Dk/bmmOL98Sl7xRK/z/MxAqdXpHLdr0xtkGzJjFOr6CV5cmP0M97lQ/G
kaNINI201UEx3kRfhzyzUzNePgfA5RGYd11xzwY0UFUcyXn6cwUBYPifq/l9Jotz
lGiaddW6aw1Ne6cd1LrTqxeC6HEF0a+qlkJPTon5RUI2XuXMq7zb24ZmkSeZJiPb
fElWDSurybMA0QktK4/ii/JMzMELYxrgir050WdRuYZLV/RPpWD74aBd+K0D8IdP
5Kh3N3WS4xkqeZvGOK1mADn2XOkNXs1BGR/s9SpjWSbmREFsuy07GyNLxvyIebtC
nZz3ke3VYz9tMlp+W/EZOeqeGgMbTBjXF4fDWs9WVbiaZ7vCoJiETTbXL31ScRev
SWUGUQvQNRQLZ2rt9j0tAwAOCeiG2ZXHNB3LgZy+9l+9ff5SeERvXOwYuzI3Zjx3
9HA76/eXa1pxldGPan2wrgie05ulP7PeKkchNXgHdyX2pRUs4VHMnm8nghtOuEP/
qdCub/HrVkAFg1QLemqc8FhfvGqwqVxalT97MAAAj4PzvaGLQPpvV08xIjf7zRYB
hg8qv0R9VdwUpbtcZn/4j3vAKk48LPx4Rl+rXPWh2JvYmoWEYYhGIXR5pHgev9n9
OdPpVzPj4StDvUceb9DvAEP8udzMduytz6GdrOy1dGWjnSAgL6Wm6slRZol5j8m3
uBMrMcM7hBbYZ0eG9InyxyMAS0HTrjK1mA6eDjE1hx8txwPN/gjIHD57xVBcoQwI
9tfYqR4Y8YyrMERck6/PPXTP8RRVEpo3q47eRqv35IzRYlidx8eLzZydKLotvfNK
92YoaxBws8Wk0IleTinF10AlFICQ/C59/CtG/8hv8fGxd0eWdhhwiLSstzFe/syO
jetQvtcExFdxi+Gos1/LdYRAFn+Bx5g8ERHVAi0WlkzG/S6jrLnxGFDf2qNTEVAQ
aTqJh/VAnLiBcOE+krtQr+p7T8IPQm3cNe3shuel8DrqhFnNHwKiqNkL9w+j3aHt
G6EmFduD38W8qe/iU5NLcRB2qNplq6FSGxZrffaCvjzho2CGEVfnaSnsatk/D++j
FJ6m4Mv1w2l5HKSMmAdrQafsH1tZaQjfiXymW9DeAV9xJLST4Wo6ya1aUCxEgGaM
nXST7NMndZF5s172b6z2VT62rLQ0k7tiW1XtHT4MNkIcBtakyB0u3nhM2PqpTsVF
wbrkxbl2GSWTlxB1lYcVXS98jNZlGhEk3OiMVrQyW9wM02vdY8zfhbyk4RwcwvDD
QwTkGaXXad5bFZStGhPsTuyjXCmr7P0USuGDj9OYCjAUaq72bwbvtaDSTriRmZMH
U8Y4sFRVpQKdKY2YOyfqIiAeS+lHiOCmmoP4FALKpcWqvhrn+i7hdSYOXjHM09mZ
BjpjVenaiF4jZOXrVUAsRQAN7tidNOytiGz+P8547GI68wsiIHr9kw6tahdW90Tz
q/w2aVwOog74XiMlO/IMA/hn6qdrsSi+sPv2OrW+5Y9Ybl9+76k/uad8iuCI3Br7
y8euzOqhepPW4Y6YSwVa6WFO3IbRLrraKs1mKsar1l1uiI7O/2lV9OvJHHh900CK
ro+KlTjkr6RfnsjsmjR/cMySlSsVX36hfLjFbdgz7CNTG7/ou1ov0xaQ4m2MsxBJ
Fk30f5Ne486Wdq3Jgj2B8ZVuUpEAPw1hbKMu1Vc3EJKC+LUiNZvB+niFCpaxiO6j
RXVmxiFx5qSu5wx+IskvWRdotchecf4QknDbyhuTND1usbnyGolFjAJQX8Z6pjY1
otbqnm/rFFWjKHq8eHPwoDBjP+/moWUcFc90I0AZuMMyAQoo8V9a1g8unoaWWzqt
iMWhyRbWKmd/ofrYmMYDCdml3VWs9GJrHrx1/mtYJWJzVjfTK137/MQJPBwQsm0S
8qPX4ZC8ZBgxxrYntoLudjqSviAxmZJcAoLdY/zS75YdVn65YZfXHTY+p1v2Kpcq
moRvDtjoi0FtpPDm2YvAF/2J2TddSButx/haT9fHyAgSoRh8VzLZX2Hor88WoIha
rs/NXY7gPJvVtX3MQB0CYse6NpTTlJ5ed9g08v4s4Ic76TIUUuqd8fl2NY1zm4hT
CFGxM2OewpSed0nvJWM/KmACsJUR4pOB02vub0Kq54OHIyJXA9TjSKa0+b5viyNG
Wd+ajDz97fgdD55WXbb1LR5uS+YpJ6es/5pf9MK/Lp4yqSg7LwJ3INOLQrBvXpXi
iyGPC3S11ivw22pQoajua3M2l7ErOD2NeXexALeX+pHfG/FAHwSV4YZ9qrp8H6wT
Ycv6BTIEAh914V66O6EOHAUkZt/EyBvCrxCx67WBvLJIaewzMMiEMZdYQyyi0mte
/fCGRgjvsjQbkXuQ6tbemsIP6N2l9mUS7z76WaBNweqS+/RknfrFn1ri/rBTxssc
p4QjIqQ0sS4EFINaEnFKlTINgLQHeFFNwOBLWCbXUtmyalgDrrlRmO1uDY0QjSFx
Zs+mUUWdUWoMo9DaFTZ8GCC5as8ji2lF4HNR6HrkP6BS5/e4Qk7cQWQ6frmExq6c
Udk/w99d5qXsR+R1ZWCjTpcn8LTV/z4avg0A7aJXchtldWYeOOFRBIyXdoRwPRk7
GNjikcUwKV/xsaEP0j6DH2a/wStFAMzo2SvkdbkaSWAf7QAYE7ahBZseSTEhu6Ip
OF1v0DBp1mdw1h8cFpn0KD//iRAuCUlLMCHkd8QrfbyNCp5aqGQrH12Dvyu3eGy7
Cmlg32W2w50GGKDwaot2FGqTAxGbIFSlHYIcJ7ec7HVcBIhroBWi/NJ/O6y8/anJ
nE1eNfDs+rnoJ0M3CGfvgNxwZxDXi8K/mLDBpLeau1xzMEeenoYKzuesUbgCJMXB
anP6VBQEoLFsOrODX2QL+EOrU545vTaujgK6OJlIHmPMlQjo5IpSIH4x7Wxhrc2P
mzk2KPPFD9ssdXur26TaVEojbAMDylmeQtCggTHGS3RwZMweNiiDblFOEDwbxo0Q
+VEyVgnD11CgeQdcXuLkXMuiGqfI7sJhbNxeYXgbKjGW4whjEtJ0ioFdF9XbbtGH
GmbZxALi0G3u/Qv15qIbeGwNufJnQrWLVk0fiXk4sJPBzxBppSHTjStqQJ5qKNLN
uxT7MrmJyevZ1VmDbWQFKLiqYp0MX0zaCs2L9yjnFxuIArvdHqD0wtRy5kfjnkoE
CopdOV6z+am8WT+zAzWebwHKBbzIGcfdzJAAzRqJJle4FFVpphfiSxO6Lx59U+ZB
sViepgG8ctan7TeB7A4QAnXO0IYwnCRuiUNswzxgggGaOe4lQJHdarof6yia9j5K
rbFOQnGBuuZgAaU2HvQC9zvZHTJGjCL3VvZ/ssU16oEspFnTVlPQ0DOSabs8QHMV
K8Dt6o0ThnpQH4GCk7WHAzSqt0AACns4NMpOfq4EX6WZHC2JrntoI1DIIdHJegt0
0IgIuAQ7biN9eUneuGhchDNt0b9wazIhKDTPt/RfC1uL4KiT428FUS2a+bZQq1qe
Hk3rTH1AOSkmdFhdwqO8169rJ9kMoQZ+Ld9c6WxrPoMoPUPS8jgXV3B080vJUnNv
p4xXEtXOpyR3GHDSP/CwNsyq4xy6quIjQFtkHWbhTrU5FguJkkeiHAkT8klnWrWk
SkxvtEpPJL5khQidTg4sdAZcLyfxPpq08cyieaUmodZ7cWWRV+DcTF0OK+Kt5xvw
har8lGrgnP8DTgsayKYRHdSgP+OG2+HGEIK4yr5Lj3t8JZH2J9qp+OrIM0DdGrlS
cwDEa1jw4RgzrX6WXvsdvnMCHvu6CwM0OenXLsAc77/JgQmRLtbuF208+q5TMO6i
BmpzknUs0uk0dc+VpHGxFIcUc5RCIsEWsDDO0fsJSufuU1V6zDPwvoVPDTqfT/R6
abjpd6n4cyjDlzrb3jiM9XgPiikRST2ezvEebakSINTmsXnhMVGWe3GmolUZmHZ3
RvenwCWjIjegd6w0ArhN8qqrrnddrKcMECumVBZpIzm4psFVGBSdFdWc9ymv8fMl
0ExVexIs2RLUtnsI7ugmkyq8W2LOKvDwQ4bbZgcZhIzqzdoVhgYZOkMJCMf8jpPP
QcfO89LZU9UfASVwpgTOPcsDmzyKFLR4nA2696V++FD7/VBF8oRfjsXtF/5J/ts5
+bcciX+ENBnfE+PH/5vlB4AMMv+/uCwdYEPNxePg11qx9E/Ey3mKmjzR8DVhUH6v
k2aG29v2TOO3SmkFz/6fRGNot2+hTg0TNA/Tc7RwnKBEuGsJKUr/Q9IAUGigAO0Q
gnBDjd5Yb0CUCOq6Z+xd44RncFwvw3aeJU7zKGGjokOt63Gz824ZqbW9u8P5SMFU
5r/G39gdTLzvYYuucq6FWdrxdkcoGoEb6XnNgBxy9fE4l/Of91PET9rK/mVZaNTy
8hkenjMlCrn8IJu6Ao4MU03K3svJrd0WMeV5DVcknx+ZMKmEko8F0DDKxUO0p2bX
ZjmEQ4TloAjIetiVBPiQqTNPDhfiOujn9OnXsUb9pwk34ta2sw0yDwVsh9q/W8Xo
igwdr6aa15r2j/KsSmTISAxT2CfwbE49LimCWF6+WAW1zchZ7JQ1ooTj0RG8v8mS
ndp148baY4Ylri6FqofrZvlVtsiq5O3m0zB2V787spONI1AD9iAY1cGecR8xmH1E
CvpH43T4N592/EQm3TCD1PRiWb17WwUh0a60bKcQlFK1GIOPsK7UNMW5mHA/8kOb
Ut/cmWZ/u3vIxkB2cFVfENqiBMUj6w4hAZCIzgImacTXE3qudAd0/XbjH6NCK9RE
RHebG+iQ+SQfWX0BkhwdR5/2Duo451ZKPTVvsu8Qmur11iSCejjVjbVOz+fLUFoE
dhsO6VvYAQw3aPKM/yDVGcBsCvUYPSjxfuhHU+BN23l+u/BwKBhznzOavEQMgSFR
cjo2nkxDyEozvZrt491m+9T+Bzk+gUC0lCEv7Jq8gwTjbesdAkVUt0HEM4ZLUXiv
aaY5jJq4Imis4obm06EnJaVHxw9QdzR9xQkbQgGS67kM+zDzvZUpeSM5LBs3piMK
lBh4jZWF1jzg9rqXJD0+iP3egmA+DA2veOWbrmy+O5bmy0sAZCCdSKhA7WXYt2nx
+Vpn8+CVKumKuqR0jKAtY2ZTvnvxcoIshR6SOKrOUpY1KQFU0mEW0pyfefIMRX+d
jt6tTeYy9x2FJy/B0wPIkUlAgjmO7FZOckhUyhQrs5x2mTOnFgU73UzkLSYoKwEe
N0C9NU4ucTbAbFAgcUDv0cOGsM5XHeN/ce7MePnnn3iUnc7F6aaUROm26/3ux/Ap
vK/BYKuvzibhM78R7SwMk15xluxb8iA8qPaYPqOBupy6ZMS8UIwHqIe6TgcxGL3K
NXZI7wBTkC2+foqWjF+h/xpEzK9SaTgI4M3i/6Z2WtbLVeULHQFnvi/XhE/5+ftZ
fpETb6pmJ6VOMON+u74UQVleCjqc08ky3ZurJMrIWt2jW8rRsVM+Z+V13TyflAzG
BwWosd03Wy1zGh0csg+rAw9UIzZJQdsTZJzMoZXP8DTbO1PzS7vUhVeLys+LpEsB
/+hwp21hw57PuXs+60vkyzK0dn2w7ShQFrjioyhWkldsnPe660Qrh7fBLJbVE+9Q
6AcTZUgnsSxv50iC/p00h3DsbnYohvlZxL5SlcKXghIiVT/MNUCp4vX/LujpVE06
fw8gmyzACiISzuMuiE5fIP7g2/p99rDXzB6GZxPgHIIbWvPJ/LNb36P9U4MDGiFB
4XlNPvdEspoTZj0ULwuSggDown46dpfi8F4n/ZhJGrI16IglHa9laAKraaqh7qKd
QTBxwFUO4cPNnRbsE9HFgIAuvQ1TRlwdT5Iy26At1RhotmHKSDf+bdN1VmOy8yec
uzi5OmlRbfP719dbDH/Y9U8mW70KiOfilNAR/WqIwneHjGCOShip4j28Z98xRowq
Rx5YDQESFQVpwISPhL06mHtjecXnW3IRfLeq9vkUibd+3/d9tx6cotIl53VI1IN1
4cz4x38zAwWAEd5igXL/EzXpohu3yCza+IhyV4giF/tzwyyAfCOZlOSM1Q4b4oGL
E0u7BoGNmcd9Zz0yhNrYZuZHEaDooSHQ0/Fo5en2+e+VVNBxUl7yHmk5y7O/fqCV
yohKl8TIh3ZH3tnPjn5SOZTLDoG6Uc+2Xf7FMCxT4E3sZXJqVBBXTubwiZ1V9s+4
4i4x3zQZu5/oFhFK0zqtSlo4M02kkB68x1jYbv63oGUSWKYBdHljaAaA2Auenqfz
nb0UxR3aW3OQCtLnCcMb1XY5vR0u4l4WMqqu6Wz0xYrCfHXpGNiAYGYGLPweuAPD
lwD7BPnTJ5yNAcWewODph0gBCC4qCkaoJ+RPOdz/mIzQU6PTAQiJStrZxUTtzk2E
aKldVIF36xVBkNrqJLQ848yHHjkW4fPYd/eO1i3E3hxPVRkV7zJ5sRGij4SXw94t
TpRLq7hcMhAAB3he8/OQ7jUGdwK77uSQoLlFvRQh3OrMR4+EPX2Xf90tyPTycmOr
jvqhVdNdt0NdxVizmRJN/QMyLstFgdGxzyeCp3fjwH67RzZSv/S1NBfejHntv+Aa
q/PnuoajQuG3dX2ro0f2dNN/zg6BQ2musNL63FeIsSQ3SiGRYJW7dMC+Z1LegXM+
dtIiNZGf/O0ko1lR+2DM2BPjbEq0OiA0ebhwKZMTedod8IScYMwkmnMsJRDpSc0t
Hho8sHmNbJdMB1EskOlFyB1G1/fBpnGsO/s2bO3j5kTLIsB17OHfC0Pa+k0409nF
32oEjiIHwGwTGjJoHGIRtTWFcWtB93U8WuZXcJkwMoG6nTIZaBaVSDzW+zua64W/
tQuKDEhtDCwOwpYhSW9GpxMzWGjMazZxs8NY6tr/49EAlwerGCY0yMU4nYtutW3x
8ajJDFwnE3Hc7Y7+CZR62sQqJH459Bu4U8q4Ewr87lOQ1li0pmjaOi/tsaQNFKsN
+QkeE7xV5VD2HtOuII1NE7DUwkJj8GnxIYoLBOTG+Sbgq7VzgZBE7qAg/EODqj9R
tCxQjNG6fuGKcddhRfC7C5e6Nfj7ARj/mo94tpoRWB94MebR6PZ8jvHa5oYmSpF8
6hlw4jsvJC9CD33KBy/nbCf22IfuvST7FYUYrk4VhxedXOsuuSYWv8xJpB1e9EiE
/PLzsLk+PyyXii6T5Q/wu8WG+7JgcZ2NnRAyfy+0IKDNezVkpgojGkn6K5k9fgZw
SAINIvGw4dnrApV+DFq+oDlbEAMWP8MFwCJkLuzOvHSLy9TOP14PzX2Voal2rlgg
mtPkYJTmIp6OYbjhlTHDUi8D/0voqJLWOdDPvUD7R5YHOwARbHWrtMD7KwFff0VD
UrTekS86imyfniLdgU39NKdBMEJNFLUpwbNDrCWR1gHtTUmpKch2egDE153um+Z6
sA5BlwJyWwP/zTwoWZZ0eNxpiY9EsWLm1JekJHhrduV0Bm/skjGd4q6AoAz82lOU
wZvGgD6/JgaEzACVULL4Oi6yC6hJ+OrW7M7egyGMZldcu+mNl2bvZaHnQ4REKiDj
aN9WhC90NEeOmMZsi/O8MM+6aIsJzGaDH/A736zvTO4qjFPjhRmhuunNYHcCs0AV
fMhGYxpQ18g/dJiAI0R85foVkBYj8QmudNi59KBL6dnZJmsoBqts5ItrxGLRhYPz
hbF2T2XbS9rf7guOcfa8syteW7YnLopdm9MGStsMr4Xtnx+yLyZLLyUfN24t93L/
jnQP3DwPr9Xgem5FQhIui3BmoxQUY9/+y4uNqQSQOJOzWL625/EEz8L66dAh7dqY
8KWMbII9e9i+PwBvKiQy0suIQ3H0ETdsZFC8QYLqealLuF3xOEVhjT739W1L+TYj
oVIu4Ry2LekhqswHkjrQwIE37+UgvjeRSOSOedDZQMBnapyIHRJoHpGVHUsYo7bZ
L1PLVutB6zS2oPDE9XjyGj2n7HsOePFh9Eg7o85iZwUzv6WLUpy5puiyBVP/3wT6
0F7IoiHGfw8qx2zqJFH3FDOCC5frcvBMYEXWJGfEM93h1ms3qX/sAYgp9U74d5hJ
U0fezOMuPVaMoFRZRfe3RubhNb1JdG1rWkcllwbb7vzPbF4jSASz5vFA9v+vE9RX
wFRPbnfgohslEws4DYbeqP7C+soZ+iLJW+/nQlN5tFOLfIoAiLJuThqWns0ZbxQy
v0SZHYTBX/qhwCIscuIHxxz3+F+OKxUjJ0oW14BGfaf0haPbH2Gi1SDN7lyGncev
BNbJftcXMlQu1K+blZjT/U1ogfcVvOYk//QVBfmXIIEhMoezsF/f1i3Wh3MK413b
4kZ3RC+42M3eQUkV+r+1M26TONNyo3Xma4nANy07tD3B0uSPpwqMelwiBdVnWxat
V2AvKNgco5xXympl9uxEyKEVQjCY1R+GmQfZsmVVPRwMI7zPQQW2Us8kZLyhLQxZ
mWokRBlCuyLKoJ84UvXGJZqBmqZ42Ggdc6FpMlAl6OBV9JlEjQzq60/tMO+1jHMW
BCLi+Rd2spzhW1150ON/J1qWsXg1rfJlTp/teSgp9YPi927C88IejSf6K1ayhPwl
TYNRcMXi1ma63fowEfleju3kS4dJ9vYGKPua50BYbBwuDmzwLVyjzu2aURQ2tIlv
7JJUQqg3xmBZKrrZaJlP6qYuL13r+6Kja7hpLezMUexYn+VekAHxuooUempjEVMV
j2OjJUR+ROEXbqYj2pSQQNo/pSNkOLabEPClWhKwlMhYNe+voB+XHZx9MPg1MFUe
uNsnfwb1iByLJ3VV3DzfWCoVJar6labWkMXYqozhk3pETKkKGXVV66VGbunnDILM
bU5VcGpJxwLYsLJlmgIshuIzeRfVZnKABDB/vlffoOXvzVaTtm3ecgMk7WBZsVdi
L227WzYW5ioreK5URO8w3ql9p8TJkm8Z4QAiYkxRXm/vOLTTi4Ms9/d4va/ocavM
EByouVUkz8hQmkFvToN3gvyQH8TMIP0pMEQmomCEZdde0vP/RV6PcydwzDpBZ45q
ZzcbU5brZSkEShmxSggyO2KdWRvVs5aep65XWK87MwXxvW7zRcqEy65xn01altUa
BxC6vQpQBbRzkZkEiF2bgVKgj00Zo2EskHIzhn3N+rickfl3vlGKffVrMmRQym4o
F8hkGsrji2QYeQicTYL88VwSA+X3qgBmFU4IaKQnq86y0WyEXo1QFWgUoVQ+4jZG
ILV6107VYtnP63bF5jRpERzdJ0Vrxn3rXwoL/OLdOCBLEbGXwyuawByffd0H/YJa
pgM+OdfZPNv7kdKlUY6zPnE3nX7P/DyyX0nu0poF3mJ1pwWrjFTq79xjNCT9svpL
3/D0Vo+w7zfkkCEP7Go4pp/fQdeZS/BuK6ilvonVnqP2lUeC/r3hrn0ZeTBvg9cc
Q3mLMKxLYUipnRxWohpJQ3brSBnz+y3NvwTieIU0uSF62Pr0tWdp/FOlDyA1L/+n
4DjunDDIMfTl2b4C/pztqUpPdTY97ORwUqqj3r3fl8ZWXfc30g9mpBQwQPxF2xhj
RWoFWLu+yyp9JPtIQv2hmqAARF/4WJH2bLKkxl1CWRM/10qQjbY6nkAs45naw2qU
A5k24LFVx6W9RwSH7vt9IS16GEpXdKZg3K657kL+SHLHDAZnhgcANTpXOHYYL0IJ
TmmsY44Ai2aEElpJCLp9TlBOXQQMkBM2pxtP5fpSIJ38ngjkWyxgDrE9vAridWSX
OPYDCbI0NWIXDTGGX3NLQMAo9tXANBQLGab47oot110oUILQ21fuxGWIYOZnmQcS
klzL8IROvJtsfROmpy5vgUFjJMiWktm2Cn/9k4Ir4b5zsUMT0pzeVdFRovOy4/5/
zbmDbiChSSc7EZoE2Xu0hmucO7v3UeE0c+lKFtD5QsG3wnjRbz0PiSh9aAC2CBBe
BK1cMbtApktUH9a4YXn6kvJaPdnpH0OqMQMTB+KmQF9Hqhj/8H/mUf3u0zolgKNx
X8/NuVrg0DaCqU8v2KOr5VcMgI6knIgwpJR39QBTF44VQgVwaKLvd1GMLSVRvNEO
+aUICvjyZmKRSBEf4y34neg3XXT5DQ14+gUDqdPdek4XM753b7qQOjHkQ3G3cONZ
fRaeLIWGe3FexpeJ5W4phGeN66D1R0VH941V/u6aDul+Oq911dhQjypFXfMj8vYV
eXK4/EOxuscDIxgCafk81SodrdC2Dt5rI+xLLY6YulLx/jEqJXL9agC6fUnVv929
JWzIL9A3pvKP8SdSlKJWf81Mrdn9BnHye91P1oHDLbEZhPuUD9iILTzMUwGlWpMA
3jogy3dZdC9wkqr8vblns+5pPxla6urs3Uz/T503ExzUxt/8LApmXg9jFgI3wDWR
tPkW42BW3NerWf0rO0imgCu9HS0CP6s8PwCXvvHWSQsB/plq0jYYgSdyN+AgO6Qs
uCVBTw3hP7xV5ZycOc1mWfQJ3Eq15K4fQxI87+nzrsf3VfHF27sckfi3nuB1QoMc
FDfzDAEJrB4jh0nGXKiQ5wItq6OF8IhOniNcUsbKiResVo35XetXHCctCr5GpBSS
GAFXH7SOy1nrpnHUbw+8oVmGQJOBIb4c2POG3fD8+Low+YXG0Up7k/iFppTC1kEs
dz/o61L/sjdLEzJ4owwuVMIN/5GHDLsBWVpqiuw9Fihj89K3E2lxVhCH7e6VlNRV
Ts3ojHblfElmBQ1joxgzXPjw64bqjFIj9tc1dGYB4cj/jYvlCt3Qr1Sx8u4oSKzJ
kS3oUuLjg01sA2+zLlQZfVSw7zz9Zs7ruK089dXIGlJaqdleL1ASAhknY4hxhRD5
yK2IP0FRRD2atYmOBytfkVgyQz21h9AWTaEq6dPFNQeXTwO9PnpLsK3xtQwvjWIm
r+JutzkxgGhJ8ZMIkZf2R9zuwBgRZ5/LU2gxmfNLG3PG5S8yl1HhleQ8FR4R3NO6
EFSqTu9FlnLaZX577kCQJEfrdKTg1MYkFVMg7FL7TZplnYoMxyKpYUBWB8cnA/Xn
0Hi8gT4jIK+9HaX2TPPr/9WhTwtBaliPia5FS9VTdFhS2y1XQiRtbgKhFZ/xKGQ4
U8nJnzL1nJ37+Zv6AP09YNViKoH19aOCoblUTUj5oeZWNOaJj+nOXAMeoslp6g5O
jpYTHOj5r7AzRnTToVJQ3nLsmoveti9E95Pl+ahbJH54RrlUWjFy9rp/IHHLyxPW
+Qw82mQJFQZ8UMrE9LGTy6MOVD1yzpREeLOuBi0/1GPkSuPfJAs1sATKvGExgXPF
MWyrv6qD+gfOr/3pZWWOarqpCqSNNvIf6+WVcSYKoFjbXjYQgF9LvAoHSFGh/Xd3
WvhXnS9IV4ZJKx3OJR4vGOnnifncwoSxLjTDm4MmFzeZU+qoaU5CikurxCBPp5il
4Q2j23ojC0zXSUNJQfbsUd4kR1aRXD8Ne1XwM+QEbsz+HToWmdvWhIMN97DnpSRB
+h2fO4rA3Qh+t9b0lOrILh6d1iEwHBggGkikP9G4iAF0fSSQuvXNvkh4XkLl+yVE
RhJ04hwXmfNT2i/wAXb0GcjPdScDnACQmSrErQBYSkPYzlyMI0qCqJu2JtDrdB0U
G6sLTSUreF/3ZdSOyWcbghR08L7nKMVlzGSCxnbid4jv/bRld3NXypW7dnZhBJ8t
NAp2qN+bsKeK1b3P7ralSl1khFrpBtu6mTeEmcBdvKkXp4O1g2KXAWA+lumoLiQU
iSjmEA0S0rQIctHFEQr7DoKcbSQflN8dSTB870apQ9KQm789Fi6VoGt9Awb9yjFk
qd1PW7HMaaJXx0ZG1nFG6y0tngxWyHAdLQEKMgrT3aFHYnDW8oEPlgfFj/zQYjdp
pFn1RKD+pQsXp1rbpXNWU8XHW2yroROwwI9FlsXbk9hu0Sq8aXXg7QD6xfO450lm
TSysGTx/PTWH6fJwOLwP5VzkLsfl69L80pPJUHPoOdEzfoinST996JD5JeCe1NPC
QPHOUeScv50D7KbJIl1CefttPZrRdb0rGwWKZ/F1GLXlTF5YUbswccOvJtq1oexO
RBsgnLrXdTxhFrTZ88FjuphOYdxg+xItzNNfGDZdpnr7PR6L5N3TlKpZZM7EG/wg
otJI1Qo/k1iDLAku+wuxgQi5h9mCNQBAZlOMjillq44m5bPWAdJ7q1rMAgQCwZ8Z
D5EgicH5MlNxk58dnvBtflp9EAKFxSnSZGxe0phPUuHZ3622FCUn6e9OOC+ogc28
P+zuZsv2luaw4KRQ+h11h8DytOPSUhccchYLR9YfDr8kiPQfetSsdH57nLvNlPOk
44TducqAPn5HcOzKFnRfWftt5d+URHUh+Zzem+2+EDuLfK200iRod3iKcBgTHNrX
XH7tbL3XWnoJm7RJwJeMGvhoSGhliWGDlJMdalGa01QLANTFwMgEu2X3/NsJJ41p
Fwf1v3DrFr2RnEkOs421HmkMTM2PiWdeiJPQ/6uu7WZs2gEV395j2TLZk5vNif0z
UZazrYhmXbtFFYfF8UpLSSXCS3Ckui2l8i3nDdO2pRQyRH7taOgYH7PHL215MBqu
ObnS+XcicSFmouINO6UOur04NFPTLdR2fUAXlSxwmR32JoLYEsHDg9inzgW7ggNv
TBM0fQ00Dqz6BlhvW7n3uZj/9kpVxNTtI7TH9UJQjOQo1fJ7WC+jzNvQ1tqvEZ+G
/azQpv58fS94kQkAZY79D7UsLEj5Vs0sH2hE7F2Zi59toMI2yXZI44vWnFpLDQ84
N90/cpTDB7i1tdYAu2wg5FqPwOnRsSASsNSmaaRibPyt0ua+8fVJ0Z2pGE72jQmU
1gkBF2fhbxG6DVvEjYJ9pX/sgHWodBUKewPDc867B2/0sDa10Lquj5kuIjiAs3+3
HERk8w82E4W4I4r2tXJXsGTD9hUUXRNlzk8vZ0TmoKO0Ys06/7X10kxdRqOTkpOi
O1kZVjO00yMbwYgwL2V8gPNHQqrKU6C0rInvDN/kn1nuXhDNDvcwme4axIjzM+dG
wU3V1/C2WQAyzVyIZ+XcDNIMgwZ9DecaKf13xM40mma9VNjp7i5yPSPXNhTM1M1R
yiR5KeTWyPTfeEkhoiTOBGkIQYGlLFalar6s5lQgrEgtY44SgG239t1Piux/68Ss
Rt2HUCtZY9OrZi9+dmgITi9iILjNF0dgrELeA+Vca6ZJLom9rQp2eo7AguiKtBe5
OjLzgH07fdX4ti+w6IyihyRJIG9ce6IB+drhDcHAcB4dvSL3/28UdFz8ga0ngfY9
Z8J14Hh9Dbj2/uZII6QpfHW24IH+ZPdx0S9ruIHSA+bon1ox5SprirKx5lKHSb8s
GWZvCWUT/eSQNan0jLDzxelHG/wWjIVMtmWWQLGYJXozwa/2s/fxhBHOFWcMhoPX
nG8NJW0VqYJSbHfrtB5nIhaGBWJO7L6I1nVzANWZthaZ5VUNYRQupj89wHNeBOXE
oKWO6VsLYpVmYnVUKJL9zM4TiMbP/Fia4hy0yayxuJ/I6Irw5+FCKP0PZGYYQHRx
SS+bmBwz7B27nb0Tn/WCOtxpgrqQBevZAxzJ4HlucHZxEoeb8Tey05pLD3B/EkZL
MHCRK9/Tfjv/wOzDbh9ro8ex+tiNsYo/Bv2waMWT38X9ckeNLK2tCChQ6At688O3
vtkXJtSBND6Pe1H9mo05KLqMBSc8k5faAMP6GYZTiphyvS5wUHSz1SmV1ptPmTkV
3UFVqTeOTgzwJUkCnhZTRyDZdKxE2YLmJWfMGmd55xJKFiyFYhyLk79W7bEIiswK
LkR3GSIpPBzc31vUEG8XW6hdHNBjWubfY9RDf4Yd7QRY1wJdOj0kZMeTReYoKRC5
9kSCub7MHWcu8O0Ng47OXH3zisgZN0h+y477gkwdUHl9M8lkDQfuo9uJjlV9+T3S
XzQVE7yaEOk5uVC39Z7aoIbfeV6LOpHp88/6SEiiWiqe2h4JYL9a6lZOritC5q/B
qZggenCy5UyhH+NAP0n3tkuj8obX6Qd/G54bmFXUiwhd9/J0a/9zmvoqn8IczkGs
YPB5NhhXItcxXy4gfSiiUDcElj+Eaw25S1dXZp6fhKGM1doxOlDcpQHV3aiDbqok
EZKj+t8Sk3MOKQnXRpGJSTzVOCEgyJgyrF+QbTywVV/Ju9Xn8Ysi4oLM9U9+VFmq
AW8uUt0c2E7bTrQvHxfgTLleQ+oVGYfNI2g8oGsfR5Rv25sscVKMuu0nECSfmdp2
fx8AGGLNfz1p/Bp+qH18W5MXMV+LffC6g4YbvWSGU39Id6jl7DF/2Hh32qiJSLHz
fvsRxLYDL/WNLsIuSxxs87848X/SsWdO7zYfXI7+vf6Pf2FjAMF/DQyFqK/WZoeW
vqqhD8DzPS6FD4W0oQIoF8BcHdTSmuYvIwDKBA/eSOBS0yqHej9lzGM2SAsPHOzL
zpGqLVjfbWFpvEZaSbldpo2leQV7FxYqPqhHfXlkl/mrwey8+V+KLoLZ10YXb1Ex
rSi2exF27mlnYKToMu87FQs0AXWp08b0fpCzl0sVI0yrqkxy62WY7JLX4KNiV8nT
dp5zFLgEQrlK3+zc1YMDJ6K9ffOUxEK2HTulOXSeHaaT7IqPJCe77mrLKkf6EANJ
KLsOZDXjYO/DPw2x0cLBUX66kz8ndoVnndRERqqqHFve12RZ2nrd+8Cttfpm4oa3
VIITslFu9yQtpUqc8DuV8tgWwBlKwjT8Fn0zI8EwqgZAHdtQWQrxkJqSfIO3Rftm
OreyQ5OXznljfolw+0e7WiW6BcuXNUYy+dcgFTKMM/4VJlAqDetHD3EIaJVMiMeV
OdUzqLBDX2C9GBJdAF2xRjJRpvymWhXol+nwd99YckalmZScfo0GYkz7oj1shu+Y
pW5qSHH0Tj2o4p67/+qY2uQuFijo1dOUGQFuec8zfCCYtjDm67judWfv2SxNHxCY
oA//f7imcnP5LR4B43aDMDmSvCtBeWN5hpUYke8dWsYsKaLhPTIZ7UmGpF84FTaw
NsXLgayt9b1bTV0x5H467aQ0GlM7ntGhGnUn1ViDpvTXcJSFcee925zIbib3DJb2
g9eYUYQ7eLrw8DEF9MnUbg7ipQcqD8of5ceXwFO8BEWyxzHSehx372lmqtEwob/7
eVuPrmWd/NyIYYI+xvPfcGVpmK1SqJY7qePmIs9HxPhi3x3BdzD0wDBNTRdU9o1s
12kDy/XYT9b8w+QPEqjlpBOOYSGc2qsSr0Wh/Nv3OZGClZo1kRWkgtI7CfH8iBDb
zftYCSnGUKj0Mvox117uchNMSflS18PjnDRtbN7G/8+yVOnhhOINsDmSqkKCR5zQ
rkxCddP/mP1qwttEX2iIF5wsTH9yZf2lXImEKbkfwaP536BGnRr4JvHZClEfTmI0
soGzC6uOUWMbELVPdTR8a/jng/kZcznYS66aPUv6QeoMnNZDtgMPcFRmuVTItsTy
2daxwc7c1rHp0EI/Eh91bRpTw8PYB7LJf2rSLKOR0dcbnRWoDGGSIARyoadAo2ny
ch9T98/3wirByls8Va44eA3sY0kYRS4JGGclTJ32rQkJR6GiKJ4Jcil66GB2lnwb
pBOreKXuqT6FTczorVu3OWRF+aRhi8lztlmO8Hc6hIv4kErkGig50+uBha2Cfspk
0Y/SyrIvsHC1YtBGcwdXDHMwDMOmDnB96Forxshtfi2pxvlod5rKfk+dUu5G8pzM
iO3XB6ogf9P5G4SbJ+2cD/7ca59YenyHsg4c+4jLyyRAJ/JarDFEDlfJPWL+X1wZ
V6er7hRzTkTf4qRDrg9cC2p0wzQQBdWkzLnJL0knKtBERME4AJxbRyB4PPyey5Up
q1EgnyQO56HsM38kq9U2ISnTpFpo8ygPc6jD3YSdAhSg+wD1pZ9sCEvj9rhM++8d
stugAuPLhmBsrqmsoWBIq6V35RBvW6+M+38F7U6dD/jrfFDhUQRhjIYtAKACixAo
+CE6eFJ1e3U3YARGeXdSgbUq9tcx7zpMnEzeFXRTYMFOfKsGDzFXvus4RasaYFHE
YTKiS9hO/mz2Xhk+QbBMB+s6HmANJQH6ybDd8PY/xya17+ny814QdxIHKYpWPVpY
rcrIOI3OtU0iPOjTAEv5uobV6DEjiwOAi3mqnbhL7XVl+V81CVDyJ8S5+hGU3IYb
477j1dlU0LN5WggF9axuxb1pNmo5BW+NUK8EWeXmQls=
`protect END_PROTECTED
