`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OeqT8b/twEPtY5LpQMO0jQofZ4+1je8dWnHxXwTbukxf5chOJkjAkPInO3RX60eo
9CHfVO0oSa3ODUhex7GClVK5aM5yeJQBe6CKGb7VLpdN2oBuzJBugp8y7cNXXXhp
bi7kSGQOkyHmgoiXxYbfc+mDvbNryKqmVYuTMO5HgTDGUATmx6lzR5q3xKSn8/yw
oCez553z9BC86euND0ARaA00Xc2aSI8NLq+HqCArRFzgZtWeNYEt6dky9BrhcrL1
Puc1Tw+jrttqJuHGyCL3ONad/B+gNJJ9Dylr6nqYPf6bhUAEaCOnkRYhw3SQdfzS
M7MGYPGxcOugGx8Rt6XVOK1z1QTTbr5/O9eIJ93z9es5JKhAaCGHhX0dFjolFdyT
ixahqc/SJ2G1WgyRs3cO/zG1151lRA7elO3wNB5tm3W7Uw4zzA1V+sHLbmqU85+I
vYH/aDRHcYhXbvEISBjqvqvohroAD10DPqJRjZ4EGrz3opTAGa1t6RBQZneVZLoN
+xOoYjbmCziqQD4+Jlt6utIHWmE0XOiOnNqv+O8NLpPEn6/tQzm6pRO3Os2N7b1R
19kuFTRlh+60D6hef0pCkosXh6s7N2rSx4CvpYW3l1lX4CoVqoCAhe+DviczKRad
8/jLFAISEGaEAWhWfpONeVwy+ZzvJ4JeOrdE29rwLvT8k117fjSk7SQlHjAX1an8
E3h6Qe6XSkGEeiA83FpHdYYDbHmOoNkBEj6VjEf3BTj8G2RWnpjZ07ohqQkqakvp
UttcnCJK3kQBblo1X1HP4cssIEBFLFd5sY9LxHGlGyn57CFC6/tsGRoK3O9nxVdj
luYHphdCURRR2o4CNwyWZUGkuSQJdj+omaeXFd7CaAylbpzMccL+sEVWhEJK1k4S
mauKB3e6ySvJ/CYlkud7pVSXkDLIqx1dFh4uqExmZs9/s7znNbLnRfw31zIy/6YF
RYR/1fHZYcIF+qHt308ob00/KgyUcESFFK4Bbr0XOeyvuTfuY20zC4oJ66Rs6de4
opqWywjnolQBKjlaeR0Mq1zuCRLDfKELWtQFypY54MM22tGQSapspa2Mphgyn2/A
Ts+eu4XjtT+57MczMm9X2udokRA0OkbiditY6YIWKa7UF5iyO62QnTY8gX6wFE2w
qOOThEAv8EkuT/fr47qFjFE9FlvmWrBownyHaT0En1tcl+I4jO6ATq2PdxYqxzuS
lM2DmuNaD5M3apOiV2XCWtLx92+PbHdpJb48RvBPwVLuTxo4lvpIT+sKfv/VUWOr
hI1G/m1MSmo7bXQ024NR3L0Xw5OXbxnt5biCJi1vzEieUSP9m9ZI8cpRdCrupFk1
0qp+RJH5gLMSVy+lLWNznZzQzH+VjxNT6uC6j+o3blnuFnIeIdxQ+zEr8kT5PEZ/
1kwdgemmoLkPQa/u+UAYga6WOul8ac/SzLwJES850XldkDoarUf8xVY0XVNAstfa
qJkQS72DWup4GYKs6/oR1gzXcBJS8eqYelB9s5jSS6453Vg8wnnmbBTsORYjUyO8
/3i4Fk43NSG1zH7pWFvljq9aR+QQ722Sz7dQxXPc9hnBdWOglHmSpcyWCPyejOz9
qr/AW3o2IY/3Xi93wLgzWLAYYxPTYaP6pbg0rwL9V1li0bHBDGgbT8Iq3g29F9dR
JqTGOGw7uymPHDcbYKPUmtgjQmiZ4rLnUSKPLtjCY7YqIsCxVtKPK1mH4qTifRDd
CuWEdZNo0fnFxNV8uFiHkzMCda/37mF/TirK26DoQAj7VbzeGAXFh/sdhtQOlkP8
jYLXD0oHaN2diP8T01i6KuQ9tQC5NFR19zvfyWItFLxxw4t3JgVJsRmfFh55guMu
xIuAjk1YOyAGXV2HJ2luN2sf6QKVfP6n/DBZnR+5MXdDvYV9s2ukQxItDEjqF9jF
jgB3iCm04XMEYzPeTdlHH4gqWv05MlrPTnW/bOLBZp7fjn4D304HXxdTnJpG/SEo
AQzN6C+oXj9i0jURxKX86tsEvTbX6BGtVE6j+ZBgyrm89incjMPWFf3yhD8VIarN
vU3D8Wbj5F1wsFsCBsCcgeUHn7ij55V0Si7Ml8k6U3W8rE/lHSzD439axZYvpGgi
uQK9Ck3NzEbaIxzfFuTPQb44tglRstKn1sqgBUU36U3jjIZkp9mOSVxut+Fr8Nxp
IRr9jS4mPinfJpi6n64PhAr5p5A5brOMB5m0OgVyHEg4nxti99irgrnaHUYKzepL
+i+UBBFNsIi7AqEoon2yp+X6Wk6niWLz8m+FV3uXakKMdui/R1WyeYEyPutjwWBK
BTdmWppN2oETazUtHG//scXE1xBI4RHUGAzBpTm749OnHoPTAmHsgcueYmRygoFO
psvPqJlHr92fFxjwGPN0UKbU3LZ5AsVU3wgGG8vBt6OZu19cPm8iGGpNzHTFB5tc
eJl6WrOixgefkezSDbDxuLwd6tKC7hWjkFGJbgxeyWJejnbSe1oQF4ao+/zU+jPQ
PNoyCppfm0lt66pwk6rS2ywIH5Vbtt5oAznZbiCvSCvnGibTy+lZq4EWbu/2zC6l
kNudwz041077rjEFd+3knm/haI/8JMwPFjFB1ahwqlEh+mhAlBgzJCGD8igWwZce
NfFSL4Yt9PUJp5kbsFROeWyN8tRoKMNeBH5wQPg+0KkR+NDQKzqOu26DJ1XNwjgZ
h0cs/pcCoHdroy9/n5twttk/wvTySQncifpO13fK6UGCQ+hrAPh24yctTEYCyFQF
75p5Llvcz/vra6fEZU0kkTIvLgXzYXYo6Wh/axXcuVQRbBGQDr/bvhkhjfMVWC0n
U1105rVu4Nbea4yxArgV2opo1VxTwwcwhZcW9DNe0kwoc1dIpLDQfv6qZyMieNxS
yD54ceNz/MMnh4TgPjuC18Dq75wYHVycd+SiIyNIiufceFJ+IlUjNjipmUM4fV0h
z1wUxA9AkO0Zbnb302sCOAawBLfAHbkbcsbAQP3c+Ss=
`protect END_PROTECTED
