`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Mw755YfIskH8uvUS3BQOH9WQAK3A4anK6OMblB6mMQlWFJGOH2ReWOysyu50llfB
ZbO6QWe7Vdo2yG+P2WDAMQ9KjqATCoOL95lVTjvmwGamTU0dPNcDeLhsBBUHiSxO
CaN3NuS6yZzXt/7Qmm0jwKkL3UAsgOPy13rEk7b855XJWjdpiZak6gKOgGpvyp+Y
1YT2Nuw0rbbqRp1Hnn2OimHQ4UCBW287K3U2+bfB2se1DluZaF4ZR6j/OjmyS1bv
iEBdwIFifIrhoonDAfBeVQoJl98C9Z2vWpoIW0luIZ3/hCnb6VECWyY/vw0ECROL
X5AY4NgjWtmqsjSvG6scpSmF6bFZ1MbGk5WKAydLU4HCX6IfKWJ+Xf/ys2K7dP3s
MCEfTwFjinWpRqq/NhmL22mFk8J0N1oCUCFh2MIFgFHv/hiZysZjD/hF2nQImmsL
HE6WXP62dXRjNDw7VvM3rVqELfCjyFMOQUWR7C4O1/G1pKXCi5MG9TygiZGFggcT
afsb3P6lKXQ6iIDA/bBuUgUHyun7EkszHkkySG6N1g6Y1ENaSKy67BaY6Rq91nMr
Be0xmVhM5B2Z0HcEtLKG7qrHv4XCwlvXmQwBmh91DY411ImXd278uqJDqUhjS8Hn
bCNzpM6X9GOS73dtA4YG62kMfJpqzSOdgioP8glZYq+jZRRyWWbEaPPS3ZPeMBJ0
BqUPIeTDdDovk/w+Wr5piQqJTVPpoBJqS+OjByDhHs26zw3MWsZPSSeYgUKgqx29
r2H0Tjcd1RqVhzXfbNN0prV/qTTtNGw867bE6eEsFnEPSys6j/52YKFWD+MlLGlt
2AXcWEDP6kUtHFVgXap4SW6mJ5aLSEpIkDbcjPaVAMYlXzmNG6IgdxZJ8OnRHNck
grzOBWhz32AM2H5lnrvF9+dsePN+NiIIHcLUIka2kHOa2x6+NarysUBa/kpkejji
7m08+karp0qeBpqbMX6b++T1KkVcoR3nScjQVmXg2DbmL8Nquvm/HOEF72Zzn2t9
mhj4jRGYXEFvtaedmZ8FHZt5N/ZO9urZzfIXmJoKT/UoYUh6tRvw40yYAYarmllL
EFaVjQusBtqVUfTS1Q4Z9rfbrBL6npoxL/qttFPC8DUFbpERfVQrzDhR4B34QMv/
lwONnGrEGm9V7p5ja7GSeOEXFAMa124mmVoS/nbMx8LZpfpFja59My/8qeNQlaJl
dT2ljcFFVPebsLd/+5eiECRvyV/oj1JmdVj79doSB4J847b8dcgTgqKHmcJG/cWU
l4CEGl+17KPjb5UwYzSPOhXdE5JmHxgfUwJxwmgOVUK9db1UKtdNfNbrdFEsqTBu
w8U9fAwj4dmEqTzvHeIFWNvu/UgDIR6c/iokUs2UFMp0bs/aRWO+WQmlptPppjzf
0d1CH5T+Z2iP2CQPlGUU2b3xqjMZbZjwRmlCpp+VDgqq0FE8HFEl0Zrjjm/8r7oq
L178RnIj+UNE9V2ZAEuRpRJnNF4OKlopE/f4/+FcpZ9uHZq64TI6L8jxCiLhvx7h
pxR+6q6AEBSlaIo0SOHemzy+VphJBqyLuXsUk8AYQzmkoOAI3tDm37cUrHnZy2ru
sIvUqt+kyJ+2pXkq4mPhuRdzwTUDQCrQuUq5skws8JaZSbf2QaSFCeiZI+IomjEJ
XxCDb/G+JaIbGVRbnW7QGPEgr75tk16hZTexkgjsyE6BRmHihijNy9ied6TR7w1U
upFChbWc+aMa07dUhHMxtaPGUyZBGj3RRKSqU28DKuRks0X8bhwjz9LRnp2BVa5p
d6LXcLKHGsx4cL6QEyW1AqdvjLVfpwAHT5KbUHgCN6tO6KT0cpzSp6R0WXvVdbfH
3C0vugHkIuLu/Va5nWDZURV8t09bu5Y7KULQwr3UdY2PmeRV6yAvi08kzLO5pZWk
sehoQHw5DMg6JmIbyGvTz181YDGKEGQpGWeEQouWA/B8pJ2iaW6J+KMM85GJTP6e
kCuYGVn9x9sFl3H86D0MU9/PY2yf3NpVsVnSceDtvTuzHm1qHvo1N4cMiHAQpfuu
781H3BFB/yd8tg0CtfbUjJG/ZU0zHmZ17s2Hqx7FQNpgfmqT4D1BgPBeUxPRFWnA
mkWxg8Ggdr3/smkAmYckAnTbD/KOeQjwNT/BLzGOO8qN6UAydGYE+i9owktTU5VU
T0VFXKvqOB5sFpIdaLTkqOjz/hZJd3sM46KNOPW1SQaYbvny0zQZnwRWbM7bhAMJ
6vt052qJomz3Bg2gp6DueUVZfscO35SE32F8kRnLoKSdbVKOdCVQ4LNS3cVg2AfS
YOzFmy+EvP1YeA54/7dEbQTYwXl4HulsGikmhwERujivjZ7T9A88kkTJmB8fnJAG
+aoVMczc2d+9lMG+6fub0nr3u08aG932y8dcLzLMWhc3VGZeacaN3cve7xLPYMMw
TZnbwOWRHDENZ/4cET6y2JSeyLwI+eg5hgiOfS59RaXzPAiQDWZZSjeediW4E5K5
AuiQMydX0Ykrp2Sf3vZVx2IdnliGxa9BYmnPMGTgpg8nAeNj9lkAl+wn8gPK5NGl
fN0h4qEtjOkF3cOVJnayP9kwcv9IveY3TOzMUEW3M3bxf0hdrxGLdJuzYBftzsBY
3yhhWRSoPwOr0KhWUS4nYYk5pvB5+9TzfRRDmd28ip1tAbX9NKjQQ/+NISh1gTT3
wZQsTbF47PN3fG48CMyaMFDbviD0Uu4y3mkNzbWOrJoFthQzA8/wJx+SwDAyJJ94
K7BUAJnW2kushQCqpzpuvFijydBbSUMyQDGD+ZeihriJNTUvZ5KyBCyahQTArG5z
LF9pdaqO47IPioGyAHwP3FAJxg3qpgUAYqMXzp2eab3axLNyY1j+uhlS0Gi+QnPg
obUvtMukiloEOpRcZjSprmHpe0VzsiWUceDsIMf7fHei/mNqbW64lEJ+OtZc1OVu
OcMLxtgspqwK0KjIfES4XV2a8IUSzoNsMj741r+GzqUga2rhdICW5PG274LIoFkk
emX7ZsRhu2uwGgWwfuDuNr6GjS1pUQyCx12PzELVciGR6aGrXafP/mDgTDNlKy7D
tZ4YeWxlaEfqTt9cJeczhw+o2D029UUVJFrIBU885B1psWnLPBP9yLB5612uJ2zq
UcO2klQtYRxckbn4V5Un6TzO5o3f9Vd/B1WvrgOe2Ui5nO3gRDxTaKfAYAgGUu9i
jihSh7jHuEWjczY2IyogSUSwzrm/aCvmpBB8ezyNGYS+IcCRrF/dDYL7ZbdXQDkF
pnCfx2g008PWMquvURlE3tzFiXXpTYNMnEpnBtzJjsTFzXnPxR9wMuhansOyr3sC
CZmNr33DnmU7lZlXu1PyG3fDSx6emyOEWADk6v2V5flMsPvd7RtmAjDM5X2Ta3PV
an48NF3uV6uLEvOjSHSbjPV0qgdh5u1RtETXHtwmEZUy+o6yWxpMwwuWc0c1lC3W
73zaDkws9Jn6bORgBYKYp9QUeBXftJPoU0rzHK1BwlZXWo1g0zTB2zkwNBzEjQqU
rXndZp1lw6xzKeqdKIKoh1AqK97FKd5Vo8OmNCYE1VmZAN/WBD3tW6myrByw0gUb
RhPCz+NRInR0Wbw/pRFE76jDUD4VTol8DmyvvIVmp1Z01Zn9kbIAW3qKqSqeaoEg
NABwHLCRDHrFGu0CJYSl/MNjgZiV/Bd9C20pK5uSGH+SwjdfBGS8hH41QxGED3ia
PVKM8Ki/NGNbuV2jLznc+dwD7NfDL0foRavZQrKAV980AjRavai7Mh5QPSuok1Q4
CMszHdP47JvqvZs6ZoSMva4gArvgVTTPU0WdWgTG+tasyn7c+RIpk8ASlmqldFlJ
M49Edt8yz+9QcLDa10/sWLU9B8vr0/vG5vayZ2rdwOuDD8Mnr80fC0yaKIAYA9XI
BSlRpu7mUGBznEqCUitJ+k/m2RUyZEatuCI6eskyh3jdlnpgd7QAtjARykcAbXTh
21z43oyyQgWrvyPECyUDz4n6piX0n6e496/tq6FoUpKhm5/1uh//gpGza5DDCpyP
Ol9JtCPttCrlUvaEOMhE/xoUh/mDRuqwqPLiHp3qDfaA+/6LokS7TOpL9d19Qubx
AVZOL3C0h1Rk4h8TFm4KTHRLAry1XBZsUiTbZnxJFxxjoE6MlqDEVymR6+X6mQL7
IlA9QSvuQmlGnvQOsMYZIcLNqmqUJFtMR/xR4hm+ZXkSsy081fJa/qHyZXPKlUza
UoiI/CIzRvfc8/XHR/70QxsI1H0D4FPollBifR5xy/HV03TBHgpW06pDpWBsDPYX
ktEir4xLi6kWEGjlcVf7dT3f92Q3aTSGjvj0zvRVy4revChT3XtoKXzJWsfrNNZK
UAg/EPvjbgISvA6ylllQiKkrjXKDklDRnsT6hg6IJqQSA2ROXlSvlBy3XfMJr9MX
Dzkp6fiXMhdywnVYDbz6tkjEa1X5BmdIv31b7JrTHgYe0mYlb8/YPC/Ct2NExjaA
EYDrGd3ufzWDVzRu+O83mJLtI9yd6BrSXGG4Mu2iXL1rlB/uDizxRtzdwSrdbVxy
ztNnDkC50QGzrwMlNhK/QFAprSZt8bpWvRbLpAVP8gRS2lyae+u8GUdCmoJnadHR
EPc5hqZqAXBsmREPKuicCaF9hONwQ20oVyzPeT/oD9/L7NUxYuO4kMtAd8CyKX/p
EIwi7VWp86N+spiKlihnROCeR46XBCe9CMdHhK/vTeo13lw9KZPDdFEWbhZptk+Z
KyZ5aH+YHj9NanXvEEUNFDEMkzkY7FOOwz/qB8BL3O/yV+OL35GNfJ+gwqj3NRwE
mEN4732ul37cj2h83vXdvwAAQzeyh6Q04Wmqezg8W5+lsAJeOAwBbwGFPg+xpZus
qk05e7tIlXwq6ijqmaT3+Ajl0NF61NI5+rvMXCE0C5HTS7gcYHpXJHookrShlPnd
T3JFQ7Sk5+kua+38PfbvSCVp+WH3nrQyG3EDwnQdbc1ulesZSsoYYKaRasega+RK
+MNWGIl13ALVBiPnbQVOaELTRRlO21Jm4UzYmJ2Wc4+s3EppBmqjAavVQxWA4IS2
8wsI9hQk64jszhA5gA5g7v1+56i1C1PAjMHCeuj8tgX0PiIjV7TpLgWo1ZELTpV1
D4iGifhXHT9iWa8qNmv3J1piY5HUCWGAHV11QVP1eQdQDFze8MTMThcEUB9Sv1hc
ERP/5T10r1gySJ4ALHE1MJC03fPgI7Y0CWUxbNB8t92ySOXSXdA+wNRDh2FVx1xH
6I0bV/wS27bL/2ah8RdO2PxB7CGxgwIsVmtNqvpDw2dHWRK6/vbuzYB8kuUOZHQc
bO1ezkPN1dH+q1VSz2xTv94L8di//TMv0sJ1JU5Fb4PucFxczzqcFvT4u9Hn8wgH
EfXw//IPLTclQgS1bt7nwxZO7yWCrcSCD7UHgjlGv1nkWWUfJx3QZ6GwYs/hh5r4
p/ijgtrZhpMGCylh29vQYmA7YAJslZfWc3nRH6Q/hIQE9zLXXvYrqamyqi61VZF7
MSmSAoCIIzax1lUtT4Qio9fwshWurgsOnejen7Rh0YxoN+5ySQyzQrK4R0oqyqe2
/vPwf6PasFcZm8klpyAPuiBsJg5tqlLm3OaC/cPMlO7iErD06o8wrr6cjjCir63p
OMdaJ3VNTo1nBShEgLy4ncVbpak8nXo9QGYggXbiYP6RMk2uJ6Ro0zSlycWgYaWy
XjwxfJX0GD2o1GatRjfJmyBJ3BvGf7sY1rPmoKckGSLGnbs1kR1CAyL/grnlBnYe
w+lvn5JvmXPkAZHNvnrYp43j4brFH2j9uSKSJGDIzrsv/jPqY7xbFdR4r6SLIJyN
DoeSJG1B6vohSRlTsrpubIGXnIrsF4E0gijYPp8/OOh4N+LSQTUIPf+Sd4tKVwYj
GAlbgWI/8s/H0+s/TojaFK+IKkPUjeK1HkBB544TRiQnjJNxlmW8Jf3iKwy//RH+
yYfCrGHZIgUcbTjz7dKDhHXhBbI82sGM/uX7XbPJWA7H+s6ASzoQfojyptgBtN4M
InNTbraBuf9w5f3S2kKRm0kFmZRtHXFpf1AFqd7CmfpapNrKQkx7OWL2ZcU+OO9u
dH+uztVwG2JDUzRLeFna6+02gxCAUSkktrHC+2O1oNlFO2IU+el6EU2BjSUz/TQx
7/JuiHFduFlih5knJEx9JxG5wM5sVNjv+0gXHmHHHoV3aXfAJJqodNXRj3SYaMWW
h4svs/zuEZRw+x9jBZGTOKl5GwUfuKuYygLODIMJD1NrkiAVzkWiPuE2irFqvN0s
6sxGitxLwjI9U8qFUqW9p2BuyJsNHtef8C798wOQ+n8r9LmVFvq5AaaAm3mr3diE
YkMlZcBcivCBRiZnVYZEhsl6XgGjvDCbdW11GWHOmrq08eJ/HE8b/WMncWVz4qKv
ESSWQ1xA4YzpWLGGtoL+uSVZXstDdWZcrx6DrSimQf/ZQZzr1GMtkDgHV1BTw537
KjB+OkB1pLpG4PpJV6IhKgC7S0Hr7qs7om7fivK1iEQARvzo+UyyWB8PRf6/E9JI
s7vCOKSfTGeTUuCJ0KzGPDuwlPRxro0xkAUInwRwY2K0cHo/jKLuQ6JFpo4aCGJd
liVT2vnKzxEgmqtBVt9oIEimacJpu5fzJniaBiUGufL1trx3bx6BL6z2ckI7BDZY
G53+nQ0pD3w3XlAi+be6oKfJn1CkPOvZxGrjbfjoz5X8arMXJyrZVMaBqOPzGk7A
Q3K/wg48zqYMNU9mtQpbnlKZb5nGcYap67DjYDKYNustXa7c4xHC4A9J9vzVDWpU
PPiwBcCMIhppWwYx2KsMaFyiEOQmdHOiIoR4fiUkeUDmVsddYAbfb/+mKbqHFw8C
oerKzwdP7NubzHf0aTyR0W5TOe+hgoH3ss0QXAbNG5UwWHlmoRsEFyKzcVb/mq1+
HIKCfGSYcw/3qCc+HQCb7b00tnXKdrWgDxKmAwNlqW9yRFRt3VA+eCgg+O+8d9Gw
239jMVwe5vHcqrho6gjZhOIsL9w3NmjHe9I/8zLm1mXxjsnjyrBLvXic1TXD8lr6
ZkFdelE1SV1NPlustpG/kS2bfGjIHYl1ZgI7m9a1rMsGVfA09zMTORuEmEIV5jJ+
nAu6Y9rpIgeG6HMbgCTOcwyprMQBAAQ417Dd3xw4omagZu8VUBTh3qrPBJSZ6/Ka
IuUMixN8849VgcOb4JSzCK9dMe1B81tH0MQFWJkCJRsx5Jas4brneRHFLEXMor1O
SfAyVkrIHpMKTA1LYqPDCXt8AZrNbSz+cB7I1aZ0esoteCjHNnuo/DoQ7cObDWaK
JTeWn5rE3E77YmEo2eMOZ5fv3BBcAzgeQJCGs27kMtjHPNa4lU1+iOxEzFyQtA9u
9cBkW4UXnWzNwhkm5h50oVOyRP95e3V4H2qMs7ZJjEM0LYVA7wdWZQ4rJLwey4NZ
Z7f4XQW8/aFbMpGh1TvcH+Lswd0f02ZtoDtpxIspquDT4l8tlvW+DwjhgzxgBEgD
IZl0mtgfoecXvN7ddVENADaRLA9SZfur3thMVpODEpnNwZ5FRKkwKR/U4XPQec90
7unCESgevoSE3OCqVbU6tCqEHGWgyMFaTbA2VnCdu5ieQuR0MpEEuqivAjFsTNCu
QO59P0jewBX3Eof+jmXw9u3ePvjbml+4B3S7QKwzgyEbEbVkTQjukZRPBzzv57RU
9bGVgQ8NcUXU4xFI9v+5F7Dkm/BXbP1GLIdXf0KFZBQlTFUbS43ZNnj6z3PM3AqL
DjP4gLBISy6dqqZt0ptva8ejJixjCVMNs7Ggq/PkRtAS56TKKGVj0NreUqjlecQ6
T4bXXCSWWrkbyVMERHRFg1Pg4eYf3SPWwbHU5/VB1vPsCyFjt/Nq7EfnibLDvGlH
0d+jKYT2EBeoZgF074WUWE4Rvwtiy0lUr6LbJ8jv2do+mW7OP+iQOs1C6ycciwWA
Xca7o857mAjlgcTQa8sd4FOUSwyJvLi6x7zTRFsfwO0Wgo4Zp6ArzWLXPZqFwYUd
UpK65Uq0bXisIt2yCV762FKlx3YE+KmDB2sNtO7nbgZnx/o02uoB4oQedYEqWCpy
z6AOsCXc/3AMAXmxsxlISn/6pfjk9FFW9PYyUhkExJpzlBuHmV4K8JPBnNn7+jMt
IFu6ysCItKa6lM3f2pbPCOeeERZpepYxzwUnBU3/hALjO8NDm7IQmwgjBwiSvvzO
ayVWNE4Pt8xs3Xcc5lduHvlCvb14lIc38ChMG8aGIcwwvppiTlp0Br3M9jTHpjg1
XrDj5gujPg1SSpjvSooPBBzBNb0ZJVPOmeBwVoV77UswZq/m6Kpbx/DIRFkKZL2V
1zDErWBBTl/cRhZvySZiRT1/utRZ4MObueI3M2mgchQLgHDxqTBJKWU20HEO3vP+
TQnwpw2xFoKK06FYy4VzlE4WCXdDYl0EssAOBZnAPCRhr7G/sHsDMQJIkvtHypHn
KDTkl5YQQxEsEsgH94sUcCONvFuHfStf3y5z2BkYOHdYWbC2N0HKI2Hesa4l1tIk
mB17yj+WDfC3DdG6aXJrBh4VL1i78nrjOJ7MeMwL4IwREXgTH7zFO3ebBzFh+oDo
DF+4YLNl4ngum/tUHzdv1JegldZ3zv6yqcr1GkwNnkf79QHeYS8Jw5PVLRMnDK4B
/dWOCC4MKUq3pU4sgUQ4Mn2q1FHsToRJqzmB0x7wWAOhCJ9pVZbBmhZJ4VmBpOjT
xHF0d+bCFzUuuChrLOGlA/zrb/bdBQ8ZbCDH4h2mvl80sjgpHgO85MaPAh06wpni
/BKgjSI46d6nS8RJNYYWDGJ2hCUc8pIIVJdqflrvqDZdl2sue8MfUXZDTiFvfnoo
cETXTvlX3hpUMri0MLhK0GJYUxV1O0N9lnobnoB2bOD1I7UHWTHv69tSfH2n4OwK
d2dX+ZMZCyYr+FNofp/wVgIEEQQRRI4j0df9ulHsWXepHTuIjsSceK0iphB0S07u
d/SkoVGMyLHkwCAqKXcb6bOHBCO4Bvgl1e5EweEWxVTIGor26tKk/owH2vuknB5G
TkUnCP2ufzTmiTKvpGKR0k92Vt3Vn/Pw7EQzRSFSi1kX0Io75IJwBinJDgybfrxy
oHN8RLSnF9p4niLcIGymhhUOe1Cy6s6dKF1b6woeJlyOy72PdlI9wNFMniDoIO6W
N48KAXKqjgdMDXssJOAjOjCZgVKVHiBpd8KqYmgT88U/G9o3jp5kw42QkY/c6RbQ
Ho0x5tDNJTI2Ee4sm4Ku9czwtBiAsy3m0WjbGCEo0WG7Mv0tabFHZr2iihKPSGDH
qylm6mDkAP0XenqxltxW8PoOe29eaGxuCDDepzdUovvyY0y0Q7j2RsE14cHEnRLx
8egXszZTiFbjVxJBkZbI5iH9VXPRDm2DMIVJw8xtyjDoKQDnoz99uf7FV/Vvtagu
an/nCadYqakH+QEBJ+JinAvSxDJcZQNzJKrmhZJm6OOQffhtkZ4Gyw4z4JIni9s2
uPbB4TA2qVQH5V7EwHcXbdPtojzGtm7dHzxFsZPestds3dVwcRY69lP4+bJ5uoZv
Nw2CIYHz/78XFsoPngRaJUdjiK2fCjDnrM2lxDoMqqj9SY9xVv385pmboX4JkIuO
0TkfeyYuC/OMexq1Ha0x7TyyZneqRCshfn5jxis4Ecz2QcDWkE8SgpHvTAEdTIN/
dYIOF4f2dU7ibOZbjBtNAa6UCuaOUivZ6nwwyCACgF+mHhz/QqTQUSZC6Xmj9tRw
ES2Tv/yeksB6YAtQCB1xP2suJBzE/ge7Lcztj7xvGbK3HjATbehcoIk/wxg7hqxC
06fSaiP+sf0gQlrl7lq7qO1pKkh05kMbkzH070l7FZO0ad2nnj0rI03urSSh316u
lOMpvWVOTi8LaPx7ffo7iLWTWeItcB/91P3tG7cHHS4sp9dx2cFykol4CkNoPAJl
YSfuCMIhXb+cKWkalTsIHNR2Yu0+CJAKCLfm+IKf2ZPyC3WlvoUqhl7PkQthNels
9sR0WEjtlU2BXBW0s5e1I3LcTdSZSzPUGEpYyrrCRLShHdh7PF2BWCDmzTRmNumF
IiEHmkoMV/FTve3k08UFhHm0OZO+TYk/b0fGCbp6Hyvqqek9YXXpwrC09ph5KGFF
aflKUXWKAcZGxygINZvD89Ae3WsvZUloWkF9wJdNSmwDC3F/Cq29QHk76NUTD/DT
ADAGks6drrEUEuYwbRpN7ebbLInhp63TGQMijNBKHPS/y7ypsujxmIlXPHdqgWMF
WcKGyg0mnBzKxZeVI6Zh9f66mhhUIXRglPu2HIKffi/FOECrjtWG+NkTsYpNu3nI
AstKXGaGDQGVHTWIsEk/OZ6o+nAnhbiXUlyVUIRdbj83i69UMnE0fBcRlqoXI0Rw
nZBJ+/O+cW0ur12TtlPNRn31Z0+F72uzhx8tTWsiSd/AFVLyZ8HH3ZsmwCCLzOXF
xVZXm0X1/GtvZ87wQV2brjbuyOWmfiJ7G1IZv4lV33Su276cCx0MD0OYn0Jx+u2B
p6nQiAc2jmQKx4NvVgz85yee+le2q+Lssff/5PsKQbbJtny8kVBDlDyccNmyQ9D9
wBUg9AyQBThtao62f9JsR4x6yB1TtzTVRspMKp+rWkxGbZHOYtOjdBZ02tVbVZti
kyASlzZUy9LflcL+VtMj0wZWcdlAlHbv/9cDospvvfY9McYjR+aIX8CHLXMLVmaa
oY8Qll2a69no4h3SfI+PT0Xi/gcqIoxiCCzMgSmxX/A1Td0UX0ZVX/QqhLUAbUKP
/BXnvtt9YDuF18msv11OhtrAOKi5pskuZiDCX+WVCLK20h0nGqQn/pEVnhkm8QCu
3ng62SOgfoKsJG+jKzFnMqNiLHNcGLmU+zQHMSLDvgWvrAddO2gKwX9CCWZo0usn
Mti3tKVd7Lq8SBX4hKFmxQtg5b63N2RrX34QsWK3L51a44XLTYlCJ0Rzkmkwlkbg
Ka1Et0dhkTJK6T8S/GWnxtNtkNMbVW/pI35kpIDxQCDnq923g3X7d3yvFZwfnSjs
FLD/KUq6oN2Oitidq8HK1vv76VDK9KKwJZA0rAdaUBlAD3hoLuNH31EULBgKkbeh
fwAHqIcim1sCZ62+md7K9dfSwjy/CtNykoJHExy82Dbs0hhKSSrnAJdWXvr4WYht
9Uz5ahEcJrsQnn2lqIa/MaZ33kOQyws8p+ixqC7AV6S4LIsb0Woo7xhnmlokNo6e
SEqWPs2DnjwbdXtdS6en2Qp9fjL+cF8s77jFf85ZrrXJdWou/4wxi136gKoIxOkh
9xI7vIa/EBOmdZUAqqxsWcSmxI0Ipg+5/L2yDd7JRieFZQ20e2MZ84yE7e9ebmON
mj5QF1crwTmKFC91WenRMgauaf7gxnwMYIQ8fMjgb0S4ppCeXsKBGKEsd6F5rozb
98uCTRUj748C4yWb0X8hzqvFf5iL88U7igbTncXfSd6jxQmjtTR8nqDt8ZP2KhR9
NANbyKZ3awN3D8SBpVpSZLHc8mLDtcnawULI52/HlnlE4qvtSEoMGCh7QV6vJuIE
u/RpkCC7+O/oVl/azsO86miCAb1FIvz/BjA3svr1N7ZukyLrBnsY1EAucMBpi0gG
m11iH6ZUOTD4rT56zMGLdoH1Xwruz4oAfztR3Be5Scm9ObVOMoaMj+ZnyqcrsJp6
kwMamqZ/K0ofva3O5OjzysCMJ9k9gXrLfUGHatPgGfSONuU+1gueCGtaEBNuvIyY
C6+4QyD9ILsFBcsqufyLc/tWefIKu/Zsff5FFh33IcMVBoH3LHGJ1i/oxSS1XZfn
bemfGRzC4wF7n/gY73W2BFzEWRGKkM4quimzEatAJ101FyK5d+z/i4sGlWfWT1Aj
9E0wXqCMWL1tlMpb5+Izwj3yomNT6p0ropasVXu59k01iiQ91uLVQHus6e3PsIdl
KqsV8pz3Kdq7RN94gMSwIXGiodnAO7uAnTdrsO0CMhIMRQSzhn+Ihmfls3mbABjq
Z7uwmb9EDVu5N8YnKwpLkyqGF0sQz81y1HyYqL8M9Duja1E3iFMpQPVkswiDr8JW
tOxS5ASFTbZnrStTaig1KlemArMYSLPcnSk0QaQ7oEjKEtcwIXt7+R/i3M/r7+n7
5ch638YKmpsY0WJ3AUrhN5rYP8UZ4gybhqxKz2XY2i16QRO8ZiSH2eUqdZYVruG6
zgMJLNR1NqcjsB+fiUIPyKOXyY/ITNUowsi+N/WvapV5UHekMmSuxX74+dVt4LI5
N4v2wwxoqriP3zN+CdtzwPRO/8S+oOLmn7a4CdEr1ISvw5OiY2vwHvL/cSthyVJy
KBWHGjrmUVJQtle+x3zMrcu4zjdYLnfLxccJ3b2Pl8mDmEHm0/NufQ60Ch1zpf0I
fb/EVFuit+ozg9bf3IgshTsVfpi/d7hbUKPF6+o0ReA8YjgIW734q9/mPTlW/BsL
sQVr2NlyWnc697Aes92QiFPa/LXBBd5TawQHR9XsnNKQeAR3fv2FqdGX5fdJKTUY
iiFMFYYC+AzjHtxZJl7bq15Dz5nqwc5B/D5mOOL8/u0YrJHD0uQcc70sVHLuHyC8
mwDrvnsvDMS/W9PQ+0D/8GAQaa93eSBOKTsOWbQ0YShW30pcmJDPGHYJ3ifXlaRY
LD/xZQPpTtmkbxtJPaPsYh+Jg3YC+jE9rEiCM9lIBluVgAzsV+4nx58ZLClYFgvX
X72/YGsV3p5b4qkpwRqZlNpyOfSr3UolN8AJ1cDBzfTpktGylAbaKY26fVaBZUwZ
TYPKSM8ZKLw3edwzmRwGanRQfJ7c1m64pG0oJUv3WoiBR2KdcjgaFbYuT21DEEiF
TtFYawKx/C1Mr2YHNH79t2qQgCn1XiSa9Vpfpffu9RiyTnJ46sWBHybGuefm8N9q
oIqvA7ttuF5vpI0UBWpKdyRJZYlCmUEfw8vdQAmPNy+h8O1X2wnvuOhSj6GXZXrl
FKMNlQVb+Gl5KuDMS8htIE93/1za2jcLagULsZgw9konX+MatFas0l+EqHoSRSRp
Ib1H4sualgtuJQjpXdy3nqiWO72Q9RvB4EbUFzIrHZ58xcR1IVNAn33Fhis1VKWL
JMH7rEKI/Irjr50B7Xz6tFStR8dlxc5KxutdOJ8vafmtS+a94zyFk/sURO9B6Uis
oYnAD60hAAeEpVJBvP0GexSXfAmmyfAbSyIv9P7H+ADoHdcrwlW1C2EfV+qBvuTd
JvodM/mmHknCCQhPrhpP/91UEg6GymYONvO4Wo9uUg8Arm5ILOe72HtlB1p1NMyJ
jFgQJhK/OSclJ1oV3oXeeIwWROeT2QmNvLCBcPsIPlFjqDwT2ADi0KUZFnHP1YPS
6ROciD7++fZ+BydEX+M3KFBj1+S6+Nw3tZyeLpg7svgHu3QVe8v0H/shy5qu79vw
VBYuW5oJnmerxQbsOYn2nE06P+vpqkdQZggLMqeO+nJjFTay7Y0217lBvl7fSZD0
0NDWwgxBUppUEzYuDDYOSlhSZi7cNmFdiMMRxv6p3J2qZgPDngsVEco3p6o7K9+3
RXL7UMZPlDFj5aRKah900DPQ5G+soFfRdR8hGiY4xqJxg22kiuC3ger3ffBFEnxw
YYbdXn4KHAWyUy9id5MU+V6nuSNVcJcxOHLmshiyowmjfK1hvnXwasjhN+UJrfeB
TTVnh3HTt1wp5+Kes8c4w1oiP9pIWdAn/JK86oGq62l16vPhs83qlQMxY71TfuuD
Y7IKbzoXJJXTGlz2DvhPOHK8LmHj2UnxXpVEziZH9ryp9rgpcy8dLAf6n5ZGqXna
Q5YicZE0d5xUiWXQ/UAFn5yikJQUc1qsIKsHMkHICrt8OwqXAdoFyz2HE0Kp9t3n
67cADgjMSlrEfifDUvCULi878uFAe3eYAlqdWC1+rYlmghQZJCIYu6Y3AU3zqdxk
JXTpEGgnDe6tM5RSQe0x/2xJycS9VJkSo0TuTfydhND4De2Ely44GDOhj8SSLDmi
nJaPT82Cs3lVbzKg2tljycZR/hnEEwV1Tb+VwIL3XF+8v0ULIicl48qoKRL/P+qD
dMy6SSMaLekjwqhzLiZbX8TheFarLTcD51akzkIJ9Owt5sgcruZxk+bZpXy++oXC
yD7WBP4LrZlBkG8MnJQYCm7Pmpp9ws08JvRcInZGMyxs0RWBrYCX/ndClrUqJcB2
s9iQlh+FsxP1FChv+PtZgA33P2DtHaGJdZsEjNdveODDKoRK65U2h5VQotqp0+jS
XN0VymehhB626+M3wp/kiIyPyVKmNSRrhq5P3+oegpPyTSrPDSX/BBXqq7WKFp7s
ChsTqAGwslJU4zpXpcaRCoO199KTiBeBgqoR28iyUdyq8z7wBGLt3O1Mw9QBuCLy
UZAh1krQPaVATCFIVovDFnv0meEufsJQ7rKP7JsejINvwRMx8Mli76jEcfPMc7GE
wpAe3LsU4LHEsoNJaKEdx+O4wD4M9DMn2gn8XD2ZTxJLV2GKlEwbCPEzHfx0k0YV
0YB85dK8QbTcfrREf8HNj/oXIRU5+VoIlw4yBVwNaeI1A1TY7cUdqaV1aGT9hckl
abUlTOSRj6G63jBhYLQu72D+U8eGWDDrkIkZvAGJQ8ELQiYrZFYoKYB9/IijtAAA
Z1aS189Q0lv/wJvdBdQKSDjI18DG2gg50TFspNf5UkO6xVUrafyylezE+W2wQ4bc
S7SEsVWtAzBuCNWZr2tqGDjmvhxSoKmGrMYkGOAyp67oD7so8t2/Emlk2SU6IVr7
yY07BxHxqJhIptT3U/bWwxG5ytzpNbdigvgxv9AH+w49jos40jXTGGAOvSd9xa/P
m1cTAwHCgHEPNYr9uZoVCVuCn/V0Cop3xW62if1yVyznBER4H9XUgaNfgSaxP7NU
qIBau2j65/Nsod0HfEfzlybyVJu2WcxdTQUSl9zpATCOyXCU3d9MmwXwyW2JLj0Q
C8jZt9NpAUV/B4WDiHp5Rx23BxiFEo//qpOzxqnnlrt3281z4+hKNSMzgAonyYAF
oyYO8aZnbpD84n66+COaB0OBvIQCwjIjUmSzmXQfcwgZOsrDLkRluif7aDAveTgy
rB2cmC6eC/wiWoYNekbk7f1WG1eehVShHzCh6rrfX1Kz1R6IqkFffuyzLxNff+lv
JcheB14BJmf7lSRNgmkDfsuslySq3gTKJkE8y1fEeHz5DqW5A0z+humsypwgf3aM
Q1NH4IihT0qXsEY7kI2BVumLFzmKZWgZdxo8d3A+nOeVFEa/ogdqRMnlDVehdLVo
vo91Thf1+FOSNzPEp/YWNaiFtq6HPm/736XedJqIkRcEOddL9vEVvGtHF5RmrIix
zJ3BCT3rF6i7+sjJL5qNhIi7qzApDuizAf8pAkuOhYzZW8z+atMEv2Ve9zupx+Z6
Ej2GhCg8qOweasEEEKfH86/bw4Xw5vpatdr3vGr65lpybxiLsM71Et4QC1GwWR5D
GGJfO0i+y7EliGpRBzgLuZUIMqXLQy/mQRXhvnli2dMrf93OoA2jx8QWxFD9Wrid
rL0lKXsBhQSuo1sNDT+cHlpUEyqltnYdHmFV0Nv3FSO6juU5KBtfcnMM9ZzCevJI
sr8jae8ph6WX3buo4lzibF3Fxo9aySxryTAHtGtC0VdF+C7MIYAa8Z4+csuOxQlm
dHMnd/9LSMdvwZvBJzB26T0QVtVcja4Duflq8IIm0EnQK7ySp+ltKdKvc402A2xm
Q+dLVFvlYYB6In7OI+GYMUrzI7ZhKX0dZbSmGWyKihM=
`protect END_PROTECTED
