`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zuj3OkUUjDBrqSjtEc5zCf+bmWmwq6RSFjge2Ub1ceCwewafOksuiOPNP9gf2b1P
LQm4uGB6oCMFyQS0cfKnDQDc3ju5adtl9kYRTmwsOAb9kMLprXQGgrnypdpqbESb
XWVtIRU4LnEd0mmfVnZR7fuOw3vDU4P1lF14g4Hnj3weU/GUBsTU9t5fiudog0No
MWcpSBP7tHE2NK4Hn0iMVTZv9kD7LPAR8Z9UEKrHPykegrUwfq023GFfx6f92kXY
j2xZmhgq5oC2Ru71wDWr5qQP/bAsjNEVO/HQR32mbCA3l6EHLNZrYB3Ya1heMpIR
XsOp3H0rdHg/Fju7dvmwq/MGG8IYJaXAumCAURTEul9gUIh72HPyTA5kC/Me7TXA
tiqJu4oLydDJacQol7yTGb2MUPYok86pC0z2TGnCfbiX/YByoTG48ESP8UVtJw5i
oYK/WDJtZFAnGf4oJuIocJQWMB9lylpZaHGwGIN+aB7A6SvX1vhziJHImKhu2Eon
70s03rWRFphvvkQZB03Wl87NSNJ7+5FBd7ve21LZYvcjv+3KM5qqYm3BFlL7X6ak
W6OTm96KeLx03DUMBi9YnICm3loxQrECGoSQ2oZIVVCsUiWVCq0AV0BBWmUmtf6f
lk8GCxfqSehXL4r9FxLIrcijvGWpMdWJeuIoXYRWcHr1J5r6S1d/GE/ghRQ/hbfY
Juy6fSsbWDQBxQD9xJpDqc4GZriWVWTc1pFE7RwekTlCCKIidkvjdEXTt0MFA8l1
vEAFu8qLkMedAwde24EpSGcUiCR4Pu8Z5J2J9eDiOaGMThZbLOZcL0ESX3jOopZe
/JDNYgGzddcJekUqDB/zPZD2Px7RrK7Jhej6dYnMFYDRC6wdQfqN1pLvVuzqpiNd
sRMMpN3jvjokxxz9JDGA2Gz4dNQOEpSWskfagSUMGr292+xgILzLTN7eCkBToYVO
IfAKrO77W1CoZgtmtvqLYjZhapOp6DfUpbcO2OV8Sw/YRwjrVbxVTRcNUW9rw56W
9Fu+HFm0P5llpIJ6T/kxe9u471psb5kTtaV92c/PgWK+5bGsqO9X+sbiMCD9D3JP
eXkGqiMxodov7uo/aC+on+4TivLTMtkJ2HeD1wwCI/OHtQgW+a/NpHjTqTap85YP
YgbURshJSOXUbGjp2X3gKUBKsJEX6ctKxq3AI9aXKbwwSy2AreW142SgzAIX8p/7
70N0ANdTbA8LXkZLMPiNjleGrrWnbI3oOwSQBiHTdzIlJdQkcW0pRmnX6FU+W03j
nFzzfeFqdfCUSZlxHRMmdSIzAsNDxTDV0tkPLHt9fpTKVMoltukC8TGDcNxet/Kf
6xaArRyMl8dRneOM31epaITNp8ILN3hnaMpmjoYBqxIHsdOObsFKcwusBkFmRHIz
9aFV5bDRg43pi5V+N1ayuvvqskYzlHHL+dE5fQkWLRzPsXuXdWqmMgYSVq/DHawF
V99EjNTrDlaap/yhH2z8v9K814CYpx9DESURpedS0VV+/KRCQpRArAkk72ba/ZQD
POvuFi5IdC4Scz80lVKauSvga6T2Y+xnq3aPFeR0h/jQDC1aludkfJkG9Q0fQWbR
0nkMDknmkBv//PuEXhJL6PFMNT1Fx1NhvOoke4IPBUebOtnqAT69B7Pj831EyZl7
zM9krtGrsFMz+2aLzqqJuZw7R+u0lGmK0dE02l1KPkrbdpMtv+/FjO3CLjGqyTzn
/eL68ianCwYbHxWQDh6vNiDMte0pyESF1oCGESPR1El0E7cMynM1DjhaEX5VTDa1
CjAEHUQ6i54WtciQFRVbvc5vU8HHhixz/WuahKXzzr34IWxq9aebhHIa5DwGdueD
fnfj0H1HdOjZ34Y0N+AgsPi91LJBYACMmP+Dc23QgQ/MNmJSwCsuoz/wyDb23z0F
TfVUA2DjKHe3SBzyZ3eprat3PZUq9cprY/9VB0FyE5W+UkbS/4PkgwpfKydHmIaG
3v/PtnyuPcsutlQgwGsqCDvoVwMcCUbX5CIoZod9PYi54N01UB2TzwSUXc/5CNaT
3gczyaNIQ0LscvQ7NntUO940hH1ea0OnCgtRXx5syAuxtY/Q9jkQwlVVZYB5li/D
f70ZQqHjNovxi69rHLOMwNZZMExkg5L0zVvEWu4KIMZJRTC51rAZmD5k6isQ1MbN
xRsdmcfKtiygb/IKHAU3ndO1kikWNvZXq8VNDmXlYqzN5OppQdgM4F1VaaiBWaOX
XhJ7qxvstdAf62DpPwMqtkKvnE4pmIyP7fch42db6Gbj7pERxKek8ylwywjNWGec
7eK7sfHAPX+DpuZhOEWeubqPwmufDFR9h6KRptT3Db5lxFaALotD7H+lsx+2459o
hYfONLzY6HsebhfPeJ+STt72k0HSLSDPdWWp/3yTx9ILBitNPZKPQBPgfWgxoAg0
P/dQ8htClBqvRYFiijcArXPbqgyv9VuP9A0UBxuMbBCEZmzreBzyStcr/59bTwos
epANKw56knXDhtaTEgCiWG7xWFstrx74wM9otC9TdRkIAxElLVmeDkbr9bDPc2XN
Tb4xlxyEGlm0jaCZ/TXeXqKpDRKXx3QmzV/N/i4ml+aHYoWPWct3YvBFO4DC/1eG
YoXAsGMGbUERhtjH3DU6YACYvYVJHCYIFDgmHVCfZMQJxVC/St4/7B+9yrovFjjt
zC2u9kd6dse2A6Me1uMiLN+H29dXUEeETw7Mlpm0wcTmEV+7a0XxIsDuFGinPiCG
wgfvAqd6KrOEHFxfaXceswlZlPhru5DJ3HNVhP6BIQgk/QJwDkiz12ejR0ShekJM
1VcOvBl68saZHlU1IcLBHvohlRUIEk7gbH8blxIqskA=
`protect END_PROTECTED
