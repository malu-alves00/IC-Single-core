`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VCKiBGMacS96aiwghmIErcp0hU5rOBARg85XahdlGQUepZvH8l6YRo+zhVKCyeab
I0M+COmnzhX7fbVKyDox0rUG7X6/oLMQfdsQ63QWAbaKEVWC4Wp/qmjh1x9chCTS
pcW0dnedhw5dL27Dh3CTmGyE2j1ojzkhavQkps3cZtRdcxZnfIQWoWAPrVLIlKnl
RH3TSYmjD5PtRDSFP1R4uU13kZmspeyos96GbEhn8RyEAzArrl2TZ+NGkbbYKSnA
FUE1P/duGP8nMQOBo2nuLt5NC87SBr45W75KVdkr9r11aUoEmPOeAtPyejbb92az
I2gpwkG4ImwJd+UvuaiTRyc3nMkxw9vCrlm/kWqKs405vdCCSM0loNe7NFpMWhfF
VimfpAV89M+zdgUhQKFUMOj/+h1Vk7LoPf65jCRKnqG01mOsQWAXZlHD8VxhRhz7
VjKlXn74sEHYxkvbd8azJB4jSUQgSCAnsEVOlm9tDTt5r0PiMrmqlh5XH3jOTHdf
gwung4LXZa8F9RkfJDlFL7Nm3/Znk48vkWNV6PJQpGWdXRqCjQ3h8cp9y4Cb6rmg
yCLKveUboc36b8egq9uo4xLKFotnx/2GHU429fyMH47KNxLvcc7k0TgeHD+K3CbO
BbWXEh1i2tF3SRdq/qKwVryflT6uteBfCw3y3m2GOD9WMJv2gtyOdktYYyM2Ay8r
aWVed5sRovuw0t4wwbSg9AnbF4UHURrU2krpN3V+l0KEVW5cgIBo5+ew8iNoeUL9
CW+LpSH5rVAOQpMYIExvL76PzLStRf7mJsKhJtSYk7psGPAEHGXjPnYDSZejN7tI
vH1a4gIEgO039zM960QzBxGnft95ebuPbm4I/xF83pmpBiVWixfuL6hxJH3REbwk
gT41J2OwnSlMrGaED5zKuJdeX/W3BzpC687bhN80pVf7OjrIrEVo34K1f/sec2OM
jmGI/bqen+DyrN3jRc8HlAt3SKNdBeg7ysuPcwg0dYSgHazdN5IwTa58nTNPQuVj
536ajSTNBfWkg4GNA1wXzoWqRb1JaBXka/EZ0X0ABAYudon4uaeiqKI06dv1DT2O
pEMFWZCrGgRmU20DYX9FvwKcPUxi8e6mNDMe2LYIAlYPEi7OS1ceSKLuY7mLa8d2
yWJISEE2/rqqcvcAEmVS7uN/SxGikuPwe7sTV8/MofK3UI1dcGWLWYRcEW1/EUZb
HebDceAfcmkTfrBIWQ5AV4+EQWtqrmnut+joQWCbft/UMcfs4Bf7mIHe3jNR980G
/K/emNLgH/DWoB6y4sS+otQGRpo2iH1XiZY0XTYjH6b9csiMAFknJfkNac3BilAM
VU4X4vSJ8Eo5+x3Tr4E3uzfCbtiDwJCg1CkWVasut0vC094OkL96XART9tZboQXO
hVjJYCZmAurV2+tu58fcXMU6bhvvWIXJGR4QPNJyJxKyi3Z2hOKizVMWsKR19brd
VkIM5TqjPQd2MXNzRNfIuSKLwcPpJzWbM/R5LxwGkL3TnpGX3BvDRpej3gOXoRzi
ISO8D2iHHATXwCORKqHbiuVeK25ZB4h3OH5buqRLVDu0kPwvWmpJTKL5wOpa6kIs
`protect END_PROTECTED
