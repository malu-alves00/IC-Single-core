`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eZUWIZNYoiYhp3Br5cSu7Oj0509tB6B0KjeVaECJrWK1aSVSEDj7o99bH/LKDXF9
olJ+iRD+mHDRIXIMkMNHrVlmEPtv/eyQf1HfsWhW1neKsufYpHQfLC3d+IRvOwpu
41+XCM458duLIC06Wa60dS6eXUGQwlDxZ0O6crdhUCeeWq5MdtYpDcPofvnrEWdB
LKlnhYG2lPzokI/kYW1h8wjORzdykdnBgTChpUaxGW7NLDXsgnGIwjL3VanRZCVW
Y+Tk7lK1dp38l+IXA5hkZuJGx2lFDPWETRZZVz/ql7Ac7A2qKigPwHqkdzpICvxX
cmyhWfiwE7yDKPSrXcK8Nghzoo3DDzBHWGKaZV05uKwqYqcF2bzHw2z7gP/HNmyQ
Y5ezqFmjXPoxb7F3DzL2I/BcRQQEQjILHy6hcp2FiCCeIzZ9LqCXfKqrpkzdXk1G
hRMLVYArBoQPyU+dIGu5UTwF5CrZPnFiM8fcqx8Y5i1gUqEJ/0qGMQew4VpnYHyg
3uM+TjJziOz48+QYy1PlyGEhQZDzPy1UlnxM1+dCk+rGN3b0cmAkgD9Xv2O0Glr5
djnKxBOsX+LdcT64jk5qpq7MzydXUdKuOe5DvU/VcFumzr83Jj+P0MU/3Hc27hbF
jtXtNyNHN7xW4uhasvKq4nil49AJs5baEZcU+aDw2wVmIgD1hBlmkuQ6OhskXngU
EkIIgBwX9pFtSCoikv8HyrPX1x5iZKkGjJnM0bMgSJlHfiiEsjTlcwG9w5rHaUBW
/Saw/A9nQxNF6KTSGNshmbmn0D/bljRYCRECicpr5/8=
`protect END_PROTECTED
