`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2TAoRZHNuf1b3+cNNdQzsz0LU4kAKtXwIcfrnqbIiPCAMlUwy9TihhMkngO2yirg
3EFnteFnzr1f2Y5V5f7p1PFX9CIJBPvRndxchwoutLV2iXefxZUJs8SgM3LLM3vp
G32jNTBUr604Bwx6tBepw/EOufBp81HMHv5wo2fqJkWYVnSFW3SJVJ8gMvKTC0At
LIx5jK+BZbQVRoLFl0UCI/lnkHfYtj8m4RBBhlOM5uYq83CSR9zsKtQNu+6lPiRT
UehiiQsuIhUVB8qdPhjcvvTzt2h9RY/hrxw+rOmwd5mnV/TrTUybYjeNbL8ffu69
y9WYJd8f0cW3+qH4n4YLf1XSLzZMZkRl+kMWl3hj5QHZyH6H058MnQ3TEOG8rGJH
XZYz4oMTGudOOJn693QxNuXnBXtrtj3U5lu4AEQ69sgRQlcHVsrwWV6hHPxf3Gsm
GM876FGVWMmtAUn1pU+1eQzZiYuYRpACetugHXzxt1mLB8tAD0AdFA+dPWSC+iPX
PNSLAwsSMS+MUgcTg33UKY8ldi+7x9DzK+klegpPb+JnpyeFkPsVrD6BQaAJFdel
7UpacwnJChjnLOztpzFAY3mUJMjFCwju5+4vu+g0rfpv/JU4Piu/kRTzIv3HdD80
ECFwmcyT+CHHnc7kYZN/GS3lFLtFxZGCvsz1sy1BP/oIWUd1p/s5SQQVDI3ngtWr
1+EWR2AgvltZaR/UrCrdgoSIPu560pkoXTE31BLYpRSZpMKdGCFTTr96zt21X5iZ
R+RRUZEzy5LJ1vGWcwfUClNAI1DROQlRase+TJlJzgz2jFm0EAfSc5wiK1wpfSAR
/MI8SKGuJf1QgtcfVHtZfhfCN+8AEIbypHaNH71JTOE8hi4St5BVMkI4Lc6CkIWo
P3x6RcUJ1LNPqJqUhBEpfUBtDp0KwMB1KqOQimdcQlp3P1b3bI3EFMj6Po2rnSOa
O8YHjUNDA6+SOqIjZvrcfK8EKf83rgsDvvUs7+VKWXtUd069l1rqE6XNaL6kLnu2
1TcT1ErjpDprNjBn2I2y+l9dC4ui/7t+UQ8QNeWJZmx1AY3MhVNRoOLv4S3aT21K
Y/u8uRE/hQKWSNXoF2+j7An9qmMJ2DWcj9eDuhGp6d4R50gVoNR3ErdIKOkhEcvE
mY1ZKvYBDfMW4gKcZNt5JajfAbdQ58DsnEcaAdYH2NTAL0YZj/weNtU8cqB9Z4nP
EqKrfVpfcz0E6mV78ypnaZXWaUPcGQgGGPysLcWJaartopwoAFO8NGyMYkN24zhG
WmceKkpaonNTSc8IjNRrfr3/tPVQtXAKpWD9eIkSxMKYtl7JtSBnQHw1wqxhTG+K
c89J2yPzSvqizPQP1N5yjDnRy1AFL6Ue8QrLBXyyKxrIHDsfLHNvu0gQNa3K4Gsw
K6nWAOD/xmbe5QBMetQBQdsNrM63gSrmmIkkFrW61Yq2ZJuNH1vLFlUs6GIueR2t
uy/qv0vDy5feummdZcUEwfdPn8AEttSU2juCpvlbbv7IMpi4+CYsV15R+lxLFuuy
gnn5cyaPI6LVxys5/AfXRqx4ED7t+TPdEKJu1XtFwnaxSYS/mq+Y68QXjHRRpLWf
Y/szOjryXe3WXeSYZEKJEKfIT+jwRLCPc1biV5YxcdyJ/XxJbahnFT1MRT7brPgP
rQxSYPPD/YI8wgKfz8eZOVSEGhizO7+JCoqMHS8huclhuqOnW05FNYAz605SnCmi
nedqleMg2pHye6chQ7lLJDzQ+OFSflr+1IedJeg6vSfOB386I7BpgWVkIghX/kKu
4Skh2wPn/uKp1zMcPbKbazYW1fkR9BHWiavQSnHtrthV3JSfUz1wqQfX2z8TS033
hM92KrW5S2ZtodTKOOACxpkYTBb9Zb4Sg6BPYECL1SvxZIO1g4oIlr1KdG7fAftA
`protect END_PROTECTED
