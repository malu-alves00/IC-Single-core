`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DC9yXf5rUsE8nX71HgiMuRxhcuFGrOsYltVFOvk13DYNG3ll4CS8od7bIVz693nw
I6QgzuIma7EkmsIMdvozQug2Ehn/88sFRO3/oxCQK8vwKmn+nF86+sc637vFzAHg
T4Z3HzEpTuKhp/SutoWmY9Q7jDyJ/xgXjn18dInPTBwVnrb3U7gPRjBq65RNMd7F
blzYdqhsMvSCW40mF1GDPtmp+eRFmh8wPbyzDUkl8a1Wu8GCof9PiGWokzoVYGky
+4yvyUTghE02h1hoZcAe4Rtmq65Cs7GLb/z+XRpktsTqfrxkpz/sL9wyq6Q4zZhh
1rqwixcik5B3mV5dBbQ+je0fXGhn4J9UHp2uzeerc1wkftAQvIWE/eCXYPMUhAKh
A0xwMf7dRpIs9sgivN+F+U1ImeaO8uF3DDpsBjcqWMgdga4i33r83dFCu74LwcXu
eNkzM2Ml1BxCodvjDMYaQ3/xvx0vWFPKTC71enUqIrvoaSBgV2zWLKtcxdU1pmVE
AXV+fflIHokwgPPiLpczW+H5HCtX5BGit/iaVR0J3E3lGtqHN3NP4UC3GzB2GwzR
Fp+YgoIoIcjP3Mo2qmpYjC5ZgqKQg78P56Dha6zvnPr53OxajBMgBYL3sRj////Y
qUUOaZpFhvwSbuZzWWKiOLTrdpqNhz+uDWUBGLAVRqMy+mtUebUA0eN9qEsvZuzK
Gfn7pqejAI5SpVlCVAdxvKbm4yMdMxLEnpognOdSHE47B/MEKr5nqC4VYH19tprO
EKPkQLRzJAglzWMjGotOg33y1GkBeeKEdD8tTRsgtPZo+76Sdd0yq8qR5mcIQ+6U
JH+o4fT9x5Z5jhrg5AKHOl130IHtItJm41c9VPc9zkv/FacFwN62xtBkXA1LARjQ
4ubvYGdXaSnNF8Cf8FvMFCTaMc3FHPUZMeKbHvj2ErweGEao+UMzwDrnC5q3+17b
Zm4fe9p/60vgMWyPB0m5HerW7M0PQ3AWEVv/6AYwQv41lN7X9vWAOPLPKde6l8fS
CsfN5LTFNubbmHZQTPtT8QmaO422DQb8eAoDWJYssGsSRNSmq9zXMnNiRNsfIRPF
0IiqLjiStbUpRbyyW4arWgUXbeeTnR9Da0oxje6VVeNv8z32V511lOFcQG4CtiQC
+33sGUWxbzVYSmzfOs53d2p1npto6oWh3nOol8OSv4LqZohiKHviibTV9Ae6WCHH
oYRk9wetk3kMff05N9DcCtznq8fQ6B3uLlcDMI9ROqAi/JvJ+o6GjyETmo0nB6ot
8GizRDIEAMnxzfl7WD7XtZwG6LxULjmbeFPIiIjjES+rJy1k1GiYW1+7IaoSKrid
3G/AJ83vmevv3jx4owTbW2mqYl3UTMiCcp70k2UbkyhZ6FdFBhv9142e/M0NRlfC
ubsRC4/k9CnpH5iGWzAzzjn9is+AM4zUIhrM/+iTjltG6lXP/GqUgm24QgBkbpTH
BCX9oSbTqLlVaDRDS5TKC2+GolLO6GtiOkO+DUYffUG2xtFcG6Lr4ZNFch4AtIFK
DqafWNPvX0rNhZF4r9koDmSrH98SFRF1F7lpnBOAhm7xTXiLm47XUkasbecy/TL1
ef2B0xDE7FQE5F0Nj/Dg6hASa8MdfXwgBSAUk+lgPMx1qBb7u9wVdqjXAP5XlWRO
8QCcadXCdYYuG72RdEnsFuxdL0usO50DFAbUa7EGXCcZ8Y9E54yw7y+yT98FKObe
u3JVaKQaEpEyE59hjCyQUZCHhcC+mg+DEN0I5LCaNjLxAgooxdN03v2R8+h/c6Wr
EmnHZIhCk1cd2wRFDS1B38OqRKNg6QS6prFg9rPWYNL0H1JmHrCjLQxTyK9TwwSX
b46t7KSrKW73PjywuXVt6SVUwpU7XOFwfaxNn2a5GCGNEkr29x/rqCrBIjeZb0IH
ePqGHMSU/mdGFKyKHKz7qCS6xzKlPqdygDD0cC9wzlkZjWb207bfp72lXwwZiZqw
eAneu2I2vdiZMwUidJADSaT+/cnvESRYX9BDzz/U9W61lCK3CAE5ZW8renhVgbqV
DxO3qjW0LlLDcOdH2JnUqv1sNJhxEFlh/ex4XyJD9/jowlEVQH5QVPhUosG/G7vL
rirLZAO5qpyaHqHwOyLYg4gs5KkIOYSQKsw8p6JJeoNVmTpqSHpv53Xjj4CUno61
eBurcISXLV5cmQdZaGiQvuvvXlaanPB33j5SNzxsMz9ox7/eTMDEkHEAYWKS5CIx
i0uEbTMdzRu+kKKe1uqaur9a1rIGH93Ibl8k4q0F9TJULXE7Ver2oF4KHP8d7vNF
mSM1r5A9pqOpLiqGCXhh9+QLZzmWetZzteLYP/UYgiBqhUDmMDinNkOFwaHBV73e
eW2kYbbc3vKAOUeUWFwcRwpQsAIgxXJlKio3FA8nFBWea0iSM2W0mUK5pbWOmsPI
Vm1C0A5mHU8ymffLwZca1/x2hQi8NUI9LXcUkgOpZzcZBuHIA9PqbpUETZ8E8q+E
0OD+9W/w1uS2a/oQ71STAxlssiBsR1VlpXWbnesPimSUNiTHH9SvX/q1lt5pNNBx
ntuM3QofAX6a07ScbsnIpA4CE+r6/li+yNRfKJKoxFOkfcacSIl3k/Bdc7WXXCVy
KsFX1IKYCP6k32dh3CfPjsW9hEndouzKBqrRJsPo2c6u88roz35InTiCrReoEIV2
8N/+F/xh8wViFVU6u9enrNggUXAjmwSUqJpGYqJrW0gHTCT2HHU0K9AfWNd3ER+N
kZKvvO4IlKe7oHIo8KyxjXqjhRWzEJobqM/uJ68Jd/RShy7QPhXeb7i7c3HuIYIi
A0+v0ga/pK8k6KqdHFUnVl9UvOVjxLVaZ/JS6l7m6jbJVtQ7iRGZaZY0iZ6Iczxr
UQWO455alJYrnTveSVBwZvruGv5Wo5twIKJjOjXIZ4qwMNkC9qYCmNMxurdn2tV7
Crv07F80SlR9d1lx7/3KLiLIwCK4KsrG+z+jf+wo+FrbPC6BvfB23P6ikM2BN5CE
9fXMh+qLNTIqImGZ/2503QEQdCSmZKHIkg+/8KezSgxKOdWTkh4PCfpSraK0s30W
/buI0UscH4vSV18Jk0pw2JEIewI9VuCrViGNP7AWeSeKAHAdOuHyx29JhXm8psZa
6vNVcTRbNMEV6Fn4c8WCIPgFkwcod48pz1PdQ3jSK/jMcJNbobWo037AebWHRqrf
oOx/TD/N4qSHFsU3eXy2SfsGm2cPu+L/oEDCWJ08FDfqQn4Vx5F76a3je4XTAHcO
W2z7cxTorBibcgOkx31Mx4dWhVbDbRINK0tRqck2xJdcq4ZFYgXVAiaIW+eHpMW8
QDKHNqq1FwWAZmTgUpT56QN4zcOTCDsDjGaxE8eGVSxFlSbHKhCrcmDwaGG0ZCvB
hdqlz776Yo8Au1v6OdbRTQxH5OvadRH9tTC/eb6qZqL9WSLn3qnYlRbvExqVeH2w
JhUFYpu0d1P725JP+CHslK7a5HSqn4kDiK4EBjD2uurvZBbn3w2697ClU2iVc02n
IzhcsEm/D8hRZ1ZFUc1RmFZ3x1crjLe3tqOEOCKDHo+gZu5yuOPqzvpAYCo/HO8t
BSKyjaJ/BfUV22AcfQmSlj77z+UCDAYwVWXfjHDyjltXWdFyGPQeq1+MrgGIgX5i
JNZcR7f37j8MH/bFWEQFyrRVOaCQKTgLg6ivh1qpUo02I72FLNyMssLFZrxh1lRo
vcSG+x5Tf236rbrOF9Nv1JF0O7fn5/SjXphIGVa+Gu/98ISZDLOXR4WJG1U31VUX
ObQh5lSylfFJPuKv5T0ZfsF0H7OjgITxF1qpxfgclIM7ebW/2pTz1bziByWSyzkK
QxaC0V2r2cGf/tw9oAZGktUitrxQ60qqV4Pz+6vAkeGEj53GN9copVMsQUlXAct+
JBBsumXSQIsy8ebSjSMm5iMsvKNB1Ap2/J80jUcpo8uavnExFrGfYQ2Juu4EQfpG
l8p7Dz16iUEBx0+9lSfmCnydbSjZ6KF0xHpddpt/ZpcIhDQgcNOwXB8LzZDQKDSS
TvwH66yZ6cgzpC52t4H5ljHcs2ZiggCsHbDScX7J4TbtSLsSkO3WsdbjMKdZwRsY
G3iHhhuLNZLV/PHhqz58lbKAO+3yhp0f2PIis/M9g5jhrDwO25oMgeTBHUy7S0er
r6OFFraRArqLX8kR2FD3hzItbM5v4pYUZN9L9Zrgopb1E31jjCPh7SXPC4ztr9gp
Nk9rriaWGr2sHC8Ng6QQUZN+gJ0XL3p8FBPFZxDbp98YZTOUmD6sGyEGNrUZ20Sd
po004cOYMKmqR5mVUi5EkwkH4hqTecOrTcxL1rcGjVEQB48sGBReol9d9SIk8vSr
MYd5RpfCWTTHYIbH44vZzc8Wdcjb0lRshUfJrrynXX+/dE7EPtIB34uuepL7CWNv
vyGkgqaK2UsiC6YyKnO4kjOeM0MW6W+N7b/NR+Eoi4WN+o7pCessm08OaD/mDYh/
pKpx/CyXwkgNpNvtx8qmjSFOD3mvpjH7xZ6gn3+hXNVXog2F7wLOHJUuqSHDBp0i
25jAQDB9WKv+Hp8kTug+BC5BYHAYHJwbO/CKw9xzOMPwYxJ0O4//dCWxLJhsF67b
450TqakGK2xwBSRnpNSBE9k/Ulr9NSYZ/ZV5MOUw8ml5BP0Bpo4FiASU7AJWTwk5
VT/pkcBIn4Xt6vlOiEPNAsVLZeQAIn2wYB7ktbOvZbGhmexa36ZkiBNPod7aGfIX
Z3kEApfzSjTrj6LlOtDcG1S8KNTrzoQ6oloF3ROg+xo7LtI8xAJX7+vCcu9lKDoj
YeV8bN3gN3FiQwxgfI6xIpV3EcFS+LYkBwQ+711xCVwtMRJA2bnMw6xTYSc85qYc
u6JE8+yrL+GuzA4sqlJeOMNX39KZnUoLko/GggEGRHlJxCScMP+HcEp1D13yxLoG
ccJ44EwyM5IU8hauEvZapIdEZbfpJtkRidm7sBFE1EZ4liAFpK4td5KQ7xdiq6YR
P3oeU3of6ymTttlgh8g0sUowWria+yeInm9d5r0udME/hlmtLou3myQ8ZWMeRgW+
Dykr9rtDG365DOW3k3fnSphga7vMK023PfZdhOSRDYuopzDIP3boT/XGg7IhWqC3
+baE3+qmMdO+AnUJNKfGdn8wb5y1ZI1pf0+LJnImAUTmbR16m8sSWZdSDttmg9m7
aW2aPv6CVN07KBRVRwiP8tw3pX11dy7agX8LQX+XAbtBqpWN+nrv+2W2TGZVXZip
Bddrlz5Ubjfh58lvOSFBD1NoI4hMbbxHl/f3aBnX5ZWwn89MY9GZJQqlv5vvK1Hc
cO1/o4Ch0CXbAep9cQiUMDqEUzRDpxVhm2YXqt7X74NGwGpsi5mpBBUxvdCezMne
yNCzt8WALXU294RHE1efjpn/iINMzT2fm+TvFYEWyl6vqTVt3S7U+B7YnhU27k0M
KAtYqaDTV7bgvY7zzRAWiQSXzcVIDlG+1XIbtMrHIkzmy7ZKmxuIOfZpQyyBEQ79
TyqtNiwwLSlHlHnWKnIaT1hZwvPkWE88aX8cJIBhSr2miWhGhnrR84Gy5Zhc778U
uBUt0pGxTiwM3mJmFSM35o5BCRiYYjhr1eEP05B0Uav8JK8gcZ1LARrRG5PUEjQq
9Xcykde089VssvQxtWeRecocVZPZrtp9N/vtKyf1/CglTpV+i9z84VXnd4IaKSK8
B3I46YsNsdFjqPHxuEyVVUIt+R5tAyfZdeU2pxDsKdfbYy1Ppmj0GGD/lka3dogk
k+Q+c9ciUihawbzS5YUjXpCKaDRJeJjzWKdocgKdbR6Dpc81X2W7JTBC2DpuWzdB
dyA/hnrgWd+pXDVwIifUDQsBFaYc9/OY6Gb7NeiqdVmORdJkrTcKGcr+YG6nyW1t
`protect END_PROTECTED
