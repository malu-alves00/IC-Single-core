`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yHfP4rLhv4F3cKc2WAeTLJEmp3E1B+onx1Kz5geuQp08PhdJ0VxlPIMCasQubUGS
8GzHQM0nZTvC45o9igztr8pc2cBpRr2k7TDnQJOugvGxaB5Ft+KkDDO8CPg0zZc3
6bFW2MfQDaArlCL02bp2pbWvpaR+aZTyyo1DQycKixDkpPW9qSOnE89pKx+w8AA9
/NPGNdnauBbeI9rvcNAprV/9fH9OXCwONnE+CW33X23mTPaukVqp5B10Y1lmqoN3
gODlgp7Q/iWsU3l+QP3zRpzt0grJ6JCGDEXi5gOdPAJenNJpjLn3qqHRhcOm1ntk
951npv4qg6s/xDoHeNAS4AK44ZCO91Vjw8aiZH2uFKPyzJtjQ6dYlR53Vo2hKlX2
bJfPY+2SqPtlKZl/CrKxMSZxfnPsZWubDGXO573iQEVJt3gvIIpTEEUl0g65ax5l
jmTD3R0yxGnHtIIbGKIyqo7vZfLd+5Omho1FWLLyfJRNw8piHOLVVqn88Ly1CyAO
XUieccShOVU2H8fmRNA00FUcHjSOrPgn1XBFlFEsHIb3SdZbxr6rXbhytAHRBGGg
wVSEC2UrVI49ya15GSzbi/W8msbzaKE2+hZzw7qd8OfTk5mNhkvs9IUtuCVHQ0l4
JDh09GXyq1eVnQG1RB5dmqOJdSc95vidi2KkG15OtNg07eyh2IvDgrpx7wCWk4o2
rMioKgGtGhUOQAiibJGWYkl5YuwgHJflQSSaAKN319e0dcnHZPyJ004NavJgrIhH
2QCrv6jvXT9HquJyHXmS4WQ7T7KyVLdHz5GV8OD1JD/vzDr3vRd4BPn00nhWc+hl
HEcQMknM25OZLmnrluOaX7GBtpxprtHPHPmmOyU7jpqOlyCL86jVC1gbbHtH8Mcq
+xgvOlAlCTRLOtjOXJhcPWjVSKyvtwWmBuqzC7fdiDlyFurv+Chc8ox5KI0qQxrk
qWtdoJhTEsh/zxz/lVD0rAtawTTQvyA1H+SNZVcQ8udzm/fAEr6EXNhRn5plki9D
pX0YdAJe/E0f/tySFy3Sp6kxTYNpSSgAmu0OA6ET1g+/Cf/cXOtLGNJZ0C9cUfJV
8BS82j6a0fLBpZ7yzcrApRPVs4UVhzRBGGCg5Rg+X94BU9KMpz0Sz5vcnpNGw2D4
jQCBcSUnInfwNM8RWOyksU9HD/x5Xn7Sp/GyXPJOlkVbaIa/M0A9zZjdCsW609Oy
qHDfnr0x45KAK7mr2RV/gRH0+sUBWCH2uqQ6uJhSdCFVIq7e5Vx1SOh0u1WUs05V
EPD2MPjMg1EzmWe8fiEBHBrxJ3IIdB0D8Ga/QtmLKhkeWXeMdlR5hHW3hW9yGpzq
cAf3UcMrKvQ4EnRU4RcfJmzXcs70ySQYlHI5Tre4IM2eYMh+USmfP9aeUfdVwAyQ
J26LUR/BRjIMKdkVWPtiGwtqUoVR0Sf625ehUKf6LzAWwP9tT53/YumZJkE3D3DM
g/nEbjj3bNpe4ZQ7uZ+ULFG+ekzrFX3SC9BhDCjGuYwmLqeT0bQyfO/FA2lIx61K
n4u0QfWUR8XuNpj5uTIJBqHA66WeLeeKqnlAmD9leBX//3VNYkd3ltO5PONE6cPK
3fq6PmASZlkpAhqW73En64eva37Tl7sXf+AGLc3Iy3GC2dqj6SVyppbLtt4sWwdI
fD1cItyRA8tSDbk7AmJDsU7fTTYMDSh13TyEu1a42yL/BT51yXcphvuMWeBdYhQI
3BtAJU233Xnzpx2INK60cOpxzfBf7s+zPlzsDj1aBGZl/mVLGftYEhl9oR+9xb4q
k03wKo2BdNN5IzM2bhZy2NfIfw3Gmob3n5ML0g4W+WggbZNLzwPJd9mcspbkeHLU
C7s+GAaIli7y6cpFOm+4JsExUEDrxaUCrlb5SIB/BuFRbBeN2D8BO//cPTg0o+xd
+H5NKXo80fqAIWYblMfgWqr8eqK6JBHQcYYXRNK0BEi6W0mjL6mqK3Nq20xqW8tI
k84svI2daR0QwnbHysQwbdnQyX+k4BD/fs1izUxkRFxCOEuOJG3PNrvBL96b17Rw
5Op+oS/S+bS+olG0WLKDnG9sMnEcRtD2fjbXXewxeBZr8wES3m+3AdhCImSf8csg
kULeMtq7CGmpVKmmvnmL0JPC8d1UISc+y9vr6/QaxwTH8vaw/kdMVU0nv4e7Bzrh
ERBg/RiwZ8Cf3mc5ewSwO7nangsHtDtOhnxsHBt3wxRb/V5GdIYWi8aeFnn2X/Ex
8VivKRwWscWnsgGdOZbVv3SaVcbxy6YjPtPFmTlKHuAaidv3rChiqgJRRYW6B5Mb
M9LLcTBrbqNywpPD7t6k58KnuhMWk1sYC9+o9mT0RPLp+wCZ4WDDj6WedpEoOgUr
Y4G3g4TbKiv9LhE7RZIwjI3bn3qL0Eovra7iXZbmDwjBmXQ7MeLOtcvEzpV9OmMl
SQNZPaFx8hWl+4rbQv/atvhf67926tYIIgnX/iN4ZDznnXNgRiHGJBpMA0WKf1OZ
Oh+nBmO3RUTAaIQ06iO0Kl+4EJL59BsvOeqy6oNNAhIP98MfrbCiQ9NI8JRHCs8a
Ek3xsk+X7Eq/5QMhVG5R46yqZU7OWS4nalTVcVfWwuyl603WiH5Wuus8z85rKawD
6lQv5JrRdJQEo6E+3b6wHLEdtK5G0v7artFwiqJN6lcS+VVxVIoR6g7QakOu5iYS
0phrTasLxH1tqMC+Y/zsx+285J2inVDxQuUxG0hCSwNkvm1izafOGmQzHb7vmoat
5aejypBY+/eVJhG9Lq3nWYF+dRhoRcG952MkeB1/9bNn9BQ4OawjPj1hTJt6CyX6
wPy7BMbYHfa4eiBdkxUMYq53+q71ZQGRaPuaT2sEXc4R7IvAbdNl5+cnxO0nuhCm
y4suh/FEmdorQDNSsd/VVOGwdmXl8J3+IjbXKGR7puXCdsMFAJZuZaAbX3PjDNYl
zch2cz4khYS/U9KMKuoa+lRAIFje0JgQkm9V0mIRyDhkHh5uWNXho8czxgVFF5XO
56iY0YFjzHcAOh7hlXUgwTgcCmBTKylFsCLSpgyErDXBTZ1AUwFohXSyymBYI5j7
Oa6iaoQzW9Q7X+vlTjLw6Lie6j0Uo0LL20ialWA1ygLqfcRfSDA/C1G7uBPgaz+o
QTAmCZHleys5v3uposL4OQWzGVG6kCLRT9Ua8AhcdRMfzU6L6fGAdYOvE2Efz9bb
/RIqL5Ljtc/O2/OP+CzTj39G/kmz10EyuQU1MxymykPtGS40fGXjJ7zOkW3ZY8zF
qDOIlg2svmBXK1jBddvJhrxGcNWw61/++HXY2+hpqED8OWJp19BrvX8O7aFjtNuZ
bFDA7gztgitj+wWyzkQIDDwUvxlr8S4xLrmVAtoLSr2sSb1hmnxnGyjsTYjKUX8I
nwsCbcLoMuLs7dGsSygtOH4e0kDY+iaCUE3pUV6tpeGvZrH238a8llqptIgSZ1TP
Ann4tj/O7VRzWxc1JVRWO6YvXvpjsS7TmaKBv4+qDMXXOz6UUokfn0uiJRuwpTtN
dXnYlaieIDp2opbO5Xzwx54jZEb/sc11gfN13arZ/xwlv4m+bD3THOwA0Pof+2Yj
NGDJftKO10Q3TKMCntKJk1asNL7y+1UVL4aAuU1m51SZ2z8VMrwVyqLo9edmF1wM
xhXxvaEF+/795ZhoG/ASK4rtQFo+REajAxOltviQYcggJUl77Oxn6GwYlvbWHMR9
k0jRoulOAph39kQD8VQU1+dwbV9xxxA4PIunuj5tsO/P7oU1hyXbDwBtkttdIwiS
iyAYJ4Ye3U6v4SEQbN6B0mjK4n1RF/ZykZ5zy9/ljkfr94nA3cMvZb+EXm7KVG82
/GMw8FWMI6SktOpGolWmSZPq37I9UC5AWNasYT5bno3Fi5KbECbyD3iYEGDRTvj5
O9hYXYC6q27igVwXJbDS8xy9xj3ktPvg7pHpjifU6n7a3iRAC7T9bwJnIaH0e6SR
uuuBCku81ParcDuh1orB09vGWSsQ9Owuz7k+PnCAt/2nKWuXlBW7Zw8I/Bt34p4f
U2A8d0txM5T+f7kax14/MFrDJKngQz/FOldf5CbSyGjdVT11mI4TpAn1tn61EmbB
39v1CEDWrYthoNM9lWW3gBoxbfH0S/svuAFgpgl3Z2leGBb5Q5vgJTdlDleQquSJ
UW6wjCqbpxGUB/w56CZFJaeHYf8QdgIh2GEi6Qdf0RBpDN+vPzr/+hN4nid+aWIV
48JpFdn0esLau+kLipAYrsfClfQeXVK4VBG1TAfpdEluoPh1ICN3blk9UKRjXaY2
e4bmMf1eT6rtP/ZcPAxA5/HewgTrdvLTWPdAQXEkDHfsIOFEKXXt88pl5ELI27IR
lRFJ3ihnYnRe81o9H873gwGtDG1Sd3QAavWAcAbpCIs=
`protect END_PROTECTED
