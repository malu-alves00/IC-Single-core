`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ATAqI0bt/PzKZv1tDvdAo5YLid8nwdzSAVfeKXSKdv86YVzC0jib12oCCnbV9ADi
bBqya/YdGSVnmZQ9gCAeDUlryrdGngZNQrMoMiZo/kFrWZljzp+xgr9tm/jjtbyZ
9HtYd/J+1wYf+8UZGbcgAdt1rPBr9gGrHNiRUe5M6YMeAU0N/iAHYTO7Jz4NLM9d
Y2Op4YZlBB0orX/TPd7oSjCR/6JkLK8P1hbjPhuG0VDpxfjra/PHGDqp6paYTWKw
1QUggWrhFMMh1OOKHn7Kwjj8JQXDXc16T5Fdks2pgV7f6i9rz2kjIc0pj2JLau9C
YVLOn+Y1q0Hxlews2uZtWxy3TyiX3uja9MKabhVDUfHhWFSBzGIQFjNfS8z5Wl2i
AquMkqdVtbXGrAtppvUuvH4k+rgBxBfg2DwP2Jjkwg9YfsSV/5vmu1fX1OttIwhK
kvMs8kLxP6U5Fj85sCCZUTG4F+ZYZDgnTHFgR84XOJptQ/1kNdy/t1noptajRGFl
9iU/6MzY7b90TcCS4UEw9ty9X1M2/9bsxb7JQ52KrSTTGY7K0+JOH+yUnw8rALSr
t92XavlmLlMB28eewMBqUHeDaaFY+12iIdJtJM1lWS1QAGA1eMHzyWJlKVgbL/5/
PpaRs3uGoJIvwPhDOUU1Nm9Jy6fnPw1jXYT5krnbnXrR0VWbgM2OhdkchnwL+1OL
lc6nniyGOaYKWFDOhJsyuJmeki/og5WRRslp2Vt/3TDKuCe2E+5Oekd9BlYBQvY0
tSXl+a9TSQajSX3/kuU6+BRN0kWe0nVRB36l6w7JKcDarg4eEssVrvoiALXRxxd3
ZL7tEVglC+jp7rMLeRQj8CI7FZXSPuUuczAD9i2dLiec/YNBmc1tSLUW7XYD3W5l
xZd46sbx9IP+Spk63I8EGmIXk3kxZVIIaJRJvKv9rpKtbCNuIiZ3Sot0Ucfb+Kb6
Y2pJow5BddMmtLpGQEzlall0PFM3gViGAdcfFifg92dQINei8pGvYmz8IymtmCnq
LK5taKYef0gaQB+WiNd31B2PHopmk3LAvJjXhhWRIF6Da/qj275I4aanNJAEwKfk
kvOjj1L5I3qBuR1gQNz/wujGyILA8HA/Tb94BQggi2GQO2o/f9mX4+g5RaqFHNLD
eQFv4Ts1YkVttB9QwKeaNhO2xllz1k1EFyzgza31tn/yotA89fCKPGVriMgOaV+T
U31K0X9NjxaZ7NajzpgbDoVYKjbb13J/mETy72eMAm+IzDJk7c41Iq1nAzi37hFI
DNaSTIPguLOaAJ9uYmluGKGtV6txILnmdagHK0nmJtNRrMrcSE+K3MJCF5EYLLc3
dFgDWkhoF6HrOk5+Q/RdUWqJyDeHtqgs67bKkA1U4FViXPTgxGj4ouQ9qkhFwB53
PnvjkdS9YlQMkMwyHB0afmG2EbX2SAe09zlzLh3d7XjXx5OzXPRkiKIkrhTV2FI2
mIzwqLfKjo7cxgvU94W8FQamANkXS46Kcw/cfjiTl7k3X2gCpPpjOfLJh6xcEs4K
Ujz4AoCgFM9bb54SvUjGg9vEg0e2e+f9Lt5wmDDfeHIqwAlnPm1WbBDUlZVAs6OX
8qANcCPU2C0GJ1+AafLBR688AvFVpeODBzyub/fASB8cP8sOK5q7n+O+NjUGAkRV
IMh3vFhIDp5WG2CImnuLzjwNIyb4zax+ajrj/1uNN3rep3vbqbjHj6pRx15CLCaY
J7SqtR93iPcrwzVj9ImFYN585RCA0Np7aX2ouddJrRP/6+nkgpixp+1ArSEUXKZc
0T6y7+ICco8BjSVeFg0eG/c4yLEtiNdosdf0T08usr+NGMhrdoEgPdP32wcC1VMY
BEJdwJqRuFVJCH7s5dgjEz0Ybfv0oc9dgWWYUGsfY6IxN8cYmC1gfnFHSemW3ueG
3R3iVTPXdtkUk/6hW8tEwLiz/gDCxoztfx0nzvayyn8NHx9PM2ryqbDERJPm+mDo
IpFUU8E/Tp0WaSeDt7pzdDfy571OLzGl7R1IK67eJEbJ8HxjpuldQfRD+X4reTSj
+2X5shxVr/i5Fyxx3M+SfgSzsB72fnBcHx9L0EulBLSaxFtYVp2p0KuZZL7xBdyZ
rbtRKTds+M/UVY7TwSlywQcg+7FBmGbU6k2a7/hKeHrJpgEpioM3b/5Ba8sa7fKn
0XhoTOZQ2HtWY9xDNk7+8ZQJFfTcVvloHiusWWQ4PQSLdE9w/JkiMWofIBcta3QG
IbUPrq8lc7x99SrOThtFtMsB/Apcc7iVxLYwiOGDHtf3pEklano+4VLmAxKq9t1N
bIUte0A0poORqtzy5lZT4Sf/c/ERtUuiN9sczK955Q5LoslvjsP+HZtKg9Z865tA
M+JHrHOGpyTfE4Zab/18xL6i7idSUZledcKhfRnbNRtRL0HAD4zkUKOps21oPoyQ
UcZkYj67O6EOfgrkhpwf+ao81+kTxWjKdiYn2zNePI8QfUMXQNZ1LxH2hWSMYQQI
+SG1JMfDHr/HhLCnfM5UC6RSRZcgW6VNc0JgtezgxfvrMV7iCvovozXFGQyV9krz
8dn2l5aVm+tXNhZ01+i1d/t3w4T9g1c8/bCZArqvfVyMcCtZTic0SMe5SP2LfIRU
GFvkd2jcUM8GXL5GmBGf8t7eqiV+n+8Jm5hSapL9qqd2xQiLIRUOOEQ1TbehlxFu
A9zP6AXgevGki5EUMoza7be2MaaGkJfxwz9euJPyJdrR6V94496HgotdoyfIuzsy
+ZJjTyhtMblB7izfqCWvVBLxjEJddjypQHWfQ8gFK7FoxIUsA4bWQAEn839tSEZt
OfbB1N1hwj53387FGBB6kEbLt/2OEvoAvzcT0dPXdc8LXZ+1PvSud/M+uGSRR4gX
u0BpPmH8cgdstqySQkUN1mm1yhhdnXTBueB4imqlUgryF8Bj3XFLC/lgHdRXFZQE
QhauSMAz6V2b74K9zdn0sQOUVZLMF4OCinAkmuf7uXFhKDnzUnu3jPItiCO8pT5P
liNuy7T3+R700cvP3fxgjR+5RJzPnnjXCME0QWVx/QxV7FhEBzLRGOkA0UwZKGsN
SIUlNf5l9XU/tFpqg0Q48Uj56IWQRCCYArTYV4ccpH2Il9qMHQ+p+7TQVKsNw6sC
A0QHlaftDmOhIAkxKZLTW6p/T9tuAxj7jGEPjzOFV0Kwty0OqQ/4inVbKklcTXju
QocXYym5kAfKf/GSb9O7lPfoLrlJzJq2YxfI+ITYKqWrTFo+ikC5GZPfKUl1v4OG
pr4HeJ9KxBqW2/LFk6C6OjFj2y6Shvf3/HKwvQ63YABebAG+hCabgyq9w16KAK/L
qibfbb9BF15DXntm2XtqNzYiVMe59L74W7FQs4nIRhZ4XejHDii+Lq1y8uv0GtSV
hwsQD2gAszoxrpPFrWBUPaWyKCmy8Cup7y2Cdrhsiy3BOWzU3NdBRpLWXrCzHl+D
hdc0GN1aYuZkBZeDNIkTE3SUUc/k7NKVaQYXtq+NRqqcJYHlFiUwC9e/eTmrrC93
Cnp6FfmPpjCYrrTTCn3mMFfkpxdAdqvRDCnIDTkT8+UFuLRZSlav+fYPVJsgFEjj
Q5SKMESDeL0B7qs+yKkDCxvp7in3eWmnOQtdibOWESiAjdHP6d008rXMIOS0JUvA
0TY/1dPyok9Wijuvvdp3NffdLfY4MOdlIjgXCKAhCe3OcX2pPcxDkCWqaxsvYukb
R+8TMUaU9BJ5iX4S6XaqJWYRLCMCDlxt/Ry0n6h4bal4JpB60eRCzYgKV+KhWqLi
KvCL0+qZ0e/FY7Le9WCs+UdaNzByMZ5Obuc4sXL4PxYz49iD9aY50Jt3CzD/CpOT
oCxWKuHSR736XK7IVpH48E6+w5mY+c3etRqdkveyl1okHWWyVa3JA5l+hm+GyAcW
IyVQFjyIVniqrcfTR8MdeQqSDiGy8UOTeGpcsqwkBkO4KyRmrdUEy9RN8ePpWWc1
y4kNN+7XiupasFpbcRxo/Hddb6AdXlk5cs3s2fM3jMifB9ujd/9eYF/xqDrY2A6R
6PHFaxvN2AN+ukhUPZ/Jie/7i6TrQ7S9MKtK1QHEzNJSWXWYSc5KOH9JKl2nPt8j
yyl8EMkfaRBKE9Jv6xmjdkxUSEKXo7gtnFzdx19ErNWskD2Zf4FT1pDJrD4pp7oM
uaCUNOShE4izeKIx4+4iebancFBYeDNFEo81J8wG/DyYF0fm3CAogLkGCZzIJogv
wg+5tkXWXXhu18T+o6J+sW6td9KyQSG+bprIsuG+CpJ7NajgppXXJaXrLtmeixXF
E88FhXMG4iStXhn3YM2fuvTOwmNgQA57ZMgshUzWsotYEF2k0mBt0rnkjZZnVEba
F9uZlaMHI3XuMhQLle1UCYQC/Ht8V5b85Nm3ymZDn843yjacEq3eDK8WS0h8K64i
JrHd+tZkKuk/iAyaP6oNiJXZAHDc0Hsp5kT0DbWzXI7ouo6pUief6SWbK8Oix0Xr
Qt8MKwG1W9UiAOsk4ZOwlwePogOL3EkBcllPquBDhczJUXsp4HT7PD1c3ey0BJXs
QXdhd3256N8BYADYu8Tg5lNy1XERfnwomKVlBhsq3LlG2EfVn9AZPrXhRjtOIdYV
NLM52Hm+7MbLTQtYVkoajdWMjGht0F7TkI3xEzpXKGiw4PsDzGsnlU3xfcXlNOPl
hz2N+EzthSy/hL3mqPP4/7jSmdIkbTULQkgg24Ds8E+SQmszZ8Wq1r2E6wq/t+cl
buxvmSqQRTL37NB+LLM8KMXBqfNOwgEw3lFr+b2TKwflLZipZCx7++omvmoTsc4m
mvya3aXz+9az6/sgLi55JBuZHVQ3USm/KjLmXB0Eo9m8TzoI2rrUKXim3WAQiSon
F7WKJKRThYRNGrmbbSQF0BRtB+bwk/wJVQNjfhaHCxe6hACO1Q1Sf2eHwCSX8Wgg
QfwjZBFI/q7Fjnjkuzy1GdxpYyc0QyGXhTWvngdXfy3f3zy9XVZOdtLZ493j800D
Sm2O9NbdlTeg0dFXRdUG+qofU/Esf+YysL4S6blvOpo3Wkz0pZ0WiuLbCvAFlL85
7ewQJW7+WOXdKxiMG7WYlHLd1ujM36YM15vufTNP4tm8wWEILryTkiAzNrh/yNqn
jYqU8VEZtY+tiehpAE5mbmkwyv/w2AMbxcX5i5eULqhmRpGf5VGiEAgN9BISR6g0
QI0F+lwMAY7fl/msJVlDv+8j01ef2rlEE0R9+s6zHuRcjV+nWAWOCg1EZDNUoa/Z
lnSFnZMMyqGmsZxbzBvTleIRTtPcO0eRasRhCnOhv4bu7zxCLhvQai+OUBnebxoh
67xmoxogO4R++XQ8Lo4jWdqC80GeBPnG51xHLo/syCVjTA/897BhTC6gB1+MHw+4
rj0InDRyHT0ox0g8vHQvZAQRXSARXRnXOQYa0EP5tm0iy8S6wk0vV9K+dfkPPK/b
Vik1XdGSkhkWVzpxybgEde13Hc875rM0sUynLGjUz7hWOPI360jChfm6+tWDCdi/
VvPn/FCV6q/qHfFTvuBbNwr6CkHxBNiLebtMbqP6oKNsv1MrhlMUcNcu3TJwRPvF
in7ntO8uTlkj5BFs/Fg5iEDslcbsG3MnveXkZGmeI4sQSgvkpaA7VNmC+b1oj1u8
VLb+9ExXbaepz8y04vrYlNpd/U6QFdRTt1Mk0wUrQnRKZoWtV/ecp6g8MtG8MrtM
Z3Hy419m9FLy4ocdYY+qEy9skvkDDWrZ4BVi4ZHwwRmnGJRNQojf4FPRBnNwYq7J
JvqvXsD/KilKMjGAhSKJ0OnNVFYnv7A3ypOiIkWkSRiapvRhRK6EJI63SCqXxFzw
T1Cw1nvvRqLLI/zn8YhAbWr29sd8QsHF7W89bfFjNy2P71Jg6qMiyx977H/pwufq
/dkP/FcjZ+C2UKz2E+LIGuQxuoLYQFLeZ0J0PceFxZOVD1JwGuu2gxuEX60ynM9m
fvltBY/yTW9+EKSUv0QQBeGGGannQV1bbzz8fLnVGzPCJVmGNYODrmE//9IC1CS9
+iF8cxflEMJMMbTjG7Esu4o4htVucSP8GPDM9pvNOhaYqDlVOk8mGe/MjcfIeXqV
tv5yN+IOBERB/Ji3z74WgGWHQO8zB+V3mFZYWjcD2yuV1kUobuq4IearPE+3NWB6
o+Nd2BbmunJS1KVwGyH8b7yf3BC1A7qkvoAqIFK+1j84QGMhHX/S8tw7PpxWebvw
Rto4f292q65ZMIdmtJkmyMVgAqpdK+JRJNyvuuOHuV09bBncZ+J8Y/3E4K2G/U8T
KbSWSA6JXraL7uj/V85em8xtd5sT1U93SYbPFEvOiLB+qnpgbFKupb5WgQ5tkNHh
CLUsdXtRtuDWienr8REIomL9S9h00Illv1gM77w8lTyg2AMzQlQW7Ja8ZyPB6444
npD8IKU6s45+E5z59x+R520B6RnvR+edpKi3utiCJHvp+a8sIU+cQj8VgFOPhg6P
WjbZrADTYQEN7ipXq11uZEjYxxth8vwiunoMTCdNaQNwIxOdZw5sSF8o7R/tHukg
TaKsh+4rCttfkkgSWlQyjphvyWmhrPSUOpfo9ZZTmzzB5t5wUluAT/b3+Rz+zruG
2iNVPJL4P2DUciS2sm+jvSybu9exTy6fKCW/cKvCXso0+jx0k1hX2ge7F88DdmuP
C6mJQb8JjJr1eT+2vIjZLYUvRLCC/gwqrCVErQxmVjx1Q63opZjthtQpwIFCX3in
dIVhInuOyQAS00z1oUbdPfTRRBEB52k+1NslwNSrAyHc6A/50dFajN6sy9P9Msgw
vJIEfHYyaYHlX00XjBqgz5PTn4vbYhLK68IqvTcUDWxAoF75mbmCSxEKn3Q0nebU
KklvpEQoDytTBuzqIaZ+0RGLuOHyA4c+bOKiR5MdKT4VD3+g1gaLLBm5dzIn0bIP
nwuJddu3v8RVEPieC7xZkOXU0hIlmgoHqC6+sS5ga2vHWuD/I1rfM4SfYHZFLpnY
cxdOtUh5aiVYFs9DIEvjH/y+7L7o/hjZ2uShBNO9h9Nm6rd/CD1AsHgkcsO2B/DP
jNVU0FWWrV6trmqYfDZZMf72iwwrfO9t53FmwM6KF6feroI2hs61WXyxIWItCShD
W0ujig9ayp2EYF09OO6NeKJ3LotGcYAQCccipxfgZjFtkvns9YpllW/AGg1NGxgY
IN6unlSl6PIaFAmMmBm3CCzwbkQz3yxTXw5JlirA73xCW2MhfckY7Br1vGm44+Uv
+io8DiDjUnWScOzDNyvHnhLysuGcjrcmmSq48wXhbxxpsZGQVrGpWLwufHXOQHrz
6vwSh1D5v5hpdog4LjCBhAXZVUXgaMpeEqNFAk7rDSJArNx5WriBv/8rBazbbqfJ
EsbPFU24+qoupr5p5XRBGG25/k/G1X+NJzoF1leQMAmUYIF5rQw0mASi36X/CVnA
LVKpKlyvXrd8LikWNImTLlNv8Mv14lYm7lrfxAjZhc9HW4JJncppop5WAtdfsEcn
NJA1w3lOsb2H2FslNqedhPfwynAOFEpR+bjKtkofLlok0FMkMNXiFP9gdcwLUFTW
PvIXXZmmOKUq3SAupvXZxFB/ZRGj6OnbssM49z/bwsKYcSsYgksnfT96D28xdVZV
4ENYoR7nysiTLjnianALdg4O6hD1TAwOuS/N0UyM8dR2BsyPyq4a6Gk5CP0kmAHI
3PiZWtYrkcX2ckgdIzVOLbGoTHzX+l7tbMNS9Ch7w0eKCeGErw7br0Ur5rqsnw/s
RUkqeA5XcWQ/T4EQV+zRj9xv1ip24kfbJO2pMt1BZTxO7SJP/D1IW6AcVzTi+4jz
TB3T/CiB0BH7kB8p3FmOB1rleQL9i2dRc8zoOw81RNEeEcxJFIypI9Gq7Nk+ZM1A
aDaEG2EK9NSkggAq15wDeWTrOcj05W9RAtt2r0ccO7abal+q/FKzA6LX/uHN6aUN
ihzfzhhvVLJ5JUnXqXu2pGHt1qUZJdwi2ECSkcp2M76kiTUCF/wNV4i/kbNuEi67
ymCZpoUJqyge9ClCsf7MBDYV88RzuYiiIlAQrer+YI6umANzNo9aRdxa++1DLkbf
Ok+soIddoY06gJwvn+b/pZ8p+DjYHXCl8ZIyaxDNj2qHECkkbXQLfQ/sgyN250Fi
5z3+/SgkQYryOxUMyYeaOyblF6eAOvVj2/gjpfkNuySGuPLgNoE2ZB7Pr9ZaPGfD
og5sM5vRXpJaba+vDHrR9yd+9H4Vl0rBi6MQhnzcoNByXGBjLkMO+Zg+EyfUNLUT
qyp2ioVeESfyodDUQmou8U8OrkpmLcsF3BmtWyuBFsd+p+Cw3E6YZXOdn89lV95g
h+laTSmbhcJ/mCX/tLb/57ft52dRbON0Dq0ZLh9Xm3M/2hcsil/ubZ+kcQ/542C/
G4//ek0DmwVzXAGqdLXwnY0PGu/ic1wbuM/WNIbTCS8qaXGsLr2Pkr6yr2v6ZtaX
S4BcK/ZcROPLwHw3nNevfXzLIaVaSSz/4tkwcGTOaz/xNTHDY8WSNKDIyosNdJRN
aloobNjlyPmoxRSdEA3dQD42viZ0Y3k21gEpDlUPhpFWTGDp0XmrV2u05gPKh4L2
vdxOWvcmyCC0SSZgcxrTYMIoMj/LkEYOfHJ4VicNjHWOQWH4AXzCqrcctzPYBoWn
klJT2s2wa45sakc+49abFy/8zwVojFpu8QTZVydK8tLRf9ffs8rjPbWq5vtiqYx5
zs7cCc8p49TFc7PQtIsKMY69ujrFjRWRobHVUfTY/9h/pBs4ZKuW0g73SZTbRehs
NvRpffSYQ+JyGTrm7X87IpI2AtxwFOmWDCzRzb5TdRUiXEcht9dsrXIhTMux3J4F
2l5TS3KYe7Kc+pSlWhYtpGbRcctBUC5Zcu17w/vHny6Cz2GsBcjG9TyjwivdtANl
0syH+5V3Y97V8ffsC3l8JsN0pguk8ZCqVKY2YA/x5ikhgxqbePo/k6l8EpHDidSm
dO+H1+4PCvFYyJGtsrjo21+IpMIXY74qWUgnTICOm+DesLg3rihEN8bwqnBHMOmw
aNDTde4DS29CKYArx3hEfpylRR1VZd5Uek3i2cCFMQqxXzBdi7k1jAJVzAQ1xl6N
lCCmfEdjXajbTfXxxSt6pYIHSl01ImnHAr6JVdnYx41T1jZ4ieWfPRYN4vi+6J2P
oHwFALkD5rupdW8SvNJhATzoMC7ZyxbOlQunibP+v1Zs7s2qwEMXVfsGNkF5kcDG
8uzaCF6P4tvR9pWQRltCiKq3Wfqa91rOovfOd5AJ35zJo297xsXwWFelDGwqElPd
ue94vF7VdTRAjViG4LS9tKCx9WtiPVJa4DJGnVH5vu9kyGvV6XaWTQIjF54Ph1Jx
Uu1OuFuxMC1xjxVH0YaF+YPkwZyFLkU6Q03A4oDHMEgbcS8u/nulRr2iKUV9/CF2
5Wvxzz0yGMJxXUn4EVtE7K52qSs5rjhbGebrpBsq6o7y+5Yl9SRxKv9QYgUWggWv
i1o/tcZCg1L1Yl8FPbcgYZDcDvF4pAW53pXuEl73Qbq5PhSWFbDvW0NwugFFpo8G
49N6VFTbPbaRyfSOtcB6xosT71LaLAwcXrAINyjO6bfVsc7yjTiaP3oWXH39VBX+
ZUF9hBy2PRwFiXOmIwKajuklIUrUzBZgj3wnGSjivPnY+OnZwurboaWwXGD0kiaP
RrJx7j1Co8j6sQHkm+tcpbuINANc0fXMrI813JVwrqUsmG6CF8NGdb2TcmtDksDs
BdagN3S0ULOuu7F7N2eWths/M21pJ8O8filxYim9nL65aYtksuRkG5VT1trALJhN
5qmGxekqpOSX/s7QYTxm8q3qrx7ZnR1lbrOoDfXqqj3zUQsUQrrTpEigtVd54lqb
JsCKLRj3AjunUMdN0iyaZlHG4K2dxj9gHwLPgul5W7vIGU/xyTpr7+vKfyiUwXYK
C6hsF3hVbgq6uHoZUut820GqAtdeM0gtaZp08ooNQbd/eWwoLnjFv0jAxGzaR/7p
xDYrU/18sVofrdPAtQcSussREyDIUBmN4tlVC7/zME8rj1/uHuBeEyb4ofA2jYys
O6yNlMKABcoFW2rpB3j43lqGACQ32LV7yvCmL8lmjCLfytQREtHmXBjX2j7s6pyf
QLlwhDAnondhUWIrogv+pdabucG5e/8vW7oxF/XAg7jH6KghM32SaOrOWx2oInsV
MgVNH5SXFvx7CLEh1u6FYYH5jxxF+t8wvJATSgflYhFfGVGqoHjMikrF0pEF5x2S
X4DxYr9dVn8KAP9pXHsbGhVaiYYbH15exL1oudFev64eQJi2/tDuJPjk3sYpQKQi
jCXND37R4XOu9FK+5z2IZOpzYjHmgkZmHkwIyGz9EkEh53c5IMFRbmYnDKNfcauI
013Nk6ps1kqzXtepgDM5n+dDhRx3L91KrahNxoZamOMpx5QunKOMwc6S8Vx+vhHp
VOmPHUivmA0VX1b44tUBYemVGi02/tQf1df18xxnED24ZmUYXwN+lBmcIq9CJukO
iL7zWf/uiwW/lY0WRqMpjs11AYvoezuLL/oQYVr9tBwI0dsDgdV7nDVzUZBh7c+m
c41puVoSMLFmj9mUl3q0zd5EpTFMemcteMCKLhqMCrx/oBnv2V3LZTS3x/QEsaYz
08gHH9CMnKeFnfxdm/k3UbD985qShJxXZUBkhPCDGx+9Cnkvul1sjNRsnHZG45Bx
s7wo+MOlAn78QnM4DGdwPr8h3DYgPW/Kpl2wyaUf0dYqe6ZX2lcrfJH2z2bEYXly
UxWgIWQgNV9W/m5XJFet2/luxp0Zj9oYKFJLabmoSvzum6YFZcZVGuvjib9J0ydP
MhZXBgicyAD6r0LsGkiL8pHA90PTpxH4m+MWNMHu8Oi/PlfiGgWBFi19QvMxXyc3
My4FTUqi67I7mt791EmUCJ+qc7RbkHWXZmWMywiuy/5KXHRhgzDb+LdA9/HwSlPB
u/vdBUfVc16crxC1IS7W7RIdDTE+EfAoZOdfgRUakrJ5LcI8seniTLuCoCOmCUWU
5QXlBLnae7+OQFUahCY98536/6/dadrvctO/k1s6Apmd0JGHWeXxQ51K9WxLF0MN
SSLYCu9sDPeEvbnWd+I3mA9xTGVTXoD2pRL0pMOLBKRjY5GABC7ZkvPGtINbZhls
JClkb9CUSOJDtV9Wc8+Kgr/ArtQ4ybNQVr/wJjVQdyjV2w35geoos7RWbK0WByJa
sw1WBzNHweLshDmCbpcY1aiMHQXBJ26M6vR5zHC9KrTNz0QPkjWPabjEbYkvcYgc
2ewn2BmSnRPoH4n0LeVLH0aBDO5ONEKrurWndbVC7qiNjminn4BWxJubEprb8nEt
e/2vIkltQo9szRg0omCPtofMHkCqaI9LnYGuVC1NuQD7SYYP9gdxZD42rBC/gjYc
404mBF+dUmvyFCaxnmyONFIv5DP315PBznar7TsLOAH6Po1SAH6cf6pLBLbC0vRA
GVUcxjtYbaZ/1FHEwY+TK8N8p8x4Yqrbq5/920IIuOUlUewCqNjOqgFo+ZlkXQo6
ScFldFSdXE0GqqOKF1yEacEBJcKbVGSAmOCbKJFmh8ESfGgdQK4QmdSIkQoMBQq1
VzOiOet/7lptwEq5FIiEQpjKq8I/AW0CKdYisTEzExUS4HyyqLfCtkajmVK+hB67
iKF2EBCVIcm2MpRZM4xZBM1twkI4aw4dHY0DMckh7f9RUqRbROv2ssrlnhsfAGmy
+VsamyZDEXFmJPORhvFb8W7VAI5c9KK+9tIWd8jt4FTZ4dPVI5FxAD22Nr1UI6xH
Jx/eLRl+V/SZN+VDR44z0l4ip9V0JqBRmJ3ZHMLqDWu14M106EPG/Bw9R0ndQh9q
PIWKKh9MRUX0zvUKeQiPSFyb684ukp9BjA/1zg8E17AItNrW6L8m+cpZhROLIPDa
2cP9tD9ntnyL2k7LeXadCLb+yasyAM/PVe14UEyDdE6L1ZgTaZ3We/ZABzP9H+7a
8N/yMmqD8Ta5TV3ekp/1yBYfvDfZVcEq6H+AhLsAnC9SAU+hi9F2KBT01jLtUnTG
+kxPzOimBk4c9+1kzYOV9ZZaZeybO52nQCRMuri8zF+BxeR9V/8fGS5LasOcQaTi
8ia052SrzkhFYB3OsdKQX2+nc6LGx+jbgzvfn0edCJPq8ZYe7rXj0AlSNGf2C0zH
rGv14fWFo7MGDIBxnvjutIze0mGI5fEhh85Pb7jcKgR/bMqYJm5KaWm9SbliV0Zi
QCHIEkV4A59APw21PJlhuiHyNzGU/s7nRoucBb4H0TJqER79F42kJHBYi0nTXDn9
fx7cKPtHVWmy8t4gr/t0QqDW/SEes6oAGRU6NYkJBHCIG8fI1LA47BClv1guQoPg
tu0H+DELyPterz/3L/cLkf9suq5eBZC0RGuNvIZ7lTOdMdA9ezdn+iqYdAMOtoAQ
Y26beFG/FGodTQk/KhAzB0P2Wrn6DkYY03w6XvsPdkTlTU+3UrSf4nHX7ks0o3zm
bInj27Tt/PNMARiuLKvzkyUWYVjehr3b1zlDCb2ThcYE+N0r4TwenXlmyFBYIA12
kpVtPm7oWT+gxPKkNS5bR4JjwwytLADq/MyRVqkwWDxOFr/ZDTDKXVLmuulzWTFm
fbnMfeaLmt1gkY7Ld84cj9jm0iWJqqje2JpVIA+JMs1OjhykzbqAQ37auQd66WgR
UY22gephjWB6caiTS4JfJxOzYGifzhjmm6CMojT88JaTrDRcX3GhxSx8OJFUNID5
G7GLH8/GHGz7UvndieDWdBTJDUPGtZ0AWyW3HjgZVvucHt678qFDJbRLuWgK/WWy
FL/zajDU2h1I8AfX4x3myEasQ0hb5qL8iAAHvPG2SYjK4VSrmYp3xdPReBT8Cy/U
rdu++MbUC+Q48jd3XNLlQ/YEjQc9vFEd2Ct85Ag8TcoYHJ1jgoYuJeEDs3sfbrdl
3cCLhsyH6SrNbSpmQ5C+UBsca7MmfMrVX0ILFpJvIKfZFxJTc86NHIRfpkg4UusW
u/EOY37XJemEdJM5AGZt+VbqRdV+OeDTUFtNIRAAg3AdwSAtU5stBcD/Die0GuRy
VgRkVQPCwX/joAZLsdLJ1sKmg0cBI6gw8ubBS56+Qf0kXoISRTUXHKbLbuG+QB50
3nKWW4+NCoc3dOV2VXlHzp0b088KSS0/ITM5Yc899WFoKIuNRyd9NosmyEj04wqT
jbE31ZxY2zynNdcZVOpLp17MTgkxXlruDrFlIg7w4ztmn7lRqqzqf/ZsLr0fyZwV
50JzmO/eZxrFfVtzi8LtyHRU7von1uh9AIacpqMYavdGxjR0RsCfXu7U12Pf7R50
830SV7QLZUYU7RMKze7dOPSnNquhP6LIrveu0TnBUcBhe795xVVEh7+1zhxU4wf/
yV5W6WyVRj+vX3emBM2NyxkZ6IkPXS7Rqgjp4IrIr1Yv8VOJzMmSm9mwtk6GbT10
4je4IYDUI9hek2OyKmdsOlCfdGd8Ee+evrldjlBt9ze+OwJqihtoJS7MW8lM+6vr
0RvdJUDJ5MiJC2XPyF2Rgbna7e4SEGK9wMLEbpIOKWWitfa+sz6rXytlN1jHQUon
nGiMz/pCprIYzO7LpeX7xAAnXJgmAJh9nkR6tzXWsr+v6bsaaoPyPXSYvzxuxi60
ZwUSMK9fua9AClTF8AlLmqto5KuJvTVAN7kfCphErCRErBnMRXuCxe0Tjar/LTCf
DDvPnkwMzMBAtG9VabZ6MpJ9pHCNdzIHf8PMuTHYUDseUup1xk/mDfeGgzbZlroU
7S/hmjG+bC3dPyRUx6nTuDcQgBIMfbW+YcuMO1TOtnTVL4LE/4mBpKHzevSyZdkh
2EBVI6+IM3uC/JiKDW5iP4uA1aVciZ+FmJIsHjpq1sVUD3CPNqGgRXY2utymCoOq
GrYIuVlEX/bmCXcRAvNqBbmpiD2JolrAvSSP1w8tC9aOqte7bpfyAM7j1tKOPThG
+bWKHRxr6zZftJ/cvRyq32heacchqe8KdOQoE/k0bDKedU7pheXF6LudgQZR9ITT
79wnBo06a+v/fXhBjZAGxCC9UMuHGOzPc9UXfxPbI2FYubsrY55OEtOx6PzFmvBL
bV0GvftYf/oYn37APrPl/gFBvriGRWaWbWtJyyG6MVS8UOHQeBHvO47kGmgUO3Lr
Zmp2VeRIfT+y1Y4vRiuPHvUXdZN4zC9PddVpm1Y5/DqAJAmvbOb+PgJTg5hMarFi
WiNfeECi3mVfKNQISwRiToVQq5IWTk6zL8XMaf1XSu67sN/Ycvm95zgCQn7iVwMa
iyLHF4bSOV2fim4+djnchCTjuVWwCvV2FKaf0OlY02t1hlw3y38KL4jFiWHtXGjR
T0NOJ10AtCgJwjlwjyr/YSoC4P27bgZV9rkyByUaR2mCkE6+PEJsbxOlg1LpIKfX
KvHIJcwFO+Dr3kA1GjB3ezXypunmS7GvLOG9uG1nKEcFvTGp6TZGG4aEhaptgqZb
I8HU1yN3+2vxSraOJj0jMH8WSfHlm/hij2C2Prg+CsRdV6eojk/VIlj7O0M/vDLD
wlcc/vkwfSZTPJvl5A44I1R1aD+gyD8gHb0xVhZj2S1S9dblFSyjW74KMDPtO7Vr
OBTDhar44UoPs98L1sklqxQ5MGqnoSjZEDV4Xcb6onIDoKTc/+x6Muetzw4rjiMN
gIhp7kjkKpr6MqeTgFUxu+D2GPoypDpVgLlDE7ArcSFCz0oWUj6TSH13ct6EcDCi
dr/xgTAPQ+5Q09kenarSDIO58LPLrVjMuIyixxuIfnURW6W72mH7XIdad6nH1txO
i7l6enk4AeG+Ojj9MuR9SwDNthLL1VYLMZMDS3FfHlqAwBiehGzINW/bIsT3Vxw1
5D+3NG1I9IXMpgu7xywmQ1T/PGRiAchBwTn92VjO+9SqdpKZGOtNPwimR6EMLOQe
UvIqacj0mBd+nmSQOI6liIDl/pp1zTyo011p2P63EQXTyI0zNQae4KFPiSnrGIzQ
iQVSLq9hnOgFtSlIQs2QZeKqqHWXU74pfCZWwxYt84JcWZZQ7Ps8n0/53/rwt8V4
SukkfuLlVihflpl3Sk13yQzTVaWcjOdSvcoK4mdQHMJW0RZUEvKUaCtJ/0rA4/Ur
XkbPoa7nOtKUireGVFN6SkKiFag/L5I15Syby9wwLcjq3It2BEVDkcCbhrMN4Y9/
Nrkr2QnhcxOs+VAu/qFWvjVbb0eO8F7oj6C2mmZFf2i/BrI2Cy6nuKFvZBg6Q13X
dh2U3P/qctKUsDJAiMV4M4j5OiwuBU99i5ZzbXuXl7gEDY1BRaNONBibbjtLjZuF
qkN19xik9CkkRZCVPzdEVcYTkrPy40ssWdYfwB+o3l+jxJuTqBzJKVNKvW5DTjnD
C+iFZAjOaatj8BMHH4Lm0KewRqHGvP86tL5d1GCQJznzwPiNcLQhibVNZiyrzOFC
JBGZcAdfSPFUVATeSqu89g==
`protect END_PROTECTED
