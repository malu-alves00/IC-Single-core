`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
x9rFQvFhpSlu7WCimKMAuu8CEMsBVPzyg4q2L/j2UBhtOZa4V4R/inT3HmXE5tfa
BjZ0uKqHRsL+k2HCyZq9c8Xn3zjyKTr6Ta8brhrlDD7u6+VsEYFqErEyOX4wxPfH
Ht6dPuYXISUdkxayBjDMGOF8JsxH8pwJbUavqK/aARYOwf5Zpq2gAYnMU3tvms/P
QYXObtfxvRhkNUpQ/vNPYxIMVVufbKsoeWIlGb+yz8hAwMlTK/aI6AmBsbKNGwV+
p4aMBzaYt3nsQdB4Tf9bLdyGXpKCPau17JT5GNdbk0ZPPKwedolsHUgJCrxUhMn3
ULAPIRiajiyziOXHEUnb5O/g/UC5pNDWjxijT5A1PhiJZz8XBGeTXE0xzNgMChAf
10t7+GecRrPubIQbfvReSERp74gyeHDhsEWMDS8Z1tM2W58xxXMCP12aaaRZPsJv
ZzOrHIQ7gM5DF1qFnstRfBkWIDdQTtiMnk6M+eoGX09xH91IBDr9d4jlZmO67hah
qyk5s8xEipg9uquEMU90H37+k7tl9AuCrRmXZ0d699gfKaqk5x27/QVE9gcpy3/B
7SArAbrMqYidFWjvYzUT/muTAa4+E7MzboU5IHrtNwbTZqKdjsF8+gtoTXViVC6N
REp1w3xKx8WZEBGz4YkuGuTtIOMIAb8OuO5BSfLfLRHLMwRElqRZV9r6X00tpm3n
VEsbzvuyzssDPDkOhjX1mUaMzRQXkdVbCDs8igq6xDUgNlfbkJTxCY6xvWILhmIj
BjrXCEDRbhWOwXmOF4uSJMEo7C64VIJy5ailmGx/w679r5WOMcbtbERcQQ1InPww
Qd5haWY6u/TVnlmSFl5dInO1qnjODHLY2ajT52Fyr8prJ5cl8jPfcvmCzPhPQ4ZL
67wU7vUJ0oRipC4ge+l1yMgAwaPjZTL8RP3wedIVoqLRzq0vLJRX75gqcFT9yIuf
VudLqzMbt2YN/eb5ex3g020NNUCc6YwTE9O5g/lmUF8Vs9CGrIs6BRb2Tn8WRooL
2bgLefuhMQ+8PMj17eDqntB4TrTqYgg/G+3k+T+LCofovqphqUUdNDR64Wvw+Cuk
ro0NVX9zd04fNDNBILE99suy+lD0apvOVqmANwymVuIlID1WPyRhhMSueb57Bdtz
h1TUYJiqam1/FBgyeRw2nxBhfiwYLy73d59TVe9H3vo8eLlNPtTfygae5Vbez24r
s02bKPUB3jX+vKsXGeuFzz24kBrrU+aG6uw+tSih2CkEGmWwTJZjY85n6ZlCpqjX
/pnTDTYXc23cJvRrNgFqnw/UZZWmJNMsFqrFrGV4FCCyCRbXNcDTZJIbnGHrRHP/
eyPHROy1oN//4J10tH6/wvd695CXj+qRy5XBX6Bn1dMq9LcLYvhTpCGFEH1OE/GL
Rntd271Eh6GM6NOU7Ho/djwtYFQAk4hiJ4CjDN203ZNYjM5dmIOoPfqxa9ugtRky
wvLtVw2noHVNACRP/BHl5SlkYGULg4EDchCO797ZMFi2WTaozQHYTCk8ghIWp+lJ
bcpI5YfGZQY5nBD0W3z8aw==
`protect END_PROTECTED
