`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wxgBNiTDfFIF8n8NIOGxWNqMmuFgMLjaxiMdXmAb2sD7zA7O//Pcs+/rUUb/Olcc
u73NIEHRyxMvZOgElQZfi7w9BzNH0cuYIUdKf9SPFxZiKv9iRzj4ge/vqRyAwk7J
IQWuVquupdKIsx2lY7mA9afySnn11V58dW8umybhM38pWpXIBrUpWCo0bzM9LZL5
+wKKtni4LTamx7T95iNPOBf/oYt9SK1khwXhNIe+RD4CGY9mT7huTo1YsoCyGPQZ
zqj/Nk2BGHN19oYie3RfySWjEf3fS1IKHSGzXHIo2Io/QzO25wsJfJY4rGuMGVJV
J3P1ZUtf+XH1WId3BF7yv5LVzVve3UAeWjh5ETbOiPuLCEa86B8mu2yMDxCeGMRW
Ndi4i4Ag6Pad4zxxDq3BF5Hba/lO86kSRQ1wh3XiHzubF3WQ/1M58D/azbhhCJss
NOrD6KgUnfPizY9IhIRbwx+TO01v1IItX/ZpruBxf5lAq9IOxaUgVR3QbstQJliW
3rxJCslyOVBpYCePz4qV8i0jC3IYEiqgkS2Hnb+MTzuQLyPlJKB7VqNg4jRZEXYi
x6Tp9A4Q9TXqgfCSHN92113tEmcPnWlME+ZFJUpTFZh7h3cN6ZOCTjKewm9PTLx2
VLo1lGpbTOmpnwSCBOcpJ6ad0Zyd843tNxPZcSgvNpgZ26dDjdFO2fEXE27NOlzN
yL6qWsqCH50Gp10hoPeYFIrMweAqf5US6hiJaE8UgdMoXK6fyuaHAZcVmGhbVuSv
PFZU248yAHs6A5eYCYGEEroH63P3uGMmset8dNBaZ26GgH0yS32wpnZfZsbiRE7w
IV2rDNTaKKc29ah4/7naToNON8Wl0D3lcZc681881hg=
`protect END_PROTECTED
