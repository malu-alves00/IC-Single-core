`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HwWXnxOBwLUFPR9ulrAENuQhbyKJoO8aXprGKSFthgq7uyPjJWHFbFPlU0WxErFE
iR5zzIIIf+NCq3hwWMprdQtE1BgnYBfhllCWmFqCTsznaV8cC8BAdgNpeMhLKuXI
FkrGHUVpZj1J3b5EQkgLSqBBipfMmLFhe+eVHySCIeSwHA0aIM6sNrhD0jIpNKRC
kLN4FmMuCMCK/4fw0jfVtbkg9PEOIGejIizCXqWPhTsbfU3ryJaX4FCPCcdKQXf4
dQX5CtISe69Sf7dyeZtReaUSWPItlACZAGfOF0xHLpYT4orwj/JuAqqEMKApacjc
MmXqIuYBsGELdedilNmKS2Y6w/gsQAoCjyMJWF8OgevC4DD2bN3YYXmPHInBXPaj
S/VIM+UpkMNnmfHnxPNAeW3QBJoxg257CjlJdVC+OirAtg3cFoaxCkGKhRJ3Os91
lClJcRVhKy0zf3RMBgvwmzawQlSuBsZ5WyNX+V3RotQAma7hJZHCuI2rw5V/VuwF
Bt1nHtWjeHkzNn8pxwGoISfsKPHTdEzo5P8gbWnWFh97erwXNsCY1Hidf8Ki1ucx
mHfGKWp3P6EO7B3GR4MHVhVX8nd8qbkia1U0uMwJHuaSF13SbtDLUUW1rP/QPnJ/
W+5TNGqEIHs7NpmXPiq3W0PshzV70VXhWPrG3dcjyPwy4Ccfp9tvBD7Tx/m7LT+/
ndbb5DOnj0e2F8e7PkWNr59f0r1ulsD3eZ+TcuJr23EKz0NT9F0kaWoZaJH2JRXO
uwf0VZi5++1Wwjtjdw5BJJQx4SxGj5uk2yHJ26TZ2Dd/GFyhwjlKHrLioKWgogwi
tOuhSQZyvUhdIKA7PK9ddGCz6lO+XJ/9l0yilfRccNNHIHaBgVR+kce++czQ+LIw
8r61T6aM6bSqvq8IGSqb+q9kPNYE8da5UF6HiF8igXlskvTwMkW76JUmmezTB9wt
ENAg1OY0qrkZ19y3Gu1Dlk5LLf7Itp3OWhjM5eiK4Q1ayuXK6r2X27dNoP6M4m72
mUSBFvhEoDxnUTdjyYY4pZ+aJg70Ok9ErXfsT5boC0p7UHxopLF+PtmBHoxcHfi0
tFebsgCZHHvEq2+Puyt5ahl0pobjvJpIaa/7fkzPNGvBRKUSXJYnzwWMf1upKccS
Wg/3/drRkmj3Yp6SK5VpW27/vQxpVNw8Xkk6ISUxPM+/cvIlOQU+ZAc8aBih3AVL
0Kc9Rvc7D2/mketqnr3X4imms6ldGovbAO7eZdEzS/QlDbgeII5cJLPqB9NRQe3y
J4EInwIiXX6LIlZpgGtKlWYbMfdhNDyZJESxm1203nkDf3NxJpd+rt6Ff5iDfxbu
5K/eaxnl52BoYQpVYnXanHplPyJP3/kRF9fkggvhEcpJWmerEIw++9S3+u+U3QWN
Hr1bZYj9eRC7YM5Fdj+qoZrxgvFT1c+dAGuG3Hg3pWggzvRsgmnKojf3EF9ncC2R
plc0FSpf7lJ7W69jIYXq18nI73dchPStGwlyvhEcJc0oSRaNNZGPzgMe4eZJmOcb
osKBIXCHkaL0B1N0phM0HoaaT546uf0Vbz0rd/TU8sHFuWBEHeOiAQwT14nSlWvm
dJrhpTtC7rN3TnkYm0CG9+9TXt/lE5FKG431F3/8btbsWKbM6lZNO2CzePjm4DqB
5Nc9cs9WawA7uHYrg7C95g09PqWSIWxjGJSsVVbF+X2+jucZb24Q5FAOVj/z2WK1
UIEPCQMlp15hWgPINJUz5dPTEGUkCZGTlS7+mBIL65c/S2piTcDO+Nk1q8PYDhuV
21nJtQ8RdTM4ILrUj3eJsFXDxmy9UhcNGwjKzq7JLuR+kJzBhFaypYT0nfzE+/Z7
3OlpMKLAADDPL4qjNkIcmH7vp+xTM17C7liAO/v0ucdePBS+2L5E4EItQVckwdO6
EjmP+8g26GmhRyS9imwfRD/vzKTRyrzLVbMAPyYgYvcgnLVsAwqiHsR5jFh4weP3
FawZqwsf8yeGKdexblJkHRqx4SCAqeQe4P5Ia0+F1JZ4FVsNxK6RLwc00VrlxFCQ
cT0DTKWTUrOXMqMj97Ss4tMS+JAQcCWKCh8OxRyNgX9FI0hIeIkbzR/uXFKXuhf/
M8ThgrsCaUAhwaXcmwqfFhsylJhbAO3CvFF9WEVvVumaseb5FMx2Cv305kcZbY39
hvqLBha6k+RcM22IcclRqK5ReLR43Axw+/6Uhlj3BZYH8eFYDRcVdKGGUoeJlA36
5i1bViJkCp5hKvDMqIU4KI2TIyRpSSBmbxlxFbXal1+cYyAHRSG1s9cjHFddX4pP
7T7zHWgPATnoWGwKZJ2Nsvkns5AGhfTvs5pQ7rHeDwyzCru0YtN1wqfLMkvBCbpC
KkmTASmlj17O3/SD2MlF/VqC17/rrv4rwV9A96LtA2R5vlMse31KjWXKnrsbqokE
wenJnsyU+yvBhLtZzQm7KD+lYZmy4HpE+L/XtHIIYr3yXlmYjvTYKYW5s7BBCExZ
HYHQzlpwG8u3vwO6QFEobGWK8BK/8h7Oek5+bhs+C3x0Ws6tE6OLspXdkOGLYh3P
B5w1YjWvt+ZwKyHYAnf+vghZsNiL767P0gFfN3ydehv5hh8t2wEQiADwYKnMC18R
DwnhL+gOfHZSkdGjMlz1PP3pKRzQyVbAiKUl91oa8gJWuzUlNbc15hdb2ihY4IXM
lzDA5BgMMzAvAvOI+wzP3uCwuN53itYpnRNKfeCY8apFT2q/pQGr+QEJUiuWsziH
tPZ46wOXPhGbe7bM4asjIZ0R2awgb8hyS9EHla5FyjHn8bDC3JHnjUS5K6FTSSJe
xN6Azb3U5lprjolJRg8YR9YnjJoxxjdvCTpmd27DsgBviS8HB7wsLY3rFtn1aDv+
OOYJbPwtz0UwAmuFla3O1jRCV0EW4xqUMgG3s7w8FiBZDYKpyu9vdMOYK34ZIwKf
EHz7cIZFznaYPyJWYCls4QczuPJpwjNWsNx6uUoverI2F8OzvsPTy3MBi0/coJeU
kqS0P+XiAw3iMaBER3SyhGXgmuaV6f+Ecv0RK/K3Oq9uTdncSgRp1MILK9OVJ/pD
ARZVZ7uDJc63REYxtlBq8yqvqxoXyCSSzf/ZCwC1oK+ohOyBTVWRxP/A7Ux8Ei3H
mVSDj72xMnIfp2aBa4CudHdC7SdOtkIDkNyfNNLpT7K5f0SglYu9nvB3UbA/ADo+
qWyjYikE2BVjOydpEqBWmyOVQ2itzetkTOurSEov1HlYN/dC2trUcCb6mv0WbCdf
WGAGJ64vmU/C+6fbKEQ8Y6ekUf1NqvNylPwU+ixzm2RpH07kHElTMqOoF7JdCtmf
30At8lrHANR0PhT+lD0F6nyJV1us5dFwkxLVMIEa17x6TGwd/g8Y1I6bQpw8DcX1
EApjF/H67MlkO1Z+v5qhKIG5ZTc12ZvPjKPK2+YZBO8Idgji/jJCmQKsCuvlIllD
MBE9OlpwDa8lEpnoqrXbCR4UVWSeMu7KMs+1ranQQ+mpJIgs3UPW7aSyb/szwYf8
zWMNqulVzEx7BfHiHHK2oIZpBS9rAidj09QAOMlFp4AV+PKbj4V6r5esQsNfk8kL
OjUPNHixgxzkG3kN0RNgTav1qP+SR04EIuPyuV3DjMaxrUo4R15CKmIoieGuQuKI
mKbwDOQME6JofRbQPpKyGMVl3uq2tOcCxUJa1vC/rvBrn8zFmRhVysjKpoMism/O
LG6u3+kA3wQ97zvSAr8yfUXe6M8KzrCfY7743k5/p1pgR7Sz/9nGRNrXGlzOtuLB
I2EBxkTBIpch7vMKEOOv7CbE6IIUCQl5lETb+51ATAM25Q80oxPredGDA7+OvOLW
tCeAsKeiYtQ/40RTKz190F5QpLXUmmFH00JP4YBTjmWpe/nbf+RBpNPsR2QvSVjK
AAEidCV3bDQBzIkqZ4ffstc4pVyiQGUqnjbtxCHoRps/BpB0HbRdUv4zAd0BgXuP
cPEgZn6qddQbm7/E0Q/gBh4uVrHH7OyfbHbV3j8sfNioKmFc5S3XpgObmpr2a1k3
Y7dv8z+hyJKWjqo7peND0UfKyEHfcOm3153P2AHumFBcufFNiGkCNF9+DQ+HRFeC
ViEN+SfqTcYR+w0vqXvXjjHnvhQ13pxkECSW8M/YAfnyTmiwLsTXlSgESnKREVXp
df9Dx1oFad0TlsIuaVgGyF9Cscnimpegf2xd7eIjig7F1lHDl7aF4FX10WBzdrQp
JCnA12k2WbqAF8D+AOWOpI/e+cghQlsH5sfjU9LJiJd+ZH9FS2bK5Kpiw2h43d2/
82vlb45kU7XntCxpGPoESmgw0kPbTYlXfdN2a/GN+Bgy2vZvu16jxJaTPcJx6bPB
+yuKirMTRt6zkgqiO9RmbmSkraZRkr4AqQkYfKtDnYO/B46wT94xeE9XD3cT//Fz
57/RPt+Mg64EynpCq5p4HsYMFdFjxc3Ur2KwFSySXrE2B6D3w5ENppL9UIe3hIU+
2KZXKQ5uK8H8DTPGlomoEZbaV029++rLjZ+Ov7wsXiGZMhRzYbAuG20d83j4hfbH
daipTtdlqCy5ccFhx+GdVJykfwLSN88TI6MZYS+xX0sz1dteTlpcTrxq48Qm/qYz
ZgR4kksBDhSjsAoJ4wXZrVC0DqedEqCCebFq5tDg2K7XQ5OLj1i7KxcNQFsVzm2V
BlDFxx3QO/3BS+cNGLhnUAEFne2ac3/xaStKQwkUkXV4m5mu62F/57ghQrh43fd0
MUt1InznV4mzhz5sdqq6h+rN4+FpKouazRKlZFtQJuHqyVImY3pw6CyHXYMfEXnK
mWixyn99xUqiBcYZOao1N/L7CTp6OtDE77KVMbcMr93/hvABZCKRqorsX/EhLASG
sGYHupZiSjLeGuzSm0nf+Izwvns6fMMG++e4emkJNbo2bcO1OUIrVc8c085ehSXA
66+6MxiZz0IGRQ8mlEy0+v2plX03/3EoKwr6ZGUgx8f17wuyrxGGrhqz0MqyavvF
2vExHWyokkxDx4Q93qG9+pvovoq2AEMpj018mZaMyMj7jo7+ATeU5Uykdjebn06E
S9wQZStQPOihOwEFg8KVNjsCabdGJGiDMpTdi8Qw2o5AYak2D7SrAiyt/6PjAGy5
R2zz0u0nqh8y2xxUallFj1AM3KuAQOoyNvXW1MuSfokOCrJ6xLsb/pjVCxaXbCC+
Oaku3auCCacvTyx44xJZs7Fuxpfoko2sK30E5b4F+r/MIyTVyBCoaPKHsEG1LqIr
uu+m92WcmagqOEn6U1ZmwvgzpyCZWL0t15ystTlkKQompMsW88PQSszzojqr/HmZ
4lDxH9bQR3a313AzLbHEdEo3kYnV2CiJBl+bBW4o1YFibB3kA0QgxpZDqLhIjS/F
mkTP3AEcC9daJPZwJ41mDchJPJSCoEMGa7qXR1gV915PbKuW2R5eQssvDAGeJIoR
cI/LOBs+6mnm5YsY8hjO4IgxP5Kz7/K3LmZce2eklLyjjMbFpDfTNXRP+N1r71/Q
Iv+K9zJgc104xEjVoN53KFi5L/aHXKVHDDz7gPwAS6rWb+OHVtZR6Sbn5HAds+oz
VJVSYKU/fGmVlb/5+Qx9+GOkogiCqoDzuOEehkzxhKSz4Y7jzYQA71YsScMKJLj+
3ybr1BOlcZMQrqQw1aKx8rLcW07o92Mk3gGdcKyGtRpsVIat6HzjK9Lg3OoTdQGP
9c/z1A4IKmvQM+c4qmhX3lVaEV6l+Q4JRDljC2RTxjeCJqGfHi0dSmaXWepAD5/Y
FCWmNHKRPfxNOK8zm2hO24VsG9rIu3VnolZeVaMj95lPRGbZJiwWYxXk3Z8KzWsf
+qB+Ron7KhC0rOpEJeDmgZz5ZVA9iJGXhmfvPfcS829nAD9tU/IKJf5vg03N9Mbl
vQZitkaiMad1LsJNlMrfIlNs9nQC73FMEVHrB34NoCfwdXL3mkau7CtrWX7rwcmX
LFzfM8lOnZLtvoa1AHDdGyomaPt1jg55u3s5DKw5w8nNwkLPqMb0BCsjwtdmLsoV
v38Nl4tl+q/bSHjyn6LNv9xJNxqleufM/jJWZxqCaC6BXBL387Ja6DKvurg2BBJ6
SqNCpi9W7En1UlJOha9XjvzgIWcvFVp5FiE12JqPWH+Bsn2krQnjHqzEJnpzyrj5
tKi2LXXxFF7Xckyrpw6SAw/kYKPOqCT0Txt1mjWYD3XO8CM05oYFMF3g0AI+0XyD
J7GuAtyoKIxWnwrGYgv+kTdIdlVupkl5LD7nljwCTtGR+Nvs9f/U4V6f7FOQ1Iv4
TJjMZszBC/RpG654jLFT98Q2/Dg17FDbl4+9LqZz1zB1EifUC7L4AasK+1n9CWFw
UlOE9OJIuezi15+R9rMi3eENnlIirqFhR1YB15kRsq59/jcYtpFXYRwntEWcvaNY
yUwwoU2KgMTmW/IK6SfSjk5/CVQYWWyaC2ZIVUHP/aD/E81EZZzCGicLYEPT2tT3
CLtx1L3uFXJM4sLvWUyTrPUKb/nNJ14w4OhkdTkQSUyvbaQUOWylL54dUf9ft1qZ
CPdC3m3mzRLDAq7xl1oxEMWI9rWyk9a4Y2ku8DDd9lZPSDLD2x1x/wf3zs18ZXUk
AQ14HmyP+JlrSzwxTc6lLZr/Dr0Dg6jlxXNlwYAKA4cgo92g/Hje7UW2wiPCOVzz
dXvnjzoFeCfVEyenj+wlVND4jm+lYDt3jDqwzuJAxhmhiEs3ZzPr8dPIb1KuRUBT
qahLp2B2dmv9gzSKVJjchyYC3x2hG7BXMB8SO71nF8GeyoVFJWFfhXrnhSNcsI9d
hMY/QmdzIsIrSrG6ei/qGDcxMAk2J1EBdVmiLGCERRCnKjvHKJCVvOIVemF8meDc
KdpR+cAaf3RRKDGHd6vCvnbdm4Vd4KBpWlwU/UvFojitwtg9atprvfrsvmjySRp3
ccqtggzKXPIIm2m7N4YPBYwM8tWW0zba9h3ivWrM4DxHMMi/WCj1nrfT+ld2RHdt
w1i8betPu6suI1A3vaufW4+aTRN8UtCj7P/E8hiDkcwiEXtKApYGXbmo1aM74ZjJ
OeOlHVX4YeYip9WU91DIEq7MGuGKmtP1chHT2FuNO7CcomyKx/MM8HgBaHxKeb+l
dQsgXOYnx7kNMFJdKZqSDUbi7dYJvFbdxv4nXnZU4T4UCKjdrrrRyhAV5aEECOwm
h+e27QHEVnHmNgv0AAOBilCSion03OLHrBD3GqqBxR0Lon1Uie0kmh/yV1Xroqy7
KGk5sv7Td5m2Iez8uPkrJsD+3l1c5z/NhaixKdL9tgsYoKhUrHyAqtB32LQc/xuX
Ts2vW4/FbvKNhHTybW0oFbleUbLRU0wJiSr38iWI05GWQLcMhwZPOtxbNtfDiR2c
YJpdZ9hBHUoiI8IAc9rX0DvVYnD0effT2x168jq5/gGBgKcgzf/tSY435jcPr9GI
JBREjsw8OylaRGzYfHgWIIj5Udap67xBmM3g+memdlt9a1oqKL/PWVxuWgXbii02
eICYQm2Ww1gBPkpy7hshjAPV7diGCf2ER3SJth6Dsj+z1hZy2jXqi5jF6aGLer/c
auuswC10gDEa1FEHEW3X6dDmtsswvm2g/xe9EkEux7m7VBrHezERGeFEaAGB4FLS
uhRs2Fy4jMscfYGLEgAa/V75DmR9D4IJrgl8uOz+qFhwCMjvKFFGBOjrHL5MII44
LS8oDuuxa/LA9537K8V4S2yElBkImnQ6Es4l2mUOweazW16hrmEfSEzJ7aMBUi5U
MQLJrOXouEMkWbce4rZRh7trAM3RlRhyxfrStjY41Z+O4so4AxfnuLQKkFnA+zyn
SEpQ1FkgQ09pAkTHFUdfMmcSOQhQkFYYNFgHn2dDhlCA9aKoPV98XOza8XnUO41G
uC+5bwRUCQZrzQirH9mu4aJzBak1u5xgR708uYi7t7x//1fCMjSeMxqMCaEG7B9f
t31256WKaKNFdaULWipVXHUjsYcIg7p/vDORvrzbWmP7ujVvuk7JG4p2BYZ/Seaw
d1y8aaJQXSqn/5baA7vcYDCcSKNw7h1FC5BnVQO4HPwL3BbVpSxyyMTKZxQfCr5k
cn9FAAbEuMMycppulDP2X+uEAQCAnQNvGxbeY6AD/2zxAUeErNzDCY7UlEOx15Qz
0/XLZ9KHmE0rAe08+XcYijKb/PVGEoDM4UUEgu/NTwbIuzK9qa5PyWAisj1uRj8/
oihhQ1f718hTWw0IH6rABjsCi8GL+hOQa1ASCPik1Kux/gUJxAYzgwQbxS/0Tetc
y8N4X6cj8hS7AjQdr+tsR/jt/5ObOI9obdjbswcBhlMvQ5Wr3YwDIqlUJ6ltdBBi
w3dRIYci+F75wsuLbO6IUauPpGVXO6W8t/LZOEVvTDrnGh5wHq5YcXcy+CFPgpgJ
P88tF9GFCjYFOPRJLKiBfdJSXj8NvgP710dqjIMtprstszygP+BvUU4bBf7DHZz3
Ixfaj+Pz+G7Y0/NhvpOmepEjEKBBLNFRu2tmbYn1qab85BqiMws+F9sBZmHXKjb9
iXo8kFvQQFew1hHOruIArldzGJh5gNCpQVlvIMSIV2brfqsZiigrjTwffQbH8aEw
Jodxfz1MOjLZksG+TjJjtSCB56XEMPCjseiXA+2OZXjH8gTvmPpjAfY6XKh17Fq3
nlbNvpN7/+Qen0lnQdLPRsZDNLCXk9kPQv85EeDvVRfRfZkZYmOzXuY7QQBRU1Yn
p95Exx8FeQl2OE27WplulRUhfCtxHN4dO44Fwgc0btsd0DGNLT9kHt5isFdTqLCM
aUcOcnl54N/ElKV7umPnxSCTDsQdgZNneTH4mCH5lk7bhIXJgz7YHobayTSniarj
EuhB9gb25LneRgjZXHoM0hAT7o+Ht0+fPGZw1QFQLL/vK1CXH4ckuJ6ksueHgg2R
OmlSC2Qni7SzCaOMjz5NyG9ZcEA8FFY2efQ0pY+JZ1G3wRiw8/dvjZE8oKhCl39z
1/Zsoy3jd8pyIDhdXjmgjuZMrkJU7MEBum21NvA2xPQRIE1duC2XaUVuhyshRXn7
QGV3MyXkps62tZpyElTNo7ySDm8HQsdpbAitM5159ckJjYg/ho31QHGJ69os3VF8
QY/E2BQIBz5nmIfFoEAeok07bqCuzi9+7QzaAJPYtjv9Z0ckeceDBI5/cmR8E5Pv
l9CrcxUdhyDGXhfnImj4zYYY7PQKbXIM393jAkHJ5YTmsG3P5rxbF8L7q2ht9rF6
y+60x4vxBTe8XdHqcBvI0yv7lN1dRfyOaXqJknaDRsMMf8nR5Ti5b7X3JgyxVLBH
RzKiIE+RfdchGJNkuSoWTqmrdXP97mzlLEhN8K2w6xxSkSzPX+D1OCwfZgSsys8O
Rc/WEMLmZBGgKcXTFFHu3Dkxkjo49b8j4j+TK5eqwdqROsCcNPPSgv2pMyvq/mhb
y0fRtj67f4+hQvWy7E75Ze4rWc3jOe229tTUY76S5Mk4y1nXhXzfllwIc8CTps/a
tVW3RcU1/X+4l4EsycQxxDYLWz74pVZOucn7cyGxmhA1J0NJ5TSuWqjS01HKIW7V
kH9Hxk51aQKvIhrCFwMqiAIHVbqRuPBzp0q8XCeJkzkCYn2uc3SLYyHXt4JveDR9
34TktoSvVqLeC7XX93UrUGkQwzXi1rOWaVGQ+tMp5Lnkv5gtDsDdVaHXWzrq6Aqn
hK69ORnFgdHHC1lElU1aoQuHf/g+D/r0yU7OxUNrs3rinpP1m6gkCpooPOBkSaGh
dSeuu7QBb5ACmW/IC2MHobc9JUAzknueJoB/unbat4G28HnQMRfoxoz59U8VTveG
NjkA9N8GaP+3nXAx5ajTWI0U6a1eTADeuOHvgukeYVqEYzcOUWd0JAkq0Cl1zSb0
oksSl+VHFZJ4otXIPxFzTHA0QiXD2BR2jGeJQrSOmuwJZNj+BJR1jz8OC3Q7XDbs
cBUsVmxF4AW/os12yvxkSZo8abJsDl0Wre3zbBRooHrKntUgVjSByEz8A389U8P3
wo3JdKRfmCkDoLFc2zsy/LE/Gk8+eZIvxmMJt/e+ORKsJVA+wFi/X3dR6tM/FiO0
hOp22iAqgy8KVrYSiTD4bDic3Z6fF2KEpRPmYdd0sGplebySX6LGIZKgMnqkx08/
iMNtpiXbXm+C7SWKsj6wS5LXorrtaMwHtOAGsU43WTG85EHYA7pFtcfgOh7XXiLL
J4ip0i645TdUmlyrTB7QqDXCkAHaGgm2E4xv1iqu1EltAFzQwj43/XnD8M4lAVnP
c6FQZ+b3314FTGpsPXB+rH4nbhsA9xrz0/wBc/AxeIHxoTQg5WAT80b8IGU8SOWc
fTrNCKQZjxNRwEj3LQIjK4hRh0DUVteESfPyAIUgmNr5KIiVn/jb4jz6D0Bc0xDH
8PoLOXTqGLLMcqGGIJoIQSWaIAIxTG8DIVH4ZS89XHWILh3grUHFTGWFpg0bZTcm
PEAEWbix3Fp29NxEVrcR5f+h0jMGfEPvfxrfjQHv4D2PLEs3OIhf0DMcPH1O41sI
dpuoX9U+WRwW+yEcWysQpM8IGv3EgHGzuLi/nzx79H/Gsc6DperzEY+vepm+uXwu
BlszCTyV8MA5xM04lnkCqdmNSPhLMlYvTbYyXYDVcvpylR8k2dgL5NPFcr+7wM5H
djIcpYG6DFgRSjfItc58w4YNzD771q7dov42yt5JTe6c+8xVk+//gK3K6I9ZFx5v
hsqwQsu/Nx/BxNzR0Qr6hVXs3odgMpci3DwCbgqOT9s3JdtITo9iKEUZBX0X3HBZ
Zv1VchwImYgKxfY/DuxNSYKCbAdtQFlOe0hTI3iqLPuM8E1R3qj3fgzxtVK1TfFw
V59zXmdG1w+fVBCRHnNM0n9OoC+TxPiQzeg5zCyXGvS+XOZVVYe8/PZNa3LKWaa0
g63V9khDzsZDjHVbCGOD2lnno6zgkL3NK/XpZOWEd5txDrMv7/noN6mNkg95fDyI
SNrITR6OCBdTJsjLvnAw4nFo8KldlQOXOGub1eQbOZKwt14KR4BMjSumYqiL8S9q
cq8S10No8Nl0AicBNyJ01z+B2RRSF1gBJ5932WzC2K6JwxP0i/cnMtUeKrFS8cqH
zcpA40lL6ehyipxoyjHmZVd6i7/VDGeEM3RhIaeDNnwZnnC8fgizjDEjcdfyC7/s
M3RoasfXrcAAdecpH9LcfiAUvUp3B95NvgMg6IIQrzmTTIlBN4tHYav1lvNPkO8k
+nSkhcTo6LjXNTC9Q4GzCZJjQX4gPg144SvqgieMUYPYp25Cn3vOw9/7J+P8m6A1
GRSW9LgUPXAlcuKcaAZrD840THXy/ggoM/q5euSHLoJpEwF0JfiruMUYaNJapQXi
j5s5rBqIa1OnNZzmnKl5aIzFLzoNW78EItfHS8CbTa7hODggF/j8X9XrO9G8yySZ
32GBJbK+ftdUxBZ8Tx06s4gz/3Y16+ibwuDnni9JEhZm6tvMTzBfo2XJ2wEpbRm4
yVkTjHdW/VVVIFcCXci6d9i25otLf0h2VLjD+CUTd74P3nv+YOyZ/fUUZ/V3carW
+P6hyrvw0JHod6c/FmL+tbuW4YnKQZI8pzRlXhkRogAy51ZEVxoHAz0MZxTcNTDm
nfOAXGqu4gu6XkrXtHtw5F5a8zVdBAlI0bxS9MUo3yfHUwZkPOgaubDJQ/4KTTmG
lPOiT90SYEnnbmlisVEETnsz0kS52Q+/v7IQ7wkByUK269JAXjUG+UDX4d4IbhLd
Xc7D7SfsjOizT1BCpfGVB4XIyc2VuFhpXx09ovBlAilxLUfw2/7FZFQ5pORY5Ebt
1amuwr+jccCKWzrGOCm0kCYR3nnJ19QqZP5AoqZbXU+c6pl7PqqpdYXNKzJ6XURR
6UAe03VfT34UyR7tnPvN6myGOKuzJafYZJd4BezFThD35T/jU4iCNuxgnpAbi9rO
FNOEJhGvfFBM8rqOnG3CNpB3i2UAIDN8oPI1JrCXfkGpbS7zlzFMI6Oc6QbbgjpZ
fma+geoTX3yrKDthGhaVIonyx5vPecuNyaMDQiuPGAEliDAMQ6miiy+wJglpfMDu
xCAsjgDS9AjyABMzahAFxdkJm9G+fFXguy4bHRdDefDhDuK4nE/A0A1jYA+4h4sb
HA8bW7CdvP2CQArLGdOgp7F+hsKc/qcScVF9gOjSdIiS6tGq+8wkvO1B2KNMdezF
cBVkpIyOSOIV6mA3/5LQPzERlwY6qhQ2qNshhqklI7dEGDccXWjDtY1LZazEjDlu
fDD/3SRAxDuPSbQye4urr0Tm/dvfFosLmLFD7BzFoE3szjkzzDEmaYZ+4Uj4Uj3K
tndIEcqgrZaxUuHzJ9UsYiZhgm93VyxU7S8J6mRvUQdkEeRFVebEncDVIAarYUNi
gIB+J/SoG+8mGaITbNK2PZKwcTR/qrOVibXiYZo+NO4NtaJ1SdPj751/EAKMuwZS
Dhu1HcAh3w5h/aELwGwD+4eJ14GauaVwHvx77IUcjrLE0833Yx2NiVEYztqb1O33
JJtqfpoCWBhYEsN3hxBMXoDYGcrSPCGJiqQncIPedZCX46awcZITUt5PNJqL2OMz
ADvxf/mNyUtLETDxHUYN4q11Gk2WFtSaoSGAKxP/eYbWTzsxY3onJBub4OZ8Wtq2
5jaGt6W35+bB6QrXjrZM6DbYrugF+KS3yMAoIYMlp3KgiZJ5J+1ILidyv4dIbA7z
XlQdV4uC+YHNhv5HteATuhKAbO777pHi1Up+zN3QpPx2/GZ0COcedOszBr4qesry
MDLH49Yr/cqNwYMwl7xXsEcy/1pvwArdVp8uK38SEupQXQgm1s2V+ST05/lSJfjZ
t42BjoWVR2upEAsYMydNfCwz2lWSozZzYZsNbS440ZVJ91jdX6HZumnECrZb6L9C
Qca70PYl7Tnm6FpYKgBulBO8REN6jyLj40KaurINBGbhr4B047zS5Dl4rlpe6GRR
48LH9tv3gSPEN5IzEQ+fFSR2QogzmknWpF/w0oxWePXXolBiLV+giv7B/a072M63
MtRgsEBtUgEwttS++rKPmCxFGTyiyj75h7PSE2P29d3NOqPpyr2rKjJu+jSKd+I6
A34cngmfaDk8eQ8qZeldVeYtgRXaHVTuOpZ/TbpW4aq6r84ufytKopIdTpHguAwW
l8d7YYWrnBBeZ5tGW8Qk0kuR3Bz0Z/YnAqgx+27/xKUWk7kSND8lPTOb3Kfc6qf8
qsBHwmQK8plGOU3MULAwoUHEjw2Rsc9WLPq2HobY739na8JCoDJw8jdtj2ezD/l7
fOZlS9WVOFrag4ohC889d/rPAdk0DrbB7tjBciuQaBJ/+pWxaPHtlWi0DJ6nOoZx
T8wfYBm5gMSTve/DQ8nAE13IbzIqtO20JYJUWzI5AMX8l6havKzs/oDjj+ijYZhR
3LBvwZ3FMtUG+vvfJOJ7TDyhpYqbfcQWBiyY3HLl5oaSJZ81zjlxoyc+UvHTlr71
0mftRDC3QiNpa8joYYCawEqj/SsSkfRYmZqFmMLLr2cUa/q34kThXwQtGiU/hDI5
QI03tlCY1GrSFgSETdZwrFNtr2HQQrA2OzYmNV0EbJaIOWgJ/EESZ/1sIRGCdybj
y6EuezPrBT7hgvyNPDYs0S0CKTULn/ecDSaI2lzvX60WX32TG3rVBmqVNM6xfTNU
Vnrluq3EGMv6gV4u1gP7gEQYUykJde0sswqjgfe0H7ITFa3kFwtIY4CDL6IH769D
XrFfN8edDSFnzYQf7+nmKaJwovNW3FOhOnrL6PNbt3ei0JGCYeBhImhNSJZ9w5i9
Qmh9ryUU945GpMIpWwr+tcCCYPWCr5AiXSGVbb7I810BQRvdrrBaSBkNor7bv3tf
9ucDgseaon1IuyXlRcrKW03GEYvFmh+67PidcvwNFmCa1PWGorFxMfdnGGU7Bet7
GlEETE/DHzAZ+eWi2rCFgIeOx+Py5MgA5wdXSFEpC7UeQMFrYgGi01vTGU8yVGD8
/c+XNTlbLecba6sYm89pqyOcVNDlUwwU4BlbrBJJdR524fD+C/I0S608CD+PG/Jy
ucfnS4jfS7gx95u8c7QMrk0G6M0JAolLIRfLaL5UbpMXSn2h66+7zfpvTCbwRo+o
MYM15x5tlbK8fTa49cLpFR+JkeQmeMVN3yjDo1qheVcNQXEpPQ43EU41Ovv+JXRh
psUFNVSL3X9cdw05phTeFdj8Mgd9fsNu8iyBHqieM9UxoOGq3j7/NwTN+WA4ORBI
HqYsZ1x/2pqurzeKD+tFbdX5lEhzafZ5ZcRpmJomVfMoGkoW04dBpD79Y/U4phVp
GMAQfsuxgPgG3u8VqDIrRZcKTXW9W3jM7I2al6KkASHiNY7IpR+lpS9SZ06YxX2D
Et+CcqVA822mBpl7UYgg1Or4kwM0DqxCR0Cbmpg7gCt+wqFo69r6W95tvwCcIqZF
/ybiCBPJM3oMl9njNQSvsQp10U/sJEgEKtfj1V5pAbLtldaSYyTXGhMSDxJTd4I+
5j3cddWMQroGRVr2VMWPIFqRzxM+DF6cKMpmpJ36dHY7uXDrn/kWpAhF9wiSFCXd
fTv7fg9s9oJsu4plqEPzLpRPAHozJXrpdDgt8Cu9O7RscAc18TY6vNsqyJ4NLIvs
P2mQQcxeTB+kMQQH3L7vPQ9bEGl1r3rAff1lq/3aKUqvsY6hGXAwOAxToA/fLx5l
7tJ451L+MKoR0p1Q8gYBQi+JacexaPIah1qxHKmOkatHNyYuju/ujZymR2Q3Ukgb
K3e399h5WtfsQ6OoXKeTdD1Q6/MGlP0cX/UL27Af6QP6Ea6TTyuKXWhaUbKkVGVA
rw0238WyO6AxCPHotuMNwDvaoVwDDAn+EMs4WukgiRrgDSHPyjH0QgPClTKXS4qK
qeJs/pbe4RK5omT7Ml6BB2aw/6qK3m0c7N2ughRI2hYF98iir2tgnniRCG1f+FTv
UUlbHOsrWi/+6ackTsGRHpDmFE4QhMesigoagoy+MzO/ve05P34JFlvkUGfXYWmp
+3B0uwe7Ly7aNZWgUFn930WuyIrHTcCIYo55kzIhYtIw+SPBNLJUYBAJWWdcfAtL
NBJ49xwpl8tHhOC1kfLLjOEamIzfI0Z/UX9conrSZHiKgKACYGkqNch+r8YlassT
VHqj2dIh+25r9n8jtfeSEJ1G7vdx66JpQlsh11cLTXMIawxrNypSUeUbip20dZ9c
dLKJdZbtWh/GUw7i7YVUMsukp5wOsMerSVSQY56Fnswa1ylN6TLgmsd42dDmA+9+
AU17JYuoXEi379UxmfkwtOAJUFCHb/kRW6WLtUggICN5E5vKr3ylonP1h3xv3DxB
Ly1Q67cNkOszHWJfd4DFghLgKvYqMYrCKyn1EeILOf8fLiR1tTiWk4Ei3dDSzB7J
Os4dxgvOXqw94U+Ka2WMoU4d5xB1G/Evq1xNzfg/yhs5c8j39pF9F0k2YZPOnaDO
IhUJqGg/RIXLB2WiNLOEUpz+QzK/sRihdP0ySpNghNRMkGakyJSJSJcc8UeGPXIT
GL+OKpdJvC4UtcgAnSF0pTgeefp8oO/ovVTd2C5mSE77azT/Nqez1oM1TNQTPVnP
k7vrfPUSquMOahk7iLXGX9h8pYDxWdK+t3ks9FWqq69lf3/hwcUbKjBsZ/yqJsSg
0IX5666moJxfes6PK9K+j/ifZR6A6WQDkZNwkGWpufYyJqMzI6SKaeR7pU2XCqNI
yAVlxiCRv/amIWK5K9MixOYAK3dMAFhL0lfPoNWiyvndANQU+F0H996VdihX4yTS
Vwm8KuGa+9hlVK/PtIADDdVVzk79nN7r2Of/fRh6RbNylgdbrUqqLeasbpw1lD/E
mO8kA5TqNzDWUqbQD1U6BvJ+GT8pF17nHU9PcOpnwaTNc6CFXujY7/u/X9O44HSb
Ojk+Hg+meZt7I/Iifev5GjriuySA1B0l+232YxDZpm+BaXWygi9sjSgnW1kpy43j
19aea7Y66sVM8o+RpwjQ2DEYUnSHZQMclmzgM2l56hnhTOZOmh4pXATmW69z5x0H
Kf03qbjTqoZvi8KxoyqwSuMspEN+bZwiVMOIYwzgTFyzBhQh3Z3zhJv48gD7ojNx
ydb8FHRUkeW0qJV/xPRGh5x9glKraeIvYzTVSS//cgSr2q3llErdJiP8pEbrvjIG
tg524CnGl1lwjssLgmrCpsNJql2oUnx27xz1oJ6hmZ7Z7rPWH4FyZxaWjlbeZd0a
hwZHM7DcNMJnu0t7R0u8fmHP7Zz9G0wxnNudcjqzKZxzowfl9rRI2nxEHp2ELpwn
xq1UaZ9LszLf4pVhFbAyrHrS9xBdHvLUYUX1h4vYQt+lY8M/IDYRfcuQpnofodqN
RgJyGUGxd6u1V5UuG9C3WsKNUDTa5AovxI2sbAe1ywfUQF6AnpS4QgVy6u+HFANI
EZKU8J7tKju7l/QGmctHdeac+PbDosQS0uJdUOnzyCdlCbtZ0K11jxc2iS+nRUgF
aa5njTUSKyMW1vRyyF7rK9JyHeudZwThBG4ofTbXuUSbqSJuMvfvE/Mz1RyfFtwA
SlkcilcAUkVa1mXOhCerdFt/9DSwlcRBIZBFY+eED7eEwgUiJKzBh3WQC9RFXl0h
I4B4uRduP0mPl+dfmpgfGqoEXHheDUvlsRWYBruyNukLODx7I1TPu+WYxSki+4qv
53ANTKwHGV64Dj3EFzSzPkk51Y7zuGdGWdMJFRL8kfsw3cZDKZsZ7ty3E2db7JeZ
AqpDTz4uD2ExPVzmKQ26RR3+dDgh/MY9wvkyoo4qQsHzoS7vH7UL2hlk7VVPn/Ny
hr4k6Ixgf4ojjKENUP5wZsDXwHHFKocyij9TncML2+RY6ayP0VMYfnpd6qviN1Z9
wDPPMFo+GZxKVSMlnPaVb6C6eeUYhM8dAFJe+NNDh5pUVTjX+yL8knvifUf1zhFe
SIlqFf26vjfE/VzXlfeccHG/O8yq3iFFcKzCk87UCwYVFBmoMBxYI4/+alDbNqMZ
8HDkTj/0HQ28SpDDiBpWdadqsJPCWCzIF/o/aze9gNFGfycUJE6AJd94CX474Me3
cG+wBjBmrf2v4VOpFXaAHdHr34LmDrnRUZ2yagigE/M1Kw0J8LzsVFkRIj2+4HKS
MI1T8kaJUTEfw2yA97VnyicV/r+tKP67PD9I1eJ9HdRvqqaEOVZdajHilevWmUYL
iKurmLf+YceWmdlt09N037DYjsFQLQsW6y3ppZONH6CjOVwC2yX7mYCBDn7bO8jI
oXwh+jLb9hyP5O2NFRZLtCj/gslAvufHSIgLjUaaqflr35lfHQ8zH1GDLybQw3Of
mZ+8L8l6H1AJyPrpsNDuDRIpdqiio5+fhYov4z4W6FuCg8yOMMvpPryBjnY3ctvF
fRxoMjmdSRQG6supcZyRmz/q/5McqTNLh2pjdhp5XcPCX9YLYHcCL8DF3b8MOh4j
I8bIoXJq13O/hq5gQZNs8dMPuGZ0EfgM0I7J5hewMIRZXqgOvnMogbStAm+nVytb
W2HmT+3Rr2bOy1TalfNPzMLAre1wER9KTb6YLf9sr77S7jGSbxVX/2f+nuoKvEht
S2zF+AZ89KkfkGDfohHle2CsdZ8iQ2VMvrEf6WztzTIcNBUxfi5YRobZrHRL8eOH
XeXI1LLCDjZeqzL2On+tASlgIWPoaouBLIkAjWUKDXYfP9UlNK0wi1IbbOdSCfrt
6ddYaQs4xWLPJUIQCl/aRixrW6SQEFCotv1RXzGbWlxyxPFRXrNBhBz6hWm0bU+k
8zZCoO0gzS47Ljr8nBR4+oiE2z4v69f5PLvTPCQQKOho1IdMBuW9W0o4C5DOuDSY
VuqqdBw1lW4A39+zmzQXLM7XOEoRfohL6sNlT79TODGrU1JVRJQOiDdohyZn7zq4
40drajLs0cbqeJYpfivfBs4PfEMtUpvHobi8/Rc5bLmrR/mL2QcFPZUKS4GGUnb1
pjSKMWwtNf4s2bzhBsaRMUKQjz3RehekQqi2NCB2bnIhjSXmaN4KZezOE0/zy2Fu
Y8oukxtNbeYNTEXkc/LFvUbgfpw3Sm7dRa7ShtKfhqWG0EHWg8ZPxfWwOQVZws3k
QrX+UPstMq6fnBbiisMLtstHBNoFPXaodtyfI+ySm8e4XRnjxyTgWMDRA5ZwVEgh
o2o1oAiIfg7zUzMnbJ9Kpdoi+Z+Mny6QiWc9q/4GFfSibjY+axHII3NZNmXNzXKh
sazDILE6zGpIcTh9mNgv5xlC8D+q8khOxDS76nhbxBlgsM0eSlK55MInhTBtzDQi
e2tohJH+lEEXY7EC4Lc/CeEP59lLxM945AdHfmwFl57BqZ1LBu/UXrnnRCNO8pH7
AcOLb11vAdT3M0uRB19aSVDaw8m3sl+1baelsjlJy6fN5yiOgzofDff3ECk+iVSd
VttS1HxbDZLYgxLKp+5lv1IfEG4QH7v7a/68KjOpHPCDVk/ItPt0mlXCHW8VRFid
0VU8e9BcqBdEpykRVKqHgpOGsNcSZ9MYG76MN07xlGIPDDReEfIeHWIkCMOLWn5w
zqqMCkEKASbVm9Hfl8GPxQjvfdejcwoq6V3IpJr3bR27NWofDbxD2c61XQx1PHwK
EiVfH7QHK/VszuM23nmVZEHUNy/jj1+WSCjE+7LqKhVrXN9xFlgrQ6zC3Z1vhvO6
isCRwFhPNSeihZmwBvzgO5VDWp/79R/JEUX94lA9jf6Zh708sN7HJkc1/bSz5o7R
0/cSiOuY7Tu8T9xewtehKvGjabS5tOs/sS0AYolHYB4eeSJcJpHYNrQi3xnakHhe
4fiYqZ3sEFE1rXyq769kzrWqidYie+VJJt3gu36u9jhDl+qLGzTSuzBp4isc1hRV
gTPsox7krE8IUikLVr8b3q/JshduQKNeRfRqrIV3pZXkgZYfxxzFg788LsWJaVFb
Dw1N/kuPfzpWItfdlcC54gWV5cJZUBmcXSqqG1oYJCb3mrdl6EDSDHZLDMycOnjo
Frka7D223T0QdOl1m9JaOEg5cVas9tSmXF9Wh3Iu40PHfF2x8eGsBtzp2cOacKfU
uhc2KPTi7az12qGpjJkYVTzSdO1wR30OqLwDTBeIlBTtn22WE/Ij6Hc8MeTJnJeS
6df7X2m54T77y7wYZ+wLrVeQz2C4Nx01SQJgYLytFD5O8EwChM1tSRhcMcPHv6P3
uZiZ2LbopHS0OFOTbupsESVOWAubNInR5CqV8qbDq++juj5qWK4mBY4mYtFt+Lwl
YOWvxDaMAApqnnA1GEi3GCD+r6k5s+qZXxAOK0jZtxGETQbBo3Tv2NpjQLKSfAx7
XB6nxrm+5caeRNfaKeVpG+Ow91XuLnVC65NCtlEO35QzjiJWrX3l4RjBfBzwvtZ/
E0NsfxCSICllfqn3sjdJrrach76KIrYkP0qp8YDdpEsQbnpcv/lr+HJe7k0IY6ZE
7dDk620ulSkvNGRdvg4o2TpuUgpFZNaWyxHPjjCGs8gShBNR3Y+0aeewEI1uAxGb
AJUXJYxNWnI0WxI8V0Lk5yudByaVi8eBebKF0ZScxX/1KrDNMV2Ci/tX9LKzfwd4
fHyp6hbUbQx5Zo9FFocpbf2mw+KVEz1eJH/mlqTMJzT11GY2XR0TJWQq9r81jDot
dINBYKAjXlr9bpy1CIr52ntpiv64MimZAv4lvyV8W1O/fRFtJHOnHFbfeQCSAzJb
Zn+XiL7NJsfay11xjQnaGiRJBykMBvcv63xco1zf3dDP/w+P+kL3NRxTcpSN13e8
ChBJogbue9PvtSoqE5+9VG3lu4tkC1+lvR+2qm7CCr7C4Xqy+3g4RhyQcA1iVvwd
ieHxVVgtuK/AQy6YxydH40X3ZjzUN8aPc2PaawF4hwWkwKmBZOh3P6q8ny8ltjEp
6DWaYJiqtGILbruHQvb282VmVz8kkTlF+vw6xmDdgHtoohPmpt6BsYFvo6xZQ3yn
czDIr+UPfNm5+y1cgnK7x1VGj7AxW8M0Z5DYDoPPk/VfzjpxMaAH7sWn7a3YHrEv
+Jqa7oWcVVfcYRaCbn3xEiIH87dMua4/MKT1rRwRp9xGTbLArEN13JafoKLEzhIi
gM2ojRpUdFORuZD/hiqRo03np7dp+wj30LvaDnwL3WnAHBxLgg4KAVC3oi9Snmr+
kvMbJoNUoggzwvjfoHvORT67FwMMde0CI/CxYlSIdvf11DSDrSt/7A9cM1zcTt71
waw8U1IbJe5b+ccffj9GwzimJtrY8jZdtzPjmVKJ8fn5bEoHzg0k0Y88/SaX3vH2
siAU2CNSZ2PpKOulJ5EKjKBqKw0x0qmIHLJAV5VOjATx15NWanZrph+Iw99Rq8Wl
t40rgkYs2zcm/zf200UDoxBdmCb2anBo0ASJ9wTfWS05+zhp+sYKx3T/l9f6MneE
6O5JYnd/MJY307V623Af15T3GM5k1f4eSRx1Ad3Z5n6ixE5BBXKoK6pUqoA1kiD5
pbvMu2vrA99W/WfaTF2cL9fcoRjU55m8mjCREeR4ldDVsp9FZeIKypoY8CZkLxKN
Nr4iY1+mGGbuofrH4i1Hs0wdYWSmYdMIAPThW5Z7GccwPA/QCBixixHP6V1zLpaA
DZRfermNycv8XBrtWvFNIrEuxKbJNmh4pSi0v+czuGTz3KoehplFovQvdHnKqfzU
nW9RLltAJGKC2pEuUQl7IIIxw9BtqINTSk2aYTp83DDM0fNSTYWddIXQKUrT0E33
xJ40FT9T4TQxYRhYP8bPp36mlJ0+g1Z5Bpjk2lON2aA5kvVHfDgOLpg9qnRUWn47
EYWqllrqJc2nJE96vNaFWgFMstqwtyz51NbyA+OOzOBNU178ikwsrQRFd8qk1YhM
bbImmXPslmf31Pq+PyY3/mPbTElQL2RzBc/d0huC0kDlWTf7VVEV0WXaI4EwQIV9
c/42TyGERFiwd5veopWosPRptbg2TFm2qjBEWyXWpyNQvKijhPT62Z5ciuhESzEP
+MywfCA6jLYG9B8av+FBI/58wqR/tEn9C/vpftPEgt/NRTmItET26pvaJw1zSM6s
qI7ML5rSv67WdX3VNPkQcAJhW1/XHsWAMDIFA93rf+G0mPLizA32G842fiQLtQIB
U+/FeEqw8NQ9wDIAokXNFsgEZ4PwXhxkcC9Tt75iEyPSfcY01vICKBQ2DDTJ2SL1
/49k38U+UN3sDLrK2b6eCiUAx14u7u5bYehdOY8Des4/MdfFISr67iuM98EZmzsQ
S2Nd1nWdpinUby5e5ajrKJ1UjO9bOmXkFra61D/sXrdLi9wVtxjwFPwFVSH1GKiH
0IbqfOpA8fA2YEeYPsLxxizBdPURKiyyVjfNay1hyVGF52X6qGwgXhyja4Nj2GRG
/V/TP+NuyNgEqQQnN1dO5mnuc1x+Mlkd17lGvlmcDeF/HQyf0g2+ejZOMc6ULBzH
zNdOr0fax9y7bI8ADX0Ms6K5v9ydTR++WGAW4Nqii75jtnVc+Z8V/ealp9a6JsLL
Zv/oTVb0YAemb7EXdQABjfjZ2BXouZheu3wKFOxmKTE2zOx0wjN3EkN8E5XxIYN5
b8tMh60ETt/TpvPsS2RUYSbbXqsEfCvs3J8w4dofhhjtC5Gm3yTJWwUvlWo4Mn0p
9C5CdGuVMoZ+lalrv9cnyA/c8x67NA62N8vJii6mxlUg2skFnxNErZAhpWFX//GP
UMuK+jWEJ7n//eTzSoO/chKfurMAA8viVyjU+BaEl06DUk+YF//NjZtW8oR66/Iv
DpL//OYCniEbWYvlDGl2+AU6cPIAUEwHFBe4Kzb0Ih/8KlKF5u/pvGhRsr6apjU8
t5XDKbsUut2s2n6BHBIKN9xC6YU0uJ/OwPDsQpl3qoIzpWQk22arY5s4VqUzpwbZ
VeWEKS1mizje6fblUtQ+cdckSs3oY5xINh/DoMAKMuTYsn7VZDUFI0yQd1DyzA43
vYMS6B1OUpuK021qS5iD0BXQaPccv6pzY/05dRPT3G/uU8RpGtamIE1oIrOhbMzp
i6VBaOYEUH9TfNwhk5pkWbdwISMzVcB2fbkA4tEOXINMOcpksh9gIFyV8wYWaNmm
b0oQdCG8BybCV4rePkRqZO8gn7o9Jy4DWafelrcjuks/D2HJwWV5jjwJt56IKd3I
uGvhS0JMMasGc011OfESRvptpewd48cfaGHVoRAA82dWvMLlwP5Swyrba7ck5YU9
99ALktxoMXYXYGvjLi8kO+VvnO67RLdEP6+E5gAGCPsYR1tHN2uLwjKEe0fi5rmh
fi59no2PN6/8e2p8Rb8X7AmozwNGl6KFeUic4C7yOwmjOEmwZbC030mW6lLk7C4c
/P0D7NM0OaBzdv5UX4fO56YSD4aYpPySU7EXUPlqVZ3LgyK6y/rwqnQbV0qBe3+b
wzPocZpUnPApz0chVGtllBiEShGqCMzVSWYMXANIhA6dIen/yaJaOnpnW6N2pF6N
v0H8KhEUvx10vg7Oww5hZJGYyXWt4AWGQRvvxrNo0qwCIg6XsWgYJI0DVYcYL6ow
O2zPiKw5k41mvG76C3oHKFu5U6WPAMoiakP0KKToVKbzwrG5v4CU+j3Zvh/0XePi
9eFybq83yKGSJl5nnk6EPl/lMAi8ypTFGJzcCzZe98EjMjMFdZGHjZLYs7+/8Xji
NWsl4XYw+vdFrldqfmEZnc4qN2HXi+lbyGriO930Gw8X1rErZkCmxMJXLxYvy7oe
wn5+wRTV4QgUc253GknxzATFL5tCBlCxxO8w01ap5hBf6OnIsZr9Uiob9McdQ+wR
rmDrAqo7jvJu2UoLj65B68yugXfmpfz9g4ETwQ5nvEnzaJ18Zh+QAERPEAblPR2d
q+raiF1FYrOTI0ya5spVUnyeCbIwdtUJC99lrBJx1anDxtnaNSoBzRr7DYwNQ8Kj
0L7cZpeulrKbxWBqjviJKpq37VYqWJILloGob4SAwpTiVhbVWQz0PUZNg7NyYAzU
M93FXR783vnfmWRJJWh+y+Ij5FbmJyJi4oITJlM3EM15JBlWASU+hY9TZfhmbgED
n28XsNLp+6DwBhUx7lWMUzxIBzXm90igcXrorN2RTgf5bTkusIaQNNwUOMVn/3X/
jsfwFxBy2NfXp0H7Fg1VayTCnQMpOWGQQ3nf3KqTDSIFcGSQZ6y/RpBz19OhdmVb
yOCY17sdFgeZ94h26V0TS4dcUkn3OHMz9sYv0hfk6oGwef0GqOVJPEhp7iewY84w
7e1rO89EBINK8+k53j+uV+Q7n8Koco2iWfGJ+7on8cGztlf/qHtAc9XVgWVJs9ep
myMKRztddtfh8OS8emTzNnIOePWjqcajGeB/DDxr8j8yb+t38p2285bI7N8SHMkY
njgWGVO84xUGcCV2vJ/+Bak5u6vc+YXu1NTr0Crhs7LUBgRD2cd0ab3/G6fFh3KS
5OjnwMvfD48SKASJW0l8anhRbDRwmPNJstfz8sOz3FBwwz32ChMklHJpuGN/6YZG
R9p9OEQCMpvWhZGh8CQihiTKF63YYCeg4eSTHNCTAy2voehfaLOmTd45+tWTL6zA
XTN3A8O2A2jHPD6xpJXLaT6DtpcJieoVEX1ZGkdNMNlQ4NkoTRMpk8AleVF+9j1d
HNzizp+Z8NKJUaQyT6xf0M4FRzQb5lnTtRKGhkqSRG7bHxDx/ho//lW5S60KVGZZ
ICTmZga3iLWTGlTF/Oo1OKZXCi6br3rXPzKUGFfFqOzZoyMVarkOvWY52ueLEEZ5
H2obk8eyLODObHmboPGn/bdWXhhMmbNU6KYPqcFlnzmXWGqvMfAkj6QU0BcjDEM2
uGibx3JpJzned2vlQbIh9GkoiqPijP6W1riO+PkxawPM/8Ac8/50Jbnc8eFacC1N
k1GyCuC3ha6pUF6LJA62NnDeLli+ISppF21D/PcWTjrsMhTV+ozLFvR9kOnRR0IL
O6mO1TphaeQqGjZlRqLVad6dMl4WtVJhOTZNYcDinkoXMzZXHnf3Jnq6KYKx5Mag
8VlVDCoOARpAALAy1lU9L3HVfd+eKbDKuCFiyveSuBwqR6iFDhDnmpx0NzeqLaNu
Eki3LzMBWOnYACc8Pks1lLkfGAqoNTIxX2IERqp8P7H9kW1tjmK3cSam2NEK7Qo6
DXGRLk0iG1BYpyiDpVlojWsG+/BB5+qN8NSAG+n1DF2zkvNuVncvVdAaY5MdXMxz
YUFup8vCAwsz15gHwKKG/HpYCDUbhCl4j7T4rt0/Sngi9oY+qmNmwuQqitM0TtbT
x9DW9+f+dg0xhgX0/1OfB8QYAyoKkIQPkGlqG3Vq+vydyffgDMQKkFtutCKgCTns
7cJO3HiyqSNk9p6cD1Vj1y8rOCfQ1X6hsH2tln8C4qrBESAaBO7WnZmZiTEf1DZG
zhNeyUpPxiKHDVG+v9IL1TceOvUHImr30G9mCwc/x9u23L7I4bBo0TyAvLN19rCT
fj6io5wg0qvaac5CAmU1/Cc2rubp6DSS4Hud6CssWXSuDxaC8tK9lHxyUTJz5plZ
8AdgrFUn/PRph+TIVicwzj4HprH5Um1YdUjIxgNi/BDaLmqItAcPOFKnVxeqXyww
5Bfn15Yg3jRZYT76pZbsUNLFJcRDQGjQNnzmwuj8yBXhYtbyu30/QLRiVwQv8vPr
YuxMP4KQNthWhxdkwJK5INqwt0htYg90mrzqGISz//WHC2tg0gJZjykLYNGzhzD+
ZBn7F6AsyZpt6Dca7/hh8bwNQeexhzJdXZCOoHL/xtWRsOK0rD1Ti0MFYs/b0vYQ
MKb7zD1MRPPZ2h74m7X91csU4lm++een3SZIHL9rSR9/8PoO4e1gBfNche6arVMD
fP7dyuO539IJrBV6cQN0puCgE6aqtpGOPdUr4JM5GefiionPOmQ7zqr1e4VeBcn0
o2sSBY/jg5GmMJ38zg2mY6V+InnzAMJ8fE5Tp4c2ovvyhk74oE7aoxND30MT/A9s
hySJjIO16pAgGetdLcQMoPPg3AddTX0BVYmVpEqtoI8fdbA1yLbwDEyE+HpjcbAb
bRxHNm3YrAt4g5Z0BInzHabvJkrtUXbmGqmcEqCsvCuMvqzvw7yotwyyUd0JI5+q
YKQvz86gaGfvvoxPSqMFStor914NHaxIEOTAfcwcXGtmJAeaodiwWYjTLSJgCbA3
OfCUpo8HqHgUsjc0udNOdkog3fA9c/RdF2qu8iT9XuIi/jRGZ9bVYgXCUEUSfbze
DFK3mIGqJN7+xciNF00L39+FxKeFycfOruQlzdUB7XV5MhMmf1FG7Z65UCAF4Zep
f1JipC2gnWazI0YU2AZglMcrLo7+L2Filpgjds2gqD7sHU43FBLhdexFOgcuFT5r
UDIULImlT2ANIlCweJctVsUwgXX01p3VDSj3ppVGTJn2WFna1vJlmMPVb9jWHKar
ZiwqvKJXt+ivjsJ1f+dKHNcAzZyD4P9zQn+o4XiDY/nI7S6VNEd1Zohsx8rU+dmc
/ecshf3cqMn2AFnXibTcsl+p32VkJN3OhfT5dIg25S0oCrKFgKzMtSE+OmWk4wQy
joYX6kKt9VFGeLlPMQQDAXL5toUmPwHMdkHf3v+rSLlPkrprjJ7k4GnKkykp+4WJ
7CErHMXlVFxTtuAfYnnJOV+VzofbL56AMPnP1kHyIOTspnUhg4U6TM6I3NxAMiY+
MhB5/bpyqABv/HyyJuzABgXNMq/CR2V4E3ittH7PHY333jzP+9wvasenujgOR7qr
TSTYBm6QWzyuRLJarNbDFtDi4DtulAP8SRlmIr35pAeFYFCftEJcNkAlUrGAXKru
ahwf1eB75UOeVg21aUVWMfZ1j1q/QVyP82m2NMST/YfRklD2Oo4eO5mfqAyNe8Cc
agqNl5dKNLKRh7RoMGk6sItJSLIHS7YbTNhNSAT7eEARclnLQzqVbb7W8OJ+kND/
yzfWuQ0/lQ7LGCcKQMR7S+AqTga5tyzKepKeqK/XUuzD11OzgajIRUb14FSSMTnF
SrC5fJSY53/vOK/H+cXu0ht1NprONIeG13YbYDwMHVPBzQ7g5sfkC1in/aB1D0AZ
HvlVEz7aJJS5U3QExZBWxOQidiGOOv3W9gGWhfvgS1GfOjzkfFemGcw0R/sYleYD
wJkFCjl3n1q9PFlHR7tnUwSmPz6qvOCobk0uiTAmWS5UYoOZZkefqVP0aUFQIZZd
rV4FUWq2GfbQ31DCV1ccvxat0wbQ0YhGjx3GIQuc1i1YAyFmXtx63W0vxTZuECA/
xM/7bZifx8fS3va9Ml2N0QxplHbMd9Stqi2+8hcbggX1iGtEIw25ppf3ZgejDxkR
TOPEF0SWnuj/GoDzHIGnDdbLQ01AFY4yvzHTRAUeCEUqY9nuhgCL4O2ji8zMlrBa
WdtKNxWpCP6juoDIjU5K87DNXvMgfX0xxrRvJSajaKtrnZ7y3GlhaJ2f9YpBA3gQ
goTtlBpOy/xlXGo7AF1reiVj4a3ciBz/mQ0afBruUoHboExHyP3RBXbdboYrG2yh
W/PwtDzrdFQkWBj5yoATsxK/FyuGuf+AbYczjsF1FCVkfc9gKRr5XtUzB0aAsO+8
tlqAKST+JSrizPbUmGDpxd7QG2XXTLXOowfkp2Va4r4IVrOzVdfhGuwRcyrVuVlQ
Vw1rWVhMgxyjOxzP660gauVCLpXxSV2wv0k7qFcjY+KOaD7UUtAPjHvQMeOve51n
fenT9+5Z167WL3NzdWZpEDsJZ9/ztCSgu3XBZjaHTBFxqWLBnaQoSQM4/hYfDLez
fRcVa5nvh6FqGlUHGUzXDgmsewS5SS5ZrDEQv6bJxlPdESgG74Z7K9vuyjhSEuHG
iX1+K8CxnKtz+o8mlwyTPYsPEUIFtUf1eJa8wVAgbOP69yZUcB9gTvAGLvzAVVoK
9TwpgG5k0NnNhyovmJAafuw2m94Dd+py/YM61a47KwTPQspEZyfUlx/2GegE4sC6
5ZmWU2m2v/UGUiOxrEcX9l176vTXWjLdlSlvSUtxnCciMjeP2xaVfW6iE7cGcBnH
kHRQsMmzKz2aMcXpJeIkK7lzPWs+mJjwc8k0faaQ1OinMLcZcfcZ8kUrQMWk5Pai
8y+QXUIJ7P7aeenUzIm9IjcNnCOieHoE1X8Dz859gysSPIjtFX67ZBJIxb85V+yn
wG2TrkCYq3XFGFavzEFXewrjwJovA/5NhQxg+LsZgt7lOn/3uapxUZvFJ9P6OnE4
X1+yWsJqzLIAH+S+3SyZZuJRtjz5P+84co1EcEm2FW6dwAhevqDVOcAjbL4Gmu1V
oqjopGZKtRRsrYm2zXVDaKtWXT+Nie9U+idhKokPl8Xb3vgjf3KWAGTN3IeZN6bl
MjpX3bgauXR10YWWu6rl+cHuHODsJ5sMMXGHgiC5g5joi5rEi2fFseOVTFXKYBAJ
BtVszs/quSnhRVKXyYnBi5kDT8tIGMv0P3BhygI6hatr0+ueRyClVBpiYfAJXZ3x
uB9/TRBEdHiZiJE7PGlug7UacsgvIRv5D20WEc93b7RPO+0s/5CvCgZEyd1vf/G1
seW+gVPXQa9btwqRu/4TiHAuqKK7zKoOC/pE8ZhwrZ6BHVwfm1ETn4a/QERdgF0Y
xAXhbSi372iJeydoHvzd2i1BmGVmPfU1LCx8VLYGO8CdB2/cW+cJVtl1Ub3lsF/k
m54KLnBcswmwu1Dw9X67m6MevFSatvEt5Yiu0fbWnTNS2EhB/v1P5y5oFF/837Cg
W5qU52MASAcyTwGd4nwvz7X05p+Kdn6CFFColgB6yi57Ic5nJrSIc+L2pq+TuAEP
fXrmKxSudq/MN3Z0ipBidp7yI1wm9aHKjbfAP41goNbowA0mf1gqMUzP2/d6/DVs
Hwo5dDaee1RNnORcnD4/My9at1L4de3vdFJhYWq2haAF+w0W8pmJwq9j42pwUjNX
dHNHVpYE9uydDFXvQ1p9sAsP7b5km++gv8SO5rpaiKPG3L7hop7HqQUr+QGoshxD
KJ1Twaa/fUn4Dvw4ZhUxFbJX40AW33IIBBRqKJjFgh+CN58DRz8TIRXwdUGMc0fU
ZjMzVVnxQPyFM7g6Ow7Texx7FGXA4zbL13DY7qQUo7ZRSxwqKjkN1kfOkEIwA4y2
KZcb3OXwPCcne2DTWDOFg6GagghrTe1pJ8rWTxYDfNOJWJna5kw6BLfUgj/GMl2S
+20/a2/uEBLLnYI8kUBcEEzkhg2Yc1K3zB1T7jaEng0l9vkns7ju1iVQwn2Z6/ws
rligrXOJmqEokGqgrIOb9MA44/JS7dWUuaAjWkRtz1w+vlPkUFttnIgGi68yCSTJ
Ljttxjn7xW44kMWJNZxoaMQPHXBt5mZR02x9I38Yexn8Dd9bIUsnFMfFFRo1P00+
5M0O1ZoGw0V6Z0w2DtCEJZbuuQTICYxSG0YXIaKTTwfQjktm3BkhS6wfFOqZhthU
K66oqaCwsXPdxvQOPyg8OhtZEqyvOjy/R/b2MtblgI4H+TFDpfzLh7678JZwkqfs
xY3XSeMsz3ZHkusHbg/haFk2M0kfZ2hSIXYtGEm5+PPis+9mTpTxq1/xQ24yOG84
0Nj18rMc/+QixG6TM647/jTThelvyIumdlM7dC0dAylnkXOlYj0bz7pHA+E+hi1t
Y8bdzYbq1KThrAUqHgAkxN/6+pzb6Nugl6hr8f+wY3JkdWMzEuaJ1XFSVUXlgLJF
ReJ/65u84AIxB21WYtkMqXxv0GLBvHtmQ3XH/mdSLVMNXbk+bC1WX1GTnhf2ZWlw
V/VCNF1yKu+BeIAHKQAWZ+yqQgrTzxPhjo4jaaPSiejAaDOxTqLILNMnj1GZdMb+
gy1lpTWLLOB+O83EoHt2+QVvoEUMAxqfXPlU+j8CXNFnHYLXTma1NLHpasLUkgUV
y+FCBcNF8u4z5kXG6/uIfdN6I7xdszydJgqOH/0KrLciL0YmLMOjCGbM+fcQoRFg
4DmrVDNOIbe17O1vBtfyAw4SENVBdY6sJDCpLNopXuD8es9UIsf1m+AbOdBLV/05
tDkiHw5grW6TcXrrjN60ELkDNFeNrF4mn4Tf2LK1Mqp4nzDsV/e7ul9XkwPcllwf
B9aVUt7uO/TLCo/by7wgxviHRED6IJj87pGsuUKLVd9I0NSfoAENvTUXj2ysUZ17
gM6wxJWpFzVrmeXzmiCQX+xWTVC3t1l2N9CQK7tYX/u7321ORMHwICnW0FMkm7n9
dnVsS7IiaHI6PDxS+iyiKITm9xWUFnaYBhcwHlOfpQgtgRBbUythvbdDgfA9Io21
LtSPRbb0kFyx6Wpia4qyY6oFXtGXuq6P/UWhPcmr351QWgh3A6UjE5jXkzkUJSGe
vGnYMObLjbdVO+5pU/NhjV+Vu1WJeEqvw3YaTgAhSmYJjPyB2t/IkXLmBczB6VUl
uGtpvSiNjFymCdE8kbB5+BqdqKsv0vbQt1SnrPp1gfttHyplb82inh2NeDHTM/Yj
KFG11I7gpM6OyFhJ4VbMVVnk9+K8gp+N0zv3TStEAZzpWEzpd8qTgvdtgNn/Eoge
GWiySSSUPUMCtVQTlxB1HaeNT3LqobCIBKuRuy/ei+yS2Mx+tSGbWgDs/YYTjxcL
KReLxduuQYNcEu1trVE+voa++Ck4vmg7jsc1ThZNi/dXdLwMyNQylyvd2+rjPJYG
tvFlKxEgMOzRta29vhgVUhL0o3I9jgIGmPJXh+hh0tMooM+qZMBfoiNeSfVSmiwc
aAlzBFGB+Uw6rU/sBRkoh6YVr4LSIKslVd79k3/zG4PvVhg4364AI+8PzYbSckmh
VR3fEATvDOHt9WYuDSoG1UgqUa95j/8DCkwLEaJn26JTVHVa+zwoQvh2VQg4FZBL
TlTwIgp+3hJdmzZNMrYBBAZfXO8upAfNKg+DUEOrbgppaX+MPUY+a/NqBnDZzrto
gAl5++0PxKZXZ4jPrgAaUvSf+b15cBW4H/x0EqOaaZcKFiDZiEDzoFkbhl0/eO16
yZ5azOQSL4XzpDV4XmaDYkdvKLzgSwLCK5z5LtAdOnTxU8yZ31M7KVK6memv3QP1
L4d9MmiGXw4RF3esR0rtUdlr2D6+VEvFaZA+a8coxafnjqeHrPjcUJAgCCY6TpzE
MLlD8TIN5Zq1WARp7Qv3+GNDpDixkckcu97+5fiJM7DtCcdQL2eHSsFiadNkEY1n
+fHprx9O9IH7fKCb8cOPHjXhbdIoMtrHIJ2iDfJ9Iq/xszuGHvvRpVgMqIlbvpYY
nvytz061UYMUr2tF9ztPiKvCgFofNK+QXXXmBP/tW6lqhcdJlSu4s1G61heqHNNh
KNQ9pIVfAxMhVLb+z2wxor4G7uXKMF4ARsisXCTEqBWB14N6dV/5S5pseSlrxGCC
vd44BFsOE8Gj9vzaoYYcnu3zYObfinGhh8YbPxFWOHpBpQc2/5DAuDIshDMhz0N0
+UttdkfbADGs0jcOWU+2vcn6xSFV9XcMLFximgw4h6HD/Dpk34p3u5j0K85iq24g
TNiO2dnIvSoHl5lR7I9l1s0NHn41zAu4PZxW/+YB0tmelfiNDjYsVPl3hFWJP15w
swQBG4inVY0nKuE3BJ73JuMq/kyvJ/7szIoAf55C+PRRQB/TPEnKtespHOr7ONdl
k5ejD5hZf8d7kSIr027l3pzIybDJ5LdS6wOqmrILbmxsmhjVrK4obqvTVh9M7xhj
ukSM6SUn/8j8LUrz3QvkgvnDFFSbcSJX3/q84/Mgc4p5eKJ/f8HF1n9+hfedD9jM
DWnBjxSUYRO0O1FlVy5GNUb0+uLbM/tqwUpMeWlrSXoQvi96tMC+kw32SThd5RKx
EHvsDrLUAizF6Z+tLZDyClm9FB4FYSTtuLVWmXlHDT/yyAf5k45pTp8AY3U6GrWr
T2NcoG65e2/udUxREYQKFRMRpOdSTRiWWT8fpzcj7JUT70RWKlWZT3JV0C7b3xVF
rEDXP/xFp+evM5GctTEQovBWzEYh7jPsaelvso2I+LBnk5GPLD02LwvWtuqcqg5B
8vHWxteggOb0C0FOcLCAU14MOBwfXikaF13DTqKvBJKAdScOsO1w2AOcIUOw40q2
Hh3EII54vbClDSrKYKNN5bmU9CrR3vToI2cZpT+fFLKH6PF0+VCDXHBeVM0iWJgg
Tl+8qIvzKuqpmRHrol1nW34ocpaUEril1eq+8G8dSoN1GrYI0lEdSneEM2K7PhFd
VSVXUAFYJNX1jko/o2hoDFYFK8dYAtdfEgl/a9TbdoHJJs4KSJhkjWsz4hej8ooV
XRFEyvjALFg1W9d1sGk92MAao/yNHMIaGvao1/KTnE4qfwj6lcb1qPnjalHxFNXI
mknW33QQGiitnDYHO7AhAgEfweDkBsYrH1K5vYac6wwzzyGGOzcRbR6fHYdOqqG1
rh2TYX7sERZIHiuzvQGU5AVGRG1GrnvM+I+hhAqVKkE24X9nOKVG+spegrEfZE6R
rN7BpC2gWgXcJZpN6sOs4xbVAXs1/eXYTIUqSPJYeYTUo1kRK43RolCf8Eu7sOBm
X5qeL+G7w6fG6zBlGFI7n5Y9dUHIRjrVkRA1BExupe4Sy+bXADjfFAvxTRu+qa3e
s4QtKmD34iIFbxv34e6qKTgXS70GItWq4lA8i/b3I0QW22FSqHMMPaE7FbhemsDG
bVYtev+h4Ck1fWG75IIIFT/7WFlVPqaiQ+Nl/wWdAUEe7IcCYtKKety/1lgsD0/9
prz0mgom+Vgod7Ru9c8UctO5oeulDOWQUknPpRLwjuE/tABnUnNz984CT/uMfTeS
WjaMYtbo8yOhboBelIJrDM0patOD9UKtWas7dW6mMvREntUTBYjTHgQhFlooVCv5
sVp/chZPZnrNOzMyR3v3QD5PS0IS9bh2HFgJ4skdqj6pw5MxuCxlQGAaYDqR/jOg
vk+GqarwXvyh7zN0jtFptW/jYzjjnfu8Qzfc1YTmTvlDFfcsumha3tIRPdMujNRt
aoYn+o67eNpjw5Re19Vg2KSyA+eNqtmihc6g35Qkef/5DdYGI8kbVU/CVy7E2Xc0
gfWj19d8BbZ9zlkFM7cnfMYvuMUAUSRdNsS+G/KhQhOmPie1WfdTTpsyDjkVaERu
J334NFGF4F0g5tgIo7HnT4GWkNgy6SpGGRJPnFU6fBAubdkqTJymzHkf1p+zaj8h
nDhLDLsYe9a7rrl0Jqs6zW8aK0wG7HiCYsWJVkS0EWAlc7fodV51FjUvpMh/e0Mj
+4wy2LHLguVO/gWHZWPXXNATHvVJMuvO6tfh6P8gbKsRPegaW5xA2xcTEShLw+rS
kGmCEnDjxhRJXHSPuZ6lcidufkVaOs1w+0pDIla9eZ0UCkycmdRL6ZT1n2nsffKN
5V9eOdAXVdq7V2ZUY4JiiztDBHMXaopVcXKhzicWNnRl5hhmT9gCqidkTBP+2uFp
YpMM+qShZMytBun1JpcNLCMFwEaMdh0+eIecZR0YsSsetfW5zowKBS76v+wPS2ai
TRrVNg7EJwK/TaIxyEZ8IUsYlKqCXgPgSrECLJcGwavyxUGMTYqVAVmPnSlSR5KJ
ckNRtSYDsbTVJDqvyi5SDTZaVZ0NPJFMMDU3gED4iimwbOA9dkzeC6HlhceMbvUY
mR8a1YY2ILjliwK+r/8FkF0/c04KVos0JsUwogKzDzYZYFiHKsx1ufqLktyiyFda
Kr4W4P+oYl9lrc85R0ke+FEXt5b+fzYMw8AQQHd7FDXgWuGeMlfIFdnRD/OFLNFO
LA4TqY9qaJWlD+EjfaVP7vFxiqjr0vLevxt1/kws2jDAy6Jr+lH19bR+IgPjuSwM
rGvuD0Nyc4ZuYDQmFSfOX3Y4Dc0OyUATFAXJ615RvUBoAfEYRufnkShtJzAIUBG+
ZsuuCQ/FjAa75pkCLy9qYTMzg49JbKGLuFvvDXlfASosSuO9IwdgZJZKUZzai6SD
XisBg31SBKiPrPSi/us39+q0GyAOtcNuCaxxgl4PrE0qWaLCwzor0/uWXGXJfSR/
98SRhFbP8+XPrHK6Kf0cGWv4jgYahp71UvEF36HCR4xkCK+G0zRB8N2pIYw5nQd1
jTKiycT1l/KcqwTnxVNuSM4rK5oQ2dU565ubkrm3x3Dn4wsSVKuRXe0D35MP7zko
wzdZ3T4QsKFpf8mSlEOAl9sB+6cXG9xgR+5PENzXBHMRximHFQ/CxDkxAx8F7VUw
9zMtMkRtQ+DXmR1HpUoja8PgjxHl/8/kZN3vTV+CkQZI3FQuEi5t5o2SLuvSHQMg
GCXHVtl1pt+3G/54W1M6kiXJn2/i2fFQ8KqzRNVEus3E77fja+prRLT1E28vVQtU
m6B9SZRRk4mfFR9oiup4nzxtfNFXfWDiCxn6VsAt7DXmjAs7Uru3y9hjw/Yr6Nb0
HYE05wFzM2Fy7y93W/rHbzmWSmpfmpTK7wLkXkKZZidVEsbPV0PFK2NsexMJBBlh
Ud1HYaVaUvU302GQzNikn616yp6eEiKCEdY+x8iC8i5/o3yzISP3hvJP1F7spLK0
QYgpK3R0+wECjRcmt0lhuqKHgdBcAm17CrIcWxHpy3vnku1Et0iyd056FwvEqiSx
/CcTxM7iF2d54TW9smJSm3NeOGQ7e2Woo+Y1WLm7H89egGCIl/2UiQ9k9xGd+gmz
1S5uS0wwDOeiorAn5Li7uYbXXYsrDODaNzEFIHdtRWVlrTCAZFyK4z4CxIPwRmE9
qtbnPkuc6rpfHA5w1CHIUS2PoaJSPnhXcTs81biO4/VLXhbtvXy0LY3FuzG8woHd
TSECSQ1VMKmHoUe8oKiZvQvuiUEFZyY8CRFANGfkLEYze+LqFApc3XQs33VMGnPx
28kEAPrm+pjzJ7eqfUwHcGNHTMRJHaDVRtN1WhPHsriOajTd4XwRhZyfl/5Yr+7p
E1OCub9WvX2D596mjZ2EIfwNkuidtI7nwnv9kTAQCq5vdeUhpHR5SXAEi432/S9k
/m1kw1PpT1+pYV8nEHUMPWwSu/Ziyx9zMmO/7PYP/pxxTcsjm/GvSNBIf6MXEWnc
5Yx8ihjga2Sj6LDLuvgHgaMTIYrJBzVC/VVviF/n29mywfewimyala1mTnO7Y0Bx
pXrWBrY+gWLS4H3cx/WVtAAVtcKmLJ1Tk8UD5+aBW5pqm95sPTuT66aOqWslM9Dl
nXVZ6u9SgCzbqt8Vj/URW8kpXtBhKpLhs3OEzWLWOyVUzf4AA6SFT96iSIl8XUox
TaA4wgsYkY2p0PTK1oy3fETGM6dmnP5LOqNSrcHY4LhuXH09IWnHVJINuQWREZkm
C5zMnrQx3Ot1dbHv3cf7D+pBO/lBL9OUScy5A4yDywQA0NDjYxK5tXJF5A4ibWxj
ppIGpDeQB3iA8FUrvpmhmBQ9PxeLgTUaTVCqO9+VDC1jU1XUIbV7PAtAQVZUdBNH
FIp4kPIWajN9nne4HD90cbT38f4nZvQESz/TZTrbNlOMsRLZC+2wu7l7ZqZ/J/zi
zX8LnwISwbKanHkpwClSVQAD29swGbmjLCb0O9a1h0rjA92FT5pfU+BEoySL8Old
6p7HQtXN+wVTsz9oYBb3jV2H2fI6qDhX3M5ekuRVrR8MW6jyXeV2dsCWKSs6KYqu
eaMF9q219QSiuZrDHKBIw7l3cPrSm95D2tZvNe6SKc2mD50uLaPP6kpG4o2iXVdM
G+fRrBXru4+8aCesJ7nsyTbXxPFVo1p2DFdfyuJEGjlePHQzdScnLZDICEjYYWe+
rO7k+X4gQBPhsJPuGlJWnUuSYka810oBUwTnoRf54v1qddYqESsp/7z/mQwV8x00
T15KytZEka5CGMCUioXiSV6fDB4OMulnozb3tOMaArWMm9zfJwGHiveKdLYER1lA
VNn41vjNxDkYo1tUWbVLrTVVmus9jDuuDCuXLc256h4MwHGL+fmXXsUXe07wvqI4
gCr1D19ntVukyFAnDpeKhGVTRX2sla1xowzyqypedUEkSClpxakf/8TOlYpoUfVL
TwjnH3LhcC8rGzr0dSW+vSUkEyc++Mf/XAD/37wTC3GB639YR7qtdZTtDvPp7ss0
VlRb4JPcPR2hoope5Q9c4OENTzicO+LIgUNUIJuebDLRNGvhr6Ggc7tRnl9gJyc/
0B9HTPYO+1VLiKAQSln79gW0q71bZiRKZzbG/bkVbKn3QjeqNyBFQlK4Gk+tk6ko
lzg3n7Y7LC8eqljw7gaB+dRL5TV1rgYmBpLdVxuXpAOuoyryD0B50d8oTfpgotXs
ugn4rCzqwKZMmp1/GjHfBzlxZd1owOFrv3ivOpASiqZC2DK9E794ctdNK0O2aulr
PTCzHv+7nEzqQgt7CLXi+1BcpgRifW+XdZ66Gton+r2hubFlaJSdHBqRZXhmYx25
JtrQbLUSMTamZAidnfsDF1nAkY3PpYsomPxxvoEdedoj0ArydfKda6DWAofvBeiz
dWjbIMsvfoixINcP83iABorhmaeyx96SKxgjf6lBahRVZ0IaSM+8+ZJHJFobxK4M
8eFrm/tblq6RaUJ7HC30Rwpn8sWC8Z3h0I2PAl1eUpzNFGWQTBl80SJJdMAQabog
z3eOLzAmQ5H8UfWjQDqpEp9WJm1wRFpLPItYfJBPxZxtjQF5MLQhBI8Msq/wG+oO
kps670yujlIFIWYX9Vnnk8wQvM9yiUHRIAkyZz9ZoDNwDch8JEBU+r6s0Z6YuWAc
fErGCirGzZZHJMrQlSHOidT+JNio2CxcrdPR/1kkzj4QO6V8jqamtxn6XH1fNZO6
ayzvlOYxLdZqg80tlVCrlmhQyAzZifpRWvmkGVyCHEnTYXs9gehEgSwrDpxg2oYK
V4sizCFuFty/X17MqJ/UvFGUzDztyPEaiA1sxNO78Zb4wqHuOPPf8EbzeBug7HYL
YMX1u3/mSPh/lpFlql5rvp/EGclAVYxc+6OGZ/kIMyyPdlXPDRbXJ4pm+BitTHAk
eHLX5l4dFiVhtwORPVe0jeQvrzrxY7GacvO4X4M15jhL+8hLM5sUbWgDjVZ2RKzi
Q+D749KPYDcQHdlMMcvV+ru7X5qfALh2w6vgc0Pf3JeBR2aAQ63UYVjJsZHPyWT9
itBa2R+ESO/D1uqRN5juAWhHZentfmsxxmBLPRTeAc7DC/p6qLzcs7FWLBQ04q3A
5Q2GwpaqwFNy86TDKy1f2jhPNwOtY01WxEHDHKx6KAkFThGQ59pFiWvaDF9oYSbc
E9zJXWXeOtuxqeM6gqhiLovA8puMfeSK8XKQRxmX3mt9Zx32X4YWDz+z9CTQBNxR
xBTQ9JUf3TqD5aZjdBenVdXSN/E0BlJ1aPf9TE5t+Vdi2kmtZNr3Pb1za0xT62H5
giujrZbQkc1CG6HpSu7n1hsaCf5YOvElTzyCnbCbU818iqWU4F/okOCUElSXc4kY
qT6na9sjyKgyGvhjtC2Im1PCFwqlnCnlzjbSmzI07mtnARP3owkHfYZVddm75Zd0
zc15xDVylS7uHr0yasbtSlPSOLmkxmCPZSYxrvR9qypkD16PsG85FlWaIzE1BM7X
zRsokZf420Imh8vDKpcz9iHBCLixymTyuP4OPlLnO7YPCvUh+iEVsrj2q+xplObu
VrB2mjZTgHH0ylRxf+qQsQzk5BEuFvDfHq6+FEASA1HvoPQRzzBq7CAr+JPKjGpo
QS9tvkzrYPgReSOgYkGimls1bIp5nlddhWPz4RyNK34bPEmAAz3A5R0yIK4isSXv
zJMOSCoBvvDg/IJcX/30IAv0GMYoKhpmlqpD81QDbqUj/FUi6ViIaoPJ/ZXuc6al
lyUyoR8reSRPb0pDwSGWTZJ15SD7LiDYfd2IQwy614CjKV4tUi1PIB4uGKgAVtEg
uY26vQ1VCM+wSdhLypqJ/59hD/Pw35Qh9I6NXL5fLRatwv0qREZBMFUJk7aVWKQG
Ipwd/+yBlekrEgS+yt4lMzvHUgloWpCfwWVKRt4P0Vbvhffj7TGcy7h0mAcmhj16
lIBsPin1XXMbWN1PzbIDO0beBNtxyb/S/NstFeg75RAZ+Z2TO0zjmW39m2qG1GgX
Rov6uGLGaIxNGJ0PQoZHO3iskzx6GAlH6C9y9QpilSpNLIO1G3kLH560jlSE12RR
HQQxLoGLlr4oS77m0+01LHVY3R9z+25oF/GeLHcP+IRygVXmt/AKg2pNyZYfbgHv
PnfOIGtMONaMUdRHruFlWiuSTpj3PLkHja8XrwlBbOjaM+CF/LvhlUBwIqA898Bk
GgDZqlkHT6a0duGdnLmYEfkPiLodxovH6y2Etz2zMlyJ+w5WdK7OmOir8WcUS2qh
Tvg5ola9mBZBPH9/n2Ejy/8q1B/vXwKPZUdJr1Ex3m0V7wryKE6eIDJ+KSvyiDeW
xn3X5r4RIXLDXZdeZCa0on9KGtGlZLrf8+q2Gn9EUus5loQng4Xt0EDQYvnolYiS
SMpzBoRcEYr3foG0jBOhYTD1lm7k+a0w+WDHIiCblRGs9HLSR2+opqD1o4BmIP2h
FnfAP/5xJlrdJptHpNl2XaffJjFVQCMPdcJ6xXFrqe9Ug8Tpb5UbwXpI+r6NMwBT
GKczbbAHc4pvLwY+g5wXStqBj+x0a14oaIWUrlzD3W/30rvnjeLzvd8Kmt+264+5
kvX6H3tXlNXqCP8pHoGONT7fwBpfdFOD1+Ox4vSLA/PQoCmiRw/wC8F5iG13CN+G
P6NQQY90HLeSxjZeH+A92kkJb5Ky+kYEgKL1BpfEZoxu8r8XN7pilQhkO7nqnPP/
bmzDEaPn47WAX2IE6ykUoCNTYMEeqPD06+o4L0VdA/dx5X1Uc/lqFlG2VqT2W5lL
VoDJMRkgWxw2ly1Q8jvFB+wldVGo5zKOihhAm4Ln8a0GOQdxWFqP0vmpvG9jPaga
dzxLQfkbnWByFFrH3+ErKMGU5/7urvNcDhs9MB5fU9gxCwozQZuXGKjvQbkx3qVw
c3foBcQXdE45kZdJ8O8d1+vouGk8Vv8TEGNoJO35MrjvLkSBVRisFNgCmHMeqg79
p5d20L7PBsOGNXj0AbuwPdvJlIBofh1WUkpHMfYe0ppNu2aJ2eJm0xRdcoB1/x0+
GksTQfs7tk2OvjS/mxp9sfNooaSSzLUA8cMmAtEdNkXf9BhDSEq2AHYTbVjXnajL
mzk9UOg9CcADQMaNjbZCtvwH3jNojajKHXCvXOzA8p6BdEdn1tDiuTnDKuYjRMI0
K4yfBTgO2oDYuoPx1aL0rp/85oQyZL5wa8cPcj+FYfash2tnSHJhGTvZuQqG9MZR
Isu9NMqHHw811ZK0dlqRDGUs95k0eWB+sFLWWjDEuc6cClHxAWmDZFM7HD8nYqWG
WUqGb15zyiJ/JL86jm4fx9cwPPTigode8i33X1qMXBRa4gY/eoCDjzqvLHBiePt7
Kv46FaQzhyGy+ndPxAt/fIm4Hi1Cjxaule/9PdDytaVfgl7LLO88ADrzOMpXrqmi
mMBRXOKrINoBUq87edoD+Le8WvYy7yTv+tIgr9KX64+mEoTGp/cFGHBWRh13dVou
lOZUj62uPxWbp5a+6nOM/t0na505sHaxAs+X2YDHkes/RFxt5EbX+WQiCB6VQd+b
Ai0JEXC7sguVKRAX/JKPMFvVUcuawarEez0wU6FnKLWKRiqIBX7cimkvia21kvcc
EY9jzQiQDAGXweaFPvaGbYrittRlG137EXAcInmtKeeUVjsL7eeWsLwL+Sl71vJ7
eYcLkixuMCsXtDpg7FJhGlYwrl6oP9d+cf4ztkEzUEjKzcONxVBGK3yL2NxiRCZf
X1qq8tyeJ2GenbxRouMxAn24rLDok8UEO55K8laOYruy67kGuVR37GmUqM5hzZI0
8XD3NXEaJvI+i5Q1MnkaESkNcze1dAMqfk9oAvB8XSUss+5ae2D64gAHriYwowtN
xb08fK52VAJ6lPPKXotxn5Eg+NsxulKnGV+9D9HS8nqS6UArHR7An4Qyvtv0CHq2
f3Fi0b/ktQ++Zd+nPv3+Bsf8k/L1wzmWCem+RnRWeQbI9Fc0y+RoIyH/QU1xoAfv
AMJHexk6pVk5Um2ID4zw6iUT/LmHaZcK96Udve+dEkEIC1DoybxzSrL0mkX7FNSX
lhPOsfLlAQAywgmBqId1/SPe8Q8gPLHAgzoohtWsJSPW4WhInvrdtot7yWrmX2ym
RBjquft6P9EbQafj+OiImhcq6GwIGQOU9mBnbwA5riYRK4zvdkpgYE8UK/ObghxG
pNl6jwhXf5hBNswYqlCnmZYFqqd6IfWxynWWy+OihA/olAo+gG2suEn+9Wu2vou5
xcdamxE3d0G4uh09StcUHQS2MLRFRJIVXuni+jTdbPbBQ3uVVlsC8rbN54ZAsAg/
9X8SlZMLP23+9v0rC5T1rnh79xyJceVEw67S4eIZtBaFdNAD+SwxGq/WTBxakbKd
/gASBF4HDKzRwqUnM7tEB0QlxmjHA4jCIJ1EsaeNQWQeAbRNllhrNq2NjeBh03Wk
UE0HPe+16v4b/VDfbZxiM/uKG7IEaUTDRLYVknRhZLqtjBOWR+lPqWOaudOYTsEA
L3Z9mViXU/n/JNA7aC18ljIxYA7B+5/eQVyPC66uusFVAwMk6cjbsQPyQGz5kNsw
iXFMlfy7/HEiEbGJ83LiA9r9GVk7mvN0x/HJc0tB+FVd0irGy4+Ed/DAXTIaVWkN
fZSw2VIN5KrXv7QGVWaHNk5PQYm1iSfRDejfHgttjZh+lwp3eaCW96G2kbaFenaw
czKoJ3ZAYxHGMdpr4iPJk6A/eBlWEJyTl4kku+zTArlb8xIOdvpAUM9JQ1QbWxqj
PCPhtCDxRJKwslWQ7Hnw9rBKrLV5bfy5LnzWAkpLjJ3B0uIfCeWpz7cMXtRbJZJd
Bk32DM1k29YB9KZVaExYitTsZulsFCC+FzCUVDy2LgEQ7GBTsxsjNTwDpXULck3B
FZECJaASRSeohaQmmSqQvo6O0CXfyBAst+cFukd6TN0mpKUN3XY1yJhZHSrjvk7/
/7+7RO1cBk/cteztSRrZgpI0a0/k0ZCrTSpsHRJ6CgVaPYRoKEXvp2ffqrG22Zw2
1XtRWQUHUpEeEZLUduW8F935BYcFzvxGHCxws+LhAEZtJkJXYPIphVDhPorfbTpd
GMGMio0NESuHmhG9+gWDZCLvt02dZOxphoNh675GkZ4=
`protect END_PROTECTED
