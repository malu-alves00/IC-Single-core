`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3dtbR0268VWAANLeM5o4y2BIMBCZbmJJLhjIRIHPR4ouHhu4AWXv+4Mqj529kbvw
wcxa8YhpE2imYJ7XCxCF4pJTeXDgmdTmrQeehhe3ECV3JwTefuxb78e5lV/QH8wf
Uc8+jVa0oosdU1UlVu4qruFDycWdKElw+I4Puj5h+uCxkmHwNlAGuAIukUdn2FEX
2nzq1kisNs/4q1UfWJUtOCZWxw+lFUCfNtNQhlRHSDiOAP8AZr3lh4Gol0NpbibR
IZxCVD5NtcTUPPSmcIT6vGs4yZXMtiCl+FMAlASIsur5YokdyD9RY5RK7Pvsz69F
B3Y9AmBW2CjQhyK+OrpANom4AKwnbYK7Y1BLk18bM9l77FaSfXNSAyuUO7hdGOy0
o8w9EmFNuFlV3HhV6auo+4sm1SbRphZ1Rc5pMjCfqIcxjUey+vJQ3RmomH5wdcVa
/yCrVzk8m1iaOM3gbq/kOz21tKXt4nZG5nPnKEsAQ9mNyv2xZkCVkQACiPsA/QAO
lli7gI2cF9/oW8VNgsRLVbaG/DgwLC9ELaTLxX5ubnpITPGu2/fZzc2vLhMXOz6+
Z40BIu4eE0EPHn3JBoi9y5mzz4UwbUByNjdxK9oMzqVm4toHex5WnpEOA4LjZS2a
usvPoxB27btzzWDTnTEfwO2UnxwFYqQ5dpc2iwTANrQRhzwuXWFy57b/jMfdpREE
8rWOO/ktrAVtd/O573FGdEr1LWZDcHMapCxeVcosr/mH+BBnNg3ofgk+bqfHgMhZ
opJIuWVE90CPvLcPKGhbnX/jFro0Rd1DsdnWR7VhDNSN4xtIxWs21OyaBepavtIr
`protect END_PROTECTED
