`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Y+PlhJdhQ2M6Z45Fzmtrswwpe7sw62VLFVmTUYcA1Ti+mRi4AolRtD50KLvrHXeB
Rvm4kVn2VHk5mNZBzNv+uY8ySovY265dgQniOJKV2JE7l6UhPfBy8dkZBjXE61Za
1lSa2z/tSu00P3YopLxsNM1OCXQwnL1rxMZR/vI6qzv3ICmOBeBjvZHpZBtUSwve
+LK9rskCIhV23S4z/Fd6S65HefgXj5UDndLgjRK+3G2hDJEM6NnfOtSnc1Nup1wT
jRUqNOPJWlE9nOvIAbY4TY+6eRRSBfXrJWo2kpAKJwOhB5YIsx3+RtPUNRfn3zAN
dAYVl+nYgeBmztr6Snx6ppvzTjtbm4RLaPQ7WL1eL/A6Aekwxn3BU08gh4dy2NtX
GC93A2kxHOIgffbDF3YPtkGh8GwduerbSgZsaFuy8R+248QjnudaDJazPcMmw1Hi
WTWPGyBD1yBq5MDW/2OPCa8k2n/6phawHdXFWr28nld/lKZxYJ/5lb5ip6Np7ob/
VbHzI8uwfiJqi88L2C9IXyROMN+uZ4MNluKIeNowfPEqYTBOT+STbOan+WMv/ws1
+T8Ei3GxOCLf3ERa86UFFw==
`protect END_PROTECTED
