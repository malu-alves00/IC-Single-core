`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yMR09vdi+/A6ofbvzPs674ge25aQ49ZKnhXCHV1ITUzeEx4BkEHBJz60kAdaijCS
e8/+Ut+TVfOj4YNhWF39t9Z47GFQr/L7327pjzDwAa0FT6P8EYSR80pGHABlqFkW
nuIwfJZvpRasT7kzLg9IMT6BxTATS5Eu8R/NpjUB8mMoJDTZbca+uhrluNQ/wNkt
/WwNVlv+Q0eAbDcsTwJNeiVGmwrENjNMMk2kA4VUfSDUaG/8tIkCbG6AvabKpYne
Phx0SBmiH4UFVnZbF5QKKwBCaGZMxJ/qstFXYtStc2EegyEmOPMyS8ravrMUqawD
aDg15HS/+J4PL6j+lLEwtBB49sw5NfIXvaETCvf0IsS1UMQKMUTgvKRzuEiEUpDP
NAlRFIhMX9W6cEOFeIbcyQ==
`protect END_PROTECTED
