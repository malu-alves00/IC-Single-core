`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RoJE+//AdWWgIJwLKRbEK0guiwp4ucUS4sC5bpwdzhzkKgUe/tijBcdyPPElm4Kx
WpDOs3f4asV56UteUtrSm+lKZ0xOf7VInCEatHJL9j2YK2Cv16lUQs5U5Uls7dil
FWdpKsMuA8ZMZffuCOqOr5E+fXvLypIGfDvcRJwtOYwT73SgE6ZoX0lO8x/mUtw4
i0PXzotfgF3HzmPbVcd9j6I9qE+CnhbQ4Uh13j56Kf36Mr7HZFGD1Kn1tre5vo06
/vio2fEEyXzzbdwNxEZuXRLz71UEAtO1f3Qds1msunA2f3CZFs0C8fdExQlaXfwV
rQv4Q9AzzhXOxoEuX6Tzw76e8Ny05px2xkKPvrNTpeICqJeDA0uU/lYg9Xgjej0V
7x7X7DZnWd0RJPMYmCT7IJhFQVmG2BxcUyBrJ+B6XPRERUf4EdifFPYMKb1Q9w4y
t23jRPZurvqN9v/ddvCO3wsktLEXmNO368/IBDDm6C0xDxrm6lcX3WQPJptBc3gR
IrRZ26qPU55qNhz1gf26XUYrXRXChKNBsYjruAuIoifwUxRln/DT1nFB41Ld/N3h
OV1i2cIs0cvlvI4mmhg0wDYCHWE7gHSD5eHkz+FzPlVcn5T8SvF/N1/byg3bMXs2
PXzW+bTQa/JgxFqpm1i9uYGrXRETvrIzk/yU2Jc117VAgJBYfICuytwK08vtLE54
DuE8H/jGTJgj5VW0R+6f591TJGdtVhzi6Pr86aRzelJOSWHfI0MkcDFCr5LnuT7Z
s92jRf7r0Eg8qSxopTbcLGjFqQ90K9pfGXJVZ5LHDbVwq/s7TsMGr136nj0kD0zq
urtOZPMArT4sE1wiHxRvBRzOZYhKnbfYwBddVSfjJhRuDgU7/088SssQGbmRf3og
GxasaN1NFrK/7jNGLmVzrrXGVClcDAIH2t+DUScA8OuplPw1GyY6asVMwVpXDxVQ
/RpJvgIpAc2r/tu4aW30saeMRiqyRZtF9FgXVZU0N6FAYs4wEfpHu95Sl4Y7QxfE
7e1di4rFQozBDTjxLuTq2STzuT0rWI9KZpbpyxaw9Y/Epul7FugBLvz3tXfQfg8c
19Lc08ARob6y/uAwo1O3Ns9iDQCm2Lu4kA0izF+/FG7h8ESwpNJ1UeaR+SSATibK
EBNUOuGbeKJM8lJPo6Rh9/O+JVSC4SVURO3cjEfUpp3vsZ9y464kC0J695o2OXEe
f3tunfPdasMwC2zGMTGQF2yzaRpq0GiBAetSua1CzUMe/qPBNllJFzriutvrMITq
J1d9SU59NDLc1M27qe4j0mBBK4ihDLhzkMn68/azb8J9CAvcVvfVtBmgllX+B41y
6AegNmd9PX3dYLcPQo1RikWaH9s4G/hdhNwj+2ZSzkLpb9KDmk5mQjw11LjZusDn
rNh+DDiy3pIyH31XyS3s4BPixwPajvu/82Me1BE+GbAPFtQbvRhZKjdAChzaXuFo
theUSrGB2FQjvK/Z7GI7t8PoBWIqZ3+9O4nXe74Fijt9fLRicaW8huJ3lLshByUt
g7DTzhlSWCwhowodAktF8SlbAdiDuWf7OHwAxAMTfJ34vqTBaWGC2N6aDa6jbnqs
osADhkct9zv32FrXTyhKsED3PbGkLZ4A9X2boTp6hdGAjykXWZRfb152Sjq2DC8n
`protect END_PROTECTED
