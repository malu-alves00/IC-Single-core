`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Lpw8mtc056nImJg2bYy64sF1xa/JtMOnFKh2rZLcxJrJf7Wv3FpgfQB+nVXg7d33
5OIEOP4zVw1K4v9bTvpj5/QcjCkJJjQjIPpMi4VftmqwMv/S/jtUtnmuHqDLj+50
KkSNsOZRmkaRybrYVXemfb6A5fJXw3PPLaE8mt27h3LBN+1Dyb2MES1jStPLb9NO
dmAhSeIgASMdnbHzWjxSvsoOWxoeAXCC7bV4estmDKcbOBeQBPbNyAFvvXM5x/DK
BMLgWPbsip7B/dn69y9iUqAOhsp+cMVBs+5WGuLxC//8lgY0U48Mlr06fk09xLwd
MF98WLitaGI7JEVrCwBTBmaulpsfs2N7x5iIudrj99U9M151/pA69MU8hrty77jM
tUX08/Ruz4pn5nWNmnvgmjo5BaRXuyqtxHiHOfcunRz6Bv/jXgEpnlfkVW9UuLwF
tchRMpELz4hckmtqY+TbE9AvqVQdLQgq+Q9qTe+a4Mu9KagCKjfKbkto7qDpQXzu
8ROogt4HlugerX5yPrXJiTHLxjiz8WyVjO95nme2OATYkJDlBawqJxvGQNVuGKx1
hRuxrmAQebhg1BlAjZR1GOuPHXQ+eUVCXlMA3H+7vB46b9c/tiZa1D9cMZD508BP
o7S0xAT9FuhpeP/HglMuFYLO5pDZ7ItrGvGYcNM7zH2ooJwWLSLD3YQKcXb5QfjE
GjT569/JV25Q8P0DQOvaOn9vLTozQoeogh2VpihKCZAR2JJh0ie/NK1ZOT/L686r
Ww8LODHnzNFVb24C+/x1CqsEW/CWpyHCBxnR6huBOvE4SmzROn24dCUjegyef4DW
BL39pELtBJ6TO/6F8H8tysQIwtIYoHTy2PGbb2JoX/LDySsTkf30VRskEHjV1Emw
uNISs098FAQ7hfolZOyJQ0pZLZ4AUC5256P3x1WzjYBYSgOIe8Nt+h5P0KZw7Z6y
`protect END_PROTECTED
