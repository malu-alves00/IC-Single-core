`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vn0iqpm9sLxFffWdT/A2x4JuV8GFBuHxC4c6ahmkz4UVXbyw87DluQ6U1Biy+CSB
Sd3Kw7pGlU9LBnCGhhDN8e7xbJ3aRXqxqq9h4MIbi/WLGWAmjOp0isH58c8XaeeY
Hjo2RYgY3VHsYyESz9Pt8AWBDTO5hN2bHu+hzNXhXCe/PBZau/wlE4ckJF6jCgLk
ZrXOebd8v6/yGoZojpIkrJzSw5xV1YHtMuq/olgSqsDEdLwRVc5xbR84zpd5j7bF
SYYDjV5ZksDJMlIoPEXS8ei0dGPbh9NQhZ6x5K3OzihebecZax7/mU7pbDkMN+DB
bdCyuAk/xl3cUuHuWoKgp3gv3yUIgJMRuO1LhKNnskIa0ed7+6o4zW1EE5e+Kdxk
ZUJfYls8I5wI3Iw+jrvQZonM1tHcDyJYJuo8nlEPkzzzrTXyZ4SlmMgjeFWIGFWh
`protect END_PROTECTED
