`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HOIxoFy9PkuljTw+AGPyItc4GH+z5f453NsfxS9WMmGIWz2q8PM53PVm7IVkT38F
3LAFq2VxtSVgbUCeAschNxlR2vtWhCBi6P+KYbLaq5lkvXnCtUbmH4+F7Ekn1FkH
PL0Szk0LRxIGPlsQVgg1w5mS/Q/nPSG2CPxtruDAIPdJtKHwXUK9Reqqphdt3pGR
RwuisDjIbmltCYtu2x7VnLBEzxknznv3mHoKm/UvWDYLMra4Nauon2BAjr7eNNzs
9waMsO9DXbIXb381+W+VQBQFE/syoaWEA4Lg8xQUJGyWjDA+DEG07+qJO0P5Ay5H
p6R5rXLEoOOOItw5AdX9GmRZY9L3ReV80BPy5+AKfwSw3vYjSwtM/B7vhSfgt0jx
/k/ZKga6Y85eNCD6HPBbLiCXwVgFwnoTBZUz64twMS/WyDRMqepAUoHojVcKMEJu
sGvZAN6JtDCqi42E1unMZPGzx6uyez4c55nnImT3t4JxEWpzl0WAFPjDbmfKyBK3
VAlKq09y7M2WgMjayaO6qEHtTuPEB+2r4q6NIAgWlfzoe93MgIMzW9ThObQx+PFm
QBLxR15WLcsEdQnM6inZ1ObrmNfsaC0vYkkrqb2afO+9YwzrVI/3yOy+wDxcg2sC
pH5IJ9gnLka6U3TldQ0CSrjQTquoFYLVJ9SVVHlpTqVd4nsWMrTfGz+hiO2DX5Ch
QRz4CgAWO0YofXtd5wSVLfI3655F+jn5HnFYpAcxXa/rUPMo+z5kMzGHNDWEXUKS
u4iUwlBMLt4dQqnIXXg9NKrXAr5nA+cRcfyecGGtR3L5ZiS/4MF/TjiAzAqTXGfv
2JOd/nJt7WzYOMS0VDP8AfYDnE3olgRlAmzqxDqkjxEfbPd2c+qa7KsE95TS80k6
kfnoL/ZB+kUuE69nArbn3oGmheHlf/seKwGnvNK9DzphqshrggU6c8YcTAITQmJy
7/71sz0bI6qWD2AUz068qqFDDlXD6ADo7ATVWj790FvWJ0y7yiXzJXHDCImsr5C0
c6JvIhxTbZ/3P8RzIqHwS2wXQLvVVKjsinVdAWnMnB2Iq2YPdaW5+sk1Xrx4I7Wc
lLD29LZJPOfQqrE83G2Hgp3/TOni+Ac7e5CIpHwfUYaH3wsU8cbhlB4tl+DRLo8g
KkWA1SfHeer5iRQSg2DNjO8G7uYiwX/zEQZFrOe3RYiemZ80e1F1vzvInBgwKfPK
DxP/Vq0INEDYnSbAz4eDay+IuQp2HmJRUymWbd9XEjgmuoFEw/Mopel9uJuvPSsN
bzIplHWpm/vp68uKz8s9ggbwFZNH7iP4mHp9imEDrkcUMToL2OBXm2U2OyZcMQc1
tFaZWx2xI+SanOOJ2yZ5+5T0SdIR2hOaC0fXwGPfZbmsg4Nw/RvET5whLb9Pek7L
eN3vsb2aYvIGkW7ZNXu1C2nmZqKFU4RMj1MdEjBOAPQSX3xIt9gTIpN7LVKOefOa
`protect END_PROTECTED
