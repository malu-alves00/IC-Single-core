`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ApEOa2wLuUg8HN+7dTMvwn5rARUDkl/Q/P69Pyf9n9D/Hbbao5HGEVLskUjPQCWM
2uujxS95Hg8YY2bqqqWyIyiapPVJE9rf1KCnh0cF35NDqiXHze0w2OETCEvS968l
Nz1sfb32jSVMhuwHrNxDVAs7fEW6nT1OyOFgPNC0Wwzqq9nNsbH6em34LGjcJaQA
3Pjpl2az1ulTwlSHk/vBr8itA8XhNOQBHIn4lwZwj4mFxSrM7ciry0VvMlCPpuL7
VShEsLgbgoWVJGHej7+DI16wGyUhA8HFuk0Ulhh0ZUBtUYnTjerYfweRNAd2nrzr
jCtI5OuWq+jokmFQZTWdgWbnFlqz2f/ivZe3BEDaiXkyHXQR6yoZhcrz0MK34vpP
r6h8wnZG3/sREgd28eVIAfedb6rqVLV1s4ac05eI7bTtptTTUa5Ic4Xl4mnsFzzp
2AeC7LMqn3CfjmKzlPyzzvwfpJMV/9l73PUvR5rGlD/0eyER73uZKib17uZe7twH
V7RnmpWudLjN1JZ9DItoHOLYdZjAjiC7levklnVK66zdoJenyPTQbFyfZVgfSErl
ckJaTY4UVK9cR5H5koZ5h01x3FMtnLcWpeKla8mFNj9qJxANEWAgFioqu0o/b6e/
S/BrH2r3q9XEdauCxRuOukfNypuaw8WXN9yLqyexIzkobvgKU5AR2y183jciWBnt
bUxa6LjnnUR/hB/cuAyTK5dXADidcMKk+EDIK8R8l6+aazy/RrmZ1Hw6Ni0th820
HsslaUcIRnrE1qJNevUUeUphWAcHZBgwv0FOY64v0wu8xHBT/Mo1LEnUj7beWMEq
W1bjECXo/7e+HoqfXOP+GEOtAMJ3Ehdh5Fj4ylyL+Ln4Jtc6gkPoqFYBU4W3r9o7
qxP8jSWfh3kkH4CCscfmFsbQ9jnqa1D0Zb/KOyAVQJu+vzoM4EEvUcIdNjhM7Z9/
I6vONiBePowZl9w+L0V9QoH6xujp3yGIw5CJdzZEfC47ylgUDi6eFt4FAlvsxp30
/IMKEea3kejbuAiMcb2vdZarIFaBj5QxKxedVb4BoBey8WZQce2o9ODorgJddb1i
Kurh97PB7kPuHjWsCg8EbFdSY5EC//zZ81jYf5FIngwNs6d6L02xPkdaxKoxYATn
J6Mmuc+mObbPrIfKGV2tk7u4iWKjek2Te2Tc4kCYDINoYWFaG3ciH5UK862MSgsH
RH5iYzRBhv/bEmeDTEuebCUhQNwX3VxGhFOGLFNqq+t2jY62UJ4nlqP/zlBLjeQd
uU6hahtNoOGI9ytki5mY2g6ttOS/2jjTDyhgt4FbvUfWvuijxarNUpWCYrRvKA2O
U2K1rsH0AVMtCn5UVgl58W64arVuzY1rbn2aQgR8gVZ/Qb9w0Io2Jl47dh5zCHhl
ORhaMK4Wo0KO1E76yKXJipXVJ5irRJ/TXGhDCcXTnVwQ796VPZRvDWPCtKKXHHZS
02ONjLUNFkCdO56j1DO9suNeNQz/LO1OuUPgzuqUdauN2MQgmCpWJqSZpBGS6Mjj
EfIkPfgpvv8gidb3aNbg1ii33D4+81Qt7einbi21YpWEChRYSt1NbYnMo3fxN9Ok
7mSJ2BFSyuXoS/O/Ap8NGfSqwcMtUYA1Bi+XYPo5pxghS8abIOx/63DcLgmwk2s+
X/sJX4EHSTuuRL0f7KTZgK7CWkHE1mcu+JgGrxVpo+yESgq/PGzj9ZPXCV89qZpK
2+8ZvHwJcOxA5Po1hUuUUVe1KAajbFK3mkeB+XrA7ofq0iecld2rtFH1fQmFgv7m
lIRdf7J9voXZbdf1AdQ/roQc5J/6jcSo5Xnjx2CFdtAlIqQeVnB1yJ8sTJc9NlWe
egof+GKzaCzmL8mjmsedEyUnuWkbzNOnpGBuvVCtigb9wD3wJxjDNSIj5E3+rz8O
150clDKOcK92pRPwNczdCqcOaHbVmAVaok38urYGa0L/Lu8kmQnyRI+H6K/h6Dg9
/TxBH826C51t0hq+MNSyQw9xLQ1TUpSv6XNwS1JVBRDnf2BG3sKJY7tD66J2rDo/
vojtPuHRAwuIwRjZi3ljZb/dF+oqqtv83EwilqVuiEVhmOctZSwYbCSI8rWR1JzI
G+rBqylmIsET25vXJbq/2aT9/ZjzSmStdnJr3NFx4HvytL5NSx/TCgFIfIEMUkS5
4pxGJvH4vzbeC9UZfOihUOTgR6Vew47Pi0/crczjdRnq4ZQjKAf1hSrsFd+h1Eu3
z1S5K1N4oEeHPkji7o6iDgFJweQw3ditxIGQIWuSJ+XPYqcY/ed4m0hLjK7pNzUU
mdO2G/6AwEUGxH3wni1VK8G3un9nKc4mcKikQ01J/lwBi9xMC6FR4Y4k1pnkqddh
Na3J9D7VV4hiAaLvddB6Y0jEfOvGr6iICTYn2+BlDFvt9jtldwv0RAYzFXkgpxWQ
sv+lC3sY7q3MA5wRGPgcWJfr2SJszSkI9lqMATLwwxXNhdIb/+gsnMCzr1fU45NS
ljD3ISLSU/GHllW2xJd1TYdV2S9m4oXT5hyqiksgKTek77p10eZ4quSSXuUgoMHv
E2acvcMkIEtIOwfudWnwehEwitexSVnO+x6fWXzc8zzka0ABjLNLzQyBu3clRSFw
1Q/VbjPVjtDutSW5VErSPaMdOlUxraa0mCCvPOamR9El7LUpBpx5UVi1vkn5s89+
w77JmS/UFE+riDLAaAbjq1SWljVV9X2Et3pMpPzLETH5OOmRjgnBHdiLVXr2mQ9u
sM7BV983tJZM3HPXNRNZNIiOaIoAZcWFmnBKU0NhgdSxxo68Y0PCkyij/3dLMMMy
/OXcXS3MvGZmwc9oIVhZPUk8fMnks3FnQCPXW40KPqJX0VLEdJNg/RtVdJB2v1wm
dffHmUnMTHbC0KBtw51gzx3y+GGe/K3C2vt+7+yxBMNVeD63ld7/kYW7kMYNuhN8
atRZ/mRJI1ApLUAIUWcGhbYZbVCJMhJOiW1pGHlw1NmXVAYzpk7IgksRpawJKjFq
OtZHzqfIAlCLvkpjR55kSIrinaBYwS6lAU1KSKKXTpDanP7jLjMw6xuYcTtAfPjE
w58I1V9R+2usF4IFHnE6OiRJkLDKoyjB9ZzOt7wXcaWLxKWmD2SE6M0FoLqtqQQJ
bmlrAHFZM4PS3kCiO4+IpzqtdiaQ2fx6H8d9hLXG4E205GnScVlnqVo1L4PxJCMi
KRUDU0zNSujSImyw6Zg86zBNh4w4l7EvgybxWeRg6zseDvBoueBVcJowISthCYLA
8PD40cNbebIlmxIMXssH1YtdqqmtPNLhKGZAZ2ZDw02suyGqNknO9dZ+/ANaTIsn
toJYLTol/dJ9ZMCPEmA87v3PjzVNE8IE+qPN33ANMUlsiDqTcyrcQcqx6SZf0+Gc
24/I58I8zwZNLYUiWZToaXsxo3IO6oek2Ez0l8rWbrT/c6KaJtG+JCzjJO43VNpG
2s3KDFvQDbmCNV8siRcHZa1BpOVikb5lUFb43oa0DjL+toYN/7HbPzWSScjrcsez
NhWmy1PeBnWr2mWhUJbVz56TvQSu0tGtETZPdHlxjsvpisfue+1tTAH2lb+Oitgk
gTgYnFR5KAFdfR7fV7Z4fQPIDqFO8UDblERVzqgZTKa/njIxIh+b3ykgnzrPOsi1
gklsUuc1UwSYUQXT+AxtAdiruSXvH41sms8U2nAFyUSzEkXHyZObMjBd0cSPPfQT
bUszN/5fEXKDXCstZiPCEYUb04QaTMGEm78tio+amKGLhtbrM255TqaANgcQt7G8
ZP/gal5pACJH7+WCuykSlDYnTK4maJizO1YwSXJcSNyteykaRRrzbvk7Qcj+uBxW
zg4Ut7O+Z7nbAM+otGGITuMd4EcVKRAg50i9cVx/uUbJqWaIbg31lO6IitwXbQ1P
Lo4d6FGm4Jha1CUNwB3HJX/sw7yArpnPEobmIlF/NxgKEizbGW4l+HZ5IZdJlhZ4
dh5eRJ8y9qt83HyghBDFuB71F7Z1gHSFrH/CCfkAzlrlYCq8pPseqtjjQxGpF9p8
WM0uq9UoKH39fn0ajzIlbF0NNSBuwTRh9vuFdjQVb6oquYjMYvK/3sCTb6GNWL4i
rOgHVQ03KpBfKVxLnjecrZNk+1T/JEb86y59Q2d3gnK8wANApI174llv8AxqUd2T
4BYwn0mZ8SqRa78C1Q2DsT932FHbrnR1haCnPb1CGcXK/zHMoPXFkRPhVIypqDAh
eg+0OiCGBHStZlOMRFKplTK4ORBUZA0I+ntJXtANh7iQcZEBl9JioijeZfMCHNz5
ZDmm43Oe0LOdV2QPnoza7wxeOn8Wc/9xYl1LEyCFe+Ur8RmvHoR4nCzCrwfJf/Hn
iR+ESIBQVhI4EoPNSe5hOImBEobtTAIeRyBntlD2bLodwyGUzfo8rTWGAsSyAXkb
c65qazOlznBuXaTWpDS55Kv0saux95q61xheOJOrA8Dn2gwkFVWiVYXUap5wQrP2
OpbNFISFDzRFk1cRlQ7mx64cwEdXd26O0V14pdzznfmd0IDHZRDZYbkYXq8BtQqX
fi0ijaW4V1h3Fcy+6z95J1MKFAsOieibemRM1PiDJq6Ad569aWtqdjbKSThJUB8p
gj0f/xZaYOA6HEoF0003tAdP/aN2ezFs5TPzr0sCxIBUSKKBABKWJnT5tLFF1MRU
QtHpeJJo/LLXVoU7FHKOdfCh8/Ho/v9GAiwOyFV6XYQXUezlacustp0xv8A2dm/U
K28mgxjfZKy68C42tBV3ZTc8ESOSd9EasLKpaq/Qmp3SFGEVySxCmTTaP7plHMfT
Jr1/X0b5Kt0K+X9eRyQeXnVJlf/wQSQkQfYKKSUsW+4/x8Z/UEg+W+mvbDdRoLNr
USI67vb39ZLQRdFQj/Q2RJ3eVNhAeqi2VM8KSSP4jx0JLwjaYEEGaJ1GXCo0yhjY
SDbPSmqYhRtKc8p6j0NkL/p2jehHOudyXbkngTDRrmKnN2PnMkuIFlj1X4eWeohu
bLf/LKVNygkF2BUX0+YNL0bTk27yPYEAkQFIH1aAaxePJN2IExn69s4PDuvQMbhK
kai9T48+6Qt0kBA/8BgfIBJggYdvmR4XrXaF6cSw7lrlVxZTZxLPVneNkSvMIQJZ
nian61P22u5IhauN++N7bWfSvT3E9i9g/rdeR/gp6UZLy1v4EYT1iu/y5UxcwKRI
jyYjh2BSOueV7SHL9sTCaBvcLM14gV4dtwXOVI9vYhya1RK70fKAtnjswtC9zGLH
RuDN0MnlvvWvPwz8aVg6dCCKKgIpNCmmcweoV5K6AUErdqJG/3mqMopR0ocCEH6Q
r/pclUov6xaa+aUsJVWyVN4NwLluYRmVIJoBAaCuq/VvaoI1vqeYeaQWULdKthKI
FMybRvo7klSBoZyX0SBla3SDH2c+FT06pjRb9eRbGmdYXjhNJjtSxPpkZwlauGTx
vVjp4jgt13m4z2gwxtjLksmodFTs0ckiUEgG1Jogo9E77Q32bNlzgzfdY8b6gD4g
FgaJp5zEtPj5Agcl7eDPLvPrBYrMfWjQ8RG2lbRkiq4FMxznc0tfDBaaZxkdh8hL
55FQX0Mvlx7iIugQvzq0PqqO32yKoUUtiU3/v0wYvV895P4hrjTneW2N9uubnbkh
SaPMOcqjbiFJHYhyd6CkZdoVzDPpn1YqInUOrFmajEJqM3+lZjBMoPn29gEClsVM
0h6ZZphD0wITLtyuIa86NrBjI/LJY1NkZcQqHy5udlYyh7L4UYUVO55EUaIqjWe9
nT73ZYaI4nvNyFD0o4jtf4qS/TCzdV2ImsZRU1CSxuiHCWIMh6HTF6bUUEHMef6O
urqGGX9dkwlEG8tc5H6adVw/aAtqtsjwFX7JI+zt/ewoyqHrEag4+dOTBmqVaIO3
aOJzgvdy4VvIJPdQJNorDdFr/+fYdMfmLBycolUb8RGdFs0Y2h9ve4uthLMd2NHU
HgFAAiq0FmzbI5alQ9KdRsegNe2vtdzS3u8LaaGVk/htxjs/JlYpTUj5l3aYX3S1
pkslT9HPPQfRKcUOJLgBIZ+bO4QP//eSsUEmRqDNiO9gdibIct6XRKBjOLJNh09M
C/YtgFr0H6CdmFs3ZYYSllKCD3ksq0JiunisGIqp809SqbT1asNGvUEF5W0dK7nd
IUAvYzJXlvsuttkq2/VOEchi93AgXDl9+gD6NqUvBQMZom7q8W/CTtpHkvNmqmpV
o7ua5ms19tTC+LjAW6irSl1+jXWQ6E1jq4RLad53zuzEn4LeDzE+u8qlVNV8aIl0
gJozXlhYvZFCVfZSZPNEk9lehxdg4WqP0gCvw2KLkYhot7HWgglpCFPO37AES+Up
cEuBEkmfVINcyPC9bChvSHmCtmv9jSEYvz7RdcwXaNqZSAKxfaHppcovEbB7NT9A
RxLnXzHYiUdR7dJ0C3qDy0m51FIZVNfNN58eOq3rQBMzRU3ubZ8onYDtE5Mx8tTm
vn7Jt69Ubv/Qi56KsWGonK+OprmVoe9sS9h2Emz/zSas4ixiXddkmM6GOK5yRlgC
9D4+tIsIKXBvpppBwCfIVOurrTXAwR9QayZU88VOMpQgcJdzlpZ08POdWFpv1SZa
xRpCuNqdRfe8dSYfpzR4wMbkAUpXxf4HYQqUedDnC4ZRu+3qhTkeyaXRqZl50JYL
FvGhBiz5wB8mt8tl2Mih96fI8dXwjfEcvwwm/wT7k2g5zvjMS0WxfqIvN9DTQAZs
Gq3ln8g16CJDjApzPu5HLyE74enbnz/McnSZ3JDMFdIcErPxamLs4D0fjy9mUpwY
srg5Oo3TxCGU52KlEmACnm18YtOQLnUntd2ZfQHD5K3IBnh0/XKZc23E+Ravghjy
dSUjtMLVc6+t3q08NtWjuBAVgevk9MNl97doA8AEDwzwBrVo/VGQtu3dOtmdk/1O
L6StkeDPQkE79sgdpBwc052Bgoak3NQpcyICGLdLUdDTDCSsDGRvnkthyEuJ41wr
+FgD4OCFvdS26H9r4Lqsf98ktt5uGiea6NeCBqGFMyKhskG4SnbVoSSGcEhANRVp
yBI4YmRkL2sG7K2mKLl0hUHf495nYRV/NMRCkuem/tqnQz79gJFM7oHaB8A3tVif
VOOHLlNgY2/I8CDj3kfAWsESNcecY0V7T7MLazDMixs8VEmPD57TrR6gzSlu9qq8
olWr09wGh+058fCUGyw/3UyVRpnQFPO5/QNqxI6Q9GWXGkTdy/3tewYgiyQ9H2AJ
Stb3stFjGDuZhSDj2yB4bIPbH8SHKqAYDYj6tWAR2MagBnh6Az/xk8ESSSH8OlgX
V7oGhDP9U+PTL5FlnIEOlPN8/oUMp/Q982LJL3Wd+vLbrBwsPxUWpqWFlrRFZE9Z
T2fTOYv+DCcQf4Vd0W85Ne5Le5MVAVZPWFjNpt+niOzZpupMNrctSCxK8Qf+2kzo
83clPXgZ+wdyN+/sKH2bA3LpiGd9y84dhY2dS9Q+DJioPCO/CLY4w3q01tqYAa1h
5H2ROaR/XvmADgAiZr/aRAurLh9GCYrsgZakz4+nfrRBO1QEPKsa1jrhAgq/OWBy
HwQk+dOVR7S+HVfA5ogKR4d8hwK1qBuUxKCIDIp9lNb86iALFhTRKoK3ZAxuT0lq
Ybz1sjnOw34yx15BrvPIwIll9DOoF8G8a81bOvifoP0EApI+Qlc92a+MbK05WduN
uBGcab0LAf5jPFmaj8K6MmJc4gEZhoHjKtTjljWJdcHzZuhKISjMbUBhJJMlU4bP
noB+NlpX5ByOOosk9fg0gif9IxZQKB7bSiSx0iyhY4uWZbYm1VY4vkNSN3drkasm
Hb0wwJDXYsnACxMOkjZTo0jWnZoeSVVhtAr8DpstMdFkHHZ2TiGYoKW7Lml8cLuL
1ZBDQunTmEyeew2CFgiwoNv8GLz+ZaqrlX9roZ7pfUWv0ZiNJVTTPV9oOBkFUvo8
A8k7FPeq0+R+DaXRm91GEZZc7MNn6YCg4pc3qqGHnyjXBdb7zhWBQdw6KTksn8pj
zc8hoLEFDGBMiOm/keObdtErH/dOqNqzRmOhx+ssgd6B5xhyOklVCjJKdqThrYy3
UGmIanoLfQMeh9hDGS9xxBpDc3PuADpY4AWyGDII5XvJMSonA7rxzgcBybTUY8YY
hnxg7ONtzIHc6vB/9swSYtMxGZgEQzwoWW9K/gHPjf0th09qWZBgmPYTyuWqmoGF
GtjMYKFdgH9fCCCbrsOfAd0m5nTe2yFFEWn9F/Smx+VgGkvkvUiq5YOsv6G6AUUI
P8s9KhpG3z43uOscx9P1+85yni5ClMW/gjudcvXXbKUt1/n/ormbysjFD7xpxczq
D2ZpCCFA2KdjD8jQv9VPevGqENr/5NciF+M3MX/1Zi0sL+SDpxryqwWY+1PGW88g
eMkXuTgCpqpGc0waw+j7fNFp/vIFK06BbB7nUSPYASyuNeo1wwAWF5IRXmURvyB5
SzWaEhxtUFwkRGOXmbrWDo3/BCMM9TZWPHGGDfTzVZeWhAhya5DTY9RDl1Q9y/AH
EQY7a+nTrXKWeqVzOOK3mJ9HA35ufgaXv3GhLkDyRW+NUR1gisfplCkt7KVev2WD
c/LKisldkNNvJQMmORmtls+emdGpq9bUrBTuh+ztxVf700Yc0nd+xPVsDFTGD3jT
qFkSe8iXiFQU1QQ2EiwfCndo5eO+8iv9gMRIVSdpQwMtLxRpELYkkiu3Ordyp1lR
bMOjJLYeF4iJRneP5TqN4JgWJios38q0dH4qLrYWLs4f75DE3CT+WvyWCA+7IhJd
8uB7f7l3qDfgc2XFWtK6ooPxcsAQZHaLf2CR6c4PO2km3SVulOGK8cz9vdoPLIvZ
rqnNpKz5XH2gytSyfN9Jha5+pIna7eval9EPdiqK3Hkm4Ifp+5b53PHhA0HjXB2p
SqtPVDNBOfis86n3mq5Dhsf1tCsLsEX1i989MgHQPg5KIXASdr/SO5qhrndn5hF+
Lmukw+exinOq1/GV3YvL8Wc8BBXYDYqq6CcnREEisAFMFFW06Kf6kaWa471BB9lz
bHRFp2SLApJYSIERy7BXnQ==
`protect END_PROTECTED
