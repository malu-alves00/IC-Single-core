`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
S815XGZttsjPHwJEexaOchEhA4KVq78yzsi8UT1Lrqw0A+mPDh/qN5tOe8UprcDB
kcECIGxgo0cTAdOJsWnxC+EXpAMRItwLjJJTEXcd8Lj3oGmm8+4X2hoi34PatUGP
6nfIlnSQxQMxC2vsgaDMsZ3I9EKK4gqRUHkYbY5Yoz9DHmaVYD1F94q8w2I2MlJV
ZT2S5RxsU2vDJAA8TojjXlGY57mu/hrGNyNZD1hf52X7rNgQ+sCA2lyOOIJx7Mfl
1WYkf07E5lDA6QSpbtCNTVYher1QKmhnlR/pHUTdVZhnrU7MExIknbog1uM9OJ4T
r38MhhdOEv0WDfQ24Dgg7wsBylOEhzhC0hTUnr8VsoQ92/5m+o0xgKm7zDraEUy1
Fq74NRTr1FfcspoWK1oCZLTjejLsG4jgIgxZIi36wxJ5X3xP5SJzVhubPjfh3k4b
PfY4M/q4trhwu+8/rquMLM3JCwvPA014H5loe52jvE0OQDLSriPmxkQYwdlibVmy
hVmWfS/IWkN9ptK2Uz0ygePoxl9rF1EgT8iCvGJ3hEUM5RMHzbKnIfWZ69jrdbiB
rx35Hvn7nK69PNog0JqSVhurRzL5Qt7RMwssL795scbjCq90Ic3PkCAwCJw3CsIA
vukYoA8acIK50yjl1YGIoA==
`protect END_PROTECTED
