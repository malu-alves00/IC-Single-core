`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KPhb+tRvHiyXsDj74VC2+rUeSjqbxyUUqTTLkTQ9S21pe+ByV9br0YqHImYe8wUE
qDIg5KIQAniMBVmUrZ0kYw0WK1+fGiccUTPNttQZWq0VUIuvTJIIwfP9O5LE0gIG
7tCdr6XqhUFDnLzaJz4eb8TgvK7Djdd6qmlxKmrB5ROhBBKL0tfyq3bgJhSbBkaf
m7oFSkkHN2TMKajZ6RI3PyGJMaVt9re3ZOYbW7IfLLrDwGqDGKW7r7wONiAvXQ9F
9xZehiMUB20lG3gmAQvbgwNujX91jjVrfGvnRQ7CX2GNt2mo0YLUVp5OMr+tFkdu
p1EnG1tDMjUkk1SKbBdeaaDioPbKwO9fTkhoOL5S6P3pXTI3T0qyOIr/dphl02qw
MPZ5z7fA+O5eEpS/Wyr/ZyXo8VUprJlIMWrBboooajF0uV0vvQG08grqr3cv2Fp8
cv2nB/dkPHagkwpTVJcM4tidkuNbFzUMn7c427vslRlabeJs5MPj+CxVBQX13ZBc
gOD7wK7kWudMZGbP1rCMzNGIrZpWtbI9jOVe7PGJ0nEfhowdH2nmJZPSloo9KYbT
d+lR34b0MYd+XTddJ+Z2lpuiVopZA8pHVAuAkXfTYcy/sSqp3i4YIsZl4QnGUpFJ
fEd+4tCZVraI7YmrmR2h5uZlmtwoCyST+xKuoLTRMQsi+wQ5pISvIfLlQC0+StIH
jqL7piPOegkGAWxuBmaXPmnaEKsEefGcHiIbzmRlNnlASCXLN5kOBNeQOhCGHaMv
GdqcsLZ5QOUXodg/IB9Bc6p2jU8+RjHZCTmocJIqyyewZcjtXbNOpPqAMZmghwIl
skPfoeg4m4TJjx2k75P4oedihDBNxxoMSrM7qw8KVMB/Rj5+TbvUhdAiER8FuLW6
WRHdqRqfnMFb6ZJP3mUiXBtbo166DqI9GHgecdJxeeQul6pr7VMqy3NginKEqqk5
q0PSDYpS1+suSuyf001TF97K2uIT0pU/UtRx1DFZgFbn4tLMWxltOQb5Br5lJfae
V3v9vzU53aFPy2z4m7qhfL/qpT4t/wO6StaRE2mjN1HyKG9anCQTrmonCreZvLFY
9V18r3KzU3ubwWrtwgY/+WBk+SQBRCXi9J2wPIpt07M4RJhjdNEmcbU7n1r5aDOc
vAz+2JutdzaCg3QxdzWFlQ==
`protect END_PROTECTED
