`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EHvEOsAO51auDLZBin2bb1JNwzyK85U7zM1YqBuxcrZiROuv1sZN8qwt85Rbk31O
e5bsQtlgE07q7tBNJpubmMczCT4MONu6LHd7qauvWTw0KTZFeD14DUQmLYA/ZcXa
QiZ3v1svR95FDS78lqMuyOCF1Ir4rDuriogo84RrTD0qSO9HuBAur1Jg2sCTjPZM
bMdeLMDGaxTS5v+rL8mhT5OGifLep2dwFdLh3f+qyG3AqKGDTPrEx6mbWDQu+VMP
RX2KXzrbK/+fPIsI7u/7+ik1IEEvp23r8ktQDK7MBpyUxdzv40h+Vpz+Abt4FlG4
98CQRCDuQHz4Gjy0hmwiDGObKDPqRguSe2vhVHCrRihhqGqVnRGpV4cYKPw+naQY
H0G8q6cPrTuG4uSMdHMmlcUPHf+fs6Jy9BT9a0xPyp3jwxBysw8EJGMpDKhRYMJT
68SEFXPF+0UQISmc2LLracZeMGr/i6GIuvCX0ShJTaVO3oCO6ZT9XOoOH5lgVVue
xwwnWQ1qcGigt2xMF3LdUVIHOX5nTfTYPxZf7B4qaJOkd6VbWvOJ6GlhkeYNKXQ/
t0R1lqA7+qQNoWIAYgx0V4puwixa1qBDTOStT+e1fVjWA4Sjv91fxU+tOP/s7Do6
Vp7+0qLGqkkn4FG0pGOjHXqLfKHg/RMOx9YluW7aQzPe4X8ExAhlDSCrRUebsSa+
gNYM5GPgUP9sTgnEhn3QFG8fqBFTCClbaUsSstFnwd2goF0Lc9D1cojnqwsLVpKY
qzOCKNPP0cDxu6yrFDYrMUFIVzctjxU3S2JXPwON8hq/bh8BmWcINY+qa+2n4GN9
Tm7P5Y1zd3yTk+5y389yJ+U2GoWISSS/LSWjiFjSYfrno5YyQJmJ3Dm03u6WkMEA
`protect END_PROTECTED
