`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PQzDGIetju1U8Gph1mL10BRBxha028rW3j+mKL+dHu4KQf5KN4EaAPbH7PlKPIEK
Pb08OC0BVonElmQik9ZTGw18Gk0LDk0nwgZV0OM1I8mUBFtnSu/zPz/Rg455iCLT
kxcACV3kQGG2IhTUgnlCNexugm8rh4l4FsOxhqoyPJySnfoHgGCEtYPGOw8ZMN3B
MCB6NLp5UylYq1hv/mePYBjUHtVr+SAuhBMPrk2Oyi3judQTt+QIde9RRYhKLQ2k
tBTvakE49hFmyw4RKgpXUMoie5PtLuCN+UGAoFh/9ZC7mBVwwn+U7WlRRVwFNfsI
GUgc/6ITzAJULKQioN1pFlzcQ1VEAYdg9vWI8bW7uxzwAWhSgi5sHcA2DhfIbgAH
HwuoBM2KZVo7wsaYR2IxzZqz0PNnC9+weezZlwmXDh8eKmXabZ5AXmL/aj3W/l1S
cyygHBptKRRS4C1eWTkViEt4XpamSud81cDyXk/Rh10YOvcYCVPXoRTjMfC1kUfk
0wrhR5gwxPFKf1MErYNEqQquqGaGezc3GEN+O844k4z9UqKfVyJhUehm8PWZutRS
`protect END_PROTECTED
