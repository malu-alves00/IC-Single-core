`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4w5U8hqfco24rFSGXlD+XiamJh+EzcRB2yxojjdFWUhZwZaO/h+WAvb2LtrWq7ok
L+oIMC/KUN6b2aoD2srjxP7lZ79YI9LlM++25EvhtZoyU7fFeuoICeOObsbEDlja
4djjxRwOLce7vnVmp77gjdd+ZkekUfOxPM/Ztp6isbTvFYvdItnP4XDlDuLV9nkf
fc911nW2of+u3nhUm9S3VeeOmvC1rN7HdjVQlzWUjmSCTCkR3JRaBjtr/VoNMDK7
RdDhim7tyP2J+snocXgch1kEJgOYJev/yinSajoc5VnGMXdVKfao8zTqBe5erxXw
SyPE7PfM9AuTaHiFOZJTqfYZqSHgiUzS5Xj4DX2hvGVN6kjP52Ni2ZvrvxFTFAZS
D6PpbCf78pcHeqmUrdBd7tN9ax3h7tyokd5cQvAWPU8tltc9apx1AXX5yCd6NStg
ij2qbl4DhLHo+dN8OXqquBp/hgK1nN4RzMBsTsOdpbcnFRpN8YsJ3yCvOtPKRx64
/pA/PiFK5djGhkZ0Q90Dpyav7Nd3y+98bvu7XJgbYozFWJKJK/L+qdZF85jS73tE
o7CnXuPaQ2940CHMQN1RpKsU2M1k5P0pNCvEpWHz2NxCDDqc3vheNHsnUqVuMaB7
tJGDNbU3iGW9WMQL/pNIPwYFa8o7qqVZQDAVkR2pMhkmtvN5evhWY2aDYHQ8Pocj
OCxttyWDiUho1/x9HRURf5XV2ZcEQObSFhDkIx5a+ndVcOHAWuq030duIUSw7/NA
5Y7QKp7/VJUwlyH2VrXRuNscANAnVqfyQkzQj8BKwXNaKv90/O8COYQXt4mwBmiv
VwYnypAGmM2g5jm5SPgd6KkQmbcOg+MOYeX8Keniyfd8BsUlLPUwfzalFBE0vn8w
6Ze2WnX9/HA1eWNPFpDGb6ZV0/+L6PyJGucFzzVEcsHEyPVnFJnk5ozxOX2kLdZN
oWhIf9FBsibaXDS8QvG74KZ8WqHXjpUhQhBr9I9Vkoc+14zuWalDufYEdQQ/VC76
T+AVJdlzrKqp5bLXLsqQ0iwgJSlFpb0oYadCTV60w5x493DQqG2pZ/z3MajFNOpU
`protect END_PROTECTED
