`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zyA++UZpswCSfRGk+8p/uc8qbt+W2qY15pgo02nvMcLoOU31BWY+2Gpzx4CPih8X
dxekh4fOBe7bIAYNhzjjGdqMo65BDZ11BFF0EkSRbc8S1mETMaZEF3obAk8tTTRL
dxhUeD+kctH1KcPaeFPymSZATOE10dXURTXsSZRPEFsmKFX34WOyb/WNsGnb1yTx
8TQVAgFWAC8bXlON138qnjfc2oBPHlOv/+IdSBPaxErEe5aAMxPlDabLRNH7ZN33
0itEoUv0M+t4jOzLrl7xWpo1clv6fEBuDb7wW3jH4dnWuAKNORwICO0QDWAd+ihK
dJYY3AxCHncj1iZ/HW+VBcK235zI02xOD+71h1+cP28QC29G+lYEmekLb9mPAgrF
t4SdWVNGoD3xBOcOv1MaZNursqWQHfwRkDekoahaL3Robz4bVOlFKekW+cAVwcb+
icyN1UL+ciCJDdlQ36hlK9kb3dmSFHdnFNJDAZ3IAMq6ge3jsnNPyeBw+9qvkFnp
ztc/TROCvPw3ZdDSRInHsD4sWAI2Dew5oaBolv9CF75b3EUylelAjZa26s9F1v3d
uv3Oq1UQEsAIM38yJskfTlHMkb/bjiUyzz3uKfQqNmqr9vjme2tRvb+33S8siQUH
6jbobGxXXUpbbjFVfb48NuHuv0lJyja/J+ellzUu5CaQkP2ppTvoOC25olvzRuH/
5FLRMIYrcCQJinFH1uGKoBwE62mbhnKHAL339AiS5tlpMgQGJtHbIdzqF78jB46h
DVPpKvHcyTt6crWunBEWV5P9desXGrITRNMESwI4oIb3+OQ692joWfLr3XoGGpqu
b4h5J/vS3PGNVNyxGZbOP2faiCahJFGX9+TxK6gee9mSVQjg0fFguq9qTzRfZ3Sl
SLEzbIulxRIJML5ZjAsRnV8Q+qxApX3AOaHECdS74AQtqJNSZx8xHbTpR8z8Ai9Z
NI6y2F3WvQKMtkeBkN7As69kWLJ1Lv1NYLN5awlbBnO21uXCae5ebIreLXr7E+XJ
RdgydNx3iOwrLFN/2zGbEEa1ioqyH1ugNjGS+/PkTcyYlTQn+IkLZM8OnOuC3Krc
ULFdEXNHw1wAJnpy3oAR0Yk9Q8cKLa+3LwiAN16wrbmr5giPfD5q1U9vvt608Qrk
1Vm0p1f5kGO111ReVC9GRgcB0ZkPfdGmlnFG8Sdf9S1RGbkV58RUtr8A+ym8HoFf
ELvaj5iadFg7M+n+TLOUr2zk1B9xFRYOFKt/AYYApP8AxiM8gkMHhQevYJntvOxF
lGcf6wdOGl890OkL3PiGcuOw1DGtTl3j5U0kruq4jTOse8wKSvXWGxE8lb7z73uY
yeSPqr/RsUaYtvPijKvXv8KWUKZgW0c3wBeB+A2JzqmJ5UKltWBztN0W0BCB2hPT
sdaCpk5bBIWoBhqLFdMD6TjpNjVwjXX27sA5xs/GbLBJT6Mr2RhgP27SaV0tVps+
kzafiB+F8tNueolMPdUHNojEQmvuPGmcEiGWtcrH/ImStIaeHG5yEQ8ZLbCYr0F3
jUvhubHJty8juHVihQBesCul891TuKHX/l5AbCU3W5ydkDwOxV9OukI0S6W1mBVn
yBZU0r20Gd9RekvDkM3QIwx/O2kxHPsIIyLGv4qagbo=
`protect END_PROTECTED
