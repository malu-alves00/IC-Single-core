`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
69DuHxR6pnQ2utYg8zT6y7ZnCEgpkTewhHmwd50Cp1gRcbNvJjrcyZc62rvhQUzP
ixdyTh6T87jv8dIuRaguvWfiFWNmwd4+FKQdQwUNWvM+rE5X+tzpfKLoAdUuiNw8
K/z6KaaFgiv1QJuk5BwaUaLuGn8MH4vfNeDdOuYD5KiJrkOalCSSmpoZT+GXRkZZ
Cxre22+xq+6JmtKp/+JdyUU7foWjJjhFnfJoPNDonky9Tp6foXV8C/UEGVsLPh8p
ova5NUMppsTg41fOpcFu5cevXWrMoycoXASqPVYFK2S2feJ7Wf+bAO4IlhG21COr
l3re8xudCtxlfoDFN/ne1wOOBT8xklJAo14CBQs0u8eMYzOHKjDI4NS0JeUN/Yyc
4xsFulnDpnuawDJSh+mxICATKYLnYJvfhrOAJhc2PNIN2g0pTl6Ggrv22NJOnPWX
YiFrk62xpV+1IJ+e5ROSOA1KJuGI5qnGCU90ZIazlbFdbfbBPeMEohLeva8//a0P
EIs7HCb514OUEjjl2qsSPpXBDqu4F1Qn8z2jaKmUusrPLTpwVVHyF1uwJ6bq9lp0
gyRFFTiZ6WZdy/ViwFfGbhcfu4dsja8eFaRO+Xjd084pHJleE7lVoBSPaFEeRiUJ
BH/bo5BLdNMqUjtLfzhe00JEwpuaOYIrey6otrCLDXi+6YVxchwvUzJPuuyOUJeD
yU7J4t9LFxGSb/PkJ+p/J4e+CL0+hY3iOtWM+481ZPA29yQUcQUufyHD8ISw9nTc
O4kMfBr+aK6RptVBYZKQSX2JuZPv1ZGRuhzIpjNU/Vamqy7aX0vJpPXhBN1x+FVN
/t6P/Rrdo0zh1we80s9gTvfBjpoUmEypWnawA2go5jbaUq8Q61mbECtBi8H4PgC4
MY6scR+pMcY+A9YcOE/nJ7AwftLH9efgmNnUpNEkh4uUkF3BwtDna68Jsdkuoo/H
kv3QZITrg2whLuoT6G/t47GiIIm3vh3huVDi+rj/xX/0XBdjDmSnxB+hfHQdjjoe
UBALMpuqUWjtuWgv3/ZuVs/p6TmEfysSYG19I6FZSNT+CTn/oH0UEr6LzIGRZJzf
m5H3WsCFiwNU1QvYBeOljqNqwbIb/R7xENvBFiAw55ABccxqF43oj5WicFejrsCv
gFRkGJJDoC6/y4+4dDZn4E/9L3ONAZp2cnv+D4kAjkusgrvIfQp2HI3a354lF3Qv
n79qSVRsaN9MzSf+2rdZt9IaNv0c02QV7zvEK/sNEFmCOe3uARRO+4+ORG63axZZ
4m+pGLzhUDPFhJ5Tdn7FyM684o/g29pCY8zu7mkbrfTxWfunN7nHnZj41GgQCsmB
dd9T1PdsTgcHsArGszECId/HBcS4qTftdR0URV7yHzRDSmOaqdPoVoxzwsvX1zab
qeDIMJkyzB1IoNqkwdCSa8n3Z0R4vQjKfT5fYY09aJL+8OOlgtQVj2Vw85wiMj5u
OApE/usNyCM06bkVu0Zvhqh9a0JMcm9CKrF2O9EVSVCVWWIOCxub3bCVH5qpkKf7
wUe1xZxd2pQ6I1ob+B7V2gAXlZsrZUSK9t2HzGU6os5glix8Xb7iOdJh1Jjid0ql
R8TQUab8vKkQVC77pRBRu6VbXjTpQIqiw9hrnlpEA6bVpCnmbo6GJs3Wf9tX3No+
RipK3NvlSnMYAaSFrV5KQETq5kaREUMP2SwDzTD4ELQyXTMICDyrJmSpHT5psI6g
KC4W3OwJwIB9fd1Tqc1WPJR+ZqXm5y/KTSh2dkTcIF+iIMHl/AripIqv32hnFZgr
nsOOv77BxYB4SHcD2KiAwhXHTNKjCKMO9J/P1ZVCdDDR9LCXJQBORh3fCR49TsLp
5HKsEwAAKVFaQcj6bURzwF8H/ZsATpp8VTXJBA3xJE2c0P1Lzgi4Ze0j/VZEnj+Z
NiXZ7wU0e0B43lrK1wcpZNdoMur3n4BYmPW06eUHNCkkXAogJowyRBoxqL8KE3Fy
4asFnKJqnBH27kMejW+YxwygCsfw0/eb0JD5u9awUVwH/jR747DP6s4ZF18+nI2g
HmRiMpHNKp0ioSzh+qpFCq4BPtrrRhNS8pewWCpDANKdH7QuJ3hINN9F0/XrDr6W
8KGA6+ldAAlts/tFR1h/2ZgfBX/bmQ27LspPzRZmrR3lkXnHn02z9u2nX/fjINb3
JNLNoHH2UrWIfjou8NI4JmLQqTukYzxL3ntUqA0L7Gz5sXfc0zujoDZ0whdwHSiy
fOOb6oRB+GF+sHSnCAiQjsc1WbPCeBS1fdNDS8abV1kNz6QGdgNKVLcvC7tSFwsC
cggeIJG9US9yJE2a7CTI+mpcRhjFSgLWS8BY/ESyAjZWcQxTPfP5VFCMtOcj/iKk
J7A2B3R6gn3+YojZNZSLRLX9RP63u1oIyS85lZn4CC3Mbd7E5RpBbokXOBZLDVHi
QZ4VhbEA0MFmyKr8zZsIy1mHJFmEG4OVYidXNCvfDZUXJo0u5KxDVvZo+MkuoG6d
crUmHMDbh5Qt07ainEBnZVQKb2qDtlb8BhptDnH/33h7+fuRUQt6WA+T6/Qt1WNS
tgn7FJ6eO1MT+cQ1NRW2KBMMMSPcKuEe+oTRtAIcBmYZbZf8yswhrFlTCyhTfv/D
U0b6sNN2ESwUfBxLRfqiOWIVnONbqTIb/NN3YzhC5U/C39O08XibTRQXtqwhwsXm
CAEwxDXR4ouyBfPUmQMeuFm/D0EqEl7w2cLMJci8yXzluRzPpSZQ5H27XS8uVgj3
7m5Cqb9WYcj/TyIkNQTDTj6EsUiqH9Xtrda+/8+atc1z4A+uo+Z/LLhPgGVzAR4I
gDqRVLGE+StPRjzaFvmg0vc2cffs4ajrOvDpyEJT9imn7jixQ0iMh4ULy+fXAefZ
j8ZiQeU5eYnQ3sxPRVg2TSKFyGCvfI8fTUp0GmUobAUJhV97hCLCRrBaMDG2Nzm4
OrMV4+6Hfm6DuDl9X9H/8+344uEJs+3W5YPTJbs9C+442kozykTycoDF66PMzvxA
W5+NuQIgoOzg0RKm1xqEYdiapwfKDmFSy98t3cqSN1AOj8mrAU6cHor77hNdeiQY
cLHxvZr63edUky2ImXRj8w==
`protect END_PROTECTED
