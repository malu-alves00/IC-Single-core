`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
l/um1lHDPf9W8xkEb9S5PkVk6sBMHdMSrU5aEJfvLFHFqhFMZ4iNOOa2OPoaYalj
uXpaPslqEtW8TawzmQw/3TSE1afdy+L+cIX9PVIrrbGws/W7hWSuTnQ5hO5m6PaI
CCwj9WmEokgBPrk1eZdfvFGSRsHowF8KsUxgkogY8+keAkAUKcR5y07jMmsSmm6f
64yC8mrLtU9G0eUFujfrDbF9sCD8SmEaob33YlaFznbdyhxisIrugiCLXS+cLWrz
UbEr4Pw0Q0DTIJICjpVp4v8w1DXiSDFpvLq2Iiymq89iVzvwncv7BR6rUTiSPeG0
hHmCoKjzZcXoR97Igbr/+B5NxqeTZGlBWQQnD46EfWDK0aMd27gtuOZNYX+7Zcfn
UlB/XXCMUr4Pd+vpZOpi5TELbDfFCoiTnYFpj1Y13HUKWZWpMil0tW+QEwxrozqQ
3vbUTGVUWEdfBEErcqcVnvWfys/3p6bi+gvaIblgvOsrHCZY/uUR/vZMZTWLCHbZ
ukzBcxAmQmTGml+B6QwcRuzT+WM+UrBX+biqhaDTZ1hGQIfoGAN5zue0d2pQ/5YL
QNYBpuW6gYjOhxUXAH6XJuwa6HRD+Sv+P/xtMwoo32aJTHLW74vcwUoIzFYkfscJ
O9LZJrmX0IxABvn9i8J1h+qQWdyuuCljaVEOLFZPUGO02R/jKUCdlxgQmO0rWEFT
5hAHJdMn42HixVgG2plxkoB1gayMegbck7xwR+BVTa/wjIGOMmVqTmMfsiAa4J4y
pdO26vgJ7OAzX2nY+BkJcxVGfVFjV8IfY1B2PjCgQ7T+pI8YA0jnUqUWZw28ec7Z
MpLhxy/W/rN1Y9qfTFjxY4CdkpgZ39CTvvwik1Tn+9YNmbWGaqG3dsj268GGLw3w
wKMVPGQDvtow9OWjhq+0reifjT0O2okI0rbf3zACowruhDQa105W+VFxNWmlVmNH
Is7FABn78OIvHezHaeJE1uI5QX6kQ73K/oFzKjaN6Eo=
`protect END_PROTECTED
