`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sI5IgNWtyRywXSsfrFpR+SmLkcc3OcHDq7a0DzWlcT2Eh499YNXfIhO8+gF8o2tC
2mOm0hy7EBxxGRQZiuCQ+QJLum0uDKFSUGgVB6FME5mwHqvCb8Z2NAEACT9Doug6
TWDtFYIgGRpG+oPpPV5NGLLGShe56KhAeIChVdQpvvNHjLj1+qvKW5Kjg2WU6CwP
BYh6a5IlyZqdDOk6sTv6Rwkq0JvJmo8k8DAROqW2a2yR1CtdjXfB2uko5Te10XrV
9wLsW0+JjSO1CT5oR5NzUveu1x3R0nmDf38i6W9aYsHrfonA98YBCZeJqv42elQP
YNJmoJYpCWMmutf3oWWHIz6PHoB5n0xS6Ae9xVoXlmAB/NxHsFjCxjSYwRtMBPWp
TkHCZMazzoBAFoLC3FZDIdlSOpmu7gb2RsvGm7R2yWBP4i9CoDB1OIZ5ZAkBaefv
3ty3jErDoXNpnqbTT+tvsbPMu1m7AdeYhfaF9GTy/N7tqvCU96CnN0SyBs6Iij1o
rSMcpFLT1vyaliNPpMKrDK+QS7YxhWVh0OfiNuLGUzYUW8ebXYwy2dov29kA1GPL
82ci3aJH8lOeEAPCaUB58lNce9mX01yhesNj6X7dtXVbbhnZY7mofEWyk+X2AFm6
1HwPUnUfu/7jT1lGJ3luiCy3ZMjRdpEuTiYq0p71U2cC+bNoXNt/+W6swqq6JP0W
vo5GaKhn1ngxHut9hF8IZ9SSzk1TkTjnwKd+L9XJpc/NFln/LBs2lchtbrK9bni/
0nmmQMzvVxDlg/FmGZPZK+3clOn7HOGjybrpsPi+v0F3OjG8tX/rhetroP/lyiJv
SA9+u0nMDQThI0hyJd2T9IpiVj57FfW/0ubAlFc10nFjOc1a7jRObjCRCnRAasCa
yiEVbNiuliXBq+xUUxctfJTZLbWl3TUFJ0w+uRfsdwxpIS2+dChIjxJQj/s8jK0m
FKjK++SB2OppL6DR9RgJ88Nucuag4kmgkUj9wVIzp7zcPXKV1Q6YzPcxxfoKAi3G
O37bZ8VknY/szDzsIOesLzSTMYrSUszTgJE22EOCnjeP2GaVCPniSAaXzc6SqhNp
Cb5GNN5xNp9XvDGUd9SOMDwpeSG/agE9ElAirU8TDU2KOWKB83CrEe7l4UTB9K0y
HnTI/4xGYfmJJchtZJpjXe+h5djMLUul6pXs0RSRZZmfHlcomBzPjKTx8g/dwFka
RA+eQl7GHqCyuRUBbgOEfPzayXX03QBG8wiSrHgB+B5xcLYe6QyH36lK0sJ3KzAA
AZB6YOcI4pk2B1mnDhh3r4SR8AY/pLSmCI+2EbFZdS+riEgg64ZMSSIH+DtcYXtx
YXsjhe3uV53wLzYCIDV/FEt76eyITGvToZGFfbrQmqZyItZCVUvLUrqElhpF74MT
8D1pvb6/I/w4Q+DzyafQEKPVY+ljn5h8IwmDl1LQwPpK7+iXive4FvImJhGLrfWR
KrS4l5RtAV+/ICIZtKb8zGzXe2wlTxVNCFK55fy7fhewLgEXZWx86hCMeJ0aJkPx
+7zoNx7uKl6/RAntGSYWrUI+UkQjXau8Phgxo4K18x9cGl5T648DGUucEcEyLcsR
OejeAKoIprfQaEJCO3qGxqvmGhfpMFtNjS7zc3Za9De1qaFALKWPj6Lg2J/svn3M
mO6g8OtuN5qzka71sE4pXFjDOHFG0pkxrRxzFlzQJNogpVT3Jl9fKkEZd/XenlIw
Kgzfn55Injswdjw3VbOhADF3PJHRfrFvgtI8/WotkHrs5APdiJqQDYuMylVAxceu
ENzUTT0LDsghAiPRpkM/7fSnLwmI91Z+ODrwiv5DHj0dK3hOuJD8Zr2ZHjsMOmT+
metObiXg85cVMIMFVk1DE65AdsafmiwwlWiXgG5UalbiDOghOWBQ18SBFuhvwZV+
OTCSv5VxtZzwfSujsTFoDyJvIdeO9osoKylH7azKos2ViH2YyIU7DW/Syo/bchU3
xvTncKX8lIMnVAz3UuYneh3Gi6B3Bn1Iz2cfRmep0qiJpJruYnRmZO6GTQDqTjiG
NJNQVRuOWPCBXOpR0Q22FA5ytnKzCxSkyPtLcbgrJhDLQd4OL3gYvI/Mj5ywJYCc
8HB83XBRaEY4QemhDcI+91RT3lqtRE942JZSZcfDRkkAPZxhIUeBsPAp1BRpycjy
jEuBj0G12IS5Ml2eBmTHrb8xhCYSARPjH5xslNRF11O5dhFOj6aDL3T5p2kiUkfN
9TO2krXNK9+uXjtrSGeo7Tso5xG9rksA+aU91xk0Ic7N1LJlT6luigl+2JxTiFPC
TtOW/Tia5yndy+lusBzwLYSo801W45mhSasm2escr2xtfF9MdxLZxOPLRj7WPA4Y
RlsmRAbwGtfUvks7I9zryiRp5R6+vpKWX7CUF1epJERMbjH7zNCsSzW0STWUn8iz
6qZdhPhDgewqpv1fNBiI5iUnwtILxoX6wou1t/M6o8EMr3i7YXvnO1XNC/gLSbyE
YqG4wkCnZ716guT5coAOHxRHmQXN9lv8gURSCGYlaqGRzsR7aC4qloxO8TCD4FFC
gaDofZdZ1dmnspFM5+kUoYmJQjuV1WhIXMN9Sb+m9imOdniRhj4ELnCYdTQbp6y0
PKVOWbIeFf7alzXNroNzfSqM/dDqPNyy7qBnkU2q+W32sENoT+M7mkN0viBaGxNd
ru3yFOL1hf/BUrTnhawPiOwHFT93WKzxBFhXlGeCJRt5Hf+eK+uOMA1NY1THjD7i
rFupGaID0z5/VvbbLXp0mA8vhCEpRKKVtFK3jO2xFcBR7chHmh8+AI+wXOQDBENo
ztRxX6RzR1qdxNzb5XrGsXxQLnkCw2oRZzhuNLfXKuaBo//MnBclZsRK//MPb9xx
n9KjNn2geALQ7KzxFT3yoaYr6WJHanXy/7QvIsLxPEKCwyYDdUHqQHzskVFYQJbA
Lz1GEI6JSXg5JKy5EdYw2t6UewGomLNq5qwE51fOQELAl4FmIxWMpmgJVjAV+20A
ynv2AX8biUWkR8J0EtllFYMbOiiDXws7oDVcz/wtQsZKkiIL7ScPYClygmaQ89MM
skGIisVpm0rlejVXaO63zWi15yoVHUNikkxgloqdfPOqS30YQuagxvnznzFFosfG
tvV3CVpkBmVEiCmagdZDA8V8iHXPTCG7nHEg8lEPayNF2WmxP97efNJ20DLBvvRu
by/ZxFR1QP0x/+7SjD8G5RSGEVpPtsShAZgual2XzBxRDLT5MD49rkg+QBFBHijt
s4he5lycLGGv0ggVyXa2up2LGEAjU2N+TNYltXyNXdBN2bZHKyTgA5bkGWSauicS
nkMHJbGrIWdlYQyzMSMB5prkIqpgRcplWmlyHOANSsotxSD2nE1fBMzYtfNcJKNF
MPM9jBYzD/5BWWXqtYWXc3gGqBdQgttbO1n9Iwo2BR5ggyNCgUsSAVqIV4FXtvWJ
tE+E7YiSXYFlt6Vv0E9tpERiyZ+/JhpJCLqmmjJrUnBtve/ss8WE1vCNf7397ZV4
Yu2iQUSQaQ+bcfOzjO0pHgbx1IufbEFB3yTVE3x3M11ceCpYy50tLiFVC/9atUys
9V11I1PyfWKe7kXGry+684tC2laAcFgImJDaDEVD2rUVS5/uMiEU+qEJS1afRPm6
3Ua5NM6OOH17ElODdW4ABgwq7hKhRhbyt60bnjzUDv+jN2eBRQdEOI3sgwUkp0+2
n5vpqnarvbXfiiMTDNaFvpy6G9E+l58ZqyYNThWjGUj93BtOOMgwUJWCvwPRHAeS
nAEXKCeZVvhSQoQXbvV6yP8pMxlXJEXwuqQxhtI3EIe5roYSFU+WCcxt5pQ7Rywe
jrfgGlMmDdPuRpIElw3BAMp9Dxonw67DoJ1kXMcKSP8=
`protect END_PROTECTED
