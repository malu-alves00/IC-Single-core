`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kjJsRwjGHnXB/VRlm1dJhAKtdCT/Rf9QSYZvo6QkYQu+rq/iZJP1VP+tQZXr5byH
5y+OKEZUfnV+7Do9+6B6VHJDAj0xuj85i6cxp4D6pBQ2p6U5zYKJfMoqu5Tkx0N9
jjktNEeWxJz6S2v5WjQotDz+dSmG6Tke3EZOrm20ZdZHGmvLdcWUDoZlOsbuFVG9
yZeMji//uNnZD4aKSbYPIaq1GohnwI3ydJcTnnGvtc7Ko47zchzTmwqYurNQOjEM
vvXKUNiKvcfVsRWyhh32iRytEvM+X8zWrKDs2/uTFEL2nutuGnK6cX2xROKO7R0E
HQYbzHmK/GysiNVbI5VMG5WdJTm2BiITTkaHv1BuJVwpifEhCgdxVs9SQpgRKvRw
`protect END_PROTECTED
