`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Cw772+Fl2k2y2ipPjFfVrUB32L1WDx6yXGTfYBCfyLPe09lqHW+M92ynHxY2GfG+
fqY5jNPr+Tk6PQV961SAskOYFtS0+wPdhcMJpqOpruwaxr28/UyxS/HW3k22Mln1
fAoh1x6VTSyrqFpffFB5DHYn/B0/tV7C+nF3AIbz9VsDKUHydyY0vf9BV0+thj66
yaUsuubzY2OfTPuta3k3JcJB020XJlt7HdTwQEuCX+4szDduQiPombrqZGm7suEM
qetA/UeKVwpp9zGF9eQjq9tSVOyvRF10PUaEPANEYU0pf1ZetV/4qBqMgIE6D4Jg
PyG5fRNVDgoXaSY8OGzRWezQ/9z82XLBYXjPtJp/O4UCo0AH2KW5WQhAgkoMv+Cn
kD+3u4NsbBsBAUFXPxTig5suLFhAJnXYsDTXBZRsgzeJY4tAgADWRfJDXok2RU5a
AS59aN/2GDvlzpx6LpOCaeMDxl2CwcnKwT/yBlvnTdXvTQPkmIFLGuhh2/ueEyi0
BvQ/b3Dt9bQjPEWWpffciQ9NC3m7T9934DURgZXouI8BiKbAiBpEwapwMHymd7lP
auyxIacJPWXF2Lpadz7W1MyWmNupnbnSmhMSdMevqkzFML8sLZ3K59YK8v0NBUMh
i1w89k2hH0fyOg47uZ5ggLr9kYY8FEGfuDFnOrhfCr/77h0NLakVaXcnyQCNm6sC
0I2ikMHJ5q8RLfv+eACQT0RPuo51snpYRn55lIMdbA8e/GvAjafgj5oZ/1CVdnqx
fvtupHkKJaE7RqaKuwabNFG535klbivAwkuLnfS05VCwO23s97oIlzA3rghDtK7s
v5lcUwAqDYDXkhRb7/RMvbCWw6Ly/n8XM921cxNPj2COjQPPA7UH+4bjoXujr/hw
yf9Ttb/FcO5nzCv832HXTlVletdQ9EmxrCSXsYzJ7u82yHarex+L9Pi2DGqLvX2/
NcXrDX+aO7bIlCqBAYXQuBAVVBTuxZ1ZvbFsALK4/TJPKrpFaCD3n9pl7t80W5B2
A/FFp0MS8KpO7jkWBpwhcC6xk+7Ka7OPCaxcXk9COhn4U6uRbsJmoZPmsb+jRSsv
muMxYwRPCjL7vmUW62kKYVFRVtxiB+VKJdsc74VrAlelV7jJ9ekQJ9L5SkX4s1uj
lKBX1DwK6CYX0lL+bomhVNA2gEAfy4bqhtwzpUnOCEsBxvyL4NYdS8eIR0r+BdNh
TjPVw7Rlm2BoeWYKu2Ysi2NmbCacIsy5OvdtOTXAhLU=
`protect END_PROTECTED
