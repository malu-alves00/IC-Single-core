`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UPYu4F0OJaw+pbGZ53aixIxMJqLG5z31CKdNyerbXxJKpgmYgNHuRbEjuYPl9r4p
b82iYtwev+pl4R+C3CynX7D85NCt7AaPvQkVHi2UfDMlxPjtHBOfV6MqvAsBBCln
VhFYUtx9AqqVVL/gfgDwXkriHUuU24556AbfM/59kAZcE64xT1w3GiLshGyUJcNr
7yh1Lcy6sKfU1oHwT8kKkPUFYkBMqZiuwm4qtUbFm6AG1SCI4i7Y4mLpbCrmH9sU
i7figrqEdND2fycen1CA4b4Bv2L/6bR5DtzCFKq4CT3g3qjX5lT38KbWpmFxpm1Z
IaVyyYV2qqD+R3aRXskEURmT1Ciir0ztFM2bhyiDXXVivqpLaBtVNIGLDwUDnBwd
jMgrSrGfqBJjBXbrRgDfCHh2IYMURgXHUWZHf1IxwiZ0Qxa943kJIcv3Bf6+Nfo3
PQg9jGUAN6lXeTHb88dDLkQqvkmy9ni8FDWZa0vtiFp/pu2HQwRSOxb1ivuOI1Ha
BN0we5lPvEibt3kSy8TOtAmfgfbODLdYikeE8Ch/pd09GIWMw6Uu6oOBRjYLXcId
7DOj33K+Ymo3YU23zZdiROKG72Afl8b5MpcwetxzS+z73FzJPZ2B0jwXJanogpAJ
L2XIGJOMbNFSPVS53IR9z8trlZUeYv9hF8FlQZBCoDvi2NTM18FqjE9/NnLhhAn/
hHOVwlOTiLVJYsBAz/pyum5ka6gZy0dZJ+Tsrw56aCO0fAAdCeWIfNNWyeqtyTtI
B/wZcyAndX0Gz89iSo00esHG55vtWJo4/wQr9s443vVvzumUm/q6mf2yAZo1iqzq
KZcHOgHGi+amdDFdbMDf71QghGKoVjT8xyEsbVyakDOn0/VlXJfz+bv9WG6qDwDC
RMb0N38iR44i8tpn5aQJ9oQAfg8fCTc8ZuSnBk8wcZTcNgWJe7M7IO8w5SCZm10V
T8NXQCT1ZyeJppymhf+0E/y8bOmi5WeOaOFl2sE/1YibD/yRul5oIvWko+3sfN17
sEhtgHadw3RpdWiIZgUFgFNyhd1nyTKsl3FZTyaM3uM9ic6WTJE+2waITkDbUO12
BWlNIeLast7jagxzKO9F8VR8xgfAHg6pZ0AW1vY/TkHCbVTnolUgJiHQlgIKfddm
qFl21pZUHif3R9bXY3QVZI/BqjAGqg7TszY2mNqK7ckULbYdvbWpcmlq4mb5vZ0g
J7P4X4y4Q+Y6YbJHiVwN5Vme6iK8ykyLf2MxN0jex2p8YrxXCFg+S89/p3wL/4qX
KBSPKEYIzuGSnD0Oe46H6GuCU5M4My+LhW52j93+6WjITYw9FRI1p3zCsY1I1H+C
lEqjhyuZLyo1SfMbd7Pe3XfvIWpNLHp6vW7l6tL7rHFTfxk736Uk2e+amjjSm7bg
rZXHpat0lQMv081j7ChBed0sx8oiwqwoR9uknPKrtxcrEaBP765WpZHIcXqF3qkB
d4wH4fBwd3V12peK87OZUqxBv1VipJ6xdBbx0d32kpw0UxevSieRX1Y2mA2JN3XX
iZqE0jyUnj9Q6i/PCWQY5FDnbZXNBFKPRjz5oBLnlf6zrjMzTzPz0k9QI2tJzrce
gfNlRIPBUuXzS0+9wQlgqn3iT9kzR2EyQOcOsbRZ4Oz4ES4rBQST1uv7LV+A0QlV
yWmbsTJDp1nFw7Y3NzOMpsGghElZo4AupE1LQl6JiF2SehFRRfNACg3qxI5c7GDH
Xk69hV83MGvbtIaBTdeJhptS7buCafonN2LBFSVTks2x49dMCUkg1vy6e9Bc4Bx2
rf0V/Q3gRId8jbBBnIxfsKar5voKjg0ABf8sEkiSFh0xJwPJ4VuDboIJlxC5LtLz
Q12Fr32vHlh3nfolE2obPfFSlIt7ZgeP0LZMj5X5/wyZs8ptepQklDQ6e2aS8ykp
ibPuDWCX3kGL6l5ZYB5hZ0+NlQuZN5zZfJrTaUvsrYkFxaSfGXBGNIGa7jJ+l9qw
85FXBjxxiXcHwwi+aVN/lRpg8niCCHEuOirHJ40s+DDY91+WDm1makgAFsldU/+7
y4mOcqHXaG6ikNVInyxIII8yapGuJ7jlC7cHjAa6h7GABCLWwlo4Cqu6i3DFnQfu
axgjPqhcENjFlP9RSD7/ts4zw5neVLmrnIHoYL3E0npdOq2Mwll4LBW9FTTONgIU
1x5yxZKGUjjWTbSDudLsF9NsDuuHYy47EulRWAHksG5hCEplXDDJdvf4YK8gkGOw
yUHgOehbOBkJcXCKeW5N4DMaStpcIeWUzxTHcDlF/f95dTPXcv4Pt596RimWhBU+
y+OfHPux+4ZDAkBYxBtrBKC8l+o0cQvdX4WFMlh+7DkvNly2ceK+lPqrA0Z0M08z
xgD3XCAEj+dwpT54DnGR9BocBqxsYIN7gNWEUaHICnEDhn5WzCG4XS0UqV12LUub
tAwdzBkzIRInhwKrkOFvB+6BprK210+9u4c5uK9Q5X4EIIwKGHtsbkrYEjXY79Xk
ESvpS4B6W37J2wEMLsEDBPLBE9J7FOjn9Q8IejAKb/IPGmYH9k6rPfZ47eEYkub/
7IKsjvP/14e3q/6gRbpzumU29Th/r9YGDPFysYo25dNuNmFI8sjrM7+/97lWY6nP
km6cexKAthf6rlbJ+yBedqd9P21LWs3ZlQxd+6lDHiRPJocezvcYgdHTZlbhPT8o
cOcUPpyad5ps47Zn4B1BKEfwny7ThV3vYQQR2WoNXeP0SBkVNwFMAGNJO+WDeXDG
9EHE3yd+O9LFmBt0PMaDAAgq4j5GBds7ogsqiGKtDQ3D/5yNWGzW3KrGf6a0mwO3
JY+XIRXrY8dgRyEEcdxDeMfnOlEEZfGQ0PBeiN9GcP30aqtwziekyzH5azu38eZc
62gQAhUX0mklU1DTsRqVViZEBiYIcT1w9sDHXYQf6yz6JHxRfM18jmcGVtGcPYTz
VsCk6JOoz9c1Yb6psv4x+WUk/BcpRWoL1Gl19+G24G7UC8JO3HaT4FggJ+r802jV
B5s/RILOqM3zZjAqaKC8gQ95Lwg1X1aiclRD1JB1HpO3yCGGtS0VFkyIM7bvrZUQ
QeEkn8UVfs9dRe4RTQkiBB1gRMn3slPdVFVzs5/eMhPv4rfLbQ9fyrvi0DBouhgL
CGHRFQrrsANg7LhT2ABFfhU8hKc9/4cfY1nHc9YWrIEo35J7f8jIeFxGDgPdm3Dz
hBbRTGdo1QoAVo50/P4IxKsZkuy2STPi5UlxxXCuUv+/2mOC/R85SiiGNde7P+22
w2kkYZX5Hs57q77mi22+sI+DnYt3+LdPa2dBx6GuCzavm7YvnPq5AplwODcu0uW3
wBdmRFoxsqYAqGMwIK91jbUrcAKHyRm1K3Vw/PICn50HaLjkC90b0GWbTw1JLX1A
+CiSIb0ElXdVTt1MEEVXA0ns154WDK3b3fJbhwG73A1Cp0EGTx/1hCptpiuHdkTa
WQpIUfWlOocpA0pep2hQ4OeWjYC7U2cP8H3nNvI6VDgAH4ZjHYa/jFgj8slHyUQv
zoNa+Vno3+D/czFztBKrqJnHb/6ku7Hk0mxdszQPtiHo11YjdBGEaHzNDcU8/ft9
3Y0hBTRuD3HU5DvRu0+HrdKDN7Co5OCAiNRQEH7SMvKi2mY35eM0GLRtuz9bU0ak
YAvvmI0PIzHm7oUAJ4shzMdcKT9Ij530D08Bg0G/H9hiL0mM89heDvsfPLR0lANt
olHk95iof1x4LUzMjA1XfQyO9QNJa5bBcyMweYRuHlnjJ9C7xLZSWpztPiOuc75w
JU4EUqrm4AieO3jlChxrnw9kmpQsMJoFt0Wjd8L2MbC1bU8euhvlj/BxLhyBQWiM
5TaYIjgGZWUsj5OEfcLhblya26uuQJFCy17hiaZPt12sxk4wYm1P2qK7oUbun8gx
lzf+7kciMZiuoESjZndESiEx270CQTi5bK8nvmBjLrTEliThHgCAApW+AgLQrvBq
7QVbO+ckHNUzJghSCn/6ejCvhzv6MrtT0cHuS3MM9fVD/tMhkHjwXawn1KL1GKgs
VAPRiZESG3w6mFo/Ifw2DZuXdYSLzhj4N2fSiTmVVdaNn/PJdHcC0+j4kEGzDaQe
2MmUHLx77IUcyx/wJWvZqGW8z0Rr7g0SDvF9GesbBF3F3j4Q62YEaYcGYsvMMPVY
L0memy018Dcoza80xX27FflQtbVUkByD17ZyDqtSI7+I+erpewScg3EHfSLw8K1h
YvBWkp0KQMflGClIZ8UR2UFSMJNKGQTM849vd0y08eWZTemSWYAH+KymgkMLTskT
qOtIwWGdehslzQv/Arz3fAfTJRiye2fBzQyuAFDir6MWn+EcbC256Crdruasf9zk
L5mRe/QJjsm1YmCAqlehBzf0W/hGKGAYuQEaBO7kp9KaKWtNUdxSvQjKzehdPD10
Rg6g9RRpzn6b3tSk2/OdeLHsNXCPOffvF95O1zPOIfN1wll4PtkD7zHRe4eI4a6b
`protect END_PROTECTED
