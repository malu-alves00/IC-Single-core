`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+b5MC/5rNO8HfmdF3qJ0X9pkHX9o3C22UvmVcD9BcmhH3BFgo1hiZyz+SrNb1UTy
+u398X9l7NlISR0AM+x0ZhL4AuzLsU3MnxwcZLTDL1Ia/fmmFDkHLiHxYbOTCh+8
BeIBelJVEQ3p225BSi+0LJEJbXMEflxKm9hOOer399wdWbczHV5qnzfZDIu/SeSo
P4IHjzCpZ5RYupLqCdDQALMoZY9n51goIdUpf5/PSHCYSFT4ZlstpUmhYwt5FZZy
tQEV94wrasEB7+8sueoAG4d/aiJOp7KWNq3+OuVXNz3HvGqYRRTmEmXQETbJw9bK
8X9PtIgZd7QQUF7e/ixo4xrfvKcvygrFmZ8JMqCxczvCij45tq+LmH2XVMEzZzq+
jwwrQYqKHfLMnHk7Zyfmbdqt5mwd7+E7v8jJz5qc9I4aNJChpfF/85+D9hfepIus
XfLlXiOsXNNOsgGZ/L6ic31PueqaNctqX9Ee8/RRXAKC1Oh4MiRogJwiwus04i4p
tRzq2HY03QJ1jC1EJ6aVvNDzclx+jAqsHigLEzdNoW3/MBsu+2b1/YobjTVTd+YK
zWbSZ9Kun/7NAcaDdfpW6wyp15ipWTo+3P7X58y77hkuMV4E+caQtRDpEr1+EGT1
naXMKNu/ooE2tJdebjnjfDuB9slCQqiZ4Gjads67Ix6KTtRUtjs5WUIsMzmVxvGq
1Acs37ma74D+jnOeHgLxsws7W69AYhILPkQftbZbFOBO3U44OHEGuAW8onVXjRCk
456GEfgbJW8ivWesMfi2WKgmJ43N96YCwSkMG6DhacqnViUgdTk2VOu3T/A/5gG7
KuqIroxgtHrms+DYeGiVywhDcg1thv4xKyV+AKDussXI/KHDRmF7K3lxk7kOuJ1B
Uu/xWTH/BeD2n+P8b52rBP3XQ/Oru3SNztDbZubUtK2a736vJN2F+AhDJCPwCUWd
6H586qgtrOmVF3TFRwe9y7IOfO+AvhewGxaPC9ODb++jsRBDAnRBc+p5n/upUT7+
eveyyRf1B8okOD2XFqykMkISPXiUS8t64VuDmzcus/LwM50PpOgeR4m06ULgdXM4
fzvcDg4Hr1ljdoYrVlxykY84e1XZSTdznXhM7ll8zlK6z3umbJZ9Lp6LHagy7u9y
3ALWjfptMFafU21xKNhjuEPKjsdDko9gaKeAcYYlzDP66BO9uozVzn9pizkbRnI2
wydhDBTTyX3Qv15zIEoGD6FTG7NouBeLoWQrKxB8yEbgzb/NWCy5ci3+56QQwsrq
e9NpfHU1Ah15sEZOEHDi69f2phCqwY7vdEYV+hUQhnZLGvFqKrxUyQGtZ+Tz8R8s
qb7a10G08UlXaOClyQYlvHikYyqMNONxRKnk+PJfjbflSe1x38ZRzW4z7N1R2/Md
ieIMGGWjdpnMTaISEZv8Va9XHHwuU8F9dXGCfL3FOe59mttKdb5iBXSiRYgZN+j4
cJP0lVjGF8GU++T3Y/wdO4PhR6BwPnjka28w5KVqpcvljiJr9blg/yWb46YNu4v0
Ij7pPpvSakP6WSxyxUiuFZmXU916YvizSf0MImqiQtRzOWdNabmA87LnE35zS0Ar
uE2dyFqeQEioyM9hEmMyVmJsVDlGXMJeRBxuSqGDAbrhJu+8hFxGrYEbugOyK35/
6GJ7tOX3BWqZ7GzY0BA330D+Qt/OnQH6+45Had8lPZ0v5S6DS4tFc24FKq8iscgW
J4t7ofgzGEgPI1V6w8TCqxtY/iMY20+roCTs3Of+VAyjn0TqYfFPWQjMxSyWYJH+
g+W7MeOX5xOOT5wiXer8Wxwpl2dhnQ5Ew8eyqyOhRMgx2xnW1pWK8jn50Jl8j51r
ZmR3QglOEZKMoC14K1KNLU+Rwyki5EYeE6BvnbyoGtcYcUZcrt7935pk93D8juHY
dywcXMvbUekNXx7xPY5CFTiB+9tnmGBNw14j11tzc73KFffJ1VUhmmvfiGcKRtQG
57dbRjDCLJAPEkXwKh1vyG2oUKuKXGavGldrUREkKXwbjeIxfPyHRog+vfRe4uhR
2Ckn3Zg96cuz1e/S/TY6Vw==
`protect END_PROTECTED
