`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bhPflD8/+f+N00r8V094qk7RsACvSJOn/AzpLpEbZFzhT/gAeIJzJYjLJAHnIp2R
tNQCkCK0FjZjiN1XPH4EToPqEw6DBhtDTfEOuvlSzp0FETDkB3pZJk8qFtH6ouy8
Sk4mfK8mFSM2YxJy0TvRR/g6+D9CTCwu1gd8WK0DUB42hLyhJNK+9VcKiopUG5cm
9zD4GxTdb5EMYgEX5mz042LxZ2QcAx0EgKwP9Dvn/1yWFCZ+YV+Yar301tJk7GYX
MG7WRm2+iNxIO9wO5fD3ADt4ywztV5eGlLMgh15Co2hTeEJgN9mxuA5sohr9Fal7
UD+R8rOG8pUZlutfHh5z6KM/ivbB6Z7rZq2YS1JFwrAQze+KUxwfta5lmY9iRI0h
GKeJSQjnvFu43rvHAlxnoUX8oWvMbQKYWw5/T3jdWm76S6tV1DcJ5FJ+zrRHCtm3
DO9/lwiOb5pNbasW9csjeRbh3J6J77b2gaBtwK7g8co78sodGtkHLjcmaPHZ0nXn
+jWJzQUYCE546hJuA13WNkQCC2OHAMK2il/1xVpY4CF7ROMHxl7Xjgj29Mw8q//D
hzIcYvugH14+CyJCeSI7F403zEd1B4eRbSr/fxdpqjih9Dr+OpWiB0VM03V9dzYs
fwpUf6ee2HoJQ2yATUB2mAC8724/DEFNhBo3MdbbELWvvy8ZPHTHO/EDp6yqHO9k
nY78Sxx3jHS3SVpdoZ+zFUOP+R7cPLTK93NRsMd/5SzKw5pRJkbWDZOXOEfyqLZ+
T0mgdK296NmOPzmxvoh1sWb3cTyhItNNRna9hANUY+qTmlP2Z/skoRzd0liDM9+9
HoBZP2Conld3Os8hUohm9BRbYXBhc0eF2p3Q1JHqUJxiJmo37/pAjZwrwN6zfNdn
I6wsNrKw3EVt282+FgWrHEAkp2gGjWPZacaV7OztgusBM8t/+WoKKcytf/sIZD/l
TbqG+QEuw1lZ1nrABUmmE9y1fiXufDLSINnf20XqNkgN3oWX8ii6a80gTptpNpAP
owwXiJgc3ArFkp1HwJ8u4Uib9UjsCJUd4AWcN/ApcLNz7saBxqiKXRkGfI4vCpkK
5Zfg15qVJG8ahvT9EIkrgFNByhwgh1IrcHNeMFxt7/68IoJBmjQV7EqzzbN+LXDI
TTPPydYNvyAnjCYQnsKn67WQ6wMWRduZ9fWwqiR2zzuPSo+ern8/RK2Y/DsxNv9/
4qiw/nb1XxWwn7j1D5QEnlNMq76pid2GX/6m8u4ins1p0BIJisIIlgR6R9keJul/
r6uE5i1NoXKqJD6sY+EIUMLU8P+KjaX3wU9gvwuB17r5P3c75zLXKP3DurOtHbbt
Fx8iGTfeHx4WKgJnAS6oH12w2r/JNSYBQPO0qeBrCUaQai3S9PFeF5FX8wQ5pvEF
`protect END_PROTECTED
