`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GH7ttO7TMw4Rrd1wqHPQ+1podUWKpIzvK3SmJcLhyrPVl/PA6AzpG/Yk8jj+l/BE
sKwVveRwrC6PzNDuhQSsqqI4ry/3y0L1jZ/RHDSvqABpVuwITBbz+gdbx1uqDIcS
GEPaWdC7gs+TvXg11vc4RYBiwe9W2SKwJRsbkuSVX91y3XC220KX2GF1vj8eQxGE
WyZ+2vurP40ENPtd6epqHlg0mKkD4WxB1VPlsFFNbqhgpRRbKpe/sXUZY47oUgZ4
EO1JXu7ggXhdKKnghm87P9HPOn1On+kPzPYZreF8H5vBcU5LP+qGHiUS+c/HBIxN
3LHRsP2VX79/WCdiuxR98HwWYv0xnBLrMLrufcd0IjzOo+0fxClemTaUhjXUQIW7
LMe8kLQRElM/Q82KOwihYQ87FgDY2GM3Akya312mu3GHs2vX4ahdAPxVdZAMRsh3
VPxQ+xxb8eUcOJWAOefPdId8ly1+QcNISDrtI9nJ99vVSNcj/PNsyfOpkfV9DEJE
pn0T78s9ml/Gr/PWKHF1t6cL3FT2bQogotCa7fd1HgY3rI8tHNVkLpBBE9fFonO7
MI9eTslz1lL4Pd8nBIVQy2mh0cZm0ULnSAyweh7ZgnWQOTrtP4+DICD9RZXAv6sS
rFNstHA9KR93LwShGPzmaUPn9+Rb+kevvqnlJUFxyqGfxPWNWcwqsySImKXzBw5p
KgdVrZQKvUi24nl5br9vIU1fJCILvPAj/5tPBD4SIcXz4BQOQ/L5UGje0n3NXm7m
vcQwLUgWZbJI2EuuO+ZyxR64LkD8OWd1rnIm7aS/yezX7gVv5JmOlN5/WoK/JbI+
tpZFx67QfNRQBN2OdQk4jKslNM879BFEdzmkrGBIFx6nDHAMdkjPTjokCTXuh6U5
2ZK5w1pZpyr0j25NXXiyXKdbRZB56RHoR1nQOcxVqRg37sDZbZGg713ufW16g/Rr
GHHffjkghGcC7Gx75ph7cp6SieK7ewjQNk1ZsVfO3WvMPB3pfMXJO05nuR3gA7bq
ihZDSxpMnJiOYPySmvlI4EEDAJy9pwDAFh6Yavvt/XJHbhf8jw1Ruw/C23tRK11s
c9MMTbj9dXWj4DFVfXrBI+CktUeweTR5m8bzxVlrBBmvi4vHW2RbX1uNStY+N5IY
QL4ZYpnhWofXNHoiiB4CCHh9wqwudDkA9YwgIeKs0jY2HFh5qX+rawG2wsHbPrIq
qEeUwwIO887ifQ9TcftPlXYRGrWLquJ4awJky32fkkLDLQg+7g3qLyH0WxShA+py
4kFapyDmEn9DsB5z1c924Bg0dshlhaIw/2UbZCCkN581IzHM9v9yG5INuV9ioV3q
nBV5h2P2fC5+NoD64t1rOEHitzeHd25Y/1EGT+clp8N9befQI7A0/WXkKvGiQbUo
eilpYJT8UPzVUBn4LbjpZk8XnMWFwnuK3LQbqJ+ipgaZc21XcEty3qto81RTNMpG
gHxEDeYFBaF1YOw7eqgKX7M8E3QBHFa/tIcIKudbvA/NOQ1kfM9eHQ4om4tq9+X4
5EV4jQDCYMrSV7Pc3zROMG9EBsknJ90qL1u2YCKE/o1tQEViTNnjPEdyCWN//LiP
b0rJ3ldfgqDdmYBodOxJbbIByWzvyZIz0aInoOOa+uXgpoCu40AksuWfX8mTLiW2
2HmCaoILhOzZUKLXQ6982V2eR46kfiasMHIyNTdYp7FJzw2ghFfMNty1JCtCLLUQ
NVbJ32CtS/HDNzblndyc4eMWxKUNlkdVs3P2dRtUX1kNUQ09j/7LnOci/nYF/+Xu
s9LfKwbeiMqYRLK4TrRBijnmT5w6n4bc5Ax7f+Op2bLMuFlMeJQRMTtHm6mnsS4K
ol5WyT9nAtfSTIFfs4dWCXdGBhBLFFMwCi8O+jTu9zeIqHOK4jqhBRYZfldA8Zcl
xclSJLcIu9ElhswaWRVdmHUVgFUtq42uYFtjYbLbjzHcoJU+P25BrIHRSI2HzwCi
lplamaUwgWM1dwi4qCHNeV1DGNKMTMcpxyTA4yR9TK+DpsxGZTLyjVTb0uuL8f5Y
s5p3YZc6+qvzEvNrY4WyTo+qOTPUdZ6b8eZjA0SNi4Xjza7p21sAUChJR7z/+T2I
5BG2sKxmtqlSRyv3N48WA6ssm+66YvupAfc5n0omUJjgY/Q+MDS2gFg7DZIg5lhD
IHCzpnkvu2dM17f39Yg+AzAHgSeQyXpnAlGuaeI6mdQIraOqn8BVrAU5qNPoQFfq
32VNAxXdwIQ1FS9XdjquqY3lfrxf3zL8z6njS7nIBgKLF9OCEA2SLZqX+D0UotyV
+Ee58zlIiHNWfQGZguBGAa+Afo05F57F9BT9Y12ewiS2Rr/dDPnHURRDq2e8fAza
Oky3z3fN0rT3NHOR23shXmEINSB8Yt/z0GWdI2EIziWyUvtahvJV1+YC2kSl7Tej
9+wYVZWwdBNuypHO17M7ylKjvfGGWi1jJK+LAg0OqtLkWMbJTgxuJM5ONSHA0UM2
1cq8/H2Enduel9Eo+dEMQnRK700h1RUWyVCuUlp+Sg+P9BWJWAVAemIEcE0a0Rcy
6hm+0lN/KhGetFNpSitoAT4mDoLgt7bfrWJqFTjTHCpkDU49xZbqSZDcVGA+MkFI
gS5GiZFz/n6m4eSPUws2DMURU0CK+VB8JAfistGFOic2fJ4bKgvuy6Ox2pTbsyEZ
gngWJmlYOmfyE5i4TRNMdGLp6kTFFJUswn7qwT626vM4WbuWbOZoUV2FdCS4KG7/
UqNTucLdno96YHsUAZrUuNmrCtTWWOEcYvncZ5VNraaNWi6GFbIBmCYbm3TfAWvB
tWwwVfu/XylpgplBgwLt9kCdyCM9VrzihY/ige9E8j1nbTgL8cc7qdDolHKUXv7V
paKHutC6g3BPo2vqUVVru8M0Wb3S6sFPLuo0Ke3LC0nQpEqqYV0wqRdT3W1nL8B9
/a4lI2HOSXslctHBEoIpXZfhZE3n+31f5p0Rgkv2s7qXEIc194mzJGk3zKHb44uy
ZarEp+SQzJqMLcA+1mR6YR4h+/N+T695Cp2vQs3MPIeF4cjZN0I9cb56Ux4LN4eh
7+dtQSlX3tgL5fRHXFPjB2gRKbmC5yiJKfRw+vEbD6eE8zfQ2Oq1T+SZVBCDbB94
6XPjBD14Rx7Uy2kNbdsNzeoKomeU1CHVgBG15nVRiwe90R3xm+raqbbi4MARgQ9/
IZo9j3Z2uV6K5zOnPoOD0xY2U8GH2Wfxa83iHXVSVrVm+AmjvE1WCqBDLPPCFc/p
7WmlY0pntifF5AGVfMUJBjv/ZxUJPrzPo2LuqcIIFhiW1tyU70eDkgAAZc+zFvx8
YniYlHjy/pPjttUg9qKUFL4N1173Pbo48I8moBmYQN1bcIY6r304co6zblOqX/eD
7mFBiGOn/SHAvVVfmZj/o9tyWoD+at7fjo7HKuguzWOAvDENoUjVO1dTlhjCoH76
XcuVKvMP4Yk+gIRF+1UNwba+M1J9b7B7tulO1qnKytja69iJoaxIlulQxeVvW61s
v88onKMV1Zru0Bfe+zLSsln6hCkKHPw3WtiFCw8IvqP387KocI+eHBvbyZQNNYR5
9c3/SNR8685lZwGIvc72K3bgPH32YV/9bRrUfJFNShxI4fHtziD2nEh/ZFT9zeRi
JfcDLJbL2PQjw+zWlZtMl2k9J1+bMRdBF3igzMf2yzC9rQrGgXjaJ2PRnDWS8/wl
HJzRTAK9fflSscFw1T6vnJL0SQF7arROl+RyeMOS1DjkZU1F2iJZQJCLbzdN6UhM
ViXZr3J0QGxrrr3+MO39JNhutfoulpt3Y5tkbR8qxYHwcYaM2hhXphhNmgBJKAOK
tBt9PbPRBXC7E8Np9KDAscPbf8TGn+nOr6wz08rwxcM95YfZCwBW7OoRhqe2PWsw
bqbLydiNdGJz3Yc6eAltEZgq4O0x24iaTxTx2ktoJ17FmF5ZDZK0g3OC52jFeiHN
k7HHxWjcZDUdnSBoelUicUBQsTc/AAPfLH1LyhtF3f/pWbhBDcR0EM6p8CPMe8lL
IUJBR7wTWvPzYoXy97s06FhLvtrHgteWSD2DpDpT68dUih11qYWH0boA3bKsKFVm
NWISUDh44a+8uaBtrAY6JTO5i8yWLPUZaDVl8FSJyyB0xqrDxYWETA4TkhCOEGcS
VCGJY2bArfaenKk/ovS+/YYgqnN2MlGC5vLJs4zKeWrHMItsZDJtZpJxJhHFm1P6
126nVdtN5iGIcFM2Ql7TWw3gEP97F9KwBs/WyeINOrkcipgjvKgG7pqHea0duB2P
VZgoIpBEK1/zcc0S50HEJ6+RvTJhxEd5cZgZuvzDL3IemRhFuWX1v1CK5cEQ0d9Z
ArIWioMwVvByLlXpP5JsU+Ka9tFfoSiaNi51A315VNNPlWyUdXUgQqDekueuptbN
KlT7NLWdftBXz/AcgwtFSeAejDr/V8OuNNBTiw2VlSblpVegb0zFlFViqb7SuOi5
1S/E/cwTRIboY1ZG8+pz7ItiQ8D+OcBD5EeXKWrKn/DLEofWcuna0S8gi4tFqriO
/xH0PuGRcUP6cPKCUiEq22K0AnZvi7miU9UzBr12mWdwTWNYjuOplnzK20ppCBrr
1oGHDKwpq9nG0TqGuBAPmosTu4H+sVfFIGnLbTOify6kYfZbrMbk8fWCo5arSiQd
hh+1eCnDCocTKXaOToFPtxV1Budd1NTnnIjMYWrEEYhDW5hitAPfiSLA+OjwrOHj
szyRB9Ii3CxVCA0XKQ4ubWLehtQLnmvYlS53Vg6hvo9zYHomICYogZb4uiEnBlJL
r+n4ix/3q8lqtp6JxksX4vmAQBzc31qbUEjWYsg/qX/NA7kyogmB3G9+9dFGpA9A
Y6k6AR1e5jk2Qak22wTBx6h0Ux5SzC+tg5fF+KDTHLirGQXyP+y/zu89ZCjgGcYQ
si/Djc4DTXvFqlwHsH81lLWjhURVuW/Hc5ZAy6NFa/UzNir0frVJbRxiNSBE80DN
lWQOfgYPq5N5TkzrhuVnWjsByyoJ3uh13SvvaR89w148sSd5EXm/paR+a+75jlhG
vch/QfOxlPq2T5szWNW3Fd1UKdxxBvtCYlb/A9mamHTloRcUsvMHlMIsWHgrIcLt
zzDtiZHBq9uoQt7AonFsj4h1kex5Hc1DXPPTRgcyFDsglpiR+MhxsKUtWmtCDJlu
iJl+swN/dTWeKX/JTQjN8ocFfzjNQiAG5vXFZoIJ0ByRZSH0gPHiiELIbm5XSYd/
vOPM0MEDRFH/D8h3IEjwCVZnTcE8KRmM/a8+EKFli4w02KVLtcEOraa3BGElGrk9
BgdKZgBdrbecbO+eY0CO1GHxvoMB3fzQisABD2WHHCr01BsCNyPoA8Xo79OYxucI
v3ADe7pX1qHBW19y43hxieuSOObvoX+m1OCqYH4TAEJb2e9hA7jFm1nqyfSCXDJL
6pt6T6dWr31BJSQ7do5+fht2U8V2mbgZpenX+qHMsSBFonxFBMR4PfETZNiNap0u
KIS/m5eHYV79Jy93hZqkuG3mVW2pdOR4DuzQ5lQhZwanbl2gNlt1OfQbpWJ6tWYL
cHP19HBj9uN2QeVd1tKxXTj5079LMApcFUjifP/FmsGCjnxui7CY4np97CQkEBmd
F1mh1/jhTozdl1dQkRx/+AT9JfUnFXUnzCmkJBQU13fcDr00RwwGcivU2TtE2NU+
MWMsTwkmgUPFP0HgSNy7E3NlwJpeRaIDrMRVtbuzJdvGwWgfLUs4FGqLUdt10kY+
O8OOpjd00fOsrJJtZWn3WPyBAPJdyCNwEz05mh6SA/lQlfuZRyW29VqpcZ6e/MoN
hdWWubY4crR7HV5abTmccFGvoEefDXkicqNrHXyPBRP0PfW5+Qfz+ZwNfiCVTNEi
T1HfDV+38kQxnZlP4DW4qeCG8TzwG4qaBz4ERWdnhW+d3L2yd3O2hX695DM1dS1U
w/HucNvN8R09FwdhxoEz6dv0r2F8+yINsJIT4JWdjeMMdCQjFxQfu7QOKxl72+bD
qoFPiXFAYx1QCccFb7usqdcoBglC7amAJYaXl4BJUgZmGitQ1I84kGevrBBWxPVS
ZMq53F3AzciK0ttLNYxKd0OYfKWEzAAqyEAYdWhGSc5YvumaL61i51L8XkBPj3QU
4lpL5CLOvaHL+sxInElSruIXm4RbExiq6uDUyy4IBmAQkqcNVFsBkzt/RznkZAF9
zKB1ppwPXyVe5kaLUCVAY3/8+TO9V7tgVA21E4DFIlidmYoaVNpPj20Xq3sraPII
PAQ6TI6ls+RHsOvFJ6UslNn5ZlGVYb7rqgBhroiaffLYpl2rm/Q6STHu3dQpUKkD
2bN5J3mBHQqsehviiiVB3W3Ja2n2QUptxqo15gYFLw7Ht0DYQNZbHOqOqld3Rs9k
ZII2Mt4uUQBOkyDxOfyKUklwLRXfuWxFmQKtfJjTl8UNqke5PlwgEBI9zN9h72gd
gAoDTMeQzlgOeIAKBz3Tzc2oR4FGZnuJK58Ot7R2YFZW8YHUS+S0DN48b1Xpz1kI
s//N+/CzW89qkwdzDNzqoEpev86dKPpMbt+ieUrOgXVLv80kAH1LOVaCdQxqJtTD
X/QA4hFRpyb9RZbhRhekN80pqMl1ckN/F6g1mOn7Icvd0jkxlljw4mANGpA//r5w
alBto74XQsjKBToppecPZlV1POXMDJZ52ovCOWsXL2o62q14sWRdOfgINrv5S20J
vBtTpWI5pzhzM3SGEjbsqZ3YfCEs7YR56H4HnxwxMW0yzJaq9+ObL6wyQyOOwWqo
jK61V+c9SgLX8Pfpv7PzvxsJwcXtpiWrQaf9etgYw8CJK70fpHyl9g5aNL0EoR2T
EIc5BcMCUQ7Zu2VxnovBCp56sJx6Txot/r02xuvjTotmG9OCWuisZWTOmF4/GHon
BehkmCQ1InHnT3/OSsdNxl5E73/zsWhuNMAclpCLqr4CYgjlyCkXPYnWNRy44G1n
g5bmKtbAnT3e9t4BpZSBkodYmUpKZvA/O1I/L78M0izM4LjVUEESyyGe3jOQnh4n
uqH2EPKzuac3TTCi0JzPhDkPa3CXn/OdSak5qrE7GRzNZ9Qz4oZNP+n5VERVGWg0
xNXksJFF1J5lwVTHJhQFCsdCY9dZyPV/ez/Py0iPb0H2wGNQdeJ/06YiwY4582Eg
VoNCu3N92wxXqI/AtT4Mu7zPiHOHY11P25RQcr2La7DNt8zxCJIaiPA37Lh3ac+1
hSyOhBnrsajpr+GYkhXu7tcm/S/N0XSvOaD6G6IEVhMgLDz7a2dWWdjc85fDcWBI
YIGs+f+yGpq3zSQtGtLAZqqMVpROdmdKYI/PZLCVepjEudjBoKreybiIXA5Itiub
8lr5YNU9GcuClkg2Moe+gX4A7H2gE65PiMHkm73630zeXb1jFtLh+b7B1GO8tLQ9
3lv/dFGRaJcrvQ+s9TwcfhU9iPFJr2W/IboyrBeZwutyDjbOyjz0WVnbOt08PMkL
vj7CW7hTMXQWxyn+iczKkjEnEbgkc18SGhjpiwZQ34I2wlbK7B98+CaESmkjvH32
iJovHBRXWkH4UvL6L2YwmOiJ0ILrcCSrRrQfFwZNkYROSIP2NR2R58xaw3R+oFhh
QHBGJZ0hmxz92CLoksMxGYlU9SgUnym5yXQH/oKjwuoZ2zSNg8MMg9fyUVc0p0bQ
kN/P+LJSVuIQ73RaVSPOMAOufzkCEHvXqUYnOi9dGNWsU1zrAocLvBxuZGXxxug9
mUEioa0Ot7zevJynO05ZG6QWe/GrP9Lp+Wm5i6CJ3L+oO7r22xoh9SpBnha9RHOB
mT6JkJvmgmnIDMNlJXEIRtLjsM0w8mCSO8YT4jnfXMYteduyO4VXHq2WStd+HguZ
ZcDRywMGNoMrdhi5qGLzeJOj6ZUY23le72X5gTPSsnFVxcvE+F37AfeC527XC7pF
oiGBC4QqI/RYGdTDKyqY7fq3YtW25ecJCjnt5haw91vIyrva7OhkKyksn9G20M14
ClXfZ0JGyHTmadYdLLqFQaBOxFi95GTafX/k4zpz0HVe7XZF3iasvvvSWLBFGT/E
ZS2t+KoeZ6gypIx3CYK5okR8ttJlgMRlpuYAYI43yE4b14NCbD/BtAXa7+MSXiHi
O9Xe49cibYgh7b7UlDYRlaM5noB9fqXA+BYu6VM6iii55llzyL4r5OQiGx00watH
6gv4lO+u51gU1n/Ogc9bxoEOSGXaFzRDewx8Eqw/LHepnNnsTPvwFfKwLdtjoQse
S0R9+BEYqjjhVDVxZU6ArqQvXMzWUEo8Gyh6qZo2TABvErL5GTjfcNmTQWH0cub9
9fb1Ld2+mZe+V1x5vVhtYmJt14hnw1MYiA4yBJ58g2SKf68YfygMsIWDcdRlc7qJ
L42ZUtAwS8pQWp+zEN5PSRC6TtlFtygEhsAsv6WGqjtBAjXxZ3/viWFknenJDDfB
mFtEOxL2mrSfgdFlnn9VwrPcODqIE011nDu3gqBYbzT+kQ1A5KVfq0ZvkkZUQJgZ
IWWwku3RXjwQBCm8RsuLYf8oxSyuidik6On5zgxSa9fx0bW+/7t8+uaYlcXT90ep
wxsAJozO6mCw7lO9ZxH1xg==
`protect END_PROTECTED
