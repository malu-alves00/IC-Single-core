`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eHrdSoU2f1CEcx5rIV4ulYwNZXLz5RBhM4Tb/gWZYcYihJjfhwM26UfZDfZu0hyP
qocwyWAK8nNitIRWSvSmN4uwaTtdfJHtRQyOecnX/+FTTOcbtKoLJWutV/o8w6mA
iNMm+NhDKy0EdztHLN3jfPLzzFsV9sYQHpikbS2wJxR1CY8XHwBBf5FYfFUkODzm
FazcCSkw4rcZBqArkAiiPZdomFJGI4hpDQnnP3f5a90L1YeoZkHUwvgi8bSRA1qo
jeHyChsXRM5oTKO/PRBwSGfRS7kWqF8AhAuA4meHk7yuzlipuCrdXQ9DORysDS9S
YurvuOsTFtr69HtR5C76iwPjhkopT1k1o5mBSRTKD6pSb0CzJF323vCzn6bUmXC6
K6E1g7WwjOchlMWRZLIM1X2zMbEUe7U4fq1DuQ47+00eeh6MkMiqIf1r0lbU9a1w
zAclkVIN2rfQG0jszQpVkp8H3gpdj4+Qw81ZQWy1F+zFkgvjXk+5pe/BYX1Ii1oa
fhx2LcpW0KzG9LIWM9G/7TQ4NnuU6UTDTzGm+NHJJ0uLe7p9Zo3iLDx6gPx18mB2
a18FG6WOhbytD3wZU2MijcBtURj+fmcqZ4/OdN3pBer6YTQ2e0jZQ7fRUgRLwWln
CR76wf2ya9/7zUKl+5dPvU+Zapn+Rxq4hnVMtuhMQaQHvXKtBlVlnAdEcgDCiiCP
fHconoZ1S29c34bDD1ESYWAcNL57PKVvhE+n/GS8aIBeMrcJotsetTdjkxyfiGdU
JdwBIIB4Mg7sCRe/F+s+olUUCS/CGporLtvFlNRt08qpIf3QFdXaTWguGRARLRk6
r3e82Whf9C2ZylVbqkgrXJUZrQlBOQOAdI29sKDs0gwIfKJ+c3C5SoYUBevD0DFR
fEVuvAp8f/3bgTjFUlefGpPm5ksAv5yIyHtk+ofsIu9KjKaYMoNvqAIA2oYnYdrh
blzNRhg8Z3nCiUBEbiC2TJFLBT2dg1dVZa9DrkFu3tvegUrxb2Q+DjbvSAcui6+D
r+0upUC4NgK1ahCse/7l7n+VyeufHo4Q+x3IByRigSJO0SPrGlCHoTPcIPe1ybmA
mP+SElTFabpOGhvGMY3v1K9aJFD4Zhq4Phih3KWKSTgko9UV6RwJmRY3TNjgZWbH
VLRFjPHqKSCGPUgxM4wL20eTygD3IBuQXkuMB0dS/IelmqeNEQ2qv45cY3V5CqnA
`protect END_PROTECTED
