`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cpZEOOfYX3/IuCSeKGujNrKoGgfOSH2GGBkZM2NaCMzHKfmuv4+ygll6VVka3A38
Zf2xa8eHj/IDAvkLGZbOs4FVxSJNJ3CdFnifo2himYDUS5xspsynEC6aa8c+/9Eu
QxQsRKEdSCXNpWvFyOW+8pqqkbTu7Hr8tKpEcpJ1gIIeWAL5gaTaduYE0CSr3Pfn
jCIYVYyHhzRoTZ4tGAkLQ/j5ljAwsZALuFyRmcSTzt5Nu0+0BVHvRZBNraLLmiyr
qSA3G94yWCaJzUbhUM+TfNN3tG0WpHCymKBc0lpW6IUnFRALIGlbLSMOdgzdoteX
T3MeKn3TnwSOn5nmXde2ttAoUB4k6svfQeXV+Mhlx/I9CNeOGC2nTpQwi1lBxORp
3wWEG/F1LNBdMwLBYCZBzt8LkObGnU79ORjLtz+ECaA+GrdfNRLvgkFvh66q6CaO
dbft+jr7OWGW/QyNHdRi1LkIPasVn0/bhZspS4teT3d6DThiUXKyuYbZoMatQeIl
6greu9jW8HpkRUtU5mMv1+iRYWZuuM3t3YtKo0PZkMcSuYjFO+0l8mL6y2cOn225
4Bzh3M9p4oPkgkGwnsEgYCxqIL3FtJpRHh7OOf7MqEpvjRp6/j/LdyYoPEdM1z9F
2hHXAwim3ndTMCC6rbPiJeDoVo/97XL3RRI2Ynq10cCnfWqhNYizBBY4sK1oioR4
kdUyYxGINVlbHMBC+xo8yQNOGzlDLCCKdWiu9lRNcYvW06sod43/op6Vz7+/nEs7
kq//cf8Evbz6/TjbygQo5ineP+yolklEphGUmnQkp/egAajl3i1iXzsc6qQLRJnw
RG0V00Vl7SBGElCFn8m8+tTyq8rW+a2DqH0t77guVpGdBDo9KmdxFuRuNANxi7bF
N7KSuVZpyCACEI3wZBWl3LsyzHgoG8+frgeJ462X5bEYli7Azg0x97HsLUPwG+zU
zBpGxCWfqqAgXnW6aq+0KIoUh2V3/R0MjVw8nDP8zkILxNO98bsRcGF2PWzePxeB
a1o7Eh/r81EZbWs3YHnCWgribQChv5Yge9E+p8FkqfaN2ucT21tH2jtxl9spfDN7
wZv86g2bpD21BOiMLoTvm923b10YZy8tpHUNSNge9tDp7CHeta98wxodHXS3DCo/
fw/ZXAVUBxG/ugN+kf31I90k5EP/LfAb8U1csPDlB3QPB+fjh6a0sKijaSapbBhE
/dOAZHkyQd9GXJeqfofcDyiHSsklMiP4NwCIduk22idHg6aJP0pqrrTOkIqda+iS
ielL3T6LYi1i/7VS59WW/OLv34mdYnbs6gFGU1I9zvMgKTHOI1YL/5QExgFhbW0e
BqP6xezhHCJqBCyxRg17t/V1RmG8doELIjMFCjsKVGTIK3hqRkSezcf7yz63L8ZK
plN81VSVmPXIYhRPVQupAdl8ofe05USE3xZ6vYOEOdDPMgfMB+PPiqcIHaNl3eL3
kdAdhVdDdLzcXfr+TYXuBw==
`protect END_PROTECTED
