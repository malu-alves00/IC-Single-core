`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pxGavC8vECsJmTFCc7tbDWbamy9ipKIhgTFsO0iHJQR9WNPiGRIOqkjL1AOD1YP/
JppDZqqRK2M0TWG4nrINZNrChKdesTXOrL1vwwErAiJSau0stvVdnu6RROhOxkO8
fCFhnr5hsAHO6m3OHYyNaM20tXh7K0u3RsLoXlEdwSdeEIcvNYUooODapV365aqt
xkacPtH8e+GVEonSJhN4x0+AwUn9cZsB+NxsGSj/gLBzwSbOnArbXYgiuBmn/3MF
KTKAk1QnfLqWxqjWEiEwdZguEpVYiyvOTSr5p6zd8R1Ip03DeviLm9zupi+oUV7g
E+Sa9DcOfbKAVn6bDUxArhggyXizbCJJhL4KsFt7ZYpqvmoM1Ru1+E78XYI4vUCO
76Rv0iDluISdIYFw2xF/rZPKWVjLWA23KwQQwzlI4ONFgbj3B5WpI/we89v7rgx8
WTvT4DcPcvtEQ7mp3yjP8l1+3KHt2BkiIonDVZ9Nia3fu1J+RsG/6YyRFNcVZ8My
SzLaOCXcDgOlzb+T5eE0M2ceC6zQUi6nbqyevdIS7RsP4Qh7FtaiYc37fh3FMceB
viPeYcIfbVIFY2KDBs1VXWKIC2jAF81Uo7oDbxu0NtXRPeV5AmUztlqLV7l7PGIi
uE4WGnDtIYQ8RjWm9kmi9LSIeZTfHqCKnAgkN20Owgxau7IcQpCHyOlMfG0u5aOm
asSIBZt80Q8hsLjeBp1t6u3V4suFMFqeRbb1pqzCAu+O9mWO9vyphS86Okhgh0m6
mJGDlnCr0nd4E9EUfYL1Mle/wLhsA/MUGIAjS0yfZDudjMUiCIRej21fxomfLfWT
4l1giz6jnbEuZCoZgmVvUnf2ndBhqGUpyy03rtk7/4bZNsuKPSegPFtbPOe4gyzd
k6VldlumIKV+Zx+iEpzMPbBk2TjYQBg/Wzuwi1WGmeKxXWbP95t5RTceyTWxcG8k
K/OWxq4pkLSJH+yxMkxHSQRACLM+TL8TU7Wx8B/yru7D9iXxCztW6L7aAZ/l4VSo
Izi5rZQ06MTDqccLMv5DbJJdQlRq+D7yVZT5RgRznDvVR52Zrx4U79dejFadqvxZ
bSkRlTQ8UFgFVJiD5511yqRfgM/AEmis/Sqky3Hjj4ZrgGRmYR0uTQ5GZr546b8i
qrapztURbJNty2rI8Og/3y4M3h0HNFBGIZJ974tar6Zm273of5EppwSJi5wW2i3h
rtvEh1IHzMF4KMNAbVaoQMiqKzsEEr21JjeoJH0IZJr3mMupA0+r8hTFA5li8ggS
j6+bRl8OOuSmoFsoDVx7/ZDiix2e56+97sQQl570hp+jcjWZADmUUUnilSi7vogf
IDmd10LnghuiEFg/k1SkNzxwFGvHeoWkQns91pFTO8gbJLmcuFlGpwZ/3dxzu+80
Sd5HXrtYVMREiMj55Q7KisSVgwynAYAVV7VdDC9UpL1ED4RtuBR6AEWDzKkha+wt
Iqt8cdEYJ2fkktyFtlN9PboJMfxzS//9IAjDZsq6yZhiJ8mAW9Z/E8Gvw34poCnS
Z1HVyX5yD/bvHF4QCPGMZsU5IiQiVeaSsVzQ/R2pvVde8AysBhMsm6PYt2BH2BF7
sjlIbWO/rFSAUdRIaJbAXy1QOKjH5P3zNvz6MxFakImmPr8oeRDOubI/gs5zxbh1
1yla6fWsLhVKSikzePnvNT1R77V+bdQgpmQmLiv27G0TJQQ5ckkSNXeVyYwONTLF
Zv/vxPFCHJiNQmxXLQg4Gz2AaFxC+6Hi5kVcNNXLbjQyboCWpFOFGBR/xdm+vnYF
AaRXw7Bam9W0Hws8+pNe9rIxml9Atmp3Oi001NAsyWLZIMjtl39XhHmclT/cVXuw
plflJX7ts7UcTkKqZ/rYmDdYNQVKiqZbr61Rsbaj461SU+VZ61Iq9rQWt42Vpgde
Xe7kbjcRka5mriX/MNl/vDrgPkiBzNfiq8Qsz3qMY9bx5oVwJHP4GFC4nz2HrAWp
Zer/C5SH7wFq9HnyR8qdk95/EQmGBuaAzE8xMp8hdpyy1viPG7Vqa8zmAAChy2VV
Aa6uaw3iE3vL0OqgzsIlRR2w6FqnzZj2cc7dN1zu+Bqt9lwqscnGYvkQ74cA8Hc+
Oa0jcqonDHgA5bouioMNu7TP6B+9ajsxqMhmjtlMn5rF44sXLY8WmslIpJlm9t/n
sd9cG64z6soJ7iIK0njBJWysWmWNbpGcIZf6N8leR49POIIZiS2q8SVR1L3NlGGf
QgPy2wHQMsscT7h1kSGYo6tVMSAmVpAWpZo5PfcnwozGSTyQ+RfIho5grKnitpxJ
FBmAzeJ0h59bzjDIPke05idVZesOvaUFIW7pEuLUAjPVfFHCHevBjjNZ/hqhduJ5
0XY0WorkfZScJXLQw1/g5C5CnXY+3i8d2YesRwx57CtLWjvUHOk/cXzqB+CB/5dR
JDtNiM4vXcxrvXMeUHqe6qEJXsf7gFt0vqWCsTH+rJbB2TpUsIi4lXuvKL47St8b
piBALCw/Axgv2pPcy5/Z4obR5i4IAEQCT5dtGkhUl7G6DxaNhoEKJWigHbrlMqYe
59XRS7xdiMVAlXDUMDmJvLYM08eC7lRYH/Te2ZfMWPqN0sxdM9pgeT6RcndruTMq
pQ0PP4qs5lrWqQYjOuDBGqh7K5GMXEz3UnxoX+c+0Dx3V94ah+c3DxnxWHnx50Eq
rwOrFK1YvcH2LR89dbrqc+HaLze7AoE2e+MaHD7SWnyioC3v5+EeGwujaH4guEWo
gNSX+aGQsxSmnL0ts8n/abjm37ms/8vDgI0iC9oh86LzuyUBFBNR0Vv21bNX1hcI
nt73y6wLjzWKNExMbwOxYfbBQVRa7JBxkaa1k5u2speWvzN34RBHCWLAwpLFmLDH
/Grz2IsvRogTd1G7YKzHtLJVeam77QadGZ3L85v5Fh+7MExxVhilgS79NOuAV7Oa
HgKr5rgYaqvmQ4dlcbjpsU/2+kVI8Z6VXIsUzn6Yusu6CKkOlHXzVL4DJ6Nj4/IQ
L/h2TXqc5+3uz3g20oFuz7gP0g0wICaIBPvli5WQfG5XzdO25ttvFha5J3/nyadC
OeudlND0//ewQ34WRcs95gJjX/QAvOOzejzE/rmi3MKaQRydweURa1gCl9DrTbtD
C9HTeOmRWk+vMQQ2ITT70P0aWt0n0EC0jwRiTVrqGOqGjHVWzzd0pJEMhHYFgoz9
JaJQd7dLchOjLfpKb5ki4+HQwLjn5yNJDSQlOVqiZJfOtnzd6bNa/SsRFASg+4tw
7LcOyfHxH0DGgsLdHhLY1f5ER4dEGobY87aLT+GL1iiSya8L4AB23+VopyMeCeWj
2NKT/sg/4l8rBPfNWtf2p3L/oVFGW8CE1bpUVsR4o2Zlfes5TR0SH9w9YjfDq/j6
j6typhEvt42RpdEjutw3KdQ0YYGe28JlZ4qb5TBnNWWCU2fAFQOihCllfOYi++aj
5WSgrOZbi5tQkeTfgFg4VH5plg0XtCVLSWvqAbguridJKbW7zCMaBiq8lFHBb5Id
0uklL6jya1QSr1U1Kqqg91EEsPluDP4F9ghb9IA6V/gVnZOiuqx/Q7TR134aKnYH
DWnbHi4wXmp3HQkE8bR15zY9a/OdqCLDvFvMi7FyLTrmhd+uWhLuSLy5BdH1b1XB
8zjFhZjABkeaCw37fk+/Q+w8RAjy0vczRrXRQh3Ir0RkT9D/c0z0HvcQ5YnmD9kK
rO2DbSusEPVzzMTWR8yDYW6yydGsxH2OU/YNfQ1tBk1UjcNzYt/iQ8zeNeu/tso7
JvGSk0r0DFrg1bjymt92pKOdJOv5suLTNJNiqhDgzLl31LT9oWxdcHiMIb2za6+S
5LnQZ223xYs3WFFzu+4/9epAm1ttW7N9CvTNB6XVhWVnF+j48Cx+b1yxgg4ajaMa
qBq+9Hcbc3Dt9CtPbimO/nHbr1/O/W28p1auUu+wJW+IeiF4lTv7uoF0VR7CYPV+
nd1XN0SdtQ+seux6a/ZlVvw00Xt0CtDgSYnizvY8YNsOfH21Av3XhRYWQZJ+ysew
D1vzzfWf7AVFqLrVqNmCo0kiy9avDNZbCMD9cVViqHqLHtn+Qxlgh8rWlDa9yL8A
lGc234pOqfUugs6tdwXUePye5YRElzqWncj++8Q7ODCoCztjsdWDrx1RhCc4AsP8
`protect END_PROTECTED
