`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
n/1xNePry+rjjGpCg9V/ZvlYofOSr8B1jZeZo5DYFplWYfs9Q8nouP9k1yfMAprB
4fFnuzDGuyLyW8B9rusvjm6Ys5TLxx9EZQeyxbyzZTkhgsHTjQe2S8oFE89+7WST
0hq3Wztn0Hfdlgn9dLvx2CAUScNxgC44EFunRatMyzx+l8YsHeMb5eS+cjDDON6v
z/if/q3v0rFwvx0WIJycaOcq/6lUNZjKcFXx+F/fPJAzVJmiamcFaq7jzCbDRjG/
Fcoc3OuBCg1ZsHzssNEk3Q2bkvS5dGN85MaDcn8kYri5+wIdlGU4GBRAA18OBerM
44jJ+kjRYIYUpfgi9qGCAOo5DrtpHFnw0yABRThsom1HnUXqDPsrYPU7CpK7ZnaC
AAPS7t9bpGCkGoGoM+NDm/lwQ2nEDNSiYMVUs7KMFTrb2AffKrrVzBaKB3qGQj03
EKlGBdnab+CffGA3vrn2ZZuNnPv0eMjsyUB519Ss6Xl10S3KMv73F5u+ZmL/sCpj
iJJ1LMuUuWqlMAIdVnJijWhOED9gGR4VMNC5bWb8b+2vxu5P1Xip94zRANCls9PH
fvS4FFYR/8WOkeBORTrGk3e4yHXeDObo+i5e182o+XbjH2/K7Ped97RUmJTfaWuq
fHigOytP4an61ZZY0884Q4b93K8bUjK7B/9OJiJbsA2/E6bTujroNI29lEIxtlxe
WyY2x/OipI1eWxZSb5gfgVlTowf23aGP+W3QcwZh1dc0VYSW9lGGQlmeJs4aJZBl
Cq004U7Bj4kx9dQ69xg1J9gIQP8cJDFXqDc5VjNB5V8mODq+i1kEZvoxHPGE8o7/
sEnN2tqWYz5CA+k9FRbMYP2vA+rcmBOdy5g6ragniVUDpS6kF147DhgXg6Katw7k
+rxcsqEPrXr+UZwGc+U/bzMYvThALpcYz0sv0nidQFlhGtIN+mf3w3iBjP41vnO5
tAjCqo6EVE3x2YPhgBLMDIStbazSrsNgLrUFsLMqIb3kJwDOdoVxAyGqyBtVJp1A
L7Sefx3LbGcS/AJNcYEWkryRDcxIQvRcfD0c4RKJJmKUkcDzLcyDtUKak2YM5Yys
zCq9md+RSE5WhYR8KoVZTU0dEL1/JU8WzqNNjPD9CcJ/iCVJhidymphWxFsbYHOC
FnuYFJARjxoU9upRegoL+cHkuKka4FqOw0r9xvNj6xCI68rxgiiOlI00Tvn1ja3V
/UkItlB75WLEHVFFokH6yS1CBvlHs7blSw0V9vYMCPk=
`protect END_PROTECTED
