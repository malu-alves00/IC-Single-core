`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EACrMuh9aql/zgvZ46dxBaWt1FIlAMbXp8FuS8XX0RJHtvIPOFPoZG9VQEPC1MCV
0X7WXH54eU/UPc+vTf/8+8L42qWRJx9FeiUY3MXTRbrSD0u6Tb/mUEn7o2HJc4vL
1BnN1DJhVBxjyqs1F11R5wSsNkF+V4ER80W59431100pkaRlCRVciqqrnw+zs5Ea
CnxeR6uF4Ij/0rE/pUf4qoKNhUPdE0lQx+4887Ok9beDKWvuargyTbkwaie6fgkp
BEFp/QUvNuRFSFN6NQhRlQ1bGZmni6HaeACzDlnZqLUN4z4vAt21DVIPpgC1dmaw
FecDXpI+so6xZiSfvZkQ9OzBJJ2E0EI9eGtJbXQy9KRiNByJaafpbNnnZvWiFAkt
/N4PJooHAjSz6yi+9YHGCHbl8JmQxT6h9dnFKVwTshVxV/IfSmi/RtdsSt+UZxZ1
F1Tbo2fFurlKQaPxu8njQvYnfrufvqebYn5TSLad3ahivLHQDC8FSXkJmGCkaJYz
pXQauq220NAyixCGDufDZqR5LznWi6J1/rQ9361bVVdhcFrOFpI9vEr5IHErjqtS
wdnceGipzWXeUHjpVz5DeulKr+jk/FHpdvDlmc1gRSG983HxXQQs2SiPP3jGN41s
HDZVDEhZxodGGVMWRsR2xly0O5nJhwPVTzDmCRg3kXaRMQ37JLttxu1KDjF+besl
RCX1yhTSUfG9A+viQYcPT+L6Ulke1+5gGEDSnt++vzTgvMaLI8cSBVgbR1wYwd1Z
Xbh9g3wIq1buuv+LsdohM/nGzS+1ntZj9Wy/v00JKEgfrPIxnxWcIZHab27bTvfO
WNJP5BPPcwYjrpY9hyhr7ZxCE/Wj2bHmhWD296rwLBm8ZLrQrJhwpK7RjQvnC6GO
fC0Hv+ET0hIRIjRWKkGRzMFzYI5qHk52VwNdEGVo+FQ5+AbIgwDE/FRJs5VdXdPj
Npx+3DIAHNZ2PKaTq2i7L9LyKD0E0+3fPCqwiNVCyYYi5TtD4LhZQ5GijjWaUzbc
8Llmb9rlnfyMXEFYNmh/MlCz55bB50LSvbJqaD+aIiRefyPTVegSxW5KHZxsY1Wa
`protect END_PROTECTED
