`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+1iXT/nGXHclVw1eA96BJ4ALEnYfKnDDxrgStuWhAVzZjM4Owyb8v8HvxwUTRIwM
QmnHEV/nO2MZ1z2k15O66C2R4G5AVmyYe4l66+Fti6xwjSVPDwGJUYdTze1SSn6R
NBRwkKwCr9A7F6sORghMDhPjpA1nq/YK9q259N8MHYe+1IWyyK8ZJLOxylatMErg
6wxKPq8w3Z2mQ4aLe+OjM1Twqn9DZYCr7Uwo91Hsx7596s8dU07+l/UP8c0VnYwp
i+/CpvyQdmHHZuXxVK35bEVarKrxkeXoToq+9wCFhpITD0FpxWvrHids19hswfQk
zonm64ioi/oAJzaOMvvZM4UwbNsKl+nDRFjIyL3hs+FtVcxDUl8kSIfoOcARno/y
qp01RQi2JX5/kjexDfZl8wiiYC4YsIKSpCP7ATbtAixPupuQ7vs5l07qWGZ8hRJY
WfIEmHb3Wmsx4pgGzFjnx9TzZQt++VMzieLne67wne6oJCEpfmjTx/s/NqIu6KoB
U4dHSrP/Ipu/pausIyLUzVUdLcag7r4jpUd8IdrGWMoFVbs/gUNdBj9DzyUwD993
/YsUQjsGZ7/xttgXjWC29vx38vM379qSx8g7UcSX4G0M8lk83wGNaoSN7n5Nx7QX
dCNbA5wqfdYyndoGO4MmWCc27E5zDytDhmpoTK/QMfEPzFj+8xq6BueDJ+hpPUPn
B7Xz1gHw5bsIKaCADBRuH0XPJQdNE402w6QP17E5bXCwueXHQ9TFNgH3YyjYshJ5
8TxXfVVu4Fs6qJSKqKnAiNBFsUw/E7yOwv4CHTpiecITazr9aY1d/DowjiekQ4X+
w7EOqesP4/yXKuCvTpbsmIclald5yoS08D2zMAnvZIkIWxTNTBy/5gEXPKE6Tqd4
Uu0/ENO6O4t//Xg1GC+H+J1XqWS5Vu++JFqqtMIMVMTSqtC/L7KO9GClzFtlOxkd
wzDOSU+V4jZDf4FqQqWeY+dZ+b8LJB6sQxyqiTtStkxdQqJyV2jOTva3D82ajMFc
oRqZjP7MU02A6K71aMN+qpJqxOylIO7iHeF3Qjh+UHfC7NMJCa/gfXAPK83CrwdE
zIyWO9PzkEa00YcN8bwQJz60BREGfAa/vxqwhVMrzJFFm5Kd+YeuSky3H/KLOkug
60cy47KcYmzxxJ4qA2Oay7v4PfaKygrOG8kY0dAjO4VKuztM/dO1vabLcJ3jk8SF
IIqOPZNtpRb3nJ6sodDrXUIKjogGkirhKab4P4XG0gHbvcB6l2Pk2tEwCZQvAHuO
bOaMRHIdHPi8yAafSCT78mPN7mH8+GDkXUAglE/HuRjL9XZ/M/j90/tNFBcj9UmU
HkrQUtTdF04WMm0S5j2OHt9K/JRwGmAG3iLwUqV3Drg+gOI+y849mRKfWXd1zMVd
oQtb0MMpMvr1Km+tKJLyUiGxJj9HIZYkfbDheIEY72h5+/DrY6dEunghTWXYWwoC
ASDZMFEXNKKl+hIomlvTltzXtrTY1sXsd7VPMo2MmlsZN5j0o8pkDwYWBqd8QG2E
e08GVh0p+rc8bSvK1u+IQ3SwQ88vGwYfoDWVwwS961YDkSv6M1wBsZM/KeYik1VH
ZSrmdl/7/2dli6bY+PNVRk9xYT0Vg01NzCMLlO2+0/wG2JYQGapN1Ityg8kh9+1i
b4DU11CV1fp9rH6YvTh7ak215FVMW93mdoXPLD5KUGFbAEwhvrETlEbMiOzvqmG4
iabp3pji7zVgutskpI+fjLTJUrJ35NPXFLaBY/fBI5FoiiuAX0BzMCfRzcpYd+FA
UFh0Qo5d39NBsaGhpuWq40zD6LGcXkvWNZfl00UBS3XsLESlmjSSAEgVk0jOTl/S
2qARm7FPyMeHwPYs0sDbhQ+Md46ddJyFyU8jCBCvKTwk/goRTs79yNiH5+gsCI3i
FFtN9zw76f3APlPwFYGevKuOLSoovM/GSRGVWMIl/b3pWhRPKzu9FvTXHbEuAYg9
x5C6l4QbVz2FD7oyg+svZZ/Tei7wpQNpvjoI+3KYXG4BhEkYk4uVf4mnvDTJ4IMs
MhRmLgoTLGPtXGY/3Grs5apEVTzfciRMCQ15/v1MN6pYrUM8U84P7QNZfiumsKCv
O1A4uTDKuJHWOknBxnsU14QDNo5jz3YxbyGKtwyy0cCA2Kzc4O+0gGuKN5/SifcF
6DNpkFtesKlOFO0GsU+3kdLpzbO1yRXD86fAD9v5tq85FqjXMZ4+mAhUYWNOpab3
QvHoXfhpd5xK07fwAPjNx8Os7syiWK/UbQJRYIQIWTSvUphsSL6e3QlA+6oju32S
3m5ILV3ArxLA7K/Wfcil/r9vcS4ELEfT0KSh0tcQaXKlJj3A6hfhKKYZsk+8/nbT
xov2JNsoFBd1wwjtSUvaeUXdnwdJWFpqEBgEYbm+byiQ1YFE43uQcM3C7qygrtdH
7RGaxbWI9iA0WVUz5b90WqfoKyAP/gASvanTmV6ZNVbHlVsaSHA2n6mHMSyFSW4a
3XkChw1Opaw2SaZfVIuDxdYNcENJVGh8awBj3Yx50jUloC+oepeGQ7U1FOvKM9Gr
4uKBDmlFgKe1szBlbFHFm8SBpFaxApAFYn8g3esZoaR9XdNcpjzA4QZgCa5GLJMx
45yeedWB8wJNQoQMOX91+D9uV/dxNGebTAYu6IDYPdFh+mgVfM5BqHBkn8Bdm9rq
4sICrkA821AA1LWCOAjJ4stk+pzsjAhaeqrFD4Lv9wrLO8IpM5n+dGGVP6hjy22F
ARe92k3spcUbDPMPaL0tnml6B3y13CYEX/eNZsci5QsA+7uj9OcicIMoJSAq1qVJ
Xv8DUJaNhLrIaBz00XdvxZFf91bJt90De6ODu2V4a8IMv/y6KsvXp4Z0/MNHrYT7
sbFDZJzJI58ktauTtZmWEEnYD0j7a9pzrs6ytG3lxreXKqBqs3tSDFCfhDmnjwYY
AcDIngIlPfaElbK0my0WKsgWm78TGFPV+KrvjFrIQndv0AbgMaFpAVRiNjfudMrC
aMNsWCo9ycKEmER4GXMggS6knYROFRXx/PqFdtMB3NTfWsLOW1j5qBCD9m3sFe29
E3B7qS59kHPQHBxnF4f56+h9qHeMtmcILx1UFCXyz70EX/jH9jAuGhLdIDCjOY6e
uuKFNhV8SKgrW88AWq5V3X3B4M0dtIh59X4nqD6Yn60t5ndSud7ktpTiv/nRullu
g4XF03xMjsg9vtyn711WnDlpz99rU12sB/YYlGvRfriTYBenE9MI1k6R9ZwxRiyx
iTm1KIsooWZVl3U+G2kBUblYhQFmaV8EhdO46jUm52cj4PMCUJBeMeGybA9NQUdI
0EIYcSPWltt1OD9oOcdRMe3JWIQabJCBi4o5v0VO62QWSu0WJBUrSn8U+MHRoYEu
/D/W2sHKjhj6ivT0Um+zMCjaDVrMfinfQoVQ4paeVqdarqwnWnO/RRNYnPNIUjVU
iSLt+kbdJ4kX1myLMMbh9+MD8hW2/tFk+kJn8HRW8fJzuqU1gjS73+72VDAkc6Tk
icFtEDpbxHqdr953kdt4oE0LRNCg0t5Xh4V3P23TYIbg3M5jqbarzHxLOG8E4vyX
erHym00IUZOV/I8bwwGV0DU2AyDuQMHBIyzPKt86tB6YLX6m9DQDHp686h7etLdX
q4QWE2KVg0WU1XNzw8m/kc7RaeBbWiISlWvlHbPjoHDSF5ujNAFpsRnzm7VBEklh
0R1FR8llSqFBhjglepOW4NliZUABCp4cyo/p+4b7IDH5PAot+kiq1kCQ+KKuK957
2NLLtb7MftQwnrlbjjnMKEZEtxkgdwVu5jG7VxfgzEN4DSudro5cWL5K1ZV+CK3E
b3EHBLDoouquaZ9MLW8gKj8F9L39i89iy/ivY76HMrGynrmZfpmUCBcTauiUX/0r
WgtxA+gDLKd1J3H+U3O73ZUfsrjlURPgRsQzMV7TCIxprfCIKaXTbxBLFVE85w0o
9omgKubPxA2+tx5cp9cP3OWc9GdcBxFHs3hZlhkKBrP9+TNYiW81QiqOgEaz3eM3
0jnTZjQhNJ1AaiNJ+Pe1Iu8MW7jBfEEVGNTZmECLnw4IDBeaCnvOjGmGUf45NDCC
N9yYsH824yfHXHJNFnSz6U1H59oKCG1ApFHWhSqD6+iEQ9z2KsvmQmSgEmCkdm4O
mruCLoeR5HmutJL2uAot+ccbtr3UQ/Gu28zjYvpPUD5Ag3FQ8E/4EvRNj9QlIFhY
HoSMu5xqTN7MdGGHLo8pzM1eByCP8/UsJ7QJPrWkxB3WXjT1xhO6go6bgKV8OJL2
EfuacHqrhjqPR25At9geI2FFSQh0JHEd4qDvjuH0V9baLZlVEhN4GgeB+nwgiVHP
n2Rxmq8e9S3Yr/CEL9hM0FLfCL6Reo4+KznWQteCh3wQfd4gJuB9zdAP15W4gqKu
vp5N8VwKAyWZ9c/nIA7MvxwJ5J7OZzzxB8Y213pvReYX9+nw/ul37T9+mPQ28bO2
gB9yhQNWZ9Y63bKzugQv6dF9x2sKRYquydcIzcCYJ+xtdGxbjEXy324xG6NUdl8R
ozlN2J9WRYgKbFiNqx9FAb0HJCyscFWkEUgahXQbTrLm+EvioDLeCKjMYiKNtTlI
4LgSyJmF0BdsPL3UuodGHK47HRzmCUs3jNEOBpqfG4Ia/hfbU7RB9j/9npxA/4BG
sPIQFcZYQfzGp0KZo2ysk5hYsPPkVTSMVZE94Db6UNIeT71Bb7MEd3ZKcsvCGouR
n8sbXKdqTbdGyEmk+Lxv6kyYPlA7Oy0gL+txKU8XyW5kdMnDah1x1u0qQAtw0X7t
qvlSg+ejr/Vj5nXM+8IwGI8QepXq+Nxn6V9hX7o1j9HjmL3aHpxCanQ4cMvsKpNC
124IvXL82yHA+6sxSZXPOb6uMiGQ59hw+FUpSR24mA7PDXM1IAIX00P44FOlwknP
tMCd7jCr4odTsWGGmzA/vPOD5LKb/mhhYOxjbXxUMbD9FqiGSP1+dbeypu0Ks9Qh
lWtJif9jWlLys8+5PMnP0TVwEf1XMU/fxJAEc/yGF2shG6lDdhq9uQUC5wIDM2pC
G28NvgU18UcePholFVECJAH0MkGZNh+AkN9pAt/Txqsz4UlOAKWOyRnEIOZTeZgB
On2whRxV3IG2X1ehiUg7bXNOWd9OCAL23xzoXiAY30HOTpREqsCDa60rtZCdYHqv
TVZrU9JDh73dTTKZO1WykrqDcJ6A6zxjrjmP6Zoa3wlNGD52mkyzEBT7XkgzgDZB
JVeRCH5MWeIoV3hMI3JJnx2CcEAPsamTYYwBi5NE/8Suu7Z8N0VcQPrmvc9uaLTr
pvKh/w+A14WYAmvgAnwDUKLnF0JGy+ssCGkSD/jLjGXjYsPuiU8fESqZetaCYnVV
EvPr3fAv1YrQlFm5eZsrqKmrv0Y1gk8qwUIbsPna/sKqf52/UloLBlo/6xFSBVY2
KkiK88eLvN09LBczUfpqqYiWieIPEkJP4pAL/dhbXyS8NkUyFeJfbh22n/UkR8MJ
vVveNkMWrGYoG9IrvS/ZQ+DsNzlEkO3zlZZkoxsov+QDAd8dgNHRiU6rFtDy+ka0
3lr48Knp3qL//jJni1yG7ACxPUI6PPrbl0NO2atYO5cgpVBXxuVOaAKIRc7ABxlu
BR2XbDA2C1vWC35JmZQtLEcZO7derthVdQsIllxg7dHUcrPS96bCpA5o3xUOIVhv
kfXJ6jaLSsKzmEIp+5PR5P9mM7GnJJ671P+cZGivmvo04DXob4z6jbRjBSJ18+3v
iuF0zchLSP7ZuWr6lIV9E2aJ7vQn23rKQRaT5OvZYvFUZi69trPWiCRDf0jnkSAg
E+bXfkGsecREYxhtH0dR/1nVSwcyWwcMQONMYy49FsNJO/xwnrH03AfsNT1Pa3zS
yop1ImcGI534GbmYMofgV+TV9bPLIbVI1sJKlqrHQzloy83qHwp41c5j1XnM0G2S
795lR5E8wgJkVXsvVVwLlTv9MWP8NFTj+fVTNU3YzfCsqe7ixw0uJINz4bgWSfqi
Evii4HwAaOXGyTWsQL/hDEN4NZ9Tsh1qNsEVgIPOZO4SuwRI5lLHWbqk+4qNore9
3YBuMTK2Fo0FssyLZbPlHjf0JXdpJ02L8Ym19h+5YbrMrkceT+sExPNtnImSt9mE
EE43DdWpNbXZZ6AR8RiutuqtEKqu3EyAqaXbU8UkKKAIEJPhdpSFSe01mqVfvPBk
J7W+2NS/1uN8VIak7ljX7nx78pryAi4zgNkXsWHraPAjmhMb7EznDfNh6jV7zMq5
tuov3DjffqXtPitj6ODJQRGh89q1vz5K9izaBHecdPKdygcPDkvZHXcCiSzBrhId
22kjcm0GGQWg5pZE0o/UklOXh6WzJxJxVB/W+Xlb4yrmketVPgo09Bur8kH65Wy/
bec+hEjNqkEFFVIbPcZLqe+saOBlwxcGHrLCkBninE01CmyOptzhJgleCHOMm5qq
0DcW+sA4nOE444UFkbMSumZJ4otwcyGLBiDJhkemJQ+kSd8zt1sE6Ey9YPLWCh7Y
TfwpXpY7OdIQ0Ou/JxT0NH4+s4wfhS2iThu4HtQIS6b8PDLNQl5HPDH597VadOL9
pXy+xfww3dHXP5fd2pTqncv75mqwRMLgfO3ZKl2s89pjwE3+0rT+o1Iqs4e1A44r
1fXGEoic7VOrWYGAstx0A5JyWguGRuY0OJ5z+nZm8E9Grr7NZtz01N7lvA/iEEkN
WAaigIXABqT3obZ7bAH1dk5X+JIXY2TgjueJERKdaGXV+hF/lK3VxeRG62J1EbWN
+irhI7/mDN+XeOCSPuOc/n31m+jn4egnQaJPyh1l/FUafjQzYXekVf5flqe1LkyC
JskXGj4jvTk5uu1twNYo3nCfLX14LgbkOuGVxVUuFIM8J3/ABBydS8i4fiwG5/c2
bGJ2Ue7NPEvdaOipXJjG/0f1baSQ2d4rkznuUZ24u9LJtQX6we4FDGQcsdyxqfG6
QAE6oflDGM4bw4C7scI6tr/lmpgMp36PcXB9rLdP6bHy5jSUqK5n33o/4K6SOGrO
M+m4sxRcLquiJSfekvL/2IDtioGt9B18gBtYHTI4mO87g5/5HLJi+VGesneF10W2
Kc+6LMP8ZGDXc1mNNTPyNCSbiEwBc7c35LUJH7rsI7T0dIVWvtgBzlIQT8C5om/o
8CGxEdeMBNs5L+9Ptb+h++3Fx9HymYtIdBl3MF+t9xsq5vcCs/BQDT4LwAk0OQ3j
dDWVOhGx1JS6SYBaTfP1ix1SprvdBnA2aBfpFHm1uMg=
`protect END_PROTECTED
