`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cejsNsspVWqnAu0GnY0S2zyVnoAFFLU8MO/+LsLDiLw10yiIwyFQTev0v7x5iSBZ
qEHdrCPlMe7tW53RB1REMTo0bCY2pjzcUL2ojWlzC4fry1tnkMnQkwi67iKTOa8t
skH3cAFTS3B0Vnd2khtY7y/1iepi55lY3An2qNNUEgQTvyj+klgHaPNAPeFTjSXj
dJDbDrW0Jzt2UaEdkNxc6xvTpcCjvXyNxfTXrqGo88v0TRj7YkPcH0xoeurg9XAZ
b+i/+sdYaig+pTaW0pSyDWBz4mPd740OFQ7A4ywVVPjcp9VIJ9jqmTkrVQRORv8l
kHtd2j0s9nGwse+P8yEmY/rkhx8pxRgn4ThznFbA28a52rrX0XE/v7k20p/AVvBm
cVNfXMHYP0psvifX/YbaEeYfdB/JTiJZ7ZjfZ6geyqgsNcrhSWNqgRnz9y1tc1fW
ga9hwz5PaNU8koDZc7YZBCVFr+x7mt4p2p/ypUQtzV3c0TDVrbPNEEp0qrUe5gT6
YOoJy5hn4d/qgamqMM9LA8HJwwelJ3+1/eA5fZ3YxWHn2JzNh9vECQMmumDA/95n
1gGsdhUCXrGnalik8JBRTRQa2yoO+XzWkUFPT+qJlmMrgBkLLMOFWxiI02y25C/Y
XXhOKgFEORe6ye6SSyAor+iiq0x22oYPkjpkbq2Gd1Ilg3VZiJz7YoS6udJTJn/Q
1c9RG9g4Y4iRvugTT9RAUSFPvnLnaIi7vPTXypxZGshxIrg+K5k6YjTU5Vy7DCHh
CjI78+AgKacMSsXpKwZS6FLlIVPU6dC0EYFggkhrkw1IgYCOSNki7Y4ZSIf5Fbau
HVBRF5h4Vh5Fur8j5IBQWCC29HExao9BBvYMsasN5M6gcAy/l1SxLYpPJNQOcKpn
DpBxuXEJtFaliDKvh0YjAmbVC/qhNdtOQTW6p3vv3QZBzNB9EoWiHipfqcoDrcvy
6Y+OwnXEL7IDfN5xVkW138qOvSw6ureG21UW/ImIEgNmFbvWGsBIbJ6+QrK1Ue/D
1wfRVTOhk7sFoPizK3ju8Jsr5iaik4WLs8Y7oquuwXc60QdCo6kaJKU5EK1bk4GQ
Alz56OfIXHhlK8W6U8+DrkGbPtKSNAumxkOL5IxncPjoKCMLmLKuYq+DmDg7z3EA
KbD47twLhDA4tG/cHCGhwl+qBg5eTH68r/MbdVxuUR9FBXQeGl5Ge3I+eIs5M3vW
FHtU6CmRNzDZXzVQFaCU1Ha9KRl71HApldWJXNj+HqZIYPoUo8qfbD5PEiaFq72G
6lhcRgkrsJB+b3S6SOlW3ujBESNI1n047A5VejyLXEi7tnPnGE+ONoK1wj+gATwD
E1b5mpJuuvjhGncXaoIp3pHdh4QSSc1MA+HpmgdDZu5kXvpw+yQbn9cyMVG+5axn
0RPCdZJcpTXkUhRIggTEmTzefE91XNjeevecXg/JiIv0GDI/7+LDw3KjPgyJAMc1
qnhW434a0ZeycPg7Ul2dfDUYEz99JtaithmdTPpLp09PYi0oy/xCZgf631OhjtGj
t3dyTSiiWDj9UHbTZoml4gUf0j0jSwX29xXWQG3Z9cY7tP9/XhmmfHDkYx4I4oby
rCxGa6bnGYETx5JQova5Y7r3XB8SOn2OXkGRlvh6F7i41D7kS9I4XZGNazfX8pbT
eeBvNVdR1gMJGDBIMV90s1zfTqLbDR95VHFzwGqZM2uh86d16HtFAe5sReVkxjF/
RfvjeIHOki32jGT9mvk9WzTe7TfIDtqiJ8K18XomnDPfOIaAsL+5FZitD5Xsoers
Nu91gup7LmNUacthRB4L/Gfqv9bKNlmz9beEcLQ9LgnIAYUjSqx+TZvr5KUTSFe/
F5RBz59O/ombJjJYG2gLw1qnnuRaHfNi0dglWmjI6CWz6sq/5N0KuQc/RTPaFe97
s+BPHGr3Nm/e+71tqkM6S4MhNwLw6GcuvA4AdmKlL3qw/C4fUj1sjoaYtIDK8VVH
6K7eQK+djGl1sy606RuAymZp4UZCJlKgygWPUPe1RtYo1iL+j+4pTyjPl7O2T7tB
m1BIBtmbNBFQ05q+CyrJMqBVqtM9MRjGjE/1HN3ppE+ghyk/X8jFCklPwOStjd01
YffF30hgjznlpDlyPYqoMGQKvfU7GYqQM+APBwfgqmynRedr4RVRWP4YrUKPauh6
UyExh+oQOn5uA4319sukUD8s6k0zbEf7XhWMrCt0FjtxJa21l3wSYjeW7sE1Tk0Z
jMbq1ykgo0G/ZNujymgWxk0BZg/VJhFrzTpEMJAZM3wuLllY+1md2M+P97l2ZUyv
HCJigMOUB/7FoposNVOgzgN/yWdrzndxea4wPZSi3MSMjR1XWzCBFBDqLcRK68+p
GzZHxwLjf+U6zizn/gL8bjQ/DXyXr6xANjY/kFNb4TOz78EhyzEcxB65+Fiti05/
7k7tmRp5qxuS9Nii4erFvjhx/VeQ4bG4hFryINRX9+E06QvoyXLvqQqr8TAw4ayY
4PJ/2vfyQZTlbfH8bVoyKj92ESr9BY5BWbyj0KgtCncaWaxcKG1uOsgx+k8EcIVU
unGj12B6fH+ixh9RW9Wf5GG7QZWTFhlaBehttEI9nYsk43QYooItsnkqBOhQRR1V
qYbR+SaPnS5VVwV35HUz6hoW9z3XAyRcV83/4lLjI4wwdG/iaHU06nZOleeH/btM
MmNpIwLbJjaYnj5f3vpila3rq4gWBAOl9CeQ3NOTSr6oMr57icysb3g2tBJdndXK
HOfirEUP9u2i2ht7dNTQWpgnBsuVTGlZymYNbYqLoeAJbH8zyrEDb4iOesy424tB
f6/l5XDfKHNJ4FVG9zMRBaCnIwMDb0KxgYn7imKfGD6MZrrS/3qU1/p5UFRV628S
0m1uUTliycy713TY7aP4Eg0VUVpIkvmu7k2xYmDNQ9CzYJHqaaWWjpZ+QlBSk0f1
ZYWNpS16OGX7DTVANo54J5XBUseRxgHUQ23/6PnZk4QYYEhmPNJ2n8WI8oH/LOtE
FbwTX8/nd6WL3Qr02RLXFj/dRw+St8vztNbQegV9yFHDFgAv7fxJLaiNv5WabTzD
F4bOR79JLbwKAuYA5Arc4xvm8aWYDtNwobDScifP797FdLSHFjwF4A3L8TZFwlFs
troRzF2wBHwEMMvnwuopmKhJL0WBDaS8ft6o+LMalXLnhptSF/91aVPuvC+qx11Y
VVgebp+h1MeM8dYqd3bNZHFix1bqomoIb63db8VdOhdV/2zN2RrhYN74ZmdodZri
eyYtFIKXYk/CRmfuXd5uZSCDi2QKl/IJQIVOzeY6dr00YJFS1GwwiFL2UhiVNwtq
/s2sJF5YrXnR7ZwSLZdhSwZPQh/veSVf2Jlm4XkQ3emH1m0YejtEaEVbFw3xjuDo
8yFicg6VJFP5MclJg34MJUFLs17Or/RjpatTEIr1Gd+qf6mYZ6lVD+d0dOTZwGWj
OdJ75t6cs9KkWbqKytKQjbEkWREty66xljrUORcj7V6BD/X2cQxbHInwhxmS3nnT
2Gl/D7X4/Hp4ZRp96OtX8bIm6SgG0dcvF+E4eS+7V2o4OZJ23jB289yh9ayHLIiE
adgicjT1K92aQMwh6Ln23N2k1En3KLBWbbWQ6v67R36Eif3rNXAp+9pyH57hOdV0
jzk9TgGxMwU6uI5x/GD7pZNfqqWGXh4WAnLVSNXlhVcFebgbfszMe+vSzncmanM2
/g46itfkQm59f/ntgu3FPa2VxJtbVHjMr2TFYcBBtVidXzo21meN0JtILOgKUxp+
+3bW95KBxA9OfOwU9x0tuvwZgyT2xcR+D+jTHm6BcK0Oszu9fGNgRnBSw5WblfB2
iToyrBWe82lwFWJJELhFyJTsQxpWoYHUewEChuztN1in311bdOLCHMKxFPuguLGC
flxJJLMNtndVP+yatK1lyw652NWZbxmAVaFpBYU9JkMZ8yS+V4Ogp16vRK8cxhnj
drEMZWRK2clbjZPv+PKASrFMHD9bkIuvITxB7vj0SeWsTkTbV5nU1zN0MqrtjAPJ
G6+M+7tAKh/gKNpjBdsf0hh4kt0J+AqLfbNVsJLIfNmJgNRgaItat9LT5kYUwo/Q
JNQgZcKVpBJwaQ8/neIGnjtZG4Fdk/bl7tCujqDixWAi6WBeNssGPqhMfLY+D818
fcg6dSlUqJCvS1jjMEpMWFyUeiGCSJpAI/boTV5z+mAgsJMc/r153mVSZ86oiMFU
OjY/U/+mNk3ADRbkWBdgJ2ad1GgQd82pZWBhxEjtR4m6tdCL+G/R94QEsMB5WVsu
xQqNj0PAz+5rWNQMNbQslO4DSBfZWJm5/zgm9r6Y65OhJJXpb+gL06/GrV5z+51N
NV/1xCMRCIJB8/DWSRbeHK5bazgISUI+Gk/MqOgfieLM7YjU1aVMjRTYjvvcqCZT
HalizyaDFSWlcr3fHGuwKQKWPIfI6m3FUjrTFdFtHvVgjkSFWayiMCTxKwB9w1YL
o68CkLMIWuMVnRznd5EF9xKMRSBCumAoL6+uuy/rQmA+/Dsc54QBV19tWH/6qwq0
UuUySQME8Q1TsNOQwgtmXOg+b7/FvCF/RMNxMwRZbSqxjoLUH//b8DjchMi8OV8s
R43NUdu5D0Jrhbu0z67ckA==
`protect END_PROTECTED
