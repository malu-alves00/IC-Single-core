`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WsSQ48z7OUosSFcbzdXb8fGzM34IkvIaU0t5Ax/6VoG/9CpnkIAc0mmYGbSnnuHf
A8TEBH7UMtRDThhHs3L1uMqPyXKDNKkBPZdHZNVV7ouZ3A8Rh5miEC8nM8pZbyHq
Uiro8mNxsOXZeFEKEmHVgA/eLRmh8fzLaSANrQm67+QwjuBX0rlfDCPTja+pLFtj
XWVLeem5DCvAN6EhE4ksNYjc2vRnWb9/S/DQXS3ODrltl0+8XcDu5AlPTrUlLInj
RgwH5WSICoqOSAdbTJLlDIyDn8U+aVMZnfhUCN5UHe+eCwtHKQdoSQlHVPKNxsi+
6CHJ4+bgoxaSggdlPSVckMB1fUAyCsHbJuZxh82RvnjAGjt0dkrN0xQzbVlNbJac
icaUTqYfcn29HNKqreP4LMzVUpScZADfyZ8llFnoXMeSU2OB1JFz/+7CVN6WjQ5H
ciNGklFdHOjfJELJXB7FF7sxbNpX33BNVYiP6cQHWIU=
`protect END_PROTECTED
