`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Kxjsn5NxfH64mMfr3aYt284LPzxqrY5ynkfIExAH16XPcliT+cc4b+Mc3VuuNY1G
fR3vHRR4HpYeibr5gFvWqU+zDKiAY7y5LsWXnEUnKpXseH1QMll/feGD6SZjR6+D
4OA9qw5bLMMaBs0BtFV3v+GvmNxed2WyczU8x7ixz6KSdu/O5F58U7egrlofkD+S
W/SgdtYWfmrh+qgpJVzaObl36xdwu7xDLxUc9px0b+8eR6Nhmre54bOBFChKYsTe
mYKdyeikHt36xQfHf3hTi6Ek/RjxVJoL9Oq/FHN1oBF0wjJraDjqxVa3goHiH0HN
CJ1SHpKA+/81/DOMoqlwGoALcD1iqHdr53N2LvKY6bCGVd41Pm/6AjLvW9R+ALyJ
B82MZp5UB1eazaAvf3ONx9WUqPSuAJwN/8QNPBUIHjgImAQgv2C/1PxYsI8OyhLJ
Pouuz3EBugE6FdNzeAOqAAqBmSewilI6Tp3dLStl6HtJ/U0sqgMhYegZRnbq7Uba
eoIHJulVEWovt4vaWJfIUfsFavROA/Oh9TfLWrKVdvYk6v10wtzPTYifISIof6I4
bL6yYdWgG3jHnhAe3wBYbmFOvzhD7S/ItAf+bYv0dxd8VuWunAYIWJcZto/vXGxQ
IJsigivrZh6cbufO75u65vBqI+rXiT+mpKaOFYNWNJ0DIoYYkK0jCp1gg+DwhaSN
LdzAXJ7EANLfMj8p++IAzZP/cdEad9gSvvf6kqU0cubR9Og3a5DQjskcUpz9Y8/7
kMh/T3tWIT5Zuo0ge3olNQ==
`protect END_PROTECTED
