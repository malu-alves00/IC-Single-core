`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
t24UCfoFRjjmIUhDsqczPogmTDDxvLwjM2KytOgjPaoC8iBXURJ4dF8jddsmuaUY
YLXP/bRwsxnXS+7kKgmEV2PrpSRIz9GERLYzNr7QiuiaT8N1hDQkoS1/hXihTeQ3
L+A5kpkc0bq+XethF1NVVKIUjg7XVXkakLQeFkrN9eS2xPX79S18ecN6cxKhrHcT
VVXRyFIAkGXfCFQovJX/0ih+NDrZ8P0hzMUyrY/C8SG0pQNR4zD+w2uch4H5F4oD
hN4kEjb46UTLero6NjQ+/1/w1PKkZFKznJoBNL+gEDqsi3+5qWUlNtarGE8pvLvx
6+62MPbcUdV7VUIk9J4l5i0Jd0rukJh4rP/AID9eFSYPnh+V2cfWLWtMPii8Ft5Z
3Vkjat+ygQLwkXhQDByw41aTFjE3z0nxblJiyIa9/HN7md/uPRw1iXjQ+7vpwqwt
5fZPNCghUeOHyJnLi2BOQ+vhFXwDxWrZpmkwIomUkTPCYRHJeg4hVhBRLQPBbWCS
dam1GIPko2/VicwOJPC2efQarkYjUV6QNiEsAL33oleSaNNIc/1kK+0zbFAdNMKZ
g7JlTJSCfcuEcxvGbCojLTStU33SMHmPAkQji7ti5pKrqUAoLy3qtbPFRKhIAKQ+
XVWvNkMgO9ua6MeX480LgBTgo9V7YRR8Z1K12UR0iKIP44qbDn+w0I16Wlc1Kxdg
r0vaOJjyRxYePADHwND5Z4kk8Mwf0iJ8H/jph48xolyzGu382b7NYMWz+ZY0FIrl
5XeJG6jrAK44MqSpgBGgyH0AG9K6a0AMy+IE1aONB+7P08T3ksut9fHeLv0rZyVW
MbhdMHxNvVKvmSn1vW4VwwEr2s4iLj3s9LwhmXIgFHGGRVZJih1VMjy9RPwOig9b
7y5IKZFizGxg8Bqif7prUyHWc9YsEjoSUx/GlYFVGQYq6BNYpfcVZJ6qf99gjZvl
DAxpelIPwbcLbDWJNrhWQh74tPuRo2VG3kI0qSt7Ufxn1XFFHBaekFP3SPg38h5V
EKlhcC3R+ZDPFFNZhp+dhOjsApiuhEk863Yk/Gp1FK1hZz3gM3znv+xOVrAZILit
TQkfp1dMGNQi297xSiJPOu3ievwhYyPN1wuYL8Wz7f6063yBQlcZeN80n5HQCoXy
jfN1PTP+7dMkRtgLMMexrwElArN4onu/aogPIRNeSHx9abxzEQbI7sW53l/SvUvu
TKbpiROKjnO808JvduaPPteVuiXqX91OvUOgNSkAjTbraD3Y00UkvjwxQpbYl27O
UkgY+POcRtThcUeTQu3HjPxQUBgSyT8rLkHx8dU/Bu8bsvYN6tAfLAFHmyd0hbzc
wRzT1kv2zEU8rzAqaL7rsD65j5qite22nUYR3e4rMfOUYCIsUcJu8Nr/DsWIZekg
qzYiDE0+IVH9563g7nWkKE1m1LdHDuwdf3De36s2HY9E/oZah5o8dJaGSYVku+I8
FeSywnb0uTcIHcKduthZZL1zrbO4S3eqL+Br1GisII5eWPKd/hbAWwFy6lVEFHKh
J/1oiw54mmigAFfFbrQo5tYM+WquUZcIYRXhyqNnXj2jPQ+nDpgMi2mM8yHcT7Bh
yJcWJfiX2/b4Cp5mrsWBJe7/hH4TJQ9wGa6TtDKDkznH2hRhAJaZYjUDb2L806Jz
hXlYF6/VZeJt7kdkNhet7TztYriNC9IiJcgwaWfZu2l5bG+dedB/Ib8WrQyZtzgV
k96Lr2jvKxEWPtk2jKmh3XCCQkmTP2xoDz+xgYAUkg6Kg3QpZgB3aY/b+8YGQuvw
vdf2Vdg0k7kQPmHm/OHNrizAr7j/1OFxk3ysGQpVO/G689A3zCxRw6BcUoy8LCtO
A0K/jTdxKBGRwtijIZupxLAGVGvuitH2QHTHVCAYjGF1qewn/yYr8thZGrlXYUXO
fgAHmP+BrlUkSzkm/P30GZ5y/mY04dT+qp9lp8klhxv6pXTQMsSNgndhffPEIWrz
ME8CvsQVGPWRLxUrMHm65jZt2EI/GHRahiqbIe5rZhIfaPzbUwxUzVcN8FkpUUJm
r11fwPLB9cyN6y8LqkpHhzeJBwvkoxLZp8fvH5F+Oc8Nd+HNtYfw47XRbmCUg4CR
aB6lYl+fF9WUD2kXQ2Zjzde0cNMsaJSuBoeDXdMef/gOneLWOO6NRm7kixV/0NcZ
9awQ4LNkWg8pNx8njnTziDx2Ub92ceH3qU6+7aWyBlbBLKWpAUvezqiQTsS9Ri6p
cH3P3ANK2o77XZ1MpguL3uQ4CpuEn5bLQTWi05xOdIhiJyGr4Mex8YvmbK+MGnTP
lEry5RJ/+cDwJ5kSVsLrJPrXPElzTMxyp8oFTLmBorZmU7HRNEeBicoZfUc/mh8L
GLJpU3xQMhefujXl+6TMJIr5LgAq6RC98KjaUooKRodAtOtGXZR8WyK4ZZcMQfbR
Z0V7ApQRbumWq7pwsTvVXr0cZ3YnyOWvGcsN2SbA4bj/VFSf6+nlgvT5uuHJhzuk
Hja+FedAoAu3rjR6zSrpsM+l1u9Ocbf7oXrE3cA+alVagqtkaWuK8RCGLSTI4Fs3
ZNuLJD3sHoDIfKogoCoAb8hhs0Qm8//2vzvbibcfW63JC6r2crP4Ljkr+q3SHnkc
nmqWJ+kJZ5mJL9zWl2lABIZDaP2TesilkCPhRFyJzmQJvZnxTwBOXox6xv5o2XkG
w1rSOBCvJnENcZS8p0oRGYTuYgXZWs7S8Il70Cq7Y1/qwrcpm0CJrH03ch72etim
+b2y+mLzRa60TSrL9b7u65XjdrwMDieIxDhBDN90b7L/K1a1SBH1rrnLZJIceW7V
fj4/SpQrBSxWdhDmTnKhfG9HkUO+pUPJlfQjpROXlYfUJAQWlfMFK2Wc4Ob6rNIj
onbfzoeHZGYfZ3cMkndFiG1o5HpC7oIdxKVxFS3iBhc+vT5kIeHOihzDyZLbQg6S
jeVDO8OfhEDj/gFA2D18wJGe0ATiWWhOwCGlV5kr9b58RmWzHpnGFoQivK2rELIc
wnoIvHISK4YBGh8VyvzHFL+FFHbmWMIPWOEJ0DxdN2NWY5D9e33IQVH0XDBqKuPG
+4bN2Z9gxkXPSq8LHDNFNrr8hTqfEUNW6A7W5xjEK3e7hdJD7gMmHDQ0pHtyvp2x
JhkqrChAYxH04Uav7IJ6RavygtNXo+Vw6hcCUEBqjFInDoBiDBCC+lb0lMtCJD74
Aume9XE9yMiWPn3LYZ842T5DWeqO+w6S4XAVsvJJiAXgLP4i+DY9yevXlymj24fk
zUtbWCFNwDwWEMjtyBgDwQ==
`protect END_PROTECTED
