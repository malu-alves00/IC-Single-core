`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kLeaW5JZAZYdc9bKgkovv5qc42aLifXUYMl9FvlQhW7iU8RGpfccu2alXu2uoz9f
ZZFPJ9zmg+CpADClp+q7MXHxyciCEeDc6P05koCUHZjfCz8U9YtciYWsX/mrwxoI
OoaBw2GE/puzW7PAkFSBF++FmB1UVS3xGSKl6PQT6KP1cXlYK1iX2rO8yxHa7ear
HHpuPQsFLQgXyp5ibLTi4t60HXxmezoDEEtJ9AwOfmvQZJiLzZMcWFdC0UGffLuh
lN0aKLZpUvmUNVkagFFJDNjreJ0V6l60zo4OCBiKvmDRylEqp6AmoXTLSNRqpCtQ
XTazwi9ZpeyvNoPKlk4BIyxqlMTcVynOHNCmjEIvxBszhipLtd47TYDTu+kJq02V
W/XJz+QdhZ4GMDMOwp5bgM4exjytJ7/ORYybZXRKuwSjJJ6vfYJJGP2T53H2CKQG
7beP+6Yvuo5DNqhbh+yXIxL5NIUAgqNPhRvxRunt0ZzfQZO/BQuC0Ehb+IRLFsmN
bSSxz7by/3LNVRgcoi9OWo0h66mdRMcSIHKFZ8NQ4Peq5nnNxKEAofbj1qBrqoZH
xfILg6WgDFVpADdoPu3FonADKC5Vgwr6banxdUhEBQ8awOHfFlZpWiahqEdKWlG0
H63R/ynfc1cR6AnGRtU5UyBAwGqzi0Hp24kyFJ1QuTA=
`protect END_PROTECTED
