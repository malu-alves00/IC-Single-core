`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
I16+TmMoGPMQXndKEg753vRGRWW1gJs/Lsb1LETVz7cDlAvAEbwBFWA1eusu9h3k
DVkR1ykTbQOYkHuIAvU6P1LfSpszoMnSOskN69Q1sjjYbpHxDw1fa6miJd1dqsHc
tLCYHDr9p6jZ5RT/vzGnk5r86M713HG2yxDvGQOsYfBo24lvourByFEpBO+BlnyA
lltiQ1KDsuplT5csImILQBvAzQRgorM99SZW+jPdK5D/HHdDNv6tf6ATLksjH7jB
JZO8WdLiuop9paerK3MF2Gm/9ChOoBhozQW9FgUwAFuGnxzlGnW8uJ+C6C/4OBM6
/HZzX7SxbOsRWJd7SxrHsI5aOvT7K/gAz9lX0PdofmFiwMn7iWa1+hUf/d5tOccj
o27taZYsUwgJtSIBkSs+LVQUuPju01RQ57szgJ4rTllQJjaGZg11+rOVdSsIiQK/
e5GpMCpwYeVgC6W7Hb2+F609pVcGiT1CugDTVv/eZ+hzm9dsOkWacsYID1D/8zCB
vf+xiS0OpgRJluMOPiOspORf50CeEJemk9ZBcX6IYvBkFIv352UcwfHHa+XW3hpv
9prwlpfUKqkw04/HttP3FQzs1Lr7emtcTqsftn/gsCmB871IRfTmL/FSap/2mhEQ
FOP297yFN60dJ9UYD3bo2a3sB/a1Uw5xRVHzxfyVYZH23nf7MHvewTTA6R/4SJCu
AwP2SnjIe9YxxyDPMPMI92KgP/yuhHSyIej/7vlNhkkIVUbd6ISmxqp17+Ec0sKQ
eXhDEEt3lC77Y53WJqfjsb1lYfHOJeOdL2TJOd6HIQwR90WsRwgJG4LSajHdmAd9
C2Y+Xjp5sg5pdAaYhs2EhiNu9wOwq/YhaT09n4p67aLYhPp2A4eZXuI0oHdQ42Q7
YNz6Hv5xLAALVGdTSDpri7h5bpwu0zCXe1MG3rTjQGrCeBBZwVlCOm8DPhNuBWzf
JNmW//m+qP+K10tpaaJgKWHtjymS955jSlNOi+ess69xYXMylaUMY393KE5zJCqv
c5fmyZEnpq7DNLFSdyxxuzn5YOgMqOvE/YhVe+XqCAnEEse6/Fbv+lEyF4N7CsCm
XfPusOorvfJ9eNOReX0dukhvwIqWxdaO/a9UyDIFHmWhPWIoZmnOAKA8EbUbK3qy
637fp2tXjFGnBTLTYUo4O53FO9BBneP4Gze954U+I9y7qEyrq5kXaxhe1YngUqoO
BP7ULjqT6G+Q374YYxZOECgIF5ioYxdq657HjB66PHghSsZFY5IHmpybi5X9o34g
zgKVCgtu9DXDcxwrdQa1kheY4B1fXL0j9Nwp7tZZGT05Vyv3oGZW9kiYSOWAtTdE
G1gCTQDpgq1Xa5HNUm3qopCgackW3YiDpZYcRCyxJL5m6k+rHdJH/QLhzbXCYkjE
IDBwP6ZieJ41mJIgs3I/HxWHxLWxkc6ombuoctK2sx5xgxduWSFKLl+X1RnWkxCR
UUJxE19jT7eQ31SRWlLJHLnYxtCvyE8BdApouWmFPi00na287GOMiJOhhz/PqND9
4qFxzIKh/QnZDo9OXSUE6Z/+XfMO6wswUOUeQFLIt6ATTgGCjwwb9rUCrLNy2dui
8lZmtjYvZESiM83/3obHD1PDwPbBopi3o07wHT77NOISOsAhqp0clsu2OXFMi+8J
0VwjaPISxAmLWdGJx2XYZ3eT4gmBssOnBih5IjusF+ejNmLWFKu4dSEiUrm6Lajc
4X3j0tV2raGC93dfqNl+nxEerM1rwt7662VL86HCuy4QqrTqmnuvZWOjd4hnjqKE
WTlxhPmIsOvOvwAog4nI49gEyoNPat8TaPjFOd6QMDLTi9c89YyBi98lskKwkN2+
0adehCkT+yZSnlNwSD4vyKUN703qSFcsyg3+5dYBnPlWkrmbMec+OererpB/7viy
J/UL+qg0b6VtdEIlJAJJ0Te6L3FEEVrBniskLHLSLKHn+dIzlhyI8nvJMgI9Jxg1
`protect END_PROTECTED
