`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dNOBZhYr2mfuPCICOR6tol4QV+XPsMaMfBfHRvZQ++uDkLL+CLKCbbT7z8PfCj1m
St13qw81VlMDoWOY7u+V4bRowEq401h2QePtw7dBXPvRv7Wyl4Cgvmrz/NLWKhy3
n6yJQatTDiz2woPYLkOz3g6h09HJd9d4PaFNNSomd5xUS4Xhd/EIlL/1Gf+qwyZ4
TcrZqn+/ff0NBYDOScDz21qjDx4naEd2sY9A22uS4ruhENwX14lByL3FrK+tiLNM
kPxBuC8rxty2RbLWQb/T6WzqnElO7pTdxpYiQWRhHrHDRBYDNvAsaseMldO4qAX9
BiWh2crcrtdab6oI203P4vJmZ4IfsNH1QjBtrjdWCBBePXadxBECe1ehhCaCJbN5
EQZ/8xziOEV0QtKJpehN9iov/V5Wt3UeEVniUk8C5cSt1NWFJYz4dzmInHxony2q
KTsY3ol8pPrdurT0aM5LxCw9cAElEjMV8H6IDSYvX3F9jsR5kTZJ1mGjH8eQzm91
hctYJf2MTfnQy2Pg3Fmjf7J53wc5uQuCBo92vCnzpMypmytYNpiAhrxZWMDEzuZE
5GAkfFJAYe1NGTlEoKErUIMvJC2RyxbQGFjmFYtkSj0/pAkktfGrGVntMp5ahOo1
gEX99VUvd7UXxwZpG0CTPVUakmz9Dmg3O3xTXPWkdDixu2nZP3RHLDSipOZuqc3i
+ai6rpbP07lH8ZHMEUWM2wdew79uaG3awfj1rfqwNiIoNzw+hlj5RndxiiS8Z7Gg
42p34GJFllZJSEHoblXZbREGFnWjuP2onvm7cbIibsX4LyofDi86YBIBYA8kkEwM
0Gzfi0qd0d15MgGMrKE05zi4v3cfrIEEPiZU/R3/LXL4YPiQz6JfWkIICNNO62Hv
qmCyJDAS7hrtx+UQU3FY7jA9D9T8RCjy1mqGuL1MQ0UEivhOvysz8d5/MGkm0Lvq
DU7dUdxzfcqAu5xIMvtjuZ94pIE92DPRewRQGlsmA+z2GK/EH+XfOGOH2bgWtvJI
mYJeKbeQf2CDcsgHHtxzDbFD0WpmTEZtill6iyLxtp+j5HjPz25LThtA7cyI7JeQ
8gaZR8Qt2rseRnoEMhkGsQKl7K/FCa8fgoYuxdFJFVY5+DK/iTHvYcqByxhixKJH
Hk5FAtI979ktaLNuHJbqL5CB0/tZ3oCcMbmyFu4DWY30tfTtVXSOOBMLtAie4V1J
uWdYbqYyh6fBTRg4iIaXX6d2oBxMKRrLJRvhfMwzq9SH8kdga9/nFYLEAooTNz8E
BjPW85P1/hCqdxeMxHQDHsfEFK0ibPwsSeNmwW/hbE1afNtF40cdBgwJebpl1hiK
nxwQrzzYRH4xp5l1ol79RA3ZF+5F1G7m8DDCCib5MntmbB6x3Wp6PvPhsIFouXSZ
GPwL5R31+SjvLYx6JGgf/vuZEHfPlwZGKiq+jXCwXVC5PCMIb/Ii1/KTPIpH+/ha
WcfYsW2nHUjbvXSUYJaLZsVkJEwhOXVG18AKcE9ev+k4CIOrIiPFq5pBsY2/kS/X
4X1oNBhBwSGsaEjGJMjGoYk249MzAu6vAADeafgObwSRzml+SG1k8pzgP7iKQqZ9
qFeVoHpJLyymfMDfSZDk77nCHWzk+mj7coKRj2W1b4srdxJRr6S8VsrlkdVyjLxY
KQmT1T9VxI+CtsWn3WWSePr2fGRnEIwwNqnc4nAM2WXE1HlU4ujYEjog9Qh+lqpF
uDB9WaEQeaM50l+iq5sHm34nPTIFna5znTzUiGpMUen5+9DHS1qU7MBKxf0tjITy
fq3tcmlmYqv6Xeh9AL8j5U7VBtIFcS2txozs2k0K+Y5FionHXD9+5Y3+cX7A0RV+
imqFDIZR5WHctP1szDhvK2qZnmxD7fzN9JfK1xsSpsJxsbVk8iLmiF0HI+UCrNl0
cSLwYrSoyzohV868Q5nseHiAu3P9YcUgMVwndH1/h/cAYmq564mZnnoLJcoJ5djQ
CZwenZQzyUOyQUn+Iu+1jN4PdVIh3ZmNu++8m8uCcxa6roDasy7LnLrtuN//oXPh
uSevZ6YfrnDtNF+U6v8mEg+8F/C0xJZw+BCGCvAqQhoodL+Ps2vk1xTcsNO3vmvc
/TdMgd8XbvxNwn59qUz4q5DxeZ+xKxgYcVje7/n5j2U+wi0ygIBNgOnG+vWx/8cJ
jXspG1lUbGOZBuho5KdYhhRkA8syY2uW4jGCVgTE99MrJ1p51W4CWpb1LdyVaKhG
cpGeLrgbcf7rSbq6QbxsrBUm6iNKQjC3wYgyrqabgmaeJPz0jABtO8BbTy85G5cD
64Tk1fmnwJd2J/L/lNuA8Fu9G/SVaUtSMBGegHJmdqniLXgD1J+4D4e4NZ0bIUw1
qBED5DYhwI2yaqRBeM9DKq1hHugl4PWHZcqO8sh9sL2PSDlvFm/m04afOeGqOwuU
f0ktcql1YnLwQRlHrlWXXKe5FJ+bpvJhgJGUFNat1/ioVW6vJm4ZZRXrq40vauRc
5meUUOwK5067wvOO39DZxc3sZFxed205NkJpD0YJJLwbHea+5jCg1IgzTfK3TKoi
u1QL8LGxAC3HLCWtVz36SytFJ9UgspC9oDatXe/Mcnt47IRjlRcP/pWnrUEsDFxE
w9RFO+5ebcnGlmT/4D3M95WFADH5Xi9SZ6qQwTLgBifIIrP57Z+VjQehDyc5SBJ+
/PiMRCA//IezGjCaSJGLwGBG+8WFqTjdEPq50kPd4skL2rqLR9PgaPZZNk8E/2OD
iUPkEu79kEHAQbngifuP08yXNzoOV023ZnXv7yJY1nehgdQ6UVn5kHqKMRGcwdR4
UsEZoPwsp/3PGykup2hfaHWJsZ15xeWf9ZlgNKrPowWRS6FASPv4kODGm7BVolck
eUDPZ00QSm9p2o51QQdvqOV75mF4tkHmzXyP+HUa/IK4pmSE7VB9XTuIm2Qa+hWH
rDcuny5gO1MG30vP2Z/YvtlGrjSgmQkbspY/YlWNAwCH6pCRNgY5SMlKXELmsmrS
8neo6VElCOvjc0gFUKYg4oJwhFtt8/PN0a8vckBWDbrW2iEvfQ9ssCeWFmVn5712
C2Kq+q83a6Y9FtPZ0M3BJJi9iKpOkoWymxNegYEfy9nDEMhZbc7pSpgVAsub+t1t
J57vU8YuIKreKf0/d70bVTpv8US1uwYJgmLjtteCNwyPNeSY7IMRdLxvY+Sq5NQF
l9N0AkkunFkP5+rDulbTbXpibLfA30rz4EX5EYjb9IkRQiTOsZPRBhgZevPCYiMT
HMep3m83CRI0HaqlMddXMcfijFNDmM90JpwSyZ/HsuL341cFPuHmOOdlhEogRGId
1XsaCQKWEWeASDZi3uzLPBrNx4UjLKDeAXY/J6czTjMnV+yccYd4bfjvfqWB3J4s
/ek8Zeyg4lJSqZ2tfC4T/FtzwYAQPJdZzPy1fbCwrQOjbaYIG33yfqRA2LWcAB+F
eG2MC1DQg5G7ywhAJ7G/2OYVSTzWvCSwMoEUdbbrVdMTTtRqlDOBLUwZzv90jfn1
yZbU3Yxr5DI3cV5+pf7Te7ScVizmS24lzJmHLrL58HbT06GTh6aASvnEt+6bFqog
n5QdSB50EiJH5v2WkYjN4lmpbUkByBPw4OSCBd0HCDNc0UQ1L1CICsfWq1QiNW9t
Bl205pl4dVLLNqKStG7MwoL3fhvkYlJygkffD/fhWStr72KBAMKCACImwZ2CodCP
KJ/ObwD8sc5N6hbRcpIU75BAOuCIUsk9frL4YBoGTtpd9wZpODBsoNLn238Q5j84
3YEJUeAyg+vL77ALGAAdgl+kBwtehAisxefSu9GmngKGl0bpBD4mN74rMhduio8k
+tUJpdHofsoleLSxgleb5Gg0+6j97y1LxfUGzIMUfeFdpt4PWur7JBgaBznj1KHL
46VozSsybPsL49s7FTZZjmlib9E6TXj/fp1HkCubpzxR7o36HBvlG26FLFHJWkzE
X/ZlAmvpZErDNVRIBbublkKiaWG/vYiPD4B5cN8c/h5YrVaAcS1WboHJCTisAKtr
05EV6vVvpdV/a4eeGuR7z4/d+eZnYvel4oA5ogjwEskFNb/g4KpddkkSEvS/2ZCv
UDIzfKOSJA7T1ptDX/KbpJnMhgVQahPpPDBLeLanThWMd5TP6onGuAwHN6s5EmUB
20QPBLVRSS0u5tk5ZJXxa+ZuL9Dx/ivgR1FkFPWOLBixZNyhX8w8EyudjsD2KhLH
URq+qZ5vw5Yco8yYHGArzcrSB/5KVQOJ4nXnqUjWi7oGwV01BQAWlWcRXBp8b2mD
1U7dbj8DR2YC5fUoZvZZ1a5V7V3Tyhg86Tod4pUDc8TIgln5w50ik5KLqCyJmpkB
pYeb8mu0C0lLE5oQozgJX0HRajlAKJZMM/zBVbrsdjSMlcNiRsu/EkGOs1k3m9gq
uZN8z4dIqKqH2dW7ccKDRzcjXpEGtNBSxybU2RrxsIJWOuZibUXX6hnNgV2D9qQG
LvY+w55Zh5sSnglyai4NAnoB3AN6b+JtwN1zgEX6iYlF/fCKx/nq39fRo2AV5PrH
59xh1lY59VY7YvgfR7IJWV8TuKHtMz27Ip4fz38be9bM6muu0RRbafDzzVB5Dl/E
9rh/5Tz2XKObm6kdTHxx7Cq9uYsE+gd0dcxjMwJcxoyVQlkjJ+c04WVkVzYT+qgZ
ZkoWj0g6Ap4cfxiL9KKpOmJrCVoQxvMB0xsZjpxPE3qf1BopsX8BR+Km9KsugWco
cTLFFCIMHIYGZlCh8NYmcg8NTWlAv4nB9W/d23XOF1eUWQMR2adnUvIivN+8j4xg
N1xxPGGB4z98DV9c1Nhf1CdKd3mAe+sdXQNCvN2HLIonbAMyS/p5biGJBL9RbYoG
rwY3NQrMjkBBEeBIO/uNB/2H+vIJ+NpBTmjEQqJU3WoSB9lo1rLwN4GjHhADLS4n
BsbDvrjxSUQJE9kUhQnrXdevv+QFVOlk6kPVdXpbruLHz7WvhPzVIvvwFTLQQwOe
ILxRVjjhcWvrYPGmOM8gCGAiZceGbBcrhYzKW/pPoHAIpniNJuig3sh/Ful5fMH9
fW4W/mJKR1yXp/vP4Tny37vmjqXw4xXgNURARvivT+vy4WCbYDR1/oe1J0o9yD+B
B53rDIbYM0uWJTIY8+c/m2FrKdqmKySAH3iVDujvDfXwWDuWBHh4RdF441tmmTxp
fLneuiq4UzoCRdukQSPgwaJzo8mBejzPyIU6hgC/yVFzW29m/jAodFgOoxBLj1lB
CcBCqwhT5wfoOPoyJNSS0NRP+cmvfl6w4VVRJanjn3wSKiL9nO1KmZFofofYYUN7
vjf775FSb8dfWne/a2nh0VdySYPMl8LOxOgNr85moRpw4wvRToZWmIStd6SG/9uY
Rnh3THAK7KFWuVlpjZWMMFhqa0Y0RGAejEosAnhJQ/2+Lw0np/W+rldKtj9p/l5T
Ea8S3g2DIzovyZWhUPAMlkO4Dg1rvw9wCD4wLn8UxHvsgTRP4ahF+xB8XyQMc/Gg
4P01kiZpj+CXPWSd/kS2IemHUJuV9SyhnxIstn+eTaZVqyMMLCQLnikUr2HxQsy3
wEWYAwqHM276iVkmrENvu7lneoh7j8a9v4ghILYBEgN0G3jNZkTmRU2W/iybGJq/
RfYV81TYoSZEOqdmlkZPn/YFsIS8NtHTdImlxomOlZGCmeTr43n7jx9NwiHP5yhG
9VXf3B77xHZXdw7IRrgo0n3K1abEvV2aiDkGUhiAd0rJrGwN8hpMR5Jpt5lbeh+4
Y/OluthAOIFoVkzLu6rgFhhyBBSxpeFjJa0lfNuquyTVfSD5n8FfiB6t3KSAjYxC
/ZYhW6AF9Gz+fuHuqMLmwRbaxeKuXyTr89rzvnJh9zcCNqTpkUnsRGLHor7+XOz3
C/zdLw8xHt5dgKLkW3UnAy6W3daSURhNcj04gZhRvMVzZCh6gcEC/L2EQfBBbQ3X
faT42MXEF21qOW4tkGsJ8A2he5RcKQLxTDa+6VE8cG21QuAce53UJ2U5ny049BOp
336qoX33SOQW7TDm/WgSlsc5prSadqnk3WjhKiwgH6VJshpGpI3/5EW3qwg5SpaJ
ltt2HMm1BH7njIyl1Hn+DTeO47IBxXnoQyAM0/GvChYdMCqb5UU+BfYqE8EXzUoL
AHmGa/IJn5+CHiaFSpx6SfbqmMxNF2OPL9KKU3/5XbJ2yazEPMA1bcpLmMTxAGRx
lE9JoTUyc4eNBq9HUXnOWiMi4ZajTBrHqwb466ZWYH1y+R8cDtpWUI/zGqtCeLEX
cBkABeQp8FVXIl2SiDnpvwp2PYJPt7UXzdDEqINdi1FqnIZ5rYKzf4zt2V8zNnGA
/TOmJ2xrRGcZfzvdMAM1QIbTByv9iF0t0dzQgV9CIwLN8k88yf7H/pIj6rQIzm+b
zLzvx2nDtS1YlH/xZhp2F3VNiElZ500rb10KFObqXMMhnazBfXO7g/wg8M6e1Y8k
t9ORfxvGT+lW1pgFXWBEWt0zYrEM6/qyYVsgH0iXRmPUGe+s1W1vwoPE7vcfPg0q
DQa42u3FTQ9839TtbPRtaYAuq2P37hzEgyQAzzYoRQft9wDeVY68hdK8OFttoDx4
29NLGmdsHmabeAH4uzLiyVosv29c6baC7ON2NChZLCkajR058UnBeUw9a4fkvLlm
CbJtXZ2BsgdFukPkCiIrTmW3/qCS0G8lAuK7g1D1+snb2Kbg+eNwEy/6dnBykyzi
Nf3LSva9nZQUNWR2+DBh/StzbZxSKNUxOPpp4Kyq2/TCop0FslmkjXDjIAYEMRgT
O1f3zmU7EU41MJ+4IImj3qjOT511SyBjMeViMdeIB0LNHPyC3IJkhUjBsE4KZ+KZ
9OpK1w0JfJJ3PkDJOqzmxh6CsPxaEYE5nmFRWMv/xAd8kCUD/OmZvHfARIFSreOk
Og46gfytVBz1ovcKlNwzG62QlqaR2bajUaEQ+tx2/L0uJOfnTYuOwiqZVwOer4ME
zIdCk8h6VTf7V9ctrJJ8MUxC12a8I7QgRFeH1Pi2JOh9RuPoEteYQAo8+WhUdFLT
vKFQX4RzscnbeL2XluYwlHQ7PxiJ8xGX6MPCcH9fqUf+hEt7wsRr/Ke/NQ7gke/+
0qSgVWsmuvLAmX38j2U39BZQgPYFbQoSeA4CfnVptyDCthPQGobtYYsSipffPeK1
Q7A180yJbhCDNxrr//cN/FILRl2udD3Ek7y6Wraf6Y9ke/65Hf/iGfzsTxI/E9g2
qfcuTyTZpqbf1zid8KgJ4uRzq/fhxa57EwHYxoEdFKhzqjezIoMciFGxTyKD3VRd
ETjOBqhJEuVeJrHNXjslCOrUO0lni77U4LYl942IrPW3BDrfR6IorBROYyMIvqYM
AS4NDfmsL/Lw4uqDetBNpyvnPTi77+T6OIJGw5/zcWXXzXfD0mHK+ZEECwi98qMG
lxT6MyhOtjUUkxhc7ahxtOP6pP2VcdzEq3lhUnZP/jhPK04auSJq8p5hvTIaclOK
Ekfc/R3QN8Q+CHB61b7xXVbXCTzZBccVDNIzwzqigO8kYube7bXMV5p5rhTmpde2
iP6nt3y2EEhQzNsC8LxXbHnzVd9H3IGfN4+H7wrGawAh5aMX5w5T5B7UIpeVkzsP
c0bdZQCBirzULqV9Wf0DUHuCTlXvTgfjXZyuu0ip7KHGsqRXJetSfzCp9tPbpzC0
/MPZxTOBC3CTGBMYpTJGEuHd4q6uo1afgMfeQJRCc8cFEw4B250CCvRbtRrxvth8
18MC7jRIEx4UCiOA0UMLLf4EAqx0NtaiI2zy3JFN5BZQ+ECpMje7nd9HjWXcP6Cz
UoEoTIv9Gwtd/ANWn+72LcnN20jDXihJuozKvIp6tYLVB/vVt2IjXIIcDw97fPy4
DJ624rraiyXXb9e5hgJShhwhpNtF3E3x3D9dI47739guED2qrVyM7gZxz8VTQpAI
NRsfJ3u2FRQUC1ulUgO74uj1FF691+7LOSoC95NTh9zrPneoCupSoij6Pr4mcO2k
vsa8T4kF9IXYR+uZDYjY70dbWecMCrS5xo7gVsfTVxJut38l9rLW/QFCLxcbKQXn
DTb8Yz6PmD2vl0w5t0RHmddcUAWz7+8OD3EsojpQ/jRThz3KYD53JxCQLiQVZ8q3
y4b51N6ux3ec+GeiE6hEduZ5QXxHrr6Qe8Cu+RAnnnPH/CLnvRUNQSaIcXsR/Svw
8BGI6op2ye/IUKOOEsKWfFu5TSYEe93Oas9HXwbai0UP/l5TWJZxq2PMfalveGx8
WcdeX39pdN7m7+Gdcgtq9KyIWwi492z4NBgH8umhD54wlrqgLoJcUw84bMWG7O0U
9Z/KHfyjpjU6AhIoiBrQFfYf4RPglELbbP+u/g915IPxLQYf8jDSHsdP+97TrG9x
wflNr3UTElpFBkJ5YHTs8boWPxFaJAl53o0DZOPedTiZJ/kEZBswd6iwkQMzwFdb
cNi+njmPtE+3fPKWWtN9qBUhfU+1aecCwDkA4ScKtr10hcO2hm3hLnpSytyFJqEt
rrNNnIhy9+9l1bXyAK+dSWYMdd4K7w5DdlQ7sUZaIWG7VSWFD84MBpXyipNnIlqY
n3sfOeZzBO83i9S4ziI2Y8cXRjctmmI0GEo+6pMvCEzXK5V150dLY0PfnP1xksqQ
g584SzrBvgE4WX6mZiMadcbqWyDE1Q/MQQFoTNBVoNP9rdYCV2XX1ZOhVKsaOQQJ
6R+JB0crWQixxr0nlE6ua8Cb3u5gN8geUHPkB2yvXdGMGySpiYt79RBelzL2RloT
lqUSt6AZV8EApknBl4oOV/r/X70C2JB4ven5nH85SczUStigZhtLH0yimImOowAd
Y+LWVh7hCbRdq5kj09C1+B4q0CH3vTGCvzyuiI09OvGGaGkcNbhdwJaoMbjgwZzD
81Ict2cfobklQrAhLGssdR4bYZkYwm9TNlOWwwOn3n1qj0ntu/0X2wjQyO7KCQpa
qXYgQJePfkNxJ3MaDhbt2EL0uvMh9CWRqnk2uer+bE4N4cvLOhY4LOVCSMofkHaX
oG02Q0RPS++6oH2g2AKI1E6aXwKp0/NMBxVdk3DcTzu8y2D+lrs0wQsg0IAf/iPK
QsB25eGQA59kWJwefqHrmxGVLpYdJfdbWzW6Eh5xKyMZVWd1MpN42rI6VVllBnd2
nd0ycE0zPKWKsYUVUIreZXrey2nuVreMZpsdBWNG21I4PzotgkESPdJigH07sSM0
VC8Xg+Qw3UJJoanZWWBk3u/vOHfpgVDNuvl5cyTcSD7tGCmqX24fv2mqyGVH9BHn
cFyfJoYxrYJlc9rAtkWvGSELzIlVKThVJ4YHmiFi4PXjPAja5xz2hj2I/yOwdp/W
Cmwd+eHW8nBqxbDlIFl8nrDROx1ArsAOQhU5Abma6buVHdGMt6xPIVG9B5GjJLvQ
/xX1n0ssXjnOv0grOSV8XTkRvDTvYldCcqdhsUqIlpLer9QsGdZB2kQP1kwkCKUm
lswqBvg2Z32WU4QySUP2wfKLduHobzlxnsw2VTQX7ptrNmK0bA3bNDY9rJwP+jem
H7Ur3cDCTMurh59hYtaYjk3M03gvmj2tJ7t+Blw+bVue/a5yrbZQo0p3ZEjbRuBl
8PKSeJ4y1sVqBFL9kJor0Sx+q0QSYXGR4Nlysut1npQwXwJPDwQnWnOKtwTY9ASf
1frk6FGiSveEqKnb0lEqn79RUDzm1rGQ2kSb5S3a3U3yvzq3nr32zKWGEXMrgvql
NNSFadb4BFygTyvrCwI0e8/vmWKDD3HuofdflrqVuVl649cANVSSCx6k0VSRPUTG
J4ZxUN/hSKZtKfeKQ2zsfrT8Qs9okZD8yCeoRNqqKl+m5II9RXMacqWhfwQUSF0j
YHkruHLpGqsMWVX0SojmE1gHa0GO1aICh/VihkSN91oiZz5QhArIQ0dXETju7dU8
XgiExgDQwPY//r62xmRTGyqhB0ia9BlzQ1HQBP+2hAb/dsOchmTh1Vd4g4A6mddI
GMJkOMT9oI9mR5NTL0Mm42/9QAXAGJPAJLmnfAvUV4VSzdT62oo9vUHClgHntbBi
aYoib5Ai/sqw4bhyzCwUz6wxsloJGmj7uVZGNCZ2IBBHQxoiKj/74kuFXR0tu0Jl
LdaRA4BL0RnJxC3xEsBMCCTR5KWxsGq0paOhG6ICcYHEGrlvp6GZHNV7eQAZg4G9
kQKJz4bQCVQ6jarbzfLWRghMJK89vIQKCCcvzHa5XmqB6f47GmgtPUlOx1tySos0
gAHAR5gJ/5OhyXHNKePMmfqkPV1TkxJ7qo33qHzg2Pn129KULro3vWv6IGB/xSZ0
OmSkstcxfixuKX31US6oPYXToATU5RRoI092E5WM36AjiZzLOy+ZaKygGwmgCMfb
CRRAwuCdbZqUOs9bNKYFqmOAbap5lF4hUfEi1OmPbFr4XYUeSvueVOGc8z4+8rn+
Oi8wynxH5tTNVof6QqZKEy/DdPT9/d7+T3Zq5dTmjRJIKXrIQDbzEoQ9wChjFF0x
plYWaL9GfhULjxWUL2MwBw==
`protect END_PROTECTED
