`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
flgBMwwAXfZML38kq9x1okRGSnSxc8D/xp9u81IslhnEoW+uOARXZ9fvhdzQYalZ
fllGXvpujloO6baHFA3M4tvrYgiYczZR3pPW1heHP+KSM1K3FC6RGyPxZ1S4UpPA
R30VgDLPE+9YX5+RvrymkjPSrheHwXVNZHXacVDDIt/LF9pdZgjDfsMg2kx/OAyw
v149h1AQ6EQVc0Te8ZYRGaLsMu8kRcA/1Vav3i4TOv3fsmG0CllVsFyYbGaiKYo3
fVJPzaTnzIysLJO4WmSRrWxTq/h+sE+MeNP40XymEGnxDvxipqJQKc9yg4KPR94B
6+oy4qRVvWZHPhaB+uv3rLfL9N8S7II7Ii7bePXSVi1q9r+4Se3H/cMS8zDjl5JS
ujwNQktijigzPhLiF1IcwQwh7mghNy6dssgvQQWbz5UmEhL9Q8FKGlZlKlNTXOil
ypwU7RinpwyE2wULiY43rvEFhy02UrfVuOVHWMkQEu6sBNT9BWCGuy/ysF0TV/WK
QL8oaErcFqCyBpnSVgU8q/F6y+TyyN3z2COKa7LdgjQpK/tm0k6BhpTFN7JBnHEB
Ysv4gM7ih+5ziWRuyZhxy3E4f/rCImWzQm4UhzMFpq2XZGKQDSyMWPOD7DXAfy/C
SVT4sZZ0YNR8Q/mCiUqCOx2sMVm2nGAQma4rXbYdLAQWEP7GbaQlRDxzmGnPCcd3
27RETjUnXqwHTka5OrdWltIr75i8eomXnjMuHPUHE4Ji4lek1L1sIuEzvjHXCvik
o19yGvuoutCWfha8R6DUv+gXkleXJWtdSEg0sVXdiFmISHOHGyfwtXOuhcjPavY8
IqvtFPj/Z7DXHxBSDSaasUfdWLOekIQ/D508ASOPcgNBWkGVC13Ythh/nJmzOiox
7outLYveSX9DPkDYgwWTNqGFQytYMgBDp3onmHfwSNn/BI6DF05m/QQgId3WuGAz
5URSDux8BWD9W+csfAzwwH0zix/nRE7iQC5f7YBkybdv3knXaJpeJwLXx30J5Km7
XImFmf//Hpit2cfWgfRwdYx8KpUFEa8gZhA2/z3e2pXOVCZXbr03ckCIO8YA4AM8
+nSewpVq69/KhfPTqeO7v71uguSfmmzmLW3iwmIJGG2ZD3QJNw3or8QEpsaZMUU9
dLnAWYd/YAGRdkcXDUNlXMuKfsUHxBp1SG5knZd+os3MIO1lDeNI7/cvSE+obIT0
NjA7+PZWhJIYjCzc/yZwvVetZmjzFWzJrn5Z0cv97wvlouJHWf1oKaKF503hg+Rt
sYiwTqSDM58N5deM5yYgv1U9It+IL06ZcH1/KjKqV2HfttURLiWEk2hZ3HlOrgOY
0MJ2yeqf6CrCxltqz4eUx9rZwofPaKX6RRA7+eTm131z/lxxYpjPK8FsjQKb88Oe
nQ7H2CiCU65vggx5cOS7U1j3rAVvJTe0uWqA3p9f5LZz67y6DZHIgh+6fy78VA4A
4/TFEn/ZujViuHjSKSOqffo02MmzuOiROosNolY3OaiYMUrcfK0E45kNuPUzjAP0
l5mLBfbNOutJ0xHgTyDsE2HSjLKqkNhZBRrB2F73S6EF0Xnhir0qpXWE8ermKEnY
k8uicjoxFC27jmL9AnJnTq7SMKtijoI4zoFMBNfgnmP7ASZJDpSIZE3lMTNVEX3C
YTHrNgpXIzRwM2c1NsQ6xKmZru3ZsJcnzwk8SFI/9oiTO6lK9EMIP2JtR4CZPWxv
n6yC39Um+HJnvKAjSDiYAe1Wg2ykaCkUKNboRA+OYa3pMR6FS7su46/QRbyIFkNF
xwZ5ZUScs1l4Ww8XM731koaOIntmZFYIBx+/lxo1TX6eDomKOJp0TFvzkhSN5m90
DVp4b+D7tDPlGIqBideleSve6LycBJAtaIx++Xid8zlEyQ5fYI548JJG2NZneX2o
VjAnTrn3GlU/wnQ9ZhNiaFmH83fd7ctVYtGTqoRI45krMJPAyarodWlBPOtkN5Ie
ICAVRAwwUkzk+uJ2fC+j0o9gamk6SFXlGkJ3/6HRtPVs2whYznG1jYqbXsNqpEI1
hlH7wVlXJY0enqN8QPW21+zrABhx8BMuW6hSQXjSJ3qsS/u7sTlteGa6RqCrReVV
hVLy9ZvVwErWgyX3PaZpYLX0KU1NJ5M5R81iUANCPvnada9cc+euGopl+l2Fe+RX
cpbcQyePAUwCwCvGnf89iWLPnCfmBhLJ1atovC317cx8lICuOq4Pq+O3ZunopOAP
LapGtHLQjlKqqadOPK5v5w+T3j03WrXIGcQ+4ImrgsGH/86+tTwZ7Zxlbjxxk2G2
9oqVGrP6yifgwqxlGffi4V2EjsPitDK4Fi63/gKOAfHkjAtxlCOryIHe17FXx1lE
sTVXP/JOxr5CwEuwJbuC5CCXLavknks2fs4Y+p0jvX7FvF/TtBLqiLFKCMb8TNES
8ybRWQ9bCbRIvezmkaQ1KR4tZkIPPy+imMv7S18WWNTPhN2nyiXZajlblwvM4oLw
t+yhhjPDXaSlxzlFCm4ej1gEdIMR6hsD9AXHZoWhuhYJv8C5Z9KDo1y810QvNtRO
qOxsy+qyoAfk67rIh0t+ZqHsN+U3QLnDIE6QZ3T8Csdam63RbnEvMM8PjoMId/kO
lj4tKiaQuJtXVt5tQuFbMdD2sgGST2NXyA3fHWcUC2WwuOfMj5WI0kZWoEbKD8MG
/gp/1i1mbX+TCVD40bA4L2xZuxlSbj9ZQXixMflkrAPsNtjsg4vhhYDExuYlsNCh
DMp9ZlmrsbpszoXhiUKMVcfskvm8kOhw59zZGo67raGyHQafEwS3kwwCsPQgq/LE
NWpReNkLVRnotCSwkzRl7pJ2zorZKyjP/qgYkZHmNCayvHRr2cqlNm7KSD20yelD
/7xAIbQyaL7a68LpotMKPSTQvUsmnf+dTOnXNt/UbzOoJ9cqsFuWx1QJervkwLFI
2isLGh8H9TLByVqgYS/YyTBmRtQYmdMj/m03MM4opsz3VOfIICF1UN2jqwISmN6S
oonvB4JkpcZdu559odUIVZBISFpGXE0dk4cM2xxjqzkhterFbtsMTiYURdLkUvq9
IUR7hqIquk7Z7Lre0VwsxEaFf0bVP6h36rGyxUkgliHew4dS7swy4I6QlPXs2H1N
MNOm3rb+/LmdBKzVy99OCbxCBd5wl7a8rOggq8Peluw9hQ8X5yY5ob5Kd8o9l8dE
8BzjSFH7Zg5My95xW5v6uMyyGdAU5LxhxPVdBu3ZwE3GFaCOizZAEk5b07sh6Xs6
3mmGg98k3GCagOmneLvUTxhCYWHeqaYjXBKUt4sBKi4x09S/mcp9HRNLWbSCnwak
ZmdZ45hMHtoOm3JjlBPC02BxJHtpU8+UCPgraFI+pNK8jYPrxfVmr1HDMvq9iysA
qSqF9YTlAKWZ/cuEdz45EkC3UVccMdN524DwL1qNArTYMQSzzKJscAss3SbV6HOe
T70Z7ckX+M0xsawQRQd7xsCoh03o/Mc5tgqgIKgDMhzs2gtt7RhMwQg8/+yLW5+S
agEz2bAm+JM2B63NkIXC6AeGHIYYKqX/kGqCJFvmYyCgPt/u4tx/tAyYDRQUm9mb
CgPFtfHOW5++vQ7QqSko9j4aBMPBUGBUotZKkSjo6HngbsQS56HpncFlLFq+WnPW
eN97yTuhIq7Vl6NBFHYUALKQjxpsDvsqVpK0PDI6cB+Rg5dp2e5tHy1zObI+8tbM
QYt59ZDqRT54SnErHRrwxRrMIbEKpB1ybT91w82elQOS5KwHpHcgGmeA2TOo041W
f1vsxW0/hUp7zJL76LDQp69k5jebGjZtLIzYx1J5rWS4YVlwTJ3IkTeDebt/v4NB
pXbvfvv4mJGCMrwrVhTDoRmd2rdmR1HDwd3oWDlOy9By1fjoQ1lUDybKCU8GSvMa
K36e4OI5tWVwam1AhIXowdnMu69WXuufqpo+H20LhMfNm4gAvMu7oB4Ch87nxFYG
qJNmg4oOD2D/pfYcQbkLCbBC+mwRaGIQZxlIi3M/TdIKQVxG2Y9feucmaUA6CSjp
tiTtdOh49F2AdkSgN+0dAFiaDE2am1vV7wv01eTFzZ+SaJ5ciOTZddFHHHiWTrx6
0yjmcDemUJvC4ph/Bplc82he+9u1wLS36ksNxtEml69AbCo5xGArgQRXpkZSZ1TV
nY8BwB/r40JZY14fKC+ZFaVDT3CM8t2DLoGS1PBVR3EKbM+9EkLC2hBI3Zt1wUpX
NwmyHgVOx78TN9BvttNJTnx6BYvBpjxvlRq+859h/9iyrQ9Mb5b73FpnqobCJcf7
pZCmZnScY1UKXOdtYT/wb5sc/hdaKikfiBm196er6dMPt1KFcQ3sMlxVes5f7omp
coi5owDb3pbB4+kisMYgaGg2X+E1R6lb/pRydhBHQprjh6ih9YQG7FMmVbd3OcCD
0RO6BIkG28ALxz1QUhMI7cOh0BnDfvLRo6dSZyGK6uGwPqEeWdcT2wHXHtCAAwdZ
LNsloA4ydSlTyz6C5Bqy0MF8RT0QCL6ABI1JE/yyborejzM00dXwJTSBbac3YBgQ
3FpYYElNsXPFMWXpsm/j7IwI+efku9Y+42OsUSabZkeKGeHwc3/e4PuPNgrZkFC9
OlWFiBYbP+lVR+EH1SpByCvlxSb8QUYgk+7U7Jym66jtM/dq0mjXMvGo61brVAgi
QbFP9VSZFuwasutGMDLf6ZMvvL9P/sK6yzjaP57vcvi8DkLiYgzQaxF99EEOOWvo
gqnog1mj2UVnIz6pmUS3yPvJ3Ll8UzTQTiIdA33FU+i3MpCx8rH4iX2BymSXwvIX
TpqIFaIBNFJPkZ4p3+To24RD91SmmjCgBo60WhwX54Df/nrAvOwdOaUynvLTHcgR
w4+xt/eWV6JkBwHTa0UcXyJIdJiAiWZ/XxlJ/f3mvsWfP2VMbQsthEvqCLcrGDD1
tvo3LdMKc0/6T9EbQSkT6Y9Oh9WIFwt5zg4egQGl+O9PyujNmY3UofluqJKMWT3G
FpstW+RlFq1bHmwURVpvQL1YuuFA1CDo//XN/w+n3JBWPVce9w5wXEksZicEX19a
qx/vQBLNGBYDPreuW/zvWz7EiXr755fW/q1iHsWQFb1DTZwDHOInCKLqnUUplBwI
+c7fMqX1737GhQjKyct2AK/H83yRDHTBx8GrNlE/ha91GsHaTSgRXRruivwWz4LS
z43zF+aCBJzAQBGwGaQXTkLI64/FEVZzUJj9eEHNy8kkZZqPRtf/1B/6hu6KEBpA
ghewwJNjYeoql6oNLo9+kNjbahOPKapM4llnNE4O8EvQWszGFLDgIzLHJZMN0EmL
aR0o+DbO9aICtigQqAVaTJCAOAFt3BH6HhFIYCAu4aoBm7b8bPCNa39WxU3ZvduK
eRnBPdE3o7Tm/bPYJDTWMUJoqAzLWlL9432nWkGMZtcSinDuIvE7oIraXXk+Ir7e
260vOaD8xzEhzX5Y4i9drv0XMCODhdC6k5aHP39G1psaWxHreHyg8YpK7nXuWS98
Y/UayJk0UpsveywkNmUvYxFWk+UqwEYztRXqGUfZ8XGl+UgksjMl841Hq/h59VJv
y2zWaot/Y0myfkRcXYlMG2Ku8ZwQ3GU6JQa97So26L57epBB1MPOgygIJ8XwBaJN
MPvZ5PzB9ddTowdVpxn9K2zlcwY30wF2f6OH/HRB5YIT9P/oKjPcRXjx1wijssAI
GWpCpD+n4jSURzP2t4J0wzFNrWiPhTbFGzsleIGVl35HrVa55nWy433WgNjPXHax
i9cMlPgIBt3t0r5pG2gcokkf5iNyQzZkH01Qak0y5e/Vjzjt0NShLYZqbGWw+j+f
OEXQTGo1uY1vuVbkG5ljkcJ0NUnlWI4KeWYIn2JiqafR1ke6j3iaEJYsqxWesZBm
MrsN9qbvqPg9rUs14Y0Q5305MAWnOq0X87M114u/YL/qgMchMDJx3/gjc8tUmvkZ
QneNWtDDAQotY7/IJCpk+6j7JIHURkGkJe2578Mktfcxtcp4VFk+WsZ5GCKaLtYC
`protect END_PROTECTED
