`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
G0WB3mTTvoHg03Tw6Ulq4oY6GbjnSIoopSFAq3pJX0HupTsFdZaLlIowInQWNXXF
UgZxJ+BLUEjCOD1WZefS0cRYmDOkoQwjhv2uL6goMLthnGYgKYtNp0ORx26wRDjS
ARo4tq8rst/X4zjJfP98KAuKCxVhWg2y/iw9m7wOIjRGZoioKkCDm9TR4H7Oyfm1
HsmoipI0Uxce1hdV29KWRiqujRWIub8olzrBU/0HV/j+x/9c54PdN7KcQEKGKhaR
PMN2Qf30iG+A+xt6LH8THgj/AXQK/UOvlT1DMnYaxDeyrpzlziDhm2J9soybmEI1
UNoDOnVpZdRSbItPgtP9XZcQ1QwdRdB5kaW/44UAeLJ5XKZSpwsBXvvNSEL2l/0H
p56GZaxfed+uSW2nn9wTSacHtvbAa+BjXOIPjHgD1DY1RQPqe4v0rPH7o5lcs7Yd
VOD9XFml7FjJ1Z4pf37QQPNcv1qevkZr3diEaNbXcLiwrz0w8pnS0wY7ShZWe7wS
f6Rh8ONdNt2CdcYsR3C7LSdDVOwaZsCNZcY/vZVCtQ6QbrvlJwZgPY9HnPswO24+
HCJyxUhLWQjiDkWYYaod/zAxrA9jblAp0wA+R2mFsWXvUx/v2tVRkNqbIUvy8BzT
oogia/ycZVK2lboxrDOsd3RuWow/WaxtR0joRIYdAnpYj3tzZ8GJWkvYDRbxTUJ+
AUPu1tDfHePw24Te2wMl0kEfJBFuz6882YfQ5si3EH7BdItRsrfWiUxZ7QNppJCl
aO2HlNas4/3YqPvdcyDOkHzVSQCNGRDSNuzFChcmioLqENqaufH1ATZ1ihXHK2bN
8i2OPIGOudO5YTXQwRhGy1bSap64HLrKRcldui1OC9smllAWFZkVDsAQgYRSatS3
4rHbhISwscYQkUNvvXzVcHu+37cNEwompaDyxutDP+eSMjcQ+rC2HCeaSXX9aQns
yfXWMZWuOgdujfU2adHjKjeSUKk6S9BF3/0Dwa+ZgZdtym/UUSMUgy122Af0S+BQ
/SK8k/Q2OV5BL75kg9CSK80bwq3tkjkKQxr2xXpoT0hNuwGw4INWksy30A16ADHk
fZuq+s24NBLlEOx95vQ4jZyapw8FuOOR3b1tMV+RkS2eJecGII0mNbfdV+/4Wl2o
p4q9EUdfM4Em/PqpNNcBmb1Vy9xYUXBzUYohUsptpxidzxMpXMRULpOXO6PaUM4W
AlghQUGN+D+n4out2MteeSCFwxp52Do0ezX5FAnsGvQeK0VSKnuuUWNT5l2LsZSe
fIjATxRo8jgL8ihB6xDOBFgrZObkvarQvtr7JmnBDxm/mt3o18J/UkrnrJMnTBmZ
VET5YhriUKMLhDkGR66aAA5PE349Hieprv6As2nlTwYC/Xww1oPavy/1TrwKiRhr
l0GuF0IqwFNxpgQwdr1M7X5qASdr50WM80O9A6ayUuKeuyWhjfe2wxJrY7Y99ZP4
UjzEVziw8dM0rjH/4eOOkSjksRqIn2d5Xx4iJHdJ5PFk02HntW8mROTalpqSktm7
s3/o+HTrmtU3gZWikYCrvBnSipBhhF+3XGBe9hL95hX+0tTY5EJe/R/SYwWysm64
vJ8c9augglcaxwMLRprCL9gj727VFHzcI1T+QvIwkn/Z6TyprEOKnxiXxHEpzOls
eyH+msmqso5hEVOGrodT2R5jon6U5qlyv5pikyxz6786Zoc6qZeW8fu/LCSMGZVr
8VZy2Y9cYj0e0ZBtRdyAtItdwzumkmMMOOd86G1NOkQXORL6gnILSRrvRCDjOUWT
08UpAYsLW1l/APt7QTpJbjT4LgdjXrdNG9tesrXR7YoDhmTI/RkzKKVOjiq7T5X5
6Ik2mwBLB1xF81uOPOJ6rrp+T236TVEqKtqe619fsLxc2vq2mi/Hxnq0HhXEm3hD
TIQHD3Sc4H3zwU0cL8uTre62MkCLNqg8v162lYxH4GaPVLDy0jTSofxxgNYcVp3c
y1sTk5urYaQGUd7P6pSV2WFIRdpNLoa7oM67pRXGEIfycM6f0+Ciiq3ZqvnvP+96
m4K2W7xnyGVCnwglHr6a5NhfZEPBdf7BYM07qukZIiCgNZOBhclbcn6ZV0rqmALt
mSnq7ajIFOfaeoUcCXOtQgtQAQA+cwmOl3r3ytnQHhBePNI6T+g/Di+JBa5rbhqw
pEi5jBOidBi9YnORBWDjAPQ3ss72bx2xK/etdL0fUUFhrCzUceSB3x7HC+hHwyMb
fhaW+W4HMxducKv/3QQLxsR1dURgd2VZ49hYkiPrESWyKrbL6xrXU7c7HxdzAHnO
ogDKxgl/ODl4l93hY6DPl2bcNG/bxdnNJ2lWZdcAbixGc/in2dqNQIzJ9IeO61f5
zb5RCQF1re908Zp5rnVMj2mOVFYjsCGDPGdhROGeXJjP7pW4ZkzWWbgNt8WNhHUo
q+z9sU5BIEthwaVZUDjAOs1dP12vtZ+KNK5K4BxrbKxiP108KnB8JVUAqOP9OdvW
GxSczCPK1SbiOAbAYKFcZengzlP27IsBItujVBHZR2cvFCNoDcdtucnXBFDuSlgs
I7owJZeYwcKuvJ3svKdx0q8q6BSCU4aDgAgQgCbtdHa9Vg3Tm/qSm64U7tdU4gEe
YhuGo2XmHZ/9iFEBLqKrVWu+Xt0F7d3E/Id7qkKu83cZQeQyb9N1KWNb4DELA4hI
rd+dHz0Kl3RkIz+1KXGhvXRe2z3CgCPu5mj7v1uL/PwN0InkWwcNTJnGdej9RL1d
zDJazvm6TSyiTeuWdpjuNLG7iLJH5PljRrr8THCQlTwGBVWqVmtNx3gjFnvGkoxC
a72z8HWOxxaeo4mFlxWFoDvSBc/W7C4AXxYLKnc2SQl2RphuuB9fI9z9Oj69qD3/
dIh5KlDQ3+bVOEXZ93jv0CLRSsHMF/F8UsqE3HRcJiWV7PT0OxndRSYO3AiJVXUo
wGNCpWlFQKIg7/B/++bZffw5APiaz6L2GmDI6b9E+bsxp4KozB+8rBwPQYB328Wj
5rM8cWHpXdy/QNNrGjrPgtk66L4xjM4CqHfgTa+jjn2+UpBITmv3ezinzHhEd1rK
b7Upm58mc1+1x3UZxMq4CBySTwv8PWzTPtOQHGz20RzDC3QkYMcp6hNwTqCLv96D
tNKksIkKlZZsiQxStC6CO6Z8ttG1tDpvdd9EpOztAZLiR6GSd24L3VUWfLl/4fMv
x64u4B8FrDNLVZ87tffo4dV9LsL33hKgJXRK2FRWfcKM706uN6qX+5fJolp781i9
V3NzrdDRjYNnNvSJB/n9o3mK4rAqTMejQmorGcBbxyg3BSS1pOsHQR/Iim2dELQS
1Gl3NMDDaI6/qp3KjQY3FlrIBBYmJv17f0k4yv33Twqw8fdhMP83PAVFBF2GtbYe
FXE8OKuZJExcsbK0WIRrsBU2KePNyutKeVcUZQziGJhnM4278QkxnOL09/6XquYb
s9vbP8LQxnvXQSwcjWFTcOVohivk+ojUFKKrSyWuU4A+CiRdtRnIj4g4wDU1/32C
ArG062bgug5KM34U/4KQrNd9t41i4V+NpZbPjGqFaBKvnZzonRYKetefo++NUHA3
oBgpXNWyXq1BC0CocnGphkyLCZTND/JgIY31z6z2K2zubm5L8B2SUq6+JWHo3A9A
BP4csSifb6DC5p1EPtSUfLp/NMnPcgsCIBb4EnYO4H89Bb+g9ZjlkypWfUYkqKXk
m1e7I7ZEBzG4VwD+yx5DSuqXjqoCGXP5KifKCY2KBxxKk6zd2miBYue9a1Qn2AAg
nm/d2MATZMKYnnmWpu5/jjSofXqzO7cue/541P5xR/PKzAKFvzjulQ32b4sOrWrC
b9x1xJYuuHnBLjlo83W9OPg4ACZEk0fqxTqoDW8o3UA1Ggmfgbbke3FKxZvz+Oai
3vKjDAphqvQRDWHGKrinOGKRTd4m40sq+JaO0Zn0IZaCtzpIOJ1MpnUOlC+H6YET
8rZLKLPuuUaKMmy4lsO99TwTdpQow51WvZCsF0RBPj1a5gbodG8Vd8VYQVdjApz3
22i1IK/AXY5PeQJw6ScOJdYDSUI01hWvHV2zqsVYp06uOBdj3cJKL9fRAezpxtCO
N4vmLUNF84vsQk9OdVKkxRXW++eCDn/mdxg/HyGk22eXgj+H2+MoNCkqEuEnRvXp
8KrDA/ukaYFZGAlgLPrs4oT3Ler8Ikk65AJoQ0spAWrgsnwdgNOd4eUU2vaCQEdz
G8IPwTInGIYTCPPIw5uuCabyvNyTKWDtI8mjT3AxSI6mjPNq4S0pBsUb0ZmYyYcp
hYd7mVWPPqVUTvPARIb5D9DN5Gdp+GO7Q5dks1OqskNXWLwJR+kUPQwVRDD8gBuK
GuVJB8kV7PgoXfmmsgNpr2SJ/C38oyFoCCUEec8TUuKxbRhYRG6imiWNisygWKR2
4Uenl7rgcIUdpI9WWwVwjOZliODDUGG8gj1+y3W64UL+kn2h6WvcPrYQkoGgfHfD
`protect END_PROTECTED
