`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ht9kXv61mxKHw7nioru16L6Zkn5zUXNI4yTNJkLqFCrAdOkYVCpWeQPn0hQ9CmmQ
TiN1uYDRv/GaTm457+QbWboJi3QJ4QAYjUlf/o3Y37dP/kTNIwMp/JIlhJ4NyKFV
szDXS7jsmtPcAO+a1RJ0bVQGEZNp6cgr54MzBLtE5vdWxz9FoNPHF5EqL1NTpE40
vGzN8MO9ldnBEUD1Q4iwSI3OxTuAnYh15wxhvARUgfJguCUtc6gu7yuzm+mKgOmz
y0IiJLg0G0MpTvqtZyFQVp1aJMQ2gml+ppF2GuXPtaUmSW/QxxbESSwgOok0aC9Y
Hd4hujGt9KgRlif1SOWTEjXWCRPyJXvwBb48wwAqoD8MKFt1AQLlRnk2xImr780o
PszH5IBPR39B5qAak0X48zi1t8ozhhsG3i9PP59MgzGa8lye8foodx4dcrlEqgzj
E/k4JO4gN6MTCXLO6cMy+wO6n8/NznVZ4KzNnpGSnveVa6L4VzLGqrX3wYTRSct7
I/2RdbUvmOMxLz6br3cYGcMbiW7xmLTzmEGCOn0CGKFws4SuzMRNPOgKPC1krFII
L/YBa+ljh2fTeNJvUcSSandSoh3GbYI8FpkLboHG7d/rN4euWykoJ9KrXZraPXgl
xxz/pPxjKwv8iq97lTxIJjcaHLp8/Og5CEdctG8qJT6bRUPmoEilCYUWYw/c+gTE
LKjUCHnY4a2XgchnyurENzEz+92ka49NrM2RfIQJvkNsdZpnHQJEljqnxp+KaJcY
93XONGSMFJAyzVCHMI71rY/ptBOFDLU8bgeo1hekwd8ka3Q9yoqZ/gl/7XGq5lPd
DZ/gJlzhpa30nuQxKVqt9+d7FCcLibA+Lgowm+wrPZVHk7c6uEVZn7iGYTJYdVSu
VfO9g4kwVe70x955LFuPp8CcAZhnV4s6KlNCXMi1UgI9DvYn9z7T9j/FVLDGiXKE
Mam0JmljG99MAbt/kyRUpv6USfAlNi4D6AYfO9aNdR7PXfIEtRwvIYngrGLd8bQh
A4acVxbdZUfntPQHGKB7sRg4/5gM5oe0gAAvICKfHB164ygPHEUcJuCmF16SCG/+
MjWden/W4iihB8489Z6mhyVgPe+c0YmBYCB+oL0WkPba0tShGG1s7+T8A82/JQTX
MUVhm7ihefoXV4WMlgixOTMfnw8ocN29KOuNTVOisNtsaiJQHBvdenjzdOhwZIqS
yNkXtB0jwysNWuV0DFgXNER5f5Qd4uyASF0i32NooU3p1HGZ4EsTwfRjXXBkUg/X
kOzzxVa1/2kwhCWPf923jDZkqyk5ZyIvEEIr350tEpRs6V82KDFLj64tOfqmkdaE
Fr6cE/shCw+BOrsL3gx+zl211CbJfSM4Oef065swvCF6FORtYswr3nvYiCRb/U4Y
tCiCB8ouHw4AFkxs0nBxFpiwLDOFOGVtK28o+x0AU3Pk5u8KgobwUUZvozgdwEuG
V0ymKD16FWQFJncvqOxSnPCzb44CUtq1Vnjji8E3pRUEfQxOGFmnbk6BGEOic0IM
OjBASMxwM3tDc+r9FNLIMOibGGqgMjlhfS6HJQf+ucfM3G6QmGWaFjAPkozvv7AG
HzJL59g1RPvnOkauhhtQP9tGWJYhAifVpqGM1J7ODc7kfmfZTKAviz4SN5BS83f7
`protect END_PROTECTED
