`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZUzNyvH7fs96REp1cat7ZcGU+PpYZzVicztr/aw83kgyDBPG6DxITy73xvdFPanK
v5/xkik6AyFBQcBscdUzp/a2gbnP63uAlyZal6ifJJn8oJxQ4Ntlq2GRqt+wZXik
IEhFmdd8DYKHl4+yUrA+Ebvv2wXwIuTd6w9qqsJP3eScknQwuFmHOinr8Hfg3Ktb
dxk6BHvhG8h3P54ApXtzAMxgiMe88OaGkAsar7bd8/Kr+i00qrskuq+jh7XlxG9Z
m6T9H7facuDVhnDLIqd2DAfcZMCX3gyN4YSYjLPdh3qyrTQg3FiDg8Mjx0siOiN/
xb3FoCDzmc+RRDv5E/ogfEmiYBy1PuSJQvXAhMVKYKg7DeczE12o0qnN/msVx+rk
7Wrdg+Vb0e4QvfMefPbBN+d+bHNySs5clndAbpYM4LynzS5lCqyqBxOFNWlUvNvt
2tvk9PZAFdLAZhB9Gx2RNh/8CCVCJzd7scQfjg3/nSXXpyTOElCbevDZDRqi00jy
jk9p5QurtXoumY0WEdZplCpAyHyWIiAffIqGZNgSZmYJuPYF2ATxJqO5PhpL0aox
hQac0kBbKtkrfVIy4e6jPNoSaChk5nXtzC41U5X7S5N1dvZHVfbdCe1xZ/4rGyJY
pTGUJC8ju+VpuFDItRDBKwiQvbVDj3WJScQRNrzHeMdBGjwrx0xk45UW1Pp8JAiE
kGFG9ocfAfkWfniQpoXEddOciSw1qtVXJQET809h8idK1kAbMKxd4gMJIu/X6bNj
PIV+CyDrC+nRcZUXcVvXFxcK4VN8yjN7EP0Jxpk8leKfNMerkNFeL2xAF2PYH1fw
Ca0mdo5JqHtDO82OY1tZ1my8tEKIIVgEJ7W9fuNcfe0rFQ0tfgpbEChL+hARPxym
Wta/7ONBSUHBpMinshcpAcmImUoM/gWWElCYtmOZ5jLXlgPKrH8xo1Pw9faDLZO5
KrFkiMlnzju0tFygduNteVqWpYUVPpVbRaHF7C0IP4+4eA2mAgbLbnJ/g2ThnRbM
3foa91VQF7SL0ExAG7BIwx2dPBHsb27tVheG+5E8k7vmOdTM7jmfq8OS8wNh4rKS
mnA4e5v2VtinL1w2YTLk9VxNz4veaUmwPONLBeRLmI/T4qwvTOCOlixaBzzcMOyQ
j/4R2cioeZVxMEBqhLSFLJg53duLJ7BoymaOzowiylhzLrvqVfzg4ToaZU40LhVF
NZe6a/uF1HuKm7MPLj8jkWwwLLJxfL6YlXdkc8jQQ2HC8qBAEXdFoTud7Y4EbMaD
0IdCRIk+h+tmvtKTw5odxLNWbmRMQho8JUzJ6YBMHj/YuYNdWE5aOo/Wm+zApWtI
QV7pV54Ce03jYt2KoFu06w0iR/OrL7U6vnPTpzZT4zn8xI+mX2aD4O3Pnazne0Mn
aqLyCwnwvr9wbePFGBtwqMQcP8gq2gWoqYEV2zuysbtkPbd5a7KbEvQQyOl1v2yK
km3uRWw7LyFtLaLGYxZkHWDvLxciW9gAPb420zsSb4aDSp/okmPxbybs0ayUw/fF
oQXSfDieEXlttZjToBbGLFGJfSOWXqG2vJqdR/fSRU3d9UA1SxDlQqBXUldgf4WM
4SDaZMAjW8U76MfPykdMPZiYBnThvn74l9nAXHUO9RxixLLV7O4cG3paK8Jhuf/B
R8Z75eGzkd2e2sEsmfJwFrd3zpApPLsoU9v9Wy4gdfvVxncs/WO9AfQ23YIVAEwU
bgMDcPxWr7Is2SZLCw7otWz0sg2Jw07QwK/50oR/ZzBwMJu6g7omt9knLfCDNgiN
+3tYTEbdBx+pYTOH2+csAHI0GxYSuFyB7myTMbOxjzBqQ6NARHdqACHceWknMENu
n4EszjWWjydP1PyfDpYkPzcaMEicOv1/fcHwSAKlSBwQnjA8XNt8dpS6SxdpW8NM
m6Uc1uFTo/FEml9F3kRsh/SHtMHLVwqlx64NDTc0pLekCc46FylMeFnE6UIBBAep
smm4Ttw/1vKPRqHxiSPRsTzX6hXhKlE93zlhB6Y6hgMkZqMdNMZk9uVCrLydPJL5
oxU3xnYEzlzKEZhCpUTSJvU9bMUAzNDYYZxvS/vbcDeFeCnCYsrGWPPAERRQx3Ie
UDE7HIOgAeMXW9lDR9TVuHUjwR39Fv5j3haMJcQJ0vsMLrKX4iE/GGBgXLBFmqVo
EZvRmLrXsci3VPNCPwaqd32kNpm4plnj9hDUUcbetAHGIKAb9kuSDguNd8M6akVa
wsjhjqPCliCEN1BaVedljJp1be3e/oqIhKDTyKsw2GE=
`protect END_PROTECTED
