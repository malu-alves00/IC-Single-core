`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OgCaguNGXBDGlGfrr/mq32SmRzfAaufx2GJ5AvkrMcmna54ykcPj7jpmvqbevvlw
EX1o3b8pODXFnBv5K3r7htE9yhtzVdzHP1uzDJFRSU4jJKvJSJCauhiSEZ5IGymq
XebqJTBliMiMHCbkZMPC7x6pZFbOOuvzmkworPNB84Sp0QhOqdA9OMkNZNhKqzRy
`protect END_PROTECTED
