`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
i3F3JwcYZlaPkSFJ2VrwQRH7F6WacJ2a8xoy2gz6sfTHqqKIIrVvAYY0MR9O7c1r
dWPq/pLGl4+FYpK/xOncXrTr1Ocm0GylW3YteRITURFvD/NaXs96S9KUqAZLBniq
EUkIIhoX4NR6fNnhn80oIBptjBXSbO9UIo9FUMIsPMh+ewsoyjqsvGxSMf+5onS2
pfprI7kkEmIWFjz7kB7Ql0SZu4/WrZda/F48sOwCugtslVsV+Ya1OlGjT+qku9sn
sOvEaYSSUAUTZPIVi7R0+sjUS8LBtwKhTR+x5LohMSypWI0s7lnJfLPpppO4Hu2F
zVPVno5NAa/T8+Fp4GvvS3waY4qWf8XmFA87ECYa6AB0mMyr++9XIkxYKamGf7Ic
ZEMvyCxrEqh9CHm90tY921SkLt4/TolZwA+m+UmIO7vqACMP93ePJkvk7+u+jcLi
KyQPwRHDw8HX4Sgm7TpXyYqhHVfvrwGfRvDXBPRtCi4cFkX4TxhHCWUIPkpOkNi+
GWcEopNZAe51SKGRTKjeR1j3ffa4IozlNqKqPxLdirDOUJlPFWXEwStNn4taN6/K
ejBxD34L7NFP5s7PDLtplqLp533D5JtGfF2fRyVh8tB1UHn0W7mG0SZ246ISd5XK
frSxEInn5GbZhOGJY+LmIg==
`protect END_PROTECTED
