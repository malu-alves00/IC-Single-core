`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
opiQIkp7x9zcaxqYqmYRHXRHbl4bjhcULTAXoFsKVSYu61obVidniuoNSl1mkKSR
a0Dhfx0a4ebL7kABolTDwbU6owtnwq5gk5DceFSdcRjIvDZzmPHCaRc0Yb3pBytO
Lak5srFCCF63yb/jIHH3vW2DrzuQ895X2Pml71gWuS2ai0LAJ4TdQDuyJkYsisfj
5Eub51lTIj05un+wFgCqdgDGNBNZCpKSr9Wqxvs4XBABmW6sfpBMCrsBQfRxM1LV
YVGQObEeRNviFBZNZ6QoM2QRiZDfYd3HWQWqTwveZ2ywXnK64w1in/VnSXvmhtgE
DcegO5srviJUtQojK30zwycp7GGEu47OUZqn2Tff5MR3vGFRRqrufGdCn9L1m+T1
M0TOUqOyH8FTSTEcGZJLch3FRd5PVgzt7WIQG8dDJSPH5XXTA+Tvrj1A7KS2wLsy
6sGl0NzgEsFkM0noXwnkowRTYNUNgN/sVJggPFMWn1FVtwkpSE7RQSA5A88RW4DM
08GLDQ0au7dcczujJMGgFMZe4EtNYs+KSYxnRlDxTiiq3qIKBtMHqMK5OK9W8mQY
hWlnjH+zxEH75nzbwm9+ara4ATFJQcRf7kZdCAxXfjXQuv5QX1CZvMKkQ2l3/097
gDIt3gYzoxN5Y3bP1zHiNxQDCzqhfAPzhy8mJZ2972Pav8WvRZ3GPTWRcj1DkzW8
83GEVkmjAsBJM/mf+fF6NrpkY7+jR2wbpe0EYOa39wGfdkyA1WLnTU38T9yZtOAf
5JIiDmIrnPvw3DP427wmRHuQXr8HsjBspq7/iCDybHUSgy+C/wYN0dsRaAWCjKcH
m8JIOxU+84QvBUA98xlaXt5cz2joRZZhZtrk/mUu3ZeAtHFEawf3j5zecImVavfz
TO86yj6uz6t7w14Va0D9LkVJRxnNc9cVflGkMsk0l4LnIUIfOGhCHL8NUfClH1gs
imQqo/VL4AdAV5Uxqoy3hsbiJmtv6ePMpiUJFeTxvYYpAaA/iW9qnkoRbbX26U1c
oB4RO3WwkOoRlZ5oaTXfKP8Qkm1pW/53GArJEkI+pkiEBEaxk3CReoXEWmvWAryH
pp0KBSdSWOsmwfKmjmDhmKjS+iKBUJHf1TCcphYQt62jVCoRr+Pt3cmnQHJgjyMA
R18EgomUYT4PR1RYKaYK1IiaGSNsyznK4gX3gD2Jd/ms4XCEn5rHo6WjAy/jfGqv
krOt/1C5ZJxkQnDULnwOVG980SqfagG8cH7i9oDK4q9Rx0UKKV8cwUj48kdPiFKT
oipnt+xlS7oZX649QqDjePExT04hXmK2h/u6+UmFb0KhRahwEWTgHicnCrQQOpYi
Cv3Ahdrvz5rhN9YjRiNms6UCGLmli7K+uBTUN+J4iHrkLiyuWqyDtu8Fia0yhSDH
7TM6L7oRNgc2q8+fNviSX6As53VwzPhOs8jSNMxy5l8=
`protect END_PROTECTED
