`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
V59UrJm4HI8kFKIhET9ctzfjo6Sc3NhES1ZUYs/WO1q7jeUxXGgFsSSHNNH6FJf1
swb1dyLKTh1JUhQzEn5MHUZYcU03p+FSYsWDeS4n9h/mnDiudS87TE1en0ySYfkN
3vosZADdQZi3CUrVX4j61mE8AtFiDf7HgTFMsU8IljC+fm7bAVniRi7M4ZQjlPk/
acljPVAkywniNr0rSmcF62ckVVpPnPUJzpS/Ba+T84uAz1O5WbFXEMLZeg03+JnI
FwxW2Xpzzj2Pchp5E9j4VsrcM7OaIpg62KwOk7kDAn9c+JdefRRREH94gIGIOHBm
uZKrqAa0iZpnQHB5rZGD1fe+uKcKND5aKYQrsFaOZeYa9eMPjoz7oHjbKOl17rbZ
pstbXc88Yv7BfQpa0BgdroOlP3dAprwhsw+uLqfJs3kwKZJITlc4B84x3tdNZuFD
EC/2eSSwBoANGMjREwlZyr8h5qFHDP/lgj9qfHKUjHz/+8g8Dmx8IAX3Y61rUX3R
QXb7lwYT8/rZlkneKXn8F8HVFJACQyKvbn2cMrfdcj2vZ9Pr7r4tIimIeh+VmOmr
Q6a+6SvXi3d6C9EAhBpAKfpn9j/Go66uEAnTQaZEf/bpltr12uE2aw/giJC9NTgK
yCk9DkSmQAdJ7LnQuzc9VvoLHKQeHt1wKYtYNxXYX+pdbKfZiHsU9gnxPMKvVL4B
udx17GcCfJJHWOHcqxqZFgw2aJn/bAjXXdgJrRXB5+A9Xo3yNe2aB3UzwIm2Q0qx
eWi/8dF8weCQcWGDAlUklwjtBXmClQ1N1isftyFThJSO0VHWCjiFtDRWiYlnmAOf
hm12HAKyLTrTGCquj2GP9Vkz6LncMyt5ci1UKYvEVqEr9z1tHeS8HPyia/FDkdYs
xnaK2XQ9DkZ0ktqsEPTaG78sTh9OBloFkE7O4DuTROf8JG4z8PcrU2zZ1jHLFW9I
7KHDldcuA28K3gqYsT9Q5vatdxf/Ah/BLPxBLxRXNJxQtEJlzFbMTbP3y1wHQcUD
k/5VnPO9yP/vk1WjSLJ16aDE3xycgeZKnoV01eLbRSKpYFcEqqiZcmdPs8RX8VZR
KjoIT7hgDTnbzSYi/SzWraYDvgndZxE9IRLzBp5GcZGc+scfIvMJQIYXQ+mf6wIA
eowXoZdbKISiwoRF9dL0dqjEycMDfTQbIXNQsqo5oI7W74K77MbtAC9WpHjMQnBb
848NoLgjG8KH/RaQn7posZz6l/gAFRfHQMJKFAgruh1KgjTVAFAPQ4bnSfrGjJ1C
Cnk+sHvlsm1/q1j8brxqGfWpNl7hgYug7XwfPYQfIuffYWV3u1d4JshOEekJQXTS
7K3qcqe8SdumIQ4l7WVc+vXzBtWw5O9qy4pj9d3P97vw/nG7+1ptrWpTLrImRRkO
qa4L/sZGYb34yebiGZXuI2IAjKqdGS1h2oWFdUwdKDx4oi99qm9kQyPgQj482io1
99vwcAJ3A532zE9YFiBMUlcsS05MTK0AYsWiVB4HLQFKdmJH8LA/lE0B8JlR0jhg
5UFubPVg2zPbczWfkGTNJTTPpcwHaG3Zb7sUAxhmda7e2511P2wHVnJNYw52RuYA
TOCenILmwQn8d7FehPs5TldcH2Jqj47mrn3ZX4U64SrVhN+tcx+Ft8oN2A2EKIvj
8usr56P8+T5eLFCZRdWXUe+lh6ASRZeu+Vp8yfSvSxBIGIhe5K1/ODPOQpwQkgtL
K4KVvp4VxL7D+PHp7jFTti6hSG/G6wacAaY4M1BVWDeUW7kLvRXLVQzDdQdDugj0
xn+TK9BQF1bsQbtkYCWMXoyCGxlrdoj7yJhRACCDGKp+v6hstObdS58gPaDgIbmE
jCegVysp0AfdWv7JyWVH8R4reb+ClGgGYAa3Yk1dDfsXW9t6mdbwkw5OLZwt1hr1
+o8MqckcTIWN4RuXrqSghlMsYp+FbcZds8R+X5s2h0QpCu/m0OWgbjTyytdktWkf
AuI4CR17xeRAXQd7U7EdMnH/NoRbO+ob2zxshLPJvfJPGI4iFE1llomSnr2f9X9l
e6hOQeWm9VpWWTRtCHP7bnJ0Nx/ov9vt2/q8TwEWVln0X4z+sBgu61QqQgaZp9fI
XV7qEY0bD+ph5Tx1GYTqpTS4GAKbj+4+d5zli5IGKJAlmqKCvsFvbhFr64NImVw4
FAteKgm1joqe3va/4OJ1iwMOxYj5LlXBfmK1DeAVKQGEDVoSb0uyxxgoSz2H1P7h
mh5zn7oVWlL9PzQFaR/YzmucziCaeFA3uiovIE1OrfIZ1yWMRRf0VqMVmbJfGpkI
Lr4hSQaVXuZ3bVaIairk0to4RzHzwKpSYojJv5mVW7118z7fy8vAgcpuicEfwXPu
/8LtitHdBBpb7hOKF4AyAglOgknNil9Fensl/RGENvZMw68jl3eLbTT9bnMcdHAr
VQ9x1rXZzWd1FFn/Pr+jQHg5u+ir1uX5A/w60HL5Q+YJ/9BDBLgv3TcRe1JCXRIt
oqEu/tsRq7SsCNlpGvbgUUcfiqcURCQ6j1PxHrEgMHIGjfnwCN55DCZEla775F6w
`protect END_PROTECTED
