`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9Wa9/xTz4ayLRQ4Qdpd/IwpBYNRM9q18Xc7x1I3k/leS3lL5iw7BNLoTMC9I6jbV
yaA3L4gHKYHd6Ni6FxUjiY4YY4/kqcGE44qN3kA8U+QZl7nbeAvZu+cDsgcpz6VH
5bx051SMU38K+TSLGbxGWZvXNSAPwD/9t6fgzaxfo8gSkxa7vUesyTvUGWk2jnVl
50fMwaOZiwd/xysTWb6ho2LipLlw0Lcva4tLn9X20N3gY5W2IrTn18fuYS36DHu1
544fDQF3pLuhndHwRaJdX7/hHEOvlCUVlPeByOkIYitkkyNVNBqmdZaK82eO8Gss
NTI9914k4iNcV43L8grA0dtAEF3gsd0dS3gA5OiDX2uemzvlwOxdO+7lueA+G0sH
hUBw99IPTT+vzn9Wa5QA9BUhioBbdo4iB36LF/aSq3YZ3mGN0B4zOfV3shzHc56W
2er0pjzoh5v3lNXf9rGjUU6EGJK/XoUuiGNcuK+vxtU7ltKC2L6KJ7MDT8mTWmPO
Vwuabluy0BLJ5Vwzm1LKYOUcR3iYcUAYBEvaKFnRKuIJ9E+qPH7OlXJxg2eOV4V9
DFdUMhyeyz/BQjGa2Tw3cnkLnoslt/p3++Em47/60mNkxC4M1nmPMPteaUK2lhq/
Qotlpfde5N6t88FejJkgYtfrSXCNuVgarbPK1iTwLZss6OMRArkT5LWT+yfy0E2l
HAlnvA6jSUXcqQIp2UhlIJnzsqv1UhiR/bcdigqB4a2AkJTo3wbBNAj2A1R84/3Z
ojHzJc7bfxqxcl0kg937mRm9Y4GXXbMsMV+qNiXfrdsQLrfTKoJRt/PTDYJp/58V
iSLZWjtc/6HLq8P5eIN9VzIv0rzT4kiRzoC7fViTXx8NwB0F0HiENYgdqTb06kKx
rR9WCe1o2Bho3aAovg/UJdUyoSt7E8i8EjC8BdgYlFJAQ2++kBfS+VANT+irWFjE
9JaGBUnY6rn2V3ZJTAWWgYoc0fWufHcw5/L+LsEAcYlcDmHZ6I+O1EHuvbJ6Qr0p
ITPeYDa67GZq6KRiOMYh6X8v1xmZcM3EBIOq2FjYBCGx3Lp+n5DzKwsRN9cg+Tbi
UvZxqEaP8e9mgBe6UnMkxMztODkSBnBvjuzcRkBsM1Y96MBi4HzwPlOgka9+1Dh+
AkeWQBvl3xEI0rVwDv/sVvza37+o8G1qDYIRXJfK/d7uvYL3a/5zZCS2PfmhxeQL
wXXtrYAY2e7KRGl/6Kge/154xazCAvEienhUOKEvoHpHluSUyxZWB1tWEPSkLulP
8ZbX6FVCvdLeTlPWrhL6j+Z0sPaaD4OPAnCvwN5DcKbCYnTXA5OW+We8G1sakSit
7FtnhiLvQK0CRJD4uJv0XHml2SDDQHgo31BlPRdVGUuaurGBTnviXcCI/P//7k7p
Y/2PiFVGUg0QBEJ8Ok2268MBRgxef3yKyBDH/WluTo1VT6UUhNnaaFZLQGcDqFlu
EOt4wpaWyhreq4CsxmEFDPmS/88Oa/uPzVQEc05TgMRNT4N4gE2uOL6/R3nGim1o
6ZPnOymTVWurCw7030UmDpH95speSHQr75M0JuSSwr49kgSqsRz7qDmYVYN9G0sz
rdrelrwv5HIWMhDlDzGa58NdI0gF0U4JH0s7SHOWDOtxAc9qYf5aZ/rAvgTkswbj
aqOOBz5+yy/CkkPPa6IWb3SF0+wkQGacVtf9H6wJ0OT0ZYYg55wA7wd5SHQ1ROUF
jR6sINfboI5QMKMZlssQ5o4GtkbXolezfO9tPc1VtjzPpj964YH4qIpQ//OLjNoQ
ODYTkrSQZ4E4Ev9bH/UG1h/shB5snpL0ySgGkSmERfdHSDoUIQ4zU/SXpLwSv/Mz
y3LpQ2a1lyiF4b/SAkAqdeFt5S11xpX91EaieIYgnFr/3AYMYZDUZ0Z2ra8O98Uf
EocScgr7A+y0A8JLhfg5z95YgIfy7c4GHpQ9UAdIZWcib07bHLu04yJjhXIz+xTu
XhQGp16tkJVjX49BUZqKX/fkSLcc+JaX2pqFlBiGnfq+pRjCpUPL1kgbnpcbyFWw
l9T6j6z/97ho/BF/gDu+/8ezM5hytE1IclpEGCknP14W0hheBVzgtMIezmc6hixl
LwyUVDo3lzER44iM6X6ac9IkwoMVWAd8pZ3f+J2uRxhS6YqIyl/y4aw4aYOOwFyi
xPwD2YDZyC+2ArN8KrzbMA6CPwQNf4tDX6vPcKwdHVxAXkL1hqDaFaVk6RVUi/EB
k1fe/Expq0GxVpJW2GqnN/u5/c9tnAa2dICTQAqq8cSITFib9sfvYvmcoLPnlNJc
q48RT6RRWWQQZUvX5XWHqfCx0dzOUG0jz5VaoCvKhf+7/zTe6ZkMVHa/NnNhfs5b
5GDvK1cAlNdaI3v002KoYV0DnLoIJpFWQwq4Qyw3X41nEusAQaQojOw18uoRhLNS
GQGdovMJBvpCqBCtT/23LfGNdRTtO6PC9rLiT4BFmW12sI1HrEIpuvgNeJirKvlu
iYop4ejawgNz98vU0YbdhPb3FPG8smT+P3p4/xQuh44nwflKqcjB/tCv/3qcd+qM
yMdJHDLJc7P7nRIwAg9Ka3oosiodiyf8t9bJZwrfETBUDji6Ukj8B4Gf7DgqgQMD
L1hy/DV0Gzyo/RDuZxRO66fP1MykAdWCK0lWFcjRUHDImEWbN2hCnBgqqQUoBeF2
o6jRoangLA/VtwOzuy+xDmi37SW6Q3JRvjW4wc0MfvlUMS5TuUE54wYdseivbSig
AoRjK/wC3xGH5I0ujVzHjxYar11eY/SWknBcg0troXZaznhS5tFcVnKbci4WFxcO
34WNK7cysLaeBZ1BMty/z01x7sBjuyApSLlSHkWPnB2fPTAUZCcPTrb44ToaXy2r
50GNmS5jWDZIa+DjvsQTZJxJK8HDdDk1G/a5lkmvPJebVqCTN3+UB/viTCdwXkva
Bp9MFXKCrdlz6Onj+u/KmAxWamQ66PF5epYUact4r+GjhkKdPB3wPO/aoVFB0eNN
igtTGre/rVQtbgFUZIviVwqdpQkbCgeWVqRDtahuDSKPZHx33HZ33fxfoq+Vr/Z3
1RpcV8PJU8XTz9g5yIQK4HYoNXMbSmfyw8DpL8PyXaXOttZbnWd/XwiDoqrT6lqV
4W+1W/iwdAwitRvu1yC8ZbepbeWh3XI5SJJopJug65nGhzJrwmsQFvEn13jcpbcH
LtqeuO0qtKWM8IAvO6sIq8UVMs0G7f2LSq9OhQrDJlx58EGwsFqZ5pWliZeD7D26
DrZOZWphxy6+5U/j8o8ps8Mxf/CTgHlLQzYTCqA9Q2PDu5XyjwmzS3yf/Hfme/6T
TcqX5XdKYYRjyUCn3DrNHMUNgXqyKBoeXceny9cRj4FqCrLi7iIPBBQlr7THzGQc
ETFm7dOrmdltyYfgjwi65xfDxnEiWwNfTA3Tto2dDQyDQzsf8sc6tGYPomORzlJ1
ZvD4ibqeJb02XUOn1pjsWpFV5ubHLv6mBfHA6KZPm7gSiyuS8Rr4CX4FeTmKM2hn
MgNzJ+HpZ7MY3FwQzarm0vfniT4Xejmo2JkFGOqIFswD70D93BxgNTqKk6YZRHBO
anwgT1UEXoHlSof8WMJPVx2iCTanNaRDwd/JvmuczwYpAmG0Gp362eZqYHMyqwQI
AxV6hcPq5WS/LyiMx5JAvfWeRzTRX4cpmHmB5l7QMe08JP1HcMuygibEFIixuukH
c+3aP3ovDdvxiRNYHaMkECxWkQIT+Jht4zBSTlgpcZPbRo6e1ag8UNRWmt8drmjr
CR5UupucXBpagm/FrrEWZiYgjAvBpUNw37LeEMg3DVay1jBioXcMhGzD+2PJKD3n
v95RCZe/r1WbWlBYgMoIK0fAblxnQ7fMsOQ1GZd5ru1+/+SbBFaORjTcgsWabTbr
u7jel+bKW3bP84JR10E7nwuVoqNJZyA7rB/0qtwJ5Nx3H1o4XbjBm4IUrg6UJNAo
vWQ23e+l859fgewSBRaRU9qLT3bVgGBVhXsl86nDaMbYvBn+PZXhzhTy4/dJyxl6
EYb9XzXPKzEEgyc2XT6gV/dWAVRd2+2/AkHJ4sH6ngpk8ekmsGyYbaPSt+rl5yhA
BgscrOvFvuf4UUa/RgxiOuIfS93EB7htnOKct+1dESQKx6S7ZS+ty1bP3Zwae+jD
48bepoB3D+Dp4Pll3eY22AzDTzwtRFrl4hKkffqVFZzLNV9c8ovojTUWBCdSsgSm
yNNr6gDQPhP8RonP0YnxEBU+evgSJZMp/zPTJvUvclFyQcr2BetOmXQlPx7fvkv+
eTJk2x4h+T7kbnc2PiFiVeGjElIQ//Zau9jcvthX6IuCXE3L6GFWL9KZ4mBRv7GN
pQ8O2xxSDAatt5aauzuy3LISLerDkxP5UdV1qRnxUMa8MHdDVcKfe51idSdOHWwv
Sqm0NaxOJ38D8u2WWQRTdKGOcqgiE7LHEmF5aBkpsrhhvFHscXOmBNgUGjy+qZZU
gN9speXKB9Z8/Q3VxzMmT4Jp/kgtSpj0IgkMaurttRzpZGIwOLbozhCuqXCO1ZMS
Q+d9qwinkwqpHcyQgiSfalWrQZ/ugLh+w4F5JDofWdPcsbu6/BC1MYqznIa1oEnk
NXdv/IFV4UHAGreYPBuuXShubmNRBNgxdwyg9mKrR5KIlzO05XBqj9GAQldU9CE+
RX5VlQuxbRZs/YYj5kO2YmPYTXLfqH/pB9jsoPNwJ4lQy6P1uSH/KREIqMkEskSa
mYjHfYihvK2puc4IuI0uPbqZYqK6swN++fLRAUgB7HMqfbNKOZ3qGPBsbrZp1SmL
HkVGpRekI1EO2oB5y8rjS/PjKSd8iaGcism7NQZ0Te8kwiF0wdQ43J7Ig+L1o0Cl
dLbujF1eLZxoyFFrKxjRnOMskBif0OdJ9dUErtr2oiQ85/pQSWZzmtCmaRIOc8kR
ehopsdS4wHiPtidrw/QL4zcNmjx3IZA6LJT0uJFd7nOtyxErhZ7gAKWg/yYd/kbC
lucAmh8MDr9z2rCIVAm4VzDkPr3DywkaQ6+9yWFlVceoDCqIL1FmDms1Oy852AQd
2vz1joXIYPQwiye8vgfzZFbhVhVTdqGTlnxd4LSfxBh9pLpyIm806YgnVuFHV+5k
eNcIJXJrSC5JQOMtPiL342K9S0nswa1hHfxNpW3GHnBSiFWmgMEV98oCTcnseaxR
3qMu4+JsUpmodAVrnyB9Hdk78SrT5w9iLWPR9ZQ2oDr4Bwt6kN32/IYfHQq+uzya
qU+nzbddgMfpNs9YRnzBtQHpRrt3bHCe9sKmiI0vLFlCoQvIV975fEzomU5WqjOl
e7NYjDb/1doDccgA9zi/b5GlFkgxgIiDu1KXiDAjK8C0wjX3529DltGymWgp6gXu
uzp91PwlzLwaEZ8vQjymRxR/xaly+lMTuwHOw4fcx6EFQzfSEYM5QWGVN6zoCeVa
yjW3anu5Ew3KKiLteCDTwQ5G0JcZmqUVD+4l1mF0DeM/5TzIUB1Y/qmuTF9kIYW1
GJ7kvpIoYM9omyXWNYt2OOeqRxDwlmpoFsM8jqjOMhaCITX0GRvSkYQstKAinmll
bKsxwWIyVrgRVtMMYH5dcA+iK9I9jg/XjL1Xr/5YiHdqoPU97+jJU+M6sNmPpxbq
+eBlsXJxmMje7bp/juT/mL0QTisaAK9fUUNVP9hQhLUpgxa5NkbtsddV+it67OF5
zuuyrlYgoeQdxsNfpH0mRBGjAScmot1BUW2TN94M/SIi8MRxzy7uiKIME3BIzMis
zFwzL78i5A8PKcfGVD6dED17yCB4pqUR6osO/9bx/DOghzRXtvWhxBvErw93Y1uK
apOOmYSSVGByGirizBiVfoT2GR1xJg6foU6IBEqBO3otyPk5JrGp8gSse8yGiPhn
V2daj5wTpfgNFRWjhSm/FHOzttaRKLHf5s6yrZbinJ0SPaZIZLwDEtnWgZoAlJj4
ZEBGZ8JDEplF7SZXx2CsviEwYjxE1d+Sg/0ck/gynH3EhodATwy68nTo2ESuOmRN
wEXooFRb/th2uAKujGXylauFmeMciXuMX3inVOpYqoCbOjBeCqLDoaKS0boF0NUK
ak3cu5nJeHCJ8OAcHqUP3Mx7tCQFAsnyAnZHR22IQn+uSlgJ+Y9EbzgO1hiyEM/7
p1uRjV9x5c4D5HRnRRa52Lyxo5yi7V50ZYM5xjVXhGG6dHxeqFHDu4Jz4neHarGy
sWStXe0l82fVGQIBmmQw7mHU1okrHUF8PRdHa+Z2/L7ven5ZohIYlr8Vj5Qe/5b2
ZRKviaLIZbLEDyZpSNQGsRbYyC/VUs/6FxqMl6XZKx0Gd6hNISQLTmx14T6kqURw
m+LrQKrtlN1QMgiBjtlKGs1pB9IgLVDfekatlmB/cNC9Un6M53s4d46XIPZ56Xk/
SflE5EmS+9LXNkMGHdaTndT5KEXiuNZlvOLQnfWnjMB8/Isw64q9xgmoFSZmqeQi
bLxIO0d6qCJJT+bWPhHwOtv5nc4g6nO4xxwkOGLbGG9/oyKORHWyMQXQh0L0w0Tg
I074MZpRQ3YtaTiT7J5+DdGku1k9DlFOMcY1BBWQUd3HFk9m3A6UzRsAJNORWT4Z
5PgIxhhDYE79pW/5VrDL57yulC4m3eepAASpNrd9qYN1G3yWSQI+pgKaH2uQ+is8
r5HfTUMrZtNjC5n7BJBDaOg8Z/b0RVd2eEumRlfVQ7I5tdQDt14xkChDD4HcZNn+
AVvEAdgeKR/jd5Tp9fIQgd+n7jTAAjAeW9Nd+iVHQMlUN3rABMCBvy0kVkdB4/3S
9Xa2IYE8Uxva0EaIk3HbP06GCS2/+b45r0+V9pSKCXb2nWTNLhCFMhuP/qxx82Rk
6PsNRhSnoyPVlG7xW8P2Ds1xMtekH1MM1/wHBsJ5Z4o4EVurBMMiMwLkrK77sxMu
pRW6t5DBYSPG3BEPBd1QeREQkKpfcIeuF2NK7jozW05QfVLGBLdUYU8MqMoSRg6N
LT5gsewxTwmk1hb6NFS8Y5cIdHNUGEB+B4YA2mv/UIU68eK6h1rTkTsTm9Orbmlp
vyAFr0QAWWbVxNKdOZy+BdauaKZkoPoOEV2zLCDJKEu/vh3KBCvMU4n/F8u+t8in
xaijLAvO5Awn6AdOSZJNRvTu7kPXApCftE/sLhfVQ1QkGfLzWsacyefIAU3PXhai
qdYeeQUgwf0+LozNAWByVd+26w1oGFZXHyPKL+KoI3yBMXAeykHmCNwKuKY7L3cR
El/T7aUKns2wn1xCF8PsX/sjKYxeIKmcJ29CHx+uk37rMK1ACke4Zu0tDFpL/F/i
ykzAp9F5637jVpVEJDWOHcSUOV1BMbg/zY8hakF/x3DPPeaCa8bj/I3Vg1Viwsli
j6nrCqce51IrquD3OhtQR5rVwCXfkEpTC0H7bzJ5hytxs6IjZj24MBo6y7NW5oZS
E011Q6pVXCMGPgbc7wUZdx1lj5IxC0ypwSBc2PCsTikuwYarjGjbSZqbcPiJ/rOQ
nRbTN4tD/OjXy24huqVXrSIuYKil3LeaM1OsQlJ8f0dBsBYkjYPI6Cq1lgdzDnMm
pj4tLAkGr4y42Jj675fRbMDvyd6hZIYgxYXjlEWdm4E5aDLhYTcgo9mwg8NcNGQW
JnUIuRInVcfwp3+Zs43weYt27PzGJH93o2LW+ICi5QJ8+VOMc55Yv2rextfGGFkM
XcFCNENVRPusaoMip2ps6NG0m2kqJQh9w/uScgScUfltznGrdZZwNvTxM+Faa8UI
xxLZH8TleH28Y7xzxBbLiVBNkqeqTqjZldSfor6UfnVrlm/EpoVn0ji780SuE15C
zES1yO8xIrhCVwPdWhNrWSNvTB6piRplqO5LrWA1Y/KDacZ6TK+HKN3T/u3rFHlr
Q23krWut8/VDiWYt355GepYNo4XcZb6LT3TprZZiqXLtGWTD+nn7ZFyKA2k9AUTU
5SIf/GE1YWQ0f0nPl6V5gTswhilxmDjowHnCZqQxS9r5BrRL7F2Ev3zcCz3MP9sR
57BAEM3nYvvU4vQ7DNQvoCtNJAYoA7k7IDcE0ZrtOpVoZv/d0Yr6OLDqRt1GrLai
eKZxn3qzMh56IytUKuMf0usMKFAC5Ofnp/9FsSKZ+nxkqTT4kXB+R/0ZWdbFVXby
yxuJGMzfgY7njIaswZKDLrDoVkyyLfjATlrAeGL9cQxAMDuZVbezpKwq73/o7xaG
ze6lb5k7t21wZxtu10UiC/F59JQ5iQch8DDGixivHmbe0BMSk6uhGIQi0xK8ZMGJ
MXn+XqGh+ycnjEEqZalw9DWkVsM/upWySqT6dBX48Kt6WNIHh+3VNys76HwrBaD5
5hYcajKfpxRM8pCd/rOGOiIiAt5nzYG+U7/H2s6xgtJ/Xf/KWkIaa1crESNwVuc4
sPF0j5kYw5HTmwOfcdiOApuVdVaw9AfTZbOAtlyKHZuFQNyHyGm9tmGqQCHU/Pyq
H6McPyEk2FX/zDRuN+kx+d76FSLvHp4epaz9IGChlsW2Xxs57kZEHDQOUzW2ckqj
YUD3Ua0t9d8r93MFtpZ2ksqFIWU+R48TJvfGL2+DvLMlQj9vYdpxEWgGHCXqSEFi
TQPUyaSW5pV7prTDaKJofks7E+JmEtptf6RKj11qd7u0DeZ0rNs3pJYJp7DDnkI6
PW0vX/BNTFqZq4F9400PdCd1XD1AYS/MYP/na9ztLyAs/8pbdKIDaFDkASHeDcA8
7bHJQyrMs/k7JYLmJTramBkSrUgDBugiGQ49/jJhh95N49wvEV3rsXrDwH3PuBp3
DU8yvNy13LvIUhwfak2BZIg/UlJte5dUiFhZD8llpijcDGBKhi7K0J904WKPI1s/
zGT/cFJmGKJpQc1vOFCKv6AdQ1HD+jcpwH+weQ6UKWFeWtqiE+358RRf1+Ra3/+t
2seE2civ11N4F/zCsTSAPL1Igk4tQUHGQ+2Qi0r5f76o+cYysC8aUK5PvkSF/cR7
3F0qmPngTIO409Oyzs+QGblM8B1+fXElOoyQf/vQnCuBONWz+N14ajBJC/bk7Z4s
PQwNVxQtNRO8KcbCXs2CfZrPqYAIvCpFPvQfe7DLpAVcYQJMbriBFHhb1TgUu1+6
0ioD0LkxS6V4a3Zg6aYhoL+bH3hDikubOk8NsDyZLlQ3OJ0nIo4kRhYbXVaLAy9I
1cpLxyq76lbcWRAXaqeXe24LSVBxj8kliHM1dHBDBPwHuPeiggZgN07bHggP6gAw
SvD+hcm1IoSVRSG0SHkWPYjflgnxIfb+ZlVZ7FjPrT4CE9WkgH2NHQV9utQvOdXf
ezyK9dBXVFltjbFCjADSbMA1lbajsp102I7tcGEeCjDNTPYoq3IlZ7N4SVCL+A+H
9a925WH7JdxFsSz9X70++/uH64JRZ4DyN3CdfZSbHC1SlLm6mSj3mslAeJjXDpIE
If+PP1jvC79Gm/x3BluN7JHnMVFOKbcOBC9LFK0nGH6mG1SLiGXuA5qVfXei8TP4
FfWyXgmvqO1eddHkm2y4q56W6REmkdD0KAScMT1Ro+ruHijgQYsYC0DvvU86YwZH
cVh4G435MvKIKoRGL7QyCVv8KbW2hL4kdYO3L5/Mlip9LLPgFMln1yCUqSRtXwSY
Da/gmiH1FPhTCMaMDHHLzOIpOMMQIH6OfLnkMkojKec8+4g4QRlUGD7UnhPd6Sj9
bAypAmaSndI27tuLSc7rH/1yrrKesWJyit5cTJuyX91Ph3hVwPeTM7zLiFMc/2Aq
dpQrMueZWLvwxID5Fnwzzi7+QMN92yWZ+IyIp2WxfV0mYMxipZydLsS4jrThUoJU
N4+X0GVItYN10gxyjoPWsjrzeuGlarkcWXryH5IIuK00VPEzwLzH9UScpn+HeEIi
TlpzLdJsTko4u4YyBuVLqJeAlWOvItxQGSpNVIL3pLRz4DfH8Qyf2eYbJ4yV2zdB
tXvLFTq4oPsbiHYhKy2Ov9emc3Now2BHQbcLnoTs9tFb4Zrs6FyzJjXYXECH8F2E
UHkifPqaFpS1WoRLmlDTG6QKPFwKXWjsyGr0g1Rj6SbQtdS7foe5ugm5iM2ozop9
EdCXDEXSMfX2EIhLosDQL3iDz9B2Nn86Cfp+f7plIj2sbvUvcZQlwCGXNBRtzhfq
4XGQg8CxMv8lDhsgl3hoSSRmEZ/vfamrW1gxUZy3qNwUckkpYDSGFyAYiExXeqAw
oEGcLKGmuP2N55Uu5v9wUx2pSbH9C/dHxh8nUlRQjppAt7cdU/9TMYVXgQTg0YBa
Wa8W/VzXLNWPIo6RGZ1BMLyDimxjEnlBJoYTnjsxb/c=
`protect END_PROTECTED
