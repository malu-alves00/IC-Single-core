`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fPWyOoPq/IVerkIkAtcUHdrfwHhGSTAwaedTCHOb23oipuTTMrDg6+mOVoBFeDmC
z2IUv4lLEeAf7X+s8KC66NjAtJKnFYeel7LWrz4FRKHfFCcAOme/b/0bp3wQJcrH
Lm7QHILu6olFko5m6u9SXnG8yenvdEE/shHZiOyTsCibOjuN5jLHQgPYlFGTbL1Q
Rho3MfK+/gobjaG/2HB5/cLNtZxU5ENShOPzk8bz+CPzcuvU8/sZ0vuT5CYWZubq
89Xv9Z17UH9lOYpMETedRmPcCV/wiQl/SLv0RHMiNNgNmH/8I6x+8IV5itcaGa45
z+UuDLwkKjhb6gUxFqFCYT5FKq56MfMqoO0Ielrq4dGfYOlsailpa30nInGQyoOb
JLPY+OE1qxG8jTrWqIu511F5rL22d5/sBDuLJPGI787K2ELiTm7zjegf6nNMjEyS
/dO4sgiqDhhnQ49cRAvT0zvCUpnHdrdh977fhJyDmOITaxT0Ir0RAVQaeU/h9Nmn
e73isMl/mTv7B9+OKPAsfeZfrY9mRHiUE84+PoL4Lqbl8v3GgM05ESS8y6xSgKnl
jYGAOzlMFEE+91bVfRgml/PuVo3NuCzBxGnA4lvDDypuLKTJ54Jw6z7iD5Yz2Wz3
FLGGheJH2/mIcRx3Cpu2i3Bho4pWcEE0+lWJhgYNazn1JyscyvbFuzTTAFTRMToe
OI7Y+hT0aFaxLREUS2tvWvyRHcQmSfwWWPlK2XOetoqcvmIALINx9EkPpep+qOXh
XtC1d5ZL4BTtJVFGKNiuilwIZfT4jxgruGrsado0V56TLiGVNMb+oaN29nLj2QL3
7+JE06r2HL6L5En0eFvcvyLeRaoqJhbbQGb71dpDGSnwa/fVexIdJMm6NSyEmPQ1
PNqYxOh2183MFXHc/6FyBU2P9i/Menixxc7JomDoeRYTCOYPu7OpvQx+cayCeGoD
e+1Wks19On3Xph5pvxrkSAKzYOFtC3CjdBCyhKGa9+TfEx6M5WyqTEu34Ih+3BfA
42NJdNf4ke8Z1geXOjE9hge4Xzi/sT82mYMVdSI6KVvQrpXEivst4I1p3W3z52hX
oqENJQ3gJnO5tGzSsLav3eTAgYe2cXgs3TjiGuOfl/FkDNHRjD7v0pPSNnkdkKV1
Rw6y+baAttTuaSVTWe6G/cHgr3U2GzMhZD16CQZpdftD/H6y40M4MjEihNoXFxBE
YlpJ8d8z1OPNx+ONu4/Ow2Loiyl0PO7DH+Wwca5ZQpI9xwhwRbGrBt7/EPo2MWVL
0JlfwWYGAlkviRQ33hGz68yCMY9P5q9zPrvkhHpuKvzyEuOTtL494pqWB76ke8wn
jTljk8wQ0I5ofaEM1sixfZWvhqUzEZlIuRlE+rQEvCXUIb5e3zmTmZh/4Iga0chM
2E13lDWhPIcD5koj+0mjxQ3JMTPQC3yW3sjOstgjXYUoM3jamGg9UyDnbONe+dKX
NbxSgfFPesQa0ccZMCSlq2XKuIXDzD1JF40BEtg0lPauBJdAcXI7JRQSd1DpGw9r
+7eR2JGCAf5HEmbIJKySkkrl6bd/znwhlcEEr708nuSM5hoI2ye4PfSIcyg37KOl
n/hWjfWaIPGL0Ylo/6lBcTYvOyaBLFU8wXFkDg7SMoM7guJKFgke7Cw/Gz0sYf2D
CFl4pKOrBxChlCEJHR8yX4IhM9bbKoYyxbfebXkMgi8G5wGrgGZXpKH1Uu0sBBmK
bH8EpyHCpETQuv0Y2zRjI7BOMBGfwZLLHkcNCpPEHvy3KgKX+HxvdDi7TqyVucSs
kMdlyLkI4gRlXVPjt5ZMua8VK7yojdpJrhW0B4URD2K2YhmwacchqtxphT5lSCO6
ejGyqMol58sJz45txjUlJHQIEADVEjOws2UmWpsQ+AfPijjWlC6A4U219BqOe0Mi
pPbU7wiEjCmdlP72EwqlQiz+d6oCyyPSw+Xb+ywr0q6fOtWTwkL/reRvoa4RqU02
FzITYzIYIQWSx6Iw1qN55NkNlFmi7vnl1Mttf5InENylG6F5gx5DeJLICFFnIPXQ
rWCntYoSh8wd3fF5kKp7M3FC4UxY46TCwg4sNkKraBumiPtC7JvjueUN2pJP/fh8
zLXRVN3kmAz29b+ymdKGdg7/3i8NlujGRaMc9Es0SBVpf5mjRJRKv0UGe0hNp77n
JwVEvrAz1Lw/tuq0qEWk+FswM9n8UQzGQE54jsr+wRBgCSmqMNqzDkOEp+FPSkf/
TDItJss75NyLlzdltW/uNzwAeR+NsoPjovz1BXSFrAgLhUJpnUcjwEyXiNc3UyEh
7DXiiBlKpBAU4rZdJFkoeHkZeXPeWBzFpQC/W38SzS0lDCdAxbGTp0KJNI2Kzhiv
fVVa0v00nxiKpC8jOMEm+P91pSbyzIky6pKjdwndxaTS8dQi7sGUL1D7LiUXLm0l
f/qGKMVYn2HF75IzW5yYC4o67OwUAFlU1PQ8BAYctK1y+RC8bEIPD/5MOUHVyjOX
yVsKevqAW8jQm+SIqKaouKYqhX+2HJr0apAlG4yfSJdXS72WJDfkWOp7BA+PRfud
Cyun6/YJ3x/zQFKVgBFjeRzKTgBxoTWuQYex3rjoG7Wd8JJGvGn2dRfoW4RrFSPA
utaDkecZ3Tpoqh3GBym1CvA9uLaQGc18EitLGY/bpN2Y2GXwbz0KvXIUhmcfKTm3
s9BBKvX/mbVl4pJgSui/YeV6y7mhtNRejij8NKnQFMgq9M9Q22CWZmC074NkwEYF
wNdGfHRtXIw+CzEnw5WhgKIbEKL/P8agRw8sUcUKKhxSKMsEpCYTsXG4b/MTPa8Q
qomLCZh18lX0RSQaKBnY8EoNnokRc9KFHY6FoTIuV4AEjAphJsDJaU9mELKhyaUE
++TYLc/cuD/XOyY44PwINUx2Er76TfO4SZbN0XSsUcKg9jKtZ0SZ/8VTZW6yDAn5
YxKZpahV4wgmVybINLQ6LeRs9bSfkAlIsZrqDwQDxpOEd1L/oyu+EEVfoVAtilRK
+A+RbV7RM7Bc6Gu4uPZ94/ygxvDzVqmB695TzeNvRLM1Ux3cvcKyM1nFaDlQVIPL
P+QczobzjLHk6gL2/9oGrFpNPAp4ngAD2G11azEc2Xm7d+KeS9jxKHHtJyoou+7/
87h2Q0EdVm3ej0NvdV43GnDrs1dvZGWXB1H1JkOj77ESvF304xKzfRDHdFleg+wn
0kNChaSXDooLbJHqAOFXp7MaWzrfji6Tiqv7RHzb3ip/sCZ0hcNJ9oA+dNhgV1CT
7QlNA6q5XkZJpthkZlZE3iKvOLGMB13HzGe5Pg6RgoHH6WqZHTWRAGmnRCwSJlX4
8txE5UMwsx2orhXajK3CtqSSV3w9uaLI6FgF1ZO17nXcLxdwgdjNzoVSwjRkG/S9
jtQIn9FwDUE8DNFO+Umk1uckSUGSUzJPOoyU50TO3ZxkHbDBg9GD7fHYb7Dugd4D
QEGJs03UwGmYPCWI+QAUl4LXyCOo2zfpuKkGHv4kQH2Zy6Wa5+rQGRyUvFv48VR/
rxjnKowpAUj+NXMnOTvYuY10kN6GL8qLwtW9f60LQrxhtpWcp1eaFSz8rcH8/uTR
q1a+LB2rvEE5rHqP92Mhqj/pveYixqHCtN+/8d7Ww960uZV7DPjPpKyexe33IhoI
fKeLrZqATX2BX8w37bdrziVUY804ovgr1kkta6sFHUp5zvANXF/BO733cb1SoQIh
0nTt+6o/PSLyh5c1kMAc2aPRUfB7Vp2kjj2pXGf4h3rn63nDfKWtLvj34kyA3PZV
aTJhMGjxi6/QtKvVWQqgEE/PKlhD1OCQo5i3giXy0xrRYTMbvReXCUtK/r3XPJgv
Jvy+oSHiM12XfwSVm0IrNzZ1S2uSPGuRdqJeTuzYv6J5q0IB/UVw+x2pXjiPQYS8
mXY93MdmRbfDkctmk4IPe2TONKUF/OfkQvciUVG5SnyHny5WqtRg7ivtg612108O
sPZ5rCing4JgcXSW+C+xm1BMoX9XuafuqNpzcU+OZvzQCG8jDJ0XWB0nMESJtc88
sFI1n9+04C7mgglQSATOev+0e+7MmzKeFbZHv1ffx5VI48a9QPcGYNFilplFSmvp
clsBGUeNwVPLWcnKpiWfUz+d6DOV2po5UthPoqckxELYzimOXnOea6uk8JMljEx1
nB16tKEa+mb6IvvOKB1MN6MUx2DOnLv3SPtn4r0uCHe79MONRwJVWyIi3LJ2eH1Q
ldXAZOel3KSFk3aLuw61j06Z5rnFi23YjqGTBCRmfPL1F9j69xtAOFBpw/ggpLG0
oNCKRkKHmrSYJfAiTalZcBUPs8nHNbQjXSKPQzxnHGr9vG/mza+vhCGZeSNWQfFM
GCKbk79OLqCwpAZ37CVH/D3uMLPS2brFMDL4ZRFe0+kP7bo77n9esnyJHCFoYUP9
viS5r/k55IN7eqDm4JGsJmKdlVxLpkgGY4mlGTUKfjtfm7axOz4Tr9noCkxJBQou
cdVuuILyh518/viLvrl2IK7lNcXtiJNDFObjgWJzgSzJsma0Aj41x1X+sN4KAETU
aTHNJFsQC/Kx2Z63zh7Vhi58igEK2B26rXDkJT2pmZ2Qcow4LSgM4Rt4aXGZ2UFD
`protect END_PROTECTED
