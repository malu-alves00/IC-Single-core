`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
i40PSAWvK0zbzUUkGYNszG2GfpqYAk0PSzGC3+OM5y48LL+ek0oTkL7aEcYM52bV
VRZLr1LTosR+hHlr/okXlgN5PnJuirgBIht9bFISzJuZhpKPet6nvDFbdhg63SHY
rdIlF8MrRLcGdDaVNgUtvlr4vzhgvltUZ48F4VQHzPbYl4jTsyrxts0zy1R6qM+U
b6xt3Pd/0GHB1XY55Ic7dTPmjuMmGqkq39grO2/YJFVetfIR6nq/DgU3W1733BD3
I0iQlrKI54GEpSj+0HnWMR0YKNwvlfz2WcGqjXJh8zoAOWFoHF5e2TTUrQZ1OV2e
yl5z4v8cLYVks5qqXZCWHA1FgBvuRcVXzmQnyTyWTUDqOUcwCl/zDni0KAYS3bgj
oKJZ9UbORcI/4oeNXPQqQw5ElWe7TMMvxySD6jSRWvEymdva6IOcn5wbWvSt+50H
oPh2Vr4R4PrcrE1UX+wpsO4TuXLvrjgp+SzCTQMiqw0=
`protect END_PROTECTED
