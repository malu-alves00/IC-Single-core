library verilog;
use verilog.vl_types.all;
entity tb_gekkonidae is
end tb_gekkonidae;
