`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BAbJ2s66VhpByNWYac732V/dGe5Vt+/6atel9/0dXseu8zLJvOkBw1CAn5aj+KAJ
vkFEg1ZNJWivdBrAGjo8CUVgp2HAO9Fz0GYMGDidKxpQtRDS22YXOUMkv8E+gOLz
Z63WujJrXkEs3fjONUMluifG87xIj4toNWmS738hhPCDwU7nTS4MH7BrxrWuniCC
XtRa4MSWUcTQBc653aQylNnBtS0dyc8qRLHNC7t9iw+Vl8O6uiBl4AKd1kirIqXW
1HEBYNsVa196NYJYJ3qRejCBdTKbGnG0UV1gGZIF/D3fYphjdwuzGMDqvkoxJ9kr
0hXm6Pp2LfFeoRuGjntcHs6D9W7QUuA/bwWLFcYBHOyYxWfBhOs8U1tXPpAWextR
FESvz7uqRcnCPhVz6tlQokDj/kYx0u3H72IrBeDlvFevkxpAfQuVQB6nOtQrV1dv
ObzASbYfE3hb2qzD+C8ticxll8meFWPffi3Qf2ogriCtL36pvnfYpqTd1ldTbeZT
1kuAZEjZeZSvuRb/lUcS3DLUm5xNWP68TSi9cVrbgkp294hPAgVI8wl5t6uDAt1X
Ia3NY4TnCjnqirVPAeDNeEeyokREWDi3WCWR+GsHR2omU77+5jYLZZSJH22B+AR7
xx9GgUxFAGb++gnWbIC92f7KCaF5+2epC/zEZkWdpuewcjkhxwCBfSIsTtpbHZYD
AxJZYyF0tpwOkG3nN4n/sR6YclgGJarRaDsxdc+cT3cWUrfHy3Ati1gI2+gS4TvK
+EqDk3UdrfyomnBnxx2pe+yNoK5XuKdUTI7rK/0b8cKcYcLqB7Ig5GSZ6oA5lqKq
fLtL5WYx+rwsa9eeLdUsaZr9YYIPZCFRzvqWZyYeOGEDURcwOfTvGUn3wgb+lfJi
/0ZZ/PSSp2qLxMtm35AZ+O73Ygau5qp5J9naakFI+OU=
`protect END_PROTECTED
