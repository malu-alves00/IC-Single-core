`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WIe/lhOZ5WeMc10uYpa1WxXF/+eS91nHJI+pBVGt6/fhSPbCAyylty4jIsnngxfZ
jksHXsymorhOnJVGK0nzNGVbeiQlf9WOXzG7boXv40M18mP3z3j51SCxfZZS5jvT
uoRsh2oSMX4CWN4p76MAgmBcr9+7CItHOmy1fSLidza74Okr5lgGoW4shiye4SMK
+Hnfv+Onl3rzv7a9fQrByR3jIdBib3zawZYuALwosiUn3rzxohLB1Xkcsu0kywXU
yhFf2EH+H+0feWNxivzkwx5yeAm6AMDEBWh3VGGxagrT8C8E2UYCVxdrIyRP1k+v
cheSCbJytuD/ekXzgqSobRyiI1OLZz/3N8pSlec8jJ6+P0LogUUjE0ZLwzP+A6fG
0YTuOR6nSpobSaeG6/pdsu5+IA19B2GM3z4QJPK8WeZzoNcHV4LLtftLWQ2/7X2S
ZBlUC7CkTxZCleqOFmrYGbw+bIPqLoLV2GC80maQgBqgbpEMercJmgZrGUsz6Fv+
B2q4UtxnDR4mLuKPXGFqfQojOZYxKtgzP73XsBKPAKWkZyp5EhYTsEw/fl0nJLqz
DTsgjyvC/OOmdeLrZT383YH3mJDoEI/VP1iZYdFJJeQZATn5pYUzhWGLF4InixAW
gjUd9JxK+ZsHHLoOej/7gp2CVZMLdib+G3smDcr7Fw5vHJGuqviyD1sE9NSBjkQK
rfYPtN8FKKyCdKnw0z4cuD2w2zckDTvXjxrfBeIoebdHZQTkb25m0jWKJoJw5Jcf
DE1ZqM/9EQxaeWiGAtJWUQPnaEXsqrOUqqnVCxAVLq76vBohTcsmkKwTsq4dxfoS
`protect END_PROTECTED
