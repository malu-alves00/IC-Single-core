`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
K9ytMZk21ayMk0L9fMJcanQbQco9Ab+Rj2tM5mZZUrZYMrBojUJQiGARaFwbP3I9
BGzWnQioxH9Ic9tek881RKrd0kw+HYxFdYEiaf9rF0TpdEL9emxuT2Cmzd4T+wbT
cJVLU/gBV+kM+IEm4IfQt038O4RS7pspm6Y53JTgfZfibasoVeFDm9CXUjvecRQk
Wkt9EpB1WsrRKgECvG41Nol5JHbhy4ujGMCIv1bD7y4/tHOMlQlraT8iRmXzj6Vw
11ZPZ1TGvwj2S2BlTqVpcTXP17E9iIOP4PNC2r3biGt25H3+MeK00VHoSP1eChaK
EsX40JVGwaCNnQ9ODyQK0yQpMHfldQXqBE/FASMeaYJhsKiSPDRBRf7vsaeMCZpw
sscL8Y3KR9Fm5BB94ESuGn664a/ka54Lj+Z2PkioKKRoLOdPgDzAl9jFckM4YbQF
PYFATelLkt1CgSaB4fPdE05t+SWicFMrNvQ9DXQBSGs4pRjzIjSQLvL/iXVLIlyF
1HTrahCwaVXBD/eqr6dOC54gTIsP1qzFz1w/Zi5iHPP5qjJFQyKHe4CfJBN8WLPe
kD6GMC69R0W3wRUj0Hi/k4W2cSdhN3ZIvI2FLtS6gUnmHmlYm937CodIfRYiDKu6
SeVlcBN08B5GEBL5yD8OSTizmM9CLfJR/a2UPiKHGSrTcIwTLx/mDOqapKF+kvvG
c9psp+H+6oss2p7F1/YP0uZnL9OAsWAloc+blAOqiWKHjm1JCQRXSUjAP2y4LZsu
3oA7W7KvcH1LTKH1ZtpiLn7ODL8mw+mwC0Fao+y357z5O3Qe99jY3N28HM7yP3iI
gzl3xH0YdqQrDi3DvvXTyw==
`protect END_PROTECTED
