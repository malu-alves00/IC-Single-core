`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
y5HCScrNKiJOY8mJ6QL0YgoJisf4vVZPKfKT0eYdF48dQEIqpAx9ToregoQsDPUk
Dqu8Yx5df3dxX4/4ZlIG32YXJQOn1pI/iuvNxJ3Eh+5XoVj6yN1kIeU1y7yk7T8z
xIglkAMvPCb+zAYKV3b9ugk2KbtNqn1/QcFwQtXa9auoCUZJ4EGmCCj9gEJgT6Lt
G+x7OToOeKOnAHt0lyabvp1rv4NLOJRdaZs0nXhGVinHoVy/yt6kyX7AjDmRV2/P
4b76sKTtuaFbXfrlWl6ccozETBhekHSB15AiRxGDOYTyq5LoON9TnLYbfF3qZsld
Hh5TGRbuEIApucIoLYVSEZn7YzMlyFwnB34+sUuQ5wYLJe5vyf05McVDDKiH0U96
5T4WW6kZCmDjmtceugnhtPpg0MLX9UGSWTAZYhS4g6f1/UDGNGWFn3BCvG8aFGMA
aia8jL3cG7KASxRivK+sXJKbSVRrcd6wJNrjUGiKJaVqG0RHBp++GxtGMOcJ1C6h
32GZOboilYZOX35PojMzfyQuuFQaP9dl3Zap21Lxysmc5ag07ItsMCiWvYLtSo9E
yDEmGrrQEpdYIS3YO73VNCTygcvKsPUB8KjA5B5lFg6AuZeTHfMNEjhkiGWyKNQF
WCVY3CM2Ltrj2XfxrzfvB+ryfhmde0vB4dpxnzAKueg/5Xf9lw1TmKHKMbeRnuR8
4UdEcZ3Q2k1tzQjAi0H9OTOontHECYcZ+C1yOKQEcM/DGfaC4yxyZjX0UdWJ6I4O
/+NiDKk9rpAPiVsPdRpNfyS05oFOiDXlkx3h7kX9jielW+hwQdxDEyOVwfophtZ0
NXvGXn+QbEBUWgt0R2CjEGveK8Idy5rMsvbiucNyjC6U/yzNq+D7//8SFQZp7/lg
Sz43vGdwipJYZeXsmEHCbERObFi20BZTP0hLt3aFW7OM4UelJL71Opa8N+bp8xt+
13tJO6hzWV1eMXyN/XA0ta1C36XzPgcRl8MuD5tTr9cqztDZJmlgCoLce3T35UCi
BaVS2aPOHOa0JELwRhBd/ljd9KjYgnGE8oIribo2qhHqcCq9ujh+vk0RaT5WjDcV
78YfifE4HO3eXmnyQb3+TDrR5UEdml7PunJa7C4Ss/g2VqJ51k4I67ZmTKR2uNwS
aUKHq9WUydItBzpTbVcFc+KRnJsTvrk2kFba4R8OveNsQQsXZI33EH8QJTmCq/kz
wxH6YHMxL1XX0BBEkKi880FyQ/nwt3FQK/TVQwT3Krck9RYUt6Zt7/7spz6v7dT4
J45+DdiZTk3YCfCI7k/kEHUzAqT4acxiwL8anE+2KYoZ8gIZoUaVeiRGKhlzzrAa
T4GRvOrJRg+fP/QMh74qqR1H4OagcRvnDtZCsrryEwOT4hHMYvBpMj/7O62KGEvS
9zYZsRqNECzGplQCl0qm3CQ/KL/gNVDyx64gZBd+rTFrUIm4EgbxZug9hHBBMxXB
Q6QTLIi0S0q1+HQy+0bavTX6N12Hu5wKlEqgTrXVQy+FA7PLEy5h/fK1BjUUbiuK
3meNGXxh989ZW/ReDk258Y/VY8lpKfSZIVzeMovVmqGHkdW64Xq2OWQTpv01HDoh
Sn0sXnGTQQTazN9275iDDodarb3BF3cEGWQ84MEvOzL6ylQNCNefRT5Ivm3lkL3w
zrbdlOL5qR6hYMUSSg3vaKZxGguPGCsptfLXCNnnpiFB6x0Nyf4JDW2RRgCuQSDM
ytI46JCs1wh9FakbIF1KkeEz5NPjTQ9TofUDJA2u95BQCx03s3oh7+n+ofK4kRHd
CN3wT5EhWIvlEZsYxDv5HNjgcV2zZiGK+gSMH2RcxDJ8Aj5FH3cQnHO6Ko6rCCMv
4IRf9/MM0hVHLUrW4wC9KEOWZ49M9NwSPaqpNLbLfgQRNK6ZXBpy+d2onBmUOxFz
TRu6iWHFxzz1dYiCKoPxl/swTIvR3iMMBjOP54jhuKA=
`protect END_PROTECTED
