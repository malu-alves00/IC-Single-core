`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LxJLUGPZ2JU8GDj8z+ciqP8H66nAUnB0ICTHrfzlU8+Cc2zRogSr87lpoz3Wdrzp
NkRAI0bTam9isavoY3/O8cnxJAqPzywCru3NUrtwm1Vj7f98zBnivUnZtu0Q+YtK
SRQO1B98yprLU1Yj1kR0kENBAlpkr9dyXK65H27IkjbnsYEziwtiRHJml/9BAbgL
gRmO2+/NIq/uh6EL2QKB54fihmhzItd/q6Y+mTGw7LFy4Dcgxppo9f9pHijOe/IY
T1eiNmo/EFkOQjXZ4gmtNfKMeP4J73VDf14irXGDpbzEu+wwRry/my3R34lowR45
gbrdtv1H8WASuB0BnDQc5RKPePucSPa0hSZQRGlO6ZIV9muGxLNg57hCvVJRNm5n
PvmCG0x+E64jGCSacQxIwPHKEl7s0eVhfyinBXItqaNaldRk4ogJsd7eTekTSBg+
rxI5yIBKb6mSXcwZx0jtLhPDbHwnMOpUA3QtY9vbXZjMe9PR64MKjh45I359QipI
XfNiTNvFvtx2tIJrcbqJz2tTbC7nCe/Eskv3BifmgBtBoNi3x+Ekus1Gegl+gcKx
`protect END_PROTECTED
