`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lkB+99brC09gyznE7JUeRGFYUntMffpMduLPkVMQ/wwzTgHk3c3Q5/quSfBW+aQ1
P1v6sBrKtRxVe9vuclT+hxy+qe3FQaUxWJUNz5X3idPjB9juHI2jdtGBtVjn4imv
FW18rLjNXEPNoYgovht6u0b1Y1UEztT1tpRd04hP52v4C2RpkqcJMT6amMX9SEpw
Ka36KHR3y4R1UbPFbj97yWgV5kxX/h+x+WOMRRNk6YZNDSGcjq5HqejCpjdFvM9V
Co35rI2ZpYDGKY8D+GTodpgKHWSFRyIQKa8M8Y2EbGNYSQlPM1NUJJHqpNF4lAP/
kqoUHCYP0eymKDzbeCDzTAywO5StBRTTSgvhT5gaaqun/bLiCJ+ArIbaOXDiz/ma
2f20CCjQrTPw5Ru4FKaZHnYFO1dZj4xul9M/+jwXqBoqIh2Col5hZepd8ZHvnLik
eZ15jRFZ7p4qIfrpGPWz/rA+Gcj+/97blheFUOAiM6YW40Qx1miRhnp+Fn4Qcv1/
xV9vJXDOkRNjkg3GqmNVeXdJhjhuwI1PYVZXJ1EbTHF7Nv6dB5xIkXDFBFhALdrY
9fdOo9eViA/d1ofJmZXY4mCCp3k/kPF4ebFVP2bDBbxV8IIK8pyZsAOAlMIf+DWc
CdE9lJ0Kjh9amXQH1i8FAUMEquEfPws8CIkn/waQTSs6tZD8tVNDCLjSU4AzQ1is
ExhfTW+QRSlpFWs6Ix2lPy4OM1sxESGwOZv+TEUD/DHrtQnWbzbnJE51LUDltqOB
nEuPI7N7HSKOugV5xka+SPqAZfqVKZV7qnwnw4UGYwPKPi9T7Kyfm39yhhGuP719
4oL+sjnIR3KetqHre0762qTjOIt6tPobxXHxs4S9yvR9N9aIoedFm2YcB9czmyoc
V6ZwQvOZVG+6zgg2W24o5K0mLuCSKMUdscPfqIZR89hGFJNG+h1pK+Qw54jWDnf8
EldWTmDkEhvPeJl2uZAG761R/AwBA7c730VZlUGwtPenUNWXGHbT9nHv9bQzHcTo
fQLdZVVY5F2z+1w1rhMBeTJTxGMkwSZ4GPFV3DcmV0abzDnJvsuBDanEU8Bl/gSX
SXiKEm2Fd2oxEhV7HvGUppHkvTg064mmBVeM0uaeIn24Wl4UyfUpEZOgQ+QtrvxN
Q+pBgNLktcHYpeGwYu6G0xRKixNEU8Y+rzI+32EtOVbP5sKWITWwSmhM/1OjuQV6
bXUHJHZSRhr/xUAHn/wytrlhtYxN7im+9czWOoAoXrwz6V9Hv5d1mvmH7XgLF9ZF
/DY0SOLgG0eFWTIMgZvqC+UGFNGwSEKR9YPKNWNkOdabp1JvABW7A75PSzJxCXpw
6+0Fx1V2NWQALhdxqoGsHRBIgl8hVJOPj71q61licP8nA8npZ+2TmqYrzkgnYLvt
PkK0HLIEl/ouTRzYa/fzdXDd8I8x8uSsEZvmhXcsiEnr6JoImrUGeMaDRjl5UBC1
hGOSiM1nXfmSefTQeMn+7JwX9Wmnq663j6WvFl2YMzgESKu2WVcEiMNRr2HSc7L4
Tlidbqr7NacEaOmINt8MoN+y0HqpnXCtHGGyRcjukfncKPReFQWFLAp6EnUNyrQS
HINeGkBkW0QbVO6cqoAXEHFKK9Clc1bGiEtXDNLeYi3YXoN21hIL3K6HMazET3/O
2jpbJIGFm+fM6fNTJLBKYvP16CG2CL1Mr13ecqfQu4qMGHN2dXx1pFg2n/gHmQsx
UHVe7zRjVe3xXTb9VDXJwtdpbaIxCIjBODUykf439ckWA+vJJXrlM5HoYIXVU9Fp
L2HOBFKyQ9XZtoDHpJWnV0M+5cejfevyPn9c+QdjO+kny9NehKhoYDRyZKFZq3wd
XHV+2H+aIs33jxvRjM6j9pveUYjAM/7n930SGxwM1MA+INP6CbMuVCZmYzwNtAC4
zFvAXUWR4C97oYmGDdeXYobGCZxwjAP8LqjIJzi6Xv4peEB1ctFZOD+rSAK9fswh
Ql0Qx+qhZx8EArDzaR8UwhNYkbDmS7tWDBlbPPb4xt/k82OWiDUE4FiJx/mRl+oh
/rv4pdEnJF4WNkgjupq6NteNR6C8EZXD6w4Uyj4WULcj6VryxcY/7uEZ9zgrfYy8
yn6eTjaPHLTP4aMIbGPxcR/tUrmoS/yh4iGki5UZtawUCAERC3ppd54e5nfJcSZm
oNHGAaT6Kh+xoXnyTpZJ4uqkS4C3Ime5z3YciaWfje7IDjniSVYomTqD89uC+3uo
2vPuDM/U06pBIvVZi4uDDLILqfyqfc9sJ7JeSFdFLQeYWH0hjCA41xrreyq3JyY/
kQPeRmUCnMYug8+O2WfaFqvHb3ejTeVY+o+oGxW84bc8JgJeJ/UzD5L5X3bSLqzL
t62aRjcYCmos1Fa7ZmOeDup8qxy42CvWJ+VTWTwDWeQ2VPtUk/p5lQbsw2rBMauX
Yx5DqBcLBLDQRPIE2RRSj51Szu2iXFyoLpltHsnxFNRByOcbseRz7I829iYMudca
yQ43YZVG6dGas+yr0d3ickRUOMBwP166x8rwzKiy11V0DNf+f1/jmguoLB1OhI9I
uWedChu38c/abiDU61lVC9sJNQnNVBmT5EogAfCOpHXm/qr274/N5afB5OBDCoKT
VXCAxGH9YbLxmCIz7aNL9yMBbetLoHxJHcZ9O52rOrp/uCeHx6Gz04GQaNLfWgm9
LEbf5RFKSouXbMiO/KRgbl6610uXINypMQXCEBJ6Gp7SLJCUIwGySLXCL8qSM37Z
aZrGvZDZBklvfiwxRe8otAEJ0xhb+MrNr81HYTFRCwOJr12C7NyeZBm68TQQ+euP
sWJrdOx/TTHyibAGdPzJoZz3/N4v8SRgcwGS89x+2j+L3+7qMvbaciyuRi+VyCiz
zCrpi4TSRRcEpECO+iW/u0oC6F8Jg3w/AuIULvBj1DUNiP985Qu/75iHsUA4BicF
bdmJQ9WIjSqHxllAuGpWg6K7uHFWzmgVvV5Y65WceaxacUvwPSOGl2noLK3K9uj8
HGrlQ6VZXzNDT8z4yHMA11UXt0Knr6vFv+ioCSCZQWOrpTxrrdDiFcHOdlP0zUV4
xthilSBjJeJLwMWY0ichMbthGm5VcaWB2cQYvhwm3k0mqqjPR3QXIEwqBpy4h3T/
JW8ah3BndKKEPJXGNNWn/0zZrhH77iG+TDL8H6crVzRtizZ6W0PK86h7BsgFg8KK
D2li4G4+JS4pltjyNyr4WzTnVBAtM5AzRPIMuC2Zb0KLY6FKQTjmzo/TnY5L9hfI
++07ldbkkdE5PfKYHhJMOBAFm0d1Bs8kAWk4zkvR3yUNQJ7IWqmE/XiSFdSu41nB
`protect END_PROTECTED
