`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZfYdujjvmJlHcUeKdJu35c6raGV/UflQcY2KUBsn2RwtvF2ITV+CKJO2g/wNcWsI
zrSjAvDFRNPLDmoTSb2dIVxaEGphiVVAFak5H8FOOsXBBOuxBQEOhBZ6FM/M4D86
b9nt8Z3L4uQWR6/C1BKlcv+deI7RBHE6Da4jw/WxlHS+K7s73HPsG1KyYY0oJPDN
RQwE0BiXOJcf7Q7nLidPOt6uSIMMyxngxJoVICJ/YNAfCLZK+66PLbtM51XkCCC2
UOcwdlU+Ax55YG5fB4y4+LokhkhGh9IONim+d+wZy4JfqzkpkJPpwRiwZSXwONKa
5FhGVb07l58R8hrZA4O8OMWfJjHguwafbkb2PdBArwF9xk4X8pPBI0nxPyGMaSZl
+8xuFDZgfE+6RSNEA9qpzhzxpH5J0yd2qDUjmTHC4J235ekRjY4/jBL8ZymYzzB/
+OI5i8NH/lduW3S1Fb1ORBljI9APvHyhhz1NWjeXQ53Qg7yDjHP/ad0AsG1/ng4O
7GLKPIICYVgTwsaYJlEKi3/3QiM8IpOq9HtZEl3vcIgBGINlFwG3/JR1MHuo0+Cg
o5shwee50w2CXQAp+gTNgziQyOqL5b0PNDfQuaQZZSeejNJDzwpeoBHh7JSObrBM
ED+OT7hRt2MyiHAMEwnuOoKgT1TnNy5XDng8qQaU6Gpg+E+1tKEDW4rREBMjvZKt
F0F7Lui9JYGcGhFsAuNKku9+H5CTTrU+BGJozORpQD8=
`protect END_PROTECTED
