`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LH0Jj2xPXUaByZFcrgpp4m6UttKqos8YCgQF3GuDHPAMbV5iH1tVrcglic4UQcHX
6tl1cV3Z+3QdRVsrF3iGjsLBhpmGi8EAjNN+E50JF01XnZQFyCbC7hgKpf1xiDWm
7fGC53OCJIyQMNWMjbo/+thVp20K9jy6D9gTNf9S3y6ZdwgJ5hpxipONaGH4xoWh
4dOhSRWl27wwiag/KJeq/RwZubswzUGQvBbqYeyGtveOPbDW3YIlI0NhkHGw/LEl
C8DvUQG010ve/4MEr6kFpU6/hB7NLMvhb11PvUAiYpKg9IJsni5SKC298Dz6Lyvz
oWF4qjCEAd/kMyrkjBFWTz342n7HF147EB8wGe2LplaCWcSdy3nPLvC2fS8ITRXT
fKUdhOGMXLQx/PqS4EBSb0ch6+Kh5ZCU7WCg3tCZ1a9c/PF/wBAx9y3D/S/JAZ/s
hawKvtzIHXl3aA6H3Z0JlYQ3WC2shjTxpjju6QwcWkJGVnjIEhdmSMC/bhulQY2U
ZGp1cKPfLV5RPMFWvgotzAYkdSEc1k2ojE960tjzr6KD6x70IdNv+jCASDwnCGfO
C47O3W/xCPyH+d3pUBKSvr786kCyCI/DddKF9KCUXBAv5i7dypApRFEx0cfrCDHw
A7XVdxwTeV8G5dBtnXei9kORIER9xtqAGnJ1NF8qwgZeWw4b4VEHTvHLttN2qxbK
+dHpv2SO9WsL15EaXvBqspszif/dr0CTpT3xu24GnyQXCWuFr05Rn5IJzBLfl8Pf
A88W6D6xZ0LQI2VHUX7M7tdMYUqSwRFuJF18HUetbscFMRAYYOv2mcmAv1Pj6wco
prCrtuO/g+XfjRTlT0mcyVe8YVOpET06PIsMO0W6urqFsz0/gg0BElA3wcihmKmF
dwqAo4g0QE0O2P2DwQEmps8GaAgZwHnnEr5C/st8tQ+DL4w0NIdVxWFTsY6wXu2y
sg+8t12aFDRCVxSVqeIvJeIPNX4sFttZDAYFGm8kF81mtuS6mFXARpIawNUbSsmP
aVoMPT2m1yND1d2Y9B/5KbPf9lq++fDowLJwAys0+aUa7s+/+Hkdc/PqdkyTXHYu
3+F+AtStuuEsmW8Q7Y4GxrIUsKyOJvKB2YbSGf++0MGJLdb/5aCvayc/GZeZlN7T
pqaik0DIQPGUNg6IDGZr7QCqgJP19FvxsVmBy0aoAaa7/oBGHW4t4huQDDoiin/O
rFtnXmRczugv67WFYOdClv1PbLrpVLa04zihmxzziC/HL8pJsB8uE9A5rVmqzuAQ
hiuCrPXnEAvQUPne6p8f/Q==
`protect END_PROTECTED
