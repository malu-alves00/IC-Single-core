`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HoBKQ+dPYx/BzsEgVEDw/J1Kf3kMC10yB4kBkADEXymEO6OlxI7TPeboxxshcF5F
coCv0z3JRsx197qvCbKTfaXJCmT2pI1r/o3L/QCrG/xHcNfj0uwsCB5knkQh1AXQ
y82PkXY+ST+mv7c3OlStcabng7C9IIBgKuiDKdFiWvMH61c9ovGWh57u03OF5gWd
au2sG8HnOnTKX78Vb3uA7AyuOy8TUyTBrhJfqZofh075Ir+Zhc2J6PaRlH0rbp30
rktp6l1st3HD/PLPzGPCFlTQx1DWekKS8av9FavWex+DcPp4FNefr//zGRxrZKWC
D6pXwk0Kxgf3x9AaK7dYkztUKZljvwvfLqukwHngaccc4YXWSEQ26aOTFxSEGEqK
qQ7ePtLB5ERFV36mKMSapR7WuJMwqKh0Nf7wu9mzARsLVzp2thVDgxhCqKIXYMQR
B6or0PiqsUcrHt/AvDHP2nkqdu4FbINxRwZjJRyVPAYLXCe0T3Hcb7Sn5UPDj0/5
SlTCmDN91MBvOgkqjKDJoeJjpPWZy9aDGiiswwBkh6+P3CwzM4FyZXzvLIYR48Nw
Vb4jsMcXx/DtvNJ7Ea7CF+gYHjhcO3GluYaZq5kC141lShS889fF6aDIgQPn8xJ4
kNbbGrPMRmtiUh3P16oJvrqoMY5d4cmk21WCsyopiZ4HyyuNEcM/8rKJs6A+piTK
A3OXC1/nDghWHZrap6iokIiuxIcW5W57AsXRS3PKxOYryWhLgbtn1TmF/BNI51sI
xzrYlgSbLREOoByoLIAMc9AXAWson5w76rbDnqYAqigDZ2B+wj5rgX9znP0zkrBS
CVdxy9ugKrX7XgTp7S14cUVsey13wS9IZPoBoq7Hp3qrGBC+dXXKH70H2/QsxoO4
Pv2Jg5IeSBcYpA2fS2icqW/ZR8I/As8q9fhbSRYHLHzZZEdEbyZwVm3x8K0FBxhq
mgiz9GVClxUy9bk1/yG0LtmNl69eSIk9IqJwRBhXFIna5kW2xUSXolNu+DA1nnvq
0xBBUn7cB1YftPgS6LzUmPB/qjQOsWzI+OPj7CZDJXwnE8UcWPzWk6XnmtLwk1Fu
`protect END_PROTECTED
