`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pRzj/UNiqZzliGQQDKK1nQwgpS6zxXxJNnVtuf86m0Ob2ykAvCS1oFHR1dKltXK3
ut8TpSFXxVFVj42nbBkurtXbKkGDo0azyLfuvZcOD4naYtsLr7YUUBN9yhcXJu1l
dD1aEys07bo6MdsLETn7iq6vN8e8OLAfev1MFh1p/HEv0/AkTWbmT7aduw2qsqXF
iCt8HIE5Wg88+bQQ0z6Ctmazs4J53n7TW5MwxCMGWGv8EjphfTQL58JuioIEc/dk
JMqDwBKB/aNI1FiIGiLFW3xIUvDLRWBtTe2iGFRD5VUmKoUiBbUU2PmZqVbcceWS
9aT10YzFiFwf6PJBWZStHk9sWA2I5WChOJE2RhAlNbrZml/ugvKV0vhIr5LULhXt
Fw2OptmoWi1XFoiOeWW3A9/SYRh7zKJp36aUSFbKe8xgs1Sq8Nt176vIadF9jKWW
t6ZTMuUkizMPxw0zfDC1nmlCTRMsCAl8mgF5uLuChi8I9PkPfufcVB1M0WJoP/Tb
iXGULHp3Vq9RzuZBv6+A4TMfjkYDHh23jgpsjNbgtcEbXM3xYM+N8toLDxDAll7x
39WodrktKV1QTeP8dszIy3IHcpjNghAbd1Tt39/if8xVssFueZnybbl7dYc/4kfP
YDa0ubCADnFyJvwUL0v+jQlm3fsfV/QZ06mX0/nbblycaZ7JFbvTYbwhhppxCSwB
dZRTqBv/ksH9x0jI0JszumRYNAc05frovcezMeltJ9xHEvl4/qxKBuG3ML8T+hvI
GPU1HuUMFk3nAxnxcLDg3ZDDRxrA0N1qJJczzwFsE4fNJjYEFCPl3NShlYWoRG72
pG6mTTHa4tTbP6NOfs86K2rFHEzSIZONCxWKpWSkohrypvUY7oFl70YbPUkNAjdc
RxCC/qkoFWQUqnolDss6c3s4WRkCxBEHHUsnELWx/ALHj2tIwxq92AdwaNZfCp88
eZ+gGL9VZqQ8VP8lYbeiV7f5xcFGQLdjkyPOQn13WgqKnQJZu0ghW1xmlashOcnm
tIk2w/xGU5F96vZyPngpgS20nOVTyH1dFeyuLo22h+eyHUH5a6RwpqcZvP+bLTFv
QEwAAX5HoOWy2s68FM9leLqbVN0f8SyAGlhQ/4Bcqrk6rCuBBhpQtqWGldORPq7m
gL2/Kdgd5sX4jNQitdmyV0Nx+LvsFMv6lqJni49DCb0+UotSnF438cphxKnU77tA
0IMYddYaFRVToXyp5O8Rvg2mOmu+c1nf+2ccGdhuM/l2rF4gh06aEOiIHkGDCSY6
EnzemswHqmkLjEcu89iGhN7B+YVzfVUXGZ52alLLk9ECRTvf+hKXJRsRRlbx31rc
U+R10Sr0fE8owkLBgqgGRpIIGS10v6q3cBPeSsSlSJ1iFxLFUo9QGnQl7BorFUOe
RV9m8sPRrwzRLotG0gbdrs75VfkKZWK2NyojA3b4UXrEuSUPaTQZEZqznWKy0Cuk
a40T9qHzjFe/INYakjUo+Go8cYBnht5d9Iy/9/EZqwc71qrXAYwgGbvWz7OK/HBm
eob92V8Kj2l8DDE4xPpATQta+KgXVqalc66AmEBZoDAWIQr6Ezye5LPc6Di9c9ff
ldLYXAkTCQ6VAKuOlThYBNMFcNUp8UFgqK53BuiPIlj72uzUAqVjZAoxD+YyCupB
Tdpgfn9FJCy944mDlwe+CLEYI1MI9p3pDGJ3rkVHyoAmECQbM8MRY5VyEgyHe0Cz
1W2DaX9HXrpY83L2BwtnSwb7wejTe+GIdnFyuC4oOrJ9YNBoca4MuAkG0RH2k8XZ
5HKE8gPqBy09VQ/ZP9xwTxyutIOXlZzpxqA/KB6BW3dGj+0kFI5iRaehqQVmd+JD
JEaz3qhlUnm3OawVSeETSOcA+A0eB5r/JO1JyvW3ZfpmZ8uqV5QkaRDACB+1kYKH
uNEkGuc/93m1XAcROZYrszHNIZ4FTS49V356qbNzMqIR8KizqLLf9RqF0O4uUhz1
SPhqIFoM+JVHpYKxmaZjKzGF0XFjkALefOk+PcWax0h+MIwDA18JhSuV37hLaZa5
`protect END_PROTECTED
