`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Yx4V4Nx1mcHoAeXQAqlpB9isXENO+lDGIQnWo0L94swSCHBRoS7MnMfbmN4l4orr
dM3R6P7FOPpDPf93WxDb8EyeZLO1C8g+rdeapvexC6gz3mUmh8esaNGzLKgPWKGg
G8l46UPg4/svFQOYFE3vHRDIA/EPlAd9nVKJ4dT2CLGyAc/KwlDYIRJNmsJTIJCS
VzD6xJbhu27hmEwTXefL/B4ePcJ/M7RmMQx/8nzGd10I0zoQ2UwM0+UKOoDzSge3
R3da4ihucVng0glVwpbg6rB6Z8NAMZ+0NpGLknU/+ZC32BflZJN7uVqjhkoDVeaA
kSxkX28oDQQP4h1SChPBv1F6hq8CtnZzQyTQfKm9vBZPrANw8DaW1Zh7tS2Hamgv
e02mpo2a9Ti1z6D/JOALKDd4SY70d16g+Ey9/W+T4Ncw7bouWqwDYhiU4KH5RQrk
3BY1DODnUO1FfysPM83LPZMj9nFszVHlt+OfL+HLFSXMVby41i67DUOChqVzRlmu
KNCn89SC7oPrKq1YWhUDmYQMq+y0MsmG6qDA5auO84dkZzFnSYSUlt4ZEX7quiyC
1xFTHEPxjDOQlY9Rz9TyZ4xJeT3Qk2AOaqdsHk9hZcHHV/BVDYWeO+BLKRQ/Fbqb
qUR2PaNUFC+K+uz+LOM5/9Fyi6ZlXWwjEBKKLVL1TT+7KhLo+u8KhT4I8yKplMJo
YlZ1gpDmmyayfvtuqnmQCubi9UkLgcY5fQcQkqbL3wTkfsI0sj3U/RWV1UQYlHov
u9XzJvEyLoJ4H17pRi2CymZWzJW1lGCcGVYCJsjCAa9QwGkkGUuQjr2HwRPTkHwX
s9iOi+DJhoJ6A0QT7LDSD37tHnxypMLkeu/B9IsnBapJl5KQANdoIMOidHFInnoh
ycjnZ5pJYv9vRajQWW3TZYeMAqA8yuR5TvTUXlRFEj4Fzww0s5sFXA/cwtureUX7
icEIXalr0Ed+y64zOzRxSKOmCFzqeTEJwuBG4s6h0xQ6CwxU0/42UFtnu+cmejho
/w75R2Xg92O00PSQi50fICxgAAe3GrdxFUFQnz4vlqyW259+TOyC39cfr0dbYzBm
ufbiODGJB+x79eqMEr9zPp6wlLkePQNs7i9kFSDLpeb6RQKCNCLY3Sp1iJn1zezE
zoUdDY3H5+aGXDZu0ekeB6nvDx7hK9YSilhbkFDEjgErikkfOJTrk6z0fx1yoKoO
ErjYDrCcmjFtxL6g1xSFkWsxEpn/E+sS5tg2YXukhA5L89kWeffshLX6Uy2rXAnj
xzJsO+aAtJEaq0LLscjRXg==
`protect END_PROTECTED
