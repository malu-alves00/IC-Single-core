`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+OO7iDVhc53zJ8p8nWAMLWwXRrlf/hv3bGoFnmPvG65sRUyW8T9Xh1DUy8DkTapk
i7kYf8ssniX7L0cn/Aw3J75avz3gD7GUNsQblQQ+43QhZIEX/6elRXZywd2FFQef
4SMxlYaIF6rt7myYEnAFKEKg9RSn1YX2K9pfcKgYyDoXWJhAkBe1WDLEBidW3zKv
TaOHOfHHEG3mukX71RfWR0CZZ92L+T3M8V75zL0SRSujF4OyvaBXREswu0Z/Wl2p
ncvPAN4Gq3ovxrIzPOppUzTvkoUdj0Grppxqpba3vJ3eo6q0LdzhqCzoTh/AeR21
W9tVO/rqr61ZG4NgedrVguiN4ucKIBj7LZRy0rbuioEnbsiiG7lYzAnXtgFPbOwr
wszMPho9dnA0GvM24uXKR2wdsTj1dt1XMkRXRsBeJuq+gbXgHjkceYs1KyTrWwDf
fejtebGtvg4ygmKZG+yHpSq9+Gyb+lyYBgXx9FSVNzZr6f0aah5K7FmwrKwIePru
5E1TXY4RxHIkpf1p2a4/Kyvcel6esp5ntoEbrEj/uPqAxI2g+hj7hZG0vdNUwV7z
Y3+AQYDROqGMnrNOmI4gzf+bMkttZoDc+dHHxh9PAZydta0qR4k650EXoNUmvtm9
941xswI7ZC/h3RbmrWme7F/ZUmX0nxwyIrdIFJ8t0VDLN7yRLpwQtl+mqNJttL20
ux7bw1AVZvFQSyWEgI2NPeUsT9cMWfJ2wj4XIeijjSbLdWjCpArn3pNkxvAaPKB8
TT9qkpqRDp7oA6grjRQjQ5AQWXqzYrS4SGIES0qdBnQwXnPRYDA3UZZp0LJ6IP9u
DCWhWviV/rnHAn491QS5kbi4YGZQplx2bCS0lc9iAnApakufPdk+ZkqKlfQ798/e
8C2XRglTkz6yaYqduyXJxbw32HlM2ssNNtCxtUFpebojfwv/a9fa5tIlAWnfDTAt
KM9wT+wFvgx1K8ruCtWlTmzaVsXM8rUOFkoFg95iRHZDgOMuK4l2tbkC6t2dZkpA
u6pI1tRLZP8M6kaHshizwSbREzM5jdYl/kGGYJyC0fu07OwkrwMVgHfgVa10suiT
sTU4KCjbw+Mt3ebMHs6zbTpyvPlZxrOsXCU3Ht7SnOKbDx4DPq8gsvkZ41cGZCeh
KiXuCNEx8dJqDsUKmbckg2UeUp/64HaCUhpWmcrQppzU7MXI6Gh4zaj6Zq0p/Gpn
CtuPbx4OB70IU1n2QGfk26jFKHHDV3/0GD9RsV25lQ9Aj6rS4O1st4X1k7iCggsj
ErsBFayGyemdqC0ebC+QHwcBRGw/VFvO1oxRGYzRAztGyopDg6kMYTDWefG6xkgz
ca+MutznO60zbQ8aMAl7D1u5/OyCTZ+kPl3ZnYq8UINXvI3uOts9n51iymdIKeml
New1xm9gAT+Z5/RYK5kAilDu30Ky0qbpSN5HFGJ4pG2a7inX1JXSenq9pvKd+BT+
Sqx7z2agR++SKifmZGNWk1pcZB9zSIDx5eH2esNI0BoSB/w12KslyjmrjpIa+Gle
uM82ouunCGsKbD834rlY7L7hY7Fzt5MJmPgBEJIr6QPOntPVa+MXoldRZFIORUNw
QOhC8miifkEms72gzJiqB03KB7pmDIvEEIkoqIVshJqUWbAnDcXN6uIRF6d6Ddld
OPqVznryMDNoAPHySf/odB2XHDEu7mdrDKskRgJPTeq+A4NjcwfTDIqUVqwMl+c4
7JOCn/PHuW42dK7Z2NlvsoxlW8xqMB/hNMFpBFeDwUQJni5V2OeyW9Pv6z/02WWR
lbXnfF4wK5GGm2pdJKVkL5sQLbMTOT0E8VvAmqMcz7VxP4OG2BO8/dYc9Tz9LQoC
W8jKJkbN0Unp4vtIOZhWGAGdsSirJxpGMXn3cnpZBOMDrXyM/t+FNpSNXjDhYroA
bB4AcAaaz4klgW5SNZQ9o3Fo9KbHYVK4+au7Z04/Fa4imzwADJ/zg43KShb4qWIZ
+eacdTU7h0w2IgO/wOsRy6y57zlqiQLIdS+9b9JyjvSCmAYSQVKBV5rGjkrpKvq4
Wm/GVLOw2Cvd++XCVfr1aveax51pyI+3WFL+SCF24yffPebI+JClEmgj2u1aduLt
N1dGE2gb8OQbeIDPFBONkt2YPHEFcl+qCW7VgOoaOy9xqd3I4JiOi1eSDhkBTMug
+TTmWx5ylu5v0ajDZPaEw6XAEq6+EE9pqp8I+gWWtWI6+WMAl/Sda1zkKYwdi0Ry
VoWL3xakHna/+BvuY7vYWlUUQN53aAL57ebS6xq3dUj1f5mfW0+CXD0TT2PNf59F
0vTixBce8yolaSiyRsp9tSoiZvCyc0o5rknU5tmP7KuAKC8a2bEwuORLXIbuAfkN
mLQkv6/fE2iRkHBMb+VOc9a3t6lP9t88mNYSSIizEz71ckbb6yxS3vnjdY5PUeti
fjnWVVfu/wQW4d/A4ONHlcJ/qL+uCAjj+fNSvn/z3JIZRJ4hTYY7zzdf24PM4pqQ
unRdlmkHd9D6ZpnzWgkxaYU09pI/6XpGY5BIoheP+OUAl4ud8YK4Nxmv/lGOKla+
ngG0njU57/sEpjBTnW/n4qJvLn7f73DpOfwRSmXGF60n4Wq2m9FirtUdcvrgaovm
NnHnZoZtLAhRWfu1WR0m0j/4LhbB6Vtj9LTtEJklgp9XwflQ5m/DeAsPMVcTTG2b
CAftPhX8n/dGa3xiYISJj2vFegEVi4IOpuFjRnijyQsjtzjf5tIoCzIZlllvxKht
MJ1uDo3vnfASeevFqPxcxb+6fO5sjC2ibBHzvt66Uq/HE3kwJ0UygVHiiFDDkWJQ
y9q8/nHKcfWE6mnHhczEbh9Y96BTS61G1HItsB2d2EeaIBAZ8AsiAWYlZyJQLgL1
oVfH/+/1WcV7KQULsNhvONMshNEfC9DIaJkATfJ/rlERpf5rZh/SWY8Epq0eOQ62
Ut47KEjC90KqLRAiWMJaWG+hIkeZNSe0amLD7HUzC9ZDKBnncJcGKqrkxBxE3vl/
YqKd9ZydbJWo8Fw1konvL8m3emsoeO8YpRKg6DMjpoAF3jVW577ls8p9TZBc3tkO
d7FOqYUMJNiUlw58RPLWF3T2CZ5sO3z2xdMX29vVvCrliJ0fCbr7yTgAIix7WzFs
aVldCeIRhwxEiW3TJBITXkdgwP0ZJ9PLioFhppN3n+jyq7g5/Ann7knbmKEXh9pO
tI6ITgTFi469U+2jsP6D9+2iz3MuMZbdXpBe9jA313HTLREjBVM0df8G3+G8xxwt
ibdnjR70bXJYXVF0E1RgNUdkGSPBpnSW/enNYhNMqR4ynoDupFJ1VfOZDn7wzD1p
emEHhOO/6eS/qvRL5aWkfvbfVaz+IE96e16uq5tcytVURUGFLD4LZMow7/rrFKeT
fli838393fWhkV9vhdfTg5SlxhU+SI+vgpLk+2wifhyMqGqnrRIRk8AbuqiTcZ06
lrudA76uoZq0xVZYQfqNE0iK0AjIUcSe94UU19Qlzi6dAV8FzxEYhPmzMdtEmE7R
+A/0zSjnjb3rbZ9TNf4qejg1+w4HdsdklgVqXQx3QwThnIjMRB725saVnhgHoFk3
3Z1ptjbUw10MoPbQ4OolgohbE1VGRdebG4WLF7A4RtH+1/6ZZO6bnPZuYNteJP00
E7W5ADd64FC1LDQuIwvaGsoUoc5h/7IQG5fTHPkBfixIRN5/Z4m5svGvY70M8wgp
v6xD5JEjcxoAwsdVVdAxvr3lcx3hO29+1emTmeMnTkqxOBWv8drrgrgQLOf06TSC
zrUqpTHgQi7XctWbqo2fpLNnQXgofUeE69/9oj3b8qfygPhR7s8jbYIrIdJtOwd3
/ZVp/ZC14JW+EtBmyIgePldmBd8h1Egu6ghRRH6MbmHPaQU6x5d7aoUgialjuD5E
5ppboXya6hqmehPBDDvgyCJk4w5cdgi83jc+4DQv6zX7jBQTzyaGgWB+3xCGWWeW
Ay171viDdXG8bokw8dZo00OIe6r5p2zUbBE25DU2C8dbfuCCbLBXVmIsWA3W042R
7R4LHwV+zwAJ2LpME+VHIkXCt02j/l1/U8WgzgMC8JIHe13iR2usZozmpxi8FP6L
RCPA8n1sPDfcIqIUKxqiOf8hvOzkYjE7C4oPJbAropJHl60yl5lhHyWf9w+ioDqH
8TeiXmC6DGObD5Qu/rdxCZPesUMzLInuA1d5i/eUxIw6maaSkg9uGfEShAnCx5Qs
e8qtMkjXJOdeSf6xIFiQmakqosrGehRdDu0TptBdUDZu73LJSszyiNzAvA742Zr+
GoQHqvXa2l5db5hxkFiKxU1uaAJXGeljXGrHjV7PeuIEifmRujVIUQCjHice4kqP
g9ajVMssLHDplFe8eo/iJexi68x9H/PXeTjXF40/OEEkmb4WDlN5vZLCHIRtUXdA
b94pFDJXRG4KUUvn9rygwRquCU5Q4P+jpTioj2E1+x3uf2HRyPLnmA9BOaWXEQ0l
KUalcLBVlZgW+IyE/hSLL4IQgPu3wdfWWFAkoc3vp4oYPU74Ubp2PrdX3q7+5UtC
QLsTtLOVOdc1lXWgcs4cuMFkkLPRvyWSJlPFLt8cbxzaPTsZ/df/8AzZHPFtP9bO
Po1etu6CZFwY+MlswNkK2eE73U+d22CIC/191I5YYX0a4aBacJbVI1aVN/GrZdhT
VOKTagU8FZNIPsCG04VJdOBLr2DD/LoJ6Da8PR+xECuqSKcrq3LXWi0lE6Ci1mUx
YGKApVlD+X1MSCPnesBtCYfhgQBu/LqHteqAEhJ2dwvyWvfCQ11EEWGdA8/2dnog
lyvQ1lAmlOHqI8dgQWl9zrBvdvQJyxDvCcoUL9paRfSJeTNFbQ2HcPAt+vN1qUR1
Kzn2JTeqooZjxQ3+U+LAKT5HBocaZCDjns8SY1yPCcdFGTPSrfSiv98bDXLD1CrI
BbVW+o8jcwQxsF6d5wLyMD2/AnGtYze4ZQKfE0BaixicbiPIAYqI4v5HC5EuI8aF
F0m25j4GwVApmdd6aYJEZuX5ekPqJpZrObkHgkH9CglCic/x6NOk+vi4XvdXQixt
UIr4TS19R9P7B85jASze9nNDWx6tw8wNj4tTJCbp0lW404PY6sGultgxa+P9iekq
xb6BUKqCc6N66VHzSMa9uvB/VVuySdHxnEJ70EODs4WvGiMcyiIYtUeZbmgjuKt0
7VQyH/xqVpzNwgWJuq685WgQEBHLkG8lderMxckDUKKd0r4qb/B3DGo8+Mv+2dZa
T6J5MTbMUJEnJh4MzotYU60XWhN8LUu8hQ+JHZt2a1QpoBpHXxqKrxj3UyDbKTxt
6Veo4oUkEa7UGscZnLk1yEY8yfAi9vrro6LLujOtvLyPp23q77ZGVqboVkESDHo1
n4SfuQsERHCgSbHowYnOckLD+Fb9+m88iqEzorvNnKUEmVbz1w5OCna3JymOWjnA
jSRThZ6QF6XXf1f1cMtxiUVQxjlFtgHUzeW6Hc3cfMqduyxK34YYPexLFESdaAdw
MzIzauzz7rhPFdDux5xwms+RsZcK6lLp12tpEqZFfTjQaPuh8NTeT72w2x7A+0em
fcj2StBlLX/2kBR+024u3wD6iF++UYDSTSctVIFXRRBGjqcLaQHVHBW4WKKoWHS7
g8vD6nRzcQT+nb1rqw4lTZc3iYB70/cv1Sa9WPw4CdcxxjtmO3fHHCiAEKbbKEFG
c/D6VawIM/eR1mlWArkLqmbj2OTrOKfxuvr5MzXxjJYPmt7aBbC6obvOO6zqzn2l
wogmNI6gN8DC2UwXvdqT3zh84JLmRy8ttshyMjw1bEEpjgxIrp2LYX2sRdvdqNkq
09S+4Ki9u90toRjeewCeOXWbZ0J0Gz6n3aMNDEb2NOeDMnCIesiYA9eA1hJXownJ
N/M0TsIaBLek5OzLhHiwBnPh8+KQqHl6OmxWeSd7oFkqjM6Hw3AIf8riWGezA7Jz
uIskEtpFgL2TmFpjwC/ZGNHjTMiIFA3J4Ib+I5nDcVEK2eozjKZ1uJN4CbqIAHq8
+N1cY4Vu70F78yF55OCFfglyOKT3raoIKnf0LFgsZHGtOjBBZmPz/qXr9TTr60pJ
DsNc8s8rVcDNU6HBsnFql78KpqqxrUt2uxzMPGMYYx8x7Ujrqxvg0Ri/9z0C1Rrz
bniVEo+uwuow08v+kjvyLjWwzFzs8YW5Iy021xKfm2zOCHNGsyZlWU5mwoIQxl0H
OVAx2mYkXuO9kBPrhkYhPoEm5h3JxS9CzbF40yT4zVN8guolQcvTx5HKTiZA0SQy
ikgxNxqX//4hk6IxHEyegwaJUH3b+fUv4xyPgOmUS6x9uNnESp9KGyqtnL0msRud
6fBuk/OMe/W7zyfEt35EqNdQjEMyDgauKcphjYEiESWhyKful7rh6d5RhXgdwQlh
kqVKKbzyfqAfWtEwg5qbo2HyraLw31O5f1v/I6LJwJo0eORBe8MfpDmlGYT9+0LL
f2HPa5UlquRYbPizrZz/Plfjs3fma/KUeLs8NwUYULqPfKiOrSkTnZSuppaVi8oe
FS1FBK3eyEA78Xt0o5UFYpo5YqGbAwM1pFU6GOQDwDCTXBkuAfvXAhWGakg5ypHa
QS3IeV0jbmiG4KlI7LC3BvqVMZcmBWswdcyuvE9EHapPuoI0wi+mz9nzUT33eSJ8
xXwd7JtcuL8/kObDauADesbQZho2htib19IOlSjg98htrcf8cUgdwl/B5MnhbJtm
9SI9G4zLtp4U3MmKrNTJoha3SlqFYPq2jhIYHFvKuUh001eqITY733B3PQopUHV/
6bKUOjui9I4onyb4eJioar32tVtHUxYnVCuIKmFv5WGnKmLjsr9p3+QqbwiHfJsc
QwTJoAOo3WLduf+Xdv16av3KfjLMhcRWWUUfclzvajPkc8fxlb4bpuqEVB8OicIs
GCuOQL2qEf599DeCs3pz2llkKN/Cm3CgXPNl3QFYYSA+nYFhD+KxbnutpYj5rQrK
ybe9LC1bfM5XhtG0nlM/1NI6vBlc0ot/ARlPn4KvQC43z5sXmXjO2Kb8ZrsgGyue
3CGWybFWeEV3UVnA6nptBXEmLJS681yJICWNvL+trgvEKY49zc+39/9lVs0nZvyb
NM7ErzYWyxwHPE4uOY+o628Fpsht+UBAU4M4qq8SsipwvBxnNg37k3WFpti5VqiE
4FdCSuTXK1J/nBHgwknr4gAR2FsIj2QAW60ZbzvTVKs0FOUq0CeZ7NRmNqs6IBqb
+6jHBR3/TencCvJPREwItU+q8jrMOhkpshfprZ9jBzSiOQuy+zaDIr9/aXVj+ka8
6B0LHabh2+rS6oqeoxW70qoFs1kcnD4CA7w/yL/Z00MBy/i/jPN4bO8zlbRzd4tz
KtfiNKD+dD5ys3r6nlB4iGesLt3eipRYW3DqRDFOF91ZtWxIcy7k7aW/0WYGx+qj
b1uJZTbxcbY5iRdzS5PI8KHidovpNbe4LKaXyl8XzB1Gd/kZmxXzW10ABpdO2bPQ
LXwW4QAJIjX3QoP3s9GdrOc5VT5xbv3AbTnUB4UWC3a8ncUy0hKMiMYGqu/i9HOp
cnt+HBEAZWWKX/LgwI8jN21U+q76BrkH2uFTdLzhp/br+C/jvxCzcs8RSBSsKKPb
XvP/4F3ZgHXEYm0ynNTMON8W8o8eXUP4LWErJOw1RVdaG1BrBT1PplrYOXMuDoqd
N1m3FDcvw6rjeyRjwsvAWwxr94C3DXIbix+Q+eT+oS2w432QrsVQjrqoG5D6L4qY
rJO9btAdp4gpfbP6LswntqlC1dDO1KsQ74n61Pk7Fh5RmDM+KvVK/TxC4rSqHEBm
HBYaXUY9K6lIwuS7cdXdoESuTlHKe4r0WKkHyyKdixoszfann5P2BS8n3WgKDDb3
mEFxnwwSRx0MunsRDS19y3NqdUEFfOVMjNYpQA/bAURFmEG1VWkFtmGkOtwSYvKI
awYHTqwUfbG0JWh2NM2S9PSkZMwO2u0xJzhgYdpK9czAXIMmiYGX4R0F/UM8hm26
t9usKngHAkTTV7RwRAnETRyNGKLLI/t7i8lkSAniED7lsDRgQTb7dCloW6/Pm4Se
E8A5qHkzvuwZYIMvQyfviMkKMSWkn2AhxFKI7fSWd3uLKPP+keUrOdDVZGyZnqNe
5lb4+fs3ycVLcxccVVzJijOd5OETncxyH+I6AQDcZs8EQ4Xe6+v3JvZGCCurADYD
XQa5gxRWvtbjckhO+BI6EBO0sLIO+ORZiR5GRcban5/7GQzXSkutqc3QboDBaRHc
P00riDyUinbcfmlzIGvrn/kcuIykzqjrwg3c57YwvCnZY8uNPYuKtOcmaDIomq0n
3+RNiPl+YXoL0SOJgysADUabU5VgP3th7OZ3QrnTLidvmbjknZ4DWMCQ9w1Z4AFe
rqkksR7rzZR8etEqLBBtKonf09bILNlH26pHmoQnzOdqxQfh2w9sgfkZ+vo+BmBz
gyRIHi2gPOqn4jE0oJ5jul4r4IQXdWPgz+JEaEswySYd5rpPG36oe/RWtvhpha8R
FiTkWBLpG6RKciPmciT+7+l6O83H4d4NZs3DXycvda1no0J5JgIB55boVO8LBtqB
o0Lp/O+RD48QMhCctAiHebPbsMFcvPqyGHIzqA44rkQr+Fbfo068FEksT1xZ5tIK
EEJNB48tjbaeD/xrDbtzPya9Cw86tN5bwwmqkPtb5kzXvEUS1196bwDDsKJBzu0w
xd33Y4lx88HnqRzuhmghEhZL9zLSe700fjuSLNSwMuyN8isHpnqxe+ch21VdFW/M
oC7NqWs9zOImuAP4XViuR6KhWg8QWn1Gwxrnz/bR38Ucc3cM5QJoHIlXjE+JjmuD
zqS5O3Gm5j/6FfxlzUtwR7GqBNN/BYMfXcDR7feI/ji3IPD5r1q2fvX45pgZBZLJ
KpQkOECU5q18/YlfM3GfTJE3TFcyt1Sf0VyAL6abyi3rSxKMoMbKwV+iUjVEXOFe
3i3fj2oQg3hOK9/dZZB79/FmSDUCYwP4el+7dWV1PerbP16UmPz9Aetx15xbk0VW
aQJRfZm8VFvjwzNbIOnicEelwvtE5z+MUV+b00uJoVe+BtytKeEcJmmo949WhMPI
xjBm5mfApJtMexczqdg5ZTCJLncmgKtLNhfZ8EtaTROluMQ9h4VnvjupFoFcX6yy
1MlVmy8ZdvSOcfHhqs87l86ZsAcTZMZL4hPO9nE0gPVtWHVE9fQN8zgeI4uCMil6
Uf695Jp3eE8VaHuyt3Zk/qwkGFKWg+mLKngFj3IFWD93o0yWIlp4JxHkO+/Lu78B
aKJWu+Onawb+l5fSpdLk8T+gY1Rq+ia1bDYOV9VM9UZpeUuLm0w4A9COG1jX5I25
qh1sBFgNUwybdj+Esfnwq+4IuffoXFtOcN3yPOXeDnJyA43UaDw3ZG21oMauisja
E0k0R+LYx49PvfTKCRkU6ZfG8wZD7ZvYvvVPO1pjQF9saTulvtI2DbEKrD4zA8Sr
aaVb5O+SsKpyUtmNzGJBKedeW3v53U+itSmzEf6Ze81US6LaRs1RWE21rm8EjaWw
UhYNhDniVVccPu8EUEN2bIiFM4T3QSRqlSocoHvzNCJlFVqtmQia7OZTFWidabRP
2kPTg2s5yJRc4UHpaVdItM8fMY5NPwn+i/NB/3w51ggjAmc0N9APsVMK4rIgvMa9
UqYCy+iq6yDFjOaBc4/WG3d4FMYx6vPyv/0VWuyaO4jjTZ1LvEdjDkDIKLMz8Q3y
ijvpsYmPFZKEQ75WLzJsfogYG6K4sWlTIfc/rQrw5ows06p8MhAsmrwqbX3ZAP0l
T/oV2S2afZEHiZ0WE7mP+VSSN9KaYHvXKTMr9amN4xtPyewOO7cEL2sNmgswjVU0
zMgBg2nn8dvhkyXa2yK6YsTiSNpPmjptkN3/NLIiWxDo4BXXq7UbazHJRgYpR/YW
UWmluC4j4tBDh/JTy6SCIcKfoj3v3gS933bGF5Rre3tyfNZBJDdElE0t7OXDZ+mV
VR9JpAOjZksNenWrd7Tv348X7w+BbkD02F0T+oY33bRqHp9r3iftsjfxLVoQnHuv
bQnGES89Chn7HVqCtM3aOqvn7BjNZh3Cw7dSKv/2X7eljx2ptiGuiRNon/X0UYYQ
IDxwm9aQ0o3bRXgEvOXVXn6siofIiuXnUmCXuQNM+en3AzsgFk6VK5DAYaf5q/dL
dR2qMO+cKbeEZoijwjreJTXWzgx7PrpHwAkAxXhMHjXTFtJEsVUUQDZ2Isrv3Y2i
dBqNne4Kpr4Uhffl2f3Jh0T+fY42lOCaoZdw3MwxyjZ0V4Clkje9TCDY20J4YWIp
Wnz/AORnwxtwYPVzac1uauVy9iBsd75Mt0Tj9goKNDNzrwgAWzh2fSEvg1V9S/PX
tb+hfM/h3gUlAKKG2/AV+j4EX71ouimMr6gkHVEevsmVxZCeQs3MU4lNkhIc0yS4
l3SSOgiex1E5T8s9xh8fRVT09eS3ngt6LeyP7hmTm3V6QVYmTIoaT5OZEv6/GvR1
A9JiU/ePhci+WK7j+pCZ73dfTFSzXVaZ1F19wb+eVuecKRKyAS9jixbMPjCcLxCt
oVqGkSSWmbGXTqHO7ofOHC4xVk5dY6Ly6FEp27VmZFd+U0vE1wJU3vPudeK/aS5Q
b6weYm2JrGEyttBIXtzva0Cgj7+GMd4ZIZutajecm+OWP38OpeQM/yXtmS1XlhE2
MryLdgLqi4jscdfiF3uYcVvY/E9EtYeqJSHVfRv8pFPRcv5+yYT0VmqHArBbMkjw
V2SSS48lBEDyOq+z4k0muz/Pz4/kH2X8Ne0aNV1XiM+P/OhPvCrFMy4WW6NWG73i
+NUT5xPkZd7DZr+C2+LerGAWixqdyN0TzOVkiwehfBzzpOPYdnK7nxiJwgHIMiGI
s4pARS+kOenmsavqxgVKTyh3E93/K1jiKtijz7D+DoyR6lFSoAVTQAaN7vGY4spx
+UFSN980cHiyAwWblXGKFcl/+xz4YkeR4bUd5MnnVTmIF/OWHvqUHUaSWJJmB/dX
NiEVtgA9GD5klSZN2+X+rmqgBgRalfS+ElKENewIAKHookbHngy4QYBi5oX9TEaR
B2MzdO7Y17+FaEBDWoBuHSbFHwO2kPnk4gypvQDywlxWoAVw/rnF8Ox9PB5tN+L4
TfoY75zh8z1lL7B2i8kFJktkqhiRWQL9iqtXbSRke9J504wuvxZ8/hHQ2GoHOLQK
oEZMfsUsvVEsrwptpieUmTs9/owe8mlPDN4M/g3LURmaM/qsykhg06YJsiKcjwI5
gsrhmPCGXkuuYHT9BDN51BK7pXXsg3UoQQ2RYRTNgE1zjAC3VFWgpFciraPv3Ppx
MoV6L6e8T33S1PJwOGDXVxOwvyjh+tCnBQfU3n80Asb41DlfLW3YEepVp1qHAvht
XHujLJHPFAqWu2Bw9GprStvWDI6nwgIGvhgTyBDd3sJU6zRnnnCBwSzjriEIhY2P
pkrJjYQvEfhrfUtrvOam9xBUKSIO1ZANZa4BLcE0K/En/g7jqd+t6zRrBFdpN/gj
lzi+PuA93bm4Ms0xPhB7vqqfpINoiI07fj5XR7NCamIGiE1HSZLxuiEHy//GP7F7
49I36pvs8au6Y/UffbhiLEEe4jjsoA3BmXzfYB0ahu4SIa193vJzNzd72ToQCuZB
TtIzfVPJB/8D6QrAaN/JRMwEN6D0LuoKqlbLevxeiRMxqeupUP8FkvMfeTOJmqQg
02cSjDBquxtJ/l78ZFmo2YFlaT4/BC9BBblFasnr7tVG4SqdDmzp/zAInYBlc1j+
2HQ1RAj9x4h0yFc0WSrf6q3en9HcjHarqQNT/LQGbgWyKDlky2NQqVU5t1qwDUt/
LDqgN/OQVQze0bDr/CePiNrwlN/Eh1ifY+ddHkb4ur+wH5iFVz3s+47e1glrXHTR
iCFp3dC4TGhhrj5FfkyFdExBqz086cK8aEcdG9lxypW6cMt4D9gNKzJACZrSGUns
UYODqcZBtP359C5XJs50odl03V4x9Wv+uaSveuOwLgphzQTp6/xRnZyUiCzoNNab
F49mUlgovh15rup6Hcr7NoUD8YpM7u+r3sgJWDjNrFEFV9F6ir/qNtNx9QbpWVTi
Wg1lzWEUo6oMWl0tJyLQM8rz01fN67HP27fcfP6yywaW5nxi2isDHfT4vkRdpUbm
kQ04beap6BJuZ8Uvxp01VPvXGdB0ScTjLTrVSYE1nBDsTQkxxe+FjLv9ja7Uyh7k
VVEvUrywn4qoIGWeGWhuuKw7CWQ9DBNB0tDiPcOQun6VSVpsMSiRLHMPiodqkA80
WuRk4lcGxkr4WUcfOctF6i7bWZhRmDoCwAyWGVb4oqvUi/I8NutLFlVocCSIZmXj
I67207Q2yjoOq0JrCFJunb8Jyy1WZYhVubYhoPFEuajdl+bxURmaeR06EE8kB9Ei
2p6rqQWOMKYa8df6VhbnbLAylVQhhQlRDEtkGZH2Td1sb4K88B6wYlROL7rZg716
SfT4yDQZ/Syuol+RNT4g/PWElnMYOvgOIO4uqXLh1dV3VyUM7n5vgbxPiv1DcFd2
FolfByG0Im3JvlEKq+2HBblZCnTsG4OkXr5eVAThHvYT/iF2NYpeWOjMNbnN2Owo
ymVqS89fVhuSt0T0MRkm5iZjSwLUMwd0DHsft8patHi7Bt0l4Td2STAYbfL8w4rm
3pIPJvztEYpyYdj2gB1lLx2aZuyMSjHd/fOC5v9ZymxWKlIPsvvY5a5F1YA1E9zm
MSS8SqGtWmKkFGpxuD1qtvQr7cFfLWaGnbzXqV//ZmwJXWOAg12eXI9KV72fjFfK
pQ0B6rzEs/Xm6H/qQ/Ta8A4C/grVghiMPIJC/1T4N9yqruRohhgppTYbMKCgU2cv
OgqzIh93BicVh2kXe/M4tiyhgp0MXj8Ur8rjNoa3MGn3wR6xGlVE2mhuLvWxhqNR
K38aOi7lutxf/V4TQfBYTOXhyKdoOFz9BY0SyFOrMbqd71WgifLNNbAswKBp1q2x
yzsdGYOBCkCc93dZCHRzB+al/M7v+C14pocBR8zk8FuZj2+H9szb1alud642Tm6U
I5Hrfmb1XVwgQDweEZHRk4ZY0fTkZnA0+ZMacRjS+k+SCBNMDxu1kyDqDNAeZMZS
hVq3A4bqmmrtllEugUREVF1ER+zefQhQLmTKdLCBdhU/yqNJaJCS/rsxD0o2fjQw
coXT1I/33SPDmmwSM+kYjmi3c0KKaLX6YuMgY147f+7BERZmZmFDvJN8o2rk1L6g
sJdshiNPutXZSFSpbVl2t1B65Ay0Iz7FIrxgJnEjHS29nG9zPsKKjjueeE59ZZGW
XNOSTuwIq9Z02PtVNqPP4yu/M4gyo/uE1ETzcKNqa+0tc/Qef6PfaXV53z2e+f6X
9IA+57COJDBUILP6Y+5elBwbzGK6qlEnTH/irzg3vT+D1Irq5d+jt1Qok9Cp6X7r
zlcxmP/w5diDSKEgz6KAe/7CNZgzLUWQCIc6AYVc+LzcBy76D6W+wiZjpzJc2cwk
Pz5vwGtA4+iwC9OK9XErV4fpgO3VoI5uqwe5mg6geIyFlZBSDCsCAOjXws7PaLFg
2fs5rehz5TEBK9QXQUgWeK7ivD+/Sk7q/U8ZpB12+yfYxifRtz5L1HnG1PRXoWzk
e5u4BOgcAYqVzZPVpl8nLWcSFp/KVNLEAZIxdQwWYIxiNzEsO9JZByHpnciUphcA
BGL2deQFDnYbuXeElpv1wAjfbmleCK5vXLjKynniFU8u8M3x5V+Itj/53od9FCyx
xPsG03pzPdhc49yrjrEZl4sli5WmGqrGeowTcUig8nKljI5JGCkS7BcWEsIG7IQ/
Nflfftjx9S56mWz5cNsV8YFj8jaTfRYr19uV7Uvejqzn1GeuC6jFNtzuV5jhDkMI
SYrSruZyG94JufoLIVSXAc1YwQyACz4x5RiNrCRqyAh2ExKEU38bYCFP5Ptor/S8
UFKZz6fxxibaqVyhBX7QN1pL81OmuJnXASdvr/KCor1hKQKCTfjh+gI6/a2aWPlU
aPeH2GiEkTnqRKsFc3cexx9AsS7/IzuB/O9PpRtaaBg9tfXPIyHXyOGxjBxAIqHC
K860w2Hzs4WBen7gKNlQW7Yv4gZm+E0tUgbOYnsNb6Tb9SLXwNCahozdbAJuCnNd
HjGH7t8ttKOJe3CxJlUY3bM7ISMZJCFoqjPsCNqjaT2mfuEFFstnmdWjz57o0ZBA
BAnGBW8V7MfSucLwBOozwu/gNJiWolIajEhjTmZrTBKcqvP/3VzG+0pGa9iH/5nZ
XEn3AnAzr8R/U+V3uqhu7/nPu4P6kjrvX3xVJyZPkIPQk7NjBTU/nEj5ID4Gm9Df
EFjmH1H/ghn1sEEduYQxP0Jp/+Ri8wHU+ItrXQA+GhjPfAbtG3xjbfWsDxaMG9sX
e1OOdaEHHSUirJHZ6gY77jKO/QX4zjlN/5BApsKiDJAVfxvJElmP8fWgcSMoHbPh
0ynkfmKuqxklWK9mmbrYxyrV3elMbeJQUHmDnFW4zHijEwHEsnyf5Ji7ZUU/92pq
V+J07auacXeoShGJsr6X79XOVz/HjEN82TqzalnpyQUmjyv0itCaHu+/bpAnagQt
Mk/oSdNaOEAmswC5wwLmXSWVt2cTZPINho1zX6mN/gHgBPq64jfPTJpRRrPYMeq/
s8r2qpBjQK3fKw8nrsDH+ucsFQoJHukFbo2+EP6kYcNVPIilIaoIagIfufigkagX
3Z9fncq9XMKAp0DD6DcU6tRTJPHoZAL/v+nSih90/I+kta/VLUxu/9bvHALPojF6
af5J1kavIuDUszhXEXSqwnKGLQyOCIXzy24shWdiY24HWpenn7N1fn48k/s253VM
6pyVBv9zfkyzpEpoKY5uPP6MAVQ4t2f1Uf9xKhb2XE0TUG8lm0KeGxESdclBXvnb
thI1n3cDaHl6cL/sggVABYso6ZyWjtfZsGGnXeP0SurXmb+Xxn4PP286/qRUe6gl
XE+0num1A5frg/pDLEClJverGBry9Wq+UjumaNATaEvKlJ/Hiy38U0qJWK9bPan5
WWzFxCyOrh5+/heMCIMWhIVSOs5rBJjI/FQnJ64aENJJ8c3kCXMA0sIjT26l3o4V
RCHBWeHVjjGD7AAT+yaC3pehMjZPwPoBJYy7sD4F92MnyTLbH4pt2D/TWwSfTVwt
EKYEMMKyShN7sibc8akT6MFepW1w4XOI3+XP1INw3UZNznacu9iGN3lPT4K4tPB6
7WygCunTgJpfYsqKlZ+5+4GPgmUR1Th4gsfeGKm/GsTgDuRU9dg4bhVmZ5EJ7HPt
TJhCJCPWNEvLwk2F/hAmv1a2KMlWcaOLjPil11yOxxTHE2MIAvD1JwTsxWpSAV5u
pXQphippHLHmLNUWX7mytEjHnhDbjOwbPiPbal9xRy07saT+aqZS/BsjaiyDDnnf
vgRDy511uGjC02xctQRD6YJtnpf7EprXQz5h0/2dak8uEOGMv3AdqK54SfswvVeA
CQ2KjBqatxUx9j1jZwqhCT6Yc6Ut4Z8FgfiQfbErLe2Lp+egNa4a3Q8SKBB4QRCz
feSnq1+cAMPrgUuTeBAJ4IWagY5k9JPaeFlgI3Tjfp4K+aTAd5LxdEkNxwJulT9Y
T7Am++NNEn2+MiYsvc+j4/L+hkpCMMY9Q9EGo/apheo5P8G2QUqq44ry2vo15MP+
ylmOYlNA+JXRWvkxq1wcVCR+sPeGDb76elS2yKltg2zs7CqyXHEwBxRyrSq5CZIg
UdXsc2XOvsJz3qSY+K2cGqzy+e12nIUu0uheAb0BxFkwH28bmuElHuxJtkrjitU/
iF0cAFY/m6ayWnBntIJm3TRvkeNooetrgJVrhfWJ6aoJBlF99/nYUTNxKol/grjQ
up2AzE1NrqtqPDubbi7stzv+99JLb3qxZ3TcKj4CtRx+kkkI4MTrDPI7/DU1XOh7
1HEyfl1LR5CwNI1NWV02hsYD+64xvSV8Vo+RY6q8iMWYf0tjHnJjc+krFMoneEr0
lNMYkhkcbJvBbXZE8Dm6+38JzTXogi92J0cIpdhShmXY+NEmrwZeEsKFp9tzgaqv
gFsIJpaHPXWfR5NCJWo2S4QgrXS6s3YhpsFcP3JZlHbpG/9wIVF/WoA76+eKwWU+
3mlfovV5/kOE+tWAt5SJRubCmSq2ju2BxevpgINGEMNqL8YqguRuXuIbA2j7OB4g
P880+wFJGUTgwROLoWXrtJWZAMSZvEiMDa9JmvcUzOgecgUFwjCWDyv8mOg2r1zl
y3X/KHpF1mrtBKRw0Q2vhZOPR0Kvate7fQGPU9QTQkB3MPRnjnCFmptDjeQviBeQ
wXlG5kRHv4SsCBWInm0QZd83JcsG6rceiUZq4Dyh9ck1Ihqt9yue7RycZCkzuCH4
4xzDx/MHgYjxdgR6rRlSvFYSEXvcgoy1r3QSBf1W0urlopcBHc+Js4XOuH1SWm78
ltPOOvzfJM8iLhde4LVvyx8ddx1jhomy5aTuoiLnJxkHHYrdopRpWKGdCCL5gHoG
qKmwRIntYPEcdSLzeWf//ytMQ2s1CIzFho2zXENq9sIsZiKhdtOzfgYJ9doysiFu
g86xpTr733w/7QQ9rIsWo7Ba3aFOuf7V9MPHRyu4vBpEkF3rumJ9VtVLkl4XeHxU
emfsh5wQEvUxtZs/aOMEF2jydcQGDhnpW7bNb+PrBrdCVRPcTGnKatIQ5JT5tMJi
gzvyscplwzw1foK610J7QfzjOlhu5nO4EdRqVo5wfmYVAjCToxCIbAbKeCNPpcbh
Sjp2Yk75csDrfaiHTlARKirWhmtOdvFI86Rx0Qd0mMDl/UpSKdL25iPr5AR/okuu
q1pjU32HbyPYhZXKwqIzSNOQHozmgytjauRYQRw64I2gHXK4+7a22TH6WEAQgrIQ
dRotY3nGISxLjVFGXu9vKiXEFzFr39hd0L0/lxc+H4JFVbtHDib7IP0Yt3wa+X+0
MYwUV4bKrVBTxucwlKxbuZO85l0Jjiw3Z3IGAof0tl7hLLn11LoJYnrWPwX0GpGr
Ivw56WKEQWB9UAfXVKa+MMHOaZRqnvYWEEsKUSCAllOaQaUeI+Pg6rbTB6vkc/nj
7hcpTY65ozNlHgPC2GA/AzB0pkrFEVSDAlQzmTvIzEX5f5ck57Du479efh2tBJDy
ZMtPI2QIXj/z7ZimjMC19DdO7vA970F0+eLrnBARwpDbvkBstnPRHlYhTnarT7Gq
QXtribFQVlXFP34NVkjq7vT5weA7yxQ2eBR8qdZqUvLaaYc6ulCuPlMnTGbYiudQ
UzREFUvVxBw2OGx0qffpE025DX8v4TBWIQeACjURPcsAot7tQZXD4uFVrVk7loZv
On0aiV2MctO7D18YO7Ph1BcoPiRoi2KkNOawyfj1nFPyiLRsThPvfAFI7Adk53Mc
KqVtnmb9agsz+kCIrmAlI05XLmg7tlo6FPPPBSCyRLe5JiP5jSjeGXB3WG2MQTZZ
8CqH/gN6j36vHsyeKQu0qo4sjsSxksZO4l/7bEdJtL0ZO8oKr2rkwj2dL7n0T+Tt
MEFweGTnfPmVzvwRtnTLxzr7UK0WcEyvMxKddVyNk/GsMtlfS57ndJvnEEFpN6Yh
AT0m/NDtFbpb988GKi7CSFqIOlptPeu+FXY6tpg6AUhZzyvzG9pH2zpVUbZ/hdwo
/IjykG7kLVQQkteBCodJm+EGlOPg1/gK+NZmEoc+kAfW2V8tgxiQ+9aLqjDLLh7o
oDfW25/YE4feJmPFL3Po4GNZbXRzQg69WbZulNEG3OhTARwg3yXM7DFmooPM1ybC
ZKtmtCNns99Yd9n/tBI581lgmVXqrnonaRX4iV2XUa5B60MZdPIROYKdq5QZn3t3
L8yXyHY84rjEY3ycROBb4a/+0nS0qst6Rqm8zMhv6JYh+dpty/5ashazdgiDPgZi
5eIrd4xEQcXR9vlEFJrxb7YKlyz6YU22LwQkjTFkgxHmPam9Dipjz1RGSE7OSHGf
h91U2L4eq5OYrSLV8ZOOLErcuvJ/4MdGhlStb3Qk7ZTcwdcZcqnH3hsj6UBivJcE
tJ78uNdKfIPOc0kkjQROc2skudIApQAKe0xCuV4a4DAlEWhNPnoaZd7EOYFB1CT6
gp5blE4ghb7PzdlQOTp/3+l72CyqcdEfY6MBhtByxTLeTCGjrOpsVB992E5TfKA4
rM55akdUXE9H0QjS13ETa+VJuIjV7Y/LAcF2Ih7WnAg/ksgLqkPRoXck5k4qI/i9
1U9XczsEK3SnpNVmH7ZPGC7k8l6bQbRLm6x6m2H56ie1xsbaZTwkSs9lwLxMDkP6
2Y+V55kypYWVUwgD0yjpbkmwu4z4s7OW0YUbuREppDSW8jgQRWcSf2XRQ3aTnboX
fjOpp5z6uVFj6Pxcyby59LyCsRrV8LPAWO6Tyo8pAVjkDLAOp3uqSTM0Aqdt+4Wz
WrtP5DfFCjtmoy4IS74ivFNzjGMEpC0RkSoHH262qU2zjGPsMK6U5AYQ19++zsfd
twDgwh8yYh2VasZ+anil+O4oUZF6i3WboGRLrxu4/fgleKPbTOIBLZA9SbT+xVVd
iCqmUeERzZSfmjL/LSKAdLoqYTuEUe4YxgMLnWRjzAC0jpiEZU6cSb5tFPWm4UUY
dpPhpDAwjk7jF5TSkfZhhSWRyqj6LcdeECH1l/mUphTrqIe0AwrDM7qHGiNm0uKj
mpNdg0Y7ZMusAPXmeZnIATWALwsjgWYH+7wlCcfMACpkVhO3wncmSkOra/9ikbRG
lDUzzE52z6+spiq6Cwu79lJuB7KTn1KMXql+uB9Gz1KeB6rrAimPY1YTgG0f1/wV
+hfnhNWlTP1glDaCvDX4ioizL9peOHsKiAper08TGv4YeaHidk2eVxnLRfmFF3J7
x/OQD5yeH7YNf/dv/A8/5XBOOTfM8LY0ECyVjNiJWd6R1xlmDNs8xVXzHjS7SeQj
7uyQGV5/5cB/Ax9451UjBmZ1ADhF3bRkZOaZydlNfNRs098QXFuk9uAV6ocngW1K
G9QvhtyKGaD+qPUJMq3kDMF28g/9qx+axwSvgAOXOd/tZiAePz8ZPW/pmEZftpp3
3xDZVdMq8LCYiOvYJNsorE2ugXJq9RjA3DQovCr/hfXOk/BHdStVQ7w7wULLMJPm
CXcfwP207DyVHHpO5G1Cirm/5Vv7uGhdrN7/5gEVo6gAudsVhyEzbdUtE/wEFhG1
2T8DWx8ZVrJdSvlvclYIZVETuVG7+N/WuBY+5tUHvLMjwx6BiRBFjArAFW/4mkDI
qh3rEdGzPU6V2Glju+Wpj3NvcrTPIXgF4lvQRdF6cCRMhAfRaSnlubK9LWzFRTD+
q69WyJ2Bf7yP6tvZkzCkanfO5geo0eDpSRyEW8Sz1lL+94L8EaiXc4SMYXg7N2Nl
VcFapXTYCaLLxsfhmHWDQ04PsXZNpZDKzJZ7KzjudCCWDnrYabycyXz7kdw/ief2
T2VkAWKvAwkhfTgtKAOznt6+v6FLWqmuBxkNPXk1w/Get5PJ6q+nB0Gy1ZjNpB5D
reWD4gkKnUbLjbxmWgf8+Ho34cf/n/YKnO2QNTpm7lPFoDg8DT1cJM+MzADNS7af
QnR2e4qDbC4Oi0rMTBNp76/sShWNshSYrehbDCByNnRjNVhPlLnFL8BAMbMCRHE3
vplFbpeeGBJBWbFR7G4n7EUJc5pTl1HolaX1DcO9UuFmgO7ibieEySkKZT/j8twv
c0JD9ypzH5piLricTmpeDUgPnvU7Qy60LfEKVpsX/juZWxZGfxVglczGgtsx2aO3
ROPqBHAuTOK+AuDAJsbYYpAabrsdxi+m5NyKIJX5zVom4lTDPZ4rlgs6n6DJkSeA
us+hm3olNY7VGW6iu0lvC1nniQUFZ1bAiYa8KLLbSbj0xbve1I7jRH/baoZdrEoR
Zu4ZNw1BfEyEW6ujQfoP9vLACQYjcWekxLYE+YGS+yU0//U8UIMQ3+EAICWXbJqX
9i+bT2mEEp5Il9mt34symLMzw8vZ9n+9F2oOyxce/KWfoGg1y2qDXHN5DmSxhR9f
mBWBES5joOIt/nTt6w34NO8g+QwuspA2lLEIak4Qzk7dqsv/LEHccEJzk//Gp8R3
4SxVYikJu3PFnrmNX6UmgYWf8QOD86DPsQiqrQE9rlxnPQcJGItb9zvKDmlfn4TR
py9IliiJnByaE/K1dxc2aWkMu0cgwVz/xqJeRVoinZh+kQfvCqWlaRAX3diDrgQ5
abU0/or2pnmNYaKvk/vWhzpDrusXzGiQxapIaXvZ0+AOwmvgSi0Lx9KwMqLwEOH8
L/sEeVuWl3JBKAMr1HiK74hPyDzl99CeSyE+VCrWLNAVCGYPruNt0mbzetgTh/BR
b2MGqj4/wxMxNPRlt5MlrrlXzhx9u3JA6Dk3as8BVQPx+hu7K867ycKtE++VPr2d
B+4UbDp1xJO6r6OCC6cI5W4W4g5ZIeAubHF0yt845NkT5TYo5HEzxAg/xj3kdQpt
N+hwrhaDyh1dFjdXXHiuWjoyOAWaK0FIOonWpDrkp/eq1A5b0UwAwA62vtFb/U7/
JrKYtieJL3oX3A5ni5aJRKUG0uo+EjVVwTs168AzeuQcdhGLMv0CDwNj/ISyvTO/
PpRnISCfGpOrGcldIEwS+0oMMZw7UaWBrRNLjrnUEdAsyQRidqjodaHmzIRMoakj
xvL8S+0Ov2cdLuyq12XaaaBRH6cPeOJPSLPZtvhmyOna08VkLTHr1XMfWOENWaei
T40Bd9iz+A2kEm1PA0VeP9iYo8Y0YXhs/gnLn1FNmChDJUEoaJ1pOnLdIHNspZJ7
oGp/iztPfhB+wIFWzh/Cc9tGYedYskIEPssW/sK7iQ8fb5V/gBNPwss8DKWv/n9N
KQuobr87IcqSmhpw9rfc1Yaa55JPTTpVoLPcQ36DUp1KUXeiQHeew4UNF7z83YIg
NPY1ykfFWnZZ99wxMrA5daT8NxQJDH9YkfEqJgiee8AyPMH71m4N5NIHoInFIjWb
D36zrbwNBB8rI1EP16TdctPmQPJIiFVnT6u51izcvSrXWsO1o+0CkcQtV20JHKxu
AK2oog972Dwnh7hVy2fW3wTtBvuMeMArg8RAFjeIPjZfcfiB6tOI497PrgJBkTZl
VOE/4OKxTSJNHB2WTCQLZSg6RD7/bm3mibFfl4LInFGvjh8ePihImAeo+eU7JhnU
J/7fTEGMuAOVOrMtCTCCqY2HEpC9f5RE2fAVY7HeM8FZ6blgAOSHXjjT+sp+dzXF
hm12EEw5hzwbe5YXQup7o2Lx6bP//Dzb/ZVVfNlZQAKzeVnHqfXxRlVwjiksj870
KuXfJ6SIZKUz7d43/yfURn/ML84DQ0MQfYPU/wz3DAxDRLqaTDh/lS2dY3KLoTvT
npZymGexhlpWZIwBklpNsq4VkGu/0DPfqdmPHW9oNABRwBR0QuBqjZVVrYAbRo/w
hwfWt8RKX6eh6bB4LSYkstgBWdL6VQnp16SDrHDXiZmhqsfh/Ccx5Ki3EWQjF1VE
KmLC5NVcjjWRXt4EtbC9E3Ld3JFzzGvsZGDeLkjwnZPhFbtjDpYaeCcfcVEMCJrm
XJVeMtZsgI9OcIjzAtMOVDGT5/ymxCuAaFejyu/cAex3JoUVF6jh1NF3fgEV2xir
MjXmuhLQZqUErfnWWLsWx8RI5htE0K0fqX8jkaVZzDC5B/XP9sG4YuGLeJNTtpD+
byLEIUkcJzOpmj5/UhuZRE6jPU3L9AlX3jjacuuiIppHRp+Z7l4VWq5KqlbUbzHj
M/XJqo7DGsrbi21wSU/oGFCUk8AtroKc/1E6ERorh/Lfi08/Ld/9QiSoKZK86iUJ
MgliR1JMANuoiYCAaHWPZWWtvBzPKBMd+GyyZTi3oOFMygcqibNqXZvre3tvVnCF
LmQIxMMV3qw6roPmbqE/V0mkCFRn7mCCvZ+1xbTOOAlYMDIyyRIbljoY54oIktcJ
nnzlo5MHafehdYLib/is4on4MfnczY/6G/0YsIydDf+SYX1So5NuWIsIA1DNJ/2W
k9aDGOAPdnunxFYMF+qPcXZ7j0lkoIbbRWXaChTYmV+cYXUjv6Poz3GxByUrJsIk
k7/97sxSIfqc2HTv0V92HDr5veSbR+4aXe2BRBSXa5gz0PnLZ/K79B/VL0sU63p/
pdQ8ScC/GuAntGuKDIALhw9cS1d+9Asheuc+rRQUDKuEjLzhPjom9xrmUg/nSPrJ
9Aj+M77OXiYMI0gTEuFjnkrSHjtLqs30Yj007TfDvjXoNG+Q3ivOrywV0uTb6+B0
ZIErySVTT8DljTCv5+u0XoFN0keds304N0zyZ+sP0ky4ekIawE6NdNtfTp67tkOP
OAgmTdO5RaRhcNQPgWusLjOXQknmunUHaIlHwYcVULrtbXiMOe+qb2F/NsxHulM1
xy1j7ZN36FVE9P0SAu+Wn7Of5mkEEwEgBXPJwP+nZGFV6AQQZyRqYXdJZv2NSOZF
BqeJjG8651xXSFqmRiU427b1ehnYmNuWW1fjewMSed85aJ2aPQI3ao+51DOFxOSs
gG/qB9u52IJRI7pE7ToyAWEPGBHtqrbs0RBDJAaVk+T6Tt6qlP75tGLy2Xi3Uuso
jEaGr1A7+Pjftdi6ej0UPL8BdW5g+abV8gs+wN1cm6CDiW6rTgLfhmw7ImFJXrye
xYNYnuRjv9yMP4uK1szgoxBB1BhN2KvOEErW0WT2miP+m9SMTPi1gMgMEz+Ax1v6
kLBPsVYUZds0hsnLTwLfL04+hAo7TC1/zGwfintvz648eHoNn6KJciyMljR0aXug
+FOVOedNvRQ/xT01GVP1UNyQdjuAe262E/y09g82ehL5iHDox/+YIneeZJz+23/u
kf3zcA1zPw6Sk/6OyiM53T/Jhu3+vpA/63cygtUjk1NLhig2Cuu8KsVAzss447gb
CC7Z5BU53L2z2dwmnFIxcbiQQNYWqI3YnvO4swzFFURejDv+ZbKUlklYqk77YxP2
ms/y2BNoSxtfBbWxZxCvC7kVtjLgtXyHPEKzFrUk3CzNQPNLZG9KYRPy1bR5/q6c
EtKALzxzRRFcn2yWaOZJRN1toUvxWeWqhk4mOGx2HN+t8w9AgED3uRBCXe5XANSL
Z1Yw2qBumwtOyXOp4ejaGZTQ/huzwgbm3pocdLEZMgbeIsdb/tzGPi5G1sgDyoPY
sYbSpWwrvR7BfkWik0d1gGZje3VDMmVTxzr80Xk06UkQrHzYbjxQ2SqrtOQo/9V1
dPpURY4YFcgKjcjwAuqvIxrA+6HxTF4bB8erfscflL2IB+RipTuEWMxQwaPrMUbF
3It6NN61MQdLrY0jUsmnvvFzccdkr6hcTvgW0709UL6NVrtjJL6e1iHZ6hzCbvIe
pyFndhdwUMZNln94EW40CF/kNipFNLjdeouwbT4jS+xEWi9AQyMyvXSb2v5Y0/hC
mlQYYRn2Lssp92eCKjApeWW2fHGY8C3qV3BXKzGtKgURenrw17QFKlyDr3czoVBG
7NXsA8GPHkfnb+APyj+HAzcz/6Qdz/KXP1k/4cDeBZv5vZt6VZElRZ0+R/D2lDzz
aDT9J21aEfDoWTb5C7XzDpHPutXGkxcY4HozudQ+BUgklYsS70MwiNG4iTGcJmFE
cHZaPbsvUqUVCkOcIsoZF4xn/8Xcz21shjdg+Im88sO+vXYx2we2MJqDB2ZLEeSE
M/VQ5MEVVMmr/tFpdWf9ROEUU63cUa8Uy3f5HSffN+qe49PSVy7LeJIQ+vLPbYVK
275ptmtJ2hIrDe2YctpRE9IM9XcDPvbvLmPtfj0T4vK6ChxFDS/Mcx94HDIEGwJN
6N0OXRq3w3rqnBDWQEvjoLGf7xqqccpD9wGrMwsibJ6Tt+gX1YOpfB+qLjlyryI6
grazUESJTD07rrFmjGnFxGNnJNfk3gQJx1Ho/Q4+s2mqPE5XL1SoLxaOQ1JhuJ2E
HiJNxfGSi5p3XBF4Haa5VFHOrihqu0ATrc06RrwZ4zX7kTJyeGbS8SejVma27iZ0
J4NlrIt0kwcmVLoxoY+urXQAmr2PKfgsl2H1IhTwOg9tWOsMKxgGlzs8JHhyeIrQ
Am51w6s96ynEY27YvAzESf+2O+0p3HpnnWfKngXyipN80VZTEhcoYU7wz2Da/6Vx
90euI6R7JlNEmRVF1gPJuzcPXYSty0oBEJHs0f1/82e69ZGyY91RPrwwqWKRdWVQ
/PprUAP8qLv5QHeAF3mwKKaNMc0pNEY17N1Nb03b58cR6so9ICEQRKAMr7CAvw+8
jNrp5LglWVR1hudpWgU/tma1/uULlRf2uW/i49SiBTcoLxTX7TO7G1emhi9XzwmK
xPsPk2LHOv4L9D6v1j4zzPuDkn7BzUc7lfl1dVMUUtmY4DGaRGl1Wluxw3ILF9sL
5EPL9AyUHaMVO2c5CAu+jBVEe0TyJORRTICdh12xy0XHXleFewHlpnu3GaQAxUjW
UFXvim8nRchi3yBG1AKAjRy12D1hi1tg8ocK8Mo/EmejPmGdKv4SBLloaBETRwNx
wVSGlIcnI2DYwH5D+7+Bo0eAY5Mn3vG92Bs9P1UmHyBCqulksSNliSyToNXg3fmw
MRIGG0JINn1RYekjq364YHFNbXHSS3DP34YKRdmjtkeS0E5s3RszMHtQ8sn32dbV
w7NxaTy02GekhXwaSZpARGm2uBugpdUy4oWviEARQqkMRGLF/Q02t4SqZNIyJmSp
xWSy/rMbJfEN6EAlYzcEsv83VPqiwm1XpZlToZd5q3fCcb29NwM2oZ5Di8t02iQu
ljV2CQ3OrFqm9s9DDSFPPE3P8Yq7wX3pnKjfyA7HFP+MzK6MnD30W4Cv71P0P5Ai
OonWEjmXScDS/3wjLjG4tFUYLwm4mZxWDQYhT8JHNXy/GevShZOpSCuiJBzoCRka
ROroPvCP300NtbFJUywc4mqdkfV8+RUOU4iqltoQ2sTZqLR9EX3sIkq22zTicOUx
yoeowxfQdha2YKYJVMt7hFYmcO4iCgtVDmXoyk7LEPmxXFArKnUd/Zbpy489QR8l
1UMaKEdoCM5RYmEhni7Fm+TXQNAyfX3MyvnDVFL85bzX/UoGDHRqoFxIE8soF+8W
gyMODUq3gdSoYJQjlhVgAeQTcNZVkd3xZkhAiAiEtAvLTwUECeAQDr+eaq41OAYp
5TalBqn/LpkMDsWxM/goradSzDdx0JqOp1NSi/ip4J12vyTCFPWExycE9HCdyK84
OXENQc7bw6RWTUjP82+zvyS3bPiPDslT70PFBDtlUaGVM9IUvOj/sTG3NEj85iEy
xczzlIt9ccerGCBqlgrLumfZxndnN6qFRyftklzM7JL5VtJZTb1JXs+TwmT93iwR
wn+4S2CWFIYQTR1DexJsbdTXk4MvXiHgCtDZTnqAzudfRdMtb2N84z3jJP9Lb7XH
xSAsnlwZHs1BuTsrj0umRMrIYkxtgZB0+93b7kwjo42o3hjCie/k/4B7G8Os9tSB
0om5oLXNIziHUcSi3xF1cyg+e9kMDa/OSksVjSspCIkimvnrSBScmCPdoP3emXUu
23kuj/FLZ+8rMWhGvswQ1ztAQxWnmTw1nwAyMQ23gDpAQHtoqKzi5iALxd/oaPU1
bEjhEzwF6NXUZ8B/CxqCDzFJCE6SaqF2aK4SUXn7VF3cSDdU3+NSYRqbKmrRD6Rz
4e5x/N+o+oM2ZSOrbzUnK0o2AD74jMiEYkipc/dZQTlwtBgMqBvZJaGAJUQl1/yu
h4zEpi5/Xydd5FPTArZA8swv9/D/Pt/+Z5SgmpDZdqSraSmzPeET088r0Cu7arMe
kRawavMxJSGGn55ukwrUCsrBqtvohC7/xy3GG164ceGMj8v+tnSvXJAgATZYOm+D
AtEzWw6TDDbSUkK7Q/albaQPu2w6vID6AuFdKb0gf6R9SOAC/YLoxYCNWz7HrJUO
PlhxF/RpkF48EEFQIyBiWb2Ow8XRS8F4k9okj4b373pP8HYl3hVBfa4jAwY7Vm3V
n/a/obbXJJEIogBDQTufIe+cvJoXHEwRUDcQJ4mvnUnqeMNVhGRIHC0RCYiHgMkm
fj/xvxXMKsuWcWo1hfYoDrKdElT1WjGfO6hD5RcrDMksc3+/MIegbWWGowDjQprW
VSxGi3nl05zFTVSBl2MgwVYjTKSjXg9v7udKh41U/cRks6pAYwbqf0zXTRuDsSXo
agrmXMavhExukC6PB8duZ0aQ/ymykiIrxLkV4kZmkCEHnYqz8eGMA5vy9aKei/XR
YAjaFgaocBssBpsG6S6P1UxW2IbC+R3kBscLuRPKX5Z1KLn1DjRHwxwE2fnMhryk
xc7b84GzGg6pcNB71/4/BkkX/ZhjLPxPI5fZeLsVHx3bWegnWxcGfdUZCKRjdhZs
aEXlncDaYa/7YLCgee5TYvlSkCp7VwDU+6G1iju6K7F4dffFB6T2BLB+QXKhzGAF
8p4Ik4UiXuFJCG7TgwMJfhf4an463FTtgx39zyueZAR5IzSVaGTkN6m0J6hpAARq
0hMO+voBOsP6WlLOVCuQBm9055+6N6/f/GgB4s7Uhw+7Mk7v9RnjjjEMoD9azPUf
fI0BcTCuDdL1hNolvJ8qSd9N5IH2ghAg9yqi92s1O/Uu7f6VLQ9yzdxYuzdxmSFO
5XSrZtbyeYMyO0llUusle8YaclDB+E0+jBDYt1pOzSec9aE6OXgsOgvaz3st/RvI
7EqQFbzxXp0Ueh8WELLanwjpx10bx4Hz3eSmqd+pxPCaVRp5/2xUL+3S5J3fTSE3
yPNQrbvP3UfjIS3fbDSoc/ieT+kkZ9PeJkoYg0xJO2oXtV4jFiB00nS0j5hOvcCk
jToqEWhZ243xlF8p3ESSXY2hLQI55jQsMo+HoghXWYe5/zPFrMu8Dpib168PZOs0
aKKD4/bQkxBcLjdkMOeG+q2uK/OygshiSk0CwJ9HGkpu1xuOoUqTs+9R7Fw4+wSx
uJGEORZf+e8bX+PW/G357/5O5mCy69GfphinaE0AWWci132cxyUegbXoGmWDsWH9
Jc1ZenYI7oLkxt8xJMiq/vQJScdwg2aqd8WSeXQlgx46S319P4bvAfHFzjQLFe/V
ddwgfBehlXTZjkDnyxSmQlw3k+y2bwuZjgx976dZ4TJRsDqFKG/eei3sgCvx972W
jiN15MsArFE6uQafVGt98gwyyFZ0JFmElt402+S5lukxID1ABDgxYC5HAF3eSMIm
Q5c0TnmzgrAZfZC1U8DwDsVv8DEeX87q3CU7LF/IFamvXJlH2nrIgLDnyWk9pKFY
QZXO97zGJJrrA3KiOzuR4R2sAWQtyQC6MKLyKzJbxeGDRrGG8+9e9WyraiFzvzM7
I+T6bM2vifwRk2+Ty3qYLwOkftju7th5RhCS+5ap3oOsgAA7/FS1eznCLphIuw14
WJCoebWtqPfFFYPc0bCNEkAQsCtVZktj7hTCbPTWpMlak9b2DjxKvyCvpFbwolme
K5eMG0QWzxoq+6c9p3t5T5oMeRDSvVIpv9/9bQEcYaoAihqeE+CdTf08Lt4O156t
ySXLPoXp+WPJotXyYdv3pSzgNM2WARtEP9wTBQmxnzGiHFZ4dp11tzDVs9Id/Biq
tjkG+lMYSlQ7y8xZuApMgrZgInNCDHfOaz1Q6ZINrqv4n03tV4Y440RJAwdDCx8x
l9lt1Ie0HhgNnpVSTtkCF84CN9cTl1Y9WZM1SimoyTQEa/XClD+HPBjERxqna7jB
ueNXinjOv9haGMVGz9DsgA0ufnB39a4CTB2n1nikmfTYUNYGh233GId3YU2aly9r
qyRvmxIj9lMG9vrWZrfDkb5v8Q93cjh1eJE0VEdLTmqE6wXm30BpeQ51PMRZbVd9
JONyNC05XmOFGTWCvZKyjWUYzjwzciTvYEFSRMAXUplzvKcszt6ECU5T4vsJXUCv
NSnxdz+VG8m4SarjiYkx0cryXFJK1U7uvC5tm6iMr1+OERVu9QQeHwAAnjCN9SmO
KgS+KFuwVY5P+RD/ekDo6F+YpwFmWc0RhsWODXzOi9ZtNShRfSKtA6TmupPZhr4R
DIA+bcnbWYjlTU85FHeT2FsznWPGqjlRma50t+x35kn8pEyVHO01IC/G0avpi5sQ
Y0nlKViSgn/l+BlKKIseAeb1+UoAIf1gMqeHDFureTqQWylq9lTBzL+yPVHORNt/
VEXFMaqJMtTv1DgY0P5WQ3eJQgbQd229eUQikVv9Lc3DRngnVUMG10w7kbTjibas
ynEEZkTHNDnrLCYqCQFjxS5P99j0KG0hMhT+i6UT6xR8jG7+L5Ze31NhbBUv6X+4
i9vOCkHSGi7mHxsSKPLA5g3XPattKVs1aaccpPoCs7xpZykb/qqRXjLpY4+BASrE
Ib6/4BG5JVntETb8SuCf0JT5VlVujLDxs0+rgApLvWkiuGTYMwCb6Sw16oT/2185
sPIVIYcMoHhhsYlgZ5zFBs6ipQSWseHjuD4X6SH+G9JsOQ3PHFyPu1AVxAkXjaLU
GpxSiGKdxAnD7O6nq3RZPTWhnCcsxk2mzPrJ8NWW5wUIZ00wEfTiRusMyyuWH8cn
CtVMB2rsEOu2V1Sqic7YY3NYH70m6MhijeWg3Q3xpdRYpvTKZwizSNSZenlPnPAc
8vs+1oQgwoojw75EHrmbCDT4eqyC1usdyR4q1JZcS+QnRmKECQ2JqXueuIp9oHcC
ZjR4opfI1ipHtqvmcM//U/1O0yTgUC+zJkWsbt0MVR+h5bBwPori9/ymZe/hepWB
FTeiymov0TmkC4nubq7kMoAvv6evib73FMOnUCQ2pcntiOskYzqQzJZ8fDsvYBoD
gJgKM+u/qpo3DcArkGs9loRWF2ZuS91AmldGUAFKLZUVJOdBUFJqnhfBmjcOzwXm
zEmENtJS8vP6AmvX3iPnk7+rC1wy/LPUli/NPQbZbNoeRhPrtlPsINI92oYEdsSR
zWLqo+Nf6Ql9TUkfPnhqaVttcYVeLaqnHFGQW5oWjjFuEyzns35Kkatmu2qyVxWX
aTV//Z5F2YzVf1p03s0raokEiR0TdtdtU3yMPCFAljAHEn9c6K/qzkBk0GcNt5IM
TNf4SBo5CwE6nyoifhHZL3AffdlTDg+KZknM+6rcJLEFc+NeNZqr3dYvIg8L3Hwk
EC46Cxr97wDdJGNGV4kiwfuFmehiGBAD8U8dCyeFidCmz2WGo1ocGeqUMtvymkRf
PtSY9APlEYJa5ilbdTero5Yc0au8eEEWDeLKen5aBnCm/NHZBASSCTumMsPpKs4E
Fde1CC50IP18BfMSm2zIM7U+9ldCRdNKgKkwRQ3xd4Gz1vY2ssQX7LPNBGC2Lplt
seSdOLFg630beuBBo1tTROdYJLy4TME9wMjJpS3XOGRda1INfO26ON1SSUGfke8x
mgIf1hH+eN+qU/iQjUDqglVr1m3i5u/vplwuvZHfuDwTbb/wTJwYVfA2YXFkuFFN
0Oi7HstY/9nTTkVSDNDDOag3lCiUB5+v3IEPRW+PtL8e4B2gS1GYWBDjAXdGW3aj
+UPQc+LEhTEF1ylBqRTmGOYM/RvWI+3dcfs2BaDGTnjzCVG+1KtuLWjZozki/ZPq
QzhhKVsFPDZwH5YZsYwkrfi6x5V/zU35IfX/xaN7OpIoqmX1zI4OvW8aHNtem5NY
hyLZqqiugkyNtzb7Sj5XOVVnbqa8GEfwCO6cVCmh690+eYrasZH2Rmax69STpV0g
F2RcHtdGZwehU5kW+mbCCBXkXVpjmt/9WXkVIPW2smS0Pnz5GxQsCxcPTMQ58ueD
XubxX1qPZSjDDMXSwJQ9MjMM5WqCb9y5XIAggEmlfQcvpXar9+GdFVlUutYVOGPY
Fi1wEHJMIw28htEvgDR5SmLIynX3xRnW+Agn8iWC4YpdOAYkgcjcClOEbrd+gVAP
6NRcHZ8EwryIaQ4QyYr85xOcWb5t0/77Y33Ldsr/Fz4Qc9ZEfn4j7/cvayEtldBB
d9Vi0zC8H/zbsQ6Dz2Pm24ODs24TKKROCPC9sTvVdvrWCpfZnc/R0ApTyWx4v2Hq
wv0JOeRXa1E1Xn6s/O1ufvHJ8Hc5B8uTZtQPCtKy17dnrSnzKoFKnDnM1cmoSyfS
PEDDKPpg++xkK7WPjQHmAc+ln7uSh9wOLZJhLWUqx6l0IbcwrLw17qd0DP6bD8aH
fU2yxgrXIc1KdBCPS08m9Eg7GsmOvTLmlzGaWOB8rHrADBnfEPDyQLRh8N6aImFs
pFo6XeT2HiRDDzoKGEBWWTIpW1Uf9mMVP3PKDhZgj5pkyenS7iHZWUadVtNRGX6T
zQ0y+un617iWft3U1jTc125j9sM7Xz+Ch3IVoXCszd9kGlj8PhWWJvqPrNKmkOZ2
kburyTzHu8AUM6N0MIxzi6nhbLWTPk3YmNvZoV1U3Y0iWxpTZ+kAknGNnZkdjXG6
fqKOb+cI3lptteKt7lDAeWGiUEMZrSWoA4yRPxKgA6yu0ciO1X6C6E6ook9UFAVB
vaaQyJGlaalYxsFRpkm+NyNpHTm/9RxIcbPY8ijpKRtNl0gl87/3QnyeEAmjLIJ+
IYqOTpM7rm+B3wnAN9VvQhziK3UXk581scIU1OEHsA7wGR9VktGv9JwWzcEtPALT
1I7UDnOR185dHIbRgtvUa3qjC2dOiTy/GF2OPmcWaq7uncP9BUr39ocVZDHGBBll
c+y+UJqah0GNQDK5iemiHqdefQFdJWCSHeDXwsUGHTGyXWA+85GCxbzEJVaQeEgY
mdzPpzDklghFt8AzkkkLd6jIAc4rgPOpWebMmHG0V8bZ6gkFHMidLHyYUppRGPTU
Y+hpBJ89fsz7sGheCk5y9zH81nE4Yv0JrVlxBeVYkMzyyyLbC5Q/JsMkrnjYxl39
2De1Q2wvbt42NDezQtXaT4tRhTUsVcvBnms186O7hNJcG5zNgxL3T2spAD0BZc88
ZEW0vlgt0r2dmnADKen0fIPuBIh0Ud+XKop3FzKgTyPRAv42lbPtsDYp+Oo26qOq
/VQiInNnnseT4YY5iVyxc3sVERepX/FQii24J5MFdMvQOGwWTWG3ftnR6EVNo+8H
I5ZzhrQZw5KOWyg07AydfEDy6jnm1ickOAC9A1RfB8czWz0wm+7NB2fP+kHHwp60
dtYKjfQFxQKjGw7RJjLMy/fYRiUyffQtFqmIXId8BXHeX/L0HYI3Xy2lyXPwIF16
dPQyIE8sq+c4tFuTwL4BlkpYJNuG302WnOgu5r3H/BhY1oBy/D7N57EQ9AQYP3ap
YXnTQTUjV23T7/j67e3DNUWtKogUM/JRmRIxs7+MEK98lTgG9/Uiyf6p1zM7hC6N
D+3YqkC7KjMKyFIUTsYkisyZm60zvyIybkd5VCfEH9DA6ANniKyD3bitI8RtQLWc
nFZz2PTdkRZ5Lq2JE0zo5t70bB5tVHHuxoQdfz/+OyoOGhJpxdG/s+AcQ8I7GUvU
Pvwbr4jC4U8lmgjFfExeKoiLCHZ4puGuQ4ZkVM5PLuSxcq6cMmzLaVSKSEGfvvNv
n9yWlC1/seTfPoHSo8QN7pvWw8/qrPSPM2B9S7XD0+gw1PAPmlFWVZwvy2G/JQ61
VqQLJwEYBKq4f4FWG0NnYxlzGwxuJtEASW4Cj3B43bRO8KCW5mfn6omCrsIPafp1
/0pLOkR7MwbIZFSWLVdgrPCKoLnHmwTy3noCIaA6vBiHsjWvvJ7py6BPe7IqG54q
2jWA4rn+eE1s9pIk7xMm2ZHWPFUgnW4JcJkXfSLUftgFlV76ugb7SC2XZ4nA3O8W
E9HaosT3OeFPDKcNIrK8hmpbkJvRQpusCSeFh/0rt5PLhDSMMZTN9lMV2X3wnG2z
Kov+rWYNqjufZPWwksFuHMSguRZ8+/pz629Qxj+D/KYFZEPn4UpVEI749+6WvV3t
nk46dlD6vAnwvwN/u0HyoaJ63GiOymrVTQj3IOtXdcsT7DJwxJsEVcoqDEgjujCT
VF8D1TgwMERh1jZ0C1Nm1EjmWuIYgy4K9LIxN26CUtp5ky1oBzVyxgbIX+nCT/0a
GQlhh9T6030YgLIQh13tEefxNtoofhqMjS8LmYPMW3zVnhXbbjDj1FbmmGSW3vXX
TZl9oQ09cohYvCyskuH6HBKHxp9uZJtlrvb0YIcT2AjUJ3vsDeXPYKrsnXHt/xJJ
QQptJcV45TCFYYf5Hi1a3LqR+oxcpzmRCLZtYGb6P+G91KzA6TrmfdxJ/cEJaY0f
i5Fd+7hdl9/9PHucVvqv2IPUQdKqwlRUBHVNXzMojbyF2im+Owf5g837Xu4PbGuY
Ee4CrEG3kZCFuv4nF4rch6RKYARw49ql5PGxVeM9YxDYIaeuqFAtWc7GTmla/oXX
xXitEylRh6R7ppmINq09o/CMkwj6w1TQm+RRUJwzmbBZb8FCK/kCQmPQCXpVnRtL
8VUwKBvf6axi0SDNuHuWPs2Zkw+FI4s+tPhR2UrL5NE5liyc2/OWDbYKZBlyxmUP
OklwbO6ahfvUXG2SxVXx66iSgSwlKGLN8Z3lbF6DzW9y6psVgeREi1PQFwkkfH+5
hh/4XiKXD2ZVy8/zyIsbAQJj+Ea8jixPjRUAaqVT5H7N5vxcJZqWp+PTwCDvrXGO
P5xaYqt40QXCDxmrAFHYBa10kn63HAHIIpDIfspVn8RyraZrdFgqd/j8+xylQtXo
j8VRs1nbiI8bqAOTZmMPiEmwwuVvi+TpEs0xtQgNK166wbm8chIcM2W165U3oY6Y
i6XFnV6fOTRFC1sMSCCTq6Mn1l2kvGT2wbSEMa1FurvwWh3n+tKwb0+JQE+mf2eQ
COUd6YTU2InSUrKrLrzdK6mFU/XrR6Mil90/bEmbSdPd6AuHOiJvSWb1LxV6Pz2Z
VYpJO4pOT7WeftL8JYKsUwMBiRNZzJbKQk032XRfJKNW/eUmfMDGeJN37kqa3Hy9
+oZItMNDYpwa+MSENWIgThMdY6MHNDwrbcaQpY3LD5qDeGGzl5E/3CVBf6iSxG7m
DUD65FQbTACKK/eB+NBJtkQiYjjEu0N0tRLgkuAO4X1wy2bhFU1qAPyTRXxRwT4p
vF+UJeV8YmNaT2lz1XQoeWiccBmaMMfJLlH4DRWFPOy0k1Ca5WlvImNEHY/Ucw1j
56mYi4YaOFr+AHUX7APfOhrBBFfu6yJdWkND1U/6lXcwtWqnBVCdwfSjGjFQ+75q
YwAdl7meyOdTRngYhdf4CClRdvdaDxwPQ8GXU0mkGx4ws9qQQnflZ2G7C1xPKM/k
MUXdQw5pfJDWI8MD4yKSO0Is0bXU02Hj7cVF/4uxIHcGNhgUTH4L3y+mn9dboUL8
bOqVL4YEe516FMVzZKTk83CY/5TWaUwACX/1efH3GRwDVKqrxyuBHdMtF6RRw4I7
cZf5BbynZWPGI39VmLSvverrjRYJwoQY1a2IjVgYeKAQQUaAuOyC9c4PxavqhqkX
axCaBydToLCGSRVkGRiq7a/erY8KFIIsX3GHuxOFOHIKpivwsxFEDHoqqr0A4b4I
GaX51qtD/ztH9QPlbz0ia5yZ27ULtrKN4zCsWVtWMTTWxoCYST1/hvWK9ViF7UoL
OuNsNP5Or8JymmGOt/TVHIhmk1pm75haGaXi/QVsMU7H+8SpN/MhMcaMiVoPydA7
azFqHlwNEh+DXFXK94SbGlqixb/Rw0MEHbUUo6n5AN0+kPTT1Tke7Nq+AUrEhyI6
FgzARIu1u/qJOD1cWuyFieT5Y2Oh3+dPWzxlS18VLwsQP258AJ12u9l9pc0Ur3I5
GlWZ3KDlJMgZEiSKTyLeSYQM7X4PMyKX6H69N1knVx4U9Z/es1BBJk4lXQsNsOD7
5Gsm0hC9Teoaz7kV0lX8PR7j+shgFNHVeDWQqtmuYz+3ldIJwM66LKDhuZ+URZ9c
4BCJSZNhTTw2eEGCqNTIdBtuRmukUcwMQR9gL+1R4DGp3BABpqNj44rN8sLTyLwt
mVljCwfrVaGHJ0fBAO8Pb8nb/USzAfYSYLYolniFB3OyUS/2br6bzqjJGZJP0Tio
UCEy6M4UgAw/wAvqeiHwpB2QebJPVT/fG4MEUfpeRHMoMHV1HudHkcj06aP5OoTh
TdsPgZ8sZkx/kn6W9nWwrm2X8pkkSrXETSDJgOI4gQomNwgLB1O9lPZaq7FfhAbR
u8iUSiPXboPYhXK6MLdu2QFx1oMg1jFJ5bpEMOrtXK1GR3+Gm4mWCEQFtSM2SxiQ
ZV63Bw15ub5RUwsYpkBiyHYYHdZjZe4e8iPKz36qwJbe+tep0EstSFQNST9/aVg+
JBdaThJops3Q/UT9P0VgqVdBwYBGluj2BQEsgZ3raVPPjvPSBqT6maK4N71hW6bB
9KpafVo5/4dUAIJ12/OE5a8eHP6bOtF3BaD0OPVJN/pas9xawlUl7/1+mpkUXkQ5
VzascgfbubnzkeKcutYKAwJ5D1c0P0/2l9jpV6cJnRetDgrtQF+JvFghWpyCwDHF
nrQrOTCCmkqke51MwiQOSzQ63SH2EGeGJeDUPQa9U+IQb3DTrXsYNc9JLkUl+WWR
LLzoXFSBW8cS15fFeKjg4jWOBRXq+akAgIrv9KiS+W+3xZzd/IoVy/3z9P9peU5z
zM07bLNAEBakWa72eG/nWvWPsLaIyeh47cGUezHYLJwJkZXHviU+iWqdmvaA0uDe
7XjMUsjtMe0B33FwU98dIWCBqA5N/UxqyPAFwI8KRrE3tyzO8ZDuyEvt9xupK/7F
80RA7Pd4sln+7kTdTHy5ga0xepDUthX6JyBVN48kJbDmKb7CB0HJwH+0jcIupeEt
J3xnMCeyzj0JXqlRUbPdHEVcbFzXuyxCp9djWgaHPSawH9sGJP9HU06BvcsEtbDR
+4PJRftPxXorBPQLH8UHmK/IoiJ3cKuAC/dN5wvEUlvEBh6J0WNzrXkp//coPJya
A0qaOd4VrzNuuYYtboKdRx4FCjwUs7UEh3NMMxUq6Cedx8d4Kzw7MtB3YOibX1BV
u7MmJgqX1c67EsXzZ2Y4agMFhIxBMnb5I34A4VFN1p17Vo2gZ+DNKiasLMT7rmmu
/D7vs1ubreWsfn/5T3lNze3kD9yvENmUVlTiHTQMldM/x2tJeUhKljEVT9mqwa1L
Qw5cg2T8l089P8kjlFc5G4L+3A1o+qx9iGC5VcugxpfIYM/MOzu0YSKxnO+IZEJ3
zB3cvXK/Ix3+2gH9gn0MNslL4H4cEt61wYrYYLYA4RbCremMb9btMuOG1DShnkJv
MpQ/vfEiyCYQG4fz8SD3G09CNwEM8S5t4YCTwO9hxfMHp4BxqG4EZx3uUdfy1Zok
W5JOdaoqoHGMKhGHHXhoINmOcyMv2JkKJ+cwTNThIgBMTxpTdUFhZ7WI9+uTmlZJ
/MKj6+a1xS5L2nnd1XjAW2fDfYw/CIeoUbHvQp6Rh5wqxbBZNhIn0ueXekCUItjc
9T6HNUIPMuDlcqcaGtUdtWiL8tn5EOG14bAV+qp6D60/Kxit48m67+yyu+/M88du
5ziPp5SuCH+/NL1iunzARVGPR5LsT+He9BG6oTMW9rDcl/K+KLUQzJSpOmXTozrS
CkjZXXx7RYaX7YhlPLZmNa5XqA8yR8+0aGYKM6Z2QXSClISAA8B8orETtipo0pqn
dag++qhsdisVHdFVS9z1WBvRxQymlI/yRonWe8xK9CO+kvuWRIdL8S2UeQ3QVFc1
Oe3pd5gAqapAIdAAS3mI4XzJp3CBkn2rSiZMev8xm7B3DqFK6afAAe3snOsFxktu
l0ujEdyJB8wbzbjXt99+h2So1LxEDuiSzg17uGnkZbNf9vzKPCclQe8VSGGi9V+D
iqrazoEQM50Fgg0U8Zq5ZqJOASwkIyZxVUf6GOUTN43xPqzJRKjJPhWgDApL4MDn
v4hFOxJFBXCmJR/BQDfFljHmFUDVQTxLaUfAbwSEeVlkGCw44B0ElygJqk155l2E
hO4VVhMmbl4LuVunk0nVDUrTqaXtWGuUo4xVsBAypLrNNeS/ONJCLGL4K6HdFPAL
qjNXacifwjb54fQwAer5uTpwLISxFnUBq8UpAeMsRFCRwQS108yNcm0GgRlKFguJ
TzyqnwF3RjiVr2H2Vey3+EPKOXzE22dCNhb+Zdc+Gm2LGhHMAs6gipWhNJQz0Fwl
V7SJCLM5/IzFlEKh04mXTpAS91QM+h7N2CAYzLwrkfLoXskSJ+qAy/AndkhZG941
vcjCshZgweFheqceRtV8VRV0mP7BAKSJAJoVRCJD1L/tzGnkShDW0NteSjZxBunB
UY/RfEG2mSvO27Qe10j0Kq3bDS72r7YfK459xBV2WhK7cTNXkhlVqmGbTwwhLxiA
/WhZN3MryMopZt0nNVM65/SQshNMN8FsoZl8ENpgP9199b41cR++QJVme06jEga9
ke6xdAHwX+moyWe51swHlTUscG4/JQ7REE+V1pITezFaUOKFJUt89PF43D1+CLSs
bHMU3W1GEdfziRx3M9BU5hAaEgOBWS2KfOQUpcCJXNLIzFS0pX5kGDRdrhUJVO94
eHT5qzd49dEqZ4EmbrWA9srSO9mX14HwdUEWVmn9q8Jnz3NYavY6r/h4Sfw1BA5G
Gevs7Irtu43NgtWU2/nKW8F3zvTWXmD1CqsaKjsl1XXF2+CPvDjy6AMsjD61Avm2
Vgfj+4u6tm2coF7sWyXJVqFXQC2MCwe5sveVJNTklKFHGomCrX1/wyvIrZlt4Gy8
RXvmeE3ST1CC8NHn8UgT09jqm94m+vp57QvB8pbUzWhoa0P0npeqs94ECYt6iHX0
mUynSRpDn1wlhNbdqbGl+s8UbqCktN61yV5xg87WYjSfxGZCdUYycKoU7wyxaQpz
f11KLt5xLBz3WpRZ8xGfL037Eahf5UYNeis1npsVt1p1BoRnZ1xANtjaAwgWD2/y
FgfK3FQkwSuulVkrkjhOEEs4IpHjVbuq9q1n8IaYvsadMWeDJk9MGsrqtaneFfj0
dG1oyS7qx7EDwPbM0xRSrQfNC75+nUpODyBMI6953i/fM3vkvkTmaih3DjMd4e1v
6RRekGJCs6HGHARmO1xEKStU2uIl9JKt6w9gBhZjKoSkYRpjNtNsIbliDgjRRBXn
6J6B9W0r54abwn3QADwCVvzlIDlD56uomJFY+C1GfkooDaVRqxYUK+ATT53r+kI/
0n1R6Z6bQ+nk7s5uCGkuGmQwc2us3+vzG92+CU6sva3SitLJCtaEOa698bVYgrm9
WTRRQkz7ViQ5SyhB1TGLlbkf2MrJhRi9R71L00jQDp/AB+PFDBDSTprN56XFoYdU
OYssB4xzadUIas9EpkF2lT793Jg6c7rNndvA5Kv2jXd/EIWn6iNiWUAESVJRGdja
f85wzDG06l3LFd1OJAtUG7LIyPaWMaR7eTyXi85OIHZ+sn5uIC+xTPI9DtIsjFln
wf0lWT45vQSG7O4yMBKh8ciu9h4rrobleGloszZhhA5xFtb3Zd8LsaUqALTocjnp
h1lozPa0mLutXR05JJw7VWKdyQifaDpxF1Bu4ZGL6U8oUuVUpAf6M89/F5FRc4nL
te/mtKmHLzbm5pI9XGCzTznntTYgrsKZUh+H5ARjJ7pg7X5YNdASxL2GTRjqqaok
WC2NxaxOrTU3Q8BlP7Acvk3FYbU5neHR0816vzdcGxnGDtPdigsLkYYOjeTRioI1
0dYoZdoJ6Yv/KOeOZ/xVAXRjd7F2QqaL3IpeDvqVdKrB0zRsx/Y3LM4Y7/VMmCap
Kkxvxn7qB6FdZc13RjIrApWPgO5bxE+AdX3PlNaTj0CQpHQNbcChAzQs2SKPZ9Oi
I9vVnd9GIlPCL8+eKr8C/ZDynoZUbjxmOY9KI19KkIqcacMAbLS0oCQl2Tk5a1Sc
r5gjORmvcHYOLqB98ctas5QY+PCtAfCBj5z3/95X5CpC+QtB1b0vQyagvyEpQ/Ox
jxp5+3zPh2RsNqtSHywyymcAcqQUEIeeIVhET0+kir25niyz1fptK7/PrKPC2YKO
GCvi4Rh2xW35D7nn9GDd1lqJoOYrQFsnV0g0F4XLYMpdOWcz/mnmfVVPPrEVfVSN
lIDUQSQlKO6z+Kbb0E4rSGy/Yn11PZwIBxNHgpB0AUbzVItO7huoSOBZEyrwyO3L
5OrzS1pgKF6/s8oRNXADsa77sN+fujKkyIAAAb1xM0naNRe1t7aYSb2RXGNS5shn
Eun0Y54nEthauUjswAn3qOsStPTNgg+3chxrJrqgjo3uAqvOt49oHkFv7EV0NN6r
JxVq7Zpn+8nNz8RkE+QrCWRTKNK4KyuvkwuQ6nCs75JyiOvtnTYqUeIGSS76wnXi
Ke1gURn2csHdAmYiTdpuFxrLqwdu0fUHqCLljNIQyV2RQOGci6Twk8SjpIWNDKIX
DqagIpt9QPLd0RQSHbdjJX7xkJoxpuJ5VlmN0Ww9xByff+NNZ/ZYE/6JLZF4RZg3
p2BDZR2fNSl0HxNjqZMbdLMSDpYcuA/4wn+kcKTr8QeLyY1bG39EdT8vm6BBuO81
VSiGSjG5Y9YoBCYi4qkT31LaGEp4kfEGO6R3hc7z8EgGby0hMU3A2VdMh20oMfhR
A540gSHQ/x/gRBR0RUcJfdyls/6I2c0kK84p46+T/1jbZnnWCgyDJW+9r2/4ztOQ
JzJC+b44bhm51YzDQejo9xY7NSDsyebbVZGurucnFg1y1yIyCTwgb4OMTWCG+jbl
gw0uqXSt4sXny6Co0G14HEkNTCfK13eepxBezsDuLhVuUffXKwVh77YaC/NhddDi
c/4V2wwhuCO4qn30rTwfoyUzpYuQDLBKFOl9jzxSnvUdNzYnvDmlQ94jj+pHx3Xy
JB/uwOR2GlHLPTylmbPOo9hx+T/D0zim2YPAK8bhwwYPF+9CFSKMfvKhgb6X3z/Y
KbdJf+VBpMfqtlUQzMvVDH5yuaEla/xa88dOVG+HTN9sZ2eFNHo5WAlMKiy2zTVP
kbgNRVmz16l6mkaF7CcC853GbaOWOGM+Sd+CIhQBCl70e0pmFHZppND2ZlWG+MsE
8XmEGq5o7sw9/U4iwiUcAzAK8zRHUoyg1PZaRfZ7wdSiTWhZq+Umn0pkAuNn2856
U9Dd/O4LaJHsjKI0Jts3Dd76ciYVDCKr5wrOtHUuqmdUZ0prGeGt2mIB/xPlfXzB
y8vhjuXgb61CirCuPQfu9FSLlMn35MMSkMUFVxfwcC0zdRyWpz+OJM/SXrhRRsJ3
/dKcy1OrpG8+3h7hIStMCP2nnL59SnDYFh75O/p+d+WDh1myFn+uZbV38uOUhwLJ
yH9QA9HGafSlLnLEHzPzBUxx4tjUnFwIE+vdzE0tR/KmprZiptObE6Ol4SvE4r85
QPLNmqwycM2zR+/bCFhrs2jvTkAFNKvNCpeDQUV4SLJrlgoXMi5W0Tc0QPsq5JnX
O4/at560ES02HJo5PEY8i8TYJUPwnkk+27E77dEtu4CLvfzyenoalxseAJc3dUzg
XZjrHsgacfw/vwqjoyc0CJCLVJXkSBRdk+naYpj+fCqteTZYFRFp3RQGLBXIVlZZ
IC+rFRokn45Pc5nc8sIyAlKTEo1x/4rawv/zsm9TbN3dtbCcBiQZi0HVpW7sH/yY
gwfQmXtJFjWGc2VLsOnSTg234mzFrmSaexhvJxMHgVTTbc5NRMmqkO9snPb6uk5W
rrmSRHHnmjzML/02C++qmKyaK0Pf+L/mPFcQNcHITbSlmScD9Qna3NToaKHHq0UF
Fe3QScvyGzSuXNZBh2wl7NtGEbAl8MuZ39CVx3VnOie/pZxBKZfvmKtSGPyY0GE/
vaLK/3NCr730x+lMchM/jAoFclcnY1nkQR2pwQoivqModFJaM0OreDTHgmfbBK0G
QGJ7GH3DWGx/btOOGJkABF8Ve6dNVb6B49RQWdGbyML7pt9PSfYIf8PlcI/faHB0
5IPOTaf73PsGOjk4rP9/viul9J2JcDH6qnOnmsCA58ODCtKPvlNCrjhFGmYPHa8n
4ohZUn6swByxjQ2+vvbYoFjZNIoJMLgrC01Tt9PUPbuoK1JzRlZ1z53WitBi/kNP
oNNyBpLPx7uRKBFZM3NebGa6dHO31EBaPt+Rw7zngdELYDLgN9GkHmazjYCXADl+
cShco/kUVmgWH9b/+kkgvmVKl40DfcQC5Ax1jVSaMtu83XqFLyISqrvrR5HI+76e
czv51ZKwi+PcDNknR9fQH842rF93Lht7Oyt/hphmo1Rfv+//WctCrnHPBpJm28qg
JVt4mZ3TMrG2f/9VCrZ2ozzmmsEVmmYkfhUqn1eR1w4uU4vclN1uHP9Cdx/mq3yx
LPNpGJdoSucBJoQNcv4MxYOB578Iqu4Gw8IQ/f2BG7snSJsNFLkUg9uAjIyb5M3d
deyjuyh+8HaXhsChU2d/OKGOb2zjLOEPQND1VlNSqkOuuUG7bZeKy31DU7vE0X18
0jffBbQwBcZliswleLnvCyoMPT9cwJcJ06Xon/CVi/UTCS5GeaKUxbWde4gRrxE1
wBcsTAhjvDq6wa00hTxC3LuMbyHmiB+dxyk3BJ1oDoZn+lWM2yE4RqxHisJgOPvj
wS28IgpNRxMD6TzfCRti93tGe0V3dKoDEZoMYIx0uUNkRdamtmQFHg/qJPy2DA6I
SsiWR1vxdHGSP+/s42r8wbGR9q1AsID8D8o7TYQidnQvIYmE6TVerqkFlZ40eNYM
1qIUyMwRRzQ5vEjWhKqLJgt295AdWPCwIpOdP002jhA98HrSy08zZ+7dRDmgQ5s9
rnW21G8mCwPYrvhi3vfPK2wnVAthF0dTrvSs78saNhVcYf19HzQHzdJJa44f/yUh
EmgEJQNOS4cW5j7zOXrTPDTfJ2i8O2hMG9/5swb1IWa8wJtCdrpbjWFNfzIc1k0Z
sE3C2r9sbD57ljyJvd5YNqxNjq9AQuzZjVbnoHVtMjhGwxGy52V9Yd1PRHBmBCXZ
L+hYzN8IO2dfoHGgm6j+IRhLiQjRb1y1Q2nCrE4fv/0HxbABYxwEH/bvsot2nYUr
2aBHFpfiDdVeoTKmlqyDPH6JrnAckgmvbl9scbJybDlXG2oNK3Uklrv5rTzOLC3+
cF7MwacSPcqSKzrKKKUJwSWL2eLLzGUVVtgqvbdDpZSJbWMNMa0fBoJ1cCNDLx4u
d7HkYB3MZRmzvBW+mzbIvoaIfidSqH2mpZ/3ZbhB3Aht53Rd+PZI8nUIUlQmotO4
DfwaPRCFbS5obfsquRYPhUaO2OvKKudZeVlKoCsm83orTjjh1kJ6O42SKwkXF6L3
3iecbcxk6y0fBWHXQbU65WU+tCsO+e40IX0329JIHZ1ZWyayIrz1RDiaoHTv3jg0
XW8TGBZtk9hoffUjyjZUCFlOsw6KHy6urwskIBzkeXC7zXYAjJFYS/WSXO/di/YW
Wb4UdKVz+9gl/0/moUJF9QdakXoebrcJp1xjsVbAyUMtdVvjj/aY7pCmWHb13+tJ
DwyY7qaV20Hb3/mM3DVhXdft6ZR/Z065XsMC1ml5KzQF8hcQAWV+aaCG3NCdnCxb
Xgkk7hSUz61NGF20uR6IyOwkYdh4mb1qfvbgz9q0ijT6GvVWsHdUynRh70bvJlMK
PUSjHH9y4RhjRUS0xrzPRl+MHHFd8mFSm02TH/pHe/GOTdawtoHwZzrqIWY/YU35
O9pyaxS2bGFHmcB5ZMW9Wg4oK2/kXlqHvxbGgar+HVZTOmum/qPP5Hh/fNZW594T
w2zBeTbVTybiJGvYia/6RDBbHBcOHgJSkuiLqbJhRqo7d3KgyMWnPSsXq6HaRmzJ
0k5tr01c7wC/+EonREHrIeovTFjpGwlEz2tmrWLxNHcVff1nrWjUyAfOxClTPdVQ
8EB6cFUfE3BGYrqhPm2cS2QhovieCmYDvy4Fz75MKXbLyzvLSLD5tW7kmq0oZ3V6
CHTBRSYsKbfLKwFMnjTFDU8e+rgNkwB2E0ZtCCV+vk9UdEEZU2GXH9y9e4aXtnJP
Esh8kImcQ/rP6r0lD7ma6Ov/dtjcNiXaU3xISr8iLX1ek+IlKafCjzSIFvh9jl20
job4/AbTvfQuX5qfuY+3QpRayKd0oaiLnhKHvwg1j6oi7IEk5rUCvkelCUtDOq9r
MaNmwP+K7iuXzElI5CNjkf54UWCPtao1BLSYhANwbjkWGeuDxsoMBVBBiuucepAo
E0GjOgxQ9jvr87zIS67H2EGlidEymh9Bct06g4Z/HBn7PnDnYLedFaMYf0zPhpmk
Joy+hv6HUhbas6r+2tU/7tAVS90Q3lm2pAl5tbrN6gJSwIFz+lZyUZrOg1+PLx9M
Qj6dvZS7++HCwAH2//EAaMJoVr9CrGtKOHNjnRQkGw/fTgrUh+oEm3F+OX9kZlfy
FkMP95evf5w8e7AapvNgaRi76S4J2T/4zBokndGKU/PHWOs8LE3amzp0hF0HumCQ
zfUqJuo5C7+7kE4DTfnX6zuJQv1CAldW4rxBfSJWIX61aizltrHhZJb5Ryem6SS1
vyTLMKqwWOrzjuAAKYK8XCMtyS43SVepaD33u3PZvthOG7raF+DfdaxxuWKXg3qF
HVZDTpTq9wohJzwxm2MVZ08Gbmpp7NDs+mMZkIHTJyTbzcQ7PGP8d/tqzHie8jEc
Jl+IKkmitfr+uwj9QA0VA5ZGl6UGQqIlIeZMvnYRNMqfu191EFYZrbKzkHWAd8Ng
NptdPPiobDRMvZIxbHs3MMwT303zgkHfanrrxKnHh3UaoCnfULWkRfW9o8ZWDtMR
CFE77lst6sVYypALtZFzxv1FVCzsz33yUya5wGcGvoYTTRH4CyYctoeba3MPgKpZ
ngieM0soPx6DgSy7cESXEQ4cytTEOxrU3rbZpcePxZ2ZMBLL05rTTvifhbyOCjt5
fn/FhcND/xDv5SgWPIx83JIoh75LNFnaryhX41xVkdDWmQZeVqHw4SnFAyyDdy6+
yhzCN0p9005hv7z2jNivCr+1zNmI52Cw67gz2iCoKdjO24Mx0UwoCL9lUbyNvpEP
qMUcDV82waijsuGarCZosTvPOJTZj6SLGVkEBQzPgXEZRzzTarPEIyEv+soeGHv6
xWBieerIxBI1IAEXEwfaHBlp19yQ2FA18vcNlGubGYuGxCuivfHeL7KN/DlfdT8b
ZRbOD34B4Epi6scVR2Pj3ac3EYlmg+adkkecAbzy1Xmoe0df8uZywyCKo6+oQYZY
pIXIVi8KvFEesPUe/Sa3dHX3UEAbjqpnMTQTdI0f6bkTWZGFPrWjGRrJD64wL73q
nBeHT1cOYP8Zgjmty9aEMMQKBUYGClGwA252NmL25km1Lcfo/iHojn6rCHz97VBY
2dwFcvB0s95sN2yXBWmvZ7s/y9aNAdambPQXbHWfUApFSovRPHDXxVicxIDpT2BT
G6PDf9HQfVGMNAr1K9IKAoB6O3HkY2nF4dz0zjb/nIBcWtvnH1hKrM56c5INLqqP
M41CGv7PgEGBzl4tW9Ys4HFWKa33una9S1OnwC3aQj9hRrkyMMQpYG5GKNMcwIiN
JvNd/r/mI3nDyh7SsdpA7wAEpe6781Z1WT+x5DZ5z98wuZSF8uf5sudypSPx8v41
z0KfaEaJ4EcFwiZ9rbmm2gzSbrSJXrH8g6nrnifrONarz0lWkB6hWuDdZeLsu+UU
ARXD8ClkajV1M1NcUf8P1uSwQwf/ohccNrR0QP2ExIvo9Thp3UPGyE9IZCzJ5lbc
i/MRbMvlN1TUdSXUMOHshdQ0AOXhh3jYquBcfYwqJ9wT3UtWMsSPHy6Otsc7QkmX
LIYO9A8oVSss8dAssAyPvZ7SdkFHNT1maOdCNjnPoCtQyKiYF3kvWva48yTSXfX5
+E62paG4F1YMICXyExsuCMIKh+ULEj+PvdCYXeCo4VhhZ00imBqtKwKFrDuJ+nQw
cSazCbH7hwXGhTfYJGpapmTQev2h1EEdkH3faMQZ2i1eNRsnrGBAmnu2dvXv7qLy
8RZA1AVTmbJYtpyc+2zCvu2uVXuLoqOaVcyKj8JbLrij2VfLSGfeBi66MWm4ppTx
29sbd3h8OjpfhB7bU2w8amBXutvXrr33sqoS9rPNhnGTns4a1kBspecsPN0Bm0ZR
6VMYKFcvrRbdgHLdPb0yqAoS/iY81dfT43XkJZyOWz0ri72KQmpucdXMJo6pclIb
0MrbQVO2DNmeXTzMX5KajbVpv0cZSOL0LDFvhcFONUfwjXgmlw835WqxGdldH4OG
tDF/KH0MxYYiSXW3+2STxmgdgSZorsksEPqtxN1yZ8IDsQzpEG/K3PyUudbDrN8F
huxkzAImz3r0btpo0cyLVV8yy4CZLBuzGNQYqXQ/rR5B2ziJOmb8O15y8kAaIG+n
caxWJsNbEFtaCFVeiBPcXT/6VYC2tbASWkEkPDfHc/1//8ZzdvSLBqggeXMobXB8
OmUIMG0m8Pi7/dOs2HUUEri5dTIdO0ShwCh8p68R4N7AISZIsTmN7k8+k+rv65V0
Hk0905bCWuZjY2tkzFRFaEhWtstFjH6JvQjgleOOMcQEuQAUm54AfEphOSTm5bC1
+Az/6GRSof8VKQKTlMuRyJwbb6oRzEHIv2fAeClWTufQkscqUHL3u1UO6nb2/8QX
rcHvY1NuKdopINc8ojuizKwTO1c/ozksG/hTkxmCc0HqNiyhLbTjnhs3mTcxXdRr
19cyhI2X5nfF7Dso9MueI2p6Gmjbo8qxIRnCzkwyqUwIT+EzudH6uiA/N23yKnf9
5k3euj9zcJ0ZCVtlEpMl0XcqyyAFG0a0oRHCAPJar3csgH6z+VxtEuDNj6zAhGCy
gO3Qy2dajO+dJjVSYIYEuhN4tOK2yuatQ2QSwHeSeqL34vEJR3qt+PPebONb4HPj
hGpm5GXKv6hihw3gO1niUY2zdvVDWw5l9ufHcChgnO0dRLY9lJi2cWWNwIPZkcKm
6sV2AjEl+xw21s6afSlBg9hOw716HnjMkEF8Bp3OmoEvwaP2JupgDXWaVd+MEqmx
Hb08YiDqd4f9euvHrfgJqODnEjlrGOpQ3lFWR6MwVrQA9EiojdqvzXhhgnedgYXL
TBYiFH4c05UWDzTmUoD5myz3wfJzusJf2qOMzmKvWhyQItJBmaVGCShDUzFpwodm
hPUOwolM9HVTpNKL73gZVOFeTyeNm86zGARXWNBGgyQS11fofqLY+PAW89sApkpz
AEVEIHM/TdNBVvlAOeLfds6Wp/O4OQIHNnyY8dODLEZnA7QUVU9kvucaFf0SQoHu
avTfUg+7II+bBGVRhvPcub+7O/qMDgbaw3DZUzKg5/CSpdbxTzKGYrwqctvkciEa
rFuvBqhVChpVU8QhJz6TIccGtmBhzUWJo0abPpgoV7wLP9+JxhzndhjAMdpr4wfG
NryQnkwpohQwKv5smqybVQ1tA9HVjTaCfg68FSx8tdQhZfn+9wR5gENh5pbbNl8B
ZIbjYT7WVI1ht1ydka7lyUsx8eUSFnhLdr3F0lI6Nlt2cugbFfmpxrmb4jZS3bJU
7mEPBPB/NeKZili3P+yqyFsOTSPWNAQfYhBG8YDfYYroMLQ/RW68zfgXNhLtCl8T
uQPeM5pXf9wAnQFoDVpx03SVvRRHlvk78QKZvinVZUMAXr82GcoJ2LNPEwJRMRT9
Q3jt3IUVVMwtnwbPdqg/LdBvyA6FdBQVRbiOroEDrVmvpypWFanzrsV1H1gB2QIi
xF7+FewcDDAaqZSNZmXWiHBDabkXWsRiIZYyaBTQd3I8HOB9LxPAiCwxVnhwWdH6
NQv3tWifPeVsyZ6hlcpYmmiPfoRJ5rL/tmW0xKkaBKHU6pV01TkPWCLOkRgi1Z98
rjqpS3VvWYlZbWP3/t19GCwkjQoPv+THww12r++Km4caL1kLpehzphE4MLRKXFGP
KEvs7NhlhSiqlXU4lkELyT2/zWJcaJmfLDYxpcakM/AB3xn255S2MTHQoAayTalo
ONzQOr/Cn3BaX8Pkg1aTugKkOTOl2EL6DbV8ImG1yTResgXqbnuMUKrdOjt6oeDG
CUXuhvSZP43g2ap9eD11vwGyWqXIAjqHk0nlu5WyvH4n4bRvUOiTwsvL23qKtibK
KVI0gcGraUKsjK8VxNXL8e3NwZP3suEBHR4nGfH4LdBnUIt7OiI8ahlnZwvFK4H/
wTKMCGCcU14tfUhwWlyD1Pk7uCHRMt6qMbHwQFBfCVKWn9NEUCVX1xTksVC2RylK
fRTS5Rdl09PM+KkQqyr2xZglv/3r7hcIyUa+/eIAzffZDK/G8ROsiSDE9cQ0LHdc
QG+BOR21x67HubuCz4DkOQeKtSk7H6dxwLblOEQeKx6a1oBpLOBc6DF2bb42GOKK
0E70Dl2vUrfu0ktmme2ffhdQy+LgZy2QWjImBelsvR++dc/fV5/I6VM+ZUrhW2VZ
5etnmn7fFhGE/1QbIEN/WxpD2n+Zwk8hr7ZuOL9uMRWKlLuA1cA+ifYlzDqbIlUL
MdjWa3RJBYcVDy6fqj86xdogkaw7wnsCAKjdVReV6HR/y3saKjxSxMQXCFAiEgBa
cbcyzY9Ub5IF/0I2Jmv9z3oNTsT0+240PCSOm6sUTMSxJORkY3OGYAuULnJiWaHU
EPd9gJQA8J+eT6mI0ZeaAkBIHa3zrfox9bjcDNy9bKAPFYbMstxL8xdpYB6/ciOl
6SwMW/ZRkiv+GKUN7/3tgpj+uNzHIqkWJvf2wpt0yn5cqX6BRxh8jbNSdwa9MGLH
hZbBsybH/1A7TKWefchJll0Ic4enVn0+j+89Dk1eSst1YawzoeNF2Xd0lLyWF4Xw
Do/kL/2Bh59ERMUjzzu1hgszAROyvl4FKnQq99dl3ngaJqB6Dpr77D3h2Zt4nRM9
Vtvu3PmAtoojUBAMMCjyc0TMNMv02z9BC7pThLwEDpHNvgvvDpBNLY9AN0+vkxra
9g79F8ZimgyWaPySMVBh7Sss6a7w1+hTrgFbhyFOdKkF82hyq9t0wFcrmBCIIVhO
MH5yyae0I5gMFy8jLEGcm5B/kIMvodPh2DbP1TLFZC9oEl7z8hpuZk2LhUxazZ0X
2AJzosSNM2LHQqTDoG6gQLDAcmdAzsD9AqiY3nWzCu2gLHws2AopZBFLyqhGGMS4
gl54vQDyjsPm/1+PhaOSGrRZg9d4DeSQX2ESCXTfxKn2jZ7abywt48zmiECMeikf
eHCWfa7talhmAQSQ86/w8EObSBCJ5eX8ICyiGhxrcLzepVzlDyP4/PFzo0IU++wS
4vOJVKOliABHp+DtyyKDD1uX5ILFgloV9JJDYFloewqm1WCJTyvs4eX4Qsw/5wXf
CfoJCveNPTvgvzUm6GkUxuyiYi/rWfz1Tp3I7YTbYCJWdEC9m3uvH6RlQR/h7cDv
06G5ommsvXsuHgnSQbvphzkyUV7WHZrmw4WzoSdntjwsS0c8pq4wWcfFhdY9CvAx
xWzqu/VcCO+r4WSUA3xYndrZxoTEQ81w4ezGWYuzD8MkPqwalhpo4l4l+nhZ6o3g
xctIROIcn01TL4p7qzibdjX6zml6YUA/oJARSjQz8TirOeoc5KNrXVWQHBXJWCRv
1SKZ+NOg2uuhEvuGlkgbX6CPlt/gggxfVkv6fXeWPE751lXHwWm1a8MsO6IuOoSo
xcf4Cfdd4Na+8M2KjQKJfrtguhzeLy1VWxYLTJw5XtdUx8JThm64DujEa1OSu5E0
6WYlZj4aoBhJrCmeEZrKIA0LhtenP5ovbmLLI3hddDRFYhHj5lFLnGUcqrjkALE2
vYSkGQBgOYS1ibONSygi4gHRJeTJhxqzBXVU0/zKwVZJ288KN1nFm68sW2d5e+5v
/DcZpv6hMhf9llhpn6u0vbGcBEUN19oRqgkgNiA3XvacIvllZFvC9wT3EjkhbtO0
jN3VefmFmIVCgqK+c2Kb6TxgI/VHGFQBEGSlOdH4D8fy77W3mRHYLRGneg6hir2B
tPomsMNd2lQo25XoG4WAjZayU/pmOGGHS3uRgFbl+gu7iUm4mI1G3FQmuLMuFCuU
ziCJrOLEK5RSLq3bNQq1KQ49vXH7F0Q15soSumA0HjCJ/VFOZ/FVaA8ZxCWW1Pv8
IOBq2v3496rLkctt0U5xQd3fYD5xKC7P8uSTm5JXVi16S5yZPJGUZm7feSNpj3c1
/pk1FA4TGMBM36yIynv2A0GocgLPVJAuaZIzTYH014Oyw71dE+FguLBarTiw4N+T
ZqX5RPG/f5kVZWmBDce1CNgYUJozJ3UaQnVQWziFW1Z2L60R5bPl+rgHWhBCEnO3
HJdTlNMunv4vHkmPlavPijLy9bOhFTTU6ZkycGUMmgJgO57cv/MbBo7hn/PIYQOv
OMcBsXGF0F3EMDUFXDXDlBVTs56sa7NLJynMgMRK86SsH535k59VxmKdJZtNQ1Gl
NuH2Q/LCJpMvutIz41VbkQzBDXoDNHEb0l95d9ZzcA1j3grCN8+EipqOzty5bgW6
m/KNG7XhiYrAUkNqLqYoA9IkkzEHGBCos34n8/ZiE3jgkRD12xN0JxpuIMe2TRGP
iI9Ehx2J3kmia9MAovonWLIoKHN9ar3tjgsnP24/2xbpPUBVNfs1SRSq+0Dk1KjD
zHB005v8yhEyJuhGrQd+g410Uez8qHFot4PNmQy62j9KcysfCeeulKlqPvaKaf9R
WxuaVjLFK/hZr94/n6YlKU+FCqNUsMqpczYPBpIm+1RFu78JGS8FrH6q9oamzhYz
Elra74rK5oVXkeK5ZkKU55rgdDw8u3Y88OkwqJurf6w5c6EXBeYp7veOQC+lDHts
1wtkuABruMU8bzrFYzkDvg9sXCtpjGGz5xW60QP/dGfEhf45+Y/awSXNDcqxGUG8
/SrwkSjkvf+uutY0YCX2SrKvxTTCqpctaU5WdWG2pPH7EuH0M4RZFWlQF1Jefmzr
J8fxBJrB5TlAb93H5iy1FpIx1rlOZPLxbf2yhb266F9t4GHKPX8xuR8Id0muUXXM
4OGr4haEo9JRGSDD+gP2VMS673YZnosGxFMlIdbEcz7DdAal9ZzbTQ5pfFMEKXPd
46RgEggkw/qPjZU27hIB6S/ocPdCcXmRvXJv3zppwI1MQInZzALvbNe2OOmI0xD5
b24poaSmfv/ic1Dgj1P1PuzeIl3UaAhRUNZSxJ7OGiSdXNKK8BBwHXr1iGcsdXn2
3ETPc9ZKZa1w5YOxrLAQXMJ8NN9/y59lAhQvuNI9aPj07ZXOt8YzN/WMZe4FKtPg
n/DHw+H07c2hz6QsmsoSFSar/KxRX5kBiUwunl7Xx5Nq2ox0E9veQTBpr/SqUVdK
k3GezWrIDqGY4Sh2lzlvLhEUVF45oX1ofQwsUw5X67mY9KYNPmPf8WNYE38x2dG0
AF721xyNuYv31zb04EPqdhHiBGBE3M+l440rBs8YNEMWNrfdPYtYoJIpvP+4MOJ0
sF9RVPVIFcJ421bWaqvaFCgF3Fma5IaYS38tqA01srzvqkNXMSK8+HN4QuAau1ON
JyJ/aYEPWrt8AYRucCa8zBNb2gHMxvJnxzfpvdhVSSccEwxWYfmKjIGMskC1U38t
tASD3udDWQhn3BqFcw4T3P81Irntsiv+5cW2shv12abAbha1PoVS7IiDaKWROZdc
bh/tjmo89TOpB5ge6T+hEuuWA3moFSI7qmKapbU0JwRyQMneH6u+PQ6j5lqcUX68
1OAfdBFpaOJ++lyNIlMExxjVF2ZjWrRaCnbz3LY6N3sX7lqgmiZUoQ8tnDCyaMGG
qm/AuQdhEjKRUpbYBuusKjO1lwBJRFkQQ3wXCk/SkYY5GXc+sBHMuzcVKw7PqwRd
/aBADmZSOYWG1ApncI1jLqKSr42+Ym8rOGFIcWpG3gDjJsjmF++DoM4/04S7yiMA
SuqfHf0yYuC0nRSL39cKhLip//KFSrV4W5/2cYwIqN+tR+bM2DTKsaLqhtBOChMp
wmZID23STxZNMvtVoUCAJo0jhIHHa2/PQohHOrqdZzY7p8UZQwJszfLWEAPZt8HZ
AIhRu/WEXibL4FaJit/mMdiATkcq2VjRX4bW7Mo8AM4mYCajogIJ942tb51/q8sH
2DuGl8BFOd9f2YvO0pCBCYBMnQdiVfnFmlTBNPg8opfA2z9cNQBHz/lnw76DSSrP
fHuyiu8AiPNlLHlChSXqPIyGEKruk5r3FQkxPRdLr6ZT8SMJt429/jRYx6tFfas+
bhI2/DRqwifjzc5Pt0ktPPXBI9jpmM1vuH8YNZnNHQvAb+wcmg79e9psZjGrhmIv
4ctRiifsLj8uN67FMRA+rAfA5bNYnEcwQYnA5rLw7A8FoqCs6BJmGl068BOQY+yo
eUBWoQJ8bkzTlHZvBIOpbbn6DFpq0Dco20cWV7eIiUXXn4eYTJLSpgxkcsqo+SZ0
5bDX1oE9fVMeynLLqxJkVchcXmXekshYY+keaX4S795piGO+hHMVFraUyYKWcFBa
ONU7wQfnmDEoDXs2dFps8/NxiChsq4u1vIpUKPsSwbDVslPVVqSQ6C//zNfIDOhM
HUsjazg7AOWtl2SDnmKq6kd2qiXicMT076P9aVR3ZgcQzvsUwJrH+SakZP0IOSdM
I0teDC8T8c0Nn8C1knJI7pbZ5V67CNwiJrTzFe7I6YMJaCJhRjH8OjpH5HBYxHkN
iezkH4XdX8aPRosDYc8nYmy+jxwwdZ+82bY8jsjNDi0+sBLAvFZZljMLb/+owGLm
jT8PTo/qmKbGpYYG1aQ7voUwb5BbnVSvGg4lcnSpF7220PqwBy5HbYIVW5TKDgrV
2QDCrM27VgSdVZT8JoUdCNGnK/1OW30f6SNp6gMPIFkoLRy7mUv9EKislYXuYrvC
4xJxoF8+FUceul2kYgQ7NivENN+Kaf+TDCBK7v/a5wYWsSVUMnb4drxY9b11TbT0
GB7QueVCqmgeci0lZLk2oHWZVCOa6vAzp6czyluVHblUUQvCWdERc55RszfesLio
jw8Us+EdmrJO6EAYeeDUeau76KScvhKaRtjVUlVIpLwz+PE3950uL2JC7FpPnQoF
MFybDnoq23sN60bLWX4/WmJ/dijBQ/7uVMKTMpanqFY4bRQrRRHiLQ3jurRnq0lf
Z4owEU1SveZoTVWFHBjnhjhzvoWFhQh1TmioFchM2vi+DghEgjaWQmsmk8ny9Izf
3HOQIwlDHkIZ4s5u9sl8uCZoaOHXEfbP4qXuiM2BFPq5y6+vzRFJljvhDjto8wNH
9nv5d6AsqJhtNULx7ip+dnU787hwj2xA+6lJXNxaiU1xPGW6ebwoexHDyGTwiWhK
p8g4aOa+AYVEXgonaS36yMZOyi83+rcKm/4OVNBJJerkAKl//T1w6VfNgcCNRyiy
clIBM2F+rYoljhy/unumXZuSjWxT/CVexqbnVPYKBFwBuYXHbeMKnUeeYYxdSbq7
Dyaw90/MlnaNqxeQiLDKGClURa+BGbbXoKKPfERwL/ha6UtfiGuqVc5CRkHp/zss
JvfCpPZO2yAmNbs9mODDKcc3WpgDEwxWSgsivRRdY/DSGO4g82/SMa9kp0con+Zv
hFZDxQoaNQS1kXtBd8JvTAjDq2QnB3tQB/AlJYdMPUcaARZK7fIEUK8CnOzr1HsM
I8a8y45qKbw+Qyf/dJx0rvdkFhYkG/vYcI8xzbWOXxeVeOJBKxXqEAiTMd8M7JQT
uBI69jadQAd2ZMNulMfNi2f6Ph5k331qE9CJINZDNiwef992y6/HmiVWrdoaymqM
s+DGju7MClEhTiwBnVbuPEETVy6HUOVq7rivjX6wcvrL/dGTSNF6AausJcyOUFsC
BHKTB/HXMSsijVTB1sBhp9pwqtriw9w0KKodqtiZIRw4hCZuM8wcqlGnJFBz59a9
P0dL12cjYn+YC4vwMy6kJcUnMqpfejypMSr3vqRjb6oXjzDMIYnFur9ZVFqy9caz
w4rTBCboEIhQieeTEsPIZvScjwPnUYOED094r6XCUAozMutXPUfNlqzSFx1bcwBz
E0N/7/699m8TaZEJp5O9wsqGTPESRRcbjd+82Px4VTgTi06UnssJFDoaLRVUOhSo
9gQGT7/Ws60auatZ8y3KQnZXCfm0i1gCJ+cvsWLRNzrDWgCC/lDrEfnIObFeO7D1
QIGJHR+HlU4uqrWdPZ/nkNFb86VWM00kmxBB268YqUQMp2kz+2ToitHqEA6pkMF+
rxkhItDz0WZc7eR+x2S9/I8G1n2P8Eo4+kLKaGISrY0j3wZ2+2KrsmPcJJ6PpZ3p
+9voDsvZM+BXRM9dhR3PDPWQdC8437wh1Z/mlTlFwu8WOhx652svbdUfGv+sYCtG
cyTrQJfEXaxTpes3nRaroY+YpRoTu70c6G9JUOTCulQAliIyK/tJRRn0AjJGdKEB
S+638Xx41evJGpBM5aiRx2Ht/hln4X4mlyYVoVS9KdK0TxR6fzNAEaxWoBMvF2IO
UMTJffUJ9ppLy2Z5lm7/DP6B8pLq6YiFkxnYM4RXI0bRlI1zhUcn/p9G9S578dnW
AfTe/t2+djPr1KAHW31d1e17T0YPrXT+wp/hvkLQhSGoe0ARFJuORdpMhTF5jebx
8RSryjJuvZTbN3cwbYOk07LjbjPmjCFuU91mfwV+9i4Cx6tDAdaKBXvlm6MfwoXW
j9QZyy2Ff21Pf6v/Ytq1OI3E83SkjjupfB8gLbsA8Ip1SvHhlXiU5utpK1BNQ5Ff
DiFemdQaasDnP+h0Q+2YrhJR6wiuYRBlQrNVjgdeznciSuhFL8ZDeOutoqgsB/ly
nqtBzcv7XlaAwafvzOnoXxGnPiEUOBZC/FWJOrqtsMgEQtt9kwQ4lig3RWlEwUW5
XuFwihVmy24AWperfHi+1apcxFP5J5ikadoDbSOO8YOQhJelwJ3Wud63s6zyrgDK
Qub3sxvCGjdHqvA7Q30zoF2ytah1XrBBnx356f7zR7wWVGZKYS/gM8mvkUe1sSoC
yWFQzXX/TNERgjPhwZfVri+WAeXJcRBRRqlmprXk/CiiNWwyr/ZgdiGGEdi1h+vx
Z+vIUWQCPWvz80Lesi/2liMwpiy43477rIc17ir/Bi5teJaZODwCCa5FkSsL+0eM
imTutPs+LjoglKU0/JZHkvX1pLRGv/wUMGaArVnwbYwPEYlZz9++oC/xWbckbSmA
mBp8BxO7gw34EC0q1q+yNYOh91KFafRl4Qw3hxEPW53mfOi6J827jI06S/NFS6Ni
6EOMCF++z1naolX1U0C//BhBl/OFp5W/j3ic6t3B4NetLLx7JPvaWaCCkMzu2cGZ
/8IXhXA2ynQDaMQFlzMVvA2MYV+p8xTiA4Cw95pEJRCsBCw3TdzwnPRYVdvX8KKy
eaFBoD2qffV3PMo4nc2UcfLFuVQXkA1NA2v+k4P57bk9zSRJe5quEUA3q7bBa7Lk
nlS46T7lHSneBkMaGT9K+VK+hwSUGz7mC3f4U/8dmFMYhxl642oQQsG/VPgKhXDF
nWpgUTQBzN9wx6tCNjGjzQyCt8b0O4Ve64xmNPczKgc6vM7RNmCQQAU0v8CHO7Sb
GkJqyQv39f9+/8bd1wSkU/VIEJeWcRXUFpkiqie8vtz10wgXuf4F/P8rswVPfg26
x+DqV8Bphv17dPuTk+vuEs3NmqpuuvNBrHNtaxNgtxrzSqUi/IokrsYYwHK8MUye
fBjHh/tNk2dkxlA0G6OirhXgReQ2b6wwSrp4M+75AgzCUJqg/XOKwyp6qwsqYqzG
+Mx/ynQolGCY4INGLi/gvoTrhUgkAyzQbWHTDZValcHe2Vm9kTpOWw0CRbD3Rz1f
g5KRR8GS1zwzTDf6ITXPrffd8GSkwFJnBucE9k1gsV4cUCh939eYHRUb3pYXfdAm
wzKOuH+FBmOzVMTtTjpqYzn4GunJKqHlhbsMsGpBAIK1CExBtZMbeuXyFZsPGypw
4SSZzKmCKVXgcf7khWafTFyLnlfiK/7g6ekGtkxwd/gTGNKKqIu/wOD+P1qCN56i
bG+aLYvEtnF8nZuuofiSMMeCZiyeIRDKf/5lV7mOfrbaatqIkMSlVK+hS2n6i24R
P7GvQCrWZqdU4anydqjkMzC1uyqk1Y6ZMsfctUvbnJvzMTnSUPawqKO94JbvLFE7
eh9f94fU9N0mpXwvMDkK4Ua/y7mlsDyFgVTOk9F/pLGoulojEiHeDg5SJLdA+FJC
YqtjKurMj8ZI1YW951+ugF97xLSesvctCwFU5Xh+XFdLCkVRhMg0oqgmxkXUQvUo
f50tytgkJ/eF3dlFI/Zd6P3P1wEoyaF5BldEPh++c2kS3tK18+/0uAB9Nj2+u2DC
L6E+Qq0IBXDtXW0nEtx2L0DYH4utQ20ec3PY0ESSEEGf+0EGbJSPfxmBAkZNsenE
FW9hYiBxyPQWo0grO4a9CHqy82XmFPR/OmGzGevRph3px1863XwFA9CYTeZ/DzrM
8YXvI+a5Q82+vRznX75EGJpAxprB28tArI3SKICWhf0uujb+UQNDcLng14Fh/+EX
MBD/XcxBSY+mMdNVS3CQaka7ow7aO0y+NsGigLHvp2MH9CExnuvEQJKtIIlYbp0p
n9jI3NtuSqttkb5KYa69CAdJSpSRe/hg4x6yyE5b6dnTV8lMBMgK9Z96F/F+PtF3
ZLl6LIZg6G5ub4hvB0WzU7i3gX5WEeBD4CtFqAu6WbMcwRiWW+YYgl70CdKIiUY4
Nqo2GTLVTil8xPL+e46mozlFyZAV41FcnYaZZTAmSjGtGvpgaf9JpGNLwlhnHXxG
dRCoELfu8+d3djIJTpUz1rTF+EjAOgwjh1x43+GMSNtxNl+Vy9p2yjFGd+p5OHtD
DEsv8M9BcasbOpo95WidnW+8y0zFB4JBpkeLIFkwr8JNqOHZ/rbVgjH3+VBcqTP4
CasKjPN3rtEVcLVIwnd6/LH4uCB1+s5rBWZD16M0GPGls0ZWdsAege4MXX29DEAl
w9MfP6JqCJd5CUVuSRvfy12wND4O2+hyu3O4NN/sXEZh8HTqHGml/9M5Ccky2S3s
1JddflFDdMMlhu3TKn4G94xrdFCbBKCWKRX/irP8z2+90Ksukpmf9OGIG3+ABuK9
+I50Q4xGyPb3k4YTGXR/An+n5w9T6VTrQNBaubKeGGcyONX45Vk7vvelktqMJT9K
WNcxVTpK6cDkg10dzYK8aiE7f8rdkyLbekRhiuaSCEo1Z2baCxY4tPJbeDZ6KjVb
OPAGQYk+FQ1kvdOJilKzsw5KkJZ4AEpl2paX9n9dkF8wZpycBiTlWqzUcUX8lm9s
zB9DnmTJQYCW3rjGA0UzRjxDnEdbjdTDsq5uR1W1UgZLEuGAysc9aA0HQ+OwnyB0
WArEcmelqCnRhtq/D17whjTB/AyhjbgmOQTYdbNP8nU6VS1iQmKTf9ri772Ahz0j
G+rjA054ZN2PrSzEjCg/iU2NBEGB9/4Xa9snYIfmP+a2UeGHs26GgwDQN0hE8/Pv
XgU3uxi6yMbVttKu66TPDrx8TbO+IeNXt8U7LfNkvlREBoQagtjnsla/d8tfS0Z0
aY/s6Lopvpy+y2055rifxb/DDWPtZkXfnRE7tsKPaGWt60BA1i0ApVA47HiB6Cu5
5IOrsbTE9LR/y443rC2roiU2ZEhzpzHCV+MdJnKZwWBgF2eBaYrU/W1fPBf5n5Hi
pNd4Y4MRWUOPYzmWAlJsqeaFFW+kdfIu+oyyMRSArTfF53w105h+FxPENsQ7hefP
+XPZlkpITs1y1x0PTfsDFG24IxCvN8+AVwhy94oneiLosTDg3jW1x0B06uLaYOmr
ZmS6K+o2UNr9zK+oPmEWu3+0FvDQISKFQ81xg+zrbrVYCnubwWlDzVZwx9DxNVuP
/5NRe+f8cxmYKMUIqVweAbQrvT3JqkfCAj5B7yzmhqHNzechjq/idvJLwH73yUUk
3rLzx3TYVqbDZYPM2c9dPUG4dvjKprFuhdsqbuOPgiqug8GPSF/Cl6j23j1SDQaQ
w/+IvBd/kw7Zlq7AFQT6cJyeKYllnMOHYmRsJUR8qi5ULijeyOMJKtXR0VX3eqf+
JD8elFBrB51R8xCosn5XpWAFgwBlFiNrarL2w0ohpLdcBujKDXWh8JscNivIOpFH
xOK7hbTk4JS+aP1lW5zJMJ0ZNmkPst9GFA02Mw6z0VxlfjkR/xXDL8/ea2zI/6oP
1Fp9ijWbmN6FqMdvwt0RbEiPg//R3NciWlYt8JxoPHXEWKaZBP3OGnAquKXI9zzV
3a8DYf6cpvvhe7xHRiDaMTdOq8MRsEY8KDzHuQaEFLkrDR9JvCF6a8xR50vYekCK
IdRfm+h7BFD0fMEht1n1wrmzxcTOmcC+IrbCOzJDDqasUyIlMZ3mr3bujHR4UEcG
1K5JVGNDHfR4yNxd/AppeQ6hXKQ31D9JUts/6RJqHbZiAsIxHmUPmhkACPcTQbaS
cJjZMwq8M6f95tX7sZ6GN8ArboLyfgIagx0UmjhK95ElHltbVCsYkDvM3W7Z0MCK
IX5Gh9xxjv4QDALbd66iOVtnolL3xR0odEGUEejY/g5IZAROj4AUMc93cBWUZuj+
syqcWmpkegQ3z0jenDglXd4gnJRGPX1byrd8gCHDcFW++tAvga8DVrxCM++DNjZP
zA6Ytz/mNjkppWUMQgzPtXnD4e76LVSY/rpF74Y19dpSl3ZlOqPYRtanqUSlM26q
PKXqmW/z2q1Au9nwrFdD+by1jq1dFaBc8KgHokcanfRDJrn5JrYzOBjqocbtR/XD
ggyBF8pmcZBHnCCjNMbekDhMv8aEo1dBttwjAib7HStFtwKWvof0rLYNq5M9wOzH
XIqlvSeIKQiUZn9aTbWb05bltP6qqxu0eftQRiVGxYi+2wJND23x6oC64bEQEpzN
Pu7y+GvAbgXmvhKROXMDp0IDFx+/K6yOog8x9eRYYdI4IAtbQY5GDR1RARdj8ZdJ
g7J/dOr6xYB8L1TycpJs3F8lRlk8Bmnk3LkU5bIhzXhNjfyNf118TQtEcPkN9R6e
waEcRF5GhFSbMuCtdsouMRtGjMTXf3CszNkbs+UnNu6jY/BGKlY2bxIdbNIVjWHq
4UkhCl3YHSA3jshMVqv3bgfTEb9wUiKb7qosDVpIZTDkXpJzIEAP9fNd5Tm4ot0m
Fv05GiN0liHoqbr1xnyOxuLblnH3wtZAn1v+VU5ggGTVHbWQXXt6kKWZQVsSLVZ1
JIWrzKspaG6w/11/dHgs/hd1CiJHc3v+x0VPmL+7LuReynxy0cn7wi5tsbA7EDTe
GgqQsJY81SbqiJyrZPTxEMyeq0b2uFbcwA8kA2EwaOwXsM0Epvzo+yD+rl6v+VDU
lWVWq6xCFradUFRg/7mH5TmTqzOUgbZQQgysFPn7V/A+2LAhft5nb3F1F3T9raby
6uTddmhNsTSDKW/5cjPefLeROyq4z+gIYI/KAUY/KRygN0IK7RqMw3fAPl8kU2oT
Wyg9YWekAbicIFAZuEmgsdpExvIQgbw0f5EcDG4dZ7qNTljEizH+tHixXa8Kltfx
sItbRwjiluy2UXTD7hFx6zFSEyh/qHnda7sDoLBBlFdXZFZ2B9kDgCopyHidXlLe
eE9F6381+ohtm+Hvs/choHmuroEZBekUAspzClhaA+d15p03BnoEkQJdnDCOebcR
Yjx8EVO234SivQo7hCBib0cJbh7vTLDnYmrW1pYdmlp2/Raj8R6AXi8YeWyA5QIV
LboBzmdznDDjrSlx2ovKiiZ081EjLvZWb5nGHl9OcCLjQX5llpGX+wIXU2Z8bpkf
QzHH/waJAbcLDJEmcoJ0Nr/0zbl2xUTSu2jnreMLxcAmO1X95/wnTy5XVnXTEU17
ZVWq+f6yrcfFTNP1r506xfjk8TBaGUX94I4lJWV/9T7icKOQrBFbPmeF5ZW6RIGn
AiH+t0FqvajwkDWKSjTSFaX5CA9isd7xSOlkPj4uCr3TAV/yM5VJry54/2Cjzy/j
7ecykIMwVtw7vwH99U78Rc7yqvlJbG4mfdCealbnOa+9HYDvdgLhpI1RqYRsFQF/
pDn5jBNGlhdwHQmjLtC5o3QwywYs/ulwyYV6q10/bCAe0EQ3G6r03nwa5Tw4iWsK
1pxVqrMXRSOpDxwlR8nmdvo8e9Y7XaMc40GJUkCzx3nRKn/yClDD480YucJ1hBgi
tNwVjXSwu0GXIEGagkbGQw7QQNxphhjrFIRwXVjJ3cBywSULBELsAcUEGYkp4+J6
sMohOTOcs3b71rzO+Q6lZSlJj3ULb8/bTGSZ8jbTIbYNn6LrAuAprQ9RLbhNMzPE
cdejeX6XHnyxk51Tp/PtzKnodIThlilQYFvu6+CeFfmJAEW10mh/LZyM6Nks5kiV
FGjrJP5PtRqZMvZJRKb5RqcuYVRR9mt+9NQHeZycrKR6ChIQYwPMnm1djYr7GVa+
iKfvTPhspDELnMlyTtZAngWiyG8MdonTv5lEcd6Yn4aScX9jTz96AXuOFJ3LVcMV
Ako0e3We9ZB/p1wldesHkUl9i95S0Xkc0/e6KYL99graip/pfF6yd7bpfB2Zxj+5
HquE7dpTPDW/4o/ZoYFZ4lRDkInz7IiZY3rVIjXODuq3bDujz9QDPmCCRnm55q/l
j7gCFg24FGUBoz3QEDqp063hKLxktjA8XKa0XN+TeZxa9FR0FMRnNJdRzepbwvOZ
nXlNGX73IMSMU65/1Z0rnORwepAaNfhLS1487imssr4P3g+oT4VHSKd1odt2Oq0W
rHpFCXCf/AKW8DOTk5RcE4Z6q+YrWm91nKVl8BCfanNWOUkSmd8FuIRk9OBPOW4u
C2HBKE+pjjh0pq//h4t//b1obvvOnnm2Pr7A0ve6wHFvFTHJwacdGO3FV7KesGEj
qt3ENeKcT4uk3btZcv/xUv02xT/makT65+v2F3TTvfrTZaZII150xbjbPnhPe9sj
50loQU5re3Q2vfZ6BruHmdd5oVPZ4uGLTPxVC3XhoczG+Qi1HLaqDkHQNea7P4P4
VdJyR694ZPTT2Cru+MI7y6R9VHvAQMGO2oQsPziJ3Cjw2Sx7Mh8BcWwVCPO+jbp9
vEmlMB4SDepO6/y4yN1GAgwWbsDt7woa18UrDOBokoINM7GGjGNkarMsgW4FZcK0
K0ppJi0SPFQ9n5NIEbJo/0wHt+MwmDArEkQTxqLe7n9iGSzraVvBvgZ9Kf1UZC4e
Y28WILBJSA26kQTsYU1gk731hoVmsAf46pKjUqLuFwCRDvQyxL5Auc89kuI/wxOR
ruKyF8ZkEAGvOIDQadLJB3NJ3n7I3blKNcRxXrRBGJIZfue/lPrQz4Rz2a66uFJY
7fzhHqYUcIlREIxV03WWxfem8P8R4iM4nPv83uaQmw2J5I18SsvuGPLk6nO34iQs
Ar6QvEHf9FOsr+yIjAsjP+D6H5yCr9gkb8yboVRXHuAoY1eQ8oz8/0eJQ2B4o9G5
U3oTgEtpmPQGb+2hAoHZuBnwdJP3Cg3gHhD17ZIP9axdyo8cCJFsrqbDRhWeBhAY
34Z64HKXrFeb+jHgqs3ggvwQMv0ZytQK/p373vaRUaatyyUWtOQriIwk/S7L8AIb
cpNmPkCPeWekT/W3cyfNVnF0TaoWNOX+h14acUbMZiS2HvMEP1OrjtPPdvq6Ik7c
qCu4J/6obS57431cQg01junMW/P4kuCKJ0yEVCGovzRjz/kOpblp7KrCZSb1A5l/
tNJKdxvAkHiWs+fDK2IkbR0vzrZ9792VfokQrhdnZqr77ruBfFik1fZJCSE0Uqt2
KvktwnDMIqbthWrimj5dK+klPqiLNfbxaQ5o0C7WBb5JN03Hy6B2WEMgFxqkxfyV
c1GUeiQJnv1rscvEk+eBFpA3SbMslTzHXhQ5rDAmIbYsOq7zl4z6UMueYXZd02nd
LCGMM7j+KikqPVPfXPdn51Aozr2YHlDGMYwsDWB8yzcP4Apr8ecOFLNV2QZ8HAdy
iudsSobFprVrIrk91KHy7jbspsG2VlBPPT+gAlGJqTAkGdl07OVjYllg8vbCG1dj
CKnfdE7hhZ23WE1dGlQNv/e/Kz2ZedBlotd3L7VCVVPF2XHtjpP/hsCkAq3HtP9L
JfVjmHWqHljK9AV/RzVNq7/o0GwLTTEG6bPnO1kSJUQpjqXt3kpdu0WoGZmnX3lf
3FH8b7MYvZux8O4o9RzD5VNxr+KF0QWYfoKy1jF/QMPsImLmyxjrjimRC6z5ypUD
+jevyjT7VfpZPnX2rfox8uwZdpt+FFr8hrwrnXIpuJaMqVJQcSrRlvLKOeCsdDvM
1AQPrcksLLOvWmUp/BeppNaLJLcVptKxj/D8cv1SkPpEu/9rWZZ3QntYCMj9PIJk
RZBIXXCadbWwm/+f0uS3yCE0eYZgSnGbIvND+RskFZR176O2P3WV0p1iL0SmzTTM
fWDCow5li0OoWPoglUDx/kC0qgh90jr9TlQ5ILvN1zPFIYOTmP3YbL9l0ZJWBypr
inE+twnmHNq6wEtdXsavIbNfQdWkHp9tZ+tgss/ILKoSGdw3XknPQAC0U7fEl03P
87oYhhPH/0lCiB0quRU1gO+KhJMUbeNP6iKkyLD/i9KITt65xSEXY4f0+n+iqVBf
S53tx52YyN8dvVwjXXHQ6K7C+tWAX21V9Wac/J8BF9g0Fv6ZvsYbsXFsH7RYdKkQ
oS05ODNXhx//Uacz34k8U7tauniKHYOIljivX2PMg1J2VRrPwpRC0yAmo/KdeP0P
3qEAWJjVM//70iUHCrdAL4zqMRrGWeXRsPfpauDaMmYEQbBUutADl4gNflTj5z5G
C86xwT5YlYpxb+zPWkhu4dOYNcr2DdQ+LimiioHWgEQ99usXZ+XY87uQVCDY53Zk
p3G9bbghEty4NwqVXav/fKroj3l9HgYIhjJZHOShxrh0h5+wkxJk3AQSLQbihA0U
wIGvfDY6fIqe59TbsQgrRzwkSoaIYYutpd+Upun/LTmUXbh1YRsb8MLjXl77bkOL
W2CDRltSLV2uZwF+j+4lXkxOzwC1rUv4RYh8B5UyIm2+m+1PzHi+0IxPWwjt4ZkC
eKzVeCtGd3ElmOzptfvD/soMMo5nU1d6HmeTmSxGudm/C8RQrWMjO+hkjKSM4Yf5
aCxfkogYiq87CAe3BRT06O8Xhq6XuEhd6s8Ojm121MJVClvBAsoFCy73vLRqbgP2
xr2rQW42iwP7rj46TC4k6BlwWL1QxDeLxtEE/BJgmHKAmYxetwTCqxzewtEzbAGw
OxuVn6YHeKhJSJK5wiTvOGD2eWmbadThHM7OfI8cE45RqaN0pk23OzBCkiyI0Ofd
herp2Pao3axTyyMUg28vR8o+KgF3QPIf2WH6AiDEvw+e+Q7VQcAklchZhw/c0FFU
iCuMt7eg0aLtZubXAPeyHkNv+dawXRh98aoli8EqVN5BSyrG9zUDVWBt11jt8ZJN
`protect END_PROTECTED
