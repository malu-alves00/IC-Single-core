`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
N8LcLx/wAkr/GSaO2C7Y8AOCGooSnd0l+oCtY+8jHkKkd5Dav7EW+Op4lWYnCu3X
VefW8GXXlEr6aldUivpaje45r8mqBRTGjRMTnRkVRUn7V5SKe29DqP7sNsX3TKtr
jSVjZSdqRHX9Cy+Nzp/KUoSzeMzYUE+AarV1aGegxx7JapOQLlhWl4qyU0XF0oWD
t/o/aIgQ5DH6cr8/JNd+wlINJJvP0eFTRy7Ltuf+5xJrHyzBoCWAGZSjnyEZ2KG7
5ECNiSzGNanrNEYMQ2hCV8dHb4lY5VqRBjB9IlU815pDEs2JuO3z88t7wfFpvX4E
v7cDjLKKYFZWFMIiNmIB6Pu2dS0FJVDE8oUYek0TaiAuP76bmdbz/IU9kdpBckRk
Rngibnl/qFkMIJidZEP0S2obTDpCix03r8U49S2Wr1ZVQ9KQcITQdVzX4ZzPXOyx
2vBULgRvih3WYU7eFCbxyiIYGtUtgUM9Qcv7wF5oO0WkZfiveSrTOa4ymkqGSto+
G7CDOuNtJOK2pmv5sdbz3bBcd+Z36WKUvEFAhj7ftLY/T/Dv7JAkEAg3cZ/UUEQ7
p5dFwPUMqFwxtBTKDSwcN8UD/agBeOIyGEVF4XP5fYYecw5yiNu9VkyzmYgay6hQ
DNGCtGv8dUlRmrACz7E7vFMHBE0sINC6qsRw5PWF355lCG8EO4vdiCh9xueDVnch
M78df2xlsq6acAKcbg+P90pW9E6Eth1p3XFDVwbEogqFyRQZIlXUx2bxVwCXysyt
pkKGO569or0Dq0AaYDffu1SBpSzjZ0zAj6VMbn2s6b45cQT4F7iI5fP9GsUi+87w
89fEdMLDZsI4qigr7akRZWH1/K5E6d3WrMOmftdXAEJOrVomGjKciJFBqZeQ8UE7
kYwMpCuSKmeoxqe5CyCkTas6cGv8Z9VkjDT03dA2lAvmVA1EIN0SuvRRBr8ePvU0
FyXkHI+EFeGHD0jkIeWm/8XvEXCXmZIlLGGT5or+Et8NHhdZfLIo3a+MWWdkv7l4
StLgywJtTm+/76aldAUOeuD+p3B1k2UOQqfoPrYVhAFvAwINMtqZ7CHWEGFj4nIX
y9G8xNljAN471qb+HrUPoNeMC/exkN/ZCNeiC2vXDZAjJiDXqgMlUzqIkatlxEXw
9F4Z43dMBlJ94ShVgnf1svbqsltG032/dFBr1bpngFLYifVzNSaB0GESetkbWDvb
vuXxdLz7J+qEyx68MIh6xoIVV/7NsWRzNjmwTx6Edv2qZzcO6csx67ESt+k5B5Uo
7Q5HhYfgnhAIRowmPoKoTNO9vD9BSAATxWWirkw85VHD4Hm0COr+xn3GivaZuzaT
lozUt1kcqBDNLim2VKGf9YtshYCrp9wcvZjw1tT7hdIJm8bY7ABF4vBkbNp/bbFN
c1mU5xYzIcMS7lR+YNlqrmFU6xvk3Wgp7iHESDIOzcJXRqthNjJtWRVyPABHLm7C
s8/EKPyS2WeJTysOkmzN1mI1Ohpei2afNYI+1C51p4A059B5Tz2MgHa99uq9cpB9
tr/0MqXisQRwKQ2K7Uilf/sUsMqzTVdJtm5ZIgcXInDC+QofPntvDRKv4aghx0vI
Jf2XAN+TnyHTW8KyySluZWpkxv7+fARzXKSk4DMD7xwmB0FZJVlQwYOky2M7eZ6Q
IXnIEV60qj77yoO6JktWlJQ9WUCYUSCGXANzQgcHtVARVKm+akZDKjMsnR3OJgLs
g/4vLmW2PdvhUjkS6nUXu/jNAeyD2RZVjokCqHkgg1fc0npdkhmvfH7gJDXneDE9
rs9z0Xua2DdoJaalENRZ4kBBeZzBo6TJKr+kGUUnuUNbaLJEaqQNlytLBCsZT1r8
JxJ0Tboo5zTQrAeCHNBt1yMqn23oHrTt7JGuzbuZ4DHHEs3lO5kaLdeOwOzcM1ER
xYuztoo9XSG7yzpihKK9TfI8tYhOOFi8BCPk1TMbRwhYrsGOZlnue9PbQ7BLRieP
2p41zIUxBcFSA+kOizJktjwfIaZHs4j+Wvn5qm5mo24XGxGwKmH7SnhxCnuObaP1
ZkTpf7wkJpmGiT+2tnGS7LuxWvo7athI4krVJSGQN+uV62QWqvQLzVEceR9n+9/u
vH1hUKn0LelotUGQGWJpZ6D38fnUe7E6FOli1H+O5U/BTN1uNXnt9YRIAP6KE9vG
2duEqvjEVJVZ8gvU+62krME/Xx2D/8pfFdmxOGs0zgTKPdrMSqfwNN4h/EKwzUem
675vT+EqnC6ujptxOsNuEaGBeRuZkRcM42zLVv8amkqdXINIO+ANpEVUXskGl4mG
VrKDR/PJqpCBECE3HMt00ODyW0xRwzRq+aNwnuiD56fyH17SL6UNzJgwv51yNIus
uuY+vkMjZzDDyrnk9pN8XujWc5mRMF4bnAus+tEvVYYFWYjPiYLu6nx1jIfrVnQT
9kVD629KdTxrurxdMeUUj6K55ZMpREIVe0RzKqMkBWaBx/xiAHZ9y/xwXtHH6xg7
h2w0NBIQLRUUnQff5rm1lSDhvf6hYOfQT4VZMlu7AAetY3VebRrugOPKGUntKVKF
7yBw3StUNOIz5NzIcmsjfA8Fr2eWkLd/uc0TnxbKjBDoQQfFMrK65rwhcZE8XK+n
zihlhyu9Bc1GgBWPzzkezUWyFvZC5tPRMfbW6KmHu+DwmtyINeeAgXvVwHonzW3x
dERQhQSyQ5Sx/YPLEW+gqEcOzNPKsrTT/N7+h4TFOmuN4zXMiwbtcsqOXJFxpQTO
2JYikQD/beblzLKpY2jRHFEEXksPt2LcHGQyjFtp0WmsMBIQXBPFxzgR+xEx2oql
LyvweHNZBBNmAdsiVfsKGgNY+xYPIyJ8Ho/jrYtLVpgbS4BVdJVMA6qKQLlFSiMl
ZP6qxj0DJy8iQuJu2esDEfUwLbObPyfTebxZ+AyOIXY4mQMpjfKdT6AmIGuvfrS8
RvmkLbbkpudK5m/T61YwmUBkrOU1GYjX7I7sogzy8iQHJs6xoG6kjbhr+OyZSxgT
327oYmvPFr3m6Oaw9fgujs03jNysk46J8JSDeb1CuYKhkvZscixATHDbCZphJDoF
cWweeBDgrFoXrfdeAxlWDsS/QH2HqoLUJ7un9F7yQxG9YD3fjIdRUQyUuhS5wv+F
Cyt2LViRTLvB/+qwc9mrQ9vuq7ZQSw6qiiMT3MzI6UKqIK1KT4tkQQ1nliD8WsYI
YLoKuDoYJ6AhXyXKmS/k6+eV+kGrbtrz5l981dK1Xg/pLK5pA8+aaZ4+bj9Zmnee
v5B/tNxg4dvZeIVaPGkPmDYmA/ujyhxNFlGZJ8nwx9mEQAWCV1fJ86poMWOZEjub
jbCejEdOt8mF8bPc8OHkWU+bkD7rGCdVfxtgMivgUiH5hHmURpWw9ROS9kgmQLU5
4kQsPofs2NVXTDeB9S5sVE+mK7TKyJoXWx5vc36Pdwkc0pc4TGE0FXBRGoBgbHy0
bCKUX9ETuzFiX2rdC0IzhsMjv03t5h/qDWQZeDc9ztX1GpL4M7Ighp90Rtr7OC2R
jlCdjVhpJyPDMyykZ/XxFuCv8c8l8SRGARPSEDWOc7a1N9dTZwO3AAebs98K1VHP
hKkKIL+BzyZUF4CIcHkpkZgXbikKbf3FjHynMteDBYt3ah4ycaavi7FwgaaoBV0+
RqbR+HBujcqvUlTh8e5JafAjixCkxES+jS2MuK1eAekbjhvzZNYICStWpJJYV14Y
M4iR74EltI3yVdfJwxZNlcH3qCiFRPDR9jJ6pQgzyPecI4L6GvQ3mXLQ8ljglO8i
LLUxFGc3/xiQ9SXdschFcNG1Us3P9fK7gmzqr6zBvlf9R4CNY2FqCFUuamcqoqPh
ztOofPgKyoxkGUNI23+Es48fOD7gsnpkBWb8UdAwnlMwHRkJq2MIeeK52AuNeo5P
5v4hNjWohYe5jw+y97ZsRYQR/+5n1fI6eXj13+3d4nU+9zSNWwjf7nUXhA2yJRlR
Xs9me0N7nGKs1m4efLMcGT/pC9Z9AVJqJWW8QcX9hRF76j5qQa3ugGfUabdYlQqX
QpOll515pAXhzZz1L+AGP/QrKkEUKp978k3NZcqCZfJlS7Ys7ihLCsZqGOC2okFf
zswA9HECMVandP1ZUQeD0DUGgAVd0oXAsSuyqmuDkWi3yJv4xSrhlqhy4nEHbTPB
/hOrH06ADHILI0sBig8HHOUshdwbTv4J/IvcLMXkhGIlYDuTk5cJlE0+0MQLSCMQ
UfAGRd6T5j+4NKouddvLOW/Jr77qE1Kjn+sTnsN61MCKSW8qoRha/zjZYw9D9Qt+
/OYCqjOJMpPV2w+uPT1ApfcyYsIl97jYZRY6zoq1/R0ZNgk/oFdij+5JjNjc/yJM
iiuZ+YRXVmumaXQyogFdGWCCO5/dT2f9UCksC2DEf6s=
`protect END_PROTECTED
