`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PrOD0Ub2GiMs4Ep38b1beofTG/+ddy6Yo+MP2Y8d47bqzlxmPQe24RK50uKOC9o7
dCcg9XnQioysvA0ujeeE/9lBWGDrGLFPqs44b6gfGb1ETN2gCjAtDZlfk74/lhx2
2hyj0HcfYq8/4+kVOEAssRjL6/7d7JAZzC6g26R76FAm59lQJjhFGjpOCatX19W6
OIfWTyKxoLAMlB9qz+8wUMOwA9ATY5mevwuvAnEANR8EY36S9Ac8kv6r0HxZ/7EL
tNso7mBg3xgQDsY5Ywvgm7xW5BXtRPx8LW98LZMmtksbnJu+nzMu7ET7O2fovcnk
hAVZ1D5FEc/hDSx3obIGfPNZoM4TCSG0QOl4QhVq4YjCe9H5Js1aUj3+is2aBsQ/
dfN0PKjavQiyep1IrFDpUZlxpL/jDwhECT71zWNVNNsfjscAaJx49eMu0xU6JRpz
dKLnwq9vluBPs3b2fsaFuq/rArLFAIgSX1n4QGEUWYYl9TmEJq/BkltkPe5pWqqP
kRps7F0lSU2673x1RXaOYo9H+E44o2sn2bg4ROCNmicoA4j2YFLdarElQxgV2kiK
GNjYFSQwVatBjatZx4LZ0XxcUcY/Fxqi+jVZel+J7bMZ8BUbqMtGh4M7znZ/bfBX
5RKI+pNJIF/gCf3U0lrZzy0BjTNWq0RcNvNIcSB5Vssj0h/v4yURUReWTczn0+dJ
icXxMKviUmYsK+g4b4fSvHhctaSM84eZGkXTAIkCji/UGlVkPYywngvFtPMs/aeE
AQuqXZovz4yyDN3fl4ljNQmRSS4NpAfOWNDoSP/YcT38asBMNsJFgGPdF1DH72tH
g3lv9WTq1qiGKlUHCW18THKt7ehw2aKE11ILGPXQXCwb8VOrbNf3SvcqLIiazCP7
WSC5FlrjKswmlpNjyFdOh2x1rNPIVcGZCxCWWhAIO5yN2DQQn4uZJRXxiX1wRKP3
E0tE0hN6YV+TeocjktLxFkTKQFhlQauSX45Ivn1DsJkiZ/LUbnRThViTiwzCdqxi
SF/Mm8xv0cFexudohtmQpXU0behTcS3kSbMzixaETrfaeEqh8tSGBg5I0BCuxFMC
RGX1Wm/bpN4aROqZHOV9IFPKAYJwcNJi3H5YGZ9AYOR/3SyAwte/EYxiyUJj2iQQ
bcawZ98NbcN+INDtCWe5MRuxLHKitFWxn6EeuRh9v2E2F9nNt+C9Z3eG/5rX0Yhw
JaSuHCAdguheFP7yZxkJcysnw1ez2ogM9tWEBHIWr+S8OYPbz6ddJA6J8gmYEqgv
q351XinY9TCOfYs7lnWTHFkJ8CFRf5WG6fYbl6CooNUAlS7XjKXd8Jd+MwvaNol1
a29F0Q9nCcPFk6MFvPrXF3IfySYMDquP+7OzfjXDyrb9rnhs8vJNTuwUrvapnlEf
ciMhkWMvadlBB+4hx3xxHjj6tdh2J6gpsiOTQcCtlsgCoQSqUf47jryNFeuWMZfg
ak2/qnUQ5VEwbGLsgUxZT3nhhfNpyepVS/LsvnR4t0MP+caUD5fZ2/+1GmOlZ5ZS
5+u3QbOTamTl6U4iTWrMSMSIBPKGn6E/S+2r8f429NRESzSc1wB/iXGCPint0+z9
Fb72DiFL2aHB2nXd6moH54kuWcVK6MHtiOn/2gHV445LK1+6+Wbd8VzFQu//qTpY
hZpMogg89EyytFC4rMY8GqAXwMYDUjYqOAf/VM3VwTznInzqHOtZ1LZVOiSjUS61
GsC/mdoNmMWCDJzZo5NKCO4YvmzK5dZrQ1FdsA4YV8FgUc6ipJhUX8TuLpN/9FMY
2g6SkE/oq3kTcsLGxs/4OIaWjzXgR9fr3pPO8sFqoekHLvKVKgqbLc9GcsuQsgE4
Tehb/aCeVdaqlFBELroTqgZv9ZPMXGX2e0ARh9GZ51U=
`protect END_PROTECTED
