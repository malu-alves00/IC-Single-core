`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YUvv0InKqtyMuNZam8AbCBkW9mxfon4hicQqfs/RcayXtuSBgvZr6l3qp/ll4lH7
THF87JxXeeH1uQ5Yn4J7sQHa/lKNgHLRoHhoyJTQ3BvOxA6Ny/WLLoZhRq6/pYP9
JDch5ZO8xPGt9xnqR40OQ6gzhMnO+pLa+fcGatWXZqpSfQa5Ipy43M5BVDdUgLLM
aeMSLwIOgvmzcpiemkvvkPWCYEIryv7T/7FqTV6fVlz3WU80lo7F3onR+cLYHAbV
nvOAm83WuwRqO2i3ffKOVClrWlWGtiqkY55DJjsya/163C7ndJpMBVNRE5fr0aJe
+5Od+xfOamuJlK4H4UFbegG2rEAwoTVWQQ6Mimte8DiH52XVbFL4RN5Ccr0RQN70
2YSth14TOltKHbfd0lNEKJCZoJtUcY8v7uUvZ8oFtSv3reA7df3dEit3QdYKjmg3
06I3jHCQoiITEwcJCwHLphz6y5uzhih7NDrZ/4NpUragsQxUbW6drjG7aLR/QtCw
EIcSw0oxDHT98CbhuxnHaa0rCkb0XQCzN89Vzy37djpahTnIsIyjweN3KlUMtaKE
EtEMKc3C3WWbyVrEA+ca7NWZjXBrth7UsyEaY0NRN6yJGU/v5b86IBoh1Uke+52o
CifVojEZvggfEczl6F/N9QR1Bd8XR/HJENdx6ha2GSZ6cRdUQRnr0E24ebOJxczd
5ZWacpmgmnzq/cwqkkXiUevJzPPHSqn6Lmw1XwfBxRX7Wb9ctQoH1jFlFHyXeLkr
2t+ObVTBAZ1g4cpQsZrAaxUzh7gEGBTNaXV/jY1KGRHeddmpL3d/C7tpwNB39zzi
QjRipWOWtqmvi8wFAwIz41weEB/6DyBcG9c+95gU87mZRgeXPAkH13QgPeXO/JJj
JPMkwk/KBUrvZx2Isbfs7pHR5HDo1BX8nKAQrDqSFgyItBYHS60fQ5XeReiBEotC
/y2H/1QsWgY9f1wjFal0zJZ1TBkun7olaJCgoHHJeY0ST2X/LIv0WPdfC0R+TGeP
cYC8kzY4fIwyXUW3uhO0UZ2xCt9NJq6vsZN/dJfhHk4HUaR1xWf4pcM8/EpgIxpG
/3x+r6hnXg3Nc7OF59ziDeUklku3oheJDhDRdny3RODHIxtgVguNfSkOg3VnOheL
kYhAsrfNIGFYTh5/XKDANJyXxSi6busqitPEs797iXI7gNvhZnyypZnB08ezfYlL
bhCJnMyflYZr/FGvJ2E9T2aiYdm5e1VtwbUAP0NWiFlfnAmCuKbJ5h9uSRag/+P+
TN86YZsjHJHljJ55QoUbCKl2ZZdINo+re847b4TY8XlYRpRWPATJTbBWVR/seHjS
kdExCOEHUuuScL297kN15mDof9+zQbkgOKTzMwqmUwvzRcfeCQohDu3TAhqnkyhb
iL85NkRnwak0FIc2AiX9eHSuEqYNo484+gCbx7W76+v/lnMHQiUrXQDRarOnMiwY
IaEuegnjx2E6CNIn/8WLbhSyQ54vKMCfaYTNc8jnwefYMfvWBDbUOyTF1OQ+r4U6
9PUzAw2DC/8izIMEw5+yzwgEsWDxAG1FC4OhlcIoBPFe6SBWSQ8WPe1HnMqtjY9P
/pNQbvxmxkD78L5BJl7yn6YyCA5uZIqbtbUnCjgyjhBiFcFwgj7Ev0jzSj0ncaMq
Obd3zc4lgiXUxpPACNnh3W6LjYnARHc4MDocWsKuWTgX4AzNFq9vYe+4QBE+FKW2
`protect END_PROTECTED
