`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
s+zyv49hhPTeVCle5KIaofBrzR/mo6hyFnC4m3hnpeIFBeDeDfkQmCRB5nNzCAhi
MBoxPmChkEt624yf5B5IR+CLlpqaGRsGMJhc4BFKax+o7lPlutYKuTRXxdGQmmKa
qVMiQxTbl9MG0VS3B93KxiTKfHO9u6NKQP0r3XB6QwPj/T0aDlWV2xHFM122mi9d
4oWAsyvpzQfqhUNWfzkY9kTXiZWydUHQyzIKFFvg6Jc7BT+GrPJ90roUNmIwkMcT
VMiYvglLgkgPGlxfs/l+9em8l78TgYNtyx2ioziXqlow6whTJE4rmah3fwI4fHDX
SRVDVgLuZ7tR8CBAGpgv/fvAWU7Ao0BNrb3i5KWHBAO3s27z2vAG7qpeJg0y+1Lm
nKZLQcjjA+YCboFj2zYYw7ynTpLGbr6JGCjUBo3p5XWtXJZRn8XjLK99QwcXmMFZ
UgZJxAMlGzA9/1sUOE9OA4tC0JKWOgSKNSJE2Nj0BxZltIjiyUfsDh8ufnCBGVyv
Pgq1qk9fUUGIfI8aFe/42VWVuAb0yFsZITWZXw/Q4R+x2MaD9PHpAtd+fDjukImy
UqX2j1fc05zF3uR0faBb8VFfKvJSDhfycNSOePUTrdZ1Xaknhq8hlQibcSkXRol3
MBC2niNPLOlFnGdNs1OysCtmzt9a5+SzUCyF1MDWL+/ZzeRkjy4tV/JynhiILMMg
5xRaA7dq6xE89eFLx/LogCxfbcbJRNX/whB+S/IdjJsElFT4GcshTKOMKzaY9QWx
IGnEedwta8iK7U0QSgxpcP+9FTgripoSnLA2ADxRQHmyvEFGqTXiI/xlXwGpgMyG
R9GScjr3IF8eYjuJLEpDdNRjUjj01D3ZGM2ONbDWlPxnEZ5lDNCD/WPAAukAmxWa
z4TtXLvQN96gXOMm4lAfLDv7h1GSZ5lGbFeCwMJBzsAAnsVWieAyGPh7kxwFtQxc
jo+fO1VlosBfDDT9xfxyRctqzACJNHS3TTqzAQliL8tOJffR4/6zgR6fZHa1vnea
qGJz4a4Xk4KYMLB17hDf5YblIl4cxAszHEzgHX2hxj2QEfmSgtALi2rg3q99aVJy
wQIkKa9hQhxhWrAV0zzKiyfjkSGmKEaIASM9e3lli6RPKhzNJ0BQGAqtFli4Isg3
OYrnbN/0ovq8g7IJYUpaMWqN+08nFtwBt5KYZmxH68fu2n26SSAbMRqvesH7l2JU
Xiu+qbqBcOO6dbX8Yjc+YQ==
`protect END_PROTECTED
