`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XGHalJQw6Tr77JYM6hnZBzDyDdpa6U6BhZ7fHVsHl9w79lA9rTSXLjEdDGHq+Mlg
At8FmrYNEiACGcF5Bo3hqpRlCghh6DGsBPp2gB/R6vxj3C2xlGCh/rum4kPD6g4f
dAUy1ZprVTDefM4mjFMlMNAh0lpw9P+MgBM2CNdMFpVoGrk/+h25FW24eB/dWXcR
veXywV29ON8UQj6o32Uv+cA0uF1zbtw5vDdQR1oUWxiBWmXLvgF6AmfUvo0b4O6Y
ZGUlGxCfPdemYp3Xohf3UoFblSlON13+yhs3W3H+etEmI/hO7KdGraf0NBzsa6/w
OmbdZyz7eDryMwt7dXgcBPwig8TM9pdu5L+ZAni3Z05OjM9pvrJ0wnq/cisURqw5
e7u8cGbQjAsj8KyaZ4rRdfzx/W8wy41FA+fjrUcjWRtqqGiuHgYGwUCf8LURyqtC
9hxy5cHIQ4ZA/uluLC5PXjI3QMs27Fi+Cgmk+H9PIcTgFJSNsJCnYNNlZMWAW6TR
0xmj8oaSROBhDc+MzsUrTioCXrmOpz5eyYgFrvJEQYM=
`protect END_PROTECTED
