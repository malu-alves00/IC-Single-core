`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2s1fg1fw3+q7XDz2Fxcb9CIskdtM1HxvOKiR4+W0BmUb9p/grn8o7eqdalCchxo6
9NgLTrxZjR9Nx0RA9/EP9iCbKTglVl2ZxUqvV605K6FV6HWtlEmf++tylpp2RxSw
xaLLqM8RRA7gUwV3ZWQDicI8xM450HhbAQkRH366NilCEDsAvdHjEwYMlVB8b2/f
HPS28uXbMwVniaDDXiNPUOCwUGJfCzEUS1xyKmPGfU5n90cS5bGYFEpzuTDRDxyD
UNnbVAiL9jUZA0vBMu1bwgwyMnamdhX+SfSmYfJXsTXblRakdqkl8w3c6ffM7xiy
1ufrLk4Ci9bo6wAsZXDsJYghBv8y231Jn326SZhgOSfTZxpZRTHCheH+bJU8Wjwr
yfXz3gl996FeGcClvrv0ruw14fzEWS0uv+UXMJTIvMTkl5BDDca7wU/ZWYmHQRPc
qKy0KEQR8QBf04cfyHSMZOeYm9vlUV97C7Oby5/TJ2RDH01rm3gEzRDFbas298SH
mm2xwHbhP06TMyU6hbmB2X7RKgWvsS/rDvTr6OWHxtdaeh5KiiR+8c1qehE000tl
V/XDUCdnFsL7R6O8qzMyohvhI5bRkhuSI1cDRnDrFUzxzxswz4TNHzHNABfKbFGD
Q5BhoOdF2qfu/EU4qUcHxFjEfIxKGW/yGRfMEXUau7BchxR4jJ3xp7Mp+MHGsssi
HkvphVf1kyPw3CxFOiZDvchzVUWpYukTOzSN+IkwLlUgckewF+RNza1Yr76wTReS
RrmSQxsgT6jJBgPp/xXSZQ==
`protect END_PROTECTED
