`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2d7CV4ZeIF66OpoL7Bvfeawo66LUoZbZ5bNIHezBei2+Au0aJbFjHqAaE/GIT4MJ
2s/cg1OXaGRTj16i3mVx59dVZ9azxfs45kYHWhgNGroTaKwC2tcbzycS5ZEnXttl
YMRjkurJqq2FbxOzrwQ6nD35mfaa5+XW0ikb1AkxS91noHWBhrVdx3q0mCoeM3OF
wxpMNy2lDbj4QZw8Gf/TEDFGmtlHMTfszrHsnSiZFmvtVZ+gJMYzDG0AYrl70Z5r
ltnBRGdUsFdmysAeJPSA+8h4wFu9mvYTH1AYzL8Nbj5emHy9HhZYNdsb5VKL3G0o
PnBUS5lm2o8n6POp6aCR/sWydcuRT5PrhH+gd+5vqiBqGIoz57x/zSG1faNfVg6p
4LNwOyFnXW9M9LYo2vVw06Cj+0Aiq89WQRtKWs72FrPZ6f3tczXiUDfjL51HOaKH
P1ZJeSFm5n3xZZjbI4T3j/SE2BVjKpI28yB8MWOis1IpzQRVzm0tjz78rztRBq1b
Yq52M4NYCpweYYwpcOWMT7ij6zzpMu86deuTx/To1MNRuLaCre9OomkkNVSQyfy0
7wR8r1AGHoK9hCCc+/t0LY5IIRYXBjCdm6rHPhE9pHyts9OaEBEH6vv70IIATNxW
6mpYOOamPnyWtcVNkv4IDzN/rGaqoSIrAnkoRoEd0veCUngXzr0rn/hPdyweW8C9
+gb/gVFsJgofkcVvEPrs18ApC9WcS+QXyap6z2X0Po49s22+yxeK+pi/f3xAmk3k
C630dOoRoemchGQ3a4PaJA==
`protect END_PROTECTED
