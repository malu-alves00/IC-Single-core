`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Pj6w+73MvN75wuQ9C8qrYla8LBhhqNhuaoehRsRAoxnerbysrseLZA9pPKmQk6LD
GteRR1XC/GVm5u31ssd7CheJEbOT8qznhm8cxv5p3vgKXjcuxUIAmX35Zsz9LmlO
Q+z/KumAA9iUEi2BWfQq4dCDL0JwnsWRieIgGw1Z0qKQ6qjW+sGOVfKOtYS2RLvY
8mwPfFa4OA6YqxENaAuyFOC00Y28MUayTeR0KURhVDKHBaw8I2ehfItJTffhK6+L
rnJDn0c00StT0I3Ith1sEna96eFK3N8cEE9w6WA44Q0PWL41rYwGUgjpHSTEn+FL
2WSKluDUGXVolnLi4R8HF03HG4WbnHewUOLqGpnIYHBfz8k5vmI329Qlr12xxP1V
o0yVZ6aaRf4nN/sQtIzC508yPTCXFbSL3YKP2WNgbBtiG1nSY6Ej4eOw+mIS5rBy
YsP9V1+M0tTT4v5AAK6VQlsIWP/cjuaneIo23/2N+6HpliB2vJxP7g4pyuP2lZPH
vblDU/TSUwabozkM+P2WJe2vO5M0MMub5WY9qZIfXHNjeID8dK/KQzCxv5RBNqCL
c2mnmseyO12MQKhri+9S8A==
`protect END_PROTECTED
