`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
G1WEU9i4Ct5IvykqtJXTouuIYBsn9vhmnjaOKxE6MWwukMsSDyMNJWDwj/KLgG+2
0IaC9sZRr4fV4sOxVPSuN9Bp+aZDw0aoaEHawYJRHlumcW+UBg7pQFkrTaDjI+Wx
dCEEUlEhu64qXZLMk+kkLlzyCkXbNCtx77VhRROeSUn7vV5KK1yl+SD9749oCH8Z
NgzPMKwBLKGHkIWzeYH9dlz8E+JHGtFR4/RRZRvIaWDn2jZd+arSu6jPOz4dFvZF
ZmyuBeZW1sTl+enpwDYTq09em87TZI8nynemMyKZPYCG+py43MTuVFfCHR5SziCC
fKIRl4okkV0y1PA+BuWzX9mu0KPSsPHt7x740Jf19pWQ7sOWkXz7emmzry0/EuB0
99mpU/taFh8awgAgFGFqWoxkVeUWEBp/XJ8ClYb1qpGaXSHZcf9Y9sD6DAmv1ubN
Lf3iZ1QdSzXOkKGEo7sPEo2EfQPRa5eaIC1gaO2kxccwQGnJTfDg51KkG0CXNnbe
cEO3XAIGo4lw7/DQcgeShfdKvWLa1b51Qtv//6li9iyasTe+AtC/R8SD7wPGN2Gm
AtaelxxgCW0Nxjkq6G5AX93WEouW+uUTQsC7wCOaSGclo2covWYlMmQVdqc07ZkJ
ocKb3+vxCLGuEJN70KW3s56D9JW2lXD/MYX4r7S0VcYHNC+RMEF4Pav+nCttIBlW
EEjj8sKiaIZZRYClMH0tqiTC0xroEYZJstOucvJHzM2wQBdTR6JoBSckN5WGYulx
rd2P3+xsONSkqrhNjagpepPOayP0yg3S+1omq6TWHWPF5fx9jMTmvsTK6xhzZe0p
5jw+ocqnPIZRK1W3kgBOTyT01u3G9CVCVKIGHT23dPYqQQVLzplZHkyY7g1vqkg9
pTrqqd5RaO+5POqNtuYshBFTRV/a1Kk7UK/LB4wokKOzYY5H0kCrY7gcB/RUjnOM
Xp1XA44O8uy09r18tfTUrfiTLDzt85oUIBdOZ9yME2/g8g+Els56AHyLb8UvW0Z3
uob/IIklQVQB/NRLXcGY8TAVCVD6wd0AId+tU3sw7eTnTfH2trZnQIoA3Z6Xm2+Y
PGLhllJJLnOguB2lSa1G8WYObyCoJXygbhubhNtjNL8j0Egw6B2Ezehlx/F73yOt
H1gEGy3wVovq2O63kQLOic9JMiXBNd5iZtcaRUguIb3DqJqvU4PrB76DKYVpdyim
KWORqvIKaumDGJuF5SfzjvsRSraV88ubN0hPktQUqQG6w/c/AhmVSEtAtE+TlGku
DZV1D1vk6vTFPtTItCW8ihESDOvCBc1XIukLValWf9d3sbr9pNkw/lRslBikTlTR
b2X3YB+HyRzJ07WOmChxRLQyXK5wvwttGcG5K4Ffal6OY8kNzNPF14QT/bXIBllU
eaLonQp5O+afgGTaoDcdWdwa3OTNWheWsPEF64NltBs4QwFsdxD533HxPuyEZd18
0x5f8rk6GLiGVSE6E6fXksu4dly92hy1+gQYu2cRfHyOiKF+OFgKdGYk985hX0MF
uC3WL6xxU1xYXGo5y7NEeJ0+WZDIYJMueoyvnLBUTU4BJfxPIZGjqDapF1SCMXda
H7B+JXHErttfIT9ZThzilrhYARTsUSlAvYv3ebkx7POYMuEH0bCKk81wBuu6CwV6
98qMkInhBR6qvkveYtoZwM++gKKWJ+UAvIq6u783mXcgYzEKFgpuNA1g/g6LpQ4i
pgTol1zQwm7Ll0T0tQHez8b+SxZ9u4R3oIDzL2bEafMQN0VT5lXC6Yu14WBYxJy0
SiCsvIxWefnPJkiQYNu1sf6Afxn/gJLWEiAzq3yYNRQl73JFWzgVE4imjpT1HikE
1PPJ3FbMVrH3fymF6aXd0bdV8+OL9TVAfnGZE2d7EOWP5yF+ELbnwKLyHSQv+9h7
bbzXhinfahc3Jj48Kie2s7sWierKldvxBQ1Yb4tcOQO54l9HHuCu1t9ikXzB4ZmQ
cTgxDDu2bgDxcQtbTLCj4jKWoze2VlqVnPQusOfMNyI5VFDb/RVvZc1VcTBC+MlY
PYgU4zaU7NFAUZl0LdVFUGJbAbz1qZxlphr1eKN1caA02N/sCmADbYHR+jTiapjz
UHcwAsSxzYOihlkfM1/lf1RTVAtU0Umu5+AqzOiwfuwapM13hggIPY68Vsm6/1DA
jCgP4HzREGW6FTny0NDNXbvBinmIC6kTbsWXBr4irfqDxN09gnDRm1WcCqcwcoyr
1GCTffF3neMXLdj53F6gGgbdJV3qDNE5lRye14NAUKmuA2Be3iIYeKufIEZhgj19
DpyD8S3ZXG+ntwdrYS3vimNF65uuQCDKN0KzbBHWBiD4AE7Rr3VZouV/W8SME0/j
6GX3OUkZg8n5/Q5rNWNJa1/PeHgWniLIljqXFdprG66MZTNAsWYUBLPnAzkOTi2M
XNaujfbAsY81HR6hBsPOqThK+jw//WhZckmcppup+pSNyQd+QHxtuQHemBohPxdj
okF1XO5QRGc+enakkcsal2gZbG5kpaXNyjd7MjhYvjxA9/WPM2TBw7t0Ia2b7CZN
QoVQ5ms/Z2sUwP+EuGfHvH/TAWiDeIAmLJ1Pe5qaJVt6EiJM+OG5rZdJoYvYLTsK
EfndvTL5BVWg8EN4d92VVdRztSyU2gAIZLFcTSTxRmmyxvyIqOtrmct06BQNXUQ7
I3Fc+VemaIVd0b9Hk5z4kQ/rTsP6bcWlrxfMvwfAfd21A842/GD6cqPQgiPvy8k2
lFq/6kSbDXVvRRAmBpPgIJ9qlOm2eCTNnQIpxqvhS1ZltgSah5eVxiZSLtslVCB0
fmvX7B6sZ7qy3NoDOOAosuIe/3ywJPiVJmjST2H5WiLfdPx6URtZCBqgBjr+1U/O
nw58TtLXrprKHE9gq2r6DQYdO3inChc2zHAp1D9yF1Kq8FkjojTaszEE1sxWvLEm
+WT/lLedKMWZzSj3/2xaayjNHjquEH3EtdUoi3/m4E+wP42XiK4RoqtSAEdlTgO4
NlQvFdPyioHN1x7XH/jy6FMAhXCsyaxVVFgmjrRYWk0KP4sypNIm0BeBp15qqeqp
CkDD8p5cgYPqEnmnfbdoq7FVa5hYJpRV+weFvxCNuLB3MdenLUPnQDpqjsKjfrlJ
glRXlA/ITh8hNRC8ps+ez/yVOaOOTJ1ywmFLde/YpbuYVAX3pZGzV2x6hHDGsUH7
avuEIK6hlxfKvf3elAxWLXfUpTMycmjVftm1TLa/gEoEXjMSsgTzgPeLsaFNmtkJ
RuxdhpKFk5Lm7aD0tGsPD2m4YzS6YyJPSVtWP70uh2BwExpwknErPu39GimcjKYA
byPsQotMRsm2/y6O7TH8IvrkzdyCyMlcJgGn4zKeImMQjUOV//6jAT4P67GAlUHQ
YeJLQAvLfQ3bmrJSUInS+IjhG64xT4dZxijgWL/CBZO24v5ssFPBOY8j3FgRKBlu
CVvWWbl1r6Mneh4vP81nzw4r8I2ds61RUqJ3hSsZaC9dEEczdDASn/kv6J+2JIrJ
B54Z759VBgl/Me+Vx4CAG+oF5PLgU/x63qLyEfllsb1ECTahrV1hCj8iIXuhQTDP
J0C9qjHN1AW+eWUqaUOVE2lYaufv6Hm6GW8i8ybW2NRzTU7jOp/m687peUs6r0No
PyJaEZuDd1q9+2EA/Gz9gUTDdggTkqrKjBDMgzOewLOkYdNP6iByXm4rm1PU1Tuk
kGh25U79+skPim5o2fjFN7ihwzn+N+p3w9DI76mQB6aA0MkNGK2hKDiAUctmTFA+
Fapil2Igy3ZOon9MEkxFj6NGD5Pv26iTF74WL6JuWCHugeGz2TybxzwwJTXbg7H0
rDECHKspxqJXIgym+yhVWkv+96IYoUBbZkyHU14kXQIEXtDKasQJRcGTYR4alSHl
ysBpezFjn0NHZatkB8EEmJlyDfoDSB2ylrtWmyMqvJoTRVZRd5pg5Ope8lZ19w9j
r0pKeRBcmkjmA/10MEUIhyFQJ1R5eaL9Qm2BS+sEaL1tIJBR2QqGc+r2a70SJmDY
QugN58h1tn/PPDJsFEDRUffBNg8CwfEuza5eoMCmvID1iWO9k0raMYQFoCmZh2/T
njZ/xhsPtfm4pCuFH2Wv0MqWdjwsgF9BUBWlugQI0MzfdTlKfePmA8ZKPMogb/ZP
o5U+yjy8YzavnFg+8t47bl8Ou57ffVzbjkkQB1jK2SaVVt1mg8ZZh9Se9l7eJhiw
3GN3qDIAKI3MZZVJrfcSMfmWziFKtbyWO/1zJ57elI27iAdb4dK6CtzFSM3p2EX3
itZzAzKbVRjdY1WOBxz5zPRxVS+QKbwyWY0ost2uORSnOppYB7/Fbhf1YCvjzis5
qrv4xYTw/iCSwmC1iTniL0PwTiE//1hoL/EjoUjD0wZsTetsRAztJoWn23pz+hy1
Gt7wKUvmC+lybf+wBEYVg/teVL+Oj68/6OsqE8G/GnnRTMTYDMjL0dC0hL/jInht
T6Qto3qNCihkgE/HRteYD3fbLMwYRPiBHqzOWmyBZN2M+znQkeiugz/EeGQPV6Un
R1wUFKrIfIRN29VHyLOaYpHIrwVbXYNSyCpfyBQad7cyDUirwLmK7YnW6e2rSQOy
YIax9Z/84w1AQvLZgyu8hPYOCwIJrXfDAnTnU2/8nibFY8ExexbBysnjgCh0e297
IWUX8jS/ps94XoGPOcUpiZaCarwsYSlfZ/bUjmaIfZV5DmqjQuC7BHHpv+XXpxcP
GfMWGIa6VZV8fLa7uASWrRks58LztKCruYsCpSFZtQUsd5SuUGLFDG/2KalbHmZj
DfxkAsUA8/htCx458tihD3fZxddp39kHYoarUBqPQxgKHSsWlf9PQXF5nYwi1WcR
L3a1iLpyOG2ZWgsjGd0XSsfH+3bnei/94LqZO5dE4fE/bjgCftVyBg+bvQ39QT19
2Aj9wqNQ+hWXoisn3UX4x5Rk2pwcIr4mgkUHRWhJJCUClG3Jsy9NttYCWa7PD5Y7
uMFo60R2cyb1nIfaIq8eMcX2tiFEKd0ZTxsd0J23P6wXCFkgqVmcL6e8b2IvfJ5a
31GyiBEDoIQKM2RIpCYC7CD6VmzI2x7Fbcq8jV4iT3Fr6FWjd83Hjx+Vji1nmQsV
s7ZmKhHsmv5BGtMWgpyNVxsHj8YGhEgBOFL2k6MdgirBVZlyLPkwBKaW7SNbMdqL
Qn/kuQfPlqy1v/M4gk5PCLvUNMhqTzu6uxwvUaIi+uZ6uE36fl2W0dXl1l5Igvx9
nZvkxiHoBUrGxvjnPDVcPyRYoEAfjfM2P1qmGb2849a+yytxkbQ6m+P+jHVKZlDL
+TKkx/eeFVhxnb/wIKdSDqeKiG2d9n3DkITST/jbOPv3XzfGphY8eq3zbr3gRmjL
AP/b26/WgkNTZBWwjYOIntoe8lbf59chlAkfDSMahIfEeAnyciY/zc8VCar0C/+E
mLwh+UwfJ68Z9rFl22xY9CxoUDHCEKefmDp8N539oRooPG7IJFZ0qDAKWb9Anqq/
2/rwI7dGvnHid67rcOJS44FR/XK89DZyX+5PZnwX842T+c6qaKffNRfVuRHunvk/
ME5R4LNI/Hv0WtjCCcSPF08JIxekwugWRPBUzv3WZKqHjlwKv90Hxr4ZQKPGftjF
7tDrnejoeHPc31IBdYIb3BrdFXIqDJtwPbwtEvK4/kTjPuILk9fgb9bt0kRxRjic
5gtso4YUTCTVl3vXR+A4iZiSSW/E3byuyOBy58mpm7nS7Bw5RTSiVuQdQbIAnuKi
+XVznyYZ93TfPxci262nETFZvYLLZVtIijOwlyXnuUmrzZhUV9ZUN8UIwmbMxTNL
9xVMnqOv2zJmwIbDLu27KX72vrocSP0JQyj8QIYujUErKG3LlFvoniJ5CshHlrLx
qiKRg+l/gPZhpzSpHoakEQOtEOhr3e9dbv2nmXH78NBOBNiPwzkCXCRJ/v/RUKT6
fiAj22IJA+r0Hwl/Rx5oFeciKirAn2cZyrSdV9xIu3oFwNp/fA0sb5hvFlMt3iHU
3V9sxFk7xCLq9cY7G76/e3Mm8jiOQRNjh78zbQeerZtNgfmEI9RnDkLWqS9cWBSW
isKkR0kdFW5XX6cKk9Z6PgSBwg+XJnG4h4tUhgk3xaBQYaQhvyzPgKL+V9x3o+74
KZI6/NG6pc4Lix0oJ9XC9/yHsWAMXhHxkHpB7zS10S0cKZUFN2XuByWdjuL8dyyO
hFW8nhmSdZYFf1LtZJqhfoXhG4KhtzSxTqYFtmdvACsSlN7EaACgtcxV0tXpiBhc
mUCF2uqQaxy8M7cr6JI8CGithsJT9ntkLfYMkm+piYhbz6Gwj5mSa+l8pDA+rpIk
e9UNcM3hUhO+UAtD1vRzshfIcEBFtEEnRtnlah9nhfLQAN5WPYeyZM6Wm+IO/feT
8ohfIiFAaSog8u8Fw/VkMbNZ4NbTyhYgYep1jnEM/dptsgUL8XkCG+O9XceIsqFX
K8wO4H+zUQrF+cKMGYWruZWGoghga94B/DGSwHyuRroevzHyilsYblY/OPwkSY7m
+a+4ne4fUlgr8Jt3XdocYPLlE7S3E3dVsHeBmwdwxAccJoo8QtbHOk3rsIIghdwO
kCFBkSQBPD0VvQxP63wHywnH45OjoUe7jKfh7eJqFvpe10E7yS9k16nBVXYUFvdk
7wrOfswAaMOZfvjtXlwzxPZzWGBklbo0y91J6scEvEgc+np23H9GP7zkBC7sxOC9
BgIibonoVhLKKs06yUZyccf4a/r1/ONjq0yBYO+1kgVTHjIkWy9n2INzv/IGf2o/
Vx6GeJDLTbk4jYkCG3QTYAXf/kD/iMeQcanaN+fsyF/akOk0x4NC5ZetF0VqTmE8
b0edoFyF6EZJvJkd1EtM8wndNofGeqI8XRRuesCJ5/4NEqnun8RhJRFt3HVVWl0/
WmMwLKihl9i+tRlFLusQDNNV3R+nzOnO688cztUIhptvdW2TpX2k3lpurEc8mOsm
N9h6rGEUNHcU9dqvwSfoY4z0I3JXB5Re79LjTup4mQOy6YYZaB8x63tJ7g1TUSdJ
e2YVU1zHOav1ZzA2zerFfsN9LdB4IMMzdIsGJMC3L8fWAhFHBpl4JaqOWcvVbu0G
/h0OnBVAWI7dR35tM3Kp1ziBVHkXNx6uDoP07BsbgNxOze+qKUKBf1PJw0zhCuS0
2EQgXZTOlDnP+C3IlpaBkC9sx2sDpsUJfVbMgzbCDSYv5SvNb+rkyAtI4uRAkIiZ
mzkC+XWCGtDUxn9DxyXHJHvFqb1qpkP0NYI/mrwbi3lvjjIQpZ3IX7oPM7FjEMqQ
q6YgUvoWrjyLE7ZQpMwRIFLcxCbqaxogV211zdZiSlByXN7UsJzuQNSrsPeGNj1M
b2LnGbRit4IciTDNpsiGCUqgtuX23iSQFolTT8zkb/KMbsamxBv9YxtkfitehMHL
9ZJdE4nLQ7YiQ1jf7BfPNB1NJpp0W2ZUnEgSnky4cOFdTrArtA2cfpkYsys8DtMr
TipQS+cqo4QmcdO838vfgPPba94bxKZ1MtxuJeSCNQs98X6iWwasfiXXF2tRFhV1
cin9WFO8iqgQwOgDJDb0vR6ablI8qwLSCxLNT5LaD0ESpph4wBRgMnhGtXcS91FI
GlIBVFu4goi4aLm3PYS+5wm/b9L8caSEHTsitmbvAD3kA2XzHJKfJ7/sPK8A263R
CN2VqSLVREMt2/redzGvmPHQeOvQb47yWHaWUEx6gyNtaKZo7x6quPqgq3rvKw8+
t4MmiOj2zlhNAh6JN/Ld/1VMzRJBoYu2qqR5fb19ldcW0K+VgAB45l5kM/OjPAY2
iDrLbkKGF6jt45NKkOykbq/J98UCLU0tN+Vs9QVLY87D75aKj3zwcgV83mZoZ717
d0q6GzZby3x9m+HnVe5gSTr5U0hvQq2uYRvZNzWVa+HF1UU4GyHGZvyM0aXo/V1D
qWTA3mM+omWJSEnadj1Il6LBVl+hlW0jGeV+C61Wxu7x0cGFxmLc4ADKDmcSpgr0
3QM30ZEHAh7JLAofl6HB5vIIur/BZjuh02/l31t3Fudm1BBS27NlRMgYhOj6i/pg
3IJ4yC5x46TD2Ct/CPGYnzrpXAQxk5vHN+eLeov38oSgJ9rgOfC3HqdUU/r58ILi
izdPNoKOR7jdzliQsOmNWmduj9sqPDI/Twz0fqzq7tPLLO9ERzd3LOJK29hhQLXg
fyQHV5AOG9WMC04Ik7lNjXDoUixGvg1dlsuEDQIEk/cYYm4ftZ/hANZV4GcEagXz
/FtNIOvAhSBhZv4tB32Pf6lwFcDrvsTYBVMTh/orDPl6SAQuaIhP19X9MIrGKAg2
R/fSmK3w8BmVrdwJ8LiEZQ6v4v2OBv8Bp/+IdYcn+61Juhc5nEGy6zaVnWqR72sk
0HraFIbgbINN0tu+G51ZsUBmoWbvpMeAjxZ1MIN7jMTwYdntDIIYQMtsnTfiXLUT
2G9jUuGVAfN3p8osvTpzMV+0Memo84YSKB0FGIBOMRSoRJ0JgPvfwBowOblxJXm0
hSFxrQvtwuILO1VU4HsktG2YVYI/NubIJbz+/9cKdINr8NFxapuKHBOqQmiEvbRT
YAsdqzv1K2S8QQKoTY6eHU9c4tiE/mBHOHbRv607K2EVa3Wn4K6FdkS+Cwe6mb7b
4r1AG2Ig2k78trNW7cn8LW5VYlzd8xhQHJxkb2Ut8H9CSLX7b6qNTzJeNBYP/nF3
Fdw7S9kUdwFNHgIn4PgIctaxU4R8cxrL6DbAK3xIvtvx6DO+urCyixIfJJbrjEUk
4Smkk8jnwrqTMBhr9z09NJPd239nTMJW9HMXMpH8IpsdLBEUs5bI5eg5WoIjN9OO
1iVYaij8GeAA8t3wV6+Nn726SGa7zcgGniKnqgIjwdyBnluxBu3f0qNZVkert/LJ
RfwBuDhqh3PEGHcuHqD0HBPvsd8irqxU0g5nf6qmbFj9x5qMNI6XSq8hkX4uszhR
yG1dOHwQatYbd0TTy1iiTTS4BuQlJB1MozEL4oukEcnnnFvaVTLb9D4zG4Hr51AD
nNaqe/mamshyoVPEg0bbNAtL09a4H7QxzRzg7UmoFJRbPaOJJE8kY63QoUqH8RK+
tuCt/KolN6eFgwQt3O5a61T5NpUA9iJ09pqz16OT/IBAagoy4WrvrdqWpzOlA277
rd0M0tpJOy493xExxCuOfSaEP3JEUW2o4NPFkYfzF2MyjYmNy7ysUya52ofEjDdm
3otJiMjV5A5WBfV8y5z0QC86J+LyjYoApcWZLSTG5OWT4zKBs9U2Y2uZyA1xQ9He
+rqEvSuP2fK2Gl5nq6m8ktHMFYSAGmTTX27Z5s/8vfUrBsBMztAxBbDbHM5x+Ucz
OmbAvgaPiDyd8MBtxn/K3eid6Ui8UxQeWiBtUIJsibNSafhyXvXOO3GhbUn9BCRu
0x34+xMQ3Hv0k/uB1Dj4Q3r+kEmgzLGp5+2SW5I+QgBo+WLUoOQokS2reP9wk2Fc
mUHvSI74wI9IrRhEqmzepmUHsN6XRlyjWD7lhQG6WIyNNFLtpGZBuz6I32lnMuIR
WQA/dC+4gqW3BSUjc9j9Z0Nv6vHyv3Fbwr754/eUSSnBE7etb2bMf9kUUtniDCCN
AlyClnmiWLKb5NRo2jpegNUlb++7V4+k+e2AoZ1dlPPTQnbPlnGnP1mtLiibx/2u
ThsSkn7mhyVGmN8ufiviGXmoy34Aa0pwX7RO67jqSkD2pyM3v+/ZG31SdrA06VlA
U675TlLg6uoWmGs+X7euNFpPmxuLhMO03/hhzTpOG0u2u/DwFhXJeyYYWw9WbXMD
q1mMRvjojN5kYJcDiOUkHGSzyxsXSeEIeUfyEOFCCSf21uvmBjdWdfEFjEchjCeu
wEZajvEYDYx6rGdHk2ArodSEUiRry0x+Oebu/jRADP/5ceu7afZNk6GBL+LNqTgP
RvXW4IOfpWkYpV5oAgKlqGlbTw6/MQ/so9VzETf5xGTo/zOSTwbDuHkZW7l28fnD
WCqzE4/jC7qN8IkJmhGhsKq5KNnOeGhCSy1Y3afSTFBN6pdHFIKc9ffNXUo5UdCJ
sqNh+4nJM0N2XTh875kXChj8cEuyGBbrGafV4mTy4DtmNHBB+qjDE+PSd3Qk/3BD
fo6QEOnqR2JEnOtEbh5mKFCuRu8GLRSDVSczON/GEuKyRHaA2lf7x5FhTHy32MsG
cDVI85mhYinZ8PcmOPv/5Aw6ZMw9yeANm0BsEMwIVbSEXlGO7K7pGp+jIpb5Y3zu
JErie2nmKg4rdwO18l+QCNkx/HFsSO1wpn2fFbMU0rZsRe46YFh3XedtyunFHWdd
YVwi9WZ8KEfcKJqmKL/GYSMOGqKn96TkPZq4QRUNL6/WrAif+/5k1OOnSj4/ZqMM
k4l5+66++Mu0YZ6Q1TUE0SibUXAGzhTgweun9YGc/MlI7XQ6c+Co+Qv8Yzzof2k9
i1Jnrfm0hyo61MdCWHUFGrFBEOrqquvDPlAClp9FNTGYWdOzCcaYqwjrcfczPNmk
R9+i+imXKG+oHce7YF+06psHlxtf73BXalLg3Nj5L9bg/inRWEFxRaCW6THzF4ws
Fe3KRiABXsr+dLgsTT6DV0VJqbr0129Runx6yvc6CvoaPZe1xPQSPOeXJds52D6a
jFO4D8fiPzPR7lWlIBH54E0EyTKgDy7Ny1NPJFaKVLEOMhDQvP3A9dspR/uFD06m
ELKko8BVNi2KIq52QNuVcI3HRJ7oIvLZEwlviceZ4nwLrrU0Zv3TZBXp37fOzbxf
OBdDh9iT1Nz/CJ/sJE7oJ2dtoS+ETpqEy1T3npoxgpcKlQGHraNZNQDDe/u/7Kaf
pe39xTti6Po0jVwarOHU2FXDkg9T3643uc7TCeXv5aUnveYQiqBFOtCs/O4YnVKB
tHIpMr6YVaw82FbGCW1MbQCUc6K6gmNblbQMF6FKX/xc3ZqtkE1LOEVsu8gDox/m
gYhR9+LOEXbu2wnfCmaQmszmORuC4gp1Wq8z/gcoc+UHF+7CObFC1PEwLi/k28C4
5AvHuD1OHQbeUOLNGJYTpV1/TdVeMpXAU4NwW8YLDCboXBaYB+F9SsPsX4P5QPI7
VQZUTwOEo0DJTxz/dagjisiB/5FQ2ZW0/LHqRE4V0QBbNJPmsdGby2cP0uJoqkuR
A6B2YaFcFtKI+mbTGyTR5hom5ZZGoB1uSgwcPLbDND3ii4l0XRrDD+apn6J9x50f
SvYlW+hsGHCFLTzk6tK5y7OFyMhkjxcAe1cy052klmzM1FvsTDOEZWkMC4WwZnub
c+y73I0yrKGdDBidWfDM2ohmJCYjvqBpmsCTJFmlqAKZ8MFJIoc5EgvocCki2M2g
LZfX/nir3I/UUrd06I1am0I8TomxzvRPj31O2wiuBbflyh56TL5bURLGpzdGlAXv
woHXK4Hhjc2SwqhbeMhLpF/uHwSdjssCMOBjbpoH5poFiy2wbpH1FbYiaLkc1qWk
fPE9YHLWPBWgX0VGNxzZl9VDq/DL/lR1LCuScuy78/nUNlnL3WAWe82QCUS3wpTi
CKH/2kSz2Ch2U00jdyawO+nDCNSbmwPDb6fU6Rjr1XPdwpsYt6sTJ7GcHJ7tHrQ1
/BY/e6c5H8IblRCp51OAlpIViscO82FbsM4Oh2NF4+RbsNVHaTqnCIUhnq6svEAJ
CwEOT6fgI0Mdyqn8xWLtOV/qOhTLRWOHahJXfL+4jiA76Gvq09px2ozP8zJbWC8s
s6DGdJJp9CdDcd0RXT94Mo4kHEuSUMHMvwQ9DPtP1kg2T/Zvwn+JlkpHwNq6u9bV
GrmtMm+tltGcvbk+/HblIHZBKQ6R9TYjG/41GPzwV3f45p7KJZ3eLrLEIzIEJBq+
d2MpCBoJnvkt0PzUdr6eQEn5DCROnZH75JRY4YrhbYTwZ1P3TJserPqL2dNeXihp
k2HMiLVn0kug1ueGDf45MBmkAfzEwSX/E7Y40M6PZzGMY+nLUNBjwh25X1DWdEMI
riMnA5WlSk9Jopqgn4jNDWabYUonqOgfMkLf//ELc/crQxhbvtspt9vvySJcPZf6
U9UCtw/PqnbYKQsyyp4OYAjiPB3Eqb9iR5jYm5OReaUGnQffPU8m4IA7BUnzBUb5
VQw11Nr0/ywbQ3MjzZnGBMXVbeQbo2TgI9LTqsC0vKFK2fk8GwFH7ZOw1Ck0y6s/
Za1QcaTd7aMcvhpE5gLIQ5WfJAIN0xC0B/WUQ9jkEmtts3G6K8UtSkANxohICmSl
71/HzD0xWL5rd4EIavrpg6zcLgtSbWYPE21q5wWRxgmpaHH6m6e5oQtNRp/HdOnl
YddmplO/x4fxh9ISkiA2kaqMDZcbz4/4E1FyENjqCjSG9TdzdRMAmcpi4V8/kTcC
EACzm/wb/FF0wRcGPX/RAi7DEdCv0MhgdOg9rOLFa4FGjV3h+MlRQoqXkEoRRhaI
ddkcrTiAjW4sjyuODJHRHgdvWgB5AYytqgUOLlx9JF9qWWc7f29vNc6J6iEYCMcM
38SmlvT7jgv7c/6mpgaPWVCTL0yV6IeKlIzb3fRPOiBZrPin4agfC3hphwrsa6UG
PkWp7dEHzNoQ0TYol+iPtNDJohBha44T9FefFdnx2kItL0YSUKQJBwVLPJIpnUKB
LKvyrny4r/H/lVH+F1JVJ1hqGGB/GBeqAaueV6j0hh0dPNdBfQpKqSdORdEhnh1q
r7dFqjeBfhR3ITLo69t/x/e82fBxfGIGPVhUnQkW+J8w7RqAUAqV5iBlqH1CECsB
/W7Dtp+0N+usFK87tOff1cT++LQf6rroFSokHCVFnmMP0ulght4zcDD0KmX8Agpa
CdSDth7nbvxKoFihJ8+hjLsTpyqOFN1lXNcXv5V43yBXO/MUcdXMa9klYbqr2QnA
Hh1qIADxxIninY1tdPOho8L7UC9wssYpr9aj5LgQrlB0rw9r1mAHUB8sLp0uVszo
Lnq5c/JxJt3c5Kxbp23g+Oj+E9FiFONVo8yHKnZOKppy4WVksO3PGHBr4mJSRzeA
X9qZDQcu2CqRZu0PQyd9yKeuszL3qoHYdzRVZxGeKo86NKhy2lnP0cxI8MkGYiI7
aOrbt9DRDLDkwp6MEvBzdjLzmNCfEjkGv9FYpO+YaNHLO6qcS4xFYu02nVUq52rD
RTTyrnMxYozx+a+ET7Dkcux/t/Th7/JPGNRSGBHouPzoIya+WRWuv0IoKLq6M0EY
SDIgJxCAYo3WgMRLjZ9gCNysFYwBnLcIjIZRoCHoSg+VtdrZ+4+OUmOPvT4Vm6MK
AY8GoLDuqAub1KD3yHAsj7OKp1D6AauoeM/Zw9kZ4zY=
`protect END_PROTECTED
