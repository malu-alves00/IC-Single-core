`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dkLa1MWS3NqudM92zQtMkI8hYq7BsKKzLW0mYxEop+mFVgXi1IXc4spb8tO15OWM
QzZm7sooVx3HE2BH/ptuKoeoq3taTBpb4uBxGjrcU+SmFeoXlrTX289VsJqR8/Jq
UqZAjQkn7/PzHmz8BXh86YK82nPa3hbZ8AMc/O+x4a/VGN1FiRUJQ9f4YjqWWduJ
GP2/udFrVhhia2LLaORsomu62A47zc7jfiqiAgHdUUzjgik4R5wSF64SU5zLfwJx
mjbU9PqMM2p1A9uf8MzMarw2xkFiC01uVM8fdm6dSvZo5f1TjYzInkZ7mfD7tmoW
2TrOIVhgLvGz9tkjIBbTWWMrHaKSRhirX+bpiqM72vlwDwMCiYukO27bbTq30ZJn
UKqG1wdcMtaBQ/pVPuqkNq4XjfYPMLKyW+oTZEKTzzvXyrEKwV+I9sIV8OXhDn1g
w1xQ0GkeLzqmjzSd/ds9fT789VsKv4fjwsoETe7CqoNADzXd6yzTZwR+uXs2OctJ
0V5FpzwGyiNuwCv5GYaPxDXdUysXnLiDYq+3untoS7C8JVjec09QmY3moXBifUSA
b+kT7R0sDDP/UY9JqAQLEqMVgUMtQYeNUbiR6eGIdguG/ONVyeUFeWm7lxNUqVNY
`protect END_PROTECTED
