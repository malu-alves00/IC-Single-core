`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RyeWgaav9k6aSnqzu1NIrHVfTubUmCtuvV4ZdoYRdGn5RqmIRSwKL9AVXmTZ5GvG
UbESrNKL6RgAJ4IphDFo2BfwSt3hPH/pBuB+RZNeqV4UaWd0zXKtBSAQLOxrhnig
NzUJUqKJXDQf6qwmYy+7w1S2e/kb8QTp3QhTgvYFmf5Yy6D19I04hIZHBWD5uS0l
Ye/BRI+A7Xd3oN1+tGf4aQ5Vn26140x11wkLJM+4XYlCcmW+NBDHMQnvcgEm6VBY
HgonbCb8pixXlio5cjuxdH+8bwEr1t6t3enEoifUi5QIvvmRHAKR4l3Xgg3MNgoO
5G00nXp+F1uCL4hFOj1JtiVMMJ9Usc2V0JrnsyaA87NYY0jkI4eT9JbUlYX2MmDQ
xzX1V8qarqAx0pQpe+dpJ7gNwZjBNlFPI5n/rX77SSck+RELFs2fFf9AZoZ1LKDU
bQsUPLRN9wzEpnMt+0NDmq7IiLXVQ1NDzWkngLEv3UXLIiu8Gi5agRm07/0jObHN
xpoUhV2O1Zt9qnblgaaDzm+Pi4qMDLzAdSZwaV5wg0hwt9BdVQqwKVC8DZ1hl3lR
cBneso5M2SN1dlsHZ/9igfE+GmjaFFrhVxHBsxj3OvE5dASmeEoUP+aGwujNQEeF
EM9f1AtW0UvAx8+o2FmeIIP3yhzM0VRuCgnJm4LVHEHCv3KD7nYjnJ8iWPikNeDA
VMqHIo7Ny5miqGwnwT3XzJpKwuqPxzSYCZbGpz4dFEDtmL+6Qbp8GrSdAdEGaWpy
BJd1NvnPC4aWNlMY0VBmDD1nX5dnIBkhUCS4QlshGeYW3G3NKUbE/0CZ9Ydf3+s1
3Y61riDYMvO9ZUjvE4alP77n/YW9HZQt7Ws3L37nV0en+rUJN3Oj5qD8UuzUJUUs
fiygRQeUaN+etJQNk9F2vzlvCcW6oNNJxjqkEDoj//I8u4zOOvYCXYHcnQAF+1PB
sghi1nx8nBR2X5UYgNyGe8B5KcwwwWS7ZX/82IAfADgcZFZfdLv8PYQx96WFnW5K
rJd0OTVobBnk0lYT4EwtsF9wSDgZ+DuiAinOqW1q33Xp2frja0f0whTe/n+22okg
UqcIRDsaXduMzRoDLlkt/63jGYd5MSUlE/SeOk+U/Kk1h3fr0IeH5ajMn+U/Fun2
TB9ZUmd8JP3k76z+vxrZ8CcbQ/WMWIXC70IrNw0d2UKWxkl/y9MliXi20eDs6oGy
vjmWZnzCDOJstynXBk3eJregJaec6pZiQG0pW/t9IzYIoVp3b33ENGtsqhvyllx8
+WFdUm6nclk7ck6EQfJg5oUmCVZ3c1oeVsnGK5CjiJm+IIxW5Lt2vNm+lJjP0aDA
0nDdo9YgGjavWyWyJ09HHLvB3sUUx1XAskHsYgPJq+Z5p6jsjDSCrYWkGWPJe1xJ
bG3I+5ry4LRjOj5EUJP2Hf+nX+Zjog8bWSB0pi2eRZtQvh80ub4sih6OqfmjtOOU
`protect END_PROTECTED
