`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
d7c+0O8rIa6cAGtNl6Uj9lmmadilhc6Vah6UgPXHRq9AhM0qa6C7ePx+yd4he6Ks
LChDBhnMFZC5iZCFXp2L6k+LkVpPg82/S+bNwS/dlKuvyPnQZgsnRRHhWsOmLxLD
FFS9Jpwq/LtC2w2uPH3BZWNIDxuXNnVM35qfBaatnCXu35RZu4wHs+WM5+geBV3l
JVzV46cDtYOiIZ6P1Z1xlYzuNa1JH8sjDWr2JXkfQHRyrEo5b8iUoLURmBaEY50l
jSZnnIW3KUZKeE/XD/bIbC9IrQwDdSePftWX2OEtf5RITn7FIL+orlKRGI6rbqgI
jXDYTBionOXWbsrB+xzwkbGnefczrArz/9PuUMMyv+8kkZOh54LmPEa3gdGXJ7ul
Xq9XRMVeZYJE/P6BI2IYDYzRBfmex2MtREaFDmBVrdAr0QhAWFWd7GlK6WpuC21C
OZbBTDeY6GGWh7PS7WZXdw/9Ou+lDmCHOT6XlDWf7fhB/e3uhoym/2VwRtW/fBaB
fIkjijuMh7mBsAMeol6kBWLHmlfTkrf/OUm3ooegpOIqDwIA0xVD+/oxu0RhCANI
3JYLIF4yr6Q/8EL+Qr7HzQ/zo328U74Nu4RUBYv08jVhWoBqBMGjl9FhbH2z/W0b
8RP55Iwf//OBE0w4P43kaQO0tjCmzgeHJlnleaYDqlN4gpl7BSOiJggcPSmsGKLl
zPMs0R7h8s2U/CvkkqAB9UanY9dvGVNiQe8GnmzjQTz1Y2BYY64QbhASa7KvC4eR
LXv8PhKtmyZEc2lYAylNL9I/bUnr81wJB3XGI971Q3q2fbr+f+pjP4XEOsWmXMDY
lYacwp35Cppmm1nfz/oroUDX0b/61f//RPJCGdwNp7mFBBv4m2592pLldNXlUYU7
EO+1XqfBqM8KJnmNfZ06StV7u3nF8FDVHXu2muL4jLUuUz0CFR2HlS51pRrb1UoL
QFPN2P4zEx7NEHFCvxafePTNoZLT2Pa8lrj2GHn3T/9fZ+SYVB197jT/quZW+Jbn
JuT8yXtYxV2oAAsVALjWiXjAo2NitGHWdKygqq4G9XbRXF/uJOvUgJMQDwikgB7O
VX9Au4gvYjlSo623fzEPUu05T60XKND4NKparZlMAM14DOdCcQty7JBAhRW+CSdK
PE734m1s5FOUxfu2bESIkjCWwmQzQOXcQDGMjRtJI/uDw+lZYx0tRHZeyipEK0Sa
a50IGWCZeVtfdt7upbxfecsX+WM/i8HCutvYvwAt2iPnr2h/4bPXtoF6ohaxWGAJ
QANdMBLCnkJKravKdiB5rkGW2NSSDaMB4Q6iN9sQA0W+l2c4kKcFkdcTwKEWW7d9
NJ5ETUa/TZpaV/i14fdxaWgj/MqUt1Rn6FPPe/23UNbFRV8bpqUlbai3ifJ+riCc
2rmtUT/56JO7setFuLOnwnJIjs6pOXd4M/E68zu84XJJsXaol/1Qa8Pc874kwyni
vtRM/9r+FYOHIutd+mBa6XbNW5ABSioNj5whwzW5sBOGaReMIDAEQQkIWUacwpGy
voSdxDeomd5YE8w2dufDCg==
`protect END_PROTECTED
