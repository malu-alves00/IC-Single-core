`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fZtzYWMss4L31Domta855z5itpQDLKNJG0oWhyiIk+1W2lxxe3dG4eHrui6D5ZIl
FMoHuRkS7ismVIx83/KbIgF7gXA64wucYzQUqLkHnpUsJxMc9ZCoL1Syx/rNdjzi
qindBeFE3kpjJHjXvnjHi2P2YMcrjQ4Vrzf4tPQhW7qWRV2qQMFA82tJTWzVQJpJ
rL+O2bQ3TvsnpM4tnuDN3+JQo8VyYEaQ5TwFDCSzkzTGru1hO1gVbf+DLJ4/K4uE
kJxj+GoCUtnadVpnQMSo1FYVE/sDsqX7fjRpPOpUX66eSdoD5CNlDdBA7wNLEJ7c
dgzhFAT4wPaRUocWUBVQdGPu7foJ1sVCmC8aSX81sX+pJ4etV6Y1ccLa5QLAGYi9
Ttz+0XBGl9/Mw1SmPodAOjPVFS4q86n0HWPeKdaZBI00STj23RC8Ih5xgYqm/nUi
8uCvkx4nyCu5OJ0aTVHdP0NOfg5vUaC1eMYb8PQ8VYk1SZJ3LyAMSJmVGfpvEg11
MU2mf6o68AH50BCYZWBO7PoG6nrM8+u+i3MyrU3uWpc+q7Ksl6SL5P90cAawMaYB
elRwu57LIWl72MCL8vOZdxhEIOvlEPu39LnTeW+DvqHjvl8vtTmcxjot0u4roEF3
ae8Ddcbg/JQ0OM+ocG6sFiWzORr+/MBjXWyjF4JjZWOw6h4o4U4q3kMEM7NO622O
Rdh3kSJdAJY9YixGrupK9gsvwI1yDLNvVuLXQsQnF7LD8iYtF1In/19FOPkm/fWP
51uxsOktRuWGbecnZ+vBJqVFLnbSaP6oFs9ACrgnpmjmKS5IIBXyVEtVbsMac5LL
zadaY0G3fWE/rw4Sp+ViDYng9Dtf6NBVLEecROyWgz/xiDP9YRZU8m2EqwvrDtwn
fGOtHv936F33dDY715zENLOAHLff9Nm/UGBL16Ed1TG9/aF6oavBLT8ZlxeoA/hy
ViOhHprM3eb015C7cm1mEiqLKTOt2omX06eEbyp5VAyvwz/hVZbg3un0/IUTy+Vl
NbfyrYdF8UEQRQY99vcu6fW8uKMfXrMoXmM47lph/0E7ygjsnVBClak2HL9uKfEB
3xFRRpajPZgSM311+0eiAPy8bZtBCff+p7YgIcIBrBtP6QxQsdATDfi/IVy5Cm9Y
Rt77vPcmsjnaYs/uEXVu2olnxYbcf2RuhOg9QohEkqr4f011W8G2zkImt/cWzvn0
DIZT3fSrU6/639xIVKbS8aEC6noDf9bhrmMwZ7Gx1Fkvpks0QJWU1nnqHgFPsBIE
XPoZGbLWRnUI+OH0ayQno0ikvhvLUsAPWPOMnvd7b2Fz0OIp50msNE8rjn7IFSlX
ti/EbfdsTZt5VKFiIjYlvMLuNmxn46Q4Gy02p6SmayHA9f6yaegqEEf+3R1tpO1w
jTRW+Iu3xyn3YgH6fdlii5M01DMH8ZT2RShieO4lWtOdnyyRNL7uA3OYQaLBYIx0
ae08YSmOSAtbtqG861anT1n/bCPCiSkj4GJAhJ4jQSOWG05wUXzMx+mqQIXoZmvb
dwLaqoMKskbIHiJxUsrW/GVKJigIABtQpMs+618LSD1j1p4rRVtzTsFdt3kHC9Yd
heGnl9LySx21PudbC/fkSvPHtv0fCFfRgayHKlDm2y1UBoSDZmbVq2ifOtcN61P3
DVe1r6BthzBfofaToo+AIKO/LKPsXFposIeV7lanEJD09i+zZf1euHixbD6ojDkw
qs3dR+Rl2hLuAC0bImNpBdkt7lUKvaRc0SgkCExLVsT3OsfGUeWm3V28N8ffU4i3
dptHDig7onWUWH8Tc3buhrUDl81XayUh6WcppxHpgRzB8nriJwx6q1fAWs2jIKaf
uyJyBP4WNADyZj7nqIrLY3rOuhO8we+RLmFOFkF1KnOPDpdzNetnSgydHyBoADvs
qp5Nva9fFA1Hzuo5ybPX6U79s34b/cf3/OBisDC577yPepnW+eh/WliEqwEQBdtM
P3by3zJxG1EiKSiTw1t7orUdUJaa6wl/b0ILlZEBqaqDGtbmvqTuQHhqh0+U3qht
Kpt66vtaOOuQv6IhstJbIP5iBxn3VyDru9odQBtZuoz9ACXcy5m2gYNwp3nQHL9j
WPm2NhEnnn3LMMZlAB3C3c+gwkei065O5gbv2jIo0mlr2+G1Xi9mr9GKYp/nyHeM
MMj7kmztYuvxMySYjgfD7afy1Uu+cK6U+jp5oYSH6d+g6mNvYjIq6Vj1JIjgkg4Q
ZA0CxgyckBXCNw6kMtGKqDqS8pUzcaooQxQGvTo46EUrs5somTOLp7HDX2xIjjbU
sJgq8Z7RZSoB+IcPcHS+8oJbnhKVkFj/WUB+7+ZIpQdrUfikfAepYcxa2EJy4kJw
cU+0/vRhWqrT1Q+VQDEYmLixjvmKOnhj7MjWe75GWxzOVBobUp1PoHLgxGupf/AX
QJRuQ9lpDE6FU9fBF2f7z8ArISNb/GavGyuxffeUh2QCx6QU1jKulBnckYEvyXj7
g0UOWegJc+7P8onvpBXln3+bwxfVRDez3sPc7XXEV3tx6Ddp+qlGfJU8IN+ma/4d
cIo3mXUM6u/5t2y50Q3YZ2pLvV0BekeRtdWil5la2W2HpJVlv1BQKZqHfdd9VJ2g
CuE791qTnArhQqpY8CB0+A==
`protect END_PROTECTED
