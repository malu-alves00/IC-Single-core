`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
t1o4fJe9qnUe9M35gsxb4t5ml2U6DeXsLKb8kDL/l1s0YnrmHGCRUn/HqElF8cHD
L1YXsryiQE3rSqDsFbf9/QG/xUwa4UBA1OqMW7m94OjTA9+ublVrcS9MrXfnsMEI
n5W1++2RIbrD6kcnqIp4YkbeX+Ucor065um7N7PZfGKdFbWEx2xImXGlVSwCE/t8
h73oWMok4cGv5P9iWPCX4mLSSpYgS86mDSC/aXugbRkEW06nNVkXTjr8YoLB0ozg
8nG2sZhePGATs8t3Z2hxIxagfi84vlyqpeDKxhIb/sYMq3vWzhq7nUixJYrA+YRR
pGpp4CYXdPZzD84100ewVGtngG+tQUFkPV7mxDoDGYiLaEBcSqwE0LZ2hC2sEKzj
AjtRGIW3948/dqHVH87wZ6B2hqOw7kW/4u7EQaKZ9MBPJy2MYHnCzvI8rGBTPUc6
VQOMUopP7DwrD6YNgLygDfE+3C66Lmcgy+3jfqxq44Cxk7EYLMDwHYlKeJLktxPF
bkfBihQBVwy33rb2/xeAttprhD1j75x3Hg7/x9A7zDUBRJsjB0twZvHeS9Hvyq1w
y00yHobRmhs/XV0ljlvmanDL7OH3uZXf5nMUCu5joX8=
`protect END_PROTECTED
