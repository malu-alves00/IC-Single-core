`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
d2f0W52031ndwK42/l5MxzjQKeXw56emwSW8olH+DYmiVrhGlZAd+/EH0QfOxMxw
lodfaa9dgBiJTJH10FfX34ggln4q9vwqoWX7hrA7brmh/HC6P46bLn3GJwqG0vBT
1F06KSxXcWroyOhfLY6Sp5cnXpYhztVEbJLASoCR0eC9Xl+oUq86m9p4nvxCPo1z
Yxf7F2TzWe8InDXUBucqRQRDvqX0qUWnpYevQ6KNOb0jxt4XfLrUKUzGeLANU5mh
moPOJT6HanFc3hYZUURnh3dG4/OM1Vphx2+FbXCj3l64IixebK0WFYEiFMqc4r/7
l0rvSU9CAgr+n4NtFbJvIWdw5kn/s4kHVmIiqDx0gtcAEkyJ/EmxgbidX+vFt0CG
w7eFJUvATWCIhMaVEqsHean2YvGmYH0AcULVEm1Y/N9xyMUqOLeL7SM7/3hJqoMZ
X7qqnL2k0blJ5O6ZPq2jMz5/HJpDFq9WYwNCNXYif//Enm5KDz4IFMEUzKwPQnRr
OXdaeDlw+i8D1oJFTafPuau+z1fLDhFl93T231vgGRHaH1IC3nJH2T82tCMMHADU
POcoJi1hePyvzHvRdW69hzr2Sggq4UBaR47Y7rnXUG5jI2u92JAq8bhZQvSmp/kJ
NLEwI00xSWvJKOFll/KM3S7xllMr3zUAfn+K71msXHNwpL6BtuwbvERyvU+HyPR4
FufoxTiCVpeQ7kBehS4+qrVccDwji7nUKddMSEgEpDGya4rB/6NsThxxl5juregT
nkmRiL6wZr9jideFND5PLoKg1oc5C5arOfl/QtgosCg0UBC8zhZs3JrwUA50SMGG
DF1h/riEQSVj4xKXFjQ6aQxHwuSoWKnSnWvHtrFSoNfyAaJIT1QaYWL978JKdzJH
SyGVye6TLx3YwdEhLYaA+mBQ05gzxtdxxtOC8Ukv1PoS+SjRMGs7BT1FfPoyylyq
JW+eTLKDc/bbhkOVJrWvO5iYtZFt2ojJuiAfifUjlqiSF8u6BTeImCc6R/pPJSvz
uXSkge3lJBeP6CzB/niipQGIsfP2ntZXgV/SxxXhT6qm+0Ozt4lME36HFgR5efDg
egz0z9JJrtJZ1f5c+zfG/rwRm6Wvzw8XcE75XJZo4MZoPOdKgUYpa90KR5wEa9EE
VgpJv3ok25UTqWPUMwNk358gXY66I+QcGv7O7dEOgUjXdcVJgW2Nl3YPNvsRUu3s
NKS48YlEmI4ZIrr0kUN6KyCT/4dvBbP0fh/d90db+DT5vPO0z4ofWc8u5HpF7WZG
0sfVfHb9wIonDUBaNDV2LWWK7OO2et14YgrYHlbQy5CaRBPQg87i+aRd/oBxpZw5
dS3vT2D8dgQPvOAy6xAwWKGFtbs4JCu1BxJaQkE4hFv5eMZ3cN7jfq1z5jXYdb9v
gOuSE13HKDH3Xiuif21ZYaRtKN1JWsTfD44NOEZmNcyemaCQObdEesKm7a4eR7Mj
7GeBDq0R4l2FMpbhr5Aw34+v0LYAiiRmEKdVIuZPLBhrmObqONetLSh0aZq/L3PC
w62w7f8QgGagQ5N8FWjKqJy7JH5ZKDq6nyJf8G7U1FHhH07Yj2VyBGuIQasEQZru
4Bjph01k2N/P8ISkx6C2ILyK7Uop3vUyrSzSSBMfYrg/mvIa83Eul8mLilgx5HVG
lb8R8tdRIdWdwffj+ZE4pKeNpFNgUMPsfAzB3gm828EIg+PI06dHyqQEiaTYG7uO
dzTPBceZrJV1qpjqjO90JOSaDxGdwp+ph8BQCHmVBdfOfnmhJ6Hh1D4sAOSXnfcN
LXAKblx++09uutRx4tR/FPUYBiR8Rjlv+JnXTJTkFd7yI1fe5q9+Hqbs77xdaEMH
1izJV9VIR21Rz73BLuhrCNoUK4dUehTFvMBKzy8aROyV2XvFkpx0+hZMmazXSGEM
f625QNHY4xz6Ar7H0G89DJGWHRbFEFm0Ztd0MH3cDeq8UNgEjlfhrzzhK4UkzvHJ
W0fJElIfti/cwVPm2kTFU2L2/1BQt0ba8+3sjFTOnpaPCioh/x+2SCeBq3iKZZDn
fRpJpuuTxGxeOUC9YICD6deB5mNDNjdXqctNQLTpaIqnwdL6/PvGuFVY2PKZviZx
41Zg1nuuECSj2c/cVjova9FsJL2yiYls1mt36c8mk5oa+GEpwui5CFUOhKCM9Kwp
HIJIy0mKv4XFI14ct3e+n0chnseIHCt7jdr0CjtOkda4xEEWzpjpM/ae+ZrdTnM5
ekxQwd1GaVy0x/5bwQxOgI8kOUa8aZsnbt3cEnWq6zzPx0gMVZj8hTlJpI+uzJzu
6Bf3Ftu6wZzrH4tgaqWp4hBq+MPex450s/Zk1ROAgIZdytsksXSLoAZ2vPYHE1iC
vfj7u8htmVRYdGYZ5Yoo8etCo9R/wezSnipao9T9VmCKxzTnVfU9iIwh9l7fuz7I
WH4qvTGUSdgKtlqXyaIpO+Zs7shCYMhUTp78MJfIQqANYaeiS8DvoM75p5pugIbw
Vvp+E3mkHvBh08b1OyzLb90lcOH3gAW1KYWuDzF5A5LG+IeiF9IPLUVsH+yVr/h1
ptua0YnENvBsRgTSRON2/CWcAtIbE4aBWOUPPwd4p4NyEcqjxyNRMKaNJ2N8ojsD
uYOutaoCPBLfCAzbEVJtyr0hi3IlqMOg2FxFkxRucv44pU0XdBCY6oY9edOPpR8A
uCjoigViFqDCW2RixP+ET09e4BSg6uFEFUdx5aTDIwfq9ZUEXrabLZSEb154Qi2e
yEpTD8dSZ08C+6b67CPlXZFdAY8SI6zz5dpX2pnF0OvStMKdMef/KoeCVvhWiymd
9MUwM68MJfR8wbD29PwWrc505HLcPg2zWRTQthfAmZdJLGJ+TsCG2qJmqA7+JH3P
c/BGfuPzRCxsBBdXRTz7M46oRWUc6ndu607Npm2CJt8PoqVV/Fs771vwSAsqPcnZ
5ig5+C2Kd5qb7LxGOHiF/Iw3wjE3Qmq6q3qzjKxFKJE/RipnGSd4ambHl8oRSZJ1
47Fa/tqR60sdr/X8506oye7SYXMvKn9BZbloQeJplTC1GAOeYz7VCJpgotca8kjg
VZXeFifghFCwFMhDl+3DDskYmR8RwdUsXHRhTkms2umHfCZfDG+TOCjUWKOcVdEV
X335tM57oi9/Qe1SMrplSkL8s+BVB5kouZmGX0lSm6aZCitk5+UuC48hm9uWFkaf
N2xsrZeLX+SN+RbFHK1nLslbV7B+EV7Co72Ak+CCVrHywPZrETgw2g89tpgWtPM1
MNWkdWc+/nb3PPNkp6H0gaxVb+TnbJQziGjOquqm/kGNslL9Zyyt97RFch4mogxX
7wvN7VUCpGeLTRAI5vs1VKBlp4bGJy1my5sxncAaZHp/w5L0R658nls7QrpNuELT
BtC3ZnKOHZrbpjOBbA9+lnNszqAH3mFB02UaQ4jEm/0AJSnUWVEoOZmA6SCQpvqL
3sPiTrIUa223wLAML7nvEbAqi53g7ZUAzW+S0Xp1Zgbzle087Hwtug/pDQ05iQa0
NfBOMPajh50J7fZyl9Zwjz+fdkd4baJysExzeCfdVJwTgjpIeToiJ3lxryhnsPzG
cL7nj1y2po2EGMMzXOrcZiCHlvwUA0Y8up8Ho4TlhUvdC6EgMWBjz0jgbByvMb4m
gvgxnkb5Lmx8/I3e1myPWUzCCXORt5Gq/g00Eh/gKqExb/KW4EerlZOvCjW1JQWl
ZakMYyjCbQUl9DzIEJXW0o5FmHRm3JIirvFl8VhJmNmpClZQBYUKr03jZaTsjTKh
CRt0oPn/zDhUfQqkvk3P9AzxQ77d8BtQheQYId5h0IR6xABbKuCd3JP6ljW6c7Ph
VSHjEPAYUbzAt6/BopHvcAjcAeS1xb03TnjV3FG9phdNhfriGOni1Umg3PLrOJ/k
rHKdPWbQqfiKurMJTqxzPdzRkPBV3osvdYzFjAhNa/e//4ODWlvh0fJGwULXR7o8
wsHOW40n6Ur0YRWFSWHamqlnMYMGeX5fhUIcMoM20z3X0eh/8pot7bZfXxPGZQ6h
PydsD6G+irPqzVncYHPRh6a87WqkCSlg3/MhUPSWQnihZBBQP6XjRJ2YY7XD3LEM
FP4iQM522Spg1FiAdKc7+//U+jqpa8+V1sXS0BbsKY1ahIyOdcldNTsCmVMV2MYW
iu9oBPoAuz8LzCzeLSLh2bQ4XtDhJDhQALnO/XGocx5ojqyeGluoo36NwNvIt30Q
sDNNxPKP2BSDAPjBoq7ogWbsKrRw9GyH/0WuKPbwkJK42C7AamIk8j9WGfwlwtBH
OiKE5zgHsJ42lXog/FyMeAAUGwTnqwP9XV9gaPM7Lq3CwDWWjpffRQU2bDQPgR1S
/pz73TIFoJcHNwbIZTqON9ROagJb5fixTe6Jrda1Ag6AIUUrjogKIjc5LG6oYmwQ
okwZ/Fy6d31HYhWVjIKSXpBIkIHnr6YEhXFIf10AubIH40fyTvfCmUZl7QntsaWZ
jZXg2ejKwQ3OYVxjxHKgzdt+sfViE+JprGoKQ5evUOj0jpSypUWyufUEa6pp8UkQ
UdyeFnu1jQ8VVH//KmsXfwoJKpYqopw4rW9xmsX/uaIMU74i9s+o4H1WDJasds3L
Ts8riTNTMhcLTQp4nb4trvbjlolA5TDZ1p8tzPBar0wpUepik0UH4htJpGMaDwrF
oFrxuUs/msOl02W3kzyqAamLeK+tqfcs5f1T9kE/fVZ6kWu7Y/5Q7RAAh5WuxT86
sQqhYfbaIBAYtoiB0aMmAPgVwdrCAwTmiHg6qIUD0OkbBvl930YH+zlgFc3LxSBF
N1GnuS2WRtGYKGSX0TX9k0mgsuTdYx08NIfsU4G/mncCqKjJdrLohZD/AFg++I+C
JYAA/G+UR8w1AaVqWNdn2phHRE4lGVn6Ch8r6AiqsxOQ+Q2/28wXg74buDc7edcb
7rJwGL80QLTKhSkrSV3AIfpVMK/eyduRs0D32vktvy86oXL3TyB1MzUZ7Jdz1HsS
IRfgO3kBYs4XnkcUVvx9fL6EMuzVM6d9gHy3YcC0yI+cU3E6eRlXm/bO2BQCC/s1
6gq922wpQ/azYJ4RloMZZL0lTbvw/ez7IzUPz+9AvdGPsS8Zj+I/lFrq81cmW8D0
NdNfRa6EHl8XlWKdHm3W9AZDwLic2nGePp95sV1Qlw9e1tKeH2hf53WlcWMruLnC
Ruab0viPPZBWkPnBtaMYj+sVaf0WJzTe9SfKt4Tlj9zAujwgbbviQkICISFUnFfM
SubnQyJAM8spPAkt0Q5iuDA7DGz+yJjmizj3B9+Eo15s0GqAUTs9y1qt8B9zbRmu
2xU/LXdnjsbeB3e9y3rNIAmW8jPdCIZDTt4bRn2x884aWmN60Z8dHRB9xbr3Z0jD
WvIuw3s/nZ9Oiq3aec3mJoEre6sHOT+hyE5g2n5d143ezc/N+vbbjZZ5iZuv28Rn
5bfq9VxazgcRS9qaLBr1HViWSETB+D2E7UjsN2lzztC82YuCiYxuhBfT+CKrGMaK
gGq17FPP8AuPwCNcgnHZCZVwaLF3oLH0DjNepZT7aYaFkquT5End5ANOWG8a/+Rz
qgsn5d5u5Jc34nTB1qOwI6f1HUH7Jmz1a9Lrqo0QJccRS3WGeY3U9c+gyR6u1426
F+hcACwUpRpn8jcym4HPns4Qkik49OXa9shvMdM9Ys06awFNgDqXx9aQsRcAhMUB
Ip7GBPWukk78QWTSWrfcuXJwKcfTYmUsikHLt2uENs66GAWNGSR330NKQsBAChDY
Dj2er0y/yCkmAkUHMfWwVCWBL8XiP8KZtjcUw1T3jJtdXT2CQK2/Cw1GNq1hYEbA
HTk8nj5yDL9xgnG0bm65vHE+OcAJCEqWl7o3qVipQB0Kbo1uGpOD2S9mTCbwDWVi
An1cxjQAgAOVPPhweugFiEYIgBYKLVwoSaJDItQx/ExUKKBXUoArE7VLEAeuFWDJ
Os9q4EcYd+LvDrFSb6FkEtu1VsWP9AArUGN6gYlU6QkXWxa8NR5C/ZgU5s2hHU9U
9m6FzNepg/H+C4EtZ+Nt0n/IhwMwVYRRMPK9knzSNkypfrxjvjk7A+trBTBLpM1R
Ick/xtUn+lJu3cREsE5v3o6XH/wCtb1xAxK4hedOR4fOoqX+vCu7eJ2xlc9TM452
IcXXrBTHHTXkEurE+r3uKfx8Sb/RFM1kX5GWlvnqr3IHb1yXyeDYYoojauxBZABL
fc5nRNoB1R6V8GuHiDON9HBFDTkw8o2VRfR5382H6LNyPCAabzvOfMVL6qWASa7F
ch480HvBavBX3dt6GdrX0keuHAPdOqz/fHR3g6vzFDCkne3o0KB4hkeb+UZqoU5m
3tZZPgKoEu5TqG7Ea7ywBpklLnnedIjI3C9IMywKvN7R/OElAGIEiBqoZ2LIciLu
l6MW+cn+7vp4W40S8cq3KROts+7gJ5Ii3RbEVziMnERzLCAUz6sUDeNXgjGb68LH
m9gaeTjqtyJHGmNotPnPO+AVx8sktWGBOH4Ma0ZF9zhUCmVzJMeZfN4pxCsOoSo0
+xIV/0wy1Kr9+/VxDjReoA42RMOKQUS8lXMxcsxttOk5i/1/Gp6C/GgXkTB+M/Ev
UexQtuQ8463tCrEihhGdLtHDRRKoYS2IKsG62ZDBh1cZRc9bwnTpNkHUNV8LbGeB
JouQ5jbjKBisnWZBYb3c8JUKsDcN0Fxj9k/d5CbnvYZzy5m7ZMIFQPPx91gqWX/o
WBiTKBmWNmsuS9Ehkv++8s0kyvglgSfhJvw15VT2Hl6XTKUsA6XGcY5A5OFrbBN+
eULkG20P3NuDmd0y++3A043MjW2gZnW/8tkaQdOEFTk+aPr/DDXCytjRY0jELmsf
hYD5F6Ef8K+JinR0+idwTbqtsGLAefd/bhWP4SHn3KSzXVOJV0tX3rRBegvDHcIB
o2F+5jSaaT+555gqmR2uhZCUy51BHh4fzf0RiI/2R/zH3s5cScUYByLTufxqzx1G
LLXO1nj3B7HTrH3/SzA3XZR2VF3fLndi77ykkR6HvMo/7s/lRJMgHMmXR1wwVLCK
Gzzd8PycKKjGelxxnTtUmn0x31o4Jqc35Z2/ilDQBAAeiFjkDmdbFPxAtMQ9XazD
cCql5tV0De+vfnkSJNrTGU1ufmUsrcZHcZ5wCJsjRoDrPXnmmA3lZ9yE/8lZjuw5
HWNIx/tqCZVNagKzgvYdb91+R/ZQYWmCkjKwkey+8d4F0aPSd10FljAr4uB96L+/
31G+IEXD0Y7hSBvS4Ddrjoo+aNNNpSDQntXla3jXmiLKQgJUyckj8grz15o+nXnE
hrtvE3j9hVePOci+Be5HmqODtlSYsmXa1Mke4rsabH886WNw0nRbbN5kwXGu6qwx
Bf70Q1dfVLtTbs4U1nWXsa+2J4cwUEmvaehE6PKQHbyjL35+F24WWPCJOEBbk1mE
/JDDp2gyuJ+HYeDTWf2wg+L8fke+VxxL+M3s3oMWu+3UX4tHFzJ9J7OJsizikoM4
IjxY1bDdLt6tcYCyeJvDIJLsAgOLEho4JY1EyqCgYzOQ7Hof3XCDMItUCap6iEcr
oQ7pHaPvU46p/iM4ZCobgaZtT3X9NK0EYtzm4bJ/SBw7MZtjMKaFdGf2PKZh0PV6
Sa3oPTbZITNL9JsF+MxibBjdSLjBREOM1ve+f/iimyGTY3WBCjvdTjb2L+YaVD4O
O/Gig+BPuktEHUVxol6wLaZfYyB20hKN3dAdbPUGM3ylUWJA8N3SWgWMjNjhnuWn
WGszQ014sZpZ79lvf286bXGDXUjiyWwKWlf+rREc0ptNP6D0GnTnnDXsnIG2p6Xv
2UqtHKKfF/TZXYjnqkU2sXvwC9qNq4k1YBHKgYTjUAlLXTJm+/5ljomjZmQnn5T2
rn5QyrACL7XRuJeCqTzv5fYTeOHW4Umj0lxfB0uXd57vT6orZoP2FZ/Ffe+Uo8oP
51DGiTfHBrznP54yAWEJn8jlxucg5++uWNsxQq864JlmOa0pT3T85rqszGsWP6CA
jJH2hkphMqVdo9dJMgFddBTiW78am5769kfKxSevy7r625Dhe1X1a4P4Mbr7jiG2
oPHK8Tosi8VlEuGZvd2EE2UhwRRjm4Sfz+uGatNKbGgbYN0YfFwYqnDtELylC89e
6GKG8fz14kXDlAJPZWauE4hYga99pTzaLWSAgsKZAkr8YOpxx/hQdC08hJ1kQuAj
vVj6FaZIXMm7a+lIZDTSiPMZhOgbYnLvVasWuFXca59+1/0zr2zWwREusgRlOo2v
klgEygkzIFFHKYEh/mFewVxtMYZbjwJBD13qTAkRwsjvwdX9ql66LXM58MLfXyUs
wCRjtfbqoHvkJ/d6nAGpMfeOnF2MjrzKAGWuhzGOIwzMLrGEl1YGO804TxVF96Vf
JS0UdUN0Zs38vuH7bI2a5n3ryyyu2gYGDBX+/gbE3jLQ3K7OXCX/gFVNfuOicjAk
C3zemxEhWJVesYRYNI1cWrnQuQF5unDVPP33DRt77nQu8XqfOCzolj++qefVsae3
nw6Xg317muGwelOJWntSW20QcXLaAdINy1f8pLFnql+AV2UlGstuer5iP6H/jyp7
kG2HeMo78rzOty1mjGufhEhxGh9dvkUqemoAgmkXA3m9a4/N7H59W2kBHkEyFrsu
GRBx5Wfpf/LW6cF6i+WtAXzAz+ARycB+WeR4gbziAoY7S4EbtGng6eL5Deqdc6xc
8XTmWKaE+FWflXI42o3TLq7eK9Vq3d/Anl3j3rO9rr5qJP5jru8zpZdBEPVt5U8x
bng3FU1TLkiTyEHLbdM4LI54Q5N1uo477HvS/eIEmTlHNZZlkXSKyizGmRpkwQQt
anCpRTxbVt0Di99W/d90zfi+/I3Yd8DYP9+Xal35HRlwAY7MWOj9xEk10DkdQHOc
1fwPoR8LjEe76s59fjDiXB+qVrjSbeIWyCqIZQx+gYi8G13VvJ3ogwG9W1ITUHF/
DwijL5HFTFXQ0vqU2wqi9WDu4Hqm+C9afSxvm16GWk7P735V1nrFcHEIEslNM3U0
QwiT7i5no19nIFeQOurch7rq8BAeC4KtEb3Q0CUkwNwdh/p9UDguHIU2E7edOR24
oFTZLXYSbmknoUyvUj1LGcx/Aur5OQ+6lr4QNbwfXAGtxb5aGaYSPG8vRixMfOj2
wCGK1jrOHhdnRZD3m89nmC5JkyQMXTnq40Olwphler8h1JrHboza8Fp3rZkm9Hdj
49wEC++7Ao0gktWI4fqd53eKvBg8n/jwonkB+XB5FhBeURlxdWzPPwEk1rRUDnPG
jesFbJHJZx77vcCIzQZgLUYiu4ViAhRAu+hSrtQqd8mBMHE5lYXvo4IvCkWmQEY/
+72hQCPC0IwRZMZU31+2gkZpLxtW6YpSRWBDfe3gVSebp2ikc4jm0BNVFv5qk+K3
IQU+Yl/aS/Aj3wOMMte1J2m69t8nPu7S7j9nfPGXymq4mFkf23JCBA2E4HXLGqVq
7XcsrKF/Zm8fJBaWOeMgfikxZ+guy8Rqov8oFajKLmeZSylvqnvsJdAminwo7mqT
brxUTDXwIsGdWK851Md7xs888B1T2a6n5FhsRbpflwxVC3q4gEeH0Un2FCuxnpBn
33W+ypjTI9V4Da455oykOravNxYBKHmz/8YNgxEFt+nHzeihnL8PZ+y4g5BJAEUR
Bjuuierf+6vNGZlGF7Arfp6QH8vcn9/T/lT0ScSRBvoS3ySiPaO4QpM73eXvdqkl
nA1hii0nbnvryEGfXxOcpKqPjV8Hzwn4CER8RY5ZrnVfnzpMQgHuJonhxKjRRyF6
z1zDyx13jTZ83WAmlycinN1T+UFFaT4pbIpkVjNOepP/BsI9cOTTJS0zsRS07PiT
5xUrEIvWLJfHd0xWggp6GVt4I3Jk3JGa3do2X/bn4rGc6zlgbHmS7AsTs/L+hB23
+W59rT1F4TMo0RrrZr/VX4eq9nErfPOID2/MH6uMo/MiwxKoA8Bv7IANkcwBDlE7
p7e4uwhlL981OFKKHDNhrW0dwtaxKlTqhVXbdadVj4Id7C/4nQNfjIrsE7z94/pz
tFSGFjvViJ9vs4XvIceJisvDROb4Ahhw/c7d+/Z6VsolxLmA4AeMNRXsxJ3A0Afz
CrbWJ8+MMwXGrn6rR2l3whjMMd7SuszuAQSZIoDHjkFEArydYcivmAvnKi2+4tBP
N8u0/DdDrqjkYUb20sgxIamGISSY37gX/8DrocFIqcs/gSAZLBgjgTJpQu45d1OS
fekdzGrvymSP9Tm3N6AjOileXZ9Oq0I1MeadcoiJfHI=
`protect END_PROTECTED
