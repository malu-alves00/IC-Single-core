`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rX04oLmV/tr3oqSq4YbmqH+pC3Rh5dsOptroaMkVZ+dmdSDKG/Xcct7NEH4g8c00
G2QiRCbCiSV+RS4sfSo+94wJVeSjTEBYGKSVKQyo2CqYDWelhsIy+PUnefE1ftcy
8KgXC0Acr3Fxy/YjMDIrpZsar0VcGTSTVSdkwMH1M/g+LYyVIKU4eRd/nOVuz/tw
1+J+pJJ34bYdtXktRkZKf4SrfaSNyZi3nQWULmu4+CbbpwCMfRDR1+2iXSNzsR+M
j9k+TtJwCYkUuTzUAQeOCZ4rz2v0aWZ1lDxtwpObLqv8rOFvLBgF9bsloxxAKYBc
QnStme+0T6L8egBf40MOrXvKOfxatrF+9X4yXV5e/rIzpj2MxkvD7PlsLkKCynVg
UYU07j8qTVOAmURpxzLkB5BgzURZlclg/BtCRW1d2nVENkWs6zIXdu/+0IaKPK4v
18CBdLQO5moFXvdmkkwuulfzWMrAFhnR3FWoZl37dPHVzZbzA/OEDqaAwgYoUBW6
Bqpa+lQ6pzbaMknT7m6cb+2fIxkq5PjYQoKk88+brmM3Rp9l7ivhq7O3N7RCQogR
JKUaz3GKvx72VQx4jtHiOnId5muQYEbMrihN7+i6fqIeodSl6lwEAzii/YQivMgL
W/sHmJfHc5iuD75H2C4II2s8QBRy65V1bzp/fi+WML3RmQlOfsneSdZu+RxoJihC
3JHx1e649XZR/bNh4slOd9hZZAByhBhhAVjZNEoTU4FYk3RGahKO5wbwuUaO276y
SIqpPqaxv5a4MsQxJlQfkA9lfLKrmBkoG4BLni1HIvBs7ro6PYqMN3MJsgxx4x1V
K/0WG7WIanWxuPtwZ3G+LxtjJY9FSDSQjOxviUdKkTusq/yOnOuBLwdVw7+oZ13o
wB66OSdoz/uGDDBGCqYOh5VfxNbKCvyQU8pebGjVdFhbebWdjE1Zt+MxZeXt+0Ik
13A6Je2cyN9ex/P4MwsXByiasMHtSvYU44dIBj75XqDSlgIwCORpZmbkVt4bGZ/w
KXBj74owvVEHIKO/Bk9nf8gxsp7botTWrHVFkGt4slImvbzA+hAfCpvBvorhlgHn
OJdfzeFoeXVff2H5pFJNeqQPRokTH2pM86cP2aaEg1XWjV8mGR2Rn++SwYSQaLWW
SoUbdiw78BSmKWskaHVdYpDiqtoG265tQT+FxAoh2+6ujIgvDQVeMK8aeYVGYBIw
oJGW+qCAAmjz4BPX3PP/gpGFql99/GARXus8aXC3vRgtyzkVgiSaGvGmeZjHn2hv
xLFiG6wPhcMEDj3WsqmgzeZDlhaHT0s9x1V5rep01SziFsON/LoiJiAd99vunALb
hTiQ40/XSH7mKZlhWKx+rPxpAqYjXO17Ip2fDdfqVIu3v69G7wjrt//iIJtTTbby
rxcUw/aM+uaERXyPxOZSXOzbAnZvMv6ThB0sO3WlNN58v8Ob58VMBrDmIgglPcoU
gPPQf84L7SXeXx584bAEroS1kv4TqwFW61JsqRzF7kD2r9eGa6jmT2QDM9KIuk6u
ZSJr6crPGOj8ZOyPbYNgnTBqgjAyJeM+lWu+YMHGlfS/23YEy1jC8OvBFmT4XkUE
lz/kftBdv3HF0sAL+ikJ9bqIP8N7U6iPtfI4tk/SdhXsCffHIdXYG9Ans4bNilcl
iwiZapbuWDaOGm+un995768g8A6Rc90MnVetLBbLKlilORei48sa9/2q9cc6MycU
ZdTbBUWTaBtlsQYcPOib6LGrlFOwreO/IZcQ+yU8JXg=
`protect END_PROTECTED
