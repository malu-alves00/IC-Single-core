`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YAi9Lt1yAadjeK0aF+ufyUbmLh75SLuz+i1vUUct/LzR5Qks6jloI9vipQaGVsCR
JhY+Xs6Zovjpj7DW3qTfYgpk0Fq5p0M4MD15h1jfJypbU2UTI0Wj/KdmAFtAnSMD
Dm4MqZ++eqLuF5JI1KabANTcqQqYmozNBJtjw9MXkqmRNSJTOPOgpvdasK8ics7r
hKKI2q8ayPK8xbs6NvwSu5pfrAdwhdd6f/X78H+vGN6DKtQBUNY07gdHq7+0fWBu
j9dRmMucuJpzWUJAMmul6Z8sJ9DTxuqO0wg/Dl1ot2vzCpjMP0+H5K36RmJ/DMwc
nRqY2kxI6E83W7Js8vEwIUuXwKYqzWhojBmUaHzUkr7QLVxU4DUTIa+rXeVfdGdL
esqsanKk0PWxBjikRjiIx8kcvJmM2rabFJy0WHaA8OMS6TmKARXrVhQkD0Z5G914
+oZz/kog3tqQuNWVFp98rrOoACnW3zQz6BqRdhKQ+4jiDKqn+HevSfIIeKw96dIp
KC8pvUjnRgdbUx3ppj0/WHcvSW73tzs++010c6Hl7Y3jrKj2zse5+8jBt5QWNf7O
dJkjTatilYiK6a6Y21h3Py35P5yRUY+g/zEYD5swtrB/lZk6pGcYAG8D0EPwnRKn
rBbua3dsDDplDiaJFu/5aUiK2sDWJ9ovmmNSebiTHZOKuh1qle0PmVA9MDZXKVft
sPewUJVfdGShtX6iPpsiW5rMaU5PqVJnCUlcA3HtDGhwEANEgRqAoKB+MPx8NDsZ
OYjaZFDIhkSWMGEtLbdVVOe1r/acR4yII5N+XwpbOnN0f6aGc/JmlNixfyMG8/v6
Aa3EMUz4Kk2dBoFP4sJfzQfbx/kfEANyjlig2U9Ol1GcXUNcQS3a0q7cG6HUs40P
tSiH5IwBys9SNJluuPUt5a/0/megy6PtJrFbHPpu5YsuRPvm/IVD2Crmlr+U06s3
1JCkLr40LF19Rjrtc3ofr6F+ZgiWmfldEh8pma4JxUqcrZYppDMcAblspxUtWlNn
yy777OmcI/Fr1qmr3TLh1s9maGvukM9JQvSiVhxqFgrQB+bARpsTzIXGXNxjldBx
uf2jbQCL+4qJM53v11jM9IFS9lNuDpLTGbETOcZkricsv4Fl0bfrTvQ2x99bGqqI
NTmrUO6wSPI8tWPmSy01BxKxF50Xvdcts5cq4XIzQDkLU5DaXKMpPj6XcVpbAylj
um5E1JGDLTTAB73E9wYQf+MIKPbc1sVwQmpk+h+2omtW6Mo4UEY5ynBoKgR+VyXq
xdnYSmsDVkyQTPAWimgDlsCfGvYbopcfldLb778HdYyfKMR+kXLgFAD+prY00w5C
ZjAgmfT3ycH4rT7iAqoLOFw4z6Ir2N6ZOziZIovN42FEjQma2/VIsSc0YFdNkvyo
qB/Zmx4xjMEs8Ru07kvhohghyScF4iop2uHQNdgrx7gP8zrwuCClo1r8Oh1i8dKW
ue+bKwv2BWbZ93CkE2l9sTZwJorZGAbij2qXAmuJkHqAB9p6Zms3nsN5gMMjRxdg
ybzOdxYXti8oYOxncucj5BrQvM47FK1CO1WDDiaUOT3dXb10u0Xvq+BcjnNZUBg6
OZL5PO4VLEbN9Wt3sa8MWHkcBmZ1i2OIl91i4PBV4nTRxYXJN0Cn/5d8GoEw1dVB
x4znZ2Vos4jB9BtivBJ6UEmdgcrzXjeynWAwzheWpe8eBKuK/Q1p7PyoOiS3tlqR
w7siFJZnAOrIguw6m2tJ1yGCKkc+C0A9YIQtY7FLSMV5yo1qvPCPo3Bd/6kftS/e
b8BEfWdyhDoS9wv/sf7ym4YKSUJa9ytP1fFzqt0EeePANFyd9jV7nezGsLhH2Lb8
WzHpL/DByBtyjbwWC7KAYWVBKsu/98uB/XZofIWkho9AMQ0E5nFgwHxXlaO92Hae
u0Uf8gTF8GdNwZSfzRYfsS0rnGrdRHrwaW009s3P1Pqe51LhhqChzCiXm9jO2dz4
lWOebjZtxqxWX7aSflWS0ARbiy1bs7CsnwNAi3L/XCbUsWFmXOh297emikMjn1s+
e4/1PZCz0ET/2bENARE9iEJdaMZLelX4Tq05ngfqv5tNn32jLo1GiDcrcT0L8ZE0
2e31emld+lXm7UuFMq2rQ2pwKxaSaIlInOoPHdBm7dgdRSQD3wxhxuWwONZUI/zk
dNj+kYVGlcXm9VP/O9LWHznBaMXA6wgjkc1AVA77iJ3r3KXSkPnLTDPqbWn0CYVu
8wXSunPIQe4ViXKX+7ptk0qHp+6U0oS4g+8ZwKMWkKT0ZiB/vFKY/YCT1KwavsOM
EEDSKrsb7GAhaZ80iBR2fQctP2NJeDXqRN5QwhUuusWc/5wxQy3g52HZafSjxVdL
nAAzYRIwOA38VlArKogXCNKjmJWetOWRWrEhtgHS+DO2P0us6Y6R9CXFNFfWatT5
2U/J5ddlWUa4QH18WFs2jizv/vkLUGzog/JQ+3NQC5noBp+dILjN8+SCEe65NP3h
mJOqsBi+lDUJQPp31ll4VjuDimKt6COURHUAtZ0S9UGBrmcYQezNMsmOEsRKNwj7
l+cfHiJfCAXgkpoX9PHO6nIHhHnHuAwkMnVPhdTz9Kew3NPWISNgJl8HIxQIocxb
i2pivlNfhADUo/4VHgRATlRgW3PzVKl0DOvL1Powdb8QEM4pGOq7nnSMlzvHqxuB
ht/W30/QEB72mhAma5U5OztVmzW4OQoLqweKrxLJSi3vzXINU6lxV9ZWN6UNubhn
HvyhOUcqCVW2ZPQ4mnLTxpW8i2Jm9W+Tz0gpk9negIT5VEqSaDofF3zux5kIfHrS
J8Aub5jjDVQfhnQfk4FRgeZ/rja14jjtpVzZeUT4l5sv+5DVZjLI3G/YftgqkKJa
w3v80RPHa8wl5++aDYRxhNT3FdDzNs3eG7+ZcbAzY2mgasyLewlZt7S9oCAL1oG9
cUWgzeZElPU4nH2NrEEhvfjSL5l2XLdyfnbpa7Did438tIcHL8MN8FTT9cFLGejP
yYdYhNUyT31dL9NPy3cGeBMkcVjJlalDOLeIhyqfbwQS8IXgcePPURrneZcw4mNq
OvMQn+zzCc2wGYmkMCJdyujwISglKLjPpW4rLIMknfTe15Xs4Vv80Gp/0VqNCKY4
mcsKcY9ix5O96tlnDOs3UzeXbnfQ6UXsyVyDhjyGPnuT4vT9KBgtQ88ZzNmLN6dQ
idYW96dItDENXtlqjU5bK6sllPnO38coJGVczwxuYiM4Wi3F51smLWXMuC4nzb5d
9F2oNx8x4lvRdtp6/xm8oqJCOV4gUQd4td/ZJ5SCCmCWtCXPWcKVuLiAZDC+Zn8V
PLCNB15LsgCMi0wOwwaAMJmzEwQhu5T2Br5oI4vuxLeTkMt7RDglrYVyYUA2VuZB
XUkBUNQp3ISYknATvvnWqO/dezpnTSPHbdODwHKrmdfjw390yWaptdrlv0+Tc/54
gZknWoPZy898m6XnaY/r5VO5Br3fsPxt1bLbpMQrwXGIFC6kUMEIWbnJa21eZT5q
/lLZR6q3Mpc0bxDofGml4NSHuRTsJVmi/H8jDIu2E4J6LjmaBbkv97c/XebcjIQN
pQG7/rDwsfOTuCiIBANsQwyWOK3ssC542Pe1SrDOwxKaoWGhYuN+cFm+NVXnbhY2
30YDdatps6Ixu27I6t9D9C00dQRdvl6odIrhoj5cQYM7N82SNYmofIsHP1t429x9
68S62gn/O+fuSFBlaVbz7T6EOt9ZP3wnC0hWc7xgq5ftJdk1jGzNDoV7myGOHZYB
M63wi4ityjUGPcI8kTDI9tPUHwvlTVX38wRZNLxEXC4kmOggnm4C0cCHBiY712l+
cI6CVAnkTvwF13pvGZEV+B8Bu4OK/DJuwad6r8obXkr//4HrSPxPKmtWpcueAXNe
57k8+++ST1gVxSEHLNndza+4MLw1V7Ka8r2pmurB54HSb9v1Cbk8teBM47dj0Q1B
WklaJAxm2QysbCH2V2ldJp/gRvQJ9/lfcNXZFcISJItQJxZT9RNPFyjZLfIMD/fr
xcv5dMg9r7Wn3Ac7HhESoKZV/YofK6Eo7C7prQmD3AZeI1sKTIPBUDO9B6O2ZJkQ
sDDd3sdhtSMjmJg9fEUHcA34no3XYenct9Z79H00nLE3iay/DljV2CubJO/aqsS9
4fZcJthFdMuQGA0aGcuREj7R9gf1zrJrE3lfjOo6lFurWdzc954tBiOgWwOeN8to
EHw4VnJ23DAbPaKQI5Y9LP7CbHYABWtmOGT9Gn5eUTz4OTkw3ZGLi9JPguWF/WzH
OVl1zRYa93/pPtHPV45ZkCKuTc0xvArQFGuB1p0SX76Doy6p1q2oMRRsx4irtxeV
LcbGcK9chrf7PtEgzbCoOGP2P+QP7zUJ9B0q2uqKOcyEtcduYrQvmRZP2ttv3M9G
EncRncP48E6jYOE3nibt506NAo2ZvdKQTwMcp7Vr6J2i0bJ2IFQCyw5nSDBCAxDy
FyP7OWKYNVaDR/NLy+NFCzRqLYGviHFItC7MhL4PocqNQwzeckJEzo5G7EbE5qzb
3sX7zgsFU4vnRiGrKPcTtXAWJzt4kbk8nIKl1ZpBA53K4TN3skWUXxuPc8Ub/RoR
dJbI/0vI7nXiJKr1F0FAiG7sbUgjuFrIOnHte49ychC4JQsZe++5so5UmSkVBawG
StLcvtPyGrak2vtjm3onPCj6Z+RIwoWiWCC/yD20Ye7pZgw0V/2hw0EA7VqLhFO5
5jqsFVgPV9QPxlWu2xAUII/KsV+Eesx7wPU2HeQCU5nHmgVu0T4xAsUbfaV7S6wx
qW8bQI57I26HEyUGXQ+yO1WHpGhEefU9T6Xm+nUi+CFOE9+zqb4iSBSHK3Bxcshl
PhinG37S71GJB2rCndmgN5D1or55CSg3xgNTcLDcGWMXxNSVHDLiJGF6iyWcnaE6
O9Z4RCDYWVNt2nfEaME7AERYzVvGwS7Boqqi2EjclpSAq4uOAcJYXxvPyAIh8MR3
WOZt8A/n2MCHsSLGBer32CEydxjhXHNpJjL2bre55/WCvgGqrC1lpXQtGecBGfQj
WAqALJt3MJ4JBPpnT38Ewq+tURZf2JsCCFs4fRHaZwUxFzwHmSkFcF+4gCQAkfTF
JoIjUfmBvnY6pEw84MkClzCHn587auU9Bg2jK9YER438heiK51DugA+ZA0go3RpC
XcWjtpdG4JwcmrrwUpecUGzN5GvzxG7xtTfCoC5uC4ex43ULADdHlDM0+TALTLWV
oMH17PyKG5q02Ty7H6zyjU931kQxs+pwYQERkbfz07GiTKkn5qI/kHDXJL9oR7pR
y0+9ih2bDEyIsmHUY+mxKRY+7NdPYr6LjbSWtC6S9Sjuvc8641PsGb6QimdHDMfQ
6yRQQRPpCT9rBk/hirQa001aILIhI1lsD2QRh7zpx64R0UTwep+Hx1Te1ztG81fX
UIKVdnKbdPMycVSl0ovnWe3jEU2r48rZRtEpIeQIMfNEDC9O2jby/6QVSA8TQLUF
qUirNprB33PvmdLxmvUsm6ZexQ3WYmhZ8uWjGDLCYotyByaSumJrQoF6sjIoxQv6
fXCkbzRZMaQH8IKOWVHN4j27N6YmCp2LZFWhzDvSJ4FwPToCFNpsZdGP3gUcD8AE
OYhFTyZbTSxAVf+//SB1eFGmRxuKHjIwLmj2hiuKfgNjuPLO8q8D1xLwqKTnAo5m
W9AdC1roPg7Mf+076LRfzNMUVf51kOrQ4gPA83//jNcZfYzV1Mr3NYeIRX/orr9P
ufVw5Nkb+lQtrORkm5O1BIkbpYNak4CcDk7dxRQ7+0+P/YqePHeO0j6Yl9FEzMSn
i2nmwj6vv1FyhGLylEcej373rJEkH06b5KDKm2tJgvcqzxqE4lj0hfiKbQKgz7AF
ksw2e2/aPkIqrrW1gOxH62CqhptVi3N+LI0sDxzzePgUJR8LMyRCh6VVwaF2ybiM
2o8u9hxJcYVNE4wD+yyDG+1XrywfS8l3rqilKbNZqzch+uBDnE/Zq7Qpyxa7uj5F
1DqEymRs7FoNozxsfWG4TA53v4S+qyPkTvOVxfQ9gkOeq7cv+aie7gCvat66kpC8
0KyK98xmmsgUnOEmaLwJm5knra8ftImCYO++sbfSq9ZLuO5qOldb/f9uboQuEi47
dEukM9ljsEgXHwf/ELE5uIQoJNXZn6t22bFnp9dh8OKoQyv8TC6UkItORiH65R2e
nZGkqWC8wginkTS9vxSvkHdwSW/1J0D+Voexal0ZzJkOQkEfPoHxQkue8Q7hyQwG
SnnH+sjcJF218XYX1s+Zry7B6jU7YeaJgQ1rXCnkR9Chb9f7GrlKXhICc+JSs86d
sBqrDG2IYRO8Zqu0pOD3b4lXoXP2zBT22GvoEa1l1KOPJ5jvgXJ+TRthEaQiI+TS
jMaciJy79ZiNON29cU8Xbg==
`protect END_PROTECTED
