`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UUZedkbzYG06d92RFJyGpKOOyf6bm3EYBfEuyEQPaWrbXro4a/QkusNwAU1nzSXe
hwZA4xTDm0yWPkwFFp+FGEtDqVKMIlDFKENfHlCiTJcjgYH27/3ZlCHLHke+WPd9
opGJ5cDwIvnDDkJEQU9n7abrA+uuEhC1jM5M2Q+KuRnlnN3/Xkwpxrl1HMF9yCuo
8rlUI0cuEke64lFnV1uWdqKYzEeLsv0+6jtholCGESH8h47yH6FQ6W8JXxJ5gZS9
Nr6u0Z5RYOigsm1t8qdROPzl2cv8raUuLfLfY8QeFBZLmX9nmlAE2FaWKQSk0Prj
NmVwklgSikkKhg+DydT5LnsUp8pgJ8YdNTr3t/8KITtpMHMonDMPvJ5KnOMwYJCa
h1i+Nf9uioaVa6UrW8Ly+R4AEoea+8VdUuOrCVePQlV6AT2qfIJlNT8HnmfYu7K1
7rhBIFTuJ0IAxdoR94Gysa3cblmnupY3rzCBVWntVRSQlAOc5r4d0q/WB5B96VNh
C73UNVlAzqF2epXx4HV2in1wG2Q4G//P5oU0fr3URsd2ch6ZlOpTzDiyb/8QPrDk
UgRjUSPCnKKFvoZfbwo7RXrh69YVNcPDuEnhlFh+d2+WHOY4NRHXEeAQK6/czf4M
G/+b8Mk9o4B5G5hU0mvnL2T5FyKZcfv+YjifggfU+nsTlGI1L5KwNJMLeVOanszQ
BCO9Lko3/i+E8eTqWzkri3l8fOZqEHWo38PnWs/yZjb2CJUGeXmoMQ3nGmu1jBZc
1K1Aj60ixSOrrmEJqrl4PhHMNoUhRKQn/qN04zSjZmgEpwr5glqLwh9WKXG99896
g90o8l8wgWgbfKtxf++Ec9QXblIx7REp476/N6p1edei+yuJJia7YiH7i0nmvfoT
gI2SzVqOXAsutmZhdRh+IR6zfCPYO8xlsuEGAIHxDx90+qesGHB62FBF08x4CqbO
r1L1RLOtDfVIz6sawebb6NOxE/T08pxX6W1n3YIwr7S580sUzsNtKiKUJ1Jx4kTD
l/H48J+ovqikJnidLpu7HX6wy7Wi/P5EV6Otzz462DONd3phLd9gc8RFYRHX5lgY
A/CmEIGnTrMii10mEkaMt7BDoVXLXNUhn2GHiye5BKeL/i2HJ0DPhd9Oyo9672n9
kH1vyWLmN/wAor3JhRU96waWR2hXCL0rHhGIy6ZRguQ3S1uOuDFDzmyZBMFGHiIU
wZFTDqpBGqWfup/8sZm+mmgU6q9lRZOBywTUWENzQrCmtqTeFDKnK7yApmMTrq3w
qqBJouDCzT+YCU40hxql0YEMINHcX3gcH/lG/gdb6iS1FZESQ6f3s+PBwWwaurdC
jvHfDsJDj9D4OJEpUuLBm17gOMVpPYklU5vGqdjgN8wxdTZGChZGRi7U1AIrXTa/
++4nCroyd2VRklyy5rVbmqsq53VBZRvog0V7Xv6IFgjHC/8Gy6Xlma6CQYQy3B83
6kYqIAPbYFdMpyCv5k8inXkESvu7CMTsw/xm9tRrJ/pMJoguB1lCzbWqPFmowpgm
1SUUiYaU9y33sgKVYh9vD+2A7IJfo9zu5pKkbOWKwPqcpQ09D7rRb85F/e7pbhvv
XB28onuNLVM5eAbfv/V1coika8bxSu+KtZFhWoAV42hXOYH4K7o1ey8I+ait0mVS
wQOdVBou5W3qZvvB97Bso0oyI778YGI+kxp9nerc2+FsVN8M6EdH/5ryNuNme9Gs
tWpzb/uGE8yhaDcdQ8ONxhIoqqT3O9bwq0ZX/NnMJqWXrhjxpAinuHJZy7E/4ltc
clMG30IhK5t4FNo9kNGN+gK4gIIGj0dbMH+u10vnmkmX6OucJb7AcnHH+yJu8oy/
OZcqIDw5ahwOUqBgW6YGQLfPqdQgSapasNkjIr0I2YAgCA9jDdpp1FaXeSstroP2
GMgWY8KRrGyyJM7AHYx/zIWyDcbXJcHwbEMq2EPriFUhR8YzPq+PU42XvBzzthiQ
g1TiCJVUbzAHKutYnbN9UGePpg0quBMOaw1WEpkSfgFCOpBmUs8bT5v9+ZBYF60k
digEpXjeMmBLKRQGesMdTmM0GrETcoYWvwlHUo5ER4KtdMu1kVNDVOwJM6qrXDxZ
+TrKzmfoewX7UaKvosKKjLJf5msZwMJLkGxrNtewjBZ/uSMpmLY0K6+TrFkNRLit
UIbrcG50Pd+1f0k4rbeAWrffMjyEmV+8Vfik22uSCNMo6WO9NUCzRtu/oqqahASK
wP5nzckUCSWWC3Tq2uxkFdr31/knz+WiFSoV6c4wN2H+8oheGnoiTLE59CuFbU3R
HhYY7cTacliwkWq9tW8PNZ4M8hmGf24cCd7pHDQhlxBz1JDMSn7ElHHUjcfXiZ5h
a1fZic7aCSHOe5Dkem+IFWFv6b+oteTANoU9COEv2hbukFN4RoVVL9v/RRlP1HUk
k1nPK42Xh9PXvdWfNWv8oaK9nQtas9QQQvnkGrgorMZEvy2jC894wH6Qzh6IAe7m
+wjR4qTP3utVqXJDQQumCzl0Py9vPPHtd3HBvA+/jZPgptwFOBW6aReFy3yeDUf0
PKsiZ87j+4ic4NgCYc2vi6tQgmDslmMutwSi9uAkuFXYAF23asaB+z/hRLC/BfMA
dgT+qQ1OhCHJ9jsAdTBng14X9gCBqBmraHdNt4Ckvie2Lbc8KKn4pU0/Rkbq7fnv
YQQ9MKWRT52aFHpfdpugAD9EqC9MPzpcngosNOx/malJKceF2i4g5RV8FkqctoA5
cLasglHj97YPrZMxP2mcck5dY8VolPn4+efWmytgFPQuAX7CRjE9HYWJ5OKsVkOC
G1HjHB87r/MQEsmoH3AC2KPZbrhgt0l8fBA9mkKujcHVGV/ZP85WTi/d4efaBfob
b3wL4nJ4bMDo3HwFXo+RLX7eQdSmqf6aNTQFshdNEear0ND551Tt3LaCS/R0b+Ar
h7wNIswRAJAOC93ac5mVRB7RXVWthvmgvyXqoBo7Em5s1UfS5Ec12lCNEwj3b8PB
f6KeTY9acJSLfTsaC9t8jcogTQoWN5a4U2gc0QBt4pWVH1FmWQOBWMRtIkfkB1u6
SU7prASY1Mw55yw4Z6JJI1aawDBT23geyhoGhafAyQyE885+J9BquoLgwNE0vbKh
JPnXpTzzY9asfs0Sm0911Ytn4Npts4I4K3EV/BsXBmrtxI9AIlOmu443z6YfKBBh
6p20xoY9fSlwnNX09e9AQw/4Is0HNluMjieeadanmI5cNOSqrcyQI3upWZccloPy
zYrbkWNObUvPoqM2CNg+1Uu+82i03kOADJjKAmOsfpLaKkuMRt0TtzXNBOAwBtdh
U50hm7jxxgUeRZCsaJxOXWz8xznygHtLiRt05V+GDwzu5pofVJzhAV2ddbofq1ac
jS7jgg/RqMVeqSXDX7UTvbx3yh6NxSkVhEtv2bOlH8k7YzrJ43Pot3YQYuukLeH3
TmeFrU2AeflowaM/CvHK/v5nvBEaTOIbovez6dh5lSY3yEk6gUVfTnd+biIHieEU
hREzE8lrVOEY021V6DfZgtiz4J7hR9Zk6RcOYxVJtYVybOt0AkfM2KKMIovymxCU
PEE22qngfCglhJrt/d4VAiM16BPv4CZJN0oNsvxPrveLn95flQ9b7dJzqiUeQG7G
ckEtTGDbYadqFdQijjXp8LrSabic6patZFpn7PAjp2838kHyyVMv6AnyeSMk3l23
/bTQ1I4B1YBgc44TiN3OPDcTlMdsvftj8G7mTcMsrjj7Xv28xPKrlfyXSgYD5GXP
GnPms/hCHuu0VfNHFSWplr1YCtoXETXEs9qpJX11RH+PPBnUtc/PAZ22XDFaBKNN
iHsqJ2Hf3l6ENt7ZKNm5iPmffA3SsNQ2jFo1jLi8MH2037SleII0NyWcrC3681qO
jfU7hhU3qIn1l9Sd1FVnzH/1lsoXt7jdhTkTT7AsU9/kf1fJOugpqt8b/qOA0r+w
VmPLcNlKYrLOvD0iZDfO6ca09CGltMLkCadvHSZOn9A=
`protect END_PROTECTED
