`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lQFB/LP+RzXk4pIVDRI8rjYPxEj6/S76lc+V3PoT4hmJntuF/5oJ+hNEPnzTI4JK
Izm5a8pn8BSWAW0Y/5gbbk2/5SIbe3bRC22mpmDvOH1zA43jLKIs2QrvkSLSzJtM
6xbwb2+F8mkOmfmP9c/P/EhGjNZUBI3RY2peh6/7bDoMzPALo/aP3C3n4P624+dc
RiooDVtj1doXajxtfwSjVZBZGLGcQGh+TSUe9pCwn1hyWDTTVuklPLKLCqirwRgD
iCiFv4NpReysXvsrwCnNCccotUPjBu2pwMfMvlpmfKJnLXjG/TZ2e25LpY5Fv0Gv
2svEKwz3Oyt9S52glVdWsWN+sumc8egCvpWwV2Yaj6KAn+JO+5fFnJgWOE2P5uXU
801F884qbZnoWCONjTbqfhLHdnPPst54zDpCQUnZWKd/ZbPokR13U/xMeWIgLPEP
GKC5rdtzIXP1+o5iHU72aiGJL+AMOozR4nwmlj0usqhL8wm8t7EjSi8MWc6Qoy6D
jBCkaWr5IygG2zyfeHpBTERTDZIFG+rGY9bKVZKhxg0FWqc26st0hfwdZSirphfb
/JCPpcf14gev6lmEOTbdaCNYh+2S3q2Si3EtegKoIMHX/pNQJD37esvbR98eqMWw
rpwVOm0mCmd658BOt+azkmPbBmrXdb+bPrn5jmvKs2YPWMqvjcbmOenQi/oxuJDP
H+Oms9n9zGgPHPkM7ZWyfftLnSkl8QBdYxxBkPlBvoAJvfyrnrvpO4tK784iTf4D
gg8pfXFw88QKwgvWoq7w+yxsE+OvpgBiRDDNGB6SzCGIG9FvvFbPTWCOoS+anULi
IgYSPrHHxvOZyg7fEcCGMvG1CfEwxs8YCvKTN7I9uzvukJP97ytTmSIhnMsIaF2v
XzsIDT+ifouBiQKM3LpLm1XAQ5ZGA1d1QnXH0m3mWJIYxWNlG7YAGaOpS8zWORfi
Zlv16zkh9ivCCJs2X2TQgH/GneD486TdRUsLn+Xr7V8h3Xyt5S1x4GL7lC68NjU/
vQOBPM3cHRL2P60RSis5RMDLCP00WUJWNBhgAUL9TbBgT7Y5ZZhN8hZCYEzfnfvz
FMlfWPiLn2WijegCJdVMKhkYdj0jp9H/l5W5OXPdRhGzWCfXVocy/PY4B7m4ye83
R2eOQDzfGWvodYOsKkyWH75NxZAo0YU524GZqFuHrlAwAhdQJ5/upVslaxacADN2
2LaofCAVvFvaIzxl4my93oruZx/8e0bUEk0hUj2jv0xnBDshv0WJMjRtPnXmCPCJ
d/Wm8TnNEhOeuzdeE6eK7wsTJux9zaPuG+qv/Uw74aOoNOuC34XlbEIfJ1DxtGmB
SuwaZ4A1ZYuPg/oRLsv6mRQpgaLpKsk2W2q3C9ZEvtTAbpRgTebcGszau9gvEfVu
JjYImPlhLTLW9KdnkXMoj25jTeT64/43/Zz9MdcRFO2mg8ZzF6HOrhUhLUWmpe/w
mdGidJ/ZQbXv3FEEd1RWB3WOhHGnKFdmsaSQzCqFSloYINSN1raNsFSE6PNb4Zc0
00OfjvEVQrgjbzcxUSJP34JZR7XYrTNbgxWwdDCcmx1QDYQR23ssSZA/ZrX3R90t
rh7YCu8P1MF8kQgLXr49Cpve34HNe8g43PckekCcFIQXSCiRiFuBf52WiLvqAhGu
VNjqBWtuQCX6Khmfz5Z2+xLvXHioMvckJbN9sBoirSTmIubNF1LXNFvauBnQqkWD
nuj0sw1rDL189+nG3GwgdAycXwE2jtXWJjfEKWDNhXH7ODh4MeZdex9yWL+XG0v+
l84yr2V3qcn4Pfrxg+gZrIAyBHDb6P2CYaxrQb0uPU2ewpyI8BVSuXNVFxjv3KW4
a4MORMkinuLgdPA8IzxFTQj1nFv7uqjNI7KlmeTHWyALoDN7npab2oYDXNDxkRU0
6oyD9igrP2xgiKXjIXmFuC2VI5dazFX8uvZmiQWO0VaG3mMJWmGFFa0XrjkmW2Ba
AVAe4sxT3UweBvUBZvSfYNn1Ruwpe5xOwXu8dq5zxOeSFJ0YeyCC7jrFZR/pKRMq
vq64wVDhPK038F8TRLNVqDmqA17uue4f0K6kN4matKKMDSS9vSzSzrZVgERVUXzb
r1cC2A9P9oOVXXhlyWfq9NFhVkvjz49vgC8/vTY3mnuysQ3M4a0r1gMhLtfeYNCB
7lscI86RMtwqQtesxZiA+z0pIzKh7cXmbGv6hzeBE5itLJEEc3HJbHgpnzospmaP
KF1wESSEQZK7agFbL4361BP44kmADdnr3imZJguX2DPr/3tzaobwDMjl412s6ERo
AY7qhGNXcStEhaR2d5KychiDIzigdWxwA5B1/Dq/milJWTPga3SpUVhtWyvMbBYf
wKgg60e/PPY515sxzIarc4O7KMcSxzFC1KJhx+N9OTyYOyg0gVNV2wPwnx0WGjfw
kaKZSc6GIWFjFxcV5nhYgLu3DEI6R+44BJGwRQRNUeoGUll4bSk1XR2hb4jmR2kn
bxbYRwq313fzVFfXlfCqDA==
`protect END_PROTECTED
