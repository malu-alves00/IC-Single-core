`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
w0sURSlSz5O+NguwUxCJs15rk75qY/gM9udIrKiw6gUVVX/f5rq/KoeK1wjYVeHe
ohV1N2zPa9Cv6wesOG8JWoJdctRz9dMC03ewSU9+h7Ne7sx9m3LuUPZcsuJvwZgH
c95JnsrzFkrb0F3CxwbckrfrwirhHn+FiIJM4riQZD3hreQyKN6tMy83yGpLf1uL
nix+E8nULQMBmSW8o3v/bTtR3jRusx6AgUZfiI1CYFQg/9ZbWrbLOYABIPyDObmL
0vzR7dCQKBj3bokgO/7dnkRJzB4vIUSVwBExwEyGsQinLlJ0HvpHJVC41ueP496Y
/vTlE4+HImWgWgW3qLIUhHCwbQzfyYmhQYrR3pamhqDYi1b2NAROyrYny/lQZEt3
/AWmnuymUxyc4ojQql2YYp0Fho5F7b1oe76uNti4Uiyj/R9OO5/lQIhzc0xkVAkz
dzOsZ7sEWhD0qo2nYxlOhBpWZhoVNOTNCoToutua+1t89w99Yf03c6uxdaUCBAWD
QynUtA6NucVw6CBqK9WHoXJ1sGU4cHjw8eL5HeCawY7hhKDT6NyG+HvOuYlmqG9s
c600OLJEEwotSI+QIAkNUnbTzNfBFUdyYogONJRK0koPQ+eHMy9KyqruMrbZOHg1
EjRDpbroje3ZigZG1ohGfE8Nx4bE6BwRiGs8qL5fwJloEle83ySAad0PtkZ8cnEO
RMcqrGc5af7oXzalsMD0UU0/Ug6mMVRIDc5QqtOiSUkPHnHdW53H/EAftT/c1nxZ
NWGYcFBY2F2pqlMpKVNP4uEU4+LGhg/Yg1a+jzjIV6I=
`protect END_PROTECTED
