`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
anNwWhp4vmO9q8Ef1lE47PbXfQsTe6OYb/UVtX7983yCjTJUfXa0wANbdYBkoteB
nY1+o3cWHKfpkOUtAPkgmXPlhWibgekfc3HJI5wlUPdHWm3itm8BEoQxNMJ0k3xf
uBeGMgzDP+Qb8kAZBjl9Thd37aCnLIwYTdX8mAunm7SezfcHM51IeczQfW8Bww+C
dOxMPewvyrj1Vbp2RwwIxYE/EVpxCDoolcuqoAWmX38kfHVQbx4lJlFHdmaVrxd+
Nsxpls/fUDTu3Id06h/vbvmyZ8P8j6cIKcft8CHU0XDtsi+ZSQgmIdYPZsl9wreC
yIOa7HsPeCVZ1hGoiQk+vULz0dEpllbYKFBmxF5Wdc79U/0JVCg6XWkXZ3LYx4XB
8usTG5jNGEehJ2UPKV9EJYSq7wzK3FFhTHtGIg6aHicg7YEw9YjGtu3hi/+iaWAz
39jh+rSao3B6mQLbQgvoriabOilf/I3NRU11W9MdJ20X9JtqhvzDuSwQJpvJ0FQu
Asr04wKLkBdBuJA/Bb/IaSdLnbdn6Q1zyJp0q1REPWXzqJFTDvZ/OWTPnBuCrfKw
YmKAudFbJ2HsBqrJUIxaDVbkFAINTntNcabzgDGHaSP0m9KYWXnDFpDnhP0NQLw6
u50WIRFN1nELvdx7q5hRyVKhgJzlJBIPZVkoGb2eUJRlY7vOYeXaabRaVBDeEliH
7T3n58eJlYQA2pH2VCG/QaYElAaVZ2DxpiNkUZ+OScsNeCVgizsz0+xp/9rg7dOS
ixLsG99ImxBSoQe7v49h+kmhFLvivHMDN48Q/QLLXcfbnM/z6cWo7C8FDE8ByPlh
yXBzOj3CujzKlMWiIfpZEKoEsfsR8wrZBxhynsXWfnmKewZo9hR6ZRYRzsMBcS8N
bpaTADZkVztitwuyCc8DG/eoxEBgxnIuUNjR1U/TQ2UDUbDPlsfzGlAt+jkGRsrC
qhqi7i7jN68c4ehBYpkY/qiCr3GxkEnC/dPDgst/SksBebSCG/jo+5dD6982CtSm
FgSO5lvEN0A0SYPIzUOMeH/pKE23TtAhh2diotWATSE9uWyK7ZZPWnYbWwLnbPPI
CswpcwX258L4w2rotaXHpu9Ae8o18au0ES7fgCzkmXn0gAVyhiAPwdPmi7W2hhhY
Ucjlmi2rN+67Ru0eQiZvcq6bN4xwBf6Mty+r3JinkEJ5jFEHNKepw33pMiyT/Qqd
lr+CjiWvzNXIi8mkDdviQaNcU0JiBdzfZXoZlH1EjHdfdy72IKM2X4KeGy3EGQ0i
tpk0Amz+9CGCffrlk1H6joc+2szlY+zlzL7lg5xccommbudtpYMoj4N5lmTP1Q5S
WLsB6VaZFgOxOd0iTZo8iLLk0r0E3FlMYee6t3HrXU36lsFjKnqWhSZ0HOoOBMsp
spW1mwAh0REiMzCJJ+gph6D/fnQRlh+FU/i2ICjb+lLdajTMD08HXO9OeSP2VJSV
hAD4mnZtv+zRXAMR+p1mIeUqgTPiahk/rE0ymlA5fzoNxmFF0aGeKjaxyj1/11eK
O4WNzL9Z/RS533o7TKypv0onfLp58KmLVuD6CJcVRzrCbyNcYjwrGiYH9C483SHc
4RfIv5N71Lp5O9ane4S48HN5bhJVY/UaBZDGsX4OP79favZaTAkoml8Eo733vXPf
bigCrLhv7neLiIhA9mLC5ZvrspEAD3ef4mlXb00bcPJ3FSzr4tvJdXX27zvWH3Nc
7IWtwTWthEHTk0RYBSCXsKVf6mTCObWUhAmA12tAYv2689X57CiJJiqFIxxcNQVs
w0e5RxAx9hd3t6rI3Kd8aCrLlwSTE9nyPQjx7X0sZsPIju94S3ValhvvWPpNw5XV
QlmOmKyV7U63YWPQ1NvQRBqqRDYK3UDlLQgbRvpaO0s82Zjlz7WcSPnkdG+wzPwM
w8BtT3XPk03E2XnmkBYJd7z/YUWqXuO+6W7lGTb/LtKZFu163DV6GutQA/si1TA2
73MhMbCT8sSQzMH96rw0y0QITaUoqyBIdP7fIQVjf8kQB1oNa6hm9+atGBKq1N2B
b0LKVOGGXxiJCCvi0GWJHX7P1v+n2zy6/BSoRy0NMJNLKTtjf+rX2CocGJo5doVc
uVddJu4qmU+DBmyuqnbvk45auICZpC/btE7FS955HOXIojzKaK3aBwVflFCNbCRm
MjOLC1CqQtzCRu1WBdyHiHUdd2NAJE4R8MtvLLiZaJEkg+MTW491Vx1XG19rmVWN
VtanoyvVdXFhBk7n9ksazLIk93NJD6fcbqyfOzbS9yQjc9Xl4olkzjD854/WwkVM
4G81s5fJ9oaTYpVOkfPcaGGQ+U0asWWId4oG5jjzxgrKB95XZQpKnRABB7WFIQMb
t/S6qxPKWPrzNtC8AyXxHP+ntHDs3jPHVVIDOHPcqFBNFsyFnNzxINnI9L6G2QoA
0XhvVpgoushF2ls7J8IxAf1MPpoSRne0G0iDXyxVOAx3PNjQED9bJV5hhPeIn/nc
eDP3wkklYOJnJ9OMTGrGBqsKFibP/LqVPr0JbRgnRgYhX6QfQhPGROWjB2FajD8+
eCzqUoknCVtj4FEqmo6xrAcojA987thXiFJZT53zA4xdYB4bKrAki4oEcV7LWco6
RnRjjCOYv2SavITwktRVNnq/4lDQ3RsgRQVicrLejLVOO8o6YLUxq7SmfXtKiBA3
j2SAgSEcZ9CShA4Pq7NWNDnkT8ATryphfJdM9TTpQ7Fq6Jrjc3Tec/y+p5QOZrI/
n9uznNQI2Pc9hg8dBeWKuqDLiGUbQCtgoFwcnLnjIb9FEEFKjDdQplLd6ZgLZ64R
PRj14o6rz7fh6bDC/Qon/7aPgK78vWGhMCjaojd+xBYf8cT3iHVdxG5UodgTAHYV
1ayZe/Q5zejmleWXaWsIh4IE0cZQJmxOW2eH+Mz79WJiLM2fJyIACGrC5kpOGlB8
z4TXC/GBN6oavp6+tRJD6cO7b0kPUSEGtInvOnkABfJf3A1rr9i3iS+8cWsAivox
ronjQB6+l7+OOx9m3v/u+8pKHCf4o6PnSRMgxeqXaQBAE7sV0UT49Z3br4YytqWU
g2eyFOtdRGAvzGoRMdHicrKJRJSFICxGdjI00MimAcAqfYv4cgfxzzm2t5WlrGRa
wotj/Exed8hH+qDAP22pCTVrzwGKQCWxpsq0eapUFBlDNCAO+LhBSx+XCSyNEA5m
hClkSXUWLTuduxAg2r1smFR0hJ2/WIRlakkC3nZlIKAdfZgWMAJcbqSZ6fYgsSqC
KAk2rkGI2r1jfFnZMVEK9mSvZjU3QPbQ2yBJ/DXG6CFLKFZsi5kaJWD5ewpGBjn2
eUQs8eJnKvKScST1OW70LUzlJGVmdW/8njeIeLb0B9b//NrUjtzqkzJUkG0jGKXU
wnP2ST6/8R7kABwcIJ6t29JH+MWwZyUe5wRizPn3poKN5gy5H0IGmAZMhH4SUreV
zGR+NDplcbz0eNA4qTTELaU1ljkn2SUHIR9l3R1D1RkX9nA4MkXBVb5aEZTBzMGR
bx0AcnVs3wa4nQCKKCbxzJ1Yw/39rNez6ojql7u+PgFheHQRhvrirwDaO31AlSZ5
2jUa0cxV6AMtNDGv32eJi/FW1vAAhpA4kCvZl0zSvG84Aceup2pSyMaA3V6VZzU4
W4MkYXjiXccCREokRQzKZtbp4GXe6PrfBimZnQvmLjWLcbTj9TjX0pYRQqcm5vX6
4p1hzFa599aJ0rpEVYUSiXkxqHt7PtdAAtXW69fF5u3euAjTTjdb+pur2NSQuCGv
DF0icFCVopzdPb4p+mcAL/Tc0UTLO4etXg8368J5txDjus3gOC7/gB4o/8mVcUdg
nMyDZf5CrftavvSe72Ckjda5qIqznAbi/jcDi5fxU694ZeWpKo+tKU91b+hvaPLD
CEfEJ38uIwBangWPuGQAAR70RgIrJzLYAz0NTpwDIQGqflt8FZMqhQ3fC2Si94cB
wkUDlVam95IjBH8wn9a08jH6H+/D3OeOR/+tj1Q0wvsFg4tMaMfWFWKwm/gnvNIt
G4FJmgGeF6cdNh9kHojAF5IfpH8WT5iKJyi9r15UPiZGdtzGHg3ROJubLSQ6zj/N
UtpXkYmz2nNRSqXbpUNOXsoizoJ09Plg2eXMvWjObMTP7i8D/Wnwb/+vzara7zDd
7aIJRbRSCY5IbcbzT8cesT2VXFKw47eXeIt/siMvU1gB4rDCKWIzOfoAsjdhr9K1
bWLAJghtLBQ5yyYIvtFLArAht1xKGwfBIPTBVPw8oGFJEwzmUL8/nJwTXhHKVZIC
aOooXCDm3RbfbUxNiDanjJJfJ4d0+QpWTBGEX4RSUV7FspswW2q+nX/JVOao82Vc
LG9Y6YS9ws5RNkOBAeHXD/AHW4aYiGdqNVdridUoJwcxZ/7rNoI881INclX2+1BY
0Cm6c/xoaGvD+4TyKPRhkEijf6hPk+V/SD+hveXy2WrIMCnsY54i7iLz/Ojs3Fv5
K+18R3o/FhCvTim1zW9Yh2dZH0SCeSqdzXYLlqlHHyu8RHc35QsisMLg/8PX7526
C7GTrtqWvqsRYWoJizvWgpJ0w5RarV29MafB4UsMJfsU3f/1oLXqaIkEC7MWYuoh
QPK7EJyxzQSpwU324suJ4Qv5JIjfcsmgN63MPsco+IKTFHFBCJNR8JwQ/xJVrwB2
AY6FLLRwfaqi1h6ht04tR4RUvkEJg6wlKRHSfJNqGoqilE7ABRTNibqvh5p45e6v
XT8Q1vDN5hoXwcwNmjXWXB/M5ZTRTwS3bo6XeG6ng/nPBwsp38zT80hvkYIemBa7
IE2CYhiFx435lqEH+S7Rc9VvDDA9OnItAkpwpgkHSuAFMd8zqyvQ7WHtJ9ZeY5ll
JPHruoEmEFHZXFynDZbYwMYxY9ci09RRCMBtKtZDvd+EclQDp9Er67jEBnTudIsb
iZGXoMmv71wPCWk0TWr3pZduc1T/SAwuhegYhrvCuD8uz+yuNBE9jpxLS9uHXyOS
LhoEPAish2bFlM7FjWNl+vCx6Pr+QwiCkdi8ezz8G5g4ErjgLO9S9GfqYyjOtA+b
MwoNat0fdaxtSIE+GIFWsXLfzQZXPOiUEVi3VrS+yGOzq5R+hDmf8KOT0/XuaLsN
QPjeoyoua+b5i5BHk68sdQXIpXs/UF2hphXSSyPS3b3/HKwmZLURKbYSrKQlJF33
kOEXGKDT2/0wo9MH1GwNR+gGldVnBTZOORwMnhgez8k0dK2ImSwLBhl2Z4S8HTUL
VhGxrxwnWalc7HBcGas3fgEatq97XfIc1XkTO/I9boS4Z++Ay3Nfm1LyuGHt/Itw
THo212grf1RxyLSxq1Wg1fY7CP3PnB2HWcoyc4224AAhtCYe4Cs+Rc97x1QqDHSx
CO4hFYsvV/FzWYwwSoOoBGQEXdthlJGBJL9/cBRPPrVqU+J2SC7Vyv+UNxdyITwq
exaejIAXS04QntcbC9ESnDoEp2Rjc92wkRPsROHmvl6W5IeZRU2aFH64n9BiKPGP
yhsw+zUzhoMLSg2URLFkrTN2aVEoIzk/GIeAEWxh5Qs4zB+Xf7Ee1fv/1dGnQiVT
5xXYiPknaSEiTf5VtGmflOnCsAO60mSTlUUJULBEPl1Eicno2bmkx2XdRs1NlP/+
CXWg2LxFwKi5RloNOG9h6NR0Xa0DJZMjz7EqAk8UCBEZ/JY71YMvXAGTzO3G7fWr
XZ28xGEG3CXdd9qrm/tH65LaH2BcTGdSU2wBPNngzE/SLt+/q+kfF9hwYAozg2nj
7AHPA9eBzA959ZONEugkKaVwUYRVCuE5AazVGEbdb5IH6+pUI4/cvthiGSQiy8yo
Ezf3XQKmsuWRqG8K419TYa//Fm2UeyUWWbfQ8ywDjFoe5wZWbfZDptziP6dCcjGR
9It9c3r8eilKJcxZemRIRKwEya880gpaU4Nkw5amzWb1SB92z9YEf/ScgZscBDzn
AMFT4zej5R4gJ3ZuaOhyjuTsLaOC2ZUI6pu6xcOAyNKng6kfz0EsWq+ccF1jhyqK
n3sAD6dsZmBo+S6XF3Wnv0ie4ZpLrRTlac2056XrPFt1LfqWf82Sk/33Zv1awaBx
FLhNtLT7ckwZ5RpUx5pHvkRKzxnpUweNjnNnHMAX1YPEatoQ36+cdVGdZile48Of
9x+ThBq487LdHmf2U6vEDspvfyqqzOW9+4Cd3Wfu38DGfxBmCNmkFMPEWbnxDaKm
g8UCYJ7mBbrmBCDPVxhbAsVprmZ7AKtQxXVvpJ2T3tZOZ6P2iwVtJvZO27QV9ahi
kWnJ5Wq+cLCNCWZVLGisOe/TDQPao8oW4CIE6cluZjTD+e3YdMOSsR8tMVpmOVja
cu3sny3KCsfcZyXrfSIi76NHoKQe5VJau1nZvcBznDs/BsrirKunfoonTCp/rjtv
LPZBxrIQTZeVdsD2w7vCjMZoT6hekmkwUVvnqPNWqGTftaMkyM/8SBC4mlTMdA6G
UiVl0bQ9iPslrpnL16OWdwX13Deib2uSO+4TOn5kaDvV6NELAwfb5KlpLDEugoMj
aaa13cjqrr/7v6Ck8J12o3B4DiCFcQ+9nr1OiC/VtvxkDOl0vPIU60SHa1Iyo3/m
cccfO3zL9C/xnv0XcVGnYwJsrB7JLjvFfnlvJiH2E4HK56D9BEdT3Pg/l6KtWc6Q
TyBQoXzrDAWaeE+xBYmfRCVnQ+NhHFzz4QaN0zvACw2+nI4X5SADFj0fi0canpyE
rr4N6Q2ti82WI4vEqfQNN8KsF0uVBEjJ8zOiWneEi5FOIoJTJdq7ccuy56lPWNZL
nDfz28XOQHnaO9o+X2ExzI34DVvRlnNF6RRZIsAu3V7qq5hFMladPtbH3bKw4Ewo
QIibx35AADCTGwTi/Ig98zVzpacg0t97tjzENVsyxNRtSWsTx0k+XZ9TjWeJUHDo
8RJWnBX9taARAu1wKXhqTzsq1TFk+yXN3xTq/0NTuC+zyZvZ7cISa0udoWkHaLMq
7cLvyZmZ1NHU302HjeS9UnXnt0gn/gllSUyrwmhVq/Ybpe03CD87rFn9n0ltFFzq
WKNhj2Bo9htddWn0jzszr4GkvTO1cpUCdW7dM6HSe+Fwu7Uu8WG7gzPx2EuBkdA5
8rKjVg9lVrei3jX2gjxND4ZBABlKIokWWFAUOFE7MgnxS0cJlnKAWvF9KKyIzglI
Xb+zoEJ1b13WSoXsueeMOIBeNWEASS7ohdY4U38j2fyvw4JBzSFNDcKxBPpA0hPp
M+Xj9WFj2S0nj7YX9IDV4DsGBifuxe6bXFVRFCzuN/1bZIYx/hD35ddElpbtLPcX
Els1K349L6xSoXKL+0PNRYyly4DZRHW3YCoVPxpM12WGGmPdmODNcUmh2NUgtTQI
/6UbmXCJub7SAatPwafG9EN4REiVNtq2PnLqLlEatGK4EWmO0rG6ml35wYDOvpZj
SBAokseAXgAZVPEnb4uZRsXjRILeRIaoGX55kimgCIVbyqnKMQOkrGRPfrYksd00
9/bjF7nAhkqU3FtJ+goBr4w49kv1YCAw9J/phtzWg/BFb8CNfE6paePvlx66kfnJ
SmSBn2L+xz/syZtA9cbxhpbGx5AssQtAGAz5NL8ZwvKv9MJdn4ZN/NrTiyXvcYiD
eSPWhTwomc75cfJuoE5uigZJNPGcy3JRGExtMHL4FAJY4xHP9t4KGxYGLaA3SMLU
HMnL5vd8eAxVG17FkewL7WqG6PLRM8QRJwVtFG9F6H1N7O6/2ekjpX64qio8tuzW
hp3XOy0EOenSpiiIKqIfECaPX1cntzE0Yls1x3sEYU/ezwdi9Jxyhgl4JAlSZw41
68nVcXe07cnfZAopMFMAyg6DMY6Nr1kR8R8NyzhLkJCKQiDNQ0lg87q0fbGypXY8
uWAEXd4LI/4/noObe07Ke2SUF/PdeLLprs8Rz+hbrTZjsOGoP9mF4X2XpUH0hFVs
n20z8Lnj9xj2pSOQpiLD7OJKIXEYNcfkfwnhmu11QJy6+6c2/1iLuXiAQZ3ENxek
SILvTGFzatyWOtsj64oEe3Jd+fLVTN6hoc1gHilxmlSGGlIXlCtU5+9yOqPo2pek
jbY37LPNAqMIWOPvOp1W8NdyMfi0/X5NE/9FIRbgmdQAUqbvKQYspYTRmW12d4Yg
7D+wyW7IQvn/Vgj1dqxoz5buvphdbAkDlMdcq/AIIM5zoRqdL95rgamEL4fXsSAD
EftHgCCh8uZsF0ip/VRpuRyn+IVjtACSkTkcYe4BCw1q3xEqMhPlS64o7Q5WQDdQ
47PeRbD3fiQFJGpcsDRRq5gCMMTcu66SQy8ZAEXbAocNfpW4b7nb3U92wbtXgTrA
icpVVl2rOi2V9NrUFACHIqY45C8Tvi8mnuobd00dTMVY2eOb+n1BOc/+llTkWUyq
igZEq/CVnCN0Wc7xgLPL5HjcE+MiQiQd96J0Xh2FO5O2hftlu2bxZP/A//7ByFVp
NtsQyt/Zlp1Tl2e7BAWG5WyztHAN9R//HepPF8MnuLIMeGIWkO5waNSkgxuPlIjS
4RvjH2Uk/F8yX+wre9Fi+01evo6tKKEwL2gbjVDI1NJqfm2Wax5ICVCFuP5Q+EuX
EWBwH1IEzfNSQ6BWaTlsK4KZJTM/hySbK46QWQnx6YPm+yVtth4fp8ORNQQ9utT9
iP6HTFgVcFGAFb/IDYCKGoeqaIe4m+64L08+NHkVW4mme79jh585M0thOn+5yjEl
iicBWr9t8eESA9F5MpAxH5Z6gv6dYBi9N3piLFKK5ac6ddANQQB9va7gfHI/zb3Y
MZzdE0smN7ZWaHFaub5dkuviJM827i93zLFdk28dywWwfGvqhRevVZfuFzpy1tPo
XXEbXR/Qo/YUSQt8puJQsALJr3EllB3jDus5FcB0HqlaTo9DTzCjlxdhUdymk0R4
ocpjgxH4g831H37w1OtN9X+FR2o8vxhs7JcgOCot0VpwJtGEBIww5GY3yTc97Q47
bRqwx81YANeet/w0m24dI4TpKDO4qDBS1AEIxxXWEtvswtEaDGf5TtsSQr8B9dgM
ZPc2NV4jkpTQzsHMXMES8vpSHZP1Vk80pIe10xcLBLrtedAZDKDhKHE9bS/YHQFG
ZjMrFsWbWf6xPJcGl+UKfrau/Lb9H6e2r1T6WJnd2f868BtjmVknvToqRd3a/xxD
h174cBNpYo/RBAqEaiYxN1X5x+72rYabLctoD42NXMYCQegLVq4mf4K9HOGU22Ld
zTEvUP2P+yKlz/pnBEBvgg0J4SaviOGYaZOtwS6zManFg+AR/UZpvozuReaVEl37
mkOTTJ/aoeoQoNexONEjhJOVltMlTdAAJ/SioQ1q/aSEZXETQnhA9AREKDM5MImI
ljbCbTw+ntvVl0rdy1d92MmGe9+TPz7Sm4vvKvWRyVJpRS4/bjCtbBMeZA0FgDo9
UM1tBnxWqsOC35/p8QLVjz1F0fDi6UNqsS/Ij1imU0mTZ1q69GxxCqaPg21DZhD3
3hRLL+lmYYRC8JLldJvKnye9Fx0xxHQ8Lpp3xaAa/KAQ2g8pN4fgR7M1JHH1jgO/
DUOZoOnM8Exs45SYye3HMvjHydEixCpIVCU9pSn4xKxLF1QQSSVJAauS+FYJiDJV
163v32+WgRfS0jZQ7OlZVsXhTTO5gt/H9YF+/50YpWtia0zKCXdtmh+U2/mr4Yb3
dSmGTYYmsq0EGt0/hWvIMhvZRIOmp0OPKwoKm0QYgGIZaaZOJQIU1P05L4kXpMSu
gUAjecu3h2LZzoZGJBAK7P0ghFzFs+lkxSPgWnmwYfXjtHe9Ky7/kciIiY3+Q8pk
XJXVQnPuche0GHSeLiFEZgZFQR9umCLYo+USEtYOC1xHlD6PX30vtkSeYoR2iX1I
GtW8T5FyHv1dOX14snKZnfSFH34xF8wykzPvhEmmgY182G03yrGIfO05NGZSlkEA
qOo3zFlTiZYIrYDfWeR4Oj4KvR0PTYUhHZUYAGE5jSl6xWpRVqhdjyKSIXMONNpk
NiIqFvsC4QBxuTRxInYev7OMbTju6RiSiEhDwnpCBgzfe+ox2pyDH6XV36QEqIXq
vKVCzyo/n8kAsvTCRjFhWVFHmxBeQqx0r3aO+eu3FzQOUl1+lH5SRst/hZ1ZH0/V
3c+tJi3HKR206YMihFeYKxOOQYgIMrFntFPuUN4bFM1nl2yIqdAmz6C13Fhwxx2/
S8IRBchB5LUKJwZoreZbMT1o9jhSuxciagjbV1xe3qH73ILfdRmu53qLBqOkTI3K
BEi7ZyUfirviHoJ2ZWJhNiqY/eWNLNn+yf3VCicni3byxBl1y0uM68dyKm5J9hRd
+LJJKEO+WZCSj6pPoodsuDgfSUXWTtpe2RN5yG0GIbR+/hZMHPULjcuWagV1nnmy
/3i261xLT2KKNdCjmmfL/Sper6ZefHsI36PhObxduW0wChjFA9H1RX0J6A8kWr/O
w7DGYEzaNnqyrHHYF785He38uzLSLQJ11xwvJk52DvAxzof4FhmFBKiUWr4Pf4tf
ZAW7ztgJTBWGsJ4xQ0s/YuDVWFAJ1w0edKeGCXuMq4m45QalaSPawBrHByjuVBFk
TMqP/k7wkeiLiT1y3qS9bGs76ObdGwGsbh38f90JQV4xkdqKNxQaUi7uUo9HxKAN
dDh2zWWefdxv+TVL9IsntQjDDAG9LMUVb8eK6OzR6NPbUYqHzCuJFmpYERfDKQv7
7wSUxN3gake3o/aFwDvcpTq2JTGgV6w/58aoMPL/0Wq625VC5UtPH5lC2XHIno6X
0nBHojC0oC70eb1fjID5YLt4PMxYKaP9pgoMCS6DKkVDp8Oa1Ke5Ya+h0tUmYaQp
FfU4LWhabH3TFVLzgEj6++x87Fn62NGQ5Q9ARDoCTKuaauaVVPXUZHb93B6OzOhu
c1oShQJiKcnzF/dO2b5PItSPc02O0ropSLOf2RXhikGkkxfQL3cl11s2/04KVTG7
PMlna8nssbxT4nvXYLBX+wWNCi/BCOiETeYmJxIcnG8d2/WG8m6nMwO7uJCTMRst
ga33T1JDhktNVqFWZz+2+8ACwHy7d47oYKch46UD9+tXQiJFiclh8Wuh6Xmc3BNq
xXHi87ZK5ZudBeqowz9G/KAgnQIXtC92K+ZC2xTbcPmqjxiNEoOuiUKxDtW54tsi
dJZCH5RcasOQmROHAsuJSez1i36ek5xBCCbCtZPaw6uqRFth1bFo/WlJsrmV2dVn
5CgkDGJUKjgOUgawkmrsOHO7r/QrdMBROcfSPIthn3ct/sWi5GAkFvcJIpOZMGss
exBQZNFbXLS34JTI1y/gOyqDmkX//Y6tYLpQGXoONIbuX2nBHET5KRKynY56epYr
ZcJqaPmHNTV3Ke9Rnh9xviJIhSNczSKIxHZD6HsxQjnqiaB3DZbxL6SSslYtqBni
EJ2NZ7SO3jXhjUQ+vHr00zDuNUHOnFVmM3aAEEO7hQIG16KpytOWv9YtX9UuUY2B
4QKYGbDr84HKAyje7ndxqC/uZXAo/KIWo+bBd1ro6OqjdCjSBxm3km47wGhNsY5P
8R+WX2qQJuP6maQQ7ZziCpWUxV3bX+SNCsiL9TEmoCbBbU7FwKkbBf+bM1WD70lZ
kiPnq4onvNG/60gKbpUgdtob8M/NIzq+ZuXDND5X7lSX1BTpPGGIRSJk8LtI7rb3
2tPCLQI1Z8XCQG4W9mryBqA8QSYfezuzlFQcwuc4Ndg6rCJSRAx/YdrELx8Uln0N
V15Fvkj92tv+svrD5ypDOeTJyF3K4pjK0CEutG7C878GlWyMg0ZpS9ojVMzXW3IY
KnSiLJHRbeAeGsqoSHze7og8H2dWwO2plGe46pJhjD4GJIRUyh+4IwNYPO20iitR
JpTvVh9pB498UYtLHQn6IBbAU7AHYHxCx7JkownaC8vtWcIn8F50Kr7KLhen3TXX
eS9YTJkjlE9aGqPjYjyL2v4mSSMhWS/5OBiNqfFQoqICIJXmHZMeGMdiUNxD7/rk
SZmyycx1nCyiZGxPmNF1dS1wKkYFs7yb/2b0q7KakLTB2Xnv3ESS92reRhZmhAIs
gNdfzhEwvo4KfNQiuWXyE2o8CNfo0XMeZj7Leuefx8f+bb+iAqS5FCPXfLmibu1x
9sbAfNw94psJMn4/StKyqvV4WMOqcovnVy2YDqON3Psqm64JQxA+4bFuGfexfl6t
BHcVRjKxE/t4BE9O9mS8b5+TCCCLSQU/aRMQ7iQpEegu3JfQ8zAcRK3gdh/QMDFq
qHcy6deif4UaLXniU/ztngQJVqczfSEogNlggH/NlL4u0srjP96It8OFXmjeuWJE
FQD0NomPbxcYOeyQ5xlB9yNojPTZi1v72QEIOfy8xokxN552Eqn/mPBDo+yynTe1
w2praPTApl6uYtdHfmhCCihwBOIpEBpjYBjOsbuiZr8QD3SGNND3V7+2TBRFCQe0
9yBaVzgYGh94KxeBNoA5r707qqCeNK1xau7X/tZJl+EaoeaneGK9L5TK4uALG8tP
kHeVVH+klrR2pU4NZuZSKihc4b6WYH07d9NI5zUjn/8LHpHD1/QOVE6yr1q9CsXF
xeya0AubYWY51KsLDv0aijJq3KXMbdVzfyckmi1Z659jVr7wKqHIOym0qvioLdW/
2XCtn7bhEkKoJR1QAK6XOV/Ygxt1PsZzz92rlt67PsbPrUHHJ9LsBKYVhQVxgISG
WXcbcWhSA8H/Fkf3SrAacc359dA5My0fx9qV2aEIYejaRVDJvFirMLcTtLUKNIu2
eoJo5h33e/2/GBEfPolJlyKQ1QgN9LZqbA9i2rNiy/EPzusPjfd5NMv3l27drNAR
Bux4TmAHvu9phYJGhiwH+9thwpobK/UK0dgfnOpL/KXFdHmh8zRPJTCtV5W3r4Q8
C2W9D4V1EppvIg1P05a7TUbuiAZ3VhfG1Fn5looQomYkZcbFtr/o7WfrA+8RUnDl
kb1jjucqRoM/nOVONhDsgg0e2ZpCndbnwoCDi1UgWyXBQA7ZasnTutNn/kh+w0au
Q5IUrwKfCbDqxOg8a+SbAewG4jd037mG9/18lXW/7N8BlDwg2mq0OWYUEUbvR67U
WUPhNvVruUI/OK4U6tUZU60FlSlirrCYunCn3HDU2eOuEEpHukRT/sSbdze1gAQa
f2hVLwpKuOf1gNBg5O8fvgiOj877tVnCXOwyCUfNEMTbmQybmYQhFoYRp25qZnic
L46mOnhhz/vw2xkw8mxPOqSdsSWVst1JxBl+IvWLsut/QA3jsf/Jzhe+K69cEhSX
4mAk+6cT/s57LlB+NjOhFkKJB0wKpvyL0hlvlq/LN7vuFPn9P0as5NYmTWGvex4k
s8pV8GbW/4hv7uCa/hQBeY3p1RibnKlSHpC0z5Q7+ycLwprudAemGlPxoShh41MF
NpHHWw3nYUbY3e1JerpS7FXSc3LCiYgZwhjzh4wn/p67x3sjfgn5uMOU2ILkHGwj
25uRmwKqRDKHqc9otmsjHUNS1XsJdqYXr/2uNcQ3MIAoqCQBVPBV2T2wbI0O9NWG
004nvczQkkIEa6jAVjaEiRX0AGxA9T6j3yGQiBgKhKU+C9PtXHCcYekhXcuCE9aT
z0/uqVBBPHaYne6xNKtjV6128WXHK1voU5dP0VBpLwkJ5v5awBfUsH3nMl2cJ8BJ
3m9Xxxs3N31V8e/UNCB7635QBkBs/9gGVX4/OlPNooe+ZH1zWOlepLMFWFVZYyJL
WRxrfAw2a+yG6dRj6iwgkvepEvck+oZb6+og5iqAtp0IzkinPPwL9OHA/+x3uC45
lHS7NBsem42i3a0bv+ABshYGAJXoNrxx/niPuMAfFoomK/5iGcB8TfLR1tVHSyWR
4+Vh2ux8iI0CRk+EHUJ9O7IWaXPuNa2JrohkGDwbT59RTN8dEqjxmqiB0T8ughMo
iJEUWgSM0l3kbYX+SaqZPfsZ7lInDLBfHigW40h6S39+g4a7OkWDcA+pJZVaFFTj
L5QVL6ciDH+BwCtt5UT5A+FNHHcWCTdPxEbhfLPGYxVU+niORxF5CwzGawtOhv3v
peCjbvseuOUZVdhbEH8s3Zl9XKdI/15mvc2eYfPndJTAcqBBGC7qYWlPSW4bBgry
OsJdUQiHbn8qkzDGC5GKAWLj/TYc6CJw2KpLorPoROn4uurMPBQNI/rzrdZr8wed
YHQZxmqZq9eUZc8UcP9wqUsO8KvnoACYLyqzs1NcrXyzMWsCk0mn23ic2SeG+riJ
D0BevA87NfUriCto+KTMWmN2mwH5/SPMqWLsplAjWfCE0ujYzHsBS0Kcp0TbdGWI
oyFzKJauyZsaFlZpYVm8oRYNXzKMkFA2EAl3kn4jk0msFFHkUAryB7Z/+7QQTfEk
1z1fWxworBf9ciJ0r9dAVgLnArBcHMngLTdG30jfIrESVs8TT1QeCM4Wy2ki+bPf
5hwT7ueDEE7dy73cHhU3icedaPArWzkY2qBiLPHsCBZGXhGiH0Sl/Kogw5UzOPCO
pLx/xopYLCaU0Y/oCZpyo2enaiDhRP+V4BxbBCpP1PK+SoO2Ml+NMX4YteKpoyQJ
378J/f91uWuVKj1p/UUyClUT0fkIE4CgfKZsYxr+hQLydG7fLRd6qT02ZzQUTPgH
PmuHCUKCgBT+jr4J+9xlneoI1z19IcPoUaGOpINddFm4+ok+k9C65xr1/LFaRNA9
UQ5t8sXFT+FkUNrozoAKoHajmxtBxZfJ+1BqO9bXplHeDixIvZY0n2K8AWxxM+S6
b6Q9EybM+x5yU8ZwkXDUHihkKPM8rKPQNnOkfRJijBVgazszB9uk1EfnP/32mAfv
PSDm1OIEMuzh0WcaLxXLBQGPouGmaZXMXqNwoY9imu/+icC+pWo+QGMTtT2EHGy/
U0lmJtdPL5wP/LwvlY6fKi9+Z87Mg6rKrOqZF4YsxOdpP9I6jGh2BHgGTYzrC39Z
UPoPX7HQsH7yJSfIgvomzcTefARI6X+MaI9mq7G831LzZHjWgV5dsU4J8ilhxpZP
yWYd1U3MDI03oU8Jo0Q46x9wYx+IRpVww9FH3O1C7Pc/y0DUGvaynpzs81nunePN
doEkfgIv6VpqqjbfpcJLYLNKTcIxH+/Mfiy+VULD+nbGqCLR1EEC5QT9y48AtpAM
5Sph8F0uP+PXV5fNKeSEhwAk9Q3qvKAcDMk7bNCykqzgvnLiHbPdut9tAm5uUsMT
F0PuUlNM8B8jRhV5Q//JjsZ40jcXMnIMS9MULOKrVIIpE7BajnN90KgTwfjz5njO
fKzgZU9ene/7TwUSB0N/fSe/i86OID/8fuIcpAOlwbWGVk1PfdMcTD46AlC7fFPA
td0g2N/1fAscNdWjOIf/dkX2q6kcHFyn0K9LZ8qpBB9oVCYcSl+H1Nx5KjCH8xqo
ZB866v2r2nUnTa4RMs8hLeTc09Y9F+ull81PLHjO2pe5USTmNtEkI5jY/FYbPi/l
xeBQAqtYtTer2ZqXst8x7Pq67ebREL6bvZVpAOORXVJAUOQ9AtMCb/8b6s5yO/uU
L1GtPs1LxcYZwXzMTMC/KOSpuuDhw0cF7uBptzbhz2YUVcuDRjE1nXMZplG2hgIG
dZLruvjJdjirLNHNxT2RnesRshsdFUJdH8mF0J/x5gjPs6QbigeFlz+O6P+frSCX
TCTAcVRkTFjGxCBjielnBLgCypla4ys2RZS/8S7biYBOv7F4UZ8nyo6QqgwWTVsB
pDqbMGy0q8E6gjZpgm5KdT4LColLxXazBvxj1q8asZHiMyhQ+ZdQ0yHiJbFRQRWD
fm2Wn+2tDEYqct6u8+oQ/TBIos3lL0AsbZTkZnH/IOg33gSXWDCtlCC0zZ/fE8Rj
YrttEzS5YIMgRw1OHRfpI1VcZGCyS5jQ17aybR7DnPxWFjNF93OnKAT4Zyxv1QFD
iGlWVvVG2lgtv4XDqLiN9JW+8qtSYofSmncAbCtHsPIBc0UcHTJq5lqnlYTrQGf4
Vw7M6TsF5Jd63RfglqQjRXhgUz50fFk3WVCF5yX4njFHTokXty0eMNdaDFm8tdg+
FhCwDj7hEKuKeMVeyHoao3FrGuZs6V2j57GVqwnT4sDnBenfCdfi4jLXvQmbKOgD
6/kRuP8Yt4tEjSd3j7/K0ezTPwgKXqgoCjI5tUOgNLLSZcE8cNETJfpSvWlclhQp
Fea9BWDNxkWiiqVuwY2CNy1PuA44JaxdUxj7+2Nx0y2Q+NpiiJUZUSJMMgcakJHj
2ie01CUOtoXeQBf5IhBy/knZFbx6u/xA4k+dE+p2DLJtsw2nMSLVUF4wbL16AbA7
3jsSa8KnTc6GDS9DabO1FpR+RsSducFcsN/1iVRLhWjot2CmBs6GvDycb9n5J8hG
hTVq/P2Vi22raqGeXn1BqZ2sOdqG12y17CxJW5B13EgnGoLHVNol0qQOM3VsePR3
e5tnyBWVAShVgrTc4WQohdglh44uPrxSpid/g4D9nmUDUuKr/SAvl81UL2kgeHkz
3GyVEQ6xCskKFrjkXQYTSISGg2XGVqEwLTZ5ut7O4IMagyDY2jr92ExclK/0FfEU
NNjduTIbYp8gL1DrS/ZXHPAGS1rU+jsfqq4X252UHyLBh/qH7Bsfi4eoCw9I6JTf
xlXJjVaOnkDPXHKrvXBinbhbeWZXfpKAEnTsRx9KDyGlsLo73whC5zo34AcI6mmA
Xq2GbRAuDf6+XTmUuuHQhUmk0wJbIdu37I0EYo95irnBJRFDOWFeCiPBKU3R3sTk
AH7aIS5Pnj7zCTDKHMlpUfXOF7a7nKOWhXevDefrdx8R9HxcnHw7jluXUMVNrJ3k
hqzxy4D63wa/VdqlMUi8+a1rQP84W3CEfVJyuWp6BOVvSRbska0RBMpBj5OMK2bZ
8cHNCz7TlfcPA+2skUfaSpMpCpwzaV2ZtEQ0JY8HTRPuMKiDQsc7UClz7cD+p6ec
q2Y/vrh7dGega5oatZa3OnRRmlo/6m7LGxeYJnLkd0RQr6jyx6WsAyfkxad4h9na
6pjJBWw+ZTwFVFCfVlDsRu1vfZ9l/ZJlPYWOo1Cqq2UUWKphPiRfDaG2qSOM1Fk/
iT6vKHIakXtf2mDEGb3UwQMMMiqMEZDM7r7ryAWW+eV4cVzWBEm+X/HqaqK4ZDE9
ehGqQvuodXcE3zoYNfJQGXCsiV/jnwLpyl+j532WhNhHZ7BZ5Db/ojWC1KolTF9q
bdyR8N9nSc6/+7oPU7JKjMiA/3ukQb0ao3R4RenrbT2q75JoksAZxU7OLuWFZwND
QJ9+h1jlJyjwjckHZExOjULj06oUal7OqG5NedONydgkt7HRkzllpDyYlQD6CSCS
yfAzKr1Yp451/B7vH8rge0WTowc0lj/vSnaCqRuX/uZs8mny6SzMEHF39ZCsrRL1
8fyJAFLFJHQw07uIcPwLm3DVKl127Q6KQmRNwiAeT+WN412IWVsrlppGLgXQjrF+
DCIR8JL/z0WsWyYAmjqKrUlQu4L7stWU5A+5tBN6yoDo8tY3ZzFBrU+WVj1vjCpF
rVX7jGRJkClubvC7QBXC6TadMA5Vi3pEzhIHvpKwOSF7XqWwAAHtd2C6lVDWpB4E
BrcRI8pbI7lPseh0mOZie/6ZNnoYjEQ7IBKP/KfMsvgJo786gR748qkOWj/Jaaxj
8Rb3Py4ULHs2wdaBoYCQyjqeFW5aomXAh7jSNQWWz934WynwiSzdUZvqMFj4xMtm
TJzTWf4o2YogEfMte4ms3qiNxRLna1+Cu3IAtSG0NZDQwRY5NpPh+mU+/Rayscuz
/MaO4N8RfCfhD+K3POc72S/lvQvTlgEvQyI+bTpl0s8W24/sIlXXcWbdBCFjzXgq
GXT4Bt385460ai1UkpqsARfDaNo4m13GchPvUP1hzs7eRUDyXNja2gJvvrR8EPHl
IoBBkZsHGfBdJWX19CGUcgpB5gep75o56LzhKhFDVQOLbYX8wKouglGGvI1o3RA3
t6Di/fF0w/QYQAeGYCgiieNxCbnTGlS3pc++NN+QlWPeDQY3Q6IEMhdrGrkmBg6j
S8qG46/Qh06lxq9p2wcIyMgnB4gDfthskDl2GZVMchhcNqY6KQES2GaWuMu0G7e9
HayZkyAKZoYSKVKmtMi0VmT5qgPLbvsxjf28snCgmxiXzhIlhI4Ti5jmPqiAUlZK
OPhL+gghi8F23eOh0Caes+vkKOvqK0kiDCJet3d/EFhGW3yzFioivBmlND/wAFP8
YHhEwTl768eOmryup8ZIkhLaJ79M+uhL8UlXSotQKTeN64H0eLUF1pNzHlrhl+UO
SydDSB9eJCygnrDcYVR4iFcZs80i7V8dXXogsJCOBgnWFVS44xtFoQjYu66rDj/c
Tx10U0gp6sDNBhODzxHeuaEKUp0xQsz2DhEx8raku3fAUgTqaq9RQgXNwdjh/7t/
AOmfV1E/+PMdqNn/QDi3NlSOMtHxws3OYUOiXyDySewUOEICfFc8WjNcpM+h39T0
fFLlwQKAZ/Ak1RwIzFoFYtKkNLAUNe1NZ3/dm9kUdsHVfR0ziZci6mwc2y1RavHw
Qb0PVXku+OIo+YeVY9tjQJb5c2wzs/RsgT/EmWqSLOOz5KtdJyXfRAGqEctRELzn
vcHQgANiQ6a+6wGgk5QoJ2TDIyS4IkqL3Op1HvSzpdvP/9G9AyUgM3nVmmUcrVMn
+A5zpxhEp1DG4PUs8NAwRXKmy5qMzymDey1PrFhkAbNotqJ4XR3lOX+hEcUcRqaF
WA8LeBTbzpjM20JCxWqOtSNnMoT0ISp8+QjcCyzffuJYMUSyf/Mrrgal6hUHFLw1
9Ejsyis7dbQNVcTQCDz1Ys4mQ+eOgQ+lgsTKD02btAv37eUENKAMpzCKAPmetiJI
L9cp/Ge/gGTOCSEmF51lmXx/pBDbSJNm2CjUxXm9aKCNKhqzC0nmTCjqv60psPT7
0oF0GsD3oxemPS5MYiRs+1nTck7Pga++AAQi1EGrhTAT684vcLYx14K7CMkdNjEF
34yBASPz539QUpJ6R1WDaKK2iTle7XJ19Pk1J58VkCdyawsCx9/C5olEMdIGA4Lz
fbI7bspc1nviPpwwUTtlOrS01AqCv256K0qc5PxMzGRlB3NSsj6Le3Lty+/xZmGR
ZwB93UKiIQ+pgYI11fbXu8r3J7fjEpsmfp8ANobKRf4c6rHBGIIr+HOKK0xCY5Yc
0Paapvd8ERAsqT1p5F4bIxh02tzVDTf3OeFFIoKad844XAKraVCaIq/eQ9hZ3JWR
PGAAA80OzNgwtp5gUmS2B1acXyfwM4Qa3owR5HoEdkmBEDY4Q6uiS521hXfywxvM
HRYUOSImbEzbLqalAtNTk5QUYa+0AtNntQGjH0w+Ju3QbdkYJh1NhPclJR8l3+Nk
SCvlhPzwroGEG9DYcw4XA2aJ6lWeaVBBLSVzwk3TegfOnwlxUGn5WM67HMJpn7ZE
U++VRmLmbqoRiHAi3hTNf2fVx3AF1tmTrhirj4R7XC+jxKDIOVB3fVVbs7DvevkX
zIsYz16pmwsJ2FC/G8c6l7PXPA4tD1dC1K7xCSddDzvOCZEcBKmGVPclmT/EwoaP
OwZ+50McmRUgCYfSjld65RQVbPCEOxKbkGGAA3R9NGOPh1RLdBqM4wh1PaDvGxzT
7KrOh4DuWX80Kj7qRuXAEg0iXorpYAem0fxQqwlkPJJkAb2lcxOrDx5mNYNMog5A
nMLeAuuZ2uk9D6hR+xLcCiXXcg8jgHVyTgYGsdnhvdraDD9JBF04MwDTmf2MpYvp
8X07zNN5Nc9/b/bTttxjmAH392h34C/DjYY8QGORdo+Oia6O8hyu1VvxIbO0ldTT
CHUpE/pdnPPQTYUK3knYMJ6e6aoix8zJANixZzJq04Dt41J1F5XftVgs6x31ZVc0
`protect END_PROTECTED
