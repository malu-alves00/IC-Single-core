`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
v4+NXXEEiYVPdpZzuFoU5o78/pSsMRX0fnI4jhcMqe8FMb+AmHmUXHPMT8eBt61K
P8U/EftomlVvb94wHf2YRmuHNb6eDWXrIBw/uHsHX1T1+G1SG9qsI2/erOL1Nde3
po2nFR5ribKFnVfgrS2Pbec4gCJ+LQrDMolrkJlGmB3NIudgZ5w2z83DE4+e0sT0
Odc+hGhPLZekR7+R+zsV8KQaWjBYgmS9n3oAcQT/u7NZg5nusEIrsQI1YTNuSykJ
woptuCxcX3eYJXcpDZUhviCal2FTVto19oxBxMpgFgNFZ/AMwhrxUxIgNj2S4kBK
2dB5lUuz6EqMDfamTfLdkDf8yEITFUTo3H2k6OwXV1F8vy6s85GW0/7ygXDUcvdI
h96OaGjydx0GqxEXN16KzqGcLeFsr/oCFRfQHDu6eJutP6LyFV7R53W/2CdvTqSm
oC9nRD2wClV3R8fCwXw5rdqllGgYt4AW0j3bQoj0efIQkDjC54FwgJI/BgvCA/dU
MlJAqoYR6biBNQ9KP54fQ8nqlZnMfmGGqFMirsE0DY2r7/VQNWB2tjxVtd+eoa4O
zjW3au4vcfmN3CzgOfeZa5XwDwyhUXM9E0bj5lVnKYl6gF7wOYuI3GH2yUTeTKFw
Q/pxZylcy/C1tVhOG7NVnhOsUlV0hiOKhXWP57GrzyolX91AuZPVFzBHEU41L8Lh
Eo5nOyPsH84MVsPVlqbHSJ/f60XHyYPdB3bDVIc6nhXtv34PL47QVZETliKZ+Cwm
aoC/2o1T9oq9M6XplShuaz2/nt0VEpCj66NrcGQP8wVgen7hkx8HNdI8LeMiHIu4
tv7tb7tvMRwwTp5hHYGG//KxrWHthwEbFQqCMh95qn4z+mKgYkgtP7R13ZRzDi1e
cg9IQJScKDufYJa+soiuYfTrXrR00p8lwH+GLb1yMy25XB9TUNzqiNd09SJ5YS6/
uaGYn4leNk/u6pFPeLCluQnN/1+t8Zoo3y7G8VWE5U/FrtWPA4ShUC7psskLcdTf
DYeDkrf3m2tEPk/L0n9pwFiEhbaeswTAfB5lvMJ/SE6uYmoCsKGjZlp8X2AUnicb
X/1bH4a7jOIlkpHgFDgRFa8o+fNlkrDBHT4xB0aTP/R8JZRn3n/s5FXDHvb/jiBF
X9myCp54CXQOVGJ7+rZMB83i12gC9UR67k4VtjbTh3c0e622nxnlVp2OEr8UGoaZ
EhjQvzXJu7ui+oTI/fEtekD3BC9bLFc0+QNPuPtjX6o8KJ1lYTtiiGN0IP2Sw7eF
Jjd7+CI+2ZHHuFjxt5pkK4Osh/hCRD+FYnw2T8mkzPe58FGoiusG+s58vt5zemBh
hUKmtLLlsXnUsnCuxQj36clByky3Wbn3jTKoK96r/mPVxG+2ZYHd4c9LwXdvGMaV
OgHep4LIOG+6CYrTGrpsOZVbczhQ7CjSy1q3Z4da9Cw0+BbO19XJ+Vu1EsMuT4ox
6l9zu20TTpvIreFPvTlXKkc+5SVDYW9jT86EAONH3ZvAXff6dvyTY+OxMLrf9Ed/
N6V562nK36nR9mFFY5PjT9kHK4tI6RZPnPivfpbxni8Xwe8KWhwHYSQT3V89BGYw
X0M70qG6JjuAJTP8u61Y8VRvt1GgKrTpQiZAO5heMxcYbvjMj5Fd8wEyxeG6ujRg
sViDSTbfaNuxM8LeFFpjXG9UKBLyNgRtvQMh4pdedQ4lrFpHARowOWDb5erR2c1a
Xs09ESCtp3BnC8AN5F+rGvVUNJ0KIvXnaHur71CSW7zNiIbjlaDWbWlZnD8kI3AV
k84jdpLrtawOh2bF+sU00WpFP11VULpV4X71iGeDpR9VaFtfWe8z3Q98VMp5jGhD
rGb7FuPXzqhl8uucK7YdK5gQI3tzRwNXqi/l2l2QebHrGqUGtPlCu4pcOQraRN7w
DtsmmOjyHw2LwM4vEGzfPmOiJ58LtBpR3Ms/+w/G1U1lvi6KqkXF1oWFyQmosLxq
MQqE4AVpZNTac7++Qn/vyDZk35van2njZDKusdZZdN8pUYqHBnbDFEsCjP/B/3jq
AaBdy2Xf4o4VO9OCf7ACoXUDhzulz2NUxJGcE0OU8TSJFPcFz8UyvWZAqnPX15KI
WGVRs2zgaFh/K9IS3cAQisLHI4UXLAoylZgd6fimzSDc220MkjFDiFF4DC7PHQmH
r+JIKRi5okbZLpSxFN3vNSNbraIEkr0wENyg2tliu8UXnyVvTr8605+H7eBsWifI
ODIQJoDN9t87+gh6Pody9E2Fd7Du0/tFxHHPZ4EQuEIcA8aISKVyFIWkaNS/B3U2
/X3flYXC7JhUC/K68On5hwdqR4VPMbrh1LJFm9xgf5tWFS1HzIslH3M6g0aEFxnz
OH5ZsUFljLfaRcQemQHMMLaBRVbhVfPHMu/qbd8PA2GhrQvVjdNqPSdlT1QHeFYw
Llw2t/x39j+ovXrxqC7lxf7jaC/KDqz5BR0x5V+5T4iELkHlP+30LWsJaPOP0oVY
uUNzYa7p6QIo0V2e/4um+zxtkjNlEBx4xyHRVtmJ84YoU08/5BZLaqXFbeVn97z2
u+e3GKplPWsxwfz5r0uynd5Pr6ccTdhiGQU80h+jpwL3ewfV85im8rP0qalfZrt2
8gH2qDDfy1pftYLYbeykujnh4h1BwZHaT73zYyEh4GK7EOoC0c9IyQyPfxGrpwPI
hwcUkBkfwJhtol9dlH6oA7aIwYzV0OItLIvoV+f5/d8iLJhMe30IXkgzYH2OB/y3
wpRMzt3dkc0EnQZtD4Iu5XBnLDxiFxyVaOgKJtQg4uQdRJ9+vg+WNRWtE5izvj4V
OTzbwBrjdKJt0rlQg+Sd9dddZYV9uXXHQR7OePtSsw2FlB869FLYu7gZZkU9SHEY
pPaIrqkht5r0v62089y6BDlySrb4dMs1tYQaR4cWXHel7oV9mTAviFGdYXHXUyvr
reme1CrUZ2mBFYTRA7bliAfzAqhfZ6HPImTqWQpGkxTnAROeVwEwoe0qSrqYNn5/
MxnZB1NBml1hZRqjpXaeQ14h82h89soaGMfR+ngcxF7vqpP5iK+jXsXvXc2q4cL7
0TK4fmYK6qoEpTcIJV4bcftYeOX++WfTj25lGd3NJPTKdMIhNSeXBxKdV4SEi+Pr
eFzXyXvOkUV6igl0uuOmvvkGGrdLM981WjLO60DZ0mpNeqTIDqAbIUwByhi1f80V
y52fYp7ZX4rv7RsMtdBWPae4wbIcI1lHLdbkRAfa5d5UzPPyMQHs/6EFWBbiQTCS
5tvNIPoTaG1x6fCCfW/5SPbkFYT+Aubt0LlHKbgD1wdMfKPvKhIy4sJfnA+bQgpu
rdGREyJ7v9FqqjHwNlqUAzwZ8b/4mGrC/ZlzwBEA7ONtawBvY+n9r4onanwb5sp7
uAWa97W9O7bKH09XscEYgu9PnlCgApUiW1+WvR4X5jjbIhE8jKLAGFqTZ/5lbKMg
5cW9VkBXx4yd1R/2Zj2Y4m0cEH+h1079utkvi27qWRV905/Pj6vBbleaWfe+ZxvT
Wwvdss9SV2G9af8Xi/E1WvjP1bdNv+34a/uXyY8N/peEl03tG1AESmDQ6ejAzY3b
0z37Pa2eLnC4B94J203pzYveXt0RHq31pDZsdZfoO2I4Ko+au68QnKIZub9cx4Lw
n9D0xdeDYOZxv5lPS8QnKmprxn9flAUSuPbWCYvdDkZ3HC4jxlYvK+kOQst2t48I
kJ4Fvqss0AMPXqxpiREGFSCTbvlW2kJXkcf6P7vXVXeES5MaWV5++XRuLpdzxuO+
C+Vanqo2LbT6grkLm8+Mj/t68briFUB8x1rB3dZunRjUjuL9AJPv4yyOvEk9NJzV
jK6Oer4h4mw28Qo4uDwpMVhk0ERa/X3L18zn4gsDicIjhDUq6+o/QSzLtOLthAqM
aKEUDaa8pV6DkgjK+C7oELu/xqx+DjKZ87SP95rmt6SnD3XYS+8eytT9Iagl42Y3
/NBmHh/VH4bLmgJ6K9ufqSRjuTlctxAepMTxz7DcefY+X6oHoEGJQsea4sS7GBfz
YJF+7eCkQdirnfe70I1XzgwfjQHGjq94KlUKqN2lwunewI0zsGmEoxJfTNq9YcB2
0+01wk7/qu0GFbVukDLTKnoVk7ZT0g12E8k7ysQGo+OnK9cQoKfz/exCKW0C6WRZ
QvRLHUuQlgCTl8NWnzUlVYgVkBO/KVo+1cs0qQ7Z4DR0HkM0nC03Yqzs8cf+ZKMS
kS/IJ9w3pve9AC1K1ZCgYGjNg8BEjTXHZPgpGOKzXzI4wA9RgiS75betv60afx0F
BXVSy9iIGAhgg6443xhX4MZVBZg9a/lyYGSbMXwFkK8gEK7q51lrypbCEW4JDJwx
DEcy3V+BiR55AoFVTjfAoBoDxCN2es9QMhNGloYSTwuYWoo6grxKbK8mQiQC8//V
7uZ8/p5j1c8dgnNTeZH7bUQKneokmr2qOAO9gZT6TUzB0fACD5GJxhPnuYxyoMOS
Pml096+1l8KIiFsqy/2sQKUcU/5duUxPBdiEwflmrMMK2XqXh+tfaOiw8b53/aiw
bEpZ8aJ7q/13QTm1hqTEjSinCkwNUDPRdkU/nKGHFjUjeJNigCn0pit9cRM3UCQp
9rc3SjjdW42RPPbkq4yZnK2eN/7kezpSWopu+bbxTFxIgJrE86YTSYfcib4/YcYp
pNORx5dB5M2bDzzTp/EXgnKDbE+33uF0ZObeHoJA+xB2e1hrB8ZJG/CfB9Bj19+R
8cXKNJfn5vTj88EG1uUCM8AhK29flUBYiPTF9d1WaG8ng+DOZi7h5lirePDxK1d1
r96r65jiI5YFbgo2MB5Z8P5Jv6Yyw9byOgFu++WOCorrh/OIOa77A7FNbxpVsJuj
W+s7SGJBAE7on412ZQgplTeCGOMsDR+C0YR5B+iwU9EsXA+r5QEca7NCDzXZoanq
OZ9aNrdh27DF8Ne/xL8kkMAwjtgFaGooUiblDVv8j/EmXJHS6O3bXm4DUw1hI0yR
kdyFUm5Zv0j8ZuJessGqbHwT3sKv9cOsAEz/VniHWhoQG/Vt8zmxyMgtjzCfylJ1
TG7gUTa4QBtp++6EZXRXPPfqoFCkcDWSaBVBqkdBW7tEd9UVqnrq2CR7zEuMg8A/
b80gcfRNYqY1/FR3EFPOGmqs/MqtmBdjV5r1Yx/oStSXSbO8+895vlV65yhm1skJ
gLpEidC4sbr74GSyW39qRjDkYw+g5ANLMr0goCa69XnA0rfCh6v0Ls6K1z4trRZX
TBKZxrQVhDiEWej6Fbx8WpmMMHmaZqmYPMO+HNeE00JhJpRo8A8Yl9QTc8JRgWsE
4Os6iJF6bf/0dDKv6Z175ChI79cOnipaQlo8aGEYZHvCxSAyaP0jKD7pJ6/ENB48
/rhGpWz7NWxEyDCFI+U7yG5xFjGnjG3bFX9NtgCMWLfw2HArw/7tzjZE8SIQQyzl
1wAhqsI35oWZC7i0FpxlpkNOBxbg5K5hX20IDSo3GgqTwd7O938dHEW8XvkyBzYl
yi6wbZ1DEakLSdxDxD5xyFk9klb05AnjyfJH6BwisAVYvpXNJUqshmTWzjtWyLfC
QWgi4jHXxY9ToW1LcFiHIdh1NB8nA9GqqJJVof1OLztJgEeMnvW4ggv9hDxNwGuJ
+N1TRTM+RQEHR+dYBYPkYaQ9S3W8e+Wyb//A/sGQZ7KPAaoGzsoARj0kuz4hMDpi
98RvRKVjKE4GiiEV7BFVsgR+O21cI3qezYDY2CRT6avKRog/j34489ApD1fbJ5rl
LXoxSHQnFONiuvYziVBbZGCr+7z0q3DR745focCdJwX/7WyzCo9e+T+yglUI13EW
82aF/PSfmm5BMRyEwyBPpUbWpgaJwcVHLYRHhKt22mEqqctuTcztWX08PhDwbep/
2yjiQSMAZYGvVjqFZGIN/AJPRceu6nIQUNdLzgjS004ZUim559HRe1EbWm88Gv3a
1y0PVJNfOGa751nAQGE43fLKamBFpGbOKyUOP9JI7yFACBPpj5urDarvWbpr4tc7
sN6SBlixlxL9jXaSovIylrXiQNhifaQUe3qShqsvRRJUH4PQ1Qb4cTfeAmtIIPrT
1gTdBmoM2wuxqDZBN7td0db/7wP+k5IW3KQWQsEPioMpGbTF+LaRnDibk+w9pxSd
WIqGiScRGTs1JCt2MWNAKZ1kZWy0uZESkAADl93mMAG1eHsZQoZcfJwde+CmPGkh
PU6ByUDf/+xmROKWU2C6nLDV3oKH3XlEyGDeTgRr6Xeg0daCLBJvnBJoDeOWv26T
DxT1jBg9gQGraz+RKMSxTWSTdlo2ulVwx2iS5z5OosMoQaqD/KZ18QeoQF87TcIR
Ly0+rZ29vB7QiKs7oKR6fgsj+rJoYOSHpYE8xB8HAasLsFTnVfKmbNv94FpYPZ37
WDtsLmfPOHwtRW7A+1GlJowxI505MeQh6oxbyNkv8pphLNuBo5o/CM+SlNuzjO7D
ipfZxZ3jKan+yOgEyX5IR9LveBSHP3LktAYlk+plAhEYzMvOu9Ze9jzNBg8ZKY41
cMY2E4G8eKiT3ADUoLOaMARvfOYyX7sS1Zf5SB4BIRXfJVBdnJT2TvgLOADTmihF
bquKonQnchv/AoCrRkNyOhHsImoDoxdwTV7cfOLxboHzyKLrdipHTClPbdHZr468
03zlUVp5ld7xeJ5fFL2QHg195R9ZpgIVT6tKDcfRMLUEXmClNK4NLwfubRG88mZg
ODedboA9TUulkz2zLIiNX8Rth1kWuec9KjyuqzsjPUsu2JM1My0VmlizEpZ7pF3m
xuWCryN+XveOgxBkl08DFG7KIPo2K8gubU8te4hypeUZHjuq++Xq65CR5lKJexsM
C6P8lNEmbE2wHrBRdPDILdrYlJKMJm9lDBpKCbgfRDulePxvBTjgxVtydrq1h+Pt
NAHLj1Pm7qTqTEU6nZqQF14xqbT/b/e/UP0otvOntq660CzODWpjTeYujqQNDJmz
72hAUFcyjrQkPSD7ZTZMDL8/emzb41wx3JyT65UHUymYzN4NfSX2vD5t21JlrhGZ
iUf1Do3OZMHiW6KLePc0ou81+45y8+VLm/VrIAPGhPxAYl2kI6/3phLxTAD/2jc+
4geonqJvfVF5sU4IKeV6sTizcK7K/Fm9tNy3abO5ob2vnwj+PrBrhtmII8hMolSn
Xwa3Tqn4wYurWg/BYUvU+P6eNLRuURJO5IPMsKG5SMpQm2sWHLSmDNvClnXQoGIA
hlVri0h/hiPf00nmIW+CJx4UubETXdyTxr+R9VlOwJCy8ln4+CV6nuI41u+laUNK
r/FrJEY6aH9M230Ib9z6pClSjkQFTRQgGg9hBV39IKshcmvhyYLnskzDRhd7QSTz
zseToHSrAgVLAgfBPmZ2vTGpu1k9Sfxl/UMZHj0lde5j/HsZ5JwBnN8WgipaF7jN
CrZsRIBLioXw0BkuqVrRRrkafPh5Gch7Qj7Ig/8YJ5SGNeNI0UGnGhUX4WelcmWC
T8dKU+7NpaNcSMz3Od8Z6eWlT5mdpDwt+Rv7uXzzFqKH7K5PuSkaXT+VEJ53YhH9
AJMs9lAS9xoSFcrjhT2ck5fUl7tTvWySvWEXBoFBHKSuk3zBMXFBCmccQNaOzUpV
/wjRW91R7eldOi6pPdpsV4zEIILxG4DNfNfdrEGPhQGzOwhjpZ6YLrVGo7ZwC0XT
xg3EYxhnCt5JL5z52xtjAf8iGZjSXY0kSyq+W67Ina4kApq3y3lITAduCK8OB3By
mca75uAGIUzFBsZkyNeIafVd28jmPJjdqPimTr6QXROFyxfQ9frQ1NM8XMTntkoR
n1ZgV7wZ/aDcWCavnBjvk73wJ5rErEBJCvIExRH6pQGi/hk5nqb8VzWJ9bbr29N7
ksWVlLvxwSYaYazh9fHlJkWS9j3DYw7XnfIu5IgZD5NWv49qKxXpICgL/pPGvm/R
0/2lWAlGTwiQP7lIB9ncmID3lCs8jZiKogZuaBbbZMkDsVVF8tYURsa3T40JCUYY
Wl/DSDx9+NTYca9734LYZ8s3A8kHB50Ql1JRY8x4/BiLbgxyGwzJtKr+cZN3J3MC
7P+SjDKA4KimZdMJVqoUAVIngl9gTjhYKXLAOt6dw1ugJZaAKFNItpbOngYgnhy8
910FKd7fPocU95Ib2aZcpzIcHpSW9kxOozq6i4pGPaHJgAdf9oNmkgqgwqWYLFIj
zknbzO1W8WyNhFzzDZOflj/+D5fOkWaP1LULVNKr3WtS+GnH+faAhD9xBLmL8MsL
iVyt6KF87xW/oj1xmCbFAWjEgY+AeYZh84vCHKLD6WdLnEAZ1/e3hEo2QKcLO+Vm
Ly989nSFqdlhNM41Z8YKLJhwLALgtLFppVPTl7B6ERYcZyl3IVVTl5UvBrulaCLs
2syC/pNzyHK+1ENa4NKznGSdmAjWd9kTqo07ToOuvhq42UW83MryMTkb8NrnGboC
LA2Ia532EfG7LkJ5ggb2oZLrQjzK5cKUiKs4jXN/eTYoErZfgFKu/74gbU80TxfH
cJ2XnomZb3XrXCHY2/Ez3LjTB9Xe5tfqA/V9utG/07K762qjIKK6RvnuUwYfE/dM
wPJm44SQuXCfrCRMm24Pj871stb9XZX9zd+7L32B0A1VQn1bLqF+/JpMFNX6TpGx
BwhrietCOEBpBHLnmXaf5qoNC0xTiEnpxkbrnJQnNu6ePn+vlfzDkqEeXSPRter6
iwKX7FdCcJm8xhIESpcECGeTSbT+xB9nUvXUbaqf7vc/D65nBLBtNGixu/vwQD5V
NC+sQQrtkGjIZUhf9t2Tdnw6WHfJCp7n2KKcarfoZNIm4lD1zuGO1ijoffoU18yg
3N/odNyUpTzuKVZ92cc7WnhH4oehY9KM6ZaeRO+c3If3Wae78P6jSloC9APnKzxX
2nw+KGlmgxQeYEiDaqwe1W0fTlSnv4engkE5KvS3sFy+2Jyp3epIagcVU9xGvO50
/emz7GRHVcXn90MM5ibfImU865uA/wrK6h/xELdMhGu+nUiBLUFdlbuWXHXw3sjG
5QN49ZvbyUa2/r13H4WFgWUSsttVbH43N4QqjhyQyhMgcsvzQC+uNWWBNkcw2wZc
rv8j1fRVJkX9nG+AYiW1ZgxIOZ+lyG0hc5tlYyLpVppreUdZDXMS5tO72a8vsXSe
9v/QIZ60yTfhWTHB3qOA3V7Pfxa2ojP4YE5P4RvJtHAI+KS9is+09xpfqSDDcTQV
/lxnZCP3MwbdSfESTArBdtxpHlNDwnLbx/qIOjmPLF16qRRLXuMXp8ZwHfeIxEWv
q+Ug67QsV4MnFLaCsI2R9ByqhwtqRsOdDskNMo/59nCPRXBgG/8sNouXCZjHIh9C
HBd6ZJ/EshTE3rCkteqtiLqw/2Zj3iQdWIolvYxCT4EDzTZsovD+IZIE3DO/+Qm1
Kf/OPBaH+Y1s4CyKIcL1+TsWpkZ3gjwvLAKId1KvP1yhlrbUmEXGcOHIG18zxuqA
hMD+1atgfkmiCUBi5CxpQeH5/Z5ZqwUoBGD80QzU3LHoRxxS5BzAY/mwgXgMvcxN
lHDjaTKdIQKtWyhIn4bFmmeMSspZNDCwj0jkzLiX1XK8hftw8L88bHuY6Y7PjHAM
fNMTFOVJO4EKvontGiXKIMRLVK7nydJHpt/tfOdQ46NWUCyophfhQlchSE6F9d0i
RhVygiSVkgJW9mo61KPBX0OPpNxe7/7BmluCyckmStradTbu3Lz+yrmNXcHW7o6I
zNBSoibWHQaF899B38W6ZMq6zHHZTrIj3NBx3zfZhiJYNXXU1R7izUN4Vaz67Tkm
oajzsihe4gy7nLkN8k5LXTD1Cb0exBFCgawB6bAzO/UUIJEAx/OQZ5sMDm0sUJ6N
qUmhOGDdq9SMpuf5fdDm+apSH+MejCmRduAA1X1t5FFpJ0yH69naClYFF+Nn9XN7
erlOCnNLW/GHbDQtPFIMdlfP+aX/j6ORWBtmd6DMc6/uZ3JkhkuksF7o7E/NmuXm
wdTVVwolVto3Ipr6Edv/hhQwInrp7vN26T1Zp1+ozTjDyPedMbyeZe52PawbK2i0
RwG+bD7di/y6nsBPGYLIzkjTkgrGHdsK7kcF3zVzoafjC1upPXGyGccjViUdetPh
G821o0TszajiDrFtt2dFxtvjxOk/Zw9Gd6AfZbNCcLHGc403qcC4SMNO5VcU41hD
O2I+Th3m3WYxrkCQDmbNeLvGN8Uk5JxOKupa6SgTLms58oUGy814Mya+hXnVykfU
2FvxcZ1dQ6tUd8Z3A52IJPra9gGKcLMnlcGFnjtkxT2dZ49lM9q5Wcl4us2MMJPB
+pyzMwCqCF4X5odsewYxtTIaE93swutu+ntvcC45KaA3e2qbK0v9RDYuqTucoF0G
Bz2M7brnTrBSbdiQzMoeJKDadVDOFfMzrDQ7EqLfiR/hYhufQPDpO5R8u5lKuaxp
jGX2xUVHX9nQ7lP8N9/xvUyMpmnZ0nrIqWTZZcZ13Wdf70IWEm4tAHPz1BL6n007
+BZXKPiHoih/+2qrzbmnVgyy1BiVz+NaxPuSY6PqKj0eQ1xLINfo+qOLEODrrAQA
3TTZe4K3u+hPGtkgN3zq6LhtdzA8At/1xlBl/5dzekkBlXWCDHwt+yF9BbhGZuIa
EWFZUqJB4B/N1EQEX2JtR1aYIi68DcKwZhkAB/2qNYyLmRtMfywyu90qVMgKVASZ
tNspvGbmJzU5Ng3ICC0pS0sOut4xCX/i/Oq/kTWCaFMsluQL1ze0s+jgHe1aG7zN
I21NTjRqWeNyiIKoilbhUQE+Gm7o4GIzkUfb0i6nFO74mqcJnxScPW7bWAYoaKoE
V45dgiTzm3MpJUMIcJNzfxVaVRJo/AgrCbXXkVlpsd3oagx4o9iKUq7IIk2WB3XB
M5hwnRNHxE2+UCUDLMkccPQ+FURqFocNFXW/L+Pk8j2TUDds014BMfqX7nPO8N5i
zqUscNTyXWx8NC+3G5yFYNWImAHx9nd5VHjExZWqMN7ZGN2RyApbEfYx/e3uVtTC
uR6O0gQsLjN/gnB4B4IGog+oSLM6zZC2eOZyJzWf86ikopByr25YyKAwMN2UJ/Y7
vOJ6XzWxxLVAqh1dcMJ6gRC5PLwx5Sgf1UYHUBJqGMXuQTFMyw6mEiWSWL5G56uK
GUJDUrve0j2qZ4i4lmCdhTGpV67YqvqJspq6fE2CJe+632TKrm6DtAUqAnE2GVDS
v3FNFP7ZyDsWlK0by5jwwED98u9P/TW0E+HoDrhPuisFZM3Dnqlph7iN2T8B2A1B
PrcjYcRbBDeaDv524k6EuH9lv44HRAfPiai1iuiWI2FZ8l4U00FKYUH0HuqfzcPe
LapucgngCDZgtF0O173dde3Ob08k1dMzH7+C6duW1xgZEL9xPOuJBAykJhLjd9BN
7efLcUV8CDOIkkCvlXe0Th/K7zNywKH6o3Bq1eq6ZdKtWiXshjfTXJ3LiHJrsaMY
Ugte6bAqdIthkJGkhYM5bS/yKvBmM20SaolB+FkRvvT4Tjv/oUbncYOL49XXVqxa
s9iou8bXi+N4szNPCSXNweLgao/blMQunGHyAXQp1TUBptHEQE/M0VApvTO3ELlx
tEBLMeo+LZPmfucgc8KgA0152rSPopCjejFeM95uwDFxe3qPXriPcxMdZ76iNPzd
DAkZKP2iFAqb81tHV+tskYNrnAWNH569GD+yKGpWlfyGcVDtIMBnPVMVMv4HuCq/
D+Pvw5dBLV7ph+2bn3IS5Ejf9VxJ00AZjBYQ4fPzSPYiTIcM9A/Wec1LHvXRBHW2
qdpf+tdXydpSOPhMLE93W8aH84ox+k9sfc9EbaO+2CXgJX8B22GIkMac1ahBxhtk
62e725F9q3QHW3URvynRQmyrl1aXwFqNrKBfLmHkbI2otUWj0U4LPW7JGJJxdH60
2DHKehwohCn84EmbJqRMTuBy5UlYDHMTgxbM0A7ol3NynNwoDTNiDAY5X2uoNAsa
+rnVEFXFMsq2Yl9OHoWPtHzn1c4Gx/eI+nDfnwNsXAxGSYeoRKM+YL6VqR5I9h9Z
YmcqDi9/JtEHXhrSz7L8mxo0gv9YUs0llevQHLiGwI3iQGGsnIxeTGnMnlbYwaAX
j+paSD/6EuEiSYyx7Qfr+krBfhXO3rw81B5BzGlz/rzDRRf5xdi15Z27f5vMSyqi
S/k1IwBzqGVoaNTYxMIQmCFJgVcUOZihHgzxPgSh61rSpZnBvMSqHBWFhrJ+cDpi
DakLmTRi/9ldhEwc2I05kIaOmtrt41ilwU/7NUW/WEqS7ITrg+1fRHvyo/DhDFwy
HaEfJaub5xRnKr7OcK6LZs7uwm0uKdv0oLGgHRICEKDIFix3yblMFa5xXSyfOqh0
5vpM9YLp/9cT+E8D+KbQEvk0MpBdR8dqoMo1sWS4T2Tc1giCiYbys7tBecjC5pjQ
h95JDg2q2Lw8dgOzO4WQUNZR88TS5/La+LvxTW5n4XVcmkfSwMamkuOI3FbViigW
sb/HgL+rVh67ixZ+4OREeDUB9FPstbkiShSFRxys1jEg3LJd5TUCsZiCw+C7ran7
N7Kj9FOQ5JPCgxNgHPUKpVj1EMM45rsdI7/A7/Xfyx/17Tipt3QtKJ0giERtyibx
R4CNJ/ys8mG/uqazQb8WPaN5jS51OSPDtJeSL4yMslG9C+A7rHTACQPd/Paz56zr
ZG0waFS07a/JfbN3RH1RvE75icfU/xtHz1OL1r8/3RswEJb0Pu/Fnf6L4Wpgl7t5
rpVpJgvN6t6Gcbc5DYwkt46T1oTxIuKhwEoVyeonx2I/MuClHP7CdAOjckk1+/LF
/MQ+d4ItAuQ+P+96oo+Aumb3N9aFYuu6iyI0dLiiXtSvfFz//gQ4hLn4vAQbJ+zO
xx0Td+eTSpSLssSF0vivomD/IMCVWFjBOvgstkq2Z3cckjNUn+PezmN2NdEFLwaW
3flIECO2YrLMXtsVrL+h9WCZeNz9n0KnNF+IINV7aHCY7rH02zonnAz3Ucm8hZUb
73YQ8jK28d9oKuarB41l/LG2Z10K3j1nu/nav22kTL5JMKb1yeFbiiJ9pLt7Hn6X
e4NlzLrtMNZJvCnOTIcZj1kZcm/07IMpD1SnGa8w29nQEyokTKX1mXzsge50fy50
xeYddk78ZgI4k/AJTAhks6OAyE2wJOA0zp1XNeGNnWWRkucYuitx7TLiYBSWmP3u
ApEQOrf1VL/Kcssfp+4NFAHhzJi4ZkgWg0oqJms8dM/dXsCRiVYg9/lrxnvVL4Kh
KvD5B1VLDT0a9S4I4QLeRowlgEbKBcsIVBRylKuEcuI9tTOCvu50BEWMPGWte/+X
3edqzarEiKuvTFKRjWNv/8rk+/+LKJz1a2hOYwuXY981zct/ZTUNf0EQgunBK8NR
uWBhGZxOx5tXEzXb/VZyisCNq7EDhPrOwC5PTUNuFIRDARoH59kfICrjWg8ci7O1
BIFVb13EUVjCAT9Nqq163ssTF5caf1eDozhD6LB1XbLuLAGgs+cpIwv7OyTb6Fpj
1HR9y/eTcXZ4W/F5mvEO7eH96U6PSWgKQYmrpF7P5L7swHGI63qpdRRpDf2latyl
0QGDRaKHFTvjgDyc40mID7OYWohIMMP8TKTcomUBcPmpl5frvykmKxugXwZHHv0L
tEe4Hg605ZUiHZi8+Z4RD+3etbfqUBtA0L/SRys2zUQu3SqyksPUbnL/U1Z8hKCT
rFCRVPQiYaZi1gwG1TsoaApo/+3+ug9SIwiJ4x4G+l9YjEQd5PdBtjD6HaSgmWts
BqRODOo0erbeU49CnqgqKGsgHobai6tovU3MiWz8mxSBir+ATy8haAkdamfmAlB6
pEZzBAZxuK+nw96vZKrNkXd/Ugzp5YgXknVqoYqTdPw3lDo7LTtU60rOPx3qzoGD
F5IeFeBTgmI9J2KszBjEAGJVUoHmRzhUw+n/jv42EuGZwwZ/CO7gO0epNzm1M+CH
IB8FKwlBnazxuAD2UaLf0VUIXdt7g8lPL9G3oE+ZK0akVg+yUh7F8CyktiL4aKlk
liSUJIQxbolShYdWfYqIebFh2MRmz5geyEqOzUxv1+8a2YxG3X1q3XJ/uXUD7Kve
A+Z1pEo1n7IlCb9qsDYzbyBJlt/UIKtEPRqahFwKph+1y2/Q3fDcUdpawAGcDx2M
NZTye8gqttG2lFNJUeBJa+h9AJ8Aq13YYbWiINHQ+lgHb0kBN6Duah6ouElDW/HD
Xnewa/dMB5oWWuiBDTqijTkuuDQ/axmSSn5FPxQP6+4v4MQ2gdazbOXvIfCvBuFM
FYl397IynQeQAxbwzELANBq9NVGLQj7z7ulgMZz2jNLVcO9gLVC0xSmS5k9+zrb6
YD0ERJ4ULswTlqj850uny4i5cfdNz9/tPpPgXvL7jNzw/YJMD63jGYPxZjBhBevX
NBNhfZQOEtHpzLUYUeXOO8xVINBhIyNvNBcQI9jYAmfz+oOBrPqk1U5avUb6sAKh
IUip0BUoolySeBroU9SLvr0Z9JOZmaCaKk292vGV4DCuZ2sBTGL4uNgwIZPkSucq
p0vhhsPDbT1vBeyHwCEfn58OenyesYyJErtuUS4GsrMDpVuXoEhj5OGXPNmXXQg5
DbQ+o6LVK0fo6PR1Z4plTmjGE8J3I2H+5i568T4DIaIjMaaMbRtL36WKnaWOOey8
5xjOw/nRBHkE3iZJnxnlLrOIJw2keM+Mqwb5U2AduDwDE5WsTWzMDS01/JId8stz
7JDSsKTSb64fDSeNei5WLYRH6W8xdywyp0i9eaeq9hWMBdqkGt3HUEXE73hhJgoZ
qalfjg84SlK/lFEr83tCk2Iz2rW7owGm/xNPGnlOVZs1U3OEvwN62vDc77jAkZ8z
AhTWKUYLFzwtISuI+ZbXUmwXi61PAr3LF+rwUgd1GedgLF7Lby5kBMObtRGxGOSN
q4M5vpODvBlDP/kGVv8LTqVFzZGaNM/4KEMToeaVaoqVNQbjMbJkrpIQVzUjoP0D
7AUyJmDi/2tu+iJiZ9q/Cn1Jz1ienTPXEz920hAtpdKzowV4B0ouvSl7rB3L/6jG
729ksCsAuBkqw1H8jN5uvDI45m31EKe/5AVxTg+UQmFBUc3POcGZx8RJ62ZBL+Dn
I7u+GSw8aScvVJ0H7QPTJYrHuwRzkXtOM48A0Tm0WnapXBRIfSbR49Jn6pkLdwyE
KFapVd5ExSXU0lPUmtMSJAgB9K7Gl4j6SD3VWDSWoQ08JUb6BojL/MBWiPTb0BmQ
s05agNcqHZr/phOaVguazHgcW/LtdOHSHuCMEl88nn388+n87qSZgJ4gclkrOzfs
ANJ8ztsnL+xSl8ntcgscCVdJwkuWuJOwupAzwLHRzZHX9WtOgWqNo5VUsdc1eoYm
o6yBCVikz6gIQSEL5BjnuaUxyOvrpELqbVdwM/uU1gUaS1Ct6wVNP7Msca9jxbcM
yBt+zKUVAxswd7T/f3/o/r6QVI4h/wu8nXS3HVm438LFVudcMNLCupTp7hWyvfUl
QqkzO7PUGIF4rMNpeXCE40u0ycMJw/Q+SeWKbVD8GbzKCXxnUACtv1PHrnWaMorK
3xMQ/pkBC0xx7HKRCfEvBdC86crEp+2eGtFQmOy6+iHJ3lJ7ngNNg8bfvZW9+1tJ
H/WBIg+N3xpo3P8cbEnJZIqVWs5i24rZqbBdnzstl6myeuZ6dTm3pBNCqT0Uhas6
bS7MLnqLKrmpK7rFwDogr64eA81mFdb9bsp0bck2cMkTwAJigDwTnkZyDiEb5RoX
4YLgQfX1v+qPqZqs40UyRy6NdR5kTrQjbsNCvvH0KJWe7PB0eA2yYavz0+4Nim3y
81Z89/mjSKfwQMuXUOKYnz6Ug7skFbE4AdJ57eVb09wgHDTObOC9J1W+MreEew29
VIPuGdGhMOQC9K/bV2nkl1WB417aQ0U9qFXj+LgPjh9XU1+bPWfoAgoWPuAc5sBx
Q3rgIvnLRO7OPKn5V0c55mLlk6/hH2eyw3Z4yfFgZn3Nju3l0i4I5FEWCEkYu15g
HZXguJtOLd2lq+Qq/k6DcdjF0awWEKg4WR2VPsVTv8qEttLBa3H87tSFWJA0tq7B
ezYsMF8DYeJeVcRUoTeZVwxXrWNew+asw+kAu9EIJhBqcg6KuJ4rl3oMuopJBzy/
T9KXVqDLkXmoM/X3RFhRYreGgbAVObWThci+6tTrQLToV0Y00iIqdIvz1AgQ4IS8
XOSHjiNy/54/Z/h/xhQ62EwROzIp/JshqCVez2WARV9aR3nKuPirRCa1vL2WEoyW
TBY60VZ4qZCX3WtMooWiyS2gl6esiAo1pbYnjIdVC+Ga1nTzgavtectg3GdYcMad
m5/0a0tGGU1ynBS/49DAFNIE8AMtgn1caDjjgWAifTZmCOoM35kEYrDFVNKGuEjm
1buvxpQxEe5YmEMNcHRq9pSn+/AiMFymW5/25kW7rSwj5Sb6vTOQ25OrV9dUB95z
q7pFx21cKleVf9fL93CcCpU5JBaJgxbVZRzH6haKG00tDJzamQJIuH5pGo8r8Lks
UvjrOzBKKS1/qf4zZNqRGNX2/nF46t5SrZ5TTnxytrxxZUTI3oCzsEJGxmtnXjoT
w7BP7dCbm992EkDHkMUusCKYLC5ibv5gXd8lXrz2FYrXnLh18FABV/gZD20vdBEU
H+ifUCncQ8DZKCEFf0xboTStriM1MTvZlmWeZFS/zrKKra6zbiu4TdzAoJoiW7+6
SXbSPTspMmYIXTbs7t1uWM0zG0KJNKRqv3vzOLCtyHlyfYg96d9A+IOwnDKa+Bd4
/+QXM3oYPR3tNx5tSCGZQ8Oq3w/v74bPjRhmraVqNgXKKr+fNUcjeq6L3QTI3IFU
9QFtlwL9vGzjqevj5Fg+gtwRmB8lbZ0UIM3i1mZNO337vN01o0H+jVuperpqr1Kn
VG0cjs92HaSlmfIdnlgP7z4YBgrkSOeaEpXFiRHf+6HDuV39a0qYDpOVhf1z4p3x
ycygmk61110FNAKrUqOu2Vn9xQGn9EWPylQhOCfPtiElx61hllIoyTcvyqAIW0ja
NqoQtGM2QO5Evx0eztPFTTeVNB/RwF9xISp2fABnz2kR04DK3X2I0JK13qIiVjFL
AeoakrvF0iP6eD+/+bmLi/Ks1TgKPPBw2cnxTH0AN0gaGXJUKL9hhuleRd8jU7MX
6IVIqr9X6qAZe0IeeBu8Ss83GuuSnlB0KsSwRkyjw7Gh40ptftZaaCAHFxxAbpJl
oB7uJbigBW8TqHqy+FWxF3R+83bHbaPsyUyxGLGxF3HDcdL9F7qma13TQ3/cMRLy
tMKUKMvW9pJ162hJ3Tlw+4uPVlpTgtpi6tCGWp9zg30tLCig2pJIRWO11K8c1kjO
zrNbbFzUddjm6rKvTuqvEkdPEYk7nO7/7i/9Q6IrqUKvOd6suOtdqK0KxP2Dxr6s
IqOth8NEzkitlTWJiU6VSvJLXUeMzuxGLxRTln69YFyQIXrRez1a5Rr6LcQIyL63
e125JymKVRVr9wSmc3GkZMtXN7uS45EL/b/oxUKFBTzZ8x6gKwjR3poSGUN5REr4
qB3/cNFOeSCGbDFiNDXB9PYdlSMo/xe54CGsfxzZNLTTetwQWBlSpqrGxtj/4nXf
XevXSj+Aib9MqELdq1spCSGMCqPWnI7NslMnHBvgQ2RNxQvGYV7Uin+kP4eC1xs+
xHW89DCkskY3CyfUmMfEU4r+S142SktKuDkZT/2yfXMlBymjbY9lo3E1b857XK1v
Cl0RohYw6uuo2/PHXb9/75fSg1IZYjgEElSYGv4BiC9q25eNNxrQhqi9Z9MG/WBL
RAyEBRkG0WQ5LN74xXJ5vTf5ayKbCG7mQL7CLisUXq/IiPgwFyF0uYEIUgwEEpOj
Y/4r2zz3IZtV2jrEeuoLImiFBCstvFGJ37z7fdUuZm6S8RRJWCqjM/d3oywY3mPR
cHKZz7KWkbKddmNFIrPZhcLInxPKg2CIltzuCzueY3qckIQT0ZH4YLGTyPtCMM1h
GZlwxelZDLj3gi61j2pYXDATutncrxL4H9U3SXVcaUQ3h0sy2BkppJI5r7iLR9nI
3HMiwY0y3NM9VJ36nOzEnipalQ+JUvJkULxlcchynCfrkNYadHAs2JsvNR9aNrEn
46ZpnQCYoP66keKryCRrw25ILQLRMVuL4qnhJDoKImNcI7g9yAcl0W3Or2IYwme9
oJH06T/aAFIvSu3L2nOOljeLpqJZl7UIn5uO25EiP6gDgz3hJg+GGayLgQuEW04d
C6J10VyQ9C+uVmtWRBd9j509YZaFXae8iMMEZOb74cc4snhKuYj9DIyJZYAAggyW
YfJy7G1Shllg3durzpAegJQcz58J0VmsVMOL4JgeUBmN5PEI5SLj0VhKIAPN1gDk
xgiZf/sFUPqs9Ad0DuztR3Hi0EyhwVIBQWC9s71VJ5wR3fQ3HMQZvlr/NyoWPZNK
I8QCjAjjv6giXuoUEWc5ojewD0b1PKaDtutRcBbAZ5aydNgrgCBnvW3JW8XkVyHH
z49fa13LKZlAC2ztFT62w/G1fDTy3t0SFIZGjmSezQfaHCfdKYbtSmIuYw5FuJFD
UwQjm3FwC3Cl/spSgldNg6j2eCWxHVzAZlcQORtBJ27PemkEcyDsu03HLTQui3b7
+j9ChETxyHzFV198GqOG7Yeb6kjClE3ubgcnkk/ecEcfRj79dao11j/0ypASFgHt
TaIBGleK31BmzlcKjXYRTLlkei8YgfvVyEqDdRzd8c4ueKs4MQJBD961efD8Tzeq
4gB8AOOkwLR4wi+szdlqkcZ1XPPuc6i+hdSYeTThCHgxgj5wd/58ehCd9qGTFSlz
zeyS1iqswPh4u+AIFZkqVkNF2fHAcPj3EIyL2M6R0R0L0RYrGlQdifeFGrBEbsyU
eteJhzmTH5NhiKmBPA2lRqqw5xWnCMDXnjSWe6a/1A0VTm69ABwXVKuUndzn1ARU
E6lUnZf5s9jofNKO6hRO5rXlBsCqvnFf6fqC6BaBKNoQ84NTZSlWmtxF4o4/sMUL
L3BvlKwwKJTd59wJtlcEodqSCbGMBq2p01fRV/CQRqEuLe+EUanPy3uSJU3NbcYX
TOXYRW4e4gEn7/V6XphQXzEj1T+IXH7QTPUlI9ziuephpsMdm2qvi7VVYtao60aj
NKi1kMndNiLHfyFgLmsMbg/i3cye2DeN2AYH7yU6sovrmkKQyYoCiUBRcEKNwsa4
CzuLPzmHzAp5Aof7oHMv/W9B2dgY12zz1Dq90ta4DoMRrw84bXLMS+G/CByagZWc
k5Nj4yd2mv3fOkQ4+MjkGiPtJhSrP2mHF9XTEA3gitJvYaWFGCbTfIP/Sl3A3FSP
jEUiD2FatwihdOUO4SznY4KxuQyzBxoVPEsXJoacgU+ipx+Q67f8JLqR2RYOnzgH
qVGHyVs3JMvq8MCXsS+AsdN79Xb/kLLvGhd0/iHM6tjWnb3eVoBew+KR/oDbtjb6
2vBZKqTgiYqaltHBI01mC6ynB1z/dlMnfo+6NRbWpFzmNgw+pAOz4lRt1YLU6UI6
6NHP0HwnCKef/oGMacxiTHH3CFOxtJjsD6/3n98WqyCc7/gb/eUQan6NflpQG0R0
BY6R9rMix9L8At5NfcmIRkGPcgjFdeHD2esA+OpIyfiqZq0L0XNPRSDxBFXtfn2P
9BASgWCwnJ722YufDRtqyHrLjz5ef9dlAvF/BwkRNvsS3BQYqJqwYihncXo2hmTs
V5MI9L7LPVI7sSImIO7bkB4pqVQzRidBZWfkRH7DNSDPQQyCZURG7PdxHDprrmGo
2lRYsQmV/qevF7Hgg65kKVh39y27i6lK/loD+iUIZhTjYL1xES5+tKhJkt5IuUcm
9fld/+T6DwDdROv22ROx95+GP/ZThX9tEaDb3FUcF+alPwsoCSGxDjoLG12G5dWL
J87g/d0Fes0vAUnsjjdJbPNLgkTnWYT6zK3qfyzXxS3/C7P8fcMmdsK0frOXcM6t
3OrZT0T1uJtjTAzeKKmbSf6kg0wfpwTW6UQMgYpCgxBbSGxY6Ydvtzv7j4SFoR5X
J4GQTkkx3F+r+941FaRzAmVrxrQY9PKC8nR/EoQu1W5SrPXWuK+GCLHCFkCMOs1w
M49PHARix8LKdkJqLQr+bs5To7nMeyPQCgMtHOYANMdDOuPeMUFMtJrVi/K9LC6N
uOz5FkiUTtxfV8+OC/ls0n3xHkU1b4oC4zZ+D+kOQbSVQN4lUZSk+yM0IVOOSNv5
r/gPF+rXZ7ztXOFj735SgtGrj+ITaR4OWd61Dc+jft9VDFDPzB5Vpr9MJ8XJBFqc
M8qzEKgMatvXSgse3XiHfFEOCSLAg7zfIPqv6NaA6mLxTSizX0NrUO4LKTsLk4Rb
o48zDjcYlI9/eWnb6R1tDNLi4Z6UTsbvXC5SRy+RWRvUR3Xgknz8APRabtuG896G
/3HX+7cdVto12nf6JvKw7KNxppIkzyIKDVJyna2jCEgLrEGbX9DGkWAdX1BWX6wo
FGOg1GqXeq8xIqRukn4LVq9ocmZXc2bESafE9De5WneqvuG2JqLknojzYzsd52Rw
h76mu46i1sLu2ReoeTriE2YY23DgX+JVlB+IGUd45+erFzgark3v0dZA9z5YTb2g
MplnSiDBZ81dO6/nrxxONEaXQLv5Duim1iz+KOe0gxeaA8wDA3S8Mi9tQ8qYvRRF
yLCUEQbT9Zo5UMk9sM/s4sPeUd8388NHktGyiqIgVRwJjizWGP9IA5hVBWl/t8KI
nU0fZIzn8g8UGy/tonHWoW6aacpB9ygFWrhp11Pr9j5qzGuOoeuDGeLDIqgMoWCJ
VPPnljECDn4Nk+ZwsPLotvgHiaVWqdLF2eZ9Q50dFYtshrlyeesIf30FhuUrob10
7VNZmZ0SjSYvmf8PU5VZW5gjlxkc5MEFZ2/V11H3/6I9j2bSJ1gLxzPzslSF3Pub
dnWUBzvxG6kWoy++krSGKSFhXQBDHDuImFvYZNwJP4A91Md0DbEQ9ZrMlGQPI8kV
G3nwtDjcGBVREgTbsKNxAe6NcHuJLe5S07PMtN+gSwiY4E35qxX/Slrk/9CYwqUR
Fss8Gr8Q9HJVuACuAVuUX0ReePiKMfRwyi9MXuvLbZ4g+ZLqx8ANoZIF26uRoOEj
vkOThxun475KodYdFFIAFR7XEnQ/NDr/zCQxeYmwmC6/BsXs8Rc+I+xPWrRrLW7F
VG+zzPBQ84AiuNcqT44bsM/fUTv9hs97EcPUqsMiHs9QLGfSYvdHdqNjYfbEyt2H
3ZokiLML3ySAvPpkEEStXqoa2mJp5ZnsidLx3/4Jj4El+IkcwiwdTMB2kcRWFLOx
RD8JuFkpPKzxs53HgRnKbLrttMF5W+yEgNXh+FFCuA1ZUPU65a3C2glnk8pVRfJr
DtJjePvyLgQf9oN7tQihdYIWbfy5UuRo2T/a53/ox44k86qhdsyYnt1uHrAi6ZiW
s5WdZpSG4W2aMVEvxd8K0VqkpFAjnYowcuFHBApuTtNoey+K3Z3Rn7tUFcxIjX+d
K2CtUi6rtcc3PErURUig+sPDf4q3JlT/Dazw5F1D4ayhk/AsPoTEm+oFQ1W+Ul/L
NM4TO5PxF7Mjb0MfkNuVUgePKbkyM4gBn6yUkOamJNNfUIPuuQjq55fxnzu5FFEU
qpT5ApF6KWE7zx+BklYqXLrU7RyotifEX2rCF1oN6VmEeno6MjUBuMc+wHpW8e33
qfXjA3Mhs9H+kk2tnMIGk97KAyMNn6QzzfRaEftqO+yVjwgT/+WfCpU6vGnrNXuE
BUWW7dMkimTw3zrwDV5XoBovLKwFG3opkOI8TKJ1NuLxh6t8b91BbS/y/soOrd4d
UH86p/GQwJ550m7H1zl5knPQxS0HdSQWrUNIzxiY+KPR5ROrZ4XXXQICdoHjZKmy
R1d7o6G6cFyHFGmMbjh0FNEpDEFKhZXqXX94NH3LgmG9kbald5NR43D/IpD5ldwZ
k3fL6vuexYaq+QRiDYt0yNRgPQViq6mjOVGCLqCKrmoRlYEk+jQT5g6VoVo5oioI
A4s9KP3PUSU1Q7I6JhASYQ92/6co0OOivnUIO229v/4pomLUPFIC3C1GK7EGTKrc
QP4Dc8qZck0MU/e+yaVTOQHzRvGdYNJz/8AyWtb9DK5voWVA6p5lGnfqHHeS6VRY
77J/Yu5C+PhFj7/0cpnTIxoL1xYLr21Co/Fls5BiTHkohH5PF/+1rv+nw+ad2LNp
0fQSWtmTTwf+2/Q+5u/ux84P/jpQci3gzoTCcddcHfrQHKioRmdX21ONOBfBaEvB
AHyNt2Vf294yNdsFtiBR1DLmumg55UIrEPmkg0Aq5XXQEtztr4mKsdJlw/B3Fwfi
SwJ2mj+hnZeJIzY8JKmkIImy+eIGbd382eMN/UaZaPzzpgUhtmg1wsSKwEH74Zv6
5Hv/FoxHPVIYZJgpF65ORGpS4ZZc46PBbPdxsiYUGrlinjdE6V1kfQp1sYkZRVmp
pF1zAjUdg0n+kaOjHBCpw6WQTYYZ125KNTGOb7ZFc7xA4B01MO7E62euwbrugXgQ
HHRaud+jJUkzHnB7DvpG7lX/P3HR21VktaRv1l1rKpVu2zsPAe/MaJBYh7i1MofA
vv2aCxkLNZlWDxjLxqB1XFu2LJdEttJtSlIHbgnc0/uerlixGt5az4GcC1lPdTuQ
u8MCIkI4iaOZK7rKc1oUymcyFmniUtGCwrc0oYMNw6MZfze8fRk9io1/H1sdADEv
jWAtzRQfKdNLPZ7b/xyLaGvBbQzZfbdvd+rW8T9GpxRRPCipaKx6YWOJiITNyv97
8c8zuIOtUuOB4EqvvfnOKyIc3oEJTJIQEan68VkxEVZ2wB7bJ6DymmfCHw1F+e+Y
C3dP30p0Fb81hwCaXhCgWZvUUp3TJvr8JVxvT65no7qGxUntiJgw6BXSK1miV95o
UFNq0pEYxtt3Fi8rn3cWnx6115m37sZg2WNBudChV3zxP126GQnlzm2BgNf1uwBU
wUUJwIWf7JvrY1bDMAZH+nfo7DM01ricYQLuZC34Dh6mbPwfIMH9Xv+i/xC4PXJV
KrnemAG+L1vXVOVxUJcGlhhCAKO42HfpnHXTjgtotG4HEOqRCtvNK2lsfvB8tubO
LLqudCCk0bnQzi3ylSfQcWQk80LOj4i62vWH6EWDStqTFsUm8Iqwxubi6x7/v0wu
dyRGL8+ywe7t8V9v3TuErwah8JmziyztaDjLpsazMXa3tmBqkNxNN0a60w37IJxi
XtpUvNak4uqshJLBuRpAuDxHg6KF760gHATWpFX98k7/5+ZiYPg8vd1aG92h09bW
efLSCs9/YhUqbqVZ+ytfyZwmCz389vsOmHsHl1WuJpxMeX9lAA5/fpnDnP5+0OaZ
1ntY0uH1hFaPeLywyWHhbevZKRWHbnHxixFLUYionVg//mQqJfQvrkJ+3qAfc3Va
GoDCE+iD5AXB/odmguZaohdJQgIWOWEYfZTt/fSvSGYt2CmM1040GyHAr5wiWz2R
0o5i+12v4jFJPRbdW8yjy+RDv4bnuRBlN8bp/Apr9hoLYnEDciDLHNY7DtuYY980
WrY6DFesA8HOmksgKFoTp13CDc+oZmZMXTqY5ujLsQ++UtZ6TY7WIIIM4MSMfEnw
XBJVnrHwj6wu2xa+w1lQvy2pSRa4o01MvrvisI1LO7R8C98QQ6Wsz1V3sFruhxbL
UOwyDxrtAZ12Q+CCbdRrCxinrok7LVkzo44fsf+J2EousD84nlR+C+PZTC8HY2+n
BsNeoGSF8kmLH5pwN1PNgyWTkgPyoMehNjkGH8nk/YCTSi/pGLD+cf6OMYM86fKo
GvUw+npVRN0z4WC91sjSrLPPRqsoUrSoUFlzCgj4CNnuUN67eTwXmrs4rqr7UJlm
kx0D5mvS0Ok/xw2zuWeDAltagewyReeGx0E2Toi5Aa6mGZ40EcQqzh/6IqEOxvXl
x7myu0NuSQ1mRvLBVt6cedxfkmTzqqQu9A0n6UuPzJMsh9Ydbk89Og88EfKFQjRy
BrFjvMEdDunDR2XmrfyuOhmZ3a1rrhqbBpz40Nw8oFp4BbQAGHhHeMvMp0QDMxVK
I6eLl5oot+9mUyg7D5zbSyI1KwQ5gI66eS1q4Ve9savv3qO2gM8NSZ3lkRLfjBCB
wy4eqrpygzE2E9XfmaI5Ct0Uvsbha5TAcTxi1r6qlxfwUPFgzH2fXuCsD3mVVWdf
JK8sO9OVmrj2Oaj78HqAHKpuaMorEZAA/VaUjTjmNdOA806qPTs2lVQnJdrjglrt
srqxOXuoORMtetUhRrt68Y1R3PdoiQP1if3hi4TOJN0izQ09ta7fFLSSrw95gOQA
/0k1Vj8eUPly59OkXlphNx7IEdkgv5barWT4jkgfgL75jiPnTfVISBamZTwJWDDB
aYI/4OEofF5WDJXbJmBSGFex4j9uVkCpqvNexSXNjWJynWvq81fdcEAmdPjZzF5s
/AMos+bjre3ONDGCd2O01YuYqkRGA4MdYTGGXkjhcgxnvBWyDNPVdWc9U21+cqHy
SVDxxmhjpzgOvHnntGK3teLPBYLcm3JdBWWFiRaVOc6UwOgd4njfL64Wn76R+0jt
ZiK4XClxaq0MSB1pInki338DkqJZhn1nUsxkxbP/9Jn5syrkH4hPdmNT4l7Wm1FD
dAUN/23QGBtsIEj/0OmeM/ke0OneB6mjzHOjvuojfXsdxxK8qbeHVDWOLi3WkhpR
HHjj9IYmiFz+jaCYGAtrI6MK8MuYgMMvQqfizZI1MAmGv4+0e4pzV0KIn2Ehhp6f
DMt8umr7rfgFEtXyOy6GgtfqqO9wHl9zwsVaQiFiliEQAnnhXE22KgJoVsH84Dnp
BAfxVK+15b8N+h0i2P+8hfI1UOMW1Mqd9k51NOLiHWuM1pTVefQ33aqc/Ul9wSE7
3R0Plmp2AcnJbsYHMC8y2W1wRrckiXU+8lTrHDvj0N1F62X4LI+m0T7iAsvglWJ9
SpcXZ7Tf1dDjseguyXuP/poSICBB4U7+I4slQUhADhfmGdf644ADUQ4pYTS6IZf2
k96hxkiPczljhZI2KvnLs0fSp+wKzViyouYSkQOOqT4OvFGGclzUoMhEchDGtMpm
u61LCBigyw0x7PAIgJGRkztsF0hYfcdECUFNXebsIpS2U0THc4PR9RBz7PJGGuI9
F1otyA3+k92QOZhr4qncycZhvWxx6RDgF4qfmU9NTEyIW7piSyGNlhUd3+im283D
0E1T90Ax44GDQvUz0p5M4RxzxxWKVPGeh88L7mC1ttnsh7F1UlwWO/V8x9IXQNTv
yWlwt4uEgb3+UKTr6RcbSpa3wREwxyHgUPibnN16kpWEs1bFj4xBfFrxLSDuZYEj
P5Drx/Gi/9nEN3Qs0NreqYvSBIR4NxPra605rSIyqb14jiXvuX8FQNAHCD4YEdU0
uYJ6p3gUic5gDiH17JTXoY2Iox+oklrGcnHUv+4z6+h3pgcvpU6s3AkfLTMVn5aH
8EC1hK3syzYyBShRmNqR8nbxt5q029+JGGjmAsFi9gX2UR7ZwVBv22cQVuCcFkKh
sfaqE2iGVjkNXOfDywW881mZ8LHSSKBshFWYYZIQNMYodmsdFkGYDKHbMwPpvjMA
am0JhNM8DJC2SmBTn1e1MMjRCkEFii0ADGnaTl9khQue7cY/5wWCuzgTgh4Dlnff
thQSJGu9bi5iRCeOCLGEAhu+N9ER8THrxaCet5fqH1c18T6YX+ukE7rVb3zAeO0l
DOasdLAA16ZSfrehBZGtREqgV4gG/OkRzwOIcIvCLZhzo3ICTYDJdBnK2NSJzlF2
N7kEg+T/LnTf4ClMdmCCm6iO2coZpzqWz70Akv1ACJ7T9IcFOXqInrjZ/hD3r6bd
QCJpWlG1lDLNke5diVqmSfYHfFYJF79QTswQSmrdsD5ko4htr4eIuqIzcahcsTA6
nAm0rtNiyheHzx+7GBQ5+iuOHfWr7cdUIjVuQXeNKPAG/lnsLQODeYxALuLfedLQ
WtN8d396tc9GhXEwvomY4TNVYu7DmAuOGOI0+9WvM8Df6a1JpQS2BaK5VjTFl06S
9U1tm0VFmhtzwZH2W6rpLAZx7bekqjqWr4TdJwfZXsA3mTHThld0qnHLCinJoNcp
SfvfTWzU9YFGDSYwVEwvwN1knrH2TK33BHtW7xu7gtF4Nwry9lU0w5GnI+t14Ltw
KmoLz213qWXVJSkmTO3M5VbOkXwk690WfARbaZGBYgYJViw/wxFm5NUG5G7ELSk3
7qE39wWZQ64/jqnz7eeLpP5zcD9Gv45khCaCgoyrNvLwtK4qbjOm0ZSyeALP6hCp
HWatodSJP/S822EpK1PUY2ZsFUXl/qRmw3OC4TJTPB2GatYcN7WErmdgsJSsI8ri
/WKGtyG5u8TFdY/OKxr9/+xXfTRok04nkDZOerF5YZApvIROT/VuNbMWp2o3r4ff
yoAOJ2J8CMsHwhk3WqSQsQS+7FYixhQ/OkzOLY5CGOwmqYSwcc1b80QUiFEyqFCm
17ZrWDZn25awMSpi/brVi3DDbSqb5yqPQdJW+GAu+x5DM0P15+I1KBgOjto6EpQs
11ACJzWiQsWwlC+nOzgTJAwzpPgIG1swYqHAbriuixSQPMLsxAdrlHpUPF8va84o
+reg9AY9QkTELmu+vK1+9uhNgzIDAqI8CZ5dQhZzWU/gr7du3feC5B01bAEeCUni
XUM+0ODuROYxbgCOiLf9f506LYo7SDgwqO4cB6mjOeJpvzPpycNZfrkMgS9P6mvb
OkbDEbct1ecoXxGeKSqApmCfNxWZkcEOqlqrjqmgqUOds8ASMIzF/s4aMtY8mFaT
hMcmMrNs0nVLs4Nbo5fYc+SBJYuRU1LeRH4Xe5Nj9FeXslIbMzAULm8erIZ7tVa2
IyPjfe3+BLIwefUbF2OINwuTWGKmyp/ZTroBuOUnoJr3lnd/G+uGTh2Xjwl9jNt4
xOJA7Jrc3fSCnmpemjvkViax8e9t88+nf9GSRvNQ+F/wlETZOOA43BJonq9NsiTY
kEqxLLXD9w6K2lvebsYJKMrk5L7l6ux4z+dlE5xFdTS6EtlBk+pKq0j4v+Z8bxu3
18tX3PhB3KU+reCE37yEIqu/GQJ3pFkrSaZ6nDuIO62C8nM3WTLyfh2chqI0zI1+
f/cwncLsFenDdJLVmOFaL3G5OhWKmXTHt7zeycNlcv4fmBlRq5xA67OK+OAPW79I
a37lDVxujmhMQgrLJakdLxtJEFOLy2lnEpFoVzOqaOKaTq6/kl2Bs4UCGPFdwGvE
8LqR6cIZuYjMRQKvXE6lnu5y+wNxtwh8zg52zAd9PZTeMRC9Fk/Zpu69eQuY6MUF
MIy3cy46B4AWBhA4JSltr+6nE+KWolfOsxgevk6QvnnBy/tQmyirZvuydS/9slK7
5U3xbdLEfBsnQS6PI/7U9SWlw1htTjr//anhNCW0WwOfy6w7X2SKiu0hZuCbYx81
fuEam7LJjbGKoMUY9p79I49moiz64Qy3s6l3LUOp7jFvCRWxWJV4T8Vp8PeXw2l2
7fBsw87O3a2jBU5sy1kjFixbWBf4xKSZqltdOns53M5WL1VZpnr7f8Csi5WH6x5v
EIAesBhaxNrcBoURDNffypP6kXkfk4NtW52O3XuRgU+GG8lZZhqZxXbYKuiXfI65
aexe8P+yXQ0tJ2nvREEosJaBkhjpt7Z1HIvQ/vvUAe3QweWDulahW6HFN39vOK1e
+f7WohOJNoz/+5nFzHNKwoAMTYkvP0UdjtT4lnNhBRKw0lW8MgWIwB5Ma9N1DowR
pqCaVLF+NEsSB/0czQpbeyvIw245bPUrW+S04V10DI5RQ29yDlFZzBpIIEvHewon
7urNk7AXaVIMDAMnEfm2YSFsCruvdqY1QuIj8hZCcO8yQUwPgulOZ9xfZW5qFH94
yqE+arj546s9/kZ24fmggmMRs9q8WVHe1CTQDwWB+r/XG5KqUj4R2RQMEUNKEszZ
QpJStIp9fzmpTchndptqenuPRA54d7cl96ZYJtZ1zIcqDI+ww35Dz2JwfQgiXbDR
3Ny4+ZgtRfbd3KwFL7dcjMtiVwsGU99sD6GoAgK1zWTfM/HKJ+eSIiflQpU+23/O
Ib0GDmz3P9f9MOjVJT8XDj2MVnyBMkBVPBDD75d+x33JKO+Gl1pXkPVXKy7PKuVB
YkWnaFr5xwHM6y7diiGg1ir2CS+2tnms/k4346i8OS6Pb5eAEsjvAFygCdJ5m2DA
Bi/ElPV0KikV1+PFoqQVHlT329D1uuSTJZsDOUiieC2w+r/k3BrDorQvKXjgKYds
tnHW0/m9M3ettptmmXP83qz5J9ay3whgUFxnfJeZ1B0k3+amGBGWOw9hqPXo6owp
sPKwMUnPuuQAQ0p8YPEEerwEsWkoUG6sxcjO2zWd3xYOtCG62F6oHpio2hfk1W0n
RsvzOrdNRb68KU29L1FOqECriR02Qh/RMLVXoFtsK1cZD0YZkSHvB+Ut+GyKk77+
LnlSM/GdhgEQA9iJ6thN9pmqEYNq3/hOA5gZiNd0nH/sB4Q4qVEgB1CNy8g4c46H
fO2RSGM4fZYyE7L7Zev6HUxyfIKAuQyxzu1GjzrWAmIvxuVQo7Md5L4+6J4JIW5+
z4PHV2l2opfpODa/k7jao2iU+gRdWX1yiP2X9M3hRvDe5Tzl+SikeM3g0U3oBJt9
SjrQhjpZ6rcgW2JzknBjFHJRsrbZZEiHNbLaHjcuWgR3eVy/nZ+DoePwsqZCit7q
uzAXTTgI+oSuy9tgeJ7AYiBl8qLQDRKP0UBv5BrsCOXKhw0icyv8wYnUTqbNQMgE
nxMxiAtRT/0t9Qij/UujR6v8gtMFSIh3NqoA5eyRY9d5JD3S14FNb3kIXYCewpDe
+CXABwS1e+qVjyuMBjkLxhxKjkND1kjoemJ7yT5PdRcaKr3X1rhRlqqP+hN90vDt
o4o6bnMwnQz8O8swa3XJkGbramTqffLXv3M9nxhgdek1bth6AjtrseNFSm4m7gv+
CXCeVDBaS0XM8PhSc8rCiqY3ARpqDHgGvD/guojm3qU4ng10YHUOdiyAM2Bhs1pA
FQzClGqoikdVAhx136V8i3Fxqm8yMig6uKuOjZrpWflJHK0E54iMYUy/jBqliuAH
kMwbb8SLV/1rSTS/awIL6F/vsivpNSCU0Qzj04pxDFEizmXnZCvJ1zl2exX/Gd0i
4jGEcqODh+3VdQz766cCTDPjWYtYMMQLS+S6VQQ1G2vOYzOidpjeuaIUTbvRznmP
a36tOPyh09Pii3LqfIlGYA1s2mnNpdbr41IHl1nR5vqMNd7v1EINipEuUI5MoruV
CoUFEZwRsEhWW5AC0Y2rtIYZnX+KrJOW/4Koym0Mf4fF+XgWH9RJ50b7gejiJzIM
8pn7kY2VYmqHlHX1Q2Fz62WxKXADdkTIo2UTs5+rWiJTbQbLXa2r9+388YPYj/qx
E8Ald/HYMlPhpVEXqnenSWbybx4r3EQLVx+z2DF/7yk6+iqZJX22bGjuJVTfzqU0
raMwIgN2y0AmqcieJYiM5NrIXvyyfD2lgBP0lsuWCm7fc0y+gEPuxm4WVhL+qvgX
+oN8qXhlu/gXmLcKpW+Z8SBLpzQfOe4mkf25JUONTPxOvu8E/rzHU9XCQPoX9aN5
OChZ7wp9tZFZIzsZmVj9bu4Mcn8vo4uln9+ZMcuzzfXXGIzcwZADj+YiixIxGZON
sXd921w4cOxsusgxOUllvcrknGR0QwqnLHBLyseIaPdwS0Jw+g41ildLCkUiKEKA
2SdouLlhnz5O6kQKA6rlQR9tY0OHfH7CrHJpZYGaFJ7pQ+ChFVIoPJbRpitm10vI
IkQOMTrWs6qsUQwdLIC6SXlP1OV5tLFGa2b4drslDxkFeqs5K5DbKXnu+CNQks8v
djNCX/4tPjJ7/bjsNDGeXoI8WDgMFfT5uEIISJX83C8uYOeacDQy2Qfc5wpS5NXU
F2I3/7WRZWDyDGaO97w9POoN9O45j0CNhFNnLZ49nhR9ABnLomjrm2Nf4OE6edsj
PTVY49Op3Ty0vDESBZKMS56trjwj2EJ+aTfLBcVYdzFlIhsWvOzES9iWQaZW/chV
K1AokUmTLE6AX19yOaY0BMIEGZMlie6fh9ODkCA5wOBmPNjIbNMQv6Ie5f0MlptD
s5awKGohhrlGMci3nu55C50Zdl9biXh0Gwk/jpjtyr9156EmeBwxpQQwREhV11Kf
bJ8nrqc2qWtcP3OInIEsOJLupqOciQPaCgr7kZiVLtgTwxez/GUy5Jhg12z1G9UB
Z6OZG+cVmc9+oOlCpyKimNfX3vhsrOMesxhQcYjYJWr6ku4ZEXyYZb5+OwunV03x
NlRwrTKZm3wBr6DsFgqUxpBNjAFkE9zSBR1IVRO2aHS3+y7x5h3Pa+C4vA6ynDJS
ibPK7hXb5w6MNyYdwZU9FKheNLm8zD+Tz/TATsTbD0gaGnD2T0Uk4LlQcxmmZCyv
s4Aeg4WFh2nJT/K+DM/GlKIVw1VPJpoxpp+ZXzuPcv8cQG2xBR6UFL6Xa6c3LBq2
mqCAPWS/TvOVpAV6MyUuIYxQsg+Is9kEZz22n9YAbc801W/G7ebq/tbBl6dzFs6A
tJX2nDuqGDe1Jh3LKDXNbH6890guVIl8H6MMMpOFU1qzegy0NnfOvsqpGWrEo9hR
1Guc8g0ihbMMsvGhk0ofKzyl86l/BIv+IlquLCMJbCgzIAsS8ch8q2/Cp/5cFMUM
MeEH9at06JOKqMNMsoE7/NSB3NZyXPuO3YqRpr00HRw7pA9NhDPUjQ+dAHAw5D8v
85n3e4HNIVR4wH+sCEII+7FTaT0ipV/66FY85ibFCxjqMveN5UJCZV1UhJacFmVy
02bMJTPPxjsAiGX50J+BDzJRSSOaHbcsiw5PDVHtcVcFXr6PTE8g4tLXrCcSPhEn
7+RlZTdsh/ShfAadp27LpELGVqHaLHxsdhGh2xd7qbKVO3t1o/YdkyGkwABnTYOX
esHeMyCRdfsCuAfY7KcNbjn83JYsTpdGBvoZg+riBRGkeUqumDSLsVVOSuWFVGza
vcQPbZvZIU4myNXjUKr6lkmiV+nagrI6dyruz/rCW8CIt1FOzEQa0t5nfxo+bpz6
raAbNJlrcsSAD33dNko+/3PpC/FhHIeL1U8MCxmrl+EuXy9JTVG/IPSq7l7rV1v6
BvhekaeTlsIo3zqDpUSHRQLk2y6dK7pYva/4WE9kQpyeDz+svPDpxYsD6hGX2sCV
1H9Geiz+yiQ2Z7ECunF5wyXbGBBwfP8vAwbe6DAlF5+CW6fyPQLIZihofTcHmPvd
wfblLH9INAUw1YWB1RkoW3IE4mebeIfNflnqMg9McT1xjAoabhr6s6Ertjy0gVVl
h7t4lMEt4MZZU0A+fJMxYP12tcur1vy58DgmBjKJuzrVaFovRvdPPE+XFCgl4KeG
jTfgl9zFbQw5KVc5fVW7yVhmhbvJ9Yvu2g5mYzCG/0d1jt52y4ff4l+LkOjUevW9
Wgjry9KDisrkf87lSm9A8GFweE5ldwh74ZtAZJXKlOgUJMmjy87FOQFYbunu08fb
vKJOguV2ansivSOknAaIzRq5yui4oGF4Zxaq67h7qFfnkm8RgIn34bVNm1mapu90
yOUn65rCvhsgvdGZFyuJZ51TOZikzOeE6nOKjAhoClvbecYtiuDYP2cURdAyPEmF
bYNm5b5380JZiSCy/vUQMVjrRum+F1VkQs90hY4A+6tydu8DRD5+4KjJjpAPQJrM
qNl4T5my62ZzvvR5R+rixUoICvbpZy1asKaxRz/NAM4UFm4b8xuYk8k36ZKwQ292
hXFocoa9IDGHVrevSS5zYZTf888ljM9estL6eykSmLuzXohk9xj1YT2zADSgVq+q
vI3BC0GRxy82Mkl4AFlQr2CVq3JoGI4Bxd1o00lCwBKv7uAGbVCZ/yd4alNu19pO
OuXVM43mp4EFZL+o2W3Y//EJEQTF+QEv1aptZc4QU5XPtr9Zr6F2UfxptFkIRd8J
aTkb1k4SzioOlK0YEGjeQwbHrPODylaLEsy8Q0P+voMqX4nJExlU0xFyegikgZF6
Cf4/xfz0+DPhUOBr5jw1uDiL2EiXHJ25Kdaezm6FpF4+BAF8oNvUVvFsC790aSgK
ekLrYewWv6G18RLGI4VZrcDCBIrV/0exxS9mkSh5MjMzKwJpUL+bwxEtq1l43Tos
GroVj8J7Y/S5Hl0uhTK5u4+phaR3cwEZpIC9hP9F9x2m9SYFaPfZsMIRa/329owm
j/TrZcCHzPP/FCThSPmXmNFqSlMgflXcevpdQWgXc9deG67P3fQw/fzlrBt7k3rg
rpJ2vJ0ROF4Hag2J/HeZKtO4eXlg68KQoW6p8YfJMN0Ssjmz6uXlUJpr9iD5jb5Y
C5z8DTbET9Fp6uz6+S2Px7tIHnaefaVIiszbnrAO1N69RteqbdPUTdxxnaqKTFC5
yXG+JWDlFi95H4jr+IcojxafA7sNOj+MZ2CXylRD4tbZT2Uxny9trl8AZAAQXCNQ
mmhNKNg2DoM/Y3jtqJLh1Dc/l26byCvYTYEiuN1V23KjsfyvURq74nl7jEH0Qpe+
bJ9TMSw2JUmnfY4NUY5dd72gdlRMrSF8fb8EESOzc9sRv8jSwcauiBHFQvxECahw
MkbQCG5mPHHMJ8rt75QqMw90tBWQEElr4r3Bw0v5OOPr7Lv74kLCXJ8GxcfylKPX
eSaEJpy0yLYeREY5SyvXoS/icBZg8uGmQ0maKNl7WJrOZEFkVCe98MmGvEJssYYt
n0O+Fgs2+GNwzjm6QXClDlXO+U9V8KRR9nWr5wj2CzxpVYDnEOnzEdN4jkGhoqeI
FpBlwR3adqovc3u79TVKhTnYRSm6QYyNR6SyGgjn9LXWv7SEMPa9saPJ6EuE5gcN
vcnTHZCLPDNnx3LAp7SPK0n0tTAEL0DZJlcYD+dk6plodV5312tTo9MkEiBgrXwn
L0KN/KFKFx/BWe4+WUvtv/kDU9Y04t2Cq5srpMZBS4w5BooIjBCv+PZwexhn4Fjj
P8ceVv1vOPmxVVvrdB0aIP7P/akaOQaU++A4TGteQWc2pSFqGjVeDwjPg5+wXrBm
d0BsM2UaUK2m2WztrtB/kHweLzVxbwQYEWsZlNLgxhvDf/mYAJ1x7yHBSwp7qCwo
qmlz3NuGdZ9LmTpfgteioGX8oIx4nqTRNZ0j2GdqYYDGlAXpiLk0ujwW45XOjeiL
EEKqOK4vTGGkO0kuSo0cNSKY6Uwc5gd6F4sNivL38sLkBxkfh2DJyt5FkOpLuSbD
bEcpdscVnhacKmL1E+7RT7OfuQbCmPYmjhk55S1KS/fjhku1rbLuLon8rago4HCl
CK3+AnhQhA36tzb0rcHs1zSoAzOY7Yd5LYeNxgVgHJqEqhB1xvM8yzYWex3dU1EF
k+QHZIBbyw/bu+c0QxAqjy5B/tZR+rLj4civTF7n/HAYLinMPOpy5XbOb16MnrkG
pNZnPD2Uc3EAfB86E+9D2qUAbSzxoZMtT1BD/wZ76LFRaht2k/YKV7AGE7IPjtOO
wrdpS3tp4vlYDCIbW5qAd9L0Ud2J3g5yTitFjabGNLaSR0hkDzbUhS8gZwmXnR3r
0Xf+zsHzr++XUQg5b0CSPVxgU0gyungq1E8tB5gUiOT4QffOEkM5cK8XqxIj4nEe
yNzod/K6/T1qaouv+kFBhyHQ8gozNTwjwRKQZKgyAu+sPNm/97tMqmFUSCmsiDDw
mZ+3XSnB9/abi+2WI1yAWsoreRgp/aLqbfSSUaL5qApb/MUy5xSIaXhvWHMCJFe0
Pb7F+X+CT5ZGQM4493zF1ff7tlwjJehGU9wLsf/8LpGIgY5V1jMlLtqIbfWGoUJ2
J3xvOt+p54Y6Zp4ohTyzFyTmp/yBP0CRjtbKPFI9wEmK7xfyh/8oqqbeMqlkPjaB
vA2rNm7IV1b2NfmVnoqrw4g8hC2Be8Vdi2v4PSvHt6q0PyLaAnmdfYQdWNyKdUGM
/Cy83LxZDIeRruW49u32+RjHyGBs07hL0cHQCMLvKx7rVQQbhVVSBdMNZhcRgaJW
8o4yZPCQmSb/FZ8BBYz0JQ6XsZuIlqhC+2Us1daozxQ7dzC4HabatZumtkz/se+2
3213G0DCoxSMuDQAgzpDqsIgN+8/yNIjDsZ2442r7yOGXrTkVYRYR9g99IZJdBfk
8bqTrzx1AK86AG0mKdvpyFct6nVkPxLbpsFAjV/AkCz4kq23FiZe7l0xvbzOjFey
KbuwHgxiU4pVXfu4G6TNAr1mPzQJfC/LvqGA6L0G575qnjgXCCO0or/IVINTnY9z
WsH9Xhohv5I9ry9hlp9CPYXBWx7av71wEy4aUvbCGBNkuL0pO1fZGsro9ch5EsZB
knFFCUXJ67LovioCvMZNkzg/VTYVGrL0aMrACLCHSW5NG7YQInOReUKivtGgob1s
lyDwBVDcgdJO11G8GyxJ9k1gUy/0bIgEIXI5so4KwQKAgD/QcxawVyYrG9Wwy7t7
NIt68YWDfYY1jOXSekn6HuNjc87Ucx6y1v2tKuIGycsFbXz5dL5DYMLkE2mHOIBs
Rcxz1Fa6jRrmS0LHXsfkDULWZ8NR0C5aYoB9UkkcqRzIvNqTyr4876kXVyVj4hWH
yO0VIQpBhQMC64YwH95uZ9y2gFzssEK3h1lt4r0+/8rhny/6PmCvKYKLO/hDkjvo
/V3ExVEx59PAjKvP5OVRmnk6d3i2pKpj7yS1C6ZIKTS+se8RTjEyG2HznVFQP/jP
jTEmPMOMMwljkfCXP3eYxB/r9zXkNq/hT4IkYuIGpp3MV5SQkyxA78TwNX8hc+3h
xVEHPqR7TaMA8pRlzNqYuw/k+W+D5LTVsckeWrgdEhU59dobBZZQ5qXNS33IICrM
5agNCx4Tk9CuR7QexxVozx+GeMc7n3NG9M/aCA96/D3GBa+RV2RhzlklgszWPWJj
LAxVc07xTjijj8IMcuXRtXXEV1BmSX3PoXjohW7+pQ66xpkXC2sFoLMjzL80HZXD
9Es3a0pdLDxVYr+op1thEeJp6W3ma+DukHqUiyApMAHJD3qo2yoOF+3BHApWpdu+
ywi5ArwAtlhq8ju0NA9sonFFpgh4+BE5L2Xs6bS+O+4UATW8edYgoWU64q6Axsbe
tJUytpRB13rCXWS6sTcRd2vBZMTIfUh9AbJPOQoiEYM+K70jbrLh3GPpv/v/B9xR
5zDVUN0t7zO56YaScpuYtFtMgKaG3azn+t6qkYbuuN6RahuBEC62SXs++3CXiQl/
sAv2V6GU8ltZj7FH9BB0/DEespKfROqhQm9uONAYpoEAZ0bfcOzfURYberxBwfGE
eOllJQFq5By2I9iO2gzdvLWvNMpsWQVp9FVl+bZPPa13V8vTYfxLV2NGEOTECywa
SGfQFciQXORI8laFGNBGYbV5/oMs+wbdGGn+FUN+xAVujZiD3bkz8Sf54vBWBsHE
X8orKB1n+Mf3L+XUT4JFlq/+DkuqMagKb8qsF1zg5yb/2haqhWfpSpMB3WyaLp8M
GuXmqoeTVurtdN0yb7h7p74G7XaFHbuyp9tI7HuOMvF7FTjchQZX78A14pRxS9rU
eOc5T8kcf06Yw0Gh0h6j5izTX1452sYHPzSUpSf5GnSR+K0Sm3wV6cEemXgHq27x
pamCOATwrNWVCzQ4+WTUCxFiQM2Zel7aoH+Mo8X5LnTfGCR2NW1b8F1K/q5tXTpp
He8nVXEBgggD0tgovD7ilxGSQSglZodAC/Rg6ky/cfE2hA2fV7Ce/I08RL5z0Z9d
7VEcrQdkdxTcAH1kjMCPdacQCsP2OaVn9bGzVf1ue6sN/qD1csBnR2Tm5Ryr6ocI
BKN4H4sg/op7QhxIlnjn3nRyY1ihW4IGSgnsgwQJYH9S8qNOmFqBxraKUrmVv9jl
56ta5MaEVF+xFzXeTKYL6o8EBfUJBbEhjGvesUtDPAvpjHfzMXTy7uMI6UMtOcQ+
64cjASG14U+tR6ZTnB8WEezVBcfO5EomGICz3zceK111jtRUtNAIHYQwYiWi48ZM
f+GhVy9sTUfnHu6HwX1mj8Wso/CdSX4l8iCWx9c2SgCoyz7B7RybFEd0oMAGCBcX
S91SCS9KKGKhFNS4a68mDG9GHFwIMvoxsJuWe8jXHvI/di92QdBqoXUz+eoZmx5a
IcFz9w0vc9QKG7b9kY54jPzC1D4VAKDD/Oyizpto1Egu0GW8hNOdSqPmXu9mmXN8
TwFacekwjDd3lZFfP24SnYyI5fQ5sIXNc6dCKgk9LJW/ulorn/7CEJB7UvVFaYCb
t5XljNTaox6BQqOSf3BqNAtL4KFsJxYT3fVik2y/Sm982yh/9OTI1682pZVpBAp7
lpzuWC7cH70QpxpUqBazmD4nstDmMDexlpO/br8WII2jOpwvBEcFyx07GJo5bK5W
OSC8DO1V29sjYoA0HSJIC+ED9A2jP5PLrPsyBloq0zkEGBOyS/Y2Ki5C82lHItSp
mKfAOTsAsm18KklpYSishgTU2W7QUjwI/rm9RBQUySXfr5zFV4nH0R6k43d4IdmJ
IT2mhwN4WNQGnrow7rbegjT0fm9onmhG5o5cFVFrPnI0j237qaWQBG1A9Jz1xg8j
cBhe90PeslRCtBB9ZliZmKK1ZKgjiuMBi1aVJgo7xkcVU92ePoE89VlRKFYMVWzH
Wb3Aa7jm3Ox6zb8A0IrtGgOB8tGcrBTMwMHyyvALzsxkPY4xwBxxJlawyrG6sotO
IboSpHTHBABe+Q397HMBTkPGf6IzleejmXGcKOD+GjfyUPleKZqnLYjRBzKgu6Pg
R3ZCHNmkLSBDJtCCEf8yuwu7uwTN1aK7SmRyxv2faCrsprkix7QgD6AGfptWjRAm
C6zA0d+zq6WTLL0nwAA7/B3ilGIyRYgiWQJT1kCdrEndfQmmtF8XIksfFsDmn04E
i/bRCw10TK3RuGs62LYOFyh9YzVPp2BqNtK/1fQGjcRYtEM+5RfHUeVmZ+EKx2h2
7FSVojOdZ+sCxiopG8+t6VqbFjTQVYy9eFeaqIutWNKotBUoFMNLVsSKngzPsSfL
rin+Z0splwA0HTEw8Zo5kCo/zWMQdeK3EAgM9WSA54CX9mDayUdxvH6a/0w3ecPq
1PzRaYEaFQrCyDOGR4eYh0nkkj6nBMYhVzujypFrxOqNsZHqvbiodiTsqGoXGHC0
3NerlE05kg897njPJzrUfluO6kllHFHACL8qNhxggiGPizGf0vaqOTVAmcKbP/xv
P5d/SUb63YKG3DM4/lNmA9Q0cJ/tidCKUZpyAnRAxk1TyNbm64tWhqgnEz7uYuw7
mw9VMDmZbDu1XQ0e9gS01ZQ6bNihGmwVTFlf1VEq4B10vb+pXpJuMbNoRsCRMxeS
JkzjNtidziT/eGPkt20JR8Ugd6p+3PArjgK3t/IrGyf2xIyKckYpG85MhTFHGSWu
c3SkNDTjhMohOHmLdL1VWhIc6eJNgtTHNa4mLPtoGugBU81RS5SdDoiZKekjLY8Z
VHuJCvMi9YAN0BZN3CEich/zVSxT3/Klsksks8ASo+CZnkVl2X9Vj4rXO/rUkRRr
LAVWXlh1pNO4VEHfupcCVO4oPMoCb7l/1i1/ReOmKcLSLdrTqCznlRed/zAiPcb2
ufqldAqUOCZrsc1KJ5ZY4UKl25WyjNQpzIygbRtKgOriZ0nUYxp1KcRsEcc+d8ov
0cSwQb0faUlu4yEaAEByFqsbasL9vPpSm1HWYiH7MLkaO6KRb6LU6AJ/g9CFjUdk
v4ZcV/fRGAmmNNpIJ5YM0U3aWCa/B74EffLEtBqar8vo61/9QY04ZkpdF16inMWH
R48SBZ2Kr4v+Q8E0F5jPbLwAM9Jr14TQ8b5PQEHaEuvjZCQdg8WmlQqdgrsL/gLY
lSgfGhw9ivfu0tVS2uUvAAkGBeCD1mG1+5JjAKMUGuKLg0fO/hswvtJu3L3FksJ9
nWsKWw9ODJRSQYBk3YyP3D1DN01bpfUpNhAxvFqHZ3QgukM62MMht2cevFUwre9F
r2ikToZOm1GSNLU2ofrmNl7qV+C8wpnY9THVWloEnjg+g6wxDfOteiHWdVdxtTFD
2UIqPQ0GuGB+/W1bcwAOgQ60SaF2u5beUOM35kmoZGopON7LZy/P/f7HXJe3wzoc
6qpPWqxW36XPxitvgBOtTVOvyDogK3G85kvzw5JmZI3UYqYfioR0jT2fxOFfAXmX
/GElRBFWgoqnxQirA21sMvSih3a8PqaTDRJ6ntltVLQbmqS4zWwOc9XnqbKgKiwG
u32SW0W1lWm69HyFsu9fdtp3DQfrJIsj8YGPwibUrwVPx6NaJJJQ5uqT4+NPONpV
niyLiQMO+CElSAezAFClvAUM3IFDOczWss0uO+uZ+BWuBqFzyAutYe9uSO9vV+gZ
1iR7Kkuz1JPKqs6k3AqsHqMEkFZYh1ZZRTER3Ziu3V7WhMgSi22PH0HA2sUEPwOh
bKtXx8QrClHFI7iev7nBvG/qmpUoUREnyf9URRHDIImhnyHQYgjpk0sn+1jBhSc7
bfXkPXvJ9qCEr8ju5+yyNZDk/64Vp1cbK1z4lEpMvP5M9H7jXVde5n0brmJS/CWn
lxAMW5oinOn7MsieXYhzkz9eV8eupUNYKrQcPcORdcmFAxdk7ScUuCEvl0lmx9CQ
KRZJefu0E42o5mLiV9oyjCNEO+nWk9I6Yn0UE6wRT0H+y6dGUZDf3mxVu33P1Smj
J1gFMOMBy0nvykiW5yOx5UJlaAVsfAodaYTkEtPbuEIS5XRuXW3nwrqHdhuqDi3P
fWIcRJ+IZrHbtHqSz1olX4HkBEvAPew17TRJFU1fFg/miCXmSmM/kPGAviEiswsZ
KTU8IkdV9O/qE7qSdomAS3Y5RF0fDMI0aHGowW7s19OXAV8buIwJjCy3ZoxxEVt1
EMPcHgNcjj9JI5jiHypA7lggSmEpEieYvYF7tSXxwSlTpiy5UWLJik5ERmoSVDqL
RF7nwgHuXFC+XnEj+HHJNAvasKMeBVc2O3YRxUof7r2edzvupAyUVijzPty+MFi5
cglw9UwCrHq/XxNR2+LvoScU5E17BBDBhnSb8+HVCo6CZgBC1/ghJ3ux0MAEeB8+
cnjhsTDBLdRYk/7MwDoj4243P5cwuNo6ZJEZfcj2hP1F6WXR2zDqg6F7eWC1EjUt
+NKWrRDWjQto8Qqx8UCAU3d/JTvlGD4+YauYaUdMtwDH1qn/rgxC0PbCi0xuEIkN
a5LBbCTSoUFV1ktQr2iCx90Aoyq4Tkyr5Kh/I2k3MT/xDu/TrZ1ZxSYlH1s+QVKf
WrtlWbTvVqNoJsmVzVtM6aO1aZvVVRIhWsh3wO+di8frLhdex1IF3jmaLvE/GOkW
um3xRwIc2vqaKqL/xjcorZitYSeOBZehaLAVkKOs6X/FQxuZVH/7JSQ3n2aueMG9
C6Jc641dhui2guMApZc8blwYzHQO4NFQnpWD/774ZDO9R3uYluUp2XY3QEYQkfKW
ZYrnE0MDjEkY36Mt+OBOh8Cwj+xDj1wQjXgzXkyQweD3An0EttgGRC8wMnulPpJ7
F5FiXHkIi7kzeaXMebj9h9XJo34JnlGQ9UB808n6ovWr7twlH/n2duOfKpaD6KXU
bC6GDPvd9igIG6f2KzyfaN5RDGKnPkBCjmYrmkuJkEHlEQVWgVqZ0UYjeBy3U7rK
JdNeiYAx3qdCPA18BYGMsFDVRGThGxLYoyi0SgzbN7zkzJ/9M1CE2JT1qOS2kYPO
KtOA6GSt9bpi3rLgY5msf8DGCwFY1ZCOFswrFFNvGLBCtGzTstRGSlKt9Dtgrgl+
p0MkwjrH72KAjP6EavHblj9wWEJjoiSd1DZUbXAgA3EfHknJ5v7OURnsfP/19fEW
FuA0yGTXOAzeqZImhwMo2VpYFi2dpBD5abo2XJGUGmpQE66pEQWYm41mqlOsRwlc
/K48b1m5DlKSG5nct4Aoz1WagOdh6VAx4kdLaZFJSqjtT+KcSOv/PuIncB63VOjD
DIi44NISG0Y0cmzQh24WVW3ac7uY7bvVFDK8f7GZxfZnomDKuPLFZHASqp/fho6b
wfmknqYads3R4ZruH63nhZfRckY29YrM5TLEvO7wXUHJNjx9mbAPXl3saf4rE88o
HdBlgika4PfqAFj8WyGEz5bDGJE2qCPjplvFaThQXWY9HS/usYPg0+pmEWZ7dZQA
tBl9WarkoJHxbmYiv7BxnVSfp0X9E0OZXUlcaJgyMGov1rNcxSJFa0JejII3T36I
YMa05D/fEOQRdPUAPw2NQCVqapHUe2iUg1hEFTAtNwehenK4R5n8emjZIpN9pvcN
IUSjCK+eIwtfnIB258X7St1vgNnBoH9vADCcDKP0IIco8s/1L84gCpDFs7VrY6Ns
wWxuUY+Sn4hkA1/20QOl+zDTNubw/89fgG6fcZxNUYq/CdR2VLba7m+RnVznjfhc
fLD2w+kPer6tTcvTn8JEqYF3CPMhzEiKGmKzyQ0KSAD+ObS9yToUJuPvsxnl+7LI
+PZxr+MfdmnD3WLrvTZTn8bOccOnTqZ5E2lNQAbgqSpbQfYEzfab4OB6lhzf/Di7
3+TzaHSpuudqZDKRBfYFambVVXcRVj+QWYCwHFTQQVHNV8A9YJKL/BfcoMfqtqh9
tlQ8QBc+RfHHG74ARv614d5p2cB2iQb3gf2PLUDl/+g+nBixRfkC/JHyP5NZPsvW
O5U/USEtFSq5E8C5ZB8uGvtHuJjcryPh3hyn0lZND5yENfgw8Zh0RSXdQs7zXjRt
gpG490bdnxjk6cM0I4+JkwBqBYG97/UAgI3cp3yX8g74vix+jPn+GQBfzbTd2Bma
5Owb9RFomWkYPrQzdZQiNJmN0IxKBO/vbZGxqkoa7FsZqZSXJnsPYXk4lhIZcmhq
tQpUy8mijAdM6ceSt/wFgjVoNK8PC96kenJtzo9J3fpl8aOlYxm9I6UhLz1hijH0
hjK+RGykJZeztIWe8IU1Cz19a8DM+kYIJE1zBxk9fsby0Us7vcTjJSOtn4a+2uhF
jeGJ83GMNfjqmvIewA8hhkFMQt6JQNXn0a1vio5me4xlVoPGZgiPPmPydKTG/UtS
RCTKl+LT2v83wcn14yCx2bLtu4CxzxakcpyQgWXTXP/U6rsoqxshEpR+MgAuNRB3
zefnRW4GIHZyz+YDtB7MJmL7Mn9WvuVt5HqLHzNuQ+MgCa2Xs/MS22bk+yjjsONp
19NLs1NQ+HkcZYH0UdJ8SgTBxfgCjXpbLu/mGbIzL1bZBe6zf0i4sRz9m+P2isa8
ToRL4XdhGuF4aGpcfdcuJWJ35mDQnYpMJtRB8/J/5BF78hKUdSZdDLxo3j4bk5+O
FdlyvZAkQKHixX7GrCKbMY19wLvzQgA1IJV515bv+cFA6W9ShEQ6S49D7IG5alax
w/EjUFyAyMIr+jMx28EdfMLHemQWWp9l9eKKeG21ppod0A1kNHIN7w+Z6SU1vOZP
f9wO5veV6WmZqum+nTLpjPk9AAc1JDZ3QG/N4Woc6DfJ66jnmE5BwdbyclyOElq2
+4mqN6WeMi8R4S/x4yng7f8R8X4Hww1VYVBW7az9p59EZHLE5whtVaxGt8mWVfbp
QRpIXfmS/hrN8k+dKwfxkzAmBXzyUR2UZHisQVfQCAhSEc0BtRf22FuwFYU5g7yX
D/A95QUBBkYnnG+kjLteyL+yYc4YO/3+XFohRsAsBqmhktzoBRwjkYpkhwlXWBBi
FV0XQYCK2kjLsdTIh+KMuRHLdUKOCUb9jkwTI4rENCjKyvyf25UEWaNk/TbibeSU
YBfwGCjFjWrQnZJFkPyWTVL/xfOZuKurdKUNNtEVDPPx9TJwQeyX+j3ofxpPeFBE
ptvU3Y5+wBMu0ADmUf3uztcmhCEMahxreYTNhlIAmi++F0qCCm/5SPndpiXNJdF8
mfOV3EfvXfQqAr9TJ3ittkPUfGZQsW0vCOtzRCVW/H+YjeAKp4qUuNe2OJhHigaM
XrQb6TwKTu3K97bIbflOc3AySbIY9pjbmN+pF9Vve1fRiUCJhFd4GZRl5jDrtJ2y
JlktbV166Nmv0wsjTrM987+31cjjBSIzY3Zl74PUTQkMejdqH1zBJ+C2/0UscR4s
ZfppJaxPiWTV+LhY3LmH+9DqCVXzMYV303Xp4q6rQC5rRp74FQvP9oOpcaRjI4Zp
LjT3/zEivOK6DZU3bydIgFitXnXAl/oD9czHYubvU5TKdyaV0469Wo65MCI9kEpW
pA45ZAjVC/MS22DrPn87viyJAV+EiJB6NWOwiZxhOanI8H9peg2fO3IHRh23MXwc
Mm3he18oDJOqDOId2+FwwIY79t9Ref09r1Fb7rs++aIlW2INXM4O4Z7TetB2Dlgv
nydjXGsD4G31/a27rIAeAQlBnRIF8YK8OFVOODOtzvH5r1Spcv+EsyP+X6Gcp0E3
98PFk/SVh28YCBIJzcsjPFACXTgMuLLVa8KQ7ONgQb7d3pqFT7zQl7NP8pJFD5b0
ZnP5td78Dd3SyOT80D4k2ALm3HJsTzm0dgBF/HWAuO7Lyz6Sqxe2t8UWQ1ADK2uR
NrN0HmR7zSRqj8ia6spGKGCTXjf7xO0g5v1hRgooaJey5Ao7DimbctlOs8e0HJqo
/aYjDdGUQL4YtrHA+HgIz8rV0zkt0hzItcEY6Y5tZI/ZgFNz2TC5tAyLeNT8Lczz
sPvF0o/XpT7r3/l5vxNwhyKbJxJ30CSKy1NK59Ur+VYhZSbenwSd+bU55VmfDGU9
Zteid6mg+KTP+cfzYj9M/PTOuI4t8ID80ugofO2dnTsDIVH4Dg0ecp1+FHwJgiA8
suaiAl9Ub7WgZx3vO7n/8TWAkOtHypSHVZrhidQlayEstSd+G5LFF05aJPt9VqqT
Ppq/nCb+/3zZyOn3rqYOhYkvXC2u5FYfMLuqCQy8ZYv8AXeRsQ0w7Hnx4YcI5A2I
Eh4iy1GifrSqJV4cTZhO0L9kSzVpXE1QxEIvkIi0zSE3RVse/Qb32f3v0SpCf8gt
wTINho+2oYTSr4xJMWpvd8CSmwAW+C0+IXfQWIVAOpnxS7TfaQ5410344MczMDIB
/nRbedffqpOeFpdPz8D8VnWZ00VEmyDW8iiwxP20cg1M1aXs+ybr1CnP5G9FUHS5
QECKLTOihD/eUR+y0hY4HP8je0/sSLp8JYwN6T33366fVW/Vk1NTt6Kz7golLlPL
RochqY9bMp4EJlj2xw7kG+7YCxGTSsl4GEmx9ROIS9lk+P4JL1og7SiUMWqXgM82
CgW/3qZfSimVElrI7MD0B236gex5bzdGVjakxff6fiiXqQjL5Pg2tFZH7nKsvVoj
js91PEUUO1uGiAbahtE6gbo+YspVeQFZ5T2+n9LyXbnym8Wha5n4mR2QhcvFAluM
s7TnAAu5ZbQf8mRycVSb5Z50mG1+X35Ow833+YhuhU1XuwK/zyc5FfJ66gxMqRbQ
KRa8LDZ3fAjBq7hRVAJrCj4AU53mx6mBVRdteaiI/HI5HgpDSFurTL0xVqCmgn5T
Gynm9c9xQC9KSZtSKOXu70cIsfXeaQCmckHrcQvWCOWX+BpX8GJUQ5bzGDoizhI4
zd1WGFrtaNP/AusKZjFSu5AUo2iePQ7AF8B4FRzj+1k33IZTOj828Or8xYQeNgDR
CiKMwBswVgWxfDzpiRNu3CXKRLJ7JU2kjn2VtSaSTNW/EwN6owq7X6SNr18l5INg
uXmtGY/H7vy/KZALhmWYHB0QZaG1mrZ/PL4eEaZ/iIeUJUBQI7qxyEhimrDSucV5
knI9iYgHsvwKPQrT/T6Ciu8aJ3MTXU9EgDSkc2CQp9WkKJCjxI9GXYTv4lv/eHxe
ZQD1aN8m+WePY9bAanf/JYQBvfeSVObtSSydZA3sy3FJXQjnWi9XEwE9V9sZgkCO
vjwGEc4WNqsCWbnUKIFj9LuU+baSdLsQbWKQkQXhOYOjbpag//dUVJo+YY2bT32Z
qYc83FmsqMyM4lV+NfZ7mqxr9PewSiWK9KkFMGZTZqDOEIIysRdQxxiPOrZIaQcG
xvz3u2j/uy0lylx1h9gS34ALQU9RIa+RiYIV6qs8n3EEcI7rce8nxLRCc+m11uA9
hZjjI/Uz71SZoxAO3/EyI17JTcAs0e/fWwx3cpysUDajInCeRiGAOZjF1lDh0rn6
RusaMN7e3ou+kOGCHSV0AH1jZTrBLt6BPn6dLMZ2qPnPwGOwfiRmwNp0m/HwuyRy
Pg5sn5gqjnVcES7FhkvzH8VgM4r4LsnIodBStEkFpDwyhhP1+FHW3X2Mipbv2Vac
uRzi0huUs8XDL570IhBgSQoNHz2wpRSvW+d/XC4MId71v908RtgKKV2yuUaK25ua
oEFTlanehul09VJUc3KVmK3eWlw2OftoEzo517ZswZOsrrGWQvI33hadP9yqFJ5r
xzkU9O9XZbHc7BpeSKGihJhXleku1N8RodF0+JvmBDn2cxqUksQqw54RPHwSKrNZ
0x9qrWdKcitZZwch2xLlyHQtGyeM25is/n+7D9fGZJcaV0D9ZtJrEvp8fw+J8fih
i8YPWIzQdwaKOqNOpbImABRPpIQ/A+7bJfjbh4VQQipGMAfYn3olmOiBGvStN527
wG63vXvWWen2/+6DRwEeHwsCCzen3SxulVfRd6VALBNiJKEgXT7xLrWiZsdyf1JJ
G+AIHJbYdh4t7o0b7zXHc7qzYIA0Ngb+NoHCeE+okUDsZtKluOAey5T01N7Mpa7H
tnFjje3C6at7DUvDkuKKE19jvI5h4ZmOrx1vZbVyaOlYMnEJ1SjM44VDPlRyJZbE
iZPhuyvVJ47ZSiGLGoNi7h4fKw1BRDnMvWNiD1ozX2kiqqhV1Jw2DEedFP9S8P34
1WSATYd/ZBgY1eb+a/0UnwoqrCc+IiJf0QIz2nqvShAlEVEaZf3Ras3h742Hhku1
nq4fifKVWUouTOM4NsHqmknI/l82XhygJoGX+FloZjfkY7yRn7gxvCwdTGV662YL
+4TgnHMxpdeIKO0Vr6ScszYmLjDLfa6qTJ7medZ08+3z3auSEd8nFsVrMnJ4+XQR
9dPPbx1ISqsVcFXZUP4oIxf7NOsbsZmDsMTFJ9vvIjXeij6maTy13QEft8J9IDND
rRF1qw+EfLOPFQuKMZ69m/offx+qYlGPRbnR1tfNzsZUQKRloUg04iL4bmbL+TFX
t3qxVo4QDdJtTU+UQjrQ+q4yjYxStbyrtgRsEzOXWh8u7O+tjlko54MgrEBdZwDq
H00j4O1pVbgZaFpsrvDqNzkgE7E64oT1F0tDbjAih2t9YMRWFYMIA4CtfpnzA+eQ
Q1yB+kGvGJh6ecmFWxoZ7USrIkfrtRPV4xaQdqqgfShODfwIo0lQTfpL+2Fc5ciw
xoj3FHqLTQ0TWaaGYo9WPiSMmkbma5tJmuCIBsVuYV89AxYjVnAvZzD1P3hGlipH
JpVTR1Y/DmrvG58IZgg4rSIu37PK0xlvhIDVKnzrvrTt6tEeMK+4tqhxZRf9UBiU
BHGjSxSkquRe4rsPUo72Y21hLN23BKlyY7vRjsvlZOWmQj0x0L7qRhQ1BI5VQlkh
07NEQUoZb/R8W9ofHGkv58KUKxu5KzBaMxxsMv3JxQ1nBLg11nSIRhLz6oJowi+D
lJ4fvUcxVnqx3kclUXNk8zcArFNjdmJTjdE3ZFdgSmVoFq+TnVD2bskHJyZXdtp0
SMqcg9ZySE5mQpH/FqRlf2jx0GBFurU03cdml8B7jsgXGI+fQDY8RpS5Nw/xhGRz
GXifvkmSOTXEayh1ctecUq+KeF1Z1czkg1JGrTD/jU4xtPwefEby93o/WTeCA/0k
ORCjASNH4tAGFOb/2UgogIV/xGAojrYP9suwjmz43BOuGuUH6HVxc3qwYdGx6PCH
RSvAzcj8VDqveBC7GYgLzPDrCkFfngX6QtZvZtdINd/69hleZHIabD0nlUMTR6n4
kZa+l6z9LWhOPbILDQ9fuCxLrFZe+ha0/gGAdqZ6JcaOm5H5tqchf/sSak/OwjpP
iq8AB78LB0y60MFe0zv9LfXeb4BrtMWcvFP0RSZOMNHP5Hh0MrBe0KQxFA4tP1V/
w+zumclej4BPK1Rneu9MXiZxhoMdK5IhtfXQPlwUX0P+pUrP53T8IWS45CkXjIh4
pq0OD3L5dybdH1QTPn0lyoK98ohFvesDv3IkDIGVboNfHFOAdrK6TZUiltPOtGtP
KIA4H1etFSABrkZnWhqdWDYYsi8nr+I2mR3fjCheFQc6DC0N5phMf61mXs4KZNeQ
PNqObnm1VgyMwnBt+sWt24eXlmuhILTAHj9YupdlvEO5Ve8BzjTRNNRN8uSLfewg
BbBTGASF7R+HQ7PsKkADFx0XSoCDNFfx8QKF6I1edX4=
`protect END_PROTECTED
