`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Z4PXID3oVd7gpsj0rWEMaqozOmiSFHmX0kDsX0CF3ud+y7Yl0BGlCZJnqEbE6Un0
S2aeETjxA7LPS5GtVWMM7ayRB0JDEG7iC2au5CcudbK9XZpSJjCT8WF0K5G7YPP/
OWxVi2qvb9SilB5Z+fPPy/XnDbLlQ9zQlTAyl8bVqwPaRhmGGEQDEi7+S27197/i
8qcz70KiPBVWO0vDUjeraHNnC1ZzG6ijJcTIJ7wLGiwc6CE91l7HJxP4sYtdS+Q4
m5BR0B+40x+daagmjm7/Twm3U+leVbWGHtLFSF6AtkmbZtxUmw4cBlgNKGCcqod7
TZE7JC/QxuSHWvbJxU0bYh6OJxAeNZdmv03B7GyKtf0Lx8DG1A+BZxzaDz9wqLyN
C1zTebfqu97PpyMbRyPvTdoLHVqePFf+FL9nywxSWkibWALjoxUp8fznQrtWEHRB
QIyfkyCKQljAI+RFmn5t0WjUc2MihN8HU6P+A2XJn+rc1fE6JKuneoaYzZNBdelZ
lyTMRAEk11QCN3Ov4QfGzJ2IR25gsvQ0z+oVkv7J7/gEtO9aoaTcrAqVZ6tjt2pc
Lo27rLx5xmaUWQffqjoZiyqQ9/SdZFWAnQhWsWbfYZLeHZVDg7mJ2s50rfbY4DIf
qCmzWgpVxQExG7N9RSc+pljRYuHthtMJU7FQgZhViFGZhgfqsMvEHGfENArVtLY5
oc8oGzdjShN0vyL1xKfooNj85D5ZSLP3rqF7kB336OVAnvUCqSJjAqN/W89WmdFs
a1FqpsM89x/FUwPZKTI8h3nqHnX37sJhFE17LB7pPmvgElpzceBQleoHXJ1oRxVN
mJgQl5H+VxrtmlDeUv3nKDUTi6n88FMLaeN8D0smbKedjRtUvpTRFqbRm6MPzYwF
h8i18Re11CS3rDTudlLd4qiluYwI9x9sB/un+Sg/p5D+5/rSNAEKuIzUT+8IkzMk
8muWjPoOI3Be15YdZ+izeezAI+RBABBQChwc0ZvWkPIYF+43Xq5dfwCELVaYk4Z5
Dl5Rbsmwk+Rk0odpgI506Fub9D/8CYFvaIa+J2es3N9xkeiMQuar1WRBVzRBmBT4
TPBJNeXuWIiFp0qyI5UFeKucRXK1PAu346JLXg32bD5fITSlPoZ5BWf24vlyCr/T
cT7wffUtaQS5Ivdw4HBNlObJeuuKG+WM8be78AQHa5SUPbnV+k3Twr+BKynwUxYp
+xoRCyhvP2B2L+9yTJEcG5wF3ENGdS56wwXWMZP2fhuXrsxU3IYHUD+T82vtCOux
1NPzrBXVXzbyx3+tYACRKnsd/Ua4c1Xyi7JtFx19Lj3Bt6iNUabTMEOhNbjiC4L0
qPeg/Od5VHksUeUfpRxjqkGHn6QtyD19N7StfPRdahPVWE0Hd5NxKKAZ3ju9uUst
aBdslj1zkw5e3YAoxMmKBej7HbqGd9RuHFd0zYG/NUXg5XSUHK5E77J3OxOcf9OJ
`protect END_PROTECTED
