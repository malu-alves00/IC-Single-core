`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xMZibQcTXBU5lTznwD/k0VHFnvcpnh1lHGWdPBEyW3b8sCQjR2NDK77qCbTEJaxx
BHR93a76O7Fz4+C/zo5C81rDdchUNCena9L7H23aFXN7hrdx07jdhbW2kl6hapVk
NrkdRKS+sCxIWkec3r23V0n9iiTQhYRioOhoYlo36uo6+qLxzm6P9/xzCvbL+YKO
JgtUgUVp37WSuMhBznuvuLSwpmxBdh3z0K8siewX9CcJbP4WZtpew3CbusIBp6GO
Am6sZJFfBkIPMPUuLlAuqkFgIIYEKi8tLGbK1ORwKKD0WTulpI4N6WaAziat+5/c
smip930kVzxuoe1ovyHAtYDomT/sEJblDIO4R6blqtYxrzpqhNyq6YMLEorauX9L
Zh6u3vIuw/8Mn4KRcFZ6zg4ZyROhW1LgN0yJpoP0B0Vq1ZM5NE9ZApahzKPyrOVG
9DxSRjlS41YsNV+LkEs/HlOks4N60key+fGWuFj/GOIDSBoP7kuXBJ8uS1NPp0QK
r0+7cb3F9e+bR1pucTqz/26jnxfY7OY7FIs8S0iQ1ya2+HuvvoPqV75RM7+nsqm2
Bg1sMUYW8BBPDkg4c4ygZNdTlhP+jlWWyFiVVuC7qd8Gm4p179zWouYjV1WqijOf
FKRIyE58rkdgb6u+WW5crP1sigK3h7EHXMRndi15GTuQoIsYfdbWegnb6FInhEbt
6Mb+wtMN+XO1d3PpwbHaqQiLRiCsBVHL3sLamW3izff36USQIMPhF8jTXN08+xAN
EJLzeXD2XpIHO2HnMirPUoEpP9cnilE/COgNySlWiIDYJ/PhhOJ4IBsymWJrp0SJ
`protect END_PROTECTED
