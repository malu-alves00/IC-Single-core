`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
514wM3gX/ASc0n7TX0cqkZEVASHfCXD+jL9brhVbDy1m+jtaeMgOKFMri28nX9op
2AGtNpfq1lHgGx4RrnbHWNaXRQJN0ce3G839WhyGzUZhxfa6u9eihGTkztcnf/Lg
9u0pp/ffysyKSHwsXo1rjb4Qn6ZuWRD7yZ8k7ZxEgL7MnmiJrjLCpBh1tZ9r54P2
GWrwGva1uHxUtFgZbyIzO5l5+lAheOR6SSBIrgLGSFQr7+FHL/e4mUGWYswFdxQH
mN8qDbWrpR+xgAskor6OqlmLh9NDH/AQUElv6XYCpp+mlyfdYYNb3Ow/5Sv3LJ0S
vYBtoBiopzLONV3h5OffsT+koOPHGaLIgC18PEP69H/UpICtkDCylti+0mysyPym
jxwr+1wblduXKo1K/vv7tgGRFfK7DTtL2uCgsHvkCt8yBgw3q0cThqDvR+qx7pd7
EnvCYOUHwk3e51xjDq5L/yjrQvtTnPZUDczQ+8uHlzTG/mMGLpXUsJVii6u9gUND
alX41P5xYDYpP8piTgactzeNg3TdG7+XHWcId4E4CE8T66PZrGkPqZXn0EhNKL6U
nSDIPeg5UT3M/zLpd6dQ2wpZuBailcKUtrZzCzqNbaES2NuhILk6ctqeFyvXdvI1
ttTFBRcOWr/JC6h/XV1naAAluQDFivxX/obxr/X7MFiwQpPM/SrzPXGrw7lnDqU9
kh1Dui0a4R1gKBtd46d5B69GF7vmvdhajXXzwfQPxHzueTC95rYI6bxjELou+iP7
pexZ2QdIS92Ertz8INcpH5iir1rluzR2GUrweCJM6fd3aREhETFrZtlq3Klx+D/F
TRvIcotFVg0mTF7mElxsIIzX0aSr8u6OJFO0rl+QFoUccMvSkQtWcJ6plxS4aceg
fiXSPV9szBO9w8NJNuWPT7S4OzqNTfgnjHKkfqy7z1jKnUB68cMPGYhgscv2iid7
qDsmxkSISGRGFYKKcW3mEqH/roGftRn9gIYkQNsDfxlNd/cnH8JQwheKvve7TG0N
BvxpI/JoWFlgJff5CQESAHqdlrgL0VaX8tD7RnQeIFU+XTLdc7eNqVVIoVk/8/zO
4/fL8UsnUBjUb955RNvFeYAZ/MGBlw49M8mtoB2RSz0PS3n4gnlOUQnKeuJdE8wW
x0sdpW9RAhlqnyhZhcdm4CALD/6Pfe3x7W0XAc0aagMygLvvCcyEfBNCTiUon1iw
1iG1tfAa+PDwODLf76GOanW+tMg9FBMxItLViHqy9nLM9CL9q2f0e9JnwITNh7zq
Q++kN16c2hN0MrUUIc+5PNnItoLCbRrcY51IvEcxHSHQcJMGH4aMj8LYtLXvqgBX
u6omo8f+opo6i9/OMgzPKMzCiSxfLE/fie7otrAd/JV0szdjs/RHMEYLDdVpQVsR
XJEFrPUo7PLeHyjxsDZxx3BlTZ4O2KdXS03Aw8QoECLA3czO81OQ6geXuAixAcNw
oMFLtxOrYmKsZN6PwUoh6pCUaAxQ3MVmW4o48+LNAm/ca0dNLetxRN0u5Mgb5AIW
hvszhdxt2GYO2+qda4a/9tHHFrlhPgXUq6DB85T2pBH1WhI3wcQWXC68aD8G1ZkH
ECaHptXl8Z6wXwWlncKFA8nqf1UeApVJ2GR2HkUm9Xg=
`protect END_PROTECTED
