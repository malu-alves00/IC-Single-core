`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UfF0TY5FXRCnxr1v+cCM55mzu1qyqjIoSuY+fomPjKEv1I3kvVT4TToUZDnSlcCI
SdV7M5wDZANSfgFOVlRydptkPMZkhr2DTICX91RvXKxba8jdI2jkDA8njNM3PkDB
NTijuoTb28x2qiUf7xJ+/YDsCf0HZcPUef6ePQQvBMzOZEuLbudczaSPmgQhhgLG
7/Z0no1uM85PS6V/5oI47VhnDcGqtyRF4vT287w05wxiZK5sWNZlI/A9WYiKPCQk
1P9v2uDgt+0mrKG6clsvSZ+4APk0ecZ4W89Xgjb5jBeP4vXK6lL4w6Bv0QsoAGvW
JqPDFMzhV17jxLC+2xagOzMJZMaE6F5iSSH+oTKS0GIdpitc4q5r0ZZC6KvOia+F
qLHdd67U/s263Jj2K09ycDl7O/hQnhT/dpB9jb317ghZLeuWhch3X60VKAIs6rCb
1vLyW5C/FWOsu2L4yYrRzPa/DnMrJo/zMsO8Dxjhm14j2vpr4gx9vfqaWFWGxQSO
id147aNBv2kAyv/atsG9v8Zpr1bFygh3TzT7lR2yRydrlWCcKgHoc1nVsbfF2kjc
wQi6zpiw/dnjw0T8YhXwCY49/+OLhMvjDJ2/clLCCe8ynxd56ZnStI1W46+9R8gK
y9CU+eTFpBxlAJCTGxt5WjVw572EYp3ztNVjaQ/l2VU68vJ9nI8HRW73lIE79wlx
DjxXQpYlWDnYAnlnJKwF5q7hNyHPEj/I7PBol4v/g2iIaWg3mWM/o/JAi+S8QvsA
jvEDgFLceuU+yG8pOe7yRQ==
`protect END_PROTECTED
