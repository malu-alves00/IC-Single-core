`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8WzcLBJ2z4UdTW+4UoOu7HchPUpn/xUDTIS3Qw8ys//IW16bHv074ROeYzVVmzeh
yMB5QzbdtkN/oyhNluJbQx5LgXYvCDaZdY1ge5jf50gHFxkHM2W0KTQvRv+I1Ifp
JylGpm7Zt4ZLxYp5+QIhi1kGxUmCzCSizdiSI3ajxPr25gwJcqpmERZ8i+6bKjsD
YswdBVrV50flqWPerzukZ02z2bEHpItSOApROpw+aQfkp269WquCVVEZYVeFNBy+
H7FlPXdBqe5ovSnSodfnSddktm1ANHqSAqNLEbsbbAadKJ5/sGKKPEebxu/cc+ts
B9vhyEK5Is9JKHR0zmbmXVh2JRSSfmtsho7wIoMFP8+WBTHUyO0UVM7Twv/JqDEt
oS101REMy686gFM6IckU3AhoRwX64S66UIiTvqtqkbQGcPZ/w9cSgPGdIn8WrpOd
b2Kk6kEr9LzZ3k/VXVpmR21R0fgtn+7JplPBLwbftUAE7rEueWvIrRTAWnXYAd2a
as6kibDVBJrn4wIDPbobK+DOFFUrtAsPE2KAKkpuwSCEcRyE63UIY/EvJxyOWvxq
93L2e5/YxSuGQzXMYx9mhlY2IGlkHlM22+GwabqSw1nucKcEFTUM22jDEpY/SAuu
I+8rDq+wcHqFaDm2CnF9gMnVrjzIpxwNgxdMiXqIdUM05dMxvm5AS+WnwWYT20ma
M7ajohB/wep71LHgrmQwyEAFpm8KuxykPH+vOeQz584RkPuyWHhZ1hhFugA25ino
NssM03yfy7lNc/YIFaROGyOLjz+iy4ER9o5HX8NlLNkKjqu0zN/9y1nWB4TT4tdm
eiYseYKOlEG3TGlTCt5Jm0NtPe7Xh2FC7sW1zdbJBQwu3FKIvua9gqkljMb8B0/N
X1drrzHaEs6bVZEXnQtshyl1haHh+/vlLY+IPENGvE7dQVT5u0fMubMBDsTyy7Mi
Bm22rfTEmeYIAntd9Moe16fPuHscD2oSySN7dBwq5gXqlLNkXJ9YY8IN5TTnNVl9
66Zx3vPQd5nWAlbNU4IxKxoZCIoxZCka7iaDPhKSP2/BhCY6Hl2+kbjbCjdQcgXZ
BtlPmiAmVccweO4XBKQ1Rx2/+JKKN9U7zW/3eksDR5pK/8YBfKvn0EPft5RS/Ex4
IFurSjGrL6YeZVpUm9J6aOhflHnwVMwqs94+lBtxiHks9lQ3eHKf1T3tz4N5zbYs
dKW/tJxbLp4wSOtubK7J12xvuXhkhgcVp5j+eJlu/O8/ynDFs0dqq+F3Nk0LpamA
xQaVnO5ySBMBfLK5RswwTyECOA/lIfuoROfk687F5lata10i52G1WEnGgtfCRq06
35ecy2VNkscuxfzkGhe6BSdOv+QcGbWDj4WdvvGEyhFVblPEqElGZc/lbLH21fZw
HK/LGLY57tJNvUy0ZczsIy2H4gC5GG1eYkT5IvePWnC6BR+92OasiGQQmUdABAxk
hSvAGvl3AFsxIPQWAzflbshqcuDWbifFQw8XHPLlDTIPp52ttTD3FY7wZr63qNJb
x7XNm9FxCVjeoDuGluMm30q7evnzDrff1G3kCfkdoRFQ6NZhcSxzTGpclPMy26R5
9QO7bBg5OZgzqS50Z8Yt01AkqGD2eGqFZQe3wIV3dfQbuSONx2WputJZb6QlckqT
0fgF1JR4ygqwmpaSMfHJ0b3cPlPRxOOEPb6odpOLxuVI1ulHyh1R3/9PiTkFX0uZ
+Fl+H8gaiZw77/7LWkT7LGyw8c1F1hY0fVj1BunHCcmdmaNiRAk0qAmLYikVN3Vn
3ElfrjOyqtBET6rJe8ypoqRPf8TyE9t/7vAuU5PGVJX8iKJ+l9EYJigTF1u07T5f
DMOCwFIbZdJh3zRudF01WBnsPL9QhLOyEb5tkl/LH0qdzfLGbDQd2JwRkF3mhu35
2Uwl8Zyi3T3Pps1wPrq+ocCEq0IkVXDjej5ZFoeMy3ww1rZzWizp8z1/sZ3F+Bi5
V6iX555G+mT367QYK31fhyMJiyIcFWmgTB5DdjUPQJ86gKhOfxJaVLj+w3R2MBtk
Px1lhJwg8WxzL8vce5sMeB4upb76ZwmLhOfVobFej/aWvKrKv1MsSL9zwsgbbWl7
7qx+lVzZ4EVASRIuVuPuR1Wz6vg5EjrY27CFAtdPHxm3bCHDgY2p9Wihki9zuaPB
EEfnKAWxEjGZgiOzEXbFtzA+1isoIwIwVB2sSQbtwZBZJ/VJB0whrLsCXSRMgUDU
FMvp/ElTq9nji83yZUbBJpdEhns8D2H+jLcoxMPwIUioje4e9uELt2xVa3BQDTIK
DMpQCKtojQR/4M2vqutA8rY5ISe4T79LT6ntNMudavTPdRRskDEDqaj4jIMdr5RJ
LF50EfY5aonXBE0W2oZ3N0BPvs2gW7D9IK1MUTV0F5+eezaJemOozAW+3gd+PF3S
n7y4PNTycbDM+GkQpGv1bnEwT1ykekRIOY1nCDsf7uGTfLjreOPGtsK/cvcd8m7c
O+mBgw38dipmImGAbuWYV0Tx6ic7JXUsyaGt5ojgLbUx9IX9vlCM88M5NqjXR8Dw
rNKIik4duAaCiPadq/n9xkYSOMjm8iwL6BDkooGqV3TIIwZL7o2o5zeD4fz4GYoy
ePLQtC7gmjcAcDHa3U8OZMqb5WpLYj9+rmiHLXdnNa7nnxR33Xq3Ae2GuqgNKQGM
80kKBBIdHY5unjC8XeUjIt94YcB4dQQ4KHOFGU8gVmJH/QniJ5JXLXsrysTcD/1a
ozKMs/GJ3e1HkYw1GwIMVwNgL9j1xO2AzlIZax3NQxA3bVmJj+zEwLoxkCbIuIBI
kyyiWDwpuTs89Mh66N1FGjuAFyVC3ziOhVBfmvXksgnjPVo1aSOhnUOO1k7b/MP4
u3rxGFUStDg2ZdUGRZqa9o/ZqA8wlr/ECg6mkgOJkEN+T/GZnmr7VoQRwAKj9srE
1mpwehTFAyB9dY6wheeCcB4blr736WZuQKxwLCev9wQCAlZGGccCLna5sjDE/AlD
CucxtrwLTu8E7dfndZ0z9p+U7xqJCyZ+qj8nWHowVqgC4vCyRq892LPL6rFbRwTy
QOiNooSt0XE6LySUDh6/V+3rjaJvdTDd+M54vVkTI5he5wWDQEjvH36YXhb5IDEg
OnlVIiddnoNyL3gW5op1XKD3E6DJtv9AkNafEDYo+PmvgEslz7bK12EwbAqY8DF/
bSJBZVQ5KS4O0pgKQzronASP9lLHghVX9rCGhcxuNzwhQTQS1zfVAcnJ+TL4pYXi
45yrbuT4tkDliwun5QXR4A==
`protect END_PROTECTED
