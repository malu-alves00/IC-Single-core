`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wEGCA/jxBY1vhVhCSKrC7wNsl8g2NkX5Oqr0YsI8F1+WUS+DJ06qRw0n1IfW3VTJ
1jmdQerY1eLYNixyulvTlzHfq4189wJgO3LgAZ5PF2W+YAublCFMRzNqwAomIl6U
6gOCvAgGTg8B3behKp+RTwuK266hccGiWNejfHi36YQh5RPoV/4WcxI0zjQdvvvY
te//Ue6NEaX4XueDf8pjP9uQztXQCQJTulzF/5SN94XVAQvbeOdkMoey1c00umzG
AVyM7Aw1lWil+xNnuK+5eOkcsVv9En//9gIAm82fpKey2a+b5IxdM9fUfLiHLChS
0fCNllxFGiCQA4Xl7v4D8CFwNQC5AK/F98McHMEVfWc8QCNP+hg6JY3JXBm9FORJ
Jue2ZwyZ1lMJy/E51n8la6cq8HOw5uRcLvUSEhb35q1+I6yQTVHd2qeZQMQ6pbLL
gaJTwofz/WZ4dlut0nMgpptAJtYp5s2OHdXYYueXr+B4dwb94C9REfBRu9I+Qe97
ICv+xiex1ly45T0MiYX5h/mvUIhx5704gmhuyuJWGmrudT3RleMrFK4lfLT3b4SP
T0XY3Em7MQXbyxGruOtjlQ==
`protect END_PROTECTED
