`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5e4GoR8V35Fl4KKFY4TbGh0xpKSjDQVFohC5aQHWLzvWqhRKeq0FcZNy6AjITdRU
parxmvcf6Xd1vX6yTipUnpJlapBqwTF65F2Kz+cjghyDmKyrbUc4YU6Z/hGRgead
f61D28uPaicoI238E/p4m3j6MxjShjSzwAskj0mtIEgLinr8+0yT1wJF/DeqHEih
D7cDfWKNHB3KJQA4mjkpBzPr1BbrrU6TBFkJMtY86XN5sascjQ+K5VmPu3MTgJEk
qCrSeDubfEmQSJ7g0tdg3498XcgsEzMMm6JRZAa7SS7W/g0Ljf4lJLu1tH89EsyA
ch4hv1rhcV1A64liXRjpoLUk/7es8Iynwj1q8MIC+ObB1rnX0rw2TjjKzPy3YLZI
CTgjwutiEVY0WwC+SkfRaVKFqDp/DyFzvV2MEXNM80/XS6NRmziQ8+KEiMwas93W
mb8ZyFTkkhJytOr5rT8hAKrrUisATQhqLRBcW7+g+RvEbJr/kv8U6xXdDwUdqgOT
dvAZvCYtCueXx+BovOLwmxAAoX+otQNK0iEoagN/CWbZpMLu69QhlMLXL1cqF48j
EFYiAQ7Hm5YiRPnkgOa2xYNRSCx9s7vMSrPaWqfceh1WfExwSj7HVR+G7sz1qF2K
wAgw60hg1yRZsdEppsXBJcxgNHlxk/l2xECMHig7NuVeKmK076YobapDs/79KO0S
o9TUMwVpbfR3q27m6JHhAVXv/U9UaQOOFUMdv5HRvXB/q0Kj72o8tTGJCIT6NNXG
2D8A3dL5vlb0nj2ry16INzJ0u2YLhfnPdie2KdyzeDuuhdLxX2CFxB13+aYozuwC
`protect END_PROTECTED
