`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qIAb7DLw79ywXmE1rxDrxFs0iT5LRREP06AmTPoIuw5H+MmXOifoHrcj0G0hbzvZ
D9lW4HkQz1AxQ+sGWs22wWUU8Y1LFckzbL4yZLckjxKq+nErjHSWNqZDe6VH6Z20
M/6D2RmpLFtJAFqrPJEkGCvWMbZV33oTfic8qWPy794erSVlBxMCjHT3+tXRX7sL
hpsUVhL9uNIz0RwSIok41t2IefKWV7PXeZifWLcv7X6rFXnR2v9G7Dohw+qZlCNt
2p67WqoGwOOgn6dY6ZvOMQrjMMy8j8eVwnKvTTtqeyE8CO74cv1EBzghNxpICmKK
98PT3qUiNh30juR7jMxseLo+9OHMQrcFUVuVa8M96FOCpzY1/V0seMSFTVI9c2IE
UAS2ujFSpEnzifOl3fPoccfJgAamQE6biO86R5EcBJHWSp5YSl8WJfN2RNT2laO5
M5mncRdZ+foBub4We1hxkr5v9gejDSm2w3JkErTcpptN1Q0lveTb6vpQOypZYAJJ
ktbNw0iGPX8D4/rYQmCWzxDclLlg5dNntUX4gq2hbfOR80Td+mm0SreFgDNkNSEe
xtp5bMsofo0etSerYdbcSuK7DO9wW50o2PiSt3y2RuxmcIqpxIRt/JdlAqHW/VLc
5KNyDG5E5hFmB/cYjMm2AAXUieYhNEoAcbbbCiiF6eM=
`protect END_PROTECTED
