`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5sNVFwKIPiKawDSx+5avHdkT6n0ScJiwwxl1B5Nu2tQnoTJ7uw6eClYzORuxfo5q
U3TgyktnxUCJURdP66bE+1bpv6G1gd5OjE+NwGP7uRKcBhsK3DXMPxRp555UnXP5
TWp3IbrkFep1oeNc+v8DQh4ncY4KjvdkzSikL2BXdCiuq0uysJldXLABp+/iw3HR
TFrv6mi3/5Gq/2IjPLzRl7oW46lLM9RKGJhblfjfLRp8u9VGKGTFwd/FxX5+hISG
8byRLb8N3r6nH9ae7IY+EKLs1hNgGXO8QDGT8omzko1Sr2SRORXTmtELrLVLagdu
XRVwa4pacPJkDe8vvNkkUDamrT4j+8O7p0s8C+AJclTpcudWHuDfnonTZcKeGHh8
ZhaDT03p1ubTDDfh0nAJrLBTEThbzURbhFdU90E+vWukQKjMQJFvx2dzM8KNc01J
kOy5Q1wzu7lmLxAyFVFtfSq09+zx0+VTPhw2O7c3XlzxV2Kuuv8MFnlj1TId462Q
M+bl8sl2NwaJNriRxtfYACNsNWnDjVf2JMMq7TcJKrIfQwN3QFSsc2fvOGh3zMfX
TjquE2k3UFgh6UPlBPEBtGvUgGEQuk2Xk+it664cE3spqk4nXc4nNOW/nt7R0XeV
P5lOhYEUozkpf0zUS5MlCZE2kZDBP6qMVFI3OKan4+i8za+WV0hSLbO7i+SaffcK
Qcd1EgehYZ1WgAgQTSDo0hlDRO4yfivZSdTLRN7ssFmSF6bYkOn6GfsrIw+YCTcz
qjqEpg5iBCO/2Gy6ejv8o80CznoZcMttNpyNQzQnaGfXp5TnzIGmFD/h5DskTeQC
zAlI2FfMcANKlA7CZnb17LwxuQFtHuukQQT+k4cl1yi8BtQR9lI6Ps+r74G/S7he
UcNF1F6ARsH4xzReJrj3oJFZQaQwZY4sKLtqP+9288Vzfcg4ZCV1nWZDAmhS+LrW
cmqbpPW6ez5Sm4YBGWvZMFXr9vJC4IMXBWyaUgjlra0zERqWVRdxAvL2708h5LDT
j4AZ8s7QXrT0QVRpH5uZ3ZcZqakoFIIasPgs0f+n9+Tn7NNk5RRyFx4FAToYteKy
O2s97rZ1DOxFFWZtBd2QLVv2JAcBfrFlfjfH4jyfz1MEg2c20ySS4HXc8a/dt6Az
9PxytyfkwOZb24KOBZPU1jj9b+VhcEGY8WPuyOK2OlQUEDEafL5Vuw975MB9630N
NeXIn0MQq8GeeKo0dAkyU231In7Iay4pJQwwflRIjMNBM7wJUkIC0/Z5x2aYOMpn
i3EbK66GQRfxo6CnLryYuwIvLeXaG09dJzSfhFJgch495KfscKn2IjbAg0WIo826
kt+2dIx2W1+rIjIjb8dxuTbzsZU0DOtAOjQUZA8D9zciXOr/lc3a6pGNJLFqU5az
WeETFMHq51Kpnw3GQrHAjVrtptg4LehdBZOEOUcoyvHxoiAfkP8TYTU1OGpmAfS3
QTx5tsUhr+WCWX3QLgr3SLwWvljD6oQ4QDjqcJR+fXsqvrPg1AUhp+ES8BlvBtiR
KhYx1HrxNK3Y7Pky9ul+QZEt1Hj+1GZJqRXvhTD5Oit7anIAN8Xe9XT54D27Rbos
N4UjSBvl5+y99beq0sJVGwBtGxdlx0TdvhBBa8friPGQwIWx3CzfV79UKQ1I5aFp
3l6xgLJt0RwiBQZtGTQ04Iumzv36QPW3orGsZlCpdvl/dnQd6HYviivakE8lEedS
/rRBILP7XlIsSrntEzHnIkAU+5GTQCdTjOv53xlOQ7Ivq6lpjaJnAC7lbZjs6eC7
lMgU9jmbuYhrAXlv4Rm6v7ZxEVO7fPNGWKQrbgliVrnWK693zJwnESDrNpVgZeTA
jGtmDI2yTLtSBkuyyTxIufPIE0OvawcnIt7RcbV42xLIQ/m7xUnADb7zPhMPluvN
yp8DMmq3I1gnEQOsB4Xnq5jEupdy64747iCt467IctGBsWknTw9XQY8zkmm6Y/vD
E7xXZioTroHgFm8ThVfLFPKsBK2K0i3vxynWt+PRlIKpowy5quUiOP4zAnJ8tRUM
+Yz5Wqqn8R6gJNZqz39kulUkZRgH/c+x5HKDeuFO02K2dzDVZ7A3RMfgC7zwodp4
fus/nKUNG8K2QrAwmSr0QmrKIcaOlob/iRX1R2MZbCpi47/V/RepDW9WFSMM6XRB
d3DPZLuS9PA8PaJ7F5OhTYtUDX9S2QQUMtaIFqwBLeldQgkJTlV6zslr9E3Hy+Te
0TalBYE9kcK513L3X2D1uYp3rdkJz5McUAMbi/ANf6m793cHklr2t5rMDfiHYjpp
zBUH4xTFhtMDZFI2AiApGYZTerms93K2cJ75xoI6RTIDTP8Ph1SJBVStVa7jSQim
OI8K1TfDCy1PzSlmOVtFzB39CcIq81tcAkos72eehWJQq9b4qODQ1v3M18FdYm5/
hrdDN2eML0JuKqJmJbQmjCkoaxTe/0/PKQqE7xdzS+XNW1LIvn5aTXrBPeIDBOqK
YeVGJLNw2fYDFyVeLdl4a8//I8JHM8Ubrpbi9JNsDw/0T7/wMNAR7vuCfRGooH3x
fZ9txwWX46Xnq4fMCvp+J08W2VF9S52PUtE99WliQHMe4XGxoJixTgBRRFR2OENo
FmP0spTGR67CYVTO7JekFRj0AhXgRW6SQrypoIhMgMBYFggBcaOdKhwE4AWPQiX1
adz8BYa5Ccjx9AnzjEvAqZZFCry7WS17W1jTYLsNER0Vffb0nbrePlNa8yjo3jWj
core1t5l/gJS8mbnU5+5HPJqxT14Assl0vP4B4UkC4QZIx80tGjnJ5Yya84gS1jd
eblcT6QM19m+qE/eS5dxwhPtP9S8rgnAZEoQ2MWMRYYVM6WOxC/THdm+QZmzMfJ2
5bUyGPYuzcOo24cFJvoP9YpLoqoVCaSMTzjp+PTPQQ0jqiK8GKVEhVq8QnD//83Y
14zLhWBNh77T2SWuBF7JEhLYszokmUkTZYfec4A7JvkhzrNA2hvNRfXRteYAJq9+
eYOv58Jell+qu7pyo7tlpE4gPrAduYGNIucga0NXGhDqzTnKfGvRDOsyKIAkp01g
L40bAS1HaZ0/bpNly3lbrgyHMirrXueGP2yi8Wx0IjbFeOUdiWS4oZueitzLadYX
IXZDr3EnqRr9pRypdB7jaH7zrbH2VOwvfKpmyt6WrmB4WfeZOoeKO1pSPlpj70BJ
9pQ1/EJku2F0LctBqhZK3zjCng6sc6gUVP9C6wHpOZcMs9M4luZDoP0siNUzZZrs
l0rtk6HhVBrx7w/4F7/0Ae5GHcQwfbul55tApdCQcHdgNsApX6KfvOST8cQSxTHt
UkANvpyHOuE1rX9/2HGgQGNZa+KgLRI4aK1PLfJN3aZN8tUmhQ1VBkcnGh/4lMEz
f0tn7CpXxi1/P41fJPGm0k3SJawaFD754ZMcbS0ueW5fe4f/+07jbw2L+Ne3uE6C
xCQtouBGMYdgUxYbP38Z2LYINVr5R5fqhb7MWcU/zH4CAFXNe39KOcrRcyTlxGzw
8Ne20khzKyf2DPsvVCTUmLjVbMpFlI9GKF4k/kLFi3//eOrsPuoQsu+qjJ04uv/p
UBD46lQbt7zHm35iKvRkRdSZ570/XN/6G0Xw2w6Ye0mtSKX7M8W42njRUpQRf6jj
9cFxJiHCM/mrvpK3GGPu24PjBoZ15x/rlFixhWswmpyaTGVvx0MGhfoZhkJxdkaH
YsCbVnKCyIg7v/0ecQiW72MNOoqB0NcofsrTHM+b8ZxtubkXXDhnsQ2JI/gLnKFz
VNIwApxisRnjplulMZ1eZ2cMVb4eExJ6SMsHirOYSct7KsJ/Sr/u3W5GJMTGAwPA
6g1vvF0MQpzGsc0KATJQVumqQ7+KEYzLis8U7Yq55FIohA/AIp5+/E9gvXcKMdAr
cJ0nStvkXO5WuqcuvvLkrOELCr0XYTtkIa4YNTGLcczY89hC+OS7ZYvOpMf1HJea
2Hl4JNj95kNKPvcIWlLia7pVt+ppFuIim2cdFMqr1xU=
`protect END_PROTECTED
