`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VV+SRGrSEGhqjYlpUotKgJPS246FlCde/H6ABcMqPNe6QCTo35OcfhE1WUxgkhFl
Gvq9nAEPI1yZY/MHY92s+7Ns8gmmsg+t9woZRcLTXJ6eKi1HZJeBMaW8t23mrfVy
Bg3GGwrIKrZIrznRzZYbWfEesiPKjP2WWynmsLdCKwOv6i78gxNnQoGzRsZGTSiI
WXiuy2/E4NLb98iy89GHtlSXHkLUzLiGa5aHGyTE4zVbxhmi+E2hexr6gsdH7NcZ
5aRbZJQ3YxmbDwejAMa/3y8LknTGdg52AcJZi9P4UlqfElE1oN32RmmP/DzprKMt
eUX25eex+eEDI0aqtjYiHuQbaPsPfXzqNFfYPxhfL/+TKRboMzxoL7+t+pmCgd8D
zg185TU53Qvqnw4voBQVWWON+/m8n6lWC5WmxzoyVlzbMozBxMh1FkhBa+KlD/Nq
k8eljnPqPDxwk46pNpSQoKBYKLK53ag6VGBqAFRcnd2jYCGZAbyYOGUQv+SOa+pk
DwR/GsIdpc4aAtE0SrB521yh6xH6zfMXt3H5MCzP6sz9cVSrtAblwZTgu408BBb0
cVEd8jmGtEqtFujVCUxFf5ZcC+zawHDMnBr0ZKdw2B4FwfpAZPtcGtF6qpzo/AIy
060rnsN+GodNTI0kFNtqwCV9Nthyu2pMOIrNn3mZfAak6nXxUCQsvrLuJPo3VCf0
S5erV9pTgmJBLEhKVxCRqzHuTJkjhJF9ogSfHWMrXuZIexJsmCMvWdYSmra4GFLn
uaQF3e2X1iAV2vZ1QKdtRhVO87o/SG3yCsxpSXj2h8b+7CjRW759hoVUiDTERd5g
ammqAIQKi9MG0ysn80+nQvauK6HrUgxBXbmgTpe/miRI+OAd8gEaSCR8tZPpD5WU
h45h/TI/gr/i2BzqIjsNgjyKIzJBpktSLpP1vKGgBFKMI6sfmIDmdtX4ifwVrXdu
uDohz6kHYs4BVlTkRaqCjs0huzR1mZr32LjBIp7aM5btPVnsduvcR3ilLKaAaedn
ZS4Oekd3a3FhUERUsFZx3faSh3hYl7GXl0YjUEXp/xR/jSbCcsaymzbeQjOHoahS
8jTrBzP00K+Ka7llavKdGqf1wd3NNGShnwhwKbMCWgZYaWCKbf2VlvGnleALxshZ
rbuEDHlYTv5ozBAE4BczhWAKZSpmrhw3ZUB3V0T6NjAE5pXLyYzyRFmTVsU6vWZQ
25Ota+mshpGRQDABl5+0tPwhEadJrC0iN+iCaTkuN9Yidj72ZRCU2JH251GtT/uO
HA7lRcTRjswQ4rd0hdcpfv179FjLCiPlKqJlI7xjyibvvxlh7HvU6AtEIes8JOny
wNBMrGlpyhWDyffbtmI8QUTVEBl1MiP7uQNkgFv1zOmyVDfUb3HmOxZ0KBEslX+j
RvC8pmKgKv684TUB/viH62YI5xCMTMXHUweEc07xEsO/T8a8PwWnoiBBpdkTNqUS
f99gRsg3iJi+0gEDCOiauqG73hOJ/7FYmftCHnX/zbBwfdIU+BUvLQggQPKIxWky
eVeuI6xbRBOu/XPZ9kVoMf4HkWf+/5EYCnNbKp9Fc+OSfhwI2VFAsiGXsat/TfLC
N7vcOZvNgRCFgehM90uTrY0sgVoksCUSE/ElROlFTzll4IkoFU5vz/WAK+uq2+58
muT19/Zo6sMrGJoJEp9jQF38DEJRKLz9oL1p9fx2EkiDGJ3L+x27fLuPxCyhVRvt
W2/oL4P/hgqfv+jSQpYYsrkTRbZYYExhp0ahkZjrwQNNIWZ6KDz52jc8F5VGscuA
N8MPtg4qZ4mjBcVUdtPpgCbTlizcUtEQATawbte/3xRfmWx5u74sgLbZ6SYOJrpt
CVhEyRHdD4ZmikwEvRPRuphsKwUPSyyR9/lu2HqVrSA4WyGubtS/8cczdBXs0WDe
9UwbnCxh4k4pKInyY1WiaMBZ6FhlAQESmVrKsGnBmQcxkOF3kqC743GA4yvH31jt
NTUpozi6vwWH9uxOZKHB3mAI9849W3FxgGt1sbsKkc68uy3V+MknuSMrePutxNNl
b+DfAQ90Rx3AFeTk+/K37v44CuLgNeErwNoJ+3qWpFIGgPN3gXHhyrhqTCCN5PSC
gBBWorCeRufO3K/uwmoydmC/jf9g5NLsXbygFuX5BWX6+QjnBjjA7WSrFzO3L1Zv
UYDz+N2H/THAZOBckG0E4cxyEbp4Ay4LuWMslH//v4Ow2Z6UHUum5mw0ZmDf2qQw
213yKD8BBEUeNMBXP7LKwqbvuqWgNfrl5eF8AB/2+vjti6UxYW4cYrBeqjnE0d9M
uo6zUjfKtk+yBh0yU0CvfQyE8lWtl8STJrEBVbzBmtGhWm5WysHcv51bv+qT4F+K
jF+uKIsTrPwXRQcOFdKCZyTKOZghXw3AXgdlLkjeE/GzWnt2OCDB4LLRKNI/kVUC
9Xmk4mCihyFD759RsN5eBlFqLAGCpBZ3yNlu15guxuRCkv648elyfAm5j3w6SW52
9TK/Ws8imtQyswzSJclq5/Xt1dodqg9Jd2DJZr7BIPqH25gcaIOW1VzO3KN9NVP6
mY5OJQUPE8nCq/6Quc3yGR9RmBHkQ3zm4GiDGbHdyuhWx67Yu1CJj6uQNv/KgZjD
6PLb5b+4Va7fw+Fzv9YksM3iFXIEPEwTxQvHhd9vxXwWsjvm9wtgUqUmerOnFOvP
l2uxREMy5kZ2x5qIRGoKC8USb1NphODKCRHPYwjAteu1cWvsN96BtxzId82+ZnGM
Pl6rw6kse6u4vPZkV29qPszhVcNNdAaReWw/KgMjEg9BM0E2PK1xyOLrbX9QB+FM
plfdAgQwP1g3GsTIInLLQh5qH7Zc+D1fRS/Zc4/lSlYdci7hve5GawwV0OBfGTgn
wsQ0Z1sz1C2WUehC7UpBopCpddgcj2H3aXxpzCaUMUaIxn1OEFIwnoh/VMoZpmW5
ysIljr1kt25sqUzmOYmAv2U8GxuF6meu7fC9TIn086bCXh6MnDv2Ik9JCcO+NIBV
9wM+5ilnlS/4n8euRT3Se026DGH7aufEB5xcoAdiRkzlkHlNH7S1mgbjJZbxqIBk
TCpC43kxvPcFlOvFyg+A5M1lYtEMUVvNPo7jpdVuCbYu/y4f0w5+wU7FOwuqEILb
nAzqol7eMHKP4aGuweN/5vzp2kigFkb8ael3g3QXrOtlpI7mB2UpXsrGr23CP37m
OOQX9VGbcQmRPEVqtt7aEbJbcs8N9cMaWB675zXPXEBodS5eqkvDeA/EE9LPAVe9
3Hi+XlXB0NgNh6YNvJyCTUq0QAnmKs1rE9+b5PLp0pMSIPysCHOMBXiTilXVvutV
zdEo7uzdWNiCsOa+ZNwW+QZyPO15+/QsmqAH9hTpC3+rY21RjCYGgNUAQ747qiRR
WbmlTkgWDp/DVddgFxy3ftiZFktJvb+v+jC4uRvI7kBA5t3EsoiI55I+pBH8ICxN
OfzUwnzVZslwBB/Ul5JAv5DCykeHRA3ZN9zp8+EI3lMBLuG1Zmj6uxlbFEtuMfXX
MHfp92m9W6Jw7rtEdccyNCDi4HD+bLvRbXvOZxNJLD7V4WvTarA7gf3gXBr2EUfv
Cx4x7L8AEwNvsVCQ6r9YeW2BliOhcY04229j/ddLeX0yvo4kCXEWcqukGBax/FmY
1vqIIvHSz2L5GOYvnoz2XcoVWrTVDNG90Ef7mXeHGOPg5ao+Vd+Q3t+uGPgA3DYR
diLoT4PjMF+6bYEA5wLzTxW5cpSwSx5YUFZ8dqUrGXH46sktTrKEvnCgGOqOCI0Y
vGvwLE0LmF+7c02lgFhsmsz3vyniwOSHIgeScllwYOMSCTa4J1yEpkyXxg75OG6S
550ok3h7YWfBFMomeRX9YWf/9rR8YFnlv8BducdtSKqx+8pNgHGcsUDpK8ETvcPa
ce2VuJL/S9WgGkvmDa/pFB+ynw9QaDFZfAH/xrJAqSs4mLdr/cbrattlmTO7As9C
AlMXmNDL4fzz5CIzi3EE+RESuKZ/d5Y/gsVyplBshFAOPP6GJ+wm3msZEdNvEJKz
B6aI4aCJCv3cFK8aaEQr2H5k6u8w7sKMPfmEiaZ0fIrbQiIiinUYbsdL6a4kAbDW
ALUbfweMTmWMaLlOWDZ/Rz4JNyRv8Rl3wDOGe7SPql3vVOnJC3d5BcW5fSZUYLu8
bCsPUQBXOEtY/4acmzIV1D7jaYJbvLQz4A1C4g1tu7+n/MRZa6ObWOP9Ui9akGp8
/BLIX60mhaQAqvpQSj+Y2IEipjjsoo9AWtu5bJ2WDkYEF/rZ4U3LzzJJvTkhi9lP
n6M5FnWJz3Q04CQyUjAuXsvlMAsWb02VTMtajgVgT7Zn2YVFl9wG7laZ7m52w0vM
JjLHe8eIsuGyNfkbqxxOvZZLOEB9rRuwlbYYdln/WoiaIUR/r8h6p9lJikJdEzqB
FechxrhWVVnxOI9y9IKk+g6oVD5MdJ/BJoffBY4m2Rg9NWrH+yV7WAxsSQDlTaWR
EzyGs165gPVc88J4yUw1R0Aoy4EVpdQU6j1jkcWBZaplob8bD/yCsPlIDzf0a27f
HKB/gWVY4Av3hWDUuV/XHQKmTkoQhFp/zV+hy6TbDatUoNjjtP0Td0Cq6gQhjVmX
durDkNtRFl1YEFiEHCFzYOq0aIHoMoH15gqnJBnPmLn8IWv0nVzHqEmglDc3Bbsn
f+4ExpfEdXKJeRgm6XXfUgcSHYa3MiAPY8lR6+fcOFN/PzM/olwh9cJ8JAuafLnY
PKHElgJlm/yUodGOji/4MYw5owdZUmgmNvzV4yrla7XU7KGiIVpgXCiQXw+veXAZ
YKRH2SISN1rYmsbIVs5RgAlaYV2mg45qLaI6wt5bWDGYCKv3TfH3XemJb6Yp0beW
GRB2+fKe+8wUtxIXh32Cz+p5ZFZAofG11larOuYorxEubmOzgJFHCFKU5cItQs0e
`protect END_PROTECTED
