`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BKF0dbxMfssm6fvjRjxfjiyKD8Ewnf/bxxp01w+uC1wHS04lIni0RpzZoerpJHDq
NU1OSq4ys13Lpwcda7G3Sb31yfWPKaTxTJfjwR3D9lomgAScLGd4jw+f221cFfyN
7E1UqGbCCLY6LAZ9syeg0FSFt4pxx0zDVGlyELiZtbhsly9XeDAM62Cvngvlk3rg
mlCz8JkG7ngivAEjJkBNJI+fkKMzQil3a1sad1sdtgCHEdX9h7aMVfzageeceoE/
WAiQWV7IuLsugLysZsIX1P4B1t4YLIr3Rt1R/PCDLgdOP3nKzNg0lhZy8pPFeSgK
282+Ayf/2WB/u0UozoImfS+uLlgZFtp2xjylfKZX74w2T1bEF9qvA6UcMrIungBI
b4xwk0wn9jV/YnPDR0Kv/sTQq/C0fvXlP0Ux0CyQGru9AYLQO47O4sYkE2owxNPD
BsjhBobQ6IIp8/vfwEMR6YrmwJJ09caHDGptnHLyWgNSl/ryI2NJ+Kk0Y+aOf+FF
YJwmPox4cSpw4O7S/h6z19bi5BsdZOU8DIvlDIklcUlfpAQhRXRND71K97RHGk1p
TTfRqGUpx6lW77a28PcnG6SzPbLCAJUfhn9KdLfPGNXFyiyBetb3Qwd+xNjCpDNo
mOI3IPMA0X1qxzw50srVwvjp9mBMHDorpPwR5nP7v4TiLklvRZsDEH/RNIuf3t5j
I41/6Sb/ri0c6BtTK7OsRGIb1qZLq5XNtszX7XEl36waXvh++qOkeeM3Ze14927A
UTdNrUU1fDw8Gsg7XivkvtN/PswbnXId23i8z7m5I26o88lCPl2gGpSyfgbB8nZG
Z1Kd1EYTxe6ktjlaZT9Cl2v9hS9F0vDWi6Etzb1upR3RzuWI3tefGc+xSFiY+mBp
b/zOn7N/sxhhxGnQXVBxC7uL89xcxShWHeJkYn/buTHNec6J5GjmZrGG9tBMH52X
K7wXaBmiUg3Y6pd34eMB3gvn6j+CLAzVt4Byvk7ekAMBJm3GsYd5n9kjKa4oDtD0
DiBYEwlNdSF3slI88DwB0Bk2jDziq+ul6qd07YxO5Oy0/X47BIA8rt6PgFyJwET0
ryzMrxYJFy2ImPNcNouDNF241kmffNO//ugBImLF+kItsdKoqLLZcFs6FfD3Vo5/
bj5/MWLWFDDhBz7Hu72cZTstwPNFBrLkBeJupazz93Zw/3caadjCysySWWIVHk+F
D4IoeCdWjqVhmkwEjbimC2bwtMmJ873iiAP1KPDk9hRyRPge4ZoXMdmZYxKhOIhs
6mR3Ue+Wc39SP6YZI5pntK+FXpnbXXa60EzJPnC47tAIe5R6cvv+r38TDU4hD8gG
jl3KTyAQsOQbeO1xIa3rlLN6tN/Cwttm8/zSqeXFx8IQQ1cGRkkbsjxi185ray/p
A/10XSyPm3/uIzmCggMDkzE2x0vk09BgJ/HpkixuU3I9cseCrY5QuwxZLv4emMor
cumr3NCOhyQGsq8syyQS5CBXVvYe3IWQMgwVJMidMiV6+nD/ywCLMDfgiLL0vubU
a65eEc8k+iwyDDi5EtZuUawnhZfDhL+5ocUcWHoJq+9QW7r0qlSIonsxLPsEr/X+
Hco0+TncRJ/BlcOEt8LxDzhx9IihMHFlVDGxAEmJIh/+qVnYyPNRYec06FnMo2BM
S5e4c/Q6pNSJSOiUpRFh1uhe6rVyph93XMxm6EynHJGNHRdZ3oxHW1fM4RAJqezq
kjwzt9g2V9O0dVh8cssvoq87zpDcV6JrNRjPOduUAPVrvMjMDxrzNeKpazU58bR4
ut/xMvJDQweTN1Z9mWUhHDjpcXlsPsYxbU6nq29bhM25fe3Ju8C/Ip8flVs+PZt2
GxoFKTO7DLZklte+kp1lxA==
`protect END_PROTECTED
