`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+53lr2yvIL4xLJFypaf4nh/OfZg4W0Bi7FaZ8yV4NWEwuwRa5gEu6yZdxwezNLyA
Vc7dQeoA5r9oIArtP0hGfEIXTqFbce1eI4GbT2CdTjd4jJcJpUJ80cnm5Dhb6nq+
RE9smYDrH4t0F/tjcOEL5JpbRDoMwoKwwOBacRD11U1wsyjfeAqMLalf5HWSRW3f
7/7offTQzDzpaocxdnoZZOmBKwS7UvYwzJj+mNwIaJx0UXCNf60Jy5GHYfcZeFyU
qQvAPSQbyvMGns/sPLecz01Voa6v2FB5xB0wPo55UCZl/2RfDuGJQP0JOMYddyYc
eVr/BlpKB8nhiZhJj0do83NFcp6QYevXhNbKaTLdB4t2ihcXBzXiiviy5wR4MB7v
8RBgpuAtkIhaPRTlauFIHdBzE496myvdV/yIPWNLly07CEtxsuCeGr/BPQ3PIu5X
TpECy9uzFIzDkiwrvvd/j/o3oldYqeqtpm8u8uBrBdVmlCtkZ+CXYCb5gsY0qBrd
xSJ6zbH29mPuWE4SUvifxzl8D0AbhTgENkQOC3c1Ysx4vHrvIwwcAJ3/MkppLdDr
PkG5oeACfnMnNt54ZN8LChcCpuv1nDmcrIrQQSN22LsJn8yF/gnXCyA9AUiLduE8
dfOdEDqbVkmCHrf5AthNPEQkID1jWORB3/vItWpK1eg5HS9Sl3V6QG/EnvdUCm/x
pqtyYE/kYs6NQii186R+7UGbWlyBNGx3wIs8K8wNHVlugAzrI+PFNKEKOuiCTLDT
CSNAjfge/9a0+MHf+D3gHDVq3PUMUTjJ+ZXA9Eo+LNiSDbTMdPtIYDYtW0nXi2tu
NuzgeGimzwq/htEFlxro6bo183kp88m/9IGGb1EwiLjaINaB2DyvTcCyH8nntZVY
RI97e+wFPIsgvwsU8WuOeHAgGpXFG//le2fdN9GOEWCWhsE3CP/2jSMbIC4oP601
OiPQrm6xTtyvCaWrg8Ry5LOEbCtMqrsKfuoHRGVnHLMP6rw/PEsmklzIQ9JAyiA6
8+m2H30gtlUMRZySBYwhpOR1xPhFTUpMBfNHywAdRG2YweXxkzEi5Dpxz1Y0/Nj6
JrzSk89cobtboIJ40wQq8Og0nQwzg10elMVW83XQhp57E2v2EgE7Nrlu60nQVmPB
u5fE9Y1FZNoRQQwEXyuqDqgaX4q+8eUQ8zPE027Ok4r/wTtxyGwZ990m4nH4KdMN
5gH0wbN10eKm+V0dHwqcBdEHBJUAds/EzVDPBXCU6LnciG0XUKbpMtOjW8qyBktb
+7Phq2JE0GB9if7rFKeUENBq5wcPJxi2ScVEs17ktyQDpBh3LCW1AZb9D0Cj4GG5
P9MmYkKuvPd/sAE4MYOtjQ==
`protect END_PROTECTED
