`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
u7LvTSj//HgHum5Om30n1LGgDLqhbXOwTFePk6jxqcUBgDPoHrcdw+KZu+/aRHEN
JtB4R6zu4l3RGlheLGHzv4EJ1Np71FYMGOSEgBfM3RmNlOiFLXpK3+ZV6N7OLlmi
+6fkIw+hfzdhHSk7VeRdfTRZ/Q/xj4jCoI3FII5HWZ+drgmLMC3U+NIGcY9LkKEA
vrOZwe+IxuS1aPYECFAnM+6q3e3AlEUumBFiZmIrI+bSda7aBJizq0ECEchjgJoJ
bKzUk5UEJc+etzFhmUlNsA0v9sUiD0bbeihAW+Arq1ZZ33GDgxG69xovmeLjZDXx
sgOLI5GF5pe/DZ+7cnMelRdpEzyWAk7GalGOTmRBIdJ1Y+LJieqiGfXzgBmFfIxS
D3lMIN2h3dA5kbHwqxsPsxe2adedDkIP9xx8aML7ax6KCPqHqsnY7Ne5At/EKca2
ZXu5avHkzVpDgGhUe73HGlnWaMb55ElVSYj+UkjEbjmSw9OBgKVneIavJmFUCxCh
MSV3HvSnE1sqOQnIfS64Kh6zBUq+K61U4ilCxN9ce9ZSdXw59tT3iT5POSm2BMcX
IrSLnz20PmLk7w2jfaIJETfde/30x2qxpM1VXWLG2wb1hryUyfC1UIWOE/F2h3Vj
5rTrBjJ8Bh4o92e8ckMDSCkxxC3A2sM9yQK7UVClnKo8Uyi18cULlwzDiwDpjf1A
zyuombWhKaKrLVlOTzZjp3BBpShUusQRvIs4z4QSLpiJj5yKZV4w9THI8jWGE0ED
JPIHA2NErKUg4PxafQrP8bKlP0asxBfpSFrPSBuuXV5OWc2SSP5IQT8GoZJGZCqM
E0mHeigMd4t5qTb/CiXAKe2CkuNmWz6Lw4cUgtbZRPHVln78qVMyWI6nKqEnbMYh
cz8L48U6Hm94RohTszMbuLMscU8CoRcYdqL4E42uy0EgP3ol1uvQZQO3qru9W7U9
sVURanVjCXwgroY+WQOpyetvufH3Sf04miWjw0NeyOwuoWR8nyfM54Ph0r5fhguQ
zFWlBb/HK3e7y3U1IYmY6V0T0U9XrssfTxVZiRKeQm0Z1D19dP/oAsF6creE2vvi
PcFJbhuANCowkifd9EwWU/ZtIdQn+GFdf6fJGAzaN9FKuot8EbLKnU2OR7kBFJ98
NBLIOGPKPE/RQjai9omq22Uq7IiAaID5IkleFVaq6z/0v4GFbSko2Pa3VGlw125L
txVYexBhg45GkGDnlVM+boBa5isTJ5CYyLmXr3+ESr6KJb53OxnB3jOAxuDtYzfp
8T3YnTgBEiX7m4g1GvhzIEVBL+j/DmHxu2uCM5KCgOt6kz48CuMXcvg4xirmntFs
W8G7OTDrs8PhxaCxw21WI08mU2eCER2+CPSEHCKZbfzeRTCuFrMQabOITZwPebWG
+t7ZQyesyvpjl5Ozb+vvW1KP0KgwXCE6tYsoMmpdT5vv9ggNZLL7F1hlFZqtzq9g
135niMbZ0BsOjPgLf0Fpwhw5iwdxnQEELv7JtBM/phlNcBS2WQ+4WpKqP4ngTkJz
zSg5GAQk43QPxkAi3vegPxd1XWKzTH+VLe0u28uqs5oSDG85icjI1+O8BKgozQR2
rPdtfhY4JgbtQ4+nfiejBTUQnIMRzlTOY1i3u8XO46yht6wDSAU44SXg0qN0AC8G
1OwZJErGCapP2HGxwfd3ECms0wCqOXsefU5SonfBpyeFl20zFEpr7GV98ERd2eJp
/9XcQriji6Ggyqf92z8sdWxaFgA23QxrJFfRfnBoa5ycMcdhsQ9mzWhN45IV8pa/
OP8Qt9La2sOLNsa0oDumWBFsft58Q2sO4PVDMv36yk0o9g2bOfpVg5SpGUHoiAGZ
JGm8wY3bXoV4DEr9Iwp0y/9GNfWjxal0T+0FtvWXOR8DYo937roeBqStN1YqIuLv
Y1W6zULkdshzxKQ8U5cMrFIEbSZHLC24bM6kt653Ixx2E6gAVu6UQBbwc3k8qk3C
ejMQG6ruApEo7UMfR9bMaMe0JGlWpWrVJQPas75ais4ZGbwrIzW6ZI387PRt2H+S
tPzy6f3WUblyw7E0iG5ENeZNgjrx06WoorOsTQKibs7bkFo4/bIZEPmaL7ljsFKx
mjkvtGfZ2WrMkTmpZDSIlF/KJFnnWfrOP/Qhzh7mCOkgMcIsgL2eODdq2nqx0Gqd
0mCDgXp/HoL3xRWxur1PZ7RbDJYQw61Fh9XgwswjKTeBfbTi0eGsNfOIv2sepcvE
szOsh8GmEu4R6nluBx7Nmth5m2jF3vM/NfLdCdc03Z3xxF2qiHF+w8lGA7VSZzsR
mbK6QAgX2E1tcx0owP86ZznoWXDIRh245gjhOs2dDuMLE6CshJ0tJcaEOr0deg26
QH260X128ie9kGLiR8RYoiEmcbCxmoMTP4Vm8QzMqJU48YbBkewGyvhBwvAiwAC5
jNcEFi2lub9OLg/ovBQwn1yVaydwkIHKbwoJy6B/2kVc+PQ8SHNrBaAAoA5XPc7p
celetYV6U8w0a/M1FALatS7BNUeKh7tA+H0bRNmqvjB4wHsWsoZE/lnEY9m2Upem
DvA39CWE2q9NO9dd7NwrGGxjLxI3UsRXiQp6hTpOV0UFuLei4WtASypB8kOmyb3h
iijz/OnQLb50TcoKi25rvGa2XaVAwO7MAYGrqgMDl8JJsXAzgPQsY0NNzbebBEII
i+3wknrglXWepDqxErwd45xipdU5uv6j5pwM02M4LqI0MECxX+qEAGiOGuEHbk0W
aDDqf10UahPJHx3lYz/bLhXVBXVI69yMR66ZDPrcf3JXXwhngc2NIumbLGvMQi8C
l9ml4FsbhNhChtVh5Fsmre3lQ+E96ZdHjXMq1EwvzOkRtGTjrYGvm1TLB102ZLL6
aCOFykZUGMA2Q14lr+yN6iGnYZGzWoB5rNcrZYOIq1mLtcIERRmUltNChm8I+7bp
jav7GNjoIpe91r39xNy32R6Nu+q1OuzNtyIopn5+iSL/ZqZ+CdNyGskNBNalFmbI
k+2Wn0q6OcPHwU+ZkzSlJ0jV+7NgOVfyGJVl2farGaRvZsK/eMcDeNLeTmnnT5YK
sFzebwOE4J7Es3V5A4PcnO8FTLh0RjNDN621KOlMvhTJIBQQQ397sq9LcTVF4TfJ
UjfR9BAZSZ7fPGJjO/vwZr/rwkxTZPVF9ERi2rq/XpAdpf2svcojEDFQ4YiH7Cs+
Xx3DWCbVfxiCkcPliYOzcPEIGmxuTnJb1+p85Vn9kTiILesA27g0mbeuISgWGuP2
teZ1gbWUmTOipdUOpZAr40XJkz1FERh6R0YujXDy1D0TDxxZM0Zi0T3dTV9MaTJW
erdgdbDdT2SGmz11M/QRnWXwiXYYKQExTpy8eW2HC+yHSKzuvJZl1a+zCJjTeIZh
7aXAuY/X7mQ07maKq+Ylf8+00MLnH5Kzg0PDCzHBaTiI4t6W8qnwq6oH69DxQtaR
co85k7ujmjekK6ZIEAsGCJ0nkMR+DnqJzEQ8EoeUWuU7KEYjFOPngw+5lvw0j8Q9
g+FmQCZMYNbci1u0lb7tZXEHpxSFH7rGbNp+KzVKTPE0/LfOcob49dbBOc4U9pz8
IJJw0N2P0YpNOE/SpmCyM+WoCj0SjTuIBQTRlguu8vw3WQfBsyGvGJEZhFDDvZpp
Yq2VHyruvq4oGgttt7E+9Kp8snzRyauHiPGeDCgzHiKsRZiH9sRwlZYXnPVf0RC6
0Lfraq9NIH5nbwWvBk07S7NYv3l2ZmjSI8YwJaOVr7dvHWUL/fF2ZBtjCJ4J06mQ
dMCkRRs4B2BqZtH3n3i6AN9tusgNcPx1O2yjSunExjradMrrCFtRLPFqGCH5Vc3L
RyYNJAYGtcNYJlgUW2F8gA==
`protect END_PROTECTED
