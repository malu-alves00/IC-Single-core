`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1yOrs3hlQNOJm5QWh0Pk+YyWFe3sxd8hgT8GWwP+xY4X9pym/irSLmdw7SFJTBKn
//xkNleIjE2hdD6BWeW1MNMg5kNVjpSZlkZzHqiYOiabK9egm0oz6iBy2Uhnos2r
x9y2TEUd2p/WbbyR1PWcv735enD8cPUMuGKL0x707JXRxEy/cM1S79RgCgdXuwVv
Zoea1Bdkg6C7Pe3rmvHqJb9D1+dRpsXcyOAh/muog2KF9x+jFECZ+Q3zyrT14IWh
GBPKB4zNC1q9TEkflcvIGJmX5mfgyv9U2mZGGkXKL4J/mZAhWNlQtELZcb86lOwg
teO8uYAjhE4OaDPK/dH3p+UeTl0bNQcyFRTK8EunldEeo0k3t4Ptn4IuLoIpj+VU
MCy58trbQmTYoj7SH4mJ3aLrZ920AaBifjo8qUPgZGKF+gIJSchHojlARhXBwwGZ
cv76TsGmqyi0WEzZTXxiw+TwegYKfyAihfaHHJ2eCu9H1S94++HKaPiUUZjyID6L
ef3Q0ulGY0qw2MbyfrxEknCm+ho6vLh2Or5jrlezsNJyA2M+kaHFyhnRtH4g+O76
/cbZEVSRAqegyjvTgAiciXPAbPAO3x+OzfZJqlJyGyW+ars9zeKSU5v7fu8THnSs
WnE/LRXsUjFNBS6fJiDS4GvQwWf5OAoBZydLPh/yYaZLtR/cgyKAvTMMNN73vKJv
d8fFjg1ij5jov+yt0yecZzYTi98Fnovk/YY24OxesOwie/vuq5jdlQQ1oMSUkJMw
wvxRsblPWlyKvxV45acrgyMbE386xqG2/6VMHl9WQLAwblozhnaq+1RTmTxpmqz3
nfgbHWJ9Z2ni8f/fIRCUh1wxCkgWyz12AS1yjE+uth9dHFwv8QWt6dRa3Mz48oR8
`protect END_PROTECTED
