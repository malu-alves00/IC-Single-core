`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4uCKpFepIAaoXJGQL89oKr1ZYDAvCJ/QhKSQRfff+Ykq6MTQHFuTFWPGDKp2c6DH
MHh6urYEbq7u8QZiZLvMB8woi2S+iFjm0gv+b+keQzcrUcwRZ7O3A0nxFEqwrCty
P0qYHRIBszy2U5Ot4LGQfaavxJuJb1XPnyEANZ8aJjs/9TivE7rzbKp7t4HbvfbC
wVhc7agiOZ05uHk4jyKUiKWSgowri/GIspTxXRQqd7LaheDaWhuZ4Ytv3UmpAaO6
tX2N7hH9DoarLdIZguKQjI47Yf8fHRXwQNS//c3ZO52Lcf6MoNWRiQw+hB+JQ9RZ
c7+CgcgmdFJw+p6mVsfTYs1BL4/NleSZf8xeIFeV7G10wN8Z0UmiEzApqV/3FikH
pcFM4PUCPhhca8VNJ/gvu3qhZFSe7BNwwX2zVeB5F9kr9VsPj29DQBf0q+qSKvLs
oC9C8pNxAkZ01nQuCWaOZswJiJWfmDXPHyctY3R5ievmrXerg530HIFHUbzydctT
r61X3v9YMSBG+wQ+Dg+ZyVpERCqH4ZHTd0aR45OdWx+1bByr3WuDZsFph43FXhYo
LtiT4DYvEgrCCN+mwLW9REacXKfdoej8EDvB7tdCnhNuuYWsRdtdWfYBVfsW8/Pz
HzcdDvmJIHLx0f5EKQcvp+JZyCynDbpJZTESFAhhC+kIjy+0nV5+yqsQmbvkpXd6
mbFpHtFN9Yc+1my6n7mgkUXb9EA9q3vtZaa4XwNNBDw=
`protect END_PROTECTED
