`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8LvlitAkFI91DAUnE1qDeRYNf2/OHU5FjUfGAcMvxAwp6lQcehsAQhiJpHseTaZX
1Lg9H8t4dpzG0F7P72DKdGTq+Y+orm9U5SILpvrYaurdTcpXmoIgc/1RoUZVzxGe
PmoJ/fwXiBwPmHWqYxjHcw3JvDRgtL2dSJyV5qsPIl21VjJgOCXYatllqpjZvYMH
V5YTBG6kZuMkFisEN3IoqpCj08EBhnKYPYAgAJQ/+EO7mbJd1vzdWJrBDUiSTKNg
/vnRC8p8W12ytXPZj3X++plfqzFbgb5gbxYYeR/LHda2bek6k+ni5PrmbciIK2bi
eHiSox65yfn8+T3daKtddO0wD4Uni9tlA06HbiIYWI8fzzjatMjL6SFnHPIZO6OA
hRMknSn2yl1nWvtU1h8xGAcl5tRpkkpsWHYt70pbDBV5WciPkiyy74v+jAmUrctv
BlddzkwQ1EBh32bm0WlKuK8z3D+ruJqMNPZVQy1tv6oQyD6OSfJLYZ8ylWVoFEkb
KfKgJDKkZV44IvT31Cpyy6bRohPNe5RcFclTPsHxQ1WE1McQFaUja8xnDIn2oWUV
GLhuvN4niFxPUr1Iqp2pO6gFOr97yaAdveKTpj13PkQDs731ueF1MXn97nnHlwXh
4du4TcEvv+BaQ0ertlj9wK1EzRRbR90DtrD8Vb8ucn9jMD24cF22trKVNxRcpHnC
o4LLqNi/qDMZUaWrwCCxP4YM3FXiADcIyvf75W/QcjgQnsXmoMjpwuOmc1ZUjWeC
WfCtUfbOrziLGTyDsSHuZtUSGUj9+dQ8fC87+3Xr20eNPmFew2GZGAweQgxWEEAW
/RmFi/OcwetxZi7SY04jH3BOlvKxnZqYS0F9hQipFUnHXu+oaT2hBvz/6ePh0qJn
lnQFE9xsR1p2qGLF/fNYkPFylSo45n+r4+g66ZiR+0ICLa7cK2rOyJ2VY3ym1mIQ
kM2NariHos81K2GLq6u3fO6puy+4dWCLiqXfwtgm6TqdiZiQkOUNWinmi/fCFLE+
p0zVyxNK6G5YDx9MZAa/IAsdR2wHnbqOjuv4PVd76UAmNLXFLkrt8BTy2jzlSbMx
n9nIIZaEZmRJf9wKo6Z0QE6YBJpcSd+wd+HWDd7m5wJN/CviMmhdHvn1MzYQY5Ab
Tww7FJ39rmt/jDyMaEcs7wHJBeehCAy1uquPJ7Bqto98lvEJXnn8Ipq9/5osbW2V
1ep8spuAuXx5JtpGX3GAsnUTywXtFViNnZuFtMCi5gyAEYKlmaql96eAXLQCFT86
srnfj21lj+8C8rt1vZc2TPl7roWdviHf8oeRTB3ifXQ/e4tUFKsJZvdTeboUrN86
1PEHhVdEc4UaBucMeOHod9GpZ9cdSOVBbsoCzYr1OezlZUsGYlmsIVxfD3wzRPRQ
eOzjH8EBI+tRZX6CnymMu4JSPyDGH9TCVUJBfT/e/TMKX3E+v7G+eqwI2VJUVvpM
Uw2vaMnyoUNYvju+BYGbBN+ie15qCduUq4H79A9SjoqDuUEi5HBhlk7ThtY1AXJW
oCxa63Ea+JeImF5W6hvaSGzxlMXWbwg3r/KWmT859Ok7O+1qMGb0BPCcFYQ0KcCh
tqDrWMFGoNm5iZU4oY7eReaPaayFCTd0Wmj2kDcRQGIhmsHIVqYt9SsgQhR7L2l8
JPf3eztHfq+RBU0hfuZhXSEbTPXUs+Es9QoA1PGei63T7wWWw/fDWNkGoVKf6nxV
zK3Nx0zD0Aok+rhoyGI5Dh5Y2CMFwRcSN/5sjfeR0UTLZpBVhy+D1Sx8uqmK4kGN
URgcdz95RWnDiBfDZ18RqfxySEB6FJHAnlU09dC/c42tgRRmoxgPE32eVaijSOi9
Lb1sEYr8xpwZ0e/mChEe6/G/GGRgJr+dEQ2O/sf/jw4fH1SWKzNXipdWGGzPKZkD
rq8hR5lSdEbLpbFr2EIrvnhF1S0AIcDjMDrLEU65NyHYsq46u9OLv1LwGIqFzR5q
BRDTfoAkh+HkW+4KQJtZdGMGGSjok96hn8CNgGa3ETsD9w2uliU6q2mwrXKt4gd5
wsrUgKC0euPzxyna4oVW8GZsTke1xlDbsrfc6Hhdu85az+I2T+O9wCVBZcgdiRwU
VFE7bJJzLilOIE2zXIO1A7Nd46ETKysYTDabgh4lcnNkUDx4tZin1XheJdcbGv+9
BRXnujMvlGm6FkaK8J7sv4WKMIC21J1O3RsfQ6B9D54RwwGjoUPxNkPUtJtw/wO6
YTywbuFgVyjaqng+GLo5B6bnOPC8feq4rX8GitVUWUGhO8R4TESgGWbDnlUpTUvJ
TC9x3mSlc+l8DB0DHBFNHqpqalR7AEfx2qYtDZX0HEytHOGAKHcAWchx2zaLolXY
mtSoslLobKzomCapxKUG26dJoGEsrTBUpw8oOZ4p3eZFo46obkZdqHJk0fQTpmpS
7CV2ZVocr4BgMHdYRX+8KhtdOnfSpTNhlw5iMwb39o+0QYZyDKJKi40PN3k+fEa4
zuxz2c2qJ2qhHsEqha4gWEuwQgvmzN+t3lpwBJXUNpuNnyysX1J1huFbJe49D1jE
vSq9e0U5e/EJ9MeDtKvoHwdqeHmetrnbKitTu6+Gq1v/3lwc/7FzwFHPyR29W9KO
y/c7ioWuThoDM3y2vceAzunJFwerBW2uO3N+ajC25IOg1jfLyGKlAOGwJoqw6pfl
fAcm5xbu4DVguFhSlH3Ea4y0u1LT9WHB+QP2Wl7VOZBHSPYoCAz1M+wly0/6DBit
6J8rgCihiCdVyLTpQxaFRAeNgt2XPHfmsGXG16SCn2nybMtnTbzc35i1IIHCuQ5Q
tifgm165ARGuGvY78VI/8nASdk5kzXCifLO9iUobqnmaGNQETKecJoMH9YNzdwxs
P2eQMQRywuofZHYh/0DglVoLxvTq0odZJKYaypyAls02oH9mHxQB3hXyoLmdc3w3
rHLyq2vvVILiIVKAJByJxL3gpv5B60xMUP36U2RxyxREpgBWRHGR1U+Qcvtyiqm8
EaUDDESouc5TRsxRT539SDSQ68ubvJz75I3xqp4GPwGZLxYYCcjyiN4wV0Vy0y2g
YTbzlF/Wdr3HLld3ipMiA34sdoC9VMGRfLHTzsSmYd3IY4gmFqX0i8ck+WQz/JN6
EOZ1s2HkyMrRucmVrO102qjM298P4FaE9ceC1gpMz8G/pytDPgQiMIkceIJanUVh
18xckV4jISShS7wDUs+B1Gn3VLaW9n2fDQx0tQIdW6cbYBbQCe4ZnOeZT+bzuaL0
wEZMiInMGRRZGclrVhQ5Tqqv6/Fac+4mBuvs7QaEC0Z7OA6YZGf41o09YAwyNysH
49uQhQYtpsoGZIVuKet+7cGJWPBYIyVsuJbgjKmqpOiRy95MCY88opkVWYrcjCeH
lHvHq76FIkrHsUHalyQTRh6oSViR98H3QOnKXchwysUJ2pBNXVXQFFjWVzoOp03Y
gUUYmj0/0aeqF0i4X3hXzCS1MJj2p5MPJpVl+TlqpM8qkX4mTU9VBiUo4+B+oqVf
mv7l+RrjZ7N8WaESgBKMvGY+DjGLkg8eYsW9hid0lI0qh8k7b4BLb6BeDOwKZioH
YkT7yLYQswIDxSW6L6p4ASnmnA2/dheZy5bKnLP4D+Q3uQDtltHDiSwH+m1mGvzO
GiQskSjtLklO7W/RJPcD2FHagHLZ9ws1q9zNFbKC/rImNToaleMK7+KyOBO6J28k
iiAyKN+TUq/2vHOshxwBvMIgWmWUxfa5be191HXFeP1BPBcgpHtSE2vPZ/2Dejfb
BLn3zAHyXnowuGaapHJrlCxc3tohT51DR8RKNaRGwxStaqImVr2LIVbRu5xapV5/
ID5P4dngUdM38LiLni53Sk6kKdwBbO9BPZTKHYBlpE530b1ba6XiAFpG1+DdWon6
OPHhFQbGiDBwz61JngGG4CAMdOKjiuBuIgqvNd0RsBbwvPMlALObtGpCnojTgZbP
4d37O0qTxdBXGsqpAbti5DZFUHGdKx2yuU8NFVm1Cqxs9tppnvRWN3mNGZPYU2n4
jU7Rx3SFr6aYhoNiIqxxW1RJ9Ux67XH/3NSX9pqY3NHsi4iaNYt9/0TMhHF29CvN
qHbJaNAKuy+G/c4pcTSU90MkaOVztXLxD/nn9E3nSHd7QG0dj30C2nHpOSCRM4km
t//jn0AvscAk25DlKCrg6uxgibz1XIK+vQQn1tmeZoQycScZmETwdtf75sdaLsXd
0Gf8yFnIFfq882BSli/3jZS+RL2HVFic0NFEg2/i6zoEPtn0H06JbkY6Kpeqxt6z
Dk3XzeOQMxK5oOrrrmeo2k/BlBFIL4SKG3hlWjOVb3sTg9WSmi0Kqr7wfYjvKihB
4p8xxIYZLMGmcHz+HT26cuDq/t4f8pBH21zYI9ZwSmE3zbIbTWvnGkqq5utOJfu4
Elf98LyL8IBxStkt2jOBSF6POxpklK1WfkxzCIlFOC5rFEbStmVZdz+XO3Wi6GdJ
OPVPOnBy+K7p8n6I5i19Wi+TGX1ZEK44Yiow0IACNk+PEdEB7ArToB1tV+VMYCK7
LVx6M5M089axHi1H3jr8VXhlwz9rDVwF7uhgdZYTosgWErPEo3H2SXSAQw0z3hz1
s8jtRgEz/5CdiR2eVWJuik7z1vRZ61XV89GujJr1fVVinNWKUJgAhlDh4MCIIUpd
LbaX5LAqObg6rB6qRPc/e+dE2O9L6MB93IO1fwizwQ4ACWXvNt6dl16PxqA4q7wm
53t/G+ynea+PSddbb7w0aLFw62GcuPDI4EJTNHUYMAmxmFN3CcEABYjXSszuPqtj
6ZPIJASj6ZlGE93zZ4Q8l7ZjK8Cied7ykZNvxCsKf99S+hhfoKs7dFs3p9w1ol/Z
VIFc1bdqVnItLHdP+xKVMikzMWPr3mxPm7eBKPn57ZdIT5373yN7b1z8nYXehB5L
ycDybeJkguPg8g582GYfHc3d/wNUQxd6p2Zn2AF302N+JCC+efZQd62FTjsDa4I5
LgClupCEbq5AX5vrcN7tK0PU8NaM1nWMhIfAzd/2iwsnmszfjjyZ6sSiOYq9ENMR
sQyKBvkEsIxTXdZEgvbmSzcWJqmalRGF6QvJ0Or8eTKpLTG2xq/fgpLAYzrzBF86
Yqo2lVoysL49z3UbTAxTU7SqCilnEPHZz517YTWZFG9Ii6sclRbc3+bXBPH3105G
g8S2C3JdOmUtn/lhKs4KUDNcspeeRX5zde86ACRmQPteewohFkyocvMW7P0YTtAP
IwLAGvFq6NZrs8J6rdogNAFEMzMJZS0C89A2mRBwy149uT8J88GG9GGD+IrdA8IE
Ze2Kv/63Gb16d8DCG1Ul0AF3m2iyhz0SV34ZkWy1yGQQYVMDQ30oA4U48UavGeZk
BhYTi9CkkjFYU+HZQxDF6shh6g1/9PSAwsr+TQJ1KI5nqHNbUx9gdWDDhBmVG07h
ZuR6limK9WdSHPHoT9oxTGyh65Hu6V3nhxYOJQoO448nykC/0G7ebJBqmlFhvliQ
oB+3TVBVp96DehfydPNl0/tEU3rh87tAhRkF4kTr3NeYCEmwl62xh26SNnnV9eh5
TY74gEDT/uMWJxl5g03QZt4o2eAiIEJI9IG0OluHyWOSZUHC/5CNRPcunCFIvusn
wnp/aWwuy8Q/wuhh79ATl5/XXfG6nG+qqnNewOSNXuIyFxMKgefv/eKOsT3UWtUB
qIxvgtnHki78HlRT9uJGHgCDJIeI7A96yuXAM7xhcQ4jeHGvKrCqvgNyNdymF/zx
4lbymzi1yfV32/nhahfEDRU4+jgVurr9lCbR9uBUt7mBeLPzCnH9L7CxEhHL1/H+
bumRCQ5RV8zkOVGQ90BMIKHVHS7oyErQghbDRerWjP7PpIIH4VSVT29XGW+HzOcF
SFKj7y1We+ENvt4grliX4grqd28MNEhcIU158nHx/iC1CuF/+tbtMOM4JWt21TKV
M83MkEsDmXEa8Wq6ejLjUvEGvIJTsfhAzyfbZMrOxUJitbd7ZmYfuCFRFxx4i/+8
JDv8uvOVDcGh5zH3NkMIZowUhfE9AVyF+tGffgeNxLEGFlqKPSWmSRvtiqKsq7pU
RXBnr7zo6H1id/DouRK5wYBIT7o23axo9z1ExU4cXXZ4+5Rau+m2AObR4EJSzRx5
NUJKWpwh1Pc21LswYjaO5+fOdo1HBIULYVKGNQUpbrlt5B6+r6qqlAxWCXkCD/uw
YqkTaKG54DnFZIvJc9u/VutLyZ/cUBkrPZjHmiEICSP8X7Zo87S5PGamRkqNs8ix
p7e+jFehmrZG0iXyPdytdsO6olBqcugJ8/vS9BiNc9dcOQcY2eIg2cxkwXjhNRfS
EjrKx8Fhq2P9bsUT4hd7DWREfgzIzYMIBsex8fOc5AjwQInrCtsZssXSQdXbolMI
o2LJDoX6uSkI9sTTe1RJc+HYSHeRtXqhj4mSweSgQmpTpxePWR3r08znnNlVI+rS
aOyc0hCQUeMjx8Yi49GRDZ+1PUWM79u6aXdHlIu/06BdfGXDWQWIIsHZdlw6BTqW
4JQeZs+hD5QhxqeTEmKijtoFNLimpX0bFMLBFKXMfyShSSADE3zPTcwumHn2N49E
JGJLGhfhjnIy0e9y7QYZY0CkTAe0JibMYhrruQmWXTTDo2q5i0/hGlpgsAVlT89z
V5Fm4StPsjc8RJvwgkWKCXOY2v3i2Oryy1RU8eAZNBXUlqopENIXcfNPZqsYSqvB
nSLDCBDpc4Gkst3G70JBMDdn4qPB/eljL7Wm1IU5JkEgpEiW+78PypqSosi826vA
Pjfls9hwFyQ50/5+HHRHeEZT66gdRKmV+uCfPIOebZyIw66xLF/ttzuLh+G5fvl3
UZbcZuoCyx769RcoMhby/IpXn8ige0MDeIBUYOrU/ERVcqw8+vXLF4gcPqYTQaZN
//F/JmS9tV6rotPlga659VSEr3TqRuNEcVcfU0PWh3mdm+QF3uKe5mMBALRaC/wL
5lHB58gG7zYX28OsTfgSnGw6vMroFFftS463BBSYFyTMESqGeu8AlE5IlM7f7j32
+/llMzuC9Fin08P1BPAheOZm825qyUuPg1/GnTavld1s/z1fNyfGgOtrqHJpIEeK
WRhzV2Qos/5uthEYTetj/JOaFgOXqeJIQXx3X8AcSOBxaC1Ct+ktaQMxEXNesc9w
a8UDUdXr2bE08QxP9YXbyOeqJuUjp5HGfw4+tgZSIr0wZqLkJ2lTOxETYxPklbC1
7HaBTZuGl3CX92ROIeYfw+CxL+DBi01pIbCyzyS85cZDYB837zkjCHPjsvr9asjZ
gzhPMB69AqdqEHRHxGwXU+w2DmMu09pVTpS2rHhsXY4SrJs9G+mOxdzWN9nes4tm
8BASQw7KtO+SKdrAYbM86rIuNO3JyaJQtXDoOxX36kDnsGVoC01MA5GYHuHsxZTa
NmCRaNKze7COXNvFEOAEoTPwrXvsZXHqv9KtS2ENY5frdxY69yX1xOuXcbqGkBgc
V/mdpviix3gC/KcRihzVfTv2nvsXjlbAKaE0AELnwn4wj6NIZSIn2pZQ6c6+xAfK
XYgwSJ+bW01VbmY37MNjhzP2SzvbNNO1kTqBc5U8+DrHZ5x/sp13Iz5vxLVKO3V9
klcNWg2mxUdhhaoNgq1LcgP5u4ndXcsVjWDZiH4e01cGTerfBLkj9NttTPAipvbM
2YjgexEsBdb3vY3OoTDEj07k8LWyY7guxGfrScqYwq/YWyeIu7BzsNma9taDdNEf
76xajl+R3y4DzAOGCsq4CFCiMXFaWR8ShMOTzkpC08RcWziluzLmXlWZYuLKTVpx
s041xmI/yFhmIOlCoQliTLQJqiNc1fKK0TErfiPN5uC/a5wuPFLbZOAljvc4I6di
Y/OA/PkNBZWMon1yvyg/GDvFOpKLJTwZkmUF+omvBzRcEiV4IyxWMuLKR3XbdRWN
MzulicVI+ZQzF/lL/z7Z/Z0G5v/zHJw/TCLMRN4VOAQfw2bn/roNPk3qPD5qlYFe
NnoCPfpOrJ8vPp4IQk2cskmE/zKdHhIHaqgbf+R5NIM29enbk8jFZxA9Zo/gHlRn
r0Hk+G4X1/RGK5iIze8L7MTlUVkzqrL/B4jdeXLI9BDBSfP1lX3m4SuqXhtU4Oqz
0ggi9+o9vDsOYfWRT4VWVAHWvVv78C79ieozl90nkL1NjtvLXec6dbueiYGHV9Or
YA/gc9dps4JDOvN2SRh6angzPUs5UrxkctG8lBHxzYKxQe9uzlALcZLJks10y7nt
ypp2JnqiIN2gV9aq981Caadr0qfVI8hwg8wINwvH26qABF8KQ2gbGWl01QNu4ZyG
yGPNzPaBjNgtEsbqusHbtmEerhhFc0kbCnMVBQr6bReL/T21OOWRWHZvACknhhqN
DttmMt5/4GPHZIfzyV+tzFFMg8EGGNVBeYqT/KTmXgqRFBsp4xHb9dZuKlmqGXCT
Mr0/onABp4BJBVebYuE6F5cUC9Ks7ATmAwEOyk3SaUqSHHxCeWRLZL074wRxjmrB
gFET35cUCIHJAnwhTOsf+AtDSoA9zXQl6z0crKqLH+kSwd+yriYzyBSVgV/+7pIO
dAy/1Py8gJdAJEj+kyrc1PsqxrC3Z4fqh3tIiKrddXIZUq3jdEAta9oZ4ZakU3nU
50RgwK2B9ZIGoMwsDYu4RLByrMbYRdOTRORyB7b85Q9JkBhx2PnT4vYUI0197jgF
YlhlgdmcUqtriar2gZaz2dVMmiYKe5GlwZuO62KXXTKNh/14U1x9oJzxwpyrQuRY
oeDOLHxzcPy3FUXuPgqJa0irO7y5YyE5yNM9Pux7HPDiQOhEK8YnXED7960WZXfG
7vAOjom5V3QPjY/X86Pjgx4n7rd3B8FaxrodWTLefaXOJBAV+/znFJoN0Ljc8gwz
jsgPyRi8VHznjrISNFOqucNKvnV6msLwos3oJ4Bina8T3DzyJf6fM49qXk0/YBqK
DnHG0BLkAgoYtjwq/t0Nzmqov6OIRZcgMCquLgHWEd7Rtx5UbZ0JU2d5C+bP3y19
pZ/gQSkOuzNZB0LNxM3vOdLHOHjUjaE9Wf9d2gSP5Zvawiv9xYPGF1NNx4beWn3I
ZK1y/FjabfZEHaUQKRImoa/TefbGU+SnaM6+aaDai6MAA7VLqsJVEgEuKAXGD6ez
zyPLhd3IKN+3GiqPjHYlp68EhPuf8eyM8ngXCyVpU2w9vacYQrAPU3ijMu893wGe
fOlUye0gOWmEZ2Tq3JzyV0gSSlBFMojrf/TAFChPT6uymW65KaLMMcX2TwiHjuty
pyhDr7Sjpj8BEUXL3qsdFcoAVA1Qy4ILG6k1sTchZ5JriN17dKpIyp1xP96tpE8A
PgPRgRZ77XfkIvsdjEXjlXjXMqtZsiYo642+iYWxW9VpbPUUEj9TrIYlIYsjJs+j
fLcZgy9Vm1GkeLFPuJUfArCy8OnZOzb3ACWgGqKJllHBy43IHF2D0dqGQaA9wLxq
6VHtTGEgdRsIWQuGxyt480YvdmrVhzpBidgpSaq5EKuXzLu4EIHxsSI0QW1hj1FM
eKUAkfQ11pLthNo3hGgXAkazxn3QBvGgkweyFK3ESA14DRazjppFhyfB4M3CLqPV
OvSvj8rJ/ms8dU0u7GMjyvS2AsZGBaFJ0nJCRSFKrvDZZ47scAEfAbxa4g663zMq
df4j7z2zRc4w2i1Nd8VJiQ0FcoB3KwlYq7oLy4yYMJGehVJKZ3aWSBQA4pcCvvU6
f2DNMN86inxkG6hvHr34WFvvFovPTUp9epLZrgKl0tzFkcf28ejJjL0H/2e2UAph
0eoXxW/YA3mlh9iGrJheZvZjomDUjb5ljdwucKIZmVroNOVcrV3mVmVVkKHvMIag
sQiDrp55EQNV1Nu+tuSr+vJWqOpFcaYv8iSAaSJKJO64lmf5YoD13C4skOorJBsN
ZiQ1LSC6rVSVmeI3srth3WEcJ9F5pTJYaOt5wYgVfmgf0HksONiU/kZnwccfE3J4
BvkBh1ECWatl2wpASA5AKZBLbL4YWOvpqLMTOWL9z0/e+n3KGNxyqZ6Zp695I0MH
IEYUNszj96sMzrx+5gvOZ+NFjeGTKlrLmZKisGyahR1BflZeELxkjaR+AQDmozu7
LNKfd0+ghQC9/t6jdmHsKoSodWJw1CgKhwS90nRZszlPxtok7Kryx+24ptWAeXT8
mWi2xnTKwb3EVuVCM4LOfBIBmjFFy/pe3/XJzjBFj8EslzEUEugTlR8C3X5KjN45
jZmX3bu296nO0McE01lYPSHjZfsJQgnYMyYiS3Q4J57TLmu1BnYuNgLrAylhnp2F
/lHuKMJKq8zB3yA3d3nG1RZFMTV9g2V1Q7ihHdz7DQIqeaMoABMzTnVJ2ecFVHMF
5MireZnRtFXvxFLvu07P1qfxV8jgfyYfCEvxIDcXIpIzGxeLzn3O9Qx7JRDx/69X
1SFI4NtRNf0Y/fIKaajAvfSojxizaX6797IAT8Qd1p4Gl4fZnlSRtMTFNazvYVJM
MJt0A8H1G/wWdaQIz4XoBb+CBVk9FipL+BBIJVtrf09fEUa8hDgJjYvXCYbn+KBo
JU5joVlQ1ZgJ0+EiiLOO9wr2dW9n4kyPirV+D/M4QlmEokPLizpISdWN44fDgLhd
ezx5Mi9zh5NMXy+EIY87buTfEuMST7C3UTrAqC+8kxgxvsXj3pd70vpqiH7vj2C3
wrcA68OM0RwUfoZKw5owm/DmAaTQc5qWJPmB4sDrXwxin2HWiM6ar6obACmipem3
BcM/z9L7yr3jIGDuMM+d1mNf7rJ2NAQpsylBcahSXhYDWOq6iP195GEByvraSe7P
KrOB+OA10L5qm7K6dMWC7PH0Su/67yCb85pruuA8YvPi7wWSaFXrsSjnB1KuFh+R
kjgVwn0cHz943zoeLUdCshpN3+eGd9fmGAXSfwa2bmy1gpKoTFNUdecMKh4tROA1
1LavWvJmKQBZIM3dTih04Ac7CdzB8IpIKFH4xIqCUjLo8ofb7NJma24TgLV+TEzm
ewkqvl0vMBbrmkFQRJDrxZAe+0QKJ0QyqT6tOQmG5eSY1cQk88WufSIGkTdct9ia
Hk9/ylaikzVRXJT2YlspyHSFoLuaOffkysLSIBXzVVidINpabNXamPFdLtVmby6P
o0xWMiIhFBeU9rfjwQE9rttMiXwWJzVwmen4gZM2oUI14MaiVtnvBeh7Rh/yWn08
drNoD24UfSNQ5qWUSvA3gToKa1ayueFh/9J2Xjw+wM6DX+7BFatNHXJo446Gsg/u
U19zusnSlZ1WuzSdIdAQpW84opP4MpggcL+686ane/g4iEcxpoOmzBZV35ujlunN
xkouGbJkNkD3a91QA7zKSZzgYsD1TtzsyAUy+aNjahHhZFUlYVXANosiw6MPPa3i
1jKq7TU6bJFJKeHb9yVlfgEFKO4Xh/6/CViTXiEMfaRjdhqys70+q3kdACyhLqi0
fmxjyvvaC4Q8e3XhsDXgm5hTRckxuAe42w2mxwNgFPHgd9LE5g147kntI+CcvJ/9
ZIB3iQQkoHECLKKNqNJ8hylbjXa+0pVzR1HnZNy7YfP/tjZ/zwO2WSlLgq/Xscic
gkXJ+m2liZ071WEQb9CtFPNKldiBhULpZUeNoZ2Wxgcbr/b7gNfmAvtifpig6NDg
kKFIERlrvKZAvLteOV4dfm3Wn29SEatSdWas83ClwmCAROp/ID1pZColdzxZlJDA
4k2h0X2HCWC/MLswOIxEd9Zv8DdlbmnJxCji+e6j/mnztbC9ukIpTAtCD8JVnCKc
mfcSrRpZtfK/zsFLosqI1HNgLy5cP0lheu2lFafwwyu3jSQTf9fI4OBk0X44Ck4F
jbY/GQRnqg2azaeshyrfbVlKra26bSFq6Ria2UQBlNzaKDJqFFX0FiV5IR6GrU/B
raxHtpxfODZwH9ZMuo5WhQCFuAhRWTYkfmD0oSxxV8RmaX3//cXAakkqDan/o6ca
DgPfe7OtqB2wO/0/RzChLkwvFp9hCbeyp/MJWQFNyEONjj+oCzI1rzEJJG2O/lEc
UlLac0o65bdVM6df0kc5be5+NbL8O6030WClefyVl78GkQXdnsMOnCpfBfLJH2wX
g2h7kShMBwf50h7195c7nCLSfntwTVBBRlRznz+IfhH6tzbjSgstSdo1rllIRGlS
cy+V2JebU+ym1dU2NZ6sc00+/SBQEsuLFmY5mDvw9eSpoccoU2ZvwYsp5rvlO03t
vlRd3J1eB/EoR7mDjWQAtIj8Wv80xLzoJD3UwbIew2KYQwQY5hTh7M8cq2J6P+U9
VSM5Y7o+ODZ8553XG3l/ToxqK4DvQLiWXLdP31nlzO0aPHteKbBAwCs3kWNhtUKB
NS5+tTV9IfD4uy4pXHXBmf//B3/22pvwJuSjpFV5shumM+Lu9YLIdla0H7+lQUPe
Nos/ZeznkiNWef4UXViNcCkkvxhyA3yz6hFAbpfMBqHg9EMMgeIMczl9O7bBrtje
nlBWvrtbDIMMvdnFTQpezUKuO3r8puOopZwHyPSzq3PNnumaXtZlmZQ+8y29bFb/
uRTp16d9J1lzC22nDWdxFhC5eN6cW3HFUAqZBNHD69n8xbGRBoisTvgY5j0kQf2N
FIvoE9vByjrYqvfaEgWxPk6BV6G8Ewjqy26JmGGdjJ0mNlcITFzHluJtJDkGHdO4
m4nbSiTwBCJI/KnuRZBP2Bl6I2AXqjt0LyDFlkOnHL0+JvmqVzTq/LYbKYT0oiH1
5aw+aUzFjG7r/vn2Qwf6TQczFP2aH/ujvCtZYnncZQFfgavNW00EengXm8MGf3Cl
Q3jE/fEyvTBgjA/ZlrCmj0yi0/1R+6qCMro8g3IrSaLKDmCUBouDuJsAaYnq4eG0
tXi9mqZ2WL402Xe4KYzmln+vqXzTDsxifZAxk4isdZWES6WgGXIEIqh7j/bUpmWL
4nnbxCHL7LSgyfkPVbttxYKbQa8e4azsfRa+fHsMrErEPkPd5V0yYHWmxCrSenot
y4sDXQaLRe8MuduO0uCopqwFpFBq+JB262KsqajnWS7LF5iyWQQqnVBJ3rutd6+q
HiZZaLVAHJzMm7rOkI/pME7wwuOhOcN8WxeVykLp59odNjMKMF5fmKo8FbU9//45
9sG+A/bKR0OwrlvFAi5hdWg09lwlmkSHnnazXifQY1dtNOWwD+r819JwxkRi+ANc
1t9NmITS7AaSZEwkSj8NltE7QYZUw2XPzZNox+T213HpzaYapSFY5fbveMHx7npK
JLTZX9i1If7II5VRTKzGkWoGznpf2UN8PkK/aoyJAgTJiNbiiOF+Iv+syivc718M
X6aC6NFk/cL/vswk0gWn+fd9eBRosge0RmvOCnWfCbt7aa91kDC7gY4Mv2m2waGH
X/Zn0oU8zQdSNu0QrAcBx97qo9XJBw09SDAFG4tTjCORcRwf7l4I8fRPjSRbFFXq
31BquAvYVDK3wW+u+Y0U6j92bErH3L8m5adxB2iEe6tdvx5f33o9gyTSzhKkMaGU
8iO/xdtVTV/jfuQULHUvZavUCOnSkG+R6KLHyt+ynks+wsk2BN8EQmRD8xNBB4Cb
eN4nU2UEyrDwx8WahvGjUQqJb/V535bjFG5N4l9CMDjzB7ggRxly9QyI4aC2Ezqu
7VL5B9SLQtVzrYJc+6sAjEprpT650z0zYQpojCFZu7MbY9g0+Nr6bC94IaNstQkl
vCLZBXy24N1wB06M77jN0mTHKG18F65ZXj0kuJdfbInbw5IW3YXeZg3XgoVDg1fr
QJlVZkZHpggsCKR727fx8pgRHgxfoHbtJ3HzTpoodSoB80PlByWWLpc7O8lmkCgS
cIxJQorRp8cSJYP8Vp4tkchUepFI+jwlgs5G2RpEG24uM/IttP6SVYga31VLUmdm
1jvZP20jrHeLMaunDELSVzE2zBj0Z6fUtGJoy/luJcQ/F4evxU22kHUy4XCol9QH
yqlJ1rLO+uRvQlc6OyFgF+hi0raM3Coo+fQmRkF22Fd/YPNanmF6zYu2Ep2IFPCG
iQAohqaZOROLUrbgg7RBDjKzQ2nR6SRjUPxDUuW1r/TEOFKjmRTiQy8GnqckoiKj
aCn5vF2dxR0Qi645Nfv2Cv6lmE2b2PSfqKZE/G/hMRYXltBk7oi+k1FbeGDZRwpk
r2PLITkOosfsrsTm66NEdaqReBK50Ma9g++Tek++6RwdTRPBqzPMI758zQ+iMjGJ
+M8nRQJhYMEUN4DYG96CWyyscYpfEc/q2BGtuIY47JjvKZetlbOtb3gI6/qQ3CYC
40BJLo3VO43uo7o+Aa1rMfXL09zSRozYvdZ46EnVocaSGwF1j6e4hpMTLOoYPu/S
UgD/4ZD6fAxon9jh+qSidXnmZZvppcdWpzrukqNHPisYGJzVYheygr0Dk4mWMw9G
oTs8PjgI34DLT0dM510VZavfPd1D83iYu4rJfdiqerWstuPfk0QtQ8eWMOKRlFyb
PNwoVcz60RE/1ejAbZ7H/wtSAVXxA7z605ag+0lpMDVNFJqeIMfxDzWT38hjODJr
eY6vb19kBWzO0Z6Cnpn2JLXvgiWa1EsQfkzT2ceb1QHcotYgwwLaljkeVgt3YkbQ
1m7GKScKY6h7y0A1jGGA7oJJS9dJlLqpCeO/9Ci1QAOVdqSw/iFoT6UqbY0qb6R6
pi6sdqEjlVcJSCHtQRKu8BOqUolPVGBfseV5qlD/ve1X2BcF80Uv/I8KmBrN3NBG
EY/wRJH3XsHkz7GOd4ealj0tIOVFIJK0sJG5SteKVSN3J1mIN1DqbCDTcFLCXMNx
24YjVFlt12Ne26A2Bn36H0TVJhhUb3aDoO4P3gJRr+LiIixI+CElS4QGUuazVdZ6
KTDboO4yP6343SIuSnvbO5RQns0LHWdRyIZwETakXjccqTDWiZGkndBqtFX7qQ5l
BdyemCBBhy3uvfG4dzlMXy34VgGdQY5t04tiLCbXEQrNHIaigxPQHKXrl0qysHJH
FvrRjtlJNuWjjmgCzdL5W5xDefh0Qtquu1Lc/FM1Ml65y8aumpIEPMzpmZv8GjN9
Y5/pbZi01rA2O+2Ijp5F1lP++1SmFTKBxjB8xzPtDKUEpFWMAHs+AH1C9HcS7qxx
6FY/x7lYRRQKdoMlQdygEhvM1g0ZG/GIcPBbdQNA3cYoVq9R48aImUzflbbwrXSy
Kijeqsga9vioZDMUfIWdCEI8z0Ze/KmMqV2L9N50c3DHzZehlNWX4fnNibHXTsuF
yxN6c0bncaOp7Q3niAe/+fR1QhVg6MyCQ2kTgU7jpzrngrAL+6kxDXHjMHDOk7El
KsSaG6B5udb+K+8HvYEqwR1akPOzBSpIZ4jHYq7I7v2rEOUVgDKUevmxMZCYR5zy
uny7jX6e9RGjTVQiscUQ/zvIB0RkBRLdFs/d9Bk/ISMM8w/HUkLwVe3OCnYfds48
jt6aV9qO/+eQeB4dh+yId1SEp2ny8ROZLpvgRdUtya1csVub05zqI3qcDWY3UzCA
GHVNwysn901timNb1PW/QzggmeJGJvayZuL2E+tvJgDxwh/fcKUKx4Ei9jkppU6z
c59vJxLfm66ZTaL2Y4Sb+OoImClq2HTF6Xl3cyqf0h8zaDc0HKadxlqo0L281lY7
/5fMvVdhUnaltb//pYD4jykm9jc48ASZ4xd8+HId1DnIcQm54VXHjelJ8doHRKS9
4yCNhILSyjCvgSuonfYbk5mUvSejwJRtGZq4YdP+HWRt4hQ1zgHVMvsBpwTrliza
lzVFBuVqod08Gjjp+o89a4WMxnHer6P9scFplShRbFXPvS+NhOd2BELx5DQ6hBsl
DeJQvkl5uESdlv5wnUiWUs3TwaUe2BksouUzmlAWKsTYnb7pCYpu4GHciaWSRBYw
RdVVHA6FxU3GuIQJmReAQ2Nn/tyAvSxHrlNmLtX4NTSCXXUAFsgh5oN7Hr27rcMW
aGdwM4epBZmFhbpqIqjuxQGuRyXpret3NGXD3QNj6mSZFoEY9zs3bL8kpN34EihP
TLiwuuZpQXSMsrmVYgcsFT/Ho4YCtg60DjSZM+67PdfWxxlsz6BOHqhZWu3l3B+q
EiXVYY5dPUJlzK6eeKEZI9N/UNVLT56PQxAmiFxyxKacpf6Dcr4RWNSJMuuvUwU0
gLz+BY/zifd63NoTaP9FVntPC11c3V0q7hM4xWKMYsz95SxA2RUjzvsiUUzk+M3M
yN52i929tgJKN1M9ujBfpBiDboy/pJdQNgjUyFzfroS39fK4mpXdrEOjob9g+8jM
W4WW49X476RVAuajuwhTMOF1frlDYIp4zrDexsj++hFd+aBar23YHxaHga9Tg3eF
92BPBmegadMJs3bbA44eMPjxmvZbZku/hMvRgUJ4rRHRiKXX7dtseg5DiWw3IGmO
7BwRwajUroy5WQXSC1oYnw1xCUVfHPTrOCQvjgUBybg2KoeZrT033QNONWyS2bYV
8kNWGqoa7KIAkvZBg2BMhJ1USLm9X9u8UgZUvez3/5V/pww+6SWWAySPK/FmJbOV
bpLARfQAQPzyMwQ/nxxAtkVRcG2qIDFUJ4GoUuVQezog5vJYWtjD5bITjpN9kU26
zLP56ESF3P2gYFpudVY9EPjNr9H4ebXOmmUCmcF7tSP/w7IU99mgLVEJAFwoYgxb
wUa9gf2UlPZDTMR8Fc43WsL1u5SYRbjI7e+oSQ+pYHh+JZWdCyZbwL+kCTUPcHH/
mOq0pAo8HTsuZvPxcorbaVBRqLiFrCvSf+sH6qLtjZEIDukE4y8XHZC7m2B3dPML
EW3S00M6P4e7XsiNnNMVuz+5z2CUSbtYSNjp4bX9pFWlkuAhrEcYDU1m0fwrJm09
zJQceF3gHrSQQJYWgWVgkbldyX8w4txcyCPfc3OtujRj+HBnSSgUTdhc3QmNxrQx
Qp2P4Td0ZeaTue84P5ovu4ek0lcGAkBfxUjxe8LXY1bzFfhkAaL/1JPlYpyyPQfT
yqeau/WvVtire3Mz8YmZW3ZA6/CczePIQoXlQpQ7d3nb3kniPCyEL2BAfLNGgY5M
U2ELUt/lmX5ThLod+ypwJhF58ZgSMjomYp56OFw8bqiAK0w8BzOOBAFOfuzxycpR
hUJSCjUVDz0CGzGpOwFY5UGfZNAWvfYBE8elid/YNcdtEgp3QyasFrc+ZbNLu8fd
fqiSvve8j0GC46Nbi4SGbzKh7Xm2g61FnZTRVo313IL0DJI+o4+y0YfTU1WC99B6
sdJPOUG9/KxN/uYNtsNYj5Pfz+iBM4ar/oZVpJqRTCzdFyNLojL9p7DsJUlmglto
piftToPEym4GN14ldysKXf3mRKLTWQLSRZ67Rc8yuafbzhw03AkZ/F9d/1cyKRZ8
ZvLOqDBnZKExvrLkLc9kAc4fbgovTYDhJZ7lbxg5rfKU+k7c5CgibQ2wDcZo0teV
HNB8znNoUzPTtap/Mo9U8O3pQWyGZjYen9pXf8lnBi1nkay7lv68QVjGMsnQrNu5
tQk10LjPDb7On4hGzS4kV+t5T0cxwttdmEosWEnrq6sbUXFW6NXpPz8N1LTDxjqk
VM7GEJKYDdXXwjvWUR1inwdwop10VhiyXKo/VVZ6/nJnOaMLxTsnWrE+a+B5SnzN
5naN5Z+ZbwvK6Cwp2ByMG9RnWaveqUJ9qA90IM0E2luVIO795Z63rmu/Bk6wMxGE
kNJdsiwia8JID8PraVy2gfjZrupxvxSm47XuYobecIWGSqZNV5QB8NB8s0wo0bHU
PkCeX6t7hBt7+/vRvL+ubC09IT49iUwmYIb4d4ZAgbQ8WZymuz4W+gwS/2za31e/
VEs5TIeCFkMr2lK6YBUCWdqwGa8LEln151AN05uC9xKhpIWBoh5XaM7L3+DhKfK4
MiKcL9NwP6vQzjOAbUDdd9Uj+uKDMW9vKC3IzWdmw0QD4fXJc7b3vw6zZsvxuTFp
grAOikwsdssmNjpZOCF4axyWQWa8/o8UT94l61a9nv2csC9/w7kT6ijCknYiN4Ig
mzt6w+1pLsWKVrNAY/v6uZlqyTwzQUxE2ufIOWR6JQ+5Gx4VKqHvF4YUXP2K4VFr
A/8T72YXeGCr8vkVt89s67mCPhUJ/SnOb69gtVdUk0Ic9Z6rMYyxgI9J1wdDzFYW
bT7vQ9Ja1d5OTLwGKkzjL9+4ZxvARxEpK6Rpc5QZJl9seYk6zn/DkQGQUT47LAZT
/PKQGhdjWGox/PaH+kq9JsU0WN+lNRIOwS29j50hK/7BVU6+/XpiOsUJ5LOYPguV
5Hm5MAgB40OQrDLzA6pN00isblX67YRP3He2z95cDAIDmSJ8OwIvgP6z9P6q5eZ3
4HWqWfjeanlqLJFtDsUyARCRE9zVjvk0ewV965uSbccdil4BWSvqjxPQJ6CLfPhe
poa4iOSJl+rSGjCpIRi2chFo1mAPl7x7pqV8jrpdUI+SSMqBnVRrKoAZXEJxEN5V
XWjS67pRXLv068HaOM9jRGutThnsDkse0ImZo0EgttsuM/WLegEIw2WzOuG966Jp
wAOIsZYIsF6Dm/1PHGrp/K7cIFz7Jdn/nQslGJ4si61n2x9AzbdXhruMDxVwcdtD
b3TTmm/AN8B13KDzXNawoQ/Cj4ekXKNITKDnYLJY9gSY74byEi1q27Q2V+kka5x+
Qp3nUl1vvOzMXEY/jRoM0rJNW49kSgSHtSzLVPkHbfj4hlP4WAURxg4FaUwsTOdg
LnHBOMQkztxwF2K7Ajb7FByzvhMKOELs82mf2eG+UJuXj0tVMCZzgGg+CLH9EGnl
gyIqxemZ4e/zoSy4YacjEMOaug0u9gBFmIhurpgYcMW8ws77TZu0Z2r+vlitLMvs
yrWiH01BpOoQ5ZAZh8C9gS2pF7nzb+5X7LCWcJ374XFb04AL55lqD0cMINmYomLJ
KEedJaHeo8UEtDKzXf1UdSUTVjd7KaFKMi4SQwPiyXv+JQyakFXgXltrNrJ+vHXu
M2vLc8uNZVX9uWFzgzXltMpj7ntZfxnMHrYuZK3DEnEhledkl1cTamxwt3staVG3
7fNM47r3glTcLosyiVehICHIdV1M1svFJw+SQpTLGHwndgPceFAKO6z0Xn/wbYcl
LGqnFASl8DAEj5W8nvq9ock6yglqgIeF4sEL6eAY/2pjqNGIMF/pPCdc6fvxkoRO
Yk1Y7rQ3nNBn9e0/wb3soIRffbVbuusJmnRORof0W8ZvacVzwwPfdc9+4JpC/Xn0
X8PdDYBkNs8c7HoZySDckaKtq8ShLwGvfI70wYwjaFFpNYYhEciq6H5qpFkMTAz+
wWHVhV3VV4Y6fDUcMpINwwHfz2VQ4/IqCu4gxuWY3wOp1/RR3qHD+e0bXaZ/QbcP
w+6d+cLkNajBalvGNnZoONmht63L+pc9lqnY2a4w7tE1epzTtQ2ftP7ElsmwIPwJ
Uj3tO7PpFl3FJpEDd6R698VCPY8AW8qdbDQVmIq0zKQgp8dus32c5Vta9RWF2FXS
uMu0VIf/QiuOFMhIG8emMsL35G1C6wlx+9SnzypfDAAWePDyXnlYfknv1zSaEmwa
OZOgw1bBER+/3U6VgcjMb5ewfr3vVKR91YdqQ50F6vIbXYMYi1O3zoE1XtAfF83g
x7MVVwgPlOWWtiAwdD0pAAqoo6DFb1k8CgGD+XPWqoefltn0+twR2ze9naDvqNCp
ANJy5eie+Gefic9ev9saJieHsYWaGJBM04vJ8o0CNuC6l9dEozJgHy1BMYzc4L5K
ztN2j/+fwRVgiCd2DmprI87l7yha3bIWYaOPCLBpP86n5ttH/NwPT934exQA3vLR
9fGl2xhphdMCJs1xOoJ7riBa3OwsLYYfUS4X8Zo+Fm7IE/020iUavMiGC1Upxe0K
K9r6bK2v/Xh7PiWaRVuenPeeKnBmAeMk6tnpaGY/RmpSMES/OWr5CaE4s5R50Jry
BvdpkHhl+7CF7FzPxw3NaJb6x34TZAkzOJXeqfat7hcBKrJLbH7SKYZd23O2Xm3W
JG3XlWc4sxZsBwi69OUTkhkpM21C7VRKmQS81darrI7zh/6hhqa6Yu0HtnE0av7n
HKGarOgn8ELnY8KnSPoL5OSsTv1U8OLol21JoAFEd7Btt3sbE4MLAed824FBOdvy
UkwcmjndrTKrA3b359a5nWLja8EgiT4EoPm+mGPZ5PfDI4iCD/NSEO0G7IzQZEFc
Np/vKrl4DYGF0mx31RN7CdvsmHpEY7sh0dKLCoEs1aYOA4FK9vw/SpZ7+gXnEPfv
5DmNOJiVM1OuslQqMIVYzTUizbqpT2ehH7Svb96PFkwYuaPy/iZ171v43LbbJok5
iLQZhGRCCKwj6SJ/0J5mEvmxBsQurb4OuhMjl/K4aDfkutkxtBmdQYc/GE3nr0DW
K9GKoqtsyU8mX2dtqpeUr/gnR9huaBDUjwK2ITGA28bSd1BGeWawsiMC89aNJIHq
NOVmGZBbej7aqe0Pkkrujk4eRME3JcSB5EFwFKU6VqYefUAgbY1aRk6yjTGM2B4l
m2CMMSF8WuDD3wlldU3EGcoCyGAPn64QP8eDz3ObBn3qZL+oYtItsTYilX0kpPFG
G9ws243QXQ//Pvz6jwP/zifAaCnxA4sPfQS1zqtxsFyoHLzXBXc8w9XL9ybNorAs
STdeEWC561PP5ekl9kk6Q+k/5D2zt9GDMOM5pqdgs5JPUIAdnNOJBG2o4SKYT14N
muiK8kgZSBTFlZuMRhAvvYkzMb1DIRV4RV8RPBTbmI23j9RG5vl5EPNu7wG9vcy/
b2e+iTmmpMLs9wHwVfhF7vXX7fQTSLu76NzfmLxx7R7Uv+rFiRTgvcC0lueT89ns
gt6zV6lQmbUsr7kkUojZ3LrwUMAiQVqGJPVmTjRAWtUN6+jkcLEc1PKcX7j8kjVh
G5KJKI5tp+45o9f5G9f45hu7/LpqLnb8A5vWUmIOAU+CNec0h8N/ggtCytRiCeq0
L9MWl3EPJut53CN/QPav2cUOHUlfIJbTo7n8quYBwjbnH6PkxUcmdgn+b8Ixw8CY
mqZU+rZpZrZWURnS9rqS828znYo1omWkmGmp3Qsb5p3o/34RbJ/s4VzXnUBs/iz3
kPD0gx/ZhvViyKG68wsOthgaEudxgzUWqMKwbhbKXDCF5JXtO8CIuYAEn9T7GKO3
mYWPaR+K0IfPlj/EwAoypEEqD0Ga7ZmjQsR5mwtYKzVJn6frB8ctdK1uxOp9BNjc
LASa0tC/ktYXh3pklppj+vB8onVpZb4u4FY7TsaSfn0XTQLqnMTk7+OLT/LLq6Oy
sWoPsCTgwG5zvdoHorSmjSWSUY88C15XRuwfuG9xtponkTtF1V3kglxQ8u9HJI9g
//thFCKsTcmJ/j0HwyUtCflM+xOsgVv70oGFMvCH9j+U+oBZh4EEe7anEZqo7YsX
yX7RpVEKGt2Ul2xjc/+KElZZjjxRMcMFN2C+7LvPNO+dYt2zKphlomzEqZ4VnGMY
d5mQCGy/E/H52wnr+8FnUZ+Hs4X3QNXjh8MbyDlaHj9L6XavT5Pbx5fvF4EwW3o8
n3DAkgA0C25TDDWVpuRdob1IBAVP6dRTxqHovHvpGozUUW9Cdwywe8iY9+esVc+7
7PHJ3o7fjAikWUvvUx26TRrjI5pQVPO2sBLVaSUSa0Nt+HSzuMQ5VkLwUXROjrjz
QI2frzR59wRA6vUVfaxn7mzww0NjPcNhi/t9Lvqs1FWPQ8mpuZjPsPm/WeVq+S/i
O4LiqhN8Ws0tS2HdJeP9tUFqCXZCFHhfu7XNUa5C80MC8KBmZALkYDhDGD6PLlhf
WsSc3k4du/6NAxVIv70a+gV9P63bgkElWsp9GDdrc6SdF4GicyC2xR8wfHk590sS
4JkOkBt0VsfZLKs5v/ujQhl1Y60r2pm/bEPBnfP2pacbPNSuHu2yt24UT0PlnOzn
LSdWde80d4NqTZRSWuSOuMeWnD/iq/yTyRTOoLrDdHehu3iZW3em9B412Kseo5Jw
a6XSEcR+WAbW9d0SXCV6+F/+hdRNDVNLPd3ANIDLMzbk8crpKfA1SaAzCFpZzsMB
05Zv7tnYrdqzDWC3CMn49zY8fWSU/ZIVlu2qzM+fO3NMZMGulS0MIYzkJKhpGlbg
BRuAe4JR8ZycCDAH22aVCEMnTPF1hGcfexZiAGlDiaxoREVnb2Cn5Aza455+vcLf
6r4oWOQyM9YEZkDc1KiPN2+8TLhRAYsmrrmeNRa6oMRzO6ar7rQnjyDAkG1xuwBV
U/q2cU5EYjM2y+A/vOL6zWzKSeujbFFNlteiukvPYsiOZmyE7kuJSk8ilCVrrfHM
6Xf45TET2ot+2HreGu+d6DyrDZzkQOeC9NQZB/8JV9IdfiEALuF08WJdioM+DTfi
N0upI/WVrWRts+6mFJ4YyZCoZRoXPhuKi7Tiy8ERN0lr3v5FveMNGXR+x2noZ5h+
BwAExTH56FzCWOZdFXTVylh29yfRMtf5r9Jfqqed5w5xNdPHWNM7jMGH7vqtKAYa
TzjPBf7eAXwDmug6aUXbbDqBOJWUdfVw+ubU5h0Xz2vAjIVGod+zAe8mcXdbDOZ6
CoUWcMYidnZ9ue5SWX5oFJWKYGc1moF2nSxlCzyH80ia4+L/ThuIFqKpNcSx88nJ
zWbH61SParM2Oc65Nhw64Ho6Ib0t4IJe9Ye8K7+xnMNO951h9CYdJ2Lb3CxYu9UL
ZKPQCgRNLnJpjltidfe1uMJnqLFwszc5FBMs2XkfxGFw4+rlotde3QquWDhkanQ6
NmuVQwqfBj4WEB2UYcsWpOaNok7lgDgWcWJmQAOaMzTLfITMp973AZESj6lpTVlv
/aIlpgH787jE/4cUG38mDgOoiwRrx03NQhHM2IHztLQwFe3TjPkeZSIYk8CD0PUi
CxTS4knZ5ZGmOAODoGXQ32Fnw6e/iDoSdrapHk3px9D1Bn81wOSfmx+FJl3KQMMV
LQZj4JyujMYAQww5opYkDBRJM0jeRjlRsOzClJiBbUZNxMDGjKbZhY0FyLUfcd1Q
24KVL3QfUzWiJFbyGYs3JhVNeXf+4pmO0o6cSA+CXOdkabX3mcs0VW5xHZyjEMtQ
+7YyimnC3Xt3Hn7Rr6nmQQk7spRb+e8fVr/0AqCBtzamQusHjQ+1cHQ/zpQg/zCG
m7HzPHhRttYRpVbDeqATGgcRb1kWDjlYQZLg4qi3iVboKj9ctorqGQyBU32sYOYb
VTOvxKtyzxkRnOMZZOpOLl1XO2l5wzse1HawEMjjnx2poldRnTMIzlGK9ze5YV1R
o5lSXAFE4moHwItbWQ0xcklMa1Wr4ZwWvnbrBgWcblFuHl3AQE7UpGe9SMrLxFVx
bxY5pz2jZYgHr66lxYNAVW/gzRxaM3fPjvSYIVRzRitfSlR2acZMx+nXDFqp15jJ
uL8UZkP8WtNXBZLHpF+2mqEvPRPsUmeAjLsF3F7CnH9sYzbMQWrOJ6plmrO25ADO
R7tmleoPTPIHQBI5+yGxjoZYDTOV6py+Xyh+1eMq18XrMwzSZEuX3wf/9FKrvzfn
E+dP89vxhmPgFGH/eAMsxahLzl9HuGAYuiujEcBnd8Iy002yA6Mypeg+Gt0LPOsy
w0haNb4bSJjtI1fgqaQN4/tyl7r0KoTzpztCVoo5Z06zj7So5Cs03r1h+Pxu+0xt
tXtyvBHpF9W/Y/FnNZ+s2XoGA7TnyyVGtzffh/kA04MbX5f6ZmMO7qLVe3mjHRdZ
/xJoOTPrwAyQvRQqzV/aF9TGOdWU2a/xen8WUtnZodPG26C2px7i38nLvEM4Vrfq
pYflNtV7CXat3t/lbPyny6Moes/nYIYE3g8x0vYxyLR7QgwgMitHXnpUwX8RwfxQ
yesGC2rUsAOli8aGChpd1pzb5SPHorUrNRPCjs6gmPmrQOQKTe2+qHBx2UZScO3B
m/ID+P1uphE6ORMzRc4yuWd4e3IJwoyFADlHV2zIPfIeb4bArYmNIfnllu5aqRFP
JiAtgjcM5xQJeLWy2RIZlc3mXFZOaZgAYgmOufWi6bauTr69eKAtvY6mk2L47Cqh
7K+iMukXMf4fNvdxsRTFas3nIzFWMgk9hAU/FhXKa8CQsCFUBHR2mOQpSJ88WOc9
erA1b8nPLj3byOpvKLO/3JLq4pMXuqFHjvqlP+debuPzAPrGdXaWViABSggOjJcF
E//r0xhxa+PLx5kAmsJGHBAWPAsCY/LDcXVtUyhf1CxjkdNDPuWxGY3BkYr6BxUq
BrE8xSXURmNMdTMfb7If6rpNbb0lo9ChyUcIJJR2kF1NyBDb9Wc2NljrsQE6Qy9B
7xTqtZ3Tonylcc8BTTTLuW/eZj+pNS7FN6b5XuDrSRTOqzJKE3PjUvdSOAkdzTad
Pie2FpMGfGT1T4zDG4RVUhbUudpAcR5c4V2yEeel9TCFfZJI5la+UZyePiKhP5IH
BUELpYMBlwQetxzadqVCATClYg/n3vdMfr2/QegWmF5AO4re8GPaVkalR34emvOq
YIbGwvqD4aHSJtIka8RKdZnV03VNKw50Z8FCwSOoK+zXE33VMD724MjK8kWrNi2G
pWuzQO/g9wIh6fDIbb5D8y05qOGfpx1nqDAi24FZ34ClB8H7CeoWTt9Tso/DrMxE
FPpCdTP5iihVxFZLyGCLfi4VKwFTScEG9qbJ/S+LhN3HaXymuYdwF0kWx1282CHT
tcOM46afTOazDIw9nT8+G/vRRW75gAS5eRA/QNsC02Urp6KuEj5QnKMJaXTZ5vyJ
LZGAbLgWfE1Y9rL4IlY1Fo/UtjbnbnR1m0OqKkxyrV3ClTvxSLwiVunfSQ0uqUgo
k25j+FSjboALMHw30Wh3kQIiyZJYAPxcKdEsZ/b43qPJliifqP32fi8u9PGKgzhu
aVKD15srbsRSCW3Qx7Snlpg2egLMPRcPjrd+DqTotf8RVSysvXdWywswqPaMkJYd
U9IBNqn7H/pXAidkRmAo6EiXpNbGWyu+HUVWD9JVur3J6nmsH0HARISs3giczSVS
LuzjhWHHvZ4xTbif6WPv3pQrE7iWcTke6bynO6SfRfOZDiJFPwrSMU9Wr93BF5Uq
MkgAoEqUDXHR46nTOpkxCwmbJlM3E/4dQnzh2XxNcTHoDmPoTQLQtjdD10hqamwT
4YZSZIaXQoU5V//sVm0LUA4BluOfHGKgjfW+np4aqv4Bc2Pm+vyYG7enlvrGORh0
KZFcKtSVOty8NOGDgcSFSVoXRgAADBRD9f/SRRwrwm5d33Kuol0vl19xF3VpOYMa
SGW9qpBLUuzWttSNHHUotemVac3hxLIWg3t77OR5JHwrSOE9Z+6By1b6FljJEND8
kNyw6JczmwBkXofW5qC0oCV86jXcqODfOnH4gZDMv881A1x7ZtPwxr54zZ2282dQ
RlmI80LRMVnUYCLk+SCqm/rGnPix6nMcqPscdQnG0udYOJxGV3g3DeesbhHjiIBx
rGdiNqVcMqknb4WfimZjKf2NaysbuWD7NtL0cCjf2OYUYf+WxNFUgmcTMfwXz96w
v/JMJtNWhFkH2FKJaJTKtJFCo6cYk3cRmQwLs41Eil0guJhumhTHYYDnWpvgCS21
jU3B2OVGz+2PY7d0KOUj1nx5TFttvleu/+2HF5Q+pXVaMLxH+N8t8Q1GRXA9Jnrg
oqoQXSP8xjjJYxvSze9SBSEkL2hMWwDqI2BL70/gDUe/1Iq5ZcgFup+ldBWXGdJ5
9bdwkRp4xxmhudSqB1+ykDQtudjgrvyxVezh8hQk9jZfqCrP0I/bzizT7HEzP0Rf
uBZR28Rrx3VCS0ClZxCbTrsCNgG8vfmI1MmOiLMjRQreyGpD3/MSFIbV9YdSM94J
M4+KpnuvmeVT6V228VJ2v0RpbKUbfKDEpzl9F1JZPZAGnpGbEcbevE38etg2/I03
CJUp4w3rNTGHwLvyTYVB5BHviKoT9pi+L1pYC3uALXLHg9is73tFeR7Ct52wnHjr
QyxqgOI9EeaQ9GWiKjESkc966GwMKJO6em2zSlUsElIOOb9H9/OXqq5iUX4MjZPy
O2HBTUIlvHfj7LVRDy2mtPIJfKiJxfL5/wGcyPeuo0E4trXrqapGumQDYLOQHlUM
yYgbput1m+1wbcpEzGikvJMGwia0t4gJ4oPOcOiPjcQJm2oQ5zhG43jD7dLz7F/S
AMuBCBn4CNOlOv1fSDg/UlVZKh5/fcvcDtgfs32g/GIq6hOFfQ5irH15hYIA9ZRv
d+/bCnyT28dGjuG3enyHmZEAIo2h1huT/PPpQ4giOSpWgy564K5rYZ50NOCizTdR
9WKlMnHl5lq1OZ9fRin0CpMtDnTUOK5uc8sb44CauRxENTSd9u0/jIYSqyI3d6/L
EYU+3ikQuaFZHTQptxskGLIZythrSJARcZcvmgMPRS+Cc/3D8vv/jUJ1/dq6lFG4
X4ii1LSQ/ZT9VCH3JreGLX/aUx9HiKw8+UzdADrGd2zAen5Pfc1f33dfuTcGJO8w
qegrJ3lhF2foSwMQOmYlN1zF70OVOXdf8yZF3A9dttpxyw9E7NkdAM3UzBJ2t5kB
GDidUM2DIYThA0zE7GTUE5Rvc5WK1+pBelWVMsCtXHdaJDy/Ds06y/Z/QWms/bsN
5ExMtoj+b+k2oSNGd/XqZ7tvisjrKoL2Ul5XklBvdIUBP9iVchbQL0eCvWYTG+fH
6+NaTrND6qO6Uaoq6taCl/5QsNtnDbwz/vMJ8bMKaYUukQSt7MlzXC5PM1ugaN+X
XvWJV1DNDWFU4GCubJGyK0ZtoUx7FlhYJBEnxB40VIAvMK5YdOgigbGrrUMfB0Q8
CcoJXhf4DkcpYyvrqPDJAtknNmFrFPpyeEwYbhntGWXdoDs1fkiDkQg1F6U9kMlT
EsNwo2FuxdNpyQUmZ4Swvep++ufkJoWyK2/HQT8fCHoZVXiQ8+WKNRFCtG1xiNfJ
5Ag70VYVVQdWXMYL+1pHvocybrpWF9Sa9du2132keyLKqAuwMzlK9Mo1pEgVVeEj
VDsYwA+E0fPri1X8MMLu+eoOVjSBjq6Gr9QtV6YyfYxwRiZ9TbWSS+BvHiyxdTfo
MBflsipAzRzBTXE3ahOKKTHNOk3Lx51zirnXZSHnWMPaN7VZEOVrQENDvydx6rLH
pat9tW9mCfuUKHqOWPLboNsQneL6ABdMvi3EQrklYiMrTFyCjWbwxh7WaY/bsz7d
Bu0UwfAOAYjK9Lj7c+bsSgv6tSU/M7mFZElYiY1LnHd7I6N6pgw39Woq+18Z397m
FPp6Vs9JClFpk65mGrnh9LNF5HnZw3uVxRel1RZejlkhj+ezYOChUpA6x6ndBhTH
qD89et87jehNF6TsMsfLLsAEQ1ASAXB8B1sXbL6qzQqEH7koa2tNg1ApHhjQI5hg
Xw4m9Zat1bwdAKUSkhgRNf7ckuAmRBcVRCJxxXyNmaM1vv5v3+vxBe2bvsGT4SYN
vyeaUpDqJk0yqAMQ4qKSjq7LPdfRWUuHW0GtzGiq9CxEQt4rmPplUCcZW8AyUffR
6xRM4hz8tSaTUSGeEvr6gNokig4ZFjjehpoya3tVzXiPj6omvJ7Q/BpRDL0sRGSJ
YA+xj8jj5C/hur+Qk3zzT8ZgEJCfsoaVwRv98BGxgFEhnE5VChh1hsGtTUlQHLjm
3ttTInsRGijvISLbvvLOCkDvDXt4ziMcSUq1koTdaKxwK8SMaXtLlhkU9vpRzniF
LM8z0Nqc8SOXbtRiVH3GRzCRBEQNHfu3gfUtg6kBpS/WB4/4X6e771FK2wMiaBXH
kzoxNnn2PqlznPtMjSfTkWSfEczCweRJY2z3yJV1oaOoh0MVbMsn9euJ2qYBlp5x
4HLVkbflAh69zkK5NlDe6W+3BpOodW4dIU9sMMNDKFJM27MLxGdVNr9cZDw39wNK
XYYkfuCGQuEJMPWiygkmY9su2UlON2nbzuRWFa1AEhXfRtVCvGAVdGmF1P7MlEg1
hPQAE0Gewef6k5+xci/z3sScrLtTmPPdGc0tf5sF5XKSFsBrNCSEqzz1CVGN1gpx
T3lrc0phkoxQSbWkVJBAtUTtO7SBFXZGgnUJn0yqA7KCagWVlsqiAMqFFLxrf5KE
6DU/ScLC1nhxSg9Bo3Pzl+naJzPJD9E1zY97PpAhh3bPnjUzZEklromjN1Gv667R
pEYiW1N+xv4MpNGoNHRsE6ONhF7xPSqVuNPrBZqY625MGRQc0nfkRP54YcY/w1oB
uZ8Ol8WIc72BWhFjHYRuTsjHeWb/gck7/Vbogk/cx5FWrSl3WsXsUigVW2bfAKF2
5iisyJOtarHdDB4Mh/zlC7HLLBKwszwEU8MnQfjzsfgmR8gBL9U+51IrPZDH5v0S
xufPFcIlsK95GZJRxy+ukPXWx2AyHi89eFcZE+F9s9zD077y2Ze8or4t26FH9nUs
hcxTdfPqUAvlNoMwWkD2UIooMiJxJ/j/07v2NgnjQaa0QUiG2OYFlwjIpcMGJqRe
HTJ7xPULo++8IsSjQq2ipWXBJMTv3nzRrVAkTSu39aFVC2eGDh1ajjW/aOlH5ewS
FQQtSvGoh9naXe/DLofS7L/fgyrXnOyhCbmDJF4U5MEHrBsPxpdX3dPa+H1oIZAn
TpFlklQ5/skfpquAtoqrW/F1Ixg4PZFm9h/CkQS9wXdluL/s4diXud4lVPBr7xTL
c0wM31TRiigMbPkchFUV9ZY1uELwo+uTD7wpFIff77+beIFDkydN7xQMTvGFEh5v
CzE0rNUiEBGTJ8BknHI+k7KHk9RvxxDHrJ64tpQ9MKZcfKIkOz8tJyw4y7BhjwpB
abJEinLb55Qn5XMu7AqwHM5h/GIfZWrycRpM7byBc6/2N0hw+Igq/KZiY3kmDE+r
YM8s70yKVvqwLmRVQAAR4L+IgG3w+iX6AztoXKIiVMn7CbzCgUZjiB7VRMoyVIsd
vIbEdJY4UJtTZm8O/V5oKBvde42HvL7KLph82aa7lPnD4lNmPg3gj5HS2tTRTVOK
yWdFKtv7N5hyEgf69W56uwUin13/DxO48h/AeeVmmMJjORmXUJdl3eIMEdEUbrnl
HTwcJOYd45pzpn34uNbIgaN03uQS3z+8hkqC8vP5kVw0T7CQxV49xBk13Zm/ERNY
TkqS/1eebuM5ngT2nX2QRW6JyLQTiAFOEpw6hycNH2lyhJlaDAhMhMZ0S+9HBbCf
jgOBKM/LBz3+kP+sPYrC72WVNqVyDl/lxkaZFMohWPNMInj1uOxLvDsNAOPEJEGJ
EjzauNh7DVY5h22zx6MyWzXuxQbxzXihBBRFQ8krkouy2zJErRFxQUqCesD5mEGz
+P+15k0oRGUZco6wL1ih6u/stfRO5kwPEcDZ6DG4v6J7338cXNoBCoN4fGhBVoUg
EcTJD3IT9PtemEDDgpORwbJn2TJTowFVUPoWBa5AOBXsAM8cHFRABfCjxQ8awnpe
ZmSYY58BLjskZH7SBdHQ091LyNyP4hy/BUmWeMD4L1fMV0uEzySYVBqOw17lPgS0
ygv6tRj77Li8X/oIO4DR8InfyfDl71K6HqFZckNfVID6ox4v0/kNKq1yLKZnZtjB
/m9Kp0/t1tNAONdczF+n+0+EZawOA7hw8lD4fU0vwwY5PgLL3oMBkYuLwYyWjehZ
89Ogg4P3/LiWceV5ifK5PTqn5L/3jvLnL99Yo+byG5RivYQ5H0ORj27+OkT8AGQW
vcO6Vs/1go3pUAv8J58gA/QTu7+HeSZCvmV+pHVv3D9oeCJCw9L0q3YIUWvWJqJW
yYvG8imG+Hv4cLIUB37vxWFxnp/TbCbWa6U35QqwcdBvBUHyBewUtGtvQVu7R4Qa
wSAzoSNT3HsmXsq0ns9P86yY92iN6TqGSSIxVQchydoyTZOmgSpxsT8W8lIRhIOJ
mOHBDCYKwdDEMBxh3SoBzWM31o0uYdiSO2te/NG9ESsuwZcsXNUFcUhpMcmYXE6q
QyFN3plObvT+3EKGlT056bGUyMcdbbts+m4WDNi+uz2xASHFdqsL3NE6Av78IV76
INLkK+JLc1l1p6+vBv5oYEXkSJioUh+B1D1zyyV/JLYJelnFMSbacOqXWvaSOYjd
1FvnHpIf44+9t6YbjM5jwB+MdrR1brFaiWgKwX4d6uBrxS4ihxzp4vTiLz1ppcwf
vNagNOsrVa9wTLGtXWUfA1HsGkZ0pdawPrmgAvRTnh8lV3zSawoe8jSbkE6QqSzu
J7SN2bZX0Ngus2BJi6O9qYWFar2PKs33wtjc8LvmA3kwW4GMbPBPiHVq4tgZ6Rie
twOXQy/m141vSix1KApv7lG6Wm5K0sO0Simce2srQB0GLVbVXzob7gwYn0YnsVzv
jUmvreTTma6QR28Ab7hjGt/tbR/8EVc44vsJABaz4IUPxjqB/ah6+a3Qm0TnHjeZ
BJ3FaZD9OrBhcWI1qvuM2qqxgqC3svaxTBJbMrB2/mRT4CauCtLtpXtVBlXoxnxz
9rtDNwbIYQM+n0ddk3ahI8Sc+UZ4DCUQHdwTo4Xr0k8EaTASislVGZIg/cqFeqc9
yF6GYRTQRqs0bP4GrTcPXfCxQEfyz6q5F9PUdDBjYSThJRjc4Ifbs1/KUfdcrcqt
p8fRnJkKcOhXLdgQEIx8IkK0FTfzlz1aJoUSuEDJOPFJ8EzXSdd89mahLHWajdNG
x6GxB4/jSZO2Kb4KCkmzquvspGOVxbIC08Qn7uiYRfkXLb80sNFzMs+lE97p7JHl
naEWekUtYB4GkwUzqmjcSqFvEZZjb/QTyDlRfq3h89O4zdSiRhc20U+Z1jZUS0VB
tdBqikIEjyXFgKhEQNKIgBRXa3o7zdyMD4dnVeqQZ6+4EFapBuoVWzYEEG6ZJNA7
FtnEGuac2q+LMGiYr2/IRqrOl3gczB7TQzvji1MiNQUwaDZmT0SSNuXBSswodZyI
067bzv8eok+XCiE4A8XKjWmXPsX/IIXnbN/lf4oIFP3fgIo6gEvsoMd62oe4r5VN
FiBRwf/egLxNyojPlfxv3HWwPDdqjObYukh80Z9140ODPrDBancWQkSlCEPm1Cjc
y12F2YURYEyQ4emC4VC9ywsrSCS4Y7lemBvtcXq/xvPvEJIIoQ4hOZtdTDeWa4yK
lIDTbKFLMs6jBSatC8nb3B7+A/BsiKtQCRA04Reukrr3RJuhpUyc5NYx9zSxkI3Y
MdpplNeDg4GoexklGICwJ7NRApTdSZdDeMmI13QOJO/NvjeueMb7nvr51CAkW5sZ
aGLOAIq8rZt2nGEfKpDB6OcCcxIf4nCfZbI4fa89mcXh9aLyMoq5Kv+bgasIZ/cN
FDSGT1EdTMzxwmvErwX0YJnNmsjbV8I42d903ZtLTjiIFAqz8GrDwmUUtRRIfPcQ
nWXeCW1G26LfGzJWBqdlvDP5jsijS8ndQQRUFwXKYp5CM4OWJMC0FlN03xI4eQfg
xhfunncxu7stnyYJbZ6husOzT6ZzXyJQ0BIgs07b6phi2TBy3Pij95tE/341aNuJ
9/HxbdGt0IT3KaEu1nzyKt9FQPfB9TOq2f40EQF98x+0roSDCNuAWgq1FuRsH7pg
fIYMlwzQpAhAy7z7DaiolYFDr3lN0cZKr3+Mtaun4ePEDcLHKU7a0hwFBX0xj72Y
yVgOGRjLzsBFt9qJzuq4IGu+uiY5kvqNreCMq/Kgj0I+wbkQpKbKuyHxo2mNkVij
evEGRJmJSuLx1akiw+X/PPwyNkxYMupeVbk6UTd89IokHEAF0jkYY9Jjk+6dXyKa
QH/Vof4PxRI43oYab7XxyX9tehItGGQFBFsAmTVKkWImv9njS8ByofE8sNUvJY0C
cmwuAAbRTAhVc1FRHiGXRkVzRFc6ZA8Tg1lMzT1JKCwaVk9nPWQ3iS2ak4HUqgaB
bCea/9ytNGrlAJeJnWKsVSnQ5O8Ncl1Zkr8CqM07U9NofclqxPzAS20R1Wk9dVrz
nkU6Jzy8T1IoRVx/pG5YStz8qhO0Bp9oHZGSAwx0yWqc5FUBfcdGsQoBNgHkzNDS
lkYiVyBDkCvKWhyBXsqfsTntl9dZfDiZouvX2O9f+ilgwpg9/lqeLj/qm9YWMbB5
E/AvtlXF2EIOEI9aUs5dzHW72p0S3DT35O88ga2hqVFzxDA3lBkMT7ux3Uix4TDu
jmooCyAsLl2rHsvvfMtBF75ktS6hWV6OoX516bt5zhNibpF4KWY1b9MywsoC3W0O
j51XNd3ou1wGk+zMtJMpDSO5SizA1QBxoTBZD/2rZ7ZpB9zL8wsXb7tyf6QeBHyV
NDQ4HB/Z9i6BGSp0v83ITWjsiSGUNx1oaPL7VVz4Y6e46AGrMSkOptAEA8B8Dd+i
6g5ZBcxVmvt2GlfShn1gAyrdC8Md9/9qWQnRMmrh24hvhUNFLTMg4c4hgDZs3aUq
cyhP2gEcSnKMUqPzevol4eH7UKyU9L9RwHnXqImJjTCsdHKWQqiUYhSNnRykJ986
r6LSKqZgB6nJAyWg7oYgNKL/848/eNYkY/0BqhLQqQVZubtS+xVzmWParxsKu+Zq
LqJU6tAUOZs6qfLPZIuJ/nFM6QYEWt/CC8T7fhM0obiDNcD6bDlHkudEMYl6akGZ
d3rXwX4KDlJRMZ5kShCqfjZEwPOT0tErv7qEUsEelEGZzWmE2tLtM1/q1dMpTLRi
xLuQhq37JDhbzu9fMiY9vfkDna93iL03B77PIiVkufVybG2JWNz4iK3eZimY4kN3
MZNN9E0oKzZZ11nd9D2/W1TA+wlpV7wDiqyeoXCn1KJAn0kTcmPH1LnEUu83B7H2
QWwHp6h1v+oLt7bIACeUFR+dzpmb/93yn0hnVpjHNsbveW4fDHqTKiPDaZNVP2mU
VQFwSe6q/MfYtDOkBibHSS+CuNBT+sUrcVzTU6QwhRTSxHXqBlGsqYgIo2FSEWLP
lz5PKIWu6Z0von9xmv7KfY/vSxHbwYzBiiFPPw9eM9DOI3jRu0PhUGo4hjxHNO6i
MxhqgDN27gkY7hshi9fxDFQRwGG0+Q0Z5DHST10A+0CYIhGyLr+HZHSiijeqeTgh
/ih+XsX4zj55aIICPQ3J+DdybHRuNdUWwUOLKmNVpOTZZ+XgJ6qwu5EnQGSH0xyr
5ZAlz9YaixrmlyYc381d5Y1u/Bxdu9CtDysVCDzHpyOm/jfPl9rZNsmZ80C+xJDS
/lW742sKSNr3b92wQYAlPzkKkaNQIk5FfBb7i0gn2Ebcj0FhT7TwExMd5N0PUtWq
G3kmDVLv5sBz5mjUKicTd4P8a1A8XOWkyPV/PdeLBA0IyF4++N8CnrmESWBeM+NV
NRVIBBL+PqY6SLx4s6lCIe6tAIB4V5M3dFiG+yiLXHdLfic82LIUb4+efcXmmGo2
2Y0u6kwYQJ0n3MGRjS7flLY1ltBPGg7XUXcnCEvAqfL1UL1NW4Kc4qZPGUy8+7s6
83+PqJvR85pwi6PCr16o4pTUmwIAQl/nwQCCQU93GHnXKxAmeVdeqRxAlMc903cr
ehWJOGJcrHeggAPIVVtQ3tOesN6RPniv077koSzJma/3qNPTcOQM1uQHoX59bwZ/
LfDc15rbskirByGRjATeEic+Ww9P52PceeGJpqVk8WAPVSPnUh4XivTwmQpXQZce
2Y0D2mfmHYAtcS9Mxasl2EI7gddPZIWBeiq5GEb9oTOK724SGYtge6bBHCXiFGBw
jfB2pMsuqoAqT6hkaxRAro0hf5kc/LhEnaB+j1p712oY/80/KeIaRVEcTQDZTHe0
Sr8tY7bSAWZiti/QVloTOC0j4kSUSWBR+9UOxWyWqnlZPBQuB8tqDKVeBPGWWTep
E+IdLpCV/+ICHerewh9fc4hG9Y6Tr7WPVFZt+ZPmFheR44G0cRSuvAHHJpshicWo
GmHujYlex2RLVTANI1lvQ707vmxizJh7ZKEAkYez5bIwLUm0YEkwkQs9+djUwIjC
vs06M/mslhFqvjerD0EwYYBEszUMFCPDXOLwMe8GzKuWKQoqHBzriKtGZkOFgJYm
xAXcfJauFJAf8eBpkJCnCU5c/dHNXsrc+2K7mxoNMvq2dU1/JIhT9yLnTf2S1TC1
ZPL/MAM7c7yILmalIbPHwtzI7HoJxEDu6cbWvhjDikWFxIhZdUDT7lFmw+8I6wTR
xn3MoQCzE+l9CHJHFfppKRdLRfDWPodcz5uZ7qCrTDYTJp3qX9EaQHbnhT1zD/jm
1pP9KEy3ckuj7jZsuvysY+JkqSy9pNBjkg9xfeSsoRyZKIQMxOk4ZaI7LPz2P/yJ
3p36tY9VwBj2h5D0OssiGY1hxeLeXhh5MfVLtHdXu6JICigSETCKfY2MtCryn0Dg
09v/5FwDN7u4s0UsP3viBbdYxzTZvBtLGH1H+tFV3b8CSA5SYGZiTxH7C7VEme6r
SSu/NE5qny1WfF5ZAP9i59GKOcIKJd++9NrwfiXVzDf3WFBLaPJMfDKJCiTvrKxH
mwt4uJSaxxI3FaOSXFwz5T4lg7fcAYeuFAe3GxV2lwvkv+VrTucR4S5IaQFpDbsX
1JanT9mLIKRYinFTGxhTBBtwlLcMDTVhBe7/ShXZN3CvrwonZbncFtQ/t+UUjFK5
QW8lqIDbhZG613b6uaOzRaQIelTkBKYuvFjSdFU618d1JNyRyAeIg/GUe1f7XP78
2Wo7Lv3kd3gymA72ZbBknI3xQMYdfc4VYERTxVgANYktNoRaCV/+y4yLbUrdD4VC
BqScjt9esjjF5MBey76JGvgnsHIpJjMZGiVev4I321r+6Pr1QHkyHXdQlJl9Tosl
ubxqeQk9IxUUrIb15leXkZibnTN0X6IubkN1/QR+0mmZdWo94SwRVriM9A/VTz9O
Dy4Vgvmncwi6xh+l/Sk5KKnu8xj6XjwOXPt4Ic750zyWxT3LOFyDo39jjZ8MW3mv
gNNvGpk+gA9LKP3JVW41zRsPlWRsSTAEaCnxg6ro5eS989cLI0dPTYac3Gm2QB+B
4chW7+5btSW5arimWyJ7rpqOHx7KnSye7LotLZIRY0x32nmOsvpAFNoXtEH2I8s0
4C9B0N2tR85ZhUReq24WQI1D1H1+/0GXF7mqLKXJCs2T6ZR1d3Zuq1eEsQJu5BAF
gXJhhoMY9vhBNMGwWj0ydQUjzluS5XNfIohnVqr8QzSCvCImWvMXwwEL/AAUg4+z
8RzuAoXmGq0GN9nPxqYdtrwEt49UbvLSgy3yUwXBsk8/cc2FXc5HzH77ZRtt3z2n
uml82rLrwiB2ItRvM5+sh6d04UoDr80H0j3446obwArJ4GdrstoOutDqkHojZP8a
rROGawCfYxavnoAMNsETQbMgRxGJeBDe6tJltzVsjTFvu+JwXBI5uaHfgK1gIfFQ
bKnqDxrZUNLppKdFAaEtFrg0KH2Zz6B3UWpORyydYLfWjfYGfF4v2i0Gr6CEcAMu
5lHyIu8ihmgAHpUrqqDdwcIrDh0FSkdG2eWU562htn7+Rx/lCJl2qmD/tfrFTDa7
hBx/61G92O9/z64aQSgbf9ZxUtChqHRsF8PjS0G6aaDuQttL/ynP0AzfgvTb9k55
Y6d1h/lOoyRtgItM2xS/+SyFjATNtkwkCvDzwoSePYBh6joucR7n58akvP8sRuHT
cyNB4CiJy1NUy8CEynakRKCLEMH6zdKJMKRckxI2YMVzjzzhZxNrsynWlFzfvFSx
ToZLk+MWjeMv5wx+5AM6R9L5ORMtGB2aPKjMCQHzpPi3QDcUpNGIDixI6ewoctHC
1v1/Immg5bcZzcdtJeE0saXktaCSHBw142eIHQOFcX0GAayt5R3+0LpHdokCu74I
8y7GyJhn0qz+PUQnG0GbHEY8vpEwPw16LCheDaX4zzx9+LbHi+lyG6KsmbvWVg2U
XSzyXr8uzH5K4cTbXnj5IjR9pEcFkc0o89ad5WqxbXp4GKJtAl49ypWI5YVz5ZgZ
0dGc/9kOWnd5OJj4adVKk+jQ6AvokYT1ilDIW28D2jypuDH+0o0okYK2BpV0Zekl
LhKYJdcpK636ym9AkXhyy0eOdQgLOY6DehB8+Gf4V/aHkk3x49s+oS9ifnhgismL
VOPAzb1PDapGEGqdOKtC7uWlDUo81XMLtfwx3y2Z1mzSCLHPdsvveJtj6E4HO3y2
qfdmBjHwWL5ItOVUEyGdhDgonglloJhj0QkBMURyLo6Je5E55Rv2DVCOud/uxO71
SpF3QjBQKmdom71agDO6agZ42izxr9Y5d4aZSslQ1/UPgiuJkKoVKnuypn0M4SOs
VMfEX4Etl/Dt8SBCPoYk4t29xiyKSDrbjxcxsRMdlHveOu9lc0IHLC6PJwxQQATM
1Vou1wJfwlL98ZllUkv39aUnJOZ6rhROS3IPGPVnPszTESOOvbgLgMRBoYZnCneq
4HsXedlLgfQepuj5I6+/jgH2PGrSPbkOrGbRX4Pg3aqoB7PtatWFCdhX9DUE4bj3
8B4VuAT+DMZr+jFXHptXRltdrGKndIT/cyNI6esNDK2eX9K8jCsSc7PQV/0GarhJ
m5n+AP3o3ro9nMCAMAL0KIqWWYGaxhCXvR0kjIFtvb8FkUhKeIgZvXr0kmYflYUm
+kVM6urT1JzilzD/Nc78u859YoHo9VvoSZl173qjMfT/bqNRox9iuXtwHdN99XRk
iwWuuUyiipOca/PuEgTcOrRrYwEmJ6XyBL+VeyZ6z/Z5++YiIGJT1nQg40xrU7rI
04WiN+DmOmHD4XxIa5phOZDJURdsXFK9GNASk+hMvjhBh6YGosAp1vynOGXqY/JE
YFbjpmFzPQbIcsFRMX7s1g6RlGZdmys9V8T4qg8H8P5mWDaeaDu1CBAr939G6CEe
WICZ05Nn6ptB8zstIPjez0Ojh9+rqEzpo1J0RiKYdbKP5gcHHkIUL8SDMLC/Fvx4
2iJF+ddpIXeT5kFJIfKbUepLd8MbNnE78tMMABn8g+1x/NoTZgNTsoYtUETmGIFt
gzIwRW+3Tp7+WV388DIP4glo85kMD6D7+JI3xiMdGKj+6ysD5h9AfTAQoWf+Sgnj
qeJ4feAVbeAABRLOTwePClhh/hZ0i00/l9yhQTPaxuCbpJyPLw6CGnC1serpKBhu
AeqeB0qfq6a27JHBYbJjiIPyMKGXATbpMFq4VVUyRWXI2oCvRkppZRSiobV07qy4
SxZ+FxeR6G7gYuFFuhqnbChar2gB9yyUXPXS3bLA5+CE9tF59WDR00BspmpRmlmn
+nmzexz42aAgP7K3FYgavB5gqRzHcT3sgMWsVpuQnFdnoAN9eYlP9B5d3xoPjb1u
ohG+yimFRttbR1Rozsrgu+yxq/vOcHr/z6WVfEjUALk9A6RyjYIATuWRTz9mA/te
6323Fx9kvLFB90PnbVLjBgYNLaHLSnqaPOfDzgwiWSnpEDql6PnCLFVXRS0Hft7T
bOx1r6Ah5TNI6OOIYpLrK+AalMLcxh+7r7Ehitiz8eexuHFUmp59Kjm0VnRwzeo0
sypPkb8QHnNXw/nMqn8j1NjeYaO+SwgyBEsmGIjFcd0KmCeiNbaV56Hr5oWWuQTw
zQT8wczJSZ9olmBCOo9z+93DUBnLT61F9lutErGUlHxKdQ87gE9pqyUj7hH3sbnK
JHIX1IK2AnsUx6eJeTYArs9VJiKxODOdDiDs5RI1+OJfqS4IJV0udUfc2q7bCUJs
sojNawE9//ffzqjnJJrad77cEGIDx48sr0F9VCi6l4PqArq+iOzJB0em3dhEB6dx
CUALpeFryXzvDdoowPrkLVO7n9A0GLGt3fKFTa7sddlJyZovTDoRH5riP0Jsu1pb
cBxq+rsockl9mP5uaABbr7lO1yxFsBXAQMC6R3GmNjFYzHmiSwl2im4eIBCT0HNQ
QS6xim3Z9SCzkgEkfoyxY3hVSsLRY93BljYYj3fRPznDddjgi1QVSlRxQDrO69Nv
7HAiayy+8PvqOxRZTHlVovyGtD1Hpj0oDcdyx4LkxpJV8Swffz1ImyMC6MKQpnS4
iLSVrot7mL5BSWicuXQhY5FQ4JG94durn4144FcD7k8RErxtin75WUzSW7CN+MMb
8atl5EtDBVc59p937SEFqCW6ZmNuoqfiBXfkdgEFOoBtDEYeqwdY1vffUjZ8w68w
zTMjhYu4PVvGyVk83rlpnq+pLy4ArYjasELE1ZjL3EyQ9rFNPRwFTBShbHy0+0wM
GBMdoWkXRILsMWoWdivGEL8zEpD1wvMiH3jsVONsHEHzshT2dk9tT2E+/Y1Hbjrx
ljMBcUwQi7TSm8jXwfhUkbj+wxxZjksT8aVB1l0IXxe5h4HARbywv8yJD8KMXSv1
E8k2A3GxbukBdjB1WmLRItZyp3A526oNVTlblI7IrfGYen/F/7OWBHjr95xzAjsu
GM5aRp543p52GK5Q9W9j289esw2qjQkAe9YRqNNsmOBc+bZlbyZKfDUj/1bIyG4R
9yHB1tgyZPqQQQQk2eHvAMRENqdcOYe7LROUf76A5gBNYvcFuA2h1TGMriRbeRu9
qYsvVf52AWWiQYrW9cO2qd8UlPtjzn1v46RRQnYknjTb3M3/4vi4Tf3+RDaeuXDq
+mAtu8KKDSFcodV73teMbQGph9My5lXSlyXgHjfIc5QOdEmlbcHEEr/q7J49uE2x
IC/msmWDu/eycr4tm5zYJr6T7Zo3/7nlqgL9/nkyviB9a0v23Lcz9pSZMITELfTE
QA+FERcP3+aqdieg7Ro6b1pGJyGPi9IXY8ejdc3Ftrpw+CmrMr5B1GDCZPW2qnkb
NVV9hbZOs2V+7j3NhEPaLT7Z9gT0GLRBEeVNOheeI7IIwms5nNfM/OhK245wAxNC
NTU1sFDbA5Y6vsxP1qPxplaTqX5QkRe+8zazpdHIJYxawAP1fY6fq9hbyQBk934F
7yx3U87+5FsA3kOPB5WeKsUSmNeouXHxQmlPwWADXVqgPRQyGQMlKwLDGY1WNt9z
Ox576cbvSmdD9V5GwoNL8VgSOanOLmiIR3n3ktwJs4H45s6UjpT8QA1znG7UHitG
3FKzC0101igcVkDMKTn1ARt5AZXAMnDBqil43cDWDI5NF+tU3ECMPhKbYJ4Ao/6a
d7AE+fL4NWUdEyXhlBL/UVFQFlB3C2gEczADxMsmRjm3+70tCrk9ICMWzzbr2b85
z1+XZspKCo/5njcLDTvK+r0BFS8fyahysvmVYE+Ilw4Ij9Fh0t+BhivQ6C8pP8tP
P1s96zNa0gcmd2rLkvRynJP77UTC17h9jAE+BS/wQPstDWpsjP279U8ci/m8sG0v
QGq7DKTJLsrA7jXMnuJhzQzn8/Ki9kq+rQqJSUmeSwrQekAJk6D3wwZHZHBsIHIX
XZlitpbM36QJsoweR9M80FTt+KGobPcK+w7Sp6hZAYkrQrewXdbq8gSNXuWJR3kN
mExIBvezCQKRpZhofbd5pLnZ2kjWWVFLN1gP+N6B6LnQcZacvA2zfzP2rV1JGzpN
qzgq+LUnUN0GpGidw/gdChkUs2/AP35yNAUCtbBtABx3ozA8jJ8yQTlZQ+1TYtJk
AvihpyGvbepj5Vfm/B+kZ+r0Yl7nyccTAZbf3t+IAuYJptfHHledCM1MggmOVlHB
d2Am8MnYNHLvhbS7oYQL01tCSt2rJRWST1LMKLQQTnZ8V/T7e6BWW9ZTg9pve+V9
1JafE7J2HuSGKdqQmgDQZiTftMGmBA8NotCQY1tBO4mvJg4N6ChtShQEk133tD9k
PPwzaLIFL9x0KgECfAIXlsD/KsBrrmFviBbnDv6osinYwVoV+sxDzEc1AweOsVCZ
OdFWKNCMoQ1T+gyWAHz2blktjG7BYGkuhyuDqSghbWicV/nLLxIwLJW3l7uAHId8
ps1UlRJxyJmJX1y+KQ7HL3SvqbicUTyI+ZCKrcITwQQZeuBxSKa1ka06oVA6zzNe
VjY+uELI5FimVq6E+y7txqv/7K9kDLX5xdSyxUtAmc1q14yyuiUGSz9wNIKQfO60
qr9qeBGtHKpJtOATJPBRMNuwZA1P7qwFSEMv/ShnSiTx2UvUdbUZFhyB/AiGokKt
lEVJtZ3hmLFOgU78nCaTYjyB2eW6GjrBNqDCe51go8XsmQwaBE95/O6J9CHC+zKS
BiHtoucopPlP+t1l+qoy/rASPE8L93STS5b33IFHZ/D0FvwMxv8FJtXMXan2y/SL
tsTGTi6j1Yah0coU7pMgLMNSo7J7f135Uy7Ckhz8Eo62bEclEKR1gNtRLjh5P0NA
y0ZwjnvNdh/OE3b6OryQTNR/JhQb5aVTky85o9xUnh0trwz/44YUvGloHY7GOQWU
KZMMGrtBL5YpZpa9sOF29iPxfVs+TgK1IP90nFji2bRK3zED1aVCnrSJ8HMO9P4d
KeeDMFfGRdaCf4jlWKqXeL7/T9xNDI3sd9OGZCHIXoe0MgBTzMG251qOlFj4M2IC
EH1gejajyyA72SARtazR7+mTcMP3kp+p2Fo4CKBAV3aF0v7vqlflZZnLoNgFGWJM
6M8yI2WiaLI0VkqodHauqZyQbm21u4PWDgfhMsddZXQIINsd1o2mtRzOROKcHDLZ
XNeyK1X56ddiBetk2WUC4O4ROp59ZuWkxWr1s/xg/NSpPFsnsAbkdNBUHUwjSK+m
+V73CgTM2g3YnnHr/gQ59oRQkQ5oBAMBsFM6UH3XiBLdGzHdEvQmu9E/BwbbXtlv
UjqiA8T59JPvaw1pOn/XlHntKetAg7DyS3tB/4VH7ZvGsnZ4JwBRyu5YdSdv9mDM
DMLfz7fkdQtAMEWc2QZ4/xeXog2BGjQAgNI0IdB+obQz+1D+WdDKtaHOJ5rQpzNS
AXoKGJLMF1DkbWT5c4bSDzdEP1ZAC8BOLl437hkldx0Vc/Qs85uiFvnno5c76kmO
wzBU6eG0xjSkzSEwJBMv/hNjSTmASL4L5vcOxAshFY/ie3XtatGEgqwOj+zzg3w+
nl1wa3zVh+liAE91U0I34McI3FdNvkzqWexlab9BuVFMfjo1kXSNi879d2UfSCyF
nlHW4039CzZywLoFxiQZEdtv/oXrAtsRWh/rbOnxT0WO77kLKC2O+Hz8XxtmGrNE
MmJnqkg+IUAZo67Isz5l9KhN/RnllqlSIfOQv0NMD2MG2KAkjDVOFze0Ti3qMdRQ
R8ORCwTkA5cf09ibz0AXnl+GtfSkEVeRH5eaROgPXHBLZX+UIkrIzmZmbGxICSRP
8r2z+4xKYaq3Od7KWPOvy2ugtkEWohO+8cDZOZGEQRH0tpasMooAPtMyQ2wPDTLb
6rXyRuN9H3mI/6aTMSlZzB2UxW2SsHyNCcZDvnK1JqnFkMd45g4Gc16nqRhtWc3R
yOCnVkqrBCMUmvLdeAhXGDO73V4kG+yXAF7bVda/xYSpqjBQVfzBlUQLhEI8MNOF
kr0mtZ6DGRBybgTemX08MFfk9cq5CWitwFyFeIvUid5R4+LfoyfAAyVIRwRS+ez/
0hOenimxeVySN4r48LzKtCawHqAQKVrNJnDi8FLg81I8HHABuM/pSqHT0zImMekV
9fV6BMBermAhRxTq0mK0mZNv+I6ygeHU5H2UWCjjyg1EADcpe1cOCvIqG3k+dszL
tnrZTz5jVSBQ9q2DwdwAVs7UA7Z64w0OwndjqWjEVXI2YpW27Kro7GfPd9kjXxTL
gIpThO3gz6QyOU4GgFhrCKbnWAfdjjPBrLJi8j+LBkOeP5LL0j5brtOZ9R9l3iDi
YdR8tizu9gz6ZRgDhyqjQS7rsit/SxW1AElXRaXB7oEeNihkBdI73eWCIsXJ7XmV
daraJWg7cLhmMlN/dzerfcz3MNmiuoVzZBypOLtwCMh2iwu0BjOUI2FmaADOO1V0
4GKuW+md+or+uSAg6idaCkwWSmVxRHuOnOeNEcEMP5fBYKKz884hnpbx7XFs2/1P
K4b4KaBVb1kfnlBweOeDT3Vw8fB2NeijChWmU5mYAOpWSKZg9oljlfBl/NjT8U5k
htMRff3ts31OdiC0K1mxIteu2If8uSWI3PJrnXXBLikzuYQ/khwyY4PNgJX0oXNZ
uMoI11dVXo0WxZBXrHMBPh3cxi8hEm7gSlhdSQBaNrkPAbqfRj98jUIU3Lwty8i+
1P9G7yG3fj8AqNSSuwsnQNTmUNyzl4ARW6sukvvCV/k8TxC6kaeUh2cyMjnwcMC4
Lnr+h8KGCeXl1WCwsuKlX+PdcPRi0e0yRKkMiLLyz4E81Gcmj6OwjVx6xdMlT4oT
r8S3xf7+Rnsu3s6YNp9y9xjSC6xRu6NMqAc2Ot9WSMV/37W+57wfF/75A64GpPDS
WoNKm80CNZtJsEMUTNQNB0SDwAVRLWZB24LrZEc+DDEl7ZfwxXvc1mJbVSCv7i0f
4WFpTKmZePYKBMO9g/mKui0qPFEGXgfjMUtusK32PEsZNu4sakwET/1nDyT2r5LO
ZqVxtOKujR/y0Wwh+V6eQkSoL7a79bCVvIeWrhXmDHgdwoLpW0PKnc1/xFsmiJxz
gf3eH2s7Y6Ds3656XZcm+QfXRX2J1drhRB4WPbyQO7nRzcYVVki41WyvyYIFJSix
xOKAW/Xa2AgHEeOrUwt+L1TtBz7xwp3ReDOeU8ykFNu8yQlpAQQcFDc9KQIvBpBm
rWlcb3Q5EIGPBXDPlPktQ6u7CjECxQyQ6DgZxTcQ4WTF9aBmhHyWv5tOadVPzPWQ
CImoBPDNdzdw3cnv/KjhzgMySnB7Rp+k6gqUhH9q98W1OAENidurQ0jSmgXK2arL
QohN8d9nxbmUnYRAklw+oFaT06cgI4afevTznCGTSQuWvMtPTfcnJuiiczUL4VTX
W1O0nTulImSwaTiUlY/g000YJ0hYiMWBesl6CG1LfAW7oeYa05nz8BKIBP4hfXQa
bVppM6XJnmHKm+TRyYAerG2wTtf6rXYn9kFam8k6jFlpc00lc55+dUV7vTHKMsYK
NkARiUCWf5/hBy+zotkKI08Fi1SXOeRojjMxnlRG9DcqjQ/KuP4ybHyAcxDYvQoJ
20dLttHmOhJCgwySF3OID+DSaq5xmzLSUl4lhiPEzEjsH4Ki8lSCgmQswRXmbd+7
chDMbaRLcTiRT88mgN7cjSh2jWKrFW+ikpI0Z3kvBi4DQ2Rq08QqZe2bEjMcmdSW
3gZdfcSQ8Pvf8pRvt8D5z4RTciMs4nXuctjfRANI525iZ3EppCMfEzSvPSvEls48
pS55GmMSqfnMtDake6VesabZA+O+wwtWRg9y4IP+MSssviqcgS21WDbwODuOtLSm
lk/m6f14CUpMuZZhN4ltihohAVjhDnUsbdyQqTxVZRex6fz3J2h0zS8d9JQB8/wx
/V+nHL28H3ccvm74cvBLhIFcyK4XnHTLls/3AbWN0kJ+XlyIb5D7RIsb2FNovsNZ
RCkQsZBPGS6xsw6FLZT2Qj0C5KEzgkZd4Z5Ezm5P/PSb8lwIo3IGutzkt66/bkSo
+B8gdID+BpukAVKe4qaN26MswXvChY33ZrRL9b3TjlJj58dCvbuRvOZd/CWFmq+/
P9N87MncFT2Kw2lHOGEQmMxdSkW8tJdaZjr8GyyhKm10xGd9vMWkSm7JeyeqfwAC
Yl8euiN0hY1PLBu22OdgTTsejjZmaM8iVvSNIhLG/d5Z3xOhzRkS4tD7Z9Eix0VL
IPYn3rhM+q+1Q05uBHgKoDLLuXOjejsRsEJReEJ0kl3q2goldbEzEwCNMG+UFdTS
OczDGyE8Jy97bt5B33Kk0xAl0EdqtjADbBx/MF/1Qvy0tgi0rvdYrA8TiMjVDPHd
gOqROkzTzolx6L5/6Fd3EEoT0TKGAjRLooMiOhVOOvyboVP1vEEZF4I0Du4N8WBX
IxSHTrX00HwfJ7iHRSWgXrfwGUnJAUqxRYfWCvQrB0oChurDVIszQZHCyi56y8Lt
cebBm0VezLGWWMmY4cyixpi915DRU+0QbbX8evs4dAmmih59FFcaUEZoa7tsmAhf
ejlEcc0WXUhKXXYq2XD/lmVp7eR3oIOw6FT/mHIpyGkl5EIsJJoFH3o/Rh9YUeew
fU9y0y4M6xj0c9YrHyFXoAJGULI2Ol8MEUk67NyRgTznGZqdIUBoctA0dsVmE1LM
4NoPfBDbUY1NP+ls02qBWH4ffJB5IsDERxGeKdy71eG/eOoLHdj6nBEXw7Xno2u/
qxcnVO8tGNyYY9NHmeyERr4f56zD/R+xBPn+U16ojwn+BpUUOrn8D0EzBS4IVCaA
gcmu+g40xnj5Eo2Svc9I708YVhi9y6umz9P/tDMMtQfCJ5AQ+uZpIhUTYMl1Fjfz
9hEZZ92Nm/ZZ0/6jINmLC7j5Rtj1olFmXkPEOPsOLe/J6WyJb192UnT+TOmKyTro
GSFf0QYb5DC+wZcR4WuoxoTcJ5zfX4bOW8WBv0LbSt76gvAkHDpJHPZlBb8SY0xV
n0i6Mp9TUAa898dbtCJvNyjcLuT8C1nY/gz4mBpjajC4HF3+zkj5h97KDeZnCerC
i7yKFUvGM57JAqHs3zJdKIgRjp0Nm2XTUAGvdt9bPjyu/t2s0nDcsQpqhvaAoOx1
l52p4fPdhW5V1Sb82N/HXeqBpGacgx0FFOMXxOhXvsvyDlz+dCJWGWWlQWeLeH9a
ssRvSRRZXIgxYGmDw10RrRGFkuBekkxntno6ARDGXaQlu1heVP96eZUvTAKoitCR
fw9Pyn5GLJN298g6aLDqZZ4Dbo12FND1cmymNlARDGz6KWh7oSt7CG+yb2OHtQGC
aDy1C6IWVl/YcJx7NyBR32WpkscckCrK5BbeLKZWI2IxtMyPFdYl1tWpM4giL4sm
YcIqgGSRabf6M8Huf9qFmYyZbrdhpecbA3IRsdZCvMx7zNVa0fwfehm0C1+Te7eO
XYFazPeAtnkHIKV+YogFd5gErmx8nHtGqPjMgZ8sE1on2ZDzPyhyLa8rE5exu5rT
UAAJ+QcJSuMhHa5OpjJMzGcgfGYMD5JHs+gpGrSGWpeGUOI73WeTQeqn01JOVUDi
UDWDKZWLk88YiYrd0JVQsZe2y1fWkIYCugPueahLNQkLSOEN7+I5w2su8CuAchNx
Ju1RpqnrVcDmPBVSQUHY8vgtFL+YWrdD3ZBUCLtPo6CG8epu3gxeDEz6z315lNRI
R6aqpgfuQDnCetFQecrxiG2yPaETUGDFgLisEB/WPzxUELNEXQIbLCj7BzaOhKAz
nJtETGZ3TWFAMFW2iac/LZa3Ph5no309fyXt3cGQB66Xb4wjtpaGtAnDPgk51CC9
RGXyJLwMGa6f8poVoVAGxVhKGmaf/pvRqZPe1Hewte9CWHQhwBbPtR73xLMbqDnL
VXQ9zjXmU/FCcb4R/Mx2iuhKJhSrTIu5MLUEEW51nS5PfUNgsdjqZvYlZM4QIF3q
4bmTBpEYDphqm6ZY4GE52jXT3BLGLiJ+v0s9Sn6kFyhZObVf0l7l9igHxznaEXxc
Fd9yR2NlcHDLQQwZy5cDvXuN5GGtHu0aPa89W2Nx8uyFcq//47Ct/66kzYqtexKF
GDIO89eNrKQUwNaYlLlSNgOLGhAjrwWEk8lmnPiFSvdN7Az3eSRw+H99QXAVjOTL
EGWBRoqS2S5WK5mWm1kLPCTMfVyqW3Dl9WCAxFA+cH5mmGaFl265dYcBvhMS0fdW
df06mw5WWGv5EFmtfPcKyZCsheIv7B5E0c9DSlJibDxNrnzVcxJG3+ppUKh8Ueba
p9Gwb2NEbu7le258e2vO9sQM2BrSWax+Xnz8sSuNCymD53q7mudC1d1SiEzpUpSj
RQRi934IExkVH8jzWvrYFfCz/VHcuDQMPG9h3QR7xQnxkg5hQq0IdhEISFN18V4E
+EkOB2uASDdtgwVbK3WWpjOUdEDJZ+YbNmTOH+rj1mMSVS+uEg1vuIw1/1gwPx7r
BCdD7FLFYeIjwMPVgY8EKxmGj6txXtsZvwJgkSLBgPFoz24V7Ju5COOFP7mjHlvr
GnKyAJOBvMte/QYSbKlUD+MDsljWONSsNdVKAc8YfQtgyInT38tN+1mhm2lmE+S/
5q9688nvnAQ7R4aGrkLJCl+/kHymJe2ylXhmycMVryIVmcWkI5kKL1KGsU5Bz/hs
bk4PH2jxU7UoRFzhoIPwFtvcJKl19kKVcL6onkCjR7e7wVK+vVeZNAgD3EGM2qNJ
fEVspJBGvPFb5G09BFNII9PkoMmwmAt6JpqaJMrr4SY1PbKsbNo4YF5kY7O0T5VH
HBB+jy0xdUd6mNUy4Fn6UFien+1Mya84lAQGcYAtYroh2OG2CUOsO4w5H6HymVT8
jYGzCt9BJT6G0aAESah/Z5fB7nyAK6KmueBifCHRzkyRdMftDAUdjNvf2r+CTFNX
McN/9bWaOy7/S7bkU9D0A6AiyEbRTixXieIyWcy/G1n8OYmYkkc2mJAREyJTwhfY
OqD2vheTistp+SeWBfscGXmCtWPdmOwjR8JCFpywRGSzH5fiu+NzrFR2arLSEd4K
t3aGylcdF6pK4e9IxD/IC1QE1gxSD6MT7/I1KaABKJUjf9awN3/Vop/vZhTBWbq8
Sy5WR1WLM2g8GsN3HPpO4dLjjvMu3h37XseUQUNfk8gj61Uv9YTJ18z4iH+oGtDF
oBkm/+Dz3v9P0ygWqyCsn6/3vCIDGKGxzA2PsUmNU3fCkZhSnh3sFeXXgREiOjb2
vvwWJ/0t6UumkxF3GZlgO2QkX+pQdt4SDDP7HZaP8JgtIQ3L9sGpSnHHOgWT+Mlo
JYe//OOP2lhIJgs+7nBy1SBYbBewSFxL1P04A3RRyAEQwiUWRChd5MZ1ukPtgUPR
F/EkNaAdt5C0jEofscVmwQJc2zAIcvyLCVg+M18/BBsQI1geesWr8l15sTcBNoIb
CymTjRHF9EU7xDIZ7yUdgUlgQ6izHo2/9EfSmqQkePgdZWY63LYHRw5e1C7JON0T
OtBF7R+qCVy85iqkp3d6M2lDJkcCIKsvyPZ7vLQBBkIpIwAMpCJ/eP01UGvk8gpB
O5hgIg6ycHHwabc/z9YKUvM6EzhuvYRzUqkasBIUc4bgTOCCP1Yk82TedDydDr+3
BYKVJc3gxNi1yPJh78BI+R5+5JlSF0GxpZ1SQ31OYM9MK0eHn2MQCuvhXQhrRW0G
BVsQp4Ku/eL4abPRBVxoQO9vma8xcvqdzgxpxFnX//ysvO//fTllz3Pn7pRqX/XW
GyT9QSjDjbI3niZHF2gYe6AR0vSjObDbXZkek6bvsaIzXWZ67eB7MnUoQE+Urnoy
qWQX0x/XEepJdeeQWN09K+0pD2hoswrA/j2t42BqCcssTcNYdISlAL4DCPkl5Pir
swksaDT9JgVuHfNSBwxIBjZNt4fb4gIFeJo+gJVWv5/vYffsDRuRrfYZf3QINpAo
BxfofobN7Ui8HBTs+Lh5rmQli0oF6cAe1SvVNvo8j1YtHoJkaO/x+xnTrTBsL6E0
VbVGeux0+xhMbsVuSu+ywZ5MPbQJzxHLVFPUwZfcYcVFdqfguAXqyNvozxWKCAn+
Kx1oqIJbA6RhqXXXA6jHeXnujnexQkopTXVOzkv9gMlH0Rr4MqB5nF4F1oI1/tjk
DaoqfFOuSWjrb6UOixvOzVu+JHKq/B8tvN2En9pPE6wOtfOzEPREBDUNljRh4uCG
iDxS+nXdJvh1yGHRZlzyiWfp3rYCVrLoMmvYXT74mb7wWFq9gao0NzVoSOxgHETR
TGOHkg3ccXmQzzR8udzZ6jNZYxu+ChV7rVKPhX5VpC1IjTKvKjKX2uj3fUJfyBr/
6Tx+vUDTiJ+WuUf+J0DBYW3jgXVjOeTagXasWRrLcnNaVF0nXdhrvo0NFIVoeTzW
pijCNggJjy7vLvohF9sWzuv3va7C1FBD8XcEsec7T9/Q44jt52g+RuuMoweqsa3L
DzBEnBq7dIoBbiwb2O7YdgVZB0A7wYS4gR3V9jQr0nTzmt+4uy/C4hzqHFzadgYq
Y0JP5kussky9Zheum81P+rlyletbXU8oVMgcAkE7EMCISr0HbJ9vyljpxZWcJ5lk
b4O5Eop9iEY22LLLQDFiN9XYwb2Ue7M5wjrKeC0xi8UyTldEV3ENj9TtORhohhB+
GG9tjMIlaQfzSAmae9Qtw2KLaRUHW4loshFgi+fmBiEhu2BH+ZGcR9nBUCbnbgOo
RajzOMV5j629q9w2MtMjVLiaSvU2h+1Kg3W9DQpGV7t2sC5a4jOpP+6qDW1qgVB2
4Z7B/N5letSSEmLKDhlqCsQs0ZHmmBADKpC4HUO7Tooq1V1oqeI66IcWGSV45mVh
Zn3ynpg289mfbImA2nh0BvEjeo7cbWbL1q8kRVHukiF/4TfjTzi1ki8cOJ6As4vg
MJ+D3Nsm0PU7E1uQmHjkAcGt+AaTKIsfcR/GFxjSSQcpdGrKPP5VdBr7SX0y9oJy
uYqhk435Lu21BnCMpTUUNP09SLUZW9IEMUZUMGdKvERFZeR1fh/zV83iOfxBVr4g
hkTa2GDqYZRtcjnu3OREVE3NfOTreRH0cH2H+Qoa8XvpOWKXmuQZRCudeBP2z9Nf
A9WhA/xpQD6kqzo/Dx9RvYq5gtO2X4njbc6sbfFkJCTehdrtuSe/4ExG6jxD5nRO
2BdfFl2/K4Mc3FRn9fNqNXAVaaD6KshExd4ZLJ8xYoPN83/SCorRKg5UOJn2LSs2
HRvsS8x7eNFDx/agSEitUcrIYvCY5wBKHgMvGnq0iixqVekAn7OrmVAEVJMEbgw3
wDFrCAk6u7vphxWwUJe4uwkcYs5aBs08zPyljuXBibRiiqB71XllvLbSoSl17lWI
tMFxUnPRvXb19I+Fc1KYE/4ALzR2GaaQI3Zw3CWuqWJrMuwCVAP8PoCQEOA2om7+
dplyiGrg26LP635hBwykrlKisv1Zm6OJv0MGSGpHuesN/4h/nGxYqiSkUGCawiit
uWMORvm6NcowxydReZPxhDFCZqPRFFzof8oVe6a7owImpUbkmhXZdrZ3+qyADSSw
/1rF44gHe6UNZUyAbeDjJyG899DaeGXOqR3iwZ2eo9388eRNtBgFK2H+z3++A1C9
tlavSz4/+lZUhBmkOi07Ib27jRXuDE8xjVa+otDw13yWZUavdeRqf/TdWpAzoF4G
Gn8cj+D+NsnVnKehndsez4Jjy57vh5rJpE70+8mmLijje04zTcnr5hKt740pIRVh
NIWc1g2M9r7g7pyYeAO0HkcbpG+bUGzcflbxisRZH9tzhyb5E4bNKiifrZg3zzs2
/+QA/pwr2+/J5C0qgOlJ4C9vvKpCzXfaYvdWZEgi4TyJqodOMwyFGVa0s2ppd+wz
0GrwW1+Rn6J8RtOkJq9ZlntZRw698h0RZdV6+hSiUDQ13ADXh44s1V2QXizWLuWJ
ga4RVBlGiR9NDuoEtUQTyuXqaDBOIu7btu4NqDQr/SqS/4rc7sMIqqSF05zuQUf1
nOE+DbUK5D6DjeVy1V1TcyVn0EX352Ei8G3jY1SgbaXyYPAlKgmScU1ZXbipWhft
s/fFZLzau5Jlkr9BqoCLdLs3+T/eI92MsVOZv4oXDIXIKxgMwJx84OlMqqpN/DaL
U0j62dhnpTGrdmuBWcmGmXlaybGbJgxPFwYatgtUPFJinTqRacKgsE4yvubPIgxX
pJabWa/Txb4cV9kFlzE4bvVcWTLqqgFl3DAJOkIh50mBGclMJIeA+TfpJleBehAj
gvI+FiZDF17gPkls88VEn2/ifdwPMLilZ6vnZsNB6wq4iD0WgJ9DNSkwGv6HtDXH
nEAybRn6DwPlva1evGqWjtr1GGB5JgiKwBifERvejY8dpEYj1r3l5Mts4JXbuW7Y
MW1mK35MMme6KVgOp2+cO48JTFFxBfR8kQvF+cGdL1sVpFdZdTw9kxxALZBrbHeY
ppLOHUKLMlvUjyFxMNs83NvSOP0TYaNX0Z13vrwv26lJ63TW9HIwojMUA9ql86fp
w+6Nb7TIB1HFwCq1ra06EfHpRnn5o7iEc2wCTxNSniDlCdjdgAm9CTDbs54WVMN2
8/Iytp+n/Cj3yaGoiA1oecmnQdRdSZKnl0eycjWYhGFBr3a0NLv5u62dlUhh4yKL
L63m1XFEY6zwsKdIVkXo0GCgmYIrcJfZr6Mura+BFso1qj9bxl/PgLDRheS7F7P9
AQa6FY7Vnnuvd7I6CGq2aSwdq8UKC8qkSfCxg17mZOfdYLmHQRtLgank/Xxdc4I2
dDBG848PACFiU2Q3CLCSCA1KwSDVTW0r3wu8R0BgSAtLfj+7vhFvESUZoUBypCaf
284IWq0tb7bTxHWZW/Mh3lRjhv9NIEY64pVjSYKq0ZjGR/g9ATTRsJY5c5QsJrTj
Bbb44gyxFaX2IpqPsWLx9A6EjY0EYp3MfeiVBIe1h5T9A2cKjkh1fizJ69MOxzZK
/Gr6b+wilNVpiQ8r2FKqfRADls3dKax9Yycnsj4XPOR9njiIJPXRffafchrPJlKk
HiX/S/cMkrrnYQ+X/pHQCNJc1aYIkZjWD4QOOZMc1TG7uAxqRDLU8QeKTCXWkZVK
kPyUpolr5nQOFl4m+ZJ0Ty0ZPhfQ//47VL09TP+HFUDUCkEBZv5DohEpK5D8w9Cd
BrYYM+0DmSU0T6abPY4sfFvXTC3ao9RMiXRYMCxLuzNqfJRecHRdKgDc+J6OewQJ
xrFtn2gBJwwi6dhq2laJ4wmBqJqdncv4BdI+iQI21Jk1AJYLcC4G87fIB/XAtRZY
JMn+6NuZ+tQ/5xNxPGLSlwDn1GqBAGhJiPz44DS3LKq4UWntmGFMDMWKGhOaCdbx
Oi+FWEiyQmqVDidByzBMos2KVQ2zljP0aZMzXJcMOlFcj7L2fXXOPCyFbPU9TNEA
bySJ4hV1beRWOlxlAI1Q2GB7PhKmIgbZH4yVDGNT/tvL6/c2hHmKFQtQj918i7RJ
n04vbUuZwA+7Ui8uaObnOGInb0do+GtjQ4gP+oRaGKoeR+XX6qsG09El5dmsrZ48
943GWn4z1ol4f4g9RvLEhzU0ekM5HjQei0J/f0EMhrtqaAzI2zSh3NeMNoUExOIC
E2z/TMeS3yI+khEBEOxAjrsgaYntFB2zbM+RBr/euAM9zIh4/tvDT7B0efRTQM0l
YdY09+OUq29yYiMQl5PqFmSQENDzrx2rdDj3NKaUUDM1VRoX/gLIqAJK9ij7UgME
yBe6T36+6VP8YW0y8hzz3B/1zKlqSY4RDyxMJQ5EsaVk/b4WdI7tkOsEABVOTHSG
id3Z5aeIFHTyYoV+Kh7lSBryjnZ62CLsVZezsWzfMXKxEm1eC83SqfIcTwIc9vQk
W13n3Zd8hwcudKCwt6yflDCYCXbq4LHAUBKtE7MfG8kH02NFWi9Twqcj80pxpRzg
WPMB/SbxQbvhApN2vcujvnmZZOL7oFiBU9/C5hqwbmlW711UvprTfnbP4oYXyTxv
Lb1yG6L632pTlzeRjGYQ50WKoJ2D9yqDNd93CdKLrrtuyZv3OvFtoVcTuiNnCIZw
1YoH+QNNsZ/Lz9s+Q6lNYn7iJ6pNaUYdj5eDw7pJVwaE1KF+FhCqJrkdGWtClsJV
6iyAipJXdnmjwGvNWpaNGAn51bx7MDEMKUACDrCFikPAii8SD039vRDuTYJyzqvQ
Q1K0weDJSGfUGbERsQTPS+9lSpUrsQJkAFN2agF+GuhqichWG85lI6IBARHEihDY
zWv9MKcHEBJOQT2MQ8lSx/JuiSjMJtT3bgawpaos4R2G2t4V1N7GigdimZMHoH24
2ghxjGwAhYs43tk3ZA3Gu04sHbfqo3AGNPV2B0e0RQtwcDwOe2N7NvQ6CtXnooDO
e16tko6DVnyjTQhPQqA+6aQbp/OkyOlIoYolaIfKTILAWd85wDNjOFQK6vH/apFI
stL4JXkUAt9oTUzUQu/MrtGLtlLtpDtWIYgh7uOGJ1nDQZdxfiM8NmW71jjb9uUC
OH33K7fUY2fvRB2QSuIIzn1mfqifosY0OMyjljYNqOpWPkoC7eJw3jWHYJw2zBa2
BOfDRSzS517+o7dEVPfbWp6hxL+qxBXVz19xVSpV73YrJVMC2SqKXVW1CKzGde51
87TtyJqguq7nEmbODk+UmygU4onrXOTaGv8x/FnWXan6staMeE/X59WiBpQq9buu
XF06XFOQ7ixOZTEhzQkW9Xnl+kM+9OjGQLnEL7br3BtaG5FYZS26SWaJ+qwbuSpz
2W/q4Go554lBuXiyaWNJEXENzOnyq9aKt8+zNOVXz8oK8mdix7MU7DGIXc/4ypvg
ZgIeZTQ8NpedVeDSqzDa8hbBh03NCcgGatw1IY2LqJYQQ8HNNw0Erp5PeHVyU0Ol
30Jy3cPhiULTMZF6min8/L39WEUV37+q4M2H1iC1Otelh8PceAX4So7qhseKrmfP
gqE4nd1k7JKBXf08/WWudvfFH16RuYGqrvEmSzZ2PMuQggw/Itqy8mAffEPY3J8z
Aq7NMldWR8awNM3VVm8QSDhqoIxBlvT6P54bNDGJAxF8hCdesxZff68kG40c1VpZ
tKmgpwiGCN/Ize5qiUdl2QZW5CGCE+jBEA4kTywzjFmmKfMvJWAILAr4pHY5wTyp
CrSvT6yegcbhve+4Oxe0hs7DXNCyItP+4FxRTSGXQfWlDc3paBuzktBCC3DLVdMj
PPih0XwYvurPn2npifm/LECw+4xPmWWCpGO7/l/hM1AISPtBOLJyXzudLzgWKuD8
CkCu8XZsezwpShp985aN0T6Os27O4e3TarTP2lr3vNmDeZUMcPbt4ioiDt5TOFyl
Q4B7I/TFEHEpYbbyx64729oylIa68buDcTlAOJJlNPD2sVaK3MlVgQWIFxAY5Wgs
VdHlrd4dn4UbJ1FH7MF1XrHGMhfEXu8PGhwNhLYgYcQeWACwCuXshjBO3wGX4Ha2
EKSn+ewUAkquGhxM5Wux7xzxukO5d03Q5uqwW3GAU+GG4m39qbavhRYLxDG3qofs
B5QFwUrCtGQ8d0bXVF24O8I99ZOQnjOEKAyncqp6RxpFTTgYO6NjP+wfuWCfTr8v
Jmld23v08X7csX8GNKUfqAQA7NUlwHrL0egTL+gZy9jkeABN0g9iNdFprLHB9C0c
ZlTeaEu9nN5HRbwp2PGWE/a62V3lowj/x3PafZxW7MG0XoWb4Olb3HJZd8ls2rYh
7LIvKzgULNYG1D+mJF4+38cDmz5faqGaJid5yR+i1OS8bUtyQNCuc+bijP3AAbyM
LhLvDvSp9pVE7viJnbCNZeVWv4U2if1Q9gVZ/uNNzhyiIbCKb/879VS48219531y
zMkB9J9PTFZj7B3/V2s7L/3DdyRR9hsCdK3fAvD+WSTWkMNpCmXIfNAedgYq+RLI
BQFQVMtfEdJS4oVBBABBYqE4gvIKvOJzYMWsjq4xtnwMyr4yCvyUM3WvEMuGcPQf
rGUlgJLQ1VXHWysWOeAIR7zscDxxO257YfbWHcimMdBxX1E910JKbscTOnioC7MU
r7yQisuWUphw7GeFa0+gN2QxCXHhGoU0PAiiJh+4BTAETUTJ9JhqZnYeBTpubK7K
XRNyvcrNuxWbWsRVMpwHmhw4CpsQHpF4R3XZ/BLNTwYuBX6Jln+ovTqDq4QGEGPm
5rV0OKcmgz0GH0L3+nh0zW82vv45oD24Q02sBSm2Pq/6l7ZH/8Xh0jsyQqEeQuHz
0T27HI2TCdNuESfQtiJId19dMirM+zmH+fz0a5+0Kf8gMB9mxOWoxDfpRfcj3G2H
OIAR9aJ/DogD1cZ9IaockJqexnobU0wDBA/Cl8L46kkBOrtbth7TLv3C9FO36UWm
/L3iptLlTqm9P3XBC2sBwCsjfEntNIRQR+cLg2boamT+4GRxf43l7EtnDMiHFvjM
IZ1ykommflcfcCz4Q8OBTU4y7iSg21AV4GwpCpImXWDNTkJXWkaCDdbfjpd/z03K
h21IXHkLyxbxqBkhSOQO+a4ydnz2SuuTLYdIebU2cQT+c60M/JwFSrfK4Iv8Zf/0
RkqdC8feK8ucwPP24ZqqV9pyRNtL6h5KY02Yi9JSvlEY6Iw5YpRymn7Ewi7umyIi
t9mDxNLQI3ZNQJonRTvvTsUCl8IcE6WZWAsxf+IeNqcNZbtUf5cHTYRJOq8+PBJh
1TgRNd9VuVzfsi7D5BMkAunyxpRe52hBNZYt4AqplDY+Zr3u39sQMWOJWt4Z6d8d
TKP3fHqT+94lRaYUAKBg8x0cy2IrtWQyD+UOjl7Z0NAFZ6qg9Z5WDN1BlRgkI7T8
UEhWyEFeKUkz9Om2DQlZIv62U0olecoYClnzNRNGxTA/rg2bRgbUtKDoDovhReZv
7/wbDOfz4z6sf66DvY0Xr/jV1J934EsIqlylwJlPxjaWx7E6Gz5erdXd4lxTeTAp
uzCfkJl5XksvlYbeqA4Vmv4S3D51tzolzPe39jGr7L/IJj34e85JCsQ6fVRNGM6f
kyKrX2O/hJGeVbOTES+0mFiSwiWaEuyK7WJi2oKZQVulFy4zia/q0Cc6ko3ONK50
O6W+CzgP5kr2r1qtrFXw9Sakl5pplcwbFENjIWnub+WRigli0jQQvynlFYbW8SUI
g+1UBc2CgNxIGZVqf/gG0XxSjT0+YReog+HV12rnXKyThKPATfnQolYhtpoKJ3tc
LBtXbSLVOXkuLeawf5cis6wzGX/yqc2hhO5OSZHBUktfYjnG5goCVfBKPQDZauP5
rgNBwLh9iN6MFAJ2yxs5By/eMl5dHacby2ouXDEY7x+H95Ww0rdrH8UvYr1WFyCJ
elweguD1qPdyjzz4r0HVOIqVa/o4Ala8TUhOSQY9Z02hFmaszrX4DeIxtgu5deAj
caEPufr/JdIUJoBTq3KJJ5eSmIQ5Mqe5rEnqVk3ie+Kx11BaIdOqXoNgb58OId6e
kB+pTXksiBCCbgvCnOj1pT+0PXWsdPbiShg8Dg/TeffFd0tXhlONKvvrUqnqYJzw
IzKHZroLPxfZ/Iiz/OrojIKSBNgBOzhdnHwK0vIQlMVVeM8X9Pb/POJqYHHOWLE/
d1mmNCyHNVb52GVPxEhNHgtptMuFzb3LnRlGzxvzXKX3D9p0JFexzPJtLo8JNS9V
wzYCwK3uOEJgpUA5stAVm4Q5aPuwpI29A3J76lIowg/x08R7kSRI9HNA8BMNhloO
1Apss+qizuaxGCAtGOCjw/JLVrxOVcyL8a/YbEfi9kiK7VLK0gdYzx/EjDQz4+Bu
jTsXkvI2io8UAKE2y1DDRDr7ovCglD01bPXKqZLwKcCnA2mnIxzFnlqHWlmJIQxL
X/KxabOOui07o//ADmrefvHo1IUlpLb8impAOqb0rKEm09l9Y6n9IGzpm7fYhJkL
K59A0iI1GjWUB7SVZVkZTT0j0E5tzW/FBq8Bkqqfd6KpXZFXxJ00wMFwR18PwotY
DcxBFwQv4xhZ1F7r/uz2wu2ViyvTeZxPyQU5D5dL+pDJuegyxdWYIJuebRtLqxdX
Yg2X6aJLJhAz/tXthrRlziudarmIwmLPq9IZN3yBHBrqJtM2iB+DwQh1hBbfo89i
X+keS789e/tEm375KP21Kc8Y57ainxBbARFjamuM+xkTqccfjBYQjt4Bzi5+Pmzo
LuojMXcfwlsJc5Fpph2q6T5/1KPM0BXuFvlukUoP/TvVVL54PRyUslCELx4d3p+D
AW+7EglxMHEYrS7CB8vDVfAruoxm4foetZgqBgl82Kwg7SYSmTHzHAFaVfIsCITf
VcET6EzoHSVdoJjFJyuK8mI8JAaw8TB3xwF41+DQHefznAyULb50ND8dwlMzYST4
f2f5QG72e5GazE5u9+3+/SiEjrf/yyZK1ImCOgpD0lppOwsIUwbtSJ451VDDg/GG
0TbCoz185scMMK0Lprxdw9x9ujfpRxxTLZpHwa8nnLUTt45J7kQ1IhF63YMXVwkE
s5bJxs8b5ZCL3+RdTDMOEC7xHNt1u7HETws4hhLeED8dEF7SC6GIF255tK7PRZr1
/ut+Zs5UuB7iNVabotZPYmiaX8OKSyFPkTQcVKEbUasOP2HYf5KXeT6007dU/Jsl
m7vY4wRmpWDQWg7kJGyhRCj6FNoBy3juJEG9jkSlzpkptL/oAz7w3aoWxEWIs+tt
n+n4SimYsjWk6bTKRZ6qIZ4ccy8dWcVWVHH+yWSlSxtbrfO3E/YqbTdTPiEdsO44
/LgqmwpQTxWtYb8f4moU7oDOcDxOtyaKWjRHSpzIZqxm96N+lwjjYEqHGuCKMz+C
lNhh/UvSWD6sYpJ+H6XGp//A0BS3fdWwRFPU0Ggx0vjg/Ei8QwQf+gB3RCouUm6r
xNK/okH5gh+CzvE6wT9o+vQCZq1neIJyJglC79gMAYucIvV73i9voX7al9C4zrNJ
xkke9L5VwSn1FkjZ4lYL6FHJ80BwppkL8e9wSUrXyAHZ1K+V2IkjzP8amUBKsOSm
KkHdTl1YVl/3HXMDANUL1GDAKw8VqEL80/7fuQ8hAYG6yQ0JMPKwk/0W1KhySVWN
t9HMfHS5ecrUc+ami6bfU5QaI18fN3gbeR9sO6YYvQMSAUDadDftze2g5vdWzMYX
JyW9GG4QPwpKn/BoXn/sRghebYChA/JnaDnY1a8gIkuRL7U8mIB1GguMktancxH3
iZ/X/TJnd8iQFknCHPxcOPQWxjBs/ra30m4DlfyoLOKYLiC8YScEMvaaRP+hJB5G
4gOqGa6zs51oM550y8BxunV0i/oa2GbHFFFfGPCm13kpjdJnkNRTaUKmSPJRWoKF
tAep1EGfb0RAg3Tx81twMWNIBdYJLiZ6jHQoLi0vshL7NxnkeT71YOpjpxc0YvB/
Rl2ljjKZ+5dLL1GJddPcMQA41trS2Zr8xfHyyLOn/ElrMoGO9pE2j+65QLzYqgp4
Qmuhb+/bMBpuhCXE5xusEoMq3SWplG90xywZNCh9ftsfdJLRSQYpXUh8ip5A4kyp
E+u1Qc7k3kIiVivsIKZRn7D/h2Vk3ybnlQ4/ajTKaQL4+RnMJb0KrRagZRtVw7L6
aHA97UcCEG2sa2mxImvDedZ6oeAH/NhZ3JhxNUqgN0/sMkHFlZz7M9/FCdohIgds
HU4xF1sO6Hr4MFoe5Q/+za6Q7UiUEFI/KJK2hv9THXf2J48DhUn3tgRHfVWHvL2s
uySYfcxwKp0jqyGhiV9NOEajbA6Vlu848YcFLEPfcW6Cj21emEsdpfvseOr39EYZ
l5DbLJCRzn1QX6Me/qweufwterXEnmZ7R2ANQcby1n8q5/aGvRQqueLZ+JtFsNWX
Hc6hn6rNShm2rqa20SdVh8dTCvGFy9Ieck+2H8P8u5znlTa1g3rT+XvDe/o4rkAp
nxxhvMWisuk6H61BOsDkxr75DMvokdjlSu+9VFJNPdzS0n6tjJ+6Bfx4QECPl/PM
dkkqOO/cG7q2U6SRScOBIGxvVrdr5ya3bOaKT15fqMS6aYoGnDlj4CctFwVh5w01
sI98cUk0TGwB/mefUUDTCOz6bQStJcOpXWGIwHYRocbKVBI7N/VQH/HEyQ8S1Hkf
IN+m13snRFcuWcHrVxphgmuTPpkDLrP8/27lRYIBS+PUvEXwApAaUZNgsLeM/b+q
8Eypywm28ebgHiwBLC1V7NMt438U1GX86X3pmtMVTGlKTuq1wQHckPlblNNEEu8S
/CqwZ6RclhmEz4//KxqBWFB2OuFRK3v2Mcv4+UrKqzFk7x0UVGZqgY1uIR6b7uE4
k68Tp6eDLT+fDOvmk6tRlGGF1ud+dA6Wx99+ggxVB4jx3mUlbdr/TN2AK2KGtFPQ
+BPLPwF06+RrlzKiZ6SmaknXpeO3P2E0OSdpW9aKbgQw6j6PL0KuPkj0jrrpjcty
DVAc4bDElOtExj9geXM7ssJyY+K9IomU7loAMHcM0xgPmksbXqJGaFcuu/Cyl15Q
6svivMq5wVEEOgFxcqBCfu/ZIUbn3slOttQqCiwfRg+wjvGoz75D5BYGiexQhUzI
VIFJWwgkMqglXGnshsBFDgm5GT3NJnrl36pxChzBgX9pnIMkXwh25bn4QzKB6IU+
dEO3RgA/n7eD1FXsTtL75VSCo9MLVoYEVsdy6lgdXJYHUE4itNs7MKWDpJFQ3tbF
HeW6tkcwRHkZl3J1yXOtSA9GOgI6l98iJIZSwUB9ptZ7ChGoxxIFzX84/rLe+N5I
5/z42E81VvJvsUxCgvg5xcMELJDjen0Ep6byxiM0ehyllTQ/8XGMPCTZP/Hs5dNO
n4xUKFyDAcc7K8y1nUpoSLTmU7B2/hhoB3+KwYSL1fCmySntisy4aVSbx0BwcaLN
SYRpDC8pPXGppdwnuS8vip/coSta0LQ3giDSTsHcApdkTYc0ss85fPT4uGvZ6UKR
iHjx5I5Eu3UOF/UxOPqPisOWiQrwMvsSCSeqWCkZ0Y+wn3KvdJCqmcMJVyusB/+e
C3S5e5b4NFly3b9j8rj64fItZSd493bd3PJqdFct93MJpdmL66QW/RMlFCrhnZxp
SBqcQH77EFN8OD4a/Op0RnsGO5S56C5idcm73HuFF9l7ikLtilzBz6lHSoc/xOdV
LTPh8QsV7SvKNRD3LecSefAbG6C+1Pjx1xQhht4KzERNavfGt3fh6XFmc2gVYGEC
ST5ZXSJx6RnbxJQfiFMnoNFw2DwIkYRODaQowaa7lcZqY8xRDqVzRAorIoEj5hTI
TpILRzZrxQzyw52QjPZNAWZHIjX8Gzr/5Uu7AEHrPHVVgoKzao0bFhqk2GZzBfvX
ukqqYoPeXgHVY8SZ2DaV5YLeqdbLrfc07/X847d82n+IiFipjvHP4YCSAaQSclgv
23VHuEuRfdD82NqObuOxHGRpfm86OoL9lqZtfhNOPnK/cJ1smZtCDR7sMWkZpL96
P0HurHlf/emMazkpi/T2TYm3AdAMmz+ZDvdoJ7B1p7jDwnhLdsrwN3tC+ttz+RDs
DXARdNxEJq7ssZIDzMe8GUwq9mHNk9eFTvpQ/BjQ5vYtupP9URH5kqzei+IwDYQu
mqhASEryT0ikUyhpHQfdBiEv6zr/z40wQb2YFGllNU5Pq8f1sZzAmAoGxo/P4g+/
5j4R9vaxmeSU0OoDRtCjbt0PxAGy8ga7Mb8+s05OAqEf+njInijhZTBtAYkbdKIw
Prgwru2qzNCbdaXtjYhLuFqGDIXKer5dGD9Gmv8pMjjS+kWOV4lua4cN5D10Gx+v
dfRzDVlvu6EZGyj6nkIODxQThLzftwt2/lFR+xB3qMyNHcfPTprcmWM2dYrEmWIn
eVzTUsQOfR8FZ2WyJO/5Pn7QG7LCKlhPdDssMeh1YW8Hz+lbWC3UKj8OrVdeB+Tq
kjgJ7S8NNP0LJmfHqsj3+TyGTHa77r3ojiKXF16MBDGJNxEyMY6doRCM1tjw3d4X
/4BfgTFO6n3tIFtv5biTh/1hPMfEwbx3oztOANChIaHqOLO/9oBcgDaE/txpkdxp
BzYMxNlfzwp2vYbFV69GohFwwG/622QKR8m1o2BS4UDZh9CVXRASs2698RsGusVe
yU0QwhHsy8SopQ67gJnhK1AWVs9el9HotT6KOPysinbB/8/SoDfm+kiG6VRvqXED
XstzWe6KiZpfwYHeHrBuUOOK8WKDQ1uuJCDiy1rYr2zCzXyWHXvub6xkyayBkGI+
ebG72bDM935F9peS1AQ5myUNQDqqhewhkd6tbolpU5mmFmUspaGg0aZmPxGz3e6H
q9qyV2mf7gz9UOLzV9TCAih+bGN26zstP8NISO/VoOvrKVLfgTylKvGCG7JwWCPo
q1J7FYkprkWOo4sTQuTZpiIYTFJCXMHQ0AjhMBcV2Wf7fKpuJmfV1VQ7C9i/mdRa
uoJYS7n6VbquBZllK6mGOL+PFziBAfOnissTGv8u9xWApRZRF2arTy31pSc+IMdr
2nUJN4xi56B7t80G0LOUoSRJ7BPXYMPh3wXld59XG0m0btuUgP4nGwT2Ozjz8VcC
qiTIfrs5JZAXlp+/dQXroeuRTRLOU0BNUrwy/wbwfdZ93+3RXuWKnJ7xaCutjiHv
I8XljDnJJJwaX3whIbAPaFi6U8nBv1rPAgcS3HsR/wjUR9lkTha5ZxbCQx44Bvfz
osFW0b04e21P76uM8E/2LcDaVof+ajWIBdIqwPqHe/hsmDiA/yV8vq12FeuarHf0
PLA4Sqn0R86sLJOVbhQYHhU4XnF6D+PwTouGIHZwAd4skKEyt66B045Q6u7uhAp1
JFLx2quIgjw8IPYcvpnT+6T+Hw3/jU4ntc1TPlOqklTU6389IZ3/ipCB6SCFUwhH
VexQ8vlVqzBRVwcd5Z0xEhEElsDuUgsBZv2S1qarrnzQ5kwRiWUCoEJXiNkbsDtt
UNNh+p472HQFqmXf2ftfvm1LOmOwJN/nnIR9iBwp5WZ4WXiWv8hSK8es50ifG80V
yB5tZA3fvY/EGf81Sc3hnPEibA3Hv/MI21GZjr4VDw8WJnbneB8opnW54MaUFPE4
BGOADjz4RJTVjmh3ySdZ6Et7SluOH46V9NySkWUpbGyooR/4JGMjhthfJ5RV5X1E
3S9otV+Lat6KR2KbmoRJoHI4Gtpch5+bo7XC35XdAALgVnTmi56OZfuHY6aJIgfk
3Rn0Vt+IuAP2VZ0aKdn8r3Ftuy/GbJMW8B9M1sGx3ndDf5PDhazdfTghUyPwudES
OcEHp9ySjr/nK4ZN5FcBncSkdm/vieaL/3nLqmOA+q+3yxeCu1e5PaEq045OkLrL
NcDsJX9/FFbHBMMFoa9RTvkvf23tE5CV0y60ILFLjUS5fMkEY2Ay5hyndUgK4kYy
xwOpXlochawTvG7h2Ri5bVU7NNuy5QF6RGh3CThcItmLdFDhDS4TmJJ8ozvp9+Ub
+hKOIhmWjXrQ934qPUB7dEW9FFj6xbArLfP32K+Flv2YfX/YlLOdK2bSf90ZKc7e
qLrO68mTyERhQ62h8puD797A7OKXgOd2SR0Gidn7KOv4Thfd1mzXgP+TbH/R0TXQ
pLYLvHX0eE0k4qNbOa311zUwo0nIpVcUkqR3FrlIXnlQGtKYx6Fd9fD2AGbXcdwZ
QMYSwKu7mw73WNQHjMxxcU47rqaMbr5uqfRmFfKfN8OsH8ecJITLNjFgDj5XglKM
rlY94gUjpXW9AFniapGcEleVsFC3s83DNeNXbA0DgnD3WZqLcuOiVW/7+xyL0eua
aqC7eKU+rQD1pP8On4BEbqZ/I6L0g09FcyvGZDxNrzOvKIdwaQMoMwSN8j4g4leT
wSAESXb3z7duWkbryHXL6qioWyHuq2Fry+so31f/H4q9ehlpyVxim6iEd5fMkImq
3UQzNX97EfzJPY4b7L8CCCUjdQCJ0Fzx/w/i06MmL0mKnP0g/Fr8vSDL3w/xP7Bl
Gf5WjI+kilnoR6+LJpDHn1HjkxMoM8nJwhDPxwLDVo4Vqfn1mmjR59sWoxUF7fDh
IGMUXoTVenu/FI/Ft2DQED6T/ftJkUKymJF3LoQq98Acc0cKCBCXlIhLhCSlZvgo
aQEU/NxWslvmuso12/M7g+zwpln8ckm/CTsz5U17glPmcTdNvLjOQHVMXKQ+Umdp
mtOLZ6evbOXaORPV2MqTD1QO9nn/yVwZBNACs1lROCJsX09bpdNMxOhqaZ80EtoD
B9j9P3R+C1k/cOBfh57wUFo9nnsKVLWMkaHPCsVA7ywqwtCn2l9hVE38F1osUKi6
qeDVFPowZ08L8OMxJT38xB2mu86ijJWqFff4na6c8DE820i8Xuo97+agB69medqK
ABGqXyzXYbL3OoKbZPbPLLcaDvNanjuffHYJ974++bhdFB9VJ3Xe4AI0OdyMLMir
iGM8WSTFM6TzTEezKPkPO75ZYIZIMQJBHbiKAdBIxhhlpGHYv4oM61t792LmRR4H
UugDybMTHWPDSoUzNzmO7qaJtiXp8oY7GHyflgvJjJYxYquQug06sXtBOCFITla8
Ls3wzPx92xRulMA0onuydWJchrTKl838/oOp2SuYqXJPL6ivoEFEaQwt2Cnb82EM
beM63aXSW4Eb4o/261z2Sw50udfBcpNfNEt4cHXU6vT1DV/6O/6KyBvMV1oPjWf5
o+or1oV3+lZ4vUEvZoKhYWaHvwjIK6qiyNyIz3QXiGl7FLpJmubYNnfb5zc2aTYt
AC5exIbDjJqF6s5oIuwmBXIIjA4wUS2aK9mJYtVXxdrMlJBDz3mY7C2aBi8cihM1
DBHeY+pf1f3/4uIMGQkQgigqMknwd82IRCCIcsZz38zByBn1UhvmFFS5fAR+oKz1
t4ZOFE2Opx/81KRdXeRV13KMGdrb0TgCXlEm/z0t0tchWUL16ViGF6IzMWoz4Uvf
feFb5rJDX8ZNIU8tiCB1LJ9MuRqSJv487nd9RcX5y6wL/a0pQf5p/dTpFvWjIhAe
UcGIROFc1LNH6QFxzNsh0XVZI9OjY24qInRoX1woCvdW8H7orNUKYasYO4VwNGH5
LUbcd5HUU5y7rVYI1IskwEc+y2MYEnv7h4P6pGfqrRx0euWW/IrDzviG9moneIhd
PV0MjNxrMX/XaAqZmkrsIub/8+Miy7C7N46nj6n2ve8xec5kdAzIwoct1yJMTVGv
kXCtA7e3Qq9DTWNX4KRMVYgfq/YdMbHtFSc07vVLq9NcHE3tEPGgnKltrh+UemwK
+I3IZOFAU0sKz12JMtwPsBfQ9kfkiVkK85eGigxyCsWnsXOuOOcA/oURPM4l1ds9
/wOKHI8eklmSKauGkrU5uUKoC2YYESr6S7JpKwEgslv5pbX7uqy9WE7Bup+HAwLg
c+b2uIGWLjExukkHcbwY5sP3sAOsFJINHfNP0wTuKegCVA0zuNF7UDvXmQNWoIb6
iw29C4rnoZ1SeFsuUsiNa1+fJg0GOLLyXmSOzfEiBW1oaLsXprEKUCitZpL/ox0g
SBMJEIhQcgVyvsN66lKpt4fXbHdUsX13+wh7uo33/HZikc/nmY1bbQLkfW8diLol
RfwbnfWNKftroSVSCyzKxNvMztTtTzjwj/lcn/V6cgl+du03g3o1gc9ScCSrYKj6
pfzZ/xchjbhiNoLOUuQyEpZJdStURcEQZDYgS0B92yk5jLjhi14KHXIE5820jjz/
0ntEYzUWR4Km1T/UIPCIZKhKO/fUXl1wRLGaW0t/XB6JlU/+5Lq36Nij4kCNe2RP
zVqie1crnHJPoHb5HWrShD2gxk8h8ZEtGfQCxsoa39mNygroGw8OeWcDH3iFie8y
KoJXqLcYULQVrlTYwwSzb49+563xmkwlooG5Hk9wgSuT2QvOQw2IJX1BaPhRR0B/
D37nB5tM2qRJ3uyFEegH1ECWZNmL/ogZZs7QWzc9E63yw8LV6nwJtoPe/N/xFZty
4KLgUu42NP4NTfgkQNMNGFGUeDXafnVCFYcFqmAbtoBX0sP8oK5l00gEVemdvNuV
7xPQmR2jHKTzJQGtA5NrL83RVc2Afl0cpqdEJEWx8+fsNjSq4dY6smRt34W5GOlW
yNvzc8odRGLN/MkvEJThTRx3fNwZbnW10lz6ypXw5tXsxvd9+Hwjj9/jczwa+5lI
JX84tsEPsRRTZcnB1mJgyjRz2SrK1rmNfN5h9uzpfzaclEadtBvlABK9kxoJx2fm
UT9D6U5FNdBWMIAktnGH/vu45VIlgDxQ5s9hHL5Ff7kiUDzMXurrNaLDv9huemsN
+8FpY/WdIhZ7QDPROn026JaVeynI3/nW/s4nL7TxlbbzDjkvy6J81xqASdC2q+wn
Y1Q9YCuGNPM+NJOeNYLE2F9GSgLSkZQBBoafZfZ6rqBiLxi4NUdzK42Kus2KITgp
6yY4raUQcAJLoYx1zWHAH6ecSxRyoJs3S0PR8jRrlJpQcnHZrniE/pjYL7KKHN+C
bgCCKHol/ueuw4z/gH9QyLfTk0pAbbZKibWPslD8ay0z/dtjxclNDhkWwDlNGx/6
WpeFC7gNVXIVK/hga0ST0rak4BY5XSBotXHGHwuohIpg1zAmcREjO5HUjL5pu69w
8llLqKuHybpeYJMcBHaTXRCl3TQVrqwQDaKza/Y023UJNdwnmjQEcpMqIkxTs1Vj
d2ZR/+iPHTdQuZcJwLAc/wZfjNf3UwKJqxlgCNUe2PuSC/Yd3ZmNf3+AQMizp93n
LiXLLlDZv0M89rOSx+waBHFp5SemSTADm+8frBWVLGO0X9QypTg127t6CcRZPrWg
WB2L6M1NVqTT86gAaaCgnnmsgCUKHlmLcHmnTJ5hDekPYSNz7SkFC+yRGGJsCSAu
OKTytL2R9jAQr3XBng7lBiqn8kePQDpEZRULlzEivy/7qC1HvdEtvHCftTnL57hc
kLM23AGsbdEWeQOUfK/ARTfJGZn+FRETsubNoG96Ug2S7vpASQpNe8FBV65OHCS/
Fz+di3vrqOGeDW1Emc8ofv/moO2KkMc5EdMf8dSKg15BObl9ie5HWefvpn84Lt8S
kxl6WOuMCK0riHo8YTZ7lDQDGkUW32VUQ9bahDxiwqaG2qCYNMaCRoYat9+n2cQ4
WFQrIldvNpxRH84ch8ehbBburJTifjpmV8m1M9PrCbmU+LRtJOaFX/vd2qsDbbbU
X+59cJXA0eCJcvJSHufoqhLWu+/f3PUhoTd3/V2FmEgyTnqywC50TZO57udZUVPf
YPmFAddKYqvPx0C5ZRT/jdWVxF41ei+SgS0g7PKGDFGxi1E/7EmbBFpjGBw6pUYF
C1eaXYIfwkVHyl1Y7tm3MzdbqcyKiEWXjpYOhJn60ZA7//MPgB0XismaiDrUQF8B
VpUWGAFPNcgxTn21fUovKI/igzgTMJJ5DopBzj0jUxbL9DosgR+JH7Ua7dW2/jeV
tZ4L6Z26dSTk3UIPIdTVBK69dxfqkVOXsok1v8y/9vF4+Am2YmMReNcc4X4bR0Mf
GtY1Q+ka7CkK3sUrEdNr5e3Ui82zCWH8OfriuAIe8pNuLalCqtK1X8KNrfQeDkvg
GedbwvEhOzAHrmBX8ngiPu4p64mCOcI8GhTJPPlf7W1Mrasf7y/nfXPdsKN6egcm
RHPCk+4Or8dl3XWsaeGgUH6fw94oSSfsZWGXoeAkz813qoZ9Qw9Y9TgHRjwBWOL2
2qHw22V5Izad3qMOiW53y1oebwH9XY3phEZQ5ZfY3/Ua0uFY4/6bRR2+Q1wToqZB
WRiOBIeGInnh5mSkEiXS0NWKR6hfiuDw5Ff/A+RE1McUCu9LB//8/ZigRGNM5CEk
4x/80T4lAcRKJa7M2/5lEFnMFvF1URiVBZXw0emLdslaGh2fUvq7rDJm4NnXd7Wb
R+GmjQtGsSEpqgXCE3SPs7rKiNQ9qwNxhfJxhR3N2Z5FjeMkjjTIKIXf0YMa16Qj
oXWgKrEfgmNTR4GFYhttLa9FcOEasJxe6kywMWy4IeCaE03NXhr1eb3WrZLn0+1J
WKFnCoOKXgeO/iVMK5WqaiyT9Z8YrVkYxavo4lDTNGQcNrto4iFSQeasBkM3HNtt
eZpLk08+Q28GljmRojgOw5MDBO9Qbd7bwCR22YNeoZG+fD6sRfxD6RYGP8GYSgTm
cOxRMKUfTb4MoOUdErxa8RTKuPyxVq9pfzg35WjPAuGxpum/PCHMIyII37keDfjs
FtAua/bBGXhg8XVLStpEfUfa8/HfgkL9Zksg+2+WXwBWOGZN3QK+YNCK2/HokBKG
AvgG+JzWIz5OuZRfJWRCIuc8g0RNqXkcyCFArkjZif6p8AIhaAbEu9KsWafyL/Yu
7QtL2pHjc/KjOV9Wk8tVpjONh9uPP7wu8SYMbVytvCwjzeFBckaWDvkQVPrjLw6O
MkWL8mGqebyB9XAtkLKVEgH1JfroO8NVYVtYm4sIvzq5JQ7tEu2vqI6e8QkiQNA8
iqYln11ywV72E5fTn2mLOGNK91XvhA9MTq0E7wvA88+tOsU38AX5qYUMFwA+sbVK
m2W30QRHnim6q/FbuPx2EGF+iDmO+Y6tnEW8/3q7JKP0EaXFtYMo3rTy9dsruQRF
zQvyC4lNYDwwdsY6uBriIQFNivnF7y5hKpBFuc5q4RLTnfWTzK0+J/oN771M7X5y
K8zKyM7/UMNghrFgHpTDwkVgQpLu6/KJQCdK1bHtsDUFdbEio25G+TGL8UvTdZeK
R1CaR432E7jddjQYiW/fp7Zrq6dBb7wkYkJqUowDCqxzQ+sg/RfxxueQoZOMWKUA
zt9V5iuGuowZOWo6vgLK1HgO9tElYI22x9xq2FkD9qXsFXdOXucCQq95eZuj29ek
VvUrIYObwe1J5ZcGb8uIRjgGleOOxjTg75wpZSR7ZK7uRBg/I3h3meU6AdXGa0Yj
6fTnLjAtS5gD4h5UF7Ysu2/4yjJs9QBcJy4jmV8xjQFfDLvFVhi7oQD9IOOwv2tr
4N1Yh4U1hRP5rD7p/mM3BQTdc2s1BvdZR1sI9B/s9vqze9GvCQuSDk65gKS5jurL
z5DwG8jxidw2Ms6RbALJqQREd7Ddm6ZWMUmSzKdbJRce0nFBbpxiMW6mJUIQyK4V
CwgeaqlF1DmocRKxn6swvcURqYBgrIa2NTPf5PTFSTSHA/VAhrpfevHmLIYDIEDs
9dkUMFBQOVMotixfn34Nw+iFmvOizHAVyIlsD9WUcUOWZD7h9xBL9q/4OSMoel60
bgiJKGwYsIUxUnRCif25X6yc/wwzacH598w34+GJJMssELELPFQWZ7BIv5JPIV29
ZPonVVMqbN/VplF+x33etBPBdaOopvKNZbopw6qWW6rW8w7c2E3d7EByNifFniEO
5BzgyZoiPf8XTVkIl3+4VyOioBx3zbPTf7YzXf8yG7NjrIraInSK9WxdjISHRuN6
yDS8PxiBPdTWMTa5c5kBN1xxsWixYv9SArvMtUBxSscEW1JX6YQ3TtVDJN3Zn+RB
U3iSABRHY85QyYmdYKre4sKO7ZB23YKymWjraU+/vBnbhB5lrUa4UPIfvVVPMAf2
H28+NDrHYvmlOaWKxc5v8QUcO3Q64IW5AJwc8+zJt4rgryVOWLyAMJQ4qHJvd8Ru
KBhbFP168IhIhbGE4rSHSfR1HN8HxFO5KpmeNxu2Gj988/P3OvwpJolQx6+N7+bH
9PO/g/UYCSiNjQrVcMUVkAgAAfzez3DDALRm6kfoHswGPWq8JrS89sL/EUU7o6mo
RJDQ6UcV1TfCTsAOsse3kBf6OTjVKq3bFO+2Uoyc7liEFDk+1XDfHCqYb+ahFA6i
0Nv+e1gC3ckiuJbcZkYy6bdHv4YKEFRKZW9DCS/1kxk8UFfMSZGuQdtEP2CcF2sQ
RiCHLMoJ7EpVeSnpVRfSX/raEzMncsFbM77vXA/Fo4EZbNRG4uT2gc3nLaEwHB0y
xJgHkHSxwxQ8dWijZ1Y97uSBbKtIw0Lm74d3AoGSi26SH5QO92+ZNpIf+NVekCFu
YAGdpUYHzXbP/F/2k/Z4D/T/cG2kDhLWwfmlAAOgz1fdi7awNhWyryo74lEAVonT
Il5fxFRFc4tHgw9NLBLlkF8Z22BDzG8N22kuVvs0tV9oTPJbdBwlaFnu0/i2GZqI
VGnjpfKaZGyWA0bet30jBW0n8mceN2AlzjrC0/ppseIFm/yGqPEoUWc7l80yhwsk
0TfhFpOWKbilYjpQjvGfvpmguti5UE7pU8kFX6gwxKbM9Jl9OKGTi6m/dLc81B0X
+c9hFA2001PrRjlozyD0dsVrojmlYml/f9tGpHhVhwRyq93CumJACvKSb7TtWzjb
4NvPbxK3Z/w26WVjw7IfsuWr+oRj1KDU2E5n4lkZnHtY+ZynwOMvBD7V6RdyHV6a
sL6semGu+ogXbBq2FY8xfm1EufE3D2CUGs/RpOC33QIylbeO7NcRV4/aoza/SWde
661WH8GssYPawxhA57dqYfhcKWgntRiQjYtcD7lrdR3O1WRt45iaZSZ2wT73dhmv
B5bfCGnZT7nOECfA/EhPzLNLHt3Q0V3A9bSntBMQEZz/D2sex00YgecTCVxG05hG
0jMj083Qc6vg2LHFhQesUmzmuZWyjLa4V/jbyRzM2GrRJJiosg+3ymnIwGVdvDO1
Ybc9pTT00qQBPGD0Cma1AQY54CX07/w5eYtnTXWYonkk/nFNh/yn9SmrPwjXDoRr
Tic/nau2IN292U7eb3p+Ttb7rtVTGaFUMnnfW3euH5qaojsxrrvEthmRdIiJ6mrG
DqexbrDsJCzkPnwtiBMIAUOnw5DFIiSGQmFhzQsSn52X7JTUiav92UvRgDoLHTI6
qE9h0j1I4DShYnzU3N4fgQxNWVyU9+3tSo+tXDn5cUqEUdZ3JOgzlM1zDGT8wK+v
qMQVQPZsuDZxIf+LF5Y1kA0Rx0CEUubnb3nETAslc6gXN11QMbIS5Pdm7h/mQxsK
IMgi8uCbHit35Q0SKcG6yN3CU8nkArdwn61AZJpTXkS4bRsG61Y0HcajmjIYSUp7
maYx68qUx4Z0eAMUerqIq6J2UUyhZydqb0jh1E0GDWVzZe15KpsT08VLtIhGmP9H
ZptzqFXdgZRHjkIWgEOM5CXYazUjA/Aq6lUrUcFIb6G5YckLn5u4elXHT7rLubE4
hqHY28Z04f37bzarEIMM4+kgQFRRkSKwZT8oYU/71x7LyqjvAPRW1VbvQNPgW+xI
0ZJX1MYAGl/VmBR62QsJqrTE2J2asgAEgD+QaM/oEAkzLrpKfS78EUPqtRt/TIXQ
tSk3iJ47oOCKVs7R4k0eGL2/dvUD2DleYXODkoz0HtnYrFSE7L/kuvug+o6b35VZ
zpzbaGNlDkYPNKqsMMcEGPKAxC2to8Oe71/8JNB7YL83AZJYz6IgZAH4iVbMNaIs
Kz0A9o3n9lculM3b+HvPzHZNgFqdk/ZVUGZrhdGeZlpp9CyRc/+YmnCp96hTNHao
BgW5K8PTGAEtf5gxUmozf+wXTXaoSyJuJI4fxOhiVGV7w1GuWRjNMfKQf5R2T1P+
Wc5vPzdlaZ+7LNXTCRaFmB4S1HN4zX1wKsyjDKAvZqNAaOLLvS/Bw36ByA6vxvb0
YLrwrMgvJOGmMlIUeviHNLyRM7rDTMTpPPTGtaHaJnLBzWnNp4FpQmacPIM6iOy1
2Dm3vf0umTGX6Jf/NdY4lIpQ37wFWYaGAX2o0PUhmx+DHd2umU+p0BxHeGbSm/L1
xjrK0MgIJ12BlkGrrye81OxXDvKHjFjRl1ejo0kUB8+C0XyJy+D/nWNEXOZZ3/xV
LZOf2BRM+ArMwd/AdVw7AK1ROr1yYEWd3f0SfELf2/0TarG/R3GlXJEul6MEL5dT
a1i45p3SGRWM7B2I4/QMWWk2zpPzFo6VZhE/14xD6vO8nXuwol7WjHinhvpxYt0m
b/WA1dnkNlajTSsWqMS7T9qFFQNqONqMgzDcIwBrEe/ygj/2G7NyGFGRNwA5bn7v
Vk/N78bSFHbs0xy2P5dce32RkpPu/ft7qWQp8jja89AWYNuojcMYpZacZKn9ASgh
GgLcRUy1Uy5qQCbx3e0QJD87KXYhLqYi1zP/4jahXTpaqI5IuVb44IaBCYtViWsm
sBi6DdUxxzAhxNV/Wh9lXoPrwm7C1V1Ya2bikjm4EmxP0mFtTJc4H4W5gbDFy97q
QaseQ/nUEqyXzU6lstxi22i0oWYKjnPc55Y26COeAwPTsfssVHGgELmn4/0Noyku
B1MtPkqst/Yj22X+1n33Qe1Npoi0skiK4I4gZjiD+9voQaiiL2m0Q1sS7nR0Cp/S
ZszXyMX4Q1amymd8r6aFafU5WUR8suy+SCMPChgVhLLiCttjpB/zFsLHQI+ivlBa
OOUeUTjxQ/aAnGpUFSONGcgdMr3Od7Pry03znujE1Txu2A+EWVYe5u2xlJAFu+GF
COG5YvwPdQ/+1Wx98PhMzxpYK8q6B5owoy5VBIYS4CQVyQZ/Sv1sU7qgVljsJVl3
W7bVDui9F7F3tY13x0o/mjf8njZQ9yVINfUMtWStRXBXXmvqgeUouyZ2VNZcv4AK
vxwzLTig/NaGXAxt77JIYUxc6lCFNJjOd74naR4RMuOjgGlVnxzEsQWr8gb5zprX
owfyb+Q/L/ej4kqPr0sbBcu2TF+4OdNkIA18WnYhJIs+gakvXOQdlOwcwW2LXRSC
bKi7bBWH6qXJWdUrMZCq3vGVM7B/v18ZxSNtCNWZHW3/ZFKmq4AXye6tmCOxC11b
+GcOjaMc9LDUypQ22qSFDu9lBoziGVl1CsJwdvBB5izrjFrZ/nOA/fYRzD7+v8Tv
eXmZFrPUrgtGlVHEYZnsV8wzZBn1+O39OcSHAwvOyyAQPxonLdjQDhS+nu2nIJz1
wjMatc4miONEUR4V1ye/oxah824H0OhG/NzTNhiGuxzBT2zyyVANIYZgWVGuvbjX
3e4F8qf7kz3ZLlL2Elxlzuh8rOm+eQFSPmFjjcyBvtFAUhjU2ykBVRptZ9AjGUlG
P5I67uisuYtLcVFATLPEYNYXnxSfRrFNQ2Q/FYHEyKbvU+k/0jZs+eKgeIwKlQ15
Yyj/QoquO7NrEVET496VEpiJAw7Cc24w4AdRSgdGw39CLm4QPXg7Dhd33dnaY4j8
xeOSboDQuGMzLJgBDnhfoJ1Ju/UBc6+NsuKgtSi0BIvp71+i1xDLjW3xCpQBzrws
tjubCA2NFHiGM62+kTcgGvgB1x4/gEx5OJogspz2SNPd7jh7YzTCtMA8dL2AoiEt
tHt1y9fdXBfmr8lCYPHhMKMt1/ji9ETWR1zkcejcuGaZ3zLK9HetJfRqJojsX4v7
KrbWgNZdsTU6hr3JhTPRpA/exCJpGWCRqxVItW5oItMEblTHg8tbrZFvpnQE5AyE
4qIN1MJoUAKNq3F7M0UJ6tnQZATnRKTSDKZhOQ2Pn5TwcOIzFbX+CGGFN3gtfwd9
zG5HsXAdpEq+zYy+16vnuqrdlmgq0t1wP4RrvOHr/eJlAONFCwCrXtsyVLMljcf4
/cgZMNdEYYbEogDruoHmsmejNanohLdtg9Z7/0YsL3j3BnsjHvi4DF4suZ1kpSxQ
seBcpFNGPopEZBzt8myX6gUkAiWERyGyVgDEMNpXyOkBVJUfVruqFhLOLKyPa2Us
fWum2tO7AA/a9TUjXf6pNkiYzvH3DJtD/QwNFG5lqgH7hTSQfH5kVq2DN6MMV2ov
+Ry92Tcn0Dfwi+6bsh0kiT+UU1/9o5FVLqaprPUlRFSZIaF3kRkaBC8tHN9OP1+m
sn72XvZLoWBoG8bZis7W4C433LeMmb7F1CjN/G8h53UYDQHGV698Pi39O/6roGXP
QYsh9NVP3JS3C4MaLrm3sARcb3rWWSy3THfnsNr25SlFCMFt34wI9Zl0go8w+9AL
xudM9pmlqBu9ZGwxAtIE6YTg8MIJKeKFk5ASsp7jPtMU/cMS0z+CWPbC9FqKFFkb
L3NpIHIJzPqTLJeAdEEcUPJegtMgFkUTPOn/aaeN6IEXn9kpjk/tikpO13YPQ07F
aEd5HT4VMZMpUhKG1ENXc+x0UcCui/ngPs2K2HNgJl5q2RtdWZzyE0WV6/uUTzUV
ZTn4Y4mse82Cm+KYFequxT/35UkI6uQWnX3kQg3waDj0bed3dzNnvIXwXA3uz5sx
ND0GRqc5DpovQVm8TIpnHZF0h2mn8kJJRQYm5FuZrO+w8gA/4NmHaBIM6Cnf/nWh
aLacj5zZ96bdh2jCUEaLt6JUyvw2gWnOXSLmRLe3sPwqiPzd/0ODt/qrf7I/dkje
HW1ZLnd/q7lueNJu6OSRjOPB6VEbTe2sT2Z/z36l8ko7zpu4rB21o3dJOBfn20Nb
VVLPTWMvMSzYpdDZpp24Obtvq3PrOb5C5HAkeCr1vBMFeAtr26gLYyXAms2Vo77S
kRN/t+U31OPSYvXjiUIEqsctCrhItr2OTQDhzyaP5Xt1klJRMk/eHG5oD0FQa2QN
qijLCiH53kdy97fjSDhv1emFw3AHgcK71Cw6KzjqAYILUd16pDthrksO1Uc1d/ij
si8MAVCEZ7rErz1DFYRAiFcaV/A/ml6Yy5PX/qiF6F62XMG+knXtJ2O8sb4UnfzD
HhusI1EQA43vj5ymu2sDNiMPVMBBkbxWg55QFjE+p3HC/UZ4xP39SRJBra3yogKR
kQWzWyp7zP28l9VBGL1pMeLeThX0Kn2Tz8OL8qVjR4SUsBYkUUm92U6UYMJn3VuU
iez+pcrQzP3DCqnJABMWh+X9NWOVdw6DsswAes1WT1+3nG5H6lD1RLBZtqoNy70s
2i+AxamJHWRswvDPfso2OsMdkqfcOcEjljk+SmViE6iCahkSlWw4pw5KVxxEhWUt
w8C7lvUIUlUWrtwbBnyDQNX8e5+Gb23eDj8xL685oIQtOksr6TVxsD1DOrm+LOKP
JPWZNA3/qeha4uUsxiCWejPiTHj8I4QmEWvcKpqw4IRl2Rm5D29RfFXdbB8vEkPD
HWRKkJSAFiVmdcyK61fCdD4QI/bzmLQsdPNCSOZSnLQiTlaMrJ5hzqUSLFf5iarx
UK3gomD/htOsv1TQ9kM4/RUvvDoLoYL09WCIAXRClZ6VvbNVF1IJr+jW2otlJ3M2
nStr+uzAXX68KI2MV9di+46A6v6x8YZXETMZ7TLcU6xncjv+5GRm8G4wxO/poFc+
qEtGTlFHoU4SP5RiYw5XPUP0kLSyhGayegT1L+lKRbo187XjLWq7DbHsl1kPz3DM
96Bpt8yQoX6bHfd8saqYfrob0PP/PgnP59zyj/C0ZbjKmAUeOSanOWGlJE5jbooA
86iyoAqIjMM8jXxFatTqWYoiFqNO3Ail1kPr20oWtfkvitmmEmR/Xq9X2x0ubTMh
IOydfUsz8COJrLWgtSgj6kQYgffSm7sTRrX6cRodHct+OHZQ93MszVy4sDU0YYvZ
ExM65MX7K/zBcUr6AJFdkvUv1bCpMYjHfhNaL7WZ6vkFcUClOTXBoQM98xwj/4ir
i7OMo064iUMUx2NEwvmLmtt+2V2NZeqnzGZWwG4r5gLUUZ9y3VpQRQsotAgKWZ05
BAt6N+hGpvGFWeTAHh9Am2eT4r9RTjLF/R9E3DmksEQk2dgtuQ+0vYt1Dyp8+Ef4
a/+tQMO2gbBepNHimDAnulyRlC+CdiCTbzlRoJJrCjeHICe86+73furMXuIFsKM1
VV0PRBzwkrrRoZm1Yq/AEA8cAAesdSS2eBaP1Rh38o4gNisH6qUjXmCN61DlQDfh
4pgdpfRRhnahhPwf8ZULfJalkyW1Pq7uC9jP4ar3AtME/nZio1ci81L7rcerDacO
yJuxzEz1xR0F2FNvH15CAJf41IKDxa/G/YI9kjFmGFOdbTppGKc/Zb1Gs2NdFsiG
qLPdZrFNVT7Gbdts3WCEloLj1g15OveQZjLW1ETbBp0CB9zvNOskPa7GhjQDkhzc
zqyqoXjlbSKdxVv62TYxslOhq8cW0COhIoNRJ+7/aSD991EaTyAx87bQ5wsjOHzz
CvkvoPPzCm3ZMzonMPuaC7+s1RZabadfO56LzV2okenz100yZcUlNnmvUMCnzNnK
nwQ1QEsBHEfkCk5uzLbK7aFNn8iEp2d3QQ5/AxKNDytDCmL/2yHDizKm+3UxXl7x
yFe7ykjSL+ZMSZQdm5J5GNkkX3mTeQ9v7m5JX3oP26n2eta/zutPVn0wO+xw8Jzx
yuhp7zjSt4CxnhFJQXr9wrQ4ajeZOzVIyiHIdFSvXWj67Fi69fs7Mak8Hh2bNhOV
GclOEV/jLYy/EPvTc/hVwvj0OUFKMJQx/TCIeZUTzE1MwBu3BRMpMbv+YoWKLNMU
3nWLZqN6YSjBq4SQyykcZIL2TZ95wCW+5T7JXdcxMJDhvtxoLLxr1dzNDXiD3Aoi
OsWXbsj2BEXXCZipH2vdI9pEB7zuUxKmaAJWLCYEqYiHnq5yk1nGxz+e7ggPtJPZ
57pJNGCy1sK4RNZ2Ag2qos873UQszoTK+6IuMEqzTaEBfleYpjYXBbUGvmqtpjMn
NHu8C3iT4bDFyEdjTm8fLqQKkEb9gG6sIJUKp5/6XStXHm/0GX1LCK4cxV0JecVa
SfGYLkPo9G0mukcGdp7VdU6STFkH75GEzrntK2T4s2EVwHhksuCbbyhGKtFNwvtg
wXICC+NsQaxN7BBvJ8BJ44BsfLD0EJOxa6501RsO4byKOIUCL58TGUlW1CbRaP4x
iV8NeH0N6KY/vnneNyDtTNq7BDFSekceWBDe8BbchEtpoJWZctri+Ic5TdoFJYD3
HAHp8xFBWKACBRKyPv5l1Z1IrfjIMnbwgQuQKQnoWgZturkGIpVwRpeDFOMZk/29
KkXZ+fZejK4nDqq9k847ZPlKy3abB1T6JbPLyjLXFgg+ANYp5B9IKiwPaLagsgO5
GbM+AFitklm6vGtiGmA4gPsNt/fVfhKgfrQYsfK5stigwlY3bb259bpuDyjLEMyq
aayKEHeU5915mSYa18S6jP6H27xxJUkjtGLj1+wDm+Y9u5Pgo+VTDP8WVo3AYKiR
PTFlA7GDZjEbBtv74UIu7RvLSMKt5XVLEJl5tOWFBwPeg18/aR43Qn9e57wgm2i6
/kqyzwTbh2u7KowTo60JO+O0eLHJH6zXcuULyzUXWqk7lBm2OfNttv5pZnp8re4/
naffOtZ0fz9TjzdwnklZ4TTaCECcm+4b4y6ZJl0mAvhsJftLsezZ7IR71pKFjDdS
NAUuB3q9j6HZkQvm15kutXgJD/OFrxtkwjjsuQnEMfS1oHs2HjNNDnscIRwrEYhJ
rr+LOS6byP1cXQHXYVUyt47vncx+Ak8+e6w83D+6phaypWnEuUlmISl1ihEkUMvF
l39fwypg9WrfXMXIYkbRoEbnERjlLA88dxnKIxNCESQqUtn/HHMvNHmorlwSXCg/
Sahl4BhAtyWH8MtR/fEQb2WNd41eVPI6F3WzX/mrB4/bnM3NK9pFe09H3vXQifJd
qIfWyoTo81miZRuLeK11BZGN70Weq+FLVaz58MeLD8toPUGWbrztPELh4/qGU3pB
cvrDWKfAqV9ZCSVX4fIyeEKmUuqvA+ure17nQMm/xdTMm9lcb6dLZ0aYZj1TKoWU
2DmYTA1TkBhaivuMBv+2SaFssJc7KEixCBrncIV+QBbPO0VmQh7C/MQR5y/OAvHw
GYZ3H1QuX/8E79LU9BlTKHPV2jjaVoGK4TMwsP43P/bHzBmkVLQ1QV+D5XD5WsL5
ZYhfV5BXWbKM7kaNwbhcV6Rowi47WfhADU7/GDGzG8wFsj+zOGoqKOvMT1nPfsQQ
efYu9qg4YHgSlSXVlX7Y88HmgbHBbYFj98FrexGmLgkLq+jXOtjsxBd6tpy8teKe
jEgbn2NXuGz84Axb9KQBnzU/+xP1TSWCIiRQ62GFHhpY2/LbLwlRXHUu1ypon/zW
5OjSY34gZ3GsiG5rqiLjEoozHuctY92gcfeqdWKd7tyfkRzlhyTGz1tVZtG4RViE
/uLXFsWv20zH1hmBNPjgiXYttvGLhkGqX9lgbBtik5IlrD3yDbRqj5yC2y16bqnG
XL0CLnvRtKiW6fCYN/PnEYz+wHFH9fxWVVpcg+KU29B42E8aRXWdcgBYWgZO8clE
wali3g5ai34sShyy/mGSOo9NFin814pqZj3ZH457tR+hzd5L1swhyDYO/NYe24rG
aWGc9nxcLP3U393ZaBy/RYurD5GnHjFKFLOAVIOdNeRrAHU6EjV1uqmBpae4irLg
KLU2kfNwXO16ATbefL26qCb5po6sys+WP+l7sBT/TO12uWwkHlSx4fW5YRjdpjzC
paJlcKcB4UxGaMLynfuED3BFHPtTc36MUl/i915mW8SmqXWP5usEjIsWk15TQ+o9
0mDElgD7h1rxlT5X07imrQ4j1FeSolFUfetBA8Lbev8zc2ekoQ2IMTwZ4FzmKvlr
ABgbNF9eNu7M16nLfjkg8dzOYNZ+D2k0KkfUcLLzHXSgDw3SY8OSpqm0ohrJpljj
2M4CUp0tEOCKYHvB/bE89XmksSnYoN+aA0JLPh0gSZ1ZRPr72AwsRERf6ZO5lasb
JJont9ZeD53wgftR55i3LHOo/PrzxLn0c2j6DTWQxS6k7Nc43FpKTLhn3LzShf1q
lclbWUCoK8Piopesovvf+gOljNWq+My5p7Xirj1ZIGjNtrSCkQUgJTt8XTq3MHFz
yfsv00WsDGRbZFc6bzN2fb0c4dxH69aYBFdPmxwstHPJeDHo0WIOrsVnabNJlyvs
I5QsO4A6H+vErE4EomgmfO/rqX5Z4IKkLk9WmqJa8DmVQoMFdwkJXEU3nH4C+fji
y/SurkEffc3hG+Pbj4DBT32Qag0gYz1qJXfaat1k93eFEfGqDoSeywhY5Xnc/0uz
LeBNASd+cJb4Kn7anfPOxaBISG8PlmVGrOllTt4Sp52rY7lDfI8am7gaP7LdBn8r
1I5qBqd34GPjXolzmU6V9E+N2zdX4PfvhIFaCWW++ZtLMK0UU0P1yAt3IRfHqTXv
7oaKIJ06ClVM+nbfnULeK9ADdJef5HfCgIb3Gb/ZUAYkrttZXDk2tbDk1tLCnBdR
kHAglGDVN5KTXhM4wf9kIG0MDitaWLmLls7Bbp2ZR1sTtza1Y9vrfNQPWhDT1Odl
UKLtIB5L0xt67OfHkcTfyhMyLqQMkHLCXf+9CXlzSpw3gTgPAlNQVnn43FqRFkP0
9u5KimaeAYhJ8Ip1LnRh/lNfod6zM8KV9CW7R0IGk5E=
`protect END_PROTECTED
