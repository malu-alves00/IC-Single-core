`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
E1wl8DX0IBe/3mySzJBsZdyeHS1quq6oRYfpTZisCgi/wPQSHxiivyxBAyZLgNDS
lkPQ5Nw1Q8c2hnj39qfoxufC9cLqOuKyOxLd3SkeD4yU8YtOnpP5gaQo2jb/Yfti
9ijiZY89zuO4VsGWjVReAcuhbV/mfam6Bi8tzboNuBc2pX0T/5Fbkx+UnpDsAMMQ
CqDfO76/q6Pi1ly2xED9A1kQLK8lrsH/OeTUIl58Q0WyZoeSgK7/zjb5D++elGS2
os5WpUsruTQZifhCbyxHzejacL5Ot1ZIAPJjARpRbz5E93vhATiUbG5Kdn3Dh3Bg
X6GXEDZJ4bCZFyOjQZ5dHJT+NHHord80kdQ15HQJqqloBolf9yo+4eNaQhfDCj7V
PltXJ2IEpu4l77FJhekPv4m28S2AcD/71Ai5lyCtpYt6Jhev8w8h+40qYZKIwPuh
O8V5Aw14IvPOMpJFHvnnXbipiJZGne2HUfdZ2l5NygA7YhKp4n5/6uD4rSLvtfwV
S6X9JQH10EoO4Irat2haQJMUJokRhPd3pFe/x6aWNPR7mdKXTuXJDaNgYNcSFUCV
fceeW/M5ay/4j675cG5HAXAwxXwbBk90javr3oRgSTcEWLRMMHy8LWpLvUJamokv
WIeiRKbGThcCTZ2HlRbnwymptKDhnB2ldYlIT+Q2oYjfBMAKGom7I6amHMsgSF71
BgWAX11wzHKpv/DxERjjGM2lEVOsfQFQBz8rL4nBlKsQBGbAQ4KCgCFNsJcLDtVH
V1npxYkcI+3nE5ZbSahJi3exDNieKf0fsO2enwxTLZE=
`protect END_PROTECTED
