`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UD5YSL6qfy/eIy6XP+DtQEoJaJayy3kh6bhAhd4bUbvNhiKjW2Dr6YdhWnI8E5zu
6BQqEkaZm+1kSzUiHAXXCfppHfC9BGJGqjmgUhAey67ILrLgOaj1Jyh58rVT5hqL
NJNeJX8KOwXDP1xuAhnPIJNhHeFGUYs7JluyVuZFLiJSfM8vnsUGMCzVedV7O91y
zDzmINMg2Um6WGD+31sUfqxDqNJhNUTGGV+Ap9XO5S/AGQ2LOi1MVfUt4/jHamDn
fFdA5xFLFnTB3j5jdTpmdhrc2wJFSiTDbGHlf8Qu6tbfrgTUZ8KWroDYZfnql7a8
xQiMOPlxrhPGyoFR89CeA3JKQSQWFQ/V8Ujng732J53jqnB8rqdpycjgV71bKp10
VpOtgZesZI4KoT9rdgwtSiTu9+3eYaWigQ7OIG+06d8oe9LAui+mb/fdXhgKlVK6
IWvyBSSifumbEUxW3LygV/GoexTmXfdgD3dP5xyTCW4aPYnV3b5f5q4BNALcnFfo
uXjLBSr8a7D369PHwvHAAPuQh4hejT4ToRHiaKtCCloNP5Rh6bSQwBt4ViOSNBie
yOd+kg2LP/QCTFq2HfMTBluHhZUAX98I7LOLzCc2ZCRxtALkUKUTfSrrzAUPxW1M
cSYJa9fq3kF9S8gMDKcNYKxWh5le8V1ZNEX9w9JXMAvAuuhTIgsjjO0DTQEYEwsG
ZwmH3G6DPYB+JU1YK1ngNYk6nirdUY9l9Yn1rdVKPnLhacijxu0CoyOMkXCPEICU
mUzR2lTVgSm6u7Pt25SrlqpQkgxL7K4fem5JXAWFAqLlgcVuX5kfj9KGZ+mMFAgg
opFL57/3l8YlpkrGK2OSuHh76LomYL6w3YvBQ2PkHEo580A2n1omT8EWb2xvuoBs
F9FooNJ0WvnWWPSbE99MwQZ5hIhmivYQ6amWrGKKmkE=
`protect END_PROTECTED
