`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
agWgmiDOHPpeGf0YCjhA4vSCZ8Fi5wkXf90cKzyW5imn60giVZeSQkl5xAwQddTS
mR9FDva+fLmSUsneXsBcCUb7UlDXeJ3Gjop9lii2PGEsnJB/zP6dvmedYaF5Y2r6
U6+1D4uvbRYmsShRCl3mTF9iE+f+wtmMLi8A0sFJYESfqF7XuXD/kAvBJMxqjp6i
onBDyR1vRCrjszM/oJz6+LgS1Wd6cJiLWPR82lJQEHL2I2Zb8wN6mEGRME0xsJI8
6puInqL+o/w8lCIeg+9s2KBOaVHNhl2fquZJ9P1tWCsIWGmkDPr1lBVvqCipObSa
xpf57lkdzb4Xg/sM+reBTk0YrJVgcpOE7cZbzoXsNwksf+Y+yNc4/NsJ3VZVYKzi
c4dEAMSsFtbXKh8VAZwNu6kmI36Qd+P18uaXPPMueDxZVL2rjZDiwIIQzXinzMeA
gn5snH2iy3OiZPxTWp26Gzo6t7D6atCzf8XSx8kGZ8HdE0poXebr7f57RBWnFAI3
Kd/m385tVuI5DI1bGWJjMYFfuJ58ywvtrO0LxVUnyxUUml9n6lKtPrnURSXnL8pN
WJA2k1kBq3KC+gNd2EBpl47ySwpommGq7f784Y7/SHbUu5L40ktvxWpxOHFE+atq
yn3HZPVPxO8d1RqVSt84UeOUP/WLdaBDrHIs/zhWFak0MheLWEOyqdVQ1bWPRvj9
F5NThl2DW3zpltSwKgUtpPu3XbLiO33Z8dva1QCPgcA9V5vujRkxX4nG9gy76KZt
KnPGRGUyOveYV78qfn7UrN0orUqKrJWr1syKnd/teRtQE4TbyhrHy9fM1ob8LIOP
ZKrZL4lK3d5RcmvozYdPijRR9dPHd0gnpk7MBHQqCIe6x0uFtNQ9q4Iw9IU65g17
2cSMeJPzIj20thuqw2MkIYSz8yiiLiI94j/t6lM0cwYDv7Gpr0SmCCsDrBOINpEg
ebMbhw46rfoL7ZSvLGelwuAlYhmmTRNtQ8QqnLWe9QGEUHrBhyjxNSNi7z0SYGTG
byPm3al/fubyV4UNCUtKEnQyGCkgqEt7vYgUdnFN4fMyy8bOXIcqm6DAXAF4iPAw
/N6s89HiiYDe7sqelsgk200l2YVcyCji5vE7krp7fP6Y47X6hYoQjkrgMvGeYF3U
cwkfPHZ8tqe9e7/7ISLIGgFqRCGAELfPGVTdaYLGmgrl7xA/wQdlukyboipALETn
lPiHMWirHAbek6qacibSB1AwRmtCr1wcNP7BjGRjJsHXeaL9v/lHzSqgpr534Fk8
ThPoS5WHHI2rWO/bYdyqaJpoJKJXptMs9OaLj7tWw5GWG23mNPoRmGNTzzFn0Xj1
qnm05np9RSnsmL7ELHex768gUG2ERPett5TTYAiJ+K0I7YKeY52MO+YCXWat81+r
6j6gA0nzQjYEEWLXAhlx3Ur6xdI/KBdhVuNBFB9sBJeV++2pvGMtQ9LdZsZBRGPT
SzyCftNx076teJDuAUWvAFQ8j/qFkHIzdh/MNxl4SXGBb/7NRAVpNKmXVm+wpa2q
foJp+9tTf2aedZsEe9bnq3Kt9blqGoZE+EZzUh6N3zdJvGkUGKtEUKWVijWjNQpU
N2UcFGeqa/RCppqXmTnA6adDf08xk2goI3bFnEenW4N10OoyOKoTXEj3rdgDgQ+H
mvCo1vosZEKz8v5cHwySZHCX4/15+lW9qvmouYwq0C9veJz50NBlQbWBAzjgkmHh
BYgjNKfurOe7tR1cdcyjB+jh9/CQ4BWzfASkwaATLqw3abpAxpFwdxXtmYWw9l6j
216fzxEJBFro2LEatzkWHWt8WoCFEWyPdZv7nXdV2NWPIhgLk7XkvhcDBXBgLDT0
fp+N2MsAqOgdPlvo6qZBR8mjSacBcczO8/xqgtNaOA/zmE8uKUSpN/VnR/MJcLv7
lwvDMohLd5qnLTlxRNPsiZbC2DMMoYCb23dwNYbhidF3uYRJMGsAyxvt52g1XeLA
N0Fa51eIQ27DGg6n2iQBbFfjqCoY28ql4YYkXJK0Pt/cMT40RLUHmTsBnKYfK0/G
ia57kG55QUmiGSyv8Qxl6pj+FhB5wCsZj41LAXiH+sLBnx/SsL8ylii0VbzdeHJr
4yoCBz0rdW4wCxOJpQyi84RbAp8pwMnYt+HlfZJmCJw=
`protect END_PROTECTED
