`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sFEbuWPfNVugK0VkanNoLhB0Rdv3TDUWm5LQp//wxU+z1NmoNCK76u+y4J773jpN
Yrjj4DAXEoQSvOvSQ6VSGdkdddTIuCoJ8FbtaHrSVkwuhM9g2DE524YgKWTDfUNG
fO5DtcdmqhnhWnH/TKm4EB3OH+meOz29OzWvMDsgPRcWPCodQiEL3dYKeVmHnYip
t+ObCHm1zE4TvXqOmAKWkPu4jnXKZrSV2J0qu5P/KO4oVfBtelVY8A1ViITpf909
chPk/QVwOL6Nji59xR9AvmkReg8cbfEwzNhWxRxd3Brc8OX4WjAOm4oGcrRzsYrK
zUTBzK3zhqYoB6fr1u8i2FDfnnIf7e8TGZPrSxH94/RAQ11sHo2V8iHH8+hrJvBO
3jlqI2HBMBvsKunwmfEo5ZrQw5FY4ezGmIppfC1SPQzZu2Op7dVkvScKR3LT1ZM3
CCDOYCkoLdVPOoqrQ0z2W84ALrwVaqR6tsk94+b/G/3QltikaY09phAt8XdcU3cq
mfJIzYHXZ2cb01keokTF9IipXSfbprbvW3Z5YShqpE2XWYFucqeNvBfI3tOdFOSu
SSW1blhWOLBm0bvbWsfCgG/vCoLlvhBtVPzWtQPkZpsBZZnbncAY9sjpFdKM/gKi
jn+nYK+DIeaLIVoRm7m484U6WqSFtPvDNTcpA0zzZEVbHH4wXQSBGbI5uo7XkYLv
qJgPWZYIQ/9LNYIk2OukCtebR93kXTi+nyNOVKiEfALcQPdhYVSyMR4I/5mWuTPq
tGYfDJjQi9t7U6BEOOni6GXzD5Ogrss5cUK9qe+uEjafgZl59QM81RLp6KHQvtOe
ojNa5g7Cd9JmqhMOO4H5CC/s+Pv78FKPvzLHxEWQBLKy7o/0ZcDfjsq08PKJ+dD2
lALuqnnj3pzVZicKUw0fGWXOCzvbldfQTnxj+9KsDFkhi/He++oQfC3Cp6/F4z7w
uMX5W4/4hAVbru6dalsJG5/ESub5hMhk2fT1TmxNGY0+nR035G+66mA0Du44tua8
MxasyW27zJppbV89yVTAr9AUhm4h3NJKG3j+onFHYNyQ0n7lTXdOjOyYXTEPywAT
MveonFS2gHvICH6B0ODlcEXIvdFTF0kGutUq6Skufsj4tM/HQqG4nnk3w2K9eSVv
0SpcEAmllV5MDXkY82FTg8GN6EBiw5b+kpwuz8vY4GNQEGcMbWPDhzoQisVI0nR4
qESB8zxVxhH3iLoxrfHm4isdK6ZvouT7sfukByG2Cpc=
`protect END_PROTECTED
