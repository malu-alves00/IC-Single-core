`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BZl8vhdEb82aShZxXAw+eG1dy0+EZP9DbZ/vTRzjsls1b+YY/1z0Wt3lCiHYKmnb
KJVRW1+DxTiL/JzScC6Ys3UVn4dIHNte6Xy2BesRwc01TZx1YEoftGcsxz9l7dZY
DJKOMSbkiGWl6MbSZSBWfG4NB8ZK6CX5fGN7mlZHUzY+2g6sNqcehliqWhXtK3Jd
1Rp9Ii/B9sWdK/5X6Ym4NebO/P/8U2ZgAOy8M1/rEYIEw5tNwveNq4cxj5Ez7zMF
kPJ3xuiV+5gozgPX2a9pxNmU49/+py9aZYlqtyYztnvpLD0yDZojtBGXblodypNk
3SySsEoLfM+4iFPdCSEiKi+ZZj8+6nxce9j3iKj81BPXJRGmF88X0aSg7knFlEcK
Eh/aqgcjXbqqz86YH1M3/G2IF/1LH6Mi/M/SmrxQzooWYHmaB3VyPCnVmevqmWa1
8Up1pBwqktU1qjkNAytITEHyjQFDQMvw/ZkzIQGVAcYnLlZJJOe+n1HPzadEyNNX
9aU/UsYIy3eefFk32VAJWUzR6ApHkg4iC6XpYFxETsomu7Rbso2gSCKR255O/OEC
M8wWaWEVqnFPsBcQUbEadZMpT6ISrWpj2oaFqrTOMdbExmRml8jWvHDKmGRIrBbE
QefOC5d1rH4Iy6nNK2FQ+oigg+kroyCrfsmhNH2AiICd4mc2c3OedHkhNIC+bLxS
3v1P7shsQXT0Kw1LVm6HgXDSgGYYJD9EDie54T9hd2+Na/M/afP912Gj1ducvhLr
yI2lM+Z/YQWd3T475UKkvxoPZntFsw6/RM905xhfzJYoL2SngkKUcdmMqKpeNiz/
Myz3TJ+CdRvWGzjkcBWsfTBtYgxuzRsmmDUt5xq9NSjNFL9td22/F4p+fOl4hhfY
+YgU8n95LBuM8d96/LEwUiV+AjAzpYo/2yRwI8OPzOqWlWvbjS1bJLevNGhv80pa
igHy2HFjBIv8qNgc2ZHC+r2j9zgMDZacZ9QTusVWIbRfiVjnFRKkhP1mYDXxuRYc
a+My4Knc9R3fjgZan51jyqMsLdn4Z2x+PXnlAS5eBpfSiYrc5l0M1k7++hwZL3gN
fyViK0y/3TghJQQ4iwwhutWz+gQ4ZUEMLmQzXkdCEZIioaY7H5HQisIgRpawWWjR
JWVFz7JRyJLYKHWelfzG07N9AItF5E+Hmkn6UhgLP3Zy0KLmTgDp3c2+8WXDIO2B
1Qv3PLMofoG/MX3flw+WOTcGipnZ8iKoj4QqS3MNkmcQDEvaCqAQbDbyhHcxKKSs
YdWxaah+2HBd3G/gD62Jq0arCHJurTiuIoAAQrpReN9BE6hPA9ZpEc/20wkEUvxt
kR+j0Wf94p+g3FiESZEQ31u6Max2veP5ObqE5BIgkJPldZwxABDxkSLkIOWQRM+x
NTadXYwy4BpAw5rWpNtieDvV3Gu/AqEMzG32jGIv6X8W9DYK0thpBE0fM0sQNUyg
1Ytkf1qpCLlyPTYm9DybjghUwrl+v744lO2aVjDhPWA9o4Hm3uIExqwX6s63nWNz
2x1YIJZoug2DTez/li1z96oqtlOWrJtd4ucBP4r/tLz6FtL+H8LKTkWBH5Ifmj+1
ooOJLPEtT0NvhZ6IAW0xKIKDQeSftG61omUn8aIKEjmqDPb4ZzagSSYmwiDd7JTj
ooupDA0jNF0RqR/7izNUmxWCf3fYgdEUyfMV2PgrbEqffWqKO29ZQkUEtFrGyZT8
PyI555W80V9ALuUnnlupIlV+qi5aPbmeWyIDEc8ZlXeCKpqSCsDmhI4MgqsVRjYy
qwU8SZD4z2TrJ4IzZ3zrEGU7PKua338F5lJj3sdeijheclLcqVlqTIw3Zd191+fo
/nY0ZO5muFNH9uPiDLKfJYv1o8tIuLteTFDfHOXg6MA02NzQy0uJGlHb6npAiJG2
kkRg24VRyH7hPRiPf3tvMP2uaHwYMtl1IAA9eaAo6CUWdsis4IvIK8itk5qTsxh8
ps/AnmtmCAnf9RV4AgYpOXzcd3B3fU8c+7DGtjZADv5HOHaGKwewXN1d4PWyikmG
T97YStcf7gq9ZSZdqiwxZdwd1j35s+nFbCuJKoGNudfEl/KgLJKvI5K1mDt0nPeY
H6F+iqP3nouJFPjnN6QS4iHaecCTzA6MaBnvWhLHFPXWuvkLikSla0OPIMieSTob
tN0Zi7EZWK9AJBCrCBNC5teBG9d3tYElZqY0vtzFnD3AnNqHXPHmEbZxhwfmxDhY
sp4p+xVHmqKmessl22k9N+WrD2HqR04PY/xGI0H5ClbJY+i5HxrCaU/8FOuaAST+
6zo35XRlg1Ucu+KyTTaR2SUXNFEhaUz6Gk04EezhroT5O3NJenPvNful10mAtU88
r5dNoS9PLbJ7ybavZ52pxJBdaeXGoPnn4aOl2EwWccNyoSgtDnjfUYJPZsLKIZjV
5DFc/s7TVACeR5FllHKdKoPaKmqLNV9LgGgRitu4PoEYlacvKdea/iCM89CAa3TS
9MIEkWstquBOTNt+WOgIcQ==
`protect END_PROTECTED
