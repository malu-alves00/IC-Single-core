`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
h9XSbFMIT+gp7RwkyeGIkBPWR2GWB+jN81ote0gAptAlu6PBZdEz51pgt8bDxPaV
ECvN0s5LXN8HekF9WNKDV44WBEO2XVmvbvK/HDXPLJwHvtz/sjZtIOmvUK5mSnZp
JhRvEJURig6KvBkZ3wgBDGx7btDjoFr3h37Bl9dsYQZyEhXMMZWeaZqe2RDoT4Q7
OSTWR4WIkV5cSHD6lf4EYlqfy55Bk4CURKdI9BO+R848nD5MasAZyveytzE6XsfL
Jl/WFEDCwmRC4iDwOIAo4g4zLlQ93D188Jhzkpo3cqkrk/BgdhfK6YXn3T7F/YXB
Eyb0x0TgyZu9M2l3RI5E3m4pw0/bdcwpm3uf0poE7Ahit/LNFunpV7MngYlxKICV
e7ZG2SX0cDiNHOMxeNONzNEOy3zClm2pgUkVeeq6jkS9AaGoPDAabMhUBp/5+aj+
dC2WqpEI4Zio0gR1WZscw0gXc0zYnsj3EKpg6oOg8sTVAKsU3bcuZE+j6NLrlHxR
YQuKSUGjzfKtCqHCKwVm/jGk1SXFHyqqcVwJMFpEeg/7kzjnkxJpDeGaYWQDnzrQ
e30FmqXFLgcBjFyEVICyv+0GYhb8L3jLVQy9sU1QF8OgZC58Ugy4aXaMSgUoAWXJ
ou8I+L3pwg60LR/dvO46jdx7KJYDqhiXxaX9GA73UawV2gHXtyR4O951EuIAOgu1
y01oVb7o9OOk0w2Mey93cptk0rc22BY4sax4peekmDHalRtroOhz9YDyRHOquGRs
1TcfFCExcfpLcqCedQQUT5ATCeuA/94xp177C1OxGVya1Wog91n/FrfQ+LoFNveh
8EODcObaHXXHwp6J2iJMw4ncIl+Lf0dzyUnyoF03GOX6ocBfgByQWwGczKvXQrRx
haGYQ3AQTM3vQ7KVGIMtYr8P8Zb1lIhbc0NQGVjGHqv+cVjUE/MiI7ddESfk/ict
aX0QYV9bwgs7qsbDAkZe3Muf6HGNsloWAidP6UDWq8oSvk7N379OKZyuRuby6Kr8
cwanheH+AdbXqyUOX7K8Db58WY64JiKmfKWTrHPzAKF98rM1z6+quKW884e6meyW
UK7Y1bhY4Oyhdt2zEzEVG29NCI29CYWlES+mkHebgdknFjMu7UZUKNSMKsfM5CQX
rlABLeE0H/XRwtIHKUVQnW5C1lfzDvYA4Y7J3K8u0XsI00bMJKi3AiGGfjDlQ7AA
k1ILb+DGR442rt2JtdZpb10eD+MOa4ioFPnwngpN4TrwjhRBX2vjdC3LPuEDrNDf
y/AanBX1GIBJpwEvLCfdqa6Kfehv+ABtI/c+fxZb5l4X+xsYD5HXgfynYr00j5NE
q4YHscr4c+dUB7PM5h8sIajnvYtR6kXKx+hc9ANSUovxcVNXWmKo8xXa4qw1dEp6
e855GU8PLA9yti3087vZCUwu1Rli3EVeD+4AShA7+5m7x9eeQlSCS0bhAdzYcw8s
AWswg1ut5PgCoVNZMYjoLgT337OLu/tJc4crOjDUnhsEDFnGlmi8/wBda2YnsL06
ekNav8vH5n187UkCPPgH9ocuGEkruS1qiKvqm7rrtMMFDKwwJMKDm7FcvPgiLTtw
InsmEbp4FDW4NWM3Vu7vfQhz6dcja1jp8f8D44GP4u2FKA0VSeLnSIEWChXSUAvQ
HXSc0oLosDnRbx2pVXGDlhyfAeZy4oGIEBg14L+OUQd4n7KFFuM2X4fYjVz7IdOo
3dHDbZH+DWvyIvpwaK07J+c1z+8SSFAFpyytBbk7wR2dgd3oZb3Ex9WSXtnsh/pz
GCnyIYwnt0U1FlIA7g29iq6jsb9pYT/FB3X0OQD7AO9xYNjgWb0lLKbX0AhobDrm
NjI/K2sc2HJbn9816N2yw6VNn3hLveCqY18lkJ77rllF2iYQoHn3gmExo3IW7Whw
gqdcIFTyUJJZgT30beJcKISsC9zgcYAU2C3OO2dsllAlNh/C+TVDe50GVh1r4y4w
Bi85OQBiG3j7UISSA5ewZZ8uCrywpJ1RdL2o1e9Z9n6Q/SST2lI0OkfuU8+LRtlS
lqyxhuXl9HX/y9Yir7vRWFAfpX+ZLzYmgbz4RoyZbmAn25/I1pd3V/A2tdBv6bY2
Ax6cxrppdWamCrlrBAAmuXoFGiJUdRxBFxB+PHzX1LjfKB8Ze5MUYVW1pA+mUtoI
R1VgEnzA2518ScZxOCT4NF1A1E4PEO9YHpold3Xf3HlRWoA+zK9BdNsvlEMaHldC
4oqhx37MJuHjwjtzE1HG+VTu+ATJnXZhnpseEHeq88OfRehVzSmvUVCUGP9xeYAZ
bsibdUfpdbEIUFAtjYvPSxtPGHpC53NEFrvlghxcc+Gu77U7QqwUO7FWb5qfbctj
V2sqRFJApcHye1BgxXVl7pCQB83cdZU961ILi9XyM3bImihzdHyUS/dxSu+B/WCR
55K1BKS/palM8FsMV46mr+OrklkR2xZMaNkdIFI8YVZL1h4b3TcGlG4JfcgkDBSF
liSRITYKlHnxleXNSAVsh08cwp/gSs1WAYc8w21YONEbauYIAyeJkiMGRtEAj2xG
hR59GX/oRVPRrRL0M/qL5Gs7ZIrlZ+OdbVcP0snNwj00ed3qj7oP/uhGKK1DXmV6
TmtWB9YgcBnkU0vm6LfqVMSHHp0RDSjhwJDYX4d2bPQzEdjzT+Q1XFg6JjP5roiw
1k0AgJ/+taEpADHqYn9bbk38wks2AFQkkaBf16/gY2RMrBcLk+TFE4B2NedhPpCw
jDMNzApbucnZZgNohMu7q8KtHnz1rm4mppgOskBrmA9LBBPILNABKTZiXRXmNWd8
DCtWfzMCcdk3U7RBcK3nJNwVIG9Zn7MtfZEM3J46fc6mdo/x92Oc08ROCzLiiujn
NsmMctsIC6zuYWbTinuipb9YlbX8loeQ8uOZ8m9d4O9fSlJudJCokwvHiN/crO3G
1i8YWaLnzDhPz5iRbCsJCEZVxHu2aCPTrat1ioXQ0KRvhJTj87i4be749qOGs11Q
Wk/vZOlEvCBTvnG0ljMpbjt1lET0dQsHLNVtoGjUSeM6OgTQLX+6H+a3OM0eBBdu
A5240qWPAaeJothqJP2eW4ly4x2VrJ/Uh6CQrn9C/uttHkooARFCJL4JHZmxcIXQ
NUiPuia5CvUm/WGlfzV/guNbfpUz1lc9DAZLUX18IOT5J/q28w7hh+uPMF/EvVd8
IdFRS5Xht96f+zwIfq+fA3pbrMNaelo5Z4TWKvMZa38JQFyFfPFjXn58W2taz3k9
NLwWCa+VzNOuvXp38cyT0A==
`protect END_PROTECTED
