`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FZEfdrcJucPpQPpwMvhxhoQsbrInGCieRBqUn4YgpHeDkQQOQj5LKxE5OLLcRmLK
fvk/5DOqFx7xdtHkGRQRQBJV415ifs2bLJs2ZYVmE4eeJFrVixBhbpCzJWHeQwiQ
pPEbcHyQTe/xRvs8zmZ+WwjtzK7RWqmIO7ad1TaGhuPGxmOsKl5+PbfIW5sErvxh
gzrSKD3bxeqc03gyttnN4UMI+qVZP4y2465/T3NvF6s3A+fe9TGmyhhcxRrtEm+2
cgTNpkyhzJmsLzjdqIc2uwKl4lYX7JjdVmn4hKCowDPWJH7ysyOmIk94e+EbXWVg
NepYnMvP6UpoiImrEwzUOYKJZ5jfPf8uQBulR1qTVPsCvPnHVD0edRU0lDDZ7VvU
IutyvH5GqaCCfZHHDRtOyjChGbwh+4+OsJG4YSzaUyS8JUYl1rNMeJDG43dSPcCm
Tepjx3CrUJVtLDakYGkJBGmpYtd5xoZjrelbRi90lCVNldNdWU0+T5BmKrRszzKE
HdkbmDdtALYNdxQCjCjfXHrx3ZlgbbMFcs2Wmbbbe7cuNUTp4hQE4S2ggoxK3Yfi
7RClV5B030L2u4eSsHqELlDTchP2ZJ8s0HBzT1GGkGxxqqBcctx6MPs7TDn7qweN
jdTi365hg/PvT6Dcahk78uwu/u9l+vGFVF9OC7WbhUU6AM5YWYXEb9jA5pHhwC8M
vSEYOg2pNUfW8KtiCxxWzQa/8hPBU77Bbmze2pIss5iXs3jmWjFpLHGaYwt41b5l
BXuAbjCPyJi9cT0pY+xQhkyZVDLg9RC2q2pGfGX3CT3ceL2eb8jQr8Qa//tP7APt
579u7bpizLD2twDz9e2ASk6WGotxdUUmadV1P/24J8Yu0C9CVtlYHjWY9KqiAaoa
FThzdg3T6G4bpPAL7Yv4ZPWVl0IghNc3RhvCK2fSvJITMl6hHap18CUAYUL3Wa01
CZsllizuhhZL6USexIFld1Hqe9WA7ey7ZLJW91dW/F5hhPNjYlZe4P3zI7kjVMCt
QmhALRfaO0w84R7vapvJpVamifGERZBCO9Fpc5LCLWQ36GLrOD65f/Xm/waYSNa/
wzlCvKOH2PFtgILrDjuQhO25NXn7FgW23NlUYZajxXa2ipVdnafHlvySUbH3+GIt
0ex9sU8WFWUEUf2TQiSVC3zSul8r0al49tck6AT2+UaGoagNcrtARXlKbTjLkp9C
`protect END_PROTECTED
