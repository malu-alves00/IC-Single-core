`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UP0O//lag6pfKI8I//LZgBz1lkoDPsbtbZigMrY+9Ve8bK9YRAzimZiNubGFemDu
NQMfzHohKUvDy2FPaxyAize1BOgKSV6wVcktfZZd6N3szZfbCy/qxl04lhTi1Lpm
cPMwjt6PjjlRbPV78/j6rfvdWgEg2tt/31Fna+Q2XNniywvnaakiMYASyeC5CvYN
64rya2B2UWtTx4mHvgAxI43AeTVEcCiQPhlbvLYFpUneyEFhE9HxlNfb0WGsMXcf
xHMwDD/WusHNreBRZHqVM44UjnX43sfM9s911wRm1n7hyJvtvekbKMXgKAa/yYv2
UhEQO58Xm6FeQq4zKrTkpzcPomGMZuHQBJ/9AkH8k5d85W8EG6g9Y9Dxpk8ha1N3
hTnv+r4/Yrgamw2YTg6pGCtLIig7XPlGNcSsnifyMJM/baFkiKtRzIzd+EbUQVNA
GedEZN5yhhEV5xFt4kBIDifPtE0ScU4AcBi1tWO/Zffvy4IKrGsEaTJUVdPk+/Bv
cWc4/MccjcdBrth8lvmXve5KMQ+XzVeskWNTQ+NGWqrKOMFDr9ZCGvsXRasW275u
xC1RbhSydqOQ5GumET08NhsQdKuooEAldfj8inkkYnAQcITy6e3SDM6ZB0yCg8yq
hkNVMEeh9CJM9vBtCYD0ILvQq1PkQYoykOjlrVQSc1X8OD+qqUxSH+fZOjDdiGS+
eGq6YYWSB1FeXVpD2fobVFdJRQRmOwZXgVhPC8skQyr1eLepNCb5CxTDul+kRqcz
EgxkzqNHrEOcdtgyD+FU7nji8O5okoX3ug3kKY/5rqVZmPAM/5J0jHEu5zDcOnjm
f4Nhd6wiQZYi3l7TQqkGZeyQCqAyNJDGPJdrgmFf0o5eA6bVcBXAQt+NBeBT/+AU
CRGMY7ClRxSAIfC1FJM0HhTgYJzARWGbFopn10p226Ly5lZsQKRAHrUQMhLxDuhr
JEL6ADAu9uShTlKzSmhR7lwdIC41v6xjafSM2fXsXxmYSJfjgy53RfBw3DtRt8Qn
uT7p7wwhjRzYP6WNnWepdejF8d5Zwn1StrlxAH9PuKBs+b469GpGNxdVwH3YSFd+
mmszZrW4A1XGWgLdOaTyMYNt1MCABrXOx6OhIx0V6qA68X3uC/FxPTKuBybhTqD/
iu96o+GnjvrMXZZWfWsu1P5APbPIzcamcwpsq+LKn46fCf8s7TsUPXT6JXecauZB
TKs8rXlz2LvLdrWnMaOSuYxaJNOojyji1aOIznDKawoF2J0FEzaQObatDoeYfMYo
vRlfZAOvQP+hqqlN3KgW3sgslbZk7jjaL8NAqCDhiyYMIXfqNk50bZFxKRbh+Xg/
hPHMIkD9Yts/6fbqQeobor5yFDhL65/T2NKubvwOYk3vRq2XpCzbVO+/FPKD4JKZ
WOTlnFFvyibsHgzaJJzbGugq64q2qQ8BL+Y/hwXIiCMXHKZ+BSkxdhCVBGqcFBXX
mq4VfHsLilWECt5auZEfmtsd6Lt9PtgnVZ/yEA8uL3NREqs9qWc2DO4TFWjSqStf
6RfxFL5i1yCDKVOgGdwzxmmzaVnIpOvAJW8l9EHiIIVR91i+UCEgSFSO781IEEze
ieu+G+OohRpHTiGckY2XVooQXaO43B7dKKCAG/2wKWAyy+BOcNUUUx3LL3Ulk/Yy
fXrozxiaAJBPqDZexRyS+8vu6ntfhMEkASUezr3ZPrreDO5ReZWAR1zXlSBq82GY
RJJ116c79vUHxpAtqewSaEXAy2pMrVgf6Ry9IIzTDKXUAZoE18mUXjrqSecScOfW
sFFIMObqqKhs+kJ7XIw9qNaAbzzhj81rKkbqsofKxZTkT4WvevOqlhb9k8FWLr1h
duNcHhdlSTR9uwqA/2DeWaI1aTToAs/mZtWBl15E6NoTlzRHU7PAPE3XlfddHiiY
ROQo0cyeAkzIWy+orREH5gx0UngaOI9Pe43/bp6gT8fCA0ca2yQ+/N+j1WAWbNCJ
ZenMDYmCNyTa1IJm7/1OEi3C0lyMIWx6+rtWKSVYzL4I0dk7uANfGYYqxJoGFB63
Mb5UppD5HBt6/dd54b6KN7MR+yRQJ+MMETSSylW1/WHcBVoaBAZiYOp1o8kpqgrv
ol/g6VuMPx33nw6jX+8fMCPrOdDBwlvuLNRj7FlC6ddTL0/5MiR8cvG6b1scHnvF
ZuARZM1yA4ybEok9z4chGXdZjgZh9cC7L6/MTuQ6qGXLlTmxhQhGd+pmSF6O8ckz
xZK3FBxKhCvEPiGoBa6n+sbCbJtvd1PX3LBbdmXDYEylUyiZrLRYOxUVdov2eKkR
G/pzLdKyR5ql/fqwF0+bnop/FFwLVS8gkE93wi6pit4ULfeeZ9TG55jFKPhMqdxd
/uxtzrZWPDOCnxSOGc3mIuMWIw5UWjkJ9rf7dnCCNxlDquy2I2NuVyAWrETe43Wv
01suS0DPQqBG2tY3ZOIee0y+ES4tLQa21Bw7Gw2lxbCR+UHnbPQOswDFqF36LcuE
P7XcQpXxBC/dSiKBY2R82lHrheV+cMp1R6US8sMH/Jm6+oQBprQJFl2/hUOhGIhO
fJW1gO2G3RW9la1uTQbJ2zhK62wW67GHNee+2F1SbojHVEwf9MnmAW49NguwHjEh
YYYj/eha5Kex1MD4CPOAk2d/etofYO/8gTCgmho445CUgm36948tQm0Fq2XrlXfs
z/Cflq2d1H/y8QEd5v9LDPScQ6sTrmZuQnRto+8JD2xC+Uy3IoW+aborgdRS3Ze/
jytqDGANVLvKM9O1poEDXWR6u9vRmJWOwjOWqXHgOKLL0u8f5QBIPgoZjsQpFdiG
PTe9vzDAz/dPTnrRr+b+nvZ+3lskEGVthJcKxV+cuE4tVF2LlMjfQE6smeBbloB4
KGswNIBF8RpVp43DlX9fl47kc66sWQ/E5sT4gsbrOE6OVflIaC+/f4jBhM4NN9fO
7h5d217xq2ygSysQfExlXbyYndpmZExcKVsnYX4/1sjfToHRrx/SlXtCNFLqPiHL
0VZK09ZheObMHhio8W21hT2BH0hRZARfTn1khnNvDKBDb3MX3wd8o657SLvzUyIr
k8oALXn5xJjHSqN95OSJ3NNchx94yHP1kPlscwW1TBgKu7XHMWNrpzk0TpCHwZ2j
Gii1d7wNrASFnX7DnfSDO+VhVtX0BtGUg5pYQx8//Otj1tHnRcQQzkx4ELBncQOj
qosHBAQdkmj0UQHR7ufL7GREEBbO1ztvqYhg+C2+kKivAAM4s40xmKnvRswZCQ2I
OJpSTEsHHWnAb4dEwxkImKbD/GNlH9+zHkP+v13oECYMgZyuSzfesJguOWeq6+Fg
zJy7zfQXg0r8U/jrb0bkrFc+HbV/7vJFNv90jj7nbpEHBOPfQWnmw8uh6m/P6LQq
fW9wa2tXLAFmAb5+e38TG+rHBrcnURDSw1aNO0ARFSHEpUa9cJjPbX7GYozrya/A
eRlfw1rA9Atq/B3mMiYzw2wZwaK7jN14dV5DDIeW9/+TW8XQLnqvoRrZPh9NGDMu
RdReq8cQvgko2b5W2h6iCjwFDNwTRPCl4znA6LrQyfxs/R4tk3mnlXMk8DDaBD+b
305lNm4M7r7q160N0RUC8ar8T961Dan43HOyjVFed9fX4SGvvAybrH9k0X4z1ukr
1NEZp3B53z2ETSNxbYydd4Ex8ka3BuhWt2+yH+r78WBX5aLcZy53/wJkqInblUaf
zDiPs/llM2lf7tm/QGIxzrREeJHkbhQIF0qnz0vmh0kfbUBvUv8vHhPfl5pu5K8c
pimCGcuo9k/OX2J9WL9UDcx0D4OpjCkJRtWxBaMiFocMoLPGUO91TjPCtaqrwEkj
qKJAN08slcjUTDeQeY8XD6BN2nD+TM9Rc8U4CByh/9DeBUgRdtF8ucMxTjF5F+4D
Pu8oXi8bsJ1paN7iXXXt/GwHdbu8xG8JE8J5I2se94c+amgU82D9rGME1DWa36sT
3Frrtm0TURd9F+0ZNtum7nZDQ4bUk0RICrA5k5CdohDzfsCV4brvN8UO4m8OEMxy
p0xxD0ySLe+A+fOCxnn+4+O+ElUVxqodqqTml+OEWTL9b6vGDYQkvYcTdcNvcthy
UQMywlyyCVZsMaAU6uTCwq9JOJoPwgJpg1kW0THb3F/NHvhZL/6RwVQVtSr3t63N
`protect END_PROTECTED
