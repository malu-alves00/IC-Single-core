`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rITYszKjZQq9U8p8XQrgpKHGraGliJKxPBLiW3CPJVjcfLpHILxpnRiPnr17ECep
EUsBQ0blHIh5BX2FgVibbGVSH2wiFFFPWEtcdCC1FqYEFHKMJFElo2/fALfi4hED
c7cakUP8w7wMdtaZYF20zCr92YZRBTmnkMYyT9Pcj2yv5m/rJbcGtlo7PGQNnqKa
r65RDTOyIeWoYdQzxTd3ngtomtOnkeXzmPH/wGG5QeC6ekuJiArY5NQDenW5cQgO
sryWo9zB2uVKU5WJyvlQHAaBDqBLU6cGtRYshiqY+2/M5WQa9kS5lhCVEgMBhC2F
XPW63A8ltMbP8kDPrGDNNwwZRPWnM/36r0oIQhHs+icIANdsxrGijWj79onqFqxU
umsGrXyEdaenaB6VrIwmBXtBJ+Ph6L/GkhwhfaS0aqtr37QMAyoMRttXxXVB/f1u
fN/502auc9cyfQMOSsJa0JgZQFUoOVSYRuDNwlkJLjV0qIjhbz7rQPObq9lX5OmO
tlew15Q7ltxrOp1SPZLr+wHO4STrspTBGFmCGco3km5814pzrN4ZqgCetGyE7gsv
gBrfVnwQS1wvC7tgrpND/vyUoeNEkp6bZFyGx1d9+p7rRMr4Smgdt9301L17tjtM
Y9DSKgRnwm3i9n4chzLLijBCJysPZLqrPHHsSAZNv3EP8VGJ9QojVUov7ovV8j1O
MOpTdOTb138hBqWoqn9tU+NQM4/Kbo5MjFZ0TCzzitZO1vj+J1OufYqq08jA4CTa
GqrzfsCEZWVRT7QqJR4Iw6gHOC2w2uQWn4eJsPsesPbRiRu0Kz74VYAue4caLjFM
wQgQWBXVMGOmH1WSsbFt2X2mvBJHQEUQhzXDbUAA5XFnxm1IcqUbcWds3Uc9u9fB
slkMDngPxLhR85+fTXoB9ZEI58moC70glHcrD6fSfehR2wZnZZUsm4voffRE5hW4
B6FLa7frh/wbs4h0o9FgAvSuP+CJcn83gwUPJWJJzwofLcygTRMnOkKvWzJdVqFv
J3KNyJiTO5SCharPTUcG2/Hj59TPv4E/k6zbtv+fgt1P/ngvTp8UCNTA63pjYKSs
ctOx0kC2HmpY3MCuXkwPicI7USGS/dxBTYwKmt6TogFfgaOUxLv32sBWQ85O/ujG
6qPoH36YF1jsYg9di4HG61zpqqxv15o/L8Pv5Zq++RZlRjt7MKWOsGfD1k0jYwAd
AzLm5ieWamF8oy27EIqXNEYtfmKE0dW+RqylD2iNh3opc8aL+8vFvqChsiBOzfbB
p9bVBd+CEGON9ldUuJ3ay1AfnDSVeHXYuRt59wC0ouJ2ZRh6HL/SkEXeAZyfKhUF
52UljrwmbTb3b8+gjPZE76aYmM+wrJk8i4NnWXmIutUWY4C2//2lU2ArMMo7gQzI
DKgncm2vPXojGu4T597qpfMdzzdOMPSBuGf8fTGtDuNydZbaWuvloZiT5Md//elB
d4e7yKeXGtkYPBzBLoA57w2pWRmMo/+gHsZUnrnKqJfhy2/dpzaIxlMaoMJ2MfF2
7KYDCBg7oynEIISWnZu/90DHb/RUU9bRfS2Szd7HbiTJcMQg+zmLkJOX708JL6cs
n9Dy9ZwX5IUgg1h4VNCgiBRMv3EvvsKOyHZJlwQsaAY/G/GM0lkTTK/+TyC8/mXm
8IYSkc8hQ1tnr78VEYSJ5FSQxg77C2dbZKFR8FlUSbn01bCTXjkNgTH5zO3mOQde
1VYUQFplHQwaHT1uWNOhxIeWl9BgbhsoTz/icbwZrIHQtXB38yVmfd/dcB1bba4E
YDW2qL3BJc/f+FGDowRmCj3yvTMrHvg4ULqy9rtGix77satmvDj6Dzc6cBf1flrU
R6xTza/D8I2CepTrRey3xBpamVj/19zKSfBtJ/farsqwgsLtdWr9dfJqE/T83OUQ
POQJhUlPz4faLVySNPRZioEQVEMMgL5PBhiqoLv+E0QYzD5BU8WlT/WLaRsk28qZ
7LLVaVtCj9t1/F20b9Hb6YQ/Kw0cKYmmUnLF98POB+yBkM786musUZl5ntPs/RsR
ivOPXjdciAMKEkDpVZyFAYCxe0Zba4BB3Pk03cmq79E7nCcWhrFhwBNV1PUDTB+4
MM79yJmtXSwuy6DLkkIG0gDX+uy2KzaDVK/tBzCPzqJP8e8aKxOcr9ErYK9Y0Cs5
L0dkU0RLhSJhdM6MPtMDum5nM1p4HyhlvkuXIJlXWT6QsFyKHNff6ei5EHcdg8ch
a51udQLjh0dlIHAOtY/CG155dcvNpscp++ypP3ytsRSrS6mgMHVK7oNetdlpW+nC
FLrUD64uXe5LY0Fn2G6VglPqK4OyWroXNzHtN6jgAE4lRUuQBaYVdMj4n/DmgeOS
EwxBDMRvBlmQybE6/8Q4U0yW3573lYbT+Dl9qTHFCUBfW2Bzzii8Wqytd3TV45xf
mHBqMEfE6boZ4vM899u0+pRkxnvcMIaUxRT8UKbAjx78p4stS+3gtP9THIeE4N8w
4b22KT5H5BtWFhHju9LzgMiUxQUCpMdq9KCD5bHd1RRl5+vAP9Kk4MBuNEQP9Gi+
yvyiBPVQrrow5PWBG0AYcyzTNf2VvzoNbvO/psclZI5dcbYBzhuFvJXwJ1KHunc8
gvQnJOrxHudwcR+6WmdpiY6/B2zSiMNowA8VaCW/OjthlRIhHvPM6e9g0Ed1lTp4
6lnWcrBo5BFnuJ8FFqaJAzPWYZ/iJiYX2n351hAukl+sc5OkLNGokbflLoESKl5a
QaUQyF8cIrAo3kEBRE+8zkfvQ3NHyfEW+Dj9klSzUM5AHg0Vcx1KDmXwyU/HjZe/
2fHD7/R9pCr1S2GvYUd6sBTwG+Ls/y2/pfeL9Xv9PjlNEUMqLp6fI/jZNUf3jJ4p
xN6GIH8fKl3SBB31HBZ/XUBha42FeE4pSfPy/fxUYAdeD6d7Bkq5dgKRLbBTW0RM
QEsCy7j7OMCNEFAPpK/HLkTEUmzIhDU+h1G9VztCOZT5Ew6OxFLvc8YVAzacrIIX
E0ojPJy6u6/l5UicKdWDzdqtMngE3mNTKmIg13R2R90H0BBveV3geRwt+I708azC
uOXqRs6K3maozNqFWw+e30ZCb9WOgS1mwR51Tl0Zo2kb2gsRNjMDM8cb1MFGYieZ
R9MKIZiPnLdTwDYps9shVqn15/35pzigBi9idb+J0n3+bROBES5hHEsKSA+AYVQD
RAsv14g90DzFOAIoT5Ry+zsmzG6HgokTaKnzeYRmuesagtzgJ3zBfcZqmBCNoHFU
GElLV6354wg11StgDM/583udgPwIXIxl0m1cwwyZWVRHTk5b4d78tm9WFwILU3mw
JkoP6bcwuAOyn1Cfm4KbdIK6/POfLxUNWk/pJV/S5APbpibeAqCbaSBO5Z0yLriM
D/PxL5jH8xjp+N1K8Xe08vGdD3OgIEHF224GJratPDw7Q3ZX0bhrQ4SQQwQeMzJY
kVUY5kAFfpmPnGj9UqnmA+TY5cdNce4L5gvApdC7hU1aLdLBvkjebHBVf9cvFFNm
5em1OSbvZKUeUSRZ4cfa3oqVZwa5jAcsYiAsv4hYvvMBmdLpxwljPp1nJrB4b+eD
xNQciTzjXV0KtrK33SDbR3nDDysf5BdFl+IY6etrviPAvDVDE5AIkgOIUmdEZ/NR
MufVM449Du3iQ2rR/49qqtRsDjdXK3uZyl+s2YE94oGZl1te22FilvTDPyDdzCHF
RaxKEsxJqbbFaJg3SkjHrOFlEr6oOjkqUZnmVwP9o4c+NDFWGUVZ/hOjwV1o/PnY
mABKtiUlw9352qDwNzzsr1SYLezq1o/Xi2dbjtzVfXoYoM6Jn9Z4bYxCt+xltXxn
SxzaCFARGJjhYo0qodNi1Q2Ne0Ko2IEPedbZThiTNvyf+rAoRQk6MBiS4YHYxRwH
JKwjntmQHMoL5EK9m1sd4Ibw0qUjf/q/O0QDN182iNrKPaK3ozW8m/m+sE1xgifH
7bvtgRtUry0DTv5L14zwKQznrJt7k6IH3lfgay1aPzzhgK4e++05p4Ea0IJRsogL
+0wvy0HpowswW8TGkHKTGvm3AwGYhHE1kxUQK3UriLhwDEgK2xYieAubAqciS6aq
6iln/VuHdeCy/kSK2hxQ4aIuVL1rWhbJLi9K5r/b+kVfW0bQiVxBGAmHzylE1L73
KQ87/QZnQk8hb4xWySMe7aolaJTuS1GI8JonUHhZ0SXSBkaobHJGDEVbkV1uxUmT
AZZEMClhczKIYTCNohtsUemhs0j08UpjQOjVJxpY2jLQdRR3q1ank+D+s3U3Ywsu
h1nTjOOJep+yjwBV17Mxls+Q+VaJ6SA/RKtWtZotr6XXxalaVGxnjZ1jQ+6ZJwFF
ZD9R6v6vo5Xm38LfAB1VvtEwEJyCMLUCBjzv7gbmRpeuKGBcNQuD1xSrYYq3om64
rN5ZqtZQkoBIIiZeLei1Aa2GwRmQNPwGVkgjmKwqk7V5ALfKdFWqTLsKE09kF1R7
SWQx8djLSb/7zmJpyh0YEGdEdyKMwhptpPiUFNAniFz3SMqjwnqjSNkndReW83l3
mCrobQYoywQQkX8VwHpFTAd0yDIUS4V+F3TO+b6LXNJYu34zkpa2fU0JHpy9rIiM
qfBB+b41FvnN0uta58sdx3TooNS2+FsDYkcozj/25y4Qc7Tjlw5P0x+K8hZsJl8z
K1V3cWudjvi0Y5uoKP5R3+cs5xmlSs5HftkBgqQ1eBhYOWk8xgHEkTB9CZz6V7Zq
RrV0JcXfCLhA44U476ZbVwAZtLg3U79bew35f3VRq2qmevAU61tz1hXgTO/I7BrD
Zkqe6y8NysP3/flA1XOo6OT3K47zZsvMRYMo4OjslIT/JG4oSbpmbgcaiF8nJ1m2
iiBwc9mfPhv0rzJroKpKpjU8XWwKnZXNAvdsIS8Y3BkFP6tKu2Vxr+UwGb5a0x5S
BJeUixeIW13n9q29aTjyR53VjB5NAL6Rf2MQ3yb6Pl4G+K9i0OftYnEzQ+AV7trP
f9fPjKrjPEA+MYRIeRpEgHBMrqP9Jsxs72HMIVPEmbtJ1FMX13dMU5qY+9laI/3q
+hm16/YXvMxFaFGA1Fepvf74m2RUO8dqm6vonwJEA+F2R7ZRaBH+6hGDMz0zQd/8
Iq17HKm/rwkZK0IFEUXP9RPr3dZSUyLZCHysshPpSOebTHCtXlPF7bnDq0rNEtV/
PvryLL4Eo4sDBFPhx2XvigwvRxAOxFhJkc3MXvwqdt26wwziLQwdkPXGEjLdMj1h
peBOMepR9Y/by+UBGestBz59AcW2pWb+aAo9l3VsA1WSwrWahRDFTVugQFtIQV2/
`protect END_PROTECTED
