`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
er3xZhK8SXpYTJuyGcHL/rTxCOj9Z/t3B93Hbq7x/l8qU0RoUjWoLQ7FFMEFSMaN
gQVkL9PXAKcW1UIuUW9FYYcIWLLQ9HSY3SC+6pJX89UaqdlkA4xFc0+igIKjrJpH
3zwe0ZXynS8E6NNb6zIfRPPQunINUmLn9tpp0mvgxljvjWWkYwcX2SY0/632xKxD
pOEd2PuX8vYZ+5+5D3R8nrn8QKelHn7I033u21fclokFEfP3NiYe3xvKW6TDhVFc
mIiH6aSRlvK/ArqOlVuXg4RrKQHl3bsCmIBUGT69TcM6KBtRD4zHGxR0OGhswjFt
mL76Fm53MqH0RWRmrZ6hYI8LI6Bk9CW2C8xRfDhR8yb4drOM++hhcHZN024tzzXh
oq+XudcxK1QZQhk27IZ5uCSpOcXId+QymYtHPlmG6Vap+fDlYh9/2KhnmRgpy41M
AFwyOqqPRxjWksXZ8hSZw2IOgPQZ/G3EgHdxP0wQSaBLEUpsziaHsjLr00kpvysv
osWM58+8QLI98tKn8CS7EKgI+ell8udpYaIcVJVH7b3U8Ljmgt+ScPdz+Orpu6OE
d/e0EYbT/Ig2LHtCkE2G/KPg6IpWPFrAYTblNikYnMpu7mN+0xNaCS+rcp6TGA2W
GfGiR0G7wff5wLvWnTn8AggWp1WBfncVd+CCph8s65Bmkme57U6gZeav5XtVYP7o
JtILb09tfNsOjSFtb2xn04h62GjocUnxmSnVVdemcnMmMZfDm6MFkjxOmwXXpmcJ
vkUJfCPW97M0GymDBM/wo0Ec3XHDopBmJ4UWrqHd1A88VFl1ryWIrB8BDKwyveMX
GLXiuvlkw/HTpuFGGa75g6ule5kv5l3G/ViAgOOxT2aTpyMLXHBwOPVbvFZR9tX0
C7po7tHTcyXi1KHZ7p2bvXoqPz4mQLpNXrdjhIa/fiFQ1ibO4QI/8l+FUmotTOf/
5gFUtNCbvuZMmO30cwe9L2X21zoUi4T14oTybCWkmvH0mYLEvX8T/uG3z2N6sbr0
lCjp8g9a+ZflmvJEefNUGhHLFT9Wp7a1iOBovrPn2s1qtUTAXW5Ytha1AwgeZ29k
dmI2TbkBF4wSFzDBvoWBABJnyY8R61+TZzuEBI9FnjiYKOyqea1FUHpEmWwkUiLZ
2pfozDT96lnxAC2awcq40iiW2NFslP3NjieWNibusJvTPzMXMxZq/vasfo+tM/1p
zM3llUSSiP4vyoWC82eheAdb4sAtWBiuDp2AIiHiZ4czcZ7T8ktXxJJzgqbl+sul
KA4ApJKttG1uEpfK649s/uIoezL6BE+HrWv/lbatXAvRgBPSeyQo1O7KJL+ADhg+
7Djl+WUfehGjWYnii6Ze10UmOqGveEQ46OL0xrKEjkRINJmP4oQ/nO2RieU9dKlo
Ef7PvUpKBt8/1G+LfeIkLE39C9HYgCvoKJuwbSV7m9wTMGwLWaaJRlqnOO/hfnlu
L7515LRLRYrN51FCDBbVg6o1tFOB6AydOaPMDv84W7s=
`protect END_PROTECTED
