`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
E4qJ308ecHKPy51YUK6Xv9Bbn4xCqhgIY8bv61Cmhts5U0QW9fX9+Aq7eGqx+eDn
YUn8Kws+tkWf1iCQ3l96DWfK+uYVsT3YICNnKovI2Zxr24PeoHB3WqQqwxG4MIEh
S+HZ6r3+JWYPuRqMNTlBH3pwgE6n4fvSXCWNX5oXyL6+jEAa4Ub+GCWMpqnxKDj3
qBAc3OgesC46iTUBv/UfqsqxlAO55jtcxyNlvNdfQ+xGO83SQVD99udsu/yx4oG4
cRvC25BmptUJ1T1Zz901dECaJdYZ+KpycVhOw8t08NQfb14xLUdL4rZoj3oGPide
LO1bcm8lMK7NC/8YyyfmmL7tAAJZK6VsCVeHmrpZpBtSoiREDYGQDR8hBtBSTajn
5LS5sm2zAzS0fkFmBcqjfrHFfrP9EZZRfFg6F6rKtz5yLvQDtklswMIoe/vD4UML
LYm7RSxgKdP3Zs040NauRYuGWpLc0NRbE0pOcUTPQSlbRB6kuMc3OMa8AtO+KPJu
Lte5cUS7yzylJwI3JzXHPMDbTZgpYiBPX6UJsimhdUJ1b5axK9+fDr4FmJ6BJBP9
Vd+z50tkwR/vSzms/tlogCNxeOl58czisHbNrLTv2irRmKcl0Acno0Cm90ZJbE7K
nZdcPEKz0WxRc1P+6J874XPk3E/w2uZyYMp0QGg2IQJ+PdFE3tPHUNV82MnXw1zC
HFvDOEv/fv/jrMt0xvnpDBXvCdqVyrvHKtoZLWT3RrClwWiofesOLWStede/GgWI
WcnfT1NgF2Zrt8iLJLYaIlQqSoR/HmaLO7TKjOeJObZinkMds3hhCK/mUEwl+Tbd
PkAgKcpqfZWxCXVqITk6Po9q2l3Vic0vnULjxoDsRbsFns3X37CCoT2Re+rx4vlM
Im/lWied08G180fSd6/dsrbd12DKYDdIXxPyMZMd1hLlahsAqN0gRt0Gn5o+yiqP
KK2IAZiUQF9uk5DN7+1p4DqgmG1eQ/Bvr7Ouyp6Lo/hQZ3nu1DyjRI8Y3kkWCPwI
J/K4OaUwzzp35XWCy550Oy/zwnwvf4sKhFXfA6qmN510IW3+5JJawriy7L8U0TIB
ihHoZA1y5hki7kRdgPCkmeCgZIXoZCmHyrwjLkNz6EMAEW3dwUZHCjAHUVga0fKW
pxhoDmSmJXVi8I30OHLPwXm21HayONqONPX8DWCd7jy1wXnkl4EtVLXUcAK192+9
UT7mWmB8RGMCMjSpuFiAbu5K9ouDfZY/mhLZ+jvYV2LNTLe1vqZfy55WbUEwhUCR
vPewqD1l0pPsMc56dL9kSBEuGZ5qSYxhY/O37l9ffilSPQs87aI+456Si+6YjIIj
bgc5xCkbB/sEcd6YOQCGjQePTtd5LxJhVJO40tTD3Y6oqkT9dWicBFa/hBGi12yh
Mez9RMtstdwWHYR5+UH5m/lTirboRIalZZXGvLTucdZCy25zkjnW1KRN9KfkVIoS
zc+REWCvc8zwsl9IuZEi16sNSQyFTDwPXGM6/DKLGAuscB9uegs3f6zwi6nWJpt/
MYbT3wvv3Wpkg9nXaOdGHmRBGlPg9FiLwIzQm7uvp1Uwv163c0gFabO6om5rjjnX
gbbAtFYBtx4Fg77JFrPUhEtDcRFNan240sJjr+EoN4u8HndIbzZlehRrp03TuHT/
+0lI2lnGEGXE5/jeJV1B4KKDIoC1pq4I2rjw6W9MxDSB/oOGcKTFoEHQM0upvUAj
pLp09kLkEsKcVsUJTSFvwsaqCL7ofP7roQ/xHWdF86HxqZkrtGxY/QRMzWo+uwpI
9zK0lHrDCGWE8/CqVKXlzN1j0uX9v5YXQefRCcCuCY3MTOy+2DSE41Kap7Nnxtor
vIbmd8jiZ8B8euT3+L/6JH3LXISqRHtIy3ENqugX9wGFhMDfuULChTsdmaxaDkmd
ToDWGqFcd6+DrMaMVk9kKZKhBezDFSXwf0OcqPswFG+qMp9PESOJgHmVRMoCXGGW
PqPvsDckElsHdvdm8bNEhYbObkOG+kktlxYumcm2fMrDoju3KYT19glXKttGdZ3s
25s1h1ZiVX4WxWoSVbQC2/Qw/k6KH25q7p0pDlFiMU+Qjj44K0H3j6AEB9kQISI3
Ntmh5Mu3YRyMaDjkt9u0uxyShz7wcG8qRc1ZZ43tknCLuYfPk6CZm9KGuruZ1ZAh
USZKhk3M5K/pdT/ENbfKxM1WgcYCZgKMO0GctPaZV/Gg423przYDbLqrmtOnIAQW
gpS019+k5TvtlMl8+lg8fgrQmichvsp9uQ0Nq4DUhuUXAmmGheDQdweGZ3mpjJcJ
XO34rm8AXfuPRyv+929hP4l22gUhfI7er6DBxAoNq3x8t5Jv6MyMq2FGTZDfsW9o
eqrCSQ8H8xEW7LNkzqqXLappQTFTDluIVulVw8jXMWdaNxyiGSSVPDLjmJYs6cLu
2UiOT5M9e6XrvtVl3Xy4H1ogGDVgrmL9p1lyDE+uV3BItg6H2NehZpC19VSGEAS3
V3FPRT088ks9thUP8BFqFtkFPOM7eCKXSNu7N6aYKWlIQ/hK5dIkPR0vDoKiuCiQ
sxE3ipSZogJGI0+OtgO4puR1q2PwSW4Q2vA2mYKdo4OwWIhVwbXAkf/Kgu2dlX9c
a+GP1pqBGjBaZkWSqyH+okxweQSm8aU5CVUvqhOAXqDlIEBaD9VXmxHv6bZ/7Ap0
5cnq7QQEJ1yTg8eG9qb7g8xKTXwb9inuQe3CUlqp+kw5SfsFHXgoYkaYmCLK7AyC
SdYkPI9UYUeOUavg2jw73LWnnSRpa6dHF6H0Gu0aNumDv2XK/CWVsX3CqUGB7YST
ACWz3TQpT/Dq25ynvtNav6OrnGKTB/0k7vIvuK/0zKbe3NWl1L3jV8oXl7Nzsqff
E0u8px9QqQvp/m4ExRSfo0Fu2/LvAZUdiWEiQtUxn8Gq3h1By58pOe7V2WsFI69k
V8YIKIb7XzUcA/MDj5zuGY4sgvoAXHFNpnMo4uGrRfdJ7c4BGFk7IOzKbIOXMX/4
bujV5moGElK5R/krGl9ZZirUZ+B4rK7pjzGaALdF+1u7BAwX6uDeMLB6wat1FVEF
ecuHd6lzlPUQQLHCFm0iB815dGFTu+8j5Z5Amv4sRZd3X3chHF4OnMTbSTKmzmm8
tTJab8XP7NAKSBRx6vSxXJOjxOVamX2re6LObaebnc0G14UWIO1m05jDm7iH/sS+
uG6OkMOC3WYXiBMJ9oMVq1JbggYvj23H5RwfR0ojqN/i+6o4GaoeVCbun+g8u7hi
0CC8WNygrdGZNo4+vtHzVdfY1T/6PEIFV08+j0uA6cdKLMBrqNw7Nq7T35br4hZt
MXWUQwZo+LuPg8acj3gryAqz0Ori7xJWk90WRkvfxzkGGj6ca4Y+IHE2I4LPhBs+
c8o4uPjwvMfzhIRGJZsg/v4lvd8cx5CLfpkN4XVxPklKSTunwntcQhTCflcCPCP6
`protect END_PROTECTED
