`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Z0rH+Cqkw7pWJULW6//MFwNiw/q3rjVDlO0b3VwfVoVap+iDJdWC+IrrXVyGz2gE
ehWpyr28wHI28qlHDvHBTw13/a0q0z5WI+uoMrAJq+Teq4DHCy3IgSR5D1mAN6fS
FlLPs9nx+UwoES5zvLoAGug/9lGKYTJLZgea2V03nCBSn+HfMok2OCUU/MEs7UM8
QafYUHIm7QzGC/p3rb6invLbFt+r+U7H8B5jecHgJD88ASkkBZkRyfsUz3rFFsWu
uXNO/DT8fQDGhNnDbcOkeORTe+9TriiFz61HLia9e+Gk1TCZx8o7YI3/cF7VpKLE
NdfqSwCKRFgK3uDW7n38QZsi/2UwOIZcNT4x+/atLHJZHe5flm5bEcG9/kx0fZ1E
7KiczCbGu3lFXQB41e5XToFUMmmKaJhYk+XZBrdW+Wr8NbgR/gEbM0s7nC0BetI+
Lg5FyWoOrRovkUE3cPgdPt7+DY6hZOhkG7r6RlR3pUeiU5D1R3k17wrMxUr+OCBL
cTfiGZmpnEAg0VzAY2hNz1g7IwrotXojco6Jz8m0L0argZFbWU5G3sbbHQzscK+l
b43XPfev4cW57jfokxmXsl2EiawZc8LsgkvnZt0qeJUjkrBarh1fqWyfZdRK1t7o
pSvXFp7Jtuqgy7djoCkNLgcqEmF7oZI9tI2j8Eq7/QJkdYovWwD04Agpb93fLuOL
stoFunPt88rQNm3d4OyKJX1LkqxT6uqWeXdHi+Ep7DGX8TIb2iGxYDHFeCOCd0IO
l1cJPv6gxQT9uQMJUUapGnR5JKZZGV72Gorstrlu2Eb1dJqosw2otMlm8M/ujOKu
d21/6iSuclfq7ZVPDgVy75FUyiENj9uiDsYp7rCNcBq8fHOUSaTu7ueKDLPSpo1j
x8H6K+JzXRQgwGxZE5nZgvITlbXI2OWyICkopEq78B6g1a2TdkHunidWtU+Uj7zZ
fPp5RbrxO7CktQexJRoukfP4aFunzNSaUT6YoWp7kC+jEtKrgksktvEgYoX7w/uq
uXhopnvCpGnvcOU/+YHuhfsGVq8YT+S7KtCHKGRndYnwuavS02DarP5aqTcp6cFM
YMDC6tM4zXSbWsBIxKeNeTmhn9MfFl2WkqP0NbvVogAG0ezogIGkZSKEHttjQh+s
HsCBK89W1Yndwe1jN0riaEjogdo7jcQ6U2AeNRJuyOrtRh/oeku4cHJBCZUJa0MN
ButxTyZzUBSMoc6jv66xMY162BgqUTk7u/eQzaB0JyImiRY6ukWBGoKmDieg0CTY
g3wqEu/XGfk29SJoWrQXWOSGU8aDbwacDrLuzij4uzEtsIkSWoQwHSCybSHpZF1O
LsnwR3QqAl82sjVvZ9d4zQ89n0tO308ZVGvGzzEFsEhBdU/JckhxNp5FkunOfQdY
TlYejZm4CVZVEGX+tPgwYoBvM/Fy4TKV+cqSFq/GbhdK4OiofRCR3U6b981/Icj/
29Ya8mKLd3SOtTL+gVBCyXKPdxIBhU9yUXiLs/7X7WI72Otjp/WG/4CCW8wg2g7J
+obCYgSoFV3oQUsLFbMi88jzA0ijGf8JXCRZmyRE6GR7s3fSB5gB3kSEX9McY/zQ
ePkgZ6UjpP4yjmz8Tuv2xjc/58AkRKJzVGMCgYUgvbvx3I8hYgN3q5OKlTr4PQyv
Y4UHt7rc7jja9MrRedwo8jxnAH1e9hy8/JK9hCYVKh1Izn6y1qmWfk/R+fTkaJcC
9DhhxP95vdLBHzlII7mmr5KEOeHMUuvVHGuzWJBWCEpOF1tH/y4i7kFOueFRFUH7
AxjQzce/8L9Og5M9VbmQRnb0/Z0FEoLPoMq1PAm3ob+9ZUD6yJ2tk8G6c5fmgxqO
Ts31XlTWQXLntvedpyPtV1L2Hxd8ucWjrJUinNQ8jS2upexUqPXwT9Hx3XaYyB4s
J9rTbmWPzb3v+gZthiIZm9rGUVWxiNEZrdCkf55CkcLsvX7q9MHX9VbWSuBkNszo
lAEV7Uy7050FO0bcnVleVyJZd7NZ9d2y6qtC/pU8dxWp0A3LpH2in4Vk/Qj2Jud8
UlcSaSrgpmk+REMMNY6e0W5rmMN6q1N/6ULaBnUbIrCNZQkEH9L0rfXr7ZFso2Hj
98pt4BzAW/0/cPsWCbEgDvLNk/bRiuo4rPthPdGDnw39NjTJStFkK2QD4Rn0M9Oe
4/hm7W0/IWxoZd9D6akHoRgfXH43k3+R8+D8oEvL4deAAsxnncn0qe6jCPCB3qC1
bg31NEWPTGYRUq3Eeahmp7KLjOpt+YNEvlh4rWD2Z45DkKZE7s/9uJcc6Q5MjNu2
NZMqSS4mwzkAK2aEO9yFlUFurQy1RtZpQ3LIsWC+fUPLM1Mlb6oRskdzYSukw70R
efyJCP3ck7N4OdkjmwMuSdMIprqkA+qV93amo/Xnh8BUNffy1gIwctoBdioLlyiV
pwHZvX8GmgNwMN/6hPUMyyhOADqSPUIPynov5sCWHONz4E8yE3cYsL+r2PIKRmua
5sUWNVE8mWE1mUh5RMTc/z34B0vp9bm2+klR3NiMvf0P31wFF8pTUEC5SG0f2C6Y
ZJRGKlqs0tl8SPKeUgXXy9MQbH5V/KN20IZjaF+fiWYfstMd9osEcnQ3rmI4gcgR
TEz62qGnOGUReYCOf21OWLAUOjm64vKOUF3ERZtje6U0NVJw0DsMNXEqJ2v8i+Oh
1yrQQOSBBJkW71HyAgICj8kaE3ZZvfec6dp24ITYhkpzUkmY9GFknwJNhyGvxHdW
xy5KcI/7mU5XD7XN+nohuqPH5AlTAD2Fmx2lE5AKcSQg7j0kDFAwCmk/alRFj4dE
wRA1bqZzr2/0dKtA2HuV+b6aeMrVKG7yeGwjaMv/QHnLc5WBhVUAx7ogWpS0XnoH
rHeRVXmozmScQ2kdFvI/ez8zfXZNg2igsZY96UcPYOq9OwYWYfxCDjzPhKXgXDel
WxczHW8MZt15jdbTDm4QdfKpjwKoKw0RCLS4daZ+LOeBxtIYbVDa6FRvNl6cRQYS
CmgpSjIiYRWjcezt/i5CCPUerV4vq76uWOw+/yc1qFgfzSZ9i8gUouLqq2os1F8+
IASosL83Thw+Fn0dxTlYJosxtfMAdMEO43/Y/MuivOWndBjJMMwpbHjGvfCmlppM
sGR8mDaeUX6T7tArnDI1T+mFz6yKAV4QSWZLKbhmiskL7Tsq1PEk6J5xx6zx8AHH
Lr1nxxnptGrY/dw2007ler7gBDXcHjiP76IiszHSF7+hClr2jDFSWICNUc72qk8v
Hm/PRHWoLkzE/1IpW6zZwlUdMdv+cqJIb6I7A6EnZtJ1+7y6Tn8gvXA44uJS9s5n
2oDFDbDlgjRXEwd+eyXGCiaM8SY8Nwh8vKkH87BAdTfJwq5aJPcc7BJHPD7mR9vy
6wfPPIThxLcs16njqJyR+XoUsGKgjIRmnL/Ok0rdu8SDPo8/F1wI0bmFmJFrTSgW
5Hvj0Gp/UYAxziAz2F6sYneR7eDeZoe0kmLxTjBQYH3KwiE9zfLRDWnYio89qC7G
l/RH+dyfZBaPhkKY9EHzzajwcx6QPDe3wLIqJcsm0MYyZ0ioCeUbT8zHkdiYD9ru
wvLsBT408GSzJg8Oezm+CePMWQJ/rSd2wzGM7Oo7hQ0QkT6dCur29LTK7sPjZXRY
dkEC+nbmas/w/mvX7vc3VOYzTNbrHq225RRKjNxopqBYdmdBUXya4R31l9j/qAbU
29iojRJFg3SDKT/QLm7cF+SWo8IR92pY0WVGGd6xZDX9/rvfSKSWCzC7OGumOW6V
vAV35anrFIv4Mc/k+7bgy+CR1lssEOCgiYqu5Xeb6HFddORto6spu0o4ve1Y5deP
a97udtZix+CT466Re24lQ4qWwxGwC8KZkxAnmuZydMroh7AEuYptwKHVuq/SrDVg
2Oy4inUW81UDpLuexmrPxj3blacrlpCsv8kJSzr0cUNj7jLUKzz/V86FAqE+GaSG
SJSZokjo//tGh7j74mA7QnamuzxY/sK0jy2Xw6jE0Z8WfvZKwl1XlkT8OOIHrgwY
K1HTW6EFdHOqyHp+DC6GwRelZJTbmBtAXyEpY2kbRBWCRfqAnRismpk725N20rdj
ka6EVVeP/W20TbDDnmR4786D3SFdKeMAn4Q+EA+LSVpqcZX/Ez4A3Nw06gBPkNZ7
2leUBllmvtg5PBwLZDkhbqQ4rmKJCWhWjlNt9LXVEA3FxnPKNKUShzmzhys1Pp7A
HNDaQx4PKBMDSXAogaUFv3n2H2FNsTBLty5++GONhseYUXSnTarpFs8PlND4Bvqp
NeLol4s13ecEV/AyOEZ2UvipwvJkTyK1fyxFlAZ7LNUxjFmRc7QKiDlrnDFWyJPU
vcr1NvIkKQhsP6xDdO2KLhst8pqIp4bufx7gDWeDKOa6RZp/7jx5GaaXUhU9+P7u
fDdaRYYqMwz+mzuxq4I56+/slzVpChJ4GpU05geD1epCeSW1a/EJrHVSBcMRCZlM
K3f7vyAsaFq2kxArLKfZ9HPl30dV5ASm54vTBTdMAyrGceZuTaFoPmeHw/F+QfA7
behIhHUS2067Cg+4VjwUTt15yflzTZ8cfI9B7QTO3LVgYrimGt0WhTx13IwZN3c3
oWA2x16QWrfPwmY0qlhx1FYSPSs5jlUV11QmmZoEfnukFCaDL/msb0iFxXd8mZFd
tsQp85lhG7D6lwnNQ8+eM33wy6XNgI9U82uR10Fj2gmwjch4L5+znJu5JBOwDV6m
sbjyckcwvoDCQUwo82Z+8jqHZsI1a9xD9mBkfo7rT8DIqxy9D1AOiscOHOMKhwON
qEAPZLJ2rdGJ1BBwKci+yyLNHxg/DnJS1IVxn48Eq857qwpxRKeUG38PvyNe87ZP
Kf3WQGCYMEJsxHVE3AfGuQ7I30K7TMx0l2b1DwWK18cMraw3QxHQ/i4TBcExozjH
l/A0d9z/dx+WK+JUDdFPZhDNwQz/qBSoWXz5806dl7f9zZSS6mJeOFRXYcmoBzW3
7L3DwWUVInB1wTsVsLkL37zsi7SUFT+1ap69ESqaOdEuS4WhmEJKlo035d3PRtkl
Xc/ghKMMkELonxYYlUmH0F3z2oZdLfmLdD7tuiUBYEpEk5ALx3Xw3iKXCDn9SprG
Mf23BzHFNgpJO476Lsv7LlzZVenEpJfeAewHsxmayLw6lTgupLtAaqGZBlWuImTu
lrskNF1JxPThYPyFXlP7PaMD4xb0rELHNeo1abBlIB2uxZoypwwmEAVKMvvyiSOX
Xw2orUV6XvpCPdjLeoeTCFH5NmHQs0/UtZxb2KtpULkNaBr23P7ZwxmKaMWvXR/C
Sh+jF6ctGzvNoA0IsAnssLjnWUlZZkUZ+8+l1ttRBjFuaAg58HcqWk/4r/DFjIj0
5x5g7WU6Ofwdfn7lL9SdjHZbzgi+VfJWJGWupkD+7VJyNGj4wWrk2/5U5jv/CgY5
hxKctFOHlI3pn7dY+jd9HaIaWC9JO6dWgP9PvBmGbrYthYkzUxEQe7m3PHpgyRTv
bxYdZH8gFl69koWTqavoJlR9RhU78QvYZaWOdWHnT2mS6xjyxiFcanZxsR31dwpJ
GfCdRWN4dyeFoTVs3UN0b/Vov5D9eK5bDJ7l+zqEhackyZwrjnxevTWWtqGWElc8
zkZSSWLpylWEh7CjS5zpaA3dN99j/ePDadGCbUuJzIgHqniSY3bq+OrwshDta+vu
XVNyBMZWdiMcrF/bD+9ZX+FksgAO2XCflYq467hSDzaneQQdTASq9tf0/GhS/TBz
ZM1Shd4jUevmstoQ10jHmrbrk0OjECzzyF0c2vOEdB+C1N6ktXFhinhtqWTiOm5h
uKfmSnOCaAo2JEW1SxnxQZTsxiXurThLXz1cvGUy0pDs3TvRGciYMJa2Tg7ldZ2g
uoX+sU/NZXMwC4Kh4I8yycCP+YNnTIo9rwDGIO6QPk14XcQwMKBdBVShNxrwIvtv
kpemC6LSUbHmHD9zLR3bMS6mbNSfEDURK0hnyo8CNMCejFH8MwIvc6CFTpd9jpyQ
DmRlMVH5KacIG21ZH+sXFlGK9H044Po0zd5151gV0M8pT0NIP4Ojo5Atxsyro3JJ
aPXLjiVX/3YP99uMSql+1yHOKqXtQt0qlcUoK0uV3kRXx2BrxlwO+GBb9CeWn6kc
eme5z3oMrSzbnoLTm/U30o77QIgj2xIlUaAWiLdEz67zuRlAksJyWOmecBCDxz2W
z46w7XKR7t9w6lcymEJRsPOlAPYzspsf6M7KnlzeV4g6BNPZpqbWUnjoxugZ8dFd
63kZp7mQpvKuzltxuIGuNG+Xr7TXx30Ksc6oweAxXmBAwX/fb6Euqc7Ytw8RsdaU
dadxpNPsYkcqvOGEMzoNDCoCsLCf3yXQeofZ+SA4QAlosJBpnjTlCJqXUacU/Sdk
o4Plkz2m6ALfCMrA18GqZKWvhuqp2rY94TNQQpJCMlA//6YxnfEIHXyR7h8ewi2W
voo3778qn5gptGWMJFyOzsZzIu5kAYowrXDQdYrhMgy+nFstXkwt/l4+gip5VJix
VdzJQV8pI+NqG2l4AyJO8aIe2APNfgwuL2L+YAPjrcNmWTfJRKRWaJKMNTlAxOoP
b/kKcJE7zCyAcA9tyJlqqHIjnmgj4INda7Abiv1jw1P8wdA23BCZtcpoKF4auDdI
fvtbUtjTCzEwN+mRa+N9lUN2Ja+FBXOCh7FmOuxcvnjnzNeEi3RdLLfLqFlvlYJQ
Mp1k16eOskHAMF4ZaZZwjbx5fQMr8m8dBjeZ090NpCShfKaU8cRc1U5abSOE1wEa
TLME8B/1D+tBLz1fctBydcSsduootxjlfqr3TOX0M05v8dVB6oGPSwKadC8l2cIx
gyh1BTSQVckujOUjnLF+w7n1XybS4/cjal+afYoOtxWWZTr+04XoK/UapL3XU+0T
sgK+F5Z1EmWyQDpb3baeQAn88u4rQzxXFOwJtKmFZUcQqlwyNLpCVJChc1ZCyVf1
dJo5iNMzUeksTQ5HhO49HfukNJxS2ktEe9LEj2cpZH0X8xS8GmVyWJ6WE+aQk1o8
JMfJc5ytj8qGYm5evgZLyRb/cyoldtYtGg+NwKVyoOxyGra4O82m5BvsWTJqVn+j
oRYo1FH8w9HOLZWC1dr8gY53Zi20Vna5CSo54BKOLbqRwvic5EEWC293/4jxsERw
f1fvtPnr0CBmywqkzLgkINzsv2gyJYl/eYBpooZrZQ5HbUu5HWYAsAZfOt8W1bP8
kg4yCmVb0ZtF9u4jOnvSfEu6ikiTFoNdhRHTvy27VzpVPM8FCYqsgT1qYORZ+ZK8
Q/pgdfUNB7TtjzlTpRxUoZHMGO8RppgWEJzgX1RI+9Cqxi6Hd4FIBpQN0k2j6qFx
G7/4F/d0CcwSle0bqO8nZvjb2eZQxd1WJ8+kobQVuKSmt0DpRLa6t4UmUS3p6GsY
g6gBSxQXWjNLy07rZ2IRxh4sEUbTKmx7DN7Rm0pPfWqpjWYZfymheYrQOYB0b/5K
KrmxZGFgmVj1sG00oFZuLwhIKO3e3/mk/YLO8PBYX7d3GpoYN7gLwW5R7XxXaIIk
edq5S8aJeNNVz+FNUi4d2Vu6j8vcNnUwozCM3GJLlhFyrx1eXE3sniYxNoRsUsBu
X2M9sjckVJcmAzSPZD9SW3D5vl9ICaKAl2bMZqQ17k5hMWvcNGD1o7+OJLA4B+oz
kZ+9Q3mOZZsA45FAiiQgF+eARVCk/AjuxWEkfqqGtQl92kEPoJjBpCHDklm5Whwy
v6Stf4Zq2jsgdQWy+hP5riBRLOm0oVRyAM878OCEinRcPBsy/OohgXvNArrAbV+C
vADNRlr2ki2sx/I+zsbbQIyBI/IF3MZVECyyWfvG35yjoixwWlei6JKhls0YN605
UZKuQ0OU0Vp1XlkFj8V/Rc5CsVvjPNldvvTGHukUL/Xxse0Z0SkUC5C95qcZRFhO
JmHjs11X5YPzeYzyTcdqi9rcgJ41IQvrHV5l9Y0Pz6JYWaeVV8zDcYXHd7r9U4Nx
YDhx/shl+X9GSKV3KzxpPrb3H2xD83GUpJ7Wbuxm6GrtOx3SY91hkIabIvrcpQam
DFmj+qxDmp0OodncMU3yFfHvGF/YdsUXYmqWnphpZCWhA5MgdG4a4SZ7YG+yozFW
mcNY1TTiPED2h2SGFQiP2oVcuKSQcIDv2sbbk3HLffVBJDSc0XPEfzCseHydPIO9
86v5hi3tSCTXQQBJdVKxJuIiKFzmUUVgh+IHzShpY/cu8rO793zMx4Sz6spKDP83
LsT5L9hJmMmYA8u6+voOq8padKQjij5gpwZZhLhqpfbVoKbSx0m3ASXAPZrqsoM9
AudMIz+2beP0OMOEGltUns9+LOJvlFgT6gVCihPQSOP506wdodTUNCoqMO9vz1A+
CgkguXcBvhPXupmAk6DRFl5rDqHAo8W4WGFD+kKLB7ELA3XrKg2mFIp3GD7DRFWp
GhlVinlyuNwqyRDwkW3kv7KM0Ics7Xx8WSayBZAy1R3YE92nKnY31kchr/HBDjtx
FajslejYxcnaVhNhGXEe1Ejtl90FFBzeDNFeo4VT4oI=
`protect END_PROTECTED
