`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QHqxzlIuc2vbdHTHU+o0XLt68fAMuHMp+ryAZLmYWHiQSqm39P66cNjXdlPQ5Vf2
J6zM7heq3Mt5F5CUaX5YbFTq38CBgtl7rNF6mR+fttw8atwu+S1YIPe+d72Q5uDj
Jf9eY/NGskhJArW7c3/vOUpzfJdTEw6Ecgu6rlTHPCbDH5Fv6LXHaF2aL8evtFF+
dBlSN02sB4ADgtQkE4GUKlYQkgNRXejBxWCrrNOnPTsbDQoTZGQv0AcCUJZPWfUg
EmeQ5HCuT0Iu7VeiVQaDAJtvHN9uOKObnfQPtI6JRDF/jrBkqKikIipOBUCiw5fC
OxKbG9tqNZPCtP3tj/hfv5yLXr6xLLWT/CMBrlpj5Ttr4BWBBUUk5YPHt/F+on0h
VBPGsE+WKSacNVHrhCDMrjqEYq9zHd/DT1Oe3tt2ceCOMMNxDivRLPIi3Pp8fZuh
zCbphVYYY/GRa4NEIMwsUUSzPjuNXERcnaTk9XJOwcgENGrmrKxVnSieIphhTlr1
1dzFIGLSrewoJiZTVXUeN6UZKDhifzm0URtf0tpQBrR6SPemb6n2+13m3Id9IpUr
hhIHXV7hXKjySsVMAiTVqQ==
`protect END_PROTECTED
