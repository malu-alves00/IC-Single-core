`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HeHTHPswjHE3fHStDD5lqqasm9lIDUIypJYf9QCRh3Ibcy/cAF6QjT/QFoO/6QiN
GRsMYLwkK7635VthyUNO5pbp2OGPggKD94fJ4tS+9010z1Tm0wv5THneug4rmNkE
QNmCVjNnYWuueOifSLOIug8lazrKDOpREmnpFz78iPW7PtDNwVB7PD8Oiw5CzqG1
FPXjGNp1W8xxV+d0K40fSU4vjK0N2ibEhSTbBrlmYgRBzKHPWiL6zkySguB+DAP/
lti2RRXqQK7Xott42NkXBZT+dM+ahTyQmU4QhH7UIPAEFLW4FPPStrFK9iY5X96T
0QXrWBmiZNR6/734VMj6abUWt7QSUo+M7R5oLlq0Ns+BYmz86IPIu1LGWloGbhae
wABD2KOUgOjy/Tbg/6FZnBQs8/ZnutokMcbysMed/MFj11jFlq6q5RFVGakbAeLc
vXEEc4p5uwmcn0gNxu/86Z/NeHGYVU6DWnIDqbJOQxYqaB7oEqm1Lp1+59cWmesm
YQg7ajGO3/rtwArXvHIUEsdWb6UB9HtsN4QFeCcjQfyJFpzKwNWIUFzCH8F+vACs
0vEm8ypv+b9UVrcNQAG/w5umIbM6lhDGBCkK6gCZiqYXNxP5PkkRBI3/eDyrtjDI
8By9ndiMhP9fohYylEXaoDfBXNE+wV13tKpmOq26QaIJTfJIP1Vn420wO/dS8bOV
9E9LeNr2+4AtgklQIzo0AkjlEOnsBB1B0ZSIHVrsMcZLs5a9ibZT7UV6IJouZg/B
bT7pnc26VCKAUT4qSmM08MHYkDYQ3d5AeSB3QD98NTeLpvHowpatfIg//hzPZa8+
4hjkh+M9V0M1d2E1expDuy+IOo1oeFWneYS2FFrNoEhNmYaU7vomi7Pw7kUa+9p/
CDfm6ZU+wbvAA5h65Y6067rvPHN0jlQYyvXNbjpOfgKpmCSUiMncKMZVVJuflawg
`protect END_PROTECTED
