`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RA+kB3R4RnKtI8w+O4DW8eL9iZ6agSyyT0DoRDVpGQk3Y+Bs8/R8aBVSs6v4mM9C
IpZ1Ohrxe2RrODxHFIpfUbSjcwB/JT0JvbMLlzMTdaXX0bI3vLApN/fVvqgefoBO
sb+K/s/thaSvlBzDu0w1XzDR+p3Vhltdp0SCNTcrVJN4Hv4Ki7wHutITbe+RLVof
XtOjhxw5petw9KvkOcdEBQj6v6yRN1LE0RI1OgpGWYOpq6GPUnlc4wPvkXWgIOfE
dATwcgPX6eVPt243YrBrguJHEYmoxZtGDNg4drEpkoPfIpSpzgyEVQpDMV3iMI2V
A/QiPcRTAUv+WV2VVydxhgtojkNLo8HcLuH5P/hgPF5gG1tqGtAvpWfj3hvvIIBX
pYz5HQ1tV3bKv8gMFz7fyoptucrf37+EQ1HfVqGcP2RzEliQVuachMIdJFhwFbT6
peb0yUAQQGYcQOqxj6gloNBfxDRsJeUSHzVSC9QFmZXlQ1UoRYy5NGdEw6NHrG37
wjzsH4Rn+wqQ+Ckw0ymKU2o1Y2LiuzGAM+VINsQHR9Dhzkg53ecscxwXDfvnEPFT
ezhZLxBMQC/KZfm8OYOd9NEhpFuJrL0y2WS2mzgxY6zZ+jtFac9mva+QK5L2mZJF
R3+B7O8W9853vz8clm4v13SNfAIY2zMFp0YMZMUyG920ZzhXpzfNbs8lRWb2C2RB
Avqx9FAsep732SHacfJdHuVZo4Af/IoCaHmxSTMOWba/CAS8wYwm2I9XxpjEwyBx
SG/8a+Q+AO0Sno6PQnKkADSgU8NrjJWwFBGE86aA1rmFtBGRPV6DkrC+8D/+Py27
zXwuqxEbBfJA4C8zRtnVg/DzPjT+9muApYMfdBMMbci3qSdrC5IwEVCkdqTOMZ34
1jkL0RJHeqMhhcihOphMwY+TIVr+vHSTgQA2eDLF7TqUVy6Em/ewUL8u4EhhOJ5d
/AdDWgKG6rhskHHRQ+++uyI0/l6CX2cTu+pshjxHCtUy4XYmWLoMLr3tHVXePaqA
xrxQDR/IpAsYacB5j7/KAnwgFIdoJOYpBvvoyTu3KAzrLnDbhsXIdUo73+pFIO8p
z2Ly19X7v6KKl9+7x0AzhDZFYPDEBzdl/3HgV1r61K+HiQHuP5pQNlDzSEWYTTGy
mVoAgkCnaGOBy44lXVP1hEPmDl2lq4ztNmA4Iewp5eep96jSdxf0lm5HQD/xY85P
Uk50W4nPOrUkfas3DSwJqyexDFB1EEzpIQYJiP8RrPBKD+7v1rsW3KFW+NeElbFi
ERWh0Iyxjg5ENKp3K0OCFEWmyDyw+SgihIHCrI0Hc7mzAq4qq1jxX7UdPP7xICHn
KUEzKlEGutswf2k6+r1cu0EPeMptDq3SC9ZpvdvN2pK1XVtFCwa25C87lsMtbNNu
Mfrha543yRyJXloHsNsyce6dYs/g3+BEljUjipSBsYxpGD8Ja04NwpHU9KoJnuHX
U4jYZM996NklPjT/ft9CzIW5y96W/IZ79vsqEB95gLYj+TFqm/M4Lzp+NTgk/2nz
9W/o2oy3hskP73bJb8Ubs8XbeZN0qZYHz4Al/TJEcqQb9UK1ik/+v7yQPRv78+G6
8Oyjp3qRHddafSHwX/De0gnsPnYAyYiLrzIXyg/d5SvULczj4sXqzBtnBO8/41nG
eAQLwYJNXdvGh84Asy3DCLNj2oiQn55+ht3gv7joROd8ghEl21fXOrduYuMBh0wA
6FtG+fo++ceo99GLAW/SvNZJS9HSMgegJI+8o4LFc8tS/18JZcmoXLdIPekzrnkc
U0TiJtDL+7sBLHyFcNM7KfpLgfu5F40rSAiAl5y6MkM2lbFjLPJ4QtR5ARWbGAZz
9KRkeWYwIrEqA8FzY1KeaVfAFk9EGnDxYP++x8dWEbqF5em+nvmO/Zbm0cgxt6Ko
/tX9lEixc6aM9xPbUBM+obA/F6+N5PD7NkNNlOHJtSqcseBspvJPK5lkbxU4DEOi
GoLOKfh8SSxSVASnQHQMoZ0YTL0VdakgGeFmjMmYCrKx0iib7s30xGYykAoXwD6A
veU6Gpyh3TGnxVjFM/WKQZHXEvidgXkNv4OtyjMrWHVcoCeOAaqMYVEEUX0EJBfF
Gqm3V7WFZG5BRlRn+5T//EFRyzKE2lcAA+dx67opl8cUzcxysRoqzlp6KQjzw5y3
z9J6bjQPDsvDDP+AjIoi5Ysc00sYgyC+ygEOkSP7BRZFsT3aK7ekJ679esbNbueP
3TGIT0Z4GAyrpm+Je6qPaNtG16jwWSoS7lXzjlW7DJNFSfh0f/sW7vc1CTw1t4Z+
2yoUNl697HocE0gZG0Ak4EDDJOpBirzhrhfMpqdygq57hfn91EsdJ7l0RPZx7jgB
f7+ZD6pEtcHcR+tG/UbUpEoTXvlkmkc0ERD2sfD1CIdOMtf40Ht81FJPpH/4RDun
wxVooRWcDb/b4f64ADW1hGPGG6Nqw2gM+kAYXGqDb6gPWS3xBKMqm/OBFLeDWBPN
I6pgeGqGODwCI2MVyPz8McP9tLKOAsi5E7BXBAUGYkSCWG0SUCis5d3bnYi0rQPi
89uURkYcEmX8fKu17so8Kc5dDv5f1CzE5pGDMvFC2bAhn8NNcKVaszSApFDpbsfw
EcpJHgQDNOTVdSuDTaYi5fCyevH2apJfUMoNTS1zDPp2rOiDGXNMhU4fRpv3dIwN
`protect END_PROTECTED
