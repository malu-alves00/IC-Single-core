`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
elZJspOKHG1iTR9eXKDxZ1enWYQnmYdpzdH5bBxEiQQegnfwGxcQyk2i7Iy48exC
Or0QAlpaS1kIOTxmaDI+FPVdZAbOCUMS2sOIQy97uyj+MyMQsk2nRkXwRhut37cc
AEScilxcMOzmop5wrfCurz+gWfgXkmlKRCc0BoaImHkteUgn/2dWpmlkOrP3y3kt
s4VQgF6lAdP1t+DA6ZkY+lazUnVFNLnUio1ZbVqcfarl8I/jhfOReYeYIjny22vh
XDOXKxHNDytUnBnZ7atFGMHzDNPOPCL5hzpotkh0C++ZvxnjnxUhtrWbn+jytD0Q
ee52pHaoeJTERcsq7IF7n+UCMTSwPNnDxmwExr8E+DI6GUQwqYHwTQzSb9aItpda
U5+6cXVI7PXddJ4qU37Y2pfb4tQ+8N+AJ79PVfUtDawZODAG4xgpZXvdPBkCSmoT
09T9VcZIgTyO51Fl5MemXSU6aOzPXtR426FZrEw2wDh3FayjJFMTJDbLvj63umip
MhqX7VB+4WmxkQl5v4XFJZUA0/2Gr8/E4evh1wAqpkfh7Y7NPY20ws7LILvkjUgR
ZVt5ECWBNVkcYnd+jWaUoVuvzjU/39PxL5ZGYF8QZ034hCwvSYD2dL5XPLSdW6jk
Ua5oREO+otfCn51CQMtaxZA+2u99zaAC/3mjZaEm66HR99LILoCkk/PrPF44y1Px
SGN4W54ssPzrkvDFFWelyU0KTX/me4Z2v8gHw7x2zgsxHcEVrG67+FrMt4HUgexY
ukn0k325wf78ZbFoQLLeCw4pf/ztJA/40DHChAiCKD9wimoopb/q/HuRQAcjDrGU
NQq9H1QQZwkx2kGc9Q9oboscP4njaj2X0JAoCZ0PLQL5nR4/kTHJNEerGB0s4Wt9
o9QgvFP80qDL4sKk7D/DDQ9teNT5UiyD1PYKHYNTKcZf+x2R3e9OzSrA0/dgsjHb
KykImxwG9J3t452cQqpZ+9/awkTQLXCyyl2Qyunhvn8iQEzENcHsYpmT2ZToLa4D
5OR8N8MOSgk/uK9L3s/FlZbTAip3GUFFp6x2SwJ0BQ7q3shO8SZ89W19QUSrziYO
Cmf98lbgsLkerw6FzUX6lI/7XBdXzw2fa4g5vi3RNiHHdisDzcqM/Px1MYjDBc1B
Yu16go3Y/IsbwptJUu8eyYbUcFPJ0wNXdZ1eri5/Di7shjwY73+15UQNgiIISURo
1C3H2kASRjh2T8iqNI1wjWMTedkBYvS/FgKHyfiILQwEOVmyJWQHOxbBGC+JT3Hd
KxBuZ0qgnBZ5BsAnXlcIWAfQsZWuvOyRUnISFB/pBbcQJkLJG+YQ2k9dFh3fIyAR
IJxZ6HnUJd/vdXbc+tp0Uekuc7ddA3CR0VQFQVf33os5zR6XQ1GZhyw+78Cnvchg
baTam4IOoTtaDa43qbvUVwkz6yjLSH52x6GfSE4e0xMvn+uHQxEL4xdFd8enSOoF
fx72q3KbyolAvgFCiRJCACQ/DFpS/gqRd+zDCXcyKFncZeYzX6PCSAivJ7qZF+TW
iZmGYcLOCp+HMLznUa27DuGYC35PzF7koaqZmQ9/gjVQeyojuyhzYtNSLX1Nu6xS
uxXpPJr2CKLTieygK4tQl3LZcjXFNX4kAcKVKzMiJxH9NgFtJZLdgQ9LBV/LfsnZ
HbdnJOFfSynnHGMC/PEUZ6ZsT87qWtANzUGO1B2AO3pZr6cT9M61WjiAzZmXRPFl
1PrnNIlluyepATNjvHFlB1eFJ6+VJH8z1rSAwI/IZXDZx4w1uipy5Uc3K6PgMKlX
7iwhuNPzEoAb5uLELQLw6PHXY7BfzfkaD1IDndXty+bsPmcaqmAjnYL+1sOEvjlx
0x9DQHQzq/W90pgkVrudZuQBcbzUxZI/EeXNR+Z2QI12ysGKuIUv3p8K0vjvMl+h
mt+9kfObvrzIHpJ23ypBbU0LTce9B3EgY6PKAYZellxA7JH/Y6bH8L+f/ORbXLnW
xGDoWeWqSLTQ6fbf71md4DxuFalj79vx+Wxi2vXgmNbb8jfE/R+eJacGLLhnNhW8
akCSanSQ4MenZyvRACE2nuClSUre2FLa7P7GnX3c9O1SdoGSnj7zoGZpQj6BMQtM
SlsLa4d8hl5MJpGrn1nRpSuwRNfjiH+NvuO2UQRSPfye5K6/S7i0kpSZBheRvRMD
ifr8FKHGGnckq3G5vZGmURvn+xNSVK9+9m/KQ1LejnYALhgUEW7TjvzpJpcTrRnr
70mK7KU5HEqUwCmNK8SlTS2ivncq69b8c0eQ6Bm1IQhrUfSP4h+cW7JbEiDx9AGx
aV3fQHhYSjvzOdVn935aHWUimUrIJ+Os4LlLb7GCMmq+xK2tzAx6CygrSTwACa+8
tL4TbUbUTj0yH03hToTrM2edZII9UqOwgtjSUBk9kMVm0ZotmHc6pdQlB6J45iik
xMD7YY9WiOzwypHPVwykw30D1qU5QWfawm1VeulD+xTSHHykiILp0RX4F9ENziJA
4qx34kLdBJZ4whjnuRYDb/Fn4hQe+nmrkcIaqyp9a6FnOB7NWrdc66yzuXarElyQ
PZPzpZQpu+Izf83CR568N1uLALY/6/iPvH41zuObo6zegQx9rMFSX0P8GoAEk/7D
6s6WKkP0Cnzu5UQrzHgztmI28EZpObSKDYgxSxxvg4uabjJiJlE1sHTMWv5lkrpW
Todf154N1eCG2h314taL65UghFIrtwAfFhY5QAi0hZiPnRcb1Y7D6Buo6Oc7OPyT
epacOuxHaMAb8e3yTBymBLqvjCkCz0BoMt1KY7VWHGMq+VdH2OEsKij/mYsYmPQN
aROtlbPte0CaxWPPs/pke3uj0VbExMgDp59e3Fy0PwZ8YhC9Xoy5VUUI2224bAFo
7brs+dKRNjoEyZenNJelq0naZgKJA+SpBm1RVyUzTsBdOLprOWs0Gq7pd6Mv56uj
epX5M3tSUbiUrqBIpVGkXowgA6eTQfqfjagBC2J7qeM7na/hAS4e5HnYWHrTkOIH
QDuCiY3g9NSUgTTBsmbh462e34N/pxKq6Zq6kSo4IBYViT20tiZ9mXdPFBUI1YQ2
iVitARsoQiln0YbugFSQ1z5AsQx0vvr3EAknjPHQxCNv28mskqPyi9sxrzdUH0SO
uGxtN2XYNwXn5dOrQfB4axDNgdY+U58uSefjcPGp/EOjCT6qxeq8pZeWVtbBSLG1
R5GF+eb62T1meKwH5pLsH/VskL3jMqYIVBKOC9AQQeSOhVtYsWbuT2LdWQIFDUr7
hczXuDeNbg/j1Xmfu9zAsxurjGgUiTuw5sN8uJ4AVJ7JtOQyknMr2vmGnXhCR2cu
bEfGeg/cxJmndg3g+gMN8rLDhe2KQGN3weuw9bW60dTw0KAD09iTeR/yfpgd8d/U
3sUAqeaTpvThjiwk5AbD++BLeia76xZs8mtpFPJ9WM6qIbyd8din35qYJAJ3uY9k
crmDTgf+O5wSZ61d5kevAm1fSCMfnYPhhL/KMvhx0Xhl9ytVw7UAZXAM6Zde3kEB
xWPREvm6jOkXDHleMuoQ3nAycX+3Vn9lPFAUTk8/35C4rhAHvTsLbcjO48T2ldsL
sx5puVPwu+cLFXkW34vmiJrDboVf4D8PHod+/M7QRZA+V/N087XQZ51VqduY6tbg
WG1fwZSOr2FZRPcSe2TBDSZ24zMIZy4T2b6gnANdeJl+wTVk5n1BVT3vfTqvf6nR
oL2GxZ8o6Jwkvdb8PwFD1A/P0WdBlfUMKKh7VmKYgwrbrTqIHhmH+ypVs/g2PL4f
XPTGUa0g3GMzVSuou1feZY5O6MFU2hceAXfjESc2BxjkZ+b+MxGzApiRoVWGfio6
/IwlIvgenVzb1xLCdr0ybkb9SXbu1ondPzhrXMFx8JOBvrzyUEJedDD3o37coLl9
qNVzfUephpGbYAWks6V8cL2TFjD2Y9ju0Tf/v018kzY6nPVr+YdVy1lJfZwCDlYD
WNmMR/iUqg+1/T8Dsv1b1A+YhyVNl5y4Tvv9mb6TgdEhmVUPMOJhodIamzBGKO35
72znG8Uy1DW/1SQtU4oTBIvowSb2xMfehtM7ze/H4nAZoMF4kHrJDa4asw/eIlTH
goyoubfGIExjcZYb9UfNm0KR0ddjADEqWzsNo+m9f3ftrYA3MYo5mqeay6+xOFgQ
6irsT0WfaSg7R6m08e5Jb3qwyzWI2uO/N44gnNMh+Alht+p2cfK4bH+iSvLoPlSO
TGJX8sTM0+y7HUeQfkzCfxIw+jraGTk49aBjvj9TddvIrlkL8rsUCgYAbbcWcKZI
dOWrz2prIa1rcTUmpW67nLp49GLqE+5ka/V2a4KVuP8x09Ka68r07naSrMuxj5NG
DhFOPkGBedNEzq/q92Q4hgbbfGV9HrdGUFE/PTC+Qx2d86PHix+7gHuuAomtCh8C
E50UdI+hvVoPROy3Dep7s5Bzn1+MfSNnHb6+xdrDHo3HR9XidyyL9O71zxWlQ16V
gR+YiAKV2F0VkrfX2Ft6TYp7WSWO6omTBfy5If35N7sDhT5IAyovvnFyXFj7828y
mLtkPyQdKY8vEantkZBJv1c30YqMRsEXb6MpxZqMfbUJu5NvpzkkAhCWI9i5I97o
EFbX2/MORfQC0wn4pDmuwAC94YPFhFSGPmrucTdwYDPyMzgNDKsGIvvDtyqK0736
tEx3+HAB0LG2DZqavf/2LlpZEYT4wmMm1gZaS0BibBQ1x/8IvU2IyHATVkGWzQFl
bYftFG5VGmHmRm3FNapeG1A30w6gmMD9tV3I5f60d/9fuDjyYH5EBoGbOjYZyuVC
24NiFc/wdBv28imlKUMuXPn04E1rFF1ntOQWMw766QfnrQXpeu1bW7eAkedcLPvn
ONB1rQ46Qjct/h2TwWaA4pEg7nTaD2dNinBfgQxjFjEERs6DhF1Ap+fCujKKJpY/
0hZP6WH+i1Lo81e/p4Gf0uYOe0Q+tRZ9rU8eBwweBZbnA1CKLFjUNkYg2OvPHfnq
XidqQjZrT4T14wl/pF1XyClCBxau0QkwzABpjNljuTUG6dPseLWGhSYcFG4m2dp7
knmrEyJmzzw5auUoxbuNGD04FCJegs7LF0mKPvvtNdCdtJqJZq5EJIhzL00w2rTA
GYuKTY/yRn+9pmY6gw6jEKixE4/2oY/s5MYmWRHr6NjnfSWkPYUaO1SBWOJtSYPp
eBAg22HOA+cjDwynzuPBESd6Zim3wy+BmlGSrEtCX5m2IP/RzClI1+7xdDK3ibQi
WxfuG0KELlYIeEpWFDLyy+DTtv61hhxrwiw1qrwLMR5jYgW2yEQrGa4rqG29tBVy
O2fKn4xIFGf63qQf1di3+fRglfMPGDBPhqwm49P52+psXYeV9wLK9aeZ8n6MvLio
jv3wH3MK08edxfloSBpWRmuHWllUSVzVeTUAgaY9Y2twb/A+08b9TD5YNHNH7p1O
YNn8J04UMTe4fK2NjKEI7Mc5iPiv8l8ekE5ygv1Zn6eX5g172Y4dXYOQRE529gWC
Wk2Xq25x9dQjExi08RsZkSt6GOhJyEGRgfqA8B8UlXYazOvO2RILYQpsz/tIhKSY
s//ZJaCWO5ZEerZENLGL2lYn7IuHA6GOn0ZWadW6dC+5kPBomWOl8gvnbVEnixQP
Z6BpXXaHoucZD8XBagHBkrvtw4e5q9dPu0SIUD2/vKdNeKrMp9g0wWcBWKNjCnsq
4ybi3kIDUqi2vwYfdipWl9MMRJE+FWC275A2EeWuzcNOsjYI/IocZa1oCpOrh224
W9Eci8jowhS3i2sUhwP+0YLjB8AXqhwt0hcyR2VwI3vs1AfXCMbD+3TP63lu0V2G
lV6/V5KmF/7nFyWpYWMsu4Q/lYoZDrlqMLUPINV3z7FItfcyIMbIfG4hGiIdK3MT
9QmJwYI93O6sg6Dyiq6aClO9zO/jO4l38xSvJ0ves0uSGwpfDQfMCaJ9oZ4wFTGo
gWIE0xGzIbcPoXqZBFjx2VMX2rRk4DeBVrmA3Jqw4ee7ZX5KfFJBQoqHhcTVfXiX
uaEwavcCA1MjNydGthL/1/skq+mAj6gFoB/uCCMbvaMCmNx2wRK44q/AZSpBwfuZ
K7GzCCxDqtmPxaIWNNSatN8HizRK+E6ScFlXxgcboI42VJhaDibpLWCWD01GlM1B
PbD1GhGgZZ1HC7iwOYwuEjhmtvsxoFQcXktOJAcNngpFqq20G0YD9HfhgCC9y5Qd
orhvI+8x/+svzLphqadzoAA0VDtw0pWqG6abyHvPHk4OBb1o0rN/tyDXCMCNzIPd
ufT/xodZI//lyR2yEV8kD+omrBafqz0DIPmJHOc4K6sq2uzeo3NfMJIIyqoth8u+
QWLCui1dODwEHvOtEbJJ66aSnvvS3qHFpEuHkqXzdwqewjpHu0mwtnNXe5KmOEad
USulBBrhtGqaikE0zuBRpdDpzih74TKTOEFKnMPF/Pqe3CcV1gqHpycHjfDW+Z7b
RTREo2pPIzQmtl6xh9a4mksmHRml3uH8kB9dOU8Z+DDr1oA6ATb2pQHd+4Tmzxhr
B5N0qv7LFpVToqe9fxFYSut8jE1oxJig0kX6mTntNY0TY+2GPL+/Ujh9/vcvMzwg
SG6HIUQzYKJrJk8OgmAk/J/0YLooN07vbOsE0fLrOzD8RkTNsHc8rSUaCQ+Y8OA0
71ZCjmcJi1ocCLvNse+K6Eu/+qDueGs2xFzQKXIt/t3YlASm5TcngE7wc7hu43k/
9tbxr0B0+Plo2RJ3wazBY90/aKVrl5McjJHJm5GrFg1xiO8SLKNo8px87fZ/IF8q
TKHruJeugmymhJ/X8QmFkBwniTIOrAdQGmGA80bqzxGHYy150LpiPS3jWklBVXbj
7VdfhOuvvqm8oGh3CLbm1RrAFB4XODM678h1jhgUyBlCq4LgJxElqJSfv/CS/sg/
waoHHVhRdo1aVa54ZRnBFZNua9qYLAfrmSihPj8fVGp7fkVsQsQoDu9XosCZG4dn
l4uM0JACpbIJfEdqyfHDbKqgZUOQmKENve8iiL3Xoj0NljDBdEXkQa7+nW0XpXEY
5wjtq37UVuZcTXjZeaN/s6HAefsUhLusXhtErErfWZ8s1aS2/kAeyw4CeW54pEyC
aJO5kKI3sDpgStyqKLfdK82n1VB3e5xo/O6Q9wqaRqwTQWvzj5pYkyHjdJgGStaC
lAuVxW/RdEPG8x4Q285/LqBKlb+g1gGYqtofifsoyku/i3XnLcHhTrQQFNmxZdEs
qjZ1F+Yz32ofN37BOGtB59BK8xaQdKwrfj8KLwpvUN6dDkR4qdm3MkAcPF2xxbwd
YzO658LI7PP4yUl5TyObT9Rhm9s/9XnhDaM2JcaWQvDydhsNbsVbVbeqle/GzxFB
qmr88y07hK+XO3hcsH8ZrVzb2rEZh0YBmFTLTCOcukm+rjiuDO46XW5cUri+tcni
rT8XKIOsctvGOp9zJ/fUvOuy5vuDxdLyE/hfPw6r16R3NHT80bV3kUa7KX3v4oqB
Y0NnoXXlarAW3JkFMhHBGQGOD7KK0cKum4K/Szx07UECZyf0EK3yVtMGrzY2rwdX
7vcqXyfvU567aLOHXBHN6pbE4G9nKsvO8aCv6EbOKNXip9dzj+MN2RPHP4HR6HxG
Dw6bjMO4UJs1wyHB/BAnmqhvlasOO3CL9QSlz6CF6kfvTYrdNsQNqNUdS+kFN+IL
FTNpfgSUKY/u4JTNTKcXvUGApQHMJvcp6A8KdN61LAPgQYP+730RU3b1fdgnTQzZ
J/Tk9AVuAB4+3kDv6heNbYt/DsnUQTXuxzy683KT6zfMeW7YgS9JwVkuxOaRyy5q
hmnZyxlqkyXw4VaeHxg3E0+BxyXxVcjWsnNIrujPY+TkHldAM8LSHEo1MzZ/4DGn
lxsNvyhzDDklr8t/Zj35fRqxAwjt4MtzqJhk1dmfYKXQNdhIf2XiiWaEtlXf3xwb
JI7nsD8bdZtEacCr+AOv/j0RDDm0lKEL271BwKmJlIvJOiLoGH1u19q5/AXODk+z
9M2HNhw5L3C6lSxoSzfT4QOg6G2J8eDuTlEKbUny3UC3ByFrtUFV6/OzGhvLUV6B
cokaz7uQiCtAQhWmXmTw/7/4mL/8iwQ+A9gzGv7VGjYXww8pQ6qUI6qNPGYBxqy1
wJXAcS/3U+B4+4POq+6oRyJtDJMmpXYKsyggZYPdbSPrFh+LHEC9ZQ7YYy05Y7TB
41YMogrqqsRJFrEn7H3eigUOgAePhskVDCN0SKLfiau7qsIeQW7GBUOifjvSW5uZ
6bJfsc8h2uIhVs7BV9xPa+RPZ+76wcAjKlmYynro2//wUPTFCQm2k0geBImRDID8
5jMxTpzrtVuE3qN/S1jnUlQoGlWQpa0OX2EJEJJl2z23aWRztggTkGT67zaZLa6i
9AN0avypg4ccpnMCEOERNWw405mrxCZrd9WKl8EbYgK3NZEPnuCf4qmzc6GeFvYA
E5TIf9TI0wMG0MY7vacUtbKp8BfrT947fv1ABZ7S4lvX9wK7/DfRPOD9rLBXZKLE
octkGAHmDcHUD6436rUhwqJuc2uGa8+Wo89RbcTdNlaU0aSVva+4jvt2CCBO7IzR
H8oc/L+fhD1JcE7O5aaelHScMdbVZNRllpSgLahdHvOjgRANJm8TP1zLoPa0A4qF
6tmSFtdtgEG5QUJI7H1f0OrWrl5WFAPLdpijyNTSOsrDg6WlZNjaqvF9V0BLxxW9
H2RpuiZUFuZm7I9MbzcBWd+WBwtIjGpEYk4yLCXDOs9TXm2hsEJUauRmYQVHGrEU
5mx+kszssE9iftPVcYJfSyRo4IAgUKOORU/+gAvDty0gi1zEsKgztlqat71c9fpn
HHGjztqICCQlIZkNC9hqb0fpZ0tAnA5HcZlYDZDOGku9bEr3WK8sQ1oCK5GRxfEf
36odwgTAf4dgEVTV4vxiAWgde0msDZtEU9HKIsBTYYF5kPg1VCatD9iCEZChthS+
KIBj8Ty8W0UcFEpqdv16eAJHqk+cKhgrEQcJEmo2PeArR6j0lHfpolaEtVrfX+Ch
ghQ4ko2te/v7kiuJtzq4O69e8pL4xJpAvqHiefAFRlTadEtC/eZwWJj77AN5U8uO
NBNhJmQ2Td9yGoY/7MhJHmlIDBW1LDmAtUYh6PBZznuJhmPGBKJAHxSvKFIFNZiC
g+wa5MD45a/nNkMdOpTji/mPFu84y2Vyr9AJqZQMP9QjvPrW5VTDYXVsHiXkGW+Q
zfHB0EqBk3F7mPcxj/2qyJZgqwSpT9LQXZRUPH1YFhHfEZtwGgzMDqB908GVGpAc
ObWATPg/k9ymkH46eSJyBcTE2E2SkUSWZrzDVYEYrEONPpKt+PntW6JhGqT6wCvc
JZHpaoT5ZvegQ/dgOjHqg2l5oYtkj3FegesWODCxMZowrJ/+uTqRwJU5IdgicHS1
M1dzq4HyXVPraITc4OF+h8mtTi/K2RwbyffGqIFaoVbT86kFFMjjYV5w4MJImG27
g2WGYy0RrfnLaK206zT4p5ZhVTg/8IZitzrvXwGxdS9Pn3tNgNjzI7yI1vzwR3RX
RxCTwF9dcx2MnxGuNTqwAB1+7LbdCLteAHWtsVibTfdOTuX7HDu75NL5dhITFcJJ
0rkQTH+5dHLneWva5ZbGmUQjBWsCQo/FUxojbQ2vVgv63l08OcUx0iv0tkUpndxb
4+CPjoT8rWz01A9mtwxxKT+FteRFFPUOIckR/BvoiamvnwiSS8R+TqZ3GkGxFuri
Vvhe334Q97calTu8czMfj6jzLgHPx0LT7LCdEcoo9MpmyCAdrKTH3tMHRO/LU5rV
3YWophvSteygKOtZn5bRY1s87P7HD2mcIJFB5pYhgj9qw0l4+YUnP3zkzqwey+qT
MW19UtGLsIZeBNLe+2+F2C0hc/nTaZKMo1CFwE2SIytFLTUV5EgKoqm43w2bO+Cb
y4nNgK5vsodkXoe3DSfL8XRh62Gbg2PxTsWQdSaNH8EQrY1cRFBlmlZ65W1jsQNp
T8eTi1hgDj5/OUeZevjO0AuVFwARJ+NYx9klVW8HOTwoIIpwaSctCbkbyYK8s+Xb
japotbSzwMiQiWFykabqMYslPW/Ax94ex3fYa3GnhlaO1DxPMoBAS9zu7IKEUeZ3
SJ8Mjqb/TSceveL1WTZb6DhCiOrGpM55dkpC6ca+c8GltQjC9DNwgiF3pjOSk0cj
dN5ICqTkDS3NPsb9qXE195YfrFW7iCB2FhrKfgDKDejeC79WaG2iymFThiskGtfg
GYvWR9kwpdeyKVSAwqq3MdS+Za/IC4wkWtzgqCoCaTDnfGPby0/W0iid29XAAfAJ
vsWEYQFd6O2eyz3Cv2FNMkFhnv+ARn7lAbgdMGI3KNaV8MSc6FMekAOYWvwBgtLn
QTqULtKmcGJKyEFXDW34R01xoUlwIP2cI9wPm4b7aBLxFZ2rU0jj0uiaOMyTaGqJ
CjyeWalOPSVPpWkDE/+ZDaFoTNaq7phyM542VvBLs0CiQ4GUPOXexgxaYZnEINK7
ipyjOVjr+1dIj+WWBv/c6xxY7gno3XKPwUPrupXAYvFKw5CMqM3+hEkJoqUaIx8D
7pasRbnwA7XCcW3MmGDR7jc7+OjxwMccFLm43WuVNFrpwQQB9bowHc+mC9d29Hq9
0Hdwn7Im6usmEzQZU2VOnM5oolbjqb/srYXIEljMXby9g60SNEdOBLaVulSCopTW
EeEtVUj1/ZzdjxXNtQH3HlUk41ZgRy2I7WhIzrpLZL6wrprQDRXZRFLkytEnGX1Q
WGOqsslq3Nt1VMS/c5m9GWDoYR+EqN7OCW/b0jpa4Xa5uLONQZe0C8SiU2wsbHKP
m8pNncIuYybKmAL8QgntO3RvLm/1gilBYyTivvzNlP8Jjy6mD4LxeWJ9Z+K49TS8
vIU5b7i22VQ3gle+Mr5/kWiTpJG4Mqkama3FfuZ/y3nJPJjmrwPQNCBscJI52PX1
T9viYnKgFehkz/v6RbrJ/AWc2d2gTj/fW3G/ria7d4+NXV2icDqBF8Oq5SmM8KhT
gyrh5nzCCiUck4NBJM/eIhhOQOfTw/0OIt9f5ftiytahtjBRcCpy+KsRbpWbjAWQ
JYS0sHHvIAntAHQYF+O70nuPaSQkrrh/ZiQjrH3xgE0RH2YJCiegHMEAgWkhgPSh
qeb5aqLzYl4ZES+ZTXkdCusPd9PIusw9VAnWNiqd16SirHWmJH3TUvRtr3vTQutS
6aPtNRrz+H8MSwj7BCrG/oVYTqHnExoUFHiRRSfzgZsuy2pCYyEToaWh4OsGYmef
PuxsK6gQLFGiv14Z4D9b6YBPB/UDvNd+sd+AJu2EatAI8VDNlODJAxg584MHKh+i
vBc50c3B7x9QO1rJLJc0CkafEFGza08CUnB/BYd2m6ZHwdyG0LhhVNwj6OzHYwWL
r/GU/5+ozMMaZLYtITa1GrD1FBTAJvi6WClzAqFhi/5AtMe1FwkEguptpRTF41kP
gseWN/4apXzGuy9KmMCNdcd5cGEkD9/hR9BWaJPi/pACmdWev+UPqeVpYcgTU/Id
0GDyqSg+DU7I3TTVKDv/hXoPzaWFW0+rg32r9M04ctpjjaUpNMx3q4/o07HnkvOp
1IN5//7oFKluiBGSovW6HTxGQeN8S8zwRL1C2nR6K/soJv0HmrFdsvQIKfCrW5Ir
OBC82rvUnquLr+mST363OPgvKTWHlX0iJjC8uSCrnhBFCZpmtpX/4btV4qntD/5Q
edoscD8Zzzr7b6J85VQllX+qyRm1Qv24cNPJKAfSwXv/kHHI/t1xFrzjcEdkJIZN
767h/WjdmfHhZR1/dwlgHEFnlPWIbAnZ5qzFYAypCQZWxqzYch3sqKaIi60Fir+B
nLof28dZYcOTKK5I4ziDRi0yX7zLsVNh1kdbZAnCuyVn0C2p6Ylx8y8kpfnacKFr
a/CZEeACrB2EPYmIeMKtIvCrdvZkbSeM6l5r9Z/xYMamWKlW/sz5BOtONaKct/6I
hVmdiPtV7hTXUBl5gtQU8iLBaoC712gRJyZ3861LduVyJ7UuMV5BIW2zwuJ4uBYb
CFA+DLbVzrTF2Bdhuz65KKXvEheGV+m+nzEJHNutaNfxIRBPk1mnS/i6hQuvX3m9
FIFvX3bqf+4nBXSVgaY0O39rUGpf/+WLOk/PcJdBiwpUO2SmFXloIboyNDutPLWb
QXhPDBD88NSMI39GV6eLnFW5iBhpuJWDp7ju61v5KRMj+AV20jiciiDl17bbZXVD
inuMqc1j8jT4dF98o2YcW4v0oan7uKwbIpw3hZq5J01dgRysETAnN74XJfU8CEX5
4ld2tL9nOI0t2429GEl5ydy37cM3qP3SJKd8f/0tnG9e5Y/gvhd0xEmgvgEgLaqr
e4JH7e6IlZADtKjCit0yaj+rCYlg20wTi8zxA39oniO86G0lK3EKVNZRp03TL2bn
A8GL5+D+cEpDmlnI4Pcafdb6fn5ckUGj/h8V+QiOKYUQvBeZs+TD+y7kxFhiCt+o
o76kfAQ9VTYToQua7aOV3/2hThOi5AyC1KdK+rB4XGXW/xy2zAYqKOQz9T8Qvqws
jHkKc0shVTiMLLXT3CTanxg7o1XFWUNIlQ8Xc/KEA4aVhE9SOxikig9GnqFX2DoU
ASDTlg1MiEe5BmSU0CGEknUOILwqcR+0Y9hermNAXgVUPQ9UW/WRk/uu20wqwE7J
LkJpvB8Hc9R01MV94rj//Yprc1hMkMHZ0gUXO76fsZR4TldoySz5Zfz4F4gMfTWM
dJxmn/M77SvNbh0/UHJ889LIqTuJY3j1gEUG7iXPPhbErwlAjHslanqc/ONHdwrz
JXPrTKkz7wJGsy8l3NOZpKiRINnA5GMjncnUp//rC9av/HtqHtXAx0fQ86bd9QWs
sWvNUdXbaqmHjI/24aVuXKl04Uj7tYV8/70ErNCMTlVFpqXW3EeCQxMMj24v+bnb
hi6RAB5l0k3DPx0f4z+Tln3NL6NPduTOm3ccLe70iWoy9Q94JMoHwqWpnRAE31Um
pxCCVMJtwmpDSABFgR3yj03+jIVYao4Wc0xSi+PlL/wruvTMFf9SKyXYG8Sew64R
R75U4NWq+5nA8RAzMbup0pCbyYH8HkuAjKlCNkaZZ791emX2ct0fPLL9qEfQ20vW
jgKGtTlEIath6Jbt7G4chyvptWooGdV0HntvXNMmRzMws9S6EG8pD9YpkJOcCcQr
HsB/JvlMehpJsRfNvoQXV+/OSHN+d55bwJ7nYOeAXlZgYXLxsXM6+cqZ3lxvDx9W
M9M8vAk0pUvsQqlfmMX9k2+gUJwIfungQm/vcOJDcONH45lBhhP2px6E/mvRgmv5
34f2Eh6VCMjPj0LkoAEAnr8noJirpGMWpEN5DHZQZW45EHGdMwkbEXF/QgC/fnEN
EeyN1HNcT2lO2cIAqn4hDBY2IUJeMXPxIoL5aXUA3gEi4G4TZ+QP+ZXVhJ4mL9Hi
bRj+9wWGKxKjxQLkOReycaH2bHFtFqGaSdG7tH0d9W2QsogNRLgbtb4bVgphOWiO
8N+XbLWbn7TwpA1ocDXSAtRuvTkWe6j8sTChaykiyM+0sgBXQDdL/5yxk02W1P++
vYTrNQnZACwJd70zuMvJKU9V6cheFSEOuxmQej4VRlL5UzHy8Cfy13Hgmr4A8qxU
bclDMpEsGZoVp4nwE3EkrCc5Tv1NQ2difkqoYYc0vXdwAis9WrXXPw6yxf9ya72X
y3n8akARX8r3SrZnTK/a1dATKzIP7OurHnuD6W1HlUGYPuLxr8HNxGMx8ktdRgCy
QHtbwUwNZY7S/cgWEJ33xdvPt0PY33Rt2xe3BY0CmrUmrj5CL2FhkRBER+2UJPiD
e+yfVi/rtR097tD+/LzdfFSpO8iHBcOd3MFPV6Z8GR3cprZLWWOtuO267r8lQdns
Vn12Se5jABjpx8uiiIKPBa1XF9mD7cRlSdSmjvx/i1ZEyzlIsOcVxZm7i3DgY90J
cdbp9Uc0FbCroZa5Zt32SMIKVPxGhXnbLUwwA6CSrzIXeJBlKx/rrriiXIfUQUgR
AUUZ2J8qas+UaEOU8Z9IF0knDhuRV03Z2rklOl9B+aRsT3O8kmxBC2ybOVKUy8S+
L/eS2LLKG726BjIRxCZl5YNL/x08Aho2VCTRdB6MPY0iMXeCUQTexL9PUwD6+Q7h
uGVDSxs1h4mteBEfr3QYnrdRSewkIwMc3XqBR7XxhEieawVWXKPKBT2J46Dn44vd
pyFMpcGQwoy7+Yq+sI3eNDB15XZ37PRMePhrf4dwk4A7GrwlVWfwSwD3ojnF4t3G
ZP8TqLx20sd8EqJAnuFCUhLABALwQBAAsT58zMoIZ5rk4FzlKbpdgQ1IcNTwvQ6t
TbC4RfGxcHHF6AtpShhMYb208Pwd+xYZnkZBv54/XpTbsI0F/9EW6mH2WYrN5LVH
H7fGYQH63AVdDsYgCdF+CFstdmE1ajo1ePLe+chF4kPC6cJpbNf4nestS1vAi6JO
AIzlPwfwYJbJEOqPNF+y1klSI+vfOdzFKoALnqtWnudn0VUePpYFzGGO6tDv0w2v
Z4msPgxv9TbL1z9jhKChBtrfpkzZPYZpBWxvij3HnbPsQXHOwX7J3Q7omR2ev3/P
6P5K8amfJ2KW2QM76wFtbqoSav5u4cBON4Dd+KUMyVoNu06wP31UOKhQlG+uXnd5
qwmhMd8Pkf6c2QbERcXPcLlPaShLqTNtJ7E8svu5agOrhOOj9FfQH9v5JifR1RlO
Vzj1Dc9rChSmC7cEvaQIAxQHVr40gmM+zIh6oBZieOtcRu40ETY+7tUgNCoMi7i9
e2A8Z/nFHS7JV2ekzKruN3YYlp9yQpJiSeGVPUoeL7kc2zpVIebzWvmrW93JxK9y
3pfplc4iViTESMBn5m9143RNBY0h672WxBBJ6aCgo4Uetj0s5jn/W1/SEeetUHPo
oIr02f6IXXnZmzHz4ElWmxVAgXSvhvHTIvER0weXMjkJhkB97SYRbn/7cYKGbb0e
oYEcAZVKAGWntgWH7Qak0ASD8LofFDi42zH18hxBABW9Y9WkSY5Gx7h8z9Uw7+6T
bjF+fYrKTf8B32aTJAyxGJN6Ek7pO9ptxkAjLyV9BoFdrJEFhbHgAgPRvK5ZaRSo
UUWhAz1LxtF9EjCPTfJ//XI1+weKLgN0Kq0lSXMvqPqL9GhHqq7YgStooHrIFaui
Tp9A5OnWt72S+vlDo0++eHa/EtDhg/8HSxF2kD+JR1y/5BdXAiga14fmZIV88zJZ
U4Aejy6SyHo/0FnoNNzXff7UBch5Yov17uCRQYecQubMYkQW12hs6JAOISt06sfK
ClVg2HgteSkIIiJmfn2ABoPoulqt/b6Y9t08pGnov8UBA9q4irRzJhNwrUg8pA4P
5tcoWYxijolEcnyaI0835wBi7u0aAxeoDMIDJwAyFuCvKs0jrVrqd35ihko302nJ
H32oQ+ZI7ENztSVEQyxdupxdBanaKxUGWsLkBolI2VW7lX6IBPrL38M2TRnXcQhh
ePuqgkOJNKxj6CKXD6CUCK4w9Ih7JHo25E4f45LMnd4o/bi7xKj/yt9RnUIwb42d
H37eO25o3NGT4InPp8g4q0DlBkno3v9JA9Vx48hRb0TUXaOwUSEV7DZY8TLlLle3
BrujcsyRjffrnCF/XQol4y1wQNu70l8X3iJiqKP+meOCb8pjzZdknXIMMbqTXixB
lUoVrvG00HzM8EBWW2H09DlCBVqG4rHIZ038y+VKNBA=
`protect END_PROTECTED
