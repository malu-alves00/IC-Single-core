`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oJJxTrMNKAheKdPJHKcrowj1cPRG30YVQ965Nf1/SXVL0LQkxGbbHqZ9MJmspqTl
Yc0nEkwaf8jMZ4NoLg6ICAnVnXxXKEQGORW2bS/J+qqepK5/9yqyNfXKyaXOYfyf
MvDiLdwcOCvu22vhoq6oioMvoXh6AcIO22+4VDRoP+FORQnXxkcHUNW6foyLEUro
cL56tA9pUGrYzREbVAbXpKGfNAR5wbGGF/GNZ+r5dgR4DTwdQyyVfm/GlbQQ19f7
sOKEEYnfe+E1Y0zGwla0oHno4oynRjjq3LJlvSWXexOA/FpvPUaWRCXsXM78X7U0
/wFrmaQCJI8gXf5NAJo7fyPAvx9Q55JXKEJHBnmj/MQaDV9+GALG6SsykdEJw2Id
bRmeyepRfP5DduWWSX/0rhKytpv3/FBpty8QFIkZxAhlxE0vAeXSDo5bf17EbElu
kbwQla3TLsLJmBBgDHfzZu+KFN260gZGcO7KCEPEroLvVc6ZVGokrGCQW9EMCeDJ
PVqwosfPPAvZNx7A3Q2Sm5grg2bR4Lfj8tj0hubBZeQ3AelWdtrf85b0e/n3TBla
V5Tb2a3XCZAESBjyzfXbeVteM+TcV27BMlQMOaTUpIqdkUYDwe1V5fP64BGrvrqj
o7ofVc9i/uxDocforFlaQamlYx63zaGLSMf39Bu4nZOnFBVB3qvI0DeXG1wp/lDY
UoSURIqxLENhFH2RtrFFraEI9sb3PX6rRzNeeHHJAhUvLwjYC5E6xxxJc1gnsACT
/wkUJ4dFMAIEbvF8GsuSYWlv6RB1Dv5le+Vx1K5FiN7Tqahes+kd5k9d2OXmIpLD
iTLeoT5By+5yTC0DoxmZzGk7FflD8+o827siVGwcVZy65aYW0zfIsXTxoPeeG3pT
w0VuKoqTPTXh6blC/gCh7HKC6rad+FkZxWshkxmMLF9Ddf9tvQNjhq1hssBvRx4p
ISnSPPL2Vej2iCUcsys5W9aXPWHoajS5S9rIRlRb6wZ24fTqBMAtrCs6/o4+DYWu
KYmwd5BE47/sdzAwwm76zTBj5IYW4+P76Up5uEkDKmmB/794miKwZ7l03SPnn9u7
QgdyREZUsfJh4ihN6YZLvJnvXmsobPfZ9j+p38Ig6a9cYF8oCz4+zdvWj+eGmYkG
9xjzsEtR76H8f3/rcYvEeonREoSLIwgOQnzlmdsvTzwhLvJ4I3BCQJr0MUWgtS6a
MRABqQYZlU1HtboaZkjw1zeDs9lfziU7giRsVlnvZXBQpZGC/3cqRiyzZTeqoBRZ
Txn8xdwpbcyUbOAqQ8yBD8kuVWoxfB8xPGLEQ/YfaizZ4l7NzHkT/TBETzjRlBTD
E5aCLzI+G3We88xxxhhZ/PK9IA4b1Rx7WGW0vM+7pFRPvPA8aWhRlsj3yygC1J0u
l1mIHXMvx2qF/9//E6IjkQeQPNFufsBzY5Z0DHByNPgSHRInn8oizwCHLgBWdZpe
m3YZlHmCZrbpfjghBViVgQNbZ5A8Jcurozut6m2ONLwdBNr/vO2gPglMF6I6WMRC
pHh5D1gnJyUUSrXTT/AkMMJghk7zpTHAHjx4EASE1OHDtEXod4t/AeAg+Fv2TShq
ZxDCE0+54WPJwsRZ5EEhftD42DZCv9kNnxsVA51OamBj4s9zKgNoQN2b2qkoMQmQ
oTaEGCgBrLJRLJFHtADlZtLMA5Jkv90uuGm9S7x1U4gPQFrrVU3WnfK+0ACit31J
dNBIhigDtQUQR8DwR0RAno2ZJPaGnw+MVr719MxIVmpfkev0irf9BpArDEPplUaj
bwBM+Z+svRDnx4Gkc6E0rQeeTvzVfuUDkL4Q2jZUa9dFMFfSE2rC6yugXtBSYxvm
C3NJJmkrt2KsrEwzhaGPyJ34FEtXPgiGw7DOWW1RTGgugJGJwW3TMVM8a5aj/ChH
jV3I1Vpwdi7pOopEY6rlgs9/NC4JzK28Gz9ZflEdLC7wUAEfEzHeq7dmIHVrmR4w
RyxOXFoAgJuDM2GS9/H1lIYqQwHGktTsip6UTlO6xm8jUkLhuDmhoTs8C184bwoY
fqDF27NczQxIwF7O5Tc7nMnH8bHrOibe1/lEXkIbjY1LOSTcV+ta13sV5sHyxXfe
BsqREqvujntBqzAK6kwC6EbCAyCaRbqdO1CHMVCSlBgunYhg8XmdpglfT63qgN/E
WWk/0vtLty6y38oSgwhryGvX5uzsfakoFutrnHRlaBLGYHDL2mrRRKNCL8NtL+K/
cEgKWDN++n4Z20iw9pvi8Wro9YLdxdAX1noNVGUaWVSd0DNg9+81QSUnoDPHocyo
FdWoAvYwncS0C1SLXGZf9ZgmovUSgd6j/DC8C3NvHHvak+3BzEcKwjoErF50HSFD
2hE7RYfcS8WmcVp2jC0/p67zsSTMHjV/VKR5cX101YXoQpbcE3Wxwbjf+J8+Kg/v
e4Y9t6V2nE55B0rDj4XNILf2sleBoe7RPlPiK2xkmou+PKxcD7y3sH5Y9tq8NG2t
ZORvj9pJeYhfqBaxHnyEtvcOrB2/4a1+6SY5O7qXoCdPtEQE2nL+dhcVFAK9y8eQ
piBQyRZbrTQw727oGEKR2fqTSeOqI3ew7yCeuZmTBrgNBmERSyGjz8mnCI9wUII/
g9Pq1pGE3HbeHNe02HeJ5oOwtIVmagKZJrc4aWW6TRxumaQvTpCdjYizqXWkr4UE
NLlDtbLwIJftea13Cj/My11sp2VY2k1CQF3hs2zFO2XAWzxmsQy5A3pLESHnLQZl
IDhYqVMPBUsJSOdaEdgRxOUrzq5n+d3hwdV4t32U1taz0692IUe8GVt0M2TX8jGx
92fMJksZ88GaqU701jOnrr+wM4NZHOFxslu7y+lHyXK0vO6t+RxVyUtQEzv+AYel
Ej7gMKHHrps2vD2mtV1awhdL0c26j81s0O+W4g70CSADmQ+sUjTNykmzL2byBAti
LvzZkBDi0XlKiVtW6pqkJ7Bp/E2t7udMyoqShUdcmXVP/eAPSgRrX/4KKcQzAcb5
s/C+J2vYuRZRIHxAxJjvD+fV+fYzjXnKW5NwAAD6m5+0L+BpWKDO/TcMeu9Dexdk
N9zXFwq9K3WtqGkdksDbWZ1rqGMS6sxvY2xv3sFVrz9F6UwPTZMhC9XLMYW+etpA
1XacHRRj66lWmYulkg6WZuVeKBXHXJLdq2U+83X3fZ+m4t/VvY6xBeJcX8ZlRrwv
N10idnN2A0WT7Gz2gdBo9BeWQI8ngnvGDeExoz7xoOFd9dS1vXg8q9GtGzvQ9Um3
A7PfnYs/CcCiUpdQCaGABWAx0ThUaCTnbkVioGH3bR9q0IztZzVOHh4kyoRy2EgU
kHUwJnn0t8YZtmlzRJjlWSrM6jCvyOWHdhzTZNeCMJ/g8Rydypy6nwP8MUcjA46w
NloQMylfaLQvvV12TVshMHF74MsSR9ILYJ5ZV9wRt4vnrTxWQq6RLAn/8Df6Ea2b
A1qR610A1fzEZQzrTDZpVXumpEWl/ntn1Ie+fkAl6Ll4aYJ6BMZlREOdvlt4Ay73
piq0ll6AHtR40OYRob8hOZ7CEswTE7iqlrfr/fyK4m9NHBFEDQhYmeTKpPXykigC
31KwyxkTJQxWUlZHrjcXaU/im1i2GC1b1r8Ah+QdBmP8QOT3tZqrB8NvI5Q3QGxB
8VOSqzCKSUfeIgSKZ9sZ+xoAG4FPeHSni1WShntzHstDbYMIrzHCoFGnamIS+WRs
kKtAQCmjmnMRJeNk+XH7uBfS5KnCeJtvR8X4VXoysFWF23v0z3SFg4CX9fSbIAek
u+9twGa2hO+eEk2DvPkuk3ujzsVSKCyEjjieh/WfoaBh8mcm+qS3KMIo0ttO2nhz
RDHm1nKyd+PJLpqAV7jCtrK40EIDAM3VR54xhetmsyyrOjYrd6+jze6v7o8CLcRH
nfyUmprNnJdygPCvKs8UiNkQYPYVhn0qMBu/bzmbCkK8VB9dc4+rYyChmfOmtaAP
Dxk/OXlVu3DViU8qtRLMIjX51bE70Y5lh+gzLTEZPfnCHu+bDG7J0wvz+7AAy57Q
VEc+F0jIYnLqlN2J5YyZmaS8vIfg3IcXOW36bxw0aSctr6fLBlD+MhArOmS0QmOc
DPjPecjwlc3SZ4B5F8LFnDlM8S4sh9xPjZrBwag4mVuQWl34Bw1EyKbihJcAg9d7
/2MQiDGrqEs67suMAekRHorGG6IZp1xXrxSAvCfx8IFpVRHeackLefK4OOlSsXIF
2SUwL4IbVVbjUl+7TzhSCv99Rr6/6uSCHeOiAtXotA1yfIuUlbRIOfyOTCLJKI9P
KpIimNsBKKx1Y0xprcfv36BJmgmcyILnwnKUe29r7aotEGO8rwKX/eKgfXyxP9Ne
bO4s+K8dOBsr7GD8V2K3TsYOiouPGCpq6VNREc0QkSpLalQLA3KS4HWb0XkTKv0v
8qlXLQQQ4GD9qw1oWJcYqL5AFvp3tkeIifGCxLJ15ts0fR8KgYW23wX4fGqtiDK0
TxOeUnuAjUNZVY63bGUDXsIgoatLJZXRJGhZgkevJ5hIT8IUWH5cp9MOOv1ZHrHw
+JaVQUC0ltW12w+eR9Tc7FQOjzOC+guew36yhefMef2mRd4pvDCAY7lFjJkAjK3V
S29RCFgIwBNUVlCo77f+sRnKW8WBviyOqejokXZizcTIYxMJIqTMwiuWQtVgsCb4
swDmo2OkNrclvqpOq0rUO4QfakezP4U9gDcgGZiJ+JdKHCpd5EXNhklhJ2HCpMbq
+6A/I1i1LGsm/KCf52zYbCnG6wkXgeceSJF1/AQjfSZ9xk+ok9lfU/i7vHYlbi0T
xEjTdkE15tcU9h0qKU1SS66Irm5g7N6J6OtSvDXhWCoaH0WCeRMHvPqJKmzACxTf
OrL4zrkjqFo64+c08KWxSKpmc/TLRDqw7tDyKC5hquF49jWs76SWorF2E05H0NWk
hQs8DHdPDdsUuQEgLsR/t49JG6hqTzCKY666xzLvTuuQy9Cum33wgGfPBz8kh5Bq
wCfm0vnaDLblfFs+KCUPSwp/dLGGfMVVzdmysE1/s3LCKe0AhiBA8R1sE6W1aIly
Qyw7EYC/OUUFqBK6Zko/H+BaTeo6nmiZHQHsN+gSBtfFL4ziSneoOJCAT10jqY7C
hsleh0WzUgc7NgBVoIKI1D8vN5gVUGUw9f9AsmGmSgraq58f5S2yWojWZjdK2jmf
2Gaon3N346q1LrH7xsyA64PLBj5/ULkrUDs300FyM7F3tR3IkAjL1WvVehMFU3jF
rYDYNQb0XMyu6ZiWQlLI62QAm/bCk2EVtl6M6vSNCzrBCBx/LyTgUx/Q3SRlt74u
/da4t5W6T0fytj/sJn/ZshI9UAXPHF+4ZrQJlRq9Os9Vm85Z3doE113lBUkx/OMQ
U+eEevjf73+XTIGfQUnUluudJjIkRBaaoBzHmSpBfIjSfQZDZD+2/pW/pktVZvAj
sYTVQkN3fkx/pDYPCzN39eyxDA0zwhOKNyXESdFoKgOm1JgwMBu2M/4jPt4WOcbZ
GaFWfad4FbiEEYZ7nR3WGA8z8buGE9Iu3MPKCPC9hE+k1iJZ692n1DaPdBsVAy6g
UMixo9bxmMBTfPEjFlPBnvuimH4qbFg2OyLTPs8k9WgJRU4KasO0nhMA6spw7OFL
CfGXVOVeooUWtbQuB98mbRy7xPwOcWfmTqpTfQ28X3HWU1RsVJB78eR8dh01BxFs
jorRMixqbrRsQSjTRP42oxqM14UmjdGI8baTd7ZL3LkF8CIWvtMFO2PBsM//sFhn
+WnjFVSg8FV7ipuiHvEtr6bMe58w12d5DFlPG13KEuz54xhH7Eo+MXTbmXyvlrvm
2OkPcyqrNb/eNoj1YMyO+3AlHEZshv8yxGMd9kZ3w0PsByrgVFQzH9LisenEcVJn
vZw87CSs3Ho9EZyR9PoLPdkQ+N8y7GC5saXD2GDS4/y7eiEMpJ6cjqSQMvZhZ75M
toyHA600BEvUvPqtJojLcc4MoOxcCGyiZcOpgrkBPcme+7tKuLTst4H0ncRzoUb6
C86+12+5bRRoZRd51ry3y2WpFZR3go227eoEDYu7PMtmgtQTCel2IJXtchBCJnGu
Y0H0TgJ9dtPQHYc7EpIN71R245BgmkDej4jCu+JZiQwLtAgL7/SHW+dXBMbvF8qr
xViWy+zaDajqhxDp5yN0hhI5fe5XrlW7h6AvT+b6kVtWRkerYniYPvU7v7/g4DNf
mjtcsI/LT3H217yNGdG/AaHfXwhQokBsX10hRDzXwESD15PC9VpUweXIsDjlLEES
zXcih7CCJCPSNYHZ1TfIe7o4GK8e+xgYH7i9mi1bpIEmGMyM0BVvKn/iAl1jDiDj
N/ewPbRoTyGSnqND1sRClEcLL8MMTIovVsD//4ERT3P7VRZyT0jqgwhbr1cxbJvt
k5Y1/nTmbxsFTSPWQDwPRxRLJR1M1wTwaaW9ILmtLY823eqGNq+f9OBW7n2E0PD/
K3vbSliWdhAsEFhitARu0F5dsteHiMXMzykFnNhGsf0vQUgzWshNEavb9bFvqNPR
oEDebnySoE1WxfrJVDjrClPODmsxSr5EKIZNZj/hu3SXRPn3/0sJ+5LAM/vnCmtI
PAZSgPLTXqXAYBw77ijKuLJ9XPrJvMM0I061eKape7fkpsb2bPYUN9dRgrQcL7Id
kIdqi6AjppK+hbog50tn15DgdG5+21rlUlLRzpw9Iw9icw5JCdF0atgFUinalFY8
GYSbZXtaqvrIesm/y4ZiKHVYc23rpwcSCcZ9/noe7K+BVvhFphDxx4HGPw6lrMVX
XSQSjPOMT+MWKO2NZnYL9tC6EeX/HlHVThBKjLpH3OBC5NHr55c4+QN4Ne+sf6Z2
QFjVtz829cR1DVJib7fHbZZkBM6LyRbJtr372lQK3lDIu++l72M9v/Ea/dg9IyHw
9RlczBnWeXUInfj7feRco4HhDhXVMmCNz4scmC2gkzPcRPtF8/uBoxZD2QTIb/Y/
jQu1GgS/kILzIWW5xhRYLY/bAIY0y96ZaTJawdrsrJpA6oOKM/u+4vdc7wkmcc3K
HYrb5+1byyFFpIQkcjnqQGXFbCmXODytudbSKWeQvJqaEGKkxZjeTKuW8X0wsV7l
dbzNmZ77nMfH3Ijm09Rnlg9Vv7+1qFTXxvj1AObYOyU5Jv5Oh8KfVMbIzNDd3iCd
hfGQjk4SXNf6gyvtv7g8y7aZZHdJHmLHa2USczuAXlmN+ZyYLnqb2QeQZzd68h46
yNXJPs5bgGKls+OjwKSIvx2e1Xe1Eg43pDcYEyLCTD5Rjj23Y2UlUWfTOvH4JV1J
0Fzb7i1zkogGFttcbPx1civiKXTDe85wSfaOgu+MaTX8V6LbTQZntnz+2zLss+x0
1O+A+DzY/60XmG7H/hOeS/pd1exVDQ4LYu7PK9z7AfU72+KPEsPXsZcdFZlFq3qo
W0u9zCvo1Wp+boKXIY6FRI3rRJkdemehsONpo5CNw46QW+67GmdpCGaDCspF3iDd
qtEjGcskRoMHHtVWaRplRPkmUoazfbO0pGzXVQkEuSD5BRVvq+1ZxKe9IOzf8zsH
Yh8ewhL+i3o7n+mDYbuT98NkLL1/D98gEbAjFpcv9BAQHpJZ1WK5O69VM/6LY631
NKMBrnsJm1JcFQj26e4YiWRnHArJP83UBVjFciyh7VGrU8KpQgP+jfSfZfxj4n+E
td9AAOv99TZ716LRdw2Xj5isxTT8l57zfLgW0gK5eq2PAw/Ws120PlFUa1/4nqmB
jvKp0Qnae83Pg1DlSkUvBSNgifYJ8l7OSPYhIhjrkiPJNc/+2b3+d0fVTr5YL4rk
2idfzBGNveZd8Ff3AgY0bwuyESL3I/adMm7ud2OdwxvyjoBVtaWhTf3o03qJCl21
+dXZP7Q9UdswUymZYTjOjPnDV+7GcqIku9MA8j3qSCXErC8ZXbCNbKSSlBfZI16a
vUPoDZn16TBTpEVG3SdvpK8EFCIWi68zTsUfZ5mDszfeXzpsQz1DK/nUXG9+Hk24
k01UrocPT1Iv+Cz0DbCNsnUhN9nmglLcMr3Ua3v59Z+SYsDhrm399vVh2H+dGs9q
VFMdH2h3SEHgAni2sgXVy1YE32HXvprLO/fCyCTlxasqfuXCeoGFBWIXl+xeYNlI
1D6/jQ+T3EZVFQ/urGd9Q7eKczMF/jpqHquIcPXYV1AYcehRrqw3YJLjoHUBzoo1
wh9AXx+gUrHCyS3JuT68e1o4+W0OOvIPXmPu0GW0RaFeAUjbI5DDbcIMaGH4Vwlm
GfEFFuWsD+tvjbosGhYf8RC36Z7bfxS2ht7CM2CmKOxxFNqUBbz51qK/TN/RLbqC
Inl5FOi7SW9bKABwL61G2gTdlkX0XaV/Z4yzfP/X7o3EPuodPetX+OYpi8fJFICl
S3+ckHlFpwyTBVzYUUrNHT2KHWptf67r93zfjfj1FqfMo9mDId+i8Yatmj3n8yZ+
UGi8zH8i4Jgt0aoyiiURGOSB69yT3CsqtGS9Ifq5zLKgWYdL18QOUfvnLwXduf8B
5UE268LPcvTNlfOPkME4AlpFXYx8vVGy0EAlLMQlNGe6FK/FN9XxDaQZ7ni9ZFO8
CjhVzJxLvujk/xP2FFnjZQC28ZS1mOhpWk/Bwu7OvFwSysJf2fPQBkWlSfEZ9OvI
L9vSDG+JgRSVBXX/okqyBM3zzpZEae1cbzf/Je7mGaAskg2vF1iRKcdQSPpc7wkH
KtRqPxUBVYalSQPY9lN26Ml8BRbIk+ZAcIJuCXp6iWa5CuH98OP4+VBTcMuOwUqm
9uFj1v6BTUPQ85ZnoUnw0xIGsFViWaI13H6cadIMrqqgzvQEgjhms24H0CY6lA5i
L7o9z2CXiRlf8wPFGh8YGuAlhEiWCYg3kW1gkc3au1DK03Po3P9eKWmnwDP05BYY
VRaWNNOw3SSxAtPt+VaUIsj9EnvD5ShBrbql6f8/FH9MtHtBNvPe74xsaBrSKZVd
AyPq0Qm1JP/Eyc8/ZbnP07JrFpkR6PUI5gbE0l+IGlUoMuFKJ+wot8nHXqTcuP/8
TAaJbOwGRydTOCJWVAVCEYy1SGiuHXMzry0pY8S6W7Fwv7Pl4dzeQwPF1SkLQvbu
gBF7EIBwh/6QHdEUecfvLaCp3Pw2F9vG3Mi5uC+mLgQ6/wFNEPL6xkPTH9GW9kpJ
vW/t81yVNxGRvImGckR87JFxsHo/0lwIyHRUfYuap+4k2xNOkbT0J+HShAWyVKJc
/2xPfH4QYx1s8DXEUh7ilOJFWHNppxaTuuiriqpe0tEtjnyuk66rxK6r+y8WPwF4
r21lolMPKmd+OsvGf7bQumVIxBfbcGVdMlNmEcO1RnywGwIkqA5LSXEzET7REASG
9S2piDUmPpJdRMIWh5vx/mem/TdI0wWX9AsMV5TVZl6pBXhpVU/NAvgkyVYtvIGI
wp/8+ZkgRbSMP6oWoTnEefF2DnFZXsePhOGeRqAT/n5hPaS1VOLsMAfbsF75HAMP
KWKna8MqRI1IuHcC4FKjYHr8f5e151yz+2hqSa/jslaOKn3kQu+hnrHSeUXZbvz3
aVqwydDLJiG7e4BFYFZbOZ8k3o5cqLCg6/nC2+tV3cbTFoHdKV9/XH07cNachxTB
YylzDbKG/AsfJLgq5o4Xg9NdbgeERHjx+Slcf8qfJOEb6jbU94D7GBN+Arhb7maw
oN9BlZSbDzLIlO2SLPD6NzQKh7qEnpde2OFNSnYh2xKm2snlUSzd5vr+33kFK/N/
YGrSELzSnMzkon0t79rzdV1/gmByTSOeeeR6Zo09JWROHSgtoOjMnJwDfAfVrSGQ
RBACU6LSdHAddb5kotnBfu+92nsu5/eXSRKbDB3p/HFx2XhcwEb+0eB5hTypOoaw
0Noa54zfp+YcjfXZ9oyXkS5QdsI39hcZgcsGlbaGevoMSs5bRT9BJjRN7IyKSVSz
D5M4Okg88zj2WQL9zhPccBu0qdwGdjbKxgGTNr/6n4/LWZdfLJ7EqWzDAFGhTes4
bpAWfUkkRWwHlzvft18lVgwJmavETZbG8gANd89IuHBSVC4wTSgGFffp6Xro5Dn/
kR5eRy8TGeidW9oHYk96I5ZBmAWxUf227P/Rjgt2YZWwmf45iEgoazXEtl65qqiQ
gqXAmKOQARpkdW0juSdABDm4SlimAE/K4900VTHEn4vqxKTafVuPSnOaLnefr3ma
9L4B6Ka9uXUjUoMMFiT8jFAMkV5JpzL24nEF9Jak04dkMCWvEg9hKI2j/An3ZkzO
GzrMaLaUO8qj/6Lr7evfL2ceXJMt6SjRzbCk/6qfGV4Wa+hJJJIG1zUtqiL2BrAU
UeBKWV30EcIYixsdbWIlxj1CEEMI6CaCkRyxAQJlaL8mYCxivH62wR9vFhYKaHYB
UiLvUsLF+m51iuTRrDW6Xu1VJV/ROASCyrm7Hs+N3GyiV83vsa9D+anKC5qudY6v
B17+h/ia2l9vIQdcchc1+XQKbIXYgoha7vTAIh0nfOIvc08H+k8OPAdq8MZKiggr
K+34NR7GXRgC8kuZQsHB7/q0OwzaQYo1jYq1lKhJMYj/OC5g4LppNnX/e3j2JioY
QYXeO/zB6vlAGuiJubUAcv3oW/vwqBzqWXXZu4xUd2z/NaIjUFqZe8diOzk30JaP
VQU96s8PBq4c6GPzAAFBeDbBvBKT6yP6lU7V6Kbx9T4QdbZ+kmoPMakZeD99S5n2
WW2cKfhtDI2fuOOEIMvaL8JyCafwWXt4DG8AXiMIMtkZvB8UJpOMoFBZ8NNqSoJa
/nbI+gzxn/WfUyhguhpbzdb25IhrWM09l7/7ABw4EYxFXeQD2jyBWgg2CTk52hMQ
d/i92QBkq7nX+uvA5D+3/iowDoMpap5LwdYXGyZjrtHg3KGXfqLZpSiZ6D3g7wUX
ZRsEDLUzJwI9Nh9eItugO4L/BHcswZQLs7IbuxhAFUc69+8qoowvII/qbupkWN5y
X9q18ts2aLrywmdHADeD+YkwaIDKF3eH0GB/ke4R5L1wXr4l+dGpkJADQz0xkg4F
oqB5kv1zJIoUFwicI/2CY2EHtyKcocC16ejG1423A9ZWD2ZUECVvp1TZR3MXwdVs
ht32yJo13km99y0zqtflripHx/I7KWk9ViJ9YoLo2MD1scRyLT2sOjB9M5SLJU/H
bDLOzumzvAnsb5TnJI9l+2qhh8m0t91REXaxvivfZnZg7bhLLr2f1H42p5OjYhA2
MUxwtFZ/3dBKxRWSeADjjZvJ7qu6dw06ZqCOtigtqVAGx9rU2CzMVonsZAX/o0XF
af7arjyP3mjJCTy5GLDxIw==
`protect END_PROTECTED
