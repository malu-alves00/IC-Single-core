`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
B68W3Ft0/w6jAqe2Gt5ueBwaieoK08gJMR5YC/XjZSgX5BRyJ40JZrOG4PqWbpfy
nssdz7+Si41xVB7S8EoyEcGPIJMNn0drlGkvy4lwYRa6CBolHFccZMao/e72Emce
fi3Fd4GvF5Ua0YAxUtusyIRfA4Gzv/qZ6Oik5/ugQyoxntWMJbVk1AVwgay9GU69
Oj17SQjGFu4QTXT2imvj46R4C33JZU971CYn8ZA1pUXhwajoRpdzaVKCENiK3r5u
BlEedwMxxEUfubwdJftHRjIaEdmBzVJzNW9QPkAJdFqKLQ+clGWSxS5c8Lpv08hs
qoHWYERl0+EAK1MBgG+FvhAj3zatJ3HG+swDpBRtdXU30tfU5EjLd4pTzsC0uOVl
y2q1WidewKlYnXWZx7huvFwbnSOCnNJ3rsj2XT303IGrxL+FDjmrtaxRrF6f2gB3
cC9q6larsfUEKnvlb0yR8Fpg5LJsstdMS7I+kDT34M7HozMxStCU/+MS/GBZVfcC
Iyi5HaCWJVOocPHtHIBOlxhsyoOBu8JPKYxR6iYr8ZmNgf4RIUol1oC3F76XzxWJ
E9e4O56Atims2KPzgfSCRt9JVfzmjIxfbJAHBVlz1Wn+3scjTIT/upI89k55WXkR
DbNRmfoRBbKDtyNUA6lq83rFWED0vMUNpTVdW/qnNZtJB9b+STPSlMwBkvD1DfK/
90QM2hyLgbqDzKY5CdQ/Cp9P4JLQ5QeW3lJDiHW6F33Eq/xHSg+bVPTmyUfWRTrz
x62+j8EQ7Dn/v9Wq8b/Biae7G+R/45ohWfyKPuJLXLf6wkhmy3O08Jb1+uSAe8K/
xd0RK0oWW1in2udy8hofCnk3B8yWGR39ZYgKOkcoj6eOi7k14YAKThR6lUilkLoY
Yoky9RQCS1whA2zhjLrA4ioPmGaA4hwkCC4pZKC4h0PlPyK6VsG0N0eFXTyYjzF0
dbQ91SGSqUUwI9KI0L0TchAW9DgyVnD/HOiEQgRDDYV5gJdDFICRapQHzl/RiL6m
dQ4AhA3RDd50VKhQRYHL0mv/1eYqTV6PJIel/HHPnixwJ+HijUlv83bOKjP5kSsa
zAOLYKZz3cql7ee3+hzAYkfw5tT8Dsn2doo2YqrB9sMGt4zqua/3YDVkJ/hlDyBO
rGV+ltzAJerEGRecbEyQ2dKaXsYutE5wP+DBU5ty2T6RWKR0BXUuk5Dzbcqj9pa1
YrGXA2ZTmbI7yRiiGiygyW50Mk2HhkuFqW6UNqLHkz0e7OeDlIQFyv9p3+x5xPnT
Cbd9TuDyGt3iqm3h9mEFggUdZ1dXgrZkYVjkJC61gXU=
`protect END_PROTECTED
