`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Sj1ejXdK7bPsrQMY56khsLUJTPqcZxeREM9CZbcfzzFOYz5YALRy2EtC7FKvhSOx
BcQRMmUTzDp2iniy5t0QB4lqyfP2taJwqLfGJ0vF5EwxpwmrCfHvt3Elx3pBe+DA
S59OjYTtp00uPdi6TDe2Ib1pREni38Bv8gfd1+Ye6LpHEHmMmi2tiq0o8I71NkT2
bmV2jySS9lp0RJ/ft9ObJ6bUPCx+XLHky7AqO6P/NLcaS20YDnHWGyq9aHqGxCSJ
z6Zgv8InYXuryvbSNfY9KS1imvNKaVtP4xXmStxRdVtpLYpplnmTf5JzHdlLO11y
qSlzqf6K7GTHoz7XZTIsr3xZ1lth4qUMghtJvRZyuro08URwsVl+11xIwg09LDMC
QoqGEfuyNNs/HO93+2lJ16PXiMjEQ3SJOArwpji7U9YzwFOD1IbUrwyPT8JJIPt9
BHMZlLRh3NpEGmb9qbuXLDj8NVJxHXmS2aWwPzcri1zlj7ogztomV++IkA9nJslu
zbUCE1zpTq+pf5649i1Nl92N6mEGDPT4RCPr888MxamMeb9hAn72PMXuXghJhlnm
Vj7mDRCVmE6AvL8QJEmfGuIz3yeVC16uJGWDQ9iWFyA4Ot23BJzs+OtyTWy9V4aR
FDlCQTQQp1wjpbdggnhoIQNyW//EL1oD6vq5gScZ+KbCR8JooNKztvUX84vRuOzy
jrvrNBTgek6bjbYSVGI+AtvXts249W3EQ07dEwBKMZX/kz73E6kGVYDevddgVQV3
JuRbDe5stMd2GbZ08l5UajDf3hQCKTqhkbTO96SeXbJfAPyuRLw2WcJ3mwvTStRH
kkHhPnuggm2jD/4zBiejDornV94eakVZ7GPv7fHEzx0Jhtjkp7wHPkVQdKXhxy4Y
xMZCnd2dtkoUvbPPpNAKADRFiZ1lza0budyAcip9AgLOQtAT5/n8PoJ4lumO3YCR
SNg4VPbL8UYlVrAXZ3Fybqw6CHcHgzDZ1f+7elkUp1vYlZlejrx3QflFUED98wY/
GQY9O+SK3DApp1X4dFOATsDZt5yq8UYFc9SaGP7/xMS0Gx2n51A9lc8I/aCWSDfF
FtzeoJZS0A/uyPo0RJ5RBGSl7kTVTivmGSP6Ow/Z+EQiqAB8AX2ox02js/eFLnyE
JFi5PDXcGs8RQXBNuZKpyBTb9U94xNBEUsEiNvWI3Khag+w4vFqBZxWaL5oSmmf9
W+tb8y5vS7hvbWyFZUNTQphH+XDxKy2UqCXMspabq0uLyMe4aG0shWe0CfcymnFw
jPvbbKLYvibI4UU0WBdUMTp6n+4EbpVHPxfB9kb93rq+YVJNpU4m0PKp7oMHRuWW
Yj/79bD8b5eVBnK8BujKpcgpZfVbUX9B5xzTzzlbqEJtwmJbGndsbzLlqeSRUkIa
8q82okyGz5JNLOZJ0UaNfe9Pu8rbSfpufX517m/JQIvpBe5HWbIJdfEKj4iEZSAy
pVSwCc0/uAimu6lm4jiX2vR+/lSjsJoM8faeAo/ZPS3C5XNxKwPnOjWglwaSmKd/
mAwTNefICBPjLx34lAciJySu2qnnTM1GytYV7Ogl88BHhN3+vqs/Tis+1YCQAEqK
IUgnJpBxawUXm2rgHQOOKikGkSxHTXG2ROO4/kizEQnfdDBqtTrZ5PjgQx9I+t6w
`protect END_PROTECTED
