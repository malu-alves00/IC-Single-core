`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kAci4ArnFcZmuDUJHC1whyVW1/Qa19wc0rhztRqBXjFpneGH0cHx+lkCBj0RzgO4
EeDjkV9J68bag+PlOoFEfotqzfDun+eFtJXAn99kzlRPmiImRYpsKoNIQpWqXrul
+AQ47liQ3eVUWf+th6N1wHuVUq930x7vylyIMJ3fg4rzwqdMtNDDcxdyJzQj1qLz
m1bolHFXyFbb1AOgteaHK8FMTwvDhiFMmU47feoXfMu7blBrzVuartMRi5KhS/1z
oG4yGkgGvM54PPbJ1u7Pjx9SxW9k8hMLK9Xq2PVSKXVB4KbyWbYgTtwsmgKP98a5
mwer6URVbAtN9E22ZwYr+3C1VOWx2h8nTTtiMGQsnSlqb9Ucf55T3qeE3bvnLfCW
aiLOn0QnkqIH4WpxSxM+Jguphq2Uv6a42V+Nrh58r/IB71p+ADytFwYY8ea+gbuq
ZEifGtmncoTSes+1A+5zXBHC6XFCqXJLZmzZkCEnOZ5lbTRFDdspyfP+nw8yo9T3
4eju3T+eTWkUbdmGPZuy1GJ1+ae9Sqhkm+wQKAHH+c7Q1xVerjLaG1GAfdoWfeup
hLKi4PMBVlmQ3ehQms0rCxk1usPzWfIfFt1D/XLh6nTAC/CZBii0mCxSEeut74wR
kgk5cEO9yN/N8FvVrDNZlHiah5o0mExZ1Qymr3R+vK4pogkF5onCKPOX7L7OfSrN
edSHbe9OFFWzII9THxbK+sPMY5gD/oHw7ADkhEPkS7K+6srJ5Jc/QRpUKEbpszAG
d+1yzlYBRgIR3ibK3O8ex7UD7LjDd+uqFXRURDJRkXjJYT/tTHjPcXeiIcCaR6+q
jD5aAI8kqQtkgEba0VsEFFGTGxC/Bj20fAUyZteJA6pfDrwiVQASCnJiASvc83ds
v/yXe79Au5W1aGl2n2RX1fSS7YTS0PfdSHu3aupnyGf3aZDV/+3SUwxqkD5qftN4
g6rKbVOgcIe1Clw9tlkr0A+MwWM5eiOFnzVGhKp0PiSGkxa4ehoiAU/3OhDIG/Sh
WAbcFdCsCusQt0xOz3NrmbdSmSoKX+H2rgfiPuhT05mgpUuwWP8Ijd+VbQeZoH++
3LM9b1h9pMCYWqG5T3HVAmRZC93CHvSn55G4LiujiHV/itHeYx07XlxfaKDt4KMx
91SjuDHJ5jMHBAkdlO3b54ldR80S2r94qaSHzNBFymbmDUuSpgDJQPPpio5UeNfl
ecJ3V1TNXaERQ4FxftyV5FgREtE0Sj+vjd8Y9BdLQBT5zfdm6aChxV/+KEINZUgp
9x8Hr2er61jL7KA8VfKd3rwugFKvFQpIqP06Ep/X4VXFZH2CpcjOE1t4gYXiA0+W
WX2vZwLsBzu7Va2pw+MDQZocOIO8M+p3MkoMiLUjsROgktQLTtZifUohFv1jBKqK
sv4XGk2O7UZC8ScO3TU4fhRr9RMYnfODgPkFXN2IwG2eb14oV693JFZCRMr4WK7m
GlqnL9Jy1dHFTYbr93zDKaD9zndEWo8JUBPPqq2dkCcSnw3NifjonWBirD+sL4uO
8WjEPmFiZ8aeag+kearXpzGg/b5g3J0tBcO63v3ZGr5fVgfBlQrZNR9ub/GHXxen
zsvcp64mPWhvGIvjkcN8+0mLPpXpMsuIeu6faVIE6WC00k6zfXgU+IbJ1a6IidRX
G0g/FOFWewS8ItqTKw4tQJJTxQsPfDenLyRzgFbM8KcD18VYkeOrq6XHvEqs0ZH7
Nd1GOS5cmPzhhbOs+z4OKATDDiQZM0n5IefCHB973iWd59h0IDluRheHDCFmPOgz
pyOGdEWn5/XdXUVYvnL+RG4mNyWkMgiDDMHcyuqozT/+UQTQJDlIn9/UFpI6hxER
DR1VXSrF+ZuPAGlmFE0mWKY9MwVkR041u/st6hu4/v1BIWhCvNx4Clx5y6fb1lcz
s45IvbEgvNxm07gUjVGD7WYWc2VOPG+54vuGeYxA/dIZSrGt3pSX7iMO2iB9g2Dl
Tk8SvMtQ3kAMWxy0rBIFrhI7lidRweEYK/awR0VsGco3EYJw4syOlnwRm6UNMq5W
o7WrHDJxgncMplLlvMquyai0cYytcdqpBggrQRXLnUVuTY+X+IFZhxXTTBQIztx8
Q9cVTEKUPYftJTBF6YuIRipfHVJydxP+hqgYRmRBOiYxbkP2+xR4sT8fGFOUPtTn
702+e9NpWc0K6FmqvGRvUj+K7m05riZ/yGNS7AkbylBOH4MxQaN2AeTxUgXofMur
yUmkYcHnp1cyda+RyIm7z7BarLr26LQa9kNeQ63+kxOx/OCJxnb4Y4r35Sn/R1Cb
qAoF+QK2rG/no2MwLQcvNTeb9SOfApmHAomrVH9X7YyokAQu0JJUP4oiUvziVNbF
Wl3py/Mga5Qb47QDr4saGw+K15YE5qeqI7e0Qrhfgmt1FPBdlB3uALukaSFjlMjF
BupCJ0Z+ks2pQqSvTSLlEZu84cF888AYcS76xXceO3h+jTEF5Navqwj6aEdME1kl
C0iUYuuCtg2N7+qyGsRF7jhwvKxXGSRkHhC2NNmQ6MLo5fWDbUQ8JbY0gBYPhom1
Xo9xblhfUOJZoTdS28ib55sKpQSqQYYmVkGUCoSXn/UN3hUOaoKDm7ZXxfFEBKq7
/hz618HSxXV/TQi76tt+TXv46lp9Bud4BgkAX+YZ7HZUMmuvzWp3Jibjy2EcvCDX
1/aND1BPA0NB5FGObivsxsMUrObYPInj3OxBmYHHJNArkFcOLV5G8aAJ1zWDHO3w
RpC8u5BF4f2wtP3dToP0/0hoExxHNa+jbROYzeAtDKbF3ClD1fI+Zvc4/aqKTvfs
7fLyy5V71Pz/De1iQEtwllcEukeWe7p01Zb/nn6hH62OW7xcaCvVInrGxV/LXlyW
lkfCZJM4jRwyDAMuASsgm1W+U8Cdit+HItU2oEVj4kHfVP5jF/pZjkafnhg2Y03z
P2mFbs+AuT5JivKDTSA86SS1uvv8pwuInqYxYM3GbgRsUaMxS5VMsmyRfnJP8Frj
L/UAfGnLemqjjuEZdRizmxQ/HDoeiCjT1VeRQ1C9Ogo5ynYHr9Nuk3hycCyv9840
oMhPBVNm1O17zxv5Ol6g9XN5Pt3t9I86P0wSI56uhmVx8zbVwYelBztXKVvro+zP
BTHfSqHAndMcIUQ+EfC50Qtg0d98X4/g6/2ZlktbrKfklXedrSZ1gv2Uw33jKXmm
zA2KvESN5GIuGZ/WtCNHuRcA7GvzTc9meNuYOsck3s587pZe9mcAXyWgww0FwFMm
ISbFsKedUXCsHcoiTA1g9Do7G5b0n/+3c3Z4SZ0tGbHVbcQg+10ai3uewffjySQ3
sle6HjzUa61JM+/7TGiGU2JfN2OJTmQJcliQHyy/KFNUZJOG+hx1BQpewP1EQO55
O86QSOHZen7IsbDLaP2n9UHM7z4MeHwbW8gf2M/+FvUNaGmW/gW4yU1TEhHAr3Kh
nabSLVwqMoVx3dRK2DleAzuaRAYbsnqTGuX3Q3NQyaCno2FVqadw1xpH1uU7iPsV
izPal5KieT8JUzlyKoDgSNy5ckReh13h+T7jHM3UFXsHnssF/3CVb3MeLHENYq4I
/7B0MIJ05rHZHaXnGV8e3ZB95NY28R1JOZMDz1muJBlBtTPV3aPFYBH6/ibaxqhl
S5jbItG8EH2FckQANYbDvnyXGIl8fH10mSj5RWGYm0Fxx+DgduH0kUuX4UkNumeL
x976Asn+kOldEH7WQQJfPPgnx6Tg5wjasy9Pz3cBSYNchHPo3iR9uBf+ZnEpIMfp
vVkJUbhqsOV0rsp/FH+lTCxYqKZ8xAAOzibqUyiwiJE4n5zzrC73eBjN2rwTHSvo
0Zk1JI16MhJFG7iV7w1utWsTMVBZwyF9ZZMXhExgkXx7+oSHjOkTWGeKTI6vJdR2
7L5VvWrEN630CwmuCVS0+r9KLGl8WuSNGDvWKzTmf+/siIiUXz/jlN80sTEPF3bG
FgVnONcfy5cxSSxLutMWNgOIs2zWwoBInFjQmEhcBl8OexVl0ut1ulgZ0qsjbYAF
/vrqD0ZU+vHQ5mIHr7zff2nqzgKsZilhxfNT/UKZXbXmyzcWOpRCukpYY0OeKe5W
`protect END_PROTECTED
