`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sEzPxJqXo1u45ZSP/4BRyIR4oElUmZnPiYmU7VNMisgbMAsffY4t6XJ6TSRSG9w0
QRpMLrrRwEX9uKKFdL/2P+DBVZ0EMUXAaKIFX9lZ96ySkRmm+iBJgnhL+BFir6DK
hYYhML1oaeQlQNumzlG83wSkI+c6BjlL3IfE9vRXMeTgwb8bBQN2nPqIeokQoTNV
ZaUetLC7fg7g3vMOHCIiiwdPUfFqaUebJB26xztRjvBtveQ3R3P0TOMKFzJDeX1W
lIr4DmrIjnRQBEz+eT8PgEDODfJ+mjksJZHpAS8UJvIFFhVxIIXhESoeIW2oULeQ
XsdGtjBGPlLDU/1tPlG5wQsGNqsrlTPCn3EvbW8PfoqOGD5JRTctM98ui4NYFLKs
+rnQ7kpOGm1LizR45/3UamY2Wj9AF2p1nMx9rV4kr4Ym2uUwVBZzoDZ/hAItRD6r
4rBBZAC+Psz83Xtw/yCLvopsOyAGCiRES1cyXFlgU98muXsEye2qRkYnxGyY4Lpk
lGAVdQ2+5vEJTii3SKQYP4ruxdmj8zCOWlZ2J4vHE05OnSj4TEtfs+3CiWX1u7l6
no+s43LbOuql/8TkhwvWa2/RjAnmk9aBWehCDIc5e5uX7uWW7DevChVl5T4lO9cR
sIb6S25TGrTiLCQ5MkD5JjsTD1+KS/ClbEElkWrkBhbeBw12Z4XMWbLWAJL8/1eS
9Ax8lThOa09wwC4s3iOr7ZO3yiDPR7vTV2kW3aJ5RGaYtJpGTFkdX0JlEtRcrxep
f2Jwox6pACEm3xURP4ylrCceuL2Cssh8qpsIiXA1xhANEihD3fJa1ccnGkJLeEAB
WjXYodwEFm1cNTurmr0oqCyF+W8LQNV0NQR5m+jSADp5MRJdxba4P+xjn+LG4zW8
UOPONimEsJBdbwbUPHksU5vOPzh8bIxqj+jUQ93VvR03v19CpPgXjvk4cV51DjSr
qKZ/XZyWQr3LY5jrERdMf+6OK3QfzC/kRixDkeI0jtZIKOFs5KyVIcqzVr6vnOBj
apaziqQqeLDCv4Eok+KqtJITtxWqVslAUVVhWtESI6X0IOgO5RtjoW+3OJJWQUJA
qd0I1sNCrikLnNZstMwuwjBVnnXCzLKBl5b0gs9gwMrNEqjFzc6tHmqnVLj9fqSn
j/SLN9fJ+PCyiHO49z3ZjNqhPL5oX072X0Hn6+11DX1BWnmmorvycRJ4HjYO0Nqp
ANmmc5qvdZA2nDhEGtiJdJjOowVCBiPdWNRlVk0N40AyjVXBZtIYw2FdeUYpbZWk
EAeReMRCLNdwV08hp+d0c5z5u9Crjzlk7dpvhWT9jbFwZ0oBDaSS10Ubh5Ge+0r1
cXT2MzKb65kIUlp3Gs9ons3eSsOsdFs4Hee8sgByODC71v/7K7yGVqIqB8u1rrh1
x1pPozi9o3vx4ck0e//ATSQ50T4tewFQ7dp/j0lu4ch7Y52RQvN9o5at1TGYO08B
NbTXRwjPLRib9gtxXt3R+TQrv1gy6uoiHDUfWrLnfSSdOmV7ixsy+9/PvvRA3F5q
X5W7elt98Yh3Qqq0KiTf+zXtznnltRnIJeE8pq8KARO7CsP4F2Zrk7L+vkOZDnm9
n0+6SfkcQEOVtV/N+W/7eVqPDLmyYCp92qR13hs2qPsBJKMhRRmKEEv84sNbMpAj
IgU7fZqXDVcCEZx5K6azaWiaI9hLOwOzAQUMoWx5jD7rXbumoFyu3ETRqJhyuBj2
nuYjB7/FCnhPkj7AgwJj2ew+LbChd+V+OZSQLa7M0J6q5RdRMmKnca7ZbyVS2i1X
8ydd+zb03MIJTQc50coRA33IUIMwgQiIaWxD3IF+LgZf5Sh1LSgO08hnMFPS1T9h
ArRcFwhk1FY5K+gu12qnZyhho7kkt7lA53UrRiolx7I0yjUafhMa9vKJ2GMHRbTu
tjaKaSrE2ZQNUEpDVScwbHJbHQiEgLemdQDEP78f9PRypQ3ELtovNV0GPscJJgvE
a66CnFtb4RIFkIA6I7SjH3QMhfOwRCD8MSh3+PHLqzLJYe9ZzOdUhyV231mlNgSX
f2Jd7TkLiWxdFnmxM/AYUqLLv6TJcl8N9vQMMyYTCoy+TPvBw27LaDjieCOa0YRh
gus/lC20Vp9vsaT+R+HW4F6VpDVchFFCjkm87iMMyt2NMvfW5Jfal9/R6pKaryNa
gGDEbVlnNbP/0m2rOPZx4GmYwocLqo8FrCR5sWHqUjCFBdmZyiGo/Dx0fg+6/0R0
0xC4DwDpNkSnnlDMHd5EILs97aoGtY4G8hyTV6C7gG9y+0rqgJSf8sb6bSA8lxt2
fhMASsbkpgezD+Ur7sEdhuy5qzprcL9gxze3AxUlTKZN+ZyOSgRaYmGkyVqr7Kor
RHvBCwMmCAYvZgqnjhbSjf2o9yelXLAdWmmy5sHfJ2CniK8otSKTa9r0pGJIfxCx
G/8glqeBzDnnSWjTrE4qbij+0+RCHK84f0RCKZ7JARC1Ht52T310Y0JAV+8aYcxU
wx+hqmloCHRXjaodce3gDdgxCvw/bQzTQcDWMHfjOBbFbvVW8LTDSfup6PcoJGpi
a/cL/p9hu5GoTJxJxgfaRH8SSdZcyka1ejHSm/DNo7v6XPWbwbVtCv2IIzuGxaUf
nAOQTkGmuDylteVEHahBoOpsyGSDuj/4J/EI8yFZfzEvIvyqmRRFoc7ImP7CPSnQ
gWS+zKFNj1WRSFc3AjmuoBrSfAF1leBkYz2KOMMSkbQqkTtCDBEby6N6JcMTLApL
QO5ec0kUtXxp79XkKb7fTPZMnJV27flrq+vOQrLwABf44n0kp+gRrbTHXav37ghG
pr++lFkwlCZu0hNtGyWTATHNjFGNS4JtNW1cgmWH0/UFJlgzUutq3Ag+pMAvfj7d
JahoroO88/9bK9MMyvdC587G3a1oE9x37EE4fBooPkIZ60nAuap1m687IDDrvJY8
qTobN/DcHteSqMbVkqkxWKF216ldbzNYBjoss7i4ycJdfKoZCZPTL64WM4q3lWdL
OuSOOFyZh1IOlfKp4hJGH4nqxe6i9cQdGDBkGN0F4AScs7uyJcSclCPlyfdkrFKc
6n9x0oTEd/ChzlcQkCpViV2O0vlCeT51vO+j5k0CmWFQ4yaJdpazop9eU2qefM9W
yLmWVjn0MH/stLVyFUs5s/6R2a/2uqtV9Lt3eNc1DKvr3pLDyWYV2dWmOG07G/7A
/jfVxjNUUcwqilEsH4CvVFMxOOhNBwEpnB4E5k4XIDVl2kZiIXpUfIRrmnq6ohxr
J7zYxVdbY7rSsLpTb2jXgE1xpnS4Ne6kA4wW7zhNHDZDL5kGiKTusNxvbRBUFflU
UxUuRK9u9EXYtIWPnssV60qIjQUtedyswe9mwV056OGNVxgCSCNHOmSDjDxC/PJf
W4Rb+vKlC/9jwPtvcNBv7BR6L6hPFFEprx+VI1ydmS+0tJtq1+IBsSmQ5Qv9zF2Z
FCPQjYwC/dXlNDyVTozvbwa55pYNGO/9RNHbkG2ZDKpwpe6SIFmiEGINtc4YVkyg
nEDnepPQxLkjMqdyWkqC5ceNi2789bpkvObLsShO6LayXwV4G+WeO1DsGv42ASva
zPmcQPdQkwl/94IFvhhFRPu6cpklKfydXQ7jktxr440LN97sb/hrytNN6E5gd5v7
MsIjL4GnG6Yx3KT+k51vXBV9HhMZbCWOxacBG+ppUtu3ShiFprWwIuM+brZn0Bgp
jBBE2KxommiKUqWIyMblJqGoyDsgQ2gr8H7HHX40dV1mRbGLAvH2gX6Cpxg7bWzx
H+Qq6xIKD9hteFfEq07e1sy0LERTQFvhYH09inC3cG52lXVgvhQWzS6rdeeFPH6V
4PJNdngjnioxtEqLKx5ThRWK9sGxL4m5OmsjExQZhhXtJt225uV6L5yIrrJN5MNh
+JOb1vKEY1rAn+sRzIKq3zqxDd67nEZA3HBuYpk46DmdKkVux8kbXvOV4kY4NUnE
mH1a/4bPB2Wm0au2eRKaNgUopQZYyHHPL8VZI3YsXOzL3onRIw/lS3RwzTdQuMv+
pRxyiHUTMM6MyIZBG2MLMdSKBgPNd4F9Fo/qp7B/OBprrVGOMFd+Cgwtz7WT1RXO
3xT0btIjXDfQm3oKSNqp/GGBCOyRBtc56yCjQ1O4DjilXWvxzl4iMuX9g6r8gX1s
gG69q6ANS2DjewBuGG3jHgApw6/9cZtnxFyIroamJO/1p0SLY1Huuyriko76KTL2
0DIICyXp6bEgmEW8mbzPgXDHGXdkO0FAc6k4Iy4C/GHqfbBMMaqtDIzoZ6JLW9Tw
3qLhdf90/gIFBL+Ad7ZBKbbWBdIQgp7luCplT+wRVcfHX+0GPs+JTUayRy709IzV
EvIHVHhBrxieCFGojayW7oy8+5xbxFEjXk+F4LlXKOf8CH8m2xUICgi2fPyNSTuk
OMzBA8EPaFkJqecFcRN9SkJQlWsF7cxxfqSrSnCpJCwq6EqDaXqS8cyI7fX7Itki
yGZpFlv7oJZmx+1RtVxkCVyfT0ZiSnjROfd3ZAhZ6g8/FEjSgdAzb+U6CiZbpSpL
AjqEz8c7+xuhVNolu+Fsv6prw4QzoY/SYw0XPcVyHogGa2GN5OQBBN0toF2nsSRu
r74D/qiceTzKiTufN73evCD0zEa1aULMeFYpLC8a3OEA+tADkByBYQl7vlFbVM/B
ZO/NeyNj2SbPGtiyxYRuVFy3Q2jYUtV3bkTjVau4KbrgTK9yAi0oBM6uBPAtAn1c
K5rqgCG6X0aUZf3Og9k2MB2hvdE6Uawahf8SzZidXcWu/M48KJd9qgdpOeknxIio
rH+J8MEfBqSff9MyIyPM+R+IqjIPF2UT7OXLKgW3LlYrvoqebeaBxy6Tk1wkU20X
unT7fZ4R8aKMCfO/gfohhWwyRythCTI7unC661AvhTrAWaAUssm4/LCltDlpY73K
VB0QQV0ggYG1exLV99gzhVwcURxVw6hvQUHhWJuoUlr9zC/VHH/D7UvIB1D3mXXa
IpEi49wD5rdXWf3WI02PENmdIhLRSD6jmjemS2wE4HALBydY/ybRhGZdGt4kPc+P
idDlvY0oPO4MK7JpWribSxLPy0ZNi6TVfCSYOGfQenC8e/SspcKb+LjY5EyGdhTF
1ya3T12HRHXjjL/2Fta/ukLcUc+M/XqMyidbIwbEYCqLJO0eMA3tCOUmprutK/s4
xkosnKy8bNB7nBpFCsR9g3UbLgALeGoPd1uXxZftTuLKrV1pCYA7gkrdDPaPpM+p
W3C97SiC1Tt00fziETmT0zLofGWlesV3obrQzaYETeTzY/1gQz/a/5jJ5K+IOgS+
zc+GwdGHAOTg/0jJtT2KEPflhv21NgRrhMGmLMHVxj2gdstvbezMvXnwqRAteYiP
5X/fCsuNCxYuBPA6wPTbkynJPHxsKSdatCU6yGzXxCZwLBiuz3EQmVy/kOW8SylV
gupkCQ+fxwZKtmY7b5kCyuij/3xdUW+KrnHeS9b7DSVZbJnymPO9D4+zdteSt1vF
484jHPSa98iyF/81zhZe5uCDiUzyK6HlnRs5tt3903SCaRJLWFxPzi1YP+PWxs86
aZrana9bt9QMs3Mf5nd3IQphaObbDgMeQ/q7kadE1rymk30+SPSXX5Vz4N9uGNFq
EAoTU76UQUf7DLoPSyZ9b0/UYEBGHmJGV+F68nb7TB3QAH5PYeLd53qjTIYyFQlv
t5Sh3i0UwN+ZD8XxD5iHvDfLHLCHOjMVaWiAwFwD3Z4oIALL08tR8dDBdM8079OX
qYltj6S9MnyL3YNagZ1gdQ2GZj17/vRHemrlFkHX+rUPwf3gvxiHNT76zppqkna4
mDFQVfxWC/llZiN79cjjadVBKf3LmNocAOeXdI4sJKhhn/kLj17BJKuMehutF3ro
WghjymO/fXdLP8gJLjo1hGJaTAszNuwmSf1jAOm4oHiJw0WBLfctMQgDcvkEavGV
13oBsgic4K511fy+L6m/rKSjL5X1xoQqci87PVfNJvgucWmdN/ljqiUvQosW0KtP
spQR8DcgqM/2DBfnixbAZoqQZqI96ucRIfHx1Bs+4Rs7lZk6ZUgh7h3w44MU9QFh
BjFDyFzfRPsEiveU2AhNU+cgHzGHk9OJCX537nHW7JZdtRsor5y2MYiODIFL8vsQ
/oH8FLOLUvaimnKy9vixXhelP0331DlHRF9fIm6iQ0O08Lll1LF6cM+wMJcYjJlt
0+zNMqle0wLwyStJwbJ1exj6L7CQi8lx772LhMw8VTpJ3nps2kfmNNmZ7eEozp7d
iiyjI2F88GrK7GNUOS0uC/j/jXXEsG64izjniSuk6GPx0rwj5UbXOo/sQWuT/ZhQ
c/L3FCU9M/RB+OTHZAfhL2jVoq+SCtMbzbpOjPNRBEqzBgPfqcqPeMMy+Xdq743t
/8fAFeQ9fo4mT8HRXTJgiZ8sLW3OGX+QNE4ZHKcfZqyF3kBEYXEQ/VCTECzpNkb2
gobEwX8UT5glPDNCjTYVm5KrUr5eGX916KA1tSZ+Oxgd5Bowb7YQ2V+1r0u77qIe
6RVejg/Bd13Jwq/sWC4G46LVSGJL2T3P7qSOSCmxLJbijEmrxIz9qh4LXpCRYbAe
P3Hj6W1d+QnN9T5/2AkrMdcndrley/l+vQ3mTP1UlNSkILPwZMVglWAgzqa7c/Ia
5VvWKnqgIuFsf7SiToF1tp7Sfu/+Kh72BXV2Mg2x3Acu+GgTyslmYf0cx+9um+8Q
OcRJVxjQg/QHed1Pr41NDJWaGt9Qt8ThTdyfWcCSpRKTR8EC84wXvwb4g+fKVSoi
h/GXwrIEjzmoE88oHLG+rpHSPAUKYPytcPwUU6AfR6HfHAYl4/5w6FGydvOYf7pS
3tFGfmzKKUaMTv3LkPITbAb6spfkRadprtL2q5V/+quuTx8W56kDZIr4FeVNIx9r
yH3il32NqjyoXipROrInkKqadHdlfmtIEHt8Xt9vwH2xykcZygY3Vza1Toh1Qtx1
XceU9S/bT0pb/6CljPm2UGylWK9C63slJSwqIGTa2D38ydY7rD2akVRTy/p41LUT
7UiahSwS+1m0HQXcPsTAxDVRF6j3w7KRuv8yMjr6xFJak6Wf5LOwGlUPge2sRUdN
6f9eoDNgjgFQXtCV3yTqjh6fVZJt+TiUg8B/FqFYRL1yRJG2wiOk2yMu1nvFVQHa
zvG2sRWzTcZSBBSGiigEVqzj9XuD4vALYNmzigxjE7snnrG3XseAEmiK37A4tYy+
Rxj48JidTW5k81i3D7sePk5yKNTP7sUDfBClEmBgtQCSm0A/5Jqth3F0FcUdyrn7
RLmHYAY/Yf7xd05QuDmP7YdRdEkv4MfEnGSmhakTNYQ7kIp8x8ozdD5QNL0SYdxS
vnDml9fT2jhFhUzTyS30CrXshQIdYEQxc+T5F8RrUoXUov6Ef2nvCWy4v0qvCat+
jCtg+S9bjCd4JFXXnk5/5EzUj93f2roagxs/gRB+CqEIZAFy+u5Yk4srKQ39qseH
/pRYjtqyrcDeKObdUeYROMJyC2bSHS5W+YsbP3M/IViUWuEAIkGTSj3Bbe3xbykz
6hctmOYjKueFzVIekmIjbWO8WJAJGcXlq7g/yedv8TEmG8yD4501uDYzE1UsbDwt
A1M8TRDs9k3xS1cDGDOMHBcBMKtD5CkOaqHdMh58rZZYOK4LTzHJce4Mig7cmVlJ
3/tWIo839NDRGO2SB3oJfSW/q2M9pFYDuGytUyuvRy3QY8dlKeFVXleqJk+x0FrB
IFxmPFteaR20qvs+ZfKjr3TKDbtjRfXxYVgo4ojJWubwMohVOTEys1j59a16BlRC
AMLTMOpRBo8RKZPogt2ikkPUKS8EKGg17ppbTbmh0fOYCGREgIJP2q8C3ZaaM53H
S593maQ5gFBQowFBEMVEEIP5NIc4rgCqXTh2aCqEjiK0ZPKL5+Qu8ufVF6SdZJus
9YqmZWVuXcDgsOwd1bbmwHvB78QmBtvcAoJG8eI95G8fb2VAntSuGLWwB4OpsEwN
pbnN+YcfIMmmkgDBGp0glRUlluz4RpxKnioqJ1WVlZ5JuJNS9NFKmpYasmlT2UFc
dvk2tjo8RTo9OXSfk5MTqFDjqY5i6HQK5SV834GvHnxTZ6KJjm4U2fpNS8CcV0ET
`protect END_PROTECTED
