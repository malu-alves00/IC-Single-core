`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
X1ibT/Llwp/gRaXToCVfVfVyMV7UnRJ3mVfR7zJecutFjhXIpB6pK/qWeSKg2jdI
8g/AXwgsmbOfxINDsfzfEBmOD0trdiqkBA61GG5Uv1AYT3CyPAAvc337qQeLsHZ6
XZO+N3PL+y0DOCm7IKWFQZEuDNAo1gbyJ9jIzFe4IlZ8GpGrEfrjsSAYl3KYiUqm
bAvTplcpgR5+9QokcoIn6Xk7eeXgxV+hoZLDCyipR8fEiGql9S0zhXsZ5OVojLeA
ZvsBA8X/NIJCT8GOn0MnOEKqvYGkjNDDh9sJJR5P/0XTcctK7Xk2n1GbkpHORlUq
XeXoKfZa95cIFTMWMLTBW+uWd50/SZUETtBiZCmgeDZKoVGEEOrIUsAWA14a0e/E
VJlhItMBZ1HJSyaI5DI4t//qmzQiwvZ9t5k2M01SrAVQcklxhwaetTipQ8pNkIQV
NMZ0tEZD+lOtqrv4h916LL180Pl6p5rygigGY9nFz5E3lTkTfWR9wvakWhz0f5Yo
AOpDHWGjSDaR7z3uPioMTuUSV74oIrUCpv6sBp3xQZkUHGTFc2MlKwXEaFcwwTpW
J3p4FdtUIksKUHAhKXignAmr8DWaDECR5SAFEwdyrrzdeDVlA2K9uiNgbBxEZniN
QGD/2+zElVDc0QilfLT0pw==
`protect END_PROTECTED
