`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uk+wsTdU06/SBp5Wt8RlDTxBU+4F94Wtzo48RAB3UcRPM0I3RrzUFn/fSGXmVsJj
0J6zBzqO5d1b8tZFxcnHmO3lPF/iaQ3cSUUYZ18vF68vEtbFgBDn7DLDW9R53s6C
cCHPHEqN4KByrVr/AY3H2iw48ngdFgtKn/Ha6ZBO/0Zyg6BPsEZ6z305DyTjUnsC
XD6bkgodaQ+wfye9YTq+pd3YJKQn23nYiFkILdBsLV1rkS0EVO9/tnxzflyCduV8
knGGji5NxLx+PB2e65hRuRUfbH+KPeQdZcub48FEhKh0vKSHcEyaaZ16ju4UYVU2
eQHmSh3peX0WrRrJV9lBt0bao0da+tKFaP7GFsuOIq7Ymy0BxO+JDrgOJwyuRv6A
HpF/TIZuhxlfvUFZI+ixSJFgCRwitnWLMZlSqsQR1mMNN17R1MyW6GOKPzySmkGd
v1Zn6myNB+VLb256515cO5iqYEiajJb+SM1vIZOMC1I=
`protect END_PROTECTED
