`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qZgbhiHeDbYiN/u6RCk/XfM5Bx/nLnZFbczItRServLkNqifPE/sN70JWxz5RfqY
fa1BHlzAja2s0GH5LS0b8wurLBmBTWSHDKKiA/8bdl+yWhWLUF4INBdEps/6Vzh0
FpCv2T6bo/9uCQVxF9tOyhcZlmxBYtQhzYiMFo+GRLvLkCMUFnt1MRII8AyA3uqH
liReedAphXdioJO4dC+Nyy9N5gd5k9t/P0mUoNpbEsfJuTJFnewW0xaRvESmGoPC
ltEHUeFqrlZFGKdxMlZqFIqHthy2gXJ51QeIZDFy9cx9Cgrx89OpUvVhqT43QNmC
ypd8AVclNUsv4oDKl3KGAuSeT1flfBaajMdYZB+KowsCNmxVyFA9NL5DnnozcpC/
OvTOFCXSUJ+yI/OcbO2LfA9+GkqFZEN1nlW0zLUyAjKBsDCTfFT9KzDoZnFZSRGm
TyzBJlZAckWDv1TvUSldKsReH3NIQP2Bn4W2QqXfbNFsHfT7L843ZPyNnm3KjfSU
hCO8f2IuJ5HeXRwTB+o6PM0TlqwJ3aRH1wXv+fVF1bJAI1t6CkmuY4h3RJCMkzTQ
cQlzTg0vjPE7C1rxDsSy/i7ununruaZFpeiC5GjlmuI0O2/Bfh/YbQ40kVgZEMAu
`protect END_PROTECTED
