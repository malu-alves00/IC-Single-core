`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1RwussHFDyUBOFLsjGjkE6Ngj1MHbwIBUWc50WdLyoOSjSswoSunWLh+RoDSgInr
m2aU8FozR5udqxoW2x1rfq7AdSKUcVlGlUvnNr2+N0THAXnxpevpBQ8QyRXJacVz
OynpJxextpz7YarJ8hznh2hfx/4tGPJ2gfCNtvJn9thGAMv4undfqIzXoFngpRny
RVOTs4XlHU8FylGDTeynAxZsIZlW+r0tvKAYpc3BdiKhUALyy/T0AzpYRyQwVuqS
IyIFEP0baOqGaRtQpQS3Cnf+pjuVhQpSoGpkkh9AsyTKz9UdDklaXhqhu9E77X0S
scf2m1kpsM9m6g1TjJs/icC1OCxgTLYsqLlnx7sLqDLyX3NwmsNsAJ52+pJvA4vn
hKhCY9+/NUFMUfaJeuDQ2/5ovskoTIAltOXinH7MnUp4hUJaB6Xp2bXMpCHhRwpJ
qI6yCYZEPaXeUWeF5hHJLg==
`protect END_PROTECTED
