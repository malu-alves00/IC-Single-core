`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ejvLnVNyW/AeOunF/d4cRbhEsdmynh7aQLkg7kDWx4DWBDZxtjqD6F4pTDN0m9/r
jGP+5um1J8KVJxx3nGtsbmtdpBjsLdFbF6Qv0DPfmHERpUZGYEl1NsjkUBEDZhiZ
9tXK+rG3hWabprK8ag6LwrbUj7PMKzUZwmqjQMZn9w6yorcMTN2z8wgiGtypyZ8s
hxFsgogFrgxSNnQ0aj1MlQ+QmV3M3aIHZFl1k6H66XP5omwLECGVOisVAyMmYsFm
yGuy1ypumMVQ8/r9gmHvdam6Z+m954sBNuerf4ERBNg6EDSInV8o2o+mzhJ6vWEQ
K2UWu8czjjlv1ZZfjITExta9F7cDM/cdpCO6rDm53QgW0bCDfeZqmu7tY5qDwVoU
UkQoCv25V4Wf+n+drWDQga82rMer90SuJe39bZ7qI8NdRvbQtVoYzpPsjrUkPksR
CKQdjkeXA++IFYzDfy09rgdIxcfhQ9k+BLHrw8gzq8MyjtmmTBEWe6eDwnQQAeUO
4pG3ybZVxTHYrsYuaSWzr4lSBE0TU+40KNe4/Txins9kUEq+R+8KZFn/krepygIh
GrrXFtsgrQ/UaZWS1stTN4glT+m4K0UCXwIRGUv6vAab14mE7bAfTRfYRM/bsn5I
EvWKSIJQwydIf5obtHC/osdZm9uQ7kMV+dQZmQcb8gR0OpaqmW98JawlbEzDIwV5
OXlnuU9B/8bjcc4zJQ1r0VyO3pff+rGMCizAWnqOCpzYQu2dpaLfIUQg96Hz7NLZ
z7xgvFalmHtBUUtSgjP1fkhaVYNRP4fBC4lgS6u3yK86I6l2EfEJql6EDlJOpy9K
pOjSXSQJIbg+ib6F2gOhhuGmI1d/6tCaRu5eyLqkbnzNA8n3FRZ6HHSyHi96YoqQ
Z7KDCwgcHCQGPxF3dtVH9IHodGRrCmKayyYe2k8rZa0RY7Ve3jkPLfkpNG6gfn3P
Vu9VYzHfGQ8eFjtBDiEh010860kuas6hznyUJ4XO1ZciXBsrq94FW0TQEaydXWgG
G/JAmsI1w2/TBqFDQH/TYtNfQtuJjO2YVGj61vMHGUOntCtor2/ayfMF9+QoFjhz
tajjeGaaA0/8JurAgtX8mthpY79yUH3Qth4hDz55dRr7VK/37l3SWUuOCoc4u4Fv
I4369AHJvb6FboMVVMheuNs4GBKEd+3zGxZXimyaiFcJnLuq8FxeiaZEZsdpZtMK
rFumqFt2LfmNA1TPwsES0omjHGS63I6NV6sWd4AcXg2XlPtScEzO7au4PTOsjoow
dsdxcs1omwXVQfb9Xk0jTqTnUxcCiJP+EM8MmHbywD7CMhfTuBntREzBBAw4OF30
wl/g692R3QJpGxb7MaMl/A1+UEZEnj7A3Hq7uLOkiTJLrfA2Vn8t/F+CXAROB1Zr
WXTX4QuE5wX2HqYbLrRmgDRF4bVxLupHKzUHjCjuoBLrrhp1FRDb7XLobIB66YmF
nug2xgR8pfPsW8mmDPDPS3l5lJYcAD8oJC0BqE4EjokqqMXpcCTrtIMwkV68RHRO
/bE2d/n/0YC970vfs9DXZ53ScS16llKaHWGtGfu0OoIOi9v2hmNysOxLds0VAkEp
EXwdD3lfv4dj1bRCyvJQ0XH0aTkyidrhVeH8p3VD2EVJn+iy9j2fwszwcvYExLgQ
8Ajb9xT0m0gi6/il00uT9ktw6jSgvb3fioBnyHh9JVOv6xWMcrYme2SH0x2bIvaE
1FmFlT9kgmuI7B17yn9rh2arFLpxUSpTNozH+/piwQ3tGaeQ9T/0Za2cWD1Byr05
CeHbNPGNsGfy0zqS+hvrdBfx43pP2J70W8iulhmaoeFTbLKCPPULenoRYaTHOFhX
gjlAEe7cInx92KREu2/tTlEn/zcEtUf2X2+fBVP4hmKAl2Y2aJb7tBlHQDiIOFTK
Z4gzaZ20yFyPW+KrX6YVxkz/MQug3jAFkP1n/Rw+V9/qltAsqGKczu4BGmJ7Tryg
Pc4lEeTG8zXXc7+qS4V28r3bK817a6R47OESAX+rwuJQpmorptX05czpNMwzQyQ1
xVPzm9DFk0oo6GXlgxo5P/gq0RyyGaUN4nZq6mi5VaWbTY6WvEd59cgGZ3NJzo8f
J6WwaEs04UgQrhBEYEbnbZ0KTjz0CAp8CCgVYG08IVPygrDPIEl6vfw2gGnq96qy
qnZDUqZAzcoLxqs9NZ/QMr7vk6B/L2BdFxzuarkqW6rIH/Uf21HDJR+nOpyyz1a2
dkhOMSHSCnCW+tVecasAvhipsyfzJB1+iZRh0uMR23YeAN73B/8RE58yXgcpjTr6
Wt3ZbwtHk8VhWW/1t1/bCr2FAvcq23LerowKUsj6YrUlFkZHk163myr/xMBteCXe
y8V17Xu+N00IaqpnOfcKHhoooBKdenPyxrPz+7c0bSLvXjRLKk+FHoICbfPCk8QN
+iBnJw2Eo2XN5sSlInxKvm9U7RTpDg6d4UGo6vFC6wHsQuhHW2GeJuoXMIgPJbde
OcQ1yh2AjNS9usDe2NCqUn10YSdjDganadgYAs0907r/8iU+g02HbwZUl2tMi5QP
JqMyw/rjqoY498jGMPtX9Uy8laHf2e67IGlYhsf037qgo4Hyv2F2QSfFgo2tPaal
ynKtVBXGlrM8eG6YmUEgjtKrfm4q4y4BH+/BXNbgYxXNtU0a4kqU1MhgrWzmOGT7
/mE3CuTQ9MNxcjFHzN5Bh731NRWcc/qHTS5HuvVL3sjm2yQz/vAZtyog0QG2wDrN
3+D6iusPozc1w8oOpc9DtLdNqwIfWYYWoNRDnPxfxJBeZXulRWh4M7KybQlkYXkX
ncx8aX36AzpEvfyTnj41QTApwZKmB5gCyWxR6A7piClR+tgZrCla1mM0Jgv1Geey
gY3mx/yWiu2vK0IK+iMCHW9vlmXDkz7vOIBDIZWYaFmNFkTL4aGsbELcjXw/Fh4j
0oz3N0jj54xihyqIk5ygVHyhwFNuRNRAc9fJkJjgymytzwfqO9K2hHsi03YZHXIX
eRTGJcoFGr1+a7ihsIfbL+v0cStUculCwCuSqcfQtdisoMXQwYiQc/ds7pGqyxOT
zgIXmnWJ+y2vMpbV6Q4yZBxL552LttejjGjgE9a9j+RRsqN26SdyqKGmcHBvf0iy
iAQCU9yzp9Hjwnrjv9Y1RAt6kMO4bUROvaOBiiPl6fEzHgAU5lWQ0bHZld9+JtFh
CEwslNWJl4+1Grdhacs5h90oQJKeFJbF0N5TqB6eN9K0YC4ZkPNW3WKw1UNUcxyJ
SyPGC0n3kFUoc6oS1JVkstAto5nf5A5lQtv81LFXF3pLUmpf9Mksw+k7pR/cRZB8
qjkFydzXXOyHHt5PGIz/cl8AajAlw8NQqe6c4BhwrK2jgpoem8TEDvjqSLkrejqG
1QIoVkynLoXDQv4Eo7Xny5ZMWgtFsNL3cXtQio+wJq9fT/rDQg1/Ru2ya/LxAJEa
mSeOZlfaMll6U2yXU0WjYqAPySq40YO0UswFJjORMsx0KZpd79MXsVTPc+kfte0O
XoEBDmgEvXhvccBH7EQ0+GgORjwbiPKrf/CSswNrhXqbn7fvhb3a3pAy4crhJ51A
cDCn2ZiYLdssYVIThEHIbHh33hDb0nZ3xjgtmDMRHR7xniCQZu+6rF365uvuFp0L
M7rDtF/s3EnRNNuVewm/MaY8vZQZSQeaxMGH3BfWJdEJC0g7jcPzY/xg8hI1hoCY
2oUkcje3QzkMas24Hix5tQUgBN5xoBNQh/ZqJc9nTyiN9M173Kvw0remV+y0apzT
5QRUGMFF9vXuxy6k7F6VbK3j9uCcCgkZJeM9GUQm4SrC6Zyh6JcJZ54Eutdg8Pkc
F3+x5D4DFFMnhxFfLRBnNFIfptxg1rBu/SQGAJP2gh7YvJtAkdeBAv9c8K65Yq5K
xWlPzdaXE4mlMCCZ8lD1dKu5aVdt0K0vWPvzmMp2FmqWdMITnMVniNQdqfS2kowu
5EdZWLZOe0Dt9Apf9jo5A8BYf+kTRnmHbXtmuJAs8edeogOBi8EjWfEmhI0Q2sZ+
v0DndL6X8LmVHIZB+NspcBnc3aM8bzOlFdsWDGAt8yF6ON7lcv08DxG4mKsm2ksA
rowLKagciqshrO0Eb+tldno70ulN++AZPjlWFiH8v2UVvrxBJEPQYmw/jnRnQhNH
/ty7T/Bi9i8n/2bKdpUqNgbsMcgzrrOB3jcrTm+CSHbHvAmxVx9l0IhpypT6Hxpk
6+mJ9pDvutRWQC5tr8x1xgeXDQuXZ2ODK7LAYhyl7Wn1kU/ZBBzsvCxyXHm7stMU
SKyxijbxOsQ8dEj5OTyF+22y4cU6flFj5X/XjGds6EKiSVVVfYoe/uSpqW3R3SNs
4UEjSJ4cGyyg6veh5vH/R+itk/872MaxnceR8c06bha/YpuQls9l+Qrtw7V4XAtX
lwr10WpE5ArLGj49pfcgVS+mmD9QoL6lqFUp4oCBQ/jF1hm+6uN27NptEIXGJiMR
PqPNIzQ8oGDpF1YO0luDj7QFAZ0DgVpxklztUI/PRPqtyG3Fee23sx6NdG2VXY6E
FYKa79jocje1LVbTbyE2/BjM8fGyPMyVsbezBMZ2IdXCibzFqVQtHnguJglQWoib
jGP0QgD5snHbKyiq+ftie1Igi35+HEDsUSXJJb9QpUTZo8Z8OkNnN3DEIjIPOyo8
VwUay0vyOfzKQKCX2JVu+OwXzxvYdQNngmTKe3PsvLanwIeNWSkiV0HbjxmkxAoW
KjgkGF961SFgwlzjrYuD2KF+H2zEno7ZVsTfQmPalbj+iA+FDLvgE3MNXqxXJjAS
ZiJbV1Oahsvz/Na2HY5uBYtrMm4PbbOyWvVScGNerHkg5doYpqNQcDU8sJasKkAL
B8kQq0HzUkhMr0pcS/1pA9nWJtEtZKJ7iXowBnh9rABlVyi3XrPtx3wct8O0tOVO
DUsQGUUzY1ac2woW3WbTya28QtP8QKsE9BiaRJOipC75NmvgTpgMlFrA+wRCB4UW
nw/oP2UTKskywZOliuT3eUQqI7/4yOPBjjr0A/w1iDdPtv6F9ihaIF5q3iuYf6up
njsETAvPEKULyefUwX0Inir+hHWFkXXBgwPoa30o+gwycQxdpBFkTnF69nnfp1mw
0r3IC28KS8xT4kvWY4SFbQ18GU62oDEkgQf7Xh/IYDZ9fUIgq6SziBCbHrhywQPU
7zqdKwpfYAI6WH760jK9TKyAVZLsh2ONY3qksiEWjalV+A6Z0WFs6s1mdRYWbIV0
unzHhEx+YZDNeDcQ5HIY6LFRuaUS4fpw7XWEvlkGHBA/qmKttIICHqeULFw5iiei
sbn5qk4Cqnb2LlnQaXsk9YW0ZDR7bkUPBL5p/PL1b5rB1Qx8zRotBpKCi9EWwg7E
sjC8NXhej+1OWxsfhNMz9L3tIUlAvu96b6P5QZRUKKIPpz1Gz+HUoZU2WhE4BYWY
1ipTDb2Zmvg5Oe41XoqeC8jf4ZZm72OPZqU05QTBG6nVbHUlevu5MmOXd8mczcRE
raosRY8xaeNViISE+AJru0YgBuZzkI46qw341cpF4aHP/Nz0CMFmYE2pHCDlNvAJ
vq4hePTdzwxCMstcrsv830JJSnlH2sK6iVxQx7qPMZ4WTbrx4IIHy448NsD4MJYj
rFgyxf0V5+3fkBRptbK/rp2BVXv45JwtZmw+A65Yd20Je6QWaGIHuWx+4Hnqzu25
p0I6jEXbLvTuNFChNl87ZBEcLdPO6F34T98kCR5xD7tILOsLI7Wox2Aev6W/tRG/
cXlIyuJD7slRVLHKRcqzleLcwgxcWJh0x6WAUv96VxGxiLFpBngUN5mqd1cYOlYW
jdgDypmZbmpTPUbHqGn/oZU5awJamt/mNsThaW488KH7Vww2NO6pXDUEHUX1foj8
5QfgyOCspyu+CyoI2oO0y1N/RzDlSwEZy4EOH2ggMfuNKJoLjrfFgR559MjAr1oJ
DAp8dDwkPHM50foA6k29Itsh0b3oryNdrXwm5TYSYHHgUO3u6DS4jAnY0VQ6dUfs
YL2LcEowLjlrffximnw3TaUFgWs4fBZHkAVZpggSsxJquAegRk75Z+4vcLIDBuFi
5bcHgCrHFDbEau2JBQtCqxaZ/odstpdBXd/FARTeCLpa3pkTDCoAP6LkoMOx9gur
Wn/YDNp9IPyO6SEm58dEKhD56CVK2s+Ss7k49yXu6DHX2p6ex2sqtIYhYk2KpG2F
clHh5FNjXG86bsWpfOhZbeTehHgrkUMuf0gjry0JMKTCyCdGWUXzaIQdUjSi+TNW
mwFI6QA2DhdIk58MJHRBv+gHDfWFi5i4qpWFZmpv/t7YDmkP+SgVOQ7yfv90d9/U
0umy58/nikYC5sOx3hv/8o3IPLbCjIdL7wRRMnUTTGxaWBBS3ALJdmQNVJvNL4d2
s+LE5NgZYuFjg2RCC2rnfjqhF2H1oNDX+iOdPVGBA5WWBb9bO7b4BkwkqRHt+KHs
NFliSGME0li6vnB3t7WCVJvoIqkNGaAZP6u2MhMwx3URAetOXh8SRws3TX/5+Y49
z93afvqUCbX3oO4tUReoVBuoenLRMWF9zs1FtYMoikjPnuJ5juj3y91XYNfxrPT5
4UOjP93eIdyON0OdjusXqEvLJxJctBr2jPfxG2Q8eg0SxcEEJPDXWdUOZ3hVOEyC
CQOB0j7uZeNLAuEtFy9ZZPYwDDQx/9Ar/mxoSsitX2FkQ34ggQxHoXD8hzG+QbAw
FMoKIh1HFVGjER99NvDDRogeAmL4tDZyvbZzfxSiyL6utrX4cQk/cD1TEcnD1LKZ
wlxdME3L9pGEmTUnUxx+9JqIHIi56bu/tFvaTTB/xZGknNUo7a20B8n95fXiQJ0R
vcaqAH/c/qvcgFc+LoSadDTR2OrP7Fc0Igs1lM8cXdYSN9eNeI63uF1apkP1Tz0I
tr+GZn9NAVkkvQmHrhJhPKHe/rJmRHnVu87wWZ8tlqEgQmqBbAZNf6f3FojqLBVi
ho+rMSx0MpYmrGDlut4MGOHWgR6IdjqSZEJtS7TqaZ3+ak4V94GchHQxh6G972/T
FaEqDgIDLR/zC/ErNx8D4dUoDpJI/mfwle0PkUttS2ruUp0IH8+YqULt4EUZkPu3
V+fLLC6sWBder6fqDuzR/k5/lSN1kVL4OXees9XtFx4VFU5FBOPTd+XaBtPFVwNt
iowjCnekKPoW4NMRRQrOsg4u2E0xPFkudkCr/3LP2Brr36Esi+kdbujnH9iz8SS7
lxvkJffmGfeILUM13IfSXec5K8BP1VG2MKgHWx5AZpDmw0PUSjWRTA1eZLTD6onN
1nrxfUwVdveb59ClqKxj3lDnnFh0O0ZDTWXNpurSj8P4K2rExZSN6fo+pWiDbr95
4AdTvJmf0vZZsn/Wqvo2yEVpbzsT+fnjEl1JYjxaFHiK8eU8XwwVLqiPzGqpBEkC
fcSvQJ6S98rtj5fuR43CWluAr12e6RtAgAa271nkuFSV2pVCM4UhV0NTFxAnd50U
VEcUqOi81j+xPS/3SEGqhba8SyTzAlA73cOnNr3zGN7Mlm3iKNUim4lJjg525jlu
2Fml5hhzv5JwDJESj5zokac7zuDF4k0ADyX7/bphd/HqtnfGJoXARvdb2cVzp5MW
a4ltzWETTvreiQpCoh7PqrS0jlQTN9RXHLAfj9cWkmO/sq7vc2eSLNlmLcTOw1VO
lPCHXWqhuSSoCml6st2ixiyaweYCuMM6EJ4JXYuXh8YMpRqnI1I8EQrnXhm54kOz
ka357s4tRbXbdxA5ecVJLH4pcioUajwPWo+2OXRiMLVRwJ6Q2UfeRsBTmZG/kWRI
W0no2n/NlaKUgSAo/Oa6YwxEjDZ+/SoP6knJf95F4z2hfFGkP+EGCPh8o6ONzSCZ
3+DHia/NMjffS0eomvjtr5RuYdzeaZtIqL/nenE2TIwjNB/5scvRXYA8+ZE/SO/w
vOVYCxY0R4wAlfRfB38hYIU4d72L+bEeZjtHXMeBI7YbKbFkIKi2K0n3cD5oYFxN
Upp2yJuO12IYPsnvlbvEASnpmQLFYuPPwmH2JJJ7zqTqXcr+W7xdVxT0fekH/maj
KDFNlxA0TQTKEAt+ZGtOtLeylAzVflvfgtvAsFVlNnAE1pi+FjqsJtCQmxZDLkoX
/7DOhN0E65nGNnmTiBdZLkUAjRwLSUnOyK3W4mx/VcGjAMq25IU/IxE55To6VWyK
JTCTRYvNBnyjT48/3MuDtnp74OuDlC86m5F1YPQUrGJlPt6jmh65Bh4LwVegp3Ed
ZPtbRNElnk7QTA4Tdv+gqM2YDfnI5UPBcwuppm2qMVpVC+oHI7rTLxJ6y/yEhTfV
FLMAw36Wamo1HJ5tV3tsB0xO3kYheFEVBWqYeKaIE9QtKD+5e80U7bKZpTCU8gTk
kKDxyv7rhESCy+Ac002PiYLW/Mv0yC8n3AviLZ/sqJz01k7c8OUeO8zUgc0+UujJ
th/NA1iya9pv+YtB2dYdt58E3NfxYVAke6qv1YywEjfxSSTmGs7AJA06gowCF3n4
YPeKvaSb7ADzOE8Zyg7eHyVJQMwVpnxdk0WxFqr3KrwknDUOrHx6kl5YDn0/Fwnv
b5wJmRdr6yvAil248+8GVYJFU9vMbrbbd9YxIOo1vOctEQtnc+D4D0RhW4mOLQi3
sqNCOBBN0TzP841wKLYsW2tmrhPo0dtQgbLPm1uzrX0AVoGVtPrDGNaN3n8SMEcI
i2qJdgUniYmhW1MYUjaPp0xKBESLex6KsnmsNLjwWs4dAEJ7HHtxS4Afdw8DsyLt
qjrtJlO7Dco/79K58Ei6bVANszoscz2uRW5loDFZdTQhOoy/0kgPs5QOZ2UifCLO
TLRLBBl9D/vpEXS7jAuVpC9spBSfhU1yQTWVZRZULEn4leG4x1tWv7FS0tNc3fbI
C/Mit4opxQ5aPHTavjDH5wbxtGLIZsX7CDNrfHTubp3D1IRt/HAs5Y+DoAgVRd0t
vizJI48hoVqMTHaO34AEp+eDISEPljzCCFjQifCtJBXhIIIY9lIdiNAzNuuOVG29
JGim5fZdnRWY/1BZ7hecOpE62QeIOET2RBYGERKXoItEBrzM/UOiWSr8r5dwhOYv
P0EcglluHgWLjLV7vx2u/rZ00ZY2d8FSYyiO7mYP7eSQ+V1pPM6tI5+p+pZ5Dhd3
oh0LXU8pRMor5rLh1FVge8iY9KR67HuXvRyWooHCATQDsXXxrPKNRlTJkPSxRQot
HHkwvgROV3KmLIKiH0xlmzvDXzeNHwfnHyEsN5hnkeD0XQuXzc4SZ7XOKUVHLj1S
sax0s0Fe4sT7wgE5gSt2cofQp5wdJTfjkduGkMWELG3kDk4Pm9zoADV+f712MYco
7wdU1E6+K6ronT209UJFDkvWbFw7YyLpNYnh92/LaIDfUFBCZ51BClYRVgORHI13
Gqvmm9eaginRUfmdas3PK30aEp1O/dlxzpPMl41Mz5akhcFMEJAUnBvrpi+Ty6f2
85C6vVWGnhQgszqt6B6Ro7ER72PN6IzFLLu9GJJVLY5Nl8kLoBIv5Hwdpl/B/DNW
ioxk/+25Pk2enY1J500X/efLvoxo8IpWCGsf/7pFoqzfV56mQAk0LCM/wZPHeno0
dThxxY/E2eAvllWIXssJmEy/vnaWOwHMHzRp8sATLgjNyQS8m9jI6knjEfPNV0JJ
fNuaGNNdUyvlKwzbKVfqMjWDAm9e8i7KDnV0KPFAc6jwziOy0TcQoMdeALsY9J/z
qU7mxjkVnLzsp/5RSLq8RxrARw+D1DTQV2OpvozEJyhfltnXrXp+62b94n7Z4Cn7
HR07csvEqr6J7pI4R/P8IO4nbg13RIm0lVprOofHZvvbNQdDLdpLTRy2ZFGUHoIw
swKEefNH6XpO5PMQuvtyNPYF32CwuRba388qaCR8RYtJpU46B0ZO4jUwht1GkUzg
ZtQ30u0iClDZKsLttn1qoL3nKhdXDV+ypUovGu6k81kBwTU8waqQ/tOVAM5bkB1J
gMZsSHi0UsmVc+TGbx9N3qhTcdkcdOQNjPMGl2MZcx7Mq5exUTuJ+/3h7mGYBwnA
ecX0OvTxV6CEm2jKYwpotyZwTcM++YlfGIXSBDAk9I+7sIxfLYgkGuB020kjtl5y
/iQ2Ogff+aFhXLkTUHGcKMTOBDVO4Qe4eaOHg/aBW3/N0HDEmoByLk36oQ64Tlv9
Alilr2qxKngzhd/P8wBnC+vtHJSet2yfgiqQgmrqMpXjyCMZqUXvGu028DDYEj5t
z8yLFHB7oaCC2WK7sxwDK/mtsO9FAyU75oRo0z0UWIsZUYliS3tYjJEpwGCTTWi8
8xpsY/ichqeyea4PeV0Ge5yeyNiEknFNPeSHvOYIGzm43KKsXbfgdnGjz397fwk+
CdR8LycQA2fP2VWjCwoJiNVlIMT90VXCv+NinCctN5f/pPVJqX4F6PjdFsyj7zg0
IBbeVblS4mbBRR6z1dA66I6u+oE5fOhjnslDf8/rRE0a2TebunUVjSqNqO3S08dE
huqL3g6FwcugFFRCW/fF0CEhMfUUfM1kh12/l2YpNdHYt9VOcjouI7rsvAcG4UwP
i6AiDdq+YSowiRI2ppVexQMwPJuSLgakSYFdS37Py9arynNzdfIG0Ql2ebjIX1sI
a+c3TdSk+lbxRmjM/6vzsAiK02wO3ma750ht9xUe/w9uc7r3s4pk5i7umoLL0j61
PvM9QOKSAhPEc2jjsQkp0xCyOBgRUc8k0Fcb/bfmww0rxCd+8X0+lMtMCqLKvvJV
WNa8A3FTRvgs2XKjAtp2smAaCL/9gpJ752A2U9HvZJ+KblcYYfP6za214CDMisSF
gu3S6WJymiSh9q5is5SzocZ7OXkfq7rnRZgZw21Vq5ju21MhUTfClQCN6okLMMIG
5SaDB4PNVqZ2G4IqfrS9cblXrGsnLeqcml6mSiVRUHmECfbefyaYH9UeAKZSjh8c
rh2vkqklZCGZ6jpVKuEU9yQw/AQ0Q57samTYR/ivZaW/As6ODU9RfEPxHmtbAfNq
2znZHVJgK+SABtvyWkmQb8phCtMuPBL5Pc0j4SvjTdN2AW+lYGxdZF2A4ifSRTII
T7zsqx7XaOB6wM2shvti9oCs3RU5cLTyKeKDHjeiGluLHfd0jDCEGYmP1S0T+BCe
gKfVaGPMYDP85DkI2F12xQcDellJ46mbho4EWNoQSnoisK8ivDHEY38PXJ1B2Vt6
n4govCRg+CXXaEozWMZXGbO+8shUON4lAKrwiF4OW0GNxhDLWw1KVXGuMQlByG+K
EdVK/TJc0yphfAOp0PiNtj+GJHqzIpM98MS+7VRajcvT97tTo0dkhnAMOXCnZFRg
Grv7rTl3Vqovx7JKa9sSFyY5APxk9ErXLwa9K5xDUbFIty56xOfZEW2MyCXWD6yh
uGMGgC5mljlUlPLtSX2RNSsH7Hvu3lQOeZzp1SApxsZ/SXVu+6Sub7uB7fZEMbDM
YhWsK4sKxYEUUfBKM63TpCjaubzMPaWG7ezIxSDRyzP0yohuK1VzXGmgOY/s2JlR
ToldqVxMoDBNvBIx3nNZRvkc1hOncHeU+uJD95X6BjxsUUZV+hkfv9yaMu2nt6ti
+ZWPlz1rHoc/1v8Ul4HDfK99RmpEXvHG5tE9IgNlJJCmsjnQiBYf12GfQsgxXh3M
524coUHPwPFHvAQUc4/PYgC57gvgM7QAyF1/+5RG8tRmfUDptUoVpuBTZ9W6t4r4
1sP4ME3YLXtj5l3+My5bROeIq3XPlJz982I12fm4BU7Waih142N0SeTTyx/hsg2H
Yu4SmM9YRRc2nQngJYNnlOVmBnYxje8NZfgKa8UMfI9y6GkmBVLopCM0ySupX+Of
dk6t1ER8S0WRg0oE7/qoRroW7HYEOBsxjBd9fC7gUSnulKlIzvePrFreyrvDZMeJ
5H8z5W2PpFRLRPMahBARJlbgqm66ldfvTNObrcRpkyCIY84wghcPjv8UNiuhqKqQ
s/gI0Vv40ALFcwFcHuqhoF/UC7SXm5xuDI+vTXYdoIRBqqT3R4Mqq4WPUHoYEVPr
CFsRbUMQZGj5WT3l1S/4M8uHBvolS3Pmz/fIFtTivZqlrHcmixtH1sEgnoNxQQnR
IbpCjdeJUH/7bwHergPXV4kOD72bM4iaMT+GQGrfZx/5D7fdGVGKGhiaLHH7Oklw
WVnvE5g/Fnwb+sCr6G0hmTcJtJ6jLWGWCKlC3vqV1bnp+vwCm/RGBPJ5AeowzBoK
u4fk6TWNj68cGw0FohzQ5WX/EC0xSXarBAbTI5d0JiwCjwbvrR6rrREAyW0bTe/I
xAeziC8jpzC37mFIiKfz6kwgudnzbqXZG2kGa0dKnIIi//2g026iRW1oVZJOEBOc
8BG5RNDjH4EAe4xNHyXyahZsBsnSEzXM+ect18NZUzxGv+NbxqTH2mx7XYzCmqGY
ctPk5L896sICHx8VHiDhqgg/t1XGyHTyjHnPgQXxZjPbd9tRWapBz6rIE9LXSlxx
jNXKweFVTTPC6l20vv51hCw/BKIryhrR1Vvx5HK/Xsrwl6hOb6b+3gCYmtg0kwN9
F0GPajbQDtqpwIXd+xdcTzVBcK+JZBZ6aa3LR5sTeZGq16Hi+O/SBrUaX1+ar2T3
i8nQwq6tYSKNEBKLkW880RBfE2Z2LK/ZlZlnRaGH0dRHsj2UsS5wFfQJRgLLhLlb
ITbyxCYxlLsvrkVRSoFtgbUOhC7av6kM0Q8MqZuBElt8RmPshEOkA3sJy/mUYkH/
CwsPvgSp/Voe95I3xIlpUYByMzbcY3zn794UF6T5Y9+ZKoz+Ua3ucdoJeeRiDEHn
CplJfhjNZ/+WxkQwGMV8nrA3gzMqAJTXRzxCqDsKBGAkUPFK5Uzsz5rXbOqsgKsg
CLUzLX3gpF32BA68QS2pP9ArENGJStHDJrjJwcC7CTI8RT/QqrbUAQemTgRcnCpX
K8Z7uRO0kotRXyJ5VEVAAQli3e/GzLEDmW4lXbpZj3v/snwIPAG8pXSLjFAoX++V
rHcI6/OeGsdLB3Roesk6FCoEmLnY5eLBltzkT9skUL1mYARPhVFJLkuOouqdvB4X
66U83LXvfVy2TGFAutJd2pv4sOYFhZ553rdLO4c6RVtFHHGZRKGZspx/zXlAtlvD
jlOFcmT4RgWdmw6sNg4ysQlHMgdRkiAasni9ATipBCnFsOMgIohsBLs2BMYSWzv/
iVHA8HHykmWMH93Rv5KwI3CFF4quYjTiOv+nCZrTx2dwvELXdGQ53IItY9yQF55R
wIi8uvtRDvk/mq7YHcL7kP6bWY5Gwx5B9jFPFElf/N2NOf8SZK9IGzQgV/Y0eac1
f7gKwVNzKn+Mjt/TDjdyZiAo7F5qV3XPGKtLtp3WWU4ORNRxgwXs2Pt/Tgtb9jku
ih6uNOKejfHwCGDwIqXcQOOYAGNerkojBwH/t5ERf4bze/94u6IDBqE2GJyO4xSf
6suU4VU7E0dqZjJomPO2zPp8rfnkBqYh4gzP7NDkJqdLR+Y3RURfP/7PYp3lvce8
PFi+rabNez4YyosbhDLRaQDf9uifetGysgpvbAUkUMdtvohfWI1IbWzt5F4edTCs
MMwqILGDhUXNYe/RTk6B4zSR011xTbFwKv8ZWJELals9E7A29ihBVbJiBMotCr6U
VdcXB2Z6M5C0G7uB3mAtm//Hm1hF2Bgwz1IpK+inA1xP0zlKUZK9wCZLWzKB+LmO
4UHwvloCO0981i1WXQxxTjc0xwEy22gzHosKIHRP9WA/6WkXAfkrwjO+cFL5dd/8
HLBBd6uAIcYMBPPiDVQqtf4RzICjhQWhRTizxVWtiJeqSSQPHeETuHBTBtzFhUB+
NQzd3s1xuGaLb0e+MApgVEAZxnWUhVslHYNvjSmkUzUu0D+WM81gi6FMd0zkQN2V
9rMhKRD9e5/BrkOFpRXkN1miwHXTFijD7nf3idhaxno2XTG9t5K2/HshGTegJz1Q
kxSs6lSbKELH19Wm40Oz6u+cZRd2fh5QyqOJaUmI7Q70reH6GQVUiqvJlJo8Kcso
Tq2I3DBZiyKjMhe3t9nwPts3jIBa1Qk+pR+eXmNNr8OFHOJdTGmb1OLx4Y3oWo7/
SzIJKZ/wfz18f4YMK6Mrb7wW+yr6ss8+ic/oOmm8aIfc4KwIsBvqCtRwoJtXhxep
UGLDEEsvNCeQPzL4bxM90ceEH82y8I45L0pkpO5W+mZcvSQjaMf9LQLTDeImCKfx
MdbzFYku6zuUktbA/Gt5+DIIMUbKtk3xyu8r/Y01ENudImLiD3WxSVvcd+k79Bb4
JWD+1eH1C9XPrqZL1byhLKI9IWH9iVxzJURwjfESObCLc7KZOrQu9PCdQlCQ55lo
Ovj1rBbqNEm25Xdf15x66e1ticOWzPZt+rpE3U1gFsfrnnuxTl2PrUpL3TRiLxp6
M+WWQ4xTolx90KVnaLjuni5b2PbXvEFRhN2qgkMQuoOEEQWSORHjQxj+IrK2wa6j
Le8LFpw8BfwVdlrIj/BzeO7oU4efG6fKKqkXtE92joFCPLsmulYB9rsisLUYxj+8
y/8qB8lbzrtsIk3Uft+x8ieqI5GetZKEVA0R4gvgs9kOnxYDBHdgej4e1FqtYYjb
OSIzQDMl4KSN2/DUHn239wSUJyT8u/1D8LSuD2/RqAH4TJEVXD18mnYn4W7rRlx1
VwELXRrvOfXsULYqv7SnP86QdWASCyEC7lNb9XzOC8qZu9/e152usaZ//uucWDH+
HtvsQLsHWmPK6jXbQaxAPtBMxXCk5Bf50xE4W0bOB256h0hJAcYUKisba7FBwKp0
DEdSK8hLtPOxUyBm3P2TW16d6ovXmSO4YF+hGGJgc3ueciYKnUO3HazVE94kZ89i
igiQ9un9mpr6FHU+Ti1PMxXB49MnnsmgB48c+LfZvbmJoVlX5ZBtqLm5EQP89hy/
4rWJmkxhlm+7bHS0hIxy9coONWOWv/ti+iAfVx9fAjU7KIBuQJrcx8PC89erc81k
PlgaqD+OmAzDIqX3Pbvz+YSofEzT8DOm7YU7N0AcEzSr7KhjEA7/mRE6OXdnJjxI
RD+A58+94OZlcDH6YCIQJVzpc61rwY1KsDDj5Wpptx3RkAPLvY3Q77auo+9lVnXe
mzPsI1o0X90hLBCrq9xEdvOdaRG/Al4y9JzBttIMqIA5F+5NzH+mwVoajBP1F8M5
j5idLSqciOslONUmKywVQy6MhW1qCyUPon96uE8pNDFXKXfiLNfVHkktQ+uho/uS
yrZ4cGzoACskDZe6AmasLqv2W5fbpr3QhCqr2vB1Fu2QHhuU30wgECpF4ttfqk5B
B6FTbtE1Y9L1iJfRQRDC4AtFhSDRmiw1ymc55pa5kMhFbOsIRbaFulRObH7tpndy
3vPli/4zqFdK13GOYohq7ljnW/a5mQ7Ii6SwAhnGyr0t9P78ZhJgL4K93ueT3K0W
qg46rViFWf/X6WKBTrwYS52XEDCg7plbBSNkSDN2c86sJTk1NX1ypEgdAUjOhOk+
x8iqXSaWP6Yg5TSmsQ8CZ9vJQyYnaK2Ye3ZPFxeJusSz5R+pRptE2RaueXnBghYm
BACAvk6g7vuSFSVKEUkmS4JgGGBd8Q4V22JT6lHyWuOVAU1L/2yKdpN6HcOO3GZw
G+ynx4RuMBrWWbVhIHYzlmc1LAuv3DoW/9GP3G0trI2KlEh0bdmcO+WSm355QKhZ
Zl5Xtp5XA1FRF1v31yWhlDaOij9/STmBv5wwUT/LV1lZv9FpJwwm7e0Sii9TypCK
3hb+Pm0KTnxV1mjqURi20ZxCtFQBQcyjoDSIa47pIpwi+lpbi84l4Ft5hDl4FKcq
Ycn8vlcG+YCUX1BdaSUOdxxxMBOqKrEJU7o8GsksrviYspa+rDieqIY9x47aehnw
yEtYxmbXykAVWE3rRWjYYlQW58/faqm7b6HfbCuz5odrfbhTM33NjJwdEeVKKSLO
Epaye4tR94/z7/j+jKMQRaBtdKyA5CBoiagNlQt/K8dmI9PD/IRemBok3YNwYTMk
lM8/gRBdRrYnn9dVM32qL49NiAtgCRA8HJMUgjpvlPrM1HmnwOiaHS7lNZATK3Ok
q6Esajyw+3pjvXKPP17ebR7LURlAlu86ETi1tzXHEr83RfrwRFHFeyoqzrwz8yQO
xk7FFm4xleLmTOTOR/weGt/L39sVSz75IraAMSA5pZBSGzygmvvBcQVYg6y7i/fh
O7QT6aVAFL7IB9FtU/Nt5uuQrjSJm8SOAQH8G8LyhyXZplgD+7tUFPo/tS3poN3J
BroeMc77QWt/dXSarov94uemFyzQQ2HyGo9le5MboKgCagak13PzzNDqOk++AquR
h2wgrEZSEVUb+xHwJTe+n5iLnAoKC+Ze5sgUbfJ3RfBXie6YIXbZMhMXas6wagTA
2Tvu9CPZTNo6fOnI+E1drLVaMSwx6ZDiwN/G23QDGoEWaUKqBXq42KnZWsJydLGe
pCRkSz7otGPBeewb8pEX4/nwIaRufZyiYL9xJ9r80NvI3HBKSNi+K0runw9Xbsdn
E0T2ag1fsM6wLGgCExtE4Bo4uNGM67qOj3RdeqDU+mvXTdYpqptuyqotKpU+hC6h
i1s69MW43PuO3bY71SwmaMU6gHgO3QvSYQsVvN6iHojyZH9f+M321lHy4rBc4WU+
Ak+Qz8ujPCKn+fZFzp45MI4PGzSKCl+yGr8sc4E8ePnbmGybIsBxzkEuxhgjWQR0
w42C5/4Aibcb5oDUSmyYOoTVBJ5rAgDWkOKhNxtHFF3x0mlBvPn/Mj2vf7xHreZ/
eEvXI49foRyIrQAoRjwANQmKz0y2CCD6kZuNolhieFBrUe073kYU20krXjVNrZcw
goecrwoVtY2FCONxz4FezvBhBZ4y8kggaiUUZIWbjUqUSsZY3thWqS1a5xWE7eUq
gNofnF1lKNjUd1EQvZpzUT57psmFFCBpXvwZvCsUPm8mVN+qscYOrtWevGKdWP/l
I1UiOPmUa8/6GevN8THFGvSqXqdsErhXkZHSkhO4LkJNcbOoYzrmuqBnrFF9Cg2O
s/8h847hzrYsyceZQd1kzVydsSJVmsQ4meKplYjzLtgBJL2ustluxLJzKAfgxhXg
46yYMJfVmFdkoDKUVtkX8d4z9uh4OsEP48Fd7ofISnAMg0S2FYxqzbutmgmCZ/6/
nz+v3GqspANgug0EYKayAwBYCiFN8U2N4LSepqFFD2RCWQBCZpdHQczdcakXdnbx
eQ58zaopj/OnbNVwfqtl4m3unIH7MjhqrUUv7PE0Fd6w476dheBmmA20ZNciXOZa
nZahrBQAp59t86FXc0B2eFKYejEdVY5zf3l3qaqVSXMZarMHjQCzFrrbDH0j0RK4
fmLTFutbuf6xcaJ2wKnNrsVQmhoyUikUllZ1xvn8pya4d6Tj4cLbIMDIF2Wf/yUj
Q+sO2qkmp7T1EDcYmeNBk//R4+13tBx8i/4mt5oc6EbSx9wBwKY45B0CvGbJ5fCM
4HJUX9Hbax6Fw2shN3lNpLQvvK4hcvytwi1HAOL3s7OP8c/Z7W7P4s8gbriv7O5p
bweJb7RCW3O29PLm0NYg00jH6GXrAMcHaKvSwzrGZ4TKcD8RTBGrh6w5S7sLwCzU
iYuDE0grspsMqvumDuK9ooWBrooYRKADGaHcBTsPjX3R/ow/rL/FQYC9SeMmtNPZ
mg6+8Bk4UzWTuZwvFGVc5snxh5RT9zOycvdOlay3N5GiPmlqx5adv5YxxfsV9/hO
CEEk3GnHJe0Lm3242y7gBidkJQSa9K+bG4l3Pet5wC5bRTGN3lHtLybHWCoX4bwH
Vp9WjYHOQs9mRGwS07rFRU2TH1/ZL5oszYjLpdRplv/vyyOkImZXr78njzFBT78T
3Na11Q8SAeEBuh8yzM968MpJXXSb5JPf0zLA9JZtAi+VLGbwwE1/8/iFmlXApP6j
aUP8JWrOI/VfxdMavsBp5ThNptCJe0ct+T2QKNzBi1VXrj88C+rU2Z2nBQyWEIxJ
02WoYhbB8X1bFWFZxW+w/WeNiTX5cij5uWY8flZfMSmlMgsYhq7q4pcXz0HdScIC
FyWvJfGPzRbDChZYl5pK3PehbQ5xunN9V/EU2QfwbIEhtgUTrz2ZKSEAHKNsGiKN
IR6U4xXtCIwDEymVLEEyDOlaqNGnb6o/HRd+c+UtuNPzlcUKKhkHr5yIjNmC+nmW
+JLeBPI0r5SCg29iRVEddViM9PDvEHx1mjNEDUBu/LG3CzbaydKps5+2H4pmNdCr
XH7M6jgmMUW9mZm0ij3UEbaDTlI4v2nM3XiRmrAy1WTG5FSK0olHmvlQQFO0Lqv1
dhiZwlpPFMREYBfudEw5WyxNLOxdCmCQovpgt0nN2Pqoo0uJBD6zqAfGH/I7GckV
EUpy2Xx389Q7rw5tsChovdPi/bVnhzsM1EbXNlLN7RTfzvwVM6amuE6LJSKnSrzp
AcZI4YeEq/NqHHOCaKFxE0l9lcb2TW0jRo0TV0Hs7R/vJ4Dqn+/XfhFBp1AJgiGE
1StAwQvX7+b4aRxcjRsMc4RYeFcdXVd+cUOZSyhr00gz+cj9Udi8x93tAWNLbWrj
8ondFU0DLdryk9ZHPpQfTe7VW2hfNDRSsr0ISQ9qRspu3HUEBoldwab36IgNZsm9
vPVoaLM0j7KdGvw+mB/8K5MIQH8wmANSsLWFcucu3KXJbm5AhHmsM0sjWdp4SKms
9A8LIQbxs7FI/W58gEpd55CUDa274DXyDOBK5AXMHpZBKHaWwiH8S0s/i8/rHb/j
+jUP4RIUuJO+PSPMZCOaeFgqHjHzrBt+C/YyhBjE0rWJKtpY58Ra2BEk+licWESE
ZaYtz5h9x+yOZFgUDxLKS+4m1tqSjEwZERkNsHR4bJyT5tGfpA6PuyHxGdVfQUnF
8GWNutVpC+s5RHCIu89CmeR+ArgaW1DEDXDftnGCCiY2VhueOv8GOPViep2J8I9V
9SUkQUSU97gYU4nTU8tIrbYGsaR0R//jZgjvfeJ6bxzPD9bR72DoRLkMVR24jjhr
vnnwIHTYfqfMmCZbx8WdCbWY6QmWPBXw04eu5Z8YRCVdK0KT6bqqJKvhPE1qFVpp
eL2mM0cRR7YtS5KphxEZzzvZjOoG562AIEPmtVoGek2CYsR/QwEMFz8jtxDhwh/z
HU+B1RNy3PZR2/H2lMzNEuHwHXCtPiflg5BP4Jd9A/WxPYvgUDLc0vUG8iYmUV+A
9PTXrYFEqZfgOKFZ1unfqq0sXZfHaFkwNbTIqw7ROO0zvMfNS90cLSuSfaiF6uSg
Lo2xN1+ith48fD0VfqYUPyzsz2vJ4zrYSbx8w6nhYet6wjYhp6G9D+QCzgs6CjcH
dQ4pMuoID3pWWy9w/d2ZiTudp/BfYwQagIMynVEL7zE1kFwaZcRQUGC2DFeWjun3
ttHxdIMXQOlHEoncIvOnPqfSRdR+544v+yFh8HUriIpc4yIXN8Hh4FXrKCSpS10C
gPbTbChlBNejyvFd39olT2/RyZVpJR8nuurrd/ue5ADPJNwrFP/G50reVyjd6Lfy
gv6jn1AgpzSx4EBbz5UT0be7tdGJN7JE7SSzTrsSSEvuGXFLowxWP8nPV+Rj3GQV
PRZwjhl/33afS6MQAzNb0P3iv3jUEM2WhjDB1UhVWSa+XGgZ589g8BPLmvVRV2lD
CgzeJQFxWr6yiVozWXu0JRJ0npSBj8IUYTriYAhLm0JFBQ7NODkf0lY/aq5yxrzs
hWUHRaC92Mgjiyg7THrl3pXLNIqO6aAPDuNu1IMlcyTeVwj9PdVyAJEQ+l74AhzY
XxzoiCFJzzz/H+Z745T+NaQjf3EOF9v/Az7wgySA02QXu3rIS9dG077Ni5lgQGms
MmE36wQi0PWUtI+2G0JKuLIlqCPphfH3UfwfVaRqUpvUOXvIfVsndIf+pTHHNX18
dDkaMyZaI1D5K7PJB/ScDOYmCycnf+4CrQajZ6Rl3EwXF1ahTflZlGTDGCMwFRip
YdIaTJ8dD+RInB/4NEryygtqyM3XpwVaqZ8NRHu8WFTtBOYoh5bR4bC1Wt2NeZpm
fIKDE+fsTp1umuL0vcTAGRJSzYBUPhlHOuT9Wt3oq8XEYdv2e3lg4PdrS7GBUn77
uEKmssptneKcxhNXpL0e1ppy20NDmOwC3pMQuMivAplPh5ddd5p5TIIsnL//Kkzm
za+4wvPzK/YBeuHDc1o4aRubo1sfV3N1bsaPG9CMHVLfOZxhxKqSmtj4dR36EGbB
PYho/Ez+dN+kmbt3WbHGBoetXIvWlEgKUTFlxRD6M/TfAcOLZVV//LUHc6xc35fA
T9bosilpgedNt6q6Gf9j/jDRwlQIXCB5yHt7Eg+cMBBDhTQZeqTxniIOO0Ln/U49
z97WU4nAWOuC3ENeeSt1Gr0mrGfDIVjh4S75U5YJsBZWvazIINs19ufL8t3wfJYL
dQ1pnS0h7LR4RVdWKNY2cwVskIuGmwuX6meCF5juAMNodZ/oslj6KKaS1E0l09WP
UavUl/pprhMmca1RysTONr5Orlyi/H98bc8aOeqQDdGF0aHbmzsVpqW9mLHyOh69
/DwPWfwUWmHbGBHEUfrbSD38WrNzooVlL4SYWQ+CAUwltZJMop0/agTIRPdbxsfK
BPUeZ3DdwEeWavchi9fJRMk6UN6vekaiKPX56VFfZ95GybyeWQSDFiKveBt1k4Em
vboK9fkQfHeMf9Ifzx6X4UaWnMiYso0UR6WE39nQ0ZNtPNOnE1gLYgmoOFaCGg4z
mnr1AUVY4NCsZN3EyZdWjq7Xp5evvTfT3JTOawwj9N8TFzu6o5+ZXoF4YjwZ6iRk
iyql309MXHvRlTvGUPfNwbWEnkzR/15bM0wXagn/xMtXbv3N9Rutd8Dr6jQKrxsw
EiFMPcDp+zYYDXKgfw9WbLI8Q6miLoMhr7zia/6ZFconAIATdHTjTK/qMn9lkI/C
efkOxSW/KxXQ+SiIwyvumxbBrvC0W3fqJxBIpZc2bf8mwNbO5qCj/ppTSRocDE7y
EEYQHZGHxVSsaequQh2HG3WryxEmGVSHCxmLtgpXMS9u++/EvxOg5SmQfmDxLs5X
XTS35RQSAkM6DZW//fSAnKM0xC5bQ9T4Br1tSvfsbDj8RSQ3GAbpQKaX5PRW3/fg
ykaRUpH4muo5p2TJ6oAgoXTy/RZeYfHJm3N8fqYFUAuvepj3rcQn2fWec18tTy6R
MxAxo8AaL0245UEu8e/6R+o3DVv7NfOFQnUUp4nA26c6K2+woJn3NA95UpUNhnBb
Y+61y2p8LZ0Yy0p89rVQXM9iIlXCE6PUUSv81mYlDPpr4WPS9whyh2gDJ/wl0UDg
yIwx3mv/Nd7Bse0sTF3pKhWAzaXsqqQINHo3e+M48Wd7xk1FbqYnN17wQDKpIc6B
v9Gx0Qd8RhaItijzj1VvbJMuaU3V9K0iNz0MkkzeM6ujT/j8zqFIz0AvLCZVOFas
b99hE9A+nJZ3vg7/gdyVrENxUHbb90+xgp+Gps4xMt9leedhKIv3R2wNverMxmo2
aEl8fYVK25pN8ObJWcBUrUVin7Zg1f/tfLspV6KSY/AUG1MZftlhoWAgQO4j9NiA
`protect END_PROTECTED
