`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zSqIMDmS9orHPUTBFYQqC0iUC3SiHu3YPDjimAWdHM8qzIosDa5pHYd3fgv9Sfdh
0tmy+wRu3nfcScwpju9ZL/g0REos7nICLfYSQueLhWqXahzntjOYjcKV+jKhrrCZ
MInG5YizezL2+e5ZF5BOPQ5sNrV1YdSTqsUa9Delytu+u7/EtkM1t9Ay7NTnPPM/
XtU0J7klGNUk53nlYDq2QoijMmPOA3aIWlkXSDbZrDZvmq4hsuhUOG0AVhqdDi54
ZJxjEixON4NGL2bw9P/i7levH71z+86valqFPiaXaBTmwbB2kfuBOZD7r3GTmLzD
zqlJDjBN6MhS0elPFA9StPRAX00PZDeNbSSE446J2JhmvHCc5Igg7OwQ9chUNNxv
atN1ZaM2v0n5RI0+wc5fRwGjlTQ65mMz6K02940k1u068OyPUzWtspQvVPc3tdI9
6g7puWoMC8lOz3bteZkPzXp+uWsE/SKEn6OckR4h6TVNQMhT4dvqHo67weIEgsPf
/zMRw1kIaIIs62Nlu+lvHVk1rjL6zI+mq9ppL1KrNxMGBa46cRoO9sjQxYEPgc4a
JVt1IRJUNgyzu5Sk3axNIqg65Gt1aFkkZN86wXvdn0i2JzQUWPe2aX3z7/0o+0vv
NZup/PzzW1IDlKzwfC/q94zPVdrCEK/4/gPZ0XA145n0tsqAH69P5uGfNGc8IEjj
rsFoKw/0Neh5Tu0EmoigA0tPA7lxLCeeebWbxCq/I3rEHCftQj+bHV+KFmlKmIIV
WoQV2WYZjjtZzMyEoHCWpMpgbxISYhjsWAqSWcDHVLwhiHv9lE3VEhPVTAwIR8hS
pnQxcx0ACXkSaZpeytQb1gjDmVRc1F1f2GpsR8D6c5aX+jVQVvu+zlpwtfBgp2nI
eNev4uUeFLw0cvIsL51VsM5+7Gi1e9RFyyQViLxq3dyxqWoyWvpPz+mS2/2YI22p
dF74r5rFOO+TPGmMKxwKQexIfGDutXXC1aWO9W3NJKEx2U4oq/nBQVDlJQWqsDfq
`protect END_PROTECTED
