`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nd2MVchZhPfJxvFYUDGzi607bujwTdWJjULqGpB3aoPusENa7O26F6RgseB3TTbZ
+9kN4PvCjvi9X7h4pECluUA6eWJN5fwmuMTgIB73ZXvePCHzLpZBBkSW1bwWmpQg
bGPKLM5KMQNhZ1YW5gFC0wyArIRq6tBXjTjMpkDSQwYdgjJcdFOmIFWQFHO2m1Pe
4NkYTn7Ud90ET0vbQSTfg/6z+Y44EYdzW3Ae2Lxsl59I5/bd6TwveEI5MxAqDnMb
5lFVEdsyKfUAbGtKLUUEP/sebq/wZv32gDpNCjzRUDQnUbrgTSMXylYMIOC3mFVN
WlB8/5wrCMuvhWN4EWQLEdIdfeGwoWwFti4ThsuFAsl2SLKTcWFqoVAA8ASnHfk2
WgIoRQy3P1wEntTL6JKIM/d5QpfaRZ/bSmwZDnms+Wf1vDSD71Xv0yA0ay7litxB
AEuloiY0tZWpE3Xq3twJARysO+fYVnwJvpnJ2w3luFuU47PvZJ2ilviuvnkfQuEP
WGaQo1EK7Kb7uhN8zbf27zsg6G36pwGNunnYXiOXKFwlQgKm0nvyxa+VWjAWijY0
sPW7XMQZXUgrhymC2DsqnRnK7mvRmAjqHKr0jAwP3GVQyTJ69zHb+f3NCATg59wu
hD40IBZtfBzgwrPikbCwPyE1uScGLrmI1Ky2EBLPwqiNS4jleMpYbtc/u3nQ8AqW
ES7dAyrtMV7cmFpO39GnbFAm6snc2DUMygKTNpxOF1FXeD74O4PcCGtmp+NPNcg2
PVpWpemuY5Q7ae04EvpG4aAQ6oYOaet/Yn78uYW0zvZQAHhijEK5/J+chxGFszdo
W+AKKe7mjCrltLnguK5/mUpwm1PamMD5dKXCFaKaEK1lqBmSiZHpaQvyG2Ro/BjY
4VyFVFCn8HqTyfLjfGz/VDpQyrJ/bHRInV1mAaKaIp6G/DWQvFo3Lbqc2oJJLy3a
7FeNspEnQXlRM4rd+UVgJ+i+1o+kAwRZ4Yalg+Otd2jHrbltICSZIIyigGu6TLXV
78muCeQQUpqNA8DTgCA4RqQUHCCsWMcHh1m/y00cYs43DieqcTuG262VgCBhtccX
g4bkQ6bcbVhAsOEF1WPUe30iwGrM/bIwpFpwINRXi6Lq+e+4jJbxQqHoxXSYe4H+
l3R2BkoQXuBNlZ+KIwIO2UmfkYK/6x6C5+XFTX4yHD9t16NKmMhTEIScSeLaJjYZ
G4AVoOBsfWjjd48vxfmVuQvOwTmmKhg0pNO+hSDytQQ1jeqr+4f+gsftoZzDSQe0
G/8Qi+3qq393ApPsPoZRlVuUV65+wpMD5lj/r3H7oD3QQ9Sgr2t2iPf11qJ1oHpD
fwGeTMeteL22Woq3oUpfdqB1g0IUCUaJhbYXatEXQaS9iRqIPYTEbS2xpSLZ8Yyr
/YnEKbWJzDlmUbWm8y0e1qa79B85x3eNUrGF0mXCGHyt9F4FFjHG85eUHVYnq1QM
OmuaQ3cMZfIELGuQ0sI+3CkdoTJVl5jIvk+DsbHftcZ6sfp2i0wwq8uD7c8PZkj4
hTRTg0Wr4y5eo3GHSe+Wfb0bNn1AO1ZDKpGVcNVUkXuxTE9Yxpk1+2MPUQeBzXhh
tcCux9rqF4ASrR2uRPbfgwExwNPW9J3oiCbSmei7uoHoR7f0KU/lxO8CQebi+V0Z
K4QzYh0aSyIdG+Gz5bP7rk8VtZsHiwdKoE2MYLpY49Q2LmiwIevlW1ZoH+k/t+gZ
+n6FWhDIgsQ7WImDu0y0sPdCR+yDFySAyn5ntXK6vOyv7SAF/C0VvaDnvCNDCjH5
mAnY3tefhlLZhSzwi5qqTvLFzXsRCC4WwDVyLPyBjWU=
`protect END_PROTECTED
