`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EMSNm6qpe6VcCEm4P2sndsvn7YamRutx1WhpTGc7hgtd1AXoNdFF0PQXmGIXGfaU
K8ZZDGAGVuVBo//mQf+zTG2BsG8gMDyLmgnDaUDwPfmYhqBZc1A5o6U2t9QvBHKO
+dK02fz8zMFTjicBtK8FsySr970rMkweN0EnEgCnQHRqWWzJAJc3jvrYn86miQfW
dbRv0Yp3rUMnteinCfdliXaVZ38BiT1xPoUlrHjI7TIFfoeWljZG3eFNyzkHv49L
nKXRgAfbflL4hEDISh9fUF0+cUU8gplf4XNGHcgEVHS30WWFV9nU/0GcTbZXNT4y
92ukriuPy3TN6NvDwpbudxyHWvocy7mxnTvdzLZ6lbn8un+SFX3LxSTGk/eW7P7L
vj5eDpJQan5hRRDR0A+HjmkPnZbqOX/YcckAZ6QGiL3oBNUDQmzZlgqVM3y8xp7S
Pj75i9osLfkz8IPwY8uTxMTg7doZ12ZhVAj/o2PzkL8A9OCzxsVy4nMqlAI37Rsx
AomPGvwsKbAUvKgU8Kt4j/7aoM7YKlQYmODhTKSdRx7i44FZJwSlaCBmacOx50mk
`protect END_PROTECTED
