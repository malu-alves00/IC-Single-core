`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zAoF2AbOPWpP610gjv/wRXtrumLI+Y20kVdvzl1Ju1PZ4eaoJeqV/0h3Z1nUDUVv
gGcpZ+exmzpt5W3grq4fZEob30ZPMs6wRn/8qGnmBSpgMuQzwPf3Axf6bSv//FR/
8OKxmOOLhGwKKKqBAdCaBct2+d2KydifUzz5BKKb/s8RbtK4LQ1aa1rzIBHcMhee
5qPPV7OQeKHBsHmaMyf3kZRhOb3dfBgVJxCfYQto/s8G+Wg5mnwoIDw9Enh2jlEA
oWT9v1jO1BBYMeedNUK8JI+qapta6Zh4mBQA2ZEcj0/kIVsr5qPNwa9utw//dj85
5WllWRfwxLm7Vv9YxMdPgUVlGkg+KHFxnzs3lJBryYCx+lArIDNDRuDOwmd1QjHh
kUYoZ0N5KMdplL9yRECMw6wzC1rNaahxsS6kF8ApX3bJLmsfM78AmWf0cHXK4CUK
ephjbUFYVNHIrBQ05FPuo2Sz9bnEjOr7EeJ13M45I0r1YAcDvAYJCfEcww4xTYq+
mKf2ZzRhX0zi+nji/GYMUzbbAP+6urD4BivNqlVcT7JpQ4Zo6mQX0uP8ITw+8HBV
+mrAThV3esoJliJGkvqDxZYhWDrWYiHMdiMuQhUvS7BUE55koTwqYNd3r2sqff+Q
+r0GNtKgR/HstPXVAqXld+BrGX/7OjPLg4vLwiQJ5X2LYzDqwM3A+5SgZoA78MSW
1AztxwDKH47U05NlIoW6Z+Gp8Sm2IxDJ/CG9WHUMMJCZj8OZMPHhxKaIv49LTFMj
jMi52OCLF7F9fy1b92SN3yNMe/rINxOlzdMIAqD9rWILKvFmDVPpzWyVOC8kd/9k
G02mu9+NGxhkLIQCN9DugoyUfB6ZCdHiPZU4jRllGHhP9gVcRUKUb0qqy+0wXUWZ
7kZSXGkFmHXrgsmch1dzkCJQg9FG4D42rX4F+Cy2cytbTHPSuKY7L52xlw1ZGMkU
5Ss2hKkv63Abv2cNVa+f2qR4jAUmK2UOHS/Ibs37+sM=
`protect END_PROTECTED
