`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
46BCjMrNZVx3GBR6/Mf509j/1hVe1XldnT0KUKcdfAUauNFH+KnjcISdRU2hzyBu
WLOSxSuJju40byTyd8NbYcuzbsEyIguMmnzM5Ftbe+5FUmdyle/GgrX7EmNC3QAi
sOzTwtGghxT+huduvT+h+DF8Zzs6b1lBtHVkR1z6vAPFoGZ4zeT/eKLY7C6xtPqE
m+Pv0/ano8cGgQQ15c3ySrY8u6mE1emA8f8hmVSM/2PJPgn5nJFsv6vFD2f+BZtu
6cBw6EzPliWJzWU2jMyEjAiAyMiXl/URllSKg257M28hCuh9aSLhlbiCaKhpWHaw
PsqC2Yxe7wEE+did2msjOnKbrcex+wvlpkv9EU8Qg1azNgxaaUbmceDPPF4Ur18d
U/Ro+QPjx/9lwk+a0O3h9t/qBRqEz2tjbnEkDsBuOvDtDkehp6G/hbtIlSCl4y2k
rX1965s8Zyvzjvvs2eLfSosqGRFlrLvCH0Kw/R3rIFTx2Adx3tHGOcPB6m2Vxwdj
njZz/34//2yVrjE4B8njzJzWWG3kgtTVosZ6zyRCGaef60/3Ceo4Zu2Gw8WAnH/0
vbDF7+ppE14b5eDCcR6qLTUD/3DIx4Z2bqR2BFqAum+QiiDcNKNq3+4uITGdibDg
sLoDKi4+1l2kvxE7ea1NLcBepkAJ55zb2jvmFeI+ZC7CsuQdBpoCK2e/uxlvIEJP
jxD2aW8zmSKuLu6MM8hO7pGBfglgJhbo40J6BrNN3Brm4SYqkYvBhpMoxIHWvQ6S
RpbaB2Pwop6yhm4NIB63dTSMDz2eQCbhMVVN1qQKf6u/HONnBXCWrxxyAL5PZWRF
IQt6YDjIKkRpS40/jnhgCloSXWWi9FjV7M4x0VcsG5HcZv/yVb4Y79jLs0F6jR8S
6sHrJjzHEzhtv6sbGrDuVOi5RSTF5MxMi6e83V440XZFiKNbYjp82qept9LpIaD4
9M/HSi+yLnZgmfkTCe+UCsI6BwEzPwfZXVWR91vSCXK8TOVEE4fWMTvdpn6R7JuF
tqZx8zawZVBDXJ1IdX5NImxz1gxP8zYAO9WWOSf2m59lUzunC6va+ONsDELsV5vO
+R6iATBpHuNuDOZg9I7prqy32UoZB7265f4WHPN7tAVMwsLbm3HEp5s1V3fc1exK
KymXQpIBTcJ0NRWON2K7cmaFHfATKKdbVd/sVx2Q1s/56FJMvZ2KpL1WG6rwzWEs
411jUM/qy4P1HOY3a31Egf8pf6Aidi0yAY0oU28+5wV8W0kB7fbvLb0iYgRngpdI
Bx7dsIUXGU1tvUVjgaxM4zrp90ZqLPdR9dZ4yjr1/M5mMU4LBNZ+SKQ2xdbHepii
xoNqejkIL83V8eqVf36biVp2rTvMIFotk1JVH/vLwlk=
`protect END_PROTECTED
