`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LuIyIQnadMuLVm0IlOxG5L1aeJyCtSvTM+gT8bP8cFGEqx69NVmsi2bJ5JiiUD/I
lDM1EdSQO6M6HeW/A1SmLmrDOKfVuuxQeSzXg4Mky1Y5RnsqC3QuKKRujgUwq2Fa
hNufqLbnxYiA47jkwgdFWIAhvF+Dk2dRUbqHVAVjQq6ILi6GdLfHdxzRr+om4s4G
HFYI20fYUwgiM8WOTKICnLYPAQgEC0gE2CQQBVqzJy6G83boJaZnWYeFWJ7EQPOQ
NfPsieQ4xcwFqn6i/lZQHNxQh8P9uW48uc918zYl7FGucCpM6B7aWGDi65syY6ia
cMwt6VOzT3Kn6xWHZDuSOol8XRM4Mpj4uTqCi6ygjW3RU+qA42iEg1bNN075vKfZ
Z+Ap3bbAeDq0dl/nMbxLwgeRLzNx1UzCJeDivx+DD0glCMJA729yJintULRC7oxo
cPW9/kqdibNlBxJ5L2mZH2L5PLrCCwwrhBRn6EQXlMkbYbM69Vyt5xQNC1tkwxtO
Tdio4z8SWdhVsR2P12/YHbSn9N7XL5qM0kd9geVe90jfXNNH3jiGAgm3YIFIOxPh
q6GYSlLfBAifXvKgHFWU2swxCGwD0XKcseH86ICMzai7+RiO5P7mZpPWiN6bhfOH
7gDDoiYrJ+P0xjDEGzhjw7zkCZstNgMf01MT573iQfy8poWhA6KeKe6yJ6p8Db7G
izwW5SYmec1fiWks0f3JWE3jy63/ePKfRRDRyPtrcq7VoPl10Ng7UIgnXJ/1QhKf
cVo7oglZmqht0F5fORiDSAmeq5xkx1Ak5BuQEBIamnGCNt/2fYhJdnN/NLCMUp7+
UWxXw+EbhqKt49i7TuE4qg==
`protect END_PROTECTED
