`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
a3nvXGSln82l/UR3ArY/qmo3JnsQHkN+1vLUoovt+PfttyLvIOEv+XNXolEQM2VI
sr+Dx6/yONr/ToEJO4rCrCyHsSeFFQeKagj9YbwZM/esTVW8zZI0CCOtkowbCa3u
yKi7aF83LS2u5PbpvsjJZUD31R7ZdDfsAzqkisiNNzjlAJQskYn9CYN3m9LsscMt
UXIVcB3OD+m3RlOxM1qRzL3ceNNG7O/m3+gOC0tgWO8WIz9GDwhJh45F9lW8IiEY
PAESLC8splYI3QLaXAYkQTGxwO2D5mo9njWrFdnmtUzDrjNYC7pQomyBJFjNPvrk
Dn6vRLqoZZnG428piglbfY6vRDlneg6xfGjPfvN243RX67PcophEPzZ6bNNeS7aQ
uT5lqhFgl4QuhvQeonOApgf64vH5WOVA6vXQjYzn+7DtEr7JdvYlDU3awn7GuDPY
mKJUQ/sfJK1yph1WjzAZkEbp37t8A//9scxw+T4TuAxb0NQO9mj9O3IdPvNS/5Vh
xNf6Vn+BOr1/qY6UwCa5jzAiLEPvH/i/vqGYT2JPPoUVPa8v74kCsbHyAuWE51OJ
YMLW61NAFreU5BL7kT4QAWMp3z3+14u0CX/b7fJYLItu+lW5xg6ovJiXfsDyCaga
`protect END_PROTECTED
