`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kxA4F9f93RtwsHfMaY6gvBhibQuFkgrA7qlbJKJonaqovhS/bgophUFC3OGXClQf
R7C1j6CDFJPZcO1f2XpH9SJbXJ5zQT+PxPxWjX3QHtFVmUeF+rNG64zY9RlnJrp4
VOG254wiO8pUxjUZNWjhhxU8+qqqxlBQNZjuhYWcNXztT4sq/HoibW6vQMFtfASH
5pPz3/sZ5X6pM8MI1x9YuVsRSg3hP+teZ83zh+F7qu+vidREUh4ICOiOyx+CGJqI
8AAeGwMW3Y9snUs0lInRsQKrUxPzO8SAS8IVT80s7OWh/6VR2wPF9k7xXR3bkhzZ
/03BS7ipNCzuCG2crZHsu6HPmLu3+5jMkp88PLO0B74StdisXJd+CkblungIFyYL
1jibq2sBnTCMmzLEg0sywKNkiyRnD5zBBbETs6MBTGv65c/Qno2aveSyF8ZTKthS
LMoWqO+r68rEYGK4FowAX0geHGIgU+uayE8AYfcCfT/XiLPzhlbLiTZgjwDmGc7Y
vy2NXxQQizfXlEt/O3KBGOcymK19bgZGE2EndazhLtOBoECXJYW+1jxMH6s+8PoX
eiAJCFM0EuCYMKy67IdS01SvOWVLZDmb5WU3JbvRtNUPvIffO7hoG/ZOo1cET5Hv
zyeWONXYq++O3YwlJY4IrwMox71VRSuXN+eb6VLwdcKeh9ME2Jw/R7OtpQrK43Mu
r7uwY8zR+nvSX1EZifYBmeumWhpdBoo9Md2bwFMkBNu0a5NxPpSZopoEn+BTGDEY
MPY969w8cMeBIkhbsBmXGctHQKAZO72GXleF5TIhrQYxk/9l9wqVT4nCt8pUqjbH
wlc3CQy+nn+gXJnQRVTLTBCOAMLhreqIezGyUdZ8zESbtzKrxjOits7fJ8LSdKs9
pyqRXkPjzgL+o2XRm7/Kqkz3YMGxt0ZgJUhC91eWp88Q7H4UxUTSEaZo7foVg9xA
8SSWRUep0cVLdpTP7FDzf5TLVuOc1+ju2w7GwIPtD1LMgxIEsdAkp6rQB/3s+iWG
VwEB4FIybcoCGqDPaPQ7anmSOb/XIT/oOEX2mDOgrX4AeOmkuYdkB2prtZWBPe1F
dCUBH0mKzM8LeAr0Dsz+zdTsqoGu77oVHN8TILsMIiNdwoD/EMp0IqYhYYSBz7Tz
BwvJEmqdLl+NAUhAxcG/VgMeOQR1srN+UuvsLymqAmTo9uBIypEpupIgXQ1G0D51
rT3ql+89uGfrj1SoLqBVNrzEe46IpKOjtjCCqgACcL8pLBKbllSHowXGpzkZpRMn
Ta1IR2+PJTZyyl6qfY57wmjd64qjBnQPsk4kSnCRjA0Zlve+uLQjSF37fAW3cK6q
BGxp/w68JhIkLMnkzB0Djdtjoqo9vJSsaOAessEGtt3eDtRm/LeBzwZf58y8M+wg
wQpwePXWK+uc+yIHM5QKvDC7AzjMryU6xvMDfLfuWkfEoX1GzEvv8Rr0unv2g/eZ
ng0EPylsyP5EujCiSSW74CoVVMg4xBLL53z/TyKdEtGR4H725f8boBT5oDNQIZqo
aZgUVDKYiOeULq0xA+O6XDzp5NObDQ8i+ZLGuzyLejJqzPGWkkq3jP3cnOe3+p8h
vr2SdJuPKi+Kcq49z4O9o2n45AttBcN7ae0Q/UeZX9dGi7xwg/MjGrmBqXNp71If
XDc8Z4pEhzZXF9s2WxLpuaCKIbivCdNiteelqKlUoEZ2dNuCpYjsakYjhV8YzmHa
HPi/Zoz6uf4/h5p3fiMSe0u6828/lracp71d55rDpU/5QPWIfiz6dghKi+E+CNX3
I924LFwpkydeVwZGns9CTiqgIbjGB2gDTL5nctW/jVPg7fhzq1u4FCY0CKGVkOdc
hFuzW30fi0euR07Da1Cug2OPXTa5GbGxpw8PgoIckVd5Q+itvPFTOxFNJlaoA4hq
CphydGVb+6EHmOF9V9bJWfx1xAxAJrZhEIgEQK5PXC21VvCZVQ6g3/ueFSb9XvGA
5SMeccPEmzeKmc2q+RSM7rqEP4y1X//myZ9s3cy64sZVBAKHOC24oLZreXfigU+l
lPmioZEVIPO3ikoZxTZMa/M6JoHe5mIOtyg/Vw6E7DIrFbOMHT3qm2Ur/CCoNTCj
qaTRNV2K7T4yXXnDIzzpYuuNg7/AztsqWJXysoVUMDyCptlx76/Rc2FwKUpgFbCT
Ho07QhwCGqOoDb+pIFrUjqJwyolj7RdEtKMmLmD9yy+8qmJwwvRpOKzP5KknuE2E
AyOcuCTQWGsINJ8uFZUJklN9fdCo7iuFVVlsPI9QzRauWrK1hUphQ59qBVl7WEkc
DOh5arXhAYeIXNzjIux3g11yta+Nki0itoycwLDZ1rAUBFui+CX8ckKtvVzjCQ15
jdZZbdI1+g2eHMxRQ7baXddh8ZoE22Gu6RlflDCtp6t/MIauOosrYyZInRKNmZRW
zwX582jVg84YUdv7CMqKi2LOoJeu3PduYsLnY/WWQh/NputWjzN1nyw3jNn2mn4n
JA+EhR3QxaGehklla/OymEnngbzApFpWMbKRK2DXGHVCEzd9D9fCVXtgepbZyvw3
2kw8S9cm4XE4TfRJKd0HbLfoRqkVEkFdZwCUsBZ9APWZcJip25klFW02hd8DzmUP
ok38HqzhKqso6gY5ErFAhlbw+iYhXrRKY/oHFNZPxDCxDB7UOpsNB4tmqr4zECs+
1xRLrEi57pkAx8zeAiNcdrxgp6YOj0YJ/yQMC/vhQkAV33sh7LoljfxuOBlgeH1B
xlfQqioctzIYz46p7BCWeIwWvUrKiWV6o+2lHyA+k0EmkPtcg5nT7UZOgmbzR8kD
YYJh9o8YhiCUaRxh9pG/Xupqsefut3USGkRvFYcuWIqyv9KgLA9wqDcfGYz/cfvj
5vlj0LEyJkq9Nppxho+uLBe8+YkAjfuKE3N2U1FSMjvSLZUgzKhES2qhCbCCbRoT
mzXGULsuptBy6tl26AvSiuiBhRO+XsADaax60A7KPvG+8u60FwEXFbBqUXn+O0Bl
0G36Yu1/zxHF8xB4GvTWDlPwgzJ1gA3Am0eCqwtOZcGiUshrhi5ieo62XBdZsFkj
WstLEreAGqCCDZCcAh7j/OgvzGDsMrxyfCo8eTUScH5J07aYwBhCATG201fluDSf
psEM3VRU55mKoNnhkvxNMUsWKLupxUllATra0lGFr0Dvyax3x1bOzclN4esB5zSf
lakXk/T5Zgek3hqdE/jJbbUDlghDHa3V+6RMFrs3IMjaIMTXk4ezScL5ZUDoEteh
odMG5/LDYREHagvSTrOcF0V9ZJSbmPdA3CrAjRH4JHJxel2tRdvjDS3YUcokcFdT
DTjzOF0HshzJNWc67YTSm72/b3KLeMsfxsbiBqZCDgVbkxA9riY2HrW+ayiZ3GWA
iirdEfhDMxaDfeWX+tEZ7VkjLsiuzBMJb/kSfw4DIXsbkO0VIADKdgQcB2gzhnRl
M5sLh4h6WRYo3nmM+aj8ADUStZCIy9mikGsM3JViYsidlBTY3HS/EaSbXrIHxcoD
3RT/EWXvKr4wMFZZEv8Vg7mzCA1sqUYUQAm7Wf/3stWdyWiZATA/XAem+Rhxo2VB
J8PCfRjgAAEuFh9nLAlA09u9FKhFu6YkDP7wdALbYNTYOJ4UtHnpdNy6RSyNGZmu
DjdWg1VwSXFSruhtkcMKpASX2WPI0dyZKIhMNCGIX8aoqvsT52NJ7ZE5S89P1lvs
hDZ/A0Q1v2Ph6HVSH0Sn1tCLg1y6aO+WOzcHncxbviKeb5hlN3aEzYGtKqID41sU
cS2seccnaUB4Qm5T7Mb/BLn9bmrlvGTDk2F6gIc6BwNkgg8NGjdwVy7M+sM4e1Q2
vBLSeiXwtau8oll7SK4XQXobzccq4vGPcr1GkBb6EAFd38xu5pLnwDBqS2TNuEzl
F4Qg7Rzu1qf+5yhPnvIBYL6kYZuF58N7jzVP5TCXs/7nfcyPgqZ+5KYqLW1eyc7w
JBtR7jjTtyXgsfK3FY0uwNTAOGVqcTqsA9ItXioBmsXEoJHYNRdJkgrsCJXyjD5N
cVCzSe3PsK5Y5Zss/vTiKM5guHUOJKgXZIl/Sn/MwKnmJu3oWV4ALzuUDNnw0Mk2
GBu1GAzVMXFAlsuro/xHkX2daY30GCs2GEvw0UcIirX80DmOKzq5aq+/IxSrKIuP
vTempXFqSBNh3vv6glfopXYoTpG7HS/3kgTLMYVDSeR8fjSMZvUiDzIVL7sRrtCa
q8jOeqUq09+o6P00UX7T10nDCclIYf0FR0g7lI6EDr/HhDTgMMm1mW1R3J0bMLhI
YN5VFb60CkVc1Is8pm+qu1bNsc9hNVrJbCwzdkZXQgLaE7yyka1gphTqZmd8bbw5
VNrfdqTgQjPdLusZgIZ9lydrnbltoHi3H/+tCqSAwH0zYRfnmp3FOv79V3R4GVlG
QytY7Hw0dfIV3R4gl807TqZYPIISKqbIR4VrjyRtHKTJSUf4lHCSsZ8eiCLXR7lu
gtbseJSUYJG3unRojmxehmPneadmOY6qWEV1cX1yv7qNgebJFjL/yxsRJ0cUFCEi
nhblTI0P9XikqvFWNE1SZ4QbZe5QyrXp34uzZGbyKscx2WtRUQj0ZVISOJqZf/P9
0/HXvmga5TPEt3383QCfGBCDvv1WWNGDc0Zt2a1vAwFbGPYohzkrS9JEKZ/EBEG6
OcQePJRc0lJ+IST2RRJ0nIPvxcpU3GNj94lyA1fPu4IPVomHzW2McLjzevH+t0ri
IBAGWkHlI2wzQXy0LFPdta9roGUnzDNJYtHxOyOsXjjbS4wBdnBHIiIIyfD19fJx
jyZN5fefgkbJI1399uj2IFTRHA4EjPqienSsmyTYI8gSU2pJKNIDNEMDaniHdOJq
yFrlWFIE2UXe0yECXX3JSue8nbOM4DtXczdLOQlmxNXabT3PKP4KnLcphT30MJm8
qfnWf9FnR9oYLSdshdGkqzPbrlEkj04BpEo2jDC4dE1h4Rf42JAQdz3xBX8X3y79
40Iy+Nws0IrqO9FpUohSkxmuxN547fJISUNFq6lLqcCDG6dDywJzVakoOeWnpIEK
2a4YaItncU3uWbPCIUPvn2vvQr0DPKMCViCcnwGN3uCA+FXoh6Iyyv1ZcQLhah0j
wSw5kojZ+1S2OQ7VXUsh12IBV74scdwSv0hxpK7fukdMSOMoBGRXvtk5KGwdWWNS
G7ruAiMgt5SLp0ivQGtIYe618TTcqonbDBLF/I6dNjQQoBuquzvx1VNCa2gdPubj
/TVjHFfJhzb/AEy/c42/lQXGGjlAXvbYFgAaOoPZoN+zzp6hZpqkNfsfqerq+Bji
Nbd/ykZET9DZ3WBELGxtex9BgaSvFTK817fH/Lbz3F80xZQ53QLpWBcPFUbg9gHz
it4FYujjQTGf7nW7Nu4wHfib0FYARQgQbq7oEtalunarha3CtJ7ObZVkdRqQMwZW
I35Ulu3p6MoItnhZ2QSaC3KXuQCGASgAVmXuDgf5s3jL0tJ6Xzwoqc/l8VbKufyu
3uxd5hOva1sm5BoFGr8Z6YbLT7MfzWqAd3vatkwoqfKWwKUOyYTPdJHrnIlDSvDi
kNFwpEd5ZcwpWFTVHj3Ohi7Ung7zji8WcmP0j418UKQRiDmbdv7b7QNJIRGiRzeh
M6FMrED3w40ku023d64qvy4b1S7gcEcRNuufrdgU2DODuDbYDplCHTx1zj49Uhfw
vsUXMRl41vPtq/ib4WNPpFPVUvP1MgXMU4D1PuPiG/gaL61aBLJnaMJhdOYwfeCT
D6C65aWLuO+YndWVtBcRIzrgHhzBTNchp4UWmXG/zY/AXJ+qhS7ux9+yV8SmH8qD
aZFMvqQGT0CquMHqtbXhp1RQ8Boi1HhpLqqA90eCW34EMnmKnxFJ6yZtT6GtS1YK
Fj9OhfZ3snLnC/1LU7L45ENDTHdgeQ7JZEO6VQL1Q+fduzsQh6CyY/EcDT8lSS8E
R/oQMsv4sk9BhY+clwIo3p0dIvckr4ahOEy+Vaer+e/pSs+Jk8mG+vLiwDwouOtC
ejpiM8HfF4OXlrwYsrhcHLbZY7XaRmDy0UKp3eho58szQmDLg6i2BTYeUSFD5wKF
9FAI3TgUlXo2jW3lrKPOpgpuYPNp/TH//SWckIPP9DCY69CqCvw/p2ZPtOTSNWbJ
X4JUS3y8HoISedy6e13hl11EusjEApiYRsp6inp7E3d+yOazmq1xihEzOFGDssb2
ji+t+LVYtT6hV18byvs8RXinXUAEwOnMW7frpkBSy7cnMjro4O1gsuQe/vRC88+H
+DQjx24GHfHo+tqawhVRMVC7f1BtPQD8nwfONj+xZ7H/Hb5q3ny60w2LQTOIcXzx
bC+dNRgwoxHSbKHAtQnobzr+MOTICm6lnw89UNi7ZWdJ/VseYeJlw6U1HUjkxrCu
E3Xxr2PeKDAo/tAKBWnj7nCawffaQ0OGo8yY9B/4S7OYwaD/XhezktQTQkpR0VI1
iHjP1T2gc9pMQstrttUxDMn7fAyELRKHVGnzlQ3zmOPwSjQMHWwpHkAN+kByNcYB
kuwsmkODzzb3ehxGZgANHCd88HCXfrqzSrdEnAdeGDiT1sg6DhNk6LgKwLEJamJf
pOdowbEvx1+eAwmyVxpVcmkAqsOp931jLrqWu0RnyNodJEMDVzw+m93rsoLk651R
Kugw6SNSZiN4bGfMA7iAhgFaQVKwk8cRIHao7Ky+TcqY8RPzl9MVsP8wDFl1hz1d
O7ThnftkuRtNbuoDQuse/ThuTSxh+qJX00/Z3H0SE61KkxkZ3OYIi3kY0i2s1kKz
jtmhNxymMPry5F7yxgkqrrH9j0E81tfTJUOrIGgDnGjPlFIy5H4cRmEJZ5rhgdF0
pLpZ0nMVpyHoT3IOpe7lIqYhqv/nrVRyDeaQWoq3d2RS2t1/RMucoV842XpGrK4e
hzUgHBHQO6E5BUhNtfpD/2wfPKcLkyraKjfy0aaoqJ+KV/glS2cYVcokM6uOwg72
aI76yiBsXeXpFkWtRUkovsHZq+NPyIH6sTz8mhPnR/sEESljSmuYa7epWlhs6Xdr
vyUCHgypIsx0PePhRc/2MdnL6aSgHWe/WMdSLwBCfRsgAFVd2bvkmMvWE2Z9txOV
3ebe+T0LDispRN3mBUdkbPgBZgQtpSeR7yaGjahe0SgdAEQnFNXL2BD3C8HCTOr5
XPbysqsFpb+XOR228TX+2HbiOHp357sjOk6gr3t+LP75oMU83MbPZhi2LYf8/+Kb
8Qa2oapW3nT4sqhojboKXH2DZ1aLflX1T/3ywr9x42x0VyCU0WN6enuHYoRKmz/u
59UKWOqeU0NiXKmOy+w7WGBTCZUPBYQbnCVsDAP1F2otQDSJyBIf0bPQnZTQsz5j
da4cvmJCl/YVijVfl/asZ35zKH9R0cXjITGfKIBgnqzxcfUizBTp+toVQaDbuaob
zH43pj/B+dJYGh4gyx5a2z966Sibu6pefOdzXGyYc80OpDbZ0jUdbXEFMswKtFEt
AIXKOTbK1mWUD1/I8NFgW+d1BTxUpTN0BmhuSnXVw7bFbwQlDHC5OZ9jrd9VAPZL
nFGa7/NUa4+lMuhYD1if3IA/m8AVv4R3ev8k6LSMI/Kg2u/0lNaNlEdkPxcXW6BG
7Q9UjlYIo86mulDnKnCqtbCxutb2nNSR6sF7CS3uL4KYGjlQMY5FodLkbZjKTN5S
wQGPmzL6EgmK7U6u7r9lzRy6mDajLHokVmGMbZURHxPzFXGL/2eQ99umpvT11Tjm
ehSaZcnZ7nabW3tz+obNtuVOKHIvSjTQiaSGxeh7uNXiJmU4Blygoe/qFWuN9w4o
Vdkwd7JYDgpTxauX8u462lha3gt+vpumAGQ69u0IrsyLw7p8Lw+iZPcfYc5xkKcU
8BR9ecVee7m7Z58y6UQZtnB1/JUVjGMN4+Lz3lXrnGbtXbaumVI+7CsmnDAi7xjY
2ak//Dfz2qd/qRSOlfa055r4BjMIIvly4tzbuB8hsDv1D9Bb7YZlJ3pJ7I3UIG71
eySEWne37I18jnrZx61EYcZy5/wAAzbglTVgwU285faXG9cEQY/FeDP6Qjx8srzb
EiMTPtAPNQlowJJgXcSSEzJVCQpoJA9hETJD8bqpLw7OwB7nox6lP2aEb/OdYOqZ
np/GlzpsKHYdD+2mctauWx+I12dgiG4K5E51vM1xDshQxJyRjsSS3ic1A+x6l+/h
dR+RDwLKu1awsLmPmjv7epuhCpksN0O1GLXAeQk6zZRP/V+cYf/JTvqgHUEjuVrv
15FUE99noVtClSgbeht1ag+wk1J5PuaG7iLGTHd7QlpQ8wf5/HFsXizikG3pA/D3
U3SJlfu2Vl8EJmAIW+JpKYptgjFlMSYnjN+OY09/G30oDSa/brujGmQg2Tv7XnDW
lHgzypMbgRmVpI1iE1jcuvJlGwEyOphZfO//kwz6JxW7J0Czrsq/S6t889XK57PV
iryXzuHmt6WkGOhVy34tG1e7xWZzisiZW0uCrYjhq9lFKELU+fL4USluVGxrVny8
VFRTL1NQFVxuxRq5kDXuoZkxQxiK1LVNsMCb0YL2EZqj3epmcKVu+ea0d9UxU6zh
vsxLh11MIp4CgM5N97I3UNtuuXe5YJ40ns+KKjdszs3DBCQqeRkanwrr6OMPsQzp
V8TJ506XgBRDmgMCN1YUHkqJlvxKn7M3qaV3/LK+WrPjejZMFVIlZhoNLEOL7hra
3hz7FxIp6osifIMjXf4/Qqklvtxdp7iVqEFB1yyYmhorY4R+GppiMlZX71ix16EI
cqOfR3o1k/1lC9We4POYCA2+/pmeAjivddU2IgG+23o3uDBtVt+5zk7Q/PBF72st
/Zutp/72//PXiXRJYa0nDkDM4c6x21c2CgDIfjc4yr7kCy4eXN2oTM4vmp61HrU4
ox5KLHQEI+VX8MZag54JrdOTZ70d1rx9ADXC5BRDYaPOVNDIku1YixvTUckfs0eE
ceG+zsodrK3dZbk6nbFOL+kvv80Qs8THlMB0bYoSn7pLQ3Bf003SsscANowme666
c42gZZxKbnuSVyggmLBq0gjFK9ZVWx11zHwjKcaBlfKgFz0jXfrMLAcUXiHZ9ipW
tpbY6EMASjAzH2u13NiN2i8zGuxRJdNZwwWh4ezmAeQkNPVoQwDRhLqQ/hp9T7TU
uPEg5PcSoEgfx2eUG76iL+zf5GvJP3y5s205oOonfirNsPbPzPgb5NhsKUoYbFPW
PeYdK365anxv48NNJebo3gbk4BpS8ZQv7jYV604fbm8MZK25aVa65QQdwjVyMvhM
FKrsvHLxSBjQQmuI4f4cxeUWrRCe5ZS+cBGhTv+6/A67L3hylJqd/gOqoKaljnDO
ESJ4XlohVEN4BQXZ3qyRmvJg8jqNfp29qLGCbLmr1coXbc8gtQoTTuEMYEMstTyh
`protect END_PROTECTED
