library verilog;
use verilog.vl_types.all;
entity arriav_hssi_pma_int is
    generic(
        enable_debug_info: string  := "false";
        channel_number  : integer := 0;
        avmm_group_channel_index: integer := 0;
        use_default_base_address: string  := "true";
        user_base_address: integer := 0;
        cvp_mode        : string  := "cvp_mode_off";
        early_eios_sel  : string  := "pcs_early_eios";
        ffclk_enable    : string  := "ffclk_off";
        iqtxrxclk_a_sel : string  := "tristage_outa";
        iqtxrxclk_b_sel : string  := "tristage_outb";
        ltr_sel         : string  := "pcs_ltr";
        pcie_switch_sel : string  := "pcs_pcie_switch_sw";
        pclk_0_clk_sel  : string  := "pclk_0_power_down";
        pclk_1_clk_sel  : string  := "pclk_1_power_down";
        tx_elec_idle_sel: string  := "pcs_tx_elec_idle";
        txdetectrx_sel  : string  := "pcs_txdetectrx"
    );
    port(
        bslip           : in     vl_logic_vector(0 downto 0);
        ccrurstb        : in     vl_logic_vector(0 downto 0);
        cearlyeios      : in     vl_logic_vector(0 downto 0);
        clkdivrxi       : in     vl_logic_vector(0 downto 0);
        clkdivtxi       : in     vl_logic_vector(0 downto 0);
        clklowi         : in     vl_logic_vector(0 downto 0);
        cltd            : in     vl_logic_vector(0 downto 0);
        cltr            : in     vl_logic_vector(0 downto 0);
        cpcieswitch     : in     vl_logic_vector(0 downto 0);
        crslpbk         : in     vl_logic_vector(0 downto 0);
        ctxdetectrx     : in     vl_logic_vector(0 downto 0);
        ctxelecidle     : in     vl_logic_vector(0 downto 0);
        ctxpmarstb      : in     vl_logic_vector(0 downto 0);
        earlyeios       : in     vl_logic_vector(0 downto 0);
        frefi           : in     vl_logic_vector(0 downto 0);
        hclkpcsi        : in     vl_logic_vector(0 downto 0);
        icoeff          : in     vl_logic_vector(11 downto 0);
        ltr             : in     vl_logic_vector(0 downto 0);
        pcieswdonei     : in     vl_logic_vector(0 downto 0);
        pcieswitch      : in     vl_logic_vector(0 downto 0);
        pcsrxclkout     : in     vl_logic_vector(0 downto 0);
        pcstxclkout     : in     vl_logic_vector(0 downto 0);
        pfdmodelocki    : in     vl_logic_vector(0 downto 0);
        pldclk          : in     vl_logic_vector(0 downto 0);
        ppmlock         : in     vl_logic_vector(0 downto 0);
        rxdetclk        : in     vl_logic_vector(0 downto 0);
        rxdetectvalidi  : in     vl_logic_vector(0 downto 0);
        rxfoundi        : in     vl_logic_vector(0 downto 0);
        rxplllocki      : in     vl_logic_vector(0 downto 0);
        rxpmarstb       : in     vl_logic_vector(0 downto 0);
        sdi             : in     vl_logic_vector(0 downto 0);
        testbusi        : in     vl_logic_vector(7 downto 0);
        testsel         : in     vl_logic_vector(3 downto 0);
        txdetectrx      : in     vl_logic_vector(0 downto 0);
        txelecidle      : in     vl_logic_vector(0 downto 0);
        bslipo          : out    vl_logic_vector(0 downto 0);
        clklow          : out    vl_logic_vector(0 downto 0);
        cpcieswdone     : out    vl_logic_vector(0 downto 0);
        cpclk           : out    vl_logic_vector(1 downto 0);
        cpfdmodelock    : out    vl_logic_vector(0 downto 0);
        crurstbo        : out    vl_logic_vector(0 downto 0);
        crxdetectvalid  : out    vl_logic_vector(0 downto 0);
        crxfound        : out    vl_logic_vector(0 downto 0);
        crxplllock      : out    vl_logic_vector(0 downto 0);
        csd             : out    vl_logic_vector(0 downto 0);
        earlyeioso      : out    vl_logic_vector(0 downto 0);
        fref            : out    vl_logic_vector(0 downto 0);
        hclkpcs         : out    vl_logic_vector(0 downto 0);
        icoeffo         : out    vl_logic_vector(11 downto 0);
        iqtxrxclka      : out    vl_logic_vector(0 downto 0);
        iqtxrxclkb      : out    vl_logic_vector(0 downto 0);
        ltdo            : out    vl_logic_vector(0 downto 0);
        ltro            : out    vl_logic_vector(0 downto 0);
        pcieswdone      : out    vl_logic_vector(0 downto 0);
        pcieswitcho     : out    vl_logic_vector(0 downto 0);
        pfdmodelock     : out    vl_logic_vector(0 downto 0);
        pldclko         : out    vl_logic_vector(0 downto 0);
        ppmlocko        : out    vl_logic_vector(0 downto 0);
        rxdetclko       : out    vl_logic_vector(0 downto 0);
        rxdetectvalid   : out    vl_logic_vector(0 downto 0);
        rxfound         : out    vl_logic_vector(0 downto 0);
        rxplllock       : out    vl_logic_vector(0 downto 0);
        rxpmarstbo      : out    vl_logic_vector(0 downto 0);
        sd              : out    vl_logic_vector(0 downto 0);
        slpbko          : out    vl_logic_vector(0 downto 0);
        testbus         : out    vl_logic_vector(7 downto 0);
        testselo        : out    vl_logic_vector(3 downto 0);
        txdetectrxo     : out    vl_logic_vector(0 downto 0);
        txelecidleo     : out    vl_logic_vector(0 downto 0);
        txpmarstbo      : out    vl_logic_vector(0 downto 0);
        avmmrstn        : in     vl_logic_vector(0 downto 0);
        avmmclk         : in     vl_logic_vector(0 downto 0);
        avmmwrite       : in     vl_logic_vector(0 downto 0);
        avmmread        : in     vl_logic_vector(0 downto 0);
        avmmbyteen      : in     vl_logic_vector(1 downto 0);
        avmmaddress     : in     vl_logic_vector(10 downto 0);
        avmmwritedata   : in     vl_logic_vector(15 downto 0);
        avmmreaddata    : out    vl_logic_vector(15 downto 0);
        blockselect     : out    vl_logic_vector(0 downto 0)
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of enable_debug_info : constant is 1;
    attribute mti_svvh_generic_type of channel_number : constant is 1;
    attribute mti_svvh_generic_type of avmm_group_channel_index : constant is 1;
    attribute mti_svvh_generic_type of use_default_base_address : constant is 1;
    attribute mti_svvh_generic_type of user_base_address : constant is 1;
    attribute mti_svvh_generic_type of cvp_mode : constant is 1;
    attribute mti_svvh_generic_type of early_eios_sel : constant is 1;
    attribute mti_svvh_generic_type of ffclk_enable : constant is 1;
    attribute mti_svvh_generic_type of iqtxrxclk_a_sel : constant is 1;
    attribute mti_svvh_generic_type of iqtxrxclk_b_sel : constant is 1;
    attribute mti_svvh_generic_type of ltr_sel : constant is 1;
    attribute mti_svvh_generic_type of pcie_switch_sel : constant is 1;
    attribute mti_svvh_generic_type of pclk_0_clk_sel : constant is 1;
    attribute mti_svvh_generic_type of pclk_1_clk_sel : constant is 1;
    attribute mti_svvh_generic_type of tx_elec_idle_sel : constant is 1;
    attribute mti_svvh_generic_type of txdetectrx_sel : constant is 1;
end arriav_hssi_pma_int;
