`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yBmTTXejaxaIxkFNOGfIJBmgT0az3WM/620Bm0pcU0nV6nRi1UVnC2uuprv5U6i5
8LGZG9YO33zBr2zut4sOdopHaGMZVSTypcozmJ+S/CWp6sP574/71A4l8BfM1J8U
/5oMA6JNH4SwnRDG0ATT6eq8/mIN6KN0YLR8VE1W5XJG+g4weFNq1KAGrr2j0MtX
+IMK/rwx7lzuRag91hLJsdPv2RtIOoGsZc7xeJddkJZbA4yiNH+q66DUSB7EbMg/
uz0ogV2Hy2kso5dWXguydZzo9PE1X76FcJ+ZpnNmFhg/qprONYZFo2mdtDnwzLUA
UQjUSK6L5ms6qm9GZAXSHaQDoc8zuBDyWO+qU0fLxcp8PabtKLc1AJ2a2DG0WMLi
reOg3Khq3ZHJbX8T1SMRDngHBvMikR9G2IXi+qx9xZ6guOj/LLUgSA1PwAzvoesc
UVXKAm9lKuapoW6ih2b9/bv2IPoqSlg+9c3Js2l7MN7N6b5wBYPDLlE6qLiIzJHs
AKq2vuwrvrJKaHUXYXgkwEkOLtGLa1Cgm7LvacrAefdC08pTwu5643pi8BlLgF/z
JTew/qVNWGCe5tVB6r3RcB9lnjkkk2/PCSZ5QZqXQ83k+mA6H+/vVV/85jnPaQXw
vvJYHYwDkftETnXQFtRrHUJCb5CogsCnvojqvjgmk4q/pylgbKv4mlbf8RXdBJHE
VO9f99Dk23fZBSkrxqKm0o9FgOou9ZNDWFOJt2uxFD6ucyPtJA4RVNmd4tjiSz45
GTf0AD8qHcOncAFCKoLSNAjJNfGV3GPeDoEM5j/7dEZh37sM3/qv6bH2eZxIQ1K1
MK0ef8I6Eadi0/wDvUr2mPXp7vq5WZ/n563i/+U/DEHIiD1VVq4h5ErBnMBI0sHT
K7nY2iS2XgWKujqJzpsbjsQ915XWLbncDZQYQtpt6tqQmt15RcY3xlLPFOnUdulq
YSS6+YNLB4kTJJ18gK3fnHK0wosXjSLqNDEvVFDCeM/SaVdYE72MhzSXTinWv7lj
bKffdKlCEsJDKoDz2mZJ+1apbYJp9p461Zt7NnLDP0h1D0GhF2J37oqfJM3vmrV4
abxJw4XetwvWSlr8YsZdBpf1f+2XLOgEBBeZoHEeqndZM8sRsNoBnOQICRy9sY6v
YW8JsXjb+DqoucEM56bqdyuq3CybmTHML6E1oPWKwaVtke3ju6rD8qyYiqVfqcvU
monV3ujcKk+eIn6JyKj9YgIzBfWV/hzO9SdJmyIR9L+Cqaz5OMaiao7uv0hhyGWE
Hg/KhV95odcnRRro+syTRdakYSaYC3L5icpUsPD/pWN2DzjCMjyJrH6eoH9FKkRn
TIGiB8Q4Kfh9RJra8+xln0BiC1LME8OB6oB4ikawcGgkQ5v592cYH+K5wOS1iw9I
LMZlAgxxh7vHHwj4VMuI9REoGVx/PEfrjag/DJqJXYBm53KgEqgL+JhkMUKkBf+Z
6V21FN38w/DdqVmT+bjaW9Gn21pYTdiM1cPnpZsb2eaZfZeH7oJyapm4An/G6WF1
fWtIz9kF7WEJalHbA/cXcFNnbHlQ8BJZYE/qTgMA9SSbf9z3hYikAM+3YAxpn5mx
KfDd4TludOeu6s4aj3iPy3Md7gh/oHwE0ibX5DiW0ohqVGTLLf0eB6V4X6YxZpHK
c2z2UBF+sb0B7eZGQdnnhpCXUN02PRX0nw+feWFaGxirGJuHH/f7UJnAMLA+WLMe
h5JN6mGYo8qJLRqZMBWOAo2eGEeBviIGj/MyhoHokUDPGK6eptlIokaOe2oqY/F0
9Ei92OtM9VJJvf/yn9WQudzYhgCspoh+BFDr3W+fMPUUJ6/ao1/3ZmZg8e4Pp8gc
PVhCGEyztsQUtgxQnC3/EeaWV5CQOl01RaEcpAx+NqhAcmb6Y5kFF4kqE/sK6HAE
AeYcRfFDwLuBm6S8XcWPbw72hC9d5fCUfVEqAXHNcsa+qqmAXc1LkL81nSuIbm61
mSC2hEt4x2UxiI7QQsjQS714xmHTyjtzPt6v8oDQqBg01PkHXb58DiRcS7bBKcox
vbw1Ws8Phv1Pcwnqjb8rRTnZMDjmfSXHiukE+4IcoS8rBH0gIKWMa2qZXWF2HrnS
uHbwfBWgLzkEaN9XeJ6bsQzBZDW2VHT8bVJXrXlDfmme9k4txUXJSCrYe9HgUYn+
Ewt5iQ6HO2YY5+uEOe93aDlP290ZdlCLFCgFtMmYCNIrF8un4QOd54YC03DIjnop
ZFzADG5/YG69caiCkQFOkB3sZ4Itcmtfoxw6lpUN633PBG9X6QikbmEe/Olboc6U
fIiPAneDtjCLeg3uQG7O0Z5hIk/S/BAkWl2SQaGBkTDhbm+Vdfyvnr/rqxEqh8ka
hHTnYSRtWggX8TrqorOgRepfy/zmx5EQDzr25i0JoMBjAPtSWUCBPiF1wesIxJya
+M1NtpCfimRykwVDxFp/s1r90MwQKCTGWq/ApznUFoenDtqXspL04XYFebjAlcHW
4AAnNzhk4a+gb2k7yvcqjpe53xTE5SITdYXqoYPWu0JH6+rZ8hUeWkpqIdTWiY45
i9LGB1X++njxawzDQ4UsCtRZfk48DTnevm1PGwwrohWCTiZtoppi9ALqHT9n+9bz
DaUsk6M9p2zgE3yUt9mOr/NR8k3IQ3n+vstqHxY8LHEI3CZJ6BJ922oOXm27fVU7
K95T5JKwhkK5LynHhu8dspGux+DGngfT9rjCrfzCMyAynWySJkpjTE7fGPkjLWyD
6dsvWohWi+lKLUxEWI0WwVNhYfcGzmKAwgptqMGB4JRomfleXB1+SiGTJCj7HrHa
15RmuJMP9Idzc6WGCUUAYdIYW6PGbdTGGOQuxJBz4i1SP8JKEqaGjr2HIlDD3A33
gv2RIDFeVCPQGfN195XWgjPxxgoo/PbVfgZqVQQ4Ua7bko+GQRp5BTdDRDwbuwO5
svtFggXJSgLm0+r5vbil6h7rEBrz21f9afw0RR3bLFrITIvnE6Twxj6ZO/ZcluEq
x2IMaWpRfMgLHbK3Nh3QWkbevf1+F2zGj3eNZI5TaibnLYaCWnYJujHV6pxX8toZ
SmILceecJTVSFlklEyIKK8EcpfSuhG49d2DWMZKx7gFOQm/tO2YHimue79jhZfmA
JjdnZZ+Be/WV8mxJ06HbL6vwZxKJNPYD4RCSXdFUova02HvjxMSB1JOT6NhehM0e
mA+t1/CpIz2WOUWNbebWVi7i1EfWso6CmspalNofL4dOOKHr0qqox+HOpDqsFFJc
ug9DoMl1JbYTY5yreKMxYJGXbEpIkrSL6ObET8DOTfYNvmIOCODecPREECZTHeQF
XnIx8rwOtOIxhP12BH0xVRabqyxX9HnlkA7mM6T0At/VwVfcH6SZnntETRS7KGGN
FuBPHvK6wPkWrACE70hVhqTRJWr9qr/mg33iDRdYs7qjDpVdNyT3aLwgEJTRhya9
s6z3pMJKcwHqnLUOdd8AWq2eL+3RK7QUDnBgCS9uaEE8NSEqIBpFaTWE9byt6jTd
VEJqgTaYno7TVH0V+DCwxf7DSwJ+7vXQNmLauW97HO5NMCI5scpmusaRe4CMRfK4
t0spDVLuMrWXCj3qSkkTyYh0sjoA51Nv4a/AwEkf4s9sidSMktVLDXcDYRba8Te/
LPeN8oNnazmCQRyrB9xSCq8eRbfmF6o0AajVk0BHg4exf2xiemW7VKGsCQII/bh7
Rrdy5YF3HR8qmpzONM1IfwRQW+HoJtDNc2pKZfylrBsNkYuCEwb1eM2I3jrhoEk7
A58wl50iR5RIc7p3n7jzVxHMiW6f1h0FP+99OCUcefIYsTG8+U0tBrcMXdChGp02
vNQSjN8ZdvyizCVj5W7SQNb3XR9KFwfEzj25ZqQTvPNdiAcSuFl4GSICL2acyBE4
LDnTG03Lp59Aj9XZ/no+lyziwh29XyQt2f7fgmrrvDYvE9JXr5U0eTssOyiygXzn
vVJmlwtCmJuDN0T+JWpXAA0GTc9aB+C9N/vuAADANKfPZGSwRyB3MqAVfU4SHzrg
FSIeCIirZmR6X3CdCRXSxOwOD62TQ2RRpYbzzB4ORlgnR0zbD5WUgejSvBXkfuQY
HeYPGqi/NiAfWzPOoGfyqgNf4lWoMs5AGUZxMnGt9LbYTms96RMYXHGrfI4hqftS
hBpff1laiXsLxkFzk16chSBtcjdDm9hdaytF+OhmQ0Z5gtZUwCw5QHc9FrTdHGP2
VfogQTuxL4qXqKCiQYn+hLRcj82XN3y3hsueC0aJK1qC7QTLr2HR/Np258aJMxO+
0Fj8pI21w5puzPBO7d6myDoMyE/MOdkdPgqtoSbBFUcivoWIeL2l4MspuyjAGehR
T+rkL1h306bJ74NZectZReUMHUsvCxtXarJk1Tqz2yefvxPsSD5r7N+2+klXQTkX
YFM4GFysGjX5dcF+EFqteEEOnthbkm+svN3BFmQYALulWsIFEQ/129qSxbq9ST+4
lXdDzesR5FF1uI6KvvEgARb3PmZFPcEYEimLS4L0IlX4QNtqk2X71gzOhrrpsk81
bsKpNnXa/2G6GC6ljeynaGG3CgvCk6KexuCXLvXCVefb3qxr00a9ek7UqwNjUHr7
Ig93b/ne7TBWsxcm2k8pcBufG0dqeswZTKrUTBnC+Ovg5a2f7YGs+e+DyZhKkeyu
usLGplg5NGtufiLcXxHVbQOfMCdLOTivJ5vYPCg8c0k72VbgAOKjqU0oIPJfyCFE
902n8Bn3qsGk8ahFDNfQ4jJtVuut5LJGKZCXclG6hmN6skOxfVhYxinlFS9kcLAv
L2b95y4EWrhQXqzp5896L3EU7wcbMHIaxZ+pFjAFVG/e729cAWdVQzWdMedFYqTS
1iZDT3hhDCo+YmVTznocS2I8i04Qg9SdO/2rik3dsgHcwW8PYxya3XPdbTW1n+ht
k6KSYVl6WPo7KVpDsbLt2gnGJqL9mR0NNu9iXhyEWrJyNe/2q9xhN5raU+iz2vAr
/7yJEN13BME4O8VttXtzzDo9BOglI3xhY/3B/dxE3/6MdVMNzWKF+mPTiaxRUhz1
Mle/jmi5K+IL431odBti7xjCngmOOX4VhNTcUY4w8ArfNQl6J3cVDe0jpY28NFzh
vo5nqjJUxBDekH0VnoMdYF6yOOvvqUkBUnX59sHFEq3IJRJb7iUWNq6ITEJrVixD
bILFGjjJH2SR6d7+06z0mvTLFDdkhaxoCO+Bcx+UcDgqDIgF/TJ1t49/anpP17XU
CwbxQrazA9Vd7dMAaBOGHt77Hwylbzo1zlhwcEAwGrAkCdogxJkIW4xJ/3aiqI9i
/9gDCMDv/05P9/WRipl6N6am6sP9ZB57fmIOvdtBB9z/4tkrELVSJUoOlkSbw0u3
IY9JPfHAkuclv/75idD+SU6z/qjlE2LwrzwhRQFirJ7IzC7jWlLZI/brzhHLW4t3
6FH4dZXaS94pR9eYf8hFRn/CEgbxJdKUTGnI0zGaQd41IlfqcHiujJsiGeLOWB5F
BSYPvOAwHet1om+pD8/kIlyARbu0gOUmEqSCRM01f/nMO+nbCNBy1RvUMRfTtZ2c
fxcX+2cD12Alo5nhfrBphR1Y/kfnSUyKdnGSZ7o9IXV9Mh8Ngnr2rHsAuo6/xXBW
FbInaAOYABOlUVHq3Yw6cWb8ERwELYA0K+que/zO4uzyjuu7FakG/QK1t50xM67W
Rbdb0diEyOXaJSjHl4YU4pPGaLsun49zC9W3+rBNr/+gPjn7tBm03+ckIRWu0Ucb
rrWnlxSuOaBWflBkhyG83yDD85qcaESRYP3+26f7KZYDeGOg8TbL21YwF1ciO265
MnYjk+CShMng6YWaHjplXPuMb1T+ZmamTnTFz6nQSJl+ENhMsHbudZqUAoBhqGL+
x8oAsgRYe5Jxikf+LAANyhxLSMhPBizg6+cs7hIVjCaMKunrUrEsbhrbXnV8lAAL
DNH0ErSQV0NL3W4aBgZK+NCpoKlBasjBSODKBmtahpYzkMrHsOXrBN+1W1/5aV38
h8Rjtz7wNR7BqJ9i0NxTxg1IHI+sYnHuG4h4yzESasi4g7vb2DHcglhwPNp3HJNo
24WkC7gl4878hH9XAcwpLNkpG4FGplwgrn6A3EfrEkLW5Sdr4gg/+upMzQyGmdBw
E8wwu36MOb/4trm2lAv8rSX4Bl6j15EzqvlQxpkF6jkQ0QaeOBvTaJ/hv7L0RWHj
mPa5bcMGvihOeXThnPOjPtJHFdsZUScWFfUHcsDMkLSYR0hmXiGfcpbxm2xArBXG
w9khlscDHPqm7ogkMuyXJUWvAqzvuQLJN22FQRt0Acj9079clgICNEN+S/0NAGnQ
slZEP4H4L/Xj+GqnH4CMKzcCBQLDQPPc+uQYx6oxN5iX5jWLva6FplQMfUeS0Tdl
jfmKluhXx5R195uhDrdVuQU4oRrkl35c6kFLIvgjYQS+799HAwREJn2cBGNWsjym
F+qQJzBJMO5fRQIwoRXY3P4JPGgoTet5i60EXlG0U3HysL2BuCxCWBgYAkUna8Up
Nqkofa1PJd7rjsIzL6LUex1uRHzre3LK5kl9JPHH9k8TsR4OOwvO7md2HcKPcSdO
zTC79WDRIokOygmTtwSdedumK4MwHsJz+mo3WYWUOsi1AhF4GPVqi0TxyLgXRie8
iExfxWxL+I1j1mp1+4qlimx8bo+5AmEverFYHnF+H/T9EmsWXQZ615fTaNryUnIb
Dt9SILVybU0V3Pe9b3pUh7a2ZnRwjq/p1PyB4rSeiWulwQ6g8EuRWOsTvnElkr7g
HgYwdlJoXHXGnjEj5JYt+18C8FE44lAwh83707bZuDRj19C/BstDw0s9f7anyu+D
vvCFDZgKFOcUuGTsILoIpTd0On0FpBbGNADHd49d1PfAeTO4PC/YAxYDUf4nPGmm
vn4I+Fx8sC8SnS3TE6j1F/JsC2g5AFI1rczNQuwJowpcjFvh9bfWjSStEvxERVD/
4+vQ1eatdkLAcY2OMLPoTT/S1fY6bc3h4EeiDc8yO8FtKxzq4g4VfYiIuPptIR/Z
4la2cPyP6VPqDYdcY45eW6vMJmdqtASpt2rdF3JihOJlX0cRzw0tsGlb+n6rynGG
HBcYgoWO8AQp3SrD26qbujXRfc470xjKvl1Z4bm6mFeVtFNEU9976ho8+xPiiHWp
ksr7yE/uj/ped/qM6ETTqbTkPfuiDGvk7TdYUC3LbBYW29QPR/prv64gX6eL1Odi
svSL1m7+ujfX64BIZqaHrYMXtDah1+S3b9N3SddLdriz5ymIZRD6q3RSv/2OsjwD
+ndYQP3YJ2k/ilnBxq0JYY9cUXdEkjKc5ygR98f112+dwj6osmIadqZQNndhYkpt
Gyg+DzZdvFE8RbdRuk/Mk6TGXQgCa5HbgjYPjXz8nXVJJiRPBUMdheYjZKBvXFVN
CDf7akgWhG3c1XhYK6lJMgniO8y/0FA5CxVjAsZt79RFXOqD1Eu7WRqHTptBWpxB
UTL30g3MseBcmLbvq0imYaFd1lo3dahdKs87tFTFii/7hO+Lz/chMK04V5uAVwSx
0jAyBgnb/qs2vFUc6DjDlZBat6B1paQChiVjDz7/BIv59TDQZd4LEizSrYiiqBWh
974JBtnnj6VXspNXjby+H5LEN2eX9P8qC3WAw84asOXE//qAa4cVV2EaZXTYS9w9
KT/sYzOODRiXQlb1xH6kP2JkQIeIhyhpRaMbiBL30039C8pNpBRg2Dfx4l2UraXi
3bFmVkBG384+qYCKYbkM8l9FxGcbWh6RScvCmJJC24nYlXXpCc7qm/grm2a7JCbS
kcB72bzDnJ2f5L4m4cEgBA7m73lxIGz44jIz96hKyUz5DpLjvBE7bDApNKq2nJSQ
ppNX2lzXbY7SlWLzDMNYDk2XX971wDpTpAJRZ7e8ZgSISlRNL+Phz9PvfbPzeZwJ
ahe2FO2/KuPW9fFPjss6EuUUSkUjzrf7AdWIddW90t4fOTRvCd1uNopja+oJg138
Q7U6lDyV8dIaRvF8xPTagyJ3OnS8W6I3uuW26y7UHaWWFtdjXl+vDAUcTirLNoL+
BZjpMiMIQ/1eIkNXBxed3/OX0+kxJVxRvVtQIeI89r2/2FRWqkmR53NlsFP9my4f
KShMiVDAL6Z5/B5lLYp0MSEkDfHPJDS/vg1OD35uwgnmwNV6cfsjLS4oJfYYSFth
kJov5Dl62tcwWuQe6m6cWFLdsN4NdnF1lratM5q2ImjZfwOy1c3W06sSTNvRjxNH
sdL95EEg6qOPPGVShyelyub4jw/w/rlbmaA2EnDCBB/v6dOTQtYZPgGzQVawfJEH
3MnZQDNWi8MVcXnYILEaZYiMoSjJngSUpuDC5kRyNVpW2epIhdv6Gw1K+OcSDgpx
qgepDoJdCBwMnbQ8vjaplU+af+G1aE5wDCCxjzg14w2FVkKwtZvr+mWNND2/IBPe
Lz9JMTJc/36aYxlkP4grrsHIDQYGY/4zkkJQadv0k6LttYRJflulUz/7gLMRbVJG
xgenjti0SO+GUgK9RSr2U1mLic+HENmJ6GrZltvpFH688/+P37js2c0EwucsiUjN
n4rECLyTJsikTMsOtEOs0XVZHCxEXbwl8oChzEKktFhqd58wirW7tdWWUp7x0ZNi
szyxxDRr5Kvj9XAw5tND2qGJ/JiisD3qGwn8bJmmTkvK1ZRVX06LS3BPDN5aH3WC
EN6rgXkfI2bCpeXRy2vtun5qpN22w6QiLSecg25pLqtANiC6+s1sQwc5d87t/RRi
KkXpo5LTjrkgVEPMGQpLItENvyHFAEnN+B7h4rXUliGKX7p/DIYyk2Qf7qabKjqB
eb75jV1NQUI+9i3Ssm54+3swyM75wApFSKoLrK29l31nL43sS/0POrS7jWxNLlUk
clZhGfbaM4PaWE+ZwZYGge14u9ro7cz0A6bQl9+xTk7XVfSfbUzGmmBNzI5BPWRg
9ft3nXx7WaewcgjMIb2CJmL3bPSkmttM27FCGj6O2bpl23vivhjHUS+MLYzon5hY
REO8FCfWXaGJKYl99zB24ghmPVpbyyv0F4AvCSr/nt1DDDRUNCPdP6ZCcM65nrhT
nknZKwjkVj87dKOnDnKQOxPIGBdbyU6SR7JFcYxW1SzWEf9IbfwsHuXnkvLFunXY
GQhGJXSBu6bTi6nvQGZ0rP9SciVLe4//ZQ9vXTlYe9h6CsC50LrjiqMvnw+tAu+w
PtedLEY/CHXVF/3Cpq6x4sdhXU22/DyKmuoaQkQ3GYf86QKxjVWQ+p+eOcj+ZsWz
bQnFRpKTXjgDP2M5UPALZN6NVyNX7mRs3Q0NfdDedyiuBzbfdTD4NZmOk51xWkwt
76NMnapAFka5Waq1wON5UNk3oKAfilh7sD49YyKv5HSuCgvBS8yVjx+Y7oMEYCuX
jbHH20mUEJN1UzAnpeMEM63hnIX+68XcgDh53cE6qIfNf2vh9F8rZR6WqzeCGmEx
P/PDio09GiVk9mGciNwZiGur//hMHWWhr8dQLVoJwt2UeHfYLRehl/3KZwqBNWOm
Snr9loBB9UjgPg5pPxhekP8JDN3QBzlFoW7FMon2GWBg5UI7d8ZxPpYzJGDO9FoG
KK/s/cNfUP89nDLYKD/J4cJpWNvwOaGdCdPLtRi5UMWusqDiblx10l0jAglaZjDV
2Jg+TI6B0obFvK5I1rJA7N2iiEshJ3jO3sissAQbxlzBrVWarVlR2uMd07yN5ydg
8jNGTNuQRRgdbeh4ctWN6MXRyzFcg1SZSTA1JPN7keiaLiwl2pBVNmQ0B0fFqjQL
bK89z+R476lFvp6ekQOmShet33OOY7E5I/sKLw51R2s05YXPDcKRRAVOPf+THk1U
dR1uWg1jc6Y7bZcT/955Xvb96lhuqSaPa1AaU5jHONH6ygcZp8PUhGw8f0fh8Ns7
y366TYbW/MTpg1P5M783PQEJZy9DEKFgCiJjkBWKOB09t8/vE44ps99sXcjOq1vI
tLYjQiMwFayLU9JS3Exa9u2ZRX/X0IyHVjRcmH/TVxO6l3MSVxzFVOLeGFIoHEFm
Lbr3+OWIRkIZtotFoxK098JOqOH2CfYQLgVovzy7+KSr4k0//24efpr52QbXoReZ
58rEjoLt4kduYpOzKGYg/J78ptaBcd4PHf20+tI6KvZIC1WKAaIkO/Lzc+YnCWvv
SWMfmI85Ynp//pZbn6pNGDZaU206tlyBlTzSos7vVOV7xMhVzU5JxEUa6ue1kI1d
EaftuLYxtd9/7xy56U0Q18o10YREVQ7p/hBq/Xyp5RgzPyysY7gzOncZd2Kl+dBu
6RnETWFaIR+CICRY5uVEVczjhyTPrT8HTWfChyrZfeSEZUetazubXuYironSElmW
kjfyAnM4jKKnnSD7hMRNS7DQaS2nkYPAo2r+N4BLIZPAZmJVr4VMc/fQuBc6g4kp
t94JGV9VAcB+Guco66Q71Nxs7w47mN4RV3UU2fI/pxDD0Xg9mBhPIj0Hx7lVDpOg
x0tXaqm+6uHE7fAEqp+Bd6IxhKpi+lT875pLiUdYYxm6r8lV4jw7E/2NYb7+bwGp
Cme7XJ3+ShupWvLtcDLuGclRYSDFX3jWNtqEQjrU0BwU43mOF6xTa1ziziAoND/p
8jezb3uK+HV5sCDJ0Z9UX5tpI2WJhC2mmT9tux8o6UkoFmFF3O5btkgkqCytZpBg
0SGDixIbnsmG2dgYP3Y/prHWv9acyGnpwxbkvkaJq4J3L53vJjrfsUkzX/pKI83u
RdUVnqmAGNi4iE+40vECNfWmC0qh3rn1cC6rr8RMzHOH/re5p69Trh9StC6wTfwZ
7mAJb2Fa54e+h+hF62FBlTd+MSNVBnGpbxqj6Y4wpM2UpgIteqtdgNDCJMPZCLZj
8xsnXhksWQJL3BpMET89ttNcttIHK73BoUfgfoRfaT2/4qWBYo87pk9wpvGoLmDn
g1INVBZapHSPRDysvs2zmHete65jadl2EbqQdL4xsgp9FEaR7QNwulQuhK3hNxlu
D2YxLjEbbLPTXWQX5lEFgcPbtZghoS399bwHWlCgTluBX3jMRibkerHpH5VCLS2A
/lNWHKXJZJ46RpLz5eMplxtPt1Bg3C4BvmP9RRi7dL6Yl13nCqQsd11Hm90j6JYG
JUkFpdgwqLK8uhk8xAmj+Us31oOBQqzAC1C4sUGqz6zDaUU3hNy+S3mnGukaFSz6
hvWA1WhuD9/yNyvi/CelYDOU8d+2+ROWkhV4KnH6BgaY3+oKonZxSBApnI+YANiz
Uglr2CrfShi9B2pJNQP/+o1DiNGcNHohXq8jegXcTvEVZprJMsrWPfpqHwe1XNP3
Ex0fOr3qXDtBPMx0Nlb7WPI1dHJt7wMjtskHPi1b7CclfLtIs+KHaBzx8PNYLd9o
ErcwdYpUW5f8D5xjh9U1PPcrQ3fHu/GOGjMPTXBwYzx9tflbtSPSX9GNwYAhmRS0
5xl7VjXeI+1SjZEOauTdiaLQPDCeRkPt5vxE4GSrapRKvXLF/Boc6vWxcY8aXjfD
6SE9WuYArNGmZVfiN4J3SnR2QxtTQUU7GZPlutxFKMe98ODHTt3QJdg5HlZsluk1
xNoq6+Qga9bm1L7EdqtmSSoU2bLngs61kTjuy9tZtIA36I2R+UMOKU1Au8580dG2
G33TJNaXDnhKuLtEbdkSLUKzO/PsG2GZIZbLQTntq0/VUJDovzdtJ0Ym2AZr4abf
iEPsQuwk7CShLJcaRQ9wMqj4G8XDaaR8RaOurZrO2tNxhvaQ31oZpzl3GYhoEGQE
jBgO/u/iSWDdTnmyk+JFM151tWKZyGYk0mQcTqCeMth8bsAw2Jd6c89gbkENWM0h
21SRfGvETRdJf53RZhjBfwcQNn+SiRBDa5s9ZcwkdAoGiUtidYN3hbIrb3XxXeWE
TmdBAtbuK7iYnFX90Wev6LST9FijvhVQvz9zNeoCIfKotkIi9hE0mapweCcr8Q80
2wDseXl676Dtr1vMx6E8chnD1e2KWx+taATby7w7mE4jkige0sxZJQ+uyGkGcjmF
WDirWjvi4b9wzyOrPm7uKLdKx1BNABBPTho1lCk2Hp3PsHkG2JcEMYC0yzCw+2XM
b4HaoWb+im+G0HHQ6Keiy6nPjNzQ1+T13Bqizl1lS7orjHxWHBFE1+EsBKnsKXAM
3jmtWVMkuwNMO5RaQhxpCEonaj3CZGXAJNwVKeAIwKthDkUD/a0cZC9485btP5NQ
Q5eY+gWGN4tHqvpPCFXORqXZNgMAVzJc2bE8JWMG5P7EB7dZtxdE9zGA93mtoGuW
bJVG8VE2OXupNrmgL2AJFXvBcKtZQyGWNt5JH4zG/71sOfUD3UobIuUiH2I4o3qi
NsO0ti85CwzDhelHyFF49lVneSLUfS/1x9NegI6q3w+Qf3z8qTrTFzP9TAY70b2f
owx35utf4dbiNLwxx8kwrcl44zR6Gy3qAuNzoLPXc4z3Jks47QL8anoIlc7kf34t
80q7zXpcHBQngjt9v3YQ3eoPEIbykF802KKsGpMULWXXRHJsil7ZrRlQUeHUg8Wt
fFEui9ST5i/ki1lFE7V3FNMPCrwfnOjJnylqfGWyT6X/hfKcpvFjFehblIW9e39e
r90j4T9BsiXjM8L02F3jA474EVEbnzaguzjcbpfaJ72YOXeQSwXoxY31djuoZGeo
2Er9G1tj9uWRxGOlPYjarV30yED9sIFI1lj+phsub0qy81z+g0cMgvQzysBsQPJl
536ZUTk+A73dZDbvBiXcZbdPB21CxXlrIJYGtTvfWL8TrSRvz1NXU1BcIeViQwS0
4CBHVJG7TRiXp1P0DhZ+hsH9hN3iAJ6BIjUgVT+ZKz2Y7/sOCfz2+gitqx6UnWO8
oviHRu103BpGC+jsix8zPtdYTryjGzVYZwU/7eZi4NoHLduxZ/QyBG6h2xlM+MzU
T3hnib7ObMg3kdQSMeJpT3b62AmIEee19P9/72xo0LQIKDsrH7mTp6qccHCGni8n
Pxl52wU9LrPtKeNIy/qq4/L0S12uXi+l5wEi6chSYJlpUyzmC2DqDeJ9Fnc9kF/R
OD+BB2HW6gkzUY95GqnxD0SdMjZx1I6oFznXpG6sWmuMotcZuwIV+xP4OnHRKRAb
YamNuHfpz9Kiq5OFPtnw1BWkTwOMWMeh1CcDjXGfwOV7KPcVgQiS8jh61kNlzwci
7D/amLcovlCC3jrP6DbtPmc+sUjAthpxMZZibsDY+civt3yt7o1x0EYlxt6ntyKu
P42FF0nzuxHex+zlZaIeBAKHz/Y0uLE1mklgz58F5rgfuim/mtq7yLkN0R5ZzuFF
/rrRTgIbDiK+h1KjfUsheOg1DETCiDoTEzEqW2BE3LlsHMqwzu7ks60kNpeTttC8
2pZ7S6pFK+W4YtNZm0XKx5we9NLqGsN2TOoY+wjiKpfTu1buP636o+jYh+jIkC0Q
lat7MJzhF9HhtbTpst68HUtUr0cvEmv5h+cRn3VBt8JIadrr+ws5/TZffGL4pQbb
Ot8EIbJz7+RL5Wawiu5A2MgVCw2n+R7DdSpPB2uPOeOMeFWQ2cj1hQGzVZopSMM4
K6FqCMVVC3Kp2/jTmrepE5q4Gj1lZPedekz7whIN8p0Xg7hmdz0MkC7YcM6UEjAQ
N9lGnQ+1qQHcqax8igNGxqYTfiKYdeDESuP/swWkY2MC6RHFywS1mgox/+cTVkjN
/bYDw0kc9tcsfXDzc0E7Xpd9ZJN7fy6jBxbkrkuyHdKCP0s6fmNFT+EW0u+avK3J
w7a1MEe+LsrYpQXg/jKb0wA0OKx+fjNPYqAvuTFHnwKaeHnVNq7uPbLos+ilx8aS
g3KDdiTKo2DJTrvAdoNMyi3ugX8ZwnQ29mABx7gJ4kwBxxUnUGlyAEVTBWILl+7z
3rXFQ7f34CmWSp8hOMUsSsxmeIb4Ckcw5WGdNpjdJoz20kTZUrsUNHqOG7zRQXCQ
Mc2fWITcKxq53LCiU+EWv9bGP6Ri3n0E/yjbU1GqJRO01TMmvdipRVIFDy0kHjFr
sgYR7mirho3zkzNd42aE7WJnOvqHvlpQTjzYKkXCf2ri8LdeCzwqARBCcdCaqQMz
lRrjeCmOkS8ShXteyw+CLKAVQgj4CGNpVzohH8TozcBowXqR9W7cSOVnCy+Mx0Zr
ERH6Rxa+w/FrG52eYbSvEE24awCQjSb8PsLvFGYSnAMbl8TNaGojCcFx5ddmC/YQ
+xU2TgbmH+8YucAD3GBNIpP8YlgynjN47v9IXgwg5geq/bbx0nzfOdeLUlh+3XFo
oTX9g0iKMQw/Yv7lmtGzhY6Supi3/kfYXry+XpZGd+uylFU424kYh2jnr0QmwYRc
JSpbVaP3EchFGQVXybc7ND4NfpeNlFPeNgUeijyWeJ8a3vIaSDM6Y5ugULjCtJeQ
EFqFH4jxqy/MiWxTYrFHbO2YBmZKHLlxYP+M1MPLYPcsPPmttGqqxvKaAXaYbJg/
doi/W+N25rfBqYpD+Ve1RdoslxLrh/sZPrmPqIGgS1jryvme2L7QEe3NRw+rHUXV
Woevn2T2hke3jIyePgXuO43r7xGUVTP2BY/7xlrK8jUlAUAxgl3pOLa+eyGHj0Hg
ilVAbFENHphJwo3dcf3GczRWvmADc5juZtRSB1rr2el/tD+gSrOLbyHYbSg4gKSd
2gLbLcU7akFolMdtvAFdO6/e2Ai46SR268vQYePYPY6zx3rm2+Y5CCUVuFsQMmjA
IxPwGy25BspovqLHsromfV3mf72uOxX4kAZ8559upM3eVeVl7TiNaaFbO6EO2lY7
uXsZO+0mba5wTfCVyq6wGsCA7Qh1GoPf3nvEVe5W7Cs/6LxunSfdi0/nV19KxxBi
3UhUy9nIvdcrHKYTaTZT4A==
`protect END_PROTECTED
