`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
onlKQUu+7DSnwgpHLJ8Ltj38lE/nHWSh9Ftt37Ubv23oXTVsPsxCv+C8cu2JzDkc
uIeJlLyFTbf5nfxZ0LIYJddvREzPN9EpPG8qMDY2Q1jFXpSOeAt6xI1M3pQ6Yx8g
DrLDwj6yDy3PrA6SnXFyLpD1lOAYmO6eBcRzMC/JzLahIvUHtznTO8pLzafN9Gaj
gJKHAkRn+yHxObF1D/sV+AypD/OLW/ruTq7rG0mJvXYW2nFG6P3Vuogze7Sj2mRL
dis2F4mEUW9H7S6NlOiJp9+/OLmlqIgSnkjWMDcNGenhap0cL+Fc6/wf3tS3rF6d
Js3s7WjN6U9As2y3X0DTJKNkNPwOOU3Sdvl4MSW/yBr40kL19NJgHHpkLJ5EJmzI
mTYCMGf0cwl4x7KaCHXP7tDErgFi0GJrnf+Wv9JOp5B/zhD7cOpcdsqHtVA1MgxH
NJm9ojF1zOa9fmuCi9zckIeKKZtc9aSECPCd7EyyGqiwITbgvteUfzBoQIU65U5W
smn3VCBbLwrhiQ6Rf8kwTfI99VWf+Qg2oggoY23qjpnnvMzyfyrX+XHJeyeYYZVM
a7pYSZI4pbNcinVR+RR16dIQi42q9f7dn+07ni8MIRUHQwk6FLoqpTwXE6xs6c3J
Yj760yb2OnQBfpFXRxrjiZPJIqRG4ga7n+o1Rqm+Z8M6xlKu7icNUazm6HBwF5ca
KVA8CRrpE/0f5ur5A8kY9f8iZmw2OwklYZoHhEtbVWWecOogwyCy5y0zenAaylht
QiS34H6bWAI6xPD9E1+fbx+BJk0HS50aLkPs1wj2QLNtLsT9EQwimneXWAqVZut7
bmu6cd0nmtMW56yI4xsHKGyNQj2F9S5ZLduzL12AsjeyrlCAhIJX57HMziYPuzJM
1ISHwgcXZsUCijFLLVpb3/16QUHfMqGt4uWHxF4Q26wtM5pcKH+0r1pybtIotnmy
sKtNJ5qOTeRsYB3741xWC2FDMeBaNzW2mD+5rxGCpx2CyXRKMi3J+BrK0Mu5iwDJ
7s5JOUxYGqGazXcw5g00GJhBaXGhJOAeM+bglkEaELVjR1lC7xipKsFuYKIF8J8U
hZbnMOAIU7bea71SzPFgQDfllCxR/gldedRhAjSojIC9SQiOLBj0srC4FBSoqNfO
i4DC7M+IU3j+mm8ufklCCTjdg/ISl3/vwZKZvbuUfkqMFDW3wJ/GBvpLy3teLtSY
NPi2HUerwzHDj344GmFjRMz/SfoEXtzkx1rMDutZsWskqkStunri2jhaVFDuCN/3
WDdll0YOyf4aGqsf1B879o4VLZZHuBgP8d6fIjE6/RnjctnfujlExt3Zdl3JfaRP
LO+hg+xm9Jqvg3HKGqREl72AYiZ/3N1szj77uaYFA6s=
`protect END_PROTECTED
