`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pCCirugy3fQ2zo8dsseHQgoU7TwedMpGJCg1w7hCs+bbk5ca1Eqi+iWYQuaryBYG
XaD116HIE2H/OHpPH3qmDGR3s80vrqBWsRJ7O1l3s7X2H0UkyVc9RDbtzQSfd2jG
8QnPBSBcO1d1KjiwSNXyZSJSkeF11QJu6BJkDVKcldohMr/urUwsNhc0G7vH8Z7h
YnSgcOmILSdRhUroUgTkuF2WYDhk3BE5wQb8eNssyEqUPuchDLvZX/s2n/5t09Bc
eWTNxcdJujxrPPPjs9zNiG7lZ9lqR730wiVcvR6JO2qGMxgFkBSy5FQVE2m06irx
JuEO++FuIu2PolnII1+fC21BhM/kiMMNf2O0lzIuJTSkK4vyhl50jVZOiv1u1QSz
LMsxykigdAw4rn7rOL4KlgbogltnKqQGpRyMTDxSc6xVJ+xgjLV6QkK1kL1ZXHOy
x1Uy+GSbV/UH9R455nc+BufzknoTYXhknLpDWpgObaUOZjFdoHq2DPNDvreMZ9RN
vRyr4/80YpwdMI6TQhN2iH9MDhhEYriugptsxzBHSDFTHTzXcVnNPCpzUH03kyR1
HFzKN9+9ye/UdmHMvTDSvwRLla/RSIxrdqxo6qJZXj1DCVnTqmKQUQ95JNH1BFJu
7BO/tBYvY0qJHBvO/vPvsywm+zyNyErmqw5uZYRDVaYReQZmUtNHCJfwqZU3h7Fp
`protect END_PROTECTED
