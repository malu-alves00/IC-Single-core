`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pua0v2pU3zMOp4kypc+pnsO2mFTS1aNdMHRiBuFOe9Bxu8cWAnXHCuS8YQMq3Bpp
DntHijOdgDea7EQesQ5Jo7L4HfImQD62I/6JtXinjTdq7C2ey1pVqUZVuvzrczJ9
FB4FMC8n4s9YIq5yFw5yHZRMFFMPSiwK5R7R22BmCCbPf/qcakOrj+ycduaz6q24
zwtM84EhqU4B/Yj+YG8xJDgk7ooJWYr+PGqclxuwJKYRq3n7q3rFy6tERwJTsB9N
WygMIjbtg/DHYkV2dTPCb7TkzydWJF7hVGAXjDiLuc2UxNQxEtBS8T8euRzPCisu
BtPURpr9t3Xgffhg3lhhOMcnpnGTI/4d/T8jkoJWMiOrcfA3x9+/elP6PXO4EBvK
voCzfrCM0NIF9TTDtzJooQ0ue1kJ8zW5w+vW/j4IlGTrfasxMjJml6ROKRWnE428
nfwT55Gl90Fu6olMAa4ISw==
`protect END_PROTECTED
