`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
K7B9RBKXGsuCzR4DEHxzpCzAa6DNg6OoL6hLrR+UKqqsymGbrT8f3JfPg6j1Bhve
S2uZmaj5EG88I4Y/KOt9tud1MG+24/KBcgW1b6AtxHsrJv/h0eRY7fe6nb+OVH54
qbFv5ityO7ohadE7WGmjdv46w9/L9oNb+ALnQBiSiMu9kMZslxj+DL5TcuLTXRWG
g3xUzX68MkyFgqlf56O0Ua9hafySNR/Yj70jHiA+kGjxC+gWKUm4VE9S3yfDs9qx
IFUXd1Xdwttn2tnHn1U3DRbSgAxLKx1GlH3oOysGeCoqF2L8euBoS7oIjLkfzJLd
T5sXr41STihMgfyp5c6z54sDJyDlQQdjq9c57QzJ209QMMAKAx9h1m0cDhdmgttu
8UMooohW4RUODr/asZ1Tb+aj1DWHYIg+dnrYcmT3MyLO9igoW+Wo2JgmqiNHNVBe
PR2bOQET3TaTMJEqALV8HGHdJSqdPdcM8jO+wG0uGxabJx0kpdRG1nDAjWhd6rZ4
M+ehI5rLfmuCtUJaX7wjAbw95MuUbsZ0Bz0vBa+VTpv8SFzAxD3BEpoiKfbYlWo1
rQzBn+nWQIqpZilJTFK5cSMjPAwRBEr4rQC2/LBpSm+ny86bUzhH49N32xP5QMET
Wci2rdsDMd8P5XkqaiEZMdYgeT1HRbEmUTfZccJAYR8s4BzhVcSuXRNYjmt7lnTB
D6ILwFQCTTAeNcRWRtbseM8o8nUC7PRtq5/O3jKE8E3TwP6OgpCiLOdP1TtAMlhQ
sbNxC9M9Y8Q8b6Esqzc6fZZebgWImcEgA9jxmHeLhoXk6tCVSl57Tq49tSJ8BvAg
bNJLv3tRjFUvTFK6AtD3H4NAJ/Hxq3EoAs7EYzcnM24SdM2v6B4A6HChggtYQLVf
lv9g+xx7MqL8x2UTjLUeH2ohJquK8OnV94BzSpiQ25gMMHP0v22egQMqJdDxrRSo
/OXAXs5OO+/7KCchiwtQn+92+cCB6PiNiVLP9PuhPth+4j+NTrbfd87bIA7LeQww
CpagK+C8CGShbev47A74WSXv0gpk1QqF/yXJ4qkS6y67FkqzrV59y7KcngyLhBKZ
8+9L9ZehXkKqGny8NzThJ8YV0ygfvyUp8aOQuH7KUALIjEBOKQTnuMRsMDjPdlVO
d6CXWQd61REjjaSsOf0hpW9DJXCYBr2SwZWLjsMnIKAEwTQRY+YClMiyYL+txMGs
teiaNvXdEzh57pef/bsUrtM2aEzbjQ55y5e0eSkx8omWZrUc3ticf2F74VmIIG5n
XPQzHimF1ahOAfglWSxeNPaSF8MSSTXqq2ilBCtQBdP3v1ONhIBgJPU6NBkW4pT+
TBw79tRwj94gOgUbLbZSqt0rn1n8LBHSq6fNI508k2F0C7N38OaRq8ozbmqsPfr+
U/bmiaxI42wzDoQ/37BIt9Yo+fSK+6ubojUydDpAGRE221bcK9R54qioiAgi/6Ye
YMyUlhQIZnXxmSg7HLjtVNdELT8usBJMSYkDvxdtchxxEVEUmw2284gBRnJv23hF
vdvnxlD6VTouKTlCh+OGZWr1Yu7ZWUhQOjvRNCC41sqMmlZfTMhtwx34dD8yUMjH
Y/RLhERT5AtBn56wWg158kGVcHHyB2HuUW0lAmQbM7qxZojCR5YryoNCcE1gYJ7u
QJD9ikFTUGRZX02S1qj9V0NzGrK71T6v8XeTdbtRet/GK/0StiiuXmyNPt5eNZ2I
+X0kcWaSuhcr/hS4DJfIVkxPAKYdGrOoyk0DpsZCRvEcaPIgZumym7JlN3A+MhxI
JkzSQ///IqY3Hzw30h4PVog63W+11bXkqsM/CF2ksvg1ruQraS5NiUNshElBmJCE
cvb/7GRnKftfJP83iKciE6LPzppSZbwkRzXlPOfR/snjtR8A0F7RPl1NxKM0akIL
aBB7QnCT64jaqj626REjoaM/K2hUBciIXaNB3U/zLb3yj/mBgNAtS4T4v8uoIrc3
jWt3gw2nVOI5g9/dyL6tSoQo4I9nn2dfwn01wlO0jMZ5XcIRtGenUBO8bgr7zoPc
MafRrgJMRi2UmYbzpSBtNl6Uq3h2PE/mnGHqvj3zMylHm63GyTRXbCm530QxAaYn
l8hkR6zybe9YUD+7VZjkuBzTbII9tpCz+dhaEDkICbrhIjnPgBKJPQkbcKMCV2nJ
hVyk416uCksehWlaIYvmx1ZiXP0LaSZdOhycU/0CXzs80VGdSvuP5MgPbwnboku6
IY63g0JkhScu4O7Owqt6dj9ZL+OGixf4/WQAkm03qtGHWAiYkFKxBBoyt3/RwSuo
WKM5kLCWLUZrAeeUmw4hJtFF2WM5dHeTRQ0RoHiww5nB/cSdi5lkyh5gu0/r4ZJv
6KcThW2tEqjYFyIikvvSL1Tyj00hgRfdHm4nG49hEWxbrMROhJLbygHoBtJ6A3g7
rbLRyzct9IG5WKyiwASXK8Kd4Ac6lBlXgSBf1zZdqW+PiHiEA8SC/reghkT8Rar+
GbUC3Ee8hD4VWQcCu9ySVVa5x110cgZrB5ymjGxrA+HTNwRQh5y5KhRNaG7b2Ioa
ibOKzsmFj2sZ2k+9S4HvqyUihjabM+FdrPvccNLdAAnXr9lIC/9iwVQKd9XMnyE2
NllwY64cCv2LPyEAy/4UeVE5dmhsa/aSLtxaRuukJWQHsAgh75oxUvoDM4kuN2ig
7r7j6DZPDEjgHqX42DCtm+hMK0fj13h98V1Pq/Zp4UOR9/jwBnDcRNLqkSC0miIS
GTPPZ3AIFRGp42H02PEMUWviN6RHfwA9wTRl8ZPmXeZRa0mtRInaLfg2n87yFB0d
glXsSc4TLVH/6udYstRI9xoFvqGYK1FIW1xNOoeFTPjhU5EMejs+2kTS4JWRr+ST
Cl9wxpJJ19g4GA8kEhX7txFXT4QNacUHI6mSrMEs6nxRN7C5JPetMxwfgRJVoI9a
LwsHT96V90q+t3kbTtiFx99IRsXputEf6vZymE46QPx7WJcOOyi1ZyeiTPoAmFxG
cVlZKXD9ZWOPTCnXoFhI9vVqEDH0/S3YJ0GeDMFfhn8TSpP/ZRbn+SzDvZfS6+7z
KUOHu0Yk/gUqcy5KUGIETWJLds3mkVhgoygccUBce5r7SdldZT4KvDUORhYIlaf2
Uq/bQS/LXPjXQHqoRLhqfVdF9ScNY+65VxYsPksPqTNybIanHEB5Y+2mZPWtVjiv
LTlQ4rIbr9TtF7lo4ecngzETKe89ByTGmrq8bEkTM8Z22kKDkT708dssXiAu73XO
ri4Glton4O2Ql6dGPIXRncNeKDbqbHAdEwI1ZyTGtJZ7KW92RrD0ePydOrxBdlt2
TOT0otnK8q3Jc7VX4qWJxethFTwNpOcZZd9/aaa8Ra5XQbp1XWvG+otrlrHSwr8u
8g9DrSrmrTiFbMhMj9mTs94tBY0Dl0ciPQvG0WKbSBZM1HCyW0HsTbgm8SU+QuzZ
r3g2al+ZkkwinV7K49qjTc8XSkIqGwacfpmYsem+v01UiL7u5TdBLDrT67kDRGGL
DugEQCtY7e+zKQBrKQ0sjVlCDbIkfDVWM05/H6Ig5Ln8in+sYToVLNoW91kcw7CV
XU6vDEHRXZOJubqFv91KytqH7z7RvxOunL3pQyEV7vAWZdJ0mg/d75NBk3Y73mlb
04LuwB/1SjNUmJB+Jr0XpaTEg0dpKqdIz5RJOIFimr4VqYiyk26ZNGjf3GbC/IR7
Bbpe8/h1DaJvJDXeQEFl0OH8XUlPp0CXVTIKCyW6qX70FaUCr/kifw1M0OiAzU+S
tXM1TEuIJYJV+iCFdyjS78G7uiYZ7eF303SOYAW8mQa8OzYKyVM3aTm9WSa4m7RC
6KpIakwBS5UNVY5qFmvm6Wh61OrfXYwXtdWyIi1dj5jiDo/QEqGq0UXFtho0hoSz
WZ9+P8f6kn4ZmQGcWt/75cQW3fetNsIv4fhoH6WSew/CPROyl/iKyWI5UfJKCuCW
3dWuwleISUMBaqrFwi7Hz1+GZBFfprBKHYb7YtMmnZ9QB8vgqZXPmitU71DSpU2U
nRyHQTSvFPO/kNAMlGg9CVxD/mgLZ2DHZf27XrxWxdhegGJ35wWgdbFMkHc4BQ0Z
1qpe652K1s/fJzdZ0T5HEZare0hP7YRZMD6sa4OSukh4FltZEvuGcW8zShP9XwLm
4RY08JO+SsMM1u2pF6PrTqoxNBLneB7/74JbLJfwk3a7oH/Ikd5WqweK7UNyQRgf
i8TCwcoumV58zpSh83XJ6uNwYlP+DmKJkvA0eS+3q9qOQCx1UHWBTaoboAYmuehY
ipoT/upo5W3/wHKdpIcllLW4Omfszwwb/hqobRafsdbLjI845KMriaDRhyxev2Q3
haGJXmwlz4yL4kr2d0lLg3yV+J2WWXSIQcGK6DfVfqQsObeogaiCp0MPn5MPttRk
+NXqm5ODaB2yZwPq6gpCDSINArXs6Kl/Goy4jvUbr3At6vsqLm7NGa1V5jR02VHD
fpQZ0gHx9qrBZ3F8LhrPDdXUbsnLmbeAu3KxN5kFasv91TAKn2InhCCDxoWtHwJ+
O/2s4D7QWwfoi4oYy7M1kgUbcDqVFnU8064cZxR2a3/UeHS7KYlSgBn6k6snbAom
ouZnbdNn6U7HuRTc7UMGQZYd0jItWPc+OV9wsPdjrQ8KgwPw8UueWfBHL66Yx2e1
9Vchxg/YbmuoeoHkfVO/J1bauFIR2VGDUT1lKRw6Pj3bm+y6yCWfq4fD4bBP3ITA
CurbIG9dbtMG8IUk0zdMeUWtE0Jr3oqPj/WSJDPzUiuCBG154x6pTEocVCMizTDC
3zsBa5h/JpBU/MOXFLIQCmZ+wNH8WTulWvKsyn8WruswnI1iLa5a+XLboJBNHLZF
r9BausjeOXP7atJPW/OS8IxlS7/kL7jqh72y3Q88yeXb0DWysUuk5VlYJ18QscOZ
NQewM7AW7D38e7DOqFALKqnLITG08mYU7k9f5rkVJ0nVwZr1dqvA3RodkLmx6qKw
pIRbTY/tWu/X3f7xWgE/Tu27tNESuQJLoAlxgACR5NT4zzJYi85wYBm7Fbg0Ib9p
zcJauEkeLH8iyD5r+KnxgnmXfRvWk+SgFuem9/2a9a0jH9CfwYbu27Q2QllLuRf+
AKggfVY8QCPobmlLQjDiF9YY89AN5wOTRXyiNMXryTZlQCrIjfPUr2MjBEc6VMjj
3vgowL+YjYzOwsgwTqOd3+tnx/Au3vadhlMoIdPZgpzgFmeDO2vhEy89BswflNTz
gDKFjPM2qdhbzFK2knM1Y1jswGgvEwlrVP78FQWS/L1iJaEQQThPyuYgsxePfjRc
pJY2sq5k6ZFzZ6d1ziL2CKkhV8EtX1Wuq0je7eYN92opczDW2G5mXlsHX0cJt3pg
sK4V4zuiyV5G6pTrw9Yg2i3zu0q2gANF8XXdrNITyCVM/vSSBX08JZFvG9pXMFP7
yIZr4zKIEmbAFPn4I7z9bEp6uhOGabIcO7Hetv3THa8epy0ZSW/t7ytYO97TWrH1
6amMmP4FdLyhCkwO065oHrHGSvEbXFWtp3+KBeuyb3v2WFvKXxwQ4Opx1Cqoo57H
z2qacdv4bhAXtnvBzp4npmv3MQ9QVsJ2/MxiE/Lw8GWb/AS+0mV7rpNw7mpnQNBb
ax6wHx63s0qXlqX87u7usDeXFtWPSFQ6DavLiJiJ6V8GDRDqqH/6FrxmAFW53byP
1dyTl57mwP0wopS5jw+7XFFCIeCLPlCBEsUSPbg2kPP6bZrPJ9vjyXtxSKhe/R2B
C1Z6/lf2kKkrXObIH3xG6XH4uNntYUkvbpJgTUfkuo525M962qYaO2A74DAw0pQY
/o1G1BpWHD/LvBeu+ZdezZOIw6nn2RTyyzSI/zdY9vCp6JytvMJzbL5/LNhI5tKL
oH7WMH248T1vw7vJxx284onyDGqajTS50f84JKrTp3fGDmF/9qobTFcpHYufbS9K
OCyxqiOFBR6HBFh8Q38dBbM88OLF+VCQ4gN2gUtay3JNXL8bxMIbPdMna957jfvR
B6PebQN6fXRMxGWcqtEsR7wgUPz7yd65eUiLscSTLNUnc0CTgWsNyCW460xG+ZM8
xLEtDqD9ouL7J8iZWZes1GNwtu5sRh6MoC6upS1HLT7NkC4dW7iJIuMnGJqI/wia
WUNcNs7sqVf8T3GNdgvepDRExkgvKdgt+jCM12yBa95xWjoawDyqY0bmpVPbmU2w
IHokFabl/TZ0fIYzE9sGWy15D93uD7GsoQg7UOIP0JWZKTbXJ/YV5YwzphLX/K7Y
2SMiM8z2dWfmFinlYclfH+W2mO7nbck2nMs8xY8ofgsjPj1CR1nnESSwmB3uVfnQ
Qv0o43q8ZpLg93DjXeHC0QdnNIfdM90pKGlhtlHdg5d5FgKDZQzNc+aX+x8ttQPw
km8NRPI/TDBywZzGGvzBT6Wp+h4yXM2C5HsJNkIDCLJXxFJYj/CldskwTgf6BQQG
sIQ0w/NbMAtL36okJU5cHdMrTQwq9qCUBQPPJnm8vHlo76R+9vB/Ogu0e3ZxjnhD
PflTtwE1yqWGQq2YoM/o8rKJLn6+hEZHNbm5qiAwBB5AP+j3aFbFKmd8ugLoHOtm
3y4joHLlMjuB6+5R1kLfUWsHRdZp57kVUooFPignPxyNSWRuIDJnn7vlR9BsSie+
bFIGDqalS6nkkQexN2Mmz3SOsLK9stRnF7Rp+zuaXgV6Nne8TPiNwJvPhKpmO8zz
TwZ1EuAiAbjflLdbzo2HYrHJV90/tlU19TzG2j61elGZOEa4a0RXjTmODm6wG2Te
Bs0JtHFpAV0Hq1mcKtA5ug75O1y/v2ivfDK1kXjdpRdzaf/E9hjREww2sAgAEQR9
51wCrMS+r398BaCTVdObsLUllLkIWCF+q0Uxb8baeNw+5q6BWWutj1Myx67m7+lM
Q1HAC9OTgyBPtF5Viepvb3XqXMzABGBcze1wa68uHCmpF3WHUgMra9TRtSEv5IrV
SVX/Ta5mCuKhzsaLPxYw4r+OtqhqCEV9mvKiI3Mm+gAYi8pMpkxrW4maefcu1rEu
RztA1Jg/XMCrxv4kfOhCEdwXnulaRJt1I0PVKXX5wwCPhARrIM4H5ZGWNqcCsaPD
mgHjvCuJ9EpSSa2Gltgb2vAWeGHCwc72gc09zoI3FV2fc6QDskollBdXhXRaEfBe
Q4J8ySfbCqGN1kpcOe44g8CgSrTRwdVt2SVuhiqx1aXfMPnI9pHmWQoW5f3eDlFu
V1GvVVnf7vOnNS55tyUUOZtdhK36Cemo0ZJmNpHo80XrfIXa9pryTapcAnpc4RTg
qeR1mcEmfmBVeFpl9grGoEYbKBGMUf1UUgE1617Tj+1hJ5Zq5bU1R4nJhlb+qtlZ
1D/q+owxl3skUBnzCfhsjgTpzk0AAbVej1H7PgDsA0bG3icIAzKStgsSkNoCU4sS
XPt8LW0810/ddM0WFH8WWqXe1YuGFABZGnL2Sf/JCpVkfaQndbPXJKxVCOAVwR6K
3paorU2eUOgVFrwsrScHUsqfv0agLLV4AFr07a+cEyhU21qazsgx5m3wDl+n17ge
8JdkxNz4jN2BL7mB8ycgj4fjKHlQHdu3BHxsOHfdoDgKDPj92b0hw47Ajt4P+zY8
1+X3C8ECbTZw6znPcaDQ/Bia1pJFzaf6oxPintjAjCfVWirxOW2gn8MOuPRPFjT5
KkYzWU5CRVk94HeScR81x/LJ9uBXzf1PlVTCgcTy1e50yxTsyGUZGMqCqoC8YQ6h
aLesp01mU/DkYpmFIq9N70WAXFllzwnSgzBz7lC8/9we4epo4CAOKkmt7Y+tZbbd
nSV1EBF2W4pOzIVr8cCcLGmIpGiJvQSHJO/p7NH0xxnDMS+1MszzUSCL26AEeVzb
I8itVi1bFrKh74EMGjEOlwwZ2CtcP6sInzVwyVh6dfFWwAGWe8QJjV6270xTY+7O
dcCvXjUiE1zzpHJpPHoQXnPEcqmhsAegbt8Y8cIkRO72HjSnEqql1B2H9XzMcD3s
CtZu6/sMcpG79UbPP0pgw1KXeL7GMTaPfc/Q+qSaX1CA89lynERZiDEcGu/h7mBf
9G9kBQt2rOZlNTL6t7BYJmz6l2TUr7kzLAl5R5AEvoZtem5nggMWUarxaWI1PJKp
DHlwmb00w67Jf9lscnIFSUNRu7NplU69mgzWDlOvQro5wwD/V1mWXAH6pNrVvOTP
BLtv2b8ezxXZJi3T0H7I4mZMb/a6eDf6Gxk1fmpzujiIgQaS1hP10OW76ppjfgZm
f/TI4q4xFJtbxswcTb3qo9yAJy/LqA6FoPS7I5ngV4XvPja5ENQWBPvwpfpeiYzO
MPw44P1q6PkFJkpLH7sH0bK2rmRl90YGm+Ln32ULLugN5TVrIzHGG4pSEmdaR8RL
A3lbLKuFPzIxWI4LYCgU9/8Q69IhRyWQyPYw+bRuP/2epbFaslUyGgOpO3VDfaNT
a7rqoVsFkhP51vBNAvSmaeSoMuskNv0QwwFo77bRRjjsXbfSDGk+pQErdEjw4lUl
KfenwoWqDHw6weczRKlppCykLScOkIaBopbDAgT943C1Er0bhBQzS61py5Uc5XFf
/lAtYpFNgSM1ILyjs8MbA8SCiO++w9wH/dC5MNa6MNeFP9oAVXv8uCuIIPFUOJjO
NQN6bgXZivCbrj94DIgqQu1fN2OLiP+K9/iAIWfvEw+D8SaWL3s+8/LwQw1sdBbI
zOrML9suiklo3xbmNr4ZioDyKcaxd0i2q3zCGfNOGe6bUpcwxHsSwjNOk4l9yNDD
8e2VHNFmTw0mIO62lBM9oxF5DcVlNhfUVdytxFPJ4jOHkR1Zd8oyhYmXRy4PgSGF
WDT2FJMd/sdum56qsER9SAwMszfEFzsEzCRategRyLGCtMJEC+fDaRrVRDknIMDx
GN2O7CQDF6ta8TtoyJ0frclxHGsfBgI48cJgzjRZuUzx1pN4bY2DfhLSKVTOZsmi
ApFyfIqZsAMZV7PX9tdU+v2Nyp6JEC8LsSogNsU3Wf5HU8jdNFkJwT1JZ0KMt9ns
rkaMJb/Iwkqpu7UMsNhxQ3Lmt7cAVlQzo6hPTRt/uAAgRQWX37ID3zjKbx2Wxo2e
SgKN0nRySyi5KGK+3nTya1wnFR48Rn3WysBRYApOk4uUS1EOLcGsCVA6o/twbzqh
gu4pfxALlBt34JzBF1MXjsgH/N+u0y1eklOqMVpAhbr59wIS0b/F9VPTb2YpQWIa
2Gaztyi1cVXEo89V4sZWwoufKVf1/0fMJsONlDJa0yfLPUhFlfv2bIoVsDJJa5BM
lwFr4gEjFM3VHFCZ7G33XhH9zJbnetcZd1LJ7Xhza3bj46THIwnj8sNm6JDOJ6kU
ys75M3BJDdxe1J9A7uhHgfpheg6Pk+COmlNDS4MZDzQ5VV9mzV+uy7AoSjebgENt
2wTzu0205KHgvi5NWQtmHyvIDAwTtowMZ7lRJPaZf0ENNe53GIH2CdYxv2egpvGc
YbVE46AT/64oPw055Y/6Wg==
`protect END_PROTECTED
