`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
m+/RTxGSVaiFDwQ7Ll22cBnMsmi2sIRN/fCXmHbN56oPv4KugqQM1PMSlt02wA3m
yE5NMRYOAuY5wEArkFBc7XUtB531K9AdKxFJ4MYfi9Jiq/8Mb0W+Y3S/Cbk95wCB
RN33EdHVdczZJPlF3fPEn9MYvCPBlQzfqyZz4RnsVUayIKwxxz8wnthA5URuHc/B
n+VpMsoQq+igubbOWd0z6udasw75prMtmx0BQQeE5wIW1xvlbxfKEAQ+REscvH7m
1Fd8ou29KXA7mpXGkFDUkuYhY6++jg/kEkjl7KQkaGEtu9JyEb85iwXigecNQh4L
0iIzrhADivpCJg3wDQR3uZYiAuTl5x/IpG31Y14RUsRpdXmxpwBWdphtGvlLeILV
3U7z5PuKd3O563ijjnrrffmtbeLm04xdB48Ecoxbvvy6nELd1JuAULyLhpReJeaL
gLDmqFvyiw7uRuDrm6Q2ElimVwyfEBJFxuZA9skCuYj007lz31ppivZftsWAOQZc
BP44pdf4OcZImI+KpvhDxIwNnAKaBlqresCnZLjJ66uRp482mR4WlkoessYv2OCf
1hKkvSlzqvddghD7y/TMw3wSD3rxzt6eSw53CApORU8Fiz+D7Z0M8x2Jn5x/NsKb
pvtgUcPZk3uN2YWxTCyiezbAygZSpf5t6uVmEaWDTBGsvnEXBzZ93kogoWpaAhwt
9fWqHfSngHTfLJ3T/Uc6GdgyRefMphvkpsUd+3v5Eb6C5NJ5eDmwGaH/DC+MMbkg
dcVOhqWJ/YiBzTJZ2sN6EFZL34PyH0m6z+HtapkXKNG+pJgUBg2HDUZhIwhCQuQm
szBSFa2BnhoqmuYZayeylWN02/9rIdhjodYwlXiDL9iMIu2Xddp1Z5ZJlZfwZszN
9/NKUHOicM5IKpbx6p5vKaCywgKVK7A8sJ+1LSTs1RK55I0NJa/hF49JYaaZvspa
1KITIIQxXQhjj6317dvXv+TffHp/q/DvoVVby99XB0C2u2uwSBzTKzCkWCO3EGuK
k6IShhLNiSLDuazR7qSFlgtyngAjgLXUcsgLIuxpXLmGrWGNUa6OnYGY5pR7Megi
XGLK/N8Imn7Qn5IwjjmjpNimI66sNE4T+Wo1seA/1fVmUK9xOoq+Bq5Il1SFI1eJ
Vi/Ecj5NOhHPO03wF4ruNEDE4fM0ZePMaRJAoXx8t2hob3uqi4tSyefaX1AvXaN3
PBx8SzKC44G+2Msc0f8MXSh184kBmZyvEZzNEKXr/VGqvL9KqsUNbNU1eMkUEyHC
jfHm27VD6dGMYGLlf3MS/E+2deNh2pveNuM38DzchYjHh4FFkeRUnFlKnJoe6SXm
sbh3B047CIr39kZ9qnUps8DFZj9qUpYb2BDt7AVi/gVahSFquWyBhlHrYgpkQg1H
1NwTQx0tvucUQ1sflqS7PPl3Fm5weKAn9XAcvOrAF+Ih19krDfWW/W3Ad6d4ebvr
cHEvSb9O39zYbFajvKToagXG3sJ03QBHluw3c32NALN70lUttN+iqfGI2ePlQfRg
vYvf1zdAOGl169Cq6qJH6WCkUCMN6qwArtmJm0cBQtX/xvyWrgRj2bNlaS+xyrub
2LfWWUAnNFNG8FFfIOq8+MiPL0ZH5twPVOu7pWAHpW+nNXAcZqqw0klWhZgz1wN0
vR1KVPrPCfiUldocU5xmM+bAQzlPvwIspwf1ctGC4AskPage//ocoVmfZ5yLnqAv
XdG6WmOAIVhzCBx8ovgvPKmc5vToLxy7jPGE5uSuwOAqVY1+P+2kuxzMmfQuHjkh
9uw4Oq049lhJ8Fnt2n8F0NM1kIIO06WY4M9Auc/nIoVYBEdgezbMkAtfiyB5OwoP
WefTp9C6uImtC68BTbcXcuv5sz9tUBY6wPiLqC0ghpv6hoQ5C5P8d1fzhXQ4KoLk
wzckxgpE1aZXv+P7Xwt1oRberc+5RKygXE4EBc6uFuEPYJBZDqEWX1FFOT4N6m/D
8RmdmK47MfthgWVQq+SPu4g6Ba9bQg7gZX2F0330bznCLi6YZv8xTEHpk1MPH0wR
UlU0Et2h3FLqXLy/DftkH7zluFxvRQ9ybUgBELMAJZYaDWx+qMQWl/PcsFxqnN6m
Pxgi61eZwk05cYqiOPfjbrgQM3le9UA5bfRXLOYb+03e0nJMKhEqO4Lor3RD7O/M
Woap3+l5zr7Gm8zGdfBgOsz0baGhrrTJPruHs+Z20rvFX9zTpDTYhL8LVxSSoMSu
s4UM52XEg2reWgRr2PT+yBxiejqKz2p5ExYUaEafaEG7rZDScXLG9oBK+zHexmcv
9Yv1yBYb2i+romjM/Vu8bgICde6ASev377zhHeb90elkxlnnofeDPqEu/3zmsDH0
4QZRng9hbNoWzg3V9McEFiQIzjQ4B/W5CZoOzQ3yMH8en9sJdC/9NuXn9D/EZHEn
vp/FChG5rfcdCiJbUZpE6oisxKsOqRr4nL96KtBNI4yhAgTHb/4MUqhDyVoLEv2j
XyyWljw+IjMt8UgZSjhUbA==
`protect END_PROTECTED
