`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RAt6m9/fjyAjghSbTgAT70bgCr1P3fB9o5Yfh8vJZHFLDGXHZut6E8fNJkMrq+Aw
7LtLREsGQ2sWo19xJgDtqBuFTwAh9Mrtl5lyVhy7k/3JRKXtsgTdkfOd78Y5Oqz0
d/DX0QEpU1zV75wXFMHCG8uiPq5jyvoZQ+D602T4au3blWx7uJDK/Osx/iyB/9M7
647GBONIuhTJ0e0RHF1CztGeF+eeLvoayDiojt2BRWLm7kvVhEvx7XJ85tHBROLT
ZKJ6xAplobLQmy1f7kqds5IRqUO+RgRli4V50tLYYrDm4/b6xZRUfcIQuQXlVzdX
GLrWRb5xEgxsQIqEtYYWWxTXm3rUvg4egDnooKq7jC5iY4w/OFV2Fd4kTEm1GRKb
73uuJg5Ahu+A+CcHLljy1X234/VowcfuYSaFecA8kwxpPiZg+3VZVkDEgCKuYedn
LQCmIZiVbnzjIk7fWd6/z+XzTqdkGvSDvRTU032HHLCjYi08qjzrQZQaKfmM1zkV
YGk+V1XJfEM58+fLH2rd7a3El71USZwj02wPIVigUsGqrDW0bBEkagiT6aPDm0Cq
V8o9q2Wx/yOzTiStRuNM16UNwIq7TeiiTtgDpEPjjKAvTN56K1dlog3/h+vuqZ05
VK2u3q45tfhkp8MIEEbiQge06O+uhc+/7ohoxOHFVFi9AHjUlnViAPXbzrC3daYU
mOiz3pOA5wZIlFuhCNqCmNC0srihTax+2nXsirMXgqvOEeNt/yNrSzj+Cp+Y3JBp
Ia1JRgrEQZDa9YhJ+LUv0jOO23jqzKnyNPyiAUSCegNZFITYy7Q1pCLwvz+PUVQT
qlKmjGAX+Bzoex7bvBD7EQMz8X3EVaSACwtSnDaBRb5G81SrwwlkUJ2DWKNqFLvJ
azP31u3CzlkQMOp/Bi4mCyVqoycDLFGmz1V7/oWMXSgM1WUoYscvPBJSP+mdIuhc
r3CkwMTgbSrvL0eltGzTR6LKAA62+2ENoBBqB6Lcq/3pLjxrbrGL7HZazl/pRHtO
9CkY51p1aJVDhfBVuVYjPVtv9LkTVZD3LfHSiO1S4Ak3VZHuXutQCAjBiQbb3hAK
5MoFfen7odxyBhze4nukINi1APxAuZlOqd+0gn2Y5nViMeiIXVrfSfBCqCTkJcbM
4ApHiHZbHJmwc85eTd8z4zIEne4qg/tmLkc4JoUxjuPJNfcfZmN9/2d4seDNhtpw
oWXSByoqaay++GhdPnA1+iMDQAkb9Mpn1y9KrHJ15hVcWRqaMaapiGmgw3Yk3kpR
BGxdgtA22yI+LuhPDjj/FrANo7XeAwXwTjwA+o+f0Kony6eFeSbjzJ4Ysnb7gsR2
UbuNRbZJ+Quj/QCmJfXaQ5THXwj9cZ+vQj3O39Hgqb2RMSfH4jxwzMiOicVbYuE/
U/0t/8FeseaTStJpathzpvL9/kWEw8iQI4NyWXIVBedcSaScubj0dBtaIMDAII0F
`protect END_PROTECTED
