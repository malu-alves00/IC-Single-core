`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oX7qiocxakm15Q2vWE31V+F8mgvOyicLXBzRIjQHzCrrzJ6LWD/5Ly8vwuiG8DrS
STbRNjtykOvobKJgH0cj/VsKRipn+a3+WGIVQ4RCBqULCr20ce6Pyk1ElRUkJBuC
EKKmUf//n4N949K5XXxXh/KdOlCnnomgcZl2H8HLY1cPfNzkmiyeUUyGAk3hqGrZ
/6V+Yy6ql26ryd/9RBS2n2rjSb1SC+0k4JVF63ULAWq+umhS8yR+48V9qmVRn36s
Fepwnp2gzVpXjXfFBlnrowyxg40dnVGIeKn7t4vZosQshb9I/MBO4CdwqZHG0kcu
DO3maYCv+BHv0HQMD/dZxM6ylDFy2wum+c+PhMQB/DJdrvQ04Ra7YEMC4FghdCH0
kxy+9xT/6CwiMft5bdgUHPrACgy26OYLupqH/X2wus/RkOzXAeigXJ7D9n2dmEMg
07t0IzK1rpHYJtCFaWIM60TjG18jZdbYvftmBhoA+5g+vSzwqsltTBpvFCZ58whV
rhJX7UpiaxvjELec+IaDC7+OxYpvROAjjKduehH7kEagd9PCU8K83JADnuHn+QRu
C8sOLsDtGlKr2ycBnlc0Q8bui8oMo8QxKWwaYYS46Bo+FsJ4l2rLPzQHpWPhpCXw
a1aIGqYr32M06V5rLZx+wxGSlUVxAg3b54j2H2KwXzMum2DiPHlNqmvKQWfpwztN
11zwdFflzOP7b+Flk/nS/6LvMnNjHG97TrdMXt64Cr7DfguVaFeR77Zf4seHFLYu
NOSIXVp1rnDOBz7pqzU2r5BfLVja370wK/a2RgnxmFinHKX/zVGMmuSqEbWGMHJl
GPOQIoKqwc9CsjsXAPeUDV4urkvb8MvqR6hyVr7H8A6Q+YFFuzjIuileevSIazTX
rdZGG+qsbG+1HWqxh2IA9lWdXdkHaQgY71Iw30oKpHWbpXGLKeTJnm7Ha+AqH6Oq
l5m7moXb4ELLhpFLgZ+hvxa5W+gPyb3tL98vuV4P96d/2kjfniJv4/HYDzd3nZFz
rHCRVrvwr6VM78mpVapbnWG9xGd8wusU3qTvs6O5okzrDy4uvzmGslM7bRdiZJfB
DeQBPizIasoumYL3sJac4Xo6Qor9hciTJ9RuBl6wZBQRshEDFTHeon+vQg3WrqKS
71DRHyQkEe+8kLoYhDuM/YiTt5Dud1XrFzXbWYwpEZGGfLmKfH3L7ycN0NDoKc4d
vozzJCPGn6VwryTzlBWDZurMvTkEMNDCycRlDo1u3Wlw34tgTnS0EvWSIw3qvDzZ
7krnva2TdZU4dieXRy3XNoGpD5mTuMFW/HPWibsFp6H/SM0FExTxg+d/XfC2UEEw
JFNw46MArSKPXLLevsiEiGVWiLTfyAWdxQAun9YwLgo5KOhaxQU2MQLgiZ6G6Tsp
gc+WPw89xhS7j+7gRB0tfbu7T9RjhkenmgpHw5WSly2wPbqUdpiXhqENlm3DPxZg
AaiAjhKMMWvk69Iv0WaGkgyULQXbXSVuSLPaxkKmJmXIeHzOUXUTKmTLdwkDyxzP
V7eJF2K+mcUpgQgXuXEO3LLpAHUtvJ9tpQuD1oKc3ptD1x3BrsOHlDNH/OSo3MXj
MYtVSeXCCNMEJd+5QuI6oDGhoFlJZ3ngigbk04Gemio7xR0B01BYCbY/uWixceZk
OjyCCr2y4xbj2b44l/eqPw8os9r2bm4nJa3tVP8+XmkOByrf4orQTDpha2FnFWgS
xONfRPHh5RnpIYrtlq6ciCxFe9do785BOWHOeF8d/xezvzNnrndNCyz9MJF11xnW
bKMonn43VDiJeK63ckjlXkqhBCbTJz3VJpcDNIaiemV9La6AySKSFFJkAO0RGU1X
7Dq+QpntrPS+rSFMa4V3lnHyC5vv4J0+ag3cQ5FlHVbcxZQFZzvHdVL/HvoEEmsP
MjXB4J4Yi0lqmpImRfXa5W0LQB3dzgcV2u1f5HP1+OHSUI+WphzpU8aBmgXI/Rzz
1+BZz73AR7m1jcUB5qJnQuaPlWKZsYy3EjS1I9jWJa4l8WorJaiobthA0BmbJ7Wv
dzu4KjCEF8bJYbLWElaJvey22qv7fymnuvqjlpVbz8IGfZLB+CSUDW7XGdYrlpiZ
TlTXIRODArDkSXtI90UUxpF/e7IxNgvZ0pCTPx/4Cg7Yh7LcZNfcIHssjY6kEORF
4OXqsdOnmxTLNECrSQgZ2XJUuUghViTRL6aCCpU2u+PFsYHLsBD97rGcnkj2HL4R
Dfa/gvjl/jgtcHJ0Z+RCj4p+B7wUQ4mMs1KriO+dqyDF4XuEO3OrLJpdGC994r6o
pPP7S0DavSD75Hn2eqR8bdWnF9RjCV5yRwDnPlmTE0bqF7hxVBpWlp7WotvyIW9r
FwDtAqHqNzc9HoWgWDUmIFvv7iD+1alyBHy+OP4/lbms77pTCR4Xmj7rojzlT7cH
OK8Ogep1PzKIW3vkphcQOYHjdi2nbDjiFGCKFFXIkhHiXLItTh8oREXPU19oJjOe
JdXmFSReOPuiLd3U0wXRWPH10t6y1sIUxLo59QAdolRrsPX+3rN5nzuA2+oBSI8V
sxbVcgTT5OAb/x776icucVmmHonUpw4JCP02Ro+X1DdYXu0thx14cWTiud2mbsZC
+benDb8l4Nz5e+0YC+LwVajbPQbzE85F2Vi5i+i3z+t+fFW5ndh309ulAcJz+9Fk
rtENI4CmsxC3TtuH7sM96ad94cXNLLuDxS1itaQGJOLDxiE+NxrBIHjG58dTNJXU
kZ8olIiWNnDqnKR0ncL1E+ZynSGsvuXX3lyTIBvfcUqT0kmVVI22zNMhk+n88jYW
VtTJbYjUInoXiTDS8uZZl0ihJzVQSAk+pDf8/h4prYt40gZj5vLCFzAEqI5N3QXa
Fki4b0EBogu69NkoF2WNrw2q120S7xuH7Ph11pLIe3u1N62jv7zcxzUtSvjQgSLN
jGMcglrOILHKjQVjjDe8/FLj/G2e1FRDq8v8OZdF2PdIk6p3RYcu2lcwm31zNo3Z
aoEsm1no3EbRSjSX85aqvdegWQ8ywmNF9XahQvLUqsj2p6Uv/2rnkkp0DLVH2Hsl
yhCnY2qBlvyjhbPEwY7cm2sfEds6SdtrjzUvv0ZIwOQtHbOLMh4GvbSD/r2zZEKH
4Op/Apl6Z3dHDxoqEORFnIXW7MUbAJPyQzS2b3tJMqUIAY+zsViQfBVwGlQ4kcD4
jRQKmE4qY16twQpkqXqcTPsPQlcwUvdaoBddrpXroo/uT6JlNb6Momcb4+J/LaBd
bpgXP5TzvGqL30qsLdInYko1zDWqpbJgqLzueW/f7YSoS4aJQD5cGsuxpJlmdGQF
i+fIXb+0k5y2XkVH8v5CT+pGRMHq1plpUbmYbb4LEIKSq0lwPJdjrwSX8DaJiVJA
2Z6cemfWy1Yra0m90MAqRVama+PhnZIJtWVysrS/6vGDkOpyN1L0fyZ8iMs03Qws
JANkV8nBRtCvE/7iQKXWtkUOTnmxH+9BiYRfryLoEtdjT5RjTTn1lwE0M2O1lYls
gllQrnkRq0k8DNJ27dEkNLrWGTF9tArGdIy7gZHi1+OnrD9PbYVrc8m73hm/tOgq
CezR+g+3kZiLgLxdEGp6oMeO0IH0XXqp7BDPOWWYKR8fcxUHlITwHATK55Ns1T8B
Ub5PDr09vuLD77y2xRKnhcIJcUvzWs4NUXmEpq8mVN+N0DaQBoiTKZUTLAT8e4Tw
FTeqf+WCh4NYJg82h8beCy4fbvUh854UTMK3EH/3OrHjRVZocoFQlufD8NKLPVIq
iT3qfeZmwWOS3hv1Re+ykAIWMCBiB2S98CvNnoxLJ+SzZUORTJ0B6T6h2cL+Vjym
9F6f9rLbDm21Bk+YkfmMkaQmgh1z9QZrqGIj5QPaABkitb9xEWauWLjbJ3e8/gza
1N2EBFRW9MmpcEGkxWcFC1QU6BGq+pFMeGyoHCceGW4hruj+9MZyizErbzo0QQkc
khOIeURJzPTDHt+hNXZ/Ue7SYld042K6Ct9f0RDpiCeyprNDdyxpso0HvtbipZhg
fjHJYsxIHP5OrSmfo7Bvt2TkYaRs56p1tm9gi8VYTKhzietn2bgAVea0uHl10aJk
BO5YRr57MqLuvsxBEmYPCgwxCsT3dq6HBCZKeQMSsFm6t3mFSsjv70BQYWqKt1wM
/dPpP1VqgNyWcUc0kNgWgyyyXP0HFMEQc10xh6mfMy80Ryf+9kbT83ps0ruuiKEL
TL5Op/7F1AVLVSPCVWGxLYWKUdTnsdJOJ6BV9wZWPdZuwEHof/ZBnDVYHgIJIG2H
pkRe/mp0fO+JSXbi/a84wRDb5R3B5zTB2VF3X6N0YmcDKBoro/kk5mTYT9l2HqTl
BjorQMIH2xikwlCu6yFSePTQEHd4RUWbdPzgIruKEWVqcHP+horhXvDr8kI6ZU1i
mSwk+GB03FiGvWZzhdz1mYjDpfqvipm9HsKhU7H3cPW8n5qBdc3LKRfuDEU2pw8t
ce+g24W7rBqEMXB1y1jrz3M49V3FNy7BoZ4qILcWThgEDzYNT9ZMWr2rtphNb3p2
fBtK0C6SZjo4wnqoV1oV+zPwaCyaw6Gtfp6i+LWWKPY8ZVhXcvaBM9/gqgkOs8TO
rf2jJNrRj4LhFk/jWDgAmRGXKBuxbiadwdHvKOnaYOsVnHgnSy5Or7iRcXcdsi4e
WHor2w00bSLXqjGFnLAqAbsgtkrrl9e/9sORij4DZSeY3IrteVjiZP0zdun2Llme
2QmkwF7ln/iGK+253ywJmsTUndXLQrcY4/Md013K5Un/02QP/qc4o1WmocUSDqV4
Wtb0Jc8vNVM9agY48uy3+3tCY+rXkjGEzxUL+O58XULf8s5PPyJEzSSmj2+71P8C
9sgfaC3pj3n1oDzBxliE0WVMkwGTFZedCbKoXFteB/U1mnQHFDNfou3gkq+t77Ix
aMavmuL/F0SRX/lwpd9reE4fwi/IU0X1TzNajof9o06wrQbbL72PughOzBZKb/ds
BIiyA5PNl6z/vFMLGL27GfuIHD1QK8YXyW5ojhwJHcQNYGdikFVtfTuDrEIBn/ZK
p/Bcy75saTQ14AJr7fQrpG/8IbC4PzN1KmvSBixOj2EQO7FvMy5W2pdbSJE/op14
OK0oZlYtzQ/cNOsz/PQcKRTm3Prmb8UUedAardBpq4fwxWMFFOU6G+dizjF2InYk
hpdMMusHh1iVFjm8+W3VmJtS23W9VG1Ly9j5fkVJB++G1xaPnyh4u22g1IZZ7ZWi
0+jNWLif6xgJsF+qeP5rfQbv30ClbSlxx6btk9Upzb3z3q+FPm4Izx0vLJMqD8hJ
PXpNJNkoEXjvjoMOKSd9zn1PLImfIaKokKxzUwejnJFNm9uULAnmUV4MyhVCXTAF
LTRaYNpHEExX/t55YF+ZErl4j7tTlx0PB7N9e5Ol1lvjmG+RAafEHABHtrRF7ln/
7tDAOVmJXCVqRyIN0wnyxrDCJp3Ab3zX4S703w9YsPjzgLtD3xGC9NAT7E2MJ2c/
tFrP1dpPg5tPVfqvFI7V+wlCFnnlJ/C6bjgmeZCj4nBmviyd8PrxN7hoypNuieKn
0AAUnWRTQ3FZm1UGUKbOTStxnAZ90unagJ5JQPLEHX+ssSfxxCyPSzdzV7tjzMeq
eENcK6ZgwqD4oNOXYuqsu/pP5pISne2NeTHuWMKlW2SgF9zhcAhpo/EUDeK3gElR
y4G7ryY+e41qI/hZwHNYtEvM88lCgOWes9YhlKkokfPr60db2tcUATsl5vpDekgu
u+Ralp4tKx9Qacujdm2qV7/e+rUiTZ1/zor5xdFPLIET+N8Ht3hg4ekl+pTtpPfA
unvcFDM4OF/+m5eOQWRjJAXRuYIvaj3pG7cECB5w9xsDEUb3dPxwm+gF4Q2KB/0O
KDlH71LCefLiwo+SoRt1gkxCcywdwuBvGR6ISOMRn1nijI8TxRjaSH58qoeCVrGE
5wFdnTB2T57UWRh1ljEkWx+MCW8JmuF5Q3ysFR+FwUyaZ8IwA7zE9nAKP71FtUO8
WvnYa8CV5ya8zO9HbojH3jRhji5S4LP9R3TKSd6u7NhRMbT4uaNkHgjLZ7CZISrg
iMbouB8CUVbPxH7PX+p8R0bNjc6cXsmbhhn6RS3HbGOKWlCUniOWMA/LekOpjs71
d3Fp0AvH5UTVp4f1TOTAkJx1J/+9F04lNPVX1Q+Iwob9hb6cueURNwQPr/sh5c01
8+zJa1mB/a3rggkwoS6FfCE4UF1CvystJ9JOoaNCgWNf8LNavSoEnGzAHaP5u0yK
S/iTDb4TjU5IBkLykfFZEtlavPr7hfqKgKx53QQxzt3CKDyWREHMiDCsOCwYyLHo
8bUHKYY9craEW1p3pS3W3f9mvj1gBdEZKkKzScyYyCJNAZJsLB38CvByLmTui/u1
KOJg1cvRwWJjhsxrAi3vE/RL5IEGsTn1cltvttkj43q9b9Y7osYzmMJizP0Ncv1b
tfDUImoqbYywRDsZuL2/8YQNDWW2oGEXaU05MvDz1adQNxuVPRgDGHuqpVyT6Gu1
TaSfVm6w1UseGfGzqxiYS9Il75CEYI+tlLXAJTh81jvewgFcB2oJL6P1sPPmCsgA
YnSBGLfsrmPligQzk+6sUkPS151chWnsSTiIL4+gHMfNvlYmcxM2tyDzFUDFqSdN
A+lRYcLY+oPvty3fB/owDOq1PToY0hqG4jz6ytCHFiAF13SUqM2i5SRnmJMqzyQu
og8ibQNqVKSDk/b+iDgSfRm9YeVjD20A/Jrb+Rkx8OA=
`protect END_PROTECTED
