`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DFeH40hafF2OJuFgp9qTd0HcmyMKXN1WTl7eigLR8t0cey/Ifnoa6q+CdUih+h76
vAjyv/ZF+Y7s8P7F8jC9l0FD4TCFllyrvqu29V0CfHILyzfnc09G/8g6Ngwfe/ql
YJgLYqV6JiMZEoX7gtV1stPLLz8N2Mk26utSaU8jWZmXz8asjzlpGoxDeccvSYB6
AATDVRuijwiJFWkFK/A9uGpwVJ3f7iHB0OXUouYIw3wE1cc3uXUDbzcHyneMxPJv
oTAyMFSQdS4Z0WZ8So+ZzxYv4tZkRO38lkAwgaR6P1gYI0Z31/VMYOQ0kAc6+a5X
OXIf6kkwmluLNcUkcTuP07evsY7cpquF32CXNnwgDrmmoG3XQkDZYeDXwIkLPUGs
MSsq6GM6XMPZSZCiG8V63hm5ue/L4wPMP5CRk+xMhdwOFR3UYAI9gV7hp1QNasb3
NBGonJBdjLdLSBNu8z7KHHXfsWzbNHj5o3DHnwganSF/j9JBbcxn4riqaOmIRihg
7RHyuCldgFDEPB3nxu7EQNfYFVUKkc2mqyEU6RSgx3ZV8HuSFSw91lc35oO4Q+oK
JvLXHdR5cjfpLRWzEsiIYeQAWyJyyVziZF9zJuHRYv9NTRjFQyHCNv5mNJfb1HwX
0E6ctZo+UYsRDC/4GjPMqG/2odPewy4a1be8BWxYOKv9vQ05cHPBLEQoSde0YjT/
am/qcvZkikqfXGkPT8rLNSKuE3T74EfUD0uJ//mn8zQVrAt3TrESSwaKLf9Hfd3p
LFnDCQlZf+jjwap9awG14vYfl8bLtaINY1XwmT3QYk2KFMO/QaUsiTwS8wravmch
/xC8onIvc1Ow0HMrq9G6yBGcDY17L1NVIzXcfI2LktZe2TjPwqyL+np5INwhCoCP
IG9MKPp87tgUm44bNNUeWr88huCFwd98JXjQnrqAljL0giJGBpGNsSpPA9NbUSd+
acY9HKF4R/R2hfkLoHzrttgGKGMCYmBoAwzIvrep9bD8eN2TsIXr6g4ErCv6XMDz
8t1seigOa66EAFzX+TqWKU1OnU3fkrQn9WfMO08UypZffOjnrZeP9qdJSvmdfpCl
rRYza0+Hu9yL1QiNyobXRSEJEUjDDzr/lOszpVQimz8CKLSXZAK7vI6+p2O6B7ul
Suuuelc+s4YRWOUAANEenBtqYlrfC6mdw3MJdQPmCSX5aqsoAg/Ng1YnIo0v7aOC
MmVdUbN0oWT+TFfXo5IPhQ==
`protect END_PROTECTED
