`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QGePZpsu7o50Ny+rviA8jaih8xT9Ymsv8TA2zuojBcBL7Fakr6r8ccILbLLjahDG
P2I4N/6Z9fFYxIyd3IKZ3cx8Z04udSuEJjrrnmVpfgltnBdXcmSbyKmAGTY07orV
gVr9dd2liTYwjI3UEmxy3fiuPm29+1hupm/uv7B8p7ePabW7bdAqrpe7UAfFZDx8
ZMurIB5L0W0KMII2ae/becEBZLs/QI/jeQB6H7/6yVPN7K4lOF//WKpAoqCnzuTL
Vjj1qAa15UDckfxKv68rU2I6BgcQ9TBu87PTkfurkOj8kPVTGgwJiMHEA0Y4yt8Y
5ncVMaHMwwvWI0btOQtCmfRHQ/nT/b1d7G1M7dTRKR86Oicu9i8FQxuIGtAcHH2f
s4cBmxeXbfrrIm6IcQUW5LSJMWDtfo14raQBHfuFK4u85emZ4spS3RM3YLISLQOP
r6XgNhdJO0LPXdRj6owY2+ju82+Qws9ZycXjFW14hDh9lWPbdvC4tyv0KQTbCF/U
OjG6Lsc2Hhb2JFhnRo46lEdTqmGv4cjHR3La3+E4vRIIGNbLvSj5sW+X1oredfTo
Boqa4BzuE+rkqqwk2I1ntaWnHr46yb7cMt+oJ6al3UCgSz5ICvWeN5k7B4bETr2z
rmBDk6dMh3tmTRoeLr2N4oATAZW6bkDtGd5njml7lil4lquHdAkPCTDUU7u2ELlR
heW6n5DkbydvwTM9l2YA1uDFbdHeEHLcs9qpXeR1VMXIg4nB8dun3qucDvgpSZyL
Bl7f6a4scMJTDkOh3XEBIL5bM3DxZ9r2kLFxgvUKR44=
`protect END_PROTECTED
