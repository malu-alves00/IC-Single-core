`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Hd5zKqeBrBWMRLLfjpWkmeKoWkqxeJHsvO7pyc1WOemBt2iVj0mKQtqgQ1egi+ZG
b9IcIlWSrxlcy6in6rO2kIz5tvJCCtZGU2jcKcDnglEbLsUE1maZZg4VJUHc1EhD
jgMbuUCxbPdkg/0QAbIrgNBakakigm1M2KDofbzTNUrr6HDY4VdUOR10pGvj/dB2
nbzWhm+147ftRPJcvZdnPQ8pT2xXiseOE90deyjeYgTD46fbsstGAUdGAfR6ZRPk
dhcgHyJZ3b2gx4yRNlVC1cZ47Oe4loYmSy66MZwXmwEnZNZa6UT4eWYt/tTgfBYt
cW8rIInJpS0JllYMiTZIQGSF6A9a6YTH3xm2oSAYp/8Lp568HUzydoGDnGF4JBon
`protect END_PROTECTED
