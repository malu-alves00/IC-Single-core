`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
z4w96HGAUPDM3W3SSUThxSHelcG4JbW8ZdihhVzp4tMq8ZM4c2aK+IW/41tn4v7L
cy86Qo7SElYV8PoKtPX2OwM3otSZNWtGHh4RPq/MmJWHhyMYXmLb+tdbs3aYE8wG
iqYUTK6UH5GlhgSVvIymWHCT8Pj1B821pAMCKXN721IyNT40eVJzQN/UltHveMNp
VcM3Fv4vo6mf7vhTBJNFOoMrTFAKcT2llOnpSy5FGSYF0jtDxj7pIw8H/J8QWcK4
7W8TlzmwKOmQtlAiSSaSqVln+a93eeCQ23KoNkCqch6GIDbGYrgwPh8KKSe57oWg
BtqpJKMAqXgWbZH70GQr31uaz7/fY5hTe0lHlBtdOcDb1b5tmRQnzz1g3deAJNy/
DbTfIB32rUNxFI95hUOdnOfS2CQd2nHO7hxqXmO/PqyXqcCj5T0I0xDsoR/6LijP
DGTnQphp06zymlzeImLleL0yNu5fH9XrfSc+W23xRZD2QhzEdOCUURTCcX+tSF/r
j5vSXsKcLy9fJmJNN6Of7euZNnv7aXl1Fnd5YhruvjV8xyXwisHgB0dmGufdxfM4
Ql1iZAfi+lzysf/sotsNuyY6pXpDbe+TWl2e/XHU5VW6NkHCZTck9BAF0+XP+hzF
6AbPQ+nayu/icBkzMPYd43nNBEDqesiZzdU7IZX58lC+YCdg02ROtLKT1WC8Lf7u
2plwndY+LTo9bosszaNPPimuE7syYp5NNPHGUhG8rqN2kWo2LHGMY8n3a9t/jF8W
gKZKioqINBSYjrCMgM26Y3TjDSWnXjtcDHHX/33zg3jxTgkT7griyiS3zOpzsVKI
eyxBnTypGXnaq4EXdowrJx5lputgN3/TmDTaxakaqmztDB+dTVf2U1U7g8rjVW45
ErKZl0o4JcMwcIBPi9hzEgnH6XIMug1Gh8pMNKOf2j+hJfqlldEhfy6gTfcwhLws
s873UDrQG3J0RX1UN0TZ0TgXjTWcChovAR10bJX+6EdM6Z53uFUP5Gzmhepa+qmp
A3ttFBGW5G7bE84AY8P3lmXAiZjAPG9vckkGUIl5qqSh/VJ3ObSWvORxyhwEFxJN
iq5fCIta26eA7VgS3Lj4h+XaIvvaRPjuKDJQKBT4ZY3Yk7i+s4As3+ryyysIihBj
3yPZzxi3ijn7cGkh2HCM+Fr2tS1OMVnKUopCMIAoE1iqoT70ucBv/fbKHOR7ZzyN
bNszUX8SazOGlh7+k9qWCPh8/rJc6xOC8gb1AeGciPpAhNhtxtmTIxqwJJHMMEbp
ilMudcOKkNXaxlNy3xIHMnv+wEFY7o/CA2/dTGXKgJ67Ke2G4ZG7z9tff5tGL0hv
qloZ1dnTSbevLyRNNgNyHZNOjkOXwwOEyao+9Kf6UeFdwyVM+QD+n6CJ7yjFGa7K
ExWCS0mLfcKDAP2oDLEmJIXFLvFnAgQUGXj5wDCsz9EqwCbaef9UgkooUH6oq3AY
t3seWu/lXFq2++CCyP1brsmBtCwuV2LcgfjhM0AmldjT3baSeKJWguVOiTPir0pr
j5QoRF6cW3926lADQdrAWQqJSAdiLqjGySrBzk3JYoYVlIpZC6vgER4/CfcEHZbw
gmlLI1k7Ai6ZUPGIfKTGpauPvTnI861ip4T9ivWBA5GeW6ubc9yJLOw/O2fb5jPI
/kAdJL+9c6RfDS3TQtckOKuQPbC3khz+JPgt26NXsKDWCytgqD7OHVMBg5pqUJU1
Fdy0Jb+B0qNKfVyolLeRH8oGUG9ZzUNeFMgmEWX1Oz76/tw68luxprPx8Sw7D5Vt
Is2lTffbp69JlEqtaBYVkEkXu5N3+dcWAJ4OkApP1PsN9MhwdUoYQX2D6dbvh6iC
89EFjnLOVH2DUJ150ijQLwj+V2/I7NQUSIezgyt4XMvzl9otUIQKglu2qYa623Pg
AgBPbkjEMfuxuTDwrnxlOe2LSN0GJ5RhHa+8R2zhAReB/AWYpktfc/8Y6WszjZiy
NIO3ZMPh6KoNzeiWF2cKFDbG1k93NSt7Hsd+oAeYM5pV1xHXxJmUprVyu04IDU/6
MfmoC+I7oAm89OaZXVUs/vj6AWDUP8onVLos4qJI/V9xiUfixP09yiezuDQLPpOI
XzUkWQOJ4+Y08Pn/PhqMQd1ZQIBJ+R03FBc8M20itNADqcGiUQmZ3E2YGWpBx2mp
JitXCsxMsN5KvyngBYbXzpSGsstmm4eg9MFeC0T/WKEhO7+upMGGUspB+jJirs6G
XRzi+A6rG1wIIyQ6m1WlcJs2VnS0N61De1arsZ67vek+VFMuw8xWQA7mjpJ1Cv7p
OH7TkWt+TuuDOxkby/8o9oRNCDtMpD/YNbb0bqwLzBAniTtpy6WOFryEhJ5TiEwc
HxzEO5uBjt9ONsPkrm3PuyJ/a63xsLQFuY9M1G6uZdmywFm1XOVvnaQd8Uk5YiCQ
e4uHCtIaCgz16SWRjsWrPv3f7mx5RCzYcUgV1A3LsPpwORm8EqHGYonEEnTjjW2j
zsqDUyHQctVRUjkvXqV6kAErRVIwMSwJ3kuwAR+Z3zz0+NschgUXY5lv2KgctRQE
DqgF9Gxa7GySUA7kYSEEbHyKey79UOYIoaTasGEvX/q70qY4RQwW3dE/zr6/ch8W
jp4YYcgy9riXff5i+jNqU3g2V6f054K27REriw77wTdEkkZ/P35P1iq8JxSYRK4T
HWbgXE52mnW01Oi6imjg4aZR6LIrq6P5q2WQteLwEeVN3mQsThuaNreuiQ6ONLni
hdiE84uKMYG7do3cinCTiHoDMEeZfM0vBEKLSIsY0FODDJ82tp/7vU7UF9zgZlhN
YV/uwYFx6p3l8qpawVooUE1M9EtniHViozSvf8XJsLUM0wDxC6VuuVL5zGo/fD/P
twmLWsKAcjJDi5TsCwFtV9eiCVLvvBaKyphV8JeRmJvU0rHtlGsS6SSs4HeLHfYX
dPieRbG85ZqKihZu6aCP49tjfmwQ5lHLCBtGDdtU6t1le1zviuy9/dvrF2I5q2/q
FPaozOGoMLMh690oHTxe81+2xIzgtSVEtcsgo2wGHf75Tx4nCza3NPXB/kQMNhNS
5KjQUSQ/cxr4D2fEYlZL6t4vB2SDIsDhs+bqZarFqBl+ad82mC8rOs038xDbx37t
oYv2UtNz48uLuoSD6s4lodw80w90RuYOFBFzJLq8nfTQoLOD8f2m1wwJtqS6NTtl
nWLpZsNgyfFoaLIUczfCgk/4BdVS34VXiRP3zb/fQPt0b7Qdr4f436bmH8DYRxMu
6CpXciHofZWImWiD3pyE5VNIreY0uF6QzuKB6Ggr+6ZLjYIydbqtE1M7PoK8MVAQ
Rot1QJGtp+di4xsDIoj5AsqCfHmUgOSuc5K+kHhQqgSS9uSYEpRWWPcesOGeEoeK
GxrPAZ3oPx6MqnQFLGdRQvgdFaVgdVZ8QhXv6JQj/+MwLpWvKFpcvV3RFZTcHmf7
F4ChApG1IpcBNt3rdezwZS6f6wK08cBdKnYwfRROiSva2dbB1Ozn1gmd1cezAo4B
9csvMVf5oYhHtTkFO1SXchy45Vdu05gFcJ8AgDrZwaFCpqfn0mrogHKds+3ud8Ce
o+XOTiWKLwdaTW1u0lp/DQTpJsI0JHRMN8GAgrtIEFVbhygXZBw4R+CVd5I5b6Ts
SLJLi2WII/LIrk43pOQklDbAi1unKxiUjJ7DYhG9M6/NLyPrv47ym3XIfvq1LYW4
`protect END_PROTECTED
