`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3DvNlSQvyZW9/DL7PutCgd2gK9zHbTAsw+DhRk1Z6tbh97O4UOI33SN9H8dX2zMJ
92fa/wGPzr9+sQ/5YcdLqB03GMM1K6fXKaafSvDgNGI6p2Axfzm1+JuXVpGE4fUD
1dRTjjgjr7IxXVzYmYbmGp6UES7H3bem/6KibUndBkLbNLgn3KsQQm2uniGeMsWl
Zdd98WuqOGAoeM2+KUL+6ocE3JqZn2mGYG66kal2QJw8+6k/2aEtmQN3y6G/oS99
/JCcNtJMz3a+jvAorH+oN+Bq5OUxZMsFEMi5Dzz1qAkwQUchYJrQTEyaqF50hXOT
ZJLGZ1B4gynTn2dIgFM1RCtx79YvclaqN7NQQIlH3oVMOpouCyQNB7Rfl/8jjY4K
jrsxDBJExGA4Ww1fNW0I92IoomPFMqgp6kqbI0jnWLtI7Cc+wov53xIfma4wG/0g
zWx/ZcVbrxPIRCCu5TDRMOT08k080phWBBkxcsc3BrA6u/AQoUPAzCPktaAukmE6
ed5yJc+a+Zyrlr30Gymtj62wz9+wMZ0v6Mu0srvmJavGD/5mVK1gKccztQJh+PUM
aRTVHGP4f6X9+YrW7DTB6fHFobv7YebBfMV9g0GZb2Q1PqdjkuwmyJpwemvmCeG+
e9/Ren98vFA+sxsZhfo3x67v262P0SxgNb9S6IswYi8oXOUwSmmdS9mCpOCwSkDn
ZRvn1n8PhFO2KNT+FaokhCt1xJbA9fvkJ0aIcONI0OUhUxR8KRBum6+yvYZB9Nbb
TPQx0qcIftbMPDJVd6qcHxX8hf53QB0G7gJaMhRYQcRz4nW4NGYMKSgou1GQl+Z3
euvbMZCE/CJH3yH7Rgc4eeFyUgUl1S+w+Bo6Rlle/Qg86rFNUErZo9BH/iaX6bwy
54hufur+hHgc+lQ9KbWfGpa/doLzn7JXkYKxLvhbuzh1i63aoEY4NK0C59amriRu
CvC+QFgGyPgFKT09wkRjJ69D43ZBvJoQMj3oVfybEhzB+rWDbsCIUpB9blqRlyS8
FjaCdP5t4b+QlsBxHrynAG5hDYIsljX1/7gLVfjgrTI/ei0lx2sBkR/fy/NJWA7+
eKOAHDg+S7hYAcKdjYg1+mrmrtNekXz6C4Ma1rAiD1ySCEe4LRLcuLTIgvKg6XhE
anY7FArEhq2+RIHB6Qofr+ncvuOqCH/WQwPos5dRVKJS+x6fv8qLt1wCcHagRmUF
lmEAq1C4F55lpY2z5J9WicZ1rDNcjYaFbDnCj/qg0blFX6rXKHlPebUcmbRYIo6L
xt7GLIK+ym5RdggmmgHnHhEonwnmSbD4woa9SSSgkyCSWyxtYlJ2nHBhIZBQ3Paz
UXC+K6utoZdeWGFRXuPj3eVDzd8rnRsOCCL9XOycToyeIdkDjZPKFL4C1IeeRvyA
OTYNQ2h1YYXH3EXHDLiBGDP7slVFw4AxOc0ObnnQOBNYsHtv1z/ppiiZEW+h5FMQ
hkSavqnXZya2HUZNx3ReSWsEIz/a85rl6auwqh5PZwuJmmbzQlBajlP/FuaFO3LT
cld6XX4tRQLBnx6lZtViUmLL+3lqE1i215fv1qGLSuClO2AOccla7tsKK+I6sy59
djkYXfDv7kNwvqCojot9FC0EKXPPtwcFmggl97n+acttOyfgiLYlSyIH+0HD2v8+
7JPZTxaPcY+J26wkeA0SxXTzIuclqFw1/AD+Mw+9kI2aKUmrUeLtTUZ8G6/85iiH
Pz2hCCApwfpHDN43S20G+q/vryphsghGgq/cgG5ak5eOuYXGWAkESFbpUzsDAU/Y
6is2TVVQM/aVuCTHFKJiE4qKzXmIBcn0g6HvTKzew0UKcs2bQs7xtt2CDKuQnUYn
GahA/Yj+QSL/ImjWQhlIbHISwOVK6IcoVjEVRX0vZ+C42Xl31shyEzz9BKFvz888
vvSZB7aINWTSZeM1NRb1OSTzRp9buyGn5BZBZ7leYf7e9JTazO2n9Lu+G5A5E0yp
UM6MNM3TpYLzrD1M4fGwZulEmCT1w5gwlcJ189uL0dYexdoL5MJN1pIC1+vrshsi
4P5G7/P2zgCdm0ZS0DC7usbcPQBrRHkG4XJxoMuQ3QijC7MOFOdmLJrpl9oODR75
D9jbix5IXGcoFt6qTcn1fpp9DaEccAGalldTl6xKHPrA9ftDvEMZ9kSnWOx8O7hV
/bJjfBqwK+3vAp84h2wMLrHAh0YKCgaMO6VEpA2iMRbdvEE9+ykDTv+N47HrK/US
zNZosAcfasUS7EpG+A78Zw==
`protect END_PROTECTED
