`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
brIf3wxdnLdqDiX3uc5fEegT8uq4HjbKESCxyQMlK7D1VlAxBFxX7yxn113sDJV4
s3fsZlnFZJZ3jAMr+n/bl0bAW7mQ0QBOee2fIf0kgi0kwLDmv5smsI+LDLWZId2Y
8PkaWzUAKZeLm46b7FXmIqtr6rIkknpFhBDnsnihqkWEhMW3RmhgL0gjAnnfeLY3
nfn39r2dfqs0782CQTaJRtsfft4EFRDcJQWpIE4D9wY3Q9OfO6sZnpBlb54LfsPr
/IeSZNVby6Fc0UWuRQ1kFohk57ah2VwxarmOoYrUgJQkIeR8Am6p898QmCm8dWDF
hCGmiEPLoWDQIEU8Rv1CFNLXisjEX+7GbRBlbew7GqSxZThx9aA00wX01IB221wq
UbX+1GJq8ySlR2Sii+J18r6ePBQHzFQ1oh7WhorfLQVH/L+K6EgzIWThXy+Ro6JL
p6yepLJa5OkldFNj5DQRCDZIMzJZgnU1avsHr6kqs5DAGq2TQF2VmnHPBsOCDbG1
ypkyqWM/6EtUX0nGG0M2FXgHEExW6pwt/ByXe/ZikZ/ilSnN7xC85z41DU0u1eo7
dO0g5XHvJ9l5ljmd31wGPC7XZP0zSglMIW9LqHP5I+DFeQ1F4qNCw9QgIze32TG2
HfrlJxus6Ei/tWt/4hGn4oORKrycQ0RoF2HiHq26s3WqMBDBp06M4EBhtcZWatEm
1X00R55Y3b2h8h65mhv5CXF0zTkwIqPJqaAsItkd8qrtf8MfG/Kzw2XG0Cf00xTt
vNKmiEEZFslgtJ+tOpBFne7neIE0O6zDbh49B4hX2W+Nr+pm4WNUi6do5lGmp72/
bnqlCbRLX9/Cy+7wPFNPo0z87aErxzea/7YHTMFQ0+zbBPk6E8KnD0M7z2Xs6Y35
Mabe3cVwDHkTlD6eJBKVi+4tlighRR05BdO5A+QBYDUp2PWThw0ebkX8Rgj0Lz9K
`protect END_PROTECTED
