`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
u7m5yofvN06TQJOSgmwLiJEj2SgW2l2+Mo0VjXI1J4wyUv65LkQlHhViFBeIyFL4
3mq3SK7+ZeY5Xv3FeqeuQbGSc/7UIy6US/xj7Urs0mEjRGI0TzXhUvlEiidkk9Dv
UMc9V87xj+gptAhLgotZdKvK8b5k7GKDgxoVSU4nG/BufudjDKVYs4ofMOiIjUWm
ffTgWQdcrB/q5UhK5CqePyoR8P00V8JPJkZt+i8EtN3LIkXi7GeLcvXRVpV0Zdis
CX9JytyvVWbhejcpn+GoC15J1aVlz4BCkgV/o3qYODfPqa2AZS1Xy8qu6gCW8EGQ
kbW/xedK3E8JVttQmYVPHca1/bvDmB25uYf4UlZ0LePgSNvuh9wC5krzGIncugDN
amr061ptU6g3gbIg8qUtqECS2d5nNJKI3yq2/sAu1QIq4DuS57MHyputsHncv4lY
jmBpSLOxE1BwvQOfXmCr2wYpnPDaBjShwY04MTdhWOzxnYL1eYs4nUt0SSJnrSp/
VF34wG0FXHkasidetnHDYCHombUUiw8nAti2Zb+yNZXM2P+XrIkubw8xzcGe0IAk
G3//w5NQkGdZu9Eop+Tea8DZHRDa0mT4kIeurHmB4LEC1HCPEKVkBUi/ABeUFxRd
k8TXQREtO3TyyJrzD4+ozQIPxIGC/ZAQY65AqCvCYEwXJHTTv2p+gX8Z3hA5Dhtp
3MdVzxkdXcGshj+bbfE4Cl28BpE2NDjHlKsbnMjBIlwzxLIyo63yEB3v2sGKddFb
Xo71/qInCdiFlZ3cN335LCRAzB3LKz098cW49NFPwSaGl5T+HoaPnQvgrLDe9vpV
lfluvRrE/rSduD0Hsd11Q0ZQIqA5vbz0h/GtfHFhhBpp8Fn9/eKPdN8eQLmBIacE
bLA9SMig68cvmDO9q4tCUBtKlPsaCSSJxQ9byj0Gzw3D0CdOfXzDq8cIjNm7KwS2
/dyb3C88eLLqAAnUw+cPNSVxJLhhaLnI9foT4J3fRCvkCRot8uvtamoLl1MEzHIp
zMCc7dLAPKPEyzqOumchNFn9RZwYAWqxQBCHa3jydiXEjmzHzyfsxKDnE6QQjSza
yOJgPQCfaQ0MDnTO7TjQoJZ+IrrtDVFkLM57EHP7tDMGx7iO5UId01fTT4d4mfVQ
sxN/eWtjwbv4DKbGa3xdGc+Ja1vAbOF4yIK/hPuqiVO1ZRSumn3Aipd7rD94+0us
BMGjh/pler9PTw2552WEg5O+PezuHJtjPiySPuXZr5vBrWP0mJakT6KU9wPCD6rk
K/Xvxis+FJcWZcsNHU7BOehbhuWPNS2CfXTpcBRiZydj4aT9Juqp8hwbZ4OhUnCl
C7RbudWKSP9ufCb++nRIIj9IgW+PEtGjyjgft68ypR2gMrQfZa/+gldXt88iCBDj
sx9UN/Hbah5IpXDVBYYuq6C+Q/zkyeSO2F4WsTkZtyVM/GrpAgjYoDMbtbL7nIG+
s4wAEYNf3UJhr2fsqvqrt+1sjlx3jtVgow3uJ7DBaqYUn7gUuQdMH+Rnkt76WcTW
892DLaphkJsV9BISIXPDcr8J8nO3x8M0tvkdlDxEcpHMs4Trm258uiq8sshWarL/
4xDdG9ee334G0E1xcXNQq6SsTO3zXaBMglqHEuAACtFWIbVE/G8iWdwzRCkmBaf4
ChXyFOVkM5GBMQ7TRHm4jRSRXP/VmZkIzYTONtAElwq2xXvhMpYR3nQUv+JYvl4q
PlVnL6YVYBkIN9ra7RnEEz4xcFUZfrE5bxVSpJO96amKXK3Wr2LYGnuwhOd/ifti
XzY/4ewiNLhKlfPYkBEMNZ4p973kFMOehSzOCjyYfIqmLnFrKC/WmoUlzlFzh6IP
2XuDz3MGKWbRze7bikv3tjhYPun6ea2Z0GAFqy3v3B9cQIFkbNkbhL9+SLj4X1kC
qM2Qpl0YH/nvpTdrskFwNgCsqcaS6TEsCjS+7ZpKTlyR9BFm3sx6H7/z3rFBoOK5
1aS9zlWlIoAiWltYX017/BaSlncIqBAqxfslfxibmrWXVLvVeahRV6MeANTA61/r
jenGPijeLhPbUVSZQUYHbTP14FBcT/LW+mNKYR2SKJuKxwmiRAs5mdueOGofs0Tq
w3cDUFfsYfSJogdvkxOU7KzKJIM/59Mkl3ruGCWkFkkNwBAAaJ0IvIwGQH2/MAvn
WW0vUvOldzR1s1GT9jA21/w0ydD0QQHEFwJOaEFeMzD8PsqZkWLn9ZRorh7MwpIP
x7zh3LEcotreyxXIW91zx2d3hjZHvEzqzR95vqZbdosvey8E6GHuz6CIOW4UcmAS
MT2nB57GMvGhfkQRJ8JWNj3DDjJOWrib2Bs4G8ieVYaxSL3vaCkasJ/81V0cnPCr
+GFs+jpkGwtt/elD+NGd1kS0kzg0EtmGRERELa1ZFtEimBCmCzyjAtnXE449/PSL
eDS2QjXqVJXBI2paYBsGbVinPI6/YRiBeYt9gXYSFiNjC6aDDcOBQjUd9mHQh6SK
HBbzlh1qOM3WSsOUYSKrZMZFLYg2p2h7NR0oIVnjqkTDOLBVb4FRchdU9j0PwP32
LXbLswBXbsYUS9CH8Lnyozqdc21ydSSNJpsvhi2NVGu3b1t18kgQnQPgzLRoNT1b
nJkfMu98RZ8fQQMEONM227pBtEZglUmo376sP1Nr0b0Dl8X/IUG0+6TtNLMmPNJe
`protect END_PROTECTED
