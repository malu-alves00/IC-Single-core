`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
696lOo9i2Fsm4l3XriHRZXwc0szYgUyJRK9oj0vkoocspl1JF1tShVcDfPj7Smzl
cDXaKGOWMeO9O8om+pt24WpRYLqhrGcZjEWir31RQLZh5SFXuZiq7pZuEb4BguEo
gML+eINT6Lt0IWK8uTMTsC+eAHEOPBvbqeUcRUByOMH42Sq1is/47NCDHcjCbDLr
cgXHayzB4UMlA2nXSA4uC7P51uTy/yo7FZhZXHsp2evXZ3qNkM6KnXCzI/ZfbJ2l
7RZUWpqzMHD6C47K57nr1DAjtMzd1VTsmx/L++Pwxsm+79NYR/HyGV8ehnK8I0uF
AG6kfVmVMctprJ5+vOnGa6BqUsf5A73OMXokIXX+xmSe5D/ARIKxL55Dm9hvkg99
Jfe1pDZCvSZnkCKWtpzWw/lTaHYQvTTDYZIcPYybZw28I+1EiIps5Xnde2eEvaxF
4yGBVOREr8IutTGWaXgXtvCu88AaWuG/HXMdL2eGKq+0W3U/Sn8wxGdocvj+MySF
q/nagjQx3BmvEvGwJjc/IHgR3gSTBTWB8PmvN6AoBcK2tAwrQmdATQv+ZhfJV972
sTWNh3JLFy6+DEY9NoxD2gAMQtdJnDINuSZXUy1nWKfrY2hlmeUdyspNJQzgzllk
G95LdfBjjwxShYO53NqfKATwPBJr1DF6BYjIzdv3TEzVGoVf+60yMA15mZSBfXHX
uGjQk92H24NRMjxMLZRUWIr9ds9nWbA6I2qEACtLmlaTQ1x3vFdGUP00ARtBVT5A
nZKekzPlmBf06uW+XY7RD8z9W4M06j/W7v5ChySAyQ/Ms888a79AlWj0PfLu46ZW
f/BECemaBBssV1LGdUvjTigjHsD8xXgu0pcqRDcrazoNujm9S8tRiWp3/37Ek1qF
pFMJkgiql/BtnQ8SWuc6llBxAU+aul8hGnCymWubE2OnBeccLXgyDiPg/I2wfiuq
Ucjh2EMakVeeYpVFi+rwiJ2mVY/LQxwanXM1vU1NRWfQRijlBdB0Rrpey0wy1km9
4T85QvupQg6zhiw+UGOp5mT5YWUFFWw8PSjcIdr9xkiAUNtu1MRqN4WA+jn9NkZ3
083vcWjB57fiH2RQ1vhk4OW+gYg19pAStXwywD+X2jSUl4jyYlVz2au/vWcp2a6A
8L7nsz50HHMNnmKIn0UKMKyaxa7WH7P/jQ81zFAYeAWrTIzUMhDJZIRKkQOX7P38
ZZeXEEcyW0tnaJNsbdjxPYMsdXkGl6ZwxpL7okoneBvZQdLoFyutxzUSQwn1K9gf
KZmxjavr0p9ZGMEhrTCy8JFnx34PjZcx6PyR/eUun8RIpa6qZRgxXixtwUgxU7Hh
9i2ove7uFtAZhRH+Jrizj+GI1vfC3cKC68Q4T152i53KnIxR+/zDqGUmMokI5nDO
G2Bo808rRRDUkTRmc5JwECX52LLAXNH5/biNJjzXfkp+Da/1dQ5JqCmoQRySehr5
j4zz38+U+8mgY9tIPSd5hKJJ9OeMosrTJ7IPYASUThjAlP1UbOAJtjS6dEnU1kj7
OkGBHQFE56y5xaGSSSHbyiViysaALfO/tklherz/aPIsbDg7hnb8d/ruGOQeq4tm
Mj8KRUBHWmrVbm5n4CW7r/j4U8dz9TN6Gf5wC++uPUmA7V5ikSeaCH2s+wynAEBQ
S8Dk9rCNp9hYU1C5gs0WnGpL7sOl+rE7O9D79pdCt0Uk+41glOzRiX5Zg/tH9WME
gZnsgngcN6jB9Zvxe05gAzXMZIHsG1hx/KVHIu+gJmBkUO4lmGbawM98tPkJElZR
TKpHZaFhxMPDDqqrmyq9sz02g0Zpjq+R4pT90nblt3I++jeOlkHOCrhYvf3jq/J6
JVFaI+D32nTLR4bwkM74C+J3vrZtJT39A0KKug7CfdIUYbW8kai0zSTTWzs/QyEo
xYHONaMSveDc1ol9MVDLd5vTfBPTj2FItfgCNKnKHH1rFqGEkRbsM47EDYqrFngZ
9DT0cbSK3RZvCCnpMSb8QHJBKMb9jv3uXdTzT6M5YHoGCmK5DjqQ7jpkT1GYNe9X
hugtEbZs/1Hj2fIB7/iUmCs2TGzhR/ix8HihkxrlskVVwPLpWV8tkW2+fL5Gohdw
Wa3uqbIacBvuaZksX9/0aIm5eMSH6pt4YnmuF8uhc2sP6ML9qovnjYyw3P57yqD/
loO7ITN8uaC1kPMyvumwM8ul5ZBpll8kNXtlmvT02VRNJvptb3b+s052sHVXVaxV
sVRpASZut9xj/MH3bniK/rQ89IsCSequGfcRG3KXRWrFD/D51OD4a3feT0239h0w
gtnBHo51E9rjvPhLlrcdpZXvjcPsZ8IvtWMCSeDOCJPfx0lhvnOQWeLMoh5XzYqP
325LIFQ0jw97dFACMLelA3tsLtdUH7/g9NBIJ9zP78UJMYJ04jjek+NDWrG07R0N
pYXXQ4ELe8UPqvotKY5sRIvRYquOPPt6uNiYxPGOwQvMzdNHdBrA6EE2sfUsUDfp
LAgQr//r3eGUmPIsOef0Ruupg10IorE7JEMIYTXabyaEF1mkUksea0QdV24nL4c0
ExrCh4bEbaP21hIr1zdXE5PYEXoTzBgezwmBWy1SdSvtVaqJJv1SbNsiGqVswssW
kxVa4TwCiO2iSyiH5OD7SFySEKioVb9Lt9g+phJiY7hT7rjSCWgA2+sevTdagySC
1c1s+1xVMW/diBQ4BngFWyikukL02Rc7xFd3qbVPgEaEPzsvo3jeA9wnZ93ma3wB
BrXYQr3S3wl2+I6JEXCrRwr92r3B9IHuMKb/4OSuOX7+WsAtsbs6SiLT95HSid+1
BVARPIuSgqd0sHKu4zIdUUMQkVdSnMtkHwllPhQjmKFktpDCMle505mR4nc3h3Rx
zpS1RKfyiQAvml8kRtic9FnL7daeLkKf33Q5jTtwai01hfn1//1KzL9YDIyBGRCV
PKdYNKPqBjObx3JRUhBVdSQaSsA7hTHBoarRhHahgfr6ZM0hvzfhOMmjsTxC6tHf
iAVd4pXMaTwfSK7THMH23PxwFca+JAKYgUNyGl98gYX2FkjpnEnwIjRGhDacp1Ut
v+CyrnPcCMI/tfOtOa/IpfWwN4VcOmtqkz7VUyjO8x+7nKqJXG+KDlT4W39wOE+Q
TjrlVD+dxXGOwi21sbPO47mgMlRKhZsgjRKzdtM5aL70HYl3XR/C+bDOsWAjCXrb
IWAzbWT8scb1Mmc2cSGYElAtRpIPmwGXQCrv6aOZlP6BtVCmMDIrL5aQm46Mappz
XIHQ+X5lttaQwqRxo61ErbKd75a+/Nk+iEG2PyGLaxMnY4afdFk8VGaH1ODaPMA3
e8j4mH2m5UtvoY0wyrz+6DwmRYcaGxp/Lxe5LUyzscRyfT1Cl7hFEuzJmhtjkzaT
UEH/jfEbt1Rd9Kjqv7k/CrG0AjPpUkZwcu6nclO5V6O2Fz9krKly7zw4iOuy/bnR
P8B8+nUF5/EVIauB2L3Xa2P3VxWmhhLFC6TPusFLoL++Daqik1jx5Acg3rcM8yni
Aet0PQrSf98J4MU23UtlMoGx8w4NvQw8WzMU6zAFyshua/VnLgFRAN0AtKykm2hj
ONzbEgfmXrIZ7I74bAUhq5Qw5jNVw8aqjl6cWCF2yH7ZxpG2r3wLLcgMFK1Nj3yB
u14cvUcogN29kfabfEGSOin4BQF/MBQ7pmULZChHp2hE9IkmAQVihVVvEVGUk2+k
NFxgYsf5dMpfAzh8JdyuwBc37zOPaqQONJ7KNCwz+COiJCxI5s2KyZeyT6jwjHBJ
Xt5Ad4nKfedq7A1pLRSFouDsd4rXfkQ2h+BxxGir62/aAdET/RUSyl2i/hnZxpZW
1z9X7CoSB3E4ssxs9+HcjqeDf0eS3jgbaz/OvHKDI6uq9bGkS+aiP/rFz1jpp5+y
Ara094lC+CQv3G3TiSU/6qYG+W/WvQHg3HLOdyG29Q5c8eAZE7A54sju9odph6qx
eGstyKjB3KeKJxNUs+ZgOiHIlmuWbFqakbWP3G3TAttCj3sd/uY67QJblgMZ+P0e
1rwFT72TFedBZp2edxJ+s0wL37lBNo4Ofb0vIws+jQqp1bIzHpwEfO7QBq9ESAA0
o66mURQIS7OlxYiQ9T+CYY7nyT5Pr+2t3iUDcdYuvMhyMXonZWG4Q1VqXroKe5rT
y8sUA+EE07/zPj8C//TwlU9UFEvx4FG4RAj9fomxLc5ci6A0N3PlxZaHOyv7cf8M
f2Qr3a9O70in6ZbgRS3PChnMF2QR5TVOcqvJ5SDRHOAm3o61m5K1j8RRhr2JW7Je
kWDs+ypbbL7spdgimJFG/SECWsUGWQZ7PCD5q71UBSu98/vyKXcP3VablpSXFKIf
kV4S3MufyA8vHkslSmMS9imOiD4Jq4OHKjkYs+FJVddmsJDu4+NtQ8QIcw9gsFWC
Euj0MEVR9cyhvsD9d/z4KeOxHUwg7cGxEdpCXXpJTAHlYzuBhbuWgRmceOuUvzmf
9e1iI5Oj3v85A7eMUSpSq0qJsE6yVPtodM4UY+iiQQMWm3/mcP4/g3hUUbSJRTcf
IYfElPYXzzaOM9b++nSqho9Amn6T4M/0UNCSUZV6CEjih/2c4tQTpI5Y+N3riQ2N
tLNLVt1vPQm/SYs9t8NJoDY0H9LBh9RoE/xCW1I9gVnZ2+SromweYj982bGU66x4
GV9VqtrSVRqvv4MCG0MzBfHsH9BPXJBz/idrQi7XwVN4fl6UZp+V3YqhA4Odlm3Q
InvRg0qkkLHj4hfqfjIGF4RVM5ZoGBlqWXXe7PlB3hfDj25k7xB5NL5F+eXV1ScV
TSD3suZkyNpGRDhMp0rJdfbO7IlLymlm/kU98gjyDCqtU+DyQs8I4/1zWjsF7tHe
jy4sT4JdUrtvRQtxQE95VRkJimHphwC3a91M90UmFO0J8PXYVtt+gq++GzwszhtJ
f/FormAC3o+b0y+McOUpcXU3CO0atQPjBVc8uwVzXBpzrt3jJ9Ow8KGPlieMe8lW
UlsCv01/QYILFTOQ7loUfwFgeFPwRq7zqYHSHG+dU4zRhLJnjPIxgFcaEyz/Xlr2
+Eby2rerGSiSIfQ2kCBD0vC5pMTXMBK44wTI6Y7+FATEJgrmT82wD3k8zDFWqHz6
S9m/R/uKDbbsWCvIAR7Q+M4gGE9F7+4vRh86cDCRDJ9tKxtKtBVm3rG0iE4PcbRH
bckLs/R8Hmc8VyYhS7Vw2z+p+zdf0/5FlF5HKvdjNz+CInmdemRj+hZwQqfdkKNg
acNqjdv3uIkCTKMAE/CvKkiP/mhibsuctPhQm80Y34EwgOPLVu5rA/KOz12fuf8O
5AgECgZXnVlkrYxjDRR9J2ck57S2uD523YHj0ishfYxEuUl4pbnGpKyxe3oaX/2r
axHrk/6YZWHCRRyZsy0rHysHDAFABC3s1AxGfqWtsJY0oXP05B8bO30L3P9Im5IB
mVIkmEb55ItGIK/HJ0mbm7PnCxTDLsSHxt1O+YXTqIPmnG5kuS9AoEuTsmKVWNs0
Fu4OikZcsEgM5dFntW0LKyKc5WwGLN7iZSzG86WnlKpAhjayQK4LBEkWRcnIde+k
3XQlpWJvo2W0jP2yLed5sOawCYGsIijr+fpZWW7SKjcdCj/6HNJXPDoyVSHLb4uD
CSiOrf5+OTNexTET8HXwZV3mKoptfK2sBdwSLUf6ucG20J2733GheOMa6s2JIUNM
t1YpvNxgjEwXXSLOj7WvBBOGEZ0fRs8iGL4BFq7vEA1pHBqgPDK59dA6y6epVkB+
wsR7BtYycOaaPTaV/Onlqruwa13C8fwoWhv03gGQBmLExSKhqitzT3ZRBfklXuy2
NHyCEx4EtOZWPvnp2fPwYlvLKPH8GMoJBI0tyjvsIpL8x0hMMRmJnv6RHLjs3aJp
or6+88DN3/qnTXRQCVGCPstyucNJZbyUTJDFl/XohkukdSZ8g1F5X8GL/nVZnh8J
nyFPoNZ1DcdyEH9eJU0u6bKooRntqhBYXZ/UkTZvCUoxmf1YTn0KbLueokfIChtQ
5MiD16okO2DxRq1EhNWAaDbtP+W9s5k+QXi4ykYKOK+QsWMmL1bbE8ME+XJy9DaX
NJFISXKlyo72d2oasFSbF3e2JdUqyqQ3z1FBqNm2Nn8JYuZQa4pP6vT/CX5Kemjt
1yxUDrxUI56kxs81G1S+uT48VqXqyjgSgcu56KA6Hpm2KgYhcHeyGF6r/xgllX6H
jOhn4GbCJ2+N+jp5M8d7qAUsUkNxLrYjNM0chFlGbUs+2FdY3YrGA+u+BYGgRrNB
v8fOewQDv+fmGubKOKBbV/az5LyMUf7llai4jGOEqyv6d5O2NQo9leiMf8yjBix+
CsWRuwcOA0fHnxC4PxLTg6AQSC8gghsr2RFluLPv/3rSzbs4tgH7EBU64Tn4f25j
jSnoRSjPy8HSEHfnVVBt9tXkxlie8v1/YvEumnNIkAAhqSLmpIPH7HcUik0w+ZcQ
XZygUyWY9GIox1p8/V83nnbmwhseMuWhhrPLIYS2jctCgcCzrUKPCPZefYufCmSy
47bOoo8wQRke07i8+Ice3MMfueeKFNVuO5KSy5OOxDEQ5/h+XSCYSeMdWL2MUpKu
eC0UKrFZvoJwzq0DBO6/U7SrHWbeQQoJkkRAhUYocwE+jjuRKDVmKPnYIKWQv8Ts
eu6kf3sNRbrDhOnf7cA33nAL9JVG7Q/RYcHR1rNB5wVkT10ijU5Xgt+AamFBK2aX
zXC09rloSbYmIFiHs6IFPyWa4ZXk+YQGmXecwHul5nGVy7VvYc3JCMquC7/sT9s+
eMd2utPdXIDqrf75g78woHZ0FFHoTRqel0jDoccpzXaMU4k1z4yA5uKFHwVGbRjn
djYFkwsSaQ4hFrUD1qnhpr9bOZ8qJ2KK1xn9tuL7M8UVOOD7B2lVLXGjflMLyZLy
8NDqNhbrXG9wFMmXfa6F/p4Y+KK9aBWrBIHBLVhbJhYvvMut2hjI7Kbn2QDOYVCH
iBgNY79U7d3wnNqgsKPaEYGNytX/eJppVRSXwDeKIR3s36oGNSLoNARVlYT3zvTt
50YX2VEoOAwBIjttTpwzhJjMNiv2NfgOAPTAPEQdAKN1vTJbORvWpPpqbn5vRY0/
VuslTeEAQRB16nfNYSYWa20zgj/Q/uXt9O8aqIs7DyiJ/lzYJdhK7wxfPsboxn32
lgAR//iqNdIPTMuqS+QZhuepo7nOkC7cwqTUKObzR0Ejy7shpE0brB4AFuQPaUj6
Oig7PDRO/l28BR9VS33iVGQxHa4Cw9dKIqPlCaDvTq6RoiHpQ0OneY/RN4f/oY6U
Ge3DZYneyAsH3r9GTF6CIZoqBndJgYpJAjCztppGEj3VnSBtbBqJKj6vUTmdXCCt
EE6XwpBMo/j6MFJgRvl+mn5wrx7lnMOo0+r8bGGeVHF4wOybSlddlqc4BGOX1q3t
zHXwPPIv0IutL1RX1sVYByM1T5Y7VWBfuzJfEUF5i3hLDY7Dm84XZabV6HKWyqbw
yCz2i+aPmyzdMfm63rYRVagRz1EuQxGnDxU/tG7BK7uLKcKduEvy1UCDzvjVoFLU
wH51d+B2UmHXK6GPEtszv1LDdwyR6li4OFH6OcuD5ahGG0UuvABLNTf2Ljd6B/W+
d/hS/IzGigS6OX8yTluW40lIKBElvkqC/MeNrQOF/3SNsR3/V/lLNrGjCddaaeI/
1TlPC4phWeCbtUtrRv29KuyxJ2HoH4XnpZT0KK0uN8n9XwJlx9CFnVsmXwyTnO+Q
aRjMdkJ6MHDW+PnY7636+NIRiBl4zGBBk6RXXtQLzROyi6EJILFfqDeCWzi6vXv7
MxdzBUknK4Z/9PkOWtFYh/bKBLU0RocB5PI7C3aERA4kRaUDZXbWl6AfCLOKuXS1
tYtnuMGX9H3Pq1YNMakKJ5n6oJW7R32SqPVTQATjYwPQC1qDDYegG8psEeEhxOMk
Fj/Drl4OMjvGgb4RZSm4f5U+lGG2julz0zGb8CR9+Fi2H/7EpuM/aIk9gB6uHeoQ
2OP4p4EbPSpwBrbN9KUqT4pJm5Ie2EU+Q+xJvAayjqa/zxhsgsMwzreAPnP3uGEk
T4/y+/7Vxrtj6S9ARyhu36v2HvxDAaG+/P5rhAVYm5He67cDRX/yZmDpLPRG8wAz
J4VOyF/oNOONnwDT8tpdDZ7Iu/AQmJhg4frHWftIHDlTWcLcA7jSnWM/NrecSYQW
oVieY6U4iRNfzeS33wYModBbTIhzj45mpnrxS3GADDbGsWY030CTuhY6GFlRL4GP
4alvqJmruT7eN/JYEbl3rgrUu8QcHQ2OGl+lXT3Ag5tTmLT+E7ULRgZsIDDa6war
O+4b0E62aXtQsT21x0v0UH5EFXX2iVVZY0O7SG84EEorld6TlDlZwCMEz1/eM4LC
EDy09jtqpsWhSG1RBkwCzw/JZD6/kk510uOS/b0dSROB8Ac53yyFJi7gsHZzmc8p
xNSHsOCjbYqi95Rpdwgnl/Ppx4tO6BAcvt46PUuo6YpYcju94pYgEdTcLTBlgtjA
QNjYDd96BIhsIp4sRh82aPL4mbVntnhnbwcF/0uRKjzwNPqnmTJxpyT98rNrYdYs
wELHrXDqOtQplPJpgp4fR9V8jBn0p4WNTKnszi5gubdFhBU6sBL+fPvkzF/VRGgz
kOcnr2jHkQPkJ2WjN/a6XD0TgMvHVDNEsZlZ83+W4l2i3ylzLUFNeBeV4w3+rrDL
aY4oe/JClFGSgALRERLZVNiLDFvn67gEWRkLWoST2jfjDsKik8ZO4ZOLhTcGIZPt
aKZdWqgXjeZlFYg6+VDWgsrJUKOSLsvCfKCbXUeXNpKWt009xxbMSIfg5Vuff2Ps
iP+kojpHznGWNNVa9rNff/+D3l689Zc5uR/esu8Uo99zg1jspu0b83IRdSboWtgW
ou5XMoO+oTyMFbZ3P744ccj7TuvvG9Pg6QmEANB2SD33+B9HAoqVvoR1NsqkvWqH
/4kr09hKjNQSKJdzv1ZGKB2/85IxvZkPseehvFHAYLRxTVn4oPDFYwU6rbn6JNH8
pq33dO0sPjQNVJKfwcc2bONiiwkK8B+YjmAZWRVzr4X/6CPkYvQlG/UOhoJR8pHh
JSs+xO4AisAIpAeQIfB/GelWkbUVIKcJ4dTMhf9ZmXR93rT7UaoqpC4a4Tsu7fQq
ao0tmqAl+HENGYnQbCxA+CI955zdERl11ZZBuMz0QAnspj9wsOPwWsDPeMUiKamO
tj5vJK/KmZHI9+VeBpQPCnEnWF48+Pf13zTw7mMz6632bB3x8wNdUdHVsSlPApJe
HVfjpohJJQyqvBn6mDtys8ljlohkNabsMYV2OwHEqaIz5YXhIk77QZhhoCx0IFmd
6yUA6zJdwfeAtJKdHUQD5J//HPElRY4kCAuXHsMg07AYqBefeczKU1YI36vtuClQ
WJktA4bXG8oGdLKtO8fE0n2an494mmef64KjEGaiy4sfgVOF+CBQ8Yy3UzL/UalJ
zgDokDdQ57Z9Fdaym2WmGFnoovx5h+li2mWRPabQPCP8b/MMVPL7eNjHLPGSeLbR
iLr8HWX6X5Kxv2ZmHK++/5pmu4ZMhrr9tySjwCkqLRipgrQ0voco1kVjhZwtbaEf
ARbjTVz7zzUVrLzSyIFwwIgsgNRY0ZQfircj5rXw2FXoKsYsS1PDGbzYwZk9ULxa
vwPHGD8nf2g3Wkh0pwvLVUAFSbMi2dKwK3n/MY88I8BmbZWTlhhW/gUDiu8IJx03
thkwDDX/vR1NFSCK+glB95WKWIJJueyen6IVBkISOh1QfR+LNfmkI0uco3OhBh6m
4FcMeGkyV7lX13k7PoJpsfoUwBCljZ6KzySyRJ/8owNDG7U9O3BKVB8LVAS+77Wp
INJu42P+7ZcR8sXjKfiDCqRUDlecB1MblWkHInPro12DcmJ0cEPI8ksPJ8vq0jti
tTpHlDJ0EIMNHgV9GpVdOrmCENoJV6PcvSTTOB7jO/QXs1SBe469NYVh29COuB9o
8Wb6570TkO8wvfs70/05abZca8pwm21sfU9zSIqVhQQ81ryQ35CPKGSqE26TGhkX
PSj6rQV0a32CIR0gQlls0r+gUlln2iqAz0JOyOYvFlbGIVEsWdfgWtMx6sAgP9mL
8k1EWLpZ4OhJWE1xSO4jclStjAgbwu3mFfIQ24o2NCERvr3fB5sV4w+dLcxqb2gH
aoYvmKnACZ56BZLIBadj678AyqvmciXPeXb9HvQsIKt/TEMQULMMMQC5BuiPjjvN
FtzG6vkUEymqzjEIcdwZ68hW/zNnB/wgIDd1uOmfXzKpp6DDoGgYxLEvNSMe214K
lAj4Iz7GWO+0CbuXfCyYhE9CO8nrmeeWVX9068P7cC4OaA3yr6XAok9LeKjMhZPv
vakNqiVQ0oDcKLXwlRhgWU5BwhagVHPTsoHxXWHXIXUEG0r4JXtgu/pHyyiAYIDQ
OEUBV5HgQT3escNfUVn/YnGJTgH4nzAnq0eaaLHuRVw3pqQoVMRG2ceXUmjvXCLo
rZkqFNjeXmlDdn8Sxz/5ynAxBCVtStVHLqgBZWeAAfUQTQ6jCWbL/7OpMBqguN5g
XqZPUGYLVhlao97VjAfB7KDk6GKgWF/AQB3Tm7HMJ6466VwfueZ4a+LHt4pd3SD4
/2F91xTxIzFSBmffwkayt4OaRe9GFVbOSilfvvV3J/9625+oKiNLN3tnp9UJnM3u
T9cpi3O9tcOGuR2VKVE+AU0IOfpX2yWWfQb407MBCmO6PIMWOjjyM0DTivXrq8hN
yp2OIXt470bn+CHqmWqbbMlaS+xscVweJjC+dbOxzukP/ImhoUaYMOAP7huVGmfk
m+atPaWTV6mEtaF++EMrOK49ASG3MfaebKmHk4om3rIiJIVDfZC27LPKDdkzahUa
oqqkYpoOxAys0qTbrRMDp4En84LUK39fbpsLViRUqu/Gnp+loBywO38L4mL4dWrX
h5oaBU5ZB7kNvkJ/tj3QyahfSdL0w75dtnYhwY+a9MYJ4nwatgxeXkX2CPIYvLB4
IzVnzHFn6MjFQQENb49ePcyg+y6ebWcdM9TDRbaFLkbUfRI60pJkf57eoRbOQzt+
qn1aGK5mT5q5Qi1LaXqApKVFYPRXcPTA0TH3zR3JuFmTri8xnrFXmOfw/Abs2sOA
g5X/wqh80HGEH0hqEplR2S4mnv853IkKJHaajGI23VFA5L94X9yaFBhWzFpd0+Vq
b9gd3mpOWfxRzfvMI7/O2Fww4/g1oo09jTitsowayalNNv+4VpaJM94Ax4GTRv72
MkmGP4oJIhLDXXHmXRzVNr/P0PwxrDGDc5FJy46OrNIfBx2gC4ke+z6t5GKNbl+b
vBkF+op2UJDmIVN1INaAXnOPaL9SYDpmnWJJn/bOQ7+ZHptCZLBXFdw354RX6gsK
3RRDzsto0choWZ/iaG1QswkLh9p2RAufStyFqQ0oeVZyo4RoJpvPN3xf0IcVrZ5d
G7bAdWGhjeepjbStoxboWdVimAAjClmxiBGxYo0a+4IH9OQh9cYLB4E9xN2OXRif
Rhpt/HxESs+YjiziqVRY7ZkCgNU1mwecAr331J7yvNApl9+fWSmbpurfoJz7qP3m
CAJ6/ZwEKm1Mwm+7wgFtXIVfEp4B4Gws8uognU6CPY6x8XJ/OLrbWjoHQHeX37g+
j7QJHciaN5OjTl/FHjLCD7YZRKpOWosv7zJQ0R6ngblKfvHvwXQPX70CNViaf5pz
sckQpp7WHVz7LfCsaAaYOb8V/rOZtPjNY/+y0lOdvhRrbGZQAv98W9ipWN1Ye99t
hu5KKtKFUe/D3n/gxk67vqWN8SbX838S3LhhfQKfkeRfj+U4xlWccsVJuX01Ys7L
R4FCoMy66n+o/ScKZI42NF3HP8HiqcjxfvLCGDGdljw9Tn4N+AnBxjPURJabmvsh
BK7ahpdXsiW/MfRsNe4lG0ldA5jWfekh5HKCuMzYDeh8xMqgacrBp1yXZA9WdvSt
RMTJ165E4GQSxSGqRlRIm9Qem+l9FWLDZXHywfbWdQOS4mq7Ra96bwGLako4U+ev
2zIPsAeiGnMnoTuZ/FQ0nDWJQToT0YQkoxuya4grt20M9HWpGSZ6OMlbOZsJrne1
XQ75CO54/V2p1cZBEAb8BYd9DxSpZyen+IUWzqagcMVlrKp2U9WiTGbo5cOYRsBS
zD380qlWvVpH+a4Ok7Lx9hDStyvAOWZ++T+61Z3+2uUcyPehWWplS42WlgpXh0eE
gEzURMqDg3pDX80U9f7GRQJwtpeR8f0jMWbZzzNLXbvq3WUzV7oV0CbvglEalLXW
R4yyZtZPuQXQvRtVomFDQeFV7jK344qgWR+OLRQ0GquWeq2yd3uWVYR53i38WrMs
tAS+QFs2Ae4hV5dF60CyAr/8P/+2iPf3bmtRZQXwMhjAYol7Z3Qg+6+dslEAnvW/
Okut5tOoaGut6b9mSR4bs6B48RGMES6t5/A3p/SmKJAbk9KNRSTJ3guP/hwVReU8
qec2F0u1cZOCXM5hL2FawiEeev5pjQkyJvapbcqTkL6yv5UVtsi6ZxWVxpJage/r
FgYj6oagdzV68uuBHGDotsg+fnJ6QVTv6FiODBInpWiklB9Cw+dqKHcEQaUUr1TQ
QMsI5UiZBTiux/wYkXhYpcT8CrUz/8UjhT3fgQ9J+G32zzWm6FsMJNrPcKPuYvm6
6CRa0exwlzlYRRtVa2fnW2i3s8vGAqY9vLj7k8heBHuYmhsAHE9yR20ISOS4ozXm
xhjGsBCe8PmbMlIp2ZCq1OaqLqkou2de+l8vxLPzFcyMK+v2eYHXbJmQg/uofQpy
Waf67navAWQcNzTx+AnqCJzJX7vFMEN+NJ6nvdgagH/i2ojI/nkmxGIAHplAxrn9
lG2OlojR98iTX8IIAMEkUeByP0HlKzDL8nFQFrvx/7QIHkG2jo8S7XABI7W+T3wv
8wb3TVx8OaDIUODcKwVSY6ADvaIEaJBRJ8a08fuZfI1KlXkVTdDNNht07m7aFmBA
sfhp0Jj7ARSXPl6Idctu9zHaDUXx68fwPPzGq2iTD2dLJYBSUicsqLsPTcT5xLVB
uGQGYgqOiHaEqw/QYdHMXqY+fUSRWjwmmtGFhpyUfMU48y0U6OE8u6QCeTBfkaw+
9F4fom7JMKkjIiP9bgwrcg7xRoahMzziDnL4IeeuVc6j87dDuviLp9rkUnkYzlw4
7zI6uAdi3x9IRJRA0GsPbtgJNxlr6s/v89u+PYls7Q/9Pyx5ic72OUkFQRafKQjS
LVd2yKOQRxmw5xGjWLYvDkjrVA4XkzG3u89h4dHxgKS24k2Na8ZPEEOzW9ooysoT
XjIrmG/j0uUZE1OzVkLkGbDjwpBqGDZd4uoYmkulXNVDtg/bi3nBZ/d11f2Ym5cH
6qKjoJgJ4KnVkxkW9JiWPVb+ccRcMfNLCfApasdOI9CrDAgqcwO4CzGneFQGOkj4
q4QV+fAhmgW8HD5PTgxAKB48PKOO/zmVIJ0HYhkB7HU0rmj8O58ljUSNc+t+JAVx
pKy7M9xf4OBQtmRF3RT2ShKMTaeV9jCd0qTniri0Kmw0pbeQIsf5/3hgMmEqGeSr
YEnYULfN0w4eAy/FTVhb2r1FjwoIVi1RORMOJzK3q6uVMOKdJykHfrXVwHADkJbW
njQ9aVh+4B0ULA2CUFCp6KLfEpioHlAGn00VGsW0wwJC0T1XQt5Fu5FoTbjRGa0+
wcsSvjUYmehvUvoaTdra9LhOC2gEld1WkOndLcEAxjHrKCxN45t5NugnJSqTHrno
J4M2knfiiKOeLFDUudhrrfGpDVo4lDrB8paT3a6GlFYq4hb27vm56vENjXSCvMtR
Z0aOFU4opbX4NBO5rkAmKQ==
`protect END_PROTECTED
