`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
a8tOD6pYhhDjh23ReSy43/ajBzWVyMz+19NHN8omr+rCXoNkWw8AopbzaUyvKVm/
o7e2XAhxNk4nH5BFo4qf13xz6xqR6xoPLVdp3vczbYDpOX3rg6/R/ZWAllguEDkv
mBTImxG26w87jVz7FYlMWlGdI8InE+rMm+JkglI0mmnvdeqq2P9DcZ7xZRpJMU6y
HuLvQ/d0IlReySFOD6bMjhOVwKmrPbPngU6j1U1FOVGGIA2dnSBOt33RnEZcqMoL
Alr0toBFJz2/b1fy3q9kSeL/qelN59jpnqq4F/iCy8tZzFpJ/i5B3H2N63qx2KEC
Y6+SsJ8jfTic35yY0Atw0hfij2P9/BB8QY12VcewPq/ABY+C/QMjopTnb2SwRF11
Z9XBc/ywoacOXfltoO94ag==
`protect END_PROTECTED
