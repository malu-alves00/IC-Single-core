`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
S/AZPRCNNn19Lt37DLd95jbUN/hinR36ZkWCvMVRuAHY3fDJFO/6wyIU7fMhboSK
IXjOlpq+ZebZEnv5+o0Y0fUE9/ErTEehykOPMiMhEIv/WDHc5UDfRLF+9hHqRIoy
SgtsX+coRh4AsesE4qSVCdL+F2Djq5zvXZn8j1UUO/oXzcGzzEZ6pdPW3ALUdNVX
EduAZ90GCEakGcH1Y/7d0s7FIVzKpApa2f+NixMoLCbc3yy78AYAs0zU9ZYOh/Q8
hbek57TKNjI7agFmlZsOv6eh2eacXE7EJNXaL08UPllDAv++iECFn7ovjtybiLj6
j53wsNxUzFn3/ss/vzv85yRiSom1u9IXlGwagmhkV4T+vDUT4IzdSawg89KDMbj+
yqMSuq3pjp4zKOA4E2OyYGIwGWl83sW1i+dZ0yGvbiDXc7+1tF0d25fFRf0ZxqPC
XjGGhXOo4pleqniOiOQFK66QGafG4OJk0U/4WTujIKsf6h8hfDSlOhkHMdpP6h7P
/Yb1ViugJN5jPxfvxqBvVo/hnYT2GKZU7LOzSHN+0FTxuiWTwN//8qV3ZaFCGJ5i
hxvMhvcAHANcBw0zpM6kuKdcHciNPynU2KjNEX7AK3mUVrvdvZADEPy3wAFFAfAo
mdtLE9pAdlf7LuuasP9R2WFbvTxRLUjaEZTXsXNrWhOJ15pM0+L9xVTjcCafAkJY
YCFy/voajgY7nAEGa+9dhJbtInM/MCh04l1d1dZ2T/tjJp1XHg1ugvyF7uZT1fHT
C38y4eD5RTQ5niQDT1jfN2TG4T1gFXfuEZa/1a2VYs2wc/+avPX8EhymyQOrp9FV
v5tM3LunBRwspD3uNwO3q1wLGlHVgBw5H79qFMEF9PCStfaCnKsWOSZ5bwSp1dUV
W6aNOuRh9AvU3bmEVXFT1gJtZh5tUVwJ96teBvU/jEYuFy4LvHQpEBx5IKfpySEO
`protect END_PROTECTED
