`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xSNaI7utSVNDnaHagsN5w7yRXvBOdyhuXzajNFV35uZqZVK7cDnRgF5s6DhPkTip
w2rc4LvuUv8A1IwMW3e4SS1mazRdV1OBclztMV764I7gbn72laV/7YsgdPAI1VGw
EtYQpzHnkgOpbw/5gx9UULWhjr0zFFGH+uKJaU1r2H8XhZltegmeI/RzlItU4/5d
8h7Cr76fHnA5v9BVanYVZD3mnfVQycdu09cAV3DrFrZIS3vBHot6bMy0XNRaOToS
d2RoZepGawYS7VtGT9x4Rud85o3ScVxo+V8ZH11iX0rAy9lG+7xbq0ZYeyAG14NY
NZ+uJOxbwuQyJH7DJOtXdxuCz9kSiDhyP3RPXJif5fxCMEXNizfMUfR4RJlWd5Sd
5WLFI23SCLjnkxtGqZbVqanG+RIu/zksRb989uW/iBClPkYO1eac4dTd0yJjFz7Q
RvP8At4idV6xHOcuIGOxLbf6xKBdMHeJhMXDzTcq4L7KbKVzmNKwKECx8vgcnGFK
wjnWwOZFmfYi+pA74DoEar0kFSLc5u6+inX7PImZ2Zxdoc5tgabuz5oQhf4lGENg
lOjlLVAez7HaXpzGJVI36HhQRA6od12zhzhXduc1gHSVReBI5LXSE/psnfKpo0k8
8GLhTqPaGTEhD2Y/+qocxFewaAQKLBi6VlxqNWDOUr4Rtjvxz7BKxlJFXBG4H6Zq
z9tGi071MbxwsNL31IeKetlnBiKCuv/mTKv9Fg5DOrjP1PKvXYMatIn6SPGCPpW5
cmNBOTFO2+JznJ3oHb0Ktd4e52HlvOHEFzoaSMwZPGNoK29hHkVMVi2E2bJaf03v
7ApbSXdxay2dQCHeP1Hb9g4/Mj9iFOJhw0wrvhdzfXAphgmGP9KNZdiSGGtXa8AU
3VM8sMtPN33Op6lxPQkLiLT63Y4Ql2MhRA6Wlsi0rDsCS/73gvJTROuLC6heK6xi
XLwvcHtMjpAPoxWOLsuLT1rd0YiRm5p2ANnn3t4ONFLCiDn1/oo2YQnIdBbva1ag
p2CQYIi/COJJ/w/OwHkTOx8QZSSJ9JQ+fo+voUaOZnI1f8a/u7gX9ClDIv2ognuC
+c2qNwkAfeLGIC6mcvRWZ3D7wARnQlU4YDNBTihIBnfsXIMSQ2NXY/dGWpni0408
Dw0BN2Save5JgZHYWP83ArS1HGv/y0wcrkPEH+QpwNQwfhKt3dcQzkNX9CJC2abN
ZA760gWmd46J8AXEG+wGwiARNg1I7kCIdevZU7XHd279mqivWHH7yPooencooSo0
O8cuSxKTnn/JEwdejqBJbhTkmw5ReXbp/mN7ubvWX/E=
`protect END_PROTECTED
