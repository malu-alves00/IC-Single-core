`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Kui4Q/ND3ir1EU+yKRticbj+Hs8bUmVwzl1Q+Ya4V7YeAqFUkOrw4844aJ5MEfFh
uqEZXKjDKeo/tua8nuuQab/o/9l3e/WZq5EItECXpWPtbVoTDGcI6VaXVdw8Ya48
Yf4Bc6MZcfJ7IGdYFMr1cxIptzuafJrJdiYvHgMOXMWgEgCGSa/boWyXoeTwAZSo
hFbgkpvj0S4G7Up2mBwkaTmyZ5ZEJfULqMkgODgNDlJ6y1yhaA0KXXcrvx5CgX01
bcCXHYx9wMLhZBPRWEdS8x8RiGlrG2ruKhdas/Eg5ix2xv3IpTLGkTRCvzY2mkgU
OS/116+cdeHym0IQwr+GrwCaCEkxqfy8nWMwmskmCp/O3Y0x3K1cYoJPB+uA4TMm
bV+Z4V/gmMDwKVeueDxJZ7uI1+BLCp385GhXSZQjjqiyDFHF+Rd4O5K4GDcaytn9
UOBtlmA61LiIEnAZvNkj9j6Cp6gIejeXUlrePe7R9Hz2KfYybMHXY+ZdKU4KCMFW
PWEVLi2QyMrl0T8CnyUC01xbkcE2Ls+AFBBMCOa0CdIGxHlJbPP18ipXXL+eno1D
SG+P/6bQrepMJjBYTsYdwvpbbnMBV/MdUOAz1O3hqaq0bDm7I/MgLwKAUE9Yq0tS
o+zXsN0+bPNUVwi7SG3394rnPIoa14LeLHL0bNLFxDb9qIxEmbh3KEZxBDudqYEB
XVP5JatWJGEAHZiHZ6jvgSgUkCUjGwX9WOtjLVOvV6USP+njkw04H/C6SPmv1aMy
Jk9xK091pGSEPtSyPQNzqri+l96FcwuAZl6cxZok3gzpl4N5c6ElQMzSpffAkSJ5
svn1SlLxeggAv4LOUkq/VTuytE+bISDAm46jX6b11r29huL/uZehhv0uIxmReF+q
oGVKR8nTctpWbte9+p7/01BEqoId2+dWbkVhXaol05shliM9mDApMlLoeHruJP9I
8od8S5MJ9GlX0bRfyDyYWhnCSZ9bSY1qvb+kSG7FDKj5gIebkN/Qz0y04Osoqo0I
iKi+9FWtTuJnn4sr8dIkbp7FtSHKGB4BeMUNH+xqod2OYVU4rYAa1XtEx7bGRodS
nnaLll01qXy+IhBV8AQtHsWGyffnzWMRU/6aSudRL/uX388JO5hVvI2tUsQfAZzm
gn5HRb5aoUYwGN6lfJY0Z2xBKWfcHbHQFlEFL/KfELLuwqx8qYbUAiYfoET2tEbj
RVmGZdcXMqLna3KFSBwuFaldUlrj4XgW+a7RdpXqKcK0OdbXJLt5/OGN0EvdQ7qb
s3a/aHAhHvk0GF3+QCNIMdRPwb9nIJAu+1aeFl5+LsWOPc76FrMQO92fA6RUPMVs
kL25vERIJcIEkruQ6UUzEDKvZ8h5Y3SvFRotyhVsY7LPIUsT0ePytokIl4Y4zjig
wIuZQEGALGLQsMMmEfLOeMO1Z7Qk1MXZzlqlIZJFCbwo4Sfrg9g0n6C+/hQPlQoj
QLqFQQxaiINZBo8MrlVj8xVEnUt7PNPFBHAZ8B73T6t50yznflKbpOIQZEHSmm8c
nssX/xueXxHaYGC/vqT+0w==
`protect END_PROTECTED
