`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ORFLXcoNTP/LBO7delbgwGwHDjjsrAuPUtg91NT3bUirLQlWFiwLf6/mjIcKUG4L
2UcpqcZ0Ya2iZlYg3V/VcsA/RLH9wHc2jpTnjgh0FuagO5zEGk4mePpvU3XrPue4
8TIog8l/Q6TLMrX0Kg3E+G3QlYUNgjugjSfV0AbXI37L5uIUhw3hI41daR/1j5tM
mC/IrgnVQcjRL+CV746L9/aO+I9nnH5F2k1gy6wO/04Tsbo8mv00tVdHJX7/nWBk
WxeC8xMAvt7+SB4KaTxdTQVGwOJhYhNRrrnMskP8FocYRsAumn+kuXYtlDpAp5OF
wiAFqbAiF1rULjoRqc0PYdNaMR3THujj3uHH3DYFV4nA2Q2dHqF9Vd5fm/XzkajZ
U7VOV5Sp9cRkzWg+3emGkG0TYkxO+d0fCyH7S1eOCR335iUlXHK3POK9avxjL3Se
FQH0vhGa03xsgbV5OeEwWHuRhr6jU36oO9xzA4OfHdU=
`protect END_PROTECTED
