`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
e6OI6vDCHpvxuEfol+jH11eWDt/jGJ0SXUq1HOqWhSbphsA9KfHbhlgU602ujh7S
fBNpYZEmLPJHukT6mEaE40Kk7oPX0tNSvgg9271U6ZjvExFGMTGxBIDi3VxbR8yV
+S615SnrXXc064gIImnbx+pnTCDYwFBPQxWM3jTWDnBOyze/Myc9WFz5Uj3dmdT+
HdPQv3pzz9WSu27UdFxvxS1EqYM9TZfS8YxJO8wrS/HvamqlJ5BSWCWTimOp0iad
1oaz5VOEqKogJXw0xz4MT+JWiGFDx09ZZpHv4IbgWuPLFYTxuOXn9Z4B3+jXSmZq
OCAC4C46HSpgfn1KuamGuRmEIhtzZEWq2z3Zp4FAdCueZnPCfM6savh9JcTTqgK6
wwnKUsJCfb+8oYdk2zvuRdNmV4R7EwjD2Cirui93C7zW6EWhuUK9w3t1ZCiaLABa
oSKn6wkHo5b3c75Q/6MsGrCvPwANI//M/3nPMm7wnS89AZre+8LTChDGT1/Kha7R
pHaAI5VShfHuxIXhuSooSGMEFJYBUG78qT8+BubeHp8PgMaM+b3RKpLNRTpsdlsw
6pQl7iO9a4ND8CZBSsVX5/yiK/tqxyNKwEtWSvLYD2q54Tn5orVRSppxALmMhC4w
oa/l+lfNEkLLKZRUqFTfQUXw/7hyvUxhzEAVspp78lIs2x94Bwk2433xLgGmcbpG
yZsHQwgMAcAepVWA/yKeuxXeNhaHFRf9EwkPwjT7XT1eU9us8nNoDr5aukojShby
3HY94i55Sn3wRl+PI0SM56Ni+9q1geKx6J4E3z2RDkaokmzCtH1y8Ucda9XAtsCL
dg5fSfamyAv3VlATRNjgkPhhPgs4dRQLAPRisf4/yxcF6lFTSi6QhOWbdv7lnxMq
+oZMJYsMNOWQYxWsCmgmh4YaBm42VtYJ5whykso7+es9OEMr52cQj6oTY8aJZ6uf
ql1mCr86xoKI8Ecjsixtp/3Ns+FUckkL7fu+GPSBI/PLBVv2SPe66iBaN4vNr5V1
/gwXDAmw6XBITaYpqAZCg4GgjIl9BAZDK7qwIiUJo1VCc1WqauhQmwRFpGyo8TSZ
aouZarDWgLjE2PWe9Zk0Mze559VBnYjoghXJzkVsM42O4qfY5IUhqHKEvpFXPxQI
Ya/GpnyAI2c9MA1gM/gDhXfyT0rFSBE3A4i8+gSDPcFzdUx8toQjkwcxtsuFZaYZ
C0Zj4aq6poO0nPXDZDC8MysBbPz7l2TfQwYhv5v6WQZpxSsLsYdxtiWNJadQmLSs
hYjqw9NXC6UvizvrdLOwvdGD6zkI/MjeyUoHxb8m4vxuahq3VDr9f2faTBODqund
a7CnlSaWoKVtzeB6uiibVF0+TnkKA23CcjyP9+6Zw0nEj6AjSCO6U/WImAiK6MCm
tR+p5vrAp9eR+Tpt5I9FstlWK2IzczeYJfY6H6iitLTt6Ap3IOeikcx0IxdD+dzE
8vT7likrDOsGww+CPW6jbBwGOGneP2DD+t3aWAaFtPM04wNMIc7I43L609mreCCI
h0VyHYFH5Bp2zLcCbPyMfeY5EpNlWOvCTtmCJ3zNTrXx8LB4uMluopfM0dV/lL7o
op7H0+Jo5dLh12LZ57y/QociH+mO/gFfm2+K4XHRj7obWly3r+ldh20MhoMgZJ7r
BN8YqHGaXh1RgUOzGyqc6j8KdR8tjev26hY2aGfG2Bv9eDS+GZncl5YOdLtFkNLm
cxdwH+CY+Ev7QOSbnx9aGrJo67z5T0CbEHF6f0c3A8u1nYKMJdDkgcT4/7VDVfrn
6JSV/3po9b9u2WEDhuxSRb5GK4Du5NJD0Nsx9YAXP5wOHmOUA6z56OWNpFWcKzRp
nD7ra+lPfnLxPtUkh0R4znbLqmh8R1mTD1FpCJ1bmdsmq9n39N2P/obFI2ixCxlW
TPQVqmD3d7kf/9UW0n9BDSsgubo4ZcHcUWtR8RjddU/kTC6lFNXQ+2hhNDvCroxG
jGVdjfvZEzveMPd2Mguqy4VOIVajlN0xarAxrUu57zwkcinHXjZTVpIF/d+s7hTG
E4/ebbT31q+S2/wvE2XieBbv7SveYvFmodsiyO0zHtJOEYjyOUqoB1la0sI2wMw4
Q+58wY3yOnrI5Fv54aMIZyilW+NsPKPSZBFrGeqIy3GaFWWbWBYOn6Pxz6KNqLHR
VjEdU7ANv8a57drvF1xysnDx+qxhYywHt+vLTGFz2qnD/IxwJRB2/ECrZAeXNDGD
cIf1UD2hz+h0TqYIJCq8krItoIP9bJdbG/PTkItxvnSGux3CH4PfDswHakezxH5x
PS0OAnEEQl7qNkC+vlrWsLhBPay1TcQ+WN9sYqSBrASK1bLW5Oo5iXW/jk/jEfTQ
eG044TsIM8hITjumGzWsEOXcnu6ufvdOo26qVSvdCkCOLjROtVnMdIuuKMP9US3R
9Km+PMI8nVMo/91al4FYfR2ldPC/67l/CO6pE3YW4LSBwuCQTySX7fSSa8iEkOQ3
4eaBsQbvuYmEA584scsY1aF1tVqHI/KdkNYPCz7qtORJs7uZrKbadKRtO70Ok9JW
uLXXOxMlx2mu9o4Cmwz74h8Ou+hP0CJcCelBYrjinv44fagfwcoHuuL4ra4i1NZi
TuYbbhYeobLo6zx5m33LTycileIviWZO0qrfnTcxziy1E1HR1dyk9olJhXoI+8Np
wSlAl4EwsUtvCLMx1BRGpgQ51I7IZe1Xqni5RvgyAMPch/N8YA8QSbo/vm3kG8vk
uhokZ1xze4AH3J4ySslAYps8DrjG4o8wEUsdIktMLpQ++wXdl8zL57uDzD2Lj1dE
rP5x53wOA4kH1ZZ4gip1NwN9R/J2digUF1p2zVeYwQOJQq3YKMhT/JL1Wq3VGW0k
rHR20M6fVBHxsDgggJF7akssxYkjus7xccwjw4ddpz1eku2vMnY/ML8kdcEMbPhh
Z9zOBWmH5kHxK7vmj+Dydt8yHzMgcxZkmdKfbIRBaleadKhLs3ENy1FTRkjCoLle
8wMwex9zl4LB+K6uW0BGLFC5ucC+kOjdDJAN1ieEvJ4WwuuGQGmMKhdIu1Vg8xzR
GgibGc6Li1GwLRI2jLuVQvt7e5ANuaAQkVUtridghWNMys0gmEKnl5uITeXzLhUe
3eNYLHS9xZLRpJTKRkTWC+H7dnEtzdMZsVHsWvEt9xyWU6zvDnHmtO9WTW2Jwnht
5BGhqDl272rgTBOTm2q8qMy1e3xZuT4+9j+Py6ubCqvgxDTjHOUzjhSrV+EEdQlG
GXtF+iwBYMg0zYpxqDWxfBB6GWqfIJL/k8UP6HPpBbPgAjUQxXsd7v3851yyKMVM
DITR1yZ1cFfdTOV7Hr8sP4CDF6fyjKljjApQSw2npt/meeMtoI9C76lrN8xPDkmV
waS3WGryabX8WOMcen+t67ZxdiR4NqPcPufhIBdEbqmGkRwZ9vbe+QxMk7/ct8Xt
3r908PlA0BSAo0/4hrVA0Jhmdt+DL++PFItbDzuj/4UufBL2QFyHsL+RchteJZAH
u7oBOLI9/PWCf+u7IWevhOd+785OVYkhFtqGg8ahMegMK3IYLF9nhzg/TvOAbGuU
Xm7aYH1iuvbCxSJQFqKGFAsWVFODQDU83KeAnoOU7K54dPz/Co9DESQYl2o+bS/m
dfe8nKQqyGUMJxqFbj4KLs+Xv+tjTRIS1jRbWt3Hb2okVP58gbC9UQPgRDJD96yB
HP+JuyAfPTpvs9X67uC6d2lNpU4OMYq58ctAMGiiPNX+wLO/FoenfVxr/WkbIaqV
/pSGD4F58ZN/xE4n4xYqZX5I6PkNdZO0UiAbcpFyOe5ngax+huCJous/MaOaqchh
UBGf1IDej8c+eQV/g/Zn9BAkgxluSO7DmJWpALoV16gsnWDYMS1/MHtdD1jrgZQc
nyjSjx4fvAmLDaufuDd1zIrjvayAHRdWGPBmgGTO/2VI7foQfNexJESkg4v3y8Sz
W8+QmOgC9mhIu+DUjlSb4QzuInxqpzTmmvzFd+R0o9wISsr3OZIsOjXaYf1W86wA
lDmBSXd8QHi2LqJM5q8gxhNI38VAe4jXiiT0Or6xVGNNl1Kzs+YhGglAToY5FffW
rjWVhoKlT7a7ssxe4iw9ctILXVQcRhhmnr1UmnJP0Egdihael0RpAi3avZs6dEpp
xBsJtwjk3v5a2uHTN+d/bgP1gn4gIviQp0gaWX0G2Mjl0fF1MKXI1e3E9tiS4kDF
eqAJ77n4q4n6e/nhn4l1KRgLeWbkdUD0SbjTzBOiKeeA5tdeyxIAUqUMjs3CCKJN
`protect END_PROTECTED
