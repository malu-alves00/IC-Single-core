`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZT9AnqkOL8YigKNcpUQ26ohW6Bm8dGYrggtsj9PLJ4g3pQ+DOrzuPR0+i2VApYdf
+k5Y3D8oi0qt0PbG1rYnuItGZVyKBzwreogWqn6G4P1UZxBDBmxIbJH6m7foe5mC
eGQE1Jp19Z4Ik/u73FhLCqEz8DxTE8TRuPULu8qAAK+Va1s9/utxKm5K6f/SLUzG
FEpWcjIY6hVAFl+/gX2SR5yCp68pIJwQpER9zjJlNxu+6er/T8lnl77ltOVkgudT
keeSSWcILti/U4qklTF3KNyTGgzrHQ3cYXnFbxgSudPQEdBoY+UUBjTOyGbe5fOy
DA57KfgSC9cOxM5tnGgPp4kLE8U8zxtMTVyTlmNWNbUFtw1k2AMeSF+t/89MPGff
lch0diiSXQEE+WyyguVwL4pRGjhAJeNDqqvKu/OZBjLzQCfbrWGvT00KlA30whrl
W7Q4XMbKbJ62nwjSMt0ZAAKReLRrOpIrl0fGFUrD42Ultg+SbU9z5nD4gmqboCab
37Rvtq2AIHM7mJ7QXDvlu6++00NVyQPA6nXWCrgnJCrAE9r2lChsH/wn2DDyLDT2
/mhn+I1hsznfttSAth0NfEpA2S4aUpQSWt/9FCrVNnMXJ0M2QevsdXcjO1AevIj0
zfH+UD1xLS9SONjjgK2GxFcdfOae5xInEdRxAiL902iVgNkukjkUvTc3+GDiOdKn
C96OyEt+OnAcvjI6+R9g1O0ycwyrrmTazUzhKHKAOhJvXMjnt64RepEHt1rSSmFY
uw77JpV9zu/h41+cmAhf+78lw5AxJb+gPKc5vwSaJKdpt0QvL2jKJWhnCit58ptQ
XyA+Ifjonwxfo4e6A3imD1xzEAEvHWPoTUPLSiShKvYkQo1Ip0kPxTRc1eo4ge4K
XlO1fQv14FIBSFXGTSYIUDjvBi08rxnFGFDNVeh1LOwTSxHWk9dVP+F7WUpGyrHc
xjrEzVfdoOCDIpp2fR91q8raWo/CQMYl0sfswCSqwz9hc/400dE5NARS+RhCj2Y+
vWVI4OoZyCWtiI/pD5q4a4vt5p7F7LF9bYJlQhg/6ZiFOZGbgst1NzslzsiYz1WL
lA7g8kbrRw2OZHUm6ACWS4LEqF7NFVEPxMgBjqgWcxX9Y/degAR4kIYFmEnLETlF
SL/pqOIS9Z0PUr+JIn/x8752Xo3pXODQhSlg9TZ1K/uOmAbhCfygCM+m5/bROODf
haH3UQzY1i1/WdgqlmYUEhYKDkz1R/7yEVJTAcKzKwA6szaxpSIbE42Au+9tVIGI
OjCJtvJmBT9CkfFXK9YEWoyrR7PP/8jo6T8qMGQ1TpvC1WGxxIH2H/zQ5ZpBgkBE
X3ZmspTG+bBVRv2GaUMr7fS9UyZo7VMAzlh46vIinZf+UwfFuJXIwBjudZrIRd8A
rbEYklfZnuy8fmAwAA+lqJVKK0+jUSSe7RCeeSEDchTQTNyVbn7hm/tDcilPNE6C
gBYNZccE5L6Ime83/cSxmkAXpGkEWerpi7YKOcKnIRt20y4itw+GmSZq42264324
5wQJYUUWo37+L3WAsZQy3RbCKwIrEbEpyF/JgN7m+QEjJS7626tDEksJSfID0IjS
qnRTkBBqrJeDMbRI5TBdKY9m7vG2wTsPrgEtw8+cM2ymu8iMvR981PdlmlFb67f0
nWqJZyzWWQqud0EK5sT2EOnhMa3YUxwEsiqsySxbcyLjhHlgpZMwkDNn7SCFyHk2
U5iwmd8iWnnAqCTplNFnJgKPqSMGbojno7T7VhmYZPL5UkClzmB6cepkcqngtal5
V5DHz9eRGbQOdmxdz9PkDlZ20CSaroz8bdnK03139x8HjaKBiR0R1IAqnw++AXxq
L+jmhTVC10U7C5aU9p+KVZRLzgaX+Qv8JigINeEt3dPfpqb/3ipj/m1NNTqYux9E
GjtNolBR5JEcI1PvVJ9cyod1z7/sBVH+v5olEev+/82QBXY7kxn5LCcEYoh+1g5Q
WHbFQbG/LdK+fNhi+DTnTOsLik2qBjs/DpfHgguI4FLrc76rhVawhHD/Qmkf20rV
0tBcx49TjjcEYlGu7qKQ74Vdhv3Sgt6hHV/MZgdQ8MgNLSlN/+3/Y2NUg6AFyjVi
FF71cazcC4If5TtZfr52REqTq6MojOuFl+ysMaTnAV17UWoCSwEUD+JM2X8/5MyC
3usEWNyW9aMZ6E+bBK1c1Prdjhf5gkugF5iPoIx+XwJh1XDh3SJEIQsBX4s8eCVT
V4GFoeqhcSIbGYZeCVBeFMacJ3QU7Ph4pSHLgn9AlDIX4qdO97iVTDhdLXXJB626
J70Rk2PFlqO+qfS0nyUoPS7964nWDSI7zkMzfuA5p3vVGMzzH3RG/B/6i8TccB1n
y8SewFuPnyiTnmGADWNbvhC860ZBYJqXmYC7XE1tx/H3PUgr0lkctrvzTbAW/tTL
iQaDmmkQfiJV16Fb4+LKzWvEDDOQYkeH8DLo/jU0WMDO8QgOrQw1VbJolqPyTTq9
W0C4L9C1TqfaOOxnudUK1nD0EB+wXCkfhDDw/zYqt+vcF6YXa/NibIL2LNu7dKrH
lL1bm8vihk1T2t8FjYZMz1bnax7Ft8CtaVWPQS08wxUn6F5/Ht0l1Tt2s/RwuYvb
crS6Mdbvi1KpEFDtW9mWnz/uB8bg91NYIn499FqedXKDiQotSk+eZ88tu7kQSkEU
WXO1YL3iBmxzwW53y2kiAZfpGIm1FvLe0+TKaUoDd56iTk00ZdXo0nKp7EdZIMmF
//sKYqozEAJkvC81gkJ7DRyd0Qw1Gk3vSO9TOaq/iKcJufntWBg0telITw8bx3yz
EtjjN87l4KiFXHNChHkWFqxVuXctjumybHjNC1oU26DJED2fBuyhTdfYGz8FjZfG
RTQDu+zSb/l82eXni+7CKZyq9lMBxx+Wu/BKGp4VJRUrLQmLQCJDPkAQ0Tvzxa94
1UkEaSklJU4Cr4eMB4ZZBdcE5qFjzXT0HFTA8gfEE879G69MXrf08XSQNj0a0Sv7
e/zuO6LLELP4TSbVHVta764NyMQIvtDjSwcKwEedZm8zQ/I6/cAfZZ+oh7A7/58a
Vcix1FI/KWu9Qsk/vzsmDiR4xtsE/cZt4U8Q6+ua+03BsCvt2Ro2TdshTRQWINRE
TGYUgJkihPMh27p+lw72KehtEBL9bCyVuWvK8Qyy2CWyct7v4YU7ON/32h2bVQnt
jAxL8nZBsnLluiTCa/CF0AhkGnGF8urYYskNwTIWpwrrhwq8cv5EyIq7xb/+O67c
vzvsTyoymAYKvwASZOTDJuFBkZE6Y0qkrf3oTS1SCbvZo0eg5wRL7HOLzvE3B5Ll
hZD6kLFr6LwYZjH27/qliUdrHxYPWz6tilPBxxGEOI+6XPqqV7wPfDDjxC55Q99M
Tw59WziQcKQEXDo1d7R3kbhu1AE0mOExVpTotNc/zGD+0ffhV9hAodlK4Ier0uoF
t9S3myAZ8iy4ruxFgqQHHASY5myEPA/MucZtG/k8dl0H3tZlpKrrV1/djLVK1u5a
OB87eAsKAcEZIPFN615+K9YivYEG4wzvdU7hCErDvD0RZPAP1USlRl2OU0l3XcCX
8TcDHgAATvEgqAXXWch1yPOfrIBpxanVCq6AAioDGkaVXVQZ+Z3rexLFW6yYfuF6
WnQZT7BTrWEtc7M7XjV8pGpu/egRwoEcBDi/tQJXZlvgi3fB3VWrT+b7m562TyWJ
E77vRTgXBQRpSdvbJyJaxKqmVf3TSQ1YmATbCLL/O87Wy1suLNPL7lYLdmj9XGqe
wGa3xQZpdsWj0kmDeI6Fxfv2GZPecRpKL1iRod3PmsOX3D78NZPkDqF+ek0v+tIr
qgMQA9XLYPMsweEe8LgVPk9D1KCb0wUPn6IQaY/EZV+C74tT4GxZouRMWyk/7YJa
a+Ait8dTc+l5ptzrRCZFH14ayfQKz5Nne+2NJ/euLmxy0wZ/fTWmrXi2UMfze0Gn
G6+s/0oSWkKfV3mdC340I9XrDk0nsJAMzXKSutXMT0AMBIUT3aiIUUu9Lfv5D+aI
wEuVCMytQqezuKxCJQDRrltZPOyguB8l/74xbnzdNUu9n52mz7SVJlbvnx8YPOg4
MOhIQi05heXZj5flqmFpCj7Wg1MHHVWT4X68mfZCzkMBTT3hCw9WNMYUbzZoHD2G
TUMa40STNEsWaFz5R6rwSgxDunnTefofUJBLGZ1aZHA6piwM42U98RB1oCFOR788
P5rL56Fu6gQK4l4qlZjcZMxGahEm40bv3myvbNm3DJ61Qb3z6HCbK7s4KEHa5pOP
pvKHmBb2dLgA/Glrk6XRNNLbQXAetTSwNcfnFy5WuBCMDRchwj3U4YeTUpElfyEQ
Bl6XVec0e6iz4+39olU+UxWjjJEb2diDLpiOpWpU0fSwDXVdyDJpfuyZPF3EiLbf
xLTkGinP9f3+FYu/axSxR+FpjztwuUQlG3MEC3Xne3t6ZlM2xNAAH5KBjAIWSwek
QnJIfL9WxR1WlnZqz+LBcvhtG/vj0oD4C9u3bPEkGyViDIv1GBxsMuWYd4jVJ0Of
eLk2uOGvSAousltz1xdoie26n5TD16svPf3vMY2x3b49onQj7m+Rr+AWI0A5CXwn
070fBNMcAXtA/bc44wA895jOfqvuQ7a1X6s2cXoRgUyHq5Dsrf3qxgEtnGRsfew+
LKtLxllh7CH63VXOg8qj9cgTVIIH60jY8muNyHrL9T0mzF9nxiBNLkUowv9oVr+V
uySCSr0NpO7vATquhO7cohOUBoaU2oeFjoUUw0QrqCIoRDWl81EIw+yTO+3AR2eP
WPr5anE5UXotsENPr1RBr6XxKhJPIFj33tu+ESHmnUgl1RUbyIY0v9DbJtnRgwiu
cOA0xofnTtU2ufIdmFLRXbQKYCuRHiIVK8DJQX5JbN5OowvAfFpCFiCicdBszSF3
ZNLA14uqJSWcIlLbNs+7Hjwt7vCwzNG4oYeFejwasvcCGku3a44cScIAjTesuGqr
Txus9ZEpdx0b6BXb1uhevxtgjV9DMJ7KyyGfmdzFuhFWHAa/WK421ERWJLG2Qy4+
MTtyI9QqMhX2cpmagjkutYbuuiYBaP9N/oV0YdPQCPBbwKJF5L30RqVleW8OE2pM
7pMM8tcCcBZeaaSZnW5dnYl3Et4CUuF4loXa4LWT2OmNyMJs9GHfn21CHsGYB6eW
gNSyUUknzz74A64jqfAFDMrQlYEAGzG/8xDL2MG8PL0PIuddxITUugBpDiNYb/cn
PhxkPsRzKV/XgvcxoA1muiqXKCTg5QnIUxN2TyZrn8dvxmLrYHbuZCHH3tYbppcn
Dk9TqrtPnYB7d6BuFyCfR9fP1VOMsc/uyju3afSAplenN/K0ksZp2VpN42UW525G
iIn0WGYs2S6vxiJUKY9uSeGCdKYi4dccGAKxxHd9roLFyCVhqebRs3ESVLTPbj/j
mbiS0zkJ2Lo4dqzeCxWiggLixQkFiawwDBHeW+f399bd3QH1YcSRCb6lejWkzIVw
5+wDHQrEbgCiWDo+HwgLS9nrRaqKdQqLG39zD2NaAkWVpBZsYWk17pkX2DILZmIY
oDPKWwpb7zD1FQeGHSDrkFmvdeqBJUaqhEsrmEbnFxf9Llk7Xm4Fw0f1lwN+63zF
txiZsYcCmYODy2v4C/6Gb3QHeIu4PzinctFys/LMjKjaOX+PMSSY/VCB8k7ItB9b
wiRZXlw0mvxcsMA5UOkprmTx7IsvRPxb01sr8ZQcunBSzGkLU8NZRcfzyKfiaVew
KupQcx46Jw72Hj6uIIcsExP+H7z17TAXteJ3EM1h/DuErQN1fYByIlSuz5vTa/VK
OuFNs+ULm8hVsPKrlJrD4uky9afRiKctNppGQo2/38LSwef2x/BcMZwTkK4XaRf+
GGVlsO1QQGJlNs14sCdUkGUZYMA36AFgFycq83qpLmqkdmPdeuaY5BovINEoQMsJ
YgnPugllK5Y2z5B+B6/noPVwr1hgr21G4+6eCFh7MlV1Nwt1mRb3XurxDS0y8o9W
POSmfTojLz0tTyYmTI/YxRXfPVYmJr/v/RNOcn/haanrvafvIYyEl5WT3t6nrjJw
YEqJ/uZf/EPmX+jJ5TIKUM1EH3xGsYwGIy6Ij8OS+9yGojG0NoqLyg8vdVwdL61E
4j3KCajxUugFp/m0UQqtm5O+bDxP/W5hj9r2B/VRtDtK0BXb3unuxODf6mWMUCO6
W72Y1n06HGRAzQ8XhY4t00zPLknQtQTKdwX7bJCS3lPoQmHLrDyss85EFyCMrXYw
Rc0Uosa3VCBNCKe94Y+2vad4S0plArQ5N8HZrjF2BBYa1tkZgepIWNCKW7/+fvph
pV+tMpt1PPKPNkvX38rebF3cHNPffpHJcoYuIJoOjFfo4brVEaQbIMZjVXIcKVe5
y2nZsTb1bBYfkyw4wgA6yEuD45IqoluM8ul+F4lCZr+9I3LOHFgrNUsmNS4qPCtV
Ap6ExXkuAeUozrySRDMqXbmxm+fPbo30I7PettGxccOw05gZglGQtmWxobhYPSF5
phRtpGPkeW87aVzadkdgOIIsJ0SrzLKn+K7c5CjCZ4pn5M8UeOOIu7ExvnSF7Lcw
bgdqGW6cXagHZDKP0XN9vO72JaaDodw3sQA0WQkFG87LU2AnjUpSj8BtvhwT/H3m
WfNsRibQ2MOfLICireElvne/QCw/4KV5IRefqrq4vaYzmE6pfjhlzpEeVWl5yxBQ
6OmNIw5PL1V8JWKUBxQzhbPsqOgKof/LN5DFVgfltR7xHb9BaVcksi+UzliXowE0
5Zx4RrcM/19oa+yYfqWw6yHblMNB0nnoqyiFiuZq3ZgOF3ln2s1wNSkARfachiiP
ZF6dMZtrbDjPHARMTEmtnibQVXOtYGSZjKPO4EmUZEnALAAGMGqVV/lLgjpVA/27
1Du2ehXf4TnmO6SXIU/oqUJt+OIgfoF54n+eOKl1IET5LH0GO7BA4R8uIUXF59VF
FGOeiZE11mC1OUO9qQpKttyqm6oWgxvjcqRQxS+B3gCYDXIq8pn+lBxiunBDA/Q8
wvJrnOZTmbvcuBNmXwS0GvNknR27YPtl7UhFAZxzvePwq4UCNIJcu0b8HNB6oYjR
O/36cOQ78KKPnip7YVRIT6/B5SeLRDFb9D0H/TfrvosFHSMarf9NSXhhIxGm1L+v
elJpNuYfsMM0jEKJ30eFlsL6/ppJ8ZggNGnrOKK++BuQKr9bmdNyhln7sLQMP7y7
yn3NtNfIG50J08P8HLak2w9INKjEDpRjhfDP2fkh9+qGi2VxnBIput98iMJMhwSg
yaiCe3XsZTSXrL7IHoo86gQJvBLruFbW+tYYJVq0YZnCBhRLWlBA5tH2LNzqYM2+
XkUkgTkWDvc5APsSW2fTlL1HzmxsiLgNZxTUYQZWbrHy2mz7n1OBD4yibSynQb1+
EdqYGCV9xu++bGx4zJHxFQJWejh3xI/4jpCyfLC9P1lFTVKGo2Jbl+lqUakM4T/E
ALltYF/ewlVwgQn+ntQjE4JfwAxte9zCM6Qs2ZNz4/wp67WHxL/Y9n47x6/CahYg
V/LMgVfZJ5QjkFfseoNvbTRrzbJhoJgN5Ad/KI5IRlrmMWqdTiXShchMulGNUV0f
WMOkgjnCir6ac31yEXWcpxj69GQbm4pMZgOvGadj0IBiQpzeRu0NgFyOpKIwMG0Y
W5Vvpl/DWDinwWqsFDhbv5Qa0rG9Qu7iJ3bSTwqd6csQZ8Zy8GWJnHOeC1Aso+y/
tNUFOm9/feXn5RI+ptuAhOJ4oS1GUfm+6GArGQcgqwl/qh0Azz6D9IlST+VwaEj/
kBShSAa6l0lUnXxP8LiNMyX63j9aHWAGYhsOTnktyWmqR31YlPvRKruIVrVmwwXw
1r1Jom90rlA9f2hdQF0+Dk8yLY7iYylIe6QJwERVLsK4eYnqQ1nkm7uQxGP2MZe3
s5MGvBnJpSUNXvEwf3FuO5It9Xc2gi6EvTsAJoQqBT6+BpXH+Ud1M66Ir/9YYGbQ
3GQpUWolJ/+5C6tld/2QNOiXJIcivcEQu10eqtH+lBkUtowy4Ri5RWsJwaNyokqm
VAqnLs7AFY+hwWiKZer6Y4ISkI7Omx0fUWHvVzcsquEQl9oVi4OMyWKrSteiqSia
CuO/1g2ZA/AJyAejhAY5q9I5+Neu8AvCpTettYc1c9j1P9dxqMVrTyOz4PiH+8DZ
Cc0GrrM8H0stAU5HuC96ptshCJJQ6V+Ou4pY5ipKYNRHE3B+9bsCVSzoGeHZ/UAl
HgrqW+bhFlENYGpCaT+RqngkWcT1Wk+ZKUvXKTj2O6R36NBxXYh7hkS0xA4KYZyv
v83hqo0PvxF0hhg79SRMy9PSmehlLAF2zusk/e91Q67+lP3P01Jlj/FDaNpf05O2
7Gurwnk2ZlkYr05dbb79s66GmT+uxKFvhYnwuJ9BC91sDczZAK+0ih0H39PZxnt2
4wcKvYzn+gVeKRUY5dDznGbfhZachJCvAqrjO1MAS1dBMzO9ByJa/FBvvQ8HvhzP
bVflpr+t/AjgOziUIBJbfaucSwq4gna5lU432artpMi5fgzjJAingVRxRZumFjv/
WeaKIAUR5b8F1Axj9IV1+U4W8+2sojwwVqd2wsgTufS7P3QIesNGc/TPIov4J25s
IyjO075SFaa6uNBwgNhP7SC6va1B/GvootRRWL8M18nbwSzZ80eEIfYwl12sAgwJ
k+l8ETgq3kP525EV+bvUMYzlgMiHLs34hU+sZHxpGAqOwEgx+uywMAReKUzrsD7E
IwItG+cepllrGb/Sy+e/1GDmnqqLLZbbQeQWdsfUrmZPWF/jxAG8P3dS031Z4Mre
TmiKQSTRRAj1q6rFOxL0pgaDg0XSalE4GgfVJRmQjSTq2PlXYmpadeWrA0X5DmXi
9aMRO9h5D51K9jiN/wvxyZ9oj8YL/hlumbRpouzNzCYgi8o49TUcHMBfV2ECZGaQ
NXDyGKrCDxVXOZg1/MjmBkwoM9BdzqTTsX1tr5GlI7R5UXLFPNtUx1VsqC593/Ib
gZWibv/WgU5owJsXSo4pcpzwXejnoJsC0UjBvxImHMjo0fPsvqG82LW5XBuW8aPx
9QzunhEQLqDq4XE8536tIkKpT9VTbjXTQJMjRPmFmm1ru1939CPiI1uvDVK8WuMj
q5C/VNRFJrX1oj9pDZLzy9GhSlMBY+x803ovCY8JYdX7Io+BBk9F5xBS1+EdGSZc
Nm6DK/o3QwRPmBa1Rom/gIlcdtPjq4duyRr/m1STJnahdLyN4qjwIIo5s546AA1Y
6pWCkKgsi89NcupMDGiTt3k+sNE8FBwTzVrLwtvRYRHrirVO2Oho9FclCKZ3FKuZ
9pO/pH0RKLQrGQ12RmRwqhLt3ME7Upk+kqci0CTOum3zJ1wOiK4lE65fY/BU3XoY
Q/dCjGGZYaDSQ7yH+t4i/IR/b9o1w//maf5WX7419zWEivBW6LQC/VBDl0oSn3tf
zX22yf8zzQIEyvOidiEHVxCz+ecuRqzq007+iNaW43NpFNrGwWOGN3KgcEQ2F7p2
hANfVm2QKPyZ0DxLpWAK4kl+f+mQtgqk4RuPpfhAj1eY/AFExIUDzUBVt0GybDq4
db6NKoFkmdFo0X0mtxUfrYbe1WnHwZ/fkxYyMyqXQj2yorcrT1TiVS7I2sqnIpe9
bislJbDZXzKzCVAgArKTpNHCCfRq8KvjIA1omdvKjQ7oTP1rmAtsSkjovc+LNvfU
SeL7VFCym+M94TTzwAWIyJye7EQF9QLjMK4S8hwKpiT2sP5fABkq6LNeoaa/RTZv
zCctcjI4ef9HDnKDDsHPOebjHg2HgZ9wRvXOvctR5UQVLm5du4zAWH/5vvINLnBY
FfoHGx0RBz917N3710LykgrkPLvxrJO6h9Pb+7/YpYGJKf1TXAAuQ6/I0CF25in0
m65foKvbRQ8Ex1j7DPgipeiLEI8yvlzch/UAeEOB+Yq7pJiJQfqy2qCbo3684p1S
fQwZIEysOe5OGaELf+gTEO8e7KdHTXL9D6loNEbsQnhwPQGQdC+7T1cIzzoxtD5F
I9JSTAxcTTPzlQztc6uDvPJWCHHQEmWeVA858xFwzccCHQfJyZ1bhpvMix8iN1w/
K2LTCZPcC5fVdzSdrF1t6A0IjazupH0JOEcscY6PNgcTequ+UdyFAOoGM+hhZIak
xWGbZtuv9zrvr7CG/4ueeOr4naVzSbJTcS4WwWhKyx+zuMrHuZ9w+hF2ieKRTLfY
7Q/LLw7ZnaAa6tb+xu7WpqjbAmgVtkUtQ8t345BUB1M2WSQ3V7h38YP6N7+DO3XG
EBlC1ZEFzHN1leB6g1wUMK40oF1bE1Vj7+ghdi2La3WhYfFMYBLSksJ2mjMUlLNN
tLCZNBNb4uXYI5z7aeuDu+ZPg7mAhDenh9LrWUYT/1bg2DNZLgEIKk8Fn2QJznmg
xEHlg9wyYsfLx21xNT6JbYtsJDZd6dgXUIjTiNcuwABq7CnocCnp6Lr8eGbrwR0G
7kTjgxo5xGpXkm/gTgShYbGxWowQjs7ErxBXSkM1JlHGE0G6qrNkzz+3TwTVQjlw
R+sutL5UCwmNvZyAfBqQMY5V6TkvnSFtwOmF0qEr1NkBi+GqeIOSoNqB5oAPvyMn
4qzmlxY0l10TrAtVzrJCrwJulLRjqxJbnNiOhmU/I/vLJjF0zld30xtIAydYEiIi
VmaAGLFUZNDVBU4tYe6vpNcbQd0zlxJgUD4lEuoh8r+dKjO0OWeUWerFAYTYE9/q
awIF7z2VoQ7MMJni/tEZrJsXJvfkmxc/32W/lAqHnbev8NlCR1pQ8771b//ACO6I
o6ce29gASOJKtK4GcToYC2TQkNSMwfhnR5KP51mv9FdYVZsHPZydpz2MQGLp+n4W
bD8sNnc+ZKGAtqgkUh+9YL7pZFYKxPcBBPOXkjkxw5y9iATqaHBEf/ZoVcUQ4tVB
1kXrSQ7/TWIprp22G3yqJzZsUc1LxEZFTkM/aJRto5LrcZiaM+GLmS/wh62xB2D7
qdgSou24duquzFxxZ0LWNGqQtXl3ZYAwUdyPSqh8JR1//VzXck9IjtEPehfB7vr9
nkzE/E05odZrflMiTsaZqGkDJB8rmp5IU7LpFIdabN5tjlOhO9nYchXuRMnXJ6UH
I3q0K9QnSNLyVg+N6/T02E7shzfvLTbdBefVhE0ZHiboUei9zLzJ9a4J9NaEt/7K
KHqiL8gwOg7u391841STrnRvdU4qOXDLarEQe1xv0siN5RRvL5MW7o/AOr25Z4lc
1NJPxtS9978OlhBK3NSztgxLwgbS8H3EakuBl7upGhmgbIK8hBF2nUGUPt+n7NXW
ytz4wsuL2d72aynF3zb57LXvp46AzocEGYyfRSeL+vX0avqtamBeuEryd/n+cdtQ
uzUVzW83vX4nK2BEBKO5314Ed2qUgUc/SmUK9/STUcH4TydTR/wSdC74ptMoWMWz
+RXqFfUS9hcFBYs+QETpWw6jimv2y8wj9esHuCNoMx/U5cpJGSuZcdeAILxYCsAg
QvX2W4dhbEN2EiLdl86syknltiDVgiYX1lroK+MZgF6TzDMCI9+RYfc9e2bTetI2
NriSuO4L09B11tx1CbX7kcHvJiFEz2s6RNQQhfZF+PZkTTpo9VfhI8KMpx6L6hvh
z5q8hcXz+/nlkCxhACfacYcITOvoH6jXjEFPImAqmSwicIPnZFwhjW7qFB8GohPl
bb9TXX2KBOGBYC19fZ8it2n4aAxdGVjBJW9HetvwQoz1nxmBtKpGXXd8Od71CRLd
yt923KZCj1kXbCNROi7RUD8wdoH4HOAeq5D4lp2yYkYWaRgLYn5zITgOmmVEHfWY
raGWnB3Mcaoxg+PWhTYKQH3evifD5CtZMCj0rxhSsbRZ/y+mXkY+sHYW8Ev/du+E
t5+CYpP2fD2bXqE9pdcy+Enobl6dPdGwKjD+/KLRRNt/gpU/3QzW/DkuLdoZeDJ4
MRpJ9MNzdorcyUq/spOJOWpDQZh/Ka2wBWOLlRlcWTUXrVJdDWB5fG3Pp4UU1FH1
SXNyN9y5h0Rw0B2xHDIwbUgAiqo8Gls4r+dWvl5f3UaNHTxR9P9VaeMCLlGGfyu7
+67TVA5H8/hJKN41guuriSsH28nhXvU7u9xlikJ3jIADtRrkU+OmXLyx/FTWhlR1
Mo/BewfjaYgupFBj9uqO1zubaD40xdiU/0VRPPRV82igjgM/ZyDlgEJdK6aUQ0Ss
zQMSBrwZnPx639HKdIZxdh1tB94ofWXixRXCx5sXo66fKqO5xWonohEwp5cnsT01
I8cTRRyV01JSh5S7gK/s0pofUjPglt333uKjEfFsj7MF2tWWHDhenn6CftGWTSSz
XDy66hgHa+aFzXdYcmoJjvcTjDot7pPFttHo334jrJw+vZRi+hJ/F3pgDzMyM8Bt
nTPaZuBWypHfOKa7nTmAbJW27zeRHfJSzgbrnm4CWdK1RDk7dF9TP6CAE0nksGj6
Ib6jrQbtGXvkmzL2CdRHnYaM5xRGfffK/hpowkYN7c8PHcRnrQOZRsgdD1mMflYT
GcE4TunRkvtxXur6ti/RUzcfK+uVSxek7pelbokU+qV4H/m0KuETpDkOq3C+6Qpv
8bBiwZEV07PixFYo5icJ2i1gNU2f42TriwIoE3e3iLfQXgRZwfA2IQwMQcU+XiTx
yG/r2dVotCVwf0k104Tpm/LMLmG9nGyr/Z4gTEGokSB2BqbiVhnpUFHO+O8v1TMz
9qyKIp38rTDhw0P9gfpLL0e+ceGGys5YEe0fVWAhiXR0B/HBOba5yU7kQCoewAkD
YhUBTHZhsFfEkdSKQeHN6AWNlhrgiF2fNnygdNIcSr8RJRvVMEDneuQJTZzuWFaO
4EsS05EiolGYdPT5Iv2Zr0HSl8+HSiEdcxs5UKFCbuwvZ76ze/pfg+dvvuTX1/fA
pfDMpjyhIDiHQXLkRxvJCpAGCRjqAO+7k0xa+DdO+HfM7/LyhWFml1AqYYrv7kld
fIP5MMhCyWnP5bO6SBywxEcfwhI1Ij7JRkxcJVk5TJZVICKQvAuXJUHuDDMTDBJl
vegIHCUXsfip61ApiDzL88ESITXsjcoc2V6xIiiFlLry0CADKbS9xyouB3cjziU1
GvgHXDxjvGhKSMeWlyA+ZmnsIpIFBMxvi2OT9ZgnfSZnthjUsfzHusNn1rVBCxZU
peh4OWBf+D9XqQrUKMvFTwbZSmLKqaolL2eCQBfQehIZc+0HQOA+/5VZteHs67YO
Ps801E2Vc5ovKDpuwZAbMHtxfdN63BYzdOya525jFWM6hqnQZgnFtiaYAMZgLpcV
ELETBWkCpoJn7URu64tAYdi4fcNcuyz64RZNACN1tMZCO1uK1AkRULixpJTW0AJf
Zo42XMkX3uc/77sIgG9BB44XQppL1pDkF9Om6Iu0UixiTyqvnEi9arFi/PaM7C3T
ODu2UlPRRlCs8JQZKK43N/2G500BNr9L9q1CPp36DpnBEeA3aD4qj1fzivJ8yDIn
+bLvlgpAWnHaFf8kv7sOcCvShRM4U4UOhg9Aubdqhn6Rfoha9KLO9lEkdo8QK45B
SB/wIE+eJ678DuGqOrCPrPhMoklofFRlKG4bS3IV+tG2m4ymGrgUhWyYTpnR8oG0
F897nzltaikj/l+8jmjx1cZcMdJegpLuTXcLbrWgadl12x5PJvkSeXR1nOjSgwma
soGfzgJvlpsMUIWwN/VhZZdyJPqddsUm+dAr7uf4cQkHrWxjAdrIs6pe3RdvJasg
b4qmWPrsha3xDFKOowW+q79YlCGdZESdjpf9+T/ZM3fa6fil1ksa9RL2eisfD5bD
bxXyoE0Mp0HRXBqbXYHxDoVH+ZdhnxZCFnkVJLKJuBWnnv2CFbYycWuaBpM87Gbj
tNX8tYSzEVt5ByhzZp8nndUbVyHA86TqgrIW74gOk192fgybHUKG0iJ4//0F4AYA
DuxH+aeJ01Q7eKag1zUp3pv3B+1HllMGzXrTA7WdqSYuT90kzqC+tEnDpWRRr3mA
mjWXoMO5oBLqaSiBb8YKsp4jUKbzudyEnUlY6CgA1LB7iycw4laPeSv58VI5m8i1
w5/FEc6ubbCVL/3P1Z5XAEZfXMKUqH86CYFKxFUemeixRNUTSLNTQSQkxrXrtr69
ve1TnFGZtSO7LcDI0HVo8Bo8CMPvlhe8PyDqvQm9OfS00w0gHN99qInXflp1N46u
q4WKF3dYxm+56tXkKXAxHflVMERLdW3SONr0kisXkVLBp57jNg1jSlXy5kIM/Brf
conwEFMrCq4+sCRml80Tk4V5H+0dcJaClZLWD2WLGHuJnmM+UoI8Ii89NxJKHCIS
RQfBnm3CAWF+LcseuhVh8BBsm6TJOI4rcKgH1ue5HaLGMYRwLVBQi2IlyyGrk6wV
bI/j6MzA8nRwHhdoC0bVuqMmSZI/pLgQI+ExUzZLc17UqI/sT7JGtxb3YEToeOAy
3lcZMkQPdeqsvuu5dGZpV3Bg3ncPYtVgrA4mMqPdrD35T3DlR2FgqlFzOerpG9CS
JvHrhIzSJ1wq+QCBc6TWjeGO+jrn39pxIHO+57D6SHEoSafuj1ydkXqAmdY9sN6f
h2hGWoR4fJ3rvtTnTSSIEPqblrvJaXjMbDo9Z+DfIsDGuR8DH56NqyhDXoTxUNFw
N+kdqGWqmywZDfiP9XyrvuIGwXOpA/HcX7BnL5qIk5BTtBQ3gyHV/XLC1cqk2IUw
oB0FCKHmIKPVnbxndy5+11yu9/Xh4fh+ySmAIi+3883DRt1lP8lFm1KWngufj3sM
Yg+9aWFwq6Gnswu01KUEzZoFj79fSllChRStepd3Xwx8OtHsJtMIjbLWjD1Kx3OM
EzBMnWGIvwQ1N9CNOXv+dSng+s4sIGwWUVFbSv2eNoJfOzGWh6MacjPodCmuK5dY
rmYs2MwOBBddl35Y8zoAPDnkTsm2W74oo897mWon6zkS91MXHCjVc+hpWXJdFC4I
`protect END_PROTECTED
