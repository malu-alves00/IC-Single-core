`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zLJV0r3oE4KCCXajdbcLKfT2Opoh5pnIIGQkuXLo8aZagnZZ51aypbXv5ZBhRlSZ
mWBJfl931LC+h6BvQF0bppdXi/4ZHOlk/GJks1cA95kdoLRc/n9kQeaE/FutRbrC
OpNS6JeYISWhptf+Gsj45Kncn8oN2i1Ogbwq/waptDSW7H4OoSptlKkfm3yQInjq
5k7UbJafewkqWz/3313lAEKNPh5PVSlmJ5ig0+Vhc8PteWMMdWSxTC3U2ScVZvUG
+2o38yaQHHNWNYo5IZmOa/1Q6tsW414boL9soh3kNrJPb4636LOnMRwqQc9D8SE+
1hbbq1Xb2RUOPsVXNlwa2IZGO9vcTOPGuRXiDdflrnD8tMAccw3S1lku/BzYX0AM
1yVsDXIdd5E4xbJzi+sWeouSlw54HCCJg0sYgD80/P5sXpI5KglZ3yKlIJgVUNmw
x5f1X1JDzCNjtZLrYBRVZkiymFaoVWVLOsrGcA3CxDrfK4CaBbVu+5PKTRxWvI0r
nHDofyQpDMQzCCdtogmUaF3nZYyoouEEfE0lMXfHe+Z9pMERMuCppqK2FA7Fa+SU
UWxCHxb/HIFFNY7HM2eP6nGc4Km2SQMy0x6dOywVtSKdmk2K3e11GiuAb2RoL1rT
hwUnIyRbHYZoJTAJRr4fGGDysiQmu+YwBrs7YyDzzRCB//vJroEzGiWLAYiwhFKH
N7pitIsmP7b10wlRUETYRHiGEpSp5+KN61ok5iYoF3mP6uPvqBLK9fcLsJx1vAL7
vukDzfSG2HHSp02YqKKw+xPxgUQtGeLY2q5Q7Jg2jDaST+3Gbkh6MeSU1Cd7NRJy
MYBm+zuI5/LuBFAVmhhfULAygvthMyhT2MsKT3dWIH4Pj5x0oUw+B3h6/5T/qMIE
fdM8bgxwpo0FAJsZJPUnF2aWLdk9c+0XJ46ZBvyTGfqSCIc2sEKh+lP+YUbMnjIf
s/DdpJjmkIOsfhEeiOdolx6xS38tyCz9/goBpsZbmqsGdzoOoMwXllKCfRfxgPvd
c49jo0ucXUQKDNKYtgjHAzUD8mOI4PjAj769MCQ5UYj7y3FDrXUb/CbopqeToRi5
osfN84+Jp7YaxJXVLvkjbFMpLGeqkZ7ZyMiwC1a28BQRT8MRoRMDmOxfoswgFk6E
8m3rvNwEkOYFW8dtI83RZ/n3jnn+VhftD6O3CjG+jaVsC7xuUT34l4pKWfjkCNG8
P+xuIT4StESNU0QTv0J0+2taOggKw1LOeP7X3nfFb4h3DQy864w76XzMckag6tGA
RMGW0VQkj6R9RRhABbNS5LSdvDezcu2WPAQ7IOkMbWLvlBsnaBFc6Sj1zDlR9RQl
r73/zPYj8L9Po0kotqZe8KAGM4D1aC0f0MwNuewr8wOr6vCBXACSbQTfuXtsN16B
KUBq0hlP3YjodfKoOH1B+b2WGvhI2v8hZs3Yk6wmzlOqAPwgOClaBx9YOmW7uHDq
uBrGbiewXg7cPBKBqGh5R5CiFYdA2d5a0oEjJoqvprdVlDkURhLSPs7VrSWwZdVJ
JM6m0n1s5T8eT3/Awf5XlxTEblN6u4GkoX0lrbsj64uwb+W7NAlGsOhG9FIdgrHG
zq2xsyZ1B+yEKMYpUxcQYEjCTlAkbcfPvX10veECcM7yCQj8tAeEpqnNyYLlrbHH
lbLrph0WVUx+cLiCmPtsueFWSZfd9SCgmODOKrAXh3fPoJ0zC8evsIH/TP+Q18TH
7DeuZ2YvO9n4qbydgiXRk9Juhu+ESmo2KXPbMg2j+xhqlGV8B0prMydPuJn/eX2Z
Z4UG4qx2tezEFW10ohw5pGxJgMH2+G4qkb9qCU8Zi207PqqLjlkQ88w3JMkUcatU
c2irtgeDdmS/BdQLPEfjSJMfx02qE5dgYartbXGX6s0N5tMw3GctsjY++qeqAHJz
MjUodpZ8sKhpYII4YiPXbvDB9vTYYAzl0oS67RZB2SQmmG0cRd5yeoX8OyBjPkDC
N17dNfTVhOLuTqJ0AvBYy/bogPd5xp7uvLF65+MZiiHmHGDtBiHJSsvAfFQka3k+
WI0VtpX7U6zzd1uHqWzEOg==
`protect END_PROTECTED
