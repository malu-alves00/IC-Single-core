`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TJoxqVdYm9lmHMun3kknU4q2ggotbJRLFYTLxKkikjPdRG0YEfQTseKRJ5C7SV8c
uUq+egwTHDfLmabXxcL4+tgon+8PJzh/8LlOSM1It+6B6dNA//IqYZDMS8C4bZ3A
fy+W/pd1hU5gg5UFmhhU94IKPxp7hlgfIcz7eMEzxQwZ4oR8y/MN+eyDAytxzXl3
L+2sKG1Kuy3fQj9dd8rPzQ1lJuCnfoo1NKYSYac2cfOqEhi/++D6r14kWOt/q86v
UTP5niNXoi02K12XGZc27eMPDlva87YWYNmTSVFZ1Jqi/62VBlsR10i2ClSddmC3
hi0yLkgppBNGK7eMcWnJ0CmBe508D6+3dUq5z+v0M6WXb63lwCs5TrV5Ng6+RWq2
WG3wwxNiAYn5zvMae+DLOVVdJW8xzX0yHRAzxOvmr5LYWPaGmHeOrZx/PiQqF/oi
8vPNomFJ3yMnDZ3RCvVDW7PRVdZnYnUCH0SDHQhw8tc5o4qYxlVRixhm3+5XBjdJ
iyONN1mSaiYAUKc/rPhD0RlN50woPdS4Gv4qG0N5N1OfBm88juzWr71GfYSSZDI3
ONN0CKcT8iSBEv87dcQp84tEI3OVMC6SeUpqZSsZyRj4f03Sro18AV4+zONaebGu
V0DUpmu0IZbLh3mQoW4l2tXxuh//SeJRKHHliXcMY0mRRHe6Dk97MKrFftg/q/DR
s0GiVmklrvMf/016wGv63u9kYTq+iCpJMuE6XEU8BBqQp2jrftIElM1RaXl+Fo7I
9I/5+0ORTAfeiWboLzE8HqtXCg2YqXOtXH1tsWOks9XPGqK/PUeieLHxzJqxK9TF
ifp4bq0pfFtXJF4Kd18oX/AnGBmxAtKT+x03otBxYz/wiTy47vcFvWppe3hjnda2
hdnF0R2m3veueRk/gN0mY2X8A3DVmgD0gj4XwGlh3rcwARK5NJd6ngXy1Ye4iacG
gLVc4GqUEM7VUQ5xbuXOHF6OEhWSUlfpoYAi+apyP+SDCEenCsXKH9utY2fVijwX
jeisik2wJ5R4cn1p2PxFW/nBNRTlLpMQOoypym5liCxoV3G66wORbcLCyfrZKzSm
Q7yEa+57jgQyV/zNCGzwAoQ+lJI6YtF/azPOTMf2vWX+zDFtvlt0cOGqR7FiZHCQ
tPn5EExRgae8NxfT9YJZZA2Jz5ZSavqZYvzSBYivS0eiB5Gv40kPvOjMDxS2ZM/5
etH/iM/NynznxThRMpJihPUUSzziFObOk5v1i3L3x/NhMe6g8T5ySZMnlhbZFkt7
O2HrBcCtD0CQukhWwnNn5vMP6ewyV9dEGY2ovjtOKRZBLws9GS3xTlWpD9ZWiW2V
iY7/nz4T4f92ItKB++AV/6fTguqFg1KlpkIXsewkystWHh/jcxDJpbKl+Gh4D1BK
0uRK2I0fqhfWV1GhSDF1VOYO3wxKRJ7sCXn74zoY8sjHqGmHktg7oRIZqzp97zSS
qvdKDffjyCSnyFcy90E+YBoy7Y7F3j04jXc2lSxtMarLq9GjxS82H0N9Z2gzhrcp
Cg8AFctO3hwj9ql6VLvxqCuiHSE/AH4p5Vj9qhEfOX89T/dlG9CpFnzhnIokqW5X
BG+5z6sghK81EOIGYicPiyWNWHjhc/bjswpyjTqyN3tMealPIpfEZAKqkYuHffzX
2p7R7631PhSiYLyAtrP+ZJ+QhBSt3VpGJgzKcVf1L3TMbkckp13iYT1Hr1j8qtvI
P42FSjz2IxyS8d+28wUqFMZb3aTlcu3hM0AKssF/nhoEVqYjNq+yHdBbK5yng5JO
P379YalVhDfYBxSAP+eOzIhCKmwwpvFZ1f2A0DZ3ha3T6MpRXFUFHHY/G6Ye6wvd
oJ/j8zmg6Dde+IH76W6/fmFF75iBY1DbmbPH/rvLDgeWXSnd9Ons3haE5NvtEeWl
YwWkohPaeCjuTUxS6TOcSWVstsRimIFqQ8zX2qYgE5l6y/dB9iuyiqgIsM/oh7cB
SUMInQ4PdS9fQ9DINoua+Qa9Tn5tVx+5dV75BDqEhB73sYpyfFnRjOrLKpMkRhiZ
witp5Pe6mF4ENxPKudt2WqRCgL9mBiJtZzq9iPHqp6xR9pZ4dUkHSMJ5T5GJUTuV
Si+XTCPV9zgX4+8EPL0YdSGqkZ5oZpSswDPld//2eC4v6H7GQ5fVp0JZN/WPlSPa
8xeOA23yLrfFwTogUSaVF0EVHja8WECvSMXDnr+e8j5II44lThtcIDAQ2O0yjNpK
BvCjTL6t8vhZaFsIkUAInl3JsIYDez3aj30/q9WJEBEnGs9jFC5YI4m3Afm946lJ
F8+s77WjGwgmV3Oref8RnYTXBZRjhKQUAvAi3uMWUxUMAvoODscw84htbtOhLBM+
wH9mZKzUkbgABWQwuY8qBtbtKv5ecdpaS25l8cfBT2yci1qw8g9DJcj1jFD+dST8
QBFKftWdTfyOszFhcbU9mZu4K7nvv+OFxbKQuFjPTJLvPIgU2B3AqLO3lvZwUFvx
rnYrxJ0fIqGMsmbsxj0qQB7ma0pJL0X0LajzJauMCLZxJpYRkRua8ArQylHI1+p8
4pOOjUhfSGit8OEBxk6VFTdF3/BUBpy3Sc9FpOV7GDZyooKJrnMuAb+OHKPhdgep
zf1Gr2iTeMXC+SpWp0FZ7sWnv/53XxGOx20zoxQMhqln72uVuayw+sk19psOZ16R
kR39Wyr2JcFUynn8w+JhvXNuBTtQWHwF0K+jHSu0Av90GCiKlkuaxjQ34lMReJM9
aH00m/XmMEiZJvYnKpIDZEaIp1MFsLflQEs8UZzavszDGZHPmJ32e/8p5giusUAB
G5LeyxTDazwgkiaEOSmjyJRxUHeqZOM2yjiOT10txJ53rx/YK7XMihGZIDf5huyL
0wwq8bd3ARDQjKWiA7PZB/NXhMmsWs2okvguZf2dgq/HFSYMPPPKvoGPNThhfsRr
a/40oJP6rR93RJ0yLELtIwCNBj7Qk7A4fcun9aJto4A6mdIx2TEsJQdm+73PH/rL
klnlj2Q8nPSV/jYpuLBh4XnNT0xeKDU+D8+YCIdz6EiOkaNEi47VOw3T5RLmnyWv
1l6h0q4DX8kThHf5QUml4y8uz324jCcLfOZdum1HwcLytkW9LIyE2wMtbcGOn7AH
h7d0HOMW5i4XroWuk1Lh/rbbj+1X5AHMVyx7Ns+heMkzRDniCu38G/6SM7vTND4x
m7P/c2THw8LrevADZeE7BV/veOsLirGpeMhLFlPw/O3G+DeDjr6+rljWmhL6N9F0
5RwK8c4TwnHfkfqX5oF+fkpgpSBrXxsZMRrHwHa+0E1RyVCBg06NDNiOcYxNA8jy
9+R6UTBEordH8i5jEuLPEPWcggIiA9wVZJsxmiXU+TnatdQbHvFr6CMyAx+EW/os
ww7nrqRBAiplkyAD6XzgLcBWdli4etzYVRi5lWQdyoCQDDMRh3NIKJBVLrPy90al
d6DXQcxCMyd+zB6CpQHIEHQEkSY7J0zRVUl2WUlziEBiOwuY82oC8P3SnNUYvo2c
p3v/mWNyE1Rh710kJDHzhj4EApyPt8L6NTA7tRBYKnRFGh1fHB6qDL9BzmbFk5iY
lFG/cHB+bv0Uwj2vxLMqpfYouuaGgrSzkMtZDkWLZdWSAimqyjAlsmPeQb+1UHIN
06yADHi6VH6V5YlTPPpxWvErsVXEB140UpqExa0ZRxdJalFcVfR1CjlsbbWMD8mU
l0kLigTgUz5ZZB9IGrFEqkqSKkc0jZIAiJuUmolYrRN4JloiQdAaXNTUL5A30Ole
wAe96nUkc+1cAJjf3kppsfwVuBTf2uiexX3R8/5Mlu5h7iIw1h33bm6q6lHw9mDl
TWrkZJO0t+/S24mUEbQySTxFDLeMfZFQHtwD9e24ep6xVGJhF+jsY1uKZAzkr69e
+ZV/TYV3w9En9/8EQLPrqkZr6DmwCQVQsnpstRoblD0C0hkzV2P+BUUjTk7EgQIz
9Tjwuq6yqr2Ulnuyb0So6G8VZuS3fyEMH8rrBfJIp0pAQk5FQTTDKJQOtR612Vq5
9K+Obe/ejYIQnX4Hb01gutpB88ebld2Dp5ZQYqkoCUAPssgA4d5gtmA215ZOUEui
Mz4B1iK6b2I8PcK2OUiXQJJ1CUJqiABq5YC7VR1kIKWC7/TtVSwZKeJASkcRGFg8
c03ACUo8/cIeLJ+dVYDbg4nzliM3Z1K27Ocvjc3QkdiIsxUD+pTwtQd1dDEc36Qu
hfB/OjIe3ymj/9iN/nRq8A==
`protect END_PROTECTED
