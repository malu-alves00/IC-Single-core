`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BhOugPjByYfIW2pVMhHC756Zdx5LrxtTjn7u4s6EIdwJUiqV1q3bksWF2iITXa/q
IOUM/wZRKVd4TIZvAs+BUl/rdkhIA68k6reMZuU7PgF7XUBU56z7fEummw86qDmX
zgYP+pBrFzBKqjJY0SsTRuZE4htTF1EjyM5jnYvAOTz9U/d3C6Pw3dqv2p1SFNzi
XIbbj+C2I0XlxuEgJD0FdZ7E1VhWqpwxAU26IwlZnFFUFupCSVe+/p4tP2samh3H
RiGeXbhfG04yWl2UFfPpuW69S65X0rhD/wxfFH6R3fx887oMh694bC71g1gNeKbQ
qNeoDSpCe2dDFzIwSk8uDIuqTXuf1+PzV6pkLJx7foufq2xNB+5aLJB5VMG14ehv
r2AU4C6nCqjUxoARWbZkZKhLK/Flyu0wjNsCc7X5QZrsbPxXd3/sH8TV6Eoe6yAB
kBb872fKCJ82PMbesyJLcijt0gnvLe1y8jfABXDoBFsMYfDpx3Rwm1oDj3qEuMVf
T9yVkUAW/ja9Ieh55f/D+6oUvZKIf4FMt6dwwIOvb/9sTqlrRZ0vO7Buj38+CefS
/dEm/5OxCV+Ag0xSkWjz6j/2tCvsamRXbU7cj4hE8TFimZry3C19t6iA6+E+wbag
P0LvjCw35VQghi3tzw7WqfbKlmanPVu5rqWF0fff9bXQX8g2b3wvZLxqzC4UHYVD
cA7rw9AYc/dfyYPm0dbwnYJcaK0eomY9/ej+MYNmmky64XP4fUo8qqhHrD0YiPLj
uSJJxrf0epmrNiaTkt02NQ==
`protect END_PROTECTED
