`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dauBu5q8WNxOFUMEAreOKzBO0K2xvsnE4q5hfcQwZ0k6vPUXxskBt+x8AAFso7JK
mDj0A+K9DNXGsl2LzII9arflJ6kuGVmeiTw9Ntiqb01/Ho2zTQQr/FEiaEst+tFh
zHTb+wH1ymt/dXcURURZhA4h/WbeYhIWTAgQxeU3EuPc6eGSikw6mzF7GDC/Ro3m
iZZllUGUMJUWvfBBJmJOalvB//yNOPrZ6NNr9a3qCLeF+/gAeBSr1m534hpgA9kI
pydO4qx54wqItbFhzjUGp4GEaMot+OgzT7IlIZ8nLOF/o3pCVl4cg+MWDfDu4HzR
wGPsiQ6+/lVVtnxnaL6a/PR5loiE0qFFErkJmTm72or+8SIYMhHC7tKhsCsPzJQN
/UTEvEy4rn8Bt9qGWlbaLRwCUgY+YEOyNR/s0kG80LEAcqgC3BiiG59evArXQXS+
zASYPiJJE7vN9EDu6IlBszpE38JCh4O4UZDB4orhr91CzyT7XzijY5eOI3ohpceH
qCdf/87LkmG842Q9vRzhtJuhO3l4F14bWWybQwu8wQ6KGPf1V5Zhc8FqntJpxRgT
kqK2g9I+OZZU6AKvZRNMIOieTCNekGBqGsN1xcJsocVbIRFL7vT0cSfRDd9SPsKz
itNQ+smtO6ymVBmvPjDHYuj/yrOUgps+Uwja2lTfGRPlMAybEKO+9/s0BjB//L06
8wutyncO55R7xFoyibkduyJeHzULs3kzDbHEn62Bu4uR7vA17PdtDc+Yrdjucd5d
8UMqmjPfpEk5gHCfIdb9X4y3H9KW+YkGY3VkiHHjRYqa/aKJxhiptaDfp2MulYas
yOjCs/Ka2A45OIpTK7U736GWgiJKR+/30qEZOKIlMVYzM/jy15Ljrd3C6cetTcWY
JGjXL8YUrBby3HjxavDfXy1oudsF/0Fl1Vg/3OqB08JU7ap5d43D7PpxICWMUMJ0
VQtabe9VbRAOs1b1htrZKf3WCRlTMgAtPjRoAy00cAaKCL42S2V+susRxkGYOQdd
rMl+3zXQf0/lr+3CtZUvLDY9k5ox2xFB2ujKfK7jycOZu8UfvOom4wQ7PeRrNY7g
bnjBFoe6brmytNNe10xzeFJyhBABVyFEtMHDPB+fKq2zSAFn1jet0Vd10h0gTcs+
OGlMIydlbV63e+9ry65WwEVk57nx4HsU4+L0cVbhTTXYYawIMjykiuZdm4cjPjNZ
HJ4JI/kSh43QUPNiEzcDBuN2I9E42wWaNn5Do7JU1IUFRTdPW8B0jR73yvfH7czu
F9lFtNo6ciR3Kw6C20XDhpY8LJgAqEP7Q3CppRIKQVQlmxMPOhSYqsHzfkWffGrs
HMb2HbR2cyaKsduqQ493AN8oDs2yDQJictoZ+4lPJW/4fuWHGxDJpCYAaEmDMSg8
dRhE+OmLPTr2G3Z4J1aZsR/X7UH9JM+Cf6ukNAQ8iG/1n6F0TJNWEjPNEo6TAAeU
Zlp79lM6iq5LiXvzxUqtIUwIUClhezQFnsaH8t38KIeQDft0nZ3VvAslqjVI26ke
558gDS1BDf3YAIRbLyFjf9IxgPBvdlPV4Jt5U/3Eg3RkTZDooP7rlbwvm+Yr/5Iu
JLU5ssoPCjZoIWySkNYMpwm/m2ApvY58gc53zK9V8Pf0asGR5OnpWA2Y4FjffqTS
tHDYkXHK+o4kxgg2EVqZpdffk6FTVuVgm+jF3idXSlOYCeWn1gMJDSizgfM0cBgl
i0RmmdTqHj0anSLPh/qQR7chU6+5P861YdFz1JjZeArpmZKB0eyW3d9W7YpZFfIU
+tdJoFfM/qeJ5Wq0l6SL+fgRXcyCnM5pl6Ytk81bF546EEUET1KYFnG/WUiQQN/A
oxytlnj5MhS4XOcDfMjuZZ6qlJ9p6ZP0y9zheKJx1UuHDQpB4zClZVUw/v4F4QTa
GQi5meVUdaNNexqBNJm0D8k6pa1eCu/9TVSct0i46AkeGhoGA/JcB8D+P6lTTkSU
bxpN2kUeSrnA8+RC4lr3ILrS3dQ2ibPhRqZjQvplvtG2lkcjuwluon1+OyHLv++9
3PdAZFpNNJ9+ykcBZxCSrgBEFjdzrXA1fSVFpB41uA/JiSTfloPs2QUF2Nw3g525
mboLvQtnhO1TtDz5L8/BlnffNBw4/51k16K1dc1LWz4CeY2nYdaqnVkRBiK4brE4
gvW1dyzwXrhV7uoON18J/fKI2Hl25CNrHyeUmruv/P9hagKLUyOTimX3v01qVFu2
nx911Rk03EABr4H7QgMPEPIyTAWCfDNQ2PIn3OM08EXODDDedOMJiVVbQkg3YY33
t1YWt0JVsxXCmCzYNf4N9AX8ZN4xREgwPE4/QcMj1VZ+oc30g6xliL30+iNheXnm
fs+2NMk6TNXyI5i9P3xPuyGoc1APaYgpnVVLuVMEp66tjuhHx3ZfZMhVR9C0b+Gp
3dnHpwb24chXClq6aMr4/NvkdqHbTs41jiNW4juajBtVxFXhH7XZijVPuT/D6tTS
FbT8jSZkGzuMHcPFegqZ7BEBMNvOU8Es9TYlGljv9IfKI93HttVZhOlk1TLrRwGT
Ch9/NvP+5s2GzNFW13pHoZgFFLwhnFL/ST0sWsNIke8EYn4MKr2IEqLA9qSbXh46
Got/7nvHhoLKXGZ8Qq0krOYQE7TLLyd5zInUSi94HnE1i2aynX9/TF4q/HiD+S/a
NUAXLzMNefWdjv34lXNyoXt5DQqT/mMgj40MpCFysGD7IllhmT0dJDs+XZ+zJ8ea
Yl0eSpunlj7ps3a1t5iadOQBVZDBSVgKHBERSTzL56r7uQlz8whHbSb6JwJ0yyD3
b9hX3omRzp7U+F917BMkvhX9RlQaTQ3wIZRC7o6s0tEYBKb2wwsXzCNJ0boIKtj7
7FgbckfstAty6bQT7CHcU5W6kOW0NzqsM5XnAbWqbWymi33FoHVuCSmIuo4N0mW7
fU5HazfPrWKgrUqujI0gIgmjcMcq0a4KGySjzMaMR8pCvKszn1k6EIVjMIhSPw0i
DMxxWVTsRR/notJxfk9aH6RpxiRlAfr+20PnUoj4lj1iiP0PulGdVIcaAIR7SRvJ
YMCzTwT6Psn7NV19la/Wk1YrG+RpvlnDBEt1DPYYKLCiIKTIhj1/Y4FDRavjPYwc
nzED4iULZEhsdWOxlLv+hxa6/b+x3Q2pPQmfknpLQ1TByokQIywfdJQXpyQUGyef
kacvAYfWAgdpZmAl4OcTRw9GAn/QDJItuDcdPNodP1OIdsL810n90cyQYsjmQzAS
GZu/k6G5T6FplMCzsfoEjn/NhXE/ErITcHp1HsSgpLIXHVR8x/VkQ93ny0UpJfBU
ghbn14oxs0AvafmLi2TJdrKp1/wOy+xLK12mAybkIT80SyRLYAXizHZAKCmjfcQO
2PfobZOlLYpO2BMPM1YCvfzF/KMzi/zEcTETPopeoIDgi4fUUGWp7v81nFtbK4kI
+T4SJQUDEPNiPGBoRjTmw6JCuFzN5pTAYZ5LWQ4KGxvSJE5FtVLnRyL+4K5n3aLD
txNAOqr56ZRHb40EXFh/cu60uiUmMqslLSiYE21StJqIwdBx6DPHZ9wA5FhRtU+z
MyusJ3/Dgw8vcX7WpUtWwHizjrdfaG9+hCrtvD/MDq3WQpHYwwedDsYCajA/Ne1U
eODOFrQpdbBpViFbe1hM92e2MQv7HwvL5RmEK9fndzN+yVsBZ0PolyT3yncDiz76
yOvxu71LQh9IMek2ZOIwUBjxUu8BRTCPEeFeCvrI0sf5FjBHiGtlwm31W9fgmhf5
Qm0caxkNfBgxCopyePxcmJnyfWlJs2yRAkNCAlXlHZ+mOsNEjfXNLNRcTA0506Ez
1qoBSceu2dRWfg8R/boQSfWwOi+nLBb4x1ofpki2k+i96DeCrcdDnzsgwkSp1DKT
y88QvEhP9hj5ZvjkmliDs87yqdAwqDGH9pNajYHbbVYd8D7lY57IGBaw97coeAxH
iMbtfLvQLLiVrNf4PNXzQFr4LmrVvngN5/mXdGZ4PW7NKM38laJ/1m/pm7IluXZB
YCaFQLkQCfuyX0Qin10v+UxbMH0oE7mnIbtuv4e5K+xFFM/54Rg/Iu1tflZw6Ebh
kSGLmxc486Bxjwhql0UVQDjZ+fF7fNFdUa1qLFKG+8pYBagfsFbuEq3U+pj5BfWL
FVz1mcZs8CF5MXTGFMalu9Qdugn/z91d4W9bS2zz/mI4VzULo/DQvEwUpPAsEY4l
oltAsR6pCQ0JsExSs0OSZySIpsM8LPbLK3eJyNJazrbJzlP4nEX1LMW7YDI7ZF0r
OYaNOiXgjjMCxjG3F6OWykrbi4byuMdm1m5jyS1mGbSeuYFoW7Iz0Q5XK5Hp5+k6
WeHIan6AgIuAMlGUZXhnlo07JHcG8TQmPsurag+Az47yF5NS1kwMIfi+xg0/1aGN
unwdoRi5cKcFICIab9koQ5G9kyZfZ4Tu8VQSl7GpacDmrZWOdCc2W1yl+f0IFbZs
id95LDwgZiAi03bBYSJYosb0rBwqIAX4yQ3rBVKmI0zTIsTeeyIMnGY6wPt77eSz
wZXBDf0W3Vnki9lVEoKnok47TDuHbez3OrNJqoSKpm2xlknyExijNh/pkcOJJP+j
`protect END_PROTECTED
