`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
S0hJJigsp8LwhExvDiuCeuBwxT/ivwYF7xPynRBVARapop4Rvber1oEXQkiiu7jd
H+h2+bZzMUgDiMsFhT1RKhPg0KgeC217nMhctF9tFPbtovcIVQ3waaTbY1KVWsls
buCkB0BFllfFnRFAg0wbgukMW5aVDuMs0c7eu35+mcPyxbatrn8tbFPwfKizC7Xn
fsqzX0yvwrGTTzk2V/iInUOWSCp1lQkacDLr2a1MP9GWpNtdBKfw8pEnsOmiFD77
777ypmJey8y590GTNGA784+jrFbB2cWyEAwHFpm/1qNaTwVh/ar1uplT+L/080iM
ik/xRnvwPyLaKczAsj+YWMM21ojxVBhkud70uWWC4Eh4sN8AVzkjhV2OF9pPvi9U
SjBK82uAwyhiWHy7s1aucSFspRSMsqfovXn97UAg7PU8EOBoQDvIxKrpfRUEOHeC
/eot9oA5+ZN9hY6b2nmNExCDvlD6DSwJxe5Ree4o+p4IsQ1hHL5DFJ2hDnhnQsuy
w1P6Fe6B8mMR8uXAROPGoLJ4T1htHG6S0wbFHdiBBxfzSFoCc4VvSLKnkaEKu5gI
j8lduIo20PqLPuVcnqYIwRAVwo3kJ7BsSq2M1dQdQRdr250QTPZy/TLuJJA0k9jy
Phi3ISZf40B0ume/1J7L9m5mlWaIITVLBTFrgx+JIntmIduAMjgTq3s2xgobNyFq
iWVhohx0wGBZzMtijsoqH8jBLONPIyHoP5+iT63sxYVVfnlnoeSVrEnhY/f72Q5D
2YZMIp0a7fvoBwwjoRl9gHpDUL/OI0/4DnUV6N/z9z6+kn9nPGFhcHG4C4P3dCMe
JvI14e32y3pmBK552Z6rgByS4V5QoLjkdOETJ4ATLkvOue3Wy31BLkaeV4feoMSN
NeVziT+M7D9q1CUCB+QReclzDX3ULcoARH9mztzwAAh+CcHD8JaNvhn4PYHrf+7R
itJKCGVpvSs9V3caUAi0xZOqVkK4ql91sbN4FtmPCiQ6m/fZPkUAbd6p13XzWR+/
wUckuBjo519RJqz4eFzidUugDjdeH9t1fEJP6hkqrChVARp9hqWtqQxkOe5fuDqL
4eZFi+2gEmDXhWPLIctcVvmch/cTIK71NQmsXcz1D8YmWvQj/o1Aq24MqBAZnfVI
4QMA1t4YrXrARNDfioQF9/1MaP0mnptz+w74E4eQa1NJUpuO/rNOzZ+KZqe4HuPn
FdqlFsiTf+kyX4xCuiS5stkqwL0SC5nkzMS36SJIFJxlJ4xazCt2Iw6GYk27YcFZ
7KTMWZwjZ6LwMKmubu5b+pHFewOU4ZlVbyMaSv+vENNolV4zfYUxrZg/4C6QUOb1
Ze9DKqM4qGYPSFEt4zM3F20aBaiZbp05ueL8rrQFZyvr6tEeQu9wPuNFTNvtlgWU
r8swz0LWU3zHNc/CLBsqVd6K/HSG9TOviWeSBtj7vVzErJjCerFEdUq5KoK1E3SM
JsxxOd6XRBrZFDH8MAbPWEhW/KUhSrnDaJ1kOvPYOsXF45j86iUheFHUM1TV04ex
cuhvw56okY5d5oVyHe1VhFPALIN5XuZ45aErmFcgceVb0pwvdks+wr3vutvdLUb7
qYi/0TabiaxBc3alCRhfjFcspw83S95mcD1ZOtFGp8jmCnObcbGrFMLE5y4+RAON
7qmciWTuTQbiBtQbDgCYt9aRvXRAho8mQHR4RI4c9rYAX2yUFqqGoiO3yMvT9Yax
fTlHv7iaHLthGqflbtz+fPM/4HM4N11xg/DpdaBTUPCpK1wr9PgPdRP9zhsPiiMk
WCAHALHsIG8KGaRaLQwSh5POnlfWCoziFdjSv98VzE5Oh7bDURVMPPA6Eqyd4Zyh
`protect END_PROTECTED
