`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NQjYUfBo1fMsxIbOnO+sYzAeRcIwMkEXkX+sfNQY4St/VlZaRPgHP9Y/la68tSO6
mgNdLDbp/z4MMFVub8r+LEw+zU492JNFCDcHkP9tEV2zO42erU0LZ2WkqNTAmO4u
8i6nTDhyJQqrpnVymIuZ3BrLTS/wlScK9g3PheTV6LoVC9vIJ7kqtGeAcxaEOiJA
NgVtkVyPAwR2LlyMer0OLgrjJPlaPeGnnjEIUP6JwgJ3NxtnWsA5zEhJceBmblCj
GytvWBRtuARG2RHraTwF0y1tY3LEoHDxvtfg9idoEA3UR/uIpceNySpD7f8m5FTN
+isFLDYvuNntJHiMEfDWPysqWGNzu9btMo9OkUX+dCNUC9UHm8889ku6PSQPPDmT
kid/yH7JkyRSn+KJcOsRPCUxKB0wnDjkUfbNn5yJT5zrJsk1SrH/81vvxNqd8o++
B7lXYwLzd1X2ACcwNKjkRZnvgFcSOGriCzrxNJ2M7HC1+P4aV7bADDptQ8FqwOom
+omg/duaI3j1oTNnVMF5GUzqRpOtkjdqsTLs8vc/2sXm1uA/2F6SSO4X/A6NjeDj
TOhAmZppa9eNye7RhQhupbsFjgjkcFasFjx/ej6OcTaT8i/GronZSSxEPGx5Eyij
SqYFYkKeVy2oZykSH3Y3U04gydQ3+h0i1ZvPs1flBsoR1gELysPQr3x11UB5JEIl
iGICE6wMHOD7FBJZxSDl0VF7/2Wov7/8HUJsDzy9/1vzikJveWxBRA5Q/rjuOFaE
9dZngIps1RBnH2d/fBYjlBj+XMyAFH5SDDZrhb1leSD6hCCuLjW/++oITdSs+jEn
AH6Z3uguioA3oWL8+6rPghtBTvFkmHWHZVbpr2bDhbBNMkCr7blS+TTWnOmoUwCj
oCQbUZB8gLyjU5uLL3jEIjDqwQ44n5mAprFDHoubC11CiYO+Dre+N1phHun26sjJ
Sp6ufZ2j1fHbvRlQNLTUFyAXVFf3+SRR46/X82NFD7YwDrfVyWbQRpaT38/b9J/o
STpVDDyTOqhCkBTc+JZ024fRelcvKYfeAmLZ9dfsSdCoG3DHNlbV/5bPApsq9FdM
YluW81Unvrw1DIXeSgd4F4Vb5O3Hm4MDGm5ZMKeFsD3suoy0JArX37NavTs1jR+L
NUqr1tzH5ev9r0ViGeQPjkhdvyooN+qliaNSkSdNzFXv42TWJVxUSXU/rOLknZPK
hERzZGec9jAcYa7KTERDruYvy5N44yCmeYAgJ4+9txRv169Ual16dlV+6tJp/JXW
3q8NWapzpENyIdQ8EdL5ps0x9V+p//SiUMD/2FeYRpH5WTxjivBDvO7YqAJGLL7U
7K6qd7ypqwSSpn1zvVcKd8gWXx5GsHsfQW2/llRO5A8Zc3+mIAgIVmyUAOKrM+S5
U912YsxG1DPtxoGavyxZwsTcPImhOv2GAXJlbFK2fz5rmmFqGKEtOfak3oM+1zUs
QpyZnf3eiJbaVuvYgp3Zi9gZU8R3hTRbUfB2uQeY8/OJ504TCIWMLIn2kUB7HSnk
E2/wCuAmUfWHKAs4pl7o0HkR6WblRfAOek+BSfb1L4y78XvWSAtLK++OWdker8va
gv1OshopThunO5t7ow2QcvQbnMYKNDklrWdmOUudmafYvXkfvCjdlzRo+vmZWlaI
Y+GD/ry1nJRStA4U503JlWuQbYvaIKrl/KzIeNKDIj9C4NIFM5EPJcVVZfL1wKWj
qqWeO48pOXlEUU0d67GXb94JWedWFWIXzJZXkIz+dhJ0WxAREdqeHzID7LYdyiYN
WutxnZZZ/BO5swt8OIxilZFDvs5juiZUgmGkJktqnGfBszLIQ6i2U7KsdTCSzWIH
`protect END_PROTECTED
