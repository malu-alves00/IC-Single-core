`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Jm6XA13BaN0mC4x1OLnqWdW0IvCiPBcmKjbKD/96E0VBPt9nA+E41XcnGgdcl1QC
fvuDJx0mK5T6VIPMXNNLuePvotceGnUEBd+o0VMD8Ov9rCYhruAf5CillJ+jHGiN
3Qr6QoBJ9hbb7jBcYFNFDP9TqNixZqKroC5+qlMVJpktOM8MIFmE2EuhQkV3jy6E
7jh1WD4lXdKpQWPxlizQ22Qz3hOMx8bFmWWkwuNVZO4WIVRaMkqt2b2Em5n+iYv1
RJ6GrzZ9XOJO8OlKfImLkZ+os4Rwc3DwGktCx1qp2K+MzD7uGEzCd7m5gwKkAnTM
dZTxEngpLPuQlzWU+WbZsLdd0+FQMx0yXORNMA7bnvxE0vCXcYAY8bgs5KKsBXfO
sX5r7aLXjIYqKHP46I6q9U9H1esQDA+weXNHTfO5dESV+zuZfcyKSItkaPJ8PC/v
zUGJzPWtu2d4MsJ19BdQxpGPFrrB+jL+4sxuPUrFjCGsQnjNC41+pW//1s/xZ584
dmJ4eT8qAFqLEgI3B7E06Jx9CQQXVXBA1la+2551afEEgvkiAeVsp1UsDSxpAZDg
+N3JOMZmxvEDB/Lj6ywIzibvgvNyRPUB8sred/wdBDG5BkwZ1JOf8V2Fb2naK+an
VmWWh54bIlrGfM3A7N6jiazwtKYSut9zum4yDFP7jppbcnXs0eGrVW9BTMpx4xvk
gyTHHtIVW9PjYZ03bZwynf4dQ5Qvsvk08X1rHcoG8z1xKv+oABjRodF0yyUcaYmC
eF1FpycFzkADApFRnnn8AlpOpy8rByg0gR5A4vfr/AYYkkh+cO6LbvKp4Iyr+mjD
MSYUCqqjh2VnHY99vJWA5VyD9zJSTY89uVBHfA7W3Fp1kDPRgwggHmtb9g6D0l/F
p3/kCL8gW9st0QWH9AZ9xOm7mtfaUvD26QmpKnafa5zS3nMaLPRkOjeaA0vzs90A
bLC5Bwx992hNSgHUbqrtJGnG07HUAMyQ6nNc6d6NlRRw5h6X0N9XAbGKY62yV6RJ
Agn8UGbBcggCgdDohq1LIikRk2Yt2ZJnJFYAfvt5JrJhYEvtpGoMKI8K6Q2UX9iz
OdNipcQg8HuCSJv1QA8fd8WKBIkCWbRN/cLCSrx8lvzMqufDjk9QIeDWN4jeTIC0
`protect END_PROTECTED
