`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GePlKwGTCOp1n7RM33f3+wxpLEven3aFC+xYUAywAYtPRVZ2gYfGGX1Id6qTjW/l
5X2lW+cOUpPl6hlotK0TDjN1p5M+h/JVj2lplfvon/Ep2yAuFuIMFoueU/lcEy8N
TwwFwWBBvKQ2H3zRr3orFUXwCXKLnty/uz/e6V20WLMIZkRWOpO/PiafyoYDx2U7
nThrNF7vNsKev8MmiurzStElYMkoAiaHLQdEjh560NQBEP1uJvOy0ymZiVxRB6bv
yWDg1Cui8o2XhyPnUj9k0RWVZ3UFL0+5HnBSEOsi50TDemCwJlurAN1iqLZf5n1X
jUKh9p3MccEGwv0y0u2rZR0gIUlb48znCqevJOlFLGt09IRpPTuMFAQyWjVXOrFM
Umcep6HnqVjoUxGgsha3/a+AmGtfXauj+qLUSWI/jd256ov/3q0UQAhDd1OTvtNZ
6swmwcfLv+yZgsqVe3e/gIt68EAd/VQpPngbiy+TdD4SoVp11dLMe2WHbIFgAvHA
zfouM+T+gjvM5/LEzS9H4ySiThrGu/EYyIJzkVeF8lbidRm62wDgzyHI6qoZroqk
qiLuh+PRKRYFsy6T25TpB0n4AeBeOq5PUsa+39YmtYyOcXcq1e7dVx95fnRUVNpz
c5/GwlXI6C+Eowg9nN8zP6yPCokO+xsR3g8D5J/Z/5koBt9BIcJiv5bp1slvYwrJ
skefQLJCzKC0ook4RxFoGgPOGKiYPP5I++LCeNqLXxs4m7sAL2bSgoFuMI0C8eeb
M4XFK5XGtkjJFwh+IvJsDDS365uIt53z0jvU2YPaBGkynR2KKMCBA7a+hF1icipN
e4BjfWZnG0xYLoVdmfkg0dFLkbvoQu60XZvXJaw9MJ1U89WJy3dl2Ui3rrYAHitY
Yg4V5/s1LDpIfYvhkhl8G9eh6lbJWLatrTwO7EaQeOg9h1sHDfnCTwJSwDKjn/b9
Mj3hRK6U8UwtUQbLzSpmz9igqNz5+fOCb7qik5wn0YbAoa+4ch6tx6sdiPXrnK+F
cAI5alxIIaT3LJJc/NHphs3IPfk7qxkuqVgf1wA0ZhcuqBy6bpxlh2tOA8keYfAH
m95LZNNZ/DSiXja+PY1JDcdGxhmZZ10p74ezcidVugF+yVDsOudl/tA5QLI7+h3N
xcDpNcD5qwWZLB9gxeh4lmU52um44A3da0jVbIwr9WadDEjMqVw4sdJrPcuFgS4K
Pz4za5UAEzt7HrYsCjcBlH6klM+YaQRDC/b/vi/F9kIUHs5KWLe402tAeB65vRgh
EKtqoLCIZyfrOvxAXqaqcg5B9YEqE0Ypwszb3d0fi671buOoZ8Ov6ZS6w1S/Tt5j
6HfqAdRLPDYXL3Wf5NuyIks7WpJJuuFxxlj5v1Ojd2djyE/NQY5xYnuIqf3F1TvW
sh5FQqgDVNXuwuuxZYNXjzuyE4Mgxll8JbCFE+h8rsccR+dXy+lk1Zc7SkUHO9Dl
9VX9hFI+xO6+siNsCkpFpPABALI+MEK5iSca4p5ADs1mgHBYHB021AgdyGjyZkTD
Dzr+MtJ4uJCyhp8JVbyBDxz3vc5mzSjzzz9u7W7/4m8esTa5UKhV3kh1QfxrxyFV
/oCV+6gKAr8pOvoIs47mgMVhOpXObl1/LN27mFy+UVcXKGI7C9sGHJN24Al1Szvz
U8EcMyl1V+PQiIhfJo1eL/pOvm8gLFUmTFYwUkHh+n5MZymrifPDL7QxqoBWneXg
CpnEssswybddqS0fyDCbx54gXF4oUNom7mDqRY4ZDRZBABq5kuOjFphUR5nu5g7D
pkWr99HeHWtALDIg+I+6L3NikBqyAe9bKJBsXIXCOSjBmPQnuAsdO9kB8uvLEtG+
abBoT64gs++AOsJReJQHopdlzetBFL7ngSfd2hvhb54hnOpvMgaSC7pTxO96+HgN
/RT4/k8S4lXcK5Ak0L0YqZyFcuVMI3OZZpIcsdpfScEpdtKpzLtzGm+hLIgZ5N8L
qQhGbnVbG9ggkh24IPTgcSOKP2hGvVpSNPaWYcnSK9nczQ1kYor8s24s6CBbpyrs
Rp+KjLRkzEsUWV2KYfAphXJ0CtTMSrc88V84EdmCGO9c7pc96KKvMKbs0mDjRBp8
vxOKltkys2ovhLBXp3cTggfXFyaRkbFkA9gTJn9a0To9mc/lTQhFbANhIXF0EV/y
yI2/cPIa4yIXVazFwcauCZL2mXMWrTYQsOKlnQ17CL0bwjbsMYYPRaajd2myoWO3
GcFnTF9pjIerqssZ4wj2GKD0ds1IVtySmzK7I5X3uGxnxvtpcSnBSvYGFZCb9RlF
B1Am/SCq2RYgfBtsOC0MyjjMEoDOJmBYDnwLb7IkP5MAi8+duNJ7R+KC3BZZZg/O
EWWhYiOj0VcKgKb8FkALv54L000dy7dG2ELnyBggH6PglZa0RsixILboSgFir075
gezBNhu4JUAsoqd7j7rTkhpKHcdjTvLUw10IlTQtHIX9SH8hEtbJanfZgooO3VBo
mgTPWi5xgkIXLh0NjkE2LLWAnU42ZRavsYZXOGz1M2geq02e47wKWbhHD2aNjUpj
/OveGYf/UKCSlv3ZEU1Jc6f+YUHG/3fIHqHvWy8XcXxlH+HaKN2jcISzdZpceiHE
65eQZOYph8M05RwfQwwFPhHp6gqKqxWcHxKnOKmshkOXJv+xrpEKlYbflKpC6rrX
`protect END_PROTECTED
