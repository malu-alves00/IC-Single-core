`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
D+9bzHuXToJISUh/0VsjDiPA77Sz81lK0Koum/QLEKo44eisP/sPvDSed/SFDtLc
HXbgn/mBuv8PB3cGtOaVQk7pAGx5zxO40KktHjRMQQ2+9Lbg/zY2Jx9+7KtZwDPm
FTw2kNtarRNH3ZIIO6Z3J1+GdPX1VCMFL/wt09dQlHZLBPzf5KZFPwhBLumETDE5
mrrafPuLyJ5o4CbCfNRTvtX933S2ei0bmSmLMGsgPPN2uZ8ZgLIxfdi2Qwijm9Yi
MyhaHNBSFNL3gMLMwhnGQWoiK513xi/EmhVGXsatdnujUfKn8olfhAHnfs6ZxRE7
/bI7+6nmwh2fziF2eSo0j8S4FW/+cCFb7rBx402TPa/Jj5zeguKnC6ffu4EVjNSt
tqGbbqOpjcIx4xjMXbpk8znGO0Y/RxfMEnMcPI6RpFHz7zlw56akdl2dw6KSTi9q
ruIZ87APMkY5jG1lTry9C2pWK2fgDwSdnof7yX1XpvfLgdT4Fh3O6vL7+bIDaZ5Z
wYbF5/J3aZjcwIzQTWaXR1xlZ72wOIYOSBL0IbeD2g5gy//332lJwopcTrADfIQV
XimyoYwZktmruejPgXbljtqtFmTLc2xmFBhZNrEewMj96Vx4wisDOojAiElpxIPG
/+3zY3WAafQ56JwhjTidRA==
`protect END_PROTECTED
