`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VIOVA8rn+EXnZGkycm8Jsum20QdJjaJMY7wV7Md0DbXAXnb3cm2dMui1QXvCMvRN
0WxBz34KXtLnCGSCwGTesB/F+OCmy72c38nC7Yxbl5igSm8bp68RcyMMor41OVQP
AMvh7JLzGHH1zALdSGRAhODmkF9WZjYpJXJTvas6LXhfHA7/V5CoRxqVXmH7Y1Me
BanNCYn7MULrXUYWgtf5z1JIe8vBgwj2rw2IISSTL2i2TR3m6nN7xp/+2+4zpfZ4
quCv20G343U+zBFftN5BPa2o2eAn9M/hgnTJnDgMXndJtz/X2EpaOnh77FARCiCl
qlSzzMIhDjrgxUXlTpyMkOGhvD/2gyEy8vYc0tyCRM8dqb8GS8vEr0tmYwWHIzfx
qF5Ce9gd/pELwYLfY+JdTq/n/yRQ8mJtfebWWIwsPHqq559nQUGoZpWjZr8YwyLx
BgTIEOtNQnp5nkv1oHvUdBhqeUFQJzgnT1O3hS5h/wqX+yvCBQW9J9hgk14PxaSQ
CUnoaEl0IsSMCK+AxZbIDaWAk/g08tFsu1xzJqyAGPHyAQbJYlEk/VWzqnjmyvI9
Md4bEgFROhd0+umPiCKjFmN9/I8OtptgkG54rv2szPbLGHSODpR23gGTtaBmQMhg
i1TB7klh12VFZNWOsg0rdBH9vpk8i7wgucXc/azdfGHMa2UEAgXcn9PZp8gvt/8i
uEVO79jJg7GiIEwO4ynfQXgxgcmNXlUXWZTwjq/+V7nBH/7yrEgpnG9QVkbQayXw
tRoYwvSLk8IIWwfmjfne0KU91COeSdJ4+z/AT4toxUcYvKh2We5TWpISr6kkag9n
1wfJc5mgrVKZSQ6fsnf5v6cRkLPpLuwsKS2UDWLOWhyUwz/wNtf+8Kzia8zmsQbK
TPs2hRySaop6RMMFmj0fRgt2sV1k1W3oqVQ0fovAyrQ=
`protect END_PROTECTED
