`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZDLkS/LD/NjSgzuEHxyx7j9y0Tqyg3gH+vL4NOxFaz+WYidYIRxCytmJ58cEYPWl
u8Pna2IsMChPB3fAyBmbFqDNMcm+wWTioTWJkPqvULWfei61PE4GnUNuuUhXB9BX
P70kgt0x8ZZ+1m6IRc9QohBD+HXTastqem4UWeRhXGaCZqknvo6npXrt4ShKzcy+
bCrzpJIxhErvbD76DC8ujLJ6x2LO+K//KZta5h5Ix6LRsAMoQWAE4der+DMmh6v7
bdsqHKWL/D4XH38Q4n0jY+ar9mlJj3IlJDbOQp1LdTK5bv4hWEnGEtz67dW9UgDs
h84HJ3eaaFhtgnAiXvTgmenpCq5gFZ5BM/0oFD9MqHXHoqBV/emuvgQ0rKTgxbjo
dzeTTChz4hp0YVNJiBxs6zQLOJY8nK12iZWDRQxOjeU4cFfo6Wp1YHGFEEVSn1Sg
nKvfbOSaCUTjLyns41M0sh3IAiOxGTIanCKE/hA3/jp/Z3Qb5imr7umsTSgHpmcJ
0ChErGeYu41RZ2XyTaSu3ZrPtOBRcL7b1NM+jN9Nbx7SGGAT7ULbmcI2sLrYEKIU
HNNKPtvEU0U7QQoAR74z917wexZ39IJrlIi12FQCPa7wGcTeYKDR7LHuStrZVhMy
EPqP05A+NsyTuafGVGbXbQ6zOceMm3gryrMftdcOPOLyeZw6/mcjU/LVsH8OiIEb
MSiR9jBh6sgD1yDtiYvMXVMFLa1bWupmydiPEONONoic2rJDgaZ8zaU4Qn371ceB
WqPwuLrJonvQcErJWfRRmjbCruR9moiyuZ3zuVUjdeolThYuxQ9BKnsboZx+0Dfs
aR49hLsDVOMcoWV8dpuCxidJqPlv8M2q//ws2ZWBN5GclhTPEWRGZm3ISlSmvhmE
HM9AQhgwHovaZVUlpHA1u+pEyLNcM8DEY9Lfp+2m/vyuhXerhAXRfiQQQSQO1ud1
WMqHOKY8xjwlA7HwzSwbcNhXhqyuTpAdeFQsDzq7c+M=
`protect END_PROTECTED
