`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zPViQDgs7tsUO+Wvqn/6Jg2kO52N52/MfOzIxj2CUTROE8jnx2obsYwH02PLT6+i
bKdEPKof8lrBftPvhXIWYtefOU1GVB1wqseIji7rXYEv/gRHZY1myp2Qv5llweAc
tB6n4WkRXR0D+wU1jWrtEQmH+spNtHEvLIbewE6hG0UFBpVnQXBDx7rI7t1HrUbU
muqVfdxAPdg2k4FcPqtVpjf3S4OLZdREmOMoirYmyev38m6hWQ43qLVumpOW7ndz
jHl58RgO/LQ+4nWBtmfgRedbJq22zhhD6zKOQX8Z1UN5DBKBl1vjKsREgjcz/k3H
E8RA9+n6lp03IiMf5M6yFUSkCNT4sT/lwnMBNlRiH6aUzyLthFEphZYoPlPManW9
`protect END_PROTECTED
