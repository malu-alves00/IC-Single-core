`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sEjxXn/xHgJVwu2La3JXo23Adv2skoDjcn6HfUKSssY2K1jIGOgmzeRRvgO3LUJS
7q6O62b2YrX9AsaOiknWJBl0/NW3G+LtclvKpe01Dd05ckHg4HfY4D0QQ4z0Kqlo
TlT+3Rz6v090kduKbgNLApaUjm092FjBFJQHZye8bbq4ro1roBM4qOfH69iCyftj
tEFRpwMzcdEDhyLyBrqcFOg21bBizUXk62Wcebi0AdrJHUe4nCszT8lwJOKzXXyM
xXcMfSB2Eg4oTDf8tEUYTbp2OD+aPTY4AEDIFAUrEwZ7o9SHUq9VUaXAk1lif7rf
4nARK2dwmEeinddWHIFrMkVtmwWKPwUjgdoUQfT1o/emR3i5d6vgq7n1e2Qtl4A7
cNpQCDcNPBzQ5dvlIsG4BTEsfVUsyZwl+kXs5sDmyBiuvOEejz5Hu/TOK/5V+QKt
5O0g5rlEMs1i5f1kMeddBJzrRlWCllZXpNfne0prz0mh3EQojg6mYHLECpOyf7wJ
8Y3uGGaTqrymU/KNIl926vLGKKqQC+dxkbnnp603PtQyZPEMRK3w2G+X/V9SLDZO
sr4xzzHPgj8lfZG2oWfZYCVtwTHwoJVuDApmY7xHCpauUBNc6ZaEYTAELRB47zLF
mHyRbCJf70b/vTUBsJCsgf8EPQyoE8ohzVXYi5DsH8pinPdFtylEEKH05a2U4J54
Mo+dHR3BX/aegQvUmh5Ovvn/D8GCRxdRzfxclLcFTi8MbQSCIxt0LJ7fwHk/ptri
DXwLSX77e+aGhqqNIhcd9y/fDrHKOVfL+P78z63Ex36p3H9s1x2qzBxAUa7CwHIM
BrZy8zN3KcrhmgsW5Qoxx7BE3gHNbBy6yNpCSr+EMDcvJMCclihNnynvKZsFXPCt
enCTKejCQBbxDz/Y1IRAPqxBsfRFNKIoa/z5FGIrJXI9c78TBKHEQMdlvNf8TAMG
6wWRtmk1RpCFEkzkXOTzbO3aeJQbZ3adAg+T/uoy6fDm6wV6s/eDXRARFvmxzvlB
Z9ln1JNGpU8oRrEkZt2yxCi4glc8x3JhVx0S2s1flHIWApjpddU/AmCJ+9CxflgM
t1FwxIr5r0TV8vpogzskYd08cBhk8DPqGGq6VZSe9kfdxllU3mhWvSi6Mj4wRl4A
V/DQ9ScPLxbwt+Rgjo0UpZjayLxrKZ8CKGWAocFWX2+E1dPDKIGxcVwcHGNzoYsx
4wIShwnszZHNqd34dk7Vx4m0Uk/xPhxN0NdkiR2zCrfpYtT1Lcue92UMpzhSU/qC
eh//y6QKsTIun+qHXRaQEt0mJOfaBEeroQPZ5uU3f2hYRjK1XGvM7yvQdKuD36sK
fijmiVEWlsZH3qX7SBsAYmuf79O66x519LgQzmZ5nKN2hA0kv6NVhODEelYix7Pu
u1yfNjnRqQTXZ3S4mtEVo0KlNkxa9RGhohG34PGXXocMhnOYzZXyHysZVYu/7qO7
lr8bwNliN7BUehQtonr5BfndI/pELoA9qZzE63WUh89LpOedXkVEDiTy614Y7w06
mlgjosRkC6/nhVh6WLL9l0KOq48lrw4Uk5LQLhgU8b/Kx3aQF9vPYQQfxLmOCLMs
Pt7PUvY10qXUxAIRV0NOAbyFZV6aCJE17Mt1lZhIEjw8o2LftgoDn25ybzb06JEP
A8glifYtSio3rKJXmNEcTH2vWX/ohWH57rrxaS7ZB6XuRC2ZmmWl4gEl5pqd7BD8
nBNIU7ORnn3S+GTm8M6VfweZ/ab8T0Qeatm6uqLTjYRq7GAT5KWRIm7BczdQtkWh
rFI+MDQA6YmcEljpIJqXIy07f0bLUFNDYIKh61Jj9abUMUSlKDtRDb4XlJylqSqn
aFPBlzSZur06U9JTfPgc8eCVJHXC0Du+vkzS/eimGLFOJasKYWNL8qGqzK6DOcgk
XDJDmzYuEg5KO3JvjLqz1j8L8PGvOJDUvylaNxSev5K8fV4gKQ7gjdxPCGLljjY6
j/QXtyVTP0OlivoRDlzbm/p+SQTvZb6dGl2TWLMqdsmimaNqQDpRjnGRI1aNjrTF
547sSZm33bVt1TxsUN+9z16tRvV9W/Lc8aGMEiM3m3v2sjmuRCpTyF9xyN1JqPML
H+xbPTPbRZtH7U9YRXbgT481gmEN6u3oH5JXNblRRWXgunTqCXjY7aKMe4wtwywV
aeT8VsgcVY6qE07gpfubLKikfM4FKZwJiNS9GmziqYtRWQwvsgdS/NzLWYK2K68m
IzD1BfRREROYCwUusZXePvUboXB/8W2Ankm2iRE0W4pe31MQUstpUJINulMI+hmR
jebbpjtTHl2vb2ZFUruyhjQXPZH5BtwLYTXeIGi5UvKgaTgjEgxZg25pu8FH9PCp
i7WfyP/anEtjqRmSwqWQEjKYsVgdtrNOM4RU9nsz40R4TAMU1y+MqPqzZ0MtsjA/
znynlBYqZZ94XIsKqmSPdlhG04GQFb1l4krafUQH/zMQnU+htxp0uSFHPUc5/jc4
nXf70VLjM03QvwwBKApAg0+w7WlhBQvF6h1/pTRrqVi/47cOJcv+tZNLAGAWcEPb
ie81nZrUIXOHBlvt5RwBUJMp+BFA0Jfrv7cs5mARtpRFel0/FCorVoa0iZOImzuW
e3ogTaOvoGuBYqyxs4+sWsm3W6P7ceQtw3TPenL1+TkPul8yBQHHGO+J7A28ti8D
pN01zzUnMvNENRzRQvyLBG79wPuI84E52lG0ggbhwRkqLeOg775WqkHUgXDQpLiA
6mkfUOgPKz+XaSRJLmKswP3vkb2gwzZFsx5M0Br+q07S0j5oFkt94pux1YLDfozg
7VvEAs0ZCHTy3XSEkKju/PCK2NrQz0tlf5GxXBpUcNUO/gmFzLSsXutyeGiF4Z58
mL3pWml0godz00qOW940BAYaSAknJc75PA7YqrlNDWnUtJF00AdGvKceXb57G0jw
72UhiGE3gmgDrpJhxrsqXpmkSDlEC9fqe3pyVw4B0tOV6pT/tZZjAmsAJdCJZVRl
Rneyb2DjRLNhxYjXR1t3Ep2sw9fX2Dg5ajTb839Ab1PX8N/ytZaYvX+jOpSnVSq3
kciTdIOvAX4xy9Qgj4fBH+AbvRjO8Ylfo3WRWNYWr5L3X1EAkZShTzS+wnzWMXiV
0lmq6E2VtuFmEtzjZjUw284CqxKlFuJ4sG6/aLqhmOePPx45BQ8a9eIrEikBERhM
xDmihMs6k+x9Jz7hTMP/RnJd1WD3W5a8Wi9hMF3Py4UqyZaKi6TOkLw/nVNYlrTz
SsA5Wj+LRAL9t389dk04dl4iFdmygWjgQEb69r/A5L86VtUHB123j83cfI70VjuJ
8HMq7jHoezr1OOnXQ7AJCTCLHO0oJT8dHC/Qrb/5cn4Nqg19WuOlpkmxQk/ffjnU
3rH3QUOdr9ShAltMpL9Q87rkW+ZLAgI3FC6nRFp2Wr++IH5uWnOR84qOC8CR2LCo
TkLkL4oWNg5bBruyUm9e2eUqQsDhFfYGnB3A5GA6gGTDqrGfBoMUBSq5InoM2JAd
u+7ti2kmg/s/O/LjR3PT4qQiZH17YYTGeA8ETKTBJDb7GYI3V4lyoVTUeFGQDiB+
wMhaiHWREBNVylnuycYiC+oYZ86xMEaTdMglmDzU0IXr+tz1r4QqhkbH4+vxHxRU
VXI2SIBmePP4AwcYzrP1WCzg9sUk80LzMSWSuvIvH/0R1LRLhH5tpZnPqAViSM4S
Az2xiT1CawFWu7TcdDhxUBKIKNe3tIQfrhhYjU4ShZfoXyM0ddQ0An2KAQe5+TXK
6OM3aC+Y3e4xC15orS0/ksUHfYr/w5jgJwsiwF2cfT5zshFZDxq1vuCotf676dx8
ud9GIiMvIBjpdlpSOtIl7WHOlcPWQRUuXVzDi20HPLzXVry3TPAB0PBxFZjty/8d
zPptPuCnisehaPdTq/ScbIc+VbHzyjOA1nem6ZEp1qyhPCauvm2N8foo1d1KpriO
RS1yqs5GhFf8Ho9NrqeipRw8+qKO9eQCFz686jr/v5+H4z+tKgKewItwwWTKTwyP
AMq67K/BYmo8KPB0HdPWREwiHfwDOsp2mYUvxgbjUaSUkYbkmw51awCwt/Vp1uXf
MlEPc7LjILtaThYdazfR/K59sKWpY1Cao+vGAnIDl5o47slYEXKQd4w2nchmhR8V
S6AzAOLPcJXijLR9BK/VUJMPZN2UNCOD4YLwfvKu7KvJ68s0Q0RfCfvDmCDTjKqn
6k5IeIsOcFXMbedf7DdZEZ0ACMSTE4/o9wn717gop5a62cGTMVx+mRLvR8oXAloi
MOs0v54pYjvoEjQQvcx3WbnK00VYL10Kt6iLyoFlOs6l1Uw3ye05rw3oaAQowR+A
rVwaz92DB/0enTQmDzXn6ZMp/4zf0thXTUwT0m/1FQkB1HxxaNXtAoTa+HKj2QvF
P4gooC+lNEtdm2UBIBc6DiLzG7DjLQVJTCsCpUFg6mKeihEnw612UcPFAqEbSL5Y
9MhSNocPNUNfFyWUc2xfsvxd1+h3B474s8FTBxOgCTHt6k5UCoMFDJ9VZrMqAZD+
AMYvOBBVbdhtz050Fxi8sih624cKtFFIQ232S/I5X70aN2jImZAC9TEqXMlIhZWO
SHTrqYGYpJ0exx0VHrVv37yKPHsxE0e9j8fB23N7PD/QwBlO55i1tHYcTZMAwM1N
xQiB6zZHsowkIcJGsqC6gJd2cl3QhBF1dhO6zsx78JWEw3TyaWn2di9wKNEAqnSR
5wv/iYM1LyPJP6qDvjgjoZ/3RBdw0LhvyFgmXGyMu/tazv5b9ABQ03TJkHN1triz
LHX5PjyhLJLiTzleMQPNTo4PPcU1VTyaVw+ZKxpRfynJLClt/rQiSwPsiRCrfPKr
cpVoNfOtp7m8b3+GbTVyawC+UxZlqx4Yt55rncmVwdbyEI6Lb22fz2Fy1zq9TPsh
/NV0T9jJ+wHqARPZse/nIdBfJQbiJONRqevBG72ew44+KUcRTvyEQblhqkNsSm8a
WA79LKacsL49nsDlw8bBm9qRGdPVlykKbKFwu53n6voHme7mAeyo+5GbW87jbsxw
9ifekpMKFMA1kpd4ButMD7SDKl5IaGDoQfXtQoQQpYRKGnKE+Qk1hWyn1IZoPY0t
ZYcoU48TDQqdVAoik1E19v3CEu+tGfx5PDkcAW/r7H1B+Ufg4WhL5jQXf5exyROB
SNZY1veMOTqfcdnkZd/zvNbE83YyXIeRG3K4X69dAxbnK/56cxolJ5GrxOPsxEGE
I8Ywo8hkET43eLahRnycbSlIrp6hKH1Dt02aivOQjcEy6vS0MeSoxS/UCjVzzDoX
vOG6K+AkhKZybDqkqKpQGiFeauACsFqwvnBl2917IXjTrn3a4AMYIwO6ZiTw8Fec
yXA964BZNCX8vXvRfMBuXaDG7Fn0Z2TOf5jOQhr5EJKXyLvErW8BWMHv9KZohHmO
5ROz7SoBl89l9ss2OQ2kd4KJysHMCAgPHW9sLg2l5+5nIHazNOPM9iSXGYT4b5AA
lAOtduzQKM7QvNerIFApb5FU6VFX4CMmBcUb0z53UVM7/cDTEHhZKLUNvqtugme+
89/X7OVXR4ZcV5Gvm9D1qAOfiwUvvuNKqVBUd6e0OcGAMMsptZGVZVFZ/PDPdJPp
3PZ9R0b5YWycV6lmd65T+t6vw1L18ySg/GEgCF5/HDCCqSR5wBhHd/DbDlwD2iDP
WIaahp9SZHsrHhHMPyr8Yd+mnaEUqa/kYAKBYBQdJsA5Z0QLz/nrHLZ5E2FU867z
AFnn5VpBlfja5o8yMpSUE3GBJTDcuZexfJB+Pr9SIT/HUNAEZqUVh3SHObjFwu2Z
aASHJXXea8bAPRXf7owjk8v48mcHA2lSpHlNqN+ypaUg+9Abr8GO5rggHBkdt4CN
VP2eecQViBdG7zxII4LPwEuUkDzAtwC4H/bUFv8onTIDOs55Tn1ImQkNAWqEbCSZ
EHfMnl8eYU6nka5nQbPvxCezihj0K+Kg22ofHmAKyxYQpWOwkQDz/R6Or6oaJhTF
HPyG+eND+vBS8ynZCTrGrtfUbGWTymvdm+Kp+RkElPVNHBO/WuuCL83p6Hp/8prl
X9Qhr6WwDmHGC0Onm/lnGWoPrwv8WQfm14xDQ6rFk6FeLFqFtS1Uzc/Yf9ckbTe3
Hc7bW/ntW0YnVGxpMLPaVqtCaeVkxreUHvT/wVQwFZPe65NOBID41rPQb8DTIN3x
TP+zjrTPkThGcV7MqGiukIq5PN9O5G80I48syWF7N+JDpeCG+Yw0lU9RWnf8P8T2
OB8xQOrt0Vrak4+063KbeLFhIDKupTbl0COuIqJM7sCVa+DeaYYQ/53x97+UYz9z
1mvI98FeqgXorpwi+BKPi6Kjc044Kp4yucnRnKV6WKtMRLowcM4caYrK8OWF0/S0
MN7//QNi47ZFfUzXPtsXyDdeUjxfgNF1AuafvX5/R391BYjwhgeB2UR0k0EherWR
st0kLE9NUREt49i1bAUQza/SCk62pFuDXPTkoXIW2iBsyXvKhM/2J7ZahUlXHat7
8W/4IoRIbbrKXog3C39Es+EykDZ4nHc/UU8mywmqtHTxwOo74pq9bD+baorEhHaW
SX9l+6Mx7/Ju7NxQgDWdY2D8255dGlyxEzEB6SwXuatB5ZlDD5nOzemODSxmb0rd
nCd3YQlyqVdZiRLHPFt930SaVX90lXCT7kjGD9bOQ/egkEne0vYIAELFZST88I8h
Js3GyvRdcIwIh32gSK7V8oCf4r0onNOBqXNL33x5c/3bkt0V4TpBqM5q3390PYrB
tYupWERooO35CyFnWTgqd5SMKo0YHxV/LpusBHBXJxx4t7eV3tLccOd0nse0ZD6Z
vx25LUbJI5XWSH4ExQvk3gpaXcjsMrP1jE2nBXyg0e4Oh9ciixOdRsFjjTqYL9iz
E3EvKMVzBiz4CfFc3o6Yx4SJFfQK2QghYOSq3SCwJNGSUdH4qdaYLjnsOBor/zdv
Cqxx/hu7uv8qSKF2UAkHYuLmiUpjfYEE32UReoMG5e4PJfDUmeeyVV8AkdULr6bV
kQ/k3GNXsq/r3pD9t85l9G3uqPoQxhZdphPpVk9yh8o3YlYc8rpi7uCaDzNw0oMQ
B7AIVjE7Q+F91FRVfII+hR3rt0YYCID+74u+LjMfZ2Lj3DkHm97kDVE/s3rkoG+Q
5oD3eQNGsmryHzEdqrlSp5IrDmSv0pT8ZGaaWT2ECBUY/1W85OveRPnjN6Wj+PC9
r9lKQLRltk4VSaQgRgP9iyvdLpQ+tQQ1mInZFtnd6H2tIeCrYWPcZniypxDcRHy/
Xp7BTZ/4QwtJWCwA0AT65KlHyrc9RErti352LXb980kbsEkCPag42SOWj+xyeP82
GZgfee273cT7469sGag5z/BhN89UzOHRdAnbFiWJ7tySkCZZ4K8SO91aayhTeVIQ
6W00yqrTmwd4n8ZEsseaxe1+1H5LfNL4nro1t/8TmpydoLPazBheG/vhhRwbYR4b
RLyeL5ZxF75WyQHMpsHLeZVhXFs12Y3k0JKLfKtzlwxV/X7bw1vRas26+oh/pKLX
AjLAzCaDCbdX0GdbwzSy3eZvYh7gz6QTVHy7DjMbLR4lAX2uB4RhMz/SLLXv0bEA
y7d2zdzWiMGyqw5WsrRyyzEoc2RyWUssKdblqQgrMzpty6IDyvwU2rmsBNM2RJdq
PYWuL0IzdOS6kzMv3MZXkk/nqaZDa3oMMfa9xTBIl9DDBvFaeRFUWTOPRPH5FDQj
Y5ZYRp0y33yflg+8gGq1WPkl3hZJuk29H6AoIv2/X9Yws3vLa1UXKkezMtOLhJ1a
3k775+P/TulOeSBcgRPtN6MR23wKVmYsdlsTswPgVBdjGS+jOgQS855EtnIy28fO
q+G1y+pyjuNch90X6GxxbmoPwooB4g30ik0HhmDv55aw+xC8Aun0rpJIL/s4MIti
EGYPDeuR/28+94ymuZdskrWgrY0D9GxKEtGC2FvcyV2X/5Mj0JeCJjjZEW07uJuu
RhJB8xTqmS9fJnFqfLdupp+mmu7U9RGiXDEOIeyyTRtmhITtN38J2yJOZwZKvpq9
JqahDG3fhzzHLJzLrcDzPK8J3zaDegWY+enZf3YkOPQA28CJJOJoHyw4Fj6imQOZ
v8i/8IYh53VF+jysWtJteNNc4bt8FNTxE7lHRQDPyAKfg0w3h2aDp2eKLh4mQkWy
dghNcL8GIa6hspk89/PKpeSuZzbUbZIFBexgch5w0DNk9kKafSUNvV7BRogHwWNb
YArGCTm5M4NRGqxwiwsuaR0bBg2VurAFmYUddfRawltrgtHZiJ0tjlmD04Hqh8gP
cA1NHFlzhgCgAKJicQ52kGJi0sa6m+hSE4cNYnXJpsW297IMv+y7njrt2u9zP/05
5SpQwGVrwWJeTIdT0NXMOHGaHWh/u2mr/diViRGdrlmBZLzmX3kdhm3K6Z82nSn1
669KisYgG31h7zUmy96JXWIaDwex9pKAOLe6YegjbnCsdTVQv7XocXxtkAo91lwO
4k7/fBY3/L5rVMDSyvD190IUTPX/NPye+XsbP+nQTUzZEApzhKk5jwTcSxTOwkwc
qheIuYqQK1Q6tIVNZgVT1Rz90dJx6u7QFiryXD1To6fkmRSv1wVAUT+6v0dpaDgX
HMGc+lgtbELZyCyVTLnNpZbgRrUbeYU6pdkMsWl1bNaexet22aO+MSKAXuhkid90
82IHRKITUBGiobT07WYoPTRX3vjE0bml+GsaB1jXUk0e4xzPhEexsrGT6KckiOvi
L7ZU2HIhJp8clWXR93LoHq63nN18gPVmjMnoWt+R51eQw+GBJmoyG0SA9cN0TL8Q
gOQ3VrNcSBdmNKMylcFMVoimF0JwlqWDdUpzoAoGlsZ/0cOnRQrO3nSutadL0SX4
0whBkxcwv6XYZmtNAER63TSTKVHz5X4fLLnRATqVlXbjbncBY95c55Zz8SMe5qIh
3IpomQRRIxBEKfD1hTk7jZRs4wFWSqCISqGL7xunSudQYMg9CtIvdXe9NOli3lmW
Gc6nWRvX+Ahqi1pCOSkVg/vRuKf3hbyl+AGFbD3G6Wu7FKbMPBXcGoyoDZzstKPd
pzCeVfp8sSoamrDWD4j/OPxNxAlpIRJJ2Unsaib01s0fIUN1UVHW53DV90mdSIB7
DZLR2aaN9Cf0QGk7pLg5EPdxqnVF+sy6OPdNHrBmFgTuYVsieRAk7GX/aeandMPH
BmWm03hT1mhVeoaeFXzJzdpM43nAspPRGjEe2LrMOihS8IAKVh6HYofy59D4TR/5
QSLuNPWdfG95hUCek/cbyYXsWy6TDYoI/Iz/YpLOo/Xc6S48BvBRJ+WJkBDcNwWP
WgfG4arbNgr7CZ4h1fnoUcmwphkCV69OTvgjVaaf3w6y2p3Gp+eupS2Yk49nSNo/
l/10+48GcRSGsR0hE//wE0SpeOE14qBjqj/iTzF5uXCkb6frT0omBTUrcmqGMEGG
ye6WQ6xuKaUZBwRX9PreKp1xqDm/N8yHkOz84KiVVfOUQi214rZSwo5K46dwjixP
NePx8rR+8cluGN+tpu9JRhdX2AwPB5sgH0C/NplXDNd+7wohFlFI6pIbc+L3nNfW
Q6KValpzG0sWFuuKndC+CMLUO+pRiwSQ0mfdFYUssjySJOxuuAhnWEVMUnS6J8vi
U8Zl2W6r/MRLr4s1Zbg1Dz2R04tMpXWeB3IxwoAL8rMaDixLmrLO9jg6YqKo1ySw
GjNtxHwwm90GbrdEwQLvJKSUeYPKcr7/K9i6qd26cA4krY4C0JuF4nj4Oh0nhNqf
YqlzMtXSe5IIA/tDt36BDtBlihUPjPbk75QPR+JfJ8bm1gTKop0gPdoKNml0WqXg
lmIUyOT3QhxQmK6v9UbFyfjF7AaqOWZhySyUwncWQ1PSlbiQebfoKsgRa3KlSI4+
dKlhqJgnLKiqXNDFgHDHe+ILJdrFXE1BWAi8wV1spJPM8dKhFscYnGF1Ui94x5R2
EK3oOByiIq8szcc/j8Sex4kvDpdD2scTdSzziU9z34iJcGvTaXmGY6C8XBOIoJqm
c4jo+ZjfNyPui23kJ0KhbCQ5YVmTrdVMfScPlC39dbwp5GPWxIzx4+zzgAsRglkT
nJuoRJPg2QoSVwBWLSER7PVHW4o4lV2nryd3vBoAqxeQTqDHjXQJE6uM7xaGMeU7
TRijKcNa8lTUN83dgPnaZ9NI5fyQp6M7I01fvpEtuUbjArMD/MyV2zlSmxOoXJR0
bceCDRbISjOvP6iLkQl/gm06w2TKc63U/MOiXRcpe5CgNvlhdB8RlZaO8JjFqZbz
4tNB7CaKxyH+n1SQ4SIM2Gjdnx4yGaNycuxYpa6s3YcAl7qbKtU82FNeQnZmVDH6
NGbG58Jc4Wxq1dRbV6LQ/HgAMkqyWTTXtVCU0fB+kuOaoMYCqRWpTK+5WfzqbXNd
nQu8zrMbe8MpLceId0nJuvqvLsq0F9JqstELpxEoyQQfHPHXjg9EOE2mRR2mUtC3
3++vbDIY2vHtm/8W47Xb2gjCJzq+SXgP46shVDFe9H8VrQc1t23Jr3nuEvc6jid/
B3F0S1vda3O2jYHSOl+yz2No7loPRsnRBj6EAr0PzBT3/YvqLPEwVYYJuhjRkGcf
oTbAi5HdTmlOEm4MnM3b0vcBZ2Y/TcPrYE49REzcE5SkMyzIW82jxRal+ZsBoC6e
KGS87i8wJJv7DCs1C25+dqdmyhtRo8c28WBPnJIh6APVtszGjIPH6BfsaocPdIpv
+1TTfsC96aLD1nBIJ25La8D7NDhYhzF5yuKgZenUtuymIWDkoNGq1ytD1tLcVD3U
yhoznk+NAmDt/YM/f2gRzKQIyoGnRA/cYayyQqhuN4a9SHOTnldQi7qGAOIBcTpM
Tu7tGFxy07CrI9EKih3NPc+e7rqihzva1ushLfIlXZGl1wPLPHn+prBZ/Iuz5Rzw
HLXdSBGHygJ+ENTCqi/2PQ+IL2txfcOn9y+WIIMiVj/ctcc9sTxnGChdxfGfg54k
vF9i7vnJaopkHaPJsG7K0akpPAFCeAWeXgRAmcD7pRl7ZsAaFkmEbzMnVMaxm19a
kse9OnDkFuMprI7Y/8piQHm60k9W7oRM7yJRfUXRa3y6eeA9aRMkGuWt+tPtrwPO
KvbDXJ2WXdNLjGCC9BNv4sLdtgAHMXKPt5ZbhKytJ8/0JyfLIDn/6PhkUxX8dBOO
5vBXsVBUvJJaywqH41OTc9rFswn0gOipsJ0KuVarcmNBUrVhsKXE/M7IV0Kld0uB
s5jXpLRBU8I2SyjWtBw3QeRQzje2HckLdJb1qDgeOJSdNzy4cf+vtUg03eqx5B6E
xATB+tvGhSEHb9xIhfwFAS95VjqJ4VOvONU4kmT3ofesbhq8WpqbFSTrybo+Pb6t
NTXwGbjeSlHDNURmiKsOQyM4wB+K3E3lYEerDBromdewU4wuM1ziSYK0W0c2fup1
CCp4rdn95UTjiWfr4evGUsRUIUomtjHWtXqoaDR8Qr/Y7yrFLPRLkAL04WdtN41e
kzm/aiwR3N4FP5Vs+wvU3cCbeKqTIHFhTQLa66614vRXVP4qgulAIsn/ce149WdY
vmaNFJh0Mo2FqiV7y+tEMntowqWSk0JXk/axFMhmBt4CCsW6z5YSeXiwem6WL5t0
DWQVQEizNBXN9vlIdRc3IClnOXkn9vx5B3Br03nGGdxpgpWEroD6bcX/splyOZgn
DfDEDC4t1rDBt4nGAynQNYEVwg3xoA5gQ/K9wW4IJfFuX/iSlZrmJUQ6y1TIRN97
bGO8bLFEpMYPVB2Uxsv0YBKb5R8h8UjMJ/JzHtn48C9Gu9iVgNW+tW8afkvNHJYz
664gaUE1qKOx8c/aHO4M7cE/ux2pJEBmNQorEnAbb46y2ItvRfx4tXQ9dRjQrCpb
byDqKVIcHHBcjDzSnIkz42W1v/fCBxwA/FGGiHAPWKNe+NO0wjfkO6JZlHc7xsMo
oqWboob6vQtZtX+L7BMdcoufpbdnJJ0qdeqWMLtko+M4Cl2Fdg3lz/YUo4nj6QCV
GdZ2lKV3MLL8sXIagTk4/Bq1pnkrBp6lxYchAN1/1XAJei9ByqmCdj66eVGk9q0q
P7+BNfDk17gs1G+Onjo4N5yK1gn+SBPqULVZMRF2YeyV5R/g2WaJymwLcbBi/Htk
/aMwJcEQilKQbpO1E78Q92x4J0Qinse5Tnkak3QRIiIYpCmVmdCUAJhOHB0oxtt2
d25/DvTHJSTdKSBt2TNUM0BAw7GJWrgmuDwR0FJl5r80vCGbxmV7a1RZniqWuEmR
+V8NGaufiOHX+QdCQCsNY5+9C9x3rHBQ1SyivqLNRna9BOUDvEZsVQv3/52hjOUU
Ef9w9z025rwsbNgZTdQ6UGNM3fFx86+ST3sG6rI8UyybLrPS2kuKBvPOhh+N4bXx
PyhdfL0qEpp0U6bIRDTnWwepxH8x2TzYAzF2JuVutx3fQLYda8JDeslfUN61mRlJ
obaJk5HBMt+IuA+WJLjHp9Wh/n6z6pVu07u4ENCLmkY/5Z+OyzuXxd9o0n0qcyOX
flH2T5GqB5Bol43hyAr1jTY8p2gAn8AmMQLNV0zhH9OYbmull/DjXW5Idp015y/9
RlhL0UEDZUXEMR5qf4lzlaekmiedkmBsTb8IT0x32kWipiCpxlzWagnB6zpnzPYU
Sd0ClfKumGYv4RnDPBlv2rSmBS2FiDZJBXGMxWT7CKulD4OLd4AvPttKd+D2V/B4
aqTTp6ouEV3LqVHMwHRYdS8PgcQ+SEVcBo/t4b/ab2rjRpnlPX06F/oJVTANfmfe
gUlu6xgtCzuA5a2UMHA+Nm1visXi9fL6uDEmP8MnRE+c2IYIIy3pay2O/Q9mK5I2
wqEr1MrVl5G2juUR9dWehrCJ91DnmrC/kHZwWjnjwxwLOi9++Tr6rLBNSBdLoYmM
SysEDHvbwAQsjYyGlYTYU+M6ViPEEXo/kgfxhLQ4pkViEzMP0Ghvi7Q6CIz5v/PY
sDuoKctX1uecPWZfSBefm6L6yEeWcAxnRgCy42jQgv+BARXVYsIQKFlaBz0xvfy3
K+CWDp3gSXW2wTlpxiCN4ftf6a+ICJTeUqiIwSETbHDdFLXCmZvo105g63rFTV7j
z5FFF8K675gaPCttBSepFV8Fc2IPlZsdZVQBs+RumUl9WU+gDBnXQ5lpBDLPF5TP
jGohM6iBjCMfSiwa0ZRgjPsQBdQ7BRvQrgtS4KsJx+7rckEBDqJK0fYZnBrL77vk
3zL+M9E/ck0f/Mnsq2RvIdfxwKSyl2kZf5N/7b1FJgxQyt8htb246xecACJ+lMeH
S9CoUSvB8o2zWOKZ9ayHEROF6bB4lXSRieKj8DEMxavDgo3GgMKjUGxXvcsz9JjP
YvX7B87pS399vfU8FEI7jr9OldbOLChUSbpuyCan+OGqzOy/WizctV8ZunD4qqgT
78KwqzONJTqbIGM/8oB+JDbWRgSu9pKcOzGW2/Xjm47CuAD/Pzdr8FV9kizpIxQl
1THA2RhP6ygwBLfnmNbNV8MsSwAG9vnU6y4B+7V5VqZKKk+Tn9gaKomyRmJ8iVsR
pvNliv/9QRn/DMZPIKaYk8mFAK9DfvZJyHmN3uStaWKqIM2g02D/PvmAThMlYu5J
SjV/VioUjIYo8xhZgo/RsvIqcpUNgrtpFhqKHmvrOcgmAjzglHbmddgmLkRsT+8f
4yEN3YjvxpdLR41WHzx7hduaP2CjD/r+BfLOwULMPaGYnjDZEl1X70fKPDNLFCQ0
NJKzEAGcJ+SwDuUSsoKu3mfoFaa2dhJKHNMI4cAb4Dy+OmwAXy8Vf65HWjdzq8li
/xYO4yJ0NWDYR6pzLvwiSM5odplTD3hSV/nKc8+nC3nHkyiFqcAyY3pDtcczfTnp
m8N9icVFjcAzMw8iWeXGvJP9P08e9SBM1S0MUmfXeghhrvrzMe0GJuoa/HoE5DCA
LG5T/j8emEW7rPwhS+HmcsPhZImgSiL5rI4G+uyejgGKM2sYp9y51+PYTfDCIfvq
Zo2nIAKx2wLvqMAs9en3oT1988N2gby1/3nkEuTg7IYRi4GFY9KClpK4b5ws7DBU
zfxD2Ko8oJm76JMKKY4vsteOMbAtnhOBOco5pe6rMuiO39eei4aV1SXMq6rcDmHH
N5MoBNHTRxpWzqq6q/OkPebwyQIrdhn5byIysa5w50nfzusB7SwlwQo3CI8/5LMf
Na9MqTl+ttJTfL3W6kiIYPcLkM1exOn4hdIw0fP9B6zEMt7Qw78Em7iKywUF7ixm
BibIFuHZJhmWJjcTTHd9R+Ck5rBSchg7OVpk1MBJNw9NWpi487A8SJRPSloIAGpk
WLFw9JeVd+J9i4K8z/7ba9DMkSEShGqrm84UIpKw9Sy/QECIyUpwIUU1dtDAsB9h
kd95ew5KZXiAAcfOAqEAzVI0/C1OgahUE94PE4Lz0wSXo6sy7qRc8EuA5p0VRESX
7zIyDLU4DbWfGaQvAQEuphCfugJjxKClxceOvMs/pQ0XEZBcNJRRT/KK/VxtTUV0
Fagp7kX5ww/gZge+r22hLALQix7J6fY4jASg22QNqV6eWEUuXrDaJl2fCw3CDINJ
XhQio/nuzaJ9HQBT6VnyKp/mbiQrry1eb77hXL6auPWzPQrn9RaDKfch6M7J8vhB
2jRmS7D/Fe54U6/yojsuTL913LfVae38Pi0oAUHCq4dMAnJW3JTkX6YrtuUInqAR
g2ApAhYaKTF6B33pHPMJxJdYpWjRmYjV7c5fhmJpdiZ049/9EIfRQvMrYXk4T+o4
6pWo++zNA0K6SV+syNYxP0iwOr6Ke6P+HE0ph/60gntFVvFnD9+GqUwdtfx6kTZ4
hM4yTwQW7q0PAT4JK0X8Zvz6RV5mFmI0xaRhOhCHOmecUkzQ6+SqrSSX3tdMbMsK
QkHoTNii7LPcxDrVk3CPG6mFny6APfvXwG+YiTjDkKJArY7SHAw0Xb/W8G5tJ1cT
FoOurki6k+zwXiD7XpPqGBl7GpxsdOjxTC2LAsGpI00CiDUY7MIwB1wRqrP+2mfy
8scTNDV2gHhU+zx2+cLLuzwISg8oHOOJXnoePrLs6B9UdV/BWrbYQms2y5jwH0R7
7Xb1WCiFjtgaWbXSQK2FU0JLj0bU3SkUfZL1TecERsySf/hIrXS0gMLIoahmCWPJ
k/6io5XTChvMFmb/zX22H09G14yDqdQG5MsZBCqt/FXK91URjXiBp8XTisW/7psP
p0qcc3NVdYDM/uEQMFhnnuR9XNZfF1zSd4xKgcWB3LE1okAyWGimwisqwtAhhRap
fM3V//+uRE1Z4Tj3s8y/EQGSqoT39jlLBJTSmNfHWTkZU92wbYPTZmlygVeOcZmP
vENV4qUxOAFnA4ATOuSeQneBdjc+0gpMo1V1BfEYQR9dh/LgJTCXRHxLyNF+icH+
GolPPUVEt85CfNa3WwtxAhnp9eBWM3u5Ye2v4q3b1TJFKlpkRAmjzdKYq3Cjjx2e
8Aehncb63AeGd3it3SEQTpVm5n7G7ALtdD80gBQENX2eylFbX5uJGPC3SG5tmoqy
WuqLkyStpv2y87dZZdouO3uPE6YiKg8+x9/v+GO/zZshxU8gGE3vCNzxqouiPWEq
xSJErKWuwVGQpOSUTe/KD2uGZ1npAKqNE0RoU47hmGXi+nGAw6v5SWLk3zMukr0o
rXJMk5DU/Ad/3OjD4Oe9rjXuqLnSXfTBDB89ZpTTe5ux4W9GVk7p6+OwNO/6kJX4
Zg0W+PNilcRutnL/EWCVbHq5xZ4kCDg0OfB8C0uKUJL7f+ec1PCAqk737+w+bHV0
WnI3sXpu44NLBeFltPCjUd38HvnAWk4O4FSRXNG/dPLhOmhnrXDuCBdGPOpn2d8m
6mIhU8q41ay+cKRGGegXfNvLjtCK0E1dVFSuy9lGWcyfooYPIQvr4W85zbXs05uQ
v4bdUvsbqOiM2cWCBTv00nPZUIqP0oTnESS2v7hZHMnAOFyOLfHU3FIBuOnUkcLf
h56xBs6UUmiejIYeld/C1PTew1RehtaWR5mU/VhBQcvtOODuLAhVQh3HBXwzRqPc
bWtdk6KuvXnrFi4xz5B+Y3X7EGDRMf8o34Cabq1xoqESjnsAs3T09TkZjzBdIG8k
yL4aCf4WW2lWQLxsJcrUCTcdNKGbiEKGx7j0fgvNPeEdmlbPQ9hTGQSoB72UzXDu
jXOUFfQRBPZyo3ad8AUydFsEn+QhfK4J/hIMM6LagHk4vk1pLRF4d8Kt3cPai/Li
iYJsvd9IVTs7ctoiJYRzLyl5JwyQ3zaHnBy5fRuwF24ivb2TFymjQaeALeMK3zxe
KsKNbTvOYW1CgxB1aZwRxyoArSzgRBD9oIP9cm1dsTgs6YrK0o/7XUC4KYpctNfp
4SDp/1bJTroKZ64KS7QqcFgsWPqx6VHsEKNVGC92OGgR3zyTIbIVzzWD7oi1MrYx
o97+QhWlpbywhn5jFb1pFcTj20GX811gSdATwKNJWycujsSm/+qPwcCJcAUYSCxd
2HdYQ8vGk7CBm9SIADdrtGzpBKRL+9l9Vqb8zizhWQG/bgWvdDqkU4O6IBbNhTwW
cy7tLHGru7Ys3nmZWEhSR++ENjB85VYcO6adNIU66LI2UgTOQJaIdexcYkFB53UY
ODZIUMZDuMUpmpY9QSUeu80OmX96Hr9EWHCJ5qS4EF1uPhCXY/ZTsggKNCvzbfUs
/RB8R5MnTPPoZK2Qqmf3VYoGp+t1SFj/IJsDMgkDZTFPkliKipbhoF0e2ZZeuhUw
J/phWlPsQd6/V4AjwV5FHMbpM9b5ye0vvm9+z/s6Pconjf7IdzUoPNuAba8p2N8s
tXnTn5tTld6l7G8OlZOdVVZNJ4hNUmw4BVZeLmgVBqYA6qDWGoME7KvlDX69FpXf
VJpqcmUSyyrAcFVqD28rRLHKwVUi7Tnqs3dRi056rmM6XxLHKkDAKqvNQkOVu8U0
xStnDLZGpIz2tKsHnIYsehtceVNehubthTTWX9BtGz2zy1rlfR52Wl38BBPv4cXV
x1h1WeyFLcvZZ8uP7TKSQedMihpH2RMtwnCsiuAel+AMbNRJIy+i+tgczpiKvauo
xk3zniLaWgtUfhchRw9Pc7l+93GgeCXmLLMfzrbb1+n2+Cu3G93LsmOfFvVIK8B5
B1F8VZos8KzJe5/QwXsATvJ5W2OT2jd6coH1SAxfHIdHLMFJrQwQTRZZ5l54zcru
yDUM3vALlwq9091O6aYUeNQeNIY8v5UYjxyEvgw8mM1BEq0kvkjqJtChtsfc2Wq3
FIknDas/O9S8NUo+K93Wc5midSfRLm02VkoxKNgJUAkXVbuoCYSpEMA9wUSqyFar
+3zNIyRSd/DHJ/Y0OFUwmwJ6/3GdGmy/tBfDq4psQTKmQCpkdsinomSqOh59QGCC
KVyN27SNEVPAzQwqZR50l6d6yaXOW+oR4DHB8b8cSLoo7PsE31+jJ9TDABY0HIQ8
HhLEjPDAuHk1tEPvTZihkNziRgn1b8h3Q3uu4e16zwu6qqtA6meP7xL7vw9VRgDw
DkrYdQtCkGi8Iy4yPnzRhRmrQjDUoYRcbzuTJ+kIZNH3Msga/xd6qWhccEXuJmZ5
uJDWv6Y+OtLImr07GLZZHC5pPUqpf8rnps8ZLG3J7ckej7VQVnfoXflz0olsMpiZ
V27fvetU5XqxpoVqM0duc/LF+zKYLcgJxmgymlEx+WKlBpm7nZEbQWr27noMoUFK
P9O4dJ1o6ZRmRN+MS1B2HOU5SSxE47VHchmcfbiRjE7M0jUWisCtgxVta6awwIMz
LoYjCIS0YfUu8mkIxYW3c0CQnTgtRoKs8ho9ZUh7NMc4XpAUYXgj9OMnfzx+EuTk
IcwbFni1FW9xaeNO5LWts0SpMpz+S3XXhJfq/+VmoQGBPsRimyXD73YM952NJsVs
EpgXLOY8FdNTTgp6sX2GOZYv1hRC5G0255Cjy7avyWrQPwqF5byyuJgakZhSs00k
in6/kla+pSzKvfq1PDet1zbMXSS6nxBHQOR1ZC49eiLBUBhJ/0xha/cDKTcpsBgZ
F5V4259+jt5SrJ6hkpSwzNCTb3QUGMVAfS4IoDTk5pjNotnvgBOUmZHmZ/1EZpq6
NoXlP55Yh4wyfFa1zM7lv2+S9/MyccBjcDV2SqryRpP9WOZXRysaIexMcatKRaNc
51kBkOB/dHvGm/bs5BuGXJi246FDks7pxcLnC6WVG5bP24XGSGLySy2gwBNXDUz5
RMqCp0tIGIH6JDpWGV9cqK2TE0VXWtVB3EIy526kPny6pkm+/09Up0h0lLAv/Tsk
ZFJNsmZ1TjrjZmQ9zJS9lL5a9uTYja77v8tWx8HWBVDbO9iXiPHBkSwTNEClqrnu
qUBSKhtsHKaSqYLk1E8EeNgPTPLsrmwmNUiZqn3q1UfZxAFOv35xI7tVmov0dYCA
Wgo9GMR5UC6uL3Ex8cqaITNdY5UsY1m4nxydtGD1cojQqOWOhH8RxV2zNaOtoglJ
IVTUIZK/LBVxFh61fPhcax6q3tyOOPCAIRlZ0loxgwwBoHOXFRKLOSQbdj+s3NmU
8AUXF3RoR2F2VDe2Ip7YxSai+rlSkg6XrTDYdWN+csSU4wVc/9ynMyD+EZl4qDR5
NOqNfmytpGjACR1nVW2gnlzTHhHGw2LePAJR69d+pgU3FsSIH1+vdFRyXY5Op9nH
Diqj3woln3K2fg5tfGRURthHt8HRXFi1YHTfaz2+0J1mfAYFH0zEyZVV3QyDgWqG
Mhd77tD3MPxvL3j/3kHJqAps9pRV2ZZkToXOLEKyPj3g6e0NDNNFHNvT2FNs+NWy
RFAqbMSwAVVTUEwhx33yTPY0srE0bukSHFPsHIbJEoZ7kNOrLbS6kaJr+LBHwkuQ
WlSVS/1xeLVOqNXOavpsk2BAxFRJoP/yn29jlJc2zfN/Awkq9Em2h8HkOVpA6jJ3
KioxC6oqcmZK3vFDkWRNiu8NjZJnjjTwsDunoQ+SaBO8c8ahd06c86RvzW0wqT+Y
EMK/Jc7Py7qXzOjLcn2REc+EUGh7TEVNcGGjFaYgzzd0qe1YFjiMS1tsIQSVR+T8
0Lx7xdjssrJxOYojlLA//xkLSnqFyNe+hiAyREWe4rmysVuEwvPPKl8j/b6AAONG
iksuPnFDrtYgjVYM89YBX1wojk5hSqA8G+4yfCk35quWEnuTZzbeMVf2NZhQ+fMU
5T/Ma8tBDH+4xzvlCnYQEFVyacp4z7/dhsUceQZZe0Jf0l36BOeYPe9b5G33+5Fr
Bpj8EOJ+kqdBO+OJ+/+fXoPZBRiocCbaOetwxEX/QtFiI5TQwR5stSA11Qiy07sJ
sHhVsYw7VKdzhWxySAJtzonrUUDTbvlzDTbYJYjC5dTZqrN6HjPj2+MufnGWwu12
oyYetyHxbGZVRuYoUjH3Siq0ICoD0p03gSLjAI6A9v1Q7aqOgWLadaHCVSBDsOna
hEKSvOwzy2NbK447KY+hgW+QzEgESWkKg5HhDuG4tmN9qxRYvBBxQ21F60UyDqti
BqQCM3bG+VDcnVFdU8x3xk5hJBBPcej72aZ/jwvHTtKKinzZ56PrgJ3nkOiRqB//
YXF47J9ypoTz1RFYQZpL76PuhEOXKWrXqg8SuEglONtXlfPgMsJvnBhRG2eR6Zen
FPnhlX65MISesu0wyXiGiG4CGOqUd3kv0NaFVz/kCB54cJ6UuGrmY2F01/5LUznL
6h1u+72rkvZ1kN/AgAqkUyVQ9+hHcbClP1kc+plL3CZW5WkmE6WGH5h+agohiqOC
//j9Pw6kX81QMRgPRL4/8M3zC2VO0JkBGLLbTYS6FmD73cTv6uUnqcBlYmtOtTWE
ZGAjVyItTLCeovxs8uu9f6uzpWChLf2e8drZJdJCWGvlNNxxsQ2HARsBmZfsbgd+
h9K+ZFRw0E4pzCXejeG8EcXhCnnQjJo2bHFNvgaweooEP47tipHZTqzeHSZWRwNQ
v6cmlSCiruFpIQAd1OwSHgYiQQWGu0z6vksnm3wNWYYZE9L9qFkE7Scvf7LW8xCD
VfZYmfwEBV7fk16jnav3ru4nj5PZB9ZG4sAKxwUYbaWuV591mII9M/xnfke3mFae
6fq5YB9zLK7BFEFcr0Ro1icujxQcePjpDz/GaaAtc+FlXXhKkNF/OGc+hw+ytiMB
LFM6Sr+wKRniHJyKrL6vW00dDV7ygHHnqziOGH/jEmYau/jUdh2WmtwyBlCtk6Jd
ERvM7w7TqeWZ+RsNYs8hTz3jxm+IEUmm17pZypOezPQ0L90sUlVcwbqLsMZgp7+g
0QieoMCjGaZqWSn4fQ7sVZiiMcQ8HU3iDxZ9Mr0Bxlkm0GJe6lwJtpflNFxqLvog
nysdirXnsFOuiL4VZaY35QR8vl7qMbKw3qZTtj2H5pic109lJshRmoJcIcKefJ7s
8dh7IbaCPMLSYB+HSz6R1hhDOK5qnwEMDncOx3/Oe9Bci391QI5W0fkJc4Z8iPen
mr61xZp/XbqZeU0IYm8Q4kP4xqN/HiXIp//AH8E+jM0fNqIDOSeI7S43biY4mCIO
zv9yHFExz1Xjf4vK2NjmFPBHuxBO2qQUUL2lVSGi+5CLbsNTCjP4j5Urpqy3jSTX
qML8i1mQLKYlUZdDPOHhOEzBYsusBRxsjlXR3QEvAuYx/HwtDDJja+0xmGM50aj0
FD1Hekj3EnUADKVQuOmQMVhxqAt/4YM0M/D5z/UKwbf8qJp0mDg2Nhwbd+i8s73T
SrwahgRobz77g+QZ6vF81rfLWwAeac1O42GdnyRETxIsMTmn/zbrKvRT98TXXyrZ
5aPTgzbUIw8x+WzoCMD2KQe6ixjZ9Yfovdm3loZshEP9Wor+MZbttsCdkn/tjg9B
KHYC81rl751rpgJDL+xD55VeFqY2YOtivxGVklbX10lvgFDEr5lpqunG45hL3sHE
OrOfP7b3/xIBUEbtoAahHwDgpQaA7dwTjnTsFiZPSgKGKDQk7yNfRWnxjvqBXYDv
SEDkYnRxH/b8m3C8WQKyAlI3sPVc70WcilZmMwFnBDlgXTY80WJ1YcJbRxrFj75w
MK1wwo1c1rtu479kzZ2saApCt+oOIrX91J1iQr3mV3WoWJ3Drw03RRAflHWyBmAx
pca7RlxqXYHJjrmWpSA/3D5AdSAkJalX/8UBrl0ILNJ02eKFl538yP8YsqtEiuhx
SO2bzwvAzFlKcy4ZfS9tCtrlHX5gl1ZogZKyk8FvwcqDzrsKs2CfrLZ3DqL6F0W0
akJXPG8ctyUlNJ/K2iNYVIfJfdbtVu8cfTqRd7lJQmywSXdL8AK2wTPk7Eeb1f4k
HkRwtOyniv2ugb8z33bwr9NeTCx14aBQAlv7XoaMPZrW9lj0n7yq6yTdODrSXFn2
jbnKCn8xmGCt97u1XSnbDnAtzrEvR75MSWyIepQZt9Us/cu0qqbpY7kbxqu0hJx4
8pdPvUlFwQTcKn6UaOggrvuo+o2w3MMyaVZKZYcMfZhak69eibc003BX3ZqAc1TS
SqnoOSy4S/K5dEuKDh9rI0jFd/jrASjRTK0yNHMGAC3exg4x++OmHQOhWhOY9l/3
1GNjLLUPh54WCPlih0SEw9YPWUuNWFJX5GhatSBS3tIpotjJNXe9NFfcotg4CTzr
zo9RnAzOiK0dunMLQ0IC96flnnWsY7l/lFSSNBX+s4KLlqh5lz5ixkkljImKEeFO
0slubLav5GPl0jXiAunhffka0QOTgTbiKbl3epDuatfdDIK5+VqhgY948cbaGhbv
0d5pDrWKbMzbT1lFOjvFXPq1LMDKbswV4ydMtovfxNPvix+OXupI8x46hFej0HX5
hddA7A3VcHlIWXH6qlE3K+Z7Xv/WyEF1Gb/tSJE7vHbVtv0ZMIxmI4+KckWL7dKv
S3OgjgyKhS/vBW2Vez4sRIUlNudiPpoCIaa+Hx2rpgJDwr2KRhc/2sweAElGrbyr
wiqaYuERSTtbJaX32ejxisvaN935ae21p4VuLjEeSa7XcYCoImaSCgfZjlsYSo65
yvJkjGKbByaGSpICFN+4Ja/YATGclEQ8pFKKtzB6nqLsoMYHIaj2bcDDxBEpA3vh
HBAN/u+r8XBurcEflHn3nbr3Zz5wN1YS62ZkmS1nZ0vsH7IKE2+DU5h0WZIJ6/Zz
fu1uJBgTOzHDxzkroV7WppMlkfJ2cOrNbSBas/aiudK7Zkw5KY0xe5ftaHroNCMp
oWemJ7j4HbqaUHPun1L5OjbSqYRSf0bozzRGCvpEbtJZqSSgQ5IHiNvPmsMGqYKN
hYa+hKG9w2RaLmABNpdmMMwjQm3nw1FQti0sHK2+QfPswrSF+JkvWqYYJsFCg6DT
u2sIdFweXW2/JuGgo/yrdklWSxJTVcjqDKSPE2hogDChcm3JUJ+eEuckqx3lWRrf
jh8GTS+tief66L0i4qRHjKsDk220KZcfCy5hoMT6KxdpH2UQtT99Jz1E0N89zPNR
GGaVHtrnjpWIoWi/QvTaFuqS6W9tq9/D9ZCm5bHajER7CdfRlm+2EW8Y7lcMTlEp
dcLBnZfZ95rXopYAnYHhbgLZFLBEeXzV+N885OanpRBZRuEjTJKX0QJtuC1NtiQM
DTnI3nkJKbYSJZwE1kddzHtjQdmNGZrp9ZnmznU+eKoLJN0YjhSRjzHpWijg+8v6
pl1iZl9PNClhVtNEh/SN7VvdfCBfc00NQVw/KGej/KBOPVkZKMJDx7W39lzbr37p
kRzLa/xU+gsOH4CpQWgYdZQ5mgfYDaaxZnJRIUzSX1gkW2swFor3leHIJrvwiaJj
Ix6ZKUjQy27Vfw/l77rfbnWygpsa4c6A3TDF+niVEz5cNFKLq69ZOr/Fyfw4VnRt
wS2mMEVTER5uwJInDAGxy6+zACDsqlMlh7ddr3im/00KO8b9JcHM9n2ewRHCqsrv
gfn870Otps0JoITQ/lEZsOQ7g9oXWjwq20ul+wpx+HRotuFUfDaCrKbZA8KPTDWX
vWPT8TCIUUcK647APBaOjOLqLHBUaP/g7Kx83NJJ8EmjPgOuUKnHr7U6KFkVuI57
bXYOJoXBScjq08Sh2ADY+fhK9vzeGUv2rzVyFNYianY1ntskJCS2RAkLfS7TLcfd
/efKSRkSMI9MMY9dA8KafK632i3xfDDcW171KKdIOWrhMTZ3jO96gA/NgJZ683s9
Dwqk6pL2tbG8bUWNypaIWC7JbKlW8Bm/4gSkyMMP7+sipSl+kylTgzqk7EaKzkZk
NbKWylXTO/E7R8gr/lkmP2djm2pHdzspdpEUZdWHVCH8nAIlPTfa3iADWvqT0DzN
4Qxe5M6Y8Fx6piW/iRS+SeXHYZtBFP/4geMJVJ3PBB+JI0gvbEPYo3PhEu8kx51C
7TAh7ZestdGym2lI8vchtpZBjgbBkc/qkJgKEvbWngaESGOLGNZpcW9N4UOPAClO
xbzE4hTgekQrR7WVkVi/hdWQH2puITjiyh496AJkCADkYWhRGwS2wO8Gpa8PC/G0
nS++dQ4P7Rae/Gbauj3ktwVjEG3KZj3aOnCeGsZ5cAyYK6W7/Xn1NyKsWKwE5Ug4
/YQAEY3y+dxluqL2ZE4SeMEpVPfzj1Ra0wiqpTJ4bSC30KWTb4mVBbLDOOEYXn1u
IHZ1xW9LrZ5YTlum2t7v+z7c7TXfEGnyHjnrGF1IebLUG2/B3Ew+tqgqNInL9L/o
Z/axHpbiTWhGvUw70Dkra8fzMx+IoI0huZ8yQZXOKFEWjPvoar2ysXYfOuFiSkY+
PLm99Hplbh7irYDoN+1GGU8VBa9wiKe/uRQbVluZDuGYQ09vqEZrTiVD9c7hBgf5
Bi3nNhk28/bVEwgkNuUhuejmX2JQFfbHL0psRcFQFhnfNhfViKLYKSOhtHUiqQx1
Mqs28kc1qoTCLj5bRA9gqSaQ8ukapZODemNc0tO9j43czfA6wsjtc2sghq9y//bT
RANWJd+tsMAfcElcKkXXsK8GJt+VldSu2MtKb+AVD68HZdGXh37HZJygCimtvg2X
GCb3tn3UXmNDyPJioAadxSbLbJtI/NTXTmapJcf0JFFxetpbdLIVPh160QRtwNzV
g4XJ6WAcA2uZ0ZV0uPkcfvOZiWAY/kS4l+jt6olu9QsXYv1ipnchXcXMlREekoOh
eD/LgOAesy4CvmVSQZ2022n8g9iBBfB9/MF+Yzh2mMXv0kABvdUfoKUlOr7vUWDx
HCXxmObEuOJc0UfqAc49KWlF6Qk+Mgsv48Ox7DwVvTdHx0EAyWDlzr1AJrncP5bS
nrFZaPvtfWRothzt5PRM6qQDF5IwIbJebuhJSYyPD8mjAYjRtoh+Kpx0ZFSUmPIB
LD28VCSr+bzeYpZ0Ndrtzp1WMycUoCAhse9f4pZ0YpUKanIZb+jzPkQ97FAg2rKa
7S986JitS8eqBc05XOsarJsU9H3TkX5xADHypD81QXEbrsmhAjWyIYEVPEKGw9bf
FsZNWBXgCW3GqnbNWgQxoIar308Q0vk0O6G3+oYUjD8zSSg8NEeKM3Dwg027bIrN
0cMseFttH52wI5ivo6CbCPNpRKBN2/SLhdl4MEEhSW80u+/Ub8KtxXQXR+vO/BI3
1QrSNneiETkDOXasqEcLA4Yg6nHENozrxQkHJIAdJu46sqKZeQ6Gk16eV1x+8Slo
7ookpR1QGJFQKGer78Gg7FOmNajihcgBGdZIXwc9bVDJk8qPF2okT2cz02BJVEFm
S7Hyve6OC2DAt8oyIFffsoB3ZlFO6+LnAsZ2qrtsPKWpMynx2nMdcHHCx9ubPMjw
axg1IXfZJYoKL4KnRCjUTBKfMyuWWeuv2aYPd8DNvXs2a1ib82QxLOcbOBopEPX5
70F9fWConCnEaIA+BxUck+M2t0GZzkqU5JIPlkCQ9MMlyamLeEUTeSVZyKf264Gr
MG6j+D2Rrf7VIrNdfS5bYaWBtju0z2AmqYnNYvB9AQ0r3+YJ/xiwvBd5lcs1icpV
1AAXRpYdjJCVWulSvYNHCz89CKR5QruPmE/23VPhCMnPiBD7uZrKgiKdVQg+452Q
DN3U0JAzZSDMockEWZfqjgYtg2vyDRdQAjD8bIqIX+u+q1H/NOkmq6TQeZfi0Ah0
37gbUylWCniX2kJYtth6eL2RIP7T1g/F3JDPKudUgwfT56HLP52d4eBK767BbTkf
blKgyeKe4d9rUI53IRZsi4qC2aGqHRK6b4m2FgsQ+jYsW+9Ves52us4vqdiorHG1
cVGl6uYUgUh6NiYjQ7RI/796vq0ftfuiyFomVzYHh5lO1GXsuXTIEqnDP25Dl410
5aREV6PK/wHQVmP6pPiDPSKvKSBXc3rSX1iO1r0qaMZPkOhuqudYwSLCuPXWrZ8Q
j9pqsVBc5yX3cE2s87mni9tPnpkHXkkkXpwGx44Y3/o6sbe4hd8FT0NcT1Bi/EA1
GtvoMFRkMSGuYxJdmiJm0gGnXhufR3UDB6EDcExfQP6Yjc+ZDiAoBDENu9Jwun4R
WaJzmJDofSJagk5nX1JWXmiJP4bGthdq/j+IcUVejEs4fQm/wk6a4baO2BykTQzy
JM1P0lSqDwIKQZvy2hWPw6fc7DLzlijXjfwEcMklgcyuST9feVSY002vZbhPc+9U
ndCrl9j2AEiNXF8sJZpw9T3oCRv0rlzRHgoKQ26AKAHgdxwWF10hka+GoJbUaoT8
S9ff39M2dbUlpp/gU+q/xLypRhCiYLbdNtLqUHpBS9JNtO1F8mPYcxRJGYx6grvu
uX4uA2G+TIgJe8bkwAWeLNmlP0PQKvXk+XIAFcuN9eloZFoejcL4pocodVxLadMF
4Jws15X++MXuWsyGsjE3Jilmfanbtt1dBB1guGFPkax/0TS4Y4M8a3m5OzlO6gfT
fgWx5Kax/uM2IRRfMTOP5mui8kalMPdOr4wtA4YGtGBUKbWpTw0skJ2BqlOVs1rG
kiZNu9kdda3YsBE9VzO9ty5YarRxkLO8o8muo0c8gLHID1vEfmBEhFQzk3E2xDmg
lsoXkAIZ6uRtCV67xBTlO6r7VbZVpPSr+h4O6/xmrgPSTFuYn4pICqbkQMWC88LG
L9LfH91D/dAjRfgHboQxkrwnCJfLKRtqD7xj+mUaTLPIFTVWl8z78INHT/4be8cz
iqZKdxUBxU2o5UeD7lMpNeuOu1jMMznBf/rHrMdd1Ghyxc9QIojzlv4aN1v6kqFW
+X2rSglVXTlxMFKmGHABaU8eu+h8BOnDBQTe2LjBGX6jLDy1mpZfcpMc9H6Ljxj/
ERuIcyfxhRY/halagwKN530JQq4SV4/D7OYGhlPpzl/EZ3ryPfHgW21U484MECK5
RXX0kj0iHQ0pk7lvW+sBE96qeStpCeHiNA/GSyDIij9CEv7/tcZ+qqzIP4TJYudf
qA6H04oPSaTYTrfB4FRDpz3ec1uIHV9+kxIxNvP90vKWKDEQXUiCpb18zkQOzFwd
swPIwGH7so4kfoiW3m2C3RSxegkiIqGVYNaoxiwPa/RojK2okt7aFcZZkuSYC3LI
gE0PFD62muvdYBGWBYxOoVR83JthfCq4bR+aaGs3hIiRuwyEbUp1Xpatz202wMBU
Iv4LzmtGHiH4JBzXUwOUDva9gElPrCxUIie4XcCNv33ODvKQUKqtuZpjl9SfqmWT
YZF7H5c1lV4N/Q/FBNjEF4CbP94vHcxLxV2UzRgs9T/cVs2+1a00ueRGjhCQ0Fdi
eejEaJxqSZK85K8OX37oyEWJ2tVV/lBf9ngBIoaLiKz7JkKAq8leR5kjCfciW0dZ
xMpXYe56Ibzy9aFZzS2Pi4zqcuu5xz4ZbUO/55/f1N14FOU5twbVR3K1dDfR9CXD
iPB3kDQ+fW/kowZwPZEWeusYIl5IlF0KcIlUrzp3EYAhc0l6q3BdB2Ls7I/GxGBY
I43P8Vx7xHxw/MR3YE+w5t4S1jFg8xsZVEveuIG7lNwO3XCf2yCxiJur9Zr2M9cZ
11tZjfjMLFo5xQEcShSz/ybJPa8wiTNp9UDcwS+9q5wH17mMseqf54YVw2vNzZh8
ebHZBjCSTwlfvbUw3NWPVIDeweENEGwVCLxO//DAIeS5gDD7LaTWAMxDwJO+GSe1
l/IMUNtLhXjwh1k3noweNjckqHk/x8DGvYzrtWbwOamqeilDIEVPnQC0y2buveda
6aD/TZdMiSlYmU595uPTZ2FBqS47//ThDhTp1OzWVAfztm5yVi/wiNw6OntV8TES
PLNXW1M1dAlrtMB4GvFxl98zTtsqTStchjgvDepln82WvQ2nLUzbrEss+JI0jjZg
KuGBvXT3Z9WVEZfyefgYrHG8XXfebdx0inUbmziBRG6amEz6gi1YGJkcNYyz8Z7n
bbXrsfAPUFG079yA2iynkj0vPLD883LvyBoOmEx+5FMu8PRic45Y1Gkr5L+KI8BC
SkU+sVNCCbW+FDlctrM5TxFyE30SHcHnkP5zfYgAD0mQ6/LbJ8sMf/5nLTYJc3vP
50E+HDoV0WH/zwPlUGgpkp0z9FT1iHt7vFhk0bTjVRSDdVkKPF5UsFV0Lwmld4Aa
Msfc5pbHKvyb7256HmL2DmfV2GFUICGEY8nznyBJyWd5kVqLJI1ETfs3QQAR51SJ
gH0E/cXHGI0wjl86RQhObcYOf1LYyY3DTt+Aa0akXOOX1MHvn6DppDLS8FX9euGf
moabFEge9a43xZlU8qhQok119npSqUme8X+SMcjiHg0VfGE9TkkL8WOVHl4enxf1
hjiplQTMM7Yx7hbF5Cba5xb9K9KtmtzBpVFdUi2Zg5b7laWQ4ad2fOhTRdumFz6x
OdGckiEEVVdwaPPL6hY7lU6tybBi/hLf9VyAB37B/MzYo0WnCxUZtH0GudznW5hL
KPKZVxn67F63diVyVvpWkBB/b2NQn0dGJBz+iLU8EXlrYgShqB8DYcxEFC1NJb2f
PkuOayVQze6iDBxkXumlF6AYKQBuYcPfE2IYza6GwRXPhZD9bMeBHuNvweBstBev
z2eTE/vSkkHMzr2tDtwSIZjWP4ClRf3mRd1TbSriWRy9tkBPwWTiLxSfWSSVC2MH
pjWhHGmItNk2Hkz/GU17dLq1Y2W42Gyb3XQTCSnmBuYJ+wHILo+YQqrqvX77ld1h
Ox+ZjNfRnCDd3JlPtkX1N5WOikNDmzlMdadb2U8qUfcQ+8yhgKocmMcpCE6vos0q
8EsXzkaWOL58pgSysF2rbCu2ejB1ZcWFzwC+QLeeqp5+O3AiBBMbXQkbItIBxv4H
1NJBEjpcE3IqQg51x7v3k8hdV0EYcZSsTGYEk9SX9lUwwRo6m22TruhSDVHSXGZX
muMTTqkdNBOxdQSRANjPyltOdtAztOem7qfhW8MyLmLVyb9sUk8rVeGv+ccKLzXG
trsj3UFDQlDUBA6V2xGNnQAG73AN9fBqhiY6oOrxCDi5Z+yG1d8fdpOEtwRVIqci
HDPZ3vVbkfVSsZIq53CEf2zKMzaqcwguxnHBfH7kp0yoZpamfgJLn4cqRaSOhBr+
wsDGqqPlFmxjF+FaDYsckBCaYlIqGHSnOcvUYkg2vKmbPN5Ix+649VJPlILlndaV
yCuUCF23e2n8Zrv277luV2UL4lgwRNOA8JjBzGfhYPgd4P1/MPdV/NR7fNrdVFMc
Y+XpjYT1Bwt4R8vU4xY+ysqRycljxN1VDoPQWKJDathpIzTtzmyVnUYgRYDrnoqE
WZhJ4j+gK0ubBuQH9NEVGI+/mFq9d8017D1EtuTMfDtMsSZE4i4qxKJ5v+Offygw
lyjQpYLidTatZNhBZltP5V8NQD4F1fdwKlxEF2jYGerpu8211FuI+pTwU6J5FjGC
1OypMukGfPnAY/iaSdHIBBNZSFhcz8h/6f9aqvHIcF09soKGUbd2XKh/v97d5T40
XBgavS8UBRj6QjaQgoZw523/zS+tcm/rjFqePiUtgNeHmpuqSPLTilUIDTOnMaA4
vCo2LvRMlyIpuaBFy3dknMOpRRC+SCmOcToTFgLvo1bw4q8iKMMZC2d5pvSbcF6f
n1zmWHOqajOxv2pH4KlkEPll7Y6nxmuzy6aDAIj6ez0eGw2jJ9iEZuDl9EIN770W
tyfpX7vhywUPr4lB4kXSMx1CoFdz2IiIYFMXjXXmpuFHKklEfl87YPD4rbGw014o
QUNPjlIRjINRC7PKZRo2OQfl2ChXXbpo7WwkAUoie4Ix74nPIkOKg+tpQ4CQGR+q
ZwfIcRS8jqvDM9uJzfMaa6ZsTDyQ85V1oVdf/OuF6hfjaP+nqmVnED4oo6v+v0vv
6kbw/NodaqWhIpo6yCRFQpW6jfSvxpwKBpK+TqLM/4+ugpQQYkZibYz9kYk4G7tk
zyb73DmFOg8VraeWLyWWFru6vtaKkKuz7lrHt+qBY+gFHdS9qDH1aqFgG8zuHyl/
IP2QpmLUwjjyXnbocfL+PvogYp+7kvaf7sYoiHFyVIz6I00GopzglLenvBgqNMwC
ZcuVaX3D9WHE6pYAGmnqDpvarvvzy2yrxwMEu4zcei7F/9DKfsdQ8woaPE49v0X2
M22OU0nceoHNy5s5Rtag361SXNBX2o7iG3wBQZG1P0I1Z1/LFrjt+Av7P9+yFbft
jb5daBqxrMdyMWA430A1Rik+gSkdmDQMVN3Rz5LV3TL+wTGwI/rmJIu3ErlbiRQH
e78GlOUtaTfmNbVqfmo7EsVPIHmLNsRwuKDQCzOa5BdfNDmCsJabse8o3Xm8MoPu
VHFR7anKU73My7XTDVTo+dbzeKS+A3Ugbr4dtMCtyEAg3E7r0U8ZcW6PlCxU+McL
f02AneQyBjEgNmPyC9TWO9fnJvs6wo+xmvM3i/sIrvrHPaVp5wc0tAWhSsc+V8rf
Cp9HGQdNSNgp1u1h6ZFE2CxoX+dtoEI2nULhleNuXM5dhIUcK20/RsUMXqrKa9Tl
pVNx1Udb5yiPr25owdlJlMeKKi4t46pf6Lzf0k7r+yWqQmobMnpwLxD+sU8+HTvb
y3Z0mO+YxATlp1nn9/xT8fyZgr0lOpAoAxdx728Dg9Ns95EKtf0rCJYkEllUWcgk
J1jbVuxhLCWDoxyzxk+BW55qKAWcQBGMOHhPK6FZXyQRGqA7XLsmkjIgk8yRKKQQ
4nZRBxpZHbtn6oQvhodSkDNZ9dkcrx58/9UEAPS9EcmfUJccyBwND2U7nZj0rsPW
0CoAiN9wiHvJCXinMATwf7ianAP5qF72cJQ3+DsAGXXVA3zpzjhv0qNeh1KT2Lsm
wlRbYovL3aU1OcvNprsGceiWUqFYQVJoaR/lTd+84wILLwl/oaPrf/YdCnohRt9i
mmi1NGw5CGxh3hnRSwE7CQCM8NJmz+STJqyZL+7NPphkSGC9ePSOyh7TfCiCrkHg
BKBWCFWdTWYpsWALir6d866hcP+lpRwna1pdKa1cKXxu0qPea9RpieMNRmDqYJwi
S0fNmo58n6SxUidWZDe25uo4zYGIzoBpWcEKZnbWu/0I+FOXrH+9y1zEqQcwo9LK
wKWXgwV7P9/HgtoCP32a4NLxPywBHU31yYxc0+T55oPTnlzdBHgBNs9WunMpY4rj
VejIj7RH9Wgxkk9wivOpF3M3C2lPONlqwq00QjuvcZi6d0Yz1LGvDTUfAv3w7hOD
YyM95VPoNr+NgA2eR6x9JSbO9z+JNUvUDpU+djSqEB6tMaPxvpi8l7s9HafRWKut
XuXdv1CDD3713uhdAQhv+oQrO8Gp+GYlway/P6hll3Zm+Xp91ZS4wLMf6E3D4ZBG
iWYgIU4LkgmPxraEUhUulkpzV/PrErjhVc284E+hJdyQMrybVZXhccpers2uXSR7
fbN1knoQWvFvIcZ6YuuXthlcHaDb3VmGXbkvherS3c6ht89rRIQNzwgmMPCzeqDN
XgGorZZ7nGaR1pQuWiKRZ4wQ+JS9RZpvoSchgXU9FaCDkQGIST9eT2Ebfa6vQd/I
q+0F9FSDf3fRjxbKRa+/Usxh8oQJCcS5fzTIDa9tkRhBPvWLBVVT/UiFkeKWHd5M
6LwxtGE3h/MOuyKLDPj+4LmSZTI59HWHwAlqy4IYkdgPg1Kn5fiPm1aFNrSiR9QB
Kz0DsrqvgD56K6N3JowZNQI0uPHVhq61kl7feljqsAi9mNVgvP/fMM3HQrmPjcbs
qxgka1O5d1Gs1syWXha7x+Sfo4nNGxtAFYE6SPNTUJP6totmXaFzHN/uqdPO5lQ9
c7FNEy25o3XlFZQjDfp4nhWKss0RWfxrhKajhnYJVNbLYu4Dz3czClw+ZAadv+cg
WDzTebMD/MuNFvavNyy5BUHdsMuV3Vil2NjmhXEAOwmvLzaVnXqTJV1UWg9mHIlj
WhzTWoo1WaF4DzafRWYf3BPQ+ShJwhrRGTG1s/qJCDor0ko1fDc6ZLUN/P04YXZs
HGW/mHSmbhWSjzgYLH4PpITqXKTQCf3ZckYvskdJk/LsfSa6rekm534Cb+RLhaH9
K2usUpPx/ztAPo6fXfoZMIajNWKzyZudoFlTxtw52d7QbzilPNcEijDDsQ7abH1N
Vx+TPtZFTh6ML2FnLT7olQEfogmUV76qYXuV1ovrJmvEiS4pLlXr2zNrnc0ZNUJS
YMJ/tWQgleUPy7cOsPPfW1lYniCDyUvVA1UAF7moXgWgHlrva4Op7n++8Ptmgnl/
M6ONTHMFW+w3qOOyGgRZvDl4rFpFVxIu5MZ0nfw6/Gb7PPxO1otJRT+Nq7zHPgy/
3oBkbx3fP8ptIAAcNz2oeG9EFm/zMAiHfg5rPTN+pnV+OfwGy/0O1G4x6YV4k6Rv
Cl17VERe5AYvahZxZ6JhVy0uUYAftNNB+03ufNP4vNPyVaS34hrSe1wQKXFzH7RL
6d9PRPaFXXAidwtdByCPYEZU/mXB2rDvcPQQFwowOzo1X64kNdRWA8gzzGTrkOYC
KU7ASJ66iuoERl4rxTXztTpPsz+mrVScP5ZwVYULlWLOLLR1QUbJoaBt8IUyL8Wv
5bjfKl0pOjh2/VXTmQUeBH81vteUL83Ty4mrOiI+I3DW+sCnri/I674VQjR6Js9s
XgxXYOKnygZuJpJlg5qTgLAe96n0WS/RHXi9hDGy7ByW/kXV++7oyTOxcqqHCdZI
eAcRvSoftZDVDSlR/jrAS+TJ01b70y+89BbUo2XCqCkiRjep5wlKM9u3fXY/tNWC
u6koHkPZnxXoLV+XNEyjLocJiZ29W0Vf+YXwsl+42f/w2okS2y8WYXbDIPB85XI3
SGnx0CDsCWmWOruVWPTWMXGXW02vc3WeH4jSRuJNPcs=
`protect END_PROTECTED
