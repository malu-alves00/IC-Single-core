`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5Dr1Tjj3kF10OafrNV5agTM72Cc64IVqD7vC6diIwnPyCLeID7wIz94823plRau+
wb/iio63UAwFXzuOZYYhKleWvgfLudTBbqRq6wBZa2VEDrEUkl0cKgPjyZgHtJB6
+0SR3Dqn8EuCnIBLy8c+3mP1yyLE9w5Rasnq5pamQM1bhKZt0+pkH0+do/ZiKA8Y
H0k9TAy1Qw6qJwFI/9UO2qOnIo6FU75MA+YlhvRWpfiLq7e8HEaFZPJrgc0EItmr
9aWh2b+H+q1EoDK8D77G1aW/PtJLf8HVreEUTmVXryzAR8eBXWpwAhOoQ3T71K7o
xo/dh8hVW2CjeC5Zx2WhZC14FU7ls5WGjsONaOMBao2M8+0hesDFOxNr1gb1XObm
pZC6nSoTdbGCcCgbj4iPcqgyoID1Cgiqp6WzIaTV/yiyF1cCqaf8RTeraxvx6ZO1
Z146U3E90mveBrPclzpAK5LShLelzh0M3l2UnZRMCWaFBNo1K402s2jAJ2/RIeoH
9C/swgySVEOSMGQPZ9h0mQRQPGeQSwKj1YajxGDCoz6KDI8UDP00JB/JKpjKJv5K
vFXOJ48/uwhmUiO7N6yLo4zW3Rt8s5EOcbKXQeOryEc=
`protect END_PROTECTED
