`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YPw3uG0TEpLymgfrG3SywNOtAAk0IT5NdUx68SL0A1hyG+KQMuV5Z0kDyWUqomMV
nIqJ09PmMQ5/PFPTcRBSgVCn3p6l1DiVgEzwPD4kFMtShd20I8XbZGaNQqVpid3D
Nljfb255HZ/ph4vrNFvfbc17EAL5rUhYApr30X3GGerbWl9Izvdy9R+Q/13aRt4Q
5mPItt6E6RPcVBcMpt1IqLJGANH7Gx4SIq+7y5Kf20+lUIFWOpbWobk6GlDWX+G9
P5z9ydIcmXuZU8eVBuGdJ8L0U4hmMuby1jnAfYtgLl0fjXkbRoiexQuGC6Ox9yW5
G3i+7YPIGHnO//jtpVeTEz6rD+JvpCXicNGy1Zyc27YLEFUba0aOfWGoUuD1bOJS
5zBoBi/4lk/XRaAM+Tkd7KpGus5rMhj/5VURNWjCz0W6Wy4C7N2qhNCpYOAdZsZt
pajVULS7JRDTCzxTofI+d406tcV9iHBEoJ5TVXUKVpwhVBfo21/X8VjCLDHGmo/n
FzYted3KluXtVoeBNz4nTiyTGzlyQezN9p+Nom+djU+EkNrinSRaSN9EZjpQULTF
kxQU2QpDRV7REN9VyEwKA8zKNS9BY0mAkfWYEGuDW4RnrrFhXKbqaXN/e99G7TV1
44USpmsCcQcgXMredaQIkam7PcZQVFDWGcZS61nXYTHYiegXuel76ptrhyUto2md
E2i9fXTDb7VsaHkd4QVkVOq0gXs5jywb/1M4Z0BQ+ElMof+1/5ME/aopwsRzFbRW
E8fhZqXtwZ7niQor5hF4TfmlG8AuHY6xCKIzYwqkCr8Y9Ytp/ko49CB142LC3QLF
bOiuh2sOCptxRiNU9jxoQpbO7GcS4lCr3wpbW/zNoIlhiJaTwwQIKpcQ6cfx/eN+
+RBPZ4vfi+4Xx9DF8eUM9ONqkGVqdexE7pnAHXo6KzI5IlwTb9hQ/M93seMe9I5c
MqHbxL20apfSLMLzRsNFB+e/czbN8b867eb3GiKYkdgnSjJS3Fn8h5vxCCfbOwaw
av2N+07PCZwfWlkkTnCqvaNCKmHEp/RwChLs/lQ/ftLZnd6+BVBjja9Z6eoEG1vn
V6QfEsY/eUnGIaE4VgvDa7tpWUbiKM0ayc63E6n35JM=
`protect END_PROTECTED
