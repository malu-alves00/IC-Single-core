`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8eLjPwazfHbjwJJyk1y7qqKLE7bPdRcqJjlZVqhcLIKHgSh6qzUigVHJ6l8TQbra
G38mhIlcFyGowQP/tg+gAcnIdBcGmPfb2uk2yGLm1moZJExT7P3/r4j/8khJ4xJ2
D6+G/tBrFO8xnJ7FO3bRY2aVeN6JAO2ZfsUvO46m/ok75YXJDzajMiIhR5L3RuyL
Di78UlQ0hUc90fnKCAjZ9+fTJW7qpiszVq31HCSbiOijGQjiW9dZ0wf+tCmu5rX4
sUDvbVL6wJDL3vpqMnVYC/Vr0vxXkJSJxLkShmlU6yI41Nm3DOB0Bxrjz1dUYciN
Bze6wXptK0b+ZnXJciIhYiQG4nPKyPFiiqfmCASHqbSSvNbw01dBUC8cciEZV5nX
aDlyBFfDhIihC+vqNDnYALt4xnBCDItajMQkh1TjAlbJI92juOxtL2OqXagdarLW
`protect END_PROTECTED
