`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DcoTMATs6WyrZxEw/9hvmcw4INqpf+U3MIY84tQa6DilOfd/u0YA+CqB8vlWrpZZ
msLpYpkxnBbFxVO5+gFOr1uHEBBXdTqZaBWUomruxNFxM7pgzL+paXdiFKQbmleM
MoBTvo9aybDrDt7Pa2N5j8zBe86T0QlZVtACJnUqG8H0kbCedEA7H4LRCsF6sH1J
fBaCtdUg3gRmUy6Q7NsRfKmk0bhCA/OfHGc/G8BAavI2ufhkVaPJxiR+P07wf/Mf
db2uDxEJ8X74nlZLgdFddXusnYeoqTDOH8ZwxbV4bRaC7jJoD2Axc0stXGs4wyFo
kFkicuaBYQ0oRZL3xulLA++ZfV6cBrAV6FF/mfE4TEAVZL5PutKmOtrcgU/pcZtK
latEDScKPctqpdFBw+h9scFBZsO/80GfrmM8ldSHRCVMBbr589cPcc/gv6bY71Y3
PaXKBzwBrDWycUdgW1SFXxHB/YO44+t5ry/cKt3uMVcLd6WW5dKZSZdu2hFqow8S
ZZHxoherw1lvxCc4qPfyLnMWBkrX5cdijmVBko66QWu+czxC10dQEWJ9Wb9ytwnA
Dg5l0Og3lSxYRVC9aqfQhAiLB5nNhvzivNKEq67hoArAEL5Wrv6+A3yLnOiAHT9C
h3ZlvyUApes0d7vOr581avHwoGd1Y+eKQl5yaWml57o6g8DcHZgEBUWOukxnA6U8
8BKE55/i8FnElCkWMenDHjEBbe7Xgmn3pbDlgAGBTpmrDh7RTr48FPwqsAwHRyjy
LSxC9s5negh6QGlQAobcBfC88XWa0cJPbZjdTBYDOV0Sp52DoF+j+6TwGD7X/jYF
83xCflNQ127mSURjH73HLwgWhU4ZsH2kI5N4xlcT8Qr53lASQNXfUSlDTbsJLfFD
4crdfMWU1HMYM7vHXUA4lQyoJAPFVkWFu0XN4fCywtE8ZgzS3R1kcKC1PjM005i7
mVa2CyJlLBC/oMW7kN8asKY9e/3P9S2RF5nne1QfJc3MTQW+2VQma+xIZYftx984
T2Ub/etLmvyMwdErCJb8LIHw+kfwbh4Dxle/6XUZDP9q3wSsP/39o6Wq/tX0Fv6f
875SmGBOozK7WCXVMzQZuvITPnl0Mzyvt9WrEJXrYRSvHdpJzfjVTs6nOsBb/sT0
5EBEfUKTAwiLszri+R7pFZIWKaDz+n7+YwjGT71nPiQe3FVKinAuueU0D5AEulnS
+U1HrVve0ZM0tlAWTq31JlKHfLSYNYHq5J215HOunZi6vlUI9ZPUSGlsmWyeL+om
cfmoXgROAvFiYpGJ9PWfgzZj/qKsWuOWWCN7mf1SSF2CNJc4kZPHCtRywUPLoHCR
VlV32LHEHw804XiI5/hYOqHZMaNqyRG8oQY1vchYmRKVhr7LWonJlBOxJ+B4//uQ
yTS+w/j+NjvU5zWntBGS/27rKREGZzujpSQXhb5KdT8iS6bTfJEDKw3x+FHQpJXw
378fnKZ/5xrgJlGRp777C3LZfoe1qPmvxVu/lNlIyDWhI5mBzA7m3FiMlUlfjU55
oJLx3D7oq11X0mzIm+p95T4M96HS9vgAWm6lMKigYCGn4gjA5mtrJNlysmsIN0Jr
OXzIbYvnXo4qjCTokLEsTVpT2tUiOWUxgQytSmm//LOmAE5Oa598J2dCWaZ5Mxoa
OJhFNI9u4YSdGN0YM0gFd5Ua3hBCSwuOl+yp6rkjVV48WZSluqvviBEfLHXMLiSq
f9tClknfbmT8Hk8Ap7Q7BK4usnIfjKTmMu/cjujmyca3E5rdSSKyLKo0E7bejUAw
42WZMndU4/uzycLpcDID1cHJIyUAzJWC1ZbEQLC324VxO25aS02tsFmKKqAbCTsI
3ox1NkeXkm1pG7/c1soY82f4i5k5bGj+gEZbK0DF1usIeZASCFX63YR7X1YEwUQ9
uq4m6s6fTBkvZ+tdvnT4MEB4TeYywpcmCTdzkmSOJ9tOHQ9bo/MZIQZGkoIM8JBA
0nl9nTuq9uXEdioNFEu12Ja5udYCwJkRgtryNBc7TxzjE60F1hAqSaTogcoDLLd0
OfnELM6elID1qNay/+UCR4JRoRtnk5fjAEfu3jMwtg2lPrU7PBw8jjKBDkcQAt2a
VW8uHzicWq0l3Z6C/yYVosOSUJhWodrEhWDSd7diTe0hMCzztazTBC6qj6fUx5fK
ilVlJusvCLEfy1teVUpMOF8mZysiBr4oXDfjTvPQYHs0aVqdxl9YPr34CTwWRJz6
GGo6sZdIFpjNjRAceVmpKzU402TJTDVCiipcA7r7rS0q5FlJUw9ox2bElpmd0QJ2
oCJz7uuEizHthnOjdNBnZ31+G1bWLXX9YSnBtB/Eb0MEBR9l73b/euoo6RP/AJW5
jzmwqQMODwaGTDC3NgDZOfmlCpjn+hM3dHYA4DW2ZcBHI4RfD4PoyQZvdAcgWH0L
ZHOUAiSko0Bogpql5v0owOKa81dTGQ9/7r3EjJod6JGkdAvbzzbcNKLL6XWP/9GV
kbCjsgXPZadPk6khIKmE8Eh49JURMFa/+nvhMWGpd5jPjpGcynYNAuqMCrQNd7bF
Z1dCGomXa6U4tICWajQISWjNps2bmnVvDBRlqYGBU8tEv4w5punKLZY8/BnDiado
CxaEHc6+y/qNSqsBThMNkvl4gqPQ3J08CVYqdU8nGkSCyELWGC5cS8rHz6K+nhgu
3hNoE1usN7iZeXoOAlRpRmG7ExCqTfyxpPM0P6vqlyasVbDUj2Z4ujSasyAo7aQ1
VJgoBvlWUNISJrECccF6g3ca9TxLAo9WgOCLFl3nmQRza5VPUYOWLxY8mh1Bx6B+
acyBDW3bn0cBS5URWkLk36lxSA2qeytWJCbF4MenBR8dPdUlpVrmb1yQcO2YIwBc
R8aXfYWzUhoR0tJJGQekRzi363RxVugHsRbaNmpxnMoQ2oGEgAsNhmi09h2v3+Jl
zocE3TDDRcds0oofIAY4eu9krwO6acpRFh0No9rAOnEsDZtxmXb8azIjX6CbMDCa
Xu6HoeIuHb4AyZ9UQIBKCdf/HVM+TonI2a/S6IyqwKUHE4VgrNoNydL6bPxwtWgO
yZIWEG+ObarksmNIx2oy+xEq/KPVjTfdYDQXVCPn3QDFan6hBdp9ORxbwROVs8Co
fTmGIRZa3RXhR2uZLyANW0N68KURlvzAz5ru5hndZ6H4Ye1daQ4Mu4KAy2Mfk+RB
ndYqNbtVE3DjZDnrQYC957ddkIBfK83pIqouXgp41UVqGSfmU5QOZcRdLXI7fgM7
BOBdXQrrly+9K5B+ae+2kVas9UJqME11z4Co87PBVdJSjMtrQEZ6mD0FSaNegyyQ
H9GV758KNpzt2CSkp0p29N7XVGbiSJBottPPGDgfYo/l0tSNCcZyus1EGGRm1jU4
+UQ54muGWtcAwwLexBP3QS4olyGw4+cdUBoefX3IZ9dPnJ5gV2SNw0w9Wocfwxb+
Qp6+J1CYcGhNKsAfSY8oTwgJoFYUDsuUXhhGjipOpWTjLPpkdhRJDBWpWr5W0lFy
/4YcxAI4n+T7Arx8LZYxhstmhI2e1IclQPE6CwUwjDrufgzWKdP71kAsDvJMkWBw
CeJgDY8QxyOYD0iq8EFhZQ5udxEVj/gZA5YrT6wLNsBPdn1WGG942eTMwqySzY2G
7nGqf7qymWbSpThmQOFTRk7D3abiO+BnJj7EF3sE84OaH5Z3/wWmiahIY53xG6qE
Nd9g314lRw5CUwgyLnMKDBtrq5GmNO8RgryJFdAQsdArb3agkYleZvQN/DkOzkb3
okc9PdDjtZKNnIi0PRatjUe4ZzuUXUNMh8R++QhPZ4FfJRPOuF4A6krfCmGHmnBI
VDMCfyPDvj3qslNJbTWN9uRd1p1sXLx71csMuTpnxWcaWCXqvPZZdU7f7RWQR7m4
AgpkbXjBj+i5VbEDQriYep4yrwzKfYXf1l3tmImVwWVijCL8bT0Tq9Ey4sGZljKF
Gh1K3/0vuk9KOTyrXnTimtSknBQR7NKBNiRkdC3BL7/22jIr9dv2PzsxDkFjpgXF
28XDb4eOGAhYOJEcxav0USQuc6yKpqsdbTvV/GmfTyM=
`protect END_PROTECTED
