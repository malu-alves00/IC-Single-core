`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pBK5xmkToiJacQgqcrjTAWvZxgHbcfm5loVlBFdtufzSm9jpJ57980w16tG8D6hH
h0ORLcz1gXqgDPqUB/etzb47bGmczEG3sccniX4pWof4UP98YvYILz9lc9OfgefQ
y+6uNLNa1tqCRNsj1PbYlWUe1yT6g4HNZOODvqwZkVftS4i8xfE0KgEMgbKT4DmV
c06WVGNO8QF6glIExcNzuupJN2V3pBCO6+ekzJ/8oqr0yRYNpKZeneTuSJ3ATH5L
QBw1USxn+dtK82tN5Vnlam3wuugjBWf/oSHdTQwSr2YeRvy7RygSFzvVOpFBYTY5
yMAlRpfcgbM1o3mb+4K6LDVfSWlVd61hsW8fXKx+zxc73xtuelTU07wP6/YiU3Ly
/q0OWNP587gaxZKgfXgiXucDY0U/W3Ett6XXbyEBfKJ9o2QUzEq3kW/P5rX9z8nk
5og7E6Z+FzW+T3+tN2CJLR2PYfxKIiI1uPIjtMZxKc22Oak0u9FuipoyyU3fgBxP
2VSK4CQJLUzwp3WsdqDbyJwtDpwVy6L4Vb/TB7LFuqs=
`protect END_PROTECTED
