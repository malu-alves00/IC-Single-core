`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
q2M5gWjlS4rEjOf9y+yuHHPyTE31MmS0KV407jZqWU7bpTED0JYnNqtDCSMguDAy
MyDa4fMSGLNMTRf7gtVPDxpxSFTO3keWMEmdU1oyEvhr5EWuVGy+7VEWGCKfUhl1
9cuiNRLFX8uEO5JoMxC10ZnDUB8cgC1Uxg4VPjSwQZHK77Ro1DrlHdsYr0mDK6mP
JmAu56VdMUeDi5DWI7UeI48fKIo+IUCnL83sypZWgtRVZ1iJ+OGJDEpQp2lkyehZ
2hR8fndzPmLrEB38xbAGoSfpz+a8/lNdNirJRXv7JIERSUwqQDln4HXfNPGQ4vpQ
jGFMCFAG8UtTOr7fPM3t4HtgG40ARchTGZpffQ7Ir3+KMNPVnfud8ADvTczMD9+a
hLIPXnsL4zxIMjEG3AvUM/uudZkQ0+yCWOF1CfjxLr2Sx9Mi1SmJQP9z19MXc8sA
Mt5uF9bkrrZuzWWehoZtnNX9m8EqR2PkvAw5HHAkAf9QscCM20jAqPDlUu/cFxRq
O11cBxV1U/J+CdFocu76bNd6jtQKmEHLl9OGI+0wF6wrQtVvyErIHRXEipxXv4iN
8lZ+zqAWjnzDu9xElhIM4zmsNmU2OnuZlM1votUwSJKSEiORr4vPKzOdkDG8adnI
MczIBtQr43qCcl6LNj4D9I+WaJgTXXmh8dEqcSxqzj5SbrP73nd0uGp/RilEBTp0
HBWDFVC/hIWYKSSNyHfXQhe5Cd9SNLa9s01qfJ1/BhjOq5JBVyJtr+/+pby2kWh7
PUTYPkt5WAe+hYA9Mj8XQZ0FXYg5EUICpn6BpEoZPkV4e3l6b5cZtcWjLhajBcRn
NEh9k1Mu1bpH3qjxg/bFTuPWJd9vD6/xd9xjf2A1SR2QhkyFqWFlRbh+QZpAbe/g
1UukPAE/qVaOhzyfiGMOoT9i4KgYG00c799YV52Brkf91P1sNaqLZRSdyJhxocGb
mnSqREJ2Wr50KIdMvPl48SK94eUp6MOSUBGpYJCevcfHp6C3tbrYTxPoSl51qjbg
I9UojeBgw549Tmf9tpHU3qVjVGz3PLXCyKGFsOz8Q7yK//pPT/zQ6HjSp2LpBg2c
l7P3kghfprOhEHgEEnN72SgH75N7D0gnLjDYUg6fqiqfF8O0WAIg6J4lPNe4n6l8
mNmzK1OdmGazSnMIsEYZJOtJIXimDq5CKRXCYoZ6OvOgg0s/M5VHytdOdFv8/OUv
wPm69ld8+TDPyetQnufHKZ7f9Iopf1o9YXPsPMLvVn0bDcoNOVqbf/BWbBLx0B2u
tUXDkxjQpjTt7IpAx+99ZXIukupFR6yrRSpDIJH0G7OgD51d1ZSHIi5jFKtR72CZ
IWDh+mFOSc2Z/5GLBMQUrJ0SuwElFTv9rvr7O5GOl6BvNP+5ntCh39unCRlAFuA2
NJcLlcjnVBJ7/Pq7mG1XM2DoegWuW+6tBHmdV7Q92dv7USu4lYgvArZvE2jy6yvZ
uJmYjLKf7BzTHxj7gjuB90KsmBcEGq9OKpI4spA8ImWrKIqc2FuPA8/6k4rrSRi5
c8wdtRBs1UZijUF/vdciw9dMK+prw3PT0MO0WO9M+NCrBngAKZFMgTiTQUtm1E2t
`protect END_PROTECTED
