`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
K0nc6EJJapOTtGmXvrgX89QBFaa+LrU9BSIDBJ1GLwtbPG0Cqc94HB9dY8qqYi7F
/cSr0fIfCkzUuMfvjj6tEZa4yPqfkunakS4wvdiihftZ2Zr5rMUE/ORk6iTOzLXr
7iVXv9xfPtDmqzBgBwoNHDUda+vVOiHd8UiT95Kc4DpuRsipUKr5wCfnEqNADuu4
6sm7/cJmFZBR24dMCchPIzBwEbcxKvD1i+eKka7pWD2PXODNBZk0D+wtTfTbZFHP
bTjAKsk0M/c+nkKcNvHfZ7hm32CmGzjZHKiy/UoqrWf3I7o+bBdzfz70wrkm0+5a
QfS+FaY1rXZamoaGTsM98xlIJZ7F6por8VrJnuf3odSt14/EKNumaAEfSuGCP9ex
q1KQ98N2gLamAUdOL2lyoFyQtAASMvtJpZ2lQ+AVfTuCb7ll9+lUFUoTisOumFLx
HaAI7WeutBdXv3lieabOYg0JHDZe/BwufsAWcZlpdbVj2iknniWOPKxIwP+XO2cc
pivhQRfqaouO8h6aGajSu9hfoi+ZrGWWahJp2XwwipthQo5a0+GsA0VHUIu5LR7+
4CLh8vQTibhIxo29yi1tbSvBJF4j38GSATnlQ2vUWNSQw1gdMLv4hxs9IS+1b3nl
6Zp7wNKjGeU56NXhRawnDfKlCDcuq9n2gM7Cb3ULyPLJptkqp32R8rVzjo5A5rIP
bkgBoTEffZYvxEhu4cyBQLAKHAkv9tU/gShebk3qJ2Bn39byfHsPYLIXQH6lcC9G
3M3IDdYKwDYHFkK1DNhEy5bSavnNCtqkjlHoSWF+faN/X8P0CMTg5rjXn7rRv9dI
uv/PrMgpDIgUyhy3jdYLRJ3WQMr0AiuDF9j0eJXCFkHDFyYAzg7rQOlWRXYGrWZ3
+s4u0uHjs4A39O47ZsgLhkQ6a3Y8E4Trn8NTSkoI0BU=
`protect END_PROTECTED
