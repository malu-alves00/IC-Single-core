`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cXlEShckgs8Pf2Z67WphjeFJZTHAhpALKorSLsGkiaESxAsHrWg9n/0LAsbwEIXw
r8MJASEz1qYhxnBeFxGT99cRUqLFoVSwe7WfPNsYfqyHkGuqhKfXlQTNTf3clMyy
0vw/k5LEwGByJ3UACVdJz/VSlqMsI7i2+lzlalecbK7WkKzq/GJVNVwhwRyqP1Y1
B8H4uOYlnADuP7ySNbaHXdtSxhyind7a4TP4ZbH4nNESjW22bHNwuzllt1sPPlNw
T2x6+WTpKeeq1iwQ07l1J6NO6ZKpnLrMHmJ1cSHJztRUepwvpSyHeCmWx39QSDSL
k0Zi9tqXif+O4ciMudQp6U+oW57HgcwR0xQUkJOKHPf/8CdW0/c0VjHW5+sdC3JP
xWK6ssy5T+u5sHOvOXv5cs5Abk/6iTvJB2RUeRBCkvgXa/Uhbne9gpGKuWq3u0Km
Ju8u+qQAHUDbqhYyTGB4lQOQxjAfpoXiD4sxLpc+Ko/c6QvlbXf5EV4PXYDbk/jC
vwFRZZf6n4g6czLk86bX7GOMSWh/7csFypWNbRJ2JY6/vQ0OqqjST2v8DqUv4hjo
J1y82JmDXzEjw6lrJDIT+B2gbTQPA5hyfdUyhsijUwx8b+gzccEKnrlvga/QHafy
ZaXo3c5CmSUxRRZq7ZPYLQGUvfP74mU/y+wxIDL7Fa0/Uo4hl0UEFzMDTzxReRbW
sa/AyiP2ilW1+ofcKPWYRCYNHiQ+EjE+eAKDFI2+NTkA0IBB6rk2k0Gtr2zl2rVF
Lqq3qZypA3g8sNYUrVt2BzIeQ1VUyHrckER1/Nvz1oa6x4AuwQYV1kkNdOWiY8Ra
fnefo4X8QimnswG3JlPk7XdF6AqrJbiYRZzgci18Qt6PrYM7XStoempr5b4lGKdo
RJb1hDX7BA2eXmsxSUoOZsFb52dmaMyuJODr9O1lnb6xCTXgrz8C10DBEQzqXEUq
iZ2Yqvk7ZrHmQlWpOOuJgGPOURp1CxGC46vZoRMKWm7sjCWKiewxh4kDWTpxSQFr
RjogImRXiqBntNInUyrrSOtwi/q6VrNPbFEIK9BtEF5aN7awA3yA4HDBBvqL4zGA
MKSJZGqEE/JTN8bVMdGa14B5wIp8RjGpR0f9LxxDWLk0JfWQibAtAmdAgHqbD/ee
Mfo57YLf38i0N+fYg/GI7jjMZ0gDHhh1Mx/yM3Hv9Dv2qLk/uPhhKLHt/OaXU+mm
UedLdU2HexrX5FA9Oi6Ciix744d4IIrpcP9Xq/nU7tJhbuSLRouR/HIq6DAJ5ibI
syHocv9/71FRF4VwvwvH89KQz9zybNxcbzpTG3mp96WG7bKyEpxcHwKX+osMSkwL
Ea3HRQUp8XaEK2vm9LFuNT6Z4gWOM1htsO2257cSmm5XIFPd5pDtbEwXXFCpgf49
b4ODf0FFtwGhNWMVL3vJ2A3yw8rB0ds5bjHi3QflgJxxXoMPMl/iQs23vmyUrpVI
finjpkzJuB3/vz43IdY9bGTzzXOijMmJq4QAADG337V3HWNOw1z7qf4jPISpvqSc
aNYlPaz+4Djy1uR1qSdf8rTTwwvV0A2qxESL7moeBz5Atmsse38fS+mUCS7egtZM
mWzBWGQCOlpZOm2F9oE/Dca6KQVA79Oa+FRNGTwQA/blfUgf5tbgPuNo99atGZMt
7Z9bvz554/E3DnGvIvUS8LkMFa9ZeAZdZ8XWcy3cleeGCI57qH11GU7bLLTrGHQ1
iAW48TXZT5YjBTPeSlUnonsjQbn+o6O0ktJ3uy3vlZTvydtywFXPyS6FVBQ3Jns4
Qw6x7kg1//G1MhBjQG82hc8ELCGwRHj5PzYqNC93+jS948eWJ0ngtVg/n3/AKImg
RRiDs+c3vdE5EU39dmn78C3VjjA40V/z+Lcfw/dMUysuWb8NSpfIKXqdMGBbsiKo
VDs7WHF+PpBvRkQvJVAnfbQHGuPQHOGrJijnxx2yre6wsKecW+QpDdaXG9JyZ7RB
ffj1fhoGStBu9b3awxq6oOdnmtZEXjABp4Rhd+EpMWep660srk7cgHqENyJEWTcr
n6VYsT3jiB909gIma8+bYC/5LfUTjowmDGbg1PXD+bnrDLrDyZOQ2Fgk9iLmXo7R
x6eKj8gQvmRC3QLd5kabX+w/oBkcQrKpc9TbdGF7GBvuaUVXyz96o4/VYtTYZibV
RfJXxyoeERWyeKXqDWkgyFFV2lGQv18vln8sY+Sw9nGCaebXkyYr5GKwlToN9NLP
gPnms8NJEvo53aFhb4nu7k1dP8wDKYJmv1ZVaaR/gxVQ/fZWa0P+6ImroK3eDl3E
8i8eQgcF4LQbws8bKvj6VksofDfhsKgXnq1lQDljiCYBL51QzyaGDmxUGFlOxn7f
hvaBJXrfdilAJm5yVfOmwH1ttxmR2pl5vNyOQ2GAc6rURCRMN7p3TEp7m/PeZGOW
BKslotLm3i5yhBZCzMO/dW8jo9CPo4J3jO0NVwVFtJnEj4Ip6mW6Inok4LTDk/Xp
Q52NMnGK5eyGEPe84+r5H/CZKPYLLShUEpMHTz/v5jpKxxDE3QZ6BSuTNABq6+sC
nIvTB5zVVCqBuD2EjsJpnlp66ED+vf1L6mvqBqXDMB1lKk3snfdDbqa8hgqWzvF5
MZWTVfRhnL4Bzk2yBkVLV7kz3mGtNp1AhRvPVSFEANUfjBfSMv5VBgZZTH3OCTYN
H+hDPxFsgI/byC/f3SknDdJTnvzQaeTPBDhOVt5mSvMm+S5K9T2rczoac5MwpHvD
EfR7zTJe0RNj7nhHjnvkhTaFxD4fua2DjFrTtBfvSZbOgsR9i2dUp1xMN7OSt2l8
Wl0b4fgQKy8jatQPyzoDNIm7bsGV1Qdz0K++fSzsd3Np49qMSY719P0ASpyJtAky
D9gn3yLgQlWzlm361Cg5kDUZG5NSdECZBs73Lczdtyqn958MSQYlqqclZqsjGCE0
hOynX00/ito8/2pAxXcwdJmXEr8ry0BpCs47/2MQiSApPzq1BFPd4/menzdZI9v4
6hDk39ZMZb5ioS5wrkxCrp1obGOB4nJHXSx0hAmxDyLGaLnCL12Z4HdhQteq3ESs
10zW7wMiMb40ijtrMJOXMHQ2ZU3+eGGMc1KP66TLhqzmflrU622wpjm+JZviLQm2
fHem81J1YCob96N7lc6YzjmtIMo+BeDyBE5yMZ6fqwulFqxHD2AC6rl7wNrmaPvC
TO3frXPS+JfYiwcTouUfOBIEqu5eGjkLOwlsXopdVzdCEpjWT0f/bLn5aLVr44IA
n0Ouxg+R7KuAdUNpDXGdiCa6DV8c8qwTc2WNEnCHaDOwBT/wrgIBiOiyy7tMgWaz
hg8+JGgDohK86JCFxSmM2kQ+m+XgB+hhEIv39G6OxAVdN5fxYvtjYq4iIZf8sgMt
ti5QlvcYF1goaBC7sdNOMM0jdJTKfKV3vQK6zgDQh2vQkkQgpiuBykNn3phVImrT
5V/n42XMhvO3P7QZaSpiUU3FJHHFetB1yDogVovTAT4s5BQpJIN+D69mPbTqnzZF
ufPEiIn7G5k3i+CMVflSBFSG+++1szJlnNyVmwIt02VKuHAj8wwqkwD5ZRVOXmOc
6B45lavu7loSdvQ2/Bi4kNJBrAwEg3RsEuKJiYMN00tx+8YvAw0QenW0tRXu0PBR
XDsiywy4XVV/Y9a/7JPdxgbEIX9Qwk87quX69gSODVjetZlT+k69wrANPcznEZM9
UM4DUvIAERvY7Bm/Kdxyo4XBYBFARnJKHRhhj15yY6FaKVopDKpR13GqOERaQt9R
5nYD+LgsEFjGGvcSxBYpsHLelRsZqKZS4IhjWyAtc5IHKmRQbCklbHC6xOBhnPRH
cUvGmPRoTqSxNPRZbYnMFKpa4eicKPIKIUoWW9jAQ3ACHZwPS+dHtV9vl8zKJ27w
heXEEoyUG5/OEUNGT7LI2jx3BMLzWBgRTq/UHg+d8EUt6C/nY1yDAAA6G8gCpedy
NL4+6FjRa+5o1EelHPdZAl8u3VEJcr2Ywy5Ohk3SAqhuquwILmTkFvAs/NBxjAt1
Fima6tbejbwozEYuAbTpULvezEbwKH3mL8JAq1JY8M6O/SrQRwTl1VfICJe1mpEi
IZP4ICiZMci+4gT91DJJspE5WG+LnKUNHXSEl1fFKKZGwbfxO4eE9Bh+WP2XF/Up
7T1m6YcFixG6IMl0Zdk7c3q9d8wiQHkkmQ0v7c+UGSOHdDor5DwXJ9ElYHEzqMyK
TxwpoEnTrCWLabHWVKqxomEa3kSJhq6y0UBWl4o1mZAeT6hIwME8B5Y8a46zssF3
z7VA9yGdKPevSykTrSCR+0LFwIz2ovhErroqHCRklXvihB/u4nh4aRhDuZplu7wS
btY4NpUguQgEsJOWoIaGGQ3jAv9+A9CnIV3lnzXoyzr3k7mxqKdG7UQDzb3rSW6j
YghmDPQ6HMLqgvr7X1JjG1ZAbrSJ0DqcNuIoT8/EIR2pIbsssQ6Tb9m4A8k8/oE4
6rea2wHHxtjAuPWRQHSlwBAC3n+DATSlevOXAo00tWhp5jnRi9R0SKK5/q2xmEdU
XpeVS2eZLHN12e9W1ezLjHeZe7SwADuUT8iF9JdB3y9kl6KgSa/ZmyBSAjz34OqQ
BgvlDAE0iJyUC5xPVZpzcihZUr6LnMuq+rtTmuVaqoCjxT8kGzF8va0IPymG31d/
mAYShvPlIgk1M3a9o13Ll2nkmBHdO+nUIlai5R0Shq8k2dS4KuTPbYtq/ALUYTP+
WPvgDcG+yi0A7AiuCjuixS8CJ0ZHv1jbugIf5KvJWUS6lLBzCO5CWieuBDpqR0sN
NWYcZ6tGGM7u8zcoT5kDCgu0LTa3lymGVBQ9qyqTqQPXElra4+zRxUKzSiygM43b
5peK9YmeL/eTyBWtZwYL69lHsLa7OeQcUKi6a192UTXao+mLdFEajSUpm7z9ocnr
GtMHWdWbtxy7/mT9EspX2x4tG+0Qj0us6dI+DWsZOba2qsOYGJOzm9t1hF2m9d0e
sVd7/bBSofTB0ROmcI8h6pTQCEIGTRfdunNqKHCPBa5o/pufC1TlfTkd9b16pLna
MzfkfEWmJbgL32DsmO2QCCvs7zSSah0hc4NPzYv7TavP8OhvAj2Zzd5Rqz82L+74
YqxmY7USu42snECCf1pf7kTNbHcL/B6XTGlxPvJ5JaUxU7vgCTikoDp4Y6RFoJ/V
FEq1w5sXctErmdlY8Q3+7WIttnMj+Fpo/oqfEq5lUpNoJ5RS/QDm+A8Glz0se4FJ
f8PSMCi0GsOWcDvn9HVr3qiGi1lc9iCBcZZKD+8w0TyJYXdWLKPqbugv1ZTECF6T
/24sUY6DWX8PX6rFx2Qb2bL+O+/+oa9mMfZvQN21/aX0eVcUaNpTsDAf5MIzcyF/
YSQNUYh/ktbm+YNVjsTWyiyYVgh5QNXh+SzFeNAUAWPi7sJzqk+I1ZYXHBw6XfjW
ZAXxFEesoXhgFSR6M2H1h4ZqtRgpIpB5KbZaqLQunFJgHrQq65a0GoURnd3DsAhC
4r8kJjV68InVg74qksbGtV8diSWi8WcYuvCQSZqdDkgO3cIJuPurA+lxFYak3zdW
514PYsV/hkURBYcW09GN7frpeLLH7C5VMRTczJhi03Q+ofcFEhP4T4S8IIlV11JJ
HqICB4LfKyfsQBBoJb+fanHHQiyJXn+7x/IoMzvTFg38Km3JhzZYlvucQvhDHW/b
OrPy7c+3yp35XZ1ZzCU+fejzTZTAcyXFMx6nhAPQUe8Y5ZfirVhO32zqdUa7vCXD
1WOcDWgdTA5ua6CcJzfwLmBy68HTlKDfg0FHY3tMGBbQMopMlpAfZlTNxOIJTVeq
2uDAEBwKW9Aa9eopMhXwekXrIlDYdh2WnEvrU0rWE+mno7zrZdsCS3Z5U6Ln3bwN
6RAu5VU29FUs13SRGLEX31Oj+gZORuwDenHmwseBpypIuykCPXPKHSjwdbIqK7mA
ogNe7l9JeWVDJy4f9ssHkv09rwZbgDptWcrVsKPB90QmmGm0PUzfbjGtb1iGqpZf
yaaWqTU1cwn4NtyeDQtAWHzmL6UDY5XeLJipR8x+6QpGKmVOEypbqczV6X4zz38a
6DlnYovxUsw92Rlp/8+NEhCrRxMuAw8/NE0JydD3wu7x75JtAFn0REyT6ETX8uJ8
umItUws1sp/7XveT0XTma+CIUudBZ6adpyLjE/+TNqGIlWcyJujXNGOne+MbnCOa
eFpomDqiVYmGjk1oN2kLcUFKv/Ln33Th/jCzFbnaClqPK1sGay67E2RW7FIq1uL+
m7jvdakPJ+Z6dEBSlKUOhLMeu/LyhM139nNbc0dSUsCU+hYtsjrfvbcGGPpB8f13
Ang+WhkZqN9srwin58AiqMaMVYgVNI6U8zugwWAHlhLXCmii/RcjmReboYdzKgBr
mpoECWprH0+6CAJN0Jsziw/1tjBrU23uPqd1Sug3t5LDu5x4AqG7F8zZ2Cq/Ym/m
aScYHJ9y8aGRLUAjnfl+K2ZEojQepTehHEsWm8q48IPOXXINQtO8b9t9TON+mh3c
iVZkYeHLrQMXsskxR0uvgXEpGzt6pHVoYlaF9ws/C6pOpieOOGE9g6ccU5gzvSXa
LlDEvoekI5/ApaMAdQggI5trYJPyr8WTtbWtoOeUwza4/Nfdu9nSXe74xHPzff+C
E/UrzbMVykd4mqHAocmwBWRQNT0nNMLZffG2M5K2eWAwu3ZG5mUVuAAbSJyPHbCa
hwnrbF0lGnWHqq2UAzLm160jQzkwmW5vtIOpQg6zFZmXAAozZ/Jjj/7SCKwC96bK
R1EjSj1vyGy9aLzSBPx2Wf3h9tr2o2uC0zCvg197vL3F7GfrAq1zOKJQy034hqNe
s0g5Ncq6Ae7vwNbKjVQruBfQ3oEwvxjsVc1Jgo/Q05gdqX1jqHnJGX51L2iRB+K7
sQRVh+YVupp9KqMmr7IENAs82m/zRmUKYA//N6pgCrp2If4Xwwr13v84Dda5gfRG
lrVp40xCZsXOl3oIl7Erts8l2BFmq92mKKzMuNLqvGw3oFKDxkC83TLnicvsgcYP
+2KhpuydtpHdO1UAcBiHVNLhEYaLDSOCZaxSNLvaACPwpHipVsx/YRqAdhWdhDZB
9FbnrL8D5snAdnAccEtd3MTTo7Du0UFjBIvQfrZPMHN9QISw4Ptgo20AZu6ZTrPk
STya9P2wG54rMvimU60+FfcGfFxJvhHyxOcOOW8+zUwl8VTGGWol722MvYvPCnyb
efDIzuYA1g0uAhKht8B4yr1EjoGzhQpd2iGbgQ+yq0z6h2QqeEZLyuTh65d6xgLk
sX/QGKylrpdt3Quz+L/LjWxuSEBg7NOMI7FcZc2FM5+XHS+fJ5SlhTouXPNpB0S/
atp61vSmOnKduUI9b1FjWQ+0gg/2kOCffdgSVHI4rNUJ52/ZSt6CIgEXC4oigkfe
8WEnjo//qoOA2jLTHDHSO1mXjmpL0B4CvoQuyBXO8ITM0NJIrYUNko+Ddn8+i0hm
uy4wrGwgyUq70C6BZvSv8haNCVQyvx1i1I/Qa93so60GS6GrM/SEoUw+7UlmJsHA
yNHiv8OHvDSxzDBp980M1zQSKLDVZob4FseysIdZg/CLoOva7DhvA16cEionGLGE
YtjabfAot8bYgzAh1/tJr2oWPe3XxpqnAYhXvV4wVankbJO5ky+GdCvgUXw6zchl
EL7gSKxtB+O6Aixd0Ph03jXyXhdaOIrZZ/cyxWMyGJDlIJpz6mMRNvqdOc/9792b
8CLYKWqkwNAIc6kVh1oQ/SqcZ6Lz0by/MIpbTrHBchEM55vxSq68i7iItJ+wa1O2
xt8U2P+I/DjBrsL7sWJUKU9CIpiXlz3pfNNYA1TUUqq/16yr/D38EllaEe/6EbZQ
mfIKkY6E5hSnQSBstjeKC/tLRddcA+dwcVBwUoWZlUs3zl1uZGkKTZ0k+Uk9V1h+
BKhuGXUcsJjMk2im0WXgUL1FNHpvk1zubcfpdSUIDavDWcRGxPQd7lkEY/seL+Rl
sp9LakERDZQ/dHT6XzC8H86BD375VdLJosqFsIwpYUlTr7QiCYrSu8s+Mnzf8u3H
2DjcRHECmIpD6ZIuDW3hlOOsdmoyAlnlWSxQQ+MJ0JNEhN94wFNNx3gLhG65Vwt1
92ONDKKXe6EnWDBX7b5kL60tu8n2iBW/Hlazby+Rqo5gf0Ryv+61qhNEc/4fQkbb
M/3S+SkpZG4WxQkMjsEYusySyWXz7vY5bj88FtxV7sIu8r110/6eo9Az+iaETqvj
JaAe+OrTkyqm2DhTudBPMPfJU+a/DCoVLkHMsnAvbCz+UDvUHBwysaACBgD++Y44
UC4Zo1eyu5nnS8ApjT7BqPaaTy0y/TrsUIV7BBu9e4OH2088z/2yUX4i4hKWPaDM
X3aLEqs7B5fE/R9j47Gzp7POeSW4DeA8QxNTBGqcB2gwqGmSmta4QAzebAiDGY/c
+7kXtRnELFoNu67CsCDfzwpHVMPRA8uIMmfWT9FuvtPK6+98qICPc80WoGm2HBom
UkNhXCIs1gjK0YkthMzEUwrYOa9lEbOtbi+RLB3cXd4pv+Oxw7aeL1ourZbBFJOC
exmWJMOZfsARYZmgNeNvBml/u09TQsAo9Re8pWEgDQYnzWv3Rgwst+cpTTzBeGbp
8gqFiqeMzdQhBWVTGjMrPyfxkdLncj4CxqaHbomEL9ALXHDccPxUfF5FINXCnY7o
gKZHqAqyXlhzkQl2lRdXUBlV1nGSF18out+I+8k3yxc7xF3GI9NCH10tyApymj81
6llsKe++nyIu0xGN+qx8TYHrKsELyYMRz9wJ04+SiljF8cUuJEgFOh2THQrQ+FR5
xlh/0zgU/peLdlElCFvVImlg1AvWqE9LkI7YqHnDPG6sdqbLYLuvyIZNymOUWxdZ
lrFXnPCx5Au8khHisL/ufuMo0aabyanP8UzWxLtzQKUt6+0JhGuk1nL6i2d42uCL
jB1l+JlslRRjjzY0XKgR+KJpL5IGqAg0kIUhEp+FmzlpASUEqkqBmGRrls3b6t1v
K+tyuMFGnh4bmWrztnfPT1k3J9eWNcbRU35+sZMophZuArnQa6kQj5adx6R/bacX
nXiHG1IZ8t/iDm73oX+mbwK+dfGGZDu81SAkrRGA0aR8Pd7o5IQEccVDM2r2J+6n
hl+GYm2O6uJEhMlViqCD0CuHhlb+WMD5G3OJKlBJTx6j021lB9QOS5mhPLlGIPHr
wEa0SlOuioO+RBHDezhwQy13jeEqPKWK1Sl42Nm4/H8xCY/6a0ULGKb2YB97N5Ez
MZwHl9Rt55LlzbN7aEMAwYzdVOz96M4LvzM0TKH8zMV8bEwW1jbHTtCqKbuSkyvb
UWHfO8k+OOV85BSdli/w1jPHFSJC7GgezYJ0pIm/ytEmHgSLQrUdrjfn5Iin4Ax9
xqCUxBvDKfP2jFCcumbsCoe28QGy+Eae4eLpsb3IJPfsYG66hB1d3C4mINy3Oczz
k/X06tUIvi9jCCKqLeGp3KqF5aIJBWgGopA/bx/OvcxTJTteDvCd5Aqe2hHtyBpZ
pW8MW8krVoHWAzwAGQ4GKeZymFaDTAX6CcJiX8Sfm4y9mfU343vweeQZcNlqY5Zb
6RXbL8pKkWwcTb2pV5L7x/ndMLjjN5vu9Oh9GJXBHXPeO7c/wythorZzKWD2tnUq
gkRcSglYE6E3Xin2I7v3KKJiX4eTi21cqm2tCZeWhRGLNYJJCqJ2Q3Nwya4yiWfQ
Hvh7l1tx1JYhEDKr7SdUGEq9LddAt9HzvzWWte5M4wMy0NtWY+kBayTXV1UWuhHK
0L/3NV5alBBgUDDaHrB1SK+Rktj5WM///Me3d0/zwNXnsekQHTu1OlTOZmdrA+uM
49wsnHrFmRdZus8wUs4ztSlvyYmItwhBgSunD8Nd9I/FKdgphAMBqOrK1StClwKN
8ckPm5HQVA/lOdhhUOHXPv6N+C/VAulO41AYDDnMiMmjqSQGCozqAR30TVZrg54y
539+YAJbPZZQ23TgpwW0atFMLHAulq7EJQ3HLQAtryTFCm/ZC4nKL+5/8HAx/kaU
zTybzX6T2jO9MPNIJk4Xlx9+NyO1HMokK6Eh58XOwmO13VEXmzHpSUI0gaLSjbLh
lNrw6zWZr7cTiysvGxRpVphvpMWGHZL84zr3aispfKn29b4bFHl9umZ1H09uC934
q1rBgRLEpz9vUGu57ijjiT2I2gpsAyWmZsyTruzO9j1AXSpXMFI5KUsSaduy/Jgi
AVftO0lIKnMWcxGt7g50dA2P3dLyGhvLW7RkrpsshFILlk+o0ZEBIJWEwq5JFIRR
vInCDbmcOokyij20baDABgf6H4+LDHyVNd/xdApeyOiLQo6QwOuqchRi4FR8Fove
QNe07m7K02sNznq1psEK0J4cG1i1fr+sFQEFpVluJ/a1nESsyff5kLrC1tk42nPz
zX64fDCj9W9AbSUII7p/0f1bzGpcz2cAsI+QFbSpF7gc+el3epJfdAPXUzIISh9P
s0WuZp6VyP1vXf0iWieA6kueChtktWjsu/h6Oa4aeIUfnJR+AUJNQGzgWjoysfDf
E0obrZUJVzovxKMP4nk4U9jQLBpAqZqH3jdmmhOXFZca9v3iQOPWHoLFPPixD+Dq
pKCHTkGtw+1KiwzeJEeNV+eBUBe7FU3QHjF/ybj7Ed7Lo1GUv6c05wXs/cAeaQVh
4MebamVBTiLH5ypLO8eOKpHuRvLniB/qx/z+7SkAiO8ftNyWl3ZxEZc8cgovqZsx
DXDE+hkYRV75pFg+iTp95QeWTOkLx8C4Nd/AOKp71deW01J5uiMGK75aLql8GC7+
JWAQsK8I0k356in3M5jk5cRq80Ftq8K64UG1qSHNFlKHnqjjsVrdid/wDU3T8emF
T9vh5+yZyWmHw4zPEdw7jxMhZDvIimjJU7QobU1nNZtCfMIUsgH9Cnq2zARNj9Jq
H5vKxBwC5OFeqiu5C434BgxrFoh2fxiDsiuKtgSuD/bGh20IizRp62tA4hfQfC1D
rttXlJIXrdiALk3JfKEWhU4WefOfmmRnhZRwirqSFU838xey72tQcDd4oDJLEtLj
8m3PiZXlieAntobcoS1QvOMYbj04oE9wq+dYCI3K2t3mWMnRJjFH7xtFzyhP5cNr
+Xr4y2J71F/9uJkDsWnH8yAMyVHICItURnuWH3v11Fsh+mAeIvfsCwaBAU9MB1Lz
J+kFEKK7BbsmndR9vNykXz6xdZn/2ckOfELHwuSmIluMPPvHfbpGni0nbemZdTIQ
XcXA/bccgdwEG0UPPKNaUa2tNdZF6cvSUVJUfYOd6r4fV731NEDnNs+xnUZFgT7q
JA8KtAWbT/abEdcLSc6b5p4mBFysIE7CWjjkdL7ey0kiWePz+z4HZN1UZytm/YvS
l/YEMeSSwZqdYkxw08vyW6F1RfBcaCwGPenpnajTSVEFL2io1lZfcfNaB3eUvSan
FrpLDnDmcR0+24QkcB1OEIzbrqPlJKd7Pp8aezUpzcmu4+tdz/5tH3DCRYG4k2je
4SpMLTkrzIJoTSbT6ACVKZgqxJLAIUQenh7vOsAm2wh/nQtpRX7QEM+ldMpUOqP6
N32K74/GcRdMJP2jbnUixjs/VNZtWOLmeI0AdE6ZQ3DPH0lXhU8w3NBHY2kMZdwW
UzlSQ6o/k90iEA777LMBfZ/07N44KgQjDFHcPntTFVQueWEAzLSH8ZEhE+ylv0p+
khGTcjKddTSA2/MPpsipcHV1IDilQyz/aG7OOAKh1RQupwiYYdr0aSq7HZpksjKp
7c1NxhuzgVxk862ZYbgC++hW/a4juAThkaq18Y6HCWNgrAmzzM3ejkA8k2hv9I7/
oAKSxW0E6BVqccsB8f2upDS4/0ghAFm2lF7eNXMci6GpHmXk2R/4//738gi3PLgF
G5JvzV65I4iaCGagO/YsxRdZi7DGa2yvF0iVxyFO7t7NwBMB7dh5xfCEWDqQzeeJ
95qaCCWDaSRorngQzNoQehmomIvb1qN4l9X6oQ6dWs81h+pOtB5V4K3yOOTiIh25
nKqoo/paABEyt2Fbtk0OBh0emdGRasgLAduB5Jk5Bcst+dbxVdbCee9dSGNqepGG
/Y6af6S3fNOhxJDDM67WTjYcj9ZWDN3RgqIXxWR/xlw/H70v/ukzG3Eonzom27cy
w50zlKfGMcwl876JmV60OwIEwB8CjA8yitIvgW3VbL48YWIPFxAYld42JPOvq15Q
YM2Txe76/nV2s19cFC+/ZEaG6ff4LOyLHzAePI0uHhe+GZD+R7/MuOWMv2Y2SR08
onucWKc82VKY0n6GGVG8mJihLJw26Uq2XltpQWdk95OJ+fLtwtW7c7vrCmMDeMwx
9uly/6w3MHxwMeF7ZbZSC8A6hP1lRfchAt6yb3F1u6uogZCrkHDUp1tIeLorJ0vn
cuvSCw2y6wj0AxGeUShyy+VRWkfPc2E52m3Q3gWX5IHxv83ihLog/K5hlizX/hbh
Zn/obdMypjZgXexaxrtvPZAmWnC3jyS1Fy5nH8UISc28xm63p4+3DpUivKLUkhHv
ry/YMy/N+z/LNYCO9+MFInLuE+SYYFxavoFCCz/ouY485Bsm/vlYeYiDQBr0V9R0
2FFbgYF6BfXHZy67bMjLoTPMs6llKPr+ewQQVuf585w1rHF0nEd40/RO+X7BKJsN
tvyqVhZU8zOKMpjtuWlWsZQ8prCs1fhgkw1M5OF2bG9wTLUStBxsdFpS4XwLNPBO
de86Gdopadlzga60WvsRNlckQXgx0NL6N0zKr+y+DFovLPkVJzOI1c5MerhrHyq+
DuvE/1aQ/LdSo/Cn2FE8SOsqkVK1oM89pFIxZIAnCWgFNISqkPzAMX/XMo8EDZ/2
7csurJOTTPMGvPZrrqauiLV5eE1dcv/5zk6eJ0FVhkRVmwy6aA/tVA9IDQzwER5k
OBkpcATXg4X5jY5v0gTYXh/DOZRkQKG84Yf35VhWo5cKb/hDQ3+huKhnkYRQf1FR
O1faVpJIFIrmVEdb9yPxvupcd340UkPQY0UkDrHrodBdiTodm8bbtIuPQRBrN5zt
9cu9at/6ydFIpfnitfvvX+hH8ZbPwTfiuNIjsnE1EmDYvPLr9FMEZgAYynVdEbAw
ubDrGQwszWXO3zB3pa1ENNPzNioDYvikg1GuYuTMtklJleBmsH1qeJgy6EZ6wMua
8grAx5cG1HoxTzaQk2+VHFyWnz5l6+NWUFNoCRccYhw=
`protect END_PROTECTED
