`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5uVwpLkCBU44pVTDX3ExaVr30hjlUOkS4P4UCg6Ks1A1fIQG8k9aGrxMGoc/CZFj
p4jS7t8xMIkgfw41yEo/99N5Lf7YfP5/ZQRwVllAcJkYJIIFqtZKKwPHmK+qPWcR
3iDixS8pqTyYk4zfCkp8hsfc1/l77LE8XNH1dP848TYc/OjL+CjGes5dJoqFQPUx
xud8S1jOVPrY2asOSVgjT3YRN/qejGCBlTJ8+GaRNkDiKovbU1gvyi8h2Nuuvduw
92Bd+qhlWe932sjtJrV0Q72+1TNa4DrRYwSgpZ/D2KltM5yDGO7nZOHgDzgPew96
GtFakqEn9jhtonSlocGkldgHlTnUEKClcDSb7p1QC5QTqz8WBUQ/3wIN4oCmxD9X
v1g5qCWHcxVGtnnAKM2/+6bbH3KThyZiPqC3tjv0IfGrYigeTa5/tL7MJRNPQ+4c
EaJJodc/LKvY69P4pkPyGOx3lAyP2uc22n97zbKZcCeFjWiY3KeacCUR0fLEzXdH
tCZKB/JfMKxKMaInNWdlSufRfJhDMj/k9caavvFSuMmIMG7dXAWnHkqobnv5X900
IScfvxxwJJ/5iecpY/TIrfnaPPrXgnKjZ2VMfuBgQEfRDQaA0XMmyrGjLKl/qUo5
Hp6s9qdOzr1pj9APpIExC+NaH21WvpSnHmvQDNFxqt3x9ECiz0gYbpROvOrGDDKC
SMiWIgWPeyl82BdgR45un+882XrcELAb8Jby7UmIyrmK9MzHFk4KELWWffCWWrDU
+xTJOgDNQJ2CYTiCH4F1OS3NXLWtEEkD8kHhVrGWySap5kqtCi24fVQKB5cc87vL
nPCTkH6DnhHmInQbEx+dqU3QEONKzpWOc1q2Aummfm/wHXMmRDyiokfauwY6LJVR
emCxC7V3uxDZIWGbE/q/3ltppc3LxZhn2Xl/HA0YP5o+e7TzYAsMInIbWfxGFHJf
dVFUVWqK7XGEWcWND3rHbhrEuYaSewiK9Y1AP+MnPe3few7glDaZrt02akjQ00U+
+dDe0ObeUi4aEQTLGKYSW0hs8zA79CFnUU/P9XtBmOBVLBYPh1JsGlx5tX4lGdzk
dKz1M30xVv4DuTDZ7YR86A==
`protect END_PROTECTED
