`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zHJdqMwH06rw56kStWI9m2mCnemUFga6AMGuNtbzGUBQyDuwbIGxeLbwfWKjowb7
g/d9Dj0KRbmqnj9qpVc2I5/JcoTUNZND/DPfmu8XXJiP6Rgzb+LOeVL3i29dBw3w
dtP/MAjuDcInLsEu5BYN9VfhLYC8BoRyxnGhWRVpXosQhNumgrFYRdZ8aQY1sw68
Ozs0RbstxsIcNvAH1TkceG3b2CfgkOEAFsPFPHm+rkUb2K5tzdl3Z4sy5w1wUoXX
aS/EgJvrh3kqdjHAdj3LumOhZlfTmAXC4xbn57GAz5/jARsmcMiT8kmNgJTY3TSO
vrbyp9nccJHRrnvZYR/WT3fEgjmYWAF2FrGAxatiBGjb+z3o36ooLQ5bUp5Rlv1F
S6fQLANIkU9wWVHEHN2sDfZkEHRqBkmoDNUuARdYzxmcZ3SV5VAcAHnWW9MWW35l
lJ5H4j6u4EOl2rw4aNjvH0TPDhp17WBf42YppqX80sPDc9nQAbMvAnLFtUQ8FcS/
OLUiDTkO/grYi4PVDLibCayF2SKpCZmBr8KEgCOCy3aIer+Dq0FBauLkpsVCQ2VU
FNjRL2hKywZ1azLhuaao3f40Yr/PulbKwegEdykVp+H4mG9ROv55ntVXFhZYTvOK
OhWvxLG0BWcwyCIOG1vVng0ew7yfEyUrg52vpaJMbvR1yMVRMcpfQhBfRUZZIwTt
fxHiG0UsOdUAQ7tCmb0acOkcZHX/4EKTKiK0MIlRc8ZQrukS9vZsG0PK9pyK4cTp
5tIiC7PTYWP06bPPJOCJHPuDvLYcthcZex3KITXzlfIOkt95nafyg5TsY82kSrHl
aA90ySMCRHUVEwEHaozNGlURXews8aEb92a623M5gNC0UKb/mQ/6cWlBfgND1+iH
goO5B3F6YodBahXgW4sz65RzVxeCBtqSrAfet68yfWqs7t9RhxwgQ1utyIcj7tah
2j9ILm1V88EflxOZdB8QQ02UPXSMIgZiHCBtTEhbVbWMdVIkoUoAt6iNQ9ojZDI2
EnV3F5relWgJ9xMZFSTPQ7JywZSbapTllzwK5M6IEDA/kzV1asJxfFBxQWJuxHWT
rZxrLIvqlWjocG83FZczNAU5/04UXXcbAow1mNhlj23gcX2IvkxOOmtiHt8/lZLs
BUXcigtDXZtXeUwYPkfRUiWC12/G/2HlOUdeXVSp9q1uD8Q7+kuWiilxvvREaMRG
xb4ifJFrKP6yTS0kcfbOteP8IsxQolSsWUregBjbZmPli5LK+Ly3QBsW0IMeNAOC
pT+lS/peTMgNkl7E/oWFjAWAtB6Ny9JLZf4vobSQLybzLWQLZ3YzlpMT3Nlnpeil
FsRMuW0nTs2O+x7Btdh+Gj8CSc7KNI87+QQ2cfap+FkJNGYTQ3p/kr856aFGFSgW
ad3PH3tOh/rgHHWODlDU/J/G6jGkfmtdLWUcRIAyL2uux9aEYmTfKGjxExtMmajn
G9ZW+CYY+rY4S9SHnVKU9rf06nl2alnThjR6Lpm1X6z/9KRCKkJ6BWo6ELwgxaE4
t6pNYVGU5ShjrUAsmQH3jSabwa7KL9QgIhhOQaEzAvGhPyRXfMaPTYbD2i1Cy8CJ
MY15Lhu6yTz0RE/BlDsF1X2AVN1YHadEqGflUwWYAg9MtlY5Xq4lMOINlROj4FfQ
IusoqJ2DRHQ37ohDWDNEoQ9XeD+n9BSUeoDl00ya0yDO57+1B7YfJj09FEBbLB9m
r+DcR+WreIy0iEsQDMkrCm5RtpzpXJxttMqORdmbKGaoUSKM2pLqKMJ71M4ci5f5
EkXDevYXU/rTX/A9bI6gQB1M44zRlJT43ymIcosbO5UCTBhEijtp4XNfAndyBAy9
DrlWgspOYLDdwgAlqaD0u5GUFkng+bgf493gfrO+XiSfGz6J6/jAVNQIvfhxgyT4
btT6J/qDHExzB6eP/Y+PfysP5XL4DrK6o+XZlpXTF7RGecdSmU4EWqxRsIsPQL/r
lgTImQdXUSLDz8JARaW49rhV7zXNzVX5jc2UEn6dB9vBN3ZyI6fTN/G6Ry211md9
kOGdCYqWruFkNAseSRBVFYvEBNEH88d44StnjG6aeFr3otpJlSom11DxiSlwOgJS
Mim42gf9F7nIArdyXwuwPE1kDMl1ZWLvGD1nbpu679QYmzkslGaSHbJ4XcU6VsnB
XnzDVxvU4bn27TpLbVruems7E7d4DUpPNFlja7Py/o+kNTczXESAZdEgsaa7zHG2
rTjdc+Ah+JouPqkzaDJQq2/r/1swn03FL1kOJHIqkuunlxNlb3X+IKSgf1RhgAri
mkItDwH06ao+6JyjP0hWaKadBMjOtVzsWcwNEPRTYY3lQ7SWabDHoK8d4wBEK+41
Wpv2vPtD2G1OPZf/4FzxdjiyYKbZatZnZ9PwQ/MKFAF9gFRzM167f0r8Sx8hxEGf
OyYmvspVbrygBMWo/q8P82JWHcYU5VoNpJtaoeyjeNla8RRm79zaGZ2ENDS24UW8
kmHX/KwaE4LJGLtQPK9SsTWvOzG4v1/Q8I0WSB2+O0A=
`protect END_PROTECTED
