`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XeyNQ66KF/N4BTmTKAB4h9wz1YuK9QeJfvSfJ/6hgCV/Es64JDcOn+wwwUAemorA
6ce2nQEQCdGbsmBPj82RVdAeFPJM7psWcUbXOYvwjDAnoMiJd1QzjhjSGS8mDnWm
1QG8o2FJigIpsQrbFb0DA4CMbdH2MG8x8BSPQtpIMPrj3eQCz6Ngn1+2u/isiflu
AnYVe+WWnn11w+lKjXo4mNViCJ4VCTJfAwEAKWyjW9meTW+mkBcXZHvKoitItNAt
QWqbA0NMuEB1QwrwKkHAgvpe+fD/kGb7BiEcFcwmSur7bPPhuc+VW678WPXzS+nt
gVw9de8t06S5uTcHsv0yKOoaMxjj6s9vvHFvZMy9ln8g2U8xIpyQjde+Gd5aEQNF
z3ITMpavOoHNv35jKCVBZn6Xi0BxEzYNt2BR0KN5TsvjxZzsXcIWqlie+k2HRMYv
z8Nn1g/RGJMIHhFt/7kT4Y/WYRXw9s7S9Ssb2ZG35nikXw/XSc3tA5QLlvQPX5Xg
bTnWlJwQvgW3ZAYkmrxCfx9SDhuZdzNnMozRZyR1eXw/d81jzZ0FhWdzMQ/mWd0j
SxJL1dWteO4nvruT7pun0w==
`protect END_PROTECTED
