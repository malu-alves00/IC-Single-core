`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bsvtkk5MsKX5PmnlBhDx3ieiNshEV7aQXwLxGjCZzk+du7UYk/qiYfy2SoST5+72
Ic9gkHDm9RpyyPTDnZzl4Mq0Yd4H2msXtfeOOjm9BrHoUAI2PmcdOzd/EQ4hSNXX
4xKqk/o1CIKxf+qtSFROOlIGUF7rPzfLSQ/t7yzSofI2+ka5E0DxuJOL+ULuGcMM
e8s+JFKYlAZfDPiJ2DbZILxzBQmyvZNICNK4KWOGO0ar6g4lu1hyo+m9zHj47jar
b6bV82lf/yVq3T6pj3qnsYDduwbcRlsOByyinEAMh4CR5zqzV3EGV30mrN4EzybF
03yepOdRd07ZKVN7vtevF0pb60CCyfecnKz2LDCOCAPiH25IEcNTNLyM9q+87Dr7
IvSxOy/70ZNX3R5s3Wpc4xnfL5zG6EqwuN2ghgZotEmQWl9Gci/JYF7XTbHlAvTm
Aq0nXTKDHilTQZ3GHrsX7nOahLZQjf2U3Hj2z32id79HrqlkDG/o6GmaIZFCKLvb
HRJwWglfPM6CNmPPyqIxqlBZxziM7Ak1zNDdo4AEZbDcgZvbsmQW3on3loYgDkYc
0hCuntQs3t1hjjsOpCo4gBI8xUfxKTv/e0n7Yu9t5HmAZtTNEeuX6bv2wRDZ+VMj
em5goPurrxXQswmy7WHH0gK0AhTiW4uzDEZp6TeIliBpfMrQEgfgAAjH39rTRRPZ
08aD1QNTkT7xk+WZeFbRC5cqNK0GH8t17GIPAwwK4PYVu2KXcfkiwGl56LJ2mPFV
p3fvyLkuX+yPSrzBknXqZidcbqO+hTfthbkyAYpapryNhn9XHnIde5TQkHnF1NVS
FmIVfH0LhW7tiqD7ztk7DGkkJ1MA2FbhHe8C3WU2e18lBV25oJ7Bg7IIoL/oiDGh
qPfb+9dReDJvhB8cLTG1yYVlX0VW4IMkhLkep3n7jZtnk1nXfF4tFr3298XwFP1W
fnRdeo9uVFqgVyBgHs0nRY34EeDEXk73gc30RFFhfrap9rMs/ueRqc1A9p5GUg4E
oB7iu+gYmU/CuiHZ8odd2TbB3+fm4aiycxPYzCwzTq4VkspGs2R4FzVeieo6WniY
pvLHwkUPa/mxGEOU7WF6HVZZYxrwK5rBZaSmxRprO8kwOX2wUgYs4LrATjEkMUwd
APM8B1laQ5ExvL/6/FPrVMZUZgMCLGRXh24PAqbrpKr1MmJlw5O/Ei28/HnFM555
yjIqNBQbX5OYBIpkWerU1SvZl+DoGOnFVNfz+dK5G4e4Pz0F8Tnj8uf+JoISr984
xiv/HNx47uFhHOU3Cm8/QerrqTNMtb9YUqoxWO83b3J+CBc+nEnb3sKEH5Pcx1+Z
DS4t2Zbm4KamX4+5eAbi0gLkZbY4Fo7DoV2raX5XzimT/TF4YHMHPIXtUzIbrCYA
etjyfN1p4kcDIBm6/6B1fN01JxPQ8xpbQWmEVEvZafRMcqaKiljpbmCs+vVrMvxk
PR2d0OJbmJWP8atsfEmFOw8lYZ1gctrz4xoKtToBCNgnGT6zjEvMlrCliNt9B6c3
Q1zLxdzHloBRAL8frSAWWyGJr7KhneiJARmaEN3sXhiEpaGI3xR3Vz/8n/OiMYz1
M9putxNdpcuvky+8n6RgAHbD056J/2P+vhRXq4biBZkHGPGtWfPevUAqKKJnz9Dq
f25GTKvljY6gtQhrRtlcS4H2Z4AxUgyU8QKuq76jQfjLqO2IKtM58jZFdPy+8rDZ
casapr5dxqVnaJF3wzcsBQA4oA5nmuPSeHL3wTWHjoBoaRz6dpiqnfuCia493D5V
kshtnM6U8Ze1POvL46At5nkYGkZFXwFH8cLSt7CbqSv4qaj8NpAzkNJJ6b32JrfQ
4tyWMLZuT0xsRQWExeYJNZJW9AFkefdAVaersgaa9l5ePDVColCq9akP2dyPzeqL
S43ytN0Vm1G5NJx8+kZLMuIajo0RuxRjaQHJ1SdRTc0PqpjjuncAVbrS2BP0oGXa
FsTJuTixP25O4FbPaGLGWw15JXX1PxO/pdfU/NDrMTijTj/ipyV46ZpvQimI74AH
q/em3bq3VvllauYcbWMoLrzblkCDeiu5Zv8qZTTeu/OL0k3wlTAf20IotbSaNY9T
Ec8M81RK0P5dh+GCMNjFyDTTwpQCScY5sEkZQK7FHnwQgBGxnJuVLr7BH41z7erP
5HQqB4RJKpJfCJkr5QZuKUadPdi1fy5TolfAC72LZleZ9UDL4nGv7jDJLsoi5Lsm
DG5H1kFrbOaBvFEuBsSpzPZVCvuJhDz6CquC6MMs9J2H3r9ygiopEvy4X++T3PpV
4omj/4GA4Ila0i7xuu9WnGV/CxlxZKsyHpJZb0ucP7M3omaveXDNk8PlueJx5cj5
yOhlCqV933epnPsHbeAFFZQuiuj2M6gI0ehqV8jPv7aWu5eSJCXhKwignUx2KjMV
742yMILzyhAbFDM5PbcJceiD6JgfonzbcvjXOBm/syMl4YXWsSGfoHcGCKIldn8h
ooYkOcK5hS3pO4FTM2pVbiPInix9wEKwPP1Z/MuZw1CKshwNmDHrX1my1oflVVoz
IFFhzS5qYjPBBPjGFSc4gsKL5ATfpZOqYkUCNjMKtl0e8PtKkpxxdRec0wgYdjvA
J8SgyCOIhcGICrQm86WeNs8JUtug/F0Xgym07K/ZQryGOZC/HS6Af1nEvwLExw+0
yo7fg9m7MipjEMK28cJhIDCeZvpsYf4fN3DyHEP5NWng8we5foHksd2u7hVvzUtr
0F4kHC4iqFU2Jn7xi7ZF+epCLnQYm+0qXNzpfeBvpK38adedjSDfvdnJwWiMIRj7
8LpbScuhRRjXZn8ozp41qCq/7rhvGExFbnZkXUwieV/z9R+MWgInY1mZX96rSoKV
sFRCXmO/ccU8AlMjrTGwPq9N2PTRIoFaK1TIPBxQTZ31aoepvW4lR2a2Yra+F65x
yaN2aihj97N2kG1a3mVXLMLdaE/AkXhTbKDoXBgwQN5QACz0P2o2zd7QoKgsapgK
EankOfIX+ARbYk4qhXbngNx/euNuXwoeRoOY+cF0IXiOcCgytb2UtZtmQMrNHrSF
n6aDGRoutZ3qw21moDAYESCBs7Sgm15vqtoCJQua51sEgsge7XrY2+Ls7QPOgPgv
F7/WPS0QDJQ4EDtzSIIpqCbOWiq3xsP1nM4xfuDUZE4B35l4l2dPR50P98jGgAJV
hMxqyauG8CbRtYHKHkOlXIPZfQaVXxdAfto6EtHhnsgWCUQU9wj+uTo9ckXXl/Dd
7knqjKiGHHVRJrH0pfTd/pnnjEAcVUg76BkE0FUWA3lbl4Jit04QgMOvmBugHiFb
tSrWvuKvRjY1/TzytxATU4X47rDVacMaJtc3vAItpaCuNoS7Xc4Fy9WLCEFtnt9p
gWJbRP7VgC+mYTWJtQ31BlcLsrHEEhB8udAnQBn4CNnfyrtfHbFfdu+GBYDfjYzC
OglRrBUZRv9i8zqS6BYSnRxcRX26SnDElCsRvOt/+y8=
`protect END_PROTECTED
