`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QCR3vFfSyc3S2usoPYCi+oo6FJNUx2t0iYsPpV+mwObbbL5GR7zmP13KW9FAydK0
mAttyRdDfZpI0MkrkF+k/PHMHBBYpmyPzKJwzErhnayw+2a1RtkV+js+drirP+QM
5EPH1kbtSfkyd4tfp2g+YNyQNg6sLFwk1mXmwZ29hzfxKZ7jJyK4PrEMBNwziRDv
NauQID6SQupk2KqhX6SHsbwEgJs9uw8O82cc+D/igqoGnZ9ShxN4DhoxI4JR2Eu1
piTDsu87x78gb7M2D99A9WgNK1e8nKq8zxAaj1S45gwRHOnN1GNVmI3bNZUWoz8h
NqxBc88QR/IHvLDG2kwOE0unUOflv81palsc8/jnP1S1CQGdQ4pXqa9VfuuzluZO
0ZvCECbH2PnS8Pv7J986cHM3KtVT4POz+KV/i98a63kMiAnKacruOje/UtDdF2QW
GkfLVQJE3XqkLDHshQbFqowIbiHjUeyfPGtsJ5jUPO/n0OhxgtVJhHqEvwNU4f+r
9FLYUfH4hw+E7p0hCrxQgyoIxJMID00s7qxWkPKju0KSSIY1LCbRqDzjSDuXM26d
bjjp+j68+SB9ugzrncNGxtJbJsG447wZg4ovPwqFqmOyp+qIt3+Dse7KwATYAXQL
bhsNo6hv6vKy/9ATDwdkLO+de0hdOhTrsCCZZqBN+FYoIAqsX2Ex/cFt99a9mLUV
nlmbOBrzkbMyHGH+4CgCZf3O0Pb1GcNNiufgMnFHdwB2vV340QWr2bjM6k95CQbx
dzWYLcYDHLpIYHl0oHV5iD89eXKxOXN0XXa2t5f8cUbACfqEJjrYpvueRhFE65rH
L9qRHtDahqgq1xlhW0JxwmGGanvQBosBg1VDOjzT/VQCxPJBvVpPshi6jNUzI+UM
lDHY5sANL/3UR6L1SJoHTHFMjhNKlMB8dEag9DFRYaGXwig7xObrdd0a5luH2QYO
3fPXuralPZjgC+Cgtn8IDqYS8qIbMqZ+8LZXCYPpMbawcwP5m1M83Q4ZWrRnmE0s
vglGof9fDmYGcfzNjn1KizX8U1eMS+JpSevY4DjZy+3zeSEzoWo8gMDfVHx1PGX/
JpZwtLUhJo5KS3nj+m0we7k5IQBnNoMcTghXuzjEJ+UQkO2+fqj9GrkN0rCoStRR
TnxTt8vW4qSiW3/1F/+udBdBUaqaWfyqv/MJZU2RE1Py/6oyYUbb0CIUSy4wXMko
L+q2uFzuS36lpm+LbJ84YZUa9cR3Kp1GdvBVhTELVTsay1nnT3b3iAXIAWMzscZP
FIMxi9YyaEHn2xLP/GZO2YmqH7v8XDSrcgsnTfp/Yna4R7bVrlfbz5f8P/VO1yl3
sMlgup/teyiilb4vMLCwzYwTdbnsQ1AGvaavpa3t+lCP+fRjVCbSVMpFFhe9kwPl
P77eiMhikvmo8F1r9aXutLHeGhrZCvruuHImuPMq5KwXFRsk0P9v6FUEL75TFSLi
FOk/91QtvPvbaTMcdH6OMj0OmCdf4eXshq30CevEGZw4rwTQW23QfpJ++UkjBxyN
OUF9RnxNMcNDIUZnt2cN95qWfm8u2WgPXLlgjeOEeSPYk373DpnpI3Dtm1LhJ0rU
R1BCUNJw+leNgitEQUMfq43tSbjulKJi/8q71Td9iOTvPWGLWjmx5ODavEe9K5i5
ffk6FMD+UA0x7rCYI4KTbUAhpJIJii29DEHWc6A7Qq0KloNC6TWFifJIRMePYwkn
FAaj+FITtpz3HIJzNLBiDLKHtQWfpg2EDXFdYgk/K5afKWuz2dalnvxtC5pgvO8+
TLxHlgL4QzFucDmHF3AtpGGf7XPWvyEKvJKAH6FMkVPBF6kwWAFyzv2LRD+SlHrb
WETadonxL/oEGcKnObd2AkvPKTb5mRLRX+pQ1H0/zdJu71+rSDoPIZFvjfT+bMaO
le//Z1kNd3sEX1u+4bM/sKTiDfz/ULJwktZBmLdoCKNSv5aIm0Hb+4gVeq1jL7+L
FGcZjFbo91/N8yy8S9/JiM9+TrAG6ZarbP1iulj0pPWxBHAAxqlrIVrO/nRLA5p+
PgaDvfsUqR5UjjS4K8BlGJvYEvpbojNdyVX4bel6dI3+LslMnOWrLM1DF4JHZ7T/
SgpgiixC8w6Nz+ZewQHW67Sh6Rl8+kA4tHLfhtp27sUcoKpBFyGa2h/bmtAnw6cS
6y7Pde9woDnr3rH5iouDjgDX3XWIKYk558G1TYdrFJKivPbFLLp+/ZPp6NDo97J7
D0B6cPWIPVvLzMB5s91/21Po/wEr/i/ukS/rx+9IAlVgLOo9lQ0BCzuH2Z+628vk
yI4d3AJgid2HMEwp0suEYQ+zp6CbMOrlnkUtzJrrIR/jCpKB9tcVjL3qjtOdWNPP
oRs4ZYWbV0/e/rLrPIZ8U57QQgVv0rgT/zsJpbRoH6+6hL4LUEOrQaXE4uInWN0i
`protect END_PROTECTED
