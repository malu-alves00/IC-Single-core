`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qOXBevkcHK2DvJipZc+ZYtMUoyJo8nBOMInNN7DqURj/6AtjLweXgM9fn4LdxJPe
xyqcf54UbogR/pUDHWqm5t4sehqN5MEq07gfRDBR+aeM4sHPR09T+eW2UCJOj/dK
Rbq53JBZOGi48q10XeXw4crRf19O2fvPuqdBqv35YuuFktYVlcfP+kWC1ep7TkHN
NeJBSEkDQn6w5JUtE/PyyPLQO6b95/hpWkX2Fsz8c32V4sz3sJ9gfHyzfFcxYhCF
AMvhskXW1B8Srd1R7PyOQoctC4EQk8rh4ug/rdKvojl2hiCz+rK98uokUAYZmAT3
vmXOhx30hTkCXJwNPjw/CIPpI1Evtuzci29Qljo++edaUHRai6rqnZIWmyu2BZCD
Bf6/372sTY5o3+mEubuZojNT6eBA8LiHqylNN7sdl1UAIOD+v25Hhopb/68Uq0F8
e5hqOQO7Z1ZVY7dHxWvTOFUijkmXCTvBJPDr1t99UtuKkJlHcyQV07EbfE5egnKo
3BdUjK+rztXQp65M7qRicKJCnMlcDgBCaDNrcYYBbGzMzt0sAu3OIdCLZYua4V80
jnt31VW1X7bduVD5GecnM2uKdE5u/veshEavczYoj37kcHDPbvk6ht+QZakL9CxM
w4avQ8UnPzOLcBL8joq/RmfXl5QdMtf92f/5xOGyWhb4siJEWIrZLXNnKpQCsCUK
CMYvv0tcMtZA2ticpKYvFO+hGYOmVTMZ6xYqIKEQB2o9I7Jq4ngllcPY3Y4ivwUB
2CKRH+3+EQLvAARBJXAIhMp52k0FRe+26DXx088UfQAUzIfPJbyWdhxrvFyKC3yu
OBeKnhq9WQQVBw5x911Ng8Acqres/pPm+4l7UtCEjVkFSKGY7NRZEtNgcPeVthYY
xf4eBptpjCCFtNRq9gi2wTzMk7eX3iodbvkd3lDUs4CPvhP0Rsf7koK6UxFkxFOq
yBOoF5ShlsnSQ08ix8Hw3u565P0hP5g9N5c0O+9koQ/2U6eM66FptlSzpeb/pVWr
yizCjbzlpPVTNd1NPDw8IyLvg6s7glVHGPknk2A2En2JC5Sfh0gKciQ4uT61ZDEn
shuG0Zh5UIs0gvWJey572TdEjfjojMyPMNa3X6z5ZXy2De6V+b2i3X1jqSgG1o6g
hsMrEre0oPoYcUy2CYqeKGUM8zainOu9i/FyrXVyX455H6WxSovmDtHjHSBWzzmQ
lXhx6BLEzZeuMkv7iPFYe0GKiXwY59OemhAuUwwpjcd718VsZPXojUl2ovX+L2a/
HQt+/DRJ5Hn4glyxiCD6rx351+JwMqQyzUbaSDYGXe8F6FA+LzAQ/B4UWdz24CYT
hQ2z4gABDhxXXlADPsJmAQw1kuNjG7S3UnhVtxu/IOhavihLYBcP62q+PeBfc3yp
5Fw2lQiTuysNNcSHU7nXXfQj8//USK6knTxJyj5IIJGRB/YitHHGLweXyGm4LyN9
Ea70xIk5hJwsQFePFADShGGIDo1anJa0fEeOsaLf2ngzuQusLa6i9XK6UROH0uaG
WrLYj7iUd/nQ6JcgVGLjFWcnimCWCcElpOg2BeGZDT6HVnPU7ChesNiXnoeqnw3v
dXxpt/NytklhHQ8tv1V+ny/87eaicP3RUZ5ouRQbOCuHApUgewyAC6cCMHgboBi3
wZD68BjaBJNneQGgCeh5jFfvy5qaaXiKH+SX3VBNYdRgbaUhoIlBO5TMKH8Jw9J3
+fmK+5QnYnlj74SZPi/6th1qyk0LNysvQw0PkuMnjfs/luijm73rfC5YIm/5tPLU
eLvpIziEPAal8iPlcsXzp62qBkv86Kgm2kSVvN4MPJySDJaVfLKYvWTLaRs6U+dD
hOJMF8TPItq8qZpQfxFbl2BbuX7SKEmToowHnWkVVdEcYB3FKTnuEW9XVGmzv0zP
r5zmUjeKXE/3cknlChbJtg2WoqpSm7cHl1RNb/ZD9gDG6FZo1r61vKokbsrtpbzs
CgG8ZjQs1PFzcSlUt7zNR9AoTvKzHXwlcSHniAC81gEt45Pb9/jAbWzi/yLs0B09
2pZsMDIa14ctVLd3Xzen9FL0EHKptq7Ca5bNwR+AhnuEb7vA0gpMz5uF4uwcaP0Q
kTdMji235QdGRA+uojZmKFLg7iAzzi9jt9Crrey/7IbBWsNh7clBRVAegxi0NBq6
pibnqKQf8JW3IkrOXG+yRUjzbccleuY2IiW05TobbaCKEd+AbWvTAUwTQ1ILDDJX
CswEHYy4nqbPAdrFDyT9mAvR8MUQ0ocy2IQ5cEaeB2i/5CPTAIVmHTtgDxySPceC
Tte3NMAiSwm3rsN2je2oC90DB2tY6xVU7C2e61uE/7uGeMhDBnbDofs+/+pSGQFM
MjqKAjkj0iM5lVyJw3CUWfJNMbUWjTMgeqOZBH0t5RLELsQQCs9SuIeypASdw0w4
N8Iqeo+cnX+A45RbhpEWbahUUT030S5bVBKKMTyl4j+qjo6v4flsHEd0KByXbpeo
4D7WrHXADYjveKHivAPeRnYK1/C5/zQT1UsUo8c3lR/FyAwBUetKafuaoUHhgXv9
C9f8jjovjWgNmUnwDLxcRkPYc2hnDskoH643ZL8IsI4n2mOjai69/Zwe96Y9yjp9
2+WG8vcTND21ps9wI8aHoN7hW0jWyfkOKr4/uQ0zlA7ER0W9cGVA5SaeZtdcbOsu
X/AZ9/1y4jUbO2Nj8N5Vtp10E/5+eBnt7AJ67Ka+Vm/KMWfEjFgOVa2AtFLmmxeq
slK6giGt7u74sg61iPVaTNCaSINIKFihDSnl6pDY5FTVfQVDppIv/+8gkDHhIW4P
/GWMKBGMpKslzcoK05+PMEMdy2ioUNPlD2i85oLUehLOKbFXwP007gKMcRZuibFt
kcOZKgTsGXXC66KeJHnLJqH1XSoQEN7xSDW84MAt05rzwp2lfTWeRdmE5G0ITQty
x/zxyBeaDe/ODj90pZks2t+zsg1gkTQODKA9Q5kvHu+6qY8p4jbIoqtfqlofjwSn
HBBwb4l/k3+nPKcMH/P3HnJfpSdwj6ijUvZ1PG8T186I7NJyF9SFTC5n0wE75ZHJ
fM+me6rbH+v7Ee/mhVOksB3h5qoSQv21E8JpAKKzCZxPPGdpeEsnnRI05TJj3525
lr52eBRfCRwMT6woXRqzba3X+p3nn4kFOvhVcZR3rxLXmnj0iJqkwPutKCuEcBLp
904wSt8NFGLsREyr+T2qXZPe8nmREeTheZDST+7DlAQNk2dL2SusyCPQc+11NsuG
eNXtQYvIfcZiJQXby9QYLCYZnZjv+Avnw3ydJCoHhMPGDegwsUAaaCNYvQDh7CBV
0IEXup5Gfp5LwV34nWzZiyBXfLWk/wH+0awgyudU8/BNWR2VbMwpmOrtB5GvXeI2
aQ0Tg/L9Do99H66vULMw8erH7dOoXp1J+0O1pgqPwkPfJzR5Nmd6EGfDmpObHhFi
QidX8K+5DRLrWEKK4xvTgctiybmvMldJE41dmqHFSHkgzEQ/SrgK9ORUYlPmik0T
IHum2/5GwDWpGkdHckdkCAQhqz8oPIiC4kFHjhUkIX1MlK4O/pbvPHWK38z8EF9+
lMfpkmbYVRlB9DjTA5wq3tXWtx35DT/Q957LnKuag4QNTR77RipVt//pI6+G60W+
COQH+qYbGdf6ltYe26rArR3IZZ23goJNU2yOahFKuG9ZY7r4fnq16BSKHwiwCl1W
4GEntzo7EeF87UI4lPnCgw/xY0ECzT+wcc7QJhvjs40BZieiZnUMkx+bGyLAVo6A
yoPnJDtscSR9ceavdEdUWwbGa11L2zy+NNnGMlZgkjFybR507rGzEVyqWCvjCT5Y
rAfrhj+SaoNLApQ/OzHRrWznE4V2gcf14vvSgJdKF33vVH6uswnRMQHpIMwa1hAL
kjq2x+h/rS8btY6j/opB00PCuNXi6RWeg0T7R46lu0Jw4q51axPfiit09LqR3raV
PMtgzTbZJ6SFsCjPgN3F57Md/cj8OytL4/eO4TlOC176cpiP5CF+44uybo5ujMBD
wCfUa61zloydaz56uYeptskONk88Alw2BeemOsBjuVyXi+BRbwTfN56nEtmqF0qq
GeYlx8NF8Ujg0OmP/UCJNWjsiVucxRcMii2O+3ZyV110PhoI2Oc5PBwsI4NFpfZx
4LqMKYLII6bvSkYEUZP6PfETDEefb9T1f7evKIrhFYHK1fAyufJVmryNzdyLNdc5
+qxUKYao8YIcQoUXDcGif7tvy2sf4zIYxEKre5hKPMpFWVULt2ZH80Sx6roDJ0Fn
wQN29XPMS7mzBtD+k/aohpwuLD8SZQMjmJo9H3bWPUZ60Uu8RGJfbA1fub/YeabN
UOYaRH0IJ67RdN1F6DtusDZ+hCRncT7KqhiXjtv3mDhl4CVLEtKNxF/gFaMjmpRP
4rl5pOEXs0fZUpSpMavTYu8SrkpJEckOEqMnnHAmqcKY75thRFORrkDhhkVXgYTu
p82JuQZu/yL+yVWzM9QFS2uiA6fCIBBZGqcGuTwjBz2pSkoqp2GqLZKgRSB3yG3W
UG+vJaT+TWoEZKjahx8SMsHSUNTioAd4WeahyIbVfGioYeK3qH+oLLKdKVh//PwX
VG5QZ+C8DNjfQ1B/56U1rOXMbbCyrfWv7S+VkC67i3ggGbQ5dItRKVrZuY6vBFEd
gB+w/dWdhSQBD+gjDXWbNgwRiz1dVt7aRl2T3v0WEAlV9SJHNzauh4La6N6Sd2zJ
8ChRaAC/Y3CmAuMp7ceYi74YMTVjqcJWTYiFqMuD4EG4zn0PvBA7JPM88+Ki0FfG
Mchmr9DnQGxIYRux3tTu7HhJw3jO18m/fKVCBa+VUGMsGrQsF8u5TDMbfTGLRp9a
sQp+fvjiMSCKas91MqMzvENPVCod8NmG6LK49lh+43ktU1nmSo2yX+yy2BQeMiw1
G4L1AB1VGYG1L9DaKPl1WKBKRyvlICRpvDXA9Tz2etdSWAsnUISA/5wbGJoXcgCd
aloq7RX+jP5Rfl+oAwuQMcrTREJPqeHhEDHca5XPYX39LfzGZBqU0Qeyab8QLpFV
L+AF2ayNWzG/lm7MBLS7vvMQOfuOa4W1bVeH6JP8zkRD3+qj1dULxnBYipMcIAWJ
t3GqGW2+D4jldU+gXzhdELUDZ3DOY/GaMuCEj0zdfVr+pNY/Oz+uyDh3bltCljb+
ZudtMNH680hk/s8Ye3rPV/fSsnTgBJ3mLwSnpV4PJygezZvsQr6Tkpaf2p6hI7Qb
TiAGToliCSVODZG0fD19LPc4psme4CImM8Dm6P9INK3XgVQo1nYc7nnqlJYIi1vA
Yh9b1bGOp1JyENfy+SPjXEJQRrMJl6Zin1C86q29CRRY/up7hsKaAm+C9u4CnlAo
lpNaIMMM/pFbLt7XtB+UN0F3FUOVFEYurj9TzpAKl1T30o3l0xSOwUmgL6RQlp4n
k/q9DrDYbWwVuv3fB4zRYteE5PvqX+kTJSsCGaPDRQma3ubCmUzQdn2yFbNmfR4H
PI62RObra3G8KXXA6raTiG7hWs0qaayt0t4RVosXSAlwSyOfM6xteXI22+iKd1qK
NCKKU/vEj0gb7v3hPre5kvlcDCITgiUfFnaXg416rddniQFRu+US7UQwuqY6eP9A
mb6J95roVZ37M6IbzF7reZz8RqjtGZn2HIkL5OA2mzJ7NxKkLS8Y+aBAeXGoxktC
wWdiGjOeMp+HFX8XgMt+sLqGmFENQ9wAiRxUYlpDwsl8ltf8xHTquWF5Q8n3YNRb
urjhqjygJR77Rrm+588BLKrERHfra5+4G1P55Y80DBVGd2IytZ+Q7ghFiZmcw481
rTdMWUcHIKwQkCjph5E76cdFwIdxE2yY9WVJewZ4W+sMazZUIrLk6XLoBBOqJ1Uw
vhNVELOcZR7EtmiFOq9HJotxsIZdsoGkMECfXzc56/QfWBrJlgVfbJW67NxFAiQ4
2Y8yuCgVZhYTvLRuvoFYAgh4Rk39E8qTGjD2CFN3B6e43Y6ENG2RFakTFSK1e0vP
iUcTrjK+e+9CCkDHtX0JPeCGGJ9NxQP01s8qz7/LqBxO9AOvGQY2sF6+59xlyDjJ
/WRmwPjlymk8sW/BO3peJrU0auLhKu4oOoN/j6689WmZ3U0f5YoumHxVpuvEj/NG
79JO4pn+yhvF6x6KtDucVemDlhHozSPXKeIOSt9IZWgRc1X7lLGFygmaUzEXzgTO
xJ0+FZMqjDjvSRESOadkXCbAvIvb9z8xKhUvrHt6fRHG/IgigEeQSC2cH/V7iCV9
pze0qDZmOpevGhDGtN+E6P8EvEQ4orQoJBlAWoRoyMOiEH7ZB8luCdIiqR9kvA/V
MegF+QAHUkeCd4pamU8Riq3Ngez4FNJSNtY+5IPXF2knf21zcHAV45J9mKkUGcrq
7IHz/Wy/jxRGUfjCRwSLwHWL6xMIsOAAv+n/cMQuNSqyjOVWE4laxHSUqFVci1S2
ZfRe56XEQCYSP+AbTAOFao++PS1ru7arM5Cy/kStONNa3tPf/Yvn3IO5TmTYuJHK
9g9RQefxuzVGoGYmP+iCN5Rw2HHwhiZYvNmEPkcrVb8tygYKlfBwdiMV5TxWFd9W
3HwVosQCj5GmC97nhfOBt02Rt0ApF7TbNRXFN4GyTprijj1Y6vpzXEE1Nycm6gWz
FPvUv7T2uMh4hpSkmY8fxBlz/lLZRsgbJHvFNlTykxGBVEaQvlnZqPtnfavqkvC6
hob8KaIutzS/CYuw+x4oVd1t5JWHW8M1KVDeXZeIFHPIP+QcjiwgATj9v6Qv9RkX
tcWA7aW94ZE3M27XVyXPPqqLgEO1pQsETE/n0rh7UIGrz292ctidHKTEF8dPbRtg
sQinDCdC2olhXH8+NYnz//b/ESswsBwNSzKuspTMDfjYj5aNF2Fdlvz57kZTAugU
GauSK/cJwVCiVMb+7uOp3Euj91NQzt4lZshDbl87gvNt31E6q6w3Z429DniaVGgO
D9dCt1xpo+d7/6grR7w8AZv5Bj1xUPmivHFnBhi6k9xmaqxrgDF8Gp5Awuv04DCd
pyOgtjAEVUZ8IRoFK8gkXAGiXjIjuzDC2a802wSSUt9PUWW3qS/YONZDQZnkSpUS
0hhZq4rBMrsQxWI/225NL307DcwOGj3pbfz6Zj/TIE1RMlzHWXskFYAUPMqxtR8M
AA6O9Q65LqOvd49fk1YTMyPqplctbgBLIujY4anxNhVzxX9zPMWwV0ext2JbTgnl
U7pPN4jdmgtD4YAFQbhahxq0VOFDVAUpUVMBHYxC3QbBNjmjDDl3O4ByV/L/nofv
50983DLi4O6Ijl+UhtpCCQDdBDNR8PMqmb0rqF7nVOXLiIx9L9Kr/IIz5+Fxy2ho
nPPCyQCaSFGZyirBSozgD9KjkUg/Zas1utXX8xZgO536ZiD6T4vtQmUnHBqNL9U2
hx3DQhIHUAqkoOtcpCb4mcLinDC9E66C4PoPZNx3ar59wElD1OTjKPAiDSINeaEu
zvmyuNCO+8mqSu9sSq/gKqu6mUdWFlbgPnX8hVZzbsvXAr3d3ZB8KlDEdiCIzN1M
iEGwUE4rdDhRhO3xR0dHnwkY/UmTShMTqOpNuqPfaCzUor2vt4Vxam2xPwVMQT7x
Qbpax3Zlpt/n1M/D1Q4WXhtc+8gwGNoMGzWv+O/MQLd0oB8juQRm2w2To/Vbr9WC
PrjFO9yEYiBzf7u0HY+A1fCUtERcPfDy8zAq/KBTdHN5jt4SHeklgMteU7ZUCyRA
VYpEuWEq2TxpEZZ9ez4sTQ==
`protect END_PROTECTED
