`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Gy+BBzpZ0HbFjABsz4eidcSuu4HqG3/BrJ4WUVIJMd633yL3dVBrZBevL5w/SVai
TCAy854BQ0rAjIQtdqS5+gqXGjFKIca6Oqv4Yx+QxLMB9XTu6nI8E+s8kv4kRGq6
8VFWYj4yi1arlGNoz1JoNOU3Q27iOgsjke4e1VjqsKq11LtET9gFfyCQuVRTSJ/i
+ZQNQ647xKJAyNlnUOFAEjC7M+RRktzkb807ySGquzVYSAOhYtx3PBS+YkNSu9rt
OIBQrbKmZDRk6qDesTsUpqyI2RdwARLaoUzGHG7Mb6Socjs/5qHNzZdoSNoLo4oX
3I3/Eg2f6xrPmdnmASl1pbY5h4cySH8x2jZG9Qj+dOcnX4LMiwxNCPvxt63wKBWG
DsrEkkXbB6kcG8Wueoht4rEOkNlXrjR2QX1nUkDZc1yIVgwMis6I3PHp4cL74gmm
xVhx3e3JMBIlKdzzt4YJw/rcPLd/MkcOHIObw5hMULP1iTqCgP/sdIcHvgCmk/o4
TBmOCYN0qUbNJ6ivnYT+aHByLrP4YsW/qJ69lgLnTt/+sUx6mh6p3M+BQ4rft8v2
gt+zgg+5zAEYdGMXHxUmi07JHfuedm9O5hzmHAg/usjeYUj4qxXM9JrmwjWxmbmB
6yE+W76/qgItiTa1mk56OoI7k9YqDJFC8wL561Wzd6gwmfXHLDYcNXdlROWPBt13
/ULkJ+LD/A6EOH997uPp84dEvZvbdH58Djfx6cf+FslfzXZm+Ow0dtzkXI60YR+K
SIKwBC8Mvtz+b5rKcoqEZhk17kW3ccQuGNhHOco+LooND6GbmRp3G3m+POG3Bo7e
VpFagLNNXnYAR7WlLgqPDYmpjNJ2U6W+qHIk9fl7DlsjwJltvdqs/Sss7jllnYZT
P3lmMKis/U9dqEGpbOHHwsAGYaL49mAlBTRBxTr9+0xsq5j3TMlheJQUkRg7AVvW
BYtgylEI4/ZtHYkuCGOCpq7XOYubKO2SKmRT+VX3NqRESLG4giSHSsbgxgY4GcHy
fgDOj6G82s0pYx22DXMeorXUQ6JDbKo7dgxg0woS/mfzhlkRPY/Hd8D4nh9vrFMl
mjnXiYy5d9rweJs98E73wI3tyw+medpjSmEjGOQhpwBxzHRUZqGjlKnWMdb+iYKi
HhzymZ+/oe3v25+xhhUk0XtkJXQ+JdbWlpSFjShBhb3l9WPREvnXgA+WMb8ssWST
svo0CUzQ976ZjpA0slquEWQQg9Yhj6We0zoXWTmDe6s7urtiQnH9cQ18by1a/Y5w
qggu/fSK5sH7DPM94c2BEfWOm9PyrH0SqdcRYu+d4/pQ54GQ3bnlecRqDM2iPsV6
X1KF13n3uakPS13v2eRcW3yxFq3D8efCy1qlVx0WNFCNhJxFQkznPWxuY83MUD3Z
4uMbwhr96AQN/ql3MdbK6ZBiNbkWhIywA9RoQ7tnrlIFpAzgAxA/h9t8JK+qnKnW
oUdPQPuEJXS2nDEoEPp73Ly/pPcEaAedbHGxPfC4nFBg0FAxH4sh4qyw6IJmoYwJ
TGjVFu7CPKiocmD0xaBW0z55XzLEoxnC82/nXTDlSwkxsFv99/lhSU8kxj5bpNwa
JtGHsd46TngWav3lvjj5JsERe7/xFpm6L2IkXf9xKR9Cd0hnmj+MxTOhXHLT1qis
4eRRgXymcyyrp8QpqglfgJmmAyjdoXCQThvejoy9icw2L8cT5peUwrx/3CRO0RmG
e+9BmzChJJj0cBMADd1qAStKiycz9YysJf0F8dkHjuIrRPGF7Y3QIoCc2eBt1N3t
FTFfNV1vAzNAI1tfHUnyIdoNlhVyaMvqUPU/XqBrUsr385yw0eKNKN+nz5PoW6P/
Yfn9DI6LfecLFbHgrKI7fkacvDH5+kO6EThGiMrC/VLcNzW22S/1J2kaArA+Yfh4
HELdVn8G2VLz54gur9MP+FkLjLitRVQFvhgid/+TzEiCJiRO1sEvr6Xf36Y/kWxR
DrH0atcPayRnx2BsCrBoSX8NGqbJO3blrEpcMZjkCAW8f6X5Fgd7tvFshynQ+JdI
gzY44yoUE2DrBdz6LQdtZ/aoMFf3RlcL9KJqS5Owi06egulmBbZD8rLgciH04xgb
RnswkYJ/aZ++vt3wpkw7dYKphD5YzmNjYrtaKANvQHa7Ui5hO/9s80BwC7diXmmc
Gg4nIPQ0CDI5JkdLmYkJPDZGgXF4ait4pIE8uLdeSJySQZeoVXQLpHsikiUiX5CU
OmuzEi71+NRh9OBGnKJSA6KuagoqJoJQaExgrXo5ZDPTZtbAWDN4Nf0C5nkQaCVA
sZeIgjh9nSLJ/lPrC1ePaLNo4ZMCFUXoEshUdwdFXgkr6QLx7DeqnngXvtX9z0j/
OrVj+5hzo/Vov4Qso+U24EVz7LIskZg1q7o/juOjuJRBmiR1mKU2AUrxLZC4vhvX
x7FjNDQWjiltFafHuE76m9QVsWprVZBX7Ne7xQYeUiOkrBEvy6M1Z8O3NkgGJYQ+
T27fMRVwtNJ35qn6XJQckd1e+i2+iPwZufjLgauCTAuoljd6sphvOyqhJSNQ2Slf
2ZErc4C8NXE6rxnpseEVG3UdjadeKOTBFKma0zQqqZ+1ZLsHPOFbsU80afnR2WoU
IOsSQIaes+v3vsEVXT8b85Scz/lXXa68+maoYWwYvsu/HZm4HwKtiT88/2J7ixTA
Rj2284DfZNbDqVVI2DOJgiTwOTfGsDJkHILNl4lmCcY16RAIWWLvxNenbTZ1ymff
Z98mk9dgJurHpm/Vzuf1b4WUwwX/5Anzz7HrwE7eggD7sPz11oGa8K5+RoauUOUo
6HBVJ2HplyDXZlx95BJEE+MCR26FMBtjyvkrA+xox07e4XL6qEFhmU0WmeUfEenn
hnXP7cxgs6e4RxyUYCfD/pQGW40hw4Lrn5BWWgtrmWWjCBQsbz7ddJ54YcjKe/Nk
t0fXxmtdS5MDW+vf7kULe1drBKZbxIKTZKNY9UYfBMKABqCc5kLIL6qSLaGLyV7/
vqZuCOkxqn9OHV2lu6dCkYZkRWTyQ8J7Rq6kGgzDo38DS5KaHE9IFLU/xoE7j2Nl
eIJK5iDvOJ4dIZjznXR4QLjI7aEak9XNR4+D+A8M015TNQf8qs/8KS3skIIPAFbb
6n3wv2k8lgr3ygSBFsCLpHoE1xFnxc50oeVcoq2YlL+8+zZcaEGo4cvm0ZXar0o1
0m9H+9tiOAG+zB98SIU3XratCoF/kjz4nM8K9GR/Z3XHP+QhHzyC22+yUGiziZuG
O/KmGVHXxBoDnNGBkXenU6cIkm6LVR2ZLrc+GvWp2zTjg06+VBQfl/Od7bjBK+0m
51GMRZydl2hDTPiwgLTaMQEQi6OvVsm+pKBI/FSGonXom12UyFu61wrIKCqTnbdj
36RJl4KIIh5VEmP+5LFffFpJs0rIaQsSP9fovkYmbcLx1PjE1oItBISjARjbZa57
NXzuWCc7lo+uMrk1LAbOjVEpY/HiP+9R/WXwJc+WTV48JV/qgfE+O3SXg+BNx+QX
WwQeKJ20tWmWgc70fKxuX9mU0qoQAntc3Fxk8pTvUsQ2wCCBvjT7CVhXNkGGZQ6l
AiQefD5oKLxYhTdDStek2V+TuwFEqdDBH8eX0Z7IXnuhvwp+Re4u6IaEfNDsjSPt
uBKmPFohY531ct5w83t5GarW56gheDp10k5XDr5nKRO7V0SmLONTlWGTSKq+ie+5
nl6OeKwFPg1+HOD2Lrd3/vas23iwoRtlRILDNnL6Ayg1Y3zaHGJsoia/WK1aqERF
s+egkwt0Kf8klrYrD0p4su5aqCQFM8pI/CmFLWdWE1zRLWDvuDSQA6MmiTdvQo5Q
I84oDqOXyojbU80g3tGBnHx2sA5FSr0WPIsxCI9vZYbEm03Q58Uv7/rQdM/NHRaD
Pv0ND4ncxbGLzkbGrfPvrL9scJL/squGnkN1VG+StVPh9tfyBEWvYvWjTnLhWHnG
MPcfBOFKH3NJcjqQRSZuZf9roY/zEu5lgWKAKciivvybkCdM+rkY3awXkkCvXajc
j5OJH3dSDLBqM6QEmZ+jEn7Aik6SsurBABcT90FLRZ6nLISmjJs9hLAGfCmU38/H
j3VZHCxeFBCTxvc/6NxWeq3WhG+Ga/Pm8FuHXiFU9KdshPkDt2RHh335EHtLtQsl
a7odyLg5OwbLfH/g2/0LUiP+Im9Y+WIfJYiGoDaBRfIUxvtqw4C8pO76dfJphda2
oh4XCOPh+lNKa69ZB9AbaRP9dXhoGbmY9T8hbqqt/t6sinNaxwPmiftCaL/zo2if
Ao6tKj2qXn9K69GlyXlyIsjHCj2zOPckET3WVxbjDVrRYHlpizX3eeX8j+i3mb1K
aR+jG4v2KfGuTYZN3HqNdLQrlwC7z8kP79FmYSEfBuTWudvmirmp1DX2i2VaT2XB
NlAuQrW1YQv+a6fC+jGmpzYUc65ujvNajMTBpZvqV6N4nMJp9VFyJXuXj8mYkHO7
XagdktZT6PNi5YByZGM0EAgMk5HOlSyIEbI4iPzfur6dEvLpbBhPS/B2Fh0kryXQ
qDYehgd23JWZl8L6myx5bYErYdOWjuSbHLq7zEtYxa8vyW8LKXZPTH98TDQocs5+
06bU3mV9jY0PJfjbBsmN3TXWm991OMMLU1ux1BQFq/gunC5ZBkdI7dUeoZ621Jtd
g0MUlfDE/0dY2+HvXuN3VisIZpXqstL8i0qXifZVOl8bkCegapPVxSiWZwg5hxmK
vWNoL1cATYfatJcV4+HSs8bOusC9M77Wj6fyOslr5OrPH9T8zR4G72Vwv6zLo4Od
0xZcl3FllnwjGoh1ywS66dyIJ/RxtLpXQFNcin36w53MQ9yifYAAAaifVBHSg4UT
Ropoa5h1TXxe4lah9UQTNE4wPvEAKg+dFOG7CkElRa7ebN6154GDvMXfhC9jovbv
H5GfxFPN4js1M4qFLq9HozIG+YDcsgGOzM3ECAYyBV8JzK8PS8euyNUsUHewkTBT
0U26vZbEfZ84XjC775Hawjnq8FW3l3Hy3bkvegideb9S1mKY0Q+e2xJqjMTwYfeL
APlU4ybT3M4ts4nmbpMhYK2FoEGNXmQtnfvjLv8iK/HwY6f8GC7Hqred1JesDmSy
LeK/+2UfZS1cUolOmpeDRM7xi/RlwR7KcaWiTowBmsQiqTxornUkZxw/K3Sc48Qg
ydV8KaddrsMDFsqsscKOhdJGbpITAHmzII3BsSHSPuh5m+N+j3eUo7HOcuVZclhM
J1cJpR8VpLPYTFN2jsAwKUYAzXZbusFBeIXMMdIryFqOiWHbJ2X2R79sjggXnVXI
rfiHn6m3t4TLr+Ue1OlzwEmGcJLWGUIK8ZM8bbePzuy2fZMn9L7QJeVRnKzHqPPv
8Gz+Ew+8NE3RxJ7deCrKN9FIlVwsdlLeHoAs+bgwZu+VxDfIe0zNNeHGDn5MAKfO
B+p/e0+U3Ia1S4JuxEW3/ymD8WXRWVjbVHAmcIqtGoiXGxXfPlZMJRu+dA/Il8Yl
BRCOVw6BYTRvsxYeP+1+Nm/8Y4aO7Xjn53UJ69nFn/XXlfQtZhNv9gYE6lYMbKJn
B3Y6Q+3NoLBNFvzqB8ENxmAQTGet335PT02Er5DuzG2BqLEhhMhrl3alAfnE51+T
ZF3jZqNj4Q49Mcr6OZtbuwueTk5AX7QHy9AcZtbkMqDbx4bjoomtUHGNlJMlOJbs
LT7ZR1HInczLERXYSOaa8rdGDIy2zcuPe6SXPl8laj+c6fZrYCRB82pLzTlnWri7
D+FpuFkA/q1jSm14RWhEenGCfmQlsxOf7cSiP2ATUTTWeC6jIsfMNnhrFIL7RjuY
IQTQsGsVIKr2McNn9JJNZooJ75nf1aYfoxUBg5XNOcs5P2mEU7Zr9npQ6J91hDQc
Aw59bQNnnQzIQtepun3GOY0WQFjTW0HHsZB2dK5wXmZx5hstc2c4uGuWXGc5p/Ht
T8RO/lYXLMIl8QeCd1hiZZLEa5M7/IeQOHL4CP4J8JH/k0HlOO/JuvwgwS/+di2i
T7XSu6s6LpiECSmSgWFoTtNxxRqpkI/yMNut+lA+rOmJocUxy6otbKKwDqsU9/Ne
ErR+Z1vDQqyUdAx4ekZv1vh75VkFYm+lZrtBF8pbbc2CAhh/+y1MUqYG8MbN/rJk
iJz8OqQ4wkl80q9j5tHR95lcM4ulD/Oeic9f56kw5QmhkprM/Hof2KgRUDEzLksb
31Xv5wMjNDQG5YuGroEdNfqowZ8I6eLecudyCmwqusdUKoEnrfa6BQu0XjGIOpjb
o20gCNWZG35Y5XN0qgh7Fv1tuV+cfQ6vlHWhf5NyR8LQqCDea7x7CuQDbBwFjHml
DXS6l48jqHPDX0rCqROebthgY00huSpojYmRhjzB9BVb+2ih249dHr3y6TYB6XTF
hT8QZ6iOMhQQu8fVx5d2ESBMBRv9b/qQ2mweaY/u77OJRQ6MiucnWKTF54l7ADhd
K2wTTVmRRmsD2rHw7l9jp0OB4kciVWq+VkPUwfRaY+ndEq+8XkNrFNl8f9jiCNEl
leB9FZQj3lpiwqCAylltxW3fnpzctTveA0Z+9l0Tt+xvIp1VzLBkTLDM8My8j7rl
v4jEV3vc6hD7P0Rbbf/nLznfavjvmZXFXdUpqr6Uw/fecYS4VNzIPV2cdUyxFq9S
FZ42qyI/78mYuoo1MZsLpD/Mrfh2wl2bLb+wEx857+hhR4DQ4KVT/MJxSVXgrAfH
sVy8m1JSDBvw8HOki4Gq2GxSfMqAew+738EHYXVxweYkuev6Pt9XuXM7SPNM/rH2
b+ZeQP33ykq6NEF4E9uEwGsPR8boPO6nTKCdZwwlikWEBCWr7PIqbuFmDtfwB+Gk
KjkcQ2BTk+ExEvoKi9MvhEHgEbMRRijHskogsFb6CFuP50RrTrmfHUJxhEZIEmRF
YUrl8wYyqAAHQVAEoFcs6Uqf2NOTYpRnOYCo65FfAxYqMMjc3mIw5VjQVqhq+jE7
u7itfXCFnh3aBBk+PfUH/XQElMpA/H5ZVaEbVWYJwZQC2TeLosRnMMR04VxNqjXq
o3lXARWy0sqadvb5FJojpvbFNw52GSoK5ANwNhx+amdl1EVHfQXpryKWJrplm8EX
DyNYlb9w6gnIZp32vfR6hjSGlMx0RapxAcUlabwtAcJ8e4/DdfKRA025ZN4lERs6
Idm0MGy7QEp6vfktkjwih3F70RIGh0gBE+L4njAcAR02NOdSR3fBDCoGRKL8J5my
OfKqB/y9n3QutW+6ahy+gI8qWgQcA6GWKaB1y+HJEjc2gjWH6v6n2FgqMy4J3P7R
V8jWO+EKuDfHlbpYeEapofgFyMP+RdgClKNSJMVaiiRKTDt/YqaVgEoNd7Q+J3eN
AUjCXp2Dv8Y6abwudmYHFnPekk/6ZKahosP1KHQirfAH7hC3M0rG5cW4uc7FGyS1
JTopKc+CTT40CT1rVyAeBiVWBgbrkfynbbLnG7o+iuxp1WlUAMPu19m6s0Cegumo
N5XamiG73uFPIfzR3rQOA57wkxf4ZRibMAUhD/MYr2QlRhGjp00PdkYjQxKsvQhX
k16Iaul1NOkdq9Tn6fthghHHrAHTaaUGwCEhSfBc9+taWj4qSy59NHvF1v/ou4fk
rkIZ70lg8JYGzj4lUCZ4M6t23DyfcA6lglhO3DZLXkEggdrSJPMPIp8PyF3YyOSm
33sAwVROC7V5dxwxFL0OVPEWn0LB387UtSBCFxxg3GackIp/imk7bTtOyNFNGGJZ
LTGzTmd19h9BiKXOrzTiSy6DGjjMpIKfqx5FSoUC5NDRn/5d2zI2WgVyKczxrYk+
zljC5vnJLAiWBjcmKmBSW19ft7lD4K/ndcrL/kuyPaZHYxD4qfWRvYMpJ0FEK2U1
H1ANn0L4UZpi7+fWKqso/4/fcQm17TgpBYF3oUT8BoKibq+LVQANgTeS1szwkE//
zPelYR939SDBppTuTWO9Kudn+KTzZPsZwNj4pY1hkluDHSbDhyIZ+qso9+zuVZS4
WqLeETwJXRAfV6i4Xpw89PH98jDgRSu7YIOx4VxGAaPrBRx2ynRum1PBnybGIpwc
1K0yJfUQDssQ7GTAAW6QJT2/sKUg4msrRYpXUIlLrikabXckeGl15KCOiud4Egv7
rwInfPIGj7FJgJKAFi59wcrysyrHe7JpsktMuCFVGitZuC5W9FzhfgLnV1ylE+vA
Efj5Er2vR9mlgmWZD6y49CZtIZ9QLs8KFg3SnIm9Ks1XC9TGYPw0wxdI69o5vjPb
rGSW8xYVO2I9jrHwzv2R2k+uqYfaqjzmz3s2FT7L8fKaOsIrXnbfUFgcK3h3ihud
g1PhxY/K+n9DpMjYFggdSSBfK41c4JDYadw9dYmDxqrv15VMwcLspM8dDKygjyfg
SwtNb/JS+8iEm8tPpxysLvLqOEvjMAAHiF09iK3r0BH2Nt3kdg5FBr3TJEIanRmd
DiyG2/2PfJhHdKVaegwhIvzAsM9xuJ/bFzhxbrXH2gK9oQWughe+9dJNjxldQGBy
iBNZqE/ClghjGC+intR5oZiHhTPknydynMOTqXPOUGR5cgjf8WXjKFZXmVzLnK1c
dU9ph08n98AMX5EfL/R2ChwmQcUSbS62MEI699022Dmwkfz0D6GuAlpnAGUvwzb4
cM313Q8cav+93uA/z/5h9KgWEJeIvZ5VvdPraauCveV370Ou4AYNVSFmOTDXCvbL
bqu/nIdxIRc8K0K7bcSuUB0vWs2zaeukn7Y9SKKOs0mKQN8r8ARsYMqip5FEdyvW
fqrwDmjB4OJHJD8GhRH/8qJFcUik0d1gK84CsBiYupfi9VG8IR6+dOGThtS8o1oM
N+cgGFGVmeIHunXKYnTDznC03UHaqfOyUkz9vLKI4ym/SgnsRZWwDOvVT9CVzwT9
Vj4zvCLv0F4AdXwc2NdZH5IN20+VqO4wKZEZFpO+o9WKTM9FhR/wFkzn4WuzWhuz
tS7pX9ok1eL6MOut8IItxNKcAQmSvlI0OQWTTwM6L6glBMwCkyT7HebDIXYWpmN8
T2y7PYJnr7riKhGvk1YO1M4h1dIJklaAFaZ+L7xQb8LgUUDP7K3Xhjs+T/d/gT6W
KnX0CB8Hqkove1j84GHHRsIVKFKLsBsnYyR8vFm8rkyUOnyK99Cc2F9bieg2iuip
PAnO/RjIVOCT8i+Atg+M3oFqZUCy6tA+IY8OAa2bWBX1giZpvNCfncC4hRGcuDOV
cHmJmfdo6+3wTDENsgPK4iERKDAPtfhaihNI8N9k4k0/0aF+QKw41Drjl16uCbpf
l4P1WPUKZ8rv2oRzpHwa8S1AMYCsw/W2dbWxMWRfnZCShXds57TV1ItDqugq7Q++
GLDylwf6FX5W+9hfNVj7m2P2wrdUtKxs3gnU6xYohtSLGko14X8LI/OlJk6PSJK8
LgVdpZ43gxugd6xzDHthU1u7l8zguiT1p2wLIV2/Bfr3qBOg8qNOqxjG1VUAdr3M
TZE7X30wtDil0Pnwj0QlxK7LfVQXCunW/lVXCNAJam6yp3cbOGw5OkK4L/YAXz4+
K1IupQWhyK76SfGlfkiYrq6rguqhNOOCrslB4wyGxcUTPTKGQghSpL9kI8uoLaMS
9qgtNa8hty1LrkS3/+J3+y4HyDiAD3Zi57dhM1g6ahrAHR4FVzXCvB+KMz1+/MdS
k58ki4mQVOoYMtaA6RIrXFnzZm/UJt0wiZZ6Ck2XcRos1Fbvup9sh2I0hE6036l0
OmX3WvX+kWdmjahwDct6y5qvUTF6XFQWsFGzu3qL/zWx7pnHanZNUF5Hf1TyP9B2
TEFPMiMoiR13Oay4k7soIepF5nz5B/KuY+4VX3dwhgG8an5mTEh9uIp0Kyd5ijKy
cPruX7U5uMN0ZapLK4QC+uaWETNDTJWX2Vzb8ZK3JtpLtZgGMwXJ8QIMmuAPlMWj
8xZ7EMYpsRl5+A0YvMIvjECwnu6p9O/be/1FweXNsum3ZjZ9QnwS0swAivKDB8s8
/X5bm7eMNfxp4ck1NzIsYlDvqCAfruCokK5FkZrXLZPn/P9zNiIApt6dqQPZPSXA
covXqCkoF78osSvEBfrmLFbwtrFMJVy7GDf1pr23RAKgc4raEXKMCJs5jzZwggWF
QrwHTdij9KV9yBHFbudFaReKjM7iZYxUQZVwRHkyomvgvs3b8RBnh8ITp247AUQW
MbV4dVCHL0cEXvGzgJffPdcG0b4opDteeq6rRNlqK2UgvPfzbMgldYMU272J5cuK
UB/e7MwXQtjoFI90ax9ICl3sQgvMdCp9PV7BTdA6S3JVUsaFPsy8h58Csv1lt/Os
0OSltnU0oMH+xkjwl2yENwqx8H6A7GZPwwMeXsmsjtcNRMWA9AIav1si/nxPvrSt
8+XIf+VIjzzLmbZ4KXljCA9KxSrrrVKMzoPWqO4Dq26+eigMizl+1wrVy8C2GA8l
Qn9KawoOPv+PwW+WI1xth+4HLLQXTm+f8zUgilNqXYLWaJj6dGOwblqXWc88RmiH
ze5nX1jjy8mBC6vFDvFk2hkRB/yHSQZ54DhmXC0wqxReg/cl+1xnaYgMMTAOBkJs
vJ0r/rUHvoL4grbQGBegH9zr5LsgEQMtuQj47W1nSqiiP6Ne0X4r83ZJ56dj3Qky
8DO4nzJDsAbklXxvVfbdvHXF85mh1rLEmczKoldx8ualFnk7H0KhqumfqYxU8BXb
4DHUnhRPisEnqL8O0zoNvXvHkfjSwJADC2gFFuwyrnVsmgsijNg6BWKLPi93TVlE
dPSttsGQYdbaI2liCB7G+2t+R/0cmXhaI5W83M+r8pxmXv+U5/LzPNST9Yj6n47r
DWO/9OJKvORQ+BiXPuARTaPraHAnouyotpSbEdDvVDp3VW+/vlh+cmXK7FHfOCL7
tgQu9pKXUecC5yeE0YpC1XS/wWaCr3cKjDcfD/OZ/xnXqKuhicjqls3qb+l7k9wX
bpDbPoWCdtQ92J9bXKCKVtq6vmjg33yI1XuPiYm9V7WGAhLfzYXbVpKoMroioeyd
l0Lu9PD8S/raJijVeoXr/jqjF3tcIPqE6my7RWtvzIKQp7D+Cudp/x5jkPKZh/WI
/k5zmI8w9y/HIUKGAHOxNM5V8ex1Brjtmg7jNBLeoIZlhtj/aC1HSVT6M2Bafwbh
lcrI8BvDNyLO4adz9RSO7d591q9NAYjp7BFOQ3iE3a46Fdec+HvK2Jqi0CiByj/K
zaQjMbur6TBr9EOBlwysGnP2OZXf29kGetAWut6Dw5ApWoQfNwRWaPsl/cVzr2bg
BaAYydzDLoWRcvgwPMpBEMhxx4je3WMLabWqYM/Kq8aQ/gNTExq6mlx56mHnHFLX
vfiveY1FhvrrAch3qcW+TcByXiTyDRqOyQqZ2xdKKYlj5t3/w61Ykpae1DHGp9wc
VTAd7ae7WnSYXM0KmFruZLyMD70iBe9+4dA67nGBmUUGHt5GGARVtLWt9X77bfv+
VjRx69s8qlYIW8Xdx0czGdf+ZgwKFzC+GT+sDLYfPDGv9vowV9gots/uRUqfiRLR
dkCX3AYmeQaQ0ihMdv6nPXnUhiuP/Oq1rF5dh3NBdkOE0ZVDKEY/hu0iwhwvR5r6
Vjlj1ldffe486CJjKXMB7qB5T0lyhooh8Y8kyKw214TzPJol2djnLs0x2Cot/jFQ
u35HuaAptoOXpSt4L0IeeRRQE5Oqw4UBR0VkHTVWo6eTYfN9mz4AX0toAVswVdPh
9ifGEYIhfXxGHm7cdsQKVj6Sr/gbQZQZEf1t6nZv4MMKaguNio5nrhudVFFCtviW
vwk3+ZtjpdglfLiEsYx5YDF1HjUYff75EXal0v8HeczcQyjTnv6sVKQlb0ylqGZ3
HaFqVM3kZMOuLPuc87iDeyiwz8HkuAPS4t7TIIhuGciu4rJaZp4AzJX+T8Pi57V9
UR9/BWxiGkEGe8U9RLXjWLtm06Ap6V+qIH7jjwVliA3kz39QKDtOWUsrGxCBgH5O
PTUgIU2xYuaZm2uOGS7FzjbiCAu/KopKPujRLFXAG7+htCgVAPdO9OpCg6TWD4sA
qGlyr4Z6wpaH7vHFulmiR71rQPrSXwLPOiAZM37jdIjxPqgTUtw+LzJMT+pZbGvT
H12INETtycuQ7VO5HU2pu4VIimjHaUeaCxby1y6LYponyLVlTsyoJFTg6ui/RAKg
jiWMqCC58CZe5WjiPlYuj1DODwN73F1Nzf88nSRaVh25FaypQspbDeEKpPWnJQEL
Jf3jXCwas4wrky6RdIl+mugBcJFyIuaUHPXVjlOi84kHYAH03xhc0i0g0lJ7MzgL
b891HWCIlhtjCWTcSxuvFxwumhE2Afq5ruRi0YjLy7n+IDJK5G3kP01lwTbenX/N
gNSCEhqeWImZzlsgzy0dLmCMElzoVoZm0mVyzJSTXR4bKl7CyQ/COlZYtSqyO9ba
3VsPaTyRMhSPOblCQ1VuPCahJ2iASI65AGcs04LCZCYEAGD5BeDKPBU/Md14MBjL
pGnAnXMpYrkJ0HYONcMS+A==
`protect END_PROTECTED
