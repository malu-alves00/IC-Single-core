`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ihuAnEUPQzD9Ce/vdEk5jToDBC0Xl522r7WA+1qLWdKKeurCyg04Rhnwmouu+9x0
eC/Nq2pTP3fJPqW7yr1j96/kjrnepGUN4bfk1iy1S2uvHG7fexld5V13cM6rc3db
joDDwMqBl/cmd3Ppaa6Io8VQcx4s7efjUBG8eQoqvrw5GZ/OaLpYSr4X4zxeyWR3
/g/rs2I3kC6rlcKiKu1/Gts2sADNUX+PoPDldCQgN7G/iqxqY3qSjRB7SG1kUyXp
JJaa4+b7EoE+b+5KEG5mhGfVnNFCP7v8rnqz4zqSm1EDPbpNcyPIzgCFsy7jIoEa
QtrhdlXuhCf9E8iGtydVijwXcVa2j4Q3TPlFrD7bNXJPKCTK/MNOvf9YMiQo+7xZ
WIeHYiEjOPRN9ytXKRI4ZtZ23doTAvbC//BTtt2T3c5JGiXrJU9G0UF3CcPAeKJ0
o7jLS20vI2M4BrVn5cxS5hmbyPoAdGlP587HVw3KxjELmm5LptzYJLl6yV06Aruh
Kr3NzabJ+beqXT5OWKEvpsVPgXikSZTJ7SgSabNBe1N7shv1Je0ioydR776inVv3
rL+RFsTwYHJa8XzhN+R0GVDUSv2ZZc6DwmyMeJWklh3YPIlksZPlTtmLfz1u2REp
wjYgkHrU80T7X0FM7rYXR6SkvWb8GHq0mBi/2LB4nm6W+dCeoRAFdUQWD5CaXNAQ
/qbFos7sbF7aGUHe/WxIMzLYKY8/315ShCq8yf/jq8QyP5E7VM71n94VL65mdkja
XwAeO30KFtUBfkhyCGG5XaUrY7+DSs6whYl2to0WV218Undur2GUGYGWvV68ZBja
MP0kV0wg1tOkrukH42JPTq3bROUvWJZ4trPYxBBIZX/BJAhZ1OI8/UtR6ajLeRXA
ZkeQl6wg31Vm4I1ufZ6Wcue3g6mKDJ+AHyz2GAx8Ib3L861+WvlBI618epYrwSpQ
l6Kz+kxoB4AD9yExzTdZxKsnN1Rp8+VxZtBGmc9eaV5jt7BrJj0ZXtreQvqM7FRB
B9jhcurk6VcQ9KNBnuwyLkcMcMm9MILDA2bUMQayUfsfgegpKK1J3JNhQGX+cjIO
sILIz9fu65b4qdvVTE4/7ejDAWr+W8dIBB3OC/oblUW/kfiBpM0GtR98GjYN51E9
OzzUGVfPnFjN3C9iRK6iuO/v3z5QkX+Nt6s8XQExD+GLYwuWdHgGy9kbpWD+Qxj4
PDIiR2xHs7cVowlOnJkgPda5KAilfvL6zf18466rYqtLfWd/eNAMApMQF2ErOvk0
ENU5eVSDsU+h3qIOkXLgnjmPuXf5psWff+qYsetkQOjDZ4Nl92QWFzCvAL/swmpy
jg5XTNXeA4G+VEMku7N5HyrTQ1x9DvuAy0XV0xJ0vhegHbB1aOy2BW8/EmeqdB2d
V6C/Gi1tDQqqqxSvtTKovnUUuyp+HGQ+vL6B6VWYu2kK0sajLxRcySWdcGsNLdbr
`protect END_PROTECTED
