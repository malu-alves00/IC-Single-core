`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Hx5QLBp68c1xROQVJBEenEOOdpfDzYg110fEbBXDVugDaFr7PquWixZXHlTxCrMw
8VU4pMFFmwwoDFLBLMU+lEWeHBLpx+3gcoUG35x1/Qjc5pN7X6ctazrAmiIN1pMT
cDy6TLwMppCRijtkHsSYgE43coH/rTFv1geBJXCZXz4dOi/Mv3F7kgCpgE3LdKj/
rwS8zC9f9sZYkwdzJAVNWVc9XbhXEtpGBHY8AMfaTfV02qGvs4P8lJJp24mb8T5M
qdTvZcfX0yTpUQS9/PDESIIhQsHaL54R2enKqPulUpQKCuCiBprgg6Z/Ev3aQDh/
shVesXawh9GEbeZraA6SmMuNO7ez9xOzGjMmB8/z7boBWIskbgCWNF5bfpex92x2
1LvCSjmh6ZCvSoA5w9nLjbNyOj6uCv4RG9Jgph8Ttj2oJxjv/VP7ekal9qEutc0i
abMJXXWerIQIoHxdvBhgz6HScW1bVpnd/GxnU1ZV7yOHSm3A8cqQtnxfJXPW0cbS
Fl0w4dy8/bohx+yslkDRbdyQtdAnCPp6ydL8Q9P9GVJeY2ouGjvre5Qtyt3qu2qL
8UfSOdCPLQ01+NSsauE9+L3RgXNcOPYp+mabcY4Y9E3wdKYUI7NsTFZUSQ15MZyH
1HYRprLDfBLHw6OdN7IZxOT28pnueZICJdUeYL2WNqG7mdNxXgC+sVOqEX+3rLCA
sDSXHP5DLsWJ8AE2VQv+iaxmd+TChrkdnNxy3F2fSK3HnkcMG4kvTDa8NcDXKXKG
Oa0uu++2UAfz45JM5XbqQ58ts/3N7wzfSLT0zzC1va6lQFbx6K3Z4JZg4LbTQy/k
0iGd0o3P8OZ2wTK/8mNoCIM726gLIjNXVX62kOJmL+xPxs+zjCMhBcKFvSTTxMDl
9Q3mpt8lhVgMC8Nqc2Xx2tvAmO02fAQeOjc7SFIkbb8DCaOMChgHstnASgX7HRHJ
EUWMYOqPM9r1BXracAcx4ji6EhQOubsfY2/JbjSeHs4AB8Sld7UtStaqUyaEheJr
sI3vWlTIghLb1HXJpZqsZENkbyvr0WM9Jg6y+tsgf8EpyIlxITVwnqFY+ZT/8JKW
r77BOvBi+rZ43haAp2fSqe7eQJsdqA/HINLyDaXvDUNE/g6nTKdYYxcEhNCSr+C3
NTIDnNIrkNbWUW0fhCrDZQ==
`protect END_PROTECTED
