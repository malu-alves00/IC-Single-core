`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
txYnwJbQLwhH2pjrlmDhIdekcXgs8EUqWnRArrFWr1umkA8tyFcNpZPwoEKPuwuZ
z0ZrfFJVP9CCx9OhSAdVpUuCtCI8xharI7qajdqWFgqo/UGDeaumsEB78xgLGkf5
YXGR7Y2COM7+800GffgKm2nocYe9Nz3lnUzbXH4/41xzR8mXgnj1BkSK6R1pqQQA
SyNsgYnSulyg3hvYOzJFRhL7MuVcc3zwGLhZwidV+7pEET6jsSpQ6nC8Khz7Tsiv
JuvPWLlim1A2J2yxMuymXdFeXWp2Gv9GF137+R4XAJWJq+nZmwVaB/9Any/2dr63
Ab+cXD/mto11etG52YvxBk6TJNp4Xej7hdD6kYAHklgs32IX3lr8+9g0eWfS2wyJ
g0hqq0vB48dt+iHyXYSgRr0bkxbGWxo53qmOH78amtDtuS/BxDgpJKNR559TMEUU
J6C/F9uF8ooI+7fGuVq1ZUJLObeCnpjmPggaPE30VnQkjDKe2xxv0kLbEaKG1ED/
lqn0Gw3vto5Qv0aA/yBay0fDxGUIr1maT/SdrUMKrs6uDvQJ3HBB3wndzDCsKKly
0uM0U1r412pf6Nqgq0g80uuM19YX7TIshH45UOMx3uSufbWK5+JOnq52ioEILYpm
WfyOvY3NChpF9obsqLNtDLsNRRdbVVJXXYlt8ehi9dljpoXRo0pd57pau/h692rF
/igRl1HEXg+RTZM1RY21gAuh344JD+wtE0nAcyUzXkaCX2OEtAwa9Io6W05Eh10c
KqwbgBm2tAQrolJB2MJeYBv16eOxjgKRCTMLUA1kkWsee0e2J9DKlxfUPE0JzbTU
F0plQgto8EKHQ/qGy7VkmUpl0G6mGh9oaN5XXqAuUry734m0FL18xACz19KwxbN3
dJgAFGxX7MlZH7nbBZvK13SCvELFiDeeW4d/ZYzgVimoRJ22ou5oMvQ9+hDpLGQF
8YrXIwrTNtZWv6zNihOvrY+/cUd63eovAbFDS42v/NiZBFpjB/i9Bq+ynQeIC2lQ
8ojbYTaIUhng2WPdXnANNZPg0BJ7+PRkuPklGv5z2En0j+cUI3LU4KONNXadnxwN
3HrflhI/TzvoJRZwkIeLSUdiwT42fM46/6wu0UmMb25kI4LJj+mXnDCELMYRmmRF
iKSxVdiDxQ/WucRUUGGdN5zsTB0eGGvTFfrGQJpqtyWEAhwr+V7pqKTryyxpcI+x
gXfG4Au3Dqg+r53YiGw5+Le8hsLPE54BwtlAlesZTfmnpyiCl3PH/Qj44rpAaf+w
jH+I9OtNQOLxFR7YhSApwDj7NsciaWKQ4ReOL4kU0Q+BS7VO91UDqZt1774syfHA
pcxxMS/qyfZp4NdkoAhGkHD7WkpmuPDDYpeEYC00IfHRv0UBLahIF5DxxCX02f9R
bCb3kGJpTSsGAFWrcZ4SFO859t4HZvjeLaOUlwLz0QdnG9e2dT2+y8qOmtOEtKba
1ZHsRnn95jkzUlEWLj4klPRYNYjL7HEVT/4z9NMmrtJlHIBnTfspidScW3VnBchd
3Mmo+s7SbGovL6grqWoZfTmVv3EzKXFGTfJ7ul1+nxHuILNSgnY93wkGSab5Yk/0
jHHKAJ8T4FGlVw3f7MpuFptru+VAC2JVhRUzpf0RGUWrQ0ASWDjpwRrPkasWCUO4
0swZCHpYFCS2eqEzFTp5Aw8GWbEShut6U3UtwAWs6J96KokqQjjHnsPnH+1B+KHe
5koZZo/fAVcPEGICBHFL1kZBUDRcgRgJWN5KN6A4dHr6OSZQkGXrgIyqLjOs7Y7g
jU3lIoTfTQqXYDXl4G7hseXj31wy+dmb/wWoR6LVTyciSmb50Lu4FFTiQbW3TGyO
HhuGUeCZyFhO2LxZeTrT7xTIXtmkGB8yT7vCwTkbA4xG7Zvf+MGHRz9c8yUwgHwz
fosw1m1ORODU+gic3g28rONiKaqtd70KI7pWvl8+gG4b/HhgXOTWYZCsv5iTMh50
9cMjM440avmBVObiGWsUH19EnhH6TIdTPSRgVsxw4AJlGM8+S9uUxUwxj0kO+ire
USmNEQgWSC2O/4V1EsUki2nhCz79k0oZhvClG0dGhiU38mOENWTmarmMrPP9qU7s
1n1VIwFrPqpG66uO4GrFsvKRtauY8pcMw+8hO5bSkAy5emPgdzYP66IU3Uulp2QF
jUarS7TqtxWWbXGM8aPBjW/u/0ezUsIL4mXivgTSQYkm0ns7lHAXj+KmeIQc+gsm
N00zxLaDySk9w8LF3OnLiGeS1sfol7SeWhglv+l8zrlQY0b7arUGmPn1O76lPyqk
SMBf+I1g4K+5jKF5foWhARh5mhtKmN0IVLILc13p1r/JuF0fELSxp/q4CNqLKx99
Lq6psawOWxC1g3JFm130S7BOp7aIPEzHJpf8zt0K3SO+ctrSEe9LJuxYOYiaVf7o
FgOMoJ/3aan4ZMhN4wTu3hKZbsmDs7JTTtUyVLJru89EyUIJqRweaYSt4ASRpcHH
7ZFJNW/Q2pmDRUNQmonJye/i85dOsf+7dhAKwUsSHZAJGdKUlBVokrBbTDcwRiQN
I64sQALPqPXNP0clEBQTsVOVNHEr6yTN0nziWJamxt4uoROf5q0eUeb9q7sTyQlv
4fvody9p6q0DSPsvqk4EsmwL3cmvyt3x0AiZC+ZEw/USATWUamB8ESEwmKO/5Qzb
wFaS6i1E5edP0iI+vb6uMaQCfgpfDJwjqbE4stDUrhJ8lBRBnI1Y6Lt648vluFTG
9AxYstXri96ElLmV28PqVeYdBEuzj2LAa4y2OdptjxcpVRdp7kBRj1Coqgud3wK2
6fcgRnwUX0/tEBxXetyvn+sfNSy/o2VbHfd2oRX5Db3g3c+DpeFXMSQYB3XAOmI7
zG+4z0uJYNqvnJv8tdRAe6OWntFSUNOiJ06cO+UaOWdAihk7qFjw/G/oluzLkOdc
OQMN7lvRo9f+vcz1MaS654PWieHfvgyWc3TH3A2x/PjHi9LRux17kLA+6KIjX04S
rriD4PVdFKbdaCOlmOoCIoGiZZkKO6rMNSIjFQuoo8KUx6eAIK/P22U3XHNdslj/
5fx5xGDl/IASod+cOp17kTi8O4gDidH/6n17bQvR9ESpnWK8FfuGl0P/0qnvrMhr
72mQJeTLcI2mWYrAsPCE1eeeTN1MFsSejCB/RtN52LzIIKM1BsT3+Fg66JR/CJed
+ZYNlGotcpftxfmnVwS9wcHyQu2dkfMTYhl2p+ELTusglU/+JRBIsBlRvzW03NKO
AfnEF/JNrzy+GgFG5/c1hpPgS1Q5/+6sPylaC1Gb1VlY+ZdXIF6TzpOHi2QKOP4X
cRhcFK5jP5PND5LkKX3G7fTLHAk7VoTw9N690+bX1BmrQIslxAsnzNWML8B+rTtb
Qy4cMzxMuQIo7CWCXjTB/iN6OS9jyHT1Pfn9eIWtF2bH8XbphXYLQDK/6ejNXGqp
B1K/geO7ZLT8xvt01BoTQrBrpsKeJFtDGLwgduSLZM/DfkmpiLIlIOM20qIs2s7O
0S9nvNDMCtEhM9THkcLWk1hqVZXPbNsa8yXlnSYdvkx/FMc6tXdFWkGPTyw6jqWb
E0/dJefnMjvozi0WD4/A3sEkQnn8qtQZqsEqSancF5NzSyYtZVs7IZJFlRZpblCu
5MHLI7heWruC1o3CgqbcGgh7TRuG3Dj2lIYbXJltcTmAmlt3R0FtfsaNSXQl6Nox
TXOu644aD+1KgIeSM2RCqO4OJ8Qy1KpQiLeYEMbl7CNPD1edZEW1IGY8TpsZSCcw
r7CryGq7SJ5ohsa6fzkHU6sEeVx/ovrKxZegKtayRFJML1HBmK1s/kKvI7A5roXo
aMCzzJIwtMF29rTLPUbE68ruW4gHMtmA9SvWwWN8uAp43PbPw6WhvkNSw7AB4h6U
Ecp1fHVnW7owx17BrkyiWCC/wz8dei0ziRQHSjFOSwx9LWFjWtvizhJvINJx+iuI
gnm+eGjGRXkKWgaWMmJv4H92tfy9A2/POiHnCOl5xHEsobLlnDdYFRn5WXpmMJba
GqLFhBbB382lDaJRazfh5THz4oGMDJ1EksSJeWq3SIFBo7Pq/miXjDlTyoCW3tgF
qHAuqEzgTwf4ZNzMuX0XCDdfuPL/na41OsZzUxUh2je0NLoilO//0d7kFQ3UBSaH
5dhL9XqWYAXMPi3zy0kDsGKpSmbdbaqyEwNLPIewr2UkWwk9wC+OqQewaQOXJr8L
buGJSjb+t5FFksFgh4goJBwY+GjxRdYZbl6ig6NKkWAG87xJsFbIcdSsIQo6SfQT
JB32UB6HG14HxwLykTHVKKIbQo/0br6qjIG3dhEb0i+zkjExB6hArXad1r5iJGZH
8OerOwiGXPgMV9d8aiNrDH0Z68Qo7Nh8+7izggvVuxkNOtEkUSitVfyuwnGzhfHE
y5rT5JQ8RRuQm6VVi5nUYuRekfR6tG2zlgpy3ApY+QeQkZXmadNc3vL4kEjsNDaK
VNkcb39twgA7s1lQ4jeV2KAYhVxZdL0/FT23zmT0Bj5f4UOhKcaNuLrqukHEOoh+
RJVx5+LYLWnv2Mj422RQ6rA19l5Q9MbPDzvHzN8qIw/OC7w6yqpoipsKiWEQONYP
JLPHND7O0jaVUP0JCl5LdVSh1ELH3pAALuWR6QUiuJWT6bQM3C2pXc8Zwod9ZmgH
tj8BRiPAzoo3GbdHA4zrpYWWl5ycZHRTd6OpdZPNFZueDUA8+5tqRVOFlaZUVZ8A
FFumScVrlFzxKPkmexm8sSEaeeQXU7lMZua7QfNCEQUGZFsToU3jLqy0O9/0OfLz
wKhQokwGtCfT+8wlJIckHmAi+zlZ4AB1rwIwYWE3uPof0Wo75ctedPvfMJGRlb4+
gKbz0hnHDU0Wja/79q5L3eEypB/P/609WuxVbwVTsc41GbGmYcziUt1A8/ts6x/t
PqA8Mwa2fnxlqSvMEQCCwUd6PA+IpjzT84QJjfiV2yJ4JXhynU7+kw8n2DqMjF3s
WVhlYpTl3Lj+QYIATzyHQYSjkWFZCye8tOPM76KjTHzuYkjD/u37pZkgS5ToUluH
wRAXzNtCGfm551MCY92G+j56xLsQWZ4safBNGveA7ZqhGz952c4X8PLo2mdQgBbZ
wNTaaMrOMw/qWuq5ZQnAZ4P3lzMGpWbfNksDpIgnegGB1G53SO9lI6KFtu4hRn8B
asw+EmHCBRYGDaSw6XUIvFyeAUXaR77HYpl7fvx+4UDtbiRfzt7tWUWgQXV70nMU
LSqE8bZNTsaUCVyhXsk3HVe9FPlVUjj9fEEsVGIxqG7Y9gA2KD2qUiqpwZQdIVPs
gSDOIi9Dm6ZBYbZoTmDbKjcynviBQ69tXZKzU8dsnuW5JIkLmof0lMpK/ullIfv/
j3Cvs3aGjrJ4bDAnaAZ94X2eaDO2HWLt9e3ajb+dSrOCLm8bcSZsZNuBnAUbzwO8
8my/1QYKmZq2hECXci83tl80JHpzA3HeVfzlkHLT+Y2YbFvjuXJN7w97ltBXzTAp
eX5moyrej0ZRAKKtdlnhqtDU3kegeyEhvrgRaleLvSCLk5CTOMeB7oeZWvZMwUdB
8VxZWXk72qVPE5ZXJfX4jqacNSikhZteKpIc4d85fv46HQflk8hYffsUKZVX0701
vP5PJF7ICFpfyVJYgBij+a57rLD9A2krRjWCXdfMVGuCM3wZ2ls6k8QbE6SchrCU
1INMo9n+BroZvwtcO2ZQUmq1zRH4+KlRTkDXCFct/OMurUdVXEx/nfhljV9flK26
zkN7T2bkACxEqxmHilP5I/6BFhL9c/gjjIg+4ppuPSQbeWXne4soIKuDvPT3YjLM
Zxz4v7lMHmLNlQMsybOthr50gxpV82MskWauNxf2Kb0JXZg1qQSXupaO+m0oyVOW
mwyttY4BYpWI1VCwXqykMKW60WbS93geelC6n4MhJzzmS1InVxC2sqRaY47Mlgip
0TT2MgxadFGgEwxSu6gl2+8EFdE0eDjRQbmghWMoGsHDs84Mj+eO8wi9bjMMs23Y
Civw65CXOBfepMN/kUzt1IUOVi2DPOpl8eyx7taP36XuXJ+uiYnzH7heBQJDbCXO
ws0sQooeTCvxbF3vg5j6G2vzA3Rgljo0FSJtKOSVIw+LOUMnlb6Qq+S2deutEn4D
y52vGeHXeEksiq42qCt9Hh1uYlhEDTEqFtpcr7/IodtyBvSei62w9qb8pLx+QzLK
MkP1BFZNdGT7Oxuc0OA37ILybbyY5wQxpBDwpyfx6zSu3InVNggpWcL+gTlPlz5D
7G1HZCDcSXTDLIN4LlMNxj0d0IInmQfl99Kt7zKpitIUoEe0ycMC7yem7PhnnVRq
Q8epABfPFSGtwHOPSSGgBDyNG9E2sQ7KVZd31DRQj9bn248lW6L2P6M4LIYubgUN
cDjM3YBp6OV5OR24x6bobqhym7zZ64KJFR91UUyXk3mqRLZsGX9UFic3A/Bqlgxs
jTs0x3vnlu6OeWbFU5O2JP9geNXNmoFzOf0v9pomT5Z2t2ozi2UU5IVFwdYcMdUI
`protect END_PROTECTED
