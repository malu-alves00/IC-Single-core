`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
R4XcUjkH+x9YjK4WkY5YNg+mUo+CwC7CiYfJyTlDkollUfeZ56hTPi5bOKHinpCF
Jr1uPQCm+cqJPEl4D0K6sFVEiJMSfjMGdjgNtMk0j8OFKJVrPkfQ9Y4FLowIPsMa
iWKFJ/2CWwWalmt9J2ivyuqYCGXuoPN1oljdG+4Om4B4zY4X6tWHrweRq5N2frBL
BnkGlEAWEqSWKl3cs9Jt0nlb2VWpF1s7JwMDRyo0zHiKGvbSwZJs1cZbCian4GI1
VzpAYoVBoQ0oHD9ArwohIJkayvZmfqw45B12AQKVx2/8mRml8yfN8O0YOIG95O4O
S/3LAKyaznw56W4Ui4RYSR5CYk0l7F0965G9juLx/5N/33tlTGeJAv76pkzUuEBD
OwP4xVup48gnuNe00L7MmraoTMY0H3zab0TG2uupSYeDduIK28Xk86UFpLMwNUEW
uSEz407pQXZA5TyL02AKmfue2uWnGUQR2X035gxKQjuk2wgQ/rH5OtD9uidKb+QL
6yopIN2BZTUiNkQA44qi1y+JG3KcYdaPc9g+DgQ6aAAQThoT7OeLWkMFkIMcV+91
ANp5wJahSiEQZURMwOp67Zjs1b9zTBCQ2Z+lLqDphu7jHOAgKtZRMBgDP15NHdIW
rIjoV4F/hd3EyoO2IT4nwr2qJgQTUgErcfTMO4nSl1AnwWXYIRpvTuHUutIKZ9sS
SBOsgofaHTEi9bK00pE0qcix58oqwZZf25chf9KOAHwv9wKNiy5GJR75UF7MI+Mj
Sr4tKlgZUqCF0n07v3vCGlzc/8PkRpNSnO4rZ053hjiXs5xegxFOiJIrdSnBBJtR
EbdQL8dYLTJsNc0rsQvVaeWa3fcY/g/TdHnXdMCs6CY=
`protect END_PROTECTED
