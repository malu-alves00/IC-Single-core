`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xR+ST86Bd3mMRrLdDdwUf8Wp7cmqGU4ypqzwf1ctL5rvrFmsLTNNsJuOZ1Wp4C6W
8leYS4eTWVQeenXjsVSCs7q2vlhHTfn3dczUfSg+hwgojMC2QYPNdTQ+LeFxSndY
V0UjKCKLZdcN4zqjwSLjg+re95LUZWDme5Tmh3qQqjQGUNHbiW9ErAsMCRu+KwzK
Hipm0aoUDSFWHKSOqn2glIJ2NTFpruS+P5En73+tbXOUu795UGjq3TPdhf52hWLq
trVOGY2/W0j0tx8De6vQ+LcQb2Bta59ledyDA2c/inOhMYTbBN05tqOS63lWujXP
9VZhSzLvro0kFCeSkRWJ6zhJxsQ0Sof5+DbkOzS5+3MrU5ZpWL/8b6HZ9ZcuhMy1
5mP3ksHUjRQe0rhUTWXx1OfCtt6NlX2K6XvCcPXDUNpx/NAZCOfszNMdFMyEY0VM
Elkqj3yEZKUHAJnJ4Q4NtpRRXtgti8XK8HrW0P4DyGu84Osm6Xw3mxLVdNxc8zqN
7TRuICIWHDJcknRClvqAIzrNO+IZ0+YqA0WWBf57Buc+ipfOipgHInEJNCh5nnld
8Ylv2H++8dA8T3INVWmxLqx/VBg4c4gA+LGgTPJAGl7N9Y5w7ykzqUiStzCt5bYe
N+Q0O67ufDfLf+LoolPPXEYz1BL9D/RC8RUVCeNJvtkPFwQnElWcar26VIcpiG2X
qsrNkJfGZyzMbLJItffL0f3WQ+vBactIkWfOa4KuavvUdFYGgwhluW663RgX5ERO
cnjl93YW3+F1h9eiHVjlN/buQAcMaOmGFdaCqbr1GamaySGcQXhl3ospoPsavBW4
DlYfeLLy+NPYFJAcieTYJppLkmcCFjY+l2QoEWrIOI5Xwf0WI727dcyMm/GwM3+c
C4LWwp0ozWrDvR8tV6Tj1O7H/hnWdbEPUTqJoavfiygbmJLZYlYRkFcZuMdijK9L
pxbxxOb6t/F3t0yQ0fTr7jhHOImdtPg7dWvqZZj3zPNvpX1c3ZixkHfWArK29rNR
78BPi43j53fVBgTbFyZDOr4jj/n+BM4c3WZfddUNELFxe0iMdoj6PmBfwlnAxpqb
eYHhgms74sC29aM+QgPDay2SwhuPlI6MS5qYVkdMVNEnJjjgL6Zh3B/mn3tehMFM
gxWFod+L6ZpnktCQ4ye8ncIxDDqX5JjAtvjW11tGGcCqtReMaoMrms7WW/kEvzXy
YZf2OkzphuAqfGdbx7eJIprTiFuHnhzOug8Urba+PYQKyEwBYpNawLnmXr5vjoxR
wuyWvyRXtpbfGay/v9Tv2KsVuwAl8iEkEf1P4vbR4YHBJi/CJcCapuI1HPjuAh+8
C3ZgA+JHCjTnbM1uTJU5ys0YknK3o78PDad2Q5/yi8QAXwwzqVvgpg3pNY1Mcf0l
oh+dg9hUWzf5Fmm3f0nHPeHVPGN1u5ISLh2Kg3evtlQRS/xaL8heIkx0b+fKjnsl
qbVQhH9U0ehBZjozCJkm0cH0jxQa2IjNF9n2p15uiEBeSSo9G6HQLMVtCEhpMPG/
QnmCKqBf/yYUJAf/rDJL+1u+L9QqsxZ6+vcvcpxeS7l2Xj7uuCFsu9+ugUwm9I/h
oL6DtBISf7IIC6NMBpGxz0ujgJK7ytDuXPAflzucvGYVeffOogCwmrpiKGTUmL94
VhkRWqgVdTCDRzbGQuf/MJXafgjNzAIAD4ceukcabMG63FrOOeH+1u+SiaZhjAX7
m46LGbm6wAmHbLOd7LM9eZh4qYyng/6aI+Xjir9+Ae9sGv7rBxE2PtUbOTafmZ/Z
TXLr964TEp6xbODzLlqyiLdqJsWEf/+yOLOkb7l1ii+QNL67K5fOt33L9KXdgPLc
nRAPJWFk90sZRnSvA7/inlkg1doamWWIGFPA/LH4oeXPqaHtJJrPHnotVpspxRGl
3H29Iw4ZTrg1nBvnZq8xcNNKQyiUX2ES1l6SkyNmve2JidSmH5SOvoYocDvzL2Od
2A6zuNCd//e49JN3nZQhEl/1gVZOg/gvGTPaKKOUuqxmsUeA9fo8uSPzpxlXG56S
5hj0T/HWU3lIopBkcGz12SybBvKl2RBjpDTLeyJWAN1UHpKaJQDWJu5fc6iz/xom
iNgRGxrFqncczPF3JrmAvt+1QtqzbIFcCJPWDE+nYuKyk0wfV2pED4RZX7NrpPQb
zB4nJiTT+D04mI+8+Ik7YvOmUAyQXflhZWfw7N7rWR4U9/mDZ8lky7blFYaMH2Yq
wdtSCPeyWdlGWNFwbzCJo0VSEY/tvB71u/70e+eChuLRUC2oK8/aSZjQTJwyDWBm
L0ePAZSqQ7j+lQfyme9lJykOHinrQqHCKD/Ct/MR+KLYsVFsHOxqOgsenZgdOdhS
Gbmh4XLGH4EoQV34EBPKqvmrg+NLW9lqN7auDdgSLNw26X8fDiej8uQVcXiez37D
y9OP0qeHrky9jP9pdHMUz/171CbXJd/6g2YQ2EEt1RJoB/LTcXQX4LBYGXsjA2cd
Gnwa4DPwA+VTaQJ9lgXht5nZUMsa5w3HawtBUmQgxztBMQKN8vvFMiBobS3t69JR
AOYkchAisQs/JRTXSczWMnsbkue1hBHmUDpEkMTLcF8bGA8gR2eRwLB7/OaWEWDh
OIR0HcBcJhesZc7jjiDYdwJGkrvE0KNNFDVzqv/YMWDLgS598VStErZhEXjMxrRz
1mD9EToXVTaIM9G2UnVnLuq3iEoQuYAm72ugrQ/4SVW03Xe/ZgpJ0sMhwRJsRnwO
i/kZbiRqN8XFaVIOyMeBcdHeck/GZLNRj4r0qBVGbVglEQzMPSUWV0MB6AlT1lAZ
dI1A/csoHUOBnvFOFtnf7J5ij/p5G+u+DyFYOSFhjcqewBpCCjeKXsiUeFXp2j/X
`protect END_PROTECTED
