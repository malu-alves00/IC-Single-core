`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+OQy0d5CRB4wfvInL0uNtz2kTmBYMq9XBimeHsCy1iAWqLeWr+a1pvzajgVraE8Y
grw9Fj3EqXgIZQ9RTIVxj6x0EyKhnKdBLfomWJ5Yg8Vx7vnpIhTLDPzEd8vRWe0c
i5kgvv3GdEdnEGtKayFHEqILb0HXeeF/Et2bKKkhKu7qlPdRrUpvX3fmXA63H0XK
ikrTVJtueQqf8luIi9gffFnQKRCcuYatTEUkJ/oZ077uOkT19nBndFJzW5ot8Uzm
rhcY9A72NN3m+JrG+wcARkMPc4MkLaAs7niCDThy3ENbKKQJp2Yb4uwsP0dnTun2
u2AsEQmoT9Bx95HcRSpAuWdmvP4Rs0VTwjtKGYbXH1IFgrDorPoGbBZD3vAfXOdk
l2d7x7s48mqxdtJZzn7tKEhYTYNG5kSq2ikxTl2gczSyqw9AEfJGrBicp5wnWBaF
HkpICpPen8CrMHw7hS2wdAIMC6MkXmuyafZPhlBmQx9xVpN5T3DdZNV80sPvh0VM
2tt9G8oO+qoMEReSb4vC+ZjRTACnAo3/xFRG7Wev036jC4PgSQycQS6D/5qp8lcL
kHr19x9eINy1ow/5aBeacynfZG4BZMjsy71F557OnlruqZmlcvHXqlBCLEYJVH9I
GuOWnbFiLUVHrsg+mQJN6jLcBdJvzqaGckOhRXNDmWUQx1Elw+j2YfEkjmpTIVqF
Ja2KxWJwVtPabHtOk+co9szonplCIYgVBkqEMxHuvHf3QpomhqCGq8a/JPRDTu57
3VRupf9/WmT2+i4Bmnl9B/sct+iCQWsyhYm+4GcO3o2nGascHJ3CVdWjjoWviGKE
5ix8D0SZq0AISyfbIJzWQznNN/rRd6QXvhq70goq41H+s8HifsxYeMMUJGZvtWQl
cdm47ZxMGdQ6GUMso2LjyOv9g+8PueUEljBKtSMbWt7bKIsyuKmuLQUQNR5oj645
qoNX4hw25vStsuzuE0Lj7DEWHLPlbUljuKsvqTSo1jDXBa/Em+SVBAbVlgfHO+fU
FsnILX781puIkCjU7+25mPBQ6v8p9omr+6JCZbeCdmAJdRkD2YmL8BL17WreYcjY
9fW0uC5VxeRo5FRhWdLSK47Z64LvzxZdJBYJvf9X52eJ/v7/mpmWPJKxPBCkT9fR
/fYRCt8tgVw3sysJYETEh9FsUlPWsCdLLwd5ahTQ2QSAHudItbgPHX8J+JUfvri3
uEaHfeaXycCW19lxCr+SNnLUkiz96yPyU/iaZFKh0P4vTvpPVq7Rg4S9hBtq0B9O
wGGwgoKjn2sm2vo73Ui5Vxf3PTgCek7zMrCySOJCRNewxT1rxyEqeHznb44oE86J
eyzu1UFAEPSkaE/5avPoi6SNN4fdxY4CHzrscvZFU60jHrQahqn/Pffy5MRccBN9
Sbso5IXGF7CZRYc0BWykxHW0pU7EAM1S6vEl0rOezoJeiIM1uyOVQZJAsnrryLNJ
0HNm47dKpuU4+TPhvjxQso/BS/oLWWU+rUQ6pyIpU05ZBYPs6IjFnLUi2Gmbi1CX
L9uVPbPHdSXEwbBJVstJTapZkD1OCUlZImn8Oke0zeDZcoBZCv26eQib9KAWi3un
z4LFIQDV7iSzOLOED2ooh0f8/4Q9TUGWvTRtlz6im2scgg+MHfFRTpeCB4yO5t+2
DtdEVIbx6mEF5kF7dMBxzxCN4LPOf79w4wICC/oCC3kEQEtlPVEz3mRX6CUHysXy
hYuht7oIK4D0bbmG7lOBUvc7xiX28h+FQnluBhSEsDXtgDQnta1HL8VT7BKafdzA
mTetD4O2dN5NudPRKG7XNHY2C6NGtt9Tha5imYcWS01JLFPEYc1nbJFiMXcDMHtL
w2fQ5XrS7lyprdAC/vWVDaoumygN0qnmh2Nb/RYS2EPSkokMj4MPxqAgyC7hMJ2k
e+CHs/lrC1QFNfX2NYzBHVJgjRVcGUSVe3aafpeFi/eHJUDzpuw2lcLsrfsy9ZCk
k5ZyjsxMvk2cQI1h6DsMnUazSaZ+/wv3TeUafoMdGX9vOtJ2oCgl9PoqlL7y0sQN
4l4FgWnJoX3JC5v8FgsIFHHVNYDvppax9pvOqUk1FQX+62kApwzTwkHeREMeyqQI
dwlPz5XF6Qp3OZc0b605IntMG+v3qX276x6SYgVx8h1wIx6p43FppmoaucsG3xsl
azTRGD592Q91VWQ4O9rDDpRs7ycdc4q1g0aQwEcP9kkiJYZbxQcq8dz+ZQH/bUg9
Zc1gabeDcxmtrO9kMqNKzpaj3YcLzW4HBf1dM5jVa0BZVovWinLtcGr2eV5H2XKN
wORsUfnKwlgjO0gK5j+HpBQhdV5ULiTFT9ZLW0wvEQJefqRhRNKmpGBAlqIu9F/7
rWXxrFz2SPhnKkzVNiDmo7LL17SM57MMM6q1NTh8TjSrlmDMZ/4ceRNSmVnM6aT1
wfNHcsvhw8kcwMK/YfhuMpBlvtdegE6rXc4keK9rwr8xBCBTNzXylGNj5rpWsxer
cqyV1Xbi70+EAW/GHDNoCE1F/xOjgByvJri0f/FmbVnx4SCK4tgmfsayYwMQbB/h
GUhzLStFsYwUri0K+wz3Fs7G5qKbfRCCsXANJBKRxMOxyx9DFqKSacobL4OKLV4l
Jwqx13qMXQOZytO0Nnrzq785EW5XUKHbfRMTy2Q/LN4SEW/5X7+JTIpYH/h/JKHL
rWsYEoMkPDotDf5dmP8B357n74WQ4UejFlRthxR98WJtozdUeO9YRhPANedkKFuO
oBt/cT+JyrIEwJ5WT+DtzgW43XZIPpWGELzJHN4O+sIcisTBxEOxa+IiYrewT7Gs
GRKna7YXkfp01hynu6S5H3kB0lO6KakR2u8IxmIYni/Id5Y/7D0gJmnUeAMSapsY
jADmEjf58T/JOoy6XCVuyssxx6BhUrFsrfk40wxYMvEKg7vSq+KWL9R0674A7TSY
rQUO6tugTfPZfInXc0xCbMeB+ucK/EzkKR8Y4cZVU+abwZDZHcbSAC1jss1ViwUr
ucevxqxRGcWVIrvxC1aJ0YUyyTNNlxjtrCUJGxksjap2W1U27MoyjgNwH7tEAH6N
TlBHwjS+9vKcc+hCOxMp13y4uyScszOjRs6wZvtFDfuvmu+SIOfoLciw2FvJJBHb
SBbMzWqaQOvWk8+jwjeIMZXPckWkmeT4JQfFKnjkmM8sE/d021oZ4Nxd18ioMFwA
lsHYwULdtkqXxr8Yqecl+GYotYwPgTr/GsNtK9IMQD2Nis2z/elpth5dEd/PXpuz
PaHHTOSX52LuuVKDhcYHwJqrYt6SclnV7nUscMl1jP14FH/fZ7nw6ul1dCVA8wVv
73sm/elYhTvBXecAicMkJKuNvWEEE9isXZpVqwBqgbpNLWbFdYod6Rvf32iPJksF
Q42QgybYOvkwSxmbsk2mFDWgTorILH3/quSJLUV6baUCWZV+avnoAnVuJef0fX1u
zo/btPLFQWM4Zzg8dB/+DoXIXlE69Fj7Qy90b7I6iYhaoUpGzWVbQnj98BHew4sb
Ykerb9/Sr4c1TqRZ5te11ic9yZfQQ54eVqV5KPBG0hkXWS4jboOXhp6Yw7TjOjwJ
ofOHcAuc9ltkRkD1l0IqyMdBVh6tc0G0Po0hjZ/abP6MtW2RM86AjiaQ0ms4tFjO
bzjZLbZXM5Q29pnGIZ0KEUIVIcqBIItpq9GzHto5RzLOR1OxRAWxndcgqKx2wASp
SWQh8ddfsClUmgRycTZh+uJg5L2jI1y9kZ/qZjomWUCq6pqZMUfrovXNRkEpQrmr
xuKZ0NnwH9Kqx6MjQR46hlX3OaYSsEfKP04LmQ4fZ2mDKKrpEsH7r609uKEiycr3
KwTipO+wSKx2woGLncx4wsab2BeuTz4iIxnwx10cRpP8Larvz7HNIdpxWGz9s6Ue
NsWQhNYqbQL1qcXA2If+m4RHiHem+tIYVB74gDMx1uVi+PkjRPonh1Yk0u/3lHNN
eIqMchTgL5kkCMNtlvQ+pzQ+VQ6d3D63ct/HYqBdNcgktmvoyChumLuuY3BQx1Rf
KvBP50+c9G0LeBHLetNMYxfKqpaig6XqGdYQ/n2aYwFUCO0MHhQ/fpYPFIut27uC
pudAyIAJFVx0bjPMsOZBGa3TKQR4dMwUWmAGAteG0Bf46IKfXrbQb74xv8kESHTS
EXLLM/IGRW94yZNOoB4GqQ5/s3mHiaLgGC2BreWw7a8GNTxi+6c2buBgGOZZq3OP
sWNyWNq6Nz80Zas/AdOaLm74dPy4+VySdAGA+druaPrY9M/1xzerNCryDQxk7C0A
8Y0Pz9aEvv3hv+yGvotd/Dz4gPKSir3f6EiLrSZNFE5eDEJW5nJxpQY26wPkef8i
J9MJOZnRsqErA6h0hhjraXkyC4QPVD7mmj3MxZa6STQcm/x9FO3GQmAJD+1sB2bY
7K2solZ+9WFNn67a1lBM1290MaMb02IGLaOfMvqR2IAwIpwQ3gAeJGGE2brB98sK
kiXxj2tHO9V0vEhjmIksbr8StAckxE1h3q1Uzx6sdbDc2GVciIW65WZrttTfjFHg
OrLNsvzgxUVxwpHaxYQE/rBNGRURVtIqqo/L/AMqVPjnMWIqeX3jEL9tNDvwGlvT
foS4nfy59JuaugKti90MAEz7QE56cYhj4Zpa0/q4vb3dGkRRjDy06UPjnSpm+Bm4
JnMsaFsiEIbfJClyqYF8zydkd9vRoeZ86xZVf3C7lcx1d6Dhxlj2n+Jm6LyZJ/+k
pwKLZo4LGYxdf5d6AmUD2wfXF60d2aZRuJM48O894ioHyB4ThcG937G3bGsTGYEX
oJsy8s8X98bddwRt/260pe9IOLxOJJTEwB8UalqUQYOrSzgaculBrvyCppumQz3W
iN5PAjzdknLs0SNgr9OBAq6kh9crlBLJ+GoDeuYaLJS9lnL/NFj50DXytwWo4oEe
QywDA8IFEOFYRX2Sp0rKIJG1b7JNIVIYXRSXTK/z2z1E5exgUAhQ3wim4XJ4jniQ
IrQela7Qu8KQJVTzyNnp+4JQmD8BJCmDkYIaBp4h8B13IxrbO6SBqdYDcd7dZFye
HhsS71lrZehHg2BsFvhPI27PgwnX0iSnJ+ntscILmo+mA3D7UAznzWtT+aeEQx4n
shM0DSLwFoCU2RvrHStlNiBPRjctXmPfT2hda7bytn4v5Y5N13nr7x+O5rHkquyC
dsmzkiWg1ZRrdQAenrJQzs5f6xkTrVByWfGtoss6t85RZMBSO0tc61NSrFzoocJQ
dtULe6dhv8mUJPb6SFs+QV4VY3W+H5LQU29SwBNA/3hhhbCbFL3d+9X360D5yhA8
jVjCFIuq58ObBN6Rvjub1cl5ehR9lTBK2EiirBTUvpMVhga4WPffZfbbyx54o2vG
g/AANQkU+LJjZWkAAyA0jAu6Q8RpqU16owZzkqD8NmQeE+UPpDA39H+LKpPVvULH
BsRa65x0kQhOTm0h8Dg+GI9ZuYF7epjVn2V4e+kJxv+SbvBf0EXjnxaAj3he+S/f
dmA8FBTL8/7kFj5pU0o2+r5qYJczrWi8mI+K1NYEv6kXzoxiqwPacf7IYFRNQUW1
35/69lpTJQwYErd+/in7GRUBOFiHBPXs4BOgmVSmb8aHJPOSgPweSkvyUj8geDIb
Af1kQkK3q0AakOe/7wi2StiCCog0GnLu0ht+qtOUW6VX69luPgQ0LJUfdHs9wI21
us/p2rxq2ubIqr1SLpltW1fcmrRP2IIYwrrCZuBb9jc+nDzJLhB30Yv7DbeBplW5
VHL3GyqCNSkxlJt+TJQGtW5Bxi6dbdILIGZ/ITwQ6fa4/81v2+rSEQPkcSQD1Kjc
8mYNHLRM0nFWlh9G7t/eOtqPXDSUFpUi6I20FZAKkiuJloF4dXviksQOVtzExCua
eo6Is+qodu9Lt1B2His/b8KtY6fS/+05SxELJwGOiOf1bmjwKCOB8o9v1a+MbhK3
oLTlPBcBhLK4TRV74Xsw9EBR60OSIz2uqcQZQBrlEqm6aux31D9dLGrGPnMRZGez
IpZ1586pJNbsNwQuExhMJ2zIfNzZfXHomgc2hpaiW0X/msNQS3rgNiI7Yse4J8Gr
WOUbrGOPlOyqHVpIX5rNAkKhdao2//wtom0dLL6ltCZYQbOVYsIlmFYyAyfznSps
bm6uxO3NLwprbaFZ9uNKX7fMvJ0yAD8IroKLZMMagDM9O+c5Xpq/UGT36ZcrNvnd
Djjq8xgZBWy2FeJrpd2W0aB4XbBX18jHJS6DmCLsFzpc+Va53fW/GJ5HTr61zaw8
5yIyEnfFeMV5DBouHaxLZDksaI/O8Djbipk5pWZ173mjRRR1yQnbOsI25rqEjG91
af24AOyYQAsO/ZVtQCbNBomWZO2i+QLL6U8QiikRPpOLTUn1IvZw7tWxmBIuUgMo
Do1cIB/62PIXFEniiDKsm4ObQdG3ppHkdNPytzPyE+EHPvG80pF1FbzPHNzc/dZC
OgqtE4erCTa3VVdFJusqwWxadBV9ixDBACOQLjj/aa435kLNqFYhw+1OsaI2glwl
NkbCwU6xQUG1DaF5rn0riqJAmtVcxKvwn4A00lbbfVG4UX1RrDm9iUz8iaWMXSi+
cqy2DjFKHsfwwGEeXZopXTlJfRqoTfYb90kBL7/SzeLAScbKuhNStlZ1wNmGJA3v
i3y8NAIb19Qdxdc60STUCUT1kynOzxQ9Fz53wsiskLF4JRHhzpHikNePSN3LEMVj
lvHG2ZvofFes/VYNwpAkoWoaCpr3EqX1XOAcC/oDw8hPQRsVzJkYSXBaKdfMwbt1
uGB+mbfDcRA5JNfROLZTtni6g08FV0l+R0/S54wzcAlPiELSto+mEd4vViAskIpa
LY+lnYj4wYXbZrTYSWPPDCcw95obCr01k5EOqa+no/79H7SfiGEH3rUBQ0tYbM21
n3TEPx62+J3Ja+zBHY2WxUS5AaJeD+eOGLKSlr8hRKtMUsCC9T3blb9M+okj70fw
PfjLmIiBs3bIgjIBcgyrJiIN2JhCweNyFpp0E1X4KsRFQ6pfbFhPmI2BHzMPIY9r
RreCU90WiKmISNzzFjSMCdkxj7wM0YmTQcSg1DdpqXnKm8mbAU/XF0bb0AOkZl+j
yU1LPVVMptQsepUK+5pTyeWNbPBJIraEFw1PVYjzSuLeCgC3dfvnsWPpuqkj7ruN
2dCDhFkPkq+nlXz4rvcYXazjx3FDkHWAHfX346WmlVylOwn1fTHhQ/eve64JfIpB
Ncir/7r+L+kFICxmOgf2AiBeTHY6KheHol2Pc8SYka6fChTlhjCGVver+WlxbaQB
/gnLx4tFDckttTWoU3dtAdIVpTwcPddjGGbXQNuY6avEAaC78LFdeJi29V9oOvPs
9y86J1BXHfTDNCAPYV9e7/jlH3ZU1A5RgmJdDlYGDjYNBwClqJGsXGmStiGOItYI
Jgafx7WJuyGzgH5aHlOfDHaq29edv9yy2au6//rIZzc74PkoNW1F9K+PVr0Tu7MF
rO8AhaBj6W4qwd+NEDvLIvRPUHaNz0TmxRl3W3Q3IGCFPZmFLvclsZeawE/V2RlL
Z3udpZDDdx8UMEdHDoRDm6QN9IrRNhQ/HwY5m9kP1DCKzpTxCbdctc4/XvQpb87X
/lLWk4+A/m+tEeofhCiqfh6bo8Evas0sSv0iXE8SxJM1/eXBn7HWbGNmsRqggYHf
BP0WO7OKVYqXu0C4oH8orGVq3YGm8AnXwq2FEj2mdPiiThfO0jExviTArMQ57wF5
pOZcD5wJtsi9kkFXjTmTsXlJBvGGjSFS/nS9oQ39vVH3OnyOA8vzNnh4IoacKmey
zEdKpbIJ1ym6P9ulO4IyuD3owMeYpTEPK2rwgmmFkvlS0Ei7SNonatVwLHTCQhl0
cqbpgMSef8qVFKr2m2V5AguEmG3YaTp/Q+dpIAUUWYuMmIqIONNfnE6hSpReBdsA
2ikOxI8QgZ9tEZE0z57p6kDQRbuFHOXj7IDg/7JTQnlw9bCpoZ3kFNukFxAHapEy
e7p7idkua17L54RJO2C9SSq4fwdddZoo8l5n8fsh9BpYBMdCeBjoRXY7a3P6nvzv
cYXtLn9gxMxzCszPxlgKgZEB0jT+PS8I2pZEa+iczt3WLtWOEI2BlSC2Jfbrz4J7
otqRQpOAYk9whakV+s9rN802slJEwFnjynEytcJ+HPGfYNXxfwk7B29Oe1ymUfdJ
hiHVmfCjejjDKT8hjg/n78vNkNdED9r+zv/8zkkO/f9OzW88JGoB7rRu87lEq0Rn
BhVvYCqz+XHTre6YYXZLZOevt4J3Kxttz6nJpCsfJBjqo1qgGtavt24WyLcixacb
kDA7+Epj/QD2OqvTzPjs3HeHXRzs+SiD6JHKL5hAQ4jPH3Z65/wOU9+8JUn3pVY6
/QXLhc0hU8VUdslV0zj0Z+DRcKp5RKZKSxAhOgNmrvQvk3ZDhnPsL9B91rHYg/r8
UNWtRQgSIRtmzuGeCqaLEGWFO+XX5SK3jzirmewQeZ8PosRMpQi8lZNOjAP8wOES
f7eVvKNFK+5ahoatUjdM9INhaQFm6dg5JfXcLHgx8mBGxCKlELS/xA7Jxjndql+i
Ab87XFBBV7plQJvnFe19MlpTWf6qgjgUQQy5J1VSOmUzk5HArWzzfE32r/Trokti
6hfxn/+roPpoLRVQRhLF99bqb4GxJzwsuxyDLkCeIcwG2s5CQKq6vzOoYo6tPosH
I02Zz7MdKTmEcaXdMEG91F1ajPJV/9Wi6Zf0XvAta/gAeUcAWGmvfnI4sWuqXi2j
mFWQQNLylEAI0H8bArgGuR1BOMdQU/Rsdibf5ryj7M1/rqMo9PFUnPcDdrY1RWex
ntKOo3NPy97ZUeMeKsnsEZyxjb2zhmLs9ntmmMagg4w0ekdESa60d0LekAnrIWfn
T4QFC6fXPabdztoAU7lvkZysLbSixGNOYbHTdC8vVRRJytn0iFznPYe8kWlcrFaS
EkqQovPInS3FnVDVsncqtkhghzqAlHnuQuOznPtsb56BXjAveWJpPgN+tKkl1UKf
pUBFtwPLRFqdVfqvOXN5LCkHAxliHT++PGR1zbw4dR5629JyBebxt5hiDfySOeVH
YA41o+wT1jWquor0DdrbV1k2B9MbLt0nuF+c77SIYu+k/WUI6SmvyI8vxvhmaVRT
1GgZnS4cXeuBVeusZdK2VsSWS65kAw1pq9Y4k6q92mBCZVX7c32QFwJZd+xTBPQL
RpQ8hx3IajQlg9jnNLaDPxFo8NmC+SnNcMG1dxtQXFq58Wv5zT6aKjnrgk9SGR3v
HEPz3zXJYJRI0iem9ItIS8a4pfEvr3b4ldvM7jXGjeBrBZDtSo8ztvDG1NCtXC5k
cq/gh+STh7X+iVTY7QpKxNWLn+3+98jVZP4h4KIZfE6mOZCjDMPNi+qdEJc5vMfL
yIVk1LGncCXjK32KEIOP4Ze1jB7aYFGtZ/Tf5aFJqAdUG4FOxzeuU62k+yXDLD05
Fco2r3RdsioD4f5IaHgsWhWrc5tLuh7+sgyzopfNWDnLWO6r0DEDA8EjN5ADY3hH
wBE4KfKX57GCT1FP2rn60XaBBXu38IZtapPBheiBb8kLDxvTAJo74avj2hpkPdCs
kdDqKWim1QCP4MAJkIHOp6+2uBTeKPkQC+Rh+VNA4b5JY5KipoZVAftoMvtX0XrB
PpnSOAjGDy7WPcSl4+BiejtL30kYc6gxhIFwjraGfgcCqn+iZBRJ8+ge4if2xV6M
HCMb487S5egD9mMRWHYry2DM4mPcr0X1bHyW3G8iCJEEgn5Q7TWncpTYV1hk98AH
YLY6cHX1ahVWKzpy33E2d6Chx+xLQxshpHVqUL77YIwQt+oOlfhIvOtDCZ1hFnHi
M/A4gB0Q1sflw7I7r6+B8JmdZSZ7DkUVKvzCOcOm6YDcpC11wnLFhT5S/dDjwuSm
asnHvTZaav7zLz1MOcQsbSXA1CyWaJFdxCVpVYxEoKPS4U3fkr+UF1ErcCuGxmQJ
aVGSn6d6TlOa9s8MvCgxmtBOVS/5feDtl7TL7RqwOkmSgJyV1EesjVIJkX60s/ds
u0SUQtkLsYIccukE3qYFGrpHqvvJsHHwEkks6V1h0byEzBjNVbxwn3WEXiE3IG0I
D4diyELzXhjg+blF8PoYEhTMlbZEysFr0jFSgJoUJW7DPEDNtZED/0TbmMF3W+IO
nqCZR2COsLR/oM0YdmaXhPPym/lWOmfdx8FTkHg5WcLq1dxyMBmKTixcaY27kCcj
FxjvfvZ7T4gcH2ojuTbVkN7NyXRiwGLdNz1j/e7bugTn9YHqO9IHh1v34xMkZ7fP
FkcKBBRldtw85DxWl67yJlHZ6gda9ikIjTB7dRouFgq9WOwdDMODb4pbxtAVgf/c
235TbakxG1Br3qylsid99SzKQELmrr9hgWlpnmoSsfUvzfSqlWMMV3QbknvAUFFm
Zx7N/HLUjgKgrdEKqjjsI4x47J89IGU8648CfhM21Eh7CYklSLD2GiXN/+O4kGk2
5a0EttISaHel2K0TfG5jbE1AZqrsASYADC43iDGpjN1NKmixbU8H+UpQpKEUlnxK
8K4NGjZVllwtHbfAtOZ1IRl6CEYWOcP2EVv7icaGS3WmWBR1yWWmbRuyKR3NTCee
uAC4bCNccy2CZnU4M5KV11d98RGXP/MH1af72duHD5zVW7TCSSiHnwqvS6RVuh9K
eTCssu4GVshSssK3nLovjgmGhqitlfXQ2Oyh9cKprYdTF/LTgVnBcP2oTjhd5WBX
F13sR0sZvsRfvaSZ1tX+HJXASokIrabwGrKg9heS5cZhxO+3tb2qqKjsLH3uTgqR
uIqtvIXWE3upPoF+a/obPnRIwwxZOCIMirnik69Oh4rBRorGa6xsPwcFFPk/rG6P
YXbmFw/usfWqQVUS+Qj+N834T0B2oWRpo6T51BSA70HWQXisK/pmNAg11EuPCYcO
xN0UAIaL2XRIJYLIz9FqsIfaCItK9gZC7k2ooj++lXc2wPvLyCvj6xp+9EsznjuR
WpmLUnAW0KrEDUV1IiL0trSd5oxSIMgOgUeTZ4MBXrd8JiJX8fJqFdYymAIgueqw
rtBZ7xukF2BBvAqodowYbSf8jtkjsc5fK1b4RcUCbyOnOi8G81XhM+c8AvwBDB4n
u2ptBh4CH1dFMYnmQZJdoNYoLF+kMwUDRNyoicZuX0VcwvIJ42HHzm+TteapUYv0
+mFiWS0aptsyjK5X9YtF1nWqhskUPLyZ0Z0CMVewZbMAeX8VUiWPhawf5djCZqsh
zaBPWIoqjCkT8YicNPBLxPj6NxLaClLxnJHjxpgcHzt6L9g5Pc7cc1pMGMeMccOR
RloDDEH0Hon/XfuKf5xtYSoSU9Q/Q3OPihiV9PqIFqoJaorbTAuFhf/WtlPN8gpn
EM4ne0ZjkVeYs4MNbGKuzwRAaPv+Cx30sFstyjN6C3qrUVcXX3fDkB3GwgmDo3sT
ICj9twk4mzqwXcQptPs4Xyn5MvpW0vkuVvEORT+nyZSOrlQcMzTaJwADvV8bdbSD
W2tWh0AFxA0wFnUZaihvEg2/74M4eyz5qSm7ax9MkjRFnbS4sxMwvvpuM6YeeMlz
KrbENsfESjzscih0aZRU17cD+/N5vYIV/6YjOKWV+/92/fPyGkcH3GGBEpHrYqRk
md419jMaZl4tj1WuHPeZud/cUROqhsKKqlbVPdczGbsOwOXRapvaLOT1ijIkN83R
DTz0pvYPgTiYoXyXL32xgWc33Oh79lJDT4IrAj7sZy52z1HUbX07P5NPhV2WB0ik
lj8nItsXGHSMLZ490cc3f2yph+ZYTCX4eyA8yWEpxQXLf9RKKlzfzfc+UyuzUbZM
aJULH7W8Wv84Q9gXM+k7vrLSGCi8JC0oNaNtHqql4HCym7mpYtw6Lw2cWaSTH3PN
Mv7xoxL7h/EPZp6ME5xIHO/t7+zJoqU5SBHeSJe2AlXpD8ZQYSHPc1eIMBvrZOp+
XHCetw281plky9dryNGr4KcrIc+4Me5171yuPgocol8A/piRua2T9pFoDXveAW8N
Wk7eCVS/5OB8KzcJ4faj6aZ9DlJMaeeS5/ZO5yV8i8frtEcQRZ1FSvVNr9FXFJ0v
uB+nGJ+2xcunuSld/wT+A6WlDr9wew+B4i1JvuJe+HDmnOATN3PZ9P13XiehI9oN
gW+JUqdX6Oi7IRSSAUMjv+U6uF8/XrncndNWB60ujk/TXNTludH5oeuWd6vzJc2z
N2NzYyZqDwaupTLceQb9y6IW4c5x+mfXskopabYN+CB5326yzS3sbuVUPN8ye/fS
W7moKF1bV13g5S9xlI4EnAOZCy0hrSao6m8lYrFwwgxDAvEjrGNuTim9eSAhKNS8
Z+muD1ZrWmalUaEpVQASNJZKJIpXMAMxTozIZUSQGwu+/2amSQUkHUa9uZJf8AL9
FtrC+RWaLh+IlL1C9XGg14LZd4/ZF3P90w6rbSpHRAWMf51ccVdWsUKJNEG9/qhI
cux9JixSgZNJuUsMRjeCxy6OH191UUzMlaPfR8HpYYseMy98+R/rEv824rqtbuQb
814Cede9yChWE0iUmbp5Z5H6ZV5Tk1FgYof1y5ex8ivvnZW76LLhDXR4+Y2JSnSP
KsOJ1WaNArSqBxOlFdhzjhzpRE7RAoVsh1l1yXVkE1d/6f7WVzv2/zo/y8Cb/Wqq
VSTXbiggkBzLwC5Duugxo7P7KKXmoTJZX5FINYSiIqlfnXrs2xsDezAyR5MCKCVU
bKIQbt1ddgTZb3Cwv0k7fKXbzU7aWyO1Ony4KvIGFcp7OwVa6fmCW03dq2OZe5/1
jGRZgDhEG9kxpNLrInUjM+RvJS7f1hgy0SZHQWHLes4WP8LbxHjzsMMXJbGvZvew
k9TaEBZ9MbglbYshmCnguznWkaif1HO8pI5RZzvdOPLu7OsZtGU2D2xBmy2hlVAj
JgSUOZOyOdP0wZSGyYmTOZ9laEfB5t4r1wLvMIcfcP61YmVInyAZASU1CKEwnffN
rTHhTKvlLe1aAEs/tT7ZWwwNE7HAc7HPGVTVsW0EdCjsAmg+Yc+0na7xdjrgkJ3U
BBX84J6e3YA3+pTwcoVeCBzg1P/joub8qH0uk5ZxCbAA1anlJwgPbckjulMb0O9c
YGA0RqvZsCoOtWhi4N+hvHmGQzkutLpU2jjrgX0cL3m8oB4XU6INfDaYm9lEWujM
2m1fALsxjpxgvYouikvhefR4lkAul7o8HGHk5hVPQ7BubMlhgmdcKMACmZmk9YaH
qiOBkyy7ZczrNtZ9xRLNlMJ2fnsw6eJWEN9aD4RrkxMyM/R82h1Avc6bTM5SbxfC
+zkH/9YGJKV8Y+8JHaaW25HoZlW/e+ZPZU1sqcoVS4gIrXZf2BMm3tAkRoKhgokk
FaPv7w5hEpTfUQMsk0tFNpragqzYeLpF69lCRweDuZRc5poBziNByuoSVWlKr2JN
MuHu4zq07RK5gP/8VhjzOe/wzBigTF9/NL5WyA/xtytmoDhwfQgWbe2Q6Yz6JQv1
5knNi45UrE+y0tU6xFdj5h6Dkkr8WMR6j0vUZvDzhrekHAeJY1Y4ogIcHC41RbU3
C8K0bI60z37ZFOzrrjrnOFV058RvGu2qNuUiGiIdS8Uxb9tmOx7gr84D9XKU19BU
tYf48UYOVEXvhWlP0lEuyUxcyzI03E1+IRl9q70G5wa4tYgXBr0Uqch+QAxYbWtK
zmPCaKrOrTL6MZpkjHeOj3X3mB3C9dvFR2d7URDpgyjhXeqg/2rPOMj79szSlTKf
3dN28MXQFyvEzcpvQDMbl16bcnf3BZRMQzk2tH3DVIYwUqh6EtaTSchXpNoC+WFX
vYcUOzDjdnXXrys+hD1azniIn7UIGL78qEDQPkj62lYYz6S2WnPCSPWmmZnDst94
tGdmb8xLngiFR+xb87wZjb1OnvhomS05ZklRHIaCPkkKVkS7sxzVOVKXpLEAPu5h
vKIl0kP0AjzctPWzTdo7R19R321x2xdiwGDPv82NSlkbccLF/Xaypkdstvg+z3de
1ITdcx4DRjaU6qw9Ew8eE90pEnaHYHZYQ5qBSCbFSrzDkLBrCAhcWPVoYmm0IOfN
21+LDlYdj4+kGyI54wR5NTmf6gkHXi9BnQVLIvesyHF7aowDic52M5x+g95oKg3U
9jANmkCvoGu9t78VS3Uuy7/vAi78B4hpFAVM7zXdFco3SYZLOESoyOaYGSnoR/0e
HLM+hRGNnq6OwGA6GOesINp+Lsr8hIrvLoBUsU7+coYb881ZlWmN4xUP61trK3DM
zT1S31OOVyV/9yXA3t1LO5lAGrXHWuso/Ykm84DpnhSGEtFluFickii4QzuSP+Pc
BpJ3ROmmH8vJ1Miy1n1j0EWB/8e9t7hJXBzvezqik2I/MKhfZaG20BfQXTUdS9JU
ViYputW477edmuGuV4Sd25soKEnFNK6L6qUgdgmg1fYdYfQhii6NiHNwc7hORRT2
EHxgB9YNJSE3TiwQq6cyIY8oHt0dFNlqcl8hKSq7EIGHPFlQSox2Zbjy4xmzeOGi
pZ8HSpgO8+P3Oy7i8tmKf54qrgNQfxXhj1CV1x7kgwY3gaov36XY8xX6+vuco7cT
PMvNVVLIF9TMm8hDwAsvkPCjHOOr2jXrgOuQOoqeMtadtlOWxMVtB2q3Y1CQkxW3
0REZtWzIlNZe0Kd/xqLyz7H2blfhxSKayItT69pLDZBFP3zjN7+4jkBOHaoJ0xcy
KbRxcaDbTCzJvf8VKuRoT9qrc6WCqme4joMxzFjEftI3hm7awkf55BC2HsFAYVxv
vIR5WEH/l2RjiKQflVtXeIyEJxDyq2qkWx+yc/HhMqu4DJRwJNsyapzbkrXS+RkZ
G+W35X4NK+ZW/Kaqy7T5foSbcnCeKfKrmCiCHJw2UgLBOf+XJt3TJVhgB/SFhiUm
Qq4G6+hnrVW4s6wJrDqndNaAjqyAdS/Ypf9N18oIFMz/8ufl2blvg8zCmqyQIb0L
TDW1tdA4xSXd5Xcl0e3n3ziJ0heUvotd+6V0GCkPdk/DXDSB7ozRjle0sEC9Jrxv
9XMYV08/G+izirLCofFlj67P3F7j8FOBMxXECPYT9TOoIXi4IgIemZiHjPBBpzKR
b9336DlE+ZrU7+PEjHDNoSkbUz7Op9F2hVCdeHnfr8ofjDXmX4UKxeMh+XczMWRp
MOwJaS+Ed9MqRItTJEqLfl2PLX3JlllBWvr/9WKvZAjOWqdxcji+x452mSerjR/5
1pGjAYlu8Pfd7gIa8gml5rfIus8k86IvVuklvPD+wUqO77NQoh6LLJgCo6y7/c/P
2bFzUYY5trwVZzvEx4kQKIcHOM8QYku5pM0b7fqFwBgNYBBATSdiztGNJ50Aemka
rWTyk+xGJoyxXutJZ2CW4nYkf8JfaKClXOtZTnzSJqiWrvalIC77QEiAW4BpBSKs
QRbaeCI+dWM1xX1LObtKsHOiNXPAVijefjcUp2PxBFDzItp5BIZRvkegtpPXfUvT
tGFsUsdE5r6A1j/2SXoTfW7dfLoyywPWq95nVRynPqkz7hyaNk/Q+hoONWOz980A
ulhImumPX8oM+WvCXd9exzC4aU2FJjPC84owHZvL65wiFSfWlxc9ruZ7WRGBjZkU
bVebZ4t/VgEDX61viohVkD3r7e9jO8IRhkyb66ObSOPWXBaLJ/3LHQXEedh/UNLl
oBihKbC6aO2ygdktWSWCGjg1/z+PL8ozHauOBRgiUGeS3jY2uptDOFIUHxxKzEEI
/9lk4WUvFL34S5WQMqBaZwIMDPaedcqb0uIhby83cPpeJxEwGhfwFSNw3KhwDtyy
NjQTl+wjVru8A2v6p83tmkV7D0IankYIban94pAaU7Bb5Cqs0Cf0/HSfuSlIPOGQ
pBG+n6eQeVck5zAn6LcZkJnRYXhqU+hrZSD9ifMOmhPHhi5+GBhQUueoVaeIdQSH
7ss9GlXkVnEx+m1GGoRdbc/Y8srW3+W9vYzj9GIfKXYG5a+wwOHPjIWsXSFbFa5c
A3CZm0z9thfw7jF1OqCZdbbq3owpCv4WiKhU0bO3y4dY11/SMQS3MPRTW8uNKxKj
mzsOsTuCvrBZyRPdWriMBIW+L2WBMVNEufVnA5wl3IlNDHxk+8ZyO4R7X3TiBZW5
r/5/WBBzsaHf9swqihV4S6prLrSKvCwQJNEQnzBi5WBPFFOWIXiDBEVOvgpz36fC
X6RP9SC9FinOF+9lr1HL4TAmYn7X83+5LqymJSbmmQXRi9ld5GozQHjFyi4Bm90S
TvDfPzsdXLZVNdkObqkVup/mnW0AWyb5EHADalulYPsjYUvaG5lpjcSK3QEnpnwc
k5HtVq1Y22HxaWylQO1Z3wn1bVnBQwD55gpldzj9PObiNRPcVCEF8Dza+BrMkRub
OjcxPLC09cZF25GNZQSpNPqQBdK4bbYIk9J7rskM7Kh7Z/c/HzaIhLAEbQcpZ1d9
MnAbg8vCOSx71kenZx6ffRwflBxmxM6QHudNKgrSfLMxUGS1DpFbpDtnr1PLgL0P
5GAr2RPqWwhsb1Cj3UWApNH3tAwtnMTPzNbYwt+qo/kf/fDTyD4++pyf7jrqISIq
+Vw7UFG0TR9PK2AyDIINM5kb1i7CGbcjrxDTfoyUr9SIq4jBSAqv0L3DKqTi948Y
UkvowXlWAhj74AFVmAp/6XC40TobuvJAYzrpKQhrIb71DrfRpzvjg38Lb7V0n9we
jG3OhxkKtQ881DEV2OdxSQM7v7UkDWBZkxP9gVM/JMGNl17CWLmu/jqpZy31ReoW
jYzy44D2YwkmmpWhRxNtNeLgoWkRFZQzj+ySaJ1sIwHosrpsJTQgYS22XD60pn1z
ypzpd+ecaNEyy2zJRmlottMgTM8GLdm45cjSu8KOUCCMlWpf1L7UmTb16po+gpcz
ohXT0Hr+gYFe/hWl0iZX4rV5r+ZflbPYDmzX+miCqruNQxi+ULYo40iTWoWCbpeC
3dHzP8DPXstPTZ5vM6BozXtKM1fcdI6tZ2kv5Kz4jmO66VmyecLd8QVBQCHay6uv
ISsURq6paXDL0pINbNE/yNFEjerTlgL0MCjiS0NCv9GkucFsi9cBLeba7p4C/4b6
tNCTlOEwhiSF91pxQnhAPDAiBVN3255pyUCq3CbIEMXkrqowSl1tdGOiMQ1CjU63
zECWovjIl1D3ciidJt4BuXpPo0fSmiSUpDyRCV7Dnqee8Rs/1F2N9p1TdG2oSSf3
9DfYlhpIB0JiGo/cKV5Fdb36u9Tjx+U36p1z4sLWRc+ShvXapka+m5CZbLqdHzaU
rQl744G29dRuaPw07gNQaHvWL28wNMgR7/ugNhXguTMSbARUZkagUbGnyg+9VetH
nefINseo3vAdhUDJ6yXhwBHs887UFABglV0onMBWpdN06HQ7Ci4varfs3MD9fubK
QJERxfD7Q5fxGfpCjbvjwMRDxZ+gSBRhMKwbXdmwUvQQApF5Ti86MrBKsyAJGcQo
1MYsTz+WcMEMA+SM25X0hzC+8OblR1s99CaoKtgDNVeKOJ5cTpIKvxipKUKx3/gd
FYH4f1BGnmAYtG7lxHJRLrjj++G9qexlNfggYbiiSl7oob7EUe0ohcrRz4Qb/A8p
bCV/fTSOeBL6F1+UNuzRJkXhi1wQxn6UwCnJBYwwxeSXUVG2hTN7/xJED6OM6vO/
kXxYmJCPLqjV3t+wTvAWMfBZOG5vR081Mznt7my2ryfgd6NdMEG2C/d+xMY00HUY
9TM4Cmu7CSRUPMYqnkpKUJEgvqoPgvmsRs+iXNLt9AMdK8wO97iycFy0DfIsP9a3
Kwg5g3t6gcpBpROKeBlHKbznkO0qINyFMADgnM8Hqe2cKaeo0at8KDbjVlwfTWjG
8k0eoEV6kHqm9t8hObLij2NT7VEMmobLPX8OvshXoZs7BfPSVVve5/ishdGm68jr
T/FyNPls8se4ME9+uZ3WnO7XG6QCt3yhIdmzkyiz0GsWXXjJc+Zb1JolLOo6T376
cCgRJak6Kbv/u6pB0uBKeh6wmxQjO0FHe3QsognybwPU0W2AO5/aYqKHLNcd0eqh
2F77WfDF+BHJZMxIrxhigXzQin2yw0clA10rl4S8O6A+nXhj9oafmMVUoTVOYZjE
F9O885jBWmspg4KbmOKzmR3V0+AuYYuaBegqWXXWDR8gWWC7UqKPBPPSxjw9tjKO
qgQGF9VbqNs3iiQQTZTU0LOSfGB+iw83Q2yCI97MWvC95zGYbiwS6f9kqN3XqUhT
UTSdc5E7NWZDH9UvIQJk6L0XNa4XofISEwOL7MfdM8D8YwaGlOkvXhx5IGY+SkO/
+bA2psVHb9bfd17YskwJzSdfhSmiKTomp+Jk9R4WkW26y9KklpMQC+V/WxJ98HzM
Hm3F2O52AFBG71iSflshvZRkuVZR3B35p/AKZDCaslZ0ikWkrF5TaNRfyZqLbOOj
i5SkpIZs2r3D1jvdCHZtrGHGxUal/Iw7XjYYHZu8mscvUzOqqc0OeYkTItb/bVYr
LWObggI7lCjRwQGq2xS1CPFNb8Oe5h9jn1Q6CBdNN0s59+6LFKIpD5q6WrzU6Cit
gz4IlEc/0xVG31TW2SHuldq4ugCelanYo/AxQ2TzHgBmnL1RZ8wmblP/4J7KwWNE
lkBT/UHmtn4VlGkrIM/3cC31thXFZUFCwaa509LHtUg+0VharY6jSlZTeXK+Fwz0
muYnF2D1XUfuJAryaIPPwcCNZrcIc12QHeCuF165b4ey9//vbMPTlr1oBfZiAjDQ
6nA6aiWyyytE3mWhvE8VA/ksJzok57X7KYv/EF3VH8bWl/4de6Jsrne40Q61aUoE
Xt6YS8613P1fDZOAj/CuZxgu5a1IMDB8bp5lb0+hEXjZ2CqCm7D9x5atWfUgG6Rb
KSwrEzYC+9WCVegSy/6wQxTeYXLFFxqByQ8Rq+mDe/kOzVSOv0rDHtgmcPR8mcoS
0qwdBnvuRr56ZTrhOMuGEyMBWPenSAsTBtpOrBW+Cg8VHmhos46LvPRgms6Pd6Ei
q7D0fD1J8pfZSvuOa4MoeBla01Nmhl4iYfJYnmZS8dCagLk2Rirw9WK3ytrMbkE5
Oll9cid97EuOsqUMKXJ9DXxTqacnPOqzfqxK4wYquQ+I5HQ40dXxNqIfi9AnvamJ
ShUvrbkTM+kmqYuTm3GLSA2D7ihQpfyVi//M38SxR2rVYHt9FCqZ9F0LrHySLuET
mp97jnJeux+dFCIS6O5zpD9VPThc5ObkNsh56uSEQr3DWozPwqPpnC0etlaX0iVq
SIHFcHkG0W5KINd5CJwLxzLnPmW88jiHunAE+5Adwg6RWDGT/wPNxiEEbb+pYDYK
WdaH1FgaTMk8zUZngWTPlcso/CwO1UHy+Y8fAAtXpeB/BMueyD9pGCKv/aEbh5FN
w3paHzJ1/Wnxg9B5KktgmNPUxLJVA5XglT12xWdRzTNV0yNmi0SB5yzVq5OR1162
JoX6bjc8M0UAZ/2otlcgJ+sj11vDbm+uCG/dT02dOuNepj/02q+2sa6PbaorUPyA
LEVC9y1tjG8rs1vFf3U2YXV+EadlZQOvPHqLw+I475DQqnw02lyA34IKPhzkDRSR
ghvhtE7xOczh99TLYTvCfH9KCrVlouCuCLH3LY+kgpOJv+O6asNCtO4KnjE0AyTC
3Tqgq2Y2vpjKloi/uVCn1XU4v9k23oNPvh1G4Pulp6yqeDmjaUTftlkJCKbYBXUK
5ZCRgO/4xSCEygX0369FL6OUZRPtuskZRRcKtHQQ0QjL7l3bbs/Aqgs0YQWKV6tT
/NgskrJ56+pMoV5f/E8kcQOy9yRs/KzHH/kIZv3fygPK3eamYWVIqqOASPIjku0S
BnDsJpiv7pnJ32v2HLuji3LoUtJT/rpcGAYW5TfiH0Ntkvc7iveEYcDkn/nzH1BA
koLmEHWXUK4w/K3YHTwzSBGrbs1F/TFzOtJTE10rkdqi7RH0LE/9QKQvca/S6AVP
Kui9hWHNQA/CpU9qCGFCPDw8GgikhcLr9+FdSLAfjK0XRggMALQCzyKQcRFgp6pL
7qI11x8VkESLUPmNj+Ruw2Srzv+lW1S57yD3b04JF/mwKOcWtgB9lN+o/ZlbGeUE
swMTvEVaOzcADB1I2+7bDP6vFqc2S9TEAkl7nrBJa4M22UThZPJHUZfX6dMzhvtF
uVLyuwg8YQahoLp5g4dtpRbyVB7xGgUN/EaDahxiIEaaFEZvmiNaqHejbBEio//x
O/L+Yg+ckv+6vxh4ex7jtHnjFXyQGRh1Iy1h4UCj+C+HYP8HH6ssRPQFWayrlUm3
jW/H73nBhb1GKqJH1jWWIljX4mm1VfY1ahFKbaFxeMhyT5BcGkTlry7J+Y2a5Jns
HAc0HORkkqu5apJ4w/Vhj9QTjtA8+ybWbbHR96t7zHb+zOtBHb2thkTcL+yvtn2d
VxkWWiWex+qHlQmQ5gIaGV/hgHP3t6zCPJRi1fmZkbsNlwy+9r638xAMuaZxa4O6
oWMwBlHRGFCnEyCtZXDC+xF4k03GtSSPPiMkb5JODyeNkeBK2dCzxBOvVY1pXXeM
GbjNFSB0Qgqm6ZQT2cOQlfgFH//Q8GLRLyZDTTTfMCcLn17uRAcvXN6XFGGP3XW2
rdfFoHrOgiJU3wblZ8aQQE4CB73XP/60pvOvIAtcsa67nSIFVKqTt8wWt/aP5r9F
J6coovkbVSVenFbZ+ynpkQLeTn6Smy95XuczRgqc0nJfUwxEyDhcm3fYEUf8zTrg
/0ta3a2uOJjT8afqW8lNpIvm99Z0bWji+EvDwWeqq/J+eVja/d7C9tln735Cex+q
10px0YUavF935aETPwAGoeH4SrWFIB1liq60Jvo0CGHwpTDUD5LyBc5wjkFcQMX/
x1gXKTNJC4FXotqVPYq/kOl5yZk75LzvLICF6hnrVfGKGs/xgi/vIa5TrO3jEbLw
hGmff8t8eVO06AJh9z359eL9YvqhfenHa5Pxtofqu8iy9Gdeacdsoe0VQ72XRpAI
g4Mgqj+NueLQuTax8Qw0yE5D/IDSk3FIcAA3CjwdIdTB/+KYkBi455sFeTwo28sW
zZxYO0khuMeU7BYWUFxTyqcIUYW36FsKyBAgAhBcHYCOLizrhetWKs6mdjNB7ifb
Cngf7iMAeRykMFTKeeGYYer4LmhNQEDmNY7rMTfwY9cIUuioGiaTEGj1K5um4nzn
quQrygbc7Ra7vnmxxYJnfua8k7HMX9Zv0MZV4YD1qPh82voS7KR1eUep6NzpXoZJ
X1ej7tURSp6iiqINDaTmu7/XH8S6AVsqRTDUvInua+Am0OPmDHbk7JzhEadnyM+O
Awu1gUQsFcn0mx4nXQaaTzdSNWxqxA6+S8HU/Vc0ajOLZIhu/zca+YPZBPGRcjMs
o9q6Dv6tnIGmfZDIb/VYKCRl+k/m4d0846URl7r4k8V5cBpWWc6ukb7Oy65Kh+XZ
/psqujGvexE3KX2fYcoEygj5ifVfglCqU7X5lfYmkc7QGiJ3CjkmqHOrGGhvWMiw
6YHMnvrP+oLaGQI3faHI0LK3sJwFe15+M1oWriyEQvxGglUzcDsXZFd7j1cA0jE5
jxCx83H98IE/iUoKz489a5kB7ZGxwEcjPoObRU6K87LidvBNgUdeD6LRdgl47Bpe
Pl1/B57P8V6Nyz9LtTnxJKjtcRbcoC1IofdsSKJNp15gXY5juljo77GQw1XgI4N+
jRY8uCnft2dQ8tMeUCf97ENSGhUFVJp7tE+5feFO+1r/mD6kOHXN6Z23g5sa8+GM
4ShDzibw/O3qtSCzl6tpflCWID81rdJ+gRtF9sX5SJmHJ7YyCjTrH5ZTmPVMkQJP
qX+djANHQnrBwSoJDyOXM8sO8Rofjg3pejqlE1p8je/ntJAdQMXd3D8YiTyh7KNS
S5+lSjBuFf+EozS7w+q9DopiB2HHlzYJyi2le9rl+px6NyTzG2ziNYfM3gPCbIBG
LTAFtR4miNpeM5BuBMUcrlF9vLcHg9XOkecg7nfdNtC5tEyBpB6eyPgLXbMWVebo
od7moH9UpGBiVWQLG/IZ39rT5JDRXoj/XOMFSHPnrCBPRWV1ggdfFNUXL1RtkYYg
b87yBEKe8zG5d0XUCQBK7EpV9+xdjCSkYv7Vuf25qW9aNPhKo9EEqfnN+KsboV+F
nWP8KBHOry0cvQkt0u4TMJnAsgq2SR4N/inFiLNEpODbdVBGhdllqhARdL/DMeWE
ysetVLUtgt2QyOqkIy+iValotYWCjOtXRX/rJ7FE2CrTYAQ6pgO86qAfQ0cnv0ER
3CXZiShH3l+GKrfxwY8eNA==
`protect END_PROTECTED
