`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8RFZTdE/PqwX88STWuBcP88qKggbtEn/gmRefEM/rD754dHd0+/4NCuhdSPzVjpQ
Y77QK5XZMMDX2N81Nwn2hthueGh9mOALoHqr61w7ydDB+pYBVgOC5VSRXC7LQ0AY
42YaP1w7u+WUGJgC6eCZT6EXAUR36NBo1TjD4Ms0x1PW64aM1k/rQAxZMmu4ptyH
a6V8Cd7poNkE9mVr7a6FzZDIgWcFQFyxHZKUWlYsu03wnsbvFXoTPoDIqhyVPwt5
Mca6Ox4xnrxaJP/+O5zf3UJIZREZwK+CbR2Muz07Wy0LeCm3Uap1nfliXqXac+R6
gSlaTVl+aq7GkSibFVxYF33Bm/7UlegykDC0eptj9Cu0dpR09lEKLufnZulGgXCk
RdDmvaz68j/Td0Y2onev+4xHRe3TfkYyPhF3f+XnQ5s9tfOrMZuuhIFTHUHRv63X
5oQN64fKYW56fzQgbdUyDmsqMAZ7Z+SGQlE0a2P9qkHfeLmCkwSbY5K70/eqKV7d
hE3OeHWnd8Jpe2H11lLYnhNUnttSPmuBYDDj4EKloZQJOkCPH+4wu9+i8sbgHphO
YWuAnc6eltrFq4p+bXpKMNZWSdtMOtesCaKmhq0HQT//njGeHaLEOjj0R+b0S/i5
chAg9njdSr7/pRiOTkjXopUIRFmucDdgWcmK3Vk9aI7JEiW20ftQ5zxHwBblSTtz
XCrQsAKfnhNr/W50Jd8weEi4nnBCH/vNyrA8fHUS67bFcp7b9c595l+r5u84+jnp
bJ/EdjCG7T6Ddvf5cepM5973IKLhBcs8WxJt6qLIDr/hvaYqHp7ZuT+dULOX24WE
0d0KjwByJ4xwYM0P5MtrkZnYZdtCBYMUERO9X3NVGRQeUTZpf3dqmyhzKTTgND1i
Ch4VKSw9CSJEnt3Jc9E3JynO3Ilc1MgynUSO28kjgvb//x/PyPLjcHVFvHBY6F92
4M8979ehtaxSRRznpz926x829rFY5nh6QIjaMhC6+4zYTehI3W9Hiw7ahqHeubvU
JeVV5Z3p8yW/bzIwpa9VokuIetnbxi5kHdzorbEoBUk=
`protect END_PROTECTED
