`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
B1Co4pTvnNFXVN+ZVEzvWEV14fh40uIFqGTiMsgA3cCjaZ9084jF6507VFygI9ch
XSQ/YsmO3t4woi3XHR6TPXJ+iNNyrlDG7z2OsH23y0c8D24hrIsQNT4Jc5oa+u9N
uqxFqbSikK+SFSx2WuxleR924j+/4RU6gO35Uz1MhGUqGbFa3B+fBk+9c+dusmdR
kubwBdgulUDlkjSncHs5Ed79PGGhAOEJs/9cC7hufM3oGHU07xUxjL/6XuQjSjcw
R042trN+Gc72q4oj6vriKLpN+DAlqmFIyuDd9jliBhcgQjJMQgoNnrmSWpNt3Pv3
6Qs2y7lBK3XtW8YRyrNrlxQBgeI/ll4gffwQkL+AyColDzfvBhd3iTdiBOohgOch
yShQZ2+mhP4VTBG9KTlH79BH7Xa9nPYoRq4B1uhznPTUoi5flrn/ck+pkvzrcNUL
GxnY4c4UUS/aV1U/qqpK8lpA1spSt+j5L5DEGN6VetsEiDrfHdmw6tLKEZ3zvmnM
AqGSf2rRjsoO8zF/xnbvtl2Sl/dgF52CMqfddEmCsJNr6vOVgpoWkgkPXLRE3jCD
z3LQ60o4wp8ebt/pZFjyGqZIqvcex7Mo0g4zEO327M3mh+zR1nSPXKPoMjYWewcp
gxrjnnAC6iLPx2sXlGCihz4mu7Z5UDNgJcG6akHSIu/8wwmFYxjVDoQbQVsq379T
koo8g9NFxP7WQ0iyLsxivpn/EywXON3jk7KkpjCOXt9wUoQ/XDLMBvLbrG+2Jrtx
nKek6hse03xShMO9S9+jGOVsvSEQjc/3BKotHyHuO0TQ+V6tzpBO68/g4P5w8N5G
cq6FDTTb3CXTpgD6noYQJ/tMBDSUjU6Y7m/DyJGTFbuxUiJrEoWieXd0WPx5yrP6
6gHikA3AsuWU6aI8ODALirvPWT8/bSsrBAheU1Bouwlxl12iAWU2EY59Iqpw39c2
gsEG38LNYHl33AIhka+fj9bAl/Gzgdjx9seHYV253WkOXI2n/WbXf9BXWaprgO5L
WX+BIo81XmKo0QmEFsYLCh/BFhnHrgwEtocp85BPTlgSDYvhsG8p5lT6dzuE08jB
9o6jc6UQYem6Vo2zP91KsTlY2al67aHqzc3x3MZ6ayTpAykTDi1NUI88Mqp5Rpgt
yaZnbh9dUeAIt0ZkzRTvHggKKAtl5B8Zxr1WLeD8uUb2NPODQlUCw/XR/Cz4KLeT
BgmWUdz0iuovB9kRsGbPD+k+2NztaG4IqETNtLPdPPw6zL0CZzXSNUH+acU7g9cq
K0rvoYjfyPj0Ab0iLZmIL+rc7S4D+A+CrueRiMa9Em3fqWsa7tqPM5LA3tIcwuOI
n3lN1WG3y3CLqpCj0wahIsNtCw8tUoGqdQZDDmyNYvVaZpqaIUdz55Pw/ZPbu2b/
doBG2bjLZlRujH89GBlTn3XnSlQx7jDOq8RQ6vWz5dX8hhKrl+WU9gH5w/Kww6CR
8EOscliLDFvcjWXuVv3jAkHyz8edI/bu2dhuXmXv8kt+hz5IWEM7Wi/svGgqGwu8
4Keuq1um22aKOCrel6aqP1/DBjUKjhRZzkZ5Gx0hoisGaSbRE1VQ9pQ3bIgLMUno
WniRVfH3L10o8QYHmvdn+OcF4zx3rtk07TboN14bDeSG+C5/UfC4lpZvZ/EbUAwJ
6geV6AtRtmOXZ104xElKv5YO42PTmi2Ir0WsNy+SyirX7OQsh24J7PRCoYixKYnF
c6yxLHmfHLItEQHE63eJrJhxDcqeBRR/TepV0bSTedB/GeWotYYLEUvkfZLHq23p
K6hV6QZ9hf05GJU0VqXPIFIqloUGQaGwtBpAGypiUSKD4aUuI50VhihrmgAmhkkP
7M3rJQg1iBGzqPgdbAviOKkWwpNY2sj4gZj9XAwqKgbxzjYYbRqJzrRsuNCwV4w+
Xr+zC0lOCTu3M6PSUTMK8R5r11CO0r6A8s9U9PvRXIoy++r5PHtIr9G+RD0rH7Rj
m0Kdwv/oVXdB6/5Pb/40wY7uI6PNNwhCBlLFbHfQOiGIbo7vlxGaUGMeNdruBX43
IhNCr8ggWuBYaYUUxNmtrlFpTW4Zj1CD6f4/dH05BGc7Ow68KVHxh9aUWv1seuzm
A+8E09r3k/LYPakBoXeo+5D5jXkM4Qii7ha+ODv0l2luC3zBG6D/t/D9SHOf+nNH
nVasHm2IG36188qEpcHmr8+VHgk8tBKTXR7BKjdy6EFa+k09k3zopMi8U7Hl4l5x
qAixhoV9+EuLFMnPdzcSuMfEDjE0gSYr7Ism2WS+V8YD8dGV4RZh1H+bsY7I5a4m
O/cFdeoZKV/u4cRY1iYM9/7jT+3QXwV+gC/mwcsrmBRWjZq4Q5OSOwHrT+Dy1fC/
gy2fbWiu8AbMGu1/M3Ns9OvTM4GwHbIGiwKYWrcg3j3iKKdetO7qPJsIEe0lfNfl
aIzhgpAckdBtDVCXS+sBnLx+n9ucMRHbOk/3Eda0PeALzpTZfXu4V0ZjV/Ry6FDp
TAYVnVKCuW1AfI5xP41Bas2fJpVn5MjkmOYPivX8OFqaD/pYoTlkNMoQQqys29Q9
jIQMwTVd7wOxgLexUFMzESdreBFXnNgVTkDvOU8oE3BhfDUoIZFDlGxN7vzusiYK
3F//NNOPqXw/pMjCU0ExiGFK85nUjZxLVnmapP2TrSgPihMnOeLdkHvAFoofYjfn
iOQ85R4Wyev160NzjN48BQMNGyEsanUtEwcH+cIbz38bAVdiqbQEeQXM0jwLuuwH
E2VZif3ReUh197+Nusaib0So2I+zHPod27yjF2WV8y2UakZuepuF9P2O/zHY3Yzn
RPXQpVbs6IdkwNzErhsKSFc7MxNu3sx7A1xoAWG5Zb29wZfBVxXPmux8Ri8O8qut
UN5FEd/2FQYwtwSZdZi2gW+lHc77wxA+7b6/kZ8LBF9/j9Ev31hWyJlV0tnzeaXN
0BnT0t+/uHElr2PJUl97FYNQVIQhTK3zRpb32tViXegHpvsbbio/6Ooyf7IXOwnT
/xGf8ZBh/UJHdu3rQVqD52Xp7U/BFZ+MEFfj8HIO5bmoDuvnbRcn/FQlPlQSY5Qq
i6qdBBB672OhhFfq5PVK+Mw0kLhnRCeTorX2yN9xaMKN7Ov3f3ihCzb/4Wq+ySp4
+wg7KIutMXyxFSn6tpsN6oa3vYL6s2P1J0wqOES1T2RM6vpvDDrzBv/VUwh8Ulj1
cB+dKk/l0KY8qoVozTIRkZ/ZRa6sxQKBfLWT0AL9xHQTQNHREZPkYli5gc++bNYS
QrIkOn9nk5RKlpYwQ1wBVaiGv2VFSIIgelaTkzRoZoq9/o0tb1E5v7O9jZiXdNTq
Eyp7xLsmYfr7gfM1bsinhZxof/RGt0x3wNvovxjzJD1a3BPyD7VzL7Tgo1WruxQm
atPzOoazrJC4ywxpW3iyXMb2kfPw9PGJArhrtpm7FkMEGRhlJ+/wMtO6XZR5rFJO
WSTO1jJZIO9uy7/SIb3/AWY24vn8MhaTZWdoxZ5f4gAFpuLQzLvVagp5RpN+YHSv
`protect END_PROTECTED
