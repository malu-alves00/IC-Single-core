`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
T57Jmgk08kqqOMLqAxru0bJr5sjc/+IGW9tKpgFiqQf6VKhETonrhpN+W/5cq164
Wr9/gaOafridLNj46fBZL8FWNGQv8+VcQoUO9DtxQY3B/QZIN+Psf7SNdbhdm3jQ
8ZSJwRDD8b8bM8S8llqw+acDexAPVmmm2+engP128L9/gqj+E8tHyEA/AXiyUf3r
VeHUFBxlzvH79ukVFACXl3TkQ17zf+/ourTvT+iOPV3JSs1V5ajqHJBS6H9s1Ucb
MX3ceZxyvjLEoag1TBzHwLZfvAeAVZQE3S72b3CF/C+RQH7Cn1cbLj+UhuBQmfch
tg5GcivbP+FmIya1awPyQuCVPZL309Y8tgD50MnEg3X9EHgpBHuXFiSiMsGmf8Kv
ga7EwdRkrTx2Zaww1IlzVdjwOl+DDz7vu4P+cT3l3qBcBXIxGpODD0fru9YWhTO+
9fjAJr4nXX/+/0e+p5iAwxyiUUsVexiexjZ4vhMwApx+1/Sz7AQPjih/sgFz+JyQ
oE131lMKhpjhQEnBf7VjHkNoKKqnGM/5a4MNsUYWnpp+zCWRR+9aQc3p7NmT5NjA
l9i4DhVd47m0ynkA9I5lz98XryDn8HPKui4XtiH5F0s4WcqbqIXVu1ORjNwVtI7d
/vuKBVem8xRFeX4foF3vXOeO+/hqInytHbuhrCnmd9gA4YNGD3I6a3cp0DOV/0n7
Tl2gOmJr3bLYV4B4XBxtVxaY1upJiRdJThSDEFDyU8V+Ep7msUoiRlnC9N/AhrhQ
zKCo7Gir61ISxW5v+Mi/bFzQQyv3kVQwdDEP1K4Bcvy1jtBMpC0Iu54e2yI+k9dz
87d45nJ7bQoHjMC0CeXq5hPBs+Wofcl87mnkFJUQ2qDW641VTfNnVtgGtDQMy1EH
`protect END_PROTECTED
