`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
G8boFZW4rYjIqHkXXuZ7Joi6EjgbxDh8wy4V5XvpFf9meJM96RpLnOBhvRs3iSdh
TRcrfnBxjVdid9fqRDuOVN3+nlY0sGpAPBAO4b23zwH1MnAfPaa461B9p5ydfEk+
vbrN8NS8dJIq4D60zYQNUBZQzwUq8/aZe+czhtNeHXMZc0Z5V4hVGDGKZ6yrQJzQ
/68b2Vw/HYicSxz7zTHsSbgi76JsmEiKairEVMwBEKr43WlSaPyw8Ko8vrekkqtb
/f9ppkA7QRLqNIlU+Lywc1X3y855NRLOELHYmbY1MA4KfvD4KZ5VwrGdDPkUOzfA
0NXiB/A2rJ0fHIG9RySLZt0vCewlx2PECLLFAmwTb8M43H95XhNWwlfYrQOZ/tm3
6vFpnKPKGBC36Gz3pa6g6ev7WA3sNeGH2TxIUgYKaLDDWGMOqkCuab5XPuTrQQik
K/nVLnGkpImzcCR1ATUR8+CM5V9au4rj8p847XtMC/gwmwnFgB3p2nS85+ts98Vh
uRaXE8ZBOIk+tEjukVKdPUZ6PREicicr2kgAyE6TYSL4qATPYL7kKV20SPDpUgWw
QW1oc8ixwjwIyEiNEnPdypt8Kg6j+6KCNSBEi0sQma5K5teuMadWz4yNsK5+3xXK
zKyVoTNkzPGt6nM800uE5UE35XeShWO9YGXwV1iDGthXwiGa3DXIuYPhlOQt9ZMl
qUKa09VGWLBzlBqxbwTbL48ucJ358q+Z9o6XS+gJIYMnFwiwUEtMOch4ttzcPjYI
n8yxeXTkepJiQFsGAgLkdXWh9QGKmTG4LHydJJmIJwHBTasDp9w0jlC0a/iDqgCs
pAIWmrE6lUduCjk3v0GQ1xv7lhR2xsRn2xE/xul4aQIAgpfmAav3AAYr9abPU42E
ukvnNqco/qgxDNlZZcQt4g+uG2AUJ779do1iwHR4qf6LmDfT6qYXqQdmhQxVheM3
rAx6yAr9MVrA+4clsQgcy2zKZqE0ZB9f+6BU5DcgrIR6YyfLiIH7PASkVMVZklfl
2Co1eJ3tdvNBbfXLKjxvA9WNJxouDxKTyg7/C43xT1J7pqkNVmrVEMwkWiHizEkR
QmX5W+qjBMLbBQLK715+F8QIzzIKaeOYb5CiLha6NnWw6L4MriJVHuQ2uZzhSMBl
WsTxFJzKuLwFysTLBQ/OR3iD1drKH5CSsSyNLgAR6q26cK5WdKzi6nlQWOHmYEdJ
rxpEatdzFXNUxQQsuxq8qi80556E4BCtSQZIdDJd4FbJmpEWA1kjVE1BvaVt0Dcm
NRAi96QqhOb7MDS4KWwINkh+zryFuk7GazYKStD+RR6cjSXyRUqp5yOf3GazInT4
xbRqZaLrTeeNF0NGTxPfVXRjckKBNR4r2aIMs/j4wmJsFxLLO6EKBNyRHBokN7nU
lMrTkxoHm2tYBOKccXcsxN7E3RxWe6yZ7EkW0yZoN0b25HBXjhIRthe2McE4Wj14
fcVkR3lNjGO9+0woseoNH5+OTVLiNgP7TnrlYbKLraIwkzoMQVfvqaH0z6EhzzG6
3u2mgVwol70RcLh8eDzHFvBKhV1YQ8trVBWLUYTFcadiJUg/KEUkPRE44BrVtplW
IQ10wKIb2KfnGyjKsRJiGR6aXKO3co4CQYptDwOZJ8GVFiMcdEBLGuwewbGE968n
7J40+QmOEBntB5b8S2PkrVVTM16eQImEgt2Ouz1Vr2JrfLXL3WmOW2E3+boUeMhd
RxxhsTItLdmtPTiq7XMdxoe197X73LmL0vNajxecwlk=
`protect END_PROTECTED
