`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iRHn9/VqzSCXyA+jS+t4M7E2RH3O281J93O9HyBV3W6zJBvkfpAx8Y9PgYkPGsTu
vvndjRPVe+1GuZz2p3bVG675jSIqA+f/IU5JGlp43c6YRSyol9946oi3lPEjdvqD
cGIkAwfKuvqaYsO3MaVAlIJVxWwM+L5ZI46IANjCy1qUVe8KuTFhgiCDA6rT6/tb
DIjePC9B74jGJsiSVjheoXgaBfVZI58uAMfEuYCOvftz8vTuD0dN9si6VQMMrALw
YGo3WN6rsy6F2+xrQFl1OgWW2emJsiaQGEF3O9PnkBNszEpzn6pDGAYvmpMJz4R5
twGY0+z7V7dJ9dpZ+7CrAUZzYXeWKYxQ90kI3PWmK1Qhkc4AadX82/TQVIZhfZ+g
V4s8KIBUnzCiVB00TAakr72sL1dizP9H//r4x7j05yG1KKBziD8ckiojqM6lrd64
ClNJ6vJRiIaGy/a/dzSs/Kpp0NoHx/bZAc94MnZH1iieeQlGLbq5NGiAqnM3IQQ5
7UhX/r1mgXkBC3MOudt7bLdWQR/63ZVTy1TRjJkQIa4xSeg4RoNwXbkaJhRGOKMr
woj+FwVo/mRaZaCttjbbDcCMkBo92b8GUGrgJQqMMMojXVcYUaX8kT7cApVmXrId
kkgi0cLQZcxMnOgFrfuXi0I7uNoTfos3/fM5RyEx8RdOJKEhGjMr6ak6m9haF/0g
3zi480WtfgfROVfjofzVNqSgkbRFTlqu2kMc+3yRFFuRaeo+dGxR2Ixd8UyihLbF
Te+GgYj0f56XJ83/j2W/rDLRXSr5XZwhlzIwcQ5qEHFotf2CQASi4501xq/tsjwl
o5EGGvvXsRxRumkxI/oqcdPErXe38McBUbJQQJoscmKBzBPnfY4d31x6v4ebVFag
amQEolWWEQEKD/YjO3fzF88RlcIJS0Aypb9D5GsIG9G+o8lY7V6azn+cioD2YTk4
zoOE/0qcjWfGtTV+1e1p1LMxrJAEbjqjDCfcUQh/HNGRPSeJtrf3ioL3lcR5jxo3
ZROwnvHiII4GhKpL8ccfDMGU2BDmH9JYREHNEW0ypTnt6myUtT1UgBHr/CCGBX0w
o/AgWdYj/lU9e7nEWKSna83Cf+/9HYMRRWDgD6GczCXwhGiQT1pFXl0caZNGMlY4
UsV8S66qZ/NXu2L57FL/iKcCedLvPtMPIljc4XKxmtfL8emPNJnnBWYN9g/9R3uI
j1avcRkPfCZtT55c2leEFqwYJcgEJEioeEYwq8NXx8ocdzVcaltB1OszwZLz2y0H
zo+la/1d1Lq2oA0Tcx2/k5C8Ak+lgGRPFzICkPSBL7efaXqulQ+h+hbJh46p3Btf
ndGfhv3wG0avjPl5mtWfD3bUvvLAJCP4ictBfwibMla/wK742CdFRpaxcVESbkq9
FSmen6ZCOXD3euGBB0vyWUsJYjffZpUerHNp7QAOmrecFw6FHMqZaSJA61RxkPGS
87l43Bfca4uBmLnl/6WL7nlvWLNxb2eOFTcdHmxB2AbsAJiMWBq6MCJEzJLUKdj4
h553WEMhTX+Pd5bTNJmTIoIhSXt/uMLmJXmDCm+Aiw8UI79gZ/jHAq8y3gyWIGyR
EPEyZx73wpvvXeRRecmQgoZXAzoHebI7t6jc+Rul4Am77IzB1nWdYDDTsgWh1fNk
r1zFCu2Zg2e71OVE+hkmBkQSIdM0zror3ohf/VOw5dDJz5mHuMsieQwaPtSYB9vK
vAnKPDCMOia4bQd++ZTSiN/w8GNjpeUgGm3k8UcEldg+ULiPiZ6v2xwIzWdVNZ/i
GNCc86MEL9ijF1kP+Gqxjl/zYmo+EOoBDHQ4YpoeIN6dTKyKZvy0Zc7r2+SwtchB
TkVZSYkUXzoy/3j+LgIMGqPgxzQq2cydZj0iIOHGuFGkwqB1qKVMoG+ALHkAjCJ3
mIS/BHP4ahHtpbgv0q0p1qgsLD8bHZjcjkdZUwYZD3s8tTNY9sj1laxOt8/JOwja
yxZMogyN7fb8WaM3RhDLog==
`protect END_PROTECTED
