`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rXpziE4dwLzRghp4PwU7YG2M2FEh9i9ZSoPDLRptTTBcUhTQkwTYcN/Y95qpoPPg
eLRqRSKu1tckBKGpkgBWdKrTAbZuh7LBqXu7zVG23kLE8Q2p5dBnxMqqVj25YylW
nvt9A+51/SDCZc9u8mK/lPhA7jqE7nFvtGMSfI5+vtWbjumgIo1gp0Ul1EEAN5P5
iMeWrd79b7DggY9dvspsU5StYRa5dTQYPKlP5/GKr5RwgqBGfSCCnda57OJ+WutB
mGVbRyIoWzSxmzL9O7Le6hU4xX/Ba/gyg5yBv8upALzCNosTTGhHCf3LGkhG58zY
qEATWnCJofYRt1h55yc9YufHTmomnnswSuuPCphmXsGqNcHSx7nXMisXne/y4RRX
kBDE2N/utnQXXU+vSvj5d6+wtJe9YcXs9E0cSW9M3tEG2WShWNCsULrPa3N4xFMz
wnRHNPd7GcLL0lD7o2wW1jEn4UVTMtLTLEmbRiOVmHTHEobsI3ghknC8FDkLE0Qr
tRQ4QJwAEgV4Riz8IVry5WbmM+Sfa1tJgVQHSYutrta1DibYcMp5oQskh82zVHS1
KR+MHfJ9ZswYVVO9o12zbWcF1bWvtpTyd6eADJUEfGTq3wIbLhLshXB4a/IyIMSV
732NIAzkulLZUm/7R2l/fEdpZwooRtuMEgz1XrSFNR0QGkirZl8yvEnB6bedPY3w
EeW6ZNY7XaZDimAlXiU9yXtZf4SP486FyaBUSvchG909VlZdoHAFbpcwBm2W6PSj
GsuaDzMGRWnL60cZ4h8aBshw+hgK1OfnnjfUz6FYlJbHQECE486Vljit0mr9HVuG
wiNrBE89XsI5pXewKhk8VV5GfHUEJRRionAGuRB9mo6mF2DMs8tRHHGcKsptjuRw
doxkJy1iJIG2leKV73q0IBZ6fafeV0SvZn9y61AMuwAUGEQz9vD442cRyRfVIb9K
0rAzIDnP0qPt+3CgGQLHxBQ9S+taJowGZ7A504OnEjh3xYeEDkRJiFtfR5592AeE
8vb5noJ8WyHoD+jWdvLyH5erjyrcUHB1p+qRT3D8ezUbEe7ItkQ12+guGdmYX/NL
MrLy9TjVGU/oqRyhMRLuTCQwDiDtWeBHdrbWR2bXjKZAotfMLy0XXkQw6MBJqrnH
QY2+PsAdy7WUhf9uE5TWT9devulgARPb4DaBMtsh1G4QmUfMgvIWT1vcD2PMBDZo
yOUlKpOgz5HFXkplkQPyWWmziVln8reBnp5lFoBRklGR0HCsY9R/h4arQWNEph55
TqHHGA6am11oTmgEVfeu52CylFZ7fdxVJYxjo+JQxKvsLwzUf2weocxz4O05I2bB
ZeV4TFwNXJYClVTqEGV6DXpS4UBHkvKaKJu0Yxvcd/3d7c1NQz/aWhsdfuqRcmPO
K0vAc0pXW6rEx3pEWG2jWLpeIPYsO0NkZ3F9iPCwyIhtnAm1uDDcvJEFSEJUEulL
Z3pl+vwGWtJQ9H6+sT5JGrzG5S1Mj9edgfWQigoDYXc6G8vb0Uo7xelinHNeBCkF
pWyeZxEr7E0ecBVmVwf5ywvGbywBMOcwBNBYSCUGy9jyPudSNlorxb+tylK+cgxx
dA8vOllp/eL5B9szozW36kLPCSMYanxwnqfb8lk5ToRDd9jnWSXlK4Qs7Tr8+dX1
KcEjeBtUGcVj4xex6IjL4fITVHaq0b+STg1OoEmbKHN5X4tMlCTWR6WL2jBpr72m
qsEkpM0ysj0XxhA/zPCWJDFJXfeH3eW9FIb5uFuEcWij2XwXvaBpSWl0dUmBxwZ8
VNNlIypkFuUdM7VS/HTPRWbR6kmy1WE3/fc492IVQpPs9LuKeBjGcn3ntKy6FdiW
6DYtS69pOuPdaIon2f4AubsVkwoFVfeQalD6N+i8Y3h1U5nohlrWx46JXZHIXhKY
OcGGLaeZGGGjvefcdVUroatUqyKEsWnVEiDOgZiwh9jsymIm8KeIMRc1aixB8p2l
l0S7tsyPL4u7UTq/20CA3cWkzQKs1wwSZQUs0v1zwYprdKnCRkOmpIDoJY6P/Tqk
wFEkm9Vsc+cCs+cGo/6RqnNX2aapm+YfQQHL8fanTsAhIFUPaUT1u5KHBDF2tj7g
j+rcIb9zNazsil5boQkz0Ct1+QXx8qD/s3JnS4J1f/MhsHSEEC3u8wpO1SKwELu5
`protect END_PROTECTED
