`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WZ29OVJA4/LtW1WFRaoNhj3Sc85aZoYyQmL3jWTNoVs94e4ebe9QJAj7IS9C6VwR
v4BQB3azHFZUKfu0zDm51N3hU4di3zGwcG7NWfPjz2Syyf98st5uj7s7qYJGFwn6
KtL7bt9adhVrONBgXYtGaCk1lKFnsJy0HKE/FQrn3+03rA0QDOOKknabvDJAgBna
4IXRCYbzLiUtcAHH9EELINeDdvfWrOFfZNAfZeqH0JNtGwu+AS8JrA3kY7FAEzWe
WI+2457F1LxjgT2QxmnMlqfGDAtl2zXJwPXxA7B7KsRz9rQOL5fVjI+8Gk5jn0iY
K3z5wVCTAC+0cm+EpyvcF62BwbaYbjWaFScFrSoW0XVRvQUUL+RSxzQ7HI5ewMyB
iEFYXQ9YKS9emsaLR/eY3WbIKcxkBVYHEN/0Z2CDcKhp+Ud2Eqg339fBUnuqefmG
TP2t/iVgYC2Ez/kQJmW5fRgyG8q7XAWF4VMDLYLjvydionUvGh/YTc5O0ZowjVn5
UvamuuMtCWwE3zy7q247e5DUD5hU+SHnB0nHWCWtO8yhXgyDYcqpy5kYJgFNGu+B
itczEESvJ9kO3zqUx/Ss3r9B4Do/ohhy8m/P2TEvxl5Vg38AWZuDQHvdrvxgX1EX
4Oy9D30ku5iSZ5vny8zhFa+8CM/zci5SJjlbrSXt+Lv+E1II3EgoOvvnOGP86bq6
0Z5aeKsUyMyHX7xM4Mn7TPeBXW+cLihAs6BeokFiT6hAgoBcbbl1GRh01CNB5+N0
2NwCkDXqSYhcoLq8knrt2R5O4Coj8v7/h/TnEY8oYxicb1Ku/XZWB9dDdRBY4yea
TNua9YrzKePMW/ybG/v2FRra4Mlnkvj77rfmfN0ntwvKO3MSODCAam0nvY9uzwkg
rm/ygnLMETMEpKCl+RyHyxxNfv85NseXD0XNBku6Yog1rlt0AMB2mLZug+J11COV
ZhoUjMaNDrvrug+/IvrcnAEtrQJcufWtZKzlUVj7uYJdzTIywMHvoEJcixtHCk26
+Kgp60Csp6qfeNvKMUDECziZm273TmDvTVzpImI01BgyY27I5/NhGq+N1l+1q7po
Twh98MkjbJQluI36ZKN3GSWvoWZ2Kdeq1QBwe5aQvPsUVYBd9T2q0X0XbDdbQR8i
CSTUN6oEvvyndU1XcplGHK4fJ75ocBknZoFWICup1dhY5MysQKrFeXcPhruApE+i
tVczQ4zRY2kaChiTadvNPzypxVwMD7YH6/sl6PteRpkb4BRbD6XQyRxrlVTmiZ3C
bdkJ7p9H4v0ef1jzlplGsOLde4xSfbvuK6QeduV382sNHvuEJzGUH3HRc2HdQXm7
0h1fcgKk8R7xpVhCbvAjRE++ajgVRjKFQRU2Q/cImYQ=
`protect END_PROTECTED
