`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lsQXSvg2MQQs2YayUXJxKbFvnCbWK2jQDU5UxHzvIxNEUch/pSIWBcmKs+yVyBME
4JbB40/SoXKQxfbGTIVz5N1yZvTJnZ6oHs/ZmWSScQ6P4ZeI03SOACBbvjm1RPr7
/DOW0mj6MhMkkSR7lsTUDePHCkm8EriSolM77AxJ4Wq/YTEuQnj/Sd/aKEIGk9iz
/b5T1zs3QIqPh4qSg7xwUS7JDcRv1Gtr86X/Hubnm7lm96YMyXq9r5WC8vIkS6KB
l74VQJBf9mPTT/4R0clr7gH3yQDXhKKzjeNFbc4oHND3ROzUHIx8dP/ZPddebMsI
zJaNT0tmsAAGGlP4aDWNzaHoZbqv+W3UPsOMNixxcskpt2qIVnZ8h9z4mxEQx+qo
0CIv6drpYXrlM/rtKP2rSRZOyWLN0Eu7K+Jisle6Dq9mtW0zylW7i1bHGmlEkdK1
GP/6fRwWxfz+qvinzoDePazbvwqONDSh8f9Vab8FsYB+VeyjJhLV63zHH0p25hae
tT29s0TIAne/r9mb9tppQ6ts5X4JaSGqqH1B94A1Zb0P6OoFtHmgOWragaxtlwUe
rgyDfTPasRLGCZJJjSXVAGb8vhJzGIBDCqsDwCAQF54Ka0LDjpzy71H0nafTfUXP
b9tUxvf6RkD1H/feEeuCwW3JG0yFa+E/YW7YnZNfYukualI/FXTDk6R2Wu6F/7ed
QK/vCn5dEWvNWraL1HR77iWmLTgnzMnKVXmzNTg5x9KapuKCoqrjpXLQZdklvaSn
+/gvobeNze2Hmfk9m73VOg==
`protect END_PROTECTED
