`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CkfQubWV9D15h5C0svkWwdaWbyQrTWsT8oW0Mr4p2FNKHkV6/x8G701yUkJAlOBC
s2om925d1ulatRd4t3/pGeG4jvKUkHtvssE+rInG1eGPysxJCSSnGF4ycCPf66NG
rKUHL/sBKYS/hm0NR/OMJGv4paib97tZw6WZBg5PeB7ai8KQgTESLE17PbeF75db
Mi1hrGgKyniX34YWYnTtAzbvPGcyyQ2LtTS5UAG4kNnPV0kfeUjwSrumZexDHkNS
4M7tHkfBNFuF3JUaLoacu486sLA3CJCjqyGyS6FQ54y+9Yteo4uH/U1iS2F5odFn
CZX01U2iOuuLPrw6lU9kcGsY8oeak5Uszoz7JPq7REE+vlF1Pw/ROO7b67s84ZhM
W+7qgJu/As75uCmBJcUnho7mohmKi9N50VdgbiP2U7rd5X2hFoqmM31l8QDRtG0v
zEXFOMniX6u2B7RsVHdjGF5/7zY4Jk8sNBbaDGMn1gPR9Zt2ZWZZGz380FEzY9QF
8iVswxpFFP3RrBkk02YW6mWE3F0XL3WsJRtgxwSlBtzBLjyHJmF2DbZTJRh+1aDB
7sqGBOdpo0SPvx5HryGui4oR3CngxxPmqXr4vD8beVD69eKNr6I+taHbhwd3NmIR
2qwGQ439CdZe2TyHQ+NxcLiRkEMlB3082116Sbq55uFV75tTfi0iDezy7RqwpFlY
WQjbzVmyZyeqhY4vJbPPqDMLhjJWcuDCIUlDOhQmen0/Fll6QbDgyS5OB3O4o6eZ
5VCikk82LZ4fFwYaMp+p7CozuR+4hwEQtrmntCiNHCJSR+iJ34VRb518UvP3AwzJ
jL6i6SiF0xmdsqlYFrwGCg1yGmX1TCdIWj+L+hJ48QjIFmiMsHdksDvIdemouh24
`protect END_PROTECTED
