`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qJAdF0FI2nrOG+xgi3nBbf7/Oya3NeDHFeLv5HxbtnndlvGxBqZW4r7lB9Ehh5sw
nVp8rWQSr9RxaAPFlxMRYeSBrjxjQKAT3k5Kp6CkQHUezetQ1iwIHbBaxG2HeikB
eiejGTrOiw+YLmOZyi5m6YlpRVCo/MZz4qX2ibOvlYTsvSBBm5XLag8TDex9Gzlw
JuhWlyXE9+Sa2OetofMZjGCo72nvNgv6rPRod8nraNW+2ipmzE8v1l8b3uBYBxc7
PlA8/Bw/0BMu/Yzsmp70UXW2zXwJJqgB1tQV4K7st9claI01UiKgTmx+xboZQkix
C2xb41OhK1fFFMjj9pHSqyTfn6PL6a/VUzoiFjERl3jJgukUD3pPcMDOVFZVhO+b
XW6ajZm6OD56EhJmhd/VKyWFCyB1XdOqFkcPRYlixOb4ETg5axpqwCt/aQfU566K
y5nxgjB7mTWB2j0sD6/kSM2Vg8wKpNvOKOsWUCGas2BnqDp90hpGKvjMeitWuGve
Rr1JGwcZEnTGUGTCeKRoXtD5ij96EGQTfoS1qcCPKQwoD86IuKXg3Od/UQeGtfJx
Q7Z6Xxb1L8dJjHbxn+dPRRUksELwCLY/iJ2wx008WrP8hY6Lx7hPdPh1dKLB5icF
uKHUqH5XUMY1RqOLRNdiAUOE+ZILTarxg8mfCeaW2OeBoYJwh/AoO8be6bD2g4Tm
kxJcvwRk5MM7kmgVF2qWjXH3EFv5yFUvPGm8JqnhELMpdZ00btIOxKU69UZqnVgm
8cwF1QjPM2jASsDPrb9E8gM9GdUf/Om8mo3IWU1QWcEomTWRT76JS/X5bQjGPEhc
ZQBanWGheFdpTXtOiNLebajlFVLxd6CHzLRZS1yIKc85j4/Mu5A3BPvcodpRtgm8
GUaulNCA7WRb8h2PTqc4jqCheZar4oUrdSSnTT/04dJO8enyoumPqPdzEULSsL4K
g3fTt2jSp3j8Kw/EoaOh2no6i/yprhb10//g5cllcsLewy7B0ky4bo7DOuZl6Mbb
BWH8NLFg/3Tgs4lHJ7veX0uSch1nHJ/9jlqf4XVTLc6m/b58+SFZaYQ0eDkKbdeZ
L3/1R70dyhrB8fzBqkf1aD/uKk1fJveCs69T2wv7B1AKQcKqzgcdx1xNSFWjLmVv
ilD8uerz+HiHoi7GVB07IOPjPrWF1Tc5sdBSTiHexZoZl07cG+FFfvC0W2FgoWyI
GYKOwMKazPRg63r7Fu6+HYSlWkTvSKiXLg9gIiYKQFHRltJY1maoijYl0IIwcrxP
i5L0+0hiTS4CwZD0HoYBZRA/Xd4yzMZu4Pj0FNO94nno+odtjjsFgG8zBxOtio65
WKAvXQ4uJJBqAPQSCT3Ci/+ZJ+iMhBirqdC2lQilQkfQqBTSM2hAwsQPq7ecBv+4
dFTRGp0B0mM0RisjEvJjQUGV7q71VaNHDe70RV0doqlpBWkamsn/ZSiSZ3xe/8Vp
meddtRNYBEM4ZprmgrSF7uLAl1SZ+/ibXkrgbNsB9HoUDyDMx1G7FiLJRsVq+pBH
0avW8Aixr2kamj7AN9QlOK9IYvk6aWmhXrQazYKgJW/nFynGzUgc8BuST23DXlyV
20Nj0D3il3fCqwv2BmWdtQAa+W4C/O5qf8AziYVoCML+YuXd9SMqEPcG9UiHLZvR
JUyU9aucXlhnQi8mmHWxuXvj18/LnIG6ib1S613XLXffnfRU+5ToioxWfJ1VB1gS
TmU7Z3pXJe3MiYDce9+zAtu43oZMKZkhoC+LIIFp1u2qAD01siycL5l5JYQePMJN
YStAqvHDb7juXhz1AQIpJCpi46G6ZCxpTKg1ao2m3Na996lFuiX4yMz8XRtx12gP
TdWIsHf+vz057pXYE+h3OwyfQkUp8SgSGKpsKGDcJRK2rhSVbTeRpDx92LeI9HLz
d2yozyBP0zdT3ZqSBp/vQuEDmvo9rPopEH1qqXSbYuyldnT/lZ5eqwLch+uon2WG
Oo/Z2hpLEaTmZkM/KirPJ7ReWeBWY3AaxGt3zz2CXpXrixdagH4yhgAAYc5tRqXm
ZvKqn70GEy8wQVbCE/hGWpuq9tF1QM0cux7xXBXHQ9+9ZYQqlr4BcQaw9LWWoyyP
oQq2YfVCXCxroW8Zqf4WqHbN7qY4KWoWPyaRjv8ZNZQ5XK2K5XmVbAC0WguI4xWe
OAlDl8e0A4UZxiAWLeWIJJS257MuBlCQcxQvzWm/ekGYaW/IaJL+F81lEXEv9qUT
OHCG6vHUUzEa1WPYA/YsSkQisu5b9brSvewNymvHqRLa+2tl/AjIjmcl3ALiWDZt
tGjBe3UoACbO/Jo5vbuia19JMQ7hxY4A9kJ7Hyh/IdeLQ/sXwDPKRDCwy0JqsLVI
`protect END_PROTECTED
