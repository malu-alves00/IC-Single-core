`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
X/0I1Bis1FhyqABu09lN+kNlIXoly8bLaS0xLsoI+5V0ECJopZZcoHhbf3E846GL
phSwXpobG8aVeqaOTmiPw/N7uLK3igW4IiIoYn+QPPGDCzlXpoV6A4CkLicdgLjM
5g+H3IARBXAccv22gx146MBNS14zBhBLcSlG+5K7rmdJjArxZ0SaqvGYf8kxdYxG
SATM47b7B8jtVUFCpI1ugDu2jcbKrF7v/lVO4UBHJr994AwlGNUdjqSs8u2jvFsz
Q2lir3uJkdOZjOoRXSZMdqVKTezkNVCSupip2Kx9f2FdSQsYLdm54HGVbpBEoh5q
p7gimZrvZDTZPp1u/9SoLYI1lEfqlQbnL0UUChWOm95jT78ZU07zt6wr13fpUg28
OBLe0pISzM2GEXF85KCe/FXgWynxYy0Mubi3UGsN795tNI+OeJOeZfzmCWA+6Fq+
KqV+hJxfQdKLwDuqUSGOwe9AKPOf1Hgmm16D2bCbvCQqEiPp1uL3m16ud3SPUrfw
qjpTq23ire9uZKjrgmb865TFcSItTU7YIEncdigkvHASMhyZpefXUHIDztlPImww
MzlHTiWkduZpXPX+W3PE+nmRQs+nQIdJJ9aZPuWN0yzlvFQSjuHEwK50dHUJNe7L
yRhMZDl2hSGWWPpmnO5gqSjAhZlZ42F59cOyan7HA7QcaE9WeuC3Bjb23uUZQkGq
nD2dEpK2f92ZesTRDHwBcptle0YHVe/6jfiQJRSQKBpNko5aOQYulLGSXSPCrom5
g1j3rOfqduAU4gAKoPJ3Q8K90AlxJjXk4hD6jA7D8BLi2U1obvcJAkgRuFQEeEB8
t2GWrjyHvLvRgR/m9FUKV27PLk10S5qLb0bp0FDlfFpQROxg+ivCOLyNCDPTnvMN
`protect END_PROTECTED
