`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
h/XOs6+IsA40l+yhj1k0w4ZKQ/jOshFZIsHB+iWm0AMqXMg+5kHiINDhZVF6MUKA
HWgovoJFuutgUwzDnQXCRf961ex9y7tw3XzBXNcio6a9C9qqKOStvikAtsgaKmL4
2pX35VdWtw3kfBvLuIbV4KOel52JjFHYqQ6TDd7ot+FlIHmF/wtF5K7C2h3qreHw
orrQwzJfCVZeOd+WlAwCiE8gg37h/xXRlhh1fQdOadKXyJYmXRUeHsLD7+k6SDjX
QWE/bOmktGb8HXhx9o9OpU9BgLUMnZRsdUvDkNwDQoWHOK7F9Sdp10keD7B7vc+D
lASg1FNtLaLRGTtMfJIfVBk+XqBCibJblLJ26sKdWUvRu3Xmm1ddN9tSKWw6C5r9
Sxk/Xnkc81HzFCKGr0qc4BrasmrIvgSCnd+HhFbaWhPRt1AuUIRhg6d06GjMl3pM
kRbGtSHjPxCIhnIG4q50wE6YMGjyeFZf6Z73PeiGMpk1tsnDHt1Cv0mLqc19RuNm
1v/09pYszbGQpZRrGfYglsKy8iT0CB6UPwSIdXgBvSr0FM6vI2tj3YXwImpLw2TJ
MT3xJSQDCOLrBWc1ANzmaxfoDSF5wZWrMKNawtk7jyMyQbpvYssk3NqjXwA9Q7k6
rph2qac/DElD2I2UU+mzDLF9wq+VGiIyswURXInp/iyu0D2Oz4E7xEVK0cAEWl3K
AJ5O5ubN9cezGD1N0bSDYQ==
`protect END_PROTECTED
