`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HvVqZ8NdAThBSPU2n3G/zPnPyDAxgRhnoZkgIqOxKZGaYC5qx1A65x8r6+INxU1M
PU2MOAsd/sb1/F0uGNOgbjgFv80H2v9wTe6cEudhXlg2aSqdz8qSpXvtPRO0w4by
D2mqhwVwHQBaC7DQ6vtlWP+eZQrjamLCT34N5a0payxcaCcJN0UirBOTrlm6Ezrp
pyHik8tTALJRVxvuVLpGLOHfrf2KVyYHbyby59zERLZSjpakR/yir9u/doz1wLjx
f22bavwbZwT3nrKCtPolTMJnCjF/CXpoJOU6jwzEe3UI25Vow5imt+OroXnQj2Y7
0m3Tz84GSKu2u3eTTIpe4Jb29kwJYP8PvwFDj9i8Zsip2RLIPk+1PRyjCEX5j/gX
OugZCUZi2e3jbf0AwcLOQaUMqBDO36eRUV9WatxW2ee9tiFEhTh7JJxkha9wMRuU
5yK4swCXV7FoqgmTBtqd7Dh6sOzg38m6CWS45930Vkb+mhbaWffLA+J/wseLyd+y
U044VSbEU3DipZ0Ro+W2x4yyc/cBzYORZpI9oPatChjPJy2HHh/dWE+jUSNZdv/z
85QIRQPoL5JSS8G+uNghRyNB10C/MI8SWAUp/NBWwF3E27J++9o4LCXMcRdRw0R8
ZZK+nUhfUhlqBaizkpVU2Q==
`protect END_PROTECTED
