`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
I4rf+EoLpk03WGtuXo+iSU+JHUPiafi90mQIR81e4mdptIkYnsHkBWqoc6dH+pDw
r3TvUYB5Gg40KP4/gsYI5LL9WUgYI4J3TbangmKRN/4hKm8tnsRkmW+ExjNHr3zR
fKwj1exugLsc3xufF1VVCusmGpPWWagy2uhtxgZFDL7bNh9qR56/ofZSwTxcaMet
1u85V2sQdK3IOc/r3ZohrJY4WnkSAuJqKQDxbd6rQ/bDwNn9PW/K6AOhCQx2QIMM
7SE2JZd90j6d1nzmiSO2to1qVz4uMgx8t3paL7sVx6MbagaCgs9GRG/KYUuvS/UL
pPase9jLMzxWLjtu+caObjFSZyUheTNCoeehyzrog1r8OIMJm8D2kgNC+27QEczp
es7AWZVbphMFymVo8oqnjbCskFWRJsZHlAQ/oYHXlv0cQ1PbjaWFtTjsx9G6rQco
v1w+9jOZFrFg+nTGb1S+pS0jX+Y6jZaaxoUHCNERcH1LZyvtf6uVXG011jyXHqma
ERTfBQBVTKUfNuUWqsDhZkwaEbFtASXsyPRR4SasDGTOQgbb24TsDJoZW86cOgB5
FE1up4jFpjWy7+DcMtVLLwO7rVEtYYaqXYKxJKXzSgh1+n1woztYEieOcckJw6Ge
1/VRzVpOrNN0ho8pAR/LKoqhcdizl4N3HXBDlhJkhDQRc5kHRJD2B79uNRm+ERRf
yJ8IsJDF3tBIiJxokXZG0jsEDMkVJUeuP7nGTRInh+MVzDZXJzxuvPqRlwv6ytto
oK7KTyEq74+kKpJmLcG3gCcx0Jy/iarJ60JgmFduQn/Z+uzUM9eMMEDVJ4EFhkgI
lYaGf55sen73halo5B2uUpln6JHquunExivU02kx+nIeH/8kq7DVK60Eu76vUTI/
smW/V/n/UxhW0pZRNS2ib/WNpux/WvjAQcEPMhCeJf831CkrPsqLwzDxGBedDhkV
8dzakyGZvMmFt3q9lkimip6QDGYyyTZmbOMK6uu5t06qweW8Lr3ljG7+w12rZg3Z
bc4WCB0XGlC2omGgk27ITVqlp5Nn7+y2TEi78z4+7GIx/jJHbHukhlKGrpLasqFe
Lx9sZXyAYjt+Hg0JKYo6o51GggG5iA+OtQWV7BFxyfj5gsor/BbpIKu3njGJKERZ
197EIMQtDyatEMhOhKqco2UJMYGr/XlpBHhjhTx5TFBbdNxMD/pj5Qbt9wONgvDm
81i4czUfIaUBJe38d8WZMJMdikOySoY4piIHe6Cf/7I+TirowSSQpRYufi5dEcLj
xWU6pmPRny7fsvnMeVxWciz4FHydl8vELoVMT7dV0hiUl870y971OhNzMl7Q7oJZ
STdjTzPz7jw+YafbXaazIg==
`protect END_PROTECTED
