`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Lv4qMXx3FwjIfZSOYwEPmc/BBEnaNe6BYjC8WK9Xi/keOQziq/RvwBComyKyA+Oa
FXTHb6mYkYNbk0XqwgLNMDHjZTBG+rAJdbdZVWLsOazzfYLJ6/NMLoC06rjqfmoM
qyqLDtYajxt0CX6xlROsDhKhOfujhbTIdILt4b0qSKE36HVTr70Sdos7/UOjkg6x
inrSFlrG7bSWNtbvTjGdh6WFcaLeyXwqHVgHsAP++k/ArqdzJyeeD00LE3ysxvoC
XqqAYhIic57X29aqq3Yy532uwHY0Csb6vCqmLxJFtWuwEGtQruftFy4CyGTBiioh
O1ZLA115w8U4mwIdSit25Mn00iWzkdjFlXdKLVHq47ns5Vn8IW/glU6dV/+zNG20
q0xpdtfeJ6XOSK6J7SNjo8gQ6Fai2cBxpm9bZcB7Wu//gsGZqFUQGYkm+HeUfN9b
duQ0TFl9TVNX/ZG8oBXsVsXp99yFcRRwzCZw2GXqYOxVtlZvSzOy+5Ghe4An07RQ
xVaFXsS/Tdna4LD04OHYjCeDFNUTXwlagNZERz5XY1g=
`protect END_PROTECTED
