library verilog;
use verilog.vl_types.all;
entity cyclonev_hssi_rx_pld_pcs_interface is
    generic(
        enable_debug_info: string  := "false";
        is_8g_0ppm      : string  := "false";
        pcs_side_block_sel: string  := "eight_g_pcs";
        pld_side_data_source: string  := "pld";
        avmm_group_channel_index: integer := 0;
        use_default_base_address: string  := "true";
        user_base_address: integer := 0
    );
    port(
        emsipenablediocsrrdydly: in     vl_logic_vector(0 downto 0);
        emsiprxspecialin: in     vl_logic_vector(12 downto 0);
        pcs8ga1a2k1k2flag: in     vl_logic_vector(3 downto 0);
        pcs8galignstatus: in     vl_logic_vector(0 downto 0);
        pcs8gbistdone   : in     vl_logic_vector(0 downto 0);
        pcs8gbisterr    : in     vl_logic_vector(0 downto 0);
        pcs8gbyteordflag: in     vl_logic_vector(0 downto 0);
        pcs8gemptyrmf   : in     vl_logic_vector(0 downto 0);
        pcs8gemptyrx    : in     vl_logic_vector(0 downto 0);
        pcs8gfullrmf    : in     vl_logic_vector(0 downto 0);
        pcs8gfullrx     : in     vl_logic_vector(0 downto 0);
        pcs8grlvlt      : in     vl_logic_vector(0 downto 0);
        clockinfrom8gpcs: in     vl_logic_vector(0 downto 0);
        pcs8grxdatavalid: in     vl_logic_vector(3 downto 0);
        datainfrom8gpcs : in     vl_logic_vector(63 downto 0);
        pcs8gsignaldetectout: in     vl_logic_vector(0 downto 0);
        pcs8gwaboundary : in     vl_logic_vector(4 downto 0);
        pld8ga1a2size   : in     vl_logic_vector(0 downto 0);
        pld8gbitlocreven: in     vl_logic_vector(0 downto 0);
        pld8gbitslip    : in     vl_logic_vector(0 downto 0);
        pld8gbytereven  : in     vl_logic_vector(0 downto 0);
        pld8gbytordpld  : in     vl_logic_vector(0 downto 0);
        pld8gcmpfifourstn: in     vl_logic_vector(0 downto 0);
        pld8gencdt      : in     vl_logic_vector(0 downto 0);
        pld8gphfifourstrxn: in     vl_logic_vector(0 downto 0);
        pld8gpldrxclk   : in     vl_logic_vector(0 downto 0);
        pld8gpolinvrx   : in     vl_logic_vector(0 downto 0);
        pld8grdenablermf: in     vl_logic_vector(0 downto 0);
        pld8grdenablerx : in     vl_logic_vector(0 downto 0);
        pld8grxurstpcsn : in     vl_logic_vector(0 downto 0);
        pld8gwrdisablerx: in     vl_logic_vector(0 downto 0);
        pld8gwrenablermf: in     vl_logic_vector(0 downto 0);
        pldrxclkslipin  : in     vl_logic_vector(0 downto 0);
        pldrxpmarstbin  : in     vl_logic_vector(0 downto 0);
        pld8gsyncsmeninput: in     vl_logic_vector(0 downto 0);
        pmarxplllock    : in     vl_logic_vector(0 downto 0);
        rstsel          : in     vl_logic_vector(0 downto 0);
        usrrstsel       : in     vl_logic_vector(0 downto 0);
        emsiprxout      : out    vl_logic_vector(128 downto 0);
        emsiprxspecialout: out    vl_logic_vector(15 downto 0);
        pcs8ga1a2size   : out    vl_logic_vector(0 downto 0);
        pcs8gbitlocreven: out    vl_logic_vector(0 downto 0);
        pcs8gbitslip    : out    vl_logic_vector(0 downto 0);
        pcs8gbytereven  : out    vl_logic_vector(0 downto 0);
        pcs8gbytordpld  : out    vl_logic_vector(0 downto 0);
        pcs8gcmpfifourst: out    vl_logic_vector(0 downto 0);
        pcs8gencdt      : out    vl_logic_vector(0 downto 0);
        pcs8gphfifourstrx: out    vl_logic_vector(0 downto 0);
        pcs8gpldrxclk   : out    vl_logic_vector(0 downto 0);
        pcs8gpolinvrx   : out    vl_logic_vector(0 downto 0);
        pcs8grdenablermf: out    vl_logic_vector(0 downto 0);
        pcs8grdenablerx : out    vl_logic_vector(0 downto 0);
        pcs8grxurstpcs  : out    vl_logic_vector(0 downto 0);
        pcs8gsyncsmenoutput: out    vl_logic_vector(0 downto 0);
        pcs8gwrdisablerx: out    vl_logic_vector(0 downto 0);
        pcs8gwrenablermf: out    vl_logic_vector(0 downto 0);
        pld8ga1a2k1k2flag: out    vl_logic_vector(3 downto 0);
        pld8galignstatus: out    vl_logic_vector(0 downto 0);
        pld8gbistdone   : out    vl_logic_vector(0 downto 0);
        pld8gbisterr    : out    vl_logic_vector(0 downto 0);
        pld8gbyteordflag: out    vl_logic_vector(0 downto 0);
        pld8gemptyrmf   : out    vl_logic_vector(0 downto 0);
        pld8gemptyrx    : out    vl_logic_vector(0 downto 0);
        pld8gfullrmf    : out    vl_logic_vector(0 downto 0);
        pld8gfullrx     : out    vl_logic_vector(0 downto 0);
        pld8grlvlt      : out    vl_logic_vector(0 downto 0);
        pld8grxclkout   : out    vl_logic_vector(0 downto 0);
        pld8grxdatavalid: out    vl_logic_vector(3 downto 0);
        pld8gsignaldetectout: out    vl_logic_vector(0 downto 0);
        pld8gwaboundary : out    vl_logic_vector(4 downto 0);
        pldrxclkslipout : out    vl_logic_vector(0 downto 0);
        dataouttopld    : out    vl_logic_vector(63 downto 0);
        pldrxpmarstbout : out    vl_logic_vector(0 downto 0);
        asynchdatain    : out    vl_logic_vector(0 downto 0);
        reset           : out    vl_logic_vector(0 downto 0);
        avmmaddress     : in     vl_logic_vector(10 downto 0);
        avmmbyteen      : in     vl_logic_vector(1 downto 0);
        avmmrstn        : in     vl_logic_vector(0 downto 0);
        avmmclk         : in     vl_logic_vector(0 downto 0);
        avmmread        : in     vl_logic_vector(0 downto 0);
        avmmwrite       : in     vl_logic_vector(0 downto 0);
        avmmwritedata   : in     vl_logic_vector(15 downto 0);
        avmmreaddata    : out    vl_logic_vector(15 downto 0);
        blockselect     : out    vl_logic_vector(0 downto 0)
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of enable_debug_info : constant is 1;
    attribute mti_svvh_generic_type of is_8g_0ppm : constant is 1;
    attribute mti_svvh_generic_type of pcs_side_block_sel : constant is 1;
    attribute mti_svvh_generic_type of pld_side_data_source : constant is 1;
    attribute mti_svvh_generic_type of avmm_group_channel_index : constant is 1;
    attribute mti_svvh_generic_type of use_default_base_address : constant is 1;
    attribute mti_svvh_generic_type of user_base_address : constant is 1;
end cyclonev_hssi_rx_pld_pcs_interface;
