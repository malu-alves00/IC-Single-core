`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wIcWP+fYnvI6vuibbOFfKuEluNQqMLVvFVJdge4QkfWOWC02GpVB7dElnUOvj4wF
tKljp8pkfnFNN8GLNlPSs9ZLJoA7c7QzQOb0jfu1J19GCexSxGN1QVNyhFH+KbY3
q2z5KVtJ5XFzjorpeEK/oLI4xH4jdY4x8+7EsRplY5WezhWm1Hx1mpppAsa8faXn
YF23inio3A5zK1lo+FZd9nr0Nq5cqFGeyzSuEdAdFoVUmo5svRQBrePup0V8MCH0
2rLL+5Eo+ucS76y6e5eeltESN/mNghNZll6WvFsjdFaJ3bczD2+KAY/hrUoGNzfk
Z00njZKbGYywApuGpLxynp7VtUo7h70p390Y6Kj1vtvdZvtue/LZtGmkT1ckiprw
MS56Or57l0/wq+1A7RE3+uOZD4exPcOtB8Irxmb2h1NVO0CAjr7BbJnm1/Nr14mc
AVgDh5pYstyjVzGbSuxiPor+mRB+o2AVGCqoQEyS89EwlPaznEhT7dq7f/hP88vB
Ub1FooLAWO54Lr3iBOgBD6sFAk7BlAM6gGsy//KhXMM3DwGL4yEdIRfX18tYBN9U
OI8S6vQtspGq9dJ2401d+SnK7upSA34CSQQBhKxDXEIaHyFeJ0c2kWfRQkA6SP8P
KXpZbScN8mLQ/SoHQsemvYIrRUU5VX1p08lzTqm2JY+Qu/ecPlxQBweJRxXdoFdt
er1kFRjWE+/jwhUzeTLPuZFIln9qnczRuXC+qGLy3BnU0P/8T1WPj7wID+fdWWiU
DlK+H115khuvOYhwzrWzslyVwoO/TU9Iply4G/TgPHpHq3zu9Di5pNw7/tbTRtXw
hsWzNmcTkRpbNelHqoLgrXj286IXTPP7B1Qv0HUcFrD50uMUQnJj59bxmULwN2jN
JRnp+Kki4OQh4+IhF9VLD0WuMSRdpgEnlZXpLeixMxT5ryOThHe8NliCEjaQ8Lqw
NOqmBBQuBIe9/L74vob1szGguSWZPiKi1iN00xb5IJomWGinH6Ilcv9Ac6V8w/xz
aSBcufmzq8P9lQvplB6Mda7E72r7Gljua4IK20WSzbNx06ce+PRApYy2D0w4/9Wx
wJmshQcYKApWO+4Ylb3Ci6pQinxTc675CmOg6zVDwrs1IEFIt/cl9dF7lvgxs7wz
wSlg9Q5Lx7CpRd0oLAEs65tJVzg1inkXrajlghe0zSj7DHvdJQXicZC7KIOuZ7xw
TQjhO9f7Ntu4ejxttRXw52z0+ahzfqnoNyl7oAFOfGa0er5a+7zR64GTX5xKfs8i
Bait+YEh/aSWpxFDdj+wC1UlAG7kPKnFvgzHcD0BezjBMprgc2UT9wZsdH6UzfKH
YsMiazScy3P18ZEf16SK8s4or2CQ8Dq1QztdKTbggrJW5fDH2Xox3cpO6itseTkB
VZ5jnh6YgW60uz8HWZ+7pTuUaUngYie6uEmiMiKB/Q4i/auxaW+ANtNVgO8oEamf
YYBCadLkmHu6dI0v9zXZkCC9RmUaLmsvvaNtGLjSKgWkFKpWVbih5S3dWv97d5aB
mmybV8ADk1MxnzvF8gJzZZ0TBKX6+ZPiPZEgANaQEn56yd6dKVQFCMjso0YzRz/l
id9lVnQUhhhXNB9NOZwQC8UNB4CcbBjMLPnxXPir4EwzSNRdOfq+A5GotcZH7yxb
pse6cMvNSIu0RzckSV0qgPnqfHbCNIM3wMkMKFprefviiD8p9VEAHyrmAIpr52Ri
BJo2HDwFRelSsXSaeDTrZZYREYgIzZpyDLhHGmlz+R5U+QIWYMmCIO1zxKzl3vrj
f/HQlxsCSwKGBTGdwLUGQJlupv7ozKoJEv/AX7mEHywg4p0PIHBTzIBzwsOzqF47
gRgMgZSkAOpqZxylB9AomgeX2TBuUth4FEGaJAeidjT/R13IPQNn3BTZvRUoIGFz
ewfPuQQ79HhYqVVq1nyK2OUrdasrhKvs+4YINC+qgda8oirYah6XHP7RI6JttePC
y+kvcZcQsn8rNkaCtqzRSbGmmi265bj9LtAXXs5p8PPToUT5aAc+aGQCDiLsRUif
lDrWyQnFFFEuw/xYVrdsA9AZ31sTU+n0PkWivJZgjZaQNti3KWNWOw1Joa1VWSpc
Or7qu5g/lsrvSGMa8J+lPGqpefkja67N7hHKnKx2FNe5KvoMSrCDhjh4Zih/O1Hc
kLlW0+nOe+7DFSRDYJfX+t9dEtPeL4wxb2geFx8P4LhJvumE97AHbIuRUzI/jjrU
QyhrKgIlM9Qt5OMDrV7A6zEW8b1+gc9HEONJ1SFNHAE21dm6qiBgJDFBzQoIaiYv
f4zP7cwUwrm5JeP4NinodTqDBFJS8bUmsK9ZQpiihb/Cqh7YCgZN34wtclpmTCGE
VAcJj2MtKzCT62lQS1/TigiMqRxllMsmgK6wejgoHlrNCiFuaKG57U8BGJRsx49H
36DTWny1tSiWyMwslOsokg==
`protect END_PROTECTED
