`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JeHMrpW17nEiJWnULCWdDrJY2LgInH9P6GvIcPiTR7/Xo+MBO1BeB5PwSr9QAp17
9jhf8/JR5rhx8uUOFmXeWyPW0iikySfU7Vp7jjeIAePld7CpiE2vB/h+mopwAHIy
1JTcxz+1uos/ZadtKRCPo3mJ1GEeY29mR30gsM6Go95HLlilduGNikVjK7pFiiJD
+zZC/RJwQlWwPqx+kNDA9Gg3TpIQ8Qu0kMsjjRXTZcEFPJqO/b6vV+ZldlGwjuR6
hq7ASXvizUhtS9btGkhPO0zR3oc60BAqhuMcWpU6hc3qXhmLbO/xevunOmx0DvIt
tIDX/YTR73x+YLgHuk3Ckb/yA728wzZxmqdN12536sviEkF37bAuKes1FIg5SKSm
6USXsrBQQ5xnGMMV6Fo8keLZiblN+F0Q4s3vBXkdGZsRLCgz0nAqdFNcxFVc3D4M
+APG18uDsTSXNNI99xnPI4hiJzadcXJeJjyMmWuAe/speZkRkgVo6z/LlKH2Ayiy
TKbQ2jNPz+6YtWqnhdoLNyjzplXH5Vb7Sh3JOhZXfRDx/H8Rr5d4OAlXGeyh13/G
4R7BvYBalmiKjmwn8fPoiz0Ut36RWNDSPpHiCW1pz20wWAmMQ7oE0osQ4tdZeoDJ
BxdedqHCv8UI2KR7vk3zSGCrpm50/NmV60HZUSeByQIhxEFdfLsiuPWZel7Y+l7j
WDkNT3usThITswLwTCoefUyF8pySltYlzLUsIdjOvFn2oUFRKUjhpCmBlKZAkm8n
IzdZ6Tr2+rzNgUiDM5R2om5FHEVyn898k9s8+G+GYf2FwmcBBSnqNIFzFj6Zl/l2
fZjUbAFktHmgQ5oHlOJUxvoOs/i6zSHhXGgrfY0wHOQSbIINQjCxjpA1UZj/KDev
I+0GhJBCquka3hjf+NTbaAzBb9naXsppr8pJ+DsYw3+vh2ZoGb7MoPQ7x3iCU0Wt
VHQmJfXKX1R9y3Ee88IeqDp34Ci8FBxa0Y4wy2vrikYkG3JHQQuI0Ty020DJ/DE7
xLhqj5oPhVzV7F/oYis+AFNUiv34FKanAjuCUgCNGZ4U0I4iKMfJRZb0GXv1ZIe6
pRq3c6VIucS7I/ZuWRYzlJMZeo2/1FGpudyXcHXE3v2Nu9UY6uaOiD79FYiaei1U
RMGRJ58PNpUDAISF/oWk3IpEje/NaLPhNdgMNU5EGpJ0AMHhuUtWnYSehKLVtEz0
NMB9LbcTIqE/aFEs0tFlmZpyWGC+Awlw2jznxY7UoXyaOmigYiPY659qZtPrHQCD
g03DeCwIOfutRhR/22fnGLN5kYcq29SNmUdRrZ12mB3Db61jK3asT7WTmms+zSvB
0w6ZgL8aKVW2Chj7/BnpQtfTPCB8jxFaLWfqPUy5sW2G7xfMhdv9H+TipzKWkrRR
k+kNjz6dUstn4CdlR2/8Tw2K3GjrWE/jcVvzu+Zutv52LTo9OszSulG1eFBUHjTd
eV8oQAs4Nbqfa41cS5mvzyXdp3zD/07F792tbSLUJ+qC9jtyAh+HqcEvrXZPwvNy
wes9+lSywE8OFECi2dO79GyfeL3p1P6IGjGT6RmFRChKIolgg9oal8aWvwmkk/Ll
2Ysu3GFiOvBvkhOxfmtoX4bKDmRCeRaQQCuQP82YEjSODjdQEZdEbqOJpafOCCCE
UElIjMTOVoZuyQcZH7gcnpt3Okkvc+LUDDUSmNKQ4dLsKpsNKrbqQpWfv/+8nvn8
N7Kd3Vv6zdOBdE9ArO97IjfmdgyKfQKYIJqn+rEGCwggSeNEtLuC75nS3YQlrfou
wRyIk9i7+CUlRYFWPZSk97l0E0Z1qplypxGNIxI9TiezW7hEqkaeoLBt2E67nrZv
PWemxQB/PtKrrTHk5+q6bX+E2tpu9FTg6h9gpK39kK3OmHL69nf7d5RSWKX/vdOM
A5KZlyXkJ1xlAbdx6no2BOxSILj3Q2PU6TRVkseiUvLT1mhOcI1RKzUESms2DC+3
PKtOJuitxe19kQ9uYBTbxVMn2zaurMkfZMRQf3aBe7Reweie0B4fxjp81M9FjJdm
zLpPQoQ2ZoYPge+Lq8fCFbPMmqcUtIkVhARcjqvLoqZOIX7Ucs4IO0/pA34uQ3Bp
wzRg+awrw0Mw/9nD+ngbVz+u9X9NC3MTKGz7HH4zReVLea2P7YOTiV2yI+IMNCvD
t4yllH1MpX5wb6USEvHARrKrgW+0AOiQ8DfsIYet3Xd9pgxjtmvSWyYof7gVeWxE
i1iXBeVglnX8xXcglkh4tft9VHkG6QZltv/Q5viyMR+oIBQm/Z9iFGCuLcM5AvH7
4sY9fl/6JIhz2FTygYJWKU2p9pBvgYYlj90MyuANIsOq2XYzrNsD9GqEW1O2q7rt
bMdnMgMXlJ3DyVWscZzjtAUAkPEO2dn5rB+MeiYIGdJiHba7sTeVKNl4P6mevBK0
OB4X9z9L2dkb/kN5gpCN0d5r/PQIG30qOARgEKpuJvEav+yOq3KkmbvWL1vPqcu/
Sl2+mo0X8Jy3qjSmOx8YvXaJwPdKrpWB0xu47V10nQJZk0hqkNc7hvbFTT8WULXr
jpMaHY3I4L5FygsCpK7B+VW/9SZGqjXyH3QWgmOxIu8XYHKJH/vmRgJPgMMSAvvh
dJ66lQHGoUOh2qyWZcsnFlYCVmkyJisPa9uVeHnNCIorjCOFG7yXxByKIxZIc++C
mooQDKYk3YAwr7AbBg+hynuSyPNF8DZh6Y3qP4ENOfrciuESN+vNe9Q6go1E+5co
Tq/HPNaGOrRz6HC1UfvcDmpikrpDpuprVAyS/WFeT7kA30TunADd1rU67hg3CmBg
3QU8xeenIEBZT/CjuWVO56DyggTljjDuJNvej0C9oRS7f0alJWlm4vQzhkKrM56K
eXuVmUjqsJ+KAZ75PQxxSYaEj09KXP4QvhS71iTfXCOJ51OD6hGBs74XXSyyGcVK
vAdJF2PGZlphbaTO9CCgyEUpC6h4hFwMaHgLva/ssM9oUnH7Bh88FqWtBRzDKhkF
`protect END_PROTECTED
