`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Da89t8JwerHj6a2+e8tasTCC1XvWCUr3q5y5nuP9i1owwnmLUFxA7J0My7r9FXZJ
DsnR37aIB940fYWQ8ZBnLF5d0hf/bqwpgyTlXT8svbVsOz3AvRHH79v54yX+K63o
CQan2CNSfZHik2rfEMK25AnB0SyUONcUSmUiq2o0CIL8ymzjNBWpWlGqiwrnVxes
J5gyIHn/VYBYDrZM+itxMSoNvtVVZYAYTAE8XwnsdoNOHbDl/TCBN+o5Ai6iPYUq
Hz2beP7uErlc2I2rZDj24V1zZBqxeN1/LHLBJF2LoMM1eWlSLpNxG6JtoS9i1lTX
zSBbl52VPmvplGzX5PC++koni2V16qsBZvFEfRoZSlBSQLQSe7XaPpOKYFQAETyM
MWJm//T9WdBzqmN0yhx6FUkniOpPaU01BlBKmHE5DAB8TJ/5sA3s85SlUYqc94f9
FXcxsXPHVYlaPiumxwZLFsyDvUotZlEd1O8hLHf52k0PpbjWhxPG49CnItOccH04
gUUIaPbjTr2eZyqUF7YuV/AULl16ChCFGDoQ8VlZm88ECThMNKGMVyRDbUbVGBba
WdEfOLniT5OyAxkNQS2I1XxyHJQyug443S/r9EbsVAHdXqi5E6gVsILvxmLylZe5
Ys68DoX4ocIipuuwiu4vFXpvNoGuIbIvSdBZ0sQC0w/+W/D5Qh82j3J+N3avnvjU
DWu7lAtue3bNaFVGLNl8pABI/tR+qJ4Fvyq27OURnyoMHA3Uc3lwRI7sYTiEUiwc
ZDNAuZoEFfeELDe77DZEqhM5bXnf3+ES4RSINN9Wg2v0QpCATX8F4nDxzYa49pPp
xQO8HcvoPCe/cRC7XiTFyGb1rO6VgJLN1mdGZ7IXFTFSr2woZINfcXLVLk2cjcP9
g4yusE0xzQ85mPa+TZUFGAdnYW1C48JJVZDqcETXY2CLxPWVE+q/Zn6S3NUNTnCl
N8uw9NYzWpb1ZYT8hKXSl8EI1q/CbiYl9Anu3ImytRg23J6LlauSIYsc66g5fC5m
SwK7iLXJjK8+BTqj843CishmMxwj+UPrh2ciW/7NEz+hWO7XrcPl7v23Fs/ujOjo
pMcG5Bbbb/sceIl63l8CZFBGaXm4RqVhMEOA+mV8x5X5pfkRhpQwyI1rhP4es1L5
GBP+IwaC5Lh6pIwupm18KKN7zf9vZ6rDdPwZjUOg6ampGJL5cSwxobgxvHT6PyIO
SnAhr3sL7bPd6L2fQuWb5ttHhpM9dZtzQGopx/6iG/ItrH5FhHvFxTRZR9E/W3A1
gD/HeY8/mcQgPeAxUXu48DMo7wruoyLcmlbUhP/j3lePkjJfV2HxpGaNb8237oxd
I31Ijbq1YJfXxocgtb3NlO3/9JVO+vu1DbtzvWzO8UFvJuzB8OYeGzTUOc1VH6RP
auDrOLEU9K6dV9CL3iy5zwMkPjtWaK+/mLKZq53UrtO1eFC0AxAVezFKG39yNXEW
r3/Nrk+ODuX6gmoQ8N25yRhuGrkqfYSz1SsHCx01npU8WEx9f+g8+RL7EIRunAc3
UQJsQepqO01z13GME6P2JgaITnBAURIwRtXbQjPLTYppXe9NS9/hyXSnAiPyHE7a
BJupvwgYSmC2j8lLpkaen3mpbNZYr/PR1krWAa3qm2vjsTMDJcblFP0c5gV6b04T
jFOSkOCmbQyaRaTWbgUSrkistgcw/H9HTrl4yKpji8AqR8PTdgunjMphh77O+8xI
xLixG67Gsyn9Odtsy9SAEWYufS+52hUH70yEJ2o/Xoy/TRLo8fRMK7d91YIahjQ1
mMA5zZ0+JyX0sITHM3+Oh4W/FhqNHgatw7dUxFJPeG2L6m/I/wdMhOGjqxvM692d
cU9sGkXPgDb4toPV3j20wXNoAa26Uw+3UCzW7QxqqdinBSYURUILrAt5vh5iG+qW
zhMk6kCTKuwqwrtQ1KHeZQwFHZPSGzSYVPyoUICNw+vuHPH0r+V/SWspvyu8c/va
iEr5/KHFHluVYYYWYJ+YOMciLEtBMHuXI9bULfgv06xM5+HjEf2UKJSaT0fdScno
4n1JxM7R8+d8DjWha65CKkJ4g6EQtqV8wGFTfBgHddHWnCBI1Y51wOn8atwDDEMp
txa6W9Ky4B7X5tV4dyHWRqRQGQIJJ5hnqHXjS86zpd5+8dgd9Duf56G1iO9M4ZPm
hEJ8/f2/M+ADT+ObIFTJdVqZWL4keTTrKJ5B644i1NYVio2y6OyZkm6T9LPGxOG8
12y7JsvnC28pE+nefz3sz+JTakr6tZz6krJqAAKq8mlTh3kpe/NYCsI1BV5K+uZk
/+f3jEFDu0QvuMMuDshLZ55fB2DuVdaHzo73Cfc9eyQAZsL+j0HSQv6U5auEzh3/
wSjfKuCr2d4ZnHvNs4Ok/MPjXmiuNj8jlnjB1hdtBJ5UHg6GtJzqKhGXjb4Yo4nP
9p7Z0t2kN68garYxbbfR8vLiP9WgmBiTdzcTiirqI4GiD2ZZyxOL+F1kF1al8Rfx
ANr/zS2nSEogpS03hNqKAUONYAnAsVfApLF7oAxpZhmiC46/8l1wHAHgcwiUU/F0
sms51XQ8d8IHvpSd/jRqefB1NtSSl9nDZdYL46xfWaNE1diAx4lg4fOPAmqA4upX
AHh+YTibu3jI7rkX7u8BZ9rkccC4w9HorTm0EFFVXgZlR7wrmarhf6Ng5hdMM2RL
sZCi4mnQsCLNs9jKZPefKuxsg8dXeXZAsW0/I/ZZsWzKyq+5acEIazJoPcR5kkqD
Y9PjU8lvrh0Y+IoqGP4kdpdvpAskHQYKLYRo3b9gF7Og2a1BFmcdKKmdWznwNndq
K5KlgM4G96wMyNI1X+VL/HQOQcnceZjck/xahnVueUj4tbdFJbDbKuWJANgKtFme
r+6GZP92KjiY+N72WrrXP3iHZrrRdV5QWD2CaZFpX5ghTbto43RjUWpsz+U+sazD
AoWKKSyUGtkZOv7a66RKfIkTphi6lbwlg7TfVm5EwKQEkvAmQ6c3D7OH0GO2VsUb
/v+WawgCAQuRonuwl6P68k+CMFnm6W2ULb/XjowHVg47Q9y9frRErdRIQv4eo3Ct
1dazbyoKGFnSyaaMJA5MQDzihWLTZe18ppnWQQgzAmOFDn655b1ErK4lDtm4hh4d
xW0YXyFzzIsUFezDT73ndLR86F7MWQsCLXxKX3j8otCb6majjn2+Bl6kCQkVkL9g
XtzXM0vnYGGocHm194S8EdCwXHlase3KAi8QA4rB5qdI+2GxlbCQG36GsT7CZcl5
VEKgwS+UMVrE0bHj68xJecLPUuPD18tVKzPY2mvEpxFJHb5ZSVD6YXEmNnzgEJP3
YXtCa076uhgrKntOuISc/rpllzCvd+uvGG5ldhWpkRVA50kwULX0yBYOtytzTwaj
9YSqOy0V0W3bGnkU+fmUrdqEFhw4ytUtpxHH2xyIXC+gwgkrCnP4EmNrDtBszkl3
oTU3IB6gp9+tLxcH5p7DJ+v2Wi17KfBsiLftLB8hPawwWSqzWgmGVZ84VMm5/2J8
5J0Shn9DIri+QUzh4I9zviYblG5q98KIOJ8+yey2IouPkILe6pr+YPPIz0/AgRnh
Ehz9TsDhT1jN7Pt3X7Jsns9byg59YikuAoZMtuedcuNWWgg1plq4yfIXheMTksjZ
7SjvRIIQIRMWt83Csd+cUS6EGQ6RQ93FOuByn2Oj7vpE6PdYOPPaw4+qlFWQ1FJd
p9489IR2+eaBISOeGtliw65flkwaiqP2GU+ajLVjBBPNACuwP7GCeSAp5H8RnEK8
LR48cTP1YuhLbVvK2to7OZLZSPsG7QLGy6/ualT8xv6RREjQnOXl3fEFFp/qJhyV
DRb6jlRUMmqESMVesitbDfD+qRwVtfTa7OwsSgEX4DO511miPQfmUtLvbHTolw4a
vSqXjcIJbjpHCPlHa0Uv76F5lj79ZaVDUidK/XdSxzfTWcRABaOXtWRd8EOBtsvi
+EWeljgZbOW9vHOZKS96M46+gGMKvL0n2de4hfwzlns9Olm+UQhXjyoWzQK5961v
ohFEmywfyQxATBKAk4yuVzE9OFQ10J2e7B0qaJUm+wbnF9tbGyX/MTDcdctnCdni
cXL2L9XsF13ZDBJh9Y+3sh/Cw8Uy/js1pbs0Ct3WCAd5je7QRsgXowTWniq0cRFi
HKsV6QCUQj1ms+i8icY/u1c88hmdBW/cRKeSIGQued9fM8P5x6F2aoDARyRSTnsw
maGvCNg336AHzO4GAM+xmJUikg+KwJu1C5PDG3VWHUDCzRNH24Dew9sM0cBYICFO
0jbUSprkDVW3t4MWiRHpKmQHvRDs9Uojh9ZVHreOJumW+EJBniENgBNlic1OkxEN
VwfVF260/I50sAJYv8ZYqH/ugBJCK8a3IhTU8lrjS3f3F9pdkPq1C6BCnmo1pLaI
F0rZ/RgZ6n3GOTzTVBDJY73RX1Rhw26gTStKeH+HfvRDXVjqr2DpQ+dXZ10NzFoh
DClwE/Wn7B4rJpwf8A+upecUn/5/v6I9271ZMTDqw3Q5t9XLtRqM6bqXa2nPFB2d
qVOtDyGasnO4uEPsnPCXpceKH/Pju8skv4JCJxB9gc9CbzSIyHQoa/svP9v/XTDj
LCFcVFh7LbbcDmjNtTytv+72dyxy5MPDg41pJI7d/H/BgBlm/tIEuPNUcDTcUu9O
lTapPFB6rQ7p1xToXjw0/Sqol5bpLqJrh1rvDsNcAxuqsyKT27JuRILujOIkR9Yh
rDLCXjOjAtg4Q1tVCZ1xJsqZqhPhkuoGe5a/ItXtiADKT8fdjCwyn+lKy4a/2QS3
pQhg64WHejRc5kfjszSAp+udSsNYtZlGFrpQmrAwYFXJxhqWx5nXv2MOQWw/G0cq
9Ox4dmY5Mqbcm8/698f7jmcqlNKyciasw3aICxfBz6COZtQdvyrSLWpNS9zOhwJS
RQbwDUlqDJZTKa0KWlxCv66HiAivTtduf5qECsgnOa2E+BcP7XEXxyso/Jr7ZTuJ
yyD4KhwdkXkNde84UpHPueoOM0lCzsDNgmZ8Odfx5/8vdHcsCWCj9aFzAfN+IP5K
xuW6LWGz4TcSa8c2cgSSVW09WyQKRXPXk+AKTxoiQLtUw4IKvkCIriRIaI/AxSmw
t46dAiP43VO3YW1LDCDNQhQ7YlzRsLo/PlluaBHZXnqDZGBzaR3mih4IIc/QKuKH
7gW6nFo6pcZUYpUlbGw/peeGi6YQdokahBR9ySNUpN5rp+p64A429pmVcRgwhB7z
ZPOoRTGDJC8xy98IoUXY7fDAHxcwZ4e1wvLU6g/nyEMiDXmvGX6XAX/FVlZs6Bem
hvSwzX0yJ8UoQwUVd3fwmqj0Y159d1qb6S8Rz766bRThi/59BZl5CN6Ifq2WBGIL
s4EbDWgBGgZH+uS865KK5PbmeAnElF90t0EDfmZiHBQqJgbxj0QhwO1MAEnA+BW2
7tR4bK9OKgI4Hm3PFn7OtBAdIFqLBasAa2nxVazU5K1YJt48+z/edLY+Y1xY3G5W
/xhEFsLlzT6F9C9F41WiP9bfIE3ikfPn1aHDjwNj+w/62VDBforSUpSeCM7L8xn2
vTgT+wEHxMcP4HCT/iYUCEFla1leTQ7OB1E+MxIb6pr7NQFxYAlK2quNpKJxlJXm
DB8UgSGI6ZvbfU/HFQstFnZDUUafymj9ck7z8KCV3rGx1c1moRXxwVQK4zkpnrBa
VjXeh3VlC/HNLYYRkh2yWCduIgHqCvl+FLNGQhF7ZSyjYmLp/vKjxsmesct9W13t
6sA0U1he8wYlGVwR6W+1dzlNUUPZHcbnDXzvcrKaXrrbcbbthstrmvXOroyzH+Zd
GTX1xme+4fpsdMJ9VuqyNsKHCFG+hU2t4NzzQX/6smdomcFJId7D5k44+ow2OYhf
GIIS96IyrwcrrA4TItqHzJVT4+0w009gHV19nhEM4bJXdo4OICvv2L6pLT4ileJg
ngOesyJbOE2atH98rFtcKpQQZLB9A7pjRCSeRfPmMtljf4kf6JxDk3egk50EsIgI
54XOdZyeGafYIK1zqjoZnLNxsFdTNMQWXXaVWM4Btfl426LM252SdGA9JNf7jx1T
UvxvDBB2CTxz2pRGK1hWVfvvXwAj6MO6cuyGh2uY7m6MqbQGi6UVeNv/bUT11+sj
1dCXBjbLVsCRPbaKNer0HhfJ2oriOWuBYtTJYoLQjk5GTakO0Malj2DkE3Ch+NM2
TPJaCZQP4LlvnfWq4wLgq4zYp/MObb+h5N9XOI2r5PSHRy6XcFR7XiRpHji+CJjs
l4OOICTYn6kBIk2Du5r4YR4dn+Rj7WYcb7gJMDZY5Pr3d4ufXdixfCbewLTz5yfH
K7F3dhf94IyTpVi2vAbi1SUzXLTb+gRjc7EVSHO/Euay/SHQ43GiM4yFeRaU16Xi
dEAgZJJjnnCuF4ap935/emhE4F/fZ44dlZiQQZa2unEDb5d1W419/dJ5G9jL/0GS
oX6dmplSmthTT4PvwbVjdWdiLJ6gUotDt5antih8eluez2+HeK10DISnbpXWSBIo
H7rK3SR+sg4nX64aUnY1xFZ53JQGSQnzYYawsiZfTlCOM2XjU5cheA/8idtEK9A6
+1NMH2ikeDywhgITLHD1txim2tKqOjhJFUMdFGuw5c3SaKUn85LJqBqhNehY5jVu
ThJ9LgofG2LXhQqwiryBroz9y54zB1K7quFB8jgwASTFPubVsPEBv6f6gl4ZOooz
frTCJAFtC2kS7he6gMOiX9Wwi2s0/tUb2aimKH2Vnnm1Dia8QH9np/ltgfe0Sk4n
Mcu3i9W34MsAEMjqqku2SWHoa2CjfFuPDMy3qTg7fC9b0nUulgJj4uu6/sHndiqK
sqF3Y01AvcrMkoJqNroVcF0se8KjMnzUebv204CMA+TutmLpq9+kupV7IWoTNcFn
cBDBBJ5PfXh+rQgzsOCtOF5E40L6/eB7cgNhj5+tU0xEb0bfNFcFmftEnwj0rFbo
a9s/5DzJXNzUcILPm8NU//8IhbED0WMQ35zZbSYJc7Yi7EjVJro51Pd+rV54RBku
QA13veTpXX/DXMvXsDxDkKDAhpaX/jAcQrzqhgFMPYzyNl61tcSR7xG88pjqDuwh
hvqSTnscKAs/0dXrw/nGORXygThiOmHPJkRxPOInTefR169HCzbdCzU6TDdakNl4
heiOrve0sXM+neIh0Rr6jdqrmMGPdo/z1kDbfO5GHous3A8bzxIRZMu50Xx+4F7R
6gstZwMdU2zFmEWMPwsO2T//nstgo8amUrjAnvApmeGogpHqGDHqZ4i1fd7sc6l8
gsN8SFithhmBWl67mTXKxHQ3o9ue/jEHY1Gsbi/wwm84GWvamNH4CjJDzpR8wsLw
5N1ImIpZ/us8uEPkSXcOIAobZAqxrYjK/yxWOTmChAPPU+hX8qQp/474LMunIT67
0V0gUFrMERMfUDcd647LDryzDO9J8looquZFl9ojow7syJhzRDxE1ERWiMkpASQn
rmfw3hOZJPT5IJU/0Ho7wzmdQ2HRjxZF0++zJ9/l1dM+chfexuznmtgJ5GUWVUdz
VSUEwu3Mc55qF/zS5WX9xRqkro5tSQo7e8c3cVj6ROG2fOh1PPq7Op+6xAjycd1V
TtmalZRm6YbEEMDzeoGgQC0qH7KYDynpUpZrSH89gGIC6GMCfpukEJevSeJPkM7S
wNppZTyMdfdmIr7IPj53uvVmB4WMPRN7SaS9jKOjBzP59PBG6h67ubxFfDndQdKv
UdZpCySzaVCWSgDN+okwYdVUPEnaGcmULRmAYEsTkZN1vnAnxfpCC5fGyoLQzYWK
Eu6eJnOHrFJe0ylWqplApyZiq3jmqw4sNpbHMTsUJM2BetpVfMXtIUzSM/I3/lb1
6hOX9isrVEehA6vkpjpaJtXMSFSgCIZg2Kh6hZvz8an3e9h0Q8MnvHe9q8EZlMmQ
tOJ8SVp+koYmoa0XNGWzQEvRSoYesPU3zYFoLqoyfKDt7fnydc3zvz9gOC3gynst
OVTHNDd2WdjDzoHjvEfcAWOX4Kv74hLi4T4L79Cmxwz1S7aJ77RiW2gQgM3iJegZ
CNzriTy3BV04ElevL10gLeTDp4biiV8tG5wP+DI2Z1wTXT5QOe7JWG5gzE9nRi5/
tHanoYh0t6vJM+R3dagV5U5NM//t0WEjCnRQOqyfHSdh48U1oumirxHAaEM4BURE
69EiOtRMbVEV/rDD0MKa8sr4Rv7/NcRXDf7tqXgglttmz0K7Cu2NeSjfZBXzrttJ
/8ZKVQPunHrHk+UT7/I+UTSh3vZ8HMPypRxVeRvwvZywgQzCo8cjt108wH1m4iDN
EAD81YCl+peCj9fMxSBiwdS3xaHjQISv/32xA+23QiBcLcqhuadytWR8WkmN85DL
Wlb1OK8D7Yedspyu+9xwJK22Zam2xeko05NsH4wS8hadmA0Cb+Ejfy3U1bfUPevm
KazLlbrmOBbLi8OWCjL6FNNyv6NZCg9yTl4wV8I6ap+AeEmW1UgkZXqLBPL0eaax
B0Zj/OlfAc1fmGWRrNVhFdL3NJ6TkG6DpcRp4hJ5Gki5SMEmG8geoWzp1/wYfn4f
fIKZ/yXJaZxicgoFC0BZSsQfuWp2zsPA8DGWmXpW84RJEDOrw4suE/7FRua6acGg
t4h5lL6nlJtITVbf+B9fhWeTTVAs1zqvJaNI7uL1r9ljE8w1+SOssK1FzQBIwDAz
lEKge2q9HDmbpwHEljxofF/Fx0nC+uCzyX7bX/NN8U2d7SMvvg8tK3WBbYbqveMD
M1TjY/xBxOLN12l1H8DAdkbx0skadcc2FcMYNC3gc0pCozCPUizeiL7BSCMIj2uc
0MwaW85FRqvzya2I53Ygjuro0ulPZQkylT45Yu8gdoKq7KXYOwzgJ+OxvyQayKQJ
9Z0a0uG3eB97GdWdX4JFiViWPTHpEmAZl59jACgr03SEhV+oFWmXC/xjnXknk7LZ
ZxUjZYxrmOA2/gLPFvMnq4ZVRiqJcyY84hHr4GzLmjvlzqbNfCiduyraM0m0lQMR
ngfxq42/ac62Wq4s7Wfyqq+S6Z4O+JFoae3+sidUq27MgCLwGGCThsAAlM9Yk5Ez
Fb8NfhfjHo6oUGP/RoFQM+2mcOtSCkvmyhwUB5AYM5zzJxTEWWktq7xR2xRMo+Pr
oL/GsM0KqvP/hnBs2nhj5T6tuV5N+qDS+Pe3e72qL6XmIrNBMSEwtTTZ/eEZjBpc
8F1vJMUGLj2TNsDjrOPDFTau2n7ckGoeXXdPWTHVtnqQjptyv9R+Txwq2M3Qy2yn
fr4lD3TnSUSiD9obcfO6tc2hsxzrgcQJFxAiN0NXEjQSgQpuzc93j5HnQqhKOYZV
Kq/LMXrqh4Gk8jwAlEWre68LY/2nrpYU09Y6YnOSF8UXh7t1tJJnJoXg9TH5XLmX
jOaS7X9sfX1AnY3S6BxaK0DChLn5eNgFVkmk44ivNMAzaVOKU4oQdmfX6JiClvC5
+dPh6/KDGSWAYRZTfgETNrEQ4gQoOPci9T+r7vNVJ2kRtvD8rBrecknAmSkHI0PQ
+rMogcjokurf59D0um23SsmoDBodkKZdWlp6/PsLI40NoppkhwGXQX8kF1V8pY0L
FD0jrzRxdT0JaXCUzCKF90yhdhZbE0alzLwROPaym5x+/tLc02xduhAm8+b/BA/a
1rm38STOM7sB3saZXTd4/+XAKcMqXFipLMrra0WYPR7ouudb829OiQE2nbgr1Z50
iaTJi31fcHnh+3tdTmmKcUAKvQpHJkMYuA2xMfYYRrirz4nokV4p6e92exE3TWYe
sxCCAVKz5YZkgLZeYFW2u098koFeuS8AEGkbT91OFB6rjepWnydup0qu5bqwnx7c
eW9R3qmGpM8CuPez8ADiNnixToc7bK6ZGG3jStaGc8QaWkaivRCFl6ytAX2Vw4c9
A/T6ChVZMtsti8ZTNj+ok8yTH/L0NW4LxvAKv3FEh1KmIwHpCnwOkL2CuybTmlFu
fqXU1Q4TAeUa03b58DRPfU7KPe499fKpd7KatsPf8M6T9+QDueY8BNSas3ymkqxg
TUQbxmEwLgqSDuRxHDRk/gRblapWdEw3LdNNTbjt+24/86zI7SvHIgt0o78sTuEc
Z7ORQySAa9GUXeJTeE+lOVLtpLZvzxnuqb88SxXVLciq5avS89XIH2BdDEX+xrZo
Iw0km0bbQGOFNMO9KsDLtQBv2ultz5YAI2tuh31QeShfexuOBLLrygDX+JFlV0Ks
WFZEIMYh4Tr38MgrFgEPZzhuSGSDNOgkZdAxJ3qiLHd+l5DNfe8/ec/yH4pOLlA3
ZYw7oSsZnqktIkJ9/LkT+8YZutdHB67A5zCD5iRWWt2dAvsFt9Zx3JAiDhaNVu2A
ydUywM8ySI+27QccAr+Lg9uj27a4afaie6fjXDVq+a5jUl5dX7+EVcLwkkudj08t
RmYSTDjKb6cF6+WEsZJR1gWx5NqJ9ehFxn/gCrnS4hm82o2Y6zaX5ruieEOD67W3
ECKYHShhi2FURHC2af4ZAnu+i/x0fuvpTlJLG1o1nqwtDAR5horT0HTrABYui5sH
bKL63oqrZafHa5rJafhdT8xdAWVQaHCkbBexCQvQ5YS8A6IH2HszD/WcAV1wxiOO
yvO3zwPwUPafbp20I001xwQUCfvmZdxRAdYONcuSPQp945k6rXAUbRzOSX1C3Bu4
couCfbFlp4fi60U5BxeMfXdrqwksC7R3S6QF3V7H4j4/q8qoeisaP8NjxxVPrb1O
l0dd1olCPe6kZq+mNOwwRgablhI4XnHSpCxOBVqV71cyKNa/pgzIx0FxLnPCPLlE
YwzuoBiu16BtV9hqAWiq8u/kZSxdVsLXKSPm3nI4iostIeHNV6NhqV+GdpN/m2GG
FIcfckgFS8U7fzZvFI714HA66VJuYKo89Natmuo+45zwageQE+5ttWpvsZiNmxVq
0iI2oUbzw7hdhUGk1rgcc5k2e1+r2djNHUEScoN5MnjnvYO6gcnIbxse43Q7PsFS
5Nz+1bB3/hbQmgf5PLzA6Sp/E1/ywBqtC/aJRjxrPFXOeOEQXbx3paUaa8egvLS6
92CkJlN9b6OEfoc6K404n6dAlD7YA+kE+p7frfn6+VKg+qANhb20kimPGldBAH7e
BEkgRoWUC6mPSpz06GdFoAtguBX1W4P97YbsZRFFNravJOCvc1d1Z5Ooy3CrlVKT
swP0nnec9UCzfvl2+u8eFj+GO0b/mINC/IIMg/TZLatL2nwyz1HTpK1VmjluXI+9
8Ww5xDPyc7+qoFN0B+a86nyIvVBKE8YRTzg66JmI6SDInn4l60bh3DhR6OyY0KqP
8W2fNDYSXavBGfATQmcT6xPdEkiB1da5vB7p/iY48APS7aLrFbqH3y3BsrYGIL/D
+dpLNMYyxjZJgPcer9zGZokg/YgHVHq6Ml3UItjHKygWvuYJMJwWyoTYrevnJ4m+
dZXf/PYC15kqGK0vzRSdpabDZ4iKgy4vl//dpt/OUomVb0PS6ZiyVWqnHBvly5Z3
ZA/Hqv3/ojDuxPNFbdQg9CXOqJ6uVSEb7RCC73YxlGyuKVOzmy9Ys8qnrqKajkyI
hUseVHM7+mBorJGoYc+1E/CRNDwFZZ7tYFhMz6aEUy56AHA9a9iNdvC7HqlZvyRC
tuw2pOjFzqX13yV0PuwZXzNqDI2BZ6RyXFuIqVKYQA++wxiY/ayiaU8io69kdavJ
d79cjTpKlPHB8r9YFAaY75O18PKz+xX1MEIW26igeFKedCGhLR4TVnY/lYXGRg2Q
UNBtYLV71mq59nG9mCyrFMi6XjQG/G1eRswRydy4JDElb3eLNX7m6BqjyGz4tLXI
zG2Kkn4H5vj0ie8QMCH+qqR5PaovMaP8zoFVxj1f7DlM5OQSJdr/JhghtEC4BMeH
pOUB7Lkjy0UajHtN5Q9B84q1Stngy3jkaR0pLTBImcE7OnSsUIGP8vndM9dFBA6W
bNjBq41akV+dDn9uNb00ImkBhotxmcU4Ouf+YF5l+8/jew4hqxIqPTB4GN+R+74G
68DoltuIXa1wN9XW4tBxkn3XPugfMDNBJpPomB/07/iQHjAi8/BgdH+eBnj6U1l1
zCdInLuOCyl1oglt7BzWcwMmUnVYWTJkU+1u68IqdagqryfnQsn13ax1sF61O+6X
8oJKyXpzIye3bvpSJuGW4V+753DK0mGfHM0Xcn/Zj67GzbLJ4M5d+mOotuJLeY8+
DjbLRSFtmj6OPfB8QqvqhN+IVmfVcKJEcfSpjd/PkA/0ZCa0H0i74/LWuIIvTEBp
zbdMbT3z/HqW8TB0MB4p4/pkNo/wPk6faSV8eMswaOLxunFxGknaLrXjGlKylcky
KTzY1GuVZDQWC+mLkZeIbnBwtkMJukahVm3/oNYR+1Fxc0RhDVXzHcLq5TKba2EH
d1qAA3XUayXseKyf1+bqnrxNhlZBLOtNAkS/RKgvRtqmMU3uFeXxA6hImJT4giUK
foXjiIW3h6OyEfNFFZY3BOhVU8sw3+iCjkxQOG78dK8+Q5bCxiQkr3sytc/c6Un4
0Yfhr3zXukwYV2oK9SnVb5evfVMiHyhdw7hYkNUtjP23NVuVZqg/wJ5oYSGaRvtq
ewbjPkCVC8vPWI2vw4gEyotyfQSDpykEDoWn0gawZH4Bre0PIIO8WfzyUHNC/8EL
ny5AO8cf0BaCujDtNfB6ts2L5mcTikZ8/Ul9MC+NzjFvJ6zN7x9fZA/cAhC+kWUo
CpvPoRikTpQib20qptTTaw5/uv7xYF4g/s53b6apc8lhXfC7LCGpIlNgSrOvYO91
z43KgBMknywA76PScWA6NNpcYHrt26iCJq2Wu+COPjzcHx87bSLBJx7NY8fsc3X/
qfc/K1ffyffmvTmEglgRWos94LDy8yiLd7ArvD7A8KkdgnF3ozdSIPckhYe1EvGl
V3A40TO8UtZpU7H1JoAZwsrcQ6imjua0FNiB6WYnzR6WLjVdDPg8Es8fJfkxXynX
OMbN54QftuCUT9DwhTQF1jgMpsBnCjqMnb8OlnS+tx/T4yWNIGdqqvBKP/z5f8wP
mZejvYMqirMhJIu8XH/pBeaqylyBgzhtIOlIK6TMwoPS7OZaVpkZhMc/U0HsAGZX
dfPBC9qXpnpAJjOip8+6E2605xuB6K7X2RgrdyIh9OJSlvflPg21Zckvsqv3HkAV
5qHK0XvD3uioh9xW11Q/3LtoTH0osb/IgVJRBnLe6rg2x8mPvbPN3QICrNcvMBQ0
GePQ0J93GzfA/KFVlNq0nvUoucIP+Bctn0UqkSBIilcpRnYVImG8cIu57Y35Cicn
3Rc3ivR36lNhCwJLEdPI02HHDiPMqDgAIuOue2V4MDSAgU8aPW7XxfyfR8b//x3T
bwXN6hXCTonnliZYTXxj67ANwDq68ABnBjDkKcsYIqJvildQR+COKT33uU3q1WH0
1Efhcs2WXJrAp/pi36htcvqmaNIUICl8z++xSYi/u0wmez7dr04ZPszAKcaocbdI
0RhEL4b1Z3d2CqWNO1NL4hurqjtKSpobBuNrheG7xopTebxu5CjcHQ6yuXAct92A
ddfACPo8zUMykBD9hOW9qWD6Sy401Nge9n68vnx9jrrKr05WRjqFCrFS0izfEPjb
yX7eAOgL4IzZlXfzZSy8fiAWVC1SH5aFMDqzNIeAml5qen+8tauqEyWBSnekCqn5
g4IApr8D8eBGY1tF/AAY1u1uFm99FOf8SyriQsUj7Gz6l+rUiCct333tRzLfFaQj
AN4vREf2H5YFMNTuFZq2Tfqk8pbnhBPYnkjXcPZTy4N/YG6RqPDP9MwwIsUx6fmt
8havz7sZO96hz4kkXzTeIQH/eJwP6ikVXLOfOeUprMUGPxBtfAY+j2YC3pUbJJ15
jx65Z4MUi59hNW6JPE8CiX4rugKnCMxJXeqMEnl7CugR2oNVfBSZFtys+kvx/tBN
JeLCh47WYVpQtOI70kC/SR8kIysI/mPAb86k0kTouGRLmNaZ/1Vo3NvKSwDBtLAG
DwlpmASbY52+FnrOGmmoFSHfg+PQnlnEcG1aOvd4N1IUnYKF9G82xx7YAE+JIc4e
wcF/RON9WAHyuGQvyTDeg+rzGD97fRyfpRco8yruMFMLNbxASX4eR8dcFkz0JubF
Wo8DAcSKSObO/h0FKmDlIeIK7fLzFvDPG9kP8kMZrVty5rEpGWqyQpMYC6eJLGed
Ih++eq6OqPuJKSjWl3nN1xVmKwXmZlevw7JtFlVXXKxF+KdLOHRjP6dxcBHOPUHe
CgoGrZHSDeCe9zpU7tESYSmyQje8WgXS6XIgZ1zjKzirOE/CB6+XPCgS7fHG0fN9
mrHUkSZ5WjKeKnLSLIS7hNA+Gx7ZwbCpwHF3h0oA8nCTdxyouN3Yyl54ewz497oe
AC7Rnm7JC1ooxw1rJKIeoVbn+7y/NG9TVvmscdzQ94hhTbDqmCZtM0NhlY4ScnSt
7L7+f1g1wDbwURp+DaiA5hUomM/zrLI7CraQfvCfkx2vaQ8nOsk5BaAfr5cqQBDn
Svmc1SwMDkHSuylKdqkpU3KoHemRoAi6xsLDwC27tB9tQsAQ1AwgAoAav9mRIzoT
Q1Q2/O6h9ES6dCgN0NSi7z565uG/U94SMn/w6Z9+32hw2yXiH8FChPJ1a05lHC1a
EdrK5crdfYphd4SIZ7uRTOEirVsJgywVVEFbGpG5hm40w2/l+DOED3plimBh76U1
7IFjzGYdNGjDkeeP6ws7RBjPEf/b/IQCiabjF/FinVE+k8xXiUyEZpUB1lYtl03C
WHH90g7joaOhyLKtB8A1PCZqw0h0QT0RlbBp4cyxctwRRzuL2OiyXX+VRdbMMYdf
KR4J/BDmvOSflm6E2OuDM5ysBV4cKEZa0BXJFIS9ep++5WRBm0ZWPyb4EIqJY0WN
10EVrb4yVhXkXyQagKGkxxizyJ2gR47aDq49Q9RqLpUGpaBFmsi0O8j2JA6hCiaL
p2oWNw87snpGI03Q99K2myb6f8CdjA2aF35Wr4xa5dqoxxWWE0nX2hi46SXMWGu1
8qyRFp5kSRe1C9Bve0k0hbgx1TnJNynqijYPbO3VIA+WxEf+b2kSYUy++FA+Bn/9
5UyT0SG3mmtEJx8JYH6griUpC8Mvn5rcPQsJP/CzSid/u8tNiWKBqkU0jTPe90kP
ashR/UHfmm1f9hUEsUoj5xU6VJWo7eNvXkHaNjrtPuDlS0Zr2clcEPLNy1IsR2Gl
MrNSQbEQO1Gy7DGwriJbwUTP+QFu6fZfeDio7s2yANjLMs46xLuGyTyzJYNRXmA7
mfWEi6jTH6sDszhEVLRr4jp0HMwYQWXEpo9kZjWeojSDOnv0X7xLh3zGPCCYzfET
3MA+UGqtIsvhsvFNnlJ+H6X+sJYS5GDldGjhCP3UnLXoBxqajAYAA3wwv1vGINkX
y0zUKnu0ZY/AHQVD1+ERuBfImvWOFsZPdN71NVEOpTfbBh+ctvAFF1JyCHBPjOd4
dDh8a41kpl1XzzyWlcf8c+IYNI22d+f4sdtf9opc3VX3Lc//7f+Kr5rDJshVyr4j
jOXTPSg2nNANllOIBHJcJBkmJBv/3rQ+W8tEzWk52WXFgAEstnOGy5FPlp8XOH+7
rR+CNgC+yb/TKkjDUgpoHKvP9mrOu6HKCCL1GxhTicTs81Z6pcOh5BawUSKCBvNe
AixmHZsxTH5AdJRTFZlqIZGUGWsTKbeKRfIvnzd/Pp59m5pxitbJ2rsr0peb0vtG
HzidyVUVs/UnCLrxaw++hxS66Jv6F1pKkvN6OPMYwEBtdHzDaJqVeuuJ8FQXD10x
kxDKR9BviJUdRiEFVLdcBBsWlvupgJXGoZcxEkVqMozJBu4RwGVYCmNXnDgr89LZ
pRK7KUYAVjCRj6mxnO9oQY6VHMaqxUu/8Ag37jihk7S5jf3H7xHIfss5L1pK3dM/
u4fDZuLRPsKfUQBk4Y1Aot+71xdM8bNSDlnCqB1WQMTdOkf/f8VEMNBjS46oka0r
6c4nMHoySFI4XZaN2gGZR6Ek9Lr+r4P/lRFa4jrEOKnu5i6RbZE9/OZJpY8HAlGO
FWsQkNOjhScE00Nnlyf5OiN6Rrs6pvo2l9gkAG+nQJr6SQmCgA9CnBwPPons2JIY
PuchmPD5+aBjG2JWo1x3Q/oilyMtQAe2eodTKIjJRO8OVs68BeNOFfOJ02eTtn1e
ky/yu0MLlOkmY+ukupgM4gMlYayAEQjXuoU7eGyiGd8LejeFu2qAPqujEAUBt0YD
NY+0o40cXULq6sGQDrQ2NbHh9EJxhFIZjnPzYxztlmxVDoL5wNW/zmmF/+hMcDmp
S+aWtLWGjG2+ps7qnr9ajQ0SiGt11t0gGQkorQW+tRbAImSozYIixx5vKpRQBEAX
K9r5rBK1BHSJZ3wevnlVIesjAlCNN13lSBAks9mm0bQl0tY8YFfBVpUuypFR69yW
T78GqHyONTpwlc1N/FBeh6sRDPGOMgyZNI21tC1SKHh9q2KolEk/5gBoQ8x9Xsz/
e8sKjH4duSrF2SOIWf9logVCeMtn2oxCVnhzDdvHfcjqxHNGv3mexRRCfEC1XsN7
MkImNR7SGBwmZGS/+h0D6/9EulPO/so6IIcpoKZLcbFCsAdGTqAZI+shVzTcbu2+
uQjC2wW59esKr0oV308lEKFmJt27DSMHsjMNfm8lzc8Zh/eeO8iGZHA8NzGEYOmo
RfXb5b/g4ybJXzg3eSjTX8n7qBdJm9IJ6fLbc4cmiysIt7oE3KzItZQ/qw3d1pFV
mgbkPa4/TFhkPEfPXCjaVM4MU3lX3RywN8568aK4c7TLjDoMByys9QfRKgospBZm
HQW621q+JSyAwUfOPPcsCSuywmQJ4McyT3RVeDbwrM/dYjjBTWM1PKd/iYbrrRaV
nFs3FDhqJllLo0qBAhuaJaTaQqAV1YUqIDB1KN8g+ndPDYm1mMkcNXCkipHdCEMS
KCl6FSf6+zGptsmysjHADZeiyjbQuqN9gefAkJamynusr4Pb6Jk9+Ke2L6E+tiUq
4hnDXhSTj2Gbqa1Y4C2sBk3uo/OAAKvZhl1VC85K0UYDa4S4ydxgZFYnjTpuOdHz
0LvppO+EgsgrOdWPaW/Qyr225FBzFJ9Le8HIMk1nkGeV0W2Lj5KiIhXnoic0S0fT
ETGpavumIMm0u0rF5DTPnxOJq/W1GmRlnThIA3wK3PzzOWLu7x5e5oZHRCoKiQft
EHSs+Fqospn9SrE5T+7oj/cgx8CO6KYLk2l0Syprj5ljWHVgEBlptjVMPibj8Aj8
ijlj/J5+h7g5m2Va5Oy09GMrrJBQi7VK/eHg5m2OKx3yyGKn0LoDEe7TnOZeMxTr
qPBs8MKlw1tg4eFDSN8eRlCsDDE01AFPQCzupo0hjI7Wj9jJXoxztm/EAUd1Sy1R
tkiJLo5RudnLyHqyXTARLpnyAinQKBL8xGFDOHj1ipACPNbkBo42t6fMCnZuE5Ty
KfIhPq7QfJyugBmfaZgu29CIoI4Fchq0rGAyZXXANr2/g9gdYOVfeXTUBMVZ0/aT
4sgADtG3qDVNVl5fvTFTFcggm81H+FMXkoz7RRXeduKGPybPJx2Nqzlb2GI6D9fY
O6vogDlHWUKB7K+DUcHw+HfVrI/xQ0TTq+Gslif3zMJriZqvd6Y3VBz19y2rOO2h
5j8Svz2S8KB1cngs2TLZ+98wKXdI/BTeP+YfsuCjXr106e3bW/EVIcCe+gy3Q5Pf
bL08dS8TWsTrOCEqeQu04SOiZYhZFp5CCn3gdXqFo116pgewcT8j5X2tMEasJH8y
MA3CdxlqHde2Lv1Y71Jix5M8np6taKq7WvCd4vNrVBrZK3uS5DNLKGPXuCQKXJki
dMRAj7/neermG+jc4uC94aXfGy2C7B3yF8OvUS+VQBoCPfPmHY1oqjYqZ9mv8Su3
Uzv8AueFmk4WursiUZvdLevyfBM16b+588tnlxdmwy8njhJErpng4koZ33kO1jDM
5t2HEKws1oNNWN3NCVM3G+9a98eA+g0Vi7A7eij3gPWyozXeBAgfk3IoAzHLLzey
lB3mM5/XqDhnXSCp5YYJQRhU0XH52GHhQB7MHcmwf0y8+wZJ0Ytn1qFxKKG+6Tv4
RpXAKm2wKTlQGN/CgFomBzWB/q5qB0gkLq6/FjsqRDVarV5U6DYpDXKcqV1415to
xSLd+ATIWHBsZQmLHjJ/2WPhMWa2+huHb0TfK5WF5eocfH/rDwd7yT4frwlsgf1S
AOlWwVWvZ1Ll6FUkF74QtdyVYtQoqg1S/aqUCDZdRk7V9PjVPd9sIuDFt74bX5y4
m9JAAJKnwenlcm6EzgCay2hbMcnUGkOuATdBBVh8d6nksZlQq/eIQdznsVcaF1J5
qNuaFYuWXYCeEC/tTp6ZJLJLFbYN+Qo7ei1OlSEzJD6IKHpNc4HPSgFJxyI/s+Z5
PYTEyZPfVnBgb+x1IrajCpXrkc31xerjfw0V4INr0H/hV3Cdzopdr55M9j5PW7Qb
kLEFXY4Mt/O5uh9bSPQFva3AubZXgJSS2R2UZvkJ9TYjLxl2y+KzNUUbw3WliIIo
SUXVoGQ+ORIMnaoS07Z5TKSrZb1pYMMnrZ54K+1fG04h7i4kulbZbzvm121/Ksmu
w+StGw7u7DTtBP6UhXg050V/aM7XO/EymypY2w/YHFvV1O5g3rw7BfEaWnTN0Qs8
zllk2P9pfkvu2AhMhehZSxtBd+seJZkop3GIqQ5eiDkTcFEg/e8w8aLtPqhButZu
2RAw9goOUpbOZMecUw5SLn+jHcZG2ImYICIU1DZRP1NWY8tr7sl6gKzFoLlbipom
H0ImgSD10H7jU5yNiynM56n5ItvSp3Gn5TxM0X8/5SQnV7mcKwVTdLKS1sQTPdvU
0Svk5dcL2sBvSFXR8wVL5RQQWOb3HtqI6wVvvqbMJ0j5isOn2iF+BLjrITYdyFgC
h66ohCD7L4xUtk8E4LwGn4R/Hm0Y10h1Xrn65nrA142vmpBn3jU68VlEqBu7ETom
2K9MyulTIx4I/KtyDqVMba980doWJL5+OkjH8mgkvwpu0ZvuTLa3D/Ge0iqoSiq4
lI/J8pRkKGIINneL0pR4dSZTs7eSMO3LlBkjQGZR+DytLlssqLcFq8ufjn6FzxX3
JmAiFfC9OlvO0wVxSd1xKxlLZDsD1syMutnhcbQzvJ/XTUDs7pzryInnunTsWMIy
cABPmGT1LD9Bh/N1WH5hwaE0Y/yFjGSaQTBinIjvWoyz4+gElXqBoAVSIORj31E3
N+1B1WccT3CMkHznsGa2BMbNWuxuByBatnjw2Zg7FA+qigxOkQWBZ23wc0eFUCVq
6UrgnT+e0Ivm7zY9ZCL9cHxp7kxs03FH8zENmHPIcsXqhchLU/7rIJ/cgwV19S9r
71j/joxy0ewsxHfqEGjgW4H6Z7bVCLr+QiHOwMIWKzp2L4Kcc+GBZhvnlTo0XeZX
mvkrs9+HjBRqae5FmvtYGDfXDbrj9VFuK1xw5xVShdpM3pyp2rmnkB+I5eTIf+pS
abETY89mdEf3HySVjDOgkfnR5mZEE7eR5i0AZPHKkVy/Hm9qlO0Y0uWQD7L1FtyX
INW9DUJviCHi03bfoQFTqGDjW0znWZNky+zbe+fQtTc8ux/HaDWYVTXsS427pQcN
raRD0yi9VNETfH/k/zEdEL/ylc5RLDzLNSc1uFQ63CYSXPGePptsEnlNa4vmkmw+
fZRajxSEa80lngHtlNbJm7AMNJZfEuBPZ3sL3eVY1ocR9q0304xAJNRFV0AnGIe6
pD6Twds6QsX3xILt+CHZHu0C5W5bDLczrgIHhZ5keK9Z5uaYNntx1P3wdzcekPKd
`protect END_PROTECTED
