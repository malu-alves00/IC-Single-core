`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2/EeMpPCaYiKKX52fsgj/n3FIAoklkJ+TzFPXgsIT0YkP4FTqIJfiPx8J/uDSKbL
UbGxeKQ8P5LP7VUm+VLwqUH3BW7OBLM4MMCcoXmObaWaiMUVI3v1sEcWTKtIx/4g
jI219lv4CmjDloVlB1WAu7h1MrU1EZZye41eOdkde5IbSEu/kpoACkVaTvCeUeni
oKjWw+rc2hW7P9GcXfklzw6P3bsdgwyb+cUsyemyRl0lZYhQtiR1vWuD+ftbkGzW
tjcRQMr407BbaF38wYZsK6spYET+dRhMGRzJax8ty0b28/hSb4VgQbXSoOZNNovu
mUm+4kHEs2bfBVDLO/+oiaUOxnUToSjO8NEOAsurMENVaTMEDp52+fglzA1uFQCJ
YluHftiGK2VLFRxg9qMXXPqxT+09ZkkeHlP60uNyI+C30u5xOSdbife9c6Qf4KXK
xjwE+hqZn/DberGJxpba7SMc/fb23NlsWeaEmJ/XbswiDIBn+/pT37aJjp1gQ8c3
vWC0E4ujK9vGu8ANqJsmps254gieVQohKWHLnclvujyeqqYPshG2N1fW6/KUG/Mw
NnDK0ssaOnMpXbLPFb8N6AK3j+SQcg28QYAW7OejqKc0YrdnGzfl0exbUcV8yZX3
FNTZwA0AV5SUlT7yXllW5r+Wofk1s4VC1nDJwDn/kGZ5vnj0A90LKu07z49Ax6wi
DglM/3Q6VXvZhZo8YhfUUjK0bjLXkESe6eLOndWLbxfw6Y0UT479gE6bp0X4bG2z
z4fdIX7GfBWlFfqZK2udpapN0Oa7RF45wKLSPMBjgH0cXf3bGLI5cZyRi6u+eVy2
ogzXs8NNBRvo0CSz5b/3gWuRFez9P25EUdnmb5aEN88wE0Eu4YK1JiUJso8zUQqU
B3qD540QrVYQsvTDmU67JsG6FNxSTthhSZM63oIyniyB2NgCgYULHNASL85xEz9s
rolrzfR8rA3O8bJlw0dHkF2Y+qhD4kENwCVhC1BOqeFoS8v3gLG0b4y3ZUYYErUt
r6DYNfx1a2XGiOsYR1arBcMG0fiSbF39NKZdRzzAfeIQKemfZvkJiRafxeeoIB83
0PDFHqywl5lvYUMu6wNE+Zu8i9G1gxMl2dGX51o0c3Q+OO901o7dOHkMYXF+lo3a
30YGkb25uo1yWJ92hhm9EtqCxfAaZMcpWaJhZla9S5tRqUw6Mq/WBvVtXbCtpnxP
LKoQT1Rbzpv0sknAfQ5uXPKxnC0ybEoAX1fN/TDHhlXiTES7oea79VsPuVecnacp
wpM3YvJ2yIBWv891e/+krVh8pf/74/EAVOBd3RrBKS5ctU6yuNmsiBXEBGK5sVDb
DWCl45VwPJyZ65qmXbeGD435UYVtJ7pT6k1LOHoZ+kxk/o93qOJMPWMJCXofzvVr
yadJj5Kt2Gv+5sDOjcJigCOeZuMvEGvJHbXkJTQDZKTwnK1L5LcmLzdz5hhPwH5w
3IUM3ajsgXAg6JVbpQQLmDR9uI6/Fx0vLUOtGepeNZGqHzonfE8A4q4jOxjHNAst
DMi2sx632ecBse8OAefDEe9d//KLUpAoJL+UMxVSxB3KNoTLE7/wosUvTS263pnA
ZK4rYXCIigAIjmpExz9is0SvsL3WqSsGWA/dk52Wfj97OnhrtrtaZfefgaQBzhtS
ZP03Ko1RwX7Y93iyiaC9aOtr4q3F5Df5ZkUepecV79G1ja6TNsCfmlPjeYJmZkUM
eAzODZ1oL4ZtKQhJSWjkv6ZE+7m4lv8zN9+MwnVmYdPUVl5bPG+Dx94OUU6UiCRG
MPng2DbS1gj8SP9SpS3uMNhD+LiPoXA/Ukl6AnSHqIj0WHoqhlzVkLqXekzZHg6S
4LqcyvXg1JeKDV/wJAGuDRoFd1D6IyCfxEyWwvK/bqbVxRJsawER0hvoXFnSXVW9
6bMOLebtdlgJ2pzSWiOXAfMNSd2r6VeeLs5UNZtvMNuD5sGhMxSaKnWg7iQHVXxH
vwUmjb3ZbXoJAF9pgxz24OQ2V5RVZH0TO6uQ7fV1DzAkm49+SNfe0iB+yvBrzEFE
fRbVY4QfraPaQYJparsO0ECJI6RddgSZ+oII+Zf719jKtYZcHh4kGiW2HD2PV5oX
C65DPvWmJgo8zCUj0EuucOY0RFUpzQKAJ5crb+GNduSAeG0nsTKaLi0Cdp5Y5L2d
TZYNmpbxU/8VDeNp0xvdPqhuTz96IV4200ArhCPw7CYFuymPqmfpR9FdQcVxMH3N
drAiiH9zkpQ22uEC3IB6nR7eEHeYrgDvxpbNfwqGceLyJRSj71cXwu3LHUwMg6tH
PznVuPO0iSFDbPeVIfdW2ddJ/hkysSxm2JZNiBma2hm0NgubJ1u87KH2mdSQJgpY
U7JEShpGT390HY8+j0LU5Snoe7XQ2NymZE8MePVD46am9/T96oQkvaqu/u9zJB9n
AfvU/yqV0825q9YuKZhBUbMym4MC6aWxmjpyn9l5seCGZ/83sLr/WT5R7K/OZMzB
/paLYudfkA2TzNEKUnmyOyxRJiCeOqpYTmJSB+4a1TthvoMOreV1w+g3bQFvl5DX
NdW3gIGTKHxInxzGrm+6KfH2rQNFk0kG6eyhxAubwqSxBabEG2zoOm2urgd0NLyK
bwZ4R6fK3V4kDj4grVoIqY2Fz4rxRalesgcAyLf1vqsq23Bu2Uf0MIBjauXmma5f
tS8cTZ3l8UblhzOeSvcokixNJ4paKhJnAYCCP+q8HG1f7FP/bKpuwhjNSeKSciCf
YElgTHUWshvkVF2LLmhSDa0IDtUdNk4JDxXuqEIKsVMKlWNkUfUGX0d3Ff1dnRQe
FQbKQJvtEHH4VdvD5ZW59ohjKZcSp5SzAhynn8x3MZWHGILde4AQQBgGY+TleXAc
UAizEp1lZCPjoEPdGhhUWTdkwBAcrk6vekvVXVWZoR6D1joJskSerjCwYTgfzkig
yr4Pfxf9T7HSOhWuF1e+rlMptYhPBRghjWN7+knWR5SwnWwuunoBEX0gYsGsjJc6
UqGjmfVnG5E9tggZAuNkUOMY5WHoM6Plj/tavobfpS/bPhN4B9EehBUVOt7P6fEy
LVhrNcF4V+fM3+X4K8FAwn3SJ1h2/3mDMxysnfUomJYzsRh3wfLsm7TjV3PsRCWm
dmT4xDO3LvFGOAaIZX74VCwnF4C/Ktr25eAhEIl5FVVRgENsdgs+ER2tc1VngaAK
FotVCjoBgkPklJuNd6NsCyC6+ID/CHcZDEO4mbUF2GmdxBwjFBD6ZQPBLYlJx+8L
hSsgewNKQiy+Yt4g+rVyDsePWExjKvna9WK0IGX06IrN2bLIAMZLwg2lBFjfSHly
fYr+vmYV9I+AZMcEVquFCgWzxqYgWii5xzvcN3bO0nXx8SIFuBP4I2EwChy4cVHB
qRXenh5T093U3X1uJ7D0e1JT/Ll68irePP54vxOuKeJZmN68DTfuqsrWCj0Ns42j
6gDIanuRi392Jq8X34QBN2Lnq2RS19ofQoiwNmIRaQz4z9jR8JbKfwQHrG1io94U
8Z4W28B/uUqv3UG7df7HHg5+2xCnOu56EwCiMNGF1xlIDogpEMwf66WbMmtXp0b+
hTidXuzfXANNNpBK4zjlZK76qJe/h8lkWBePKa6j07okxaZnmTkUrs0gRDERaBNn
i/dGL41BPZnXq6m0Rx4z6tECjF4k6s7Q82gl96LWNUo75yEOKkiLFI0QZSxwv1Ea
69YXc07HjD7gBXNVK/7DE6MC4ybzO/AYHk3O6x+CkgsQLHp5FaPjr7HweQt4X0I3
3+e8/7geu0lmZ5U3wBqBFpGI8B08haUpq+AqCMZ77+KRFJQ7z8EVMPwXizFrrTEh
69b1yJUtdvwXQmfVKH6JlVWok0tJ10PTeVZNDu9pO5/vIOGGmCBONxsMyt3EwEVg
9vEga7Y4ThqAdglHV8uLdfEwtc8AME2mOr0osTBHMc07JWwGgrYbDRcndqGOe0xO
eIgn6y42S5kY3ZsM+kmQZ3ZlEwQ2nfyq2Dgf4M5pAgYL27dI6wbZNzk4rVZ5wn/g
3XQUr+0uCx4BUXy2/uAXF/PaEKu8qtnmlklG7qHYajup7g3DwpMe7F0RnsRCPer3
DV15aIbnrkLX3FTfYcYzoIHpX/2x6Gg5tPRK5K9z16nKDeqOZNnND8qFkoNyI7aZ
3+lIVFSj6QhBZDAHvDxXL8RWfQgFmUY/1c3d0XPgorwTeb0oIcAXXTlvpRPZPNEX
VGKi0XP2Ps2aS1RLw38/nc5hYbu+jOrjWD9mRMQtebxke5PexYKD/nRN1wQnmxS5
7aUt66yhOEisW+ctCwls7/hqviLyKhcx/xOaryHYYGwe8adZBPDGxpzuJeGmAkiP
pV/agSoXIaA6ZXlSczCVcLHZHjD45RjdBnL6CbN5T/wEuszGA9gKpZa5PXleg7Qw
RpO2NzwNusxrRUjZSerFCon00xjb1UM0GLVC3TiUe9bcccO4NoT1GVqWW2G6xTqj
SWYqnHZSTwSCntuOxZfppvXq51IvbJSj4QxAYastF+8iMJFQ0RpX2aZdD43WD75L
RWSe5n5CVLkGK5G+SmKAg4CExlhR59S6EYSt1+3EHCWoXoO94/lsTTtjbZTraMmI
QX7AgO92ixbVhdSuyKCFM2s1lwaNcrxTve1NxI+1rc1V45aC4F4ekV562lyMMyk8
h71gRTJDN2d54YcNC0DpViDIE80LzrJMCzxie7rSQ+SHq47x0Ic7TEA67N2tXWiP
WKyqOcae0H47HL5ehuJMLc2y2W1kpOCtCG7J0D1vDmAh7UchimfaFSlWxnz6JXMe
j71fI4q06ZGOY/udHC3J/FgNBdoPqcxg98DLgXd7Wo4vE0CL7zetmEs/FYoHwQFt
eWzym9bsw/8C1ExwqUPcRJu9AdfXY7Q2N9qB9BkBCpTwjy78mCPA5u9C4FEbfyX9
lPCLkCvlJw2BiIcotVnTVuLlNdHyNalxzb/bIM8SkrfvK41FsnrC3mJBlLaDtUS1
a+ePc3GfKmwDAeDZqii6LUJpdfUyPZN1vCKrDjN900mQk6NeQ1x7uYBYMgACmvv+
g672pPr0x+AvX+mh9cF8cqWBU+kYnUGKnnMpEaiB2gNOpunDvKeCmJwop9Zso2Oh
U0rrzOMn6nySzHvotjE4clgN67xD5SzH9mYinPOhoQCavQ7ppjxFn+iVJPGEDrM1
3krlFsmiggDiiTPfy8mWJe++/LZrZeSU2XECgkEssxwzwEews/9qDrEKk8g/Z5X5
9qZyeDDdEWVQN/MXfH8zxgeZGcC98wkH8vNj0lV7SiEjjEqcDdSIpO8saO/g7lOd
7abgfCfpcfJm19Qj8m6Xm2gv/BFNWLcHpCWi5RU6wbTAYhs9X6l0CISPcnt0PAp1
aO2l8ECxMVsxXH0KlXH9v7cCTVn5hT8FIFc/wxpn3E5HFI/U8ulqDzsimCKplD+Q
To/562OF57e+ue/ZPJN9uA==
`protect END_PROTECTED
