`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DOHebAV0u3RBzzEcKsRpWQdWIoGj6A0BfoP9tv/0cFygtTz9UMvtmDdigSrAl8+3
RJ59I6KktchnTkReW3yvX2xy82/93aj14UA7XzzXeymibABeH2Slt/qH9m3Pe3Yl
ZDA89Uwd7V8plKGrkBmM2/qDwO5hhV1TvUKyDWnHziGadIleiXI+hrrNCoWtvFQh
7BuXEwhqb3SagaoiWGMVPPExNQz7VlnYjbb/3fl9/ZVxGVG5n0MeY6MmpBSXjULW
ZpRb1idy6rRJ8kRQrUraI1sVjrfciRAQqkI93NpaozF2U1fWl2r/fDF5FmYtSsFt
6mPGVA7ckl6HHrOnoYaWmaPfZokbERzFpERapLDP7kWUYK0bWjVlhOywHmEVRt1U
pUAFQIlOKAlzYDwTSCbiH6MRWaXlspQ59MsiQU476sIFvm1Btb7d1qIKDPT7vyQE
G33DfWK5rC2di2pLA4waznyj1Yk6dv1rMfNeBBpEmyio/H6DbZvPrQjdc+j3Ht0+
NJEDDJEwBV3tk4ZQnES/YeLPgTPxfv5BbFFrwRkA7OOWqfrEDm7VZUx4qYtdNz3g
5l2CzWuvPcQZTZfGhSa8+LeCXH78BDVXZbtWGxeFKUT523aF9HajS0qzrgayiqsz
oTx/h3DD9nkLVEQ3cN8l4b2zTQ3NT27/o0L1hITxH6HxQiTU5oFr5kuKHcLH9xat
UvuNs/ScQsjY+irL91TXnvBGMk+C+malJhw4syfUbX+ljf6h6BH+tzn836G3qwNY
Jvz/jf/an45nM4iJmJFDHEYHfwoFmFlN3j2bwB+4UN51KCa7ZeIei3U7EGH5x293
m1lqbp2hjEU4b3n51E/vTPVsPZuxkvwiyZwQgvn79VPF6O8XCrtN7NfaE/Xnhs+9
HkUkKf3HjYSkpBlcWzWl9t+grGh0UMwxPjfLfE+9xlHeOVD0ZNq2dgX5vmWoia3c
8o5SSVFBsfqUn9NmwKA8gkg553+WJ7MOnErlA4/KsPies8fA06f7eSHNemXlJ404
NwWJFWvQS4Jr3fO9BjP7q7vGhBUzi/5Lfpdfwb8Plia2ZDyLOUvutx0fbl0PsLSI
VCz8L7jdmO9oHtZURRIx6PTXGpf4msJr6TZtzrGrMTL0L5gN8nYH/Gwia2dUkD6M
p3SUDwyO/g88Rj4xBbvDoVqeE+t4mkmTwgLAfa0IAqsQ8rjwnolJEFHBPvB9xy2j
2FmzLNvumT3R2lDAjtBr2QYUYo6HUyMSWaew4d28JZcgPQOcIS4P9RRV1jnb/ueJ
8Qz65PtXLXvmjkTyck41qJGUhkKKwEVz0T9b5HZtEVj04wlawHLJSw1HyntuSAzz
4rTjrUJePMjAb8MKB8sColgoYA5apGj++jG/f2CbIZoSZ7TiXd4cK+6LDu8APLTX
9scXEtsiCGH1KspOJ/6OVumlzOIrrsQI8AkxAtl/PsqlQsEyfCsssOJcPzQXggTz
aUAPCm4HHfeCPWPczsVj8w1KsAXRJ9DiLZpJSDvjI4zZ2t+3OJZHw+OYlkf+1TT6
1CyvUeQgq2/2HcV3mP0u6MiIPktto3Xkq280r+Ta+asiL1IhGgHKn0RMthWk1oso
f43GeQFYMwqr78UaflU3jAD33FVD8J8ZkKdVIZeZif54soEoBOepExBygOdE2ORw
n1Fxyqnak+zR13SvZlBmIPHU3E08JIq3w2eDTgNhBVCBxO2gP4G4LnFXIIq3yDVa
FrwtiITlONuGabmoa5f9jJovg2he9om0G9MaZ8RtyiC36S9bl3q+N9rwmfTgDbMN
WytjfVcJM//U90juzX8NziuYiIi4UnxxUaioTtgUZhlQElbLfWN+9wulKHsdhvdX
L2kjzYkOkp25M43w7+HrSZ8Bu8yTUUKZZ5LFYUSabyvMJuYXak8wCkyBzxpWVwky
g3nuQ0ZNu1zktPuoQSqawJ3nWgv2fxL2LXhlkWYKBfFl+KkeSjT5pAdp44uzL4hD
Whl62bljapLreb5PEIpEzEKEU3rGggS0aBY5GagtyMGcBukUwToOeiFR7lSoAQjC
Ml46XE+oEmAzMSh0gaemwTupSwSIwRt1M3499SaDrbJvWXKnWJRVNIbQy50Rf4G2
OM4ZAcw6ueJ1Vydznr2TrIJi2Vf811kWzCkqK9c9OCIF8KvljmS5G1wonCX39Wv7
ydym8vTuYucZdagrwDcoYUpvh4gJLlJlWO5572J+BJLFEClQqGgzwwrEbjPGBXus
nAYAY86ey8W0EoPTfzOtGFRklQ1aUKoybci6w4EiSIlWZQv3azTzTftPVgxSgAdN
Gb7sU4UmTZ3p9mo4LxsVmh0zOZS/mlcf18Wq2AVBiqKZVt0YrBHGN3KoaVLHPJdI
jUnvCtLRBHlia1ST/HIQCjMA3hxwzZhxcJwnAvGmGNfJ08IXrioaFXlw9wtutpzi
wLeK10bg8HHW9zE1HMPsverPM+xFa1qKNMoW1cPhmuWig9u2cPUlCM49xt+4i9vJ
6pnmBrsbrkHc+qUvXPSCMgRQluQu2btzvDeYP5ZGQzNpRah5sT8sQI3CjB3Ye1yk
iJB7IazNf+fsmMGOFFcbuVYFRVe3GNik1Gugvl70TTlTLr3eDFcJ8BO4uXQrpmvD
AjinsSLWSDvOZ2hEYVyz7DXMkd4jPQnPCMU+QpEzuJMbkj8EAPHXb0hxhBO3Li8A
71+qwgDA7xJNLBL/d3AEggCmGicVasR0/OCQbxfyiROAmGq15uwU9Jxx/fk+i0+Q
+93EKT+5sEbPeI92wKdO+qa+xD717KAIsPV7b9FgpaZce4oAKJM/aVf+eUqACc7O
pTTScUl1DQP5FTEkdzXpSAv2TW2uvolldy/4xW/MNhbsA8ZHort6APToZFFfXSLZ
TQUNFbZe4rY8Cq/Xe4pUK9BCkZ8pLDzzwsZ1ZBut6bc/9FN7wIWrE8cajmbMAgzS
PNEORuLlJOF5mk0TUEzD0cL5/buYrTBj6UKQcmsdPATeo+RXZPryA8Tb2oKvPuRd
cEdm8BoDgRHGlpuegwU3BBLcXjZ59IKtVjqamS4U/mU8TTXFFQY+T4+eGqClmfQb
eGFRJivHjnxk3fftG30JNBoZUVnJ18B2RPlRLCXhk8NvNYLKO8+BTV9uUvKjRmuC
PbtlLhut94O0lcikTcezJaeGAwiOxCH3gEHVEePgppdrMuXem0LKBmPiEPJLUSEE
45O2mdCWc2y8lbIil7acoirY8qtxrf9TQmvrpbaXNfPTNdo/n9E3wnUFSSz8BqW3
PqeM9M3dpfKh/p2xJju1DaLkik9uECTu2QQi0oXOSIYeJlqKHa+rrF7OMxwkEliG
BGphYOlgjkZp5vELNiyXOebhilr3gVEEE451iOEA9r8Ugtnm6G+u1sj/XB4ZLQNU
05BZJU5XxOXaXNZx9JrSPmUAT0xQjHnftgw0T+8u6k2XunBzcY2kzaC1gKu2GvMP
RmhWQXtnOPc5jfkSTZWESldTsdO4hzmB74l6TuJ9bjO9fOhkd6NHFTjcpnDEK/CO
gcihbLC3eWqc8O+3g0kzPthFFL2930zs/dRYxO03DjlHW13VdzPm5D3ydov4spxq
UOrEBa7zyDnIvjjbapNXV9X0L3xvtQTgcgZUbjSEqO/SJHe0k4vwjgccKxo1Zlml
km5355HlOdpgmMgzg837D3InHPaWOQ68fWIA93Rl7y5C+DqAQ7ODL+Lygt4TTvKi
8+1ZN/KkGJEnpUfv3BV1+V9ox3RP72UalcwG0h+370Dok5DFZWzCDpEYMrH+GJwq
LHOUxwi/fysLSZItlsiE0R3NseBkUQnX68Sm9UnNp73Gx4CzCT9Frxb7Q7LGbwKR
kHMFY3MPV7W8EyS3534Jb/pzl8QEai2+PHMbqxPwKY55tV3io/NvmlsyYB3HfQs+
bf6B2Qx4K9X5bkuY7wUgTfMkF07kU6aU1bV8hFaLdyCKpAHMMwVBhetyMMmGOR2U
UTA2e83DrBGGbP2o9A7/8CXABij0E842kdlMQvHI6AUmOfVBx3VqmHtNxwf/W8ML
skipgTZS808Jizs6HkRHprs5T3LBuy7i+v8kAHMYG5QH9yEfgqMTlHQHk8+1Oi1z
3OylwRL5znsZrjD2Y89QXuLCC6tBDo3CKlYERfSa8MQUGb5Zs8YIrYQlSFXfyZSP
7agK8TVHhalldPkHvXwnKbcdrU91QOdpwTzjI7YSFtep85N8QAxWRTCg2k/HYkVj
K/96gS6CWwi3KPe3j3wRm9lJei+loRt7/4Qs5jUBJNaYyOXnO0k3LrgslhAPHttB
hnrMoeOXqITudrji4IMA2hNS+ab4FLDOhdtk5lRtCnZD1gS60gnuuUI/H9icmK1w
QPwJsifqRI1yQRv8cuN92Tmz9JdcWv10Dg535SLy6u7V+ff6l6MlpvP50t5OK8ba
QYNErnpry2u3wncnjsdeqEEWC+RxIuS1r8lHkxLLkW6DaSXtHdHZDqpLL4L/ynho
t66AAXGnEUMvrXdhNWl8R3Rph1AvrmpfO6kB0rehdpfDZkPEymsY+aOu0wcNg1TL
mvqC+p5TPiIXqLTJc+DX8c5UW/Vfhwa1IxW47oj82MLNnyhDcHEkkGVbIkjGrxoW
Keu1eL2X9By9hqDN7hTUF3SMZnVSNCclMoQWnBwOj3X6NDU4ujV6uPtSNRYMC8oz
tE+rqToHFwsuVSDZKqKY9XwH4hYvYcHjcNoxs45Mhb1VYhHkh+lbtJAzksOIuY6z
6uMewLx+oLGoviiQ7YvMYvP5VhEdnKdUJOlBYVu4OILiK6zQt8M4z4KbcvUVHVQb
jUetvsHvRDvTSA/jeTX035ZsBWzALfZa9qBuVBmR1UQySysVSEoFnX+zGRoC+lY6
ySVDBxg/q0bxxdMl+VNSEgcVlUnKvBpa8SgSJ2ElG3EGyV5kDrLYtLfPG5ilXzZv
qy2twQaMkJZI12+l/EJEMDZe8IGdtqWv2Y4DawsU1xc4p9YUUACQboEWc98A/jzD
SW1BAH6NDlqTknocGorkTWAIdR5M5IPMO8uzMyUvSWf5qTsNgiZJd2oFPDHhEz2V
+JvTVS1rb1YRwKYB41kYCEhEeNb9F4d9aQqpA1YU/RDqWEJHkAq0jWBn7uizuYhK
`protect END_PROTECTED
