`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xFRJzPj+qcE4Y8RrQpVWYXf/xdplVfX0BZ4EHSYVYIm6+m/Mf6J/0Z+Uxc5znLm5
ERfFVLxOmFuK5msZwzWZTzKVgHPZLCi5LoDTH4FXl2YUQYg7J3yRvCITGJ/4lO2h
ODRSKqTIGIjUcq34+s4lwiV1t4RnkFA3KgcnVZ1w4GplSK3HIEwkjm0F44UrOaVG
T6gwWrnkvb+/BivCv6n5y0iKIJswNh3e657OBTaCmgMGB2/Ny5HWJXkYpJ62uvrK
e7oLp/hG7gMkySDTexaIGEl853WChU2s6XwKr5ZbmPOjtlj5dH9cHf7ENb4Gkdz4
Vd4aQ4MpY3CFpjkRqb669+Kkn2HxlUwDQQa8jn3Xun6LTAa7wc35CIc3omwO3+02
KaCWJeuuyMffIzyyqRpS5BRWkCBqaPz9+kkinfJjHYgN4jDWTkgV4nCS/D8enBXb
Xir/FLcBVILJeoy9IkB0WdD2xO7kgeKXcSKRxdrw/xv89c1Ih0CufzdxKLgnT+vM
plSknN6EXV2KGeKZKcOyaZdf/gESiICXH7LeD2hGFsn6xVoWPKpRezFv03YrGbyh
pezzwlfO2SHaYYw1ChMWKdyPCsuhjRwn7agbsUI274Zs4XNEh+2fPRkXgD80Xr25
`protect END_PROTECTED
