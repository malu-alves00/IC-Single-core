`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1GZTwl4Vmr4cOyV2URWQqu84Kai8jXsfa/DYOjOE6pltfeq0zd8agIa2kMwH+cMf
Qws6UuC2u7St0j2kSxYkp6PueIKX2vlZxtlAaMrjEZICOoCuyoXoPqU+Ey2IbNQj
Cu3Z+TDsyYVTcH7pf5IbKF/HKyffKXS7HaK+vG2b8fJkX9IlhigXyNI6QK1ZNDJf
a0Df9sooPzBhUu73iYUAGqvrHA68UEn21/iYY48fGUVqgVU9Nos5iywXeyAMJfgH
3OYDws7GUD4I/1BtfYYXi+U0lqlNs77K5Bcw0/0IrgiPKs0sh74ggy3UCICdyJWy
g+GnjQGGLA5+NGu8oBrYucGsfWu5Lyv46zepjLiDbX4o1c/BbKePVsCOM8GJY6gb
MFh9r20AffIDPN7c2V65yO6NGBF6p1l5v94mWz6QExSEtiHsye+TIUskzrXWJOYl
9FdCK2rSfQ3qSvZx1UDTvl/HbOTVKkt9xD3K8fYQJs3Nrdvz4nEJWr8pzM1E7/XE
YfFEHe1MxNUMup4rrH8hFLrgz+go+Cm6/2RfhDaL7sgSXgn8mhV9egJNCUOmC/1Q
ilGz/DlDjYcJalqdRqJTLND5JCLCYdu7CdZYdRp0DNv3odCQ3ZiZLWF/2QBV6Zgc
ofR1La8ZUbJHm7IXX+LF4jtzw84vXgnOkhVP12Bu8AUAmd9ZjpzMtzdsKAkhWaf+
WQWgSEsG74tfMP4WMK0AZXXJNMBfXgZ3xTuoY/UJo2B7EaQkt3Kc9X0fQykWc3f6
9xg758sgiH74ZBJIQKGP9SfefHARliMQT2ug4fLXc3De8sp/j5DxifjPdAqM2EBf
yE0KjGtl3sL5wRfICw0b85WGoeNT74Nu64/cFGsuKwwCqBm/d8djxdztu6QYtfeE
LGMhGtZsp05J07Za4vHxkacVI1bLkKxxE5KfNHhcl3ubNEFzQyT3nOy978CXIzWp
qRZf28UFFPjdu//iObYCNS+pDmNLfregxtPO1G0kXYm+LRWmDsDCNshCfHGvlCVQ
bm4mP0YZocrJ3hl/lk7SOL9tweLdY96aS6vRFPW550lo4sAnTCRmdcHbBdAATugL
locKD1AxgHWtaTX+hRswWHb8FSo5VirKoNCDWBuoVyemBZD7QtjJiZaGqgwc4cSq
NOgGNF4Dw2iiMwSmB7lbaiEsfgQ18tF1Dlqkz+lGIdi5mSzRbU6DohKJG2EjoOcr
idPAnHAwpLq9vlhpqZS50JPxFlAHiuqwVSdEokgquq0+7ST2pHN+6gbGmupRTj05
J7XDsOdkg+mUDMKtMcIl+rTOJbVXvxiE9yo+LEpXZleB3k8qXSoIHg+oZKVHQZ0s
ydRzFpyphVbjnS2/Qf/3nM8+1zIdLhJp7i0QRaFtexEXhtdqxgRS3UvYTgC2ixFS
osm3wUL81jatxoXFt2w98CBLvRLFqQHRfEZ1lsEBnZe72rpKYUMqgjoMk5ZL4O4m
eOYbdZuDaI05PCxWr95yxV8jblPSiX6wocF+IQzoboSK4ifwVhE1wK8cBIeD+ncV
td5rIq11+WAG/JIvVwvRwoNiRfZlMjKCRUDAS/nvLNoyB372w9MDz3zAzeY4PfDP
BMwYxld27bG4dwRgAB6gjNVh0dyg86sPAcjxstjVDFZcx1KDpZkwvX/rblGm5tSm
EuDII0V5q0xNSWNPjNWPsoRkMrFc7mipf+lXkLBCYHtFoiup4y2U6WQImrWN7hbo
Tl6qHGz3BT/Zthz9aaxASan2SAMzeU8eEnQ8ClnssfCqyAdxoSeam2BJjX3bNX4z
UnOM0kbO9TH63FqvR7/PCuVjdZr6GPVxXLIUH8+jkUUzJ0pOFx8zW9KR1zWhBG7H
q4FVR2M1be+IGyw+JMkgw9cCpRfeujYxyv8ktt441qyrX8yIo7YsKyx6hJ2KlDcC
PrbachHDD6X+M+zct/LROYIYm+p1EcTDXB0JCt+GHBkCE9m6KNeqLq0mKjfwgwgY
5VM2P5mPpG6PkFIxxinzUCjaBTsXUy2gRUoU50thBdYpuT3oBrEy7mxjdqGOF+5d
AASXHLHkwYXyKG9Um+m6CGWdxa4E7HOOz+q2T06EDM4Nm1NETnuhu858wzkYxZe6
ORkv/hXWNLGLxfbN37M9ohzIC5+5xsuBVnRVSnfcOX3nnH7TK8pYyWGuN7YbGU+8
/XOFayMI9jyBbVi0tMVbRYxsKHimYaVJohta+/lKpNUwjra6Z27Bh110ua5uaW3G
N1412QJvTI4utNZgJmk+qGHIu0k5UmYrq2zF2GXCT1k4ywlgStlCiZbElvgk6jha
4rk/XXH76P5Rn21LwkD6RKZ0jKPXq9lTR65Z64rUTZRSUZbPy1DBoDw9jbLI5YnA
WsCiHWcrcDkoNH06p/vacYUESyScDCPl2L3voG7mf8V0MOX6rilLDV/fpWNi5Ycp
Psoir7JZC9AvrUUKrIbOQjIrCFJju8UE2Npf6BXepOoGn+8uvZKl/al/FexVulaD
RfWbwP884y2fkn2X79KWvBb4e0pAKlL739HaeTtllUCQ6sI7KoneXihcDPB2qJhy
+MT1j/j4z0nwrDG2xyrEEMHiG1qQvOJsPPO9CJbo55NEsbt5436GTIZic06S4js7
pinY06JhOzF6djioy4xFqljplTZa/h3I2zYHvvl3OU+5Y4QW2+lglBsGCntDY4gH
DGvQPE7kHQWalXXxFO0/koTtMBbyWQMJwGjDjjyzZSOpeSID1hHQyhWFH6gpshvx
EUVzB03qWiMUSHKhb929et7oftjfodngTq/RRUrJoRUW5x0kjR7lf1SFlam2B8ox
zEu44dG1vqB3Rqbj69MWz/oYHsb3KuQzGPe201h4sFimy4OXfZSIECK7elBKQUzz
Um0XfaYmT6GJaxY3IGLLc0OFfRJ90+y69agH8sWdwnoCs2d6jDWvS7RSMByqzuw4
BO9///P4/+cJo6doXT4FSuR8Fui5Kne+jq1k1V3PO6G5A/4qCZALRuOLAldY/n7u
YjckAHJ/e+X7A9ixd7fAL5a+jvCwdUdAMt5+spxIVwNvXZmV31Eaa2V90j9QpZ1+
b91X9OmyQLmYWjGCC9ZKCZKzsURFClhkd8B/5GE6VN9J5jeVBG98FeY5mEhB4Sa+
aQxmb4hF1tk5YKChxFNbVQUyhuzu+7xmd8+M91UWsXbm95Z+F29ZAKIFkGTA+Pvj
r71eP3KuoOxoygUUhqs6cpPT/6FRhzh+aEzyn0kkcFzbK2gVLM4aim42Y16/uG+2
o/7wSB7ucxdAGvXMRrNfK5XFCsMjbdO9771GYA2S9kzCDzKrAOIOUc/Amhl9w2t8
ej9zSgJlm1IulAMwUWvJhUSZz1RHA7ley/hNsHvDwx2el9VGHxu5X1uadcywqybt
uAqaYP4rrry3jRHuqQXth7ScnbYnofkxd4JnWXIVxfhZXycsKbxC+h+x/6F0lsD0
q/nW+pjrwYXSpOLdDB9e9LE1QvbPbXfIW3uzSjt0Q2dYsJJCpIU+JU2Yoy0nTUaL
`protect END_PROTECTED
