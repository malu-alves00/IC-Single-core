`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MOW4ryIzp/17q/XBkk0Dg+77NBLCyapFogohK6BoiEsLvlJIwcv/gd3AJlSlL6A5
+eLflEMDkywFJFJ1jnukt/UJpWmKHTQ5g3YM2NPwETsKWYUvoeSYy26mR1b90Bz/
vOGjvqsq6SQ/0XNVkwlkiL+Qgy8YKM5aSmdt7YhTnvNl4ZlA+zMLSKuqJSeUO4tu
73LVQQKRrVvZCOL3Z5881ndYZSxESXo5+k5NmvwcsLJfTTo6BvovSq5VEPL3Jbs+
I/QjFGvNbCYy2khi4Ra96C1NWFBgFkN3Hol7qS1o16Sq2+5ilyv8gVbhGid6FXst
YOiLJUAIs+PJCo8Nukn5Tayoerc6zUcXVfDFFOwR9L48D9qgu9QhEeIGCkxUVHk2
7WbEmrVcpFR+E5IoScLXnRVAfFC1HzKSndhCYctRdej5ZHWSKjJgRjHI7CQv8og7
imSyudkJvp5GiifGFqFzI5YQucbmfq/jGtHxUkIo0fw68t3UMhkh8z5lWTYVUNMo
PkOy+9JeZ15FoPtzJSWDPGaL12bMJnKXF/RxbyGfK02Bsvjvp9BdgPSemdTLYkkJ
VTK8cotF0eUs67WRo1j2d3KVASZC5AQhvQmHw4ZgI4xtP++vCr83Hb4VM8dZKuQa
1LCxhj4xJt4vZxP3eVYiREcundbB/bFpEUfuSgrMLmjjMbsIapvqpdGnaAiojbhT
05zXxWT+20VnkJOUlWV9EUAdadvpdMwTEh3bDDGEEAaAbnvRs2ZyRgIr4XdqbYO3
wUe2pmc9SxN2lDhAxhABKD5s+PcYsOfV3/VU/Y5LYvfggqp8bSm02TCzlvvzVrEr
zv/qNLDdnq5+IEo+ODYipUkiKVGKQnGqBHkilyc7LJmDikeEX9yXCXJ3JLENQb7S
+BDOiD0eb116u9BBPRIaLY8zAsWQ/GfREfKTQ0D6WslZ0aB7wGF/2fXmjej5nhHd
+DppYy6fzFxQIeAHKmdjJVtleAERwAeyQ8dqsU2qZElmDnDCn75d73vRZWvMBW+g
khzqHusA9junYO8zMSfm+oVlsf1HGIT5UWW8DxOSjHqW1AdSYBT7+VZxelpBRBio
WKucFXHI3+XJ/1fZhMICorxtH9hxLcgvZ9XjR6eDPYdT0XF/fMsbQLQmRqNMvZ0c
TdB5RlnY0h6w7k6fyBpIQylYg8nGFHMBbyxvXjQr9qJ8sSt38SwkaGTDF5nVz5yM
4FD4f7YFg1FlIzR3h0g9VHBxCnWc0eix0ELf4ABcCZn4LGRr07+UmKxZYbS9kPAJ
GpfubVYC9cZmyXVgP2N41sj1LHM2VWYqo2JNY9KqHgZ7QznzLV6G63fzbgoN8326
lJmdi1dMYblqSN6/vgURmuwLGSycW7x1J/5sGgU/6Act6a5Tl1ED/fCzQC61zub+
tyL5GHuTndCg3JaVU4KfHVxy/udif8vj61E1L3OC3bKw8JsBbQXgownNkrX0+29n
7Ygy/pl/WE49IDBcCErgxUO6lS9UPfZ74JaXqzQETaK6U0yDafl75yAHziVzLv7R
Ii4R2vuNpY+7SapT/pdbxZxH+cLfrXhGx9EvXaCUoqI8WL64aPIFUnF+VIAhGV2O
0rTlv92wu9m6wRS06aHZoSje0PC+EnWUggawK8OFaoMng9wjtmz7SttklL3pCjhM
HoNGMM41Wxc1DdC2swqw63QQBy+xT9oHNl0mWqwebBv2+QjbkLgCvd0l9LE88fMA
pO17DkM8s7VAKc53rrCCrTqh6TEiCcP/MVxZq+khQpbIPkuntZyiCGEOl0D3N3Go
mPXamx22URt8otAYqy6bc26DXim6JNh14V15Ccpq+BzjmPE1/bqhlRjfRjy5nCHD
IG8/dcAcsXGSvkAq21gRxLqt1o4pOoCPREz8MR/UUFL8pavoS0nTs5cZBFjafP+s
DCBeYOx+tRhifAnyX1jZdy2c5q5/nRhnXiMvz9PEyK56k6Ndwi2/piVFmHwUkqhd
8ctWP+ql1t0S931z+H9dwus0ld8NEUFonW8mNjTYMMqnSq/ze9uPhO63s6j/67bh
7NnKFbXm3I/XIP2UmNafxypE7wRKFbf2DmjLgw4K/ZKVoLg0BN3UmasKDki2TB30
S94saMA12mis0AYJ7KcjIQ3bLTawiUiNDG8VjBbWSSS3Lsr0kkLSe1944tqzkFix
MWmobDOhiAX+Fy6/YLcdpagkmfiRzeBXpJyEeirFsa8RKwOdb8SsSSRobg6Ou/Ly
1d0X8Sy7vcc1T0BcL6EHTeh14jck76zpxrZXaeGYiR3yxTJKxTDAs9qJ2DB2SppB
IaP91eM3Gb91NaYB2HoARHoz7XfON9UrYkJM2kqbgqPpGpmxMtLXWKyfVLRJfG7E
a8ZeV6WuHWfaWQ1lIAdkMOxQ7Se7mZoAyWCc7FJ6NK55eLR4Hyk9BZ9jZ3HifjGG
HPJ/FqOeDLhRhMB/Fwbm3E16SKqJwoz8HMgo9vSc7YG2yGxftc6UBSB9ttdKFI/x
ecW5T/4074Xbr9aHhtquTAO9A4Moc9QryyAJAIOHtMuv9EG31dNqK9paucaXAER5
bypMzusYBxmnD64aKTYMErj0LkaVMQrnjFGOYIAZtc+3K/QMtvS1Pdz1HYBQ7zcQ
C8c6Ptj9nZshVxxkexnpJCvKz8PUYGadfMbR2Ss2OYsAQd2t4vMX01V1R3VlYiNb
e3Jiz0eVgPLnNDGpoKD3oAYMc5edfStj3T015vLDXSYTKv0Zw3A7TdqEjLMhshiA
M866r7veBTk9x6O/m7uzh3BRUfs1bFsuKWd3wYe79GV9aesQfNiGfYHW3EKZn6dH
TqjK7n6TL5j6P5yz+9iBSoBrk4JOxHkbveLIBSh2g980s+FRy4FiKuaauSmVF1mS
w3evLevMtKZhSzgMCUcxttXPhiN8CSN+z9IsHfeaIfqcysVSJrQ5JqaYyk//z3Fa
tnJcxWunQpik1ZTeKKNXrmWmxKuoByV+V1MLDynYHPaqOWIx7JArfLmhvT2Q7hvR
rFkcFRjgzgeGhXspe5IlSkVxJ4vQGm01zv7U/laltWF1MQbTO0Rp4dic/2PgyVNV
KU7JAYjjXPMqFFK3Pn6HCGclbEk7DDNElkygcbfZ688XuYImnkcl5jilUFQtMDv9
M6bOHhJ/3CSvA+2gAvBN6ichfbkBrMDo3HIxYc2ZNY5Bl5xRml2o1HVs/tEAaCxS
QY3FLHGdxH8Lqqixec9d3PDKuIu3fRq1nFFlTh42qDsCyTp6RngK/PuKHmqGSxvc
jgCZM1WvOICKsWQJ/l2S/7kR6uZtM9sfpVFAtwWitk0GVzvz7JLe9w3TllmVzJGK
KnS+hIN5oLxxGpUc0CAh68VEodM+02oQKKIXZWn5GImHOBPqAMnxRMUuhbrvRAPO
ImCMrODWVPG9TiVzQZ/gUaC6ivC3JbDB4ooFSx7DyAw5kUFS/DIJ2XP2/OspCmIP
tsE1imRv7vdqgEpgdSku5jB7p6z3+jvhDJl8zAwGsh9bS0+v60RclXhVrhidlsup
BEZAMWVD9+bLyyyNdSXODuEYYZRHcMYnC0c5eZPIkui3BU4uTcBZIU4+cX6CQ8U9
/vRfuRjxGcd+TnWuvV5V9i230pFvCUNjWbtaH0wY810z33ofAVXnlTCR3sSTZKZ4
KkMFzLL7ggqz4dRwjqzbZWFZfkA5xhn5uZKga8oyz5gihyGKPb1RbgYgoVK4ywSg
qTccLAZvpleRyF1NY8fqBgQW8PtbE41a95zIUi/tdctBDLNh8npwkogOMQnNuVrg
JafSG49VOyBMdCMzoyQ3RW1G98CuEOjxSSQFAtJaA2B1ZaZBqZjNfizPN0O2kaTW
aY0m3dfRxFyNwDKVhjUcb0+P8YOHTQxckTTN4hmqzFIMk4USCa/4BErPsk2hj+sh
btB3a6XAiZPYrGNuVjZVCrp8q6xbbaUFRGz3VBpu7VN0uS9FK4Joc3vm7KKY+Xvb
8OscxtjhMN7hCB/NKb1W4HJZ9x6MBab6yFsePdGjdUmM1IM0/5DAu5Qulv5Vc1rv
N63Ue1IDiT/aJQVGCygo6kTP35VgO+dNKajLw9zQ0R4/1/ZTW/WmfnzVtxTplhFw
KV7N4ogh5QIDC4inLyOaFGJLGSGuNPyGbyUJvKNFan9pdOgqU2wdbRVt5hWhPmIK
53DATdwKtvjAbkLJ5HRVCGx36CbcO1bH1dkSuI1PTh3Oo9tXO6KOqS6ssC0asWB9
20dTBarEkCoj+Ii1+Y4DHXeoo+2b2ePyBk2CTSJGXR7vus1J0SbEBm/bUX2KSuDL
/tJJS48Et35zMcKa3c59jFAqlkFn+L7debVAT2qAizOd5FzWJgTyt2LUDE/up6Ei
VSx4CYbI+aqIN3EsCrK1OkQaquGRL1suaOusAaT07ZEs2M2fnZCQeeKRe+I7eGdi
jtZL5QtLo3/kZi1MCPImZS5aCKmY51lRkynFbMYonZvBPfde7P3m07EN8OHOFko5
rfTbO/zn1vbR6BiMIckh8VkMrtmfc5XWbDOWXHzEUPVABrtveCv8ei4CmUudy5YH
kinmaScNeFU3fEKASGrrIatmNtbMA1pnv5Sb1V64kU6GfE22DlxNwQqXSen6J6v8
/Mqd3N83sCWw4iVTAnT/KOMTDRaDgk25mMFw8+CMXJSvbOtg1hYWE9tkdnxJAIsE
aBFkYxi/9muLh6FlSng24pb0e16aarm84xpExfb4PkkaF71UYw/BfVx1rlagbwl+
eV6YbSlJIjHDRzMwQH+WxfMgz+KXVK5CBUcfpcN9K2paHkLVoSM3kJwIhi8OLn7F
iYWxdXP71OzE488xinquXN3FosEv0DfXdWMB0vfnjotQEr6zRU94WdqDkKP86ves
u6a6rJOuZnt1dkTtImjm6VH6MUJ3pyiPSkWhm38XPx7UMVhhqklrn97qHDUF2Y/I
Elr2TvwfTQgi9osxuEKlWKnstI7CiVqJpReX0Aozc0QlN349+qUi+UA1RtwRnhyf
BWk1Jpi06sz/jWGbmEUA9MiQkEem5wnx22Z8gxOLQpMMpzKSyoUPEzenaPfgGimv
djLGWdDl3p+EiD7qlP3F1f0HiOdds/7WrRkVN7X/XlwqsYTQ2Ok9AbVo01w5nqTY
DTwKbmjwobuJLtEOZSknU4yMO82KK6z9v83Cr0p/KPHL1czstCo/q4/oFYElRtm9
rPpwO0D1mwdrTq7Liqd3zn4rwf8LsTUPaerSa5Cv9FEhUqUwMT5Y85b2TqkTK7H7
F5cw8WpIb54gwuYFSF01DuB8w/8MbskHvwRCDUtHO04de/+6mvFwht6G/LiJAVnw
VWCylBtSiNnra1QAYpL6naH8+A2+tLiirveTZxt1KnysJ9+kzigdczYbjpD4MgYs
PfQuEKJRbJ9WSIKDHVkxUvFEj2WLtAg/TxqzryGMymen9BGd0eTCDepgNxM96lQT
/9iiSI4Rr8o/lTiiBYZAu6BE27hAIoJf5qAJHZHJroIZgIkzNSN49gENOvslaJE7
CpCvA6C4fXDa+5R8qZbwF5EDSlPKSQFHiYG4ZEq2LhW+3dSwpcj/U6GL8KD34JrT
yR61HLFSwQ1G1GpNxflszUVaRQRD6ETuueMa/5J/ptuAiy6QMHqomVoogbBforwA
u8cpWJb7GTkb1suGtBkYD8jMyri2hV1EpgsfaDifw1gKk3T/jRKCJPv+B9VYLMIZ
0wweuYwHJiNU4dBjH3IrmxxNVkYwE6VZOobqvt7CVytjPXQE0Le5P/n1jH8PLaSQ
roEHGQUP9DiIbwvI/V8Cp6WO8fCD13UUjtC8OoYTdDznNbm5I9siLuoj+U3RyRpA
CP0KLV307Kn0ywQrNTtX5iK2Slfu4cdKbmVn8/UcuJbb7qyODkit9wKKay9Wsmxy
25DiUG+YndNIuA+LV4EWmfMwxQtvoNfCOnlCLJOoUyMQvKNiSoXZP93bbiMB5WXO
Y4jOe+0uSCOnBm8yjPwGXu6efgfkNHDjL8tnFIRuj0H7FG5xsvcxeBxdcpJgpSZW
3nn4rInhql/WXzL9t8tRWEyK2sKktmCt4gTH72youapOcfAnWEmu4KI6SLSqZed6
cbY4bBnCRY4KJI/qRJm5gg03EfV1b7kkNSPz6cst3I45WKvZbuYArvYFJYBEKGz3
VbJvqScWV2vXHU8KqDAQvE6dltSUNCtQxMrzGjiQmn409zUG2uWU7jmdf044vDZC
1evjs+oW+vGHAm9N5p3/lBJYVaIOncYzWWlYOCfhCA78c6c5FtQKoBXAs9yUOcR4
w3cydg8LUh0YqADfsUlPqYSmJsp2D+jippN2r9+0u82o6MrRgaiVm+ijZSwOpMVy
3gJ1zYXlIIbymBuE+OjjEdgXcNgzYPY1QwWuzRhhCvSV0q/hd+YTnt6pEF+8uA/N
zmzkks9MFdYiWU0YhLqGT74QSln0TEpHI5SIGAwCOPOkT3M6O9NXRMQ50TdCpYuv
ZLJEqsVQzv+Amcp2N8YPON/FnHwvRxtHWRP6sEcydI8oKbFQXr2ANkSOz82qcdKV
+YiEjjzj0KAuBuN7O0b8F0uOuT5YRH/cDptlJy3X6lP/6GGNjnDwxqBWgJ10dksX
cK0j93/vZ2Eoe+BnpD7H+W8lKcqv1HeXXnbD9Q+bLI7Bcikya7f6bKlcZYSOVHpu
xWXmRSzbu+bXBJKlUCqD4SBkBo+i6x88aOVxjBu6mzpEPlHZ5DuOOMGZsIWW00WH
n+CZ7tSXQxAB37s5AFKsDlrgXJvFwntTnuYvJxwjdn6R8EqKt6GcbkTYsaKevl+I
GznpcpTEiewBzflo7NZ+QjP/w04YolX6Csy3okTPo3o7WVs9zmpcP8qLFIX8OoP8
dfgAnbgW1Ga90e+VxkuowckGBmahQfWxGxZZmu5C4EvSL7rT67NvcsSJEzlUAtIq
d6I0rRsxjiAXGVDM3WfQlS0oqDu7U+CBwFFGtjvi2PvBi41jqkiaWZlP71Ful2WN
1ndrd/DZhX9ZLOtutyRTH6oKrTIP4Dp3Ji+4BihHn98zEymjfelIxxT3ccZ6C4jb
LjsWhL8Wzl9aXKQamtMiLsOD1pg0QA+VQypIISmeJhvgtrM0YNArZ7k6aKUYJi1N
HhyPwjawd9flp5u4S2eKmT2+MpmsOBD0O2t5pVS72MHXSrkBfPaWMb7oy1rLQTnL
gUuY+QHwkluoLgGwdMoLBYzPy/J2+QKvJjebtixbkm47QvlqDKSNTTicEFy5hRd7
gmZvM/3imtJQzS4NyR2XpaMltYh0m3z7z566CXunttUUgwqSx459uRpjj8CT60lz
n5lpwWKuwXql5lIt9hlLzOGR1dCeZtBV+ipUMEQYamQHDqyf3e2Tp+XcJiRdc4wu
Pzhvk8YMUovyjF10rT/kb4Xm7uHR1q1z6HK0Ock1KNK53xynms2C1vfzrsuo+aXt
FiecT8ROshnVp/yECYv87OApwW5WML+Wu3NP55yEgyoi3Q362+e8dJxqprFJMSax
VOv5BZ6LnndVoFMas0KUrKKjxIl0XeVfA93eangeLmuITRecv7L6Z2Y9EDyYzYeH
/E5eHbZ2KNV/wtPxUQ+aZgoOQXxzCaZ6S7f8n5f2RPu6tDF+z+em+ElGZea0K1kT
7d5nuq+WPXpDh9dxtpzYZQBVfT75komEfjRaxpwoBsux1Pl9hxIKriobwrLtxbJS
vYwHaxnhK1ZZ4vl0+BkaIxQ3yRkeuuW7sreYObXL0rxpcpgcj0BPMtpL5wyI0zhC
a6B7Il+z2Ivbkga0Nu7mruakkJ/ULjyEoFK8730qxIG+JOwjEDJbFiK9grAgSFwe
TLWhmjSxplphJv4cPLZh2mqjTH4f00XMsgGn6Vw77LiJzEZuaUHf7YXYr1oMJSII
W8pLF2ALjqavZ9JJILzcvN8CTpE9zdaq1Etf/NWCquncNKUjptnOsz9hQdhXrRJC
OQhzldkB19Wgb8/xVFzV/rNb2NXu+YlrUF0kGy6jnxe8SNA9QqZXBhwrR+0nCFT8
NaPGLxhy/qqMFRgoXQnPa37N69RsC5ZBUtdYQ7xswVAT7L5gRImPZbnYG29WD6X7
XJQSV+803b7qJJ9KuU11dnJB9KEsDhd3olCL3vpQNMPZu8nq7/tQjGRQ8SXQzWUM
ZsOFb/cjtHXtljjuftXQpITh6sqRiNJSdVa/W/j+Cz2B9cfokBduw8APEPypEAdA
2hQBQKJ92d/xh8fUwaJn4bcz8BmgYYwkP73ln/I3DBGDmKjW/kCpic3L/SkRlMj4
AS05YnFa+3AHactS1wQnCBnZ+7vPyyyUuVsFxe2r3SMHsAuwm4mcqUcMF1VWppt2
tVFEZQQ4YuXXy8r9s74CXzAW7BepJKXXTEqa5yCW/LHQMUdXkEuy0OGyhMvi9Xo9
10QtYc8qQ57bD1+RS2Reb74nyDS83V59FzZ5q2Sh2gcT9xeMhsLdAj2GLZgc4K+O
1gDWGhGcN2juuoJ3OBCrvPtOwRhyOHKXr1lrcMvDWOxRuB32tckPLjDygnwnneVO
VBn4B3hMrvEUoHXBO+ckdzr5eld+g97BbR05nFeqFJAp6xeWoCFOT+9RuO69XSNX
ta+fUQgLKTpDwLOyFOzr6sj8dX9eHu3DHwnbyvZF592/8t19hDjORi1vc3h1epjx
7pyVYHlNArYLXL7UZykbHwgtPBqFBrrxZssxFVxerxZ9uojKPzvZ1MUmwBYVQetM
Yxskl2cJqfl31cUCBkZin9hRUxp2X6hl6fBWmOaAFm61nIrY/NC4OVJ1//RO+9ak
9OTtl1IhcSTV2oEHd7rP4B8PjxuctdO0RAFZQwTJ+9pw31flMLxqx4KnLaFRZV1C
9VLFZLevaNtEZUSslw1M/PcYsWLL+La2IoC2FqX1hIkwFqikLZOIgB4i7WSvAgOD
8nZ4aQ7LIcr9wv7A+VbGhiBIXShlXC0EvX19bc4s/F9SqNICBzctdPpUVWuLl/xI
PGVCEdB2GIM6vt4UzHV0J2fnnthRI4Op7W2nvzv4qpwHHOyDDXdcNfQF70rmTsVJ
DPvqCcfHlS3W2f28xFBiXDXWQza1GGZM7kp58FhI/jn9tc5jbV7InOYmxiGLbyy+
j+3ftRpbYfa8aZB27w/8abTCUltKajKwlfE2cVg4SDDNbjSMrGisaUqPT3XtvODg
xvXMzfQFsq/CWfa3hYDVzewCR1rp7+4tQh2bOjArMQKia2bsoB5JL7pX0Qs7IWa/
Fo1xz43Q5B6ZFWvWh+g8V/7zHZdyNKcgQa7zeWVrsOWgU5xi837hpg++F/U7xyn8
0l9GuFo5A+A/JMJ2evmE8bigwqMrLlxrAjvI4A3nBFlogcF8jZtV+5gy9keC5fws
Jg9Ct8D9lMW6PODDnnHjU/BdwuLGPGnzjlNTYpgk0Zro3pNvm1hoDp4mAtJQxMTh
cVDnTXhFEyXdEV5DkswpOTDGpo5DZ8Wu9LiIdgdXPZVsrLq2oNCrobmkA/2isLNP
IYwnVaR0G7yb24YYNExCmmub7MUakECBq5B/FAFhTjUwulwe+JpfWEsrEu1hLsZR
9v5PjxUPt7egazcEe+5RQ5N+4GcaY9Jv12M5C0dh8Y8fmCpx5TO0potMD2igpa4C
DAgQRjyBdA3THNZbkj0RgYCPg/Q5sbN0u+HKzBLxWyTzg+f3FwaCGjGduc033HmV
c67wwgn7lpmwXQko6QIKdJerSvprMgI4NhAffyHayXaJztOtvvbk4rmWlzRCfToy
qZfn5bI/1QyZ5X5dLhSvkahpJluqCXOhOCIeYlJ9kHrlhBoqOxph/Nud/yOBRvUG
3acWvd93zxqQGwzfYkTSYv/MpQFUtJRtbiYkC5cmri34ZUd+lond0HDOxXSjGBO2
SN3dKuMGQpk+E1fgDfFMBrsyBBRUX/BznK7TaRTr/6lFwZhXsc2zHZ5leyyQaYNO
/CcuRWRyaDVz5SWebqB/oyYe1miFbaI0tm0TRV6hgobLwMfIhzqTIUI8EORuoPTJ
ExaEhVHONsw4KrxLyM0gTXNKFChbwMqa9YY1nBeKSvMhsc/Vk+K+qTA3CAVtxdDH
v7i+QeMNZENbnIKm03NlA2THoJu3xK1qDQndankaIZAkZRPKCwkI0bU++C4UOC2F
+QSABL2oVvNr/IfXEB0fkp+FDEW0hMGxeODdvx5ZCyAdMLs0fuDT0U63XQHt9zci
+pMOXieAMwHDMiEyL5EiNY0JRQpBQGrwxpylIlzekG5i4Hyr9TKMdQtT/YiT+SAr
2dQBf9zidWXogYCAtmP8gU4d0Z66B6jDv25008wOdhrylvhGxMTc4R9tWjmQAgoP
UxAijRseRu7woC7H3IlEZ+JsYnq3sdLDcSzayNDYaXxCV4XMBLh/2dAGWCXJzVzi
rjTtnoWBPUjLmdetI+xK2HEnSeeR95XganGJ/u3CgAGNbx8vHFLr2gpPHkr3sLtj
RI+fACKSp51nGB/RfttCu2D1VFNe4tSgUIAVfqsIp299x0RBlZnI4F4Hu/MVkolX
/MtcTX+2V19+S+ymSRPEY/g79+uwg8+nR4SsZioJgvR7UxPT7fhh4blUHUc7ekuc
DsTlNRDWWJQ7hAFuo+1yFZNVyu6M5krnptIvhGWxlYEZo2vqMhvxlqR3ujOzgn3s
lbfJqw0djEL6e82PL4/HRuxGDOb7O7CRvVSuSa8Ono7zQMQPprtxsBNiYVp76oO5
oqm6MTl4Rvr+iMXAksD1PzTHoJeEi8Wdckxxdi24wet77BElp6Xw3EJhh87RcOmk
acGh3TTtbB6EwtfP0hRpIpSWl6qKUha+Bx++xOOPZO359eC9CwxwkEsmZk7EFa0k
5LOK0tqmtH/b8Z+1wHLMW73tuWaFD/VN09jzphYPZaX8m0DA7iEXHmtliMiSiiXu
kCsMmFh9ocGF/mg+/MS/9BRcOIFTNhuYtxBQyX09Tv1ewNetjGG/7f1xhm4IbDCU
QQoskAIAhMkYAx4BQ5kKnf9IP6lhnDC6l6p42lG0MhbIqyWF73bD2SGlH3SrLfy6
eMPrQ8KCFlmKW07YXtJ/lZX7iXudd3GRTVDwyTzOzyzXwzUpJS3NrC+HPtTFeH1G
Q6iLorUoJpLbRft2By9m/oE5+9fZWZwZ81P/q/7Z+hVLldWHnWJRNnUsyYJiNjy6
S/TsSLJ+gU3x7W8Am62eZseNR5rB9a3bDllQJMFeWRFIhAnCmrtuaZxfQLhSaebm
B8WiNF8mmHSCo/aSnje+M4MTAo5ikB7AEyee1IiwAkv71o1RonCuAysQ8C5g2KY9
/P06y51AUBIu6WsEB77cRcLp1wsc+4djG/gzR0DczwCX9KSiQdHWI9T5DNHASC9+
rnjdx7QdDFG1TXmni3xOZQMttyxZEWGUi70MMU7XnL+ByWg/2OhbZQ38J2Nfoj1r
YX7OLQbuAZhPuTfRBGNX0Y4W3iY8dmzzSYBMhu8/5+eOa5rVt6xwnTc5vpXn1Xlu
FqjMb259eXeyFCYd6g2RdVe0UPnI3x9zQXu4dZF2PRcU3/09kk/72fUEIyp301Vq
6JnSikQzVnK9ylO//0GCh9NY+A4hhpsCB835SQ/BxD+aUxHj/LrjHJzZxf29Q7vQ
HRajKK6IpatvAMO3wxLcyr8LuCLyfOjjyqf0i901RaxWRyAdIJalRRcMgWpqOuib
bmrIrLHhReiTVdp/2lSWQOWOu8eCQCOmjR0iDagGFLKChwg994r9RAk7CY7RNef+
9VIRPASyTk3xqFM7Cc7MH1oCVoMffjBI4FNLS6lfYsWS1AEuxYS/Y9Dr0Z1XK4hU
bxSmSNwfHHMowCV5bGO05zhGwb7V4+f/yjzCAavm28Bl5sSdc1SZSxcQ3rEsqhTQ
/oEXk4MXvTUTidJXkvbe02uBjpJaehspJ8Gwb4zJxsOZLXKaFc+f6O3pMIEx+ORA
zQAT7c2NpZUgrb6ieKoS162LNSjyNDA3KISAuBU70K/9F6pKC7MAxO5vb9l2qD7r
H2yqr3649sl5w7LT5vX+MEeNb60U5Qze/ZFoKueXwONd/+dvBlrhE+sYYRH8/Fyq
rr7pTn8Ggc9E76rsYDPK7D7QRY378+w0ybnzdHmtEBJWmDqSS1IWsQGhitZU87OX
AHxp05MInFuaxTOHSv6fw8t7PtN4vPah1CK3wByEKsgyPUzmY0myiv256KTsaBuN
NX6TVeIxgDXTsp1vrthIPHzT853jd6gGkX9Ku73dDwPD0lGqaQKBdJNTxz6QTUgp
okQg9e123PPsBx2FLh4gup0ALB+SLZo586JUy1LYk8/JyzfUN0CF5epJ9gMXDzjG
eAIxK+6nVHBDWmzGyicXjzLmTFhQoJrILmyuCTPG8jSC8LzLZwYarEXE+urGrsP1
XG4aQVKPG9H1gj7xnnK9YFTdMfW+31SFccKDgSvTCwOKXCCrT/Fa9NRQGvl6CfIr
U7TEo6K16PAtr2Oy/oErIzVjI7057aUTyepyaPQtEGf3gw0isrxjrO5iSuhPps47
8OTrm6QR7ENoWAYG43dUsamDLFmwK6pHtKU+7eBTxApooG5e/voWpi54/z4pln/w
tFNJFyJUYDnRYiT3J8C5XeAa84AvZ4GT36T7HcGex9fovWLTkgLGodHXdz6iJJz5
rCfPDtk9wEYMyJmd1nAQGoeLaCma2IkjmwI7YOxqIL1MYdzUujt83xc6iccy/Orr
hoyiu1IRMS6MYoPItPrnnh223qyENkZLJkct+qpVDERSevnNjQVWFstBD+gE4jb5
fOgpoqkVs2u1nkW1smqjz8GWU9CagXXOPSqKWe/v8ixjBY/Sfhp+wB+8ePGPLNkW
UJZAq2lY4UW5IMOawuv764KnmxiBLN8oYC7m+J8LdR5WdpRdLFQlfccEQ9GCUmvO
xh99i7rlYVEuZTrl0a+K9aec+iczbhmG39Q3OtRvhG4EYh4tz7NZLR4+mY344MzP
MIWXv7yje/cUChacnG+DJYOIQf2f3JrbpXALwu4yFt3EqF0FtgxEn1quglQ9p2Ly
Q/RZQvn7pS+AeDuLh8BSiRxx6je1a0UkwsxEqwUHecEzgwviOgI/gDkw6g1OoTJX
Lj+5LuxYdnqIN1rd2Unl4OTsfIOT1DAeoXZ1aeOUEk529A97ivBNlxBevyc+gl2E
zXgG7wPiB+6tedIsVtJo1NEsMgnYgTw5GBo0/TfVwtzarms77LLaEcrocNcFOrBV
pVi9GmfFiJUCJ6rjOSytPx5MVO72ZmhqW+++EbHNSkb3Ymme0TQg2Uws6AMlIq8G
yjJPNT7syYJLr0QU6Wiyhl7XSaE3V1HF9yTwkhUIjiEn67CT2CtVi3fQBZOMjac4
P1QUgsud+CuDY8edhzQiCxHpQpJrLs6B2bFr19zZVIFXlGvSvYYXgmuQgec6N5FR
Zd/jWUAR0ZG2/ASdlvW/s7Ed2s9diOhvc7svQkCY0TfdSLg03Aq3JHwYfUyKxEfC
dTgpDBl+52cLX5z0CSKyWB4OhOeIDftdHCjY8i0urZZ81lvoMZTg2PUoaQOhEhKA
7rpIF9ZwYRiNSTrbe9wbIqBTU0tSOlJ4JChFnuSqGfv8uw04Dx9hhZbh+Dkw2SBg
zIBlQ6yGr1LVWhsmw7v6BfUAph74FoP+ghCXoZiI0la3awJF515nhUb8jcEy9lXW
L4860Nhw6psU/hlg5nDJJrJh9y1PVdc5m6p3TgC6n3qoNUeK8zU6ijkaPUg4mlTV
TdDEv/1yUnxsX4Pw+3eH2UhQuB8REymnfctHXqdQ/5tWf06iQNl+2jlLxfUp1jbx
JJvvlZQFHJgRuo9ykrkZw5qRiv4nWycR7sVuDtLVmcE/w5mbiULcYRE/UklN/I/y
mqyE+VxruZhpuF7N9lY7IMBZ8UOCWlivpaQJVQEYGMmVXzE/lOTTe1FaLmJwC0wY
cUrUvWrVTaitPH3crQcfvihEHJD3G0XmewFmL2cm9WvTW3egy387tSyW4ldOc3Fq
ihwe4Ea9iZkgciWAexRxmEr99eowVsF3acKAerkA4lO8hTkyVU9t40QzusduMSXw
pO+AOgtcP3Sx1MGcBF9TI6R8rh3+2SUqquoto6y/wBDBsr4fZubJLNDh2swMhCMa
HB+0flfg8f83QWgz7PjaEdRz4k6PpgmLFGnSBVBr3GVa7touV4/y6xBtBFIHY2tg
faRF4Sykf3M4IinBt4sLAa9Dh1in4sfHZ8LsMX4l6VTOc/MGiN1ypuThmOH8vtke
UBMjvXolRTLVqYuyFc84VU24+QfDazMjkqAFOgZS1Cp9FmL/qt0sKG1hYVCuTqum
uk8wBsdOZvOKxojH/a6txiKLhASElehnL+e82XaJpPRQeN623lZ3Be6pgi5tyUrV
S/l14nsZyGFjAlDn26KObntDZCDu/Vi4P3Hk67+OBCcnvqggd1n/+sEC01gCnL3t
x2t6LgD09iOTLxaqs5B7wQnzEymgScnYIhayFcwLRpOhccWo/Tm5ikE/388wuq8L
7NRiFxw/tR4Z9MvFJYAEhQ+Lse2v8kvkwCE61FOCDaFsC0fj3v/AseqxYAG+I5gD
G1H7IA77OlgP0Yj5EWkZRUdYHcJ+3Qt7OREyErSgcnnknkybWm3QPwYgsbZuUOg6
bim3+LPnCd1sWVORB2HCxeZKD/u+e5X6d2i8lezJpzGkD6VdMAbDSN5xKMn2QkLh
lUXYlY8vApz+fA3dI3K5mcrfxIU3OoWV9mYDXOuHdZ1fIp+AyQxk9c/COgpXiELD
DLqEUenUICX71fEG7KXJWf7nbDyYtjCG3A8I55EzFkQUfSQrWj6R8w+M9RrCV2kD
VJ9z34GBxZNocx0JZeR2Hr61f/TV5kSYPR02YYfaIekH8MnlJAW6Mhc4XW59sqkU
QGaqstlKo0VkpiPljPl1x9YmpiYxBNvd1e/ekdilKTfFJwuGueBu1iz4LXCeICMY
yAKM2KvM6w6Vr/KXDOz54b9POHC74dNUMR05Men2ibzdOTHVgwezcnGuQPyj4Rqh
yqtjnDlZ7DzbXwQc6IVNzjQT+lDk3TH8zrg4nUbfFLNMKV6XrAlWuVEzKuzzM7UM
clMdKvIn0kjkG8dhMGu21S629F+Ic1/seH5Qyj3LsAu5XPfm/K15en7NC4eSCDQH
QpGsc285ZB7z8Jpwhxrf+sv44ra7NwrN8gtGTsToQ/mZIMbdh0J4DZ63Yllyy3I4
GCOMx8RgD0dzvjs89UWrpBrJqpgAn++zz1GrOWN9/gCFxmoIPE217Bdpb0SELjMo
WMKL45aIbSMlx7Um5bs6MAR4ZCXecdl94Mqz1AyObtmjmEn3nWL8w/HK9GNhWMbh
28Ur3kOybtleRXhRkzyjdsXglKx8hp6WFbDUwZukpocdwcNSz8PIDFNshHlvFvsq
CglrfYZzPr8L4XonDETloGotu/dl7NnoyFsJa4di59xoEQ/4jVkry3avhU3Si/wN
rVTgO4ohRsmHSu//catk9k1CAPOjx4usV/itLGXOvPM=
`protect END_PROTECTED
