`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IpPI1+uq7E3Tz0aqntyE1cWhV5E+xS3SCzUCrvEnKsv8wNO5jj5GH4BwlyGADrJG
I03IX9AVy5Vd6Qa1qY7aXSqQ9l5bAohyF6ds5xy6M3GhZWF1Fyyva8jb+1roN7wP
+m2dNZpxLAvJ3CCaz+ritfWW95AsxEZNdLkp0Z6tz406qefaNSBQVXSZfqZkpf3s
rEIpGIqHiqygqL3b8xeOb5W9hoTsEP/nd8oZ7meWIVr/DpbehDyNFpHd81TXGoQp
GeaOAUNFEwdvhHWldgzr9Ri/wbscsv81RMshOSSO7SGNzJOwHB648j39Ina9RLWL
9MsDmexrzzcGpf6s4d2MGAyFlJ/+TeUeZcE0cWxLejwm8DkmCOUtC2nLFYTW32C6
yer0CWuoO3iUy2oRM4WFEvaeejD55gVOeKBSma8dgz/t2uzM8UTj4vHjTDwybTXS
lsegPsLLC/gIJ6OXpKV+G8yYaH34+6cBzfzT2SCt+BxuqEvflPHECR64/nCKO5HW
lcSNDMFlTU3HudEaiFTYREmw9rDDt5qW3T8D3xY/rH3XitxOy3P3wBriRNsmQypm
/+U/VGnOHbfIZS/Ly3B0R5rj9K12l8xTMPUn6tY/PrhMklAqMN9Rke2dK/c5UQQq
StzxYLjjMDilVaHqQ5zL41qsK93yoMGINtkxa3PwrReO9z0hbtdaAN4quhViBmob
kBcaV2cD3oKJU08YnCgqnJ9rmkIYNWddzojYljO1W1rV9bEyA4+nbZXQjrrOyq+1
i6shFCVY2HBLi08f/vrga//eEN4k8k2s9kxbYURaHC0YQlbVetqk6oekqNdUuajQ
J3WxGBCp5wKs8AftG+39fEBehB60lx3Ibi2uIt5PU8uLqd/emNea+ZMP2+HiHp50
xhikWsYyIIjHajazsoUHbN56ek8dC/XO6GweO7jjXapXJ+gV3wh3/54BT29pj5lK
rDzSoS6aEgGvClU+TyqKi9xzGufjhAdeTu3Kb8w/8++aEZ7T0xrLTp/eOXwh62+Z
DYNd1p5ooBzA8wncK0o2YlQR44auApRHXL+MmAEvM5AQTKDdlVjoNJgG54UmlTv1
y2DuRllt95vUv9JjphdaZesl3ufySeakZY9mNnUm54HZ2i1KFm8swxIV3Fhndf8G
SLCHSU88P/tl5dqTULxvojXogwZbfpj+V9CkcFiqoGfy3vULXejUn40VX35Zg617
T8gWgsChj1GZHFIahX0j73ufy+aw+YiC3yLopoNZaOdPzEwHOzgKkoFPIX185mIr
/L1WT+Zfr7w+8CkMhTbop4IWo31GilUBpZiHxLHXpGBK/WEye3UU18/WYEGnfrzD
RuirgL8DP0n6sqEOTTsylt7cO5wdOCLUp7hEfPVkJJmEfkWaMNLfkhuTh+1mF84y
p9x7qeJg7JtbIguE+fLOqQ==
`protect END_PROTECTED
