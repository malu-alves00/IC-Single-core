`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QO9AzNO4rVRzogeftdrKph0SqrO96QnJHz5M6nCgmDScqUNAxfJxHxA5kp+N0wP3
LxSz7F12jJK6grTtO6jO6JPLEBoEoBa71HU3h0W4fADNUOcXpUHkiA0Pz5pEwlG8
dWkbfU0FYvo2NtRQ38CjcSgURk/P/xGhrl1UmraSpUgZ1s6JUf++ZBY36Zv0qORs
0xYWdOUtcD3n5BLCSXujWpQDbwSAYm5/argLx9a4BUWZ9ugR4uqAmY5L8SHAgUTL
bzg+tO1r0N6FQLMw/qOKhmSCWIydrJG+4K5x+AKwFdc5WIz/CbCoXtdV+2BMcbwe
A8HF5typSFVMD+NhhA7wQxrkPYjmj1OT0im/PaqZExRi1OI3X+y4NzypscAZScRw
sZrZDZq1gI6tafw2yEOk613/sUz5l/Jt7QttFvdRMdR2CAEzl2E0lFe3rAh/8fPp
RAo9DV5ucOz+9QX6LE2poahlTW1RbXSyDJmnLGTW78/lIawztPCc0cqWah5k9VUV
ubphQkRtmxuEmB2bkG1Sr2L8drEQBGHP7JtTKbsLEFaCb6TRUejR3ivOQgj77sXh
maH9BrG+nNNC6uFloyMamNnyBkoVV/gVj6B3Ezk+Ose1Tmyow2ZWMQQ0x+sA4r6q
ub8WVgMup4yrKqnapSYDFqcvgmeU6PR8XoDKaB+HwLNESZZkxQ9XBlDGmYtSAicM
PxKiTFn8KMIx0S3axsP34aCjFIeiGgs0L06SoTIT6TpmLOEZH5wh1vAiKBv7X82S
yLAYstXA7vYYESDf4bzRmdI/j4lXBFXDVcJecPPlZq9g2XE8D5bpyzgbZRoq/o3r
EVpsIi7/s+ma9uAM9nmUHtFd7w0L74nE0G4h3fukbV9ATT2IvndqkidwFBUGLX+G
z7Wyu7Uob7iFGTW6zTenBHXhMXXE/FqfH6fBOYFTN/9D4GPl58btHQVoFfCKcTh4
M6QA/xSuWjCd4GrPqV6U94e12nHlLcNeDn2t6e4dOYejdv4eBL9JtQ7i7R0U3RkU
1kV95Rmm3LJXcckbfPVo3ZwdjL4lcSXZgjqsJKPVNBq3FX1pF7DUm5w/4856Qaiw
qqJcnDXik7To98bpoKtqkHRB54HTiI+4INJJ07/Nd+JaKOhPKkBYTVZaBeCjobVg
/dPAe8nTf4zGP8SvjN/b8cCr/7K9ADqNU1KfdGTs6DaPwI/W2UgJ7fB0wIywvuSM
dHCADi8A+QMAkgVYj27a6r1HkTgfysGqXmaGCMNXBnFeGTpDnz1kU4ii2/4RuTYo
61ji/bQXcQ4tIVlxOvTFnjYtKTxTN4TFpXVNpAzWHyc9Si8ICC/6gM5+RtXTJqnS
a8w1JlOnUcf1ucZiCQzMUV9G6pGp1rmvE2NmplyVpUq/6K29BzrpIKet898xsn3y
AD2ItJr+VtG9Jc3im7weY5Pt/IKjQ7Wt3JwPI2+6jxV8d4s87C4ibKVUnWPuUbe5
+ztdP+vtetr7f4panp1T3UN42IUsunAKcDCB2rDYvUWclXD/Sy8gjg/aDnS6Tw6p
N07KFyT9DsXDJ+ctRdw8Mg1lkpnu1kX/T+iO9BrF9tgsryXLd9VwbHEO0BI8tcpw
IcXwtk/9jngeFknZ5p2lgjeYAiM6NIcdLh7DW6RVSePnOaZ+KgsdWfKPgeS9pYET
oWMJkn+CyWpD2QKbWRhmO7gjnt456p0HZGcPjp+uIEuPag5wUcuv8gNlEy9vr+YJ
37DphT3hIuOoJeYNqCbRKcIre+RfTwaNkwkTSXP8J0HI4hLvgYDN+w5n1dHsh0Ap
UMsWSpjtNXSmNdihqp6f0GILKBX5hgag92s9LfVM1b21p8zWdo6fWJ0v0nyhWcja
nhab5kQL+VLJqFqqYkvLbB+ohPSzxckiLLrVmf+VYGL/fAnD1G1FdZLrZJ7/BTBx
oQkrbhfOjlUc2Gf9CDL19NQ0ozFeHE+b0IzTWgF0yKAQ1LKJt98oQ4dsCOk6aAMt
Q5cclibikhQLqT4Nbfp8199w06cJaXcJqCZL/sR466o9ypKFFVq5Wvf57ls/9QtA
w2PucUnxQ6HWb0tAv9YPzn6eV9DKfqHLepXEjksSrQStjac6BhnIc6vxFlM3/54/
K5mG8jbQ8OQRIWNl08XrtKD4ZSIgeZoiKuHz6lBxeui0CuB+SAcZV5a23SDoDbHN
6PvThz+MpJR/ZpElraq9lVjZZexSL5icxsafECP//3YKLLZ54uxz5UvZhcKT7b0u
bq3XH30YY6X+lF+KCHoZFaAirvfnnfzivQPnJwVloANZHy2eul1NXGSgZTVwXkzU
YG2zOEjZFImDA05u0fv95Ia8ulOoh1vV5vm7n8fpWgHKRwkIUJjIDt4KU4tn6DBZ
Q2FDfDCoBnTvLv1zwfhOYg+Z577/+FeNLGdIId9Ikud7PryjNR/77hFN4RhZluW7
+M5RCvTGnhXoVxvxGVK0a1Lcb0g40a6s3o9iCM36YrztiNHDjr6iDfC1GePF7Mcb
CcOsHz6SnbvhAyhaMFpcsn9OCcGXQ+02yfkRX5p2bxhp/hRM0v9FH0d7BUyHRAxI
P2q3WV9JOjzZGc+v1ANlGaC3cQRMC4dnTCf2hXNvs50=
`protect END_PROTECTED
