`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CCgP7wUdtRjPrnzsWtNkB2g0GiaSkijkIlu3HF+08Pv+R6Zdz75DthXNA9A8T8p9
Sbmt/AkMAkTd5GeiiPauLACdTd7hkVfpdGyGS/i0s8if9seud7jUvmI5/hm17PBw
9R9z5seD9WWRyEFviaU7Bo7f47yyZuvkjJDTrybf2KyT7dezOutoVP2oiZTcKkg9
gnjiutSizWGC5zCweAPITCoq7KcgeSJDvHjFAIWA6/F1AJYInsRIVcTKn2nau2wY
9EPWU866AHzclAqIcYHWQGSGplJDoEHdVfx3a2a+InAqK/fnYk8+e8I2HbXvvD1D
5Cu/ANDlnF9kamnJEViVyUBlRxy9+VaEGzlKPnJCjNvhatjlKkXqAwitqo/ug9Wh
whNhV03gfp6Gi7WotrwWRvpRwDW+viqXvj8GIHW+mkYF2fbEN+7BGP5Fc1EHVhop
gUrr1D98GGADYeKGwf6lBJVaPSmkiirY8OVm6XPfgVRmh6+QMJSGZ4cShpEdkL3F
/V0i/7tzvAdTZIAMBRt1HuYCeObNfZvhstvOMEYQc0JTnrKm2ihjWA4n1XjRrIiu
YgNCGIxMKmRS9g2124zy362tFzsMKWPB+xiWjakJgVaWh97u2RILXH0qCg3Atm3N
4FFr2Wv6N4bjxuWtveVtdmLTyxx6ckM+joT3OWjj9ftmPGHDmozbvmvD9SW3LPtz
QzX51WPy043HL4pVqQ76+xZnkBJMARVyuhSbwpPVF4DlNiVZ3VaN9zPk8Rws9zUq
QRZGUQ+K1yVhSaxsDIrApQ==
`protect END_PROTECTED
