`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JXw5XQavfgJt318RvLKdHDJANGJFfMNJ0h63IZPP97kSjpr+xiuh++BkxbnqQSHG
DyQRS6Sy75kuJKqRl+X9zoV7xi5rpSTnGr0SCqFGEXLdnvRh2xZDU07lZ9b9IdJ3
sIyNNgvy1gWlSua12oBpGa5vBhw1sUXFNgy5qXfkTXdPG4/jNsVNj6O6zpl8OiCw
hACIgWvjyj75FjxFoABhLKh9IuFmbDj0PWjZgAQnkQoxnGK0nUKXMAqNDfPXv1js
zTZrez+iJGuE25+eqoX6nc8isPihTbhnJD4vJ3P2fTW//zIJsLC4oXn+Z6kjDZW+
CvQItI71URwk5aBUpj/I+ZxwA8lF22RqDKLNLKuGUspRI84fcLYo1QefxuSZGD0B
`protect END_PROTECTED
