`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kfSM7bInEp54QWnchGCi3fLDDp3G+TJDm6ahHTBDndIFCTHxIf3h4T/cMmpmfNde
nVrUt2qfnAvR7Iui2Wg2dF//Ro+I+bHZkn2znRazRedWJYC/rt7qq6GLicHO6Lyh
vfhxYtUmEGP69UfBChZ8zF0cNb34YA/1iI+9Mo8MxT+8s8JK18KtmZckNvhOxqAb
cXuuZFA+luczQ2zKvZkPNLuVa+Nk0N2Ddziro81ugWiKJKeyrrsYpY0TqQNUxNrD
G+oHnPSMWdy//eDqOeUODdNypE7d97ldnAiU/cU4bxLsyfWj+YGaAZqYXwodvDEW
yxp1SXDfZerW7DsvGpw8KHRKoH5k4hVccaFy+QmL7BaSMpBowkA3vlUnPpQG1vKH
mQnhMXjHFbinb5Y2jPaR+SWgg4Z/06e4C6U7QCVM71s63pd3vTHmzil9dIEvAmAB
ACV7glHMEjDVdy+kWUl6zvj2TV4Y2DZEjqeBemRffkb5KPOS+LRbdK9A5Opt4nSC
YEjXuzO670ubcjT2QRVnYQ==
`protect END_PROTECTED
