`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Z/c1ewPd/NL/nE0qTvHGfm/+KGBgWn7b/Z/ak80MKEUa3pKyfiVp8HRLuYjVA3dd
P7Nf9eiSsObzQdJkZaDLPzS284gX+ubwM9rneNlFYZGIYjTdWxNvxZsT19N4jlyQ
6wyPdtooujziWNe/xV6Iv1aeeEeKvyX7uJiemb9i5f900i4zi7ZnWyyAH6aazReo
XUwtgFYmO4S2pJ6jEfeHwj/k/NqJxrLjGvo/7cHS7hlkxVpWfHJmBWnOgzuvhf34
FPd+QGW2TaKe9WLHpV4FwVmwKTK5JRrz1bYwtefgaibwRkdXLyB+OyOaL4xPXsQA
yJmgYMIS7e5LlOYIg0mXtiznSyNYTtgzMvntp6IQJ35rrQF2X5b345ySuCRtV2yJ
BkxWcec8pxJ0s6yZWd+SGoj31hj6fsaNqoPgqlMPAaNBVhRWjJOWLRR7YoGRPEVk
gM3jrn8ONvLFIEX93cJNM5ZJAqXLxjnz94UpyJ0ITI3J/oL7q2JygfpkNXJNLfOg
G7uHZuxNRy+fnKUwjpj0pYJ8SAaM7P1rbPNBI/V/1vby/TzUNbKxyl6s9AcTLSxc
m+Ac55RThPhpLHZIX0AtXp9YCgQ3EVtw4ntwAWvPFQSZlKlsZseUKJFB71CltA9o
K3tftFkf413LyJPQ/fiwyq90ULpw3hgT5sE8Bf0Ns0QrLNs0zBIBUEeGR4j19ngK
Uc1APwR2z3z7hbC4sGDTHbg78n5va8/Z5Ow3NUhQAeFmdgXDM1P9JLXY7HGNGUba
V5iZq/POJ2vSvNQ2IyMEoO+UkVZib6PiXm3UtgXeTUUdbrVjhHNo0cOGowz7jer6
7XNJLtSufcBbO9waoAPD9Q==
`protect END_PROTECTED
