`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
E094ywjtlE511Jw9JATeZlN4FqDFi4GDGxedDetDuaKdUxd7q8D7+iXpqqeUKsi2
MGDXn14iW880lQa9qQt0mAbTuz3u8yvTCanNW6+afFd1UdNnWB+jWgRSp7mYsKdT
srFs/jYe2xlpS5ElxkFglu1CTHAewC2n9z949xnmcX3S02l2DK6kit7z0keqOLw+
dWgfCBTJNYKB2ZN6jVCyX3kH7i/T3iH+qYy3824zLlbhXeHYrvaBQmS4z+R7aQvy
R16lW4qY//Y4gPcBr4dcP98LrzVYB17PX2Kh2DPwwnCelAYk9TZPrth4/MSg1MYQ
QfS1Uxlu9JimubEzn7qUeEh5aA9egCFHbt0KQlCRew9FOiF72BHzOTm7K36oti3W
CAeoIjmgz9YLRqU83vW0I4SoiVX3y8fqwCSG3fF5m/R6WXvQWUaLL4qsx+RBpC/m
oqmhrceCSqZzFRswHlwjP5dvK7QO4f2eh3jo/HK2VVdb4yF3aqNEOvepBpz9gcT4
IdBlw/FEfxAsH5RWdvR6vswHC3leCEQkagLCtqXqMEu92Yp22Xk+HIHFYQ/iLm29
vuml28b/63+a0yQtgqFyzEuVaYmP8vvzZsppsOJM2hLjGwqWeK6YAHr0ReT4qhP5
IkrczSjGWRTJyduTQeaUog8k6ynPe9X3/iBRDWkUUC3095VzcDEGKoxAhO3QiSEq
G33jDK65g2krNXHCva/Os8JrAv79gv7MWqbbej9TbTMTjwqNh7uw0lQObFQLJc7Q
/v+fVzQDxSU80NwLA14aEkeBkvgDjAvyieHrpgmXlWTftNg68BxIh4Pn1PkXDFQo
NShcbUwCAHqXW3QXOnDxTvqVnnoBeqjjV0HxtNl6hMfRm9P61io/gm7VrubQxelP
tSxk74rsF5MkeQqb+zCW2VvRp8mvT3eue3WoJQkUVUdpZBRNTwYrhLR7FuRAA489
MBBfP2Own1wH7hk0JyhzPrXhHnLgXeI5DUQnkuIpWD3+8n7JvZUeUV7FgCSpR4W1
5H04xwdWGMgpJj+ke7pLKnjL4OSd8+ByxcdjduV8AyaG3OmBgjW0ij74qwIHwXlu
0cDSKgLeMvxd3BuJiHK4ww==
`protect END_PROTECTED
