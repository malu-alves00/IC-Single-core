`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
u/uefeVPM1UfmDJDRvlrAbcIwvnjMd9hH1AbIsBvcSapFikF2c4714IeTEL1NUID
MzqOAIp40s27a+0uDNqZndCxRusGfibQQnX//4I7tAK+p58vBc4c0AhXGcbspIuo
4bMFoldWmQ1p0ds99SxnsBIMvdOU0NKkX70bfR/bLgwpR2QbYxBOVkmbLGgJwVE+
FzNJowaqRLHfQCaYxMZ3HUReQxN1A8eaRSzpH9naDOsR88z6oJH2Yii0IyB619M7
MYNzbPKdwSSliyLRkzIm7ZDbdRgbNgDNXThLdRImN60Uz2R8ejW3GEVkqbVF73oy
eTy4EzirOhCnRUt5MkJDDi8iRfEjGRnFSeuaS6df8FbZmK3JLumta7ZMR106z5pc
4mU8IPWMKkQqrK+SJLyxifty1o+jFBoiLGITpk1kULr7ZpNEsrTY+KqWtbCjx4p9
bx3T4hCz0t8rZ3m+bC2Y7fQsf8hvVDmH5OCDZsJe1V+0qt3Mlj51Pxvg7KM0BJAH
loMNviMLaM1HzeonrS/Gz7xD+8HfV/LvDya4Q+yefj8hSltD/wLBdgHJPoAG7hWd
E8Lr9yUjR3RKYn93oTOKGyXBFtJkO5VvtnNVcl+wCQ494RuPxGx0kEiXIGtRAyRe
9WBMg0FUR6LrOKxPILlC/KmFdQezcOOu3Huh2SuaEJW8uX3dlpPTfaS8AA7Lb+JJ
gHFJsFVAy1xBWAobV5gpDbIPBS3Ue540GK3WNNwGASHvsyifZo9XYligjzKyGsfr
IWmE/53HsdLfUfwZukSgzINWH51v6WH/IUnIILmLc1j1a6zNoGywtCa68b8s+DSU
3/QWXvBTpLTIxbUEr1LEW0l8om6wt+ZqqMnLKtwnOlJENyUb/0DZrfrwwQAnw6na
vkukfLgiC4ebhAQY6UfVfxicq97/BHQjtIpxwkmzIujo8hXZdAebmtJu63mDHVuq
87j4GQs26b0d9AF2m6bkphOlIawNKw9XsWEpzGvsRhKk1OkN8eg25WzFfEcVjhcy
URTG7/P7sNWSYnKCIgmyd7wT8B70LL3T2rGnMexzAoBAW8V0t5kaRbr3OCK7Ba0h
oJlo6TQ0OlAHrAfLDpDcaPbxF5eLtCGvc3LKvn+E8ppb6Ropi3lPnueitwa0M6qI
3sK3bGW38AxZwl9Z14tWhTPJuTBrRBIRTgKziiAh0pulq+7iIwFHAGbsHKlxgVek
Q4TDIlLC9HgpcTlqY+1YOEOfxLSZGzF2HKZ2IMvq0TN9pSthLbHGRRD+B9Fns+N9
Es2CMMIJyTDs+Aikg0ZmqbkUemoQjkj9h8EgJnJvqDvE9cd+B5miP4OX897uhLdQ
kDIbB8Hf4FsER+x6cJRQBmuZWlHsOAjGV152AOpvkee0+lymUU8OwYbvGPs/3tve
4JUZ+DHut6jneRZTjXJHmnHDpVwDwsRrp6P8OqZWv6bhZLt5rcn00YkvPmfjJ6B8
BwDadsMyQqXrmszm5nS6LbV+bmvq6jSxs3+hIsKYHwHusZ2wOQ3F3pf6eCmAc5+2
ONHiNWaBI4bJ7Ji9AgM1SAVLgUUw4ERpD/gqHcpDSSaoKySTC21xGCC5/9ExwI1b
Wo4y462euMzAS3ULKJgzFkK4/4eVBX+32YVvyRyiXK2WL8PubLH4q7+ABloqTf1c
N74EpyzVL9eWz3NQ4HEUFEHS21CZB+FmsqUEvDhmrViJg8ptCBd47BmulmM98620
Fd+oVbujJhEVbSnENNk+R5bfV44dFsG/giH9SmQrLvMAC0bSnFj+s6cr/Vlzj9BO
U0A5w65EYhDN+sZpXW/A9juNVCMrKK/nShhdU3NWA/JWCzksR4iVauApo1OdPwQH
Wjbo8exxpsAe4mPCl4+igV360plC4v6lxOVmRHGgVOAQmtuwMRAiS3D5rxqfEh4B
HEoiEcpuwxDVMEvlTwFIyM9RGq7gBo+fID/TaI5KkFVbA28Y4T4z8YAYixzj6dGl
0DaPs07QKpyZpO1sUd0kzy2D4KAPgL7JFENLjMnaN8GxKkPfNEo5spMJMoseef9p
EeSixZuZF+ERt2qqeDx7CgDWVuI3IexIRxzd+BXeDlIJ9eTbKYj3tefjbUw5A7ng
cZbe9CeGqw8ghxiSUjT5HP3bKptFNdrg6GzdDQIAJpw6Q7BIlbHLDqk5nplQRwvR
FfhVE2HkKHSF1i/rFTFheHIWvTfqyhMXf7++baNnRMO/kfMzE2wbYTHbHgjaipbV
H2ftQPqDbFnSGRJwoKHqHEmI3k5Qyuzv8cVZJkqdqmBj32s7Kvy0Zh2WhsDovJ8w
eNqYicMUiT+R3Ewf4StWL9gSqhLRq+ZBroAIipfx8id/Ewyrc4oGHXmdBnxLRErm
1lwphFQgwwEiKl6yb9zVj7hAPb3jR6CNJ/NdIQxKUSk0WuGdYDN5aS8c4HC6a5t9
TWXlsoD+barocO+dXzIJmZ1oXdxmopOdnjuKiMk/CDIH/9nfQwuNUsL2XpMwjinD
MIGB19Ud5W61CYnk6Rr2ixla8PEju9TXHIvQkZXBRZ59aIREAqVlv2TDM8CCozJ3
GRpOISpuzeRZc6AReU38A+21zr/O79GdEcVJTkZEK5/Klth9vZRJDTl8haJEn8J+
AKKAyz9z/0i1tm4aBB70Q8u2a/WHA9NF4xJ1DfM/WNRLa08BsUMFTFVN7+OkqIsF
SIS2JHGX5EeVMAGijcNavo1v7v3UnaTyoGaPmNOfbuP0qZMW7nwmP7ELUZiQKOeD
OO5QeRc85ytLSfTfH0f8vUfTcEWudyMEEqgMKh9k0gky1jvXG948HjSynz8prnMJ
7gpzTRc4DcrO36fyuN6fmG++mknJ5bZC2H7mpJPbREIvn8hm4AZBiVq24lR+tS9L
OQ4mFiXaJ7rKL4vX9TczHRIkeqyhKEXEoaMIMyBsZbDPdWMsoRpy+8jR4bSrDbqq
0xo0HecQPxYeA03qRi7VYsSYoYcKXxMHsO+IivmlDd+VLgGO1NxWnZJp3/ykTad+
Q3bDekr4iyy/hh6vex71DhMQgRp0blbd9pnfqi/1rlrsstsC2zGuOiQ+pHAWovAP
0vc1unKcuI16TvfNI3uOuBAaODcTBduoBjYhRD2l3iobOZVgR3srWSqSRvYccS7t
4gMqqEAKR/w+GeJhsM+BcX/uoOtl9Gx6AaKdWXpzwJcZ88ZZQ3aEGTREtOYBl7Dd
azD4CeOzCvlcX0IAsfshddUa7ZcYGsynMP+P/LMP4AWX6aMsrjQoW0diyXjKtSmV
TqoiX+QAoSCmLxMfIwgOfFnkCc7045glqyU/e1KQ2KVmf9R1vZj0Sj9O0CuYF2+y
zIMy0wsTkxQPp8YSh1DyEpKJjiMfo7PLPn/3RAYVIyZuIWlaPHS9FGttlmYSzOA7
WBmNIuUek/wDePFnJoLUQZ8otkXBgJaFaM+/DToDF+CAyF7g8PIdtvgx8l/3nLqJ
MBt1Qu4oBw4BJ8+k8IFTprGvVAMPb/AIRIAjh3gxo2dhpw84kqrZGq809UL2FS6L
/iiMcpnu91plvlY6YPGvJFJUusPD1gIa0f34018m+fGUTBWzr1JBj9dku0KdE/xm
fGpekyTI8y1xbhHG0ET5yuC3zxs9o3Z9xbpH4q/s7iW1nmNV9itQM0BVCTysR9Sw
LB2itHMWGynBIGDrF2kRyzXFUMhVHysl+OX8rr8J48nD/DeqjVBAKKhJpyfArfLj
0XRVVd6thZC/1JhwjeHgnFNXPZ6SpOUFWkIBJcrThl6ZPyQUjx1fvTjWr8BQQ9rg
Zu/lhp34NkkzYJMAiwSXuexLYIe7RDWTUeMlhJ8Y7eF8tyJZbANjtW5bLLqP1Z1F
/LJUwtPcM4Tl8m+mrkgM47PBiz8WLQLpNnxBgqWEOevOe/b63sYr/MQ6D9Sd6emc
SlM8IulAqaqjSdyR0yX4g3woiCl3n0KP7eHZoQFaryPck77Hz7KnpQiDznk+OC9K
TZkdJKItCGuxAjJ+dKf+ilC7XspGuC1+GUZiSnLR1duXhcm45MBlL+/kV+imMyNw
dOctpC/CVHv0an1tzjVm48BbAXfa4upKys7MFVGKoPsKQrE5QHfljTBBrWa85TRX
UrW8fEaOgVPH1usLm4aNX7on3BHLM9TOnIGIzIfZ3RvuTOwIiGYC8U+ejPg+Jaba
znmimZhn3B/qpzBlbjUX5BWXXzaPc62CDSagNC+7Z77GxbtqUfzLeysnw8iZc96x
kYaUAEPcm6EwpVrpsYYaGjmlj+YEENnKMQ5D9iCdOLKO3sgEB9Yp7URUodDTX+3i
psYfCGovWpGe5yh/hKD/ZMLGAyhDf1oTOHzGK9T+io2BjGEPLuECK8AEajssGPMS
ZludiYSgmeDmVnus8H1seXIAijlNdBDxpUykh21SaNyDI0/WTtdjmMUvFxWYd8+n
0+lnYIelT1I/h5/mWFCZ9YytyayH9/SroTsvC1KyCwu91xndQbYlyrBOzUDXhL0Q
p6POTVIjq5PimDUjpPQwjH3nmfY+jdNgqzfNFzMGdpwJ0ChBk+bqel9vbYL3EcKw
/Znu306rUxvOZzKLw3Jcazn5U2ZvZqFEKV0VbQD6fsIZNbAM5qJaIsd8j9yWABgd
9QhWETyvFCtPoLc03iJxdfi4FSbx85LJ4ncqA0uDn2sMsXDbhHejY4RfzYUWak+6
vQsd1HYC44v9kIc61U7+M9Hcq3L8BbO3goIx+9/pDPardnDGQcw4gvR5OP9t9lNP
zJhfM0kntzv7l8cbtTFRMYjrtz9LP1b7lumqv9LmR8jqd1LeuorpZRjdWacAva9i
cl7gICjO3mQ2Uck7C3nqzumvRzlsA/DSKFDB263akC23yjA5TRHm6WQ+x/G11tS8
v03XU8E76DBx/tq7nCI8p105Y9G7BWh7LwZBKnybg4npl2nu9JaOq57GxvJAdXM9
rX9/SUW8Bcdx2pG/v8LAZNtRfPn7RG1aAyGQBMz8Uc7qXGCT+Aak9/kcGP5pGyZy
zDbG7eunmMcxOkj+uvWgW/AMIlBnymFnXGQPjbv3Sm8CvEoUMvD4uvnDZGg7uVH8
uVvSSs2S9HFqVjEp06e8vXdM84pUOE/hxxYT2rD4uVLkytYvQypLrXTBv0tnIxVT
1xdlmWgCtSFdK6eJneYzQJtwGkqyKu4UzaWMXVioGrOs3tprOWh+Kw925fEKupAj
ABGOEUmxsQpL7paNQmdywm7CZkEswRWzZzqxH0/XltSlbcR90o+1YQEbG7k9VFTW
f6KfUfrQKAckQ+mzW7bptMOTZZziwA62K7u62sJ8oQHhSnZ9Qx21gCr6Mkvxi65G
XToujNerWu+mO21Us9ECwc8TEr8XZ4AgAcO7+9ER/NKHHsgjMV1YjTur5H4kj8v0
t3c26iH6cImGhIIjaY2WGc+0prW7/Qy1hKJWL5d14WXskiIwR5dYQWd8JCcLo1LW
47XquQSUWQYL1rKXcR3phBZfYJcwIMfr6qrk3+o1PKYESOfodWSCfhq6csXUpv/P
PMcPZKGUx2CINqJSmn+Uzsdkbf2dCzWu/n5nxVGVkgY+BAJqTmW2mAUzHJTYclEm
Ggi4mcEJ4nY8yirJzPv+57gpT0W4ZZiP9JaPiGneWcY1KQfSwMU3qw/iLpmAhiRs
bqkA66koS1OzyyT/dqhh3GX5+7UVS+Ps7uy9NQ3rRQm1B1CFh5eyrWTNTAyA/wS8
BHw3PPFtibNKzUXtG8kQ6o6kw+l6tNTiE+zxiYUE77jsl7FdsV8jG0qTZTHHSbXM
eNKigeizNAxYC7Rhy8H55xZfY5i7eOW/Mat/nrt0I2FD8PRr4hUUj/zgiqFEpkai
dNr2kn5YTsOljKvbq++ze5GAQAxMGu7SZJtB2VwaSLhqQYutEb3h9t8RkAXxo10G
jdWKnAFp+jTcfDatvVv+3dAdw6dGCEnbEoh7XZmasngg8PE89ylH8UBhYu5Xss1N
EtPZpLkX0qYCKSCYfhE/FSPex9mM00da5QonOAUbDbw1ucKTYuKP3HTPNSqNB5Fb
/mEzjIGCHPmykgFACNgKKESN4eT6k/TNyXVac66kqM+bar1LB4fo7V4eNrxsxvAY
EKvBc/ql2f0VGhCTr+pBn28vtF1Pf873T7YZYXx8+kEZdNa1On4mFccw80N38s2g
KmWll1tvIrSgVmMzsSIroD0O+kyCvnjEoJJ/8uhLdqmWZ7pp2/BwNr5hFskySdYW
9gH14B+utvM3M8+axw702vq4uIdoUYku50gS6yGYQng9+IDszkg2zscqnCeXj1RJ
1zDB2eMT9z1tiTlerCRMUwHGhBE5RBBbCmlgUnISoZ7/hlwiLe1rcbi1UJqjki/1
w8h13iQqrOcPw6cB3k0+xA==
`protect END_PROTECTED
