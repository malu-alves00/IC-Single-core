`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tmDZAH8+vAgfmu91X0kDyzNTGFCvyWMbTsFbm0SFQb0ZSdfA0pm9OW5Ho6G9otvO
TjCtTnOdUt/hBUn89MwzPuAt8IKR0q0fFqZ+xJxJt0VUE2Lp8aJDV0oyepLykZuf
Y8Bf4ayWijZP1pcoyiGpjRaq2QscEs80c8biKT7OTfUgKpoMWzBUQsv7XoksbbQp
Fv0/QWJ0QOR94mzok1TVd2x24uYAbk211/fXTIFKlFpbjRNuWHM/8qJSWKzosmx8
W6QgApYa/7U2kxuikyTSMFxNHahtvehrQu9Bc5gGnBPGzn0Ks5K1euYrTYSDg67s
RsE9yEZ04wuCfKrJnszKjztUbHkN7PxxutYt9xyx81GGeCBnHn5uNrrNRlBOOT01
/kmXWYfd4VuwSikIbAOdjmKc7JtEm39QX5cdpjMUnKYjoJVnMmRvV0XhexpxYEA8
2NEzZ89JvQwt/ogNb+DnpzyDgcKMDe/z8vlEOsa96oPquF0Ge+XJm/ra02aNd8So
m9mbCGGDEq5akmSsCFuS2amqgfB1BhKyjpp5qM4lfHTc9Dnve36lVXNUHTL/s2Zm
jYTd7qdHqgamnxKwI1NQiYFa1qRB4NVW0AWgeueZI5iAMYU1SgCcFf/SizgtEX6y
W91qwj4n3pWlTxYmIPKQIb4/KIxmXY/LEAlFXGbMhB4Ree85ltIbL1RxCRt81Brr
9J9xESSIM+dt0HDA4J6pfMHCsUSfq88/mhb4WDqkvMUeFbHTS2vWHWp/ndw+WAih
eVvoOK0rkKdcU/0S0xIibXY40uo/m3ddftbqT0v3BC7SIjI4Z08v8GTxFIuKBsqv
eI4Vf3Z368m6SYStOAJPaEQD2Y2IJPYoaoNNsZ4HLjO6yC1u2SCJbzoQYsMJ++9f
jg2InOG3pIK3Em/noU8myuFHB+dY0mM1Rxkv60ISQKw/DOabMQvlz4nKqhJ1xiS9
xZpZha3oa7B6KFP2ECfz9BbL3gprBL8Ox4WVEU/uuSCPQcbHk/cBfZx6beGQsUpa
8en98mLtVBM7Iuj3Laeg7wOBzqajWik0CT3j3sWnc70sUvAclv24bZGIcpa1Cbgl
ERKAKs5tAtycPxhmKITxsyle8Gzn984A34OcskaUeBZj9B7C7iNGUKZ7bUr8h6wm
JmjKmWZu8v0JNxvHd7gaSBQOknKvo1jTZBSXN7F/qFMrSeHlEHFWWl/OnZpNRk0J
OYm4x0MHZNwh2YNMxGQ6oQjSZouZNfRKOXcgrMKpriHObeJdfkkUltxYxmJB4aPF
ql5osGQvPQpy53p1t3ahKS//MCIIYtWa0SX021kfqTC0CBQmIn2nALDlMolxamLF
6rPaDWg0we4HWZFBpSdzDuKRf3ksAVLl2eIKUGcVJPO32VRjvihpDU7aXKQBsAHo
R6pqYkQWrF6ysTv7NdvFCCk+LBgH2kxcbdXozG+jpEPgwqvWJRLaDyzy3MMqRs0t
77eKB125WVf0jhyqFBMksgj1ujf8QXyx4xUe68QsZHRlTB/VpkyZAs0OwogTZfjL
`protect END_PROTECTED
