`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7YF8wg6wmlw7+JBJYcokYP11u7LDV7KryHjnrM7UaxrAf8Mhc134x9jsu/yaWZNV
m471cpArbcZY1FmUwi2Wgk8pE5KrKQNyknXWOCnT2EfGA6AGDlIbr7XQhIYkLjfd
lP9BqfK8RSzTrg6o2JOYRUi4/btVayO/B/V/MXTP4zecFugj+dpsBGYKUMWUg2nm
iEMDrs4rmhE37n+Idhb9qfQgRi7i68mdGamhiJ36RDW7XyqjOYfiM6xGu7/DwSFh
VOXmZiewIaiqxrV841ZQfNIPqmsKT7OmdBIV8EPgeRwxETOG/KOl5gSGwoWhwGYf
loq7FaDfRxW1/mU6qH/qM34lu7K/km6blopdG/me5hP+5G1cS5uzDXjU5UoLL/tP
UcILad2WHUz0LBZ+Cga35S35z4QD5P8qHLQiIU3dwvVjwb/UeK/mPkxpQyTrWIy8
UYvpweDWy061UoMM5ic6v7gd1VVpuxRLiSClE5KlkNNkOYSALiV+IzyO8FK5ZHun
kU5NVnJUv0GKCpYRZ9BZ0xIeo/W13nY9s1Q5pTXRVy8UjtKv+C9p2MiGttgd7/au
OoCS0yLKZEB0ktztXpTrLqoktuozFAjMUEmUuYMMCD7kdrbRyZufJzKIXHDMFQIb
y1nMFzLbvhSimZYSYHBepnkVG0U5aBJ2Umy6l/PA3QN009y+gjdm6C+LjE745d6/
dZebAQaBTrOnoPVjxMEVWVA+6Hisz0iZbFuQYa4q7qYOmntB/jKimrGfDSgaPUzq
l62eCtbGWL+CU3O5SgOoHvHQB9ISh3izepcHaMnQ8bE2uK8P2ayUFbdJF4LvNhyZ
DBiJrHcH+OqaXrY/YRkYIQHfdCz7cSpZBabyyIJmSJkggQtjMKn+jAGtD/PAFep2
ciYaSEKFMWMJjTCavlpk1PTNW9HEGeaonSV6TZhTbjaG2T9Wu/gl6HsXFichq0bO
uPfEvdb2RvN9VKVIjJerSBBhrDXxzD60ZeN9mFz0dgcR6FujrCnQtfxcph5MAFf4
4FqDQ+JwF6R8CKurP+wYQZm37Mky2h+vqgSR6QXU5gdWCzZjlv9QR7JF1FK6pC78
ByPkv13ePfqJcQZ+Uds7mr/tOvQAYXTh/1Evr8V+mwaA40Djg519PeDd1ynmjb8X
Pwk444uNLYsQmDdiCBOpX0WRhDxjmQrX/P3jNyjv9hC5s8XQogCBe4PwCCm+mNft
t0DF/DKS+IfkZlymwBy0ySzMS+NS9ETcElk5P3dIU+PpOEC4/gEC+Y2A+TDIqmU6
NXON+tl9554wYQ26q6taRMq4b72Hlqiywlq0Gqmc1bJes7QGIQq5XBFAPGLjUPkM
GRjbw6VbvRr6kj99efTlxdA/zo/NoPbonK2Si+kyiC66gwLGLdCg5v7E0O6UYVZl
1n5OC1T7Utyp52j0RhFAluKCZVrYPyZgIHMG6LdpG1xadh1ZgvF+y07IlfFIoFBi
8HU5+UtasvcG93g6ZyWCEWkI7USm2bwWBcATEzFH7mOGXcBY1OT6uOjI8BgRou0c
zc38z+8WnAuGn9yTVhFG+ednlzaebhgELk5YooVTkd8lTppEYeXH30yd80lxvit0
7tUCLkHiq+qJOePhLnDfH5JasQX8WGOmjTpNrgMPJ9HwPdnaPDqK/IuMMlxLTlPg
UbzJ6QFgz2EsuZrATc1ENWx2fxlLdlwwBdGwh/8L28cwNKgziOTLpljt8GI0uD8+
v0F8UXxXmG/Y/bScuXi+5vM2pgMp+/PZsc2WnqBe8oKMufhvmitmawqQCGRnQJaE
ZLV0p3aMATW+h4Ou1w+QYAKXQELoeJQBH7ikamt+5sN/0K4EpW3GwXM59pwEirbg
Lrxs//EIsNQg2qXQdY3UUjOlb3kLS8ZD8v2tJA2/gUAQKokc3TfTUGOOsabiZ7es
r9Wk+S+VcZSyyFJKQYvdGurX+P2kGpLoPdluLa+AmoWoFxY57G/7mT2+cWmEMe0M
7HCAhAE3NPnpUnhkR/DcCJJa3VnCuUGaEdU2D8ZTJ9aX5Ol/g39H3OphtLA122HQ
YEF96M5ARBQCwTbPRPywdHpXHzbdsjZLwzYaXV0Jt7JbCGa9SMkuCGLxCIqJHDaZ
IgKmePECqH/YRXdlyGrPX07tkGAgfTPozTH9u9aD2K2zUAZ5b4Zj37q9GHmlVb9H
9Cs3R37BbGcpfy/VU6hu4xGZSqpWsVkF53xwr2CdkH7dazMI/eQSsrlThzOwYovG
nWrPcewV7erng7KHlppgUIVjMDEBIJwe5mx1bkzQSQmIaL34eCOvmdI1uYXzCqT4
Wx2eUSVbqg3DvRdSTrZWnsW6y7WYFzhHaTIbzq0zjEvSVKKSVvT+wFibMDKy6spF
6fpL82ZOmu8eXeCObfLFIDgOPKcOqIK/xdKZ1cxVqBMFKtTBABuL+KqEJp9OY48y
6BJU5w4VWu9zsYhDIHMWJOz+kXC4jC+BKT7xAF8djEUuXLQPjfLWqptZ3a3TEKFw
VFBkVmIfM1hQ5wN+loo0YqUVhBrifxDCzkklaTbvGQjiYDoW5XHdoJbYOYhP4zj+
RgIK2q5ALfLLiVoVcHhrIh47wbHOVsrFlQ1KGZk13LxNwQTbK+KIVp0lsXG3d+VM
UQcQenr1rQFzfN6aiYB5IDzq1crjtg+H8yTEXkqWkwYXFR+RnfES51T3/VVgzW4x
cdR4udeEQiWrq5ypY4/4FlGVu737RHYE/q3qD4TX4WkoPxRDx5N7Za63nT3tVOpZ
pEls9HaY4AoE5jK46BDOQRW+EYUuNSh1crNK7UDt+xGDL++86H7EODsCqEQt9fbC
Rmar8Cn+2+uZeauUag/6tz3pX3+MCLE6tXjZWCMJSRB0IZfytN5MynQA5kHYR8Np
DEca1gqEBsl8aPQw6cyJSoDzKowDAEPtYAQf4Nz08kOVumQg8aKoXXbJM/SCpGsR
3kLN62R5HKL4cblj2y9UnKxq51KrJT7gCUE9mmeox4bOtMYDDCyXEPX6roc9z/px
AfXqE8qB9+RbIxL1eFeK8+kM4psuan80KlKvJbdXVlygTRY8EZOHlwEf4W31nokv
q7zVJSAQRu6sXcTi5bsIJzshp/Ks/JqIk7KWvxMB7dr3F/6PjJwpIX872oRweGr1
yZywwyh4NhM4b4tt9RUVnW6ZoVNYr5Sl3GQm6ff+5CeblbFWCe4HrMNU73HakfE3
t3QQp/9Q69c41uDc/YtQ0wrI5CkPeHsboVKPCrw1iDnuIGpBVjiyYgCsnkVHqKqO
lyseIAtTIOGsgdRpv9xIWrwZQPhMxWenJXIXxXlxScMpNJBKkNlEImrCZu0coUsK
KGagOOI819ZeANbb5M3NmSXLQu+HYZ6Z1T+kIbMe3/MPpFZ0tIRF2jhEI9LMvvDu
fNdE3kfHx4c8OWQE7D51GHtbMfA6+3LE2gZw0z/w2sUFVFkvnWMYajvA6ySRxPq8
R74kSJCNiYbO1nELuwg5RwPUgg/lME4emst9yVoTFxBrolg5RHsf63uRD7fMzllb
QQ9+Ig2A8oxYiAsUHzUD5orv62atOqx+6j6x8kWMhXhJbvGg7LYWiaW4/LfucFtk
QEuYylx7zAZKlYR9lTRrt1aojglKwYJHBJATNx1357E/1q7O8tSKnnne8/phCzLU
J3YGDl4dXyzgv3N3voHLgaj81VLvlkq7EW4rvy3SRMTMwLXWyNNKcXWURLJIC/s1
qKy7Hloic5F7GyB8Gec9ZK4629ZdXhzmeZEig/BVlFD7EBuG1zeVBb+QixMFJS5H
Yiot0+zdjKZfL7f3WTr4nBxvzpxx1pQuQ7ysmKtYab00/vvZugOfr/+cqwiHLnJh
U/sJSoHAJs4zF1YlIvsWvhBKKpRhId9O15x7dcUqIONgvqLB2UuZukDzeoUoF5TA
zkm/DYhH3NRq9m/UpyR1l3WNB38HiOdUotZupNAITQ6OztHdsbIJJUgR53NxF+RH
Yf39X6xqGUTzBtSP5ee59Stt8wQ+s7KD+T8kfrNfKnOOTwH67H+C2BBZWi/rRepl
5n7Kk0MXT7jo+CZUyFQ3YJhMGeW6TI1ct1KIEqH1jmOsAkpV8AG0BKmGdoPhoqbU
FMtVlYkkK0HaxQ27yiSDSyX8/DfNTKddMkqwRO4TeWdxKUVSeXINI3/E+mXuFGRR
EjgIcxxi8QG6IfO/59ijtJKgbimBm/AATXu+jm1T2z18HDQ0UCmvLjGZGZiAIWxw
Q/oVwhN1zEbM7zH/QMwm5RF6HYeWAnmv+Si7RHYdGhKsomkE8Zu9wEZMqz2JgGmk
qAF2QLS319zNcqSLk7w8HZ4nHwovNepl+MSbv27empIPoNtZSOe8ArECWX3HajHl
BDsi7Dnqokl38Oj0e8sziNnSTWAE4YzZgiAXyYi/iRBrWkxASP3OQoXVTtheHnjI
HvkAtxLt+Lk2VxJdHcVzOPW16j2t+IjQYNV94yK4Y2UTZndor2A5yVXp5UWUDqZu
qJU2m3NAZBP7opaBxKzaj2RlLeSho4ML9yV+1Yu0SGcsKnFR/GGXVjDZEBSoDBAK
CWBEB1b416nvnfTO1S3q4XftCp0Eg6JrfyHnwnrmeTQCKDBAHzyoD8/p0r28fqWF
WvxuT5BHEhs7augdLlZi8XP/GsjGOoApLyUKi6LJHxKhdmlIXDDs5yCWSJnYMS1H
32EkYrW/zurLXsF2+kUJV/cAvc52qJo78mGeBls9vYGkg0f9niHbLtHRg+oA44GC
Z36Her0Vw2sFRMdMMAuFEUDdbx7GvIQ3w/jrWHw3wP6xq3f/vSnaVTIgMlbhkFRY
XTM6V0m+GP+QKy1bSYKyChjTKHkD8eZs2YqMZAssqY44LdTYWio0OuxHZBjRFIEV
r4HErjcBXlpRTlUSy2Rx1HLxBBvIwjTL/T/0LD2QjpKTR0RleEmyOqhmu7dJJ18u
Lh3l5nb4zXPWHMSRJ/Ar3dQF2Bv+zHYOK1V3McgdgQEa0iWUA78tNhzHhfaRgyjQ
uhv2jhmO6rR3jvCc1Wuc950rkh5f7mvTmW1tDQLIvUhrCogq9215BgRxFX0JBe8/
FOqoGqKG8ohB4PMpVrT0jt7/x/RGRfA422KCJ3s2Tn+3p27GgngmdU8Ecv0AFRtL
vVVOlupsFs8OEft2ydgJfe3URKSAAb810sYFJ/7AFdxsLZ3kZKfxLh7kGbgZh/WU
0HVyd65vKoxfUsToDFrKJsra2Z68zzlDLwPEnGGJhklHET7EdAkCOug0UPxd56a8
f1eH7Bh8K7i1SMor6YcpV9KDkAwPzq6o7sA7EsDNc4Sm8iozVMnSu49tIBdt57GV
TZ5LJehBuPdR3mQBTW38uFtLLgiPNVH2rxKor6clWH4qflNLdEUhmBjn/+ZYJNGZ
EFj7xNc7+ChPE/XT/nPQM0dtkbf3GOnBA0EoPfRqbpTyj9cwzoXwis4zaPiGv7Mm
TP0DlZz//nuL2mHQdzrfrgc1E0LHitwPGRvMuHRhpvtrbnxuTRkooA0HGTmTzC+z
oAhmxztcOxtiYN2M1jgQ6d/SP/x5uKTqfqb/7wCj7GdnhQ6R6N9vynzlnP4JeSTO
u8J777ISv/Ga8gp0tZut6OXyXwJGL+1Ig2I85xkq/B6x000sM+EugpN9NwABrTDO
10R8F6DNX9NXwlMuIcAisZY8/JHPew0TC0z7L5FLtn+N20j2DmAaCWwKqf6loH66
yz7fyYviNJckhSi7CINaBB1gfJevnpCBZaYLld9qNtY3zUFNvbIXppN13RYA3uAJ
4H5P9efFlHG/vOOpsokmrifv2IXgbpc1xzUBbnAaICkLhjCXOHXc5W3Axvs8xYTS
hKOf3VBsRzvQZ9wCKd3DH3k39b0IuNFrDlc6aCtYDHOV0052XldDxbCuJgwtdxid
8wVieBN2Zn8ikI0j2eC7sIGGwZ3KFbhOgPhYzYEoFv/Kmh/6Be7hY8yopK34T0kr
c8G32QeVbMvzDNIH3dcMMArPDg8x4c7vek/mZ6frX5VQxEhGa7GA9BaKQRddn83S
bqA5t+WY85hCYOlO7PtRcJsZcMM1/Lkr8un0FrZxCL/AggA2t0Lg4HMBz3dor1Zz
6dUO9DbinGJUBlmcDovdM2dY4KYQyRR3kbOuJUDOMg9pCHVEZDIdPjZ98H2OGdQz
Sb2iy5ao8qNjQMMueaYVznmFWGV6TViRIBBqd3dr878DQDl11Ogo9M9W/sw/SLmu
jIqMTnHCaJUUg4ZkPJLg6xfdQ/Xtj0TShOR7viMjxokX+VwEnQbcPeLKUah0xDC+
iHPJS8gdf+pxHxPUAaKikzsTsmdof7TGiIymKaNF65FYItX9S4cd7Ku2uOtCq9aI
D/a7hZ/FvGxygJ9MWPsHohCaOECoZqMfWZ5depom57zA4T1wo622ifaRKLSeq+57
a4VrJD8wz5a2xT2pIXHYlEoWOrqbLF5Ur+NXRvhrVoulh6icR8ik0jQ87gYyfmYu
5PbwT1o9gBo22jJVxHD/Xw1IU/QBH5HWlK17PDyLKfe5aLoj0evQ18f6t6qQIQVR
GzUd76kQs1/2Bm38Xb5JEETUKyGUpzVfdc8Ebqer3MUrjtVqGpwAeXglG/Q80JOP
xkGqhaILarXyl1trfHt/gxyCkrT5z08NgO3V+3ZP68A9sljMz+Q/h7ZXv9CTWetD
I8fa5Gn8GPHsuFqxS3h/mLeRaj4uVDaNO8dAEE7ws6FJLPPm8jymhMfqscE7q6D7
D1sqi7+T+l0Jy2JTd6NgWdcw5uy7qfw1EfseFZl/WsdQEadjWGTMsIlzIJ+8ZLfB
yI/y5jRlcLW2At8Uagh1vY0WDoNcesDmgVrl8Pfgub8QfsuC/eGMXB6CzfgdU0MV
yvz3gwDhu+dsKmwjaAsWOYJWfbsjIO54Fs4a+dMxg7MBkt5NPWSHVYqhW2yyE30f
3rh1orTZzUl0UC6x2hz2NXi4ncGI1EtnaIy4X2jg1Cej2Mh0gXEc3+4gq5uCwkZs
p0cwSQaABlvIUbMnlENAPJ65ifd8G0w+rwREnw84BOcqiuQuYwUK/Lk1kP09xAhq
o+H8Amqw1LFNojsNgaTyyIEwoKh6FadWuyiBBhcEt2KUKt1Cgk8fAksKViTGW3g7
Em01sN4v+1wXVFlVlAw9KGDu0iL/ZixCaBc0b/0mEBMKNNa0Cox5W845ZjZyKJW9
fOTgRECE3CVpFTuEWKC+uUvB+zAfSLwkE2v2u/1TbzPy/UjYN3iXR8k/AdGd3KWm
Q5MR165kx+1Z4JG6ECqXMMzsRvmpV/L/hIu1cjJcmV0q5R6QdRAOMjLMKSWKlLcH
Mmx2ymbJ3806RLcg+jCArxNowa5uApzyIOaR7RXjkoaPQA6Zm8bxLKTGrhRd5wt/
O4WbsMFkTxyK77UyHfcnqoe4TFcH39GxfVboYp0XWhTseucJMpuCfsZX7YzWxnRM
mEABZ7GR/dxeKJ088U6pA3V4GjoYzOAhsA13Z5lLD3017xKNmejHCz58n77IUEIV
61U4KzuM8c31OUOkU0q22SfnGBpEDwRm27psHcemff8rxORW+3TKRZFH/xLqKK2z
9Yr2AIqp/EHLPBBnG3G9H85lwKZ6UYlURtFqs10ZowOuJBJelj5bbz1rSWbfm5iD
UFrXtFhzYID39ayvKRmqAUpfGvNyNZqgZVToUkYU+0EYno4qhlTmnwfmLSs0p1Dv
Nz05jpqo1SvRCRJvgjfPbt/X/soAa18XwznQdxciWmiVaTdA8QODeVufGihKQY2I
OMromAPobgQoyIqW0PhoekDn8R6HAIt63HW0Tdt9jzh0yzJir1A0of+uCkM5m2eZ
EC/Izb0cnFlAWUqEsFWXrHSUJLeiwfu7WY/YpLVKSu7HHxxd+1pOSG4FKqn04jqV
BVvOsa+GUIjq2cd9mwHfE+eTBA/ILeW9aTf2pb1ifbxv662ygqirTCoiJTIj64LA
NNMMchT40De+QZN4r8qNXnETrHiS01pVkxtVAevVDRd421tOF5GlJptu1NpbXcBg
9oZ3jwTNVhFthUjo++a8L0/Q8lmY3NaRv8eGbFrhABEV9+lOmcc9Jxpqu/jY2+70
gWX9SWCDrSZVAtca4krUEn2skUbQUSQMWOgLRtovfgFHF/X5QHLOES3trFommGzl
Nt3kev3m27cBpfAce4/hcqoMAKuMm99H67ZxgikV+wRJPPvUW0ZYRSHWHBd5kRZc
0tj8h70Pqpe2FVcJKtoPDknX2QgyurXWPpeqauX0XOblJ8t/FDKUQExkRs6Bbpdq
KqNFvdolwk8Z68YoGw06ahKBt2GoIjnnTI9PBNzd7I5qHZFT8/69nYe5Y+s2DZEp
cZeBIiwjf26/Wxf+fktv30kfKHycv+hSQY2WvILzVEUH6eb20garmvwbIjJ4Bgw4
pX8AtSOjLImk9U/ocPHk2kRyRfB1zofe0+k0tf9P6RL3YnVOLVLkBMHVipWhgOzx
GiRTik4IqoYjqOlX64cf4qPZH8sOHfWyr1mAUjC6R5t+xgg121D3xz2n91XUq5qw
icmeEuH2SWYUTmsU2dUsov8ggoUAe1Zp1rQz1FLAP6eDQugwUYlh6Qg7p2uhWidK
FJq1XA2YI+IhQpwpXxJavKbk6dk5Fhwl4Nl79P2j3udcm55Dg8nPlh98+KpXWx+K
JpR4/B5RM1a+GgTrCKp0NZqGZEv761wAps3QjymEB1L9cSBOHMCxTXa6jbSdUt3n
PvSgSNJ7FiMbqClxrciZc47DviqgE6vN3THACQdGrE/eF4EzIkEZ/mG1ldO9p2wE
omBpl/nIFGdSB7Y1/cnZlX6h+8Af8lRP16wdulP19+nJeYezHY/rfSWDf73WESpT
lHfTX4nE/foikED7uF185g0QCm5Hz1hNUMjGAmlvWa4Qye/S7wbE3wQgD3j3K58N
wTJ6AnhEJvyKUAE6Rvsa5n5ljbvFxscJ4ZoCT20+nE97E41kExA6v/53+4el34Ht
UyeMrCuI5DuhBm+bWk5xBV/5zaiLhHfoiF4LPufQWZhMcFpKIlrmPQTsnKeYXr0A
iB97KxEjMNJ2C47igyx92Flh3UBXpMijPpxE2zh9DHpGChMEBUaEZrmPrC6HAu3I
Q8kvHoHQ5uHLElqzAZ76XhRKsIu0PLoIA8V2baEyBp49PBfI4MF5X/lPNk6ZrZp2
p7yd5SjzEuMZy/qxf1+QPQyzXS6JqHT6GY+rfmx+2wosLhNNPTU9LNhgSnszZdDI
zLDK62U93wz9IYlN1l3bLlAgI4OoFQmpy2EuOVZRNo8B3xl+eYsl9teOtsyEUa/n
vhPF/74ha26JQVgXLIwtxUy1MJi6zesr4S0lHCpeoe86einF0F/jrb623QwT+gV1
qJdtm9OSxpoPceNFpP9DR3liAGj2TxBMEmX7shk9rD1IxaARetgHFaS2esa/pfAF
C0BTGlzeWztdp3GfCZzwCkKYexgUhdqMyxY3D5uUGK4D9SpaSqaJvC86DHmt02qF
hgwcUG/SwtnGpYT0kgNc5T1dlth4Zw5PUAM9uc6TvWOoX82a6rF/Ew6/xgyYlYfg
nMmfkSaeDZrP3CwkSR+HUXlTaIMfN8BEOUhnpZJYBuIQh710F1o1nfsd0L5ZSUJh
71fFFp9YAISVacYbmRHu5WHPddbV+UDMQJzprlH75GymWukEYNGJKReZAyfHS6k7
oj3FiqangIwLFoEfmGwpQfxibvrCnCoso6i0JPs2kCk80BAAP1H5MITyCLTSZX9f
gmi8HOueQgzo7/nQdsoDORYpcXhAdYCWTnuhXXBo05dhj5N6SPceuhgtNK2O1k3e
kNF4BXDCiutKkcN71UIW67dcd06J722Z182MHkhoD0Mtg/mW1VxzRBwOOSWl9D/V
fZbZjLjzoh1BwXggaBkq4EKUhnTjYPgwL2VpSX4BuUlbFaIOwMWSlNbpGupoiFJ8
2Rp+frFUo5xDUvTjgb90UTQZ035C01wFP+SBUuql/CXW1czr31Lco/jElbuLRsew
7SerqObV5LBy74YUsLRxPJbMy4OZTgJXB+ZafbDE/6FnRjeEsqpOiy+XSWntSYc9
hACBT6pbXiVfhFGrBf+eq3u2WAJp8e/pOwxp7iOGsi1z4H1MHzeG4XphYOFAcqu8
oikyFuZ2te86HJHk5Ciu0+dDtOPkkzTcqSqjNwBI8KDVsIRP7UI+tvL+b/zrvWTC
yONqFAXMYNp+fnVMiokZXX7pl5CfDLS6+GzNvhFlS6RJtPIJ9CpwVAWIn4v3qekq
YiAAC9CUAoOI+5NcHifIktvY0jpBGaPxtKcr8oSgKZsPNuiHW9XAJU6go1GQenkP
8xw4aKrXdnVhLwN0mqXx2dcXxE3sEGmBAoR0PZzUdqDfrOiMOqBREUt3MwDvx5p8
B44NUCd+g8emwOyTWv+RmZdB7h1rRRogKHVwC354kr3F8k/bTT1lytMn3iHxNl6f
/9PAMzvvGdZihRz9ZIMJN/ACsd8DXtOXukBOLf6MrMcZY0gWOkyMTVtUR+In2KgT
Q6ckTlrhp/WPMfG2D2hjqO8/llAlJLgxFMEHbZX2q5zQP/r2HWPdVTJ9IubIYekM
vY2S09AXhk0vBOi2n33BzgYpiIcoNktEGRgGWZ9BJes9JZRDvxr55f9Ig0ftz1Ul
cNKI0RBJ7E3CanBG1CYhnBHGqWvfHzZ16H4sSzOSmlZy4eOhqrNOyMxJtce8+lCa
Vu5W+Bo6x0xlSMGr446HsOh9o0kVlDazyFeRBsgFgzayygsXoqvTnxAYthpoFvZF
6PM7ltwIoa3/LG1JZXGt9BvizstdWrRPM7BXSCrxNDnxMFDy6D6N7PzN9XreX9k5
IWKxbDsFcUwfNJnc6Hc7da69Z/Usepzu+hdMqRXp8DlfRPdbh90RhTEMsf4wZZGW
wwnjMBzCULQjMSRyqVAU0zjJ2aU/Co7yLkpa6ww/wDGtghL2UCFAf1FKF48Ns8fS
GE/1DWozevqBgJUfM9tjSogKyQ3iEd9jV3lBWOHDZZc38LPXbiG91w1jXCkqUgJj
Mm0n2YKF+V5WXiaAK8w4R1u8xw2fsFsyhxdk4xFy5L7jYP/NpRbavstowuP2613e
zfUAZ352bi9E0Z79H6iegpqha97jqLr2BWgE0/rTOVmCdKH3c9QdYNBEF1YhmwtJ
BiIFMKcDHeug1GubAy0dqsRjor+YYB8l4xj6DjSmg87SB/B5Kaz3fkmnsDWfSut7
MUYvX8MCOFQzFK1rygVcQluzjYqBald5q/cjF8/tBEppLcCqqj5NKMJXMW2uA/Fh
w05kIQU2NFanABhMOrV+vNY70WGNzVRxP6bNEUXEFdfQHSdvgQc7W1d5s6KlQpXk
qj+MPE/7OJl5dnPPwkvrouAl5N09gLCswTgX3AyYnyGV/sBGwPd/eSptqjOYhG/c
C9dyRvEealaEFQucupIM4+tc/X5Jf6zzvte+DbJdxQjYUeM0OnFg7hDAXVwAbulB
Qz22P96SfxilWMSyf0onUp33gl9hRX/7In41GBfNzXpzrBim2VlAMPbB9WLcdUPu
Y/HJBkH/DfHAgDpFAimmeSI1y7oOWzxFaXaxupFwk/Aj0cErkZFiFhbF5rqDmSy7
INlAhRqMMWQDlZgwjRGh2i0nRH9umZCvTCXwd2G9uLbNSsIKNk5k8WPdk9s7NDi9
eYZKlZnSnOxArJKAXt3WERuvJ2Z3JEyifbu6JaFDqd0H7friJePKvgss/pz+SFu9
VFYIJhr68cxXHbc7BOfFK6uw/2iMQnPUT49v8X2C4V3RLU5Jbo2pfhkqhxg+vm98
4M6bQgbObxh7TAJDVQ6PZJIwshDluKCo58RI5JdF6Y8JPVZ0OTNS1nh/d3fYhYTK
/Oqm5P7Q4l30hP57txkuRrPe0vRlintl2IwPMPWIzMFpZ+dqNFtnKyF5w+zCrEL5
1mr0m6Alr62INxaqQyTjfqEZS45V+xAm4pEYGQBrl9OC2nW90UtY1LOxdg3f+H/F
wTmbRFpStTF6ZoB4sBFjRQVqbfugop6clEKBIqLGSo08jcJKIBEtvvYMCJWeQZDn
lzk4dkIOknhJb6c9F9uS8FlD8zgfesFQwMcB6PnX+jHt45vak+EcF1J7rvKYbJv/
F2Niiwd51MBS/4rmWenv1MSOIesB+gw9RRZWJhK//76rDIeQJWmupMbxuPctl2Xt
MZ7hs0W01DJ5BYgomrz0u+GOaqWHLXm36qwRFOhAUa2O2/ad93tnqbWCFeb/se/h
yiqkWs7Ke45BEnIX0riV6s1ZLovykIHxQ98dxwX/jW39tTR6Ku8AhZ7IgrV+34jX
B8ztI9bGDbx6ElPGXw3Spd8XCvocXAwG97eKeiNxZ2EdgpVa9guh+evybY/0SnlQ
X8b1+bTp07IKVvCTexPhqh7T1D77+pvGP4K4Sadfm2gDK8C5aDjtNMb/MEyED1DK
PK3NzcW4K46MFVbDahN++RDLuNsfZypZICP1wB978QAXeb0uBVwA15U2p/0cE9wd
ihAssXrTb8ODZ6rxJBOXY4q+Bwi34zaI8a9PfLYTFn43GBNroLtspwrp8ac0TgkF
kmH+OKpwkZOESx8lUk6p2WlBZ5j30P6IjfMygfjvHzMo0KQXEIBgH9MphoPvkNyy
ghWS9Ks6qX23SR7ZoB6AmiyI7n0ED6SWKKlwC0Ivhbc7mjf2pp2vIvDz8LzzM0b3
0+oE4dZ+IqFTzaXm6WELtv8yf+gl05/F8Eb2tED/UxqJ87eA7qr4zBcu6RPHUJPx
J5WgfiO+64tS56curav2nkjlVM5Or3lxAPg0sl0mcZMPKrFoABV/PkqMFVJfceZ0
mF4uaJqx1NwBJ41bZfFtwbfXJSH+m1zm+hGFVEHWg8BBGwuZ/g7NGf28zS+OlMgw
t9tfb2diKk2x+qpApdVD0ZDd1o0Hotsm3wJ6mW6LLlhnTw6ZTdY+NBXTf/yWe8u8
GgTkliHjmLDTj3jazBfdmkdBlONshzWc47FWU3BQh457sEyKtTZrflpy8Mh7Iq2l
RnJc/iNFw4M9TRwDIaoMCMRE3cTvqkwDY8jYC/wrSj+nkmVlAPQzXmMEwfIJ5D6i
snlkElWgJQg7OV+ptNbeQi0hTJ8jnJ4DB9C7WP6hOsYOg2AZDfk9TV3xExcaTwxU
ohOj3vlphd1S+y03nXeZuaTYeX6fP5o5Yor20TrfJGQ+/pgV5FAfkTz4lDBbnoQx
fJanLd0CxpFqDaAp4a+XWVGA/qlZ+3gdJ4UDOPfQKSRbj2T7PWFVo+EY6H8my2Nf
k/0S3x8SNf2dLOZAQYRG2nkdEBvdh1wcB9q/wM3t+YxEAHNdW9Y3dVlxOcUnRSvD
mvhrfd6vGk8AA4o9401HMHHQ/z6V0Xdz4qfjuITprhdH8LP1/NiI6djdNYKs9Jnn
L0NKbVSqopM7i4Dw6SHUDIE0tavEOC/H4x/VgeqSVY/VSe/sWkpvnQtAf+6vq5Fo
QbanYl/JvaXajP7Dmg8O5tpKM5NeKSEnBKMdAyzPoGpeXLdrgD+GsgSJVofSIGW9
umXCievkXwghdmofjXJwjI107w1kTAv/fYtbQQlL61p9bLsztnBbc9OnNnMkRNVQ
iT0bRRhx1tsVqGFDIHxOpC+mp1J6WVrGBbm1crsYKpIeu/popRS1lliQPTxMVgtU
4aMZcq3CWVATJDu/Sty/FlqGS8702HQlT8iQf6tQABg0MdMw04UFqd6ob22DlUR6
XI3dfEccfOj2XnXmjNvnJxKvuv8EuJkv8W3biOG9b0QWuuv4BG85EuFhgje7nZ9k
Af4wcUGbes9MgQ9l6PcqfL9+8UG8txpdWIXzP/k29CfKG3OI2EBpqbnQ2akLe63m
GY3sfpInHiBBI1knxodXAXQx2I3p+KiHVHaY7YffyzHCKgvD/HPSvBdoYzkejlor
MOHx4mqkdmhWCTX5wYvuBPnuSl6ECs2h+Wmxp8Hujs+aW8TXKwxHjdUSTscuseL+
q0XSAaB6ROXqdYYsDLaWaBU3S8FZ4Y/zCRn4Tt3RUQMK5XjHWUenBYDanA+pPwSt
6DuivK7gFmjS1WgbKy6jgyXL4qpRS4hUbRiySwJSkWEIKiQzH7Me4RsMCNw6Hdga
yz03YuYGwRKUzyy1jWUz4CcCFYgZWf/0nps6lMN6xNny/6hSGjA+yZ7MI+yy4QDd
ZLp7YBuAQ+pNF5uoPX3m2MajdzsanZPKAjOyBsCJIhL+XHbMCVRTI4gJP4Rz16g6
4VNLqZ6EEyXrDmd2ebuHroM9eCcpAc0DA6xzDn7TKRQV/XNmKb/wsSJM+DH7geNC
Jtu8h0MwK7SWPwpvE3xAJ8c+JHQRcnrw86o+h37/7N4deUVe8+Cl+F0C+msPBwW2
v9hZwxjNYFA3G/dORrkG1oT2qmRbU6Ruqxd4c+78Cb7efm63xcKgBu0ygobXhxC5
r3ip0hoPzmOOBp9H3/ECSKmHU1ALWTD/8FSkEfpe5sf7gnBVrnad1nGH7g13j+fh
9zJr93eSLfCMxDzzb0UAwDEZqSnFbh3oZwWkgW6RP+VVv//BhLCPaTwMNeFEH9P5
r3Ui5jsptIV7fZDVjDu17uS35QBjHDpbjjP7bSCKQa5Dtr1JKuH/+n5pYhMBbYUM
TkIj2D8lKLAxSRNSB+ZyO8LwsuS4cA0Zh/kSvsRu5FbMoNjAvaVOSS5IyYVYRmq2
9OAnP6bcLnrGsJ2WfsqSC+sy7ab5KDiior/OszZIoykylHWzUoW0ASNMhTlCr94x
j7iHcZE+Ef5G5oALGs4JNOZ/CjZTx3YeMWD/GyoMCFHBDZ6Uaz1hFSz0pbmuIG/V
u1/ExEpXdkcEDPhpxVDOH09ekl9Yl02Z+ZcidEABWbVsBjzXwUjrYeVhTPiJgmvt
ZaODLWAUO5FU5TMciVm6UECk4aq/ePRO/gqSkFA4Huo4/eR73IBO0JD/q5L+MreX
ZPlsH5/dl4QEaEzwKgOeijUFV2Z2x98g650ixq6MfCz/397m66MGtgPaAblYMW4o
gqKL6vbQzJh7TH4r1ZLOvn8mZd60R68bCXQ94+ALPYloBbit7QRu69UCxBUxJs4E
8Sk/xKeTonqs/yZATA4co+bn4ZX3qgtF6FBHSZAhTKOipgxsYsnqSapuJ8MtMXh9
6dZLoVjE/zxzkv0JOMPvn26tsC78Y2DM+rcRmo1+WOgQJPonYLB23gpWOqEJypV9
rZIxrP5mJcytrN/ip/ZkLhJM5SeNZpaM+WQkXwgVL4uzXOx+LAqxDmgYnCfgLVJl
pDeaE9T3K+tmGvtmpKeaRRwg1yhGH38DUagC7Aszk2m2gp8Ctg9fJLKyve3603B5
in/h8kv8B0/0a7uco8ML3+9wm2uRnNrMefRmvWUZ9+9tDF9ObAKq+bNiaMCNKk4Y
SZ2aTgoQVYW86lvyqETO1nRKoZq6Fyj2kLqYxD7w6YZJgXsAIlVDUQJqXEhorS/7
ne+CUOM/mm0fiBSwcpnJGRZOCCEOeHKQKwSGbDscspzR+pGevFSi1QMJOEphN/Df
6A0RmbaFEGkgcMaPRTWX3XJXqUbhDwxdbNeQ1mJmya1Hcbubv35jRRfPEgZL7OBe
0SvDRFlm+fCmoMMjpIFTLL0iQ/oTzL6oH9OtcRTL0XZgt5QmWtNuMWb3E16+LEcd
1e6zuhkWu5qTs0ug5EflAXZBNnBoEunSEu1NgKXLk/Xc18oiX98NQ1UOlCm6dKBv
n9nuzMx50Z6dcsJJ0SUCxyTmXBXG2kgT5NZexJEes/FHbK845iHP94w0ngDUlbtj
yQZ2qeh4Ux8a+GFYOq+D9nbdCaO/Ris0aFpD4/mhZLjRrpDmBNU9N9Y5NBQGwyNi
95Qy2q7AVBYIlw3ws/H/d8CbuAxX3HNzc5W+4A7gnCPxiwkTiK58f6xFleaDf3pc
gS7iPfF4+l+qG3DnZkmj1B3uCasVypEboHXUxTT5jj+Pvfg3t767A/luJnSjVJMl
U9Hq3IA10iUig6lKFwaVq0dPtk0/y/S2QyecERY7V5tD3L+zLhR0bQl6EjTAtVPR
zeni1+SBLvorlblyXSU99FW6qoIb3LsN6MIDx5zQDYDByyiTBO7OikA8r1gHRlTQ
WwCxHTer3zb738VGfYg4f+I+QlAjpwEZHUFb8dwg4zqLyKvdZephY0qBBfopOCGY
B41YpfqnOtBXKAZVaXsyQh+gdgDLcCTJcuevy1T53ro7Dr4LuDhs6OtALcyFpTUe
qmwK1Q9krUAc7cCvfazKRVw8AqUpDIFpKF8MJwqNpczXRuIlYMIHfb3l+AHy5z23
JQEuP4xpFXQWwKjBh8+IkwY5gSt3SEUg+tghsh8iU2zCPLON3pC6Z2lle6CZbFu8
Z1SxXAMEL8NSFiacOZHST8siFq6Sp2enhcbdgzxvbsX5Kgb2en+1rtqYyvYVTnNy
8AloGBrPRtEU8raa4U0rMMjSZMsP7gwE2pXPRgOiafUkGIlPhGlXCBqBhmR5Ggd5
i0OWa97Ya6x37BNEYphZbIaoIpUkX2KF0AMlfPNA21yfN3q6acoEZpMRHAzZvtcu
0Fotu0a4BVpzcOoEdN6YhnKWFWd5k09kUw7a8YyOaYRrFqDic53b98+Lpoo87lub
hPoRGDyjqMtk6KwmSlXf4GbshkxGowd8eo6re83JtzlYiseIoBLr5abxgGXHmDlc
9aBNWJplEByGXm+fAgRP2Bhyt5KQaalJlOMQ4V++OqhhcAfVnIbFcaDmKoVutyqx
MPG4A2l8RNV+wlB0nKgKIwpS2Q4nRGF7+aRh7sB3ot2+oe87HmrPm1uDCrzv/sqE
Asx2x5uqcJoIkD8QDS7NHtbXOkCHyOukAMIGv5dGeGywETiwYwOH6y3ARIcfqoQD
5ZoYWQvWEjmyXmMpc3mVnDiXrmtAaYup7774X7Ss0D+l6RrsxoI4wSDq15ZdwwoM
8ULbDHF3x54/iIXAUfK6qOAc+y229kQ7MbH/4WXcW6yDaF0AgQqk28huK1Oa/lmr
pjncd6f7d2ESf71yXB+xp+zHqvSABkZrogrPAPlBahpBVoMsDrQNgR+t+rRyzNkM
6cF7dSHSGS/okN53kpj95Y3L0nzyKV+4rwFJ4xzVu2+7o45ppY8+dh0NmkIW25Sa
GYu7MrLUXYffxVwSuXKHT/bFnI+V5MSVdd6jpBupx4jQZm+C1j17pvoyad4I/fwt
ki46KQ+ahIx0YO7drGMsuFACNPguo/jLN8T0zJAtnJiST1YZjyER423ozs/6b+TI
EX5T1mvNcgpj+oOX3Scc7t7Zf02V4lkEl8+YDR30/mj7+IOjr/Nq1vrMKYXra9wE
ZAZPFoQzN8YcwloidX3xHeOOIzmXYAHLHZYPBD9AelmaabS+hLp3h3I2Jizr8ne0
PG7FPG9zpMhoPh1+rw9uEm9xEQrRnNb2HilPbjBhWlhY7XqaCDACQabV2xhgZ6g6
wWR8rFxqKesBE7FRJJjTMX6z7iiJ8EWreQB5ZW1CLpoz+FIz2OjLa/UMoFsssT+o
4lLTpGEVtdzvgKWPrwzfq4ZKGDamgx3aXpNTZZlsmcEJN99w9ALA/ps6ZeBDx/2c
wzNdLBBexc0WH+JvAFgaUYohyIRZniTAdZHudpdTzQTuiFe46O7CL4/sSEHSByyh
9QjRB80P7MK9DfSkF8gp4o3p9AdqtNtllJo7y93PBWmjY/lqDxcRPcgwveLJP0n6
tNfNF1ZcGNBbojtyd9tG4jQkhc16vZShK+q1SEuvN8h3RXtzVT+0mcH47xlyTkdQ
lx6o1lhDDT2q2Rc0wMeViqLW0r9wLst8oL0MNKr5CH4TDiQhowvmkzCzuYWhezCm
LDlGJIHTw9ZB4JLpMXl38nKr3t8mtaQI91yHhi5XBt/iqMgii9eUtIUCtlTF5aiD
I/F2iEv5SvWogzh3rzj4bMgFOtYxiyEDPTQfsRsFaY1eXiv7N/ahsf0Yo16Me3s0
XadeiMSar+AvDTA78Nw8rQX7Jo7GjyvTjxUVTFRSEOMn8wtXD2/pRyV4eG+q9FDn
/CZupjKmbXj+eHQeYQURLpZSAPgAkAEUYA/Y83j+w/Tn/F1Uuit8R4Ig3ZKUzjJC
ShqlZFHq9Ri582zF1ZHRtDK58ejDFqpL1dogFNQIEgHCbVDV28lRWSPZcOaWMYtp
9kkDdRwfp7TsVA9glyXOwMiJnGfwRRuf+rB+FipY0sgPvtYE9iqdwj7Prl74ndkQ
9zZkNAHUvRYFYCaaktdcCHTH8l76pSxs7wPk61v6nXOrTEPhwykLSnpnktjkGHYO
lr0YJJCdALhMKuMXYgBDAD7CQMNCTv3XeaVCpXVBEvLxC/GRynPYWBVjFn2PkS88
W0Rjiegf3cWLxxAJ/vlG16ziTVq1/2X8qkYFVF3ed5Uk6jQrqKGb0yXb7yscCcL/
uadImEB8mEXI45QAIkq/QKxZd2px52bO/GYyWWXhGEKezsX6vWVe0xcOpyHUbxR2
iIM8+JweV1StpWmn12ehA44QQHoaM8lmzu641ui9FoVxzg7zq70KJgEX8patxPKT
PRbOHOc8ONpjjV57swmz1sO2h2tpu0PmeVDaxvS15dOXemjeKyvEgWCog2v9guNY
Ge0vJ/lhQ43KQZEAC6GnecLX+kGHvGYUG9bbxXO+109Zh5Ncf2svN+oP/fvPv3IK
fyeclKK3laWsYNxGbrNsoCODrbgq90yw25vsAhSwsTXir+kBUNa6ue/60LkHr1ne
o4EgatDuvvII6PbskP/5eKAr8Zh8GvSyAIiOHjd6MomNea+Dn3zaG+WNhmyyK/Vz
k4+OBqur0xX7Bn8dLZz6J3+dXe/Cr30RtTk18A5TXQ+5bKwBRPnViCIlKq4tJvLS
dfbXaDQId0VjLEU9HYG5wvHdAIIrG3vTItziKNRVzkmzID1ZOy8wlfz8eIgjbXkm
WCf3IPv3rpc3xVwYUwrUihKVqL2yDjAbKs4F2GMWY46JtWl1vZ7XawTzLY3Z8MCT
J4n+04+nMHyWd1xtuD62whLd+QoEjT6L58PR2BCkhSeEBjvjcyevtRS1A1q9j0Dm
+Fu55AVoAcoPyxx2t+YJnHlVxq44n/noMU8Iz7lFLzF7Yysbu4OtvPkyOIpk/bMo
LPIrMCe6zUr+M3o7JVfvsnHOuT9trgxHZ/lLNp5hN7ebzeO0lfoGWuQ8OxepCL7W
HCti4Gse0yL5nmrIG9SomxfTvVwY02hEo/Vsy7hiPg6N8k4HBXuuzuWr5BqF5lMM
K5rl2/IOU4DFGbQRmLZx3r4L8Qpp+reU/5xAKXG5+pgbSWvdsg3Yu6noqgQ9QLVV
n+GzjOOWv4n3Nq3UlvInEFx5Hbz8rWbPkc250qEd7leA7rD2HCR1Mb2Pjzc10JIL
tdz1ctcoYqx6YYufEpa8HGMgqHVaHiqBDswHaOJnoQjN7OSgA3LrKcViDLhI3Cpe
I6wFjxji6gf1MZeQSIyJljM9FI8ZgGQuhjzwYj95heqP9u00xHlmy2CkXCojlZX7
gHPk+AK7s7d2SAIi6+ueNVOIdB4W7z+bedpBvwwc2rltfmLisKHjgZ0rBGC2q86Z
v2tc4/lM8mLu0zfwRYuTdo2W+OSyYN9NIyRgiSldQIpnGiG4XFVfSRL3xtvCu1zK
ft9cYvHWapYjXuy8YWs6Q6IX6unCD/kldHtaZqMI/KlhloOMFhG6V/tVCekGqLyQ
pWnxu2vqX1UEDTOzoNaWvhy/F97DieZnK8DMVf1VPAbHxnfyaQ6EtWDJybDR/vAt
KfPhGu1/uIU/+XFe3vXMV4sM9iYfbmvPxE/WOYPrhtvjLbVmkx7A/CyICsEvYuAz
EJZWDs90AlnxYLp6bbjWZCfnCkkClaYJylQgu0yxuMtI2KTq9zStVdruuylSEiuC
WKHnJu3UdNmOFaNQGGBROgoEo+wWJLHflZH+EnyhCCUJM3D6+69SHoZcKtq9S5vJ
rd2yjLXTQ3r//GtgzKtpCiSXSHWSp53GWa9/pLYTZa93cJVji1JUhcHxGVMC5bfL
AW+ekEDWshnFsH+SR47RSR1wwKwJjvvvyfYw+RQPWBBos34pM6mDNxneobN+yJ/C
UlfKNCBToX2RqXh4NBmz1GmxM6hs2zzp141WtxUq0SiqfAxdHSIiQHcKx6w7g85p
N/KO1BqoxCXqFhna2+QiYFgueot/+Umfzls+9eFVRMQSKpCtpuE+g0kEdsubIPbl
LTksIfOqcZei+RL9oqTBerxe0IsRq2wcYCVKe7IxrhvA5ksQ7r65YAeqTroZsXtr
jDyMHSIj/tlZJcQrP/wcVAeIVggPWz08jtlH1hV386RysetUkk8Hp1aTveKsfR5z
mhA16ynAoJEHkqI8PvtqlqhUNWvSxpxj56gAjJOuOq7A8iOud2/HxfkSlWWu2qHM
v/+Dd4CCtE9V1qywsYH3ZD/E/x+Rg1LFb17Amvys0JxajiA5TRhKlIXPBDLTarfa
Jpc9cEKTeW7Q3SbbgmF0C0wM82ZUthnXImXMUgS7ZFXMdpYF8z011j+DjGHSPJqL
6kh7hfJeG+9CRQhokIezqQu7h8jdvSpFTAdrRfoflNQO8qa2JViEAJD+usVpRxWb
HBCEt1Qzrt1zz8lPEF15f6GA8YskMj1K+CWMlIWbJiXqZM30v8iWMKxfPpAESPvs
YyIGPUTiTk8cHt1buvWwfdnOjzbjpLFz1SgsJB1QmqWwrC61A+3+JLdl1373IuFv
6oWpWX2/XGD43W4FifKEGsEEuIrjFrGPyW2D7h/kwt4FELIXSS7AHKaF/BWrBVO/
ftG22O7WgrhogEGXdhZmgctWn7fnAn6gBTyqq5WpbjSzoC3cC4Hot2TLmOZsej5c
TTRtDhea4cVfjRhWaftTKhHtk8OUWDxlqySZmzw4APfBS/A8z3/nfar6qyvDxdr8
ItNM2vsZgOOh3/NQWGeIpXtzj4bHrLN3O6vQAyvNoxfsRg7ewwcyC3yi2Nmhz6KN
BzQ9TTqRVDX9cpHtik4PaypiK1cVpbhCulw3OQZFFTc7iS9fYQyYUXOlvn8pisQS
Nn37bV9puNYTHgY+U75GS0x2zY3HGYDoWPOMbZhQeAjBnoiaS03eY2vrUpyZkj/s
rzGOejDWLZlihYYx4P0tX73GxEXgeXkl3MYBjCGzOxMZNYtBuNbCYka/jVZC8Bcz
mAOtmsv4OSrKW0sVDFmLDtIwkHJ44E08+MN0OIEsx1QFaqMG+VwzsHv/iA2uYBiE
XneGKdEm6CLnDB+AwBqAmALjlcw7TECIHJDjJvo092+rlKvgGAEqj8q8GVKAJkMc
aerEjItJR0Oxjw2lED90jhnHCD35BIGg4xkceEqcaqrpAr1KxmlUfnAYR9Xk+AMC
mM0pIpy/+Nt7Pwaj7IZRpgLVdr+HldpjlZjs4v5UY7H6C5gAVTnP4jlx72N88PP4
LlsbA3Q5k1p2QSPzzohbiJ8KB/TmWvBDSiNM5preD5HjM5ZKMyEFM5l1InjS82jp
kmMvUedbbzXMm9d/5tJSJnWFlA39CieMuF4qzAEX9yDwr8lAqy72Se3+k/xQPyjx
HtW+ogt/ZaEbzZl976XimSITd2WHvf0aDkP2/PFzos4Mc+3Pt7OBg0yndiCFwUdT
e64S7mWn8bpycqFE+0P+KNcPEx1BMgVSZiCXzejesrVDAtZN8jHvbMBcNgEJftIJ
9cD2MI7FdgknlvkUAV50CwKiQKPka0u6HFwceWCobDBpIkgk+kjak/xLMWrEY9Qn
N40/5sVcguONs1UoO3/Rdd+ZSIyTzlo2whe+UFwm/GcippQQoFer+Iyvlw/DR5RZ
nilOGGIVb9lalpyBkAiDCfLfXaFuFQ4src+JX0CRvkh2J9cm7vSpQIn0yoTmtRSJ
GrJgxecvWYOmGDUmGVJkOQZ/AjFuSwdpbnRaZaQG12BE0rpYKAbeETzX4/yYz8XU
AEdeJI9VxXxVja3zrB9g+h1pVoSpfN+BaDp80Q1Si1BqSwqUBlEsk5Dd3SEJoB14
NOTzkHpOBXO17QiDZwZ6oLorq7gho9owrK9GsfoOHFdNzw+Lb8ZIp6s9EyzHixZb
3moDZmdSCyk1HGh2kg1cle4n8GUQx5cxQ9iOdjyHG9Si296jU1YdzyctqfDPk7XF
BbledJBICBtqGqkj5lmblX5gtQ5SrXEq9UB68CVbLKuriHuT7mlSOvb6haXWqhP/
bM4KkoN63n1chBHnkRuazMV3f5sQVAKjDwlTRjLMBhInC2Ls9Itg+MmrabGNRhSg
c6B7ShrZgJZh81OUJzTTuyBkr1QaBFu0Bl+TflJn6sicm9xXdHHh9GP3eI0vmsYD
5c1/DjMpyKbaqh6mN2bgOnAkwQjN6RyGalEIjf2ZRxirfJj0VnnP+1jZdbhNGqY/
qbHr1cK/IGzbhha0MNpE/bzs2XUeT9dp3YHwWS8UBHaPIHwsu461N0Qt3rIBmrh3
yoFy/7ImrNrGr69siXCmJ0p0NMjA6y5dQSKOhAQLe1ZawWKh50P5HKsgRqlQ9XV/
caYEntSfxgosfOgT6VIGJJndx9Acx2AvlFoH+ZRX3Ph5DjdRebuQVqC/5/sYDdcp
jhmPEYGqPYGDZrcgoOcSWLPJdua5/N7nVrZm3/ayTH4wCmmOvblfrGJv8E/9U1IM
d9NNcpNVkjjbQ71unkX7x5k4RRzvsz3OgmsyzQ4AgSIB+wwF28+mUl1JHzu/Y/0d
Lp1bGW7fRR4qwM8j8I1gi3+y9i0afnro3g3Msx19SJ6lwTQnSUnOyM9zn+vDmsBI
tZxb4iO5RAr4gII/Ge52JcdVxfq495bG28Bv3l557smKiz7VEEoSAeGmDwaKnO4y
MR9JjtNj16tsMR+kW/lep0GvdIgJehXJ8LcQcsIH8CHx4MqUTNPXwQXXk3e2NjLE
sepZ9fdK36w+m0vLTLXdlmXY54NuEkyhnFkuQJ295Rgs5Nr23DxcMFTTUvn7cAOM
4/T/BfKDk7XL+tHHdIyyD7OkWVzBi12Qn43d8hUIf/M9TcGw0sp/JaFeLlYJFI1g
hfq06VSMjEDYpwcr+QHZ3KuS2ej4Fdmh/flOawZe3g6lkbfwEQJLs+VgJcD9FoYF
XSmUySafFXWneSHXfLVwMF+X7GZZA5SrtJZJUuNPQ4DcCzTD3TG4C6bT8CSMCtM4
9gYocsFoiUp8Y+av59pJtqY7bW5e3OT6BdWh/9/nikNQF6Cw1wTtshGVlrzT69Ap
4vNx8GG9fRqbVhiJ2FBD+lWoU9vlB5jcursVSWGKHWXRQ4u3+trSGGVMCBlmU4xc
VVewzSEOws7Tdft3N/DDhNVAXSVLE6Rru52YNdLUgzcp7dICce8L/BYQbyMmdFIM
sOvs3MN3YF7GZKOCUT//LG2IYlRcpFFXcWRlfsiFT71WoAktrv6GscqKbrhIu6W7
1TVCH5lsvBpXJ2zXn303lQeFVB1HKr0TILwd8lV8H77IsBKXdpILLatWziGKErif
+MnFxq9w6l8N+gRyar2m7P10EXlB7Db/fWWGuTjQi8tUa8ZChJdrt8ICfgFQlrlx
O8ImClEbuCtgcOfkWsEiY2hzieXDO9m/IkywHaFZuI18Wt++RucjjR+YxC9u/hyX
IWH6rrLtg0WSH0Y+dnLZ3ic8WgEFHEzzdTtDBCH0H/UFLC6S9+WrM5U9DPKzapEg
fIP3FBq6jQqlgwbolu7QLH2XfDaQsi7qluNmC0/EopozNE/wcM+8MPSUOa6qGk23
ir0nIJbmWrPxRs1VUqD4GtQJ06zGJeZA6aPQfZgTF+noPMet8sUrQ7jjwLneJn10
x8iG/+ujmsFJcbqkUtlLwaTbp2w714Inn31g1kGnIxTgqL9wHCVm8ev6Gl+m2znT
D7LEImCGPY2MUJp+3R4zdBcTfKBrMr0R2vSyXbN6rEToL3y7jvNvFLtPn9FJSOT0
SJAN+X2aFQCVrlWVj26sD+UTp4oWuDVBvof/ohLYWacp+rgWR48frXxTty61nCVT
rNYFf+M8Zb+ttbWVt3ZWBTb/mu61Argz38tnKdj58kTFCyF2y8nU6nCuVcNmhjRM
Ck+OYn7AsVfPIISLUZUc9yKVmqoC/gJJwnex9fF4QdughM8bZIE9yH290d84yUit
h8kA7AwEC8OLFuri2OZrmyXSG8X3doRmMH3Ub2Se6xL2Wc4s2mwCwkIEQU46XQ8l
dtCd+HDglrH7d+q11By1piy576Gh+xyfkxcP05WR4yonU0um7je1eIuDbaffMfBN
3ukMeMCR9NrsTn/aaYcaxvqWZHSbcPSBtmzZnlhqV8TAzbNLynfJsDId8P08wxVc
9LFboafUx95Hg+kFXJi1nZwo1oMGC3GoYSNUM8koOznbGRn5RKXFSQa35+8RRPl2
fv4QIesapmwEC7EiatJg6KKVZHeJU+DM+Y90Q5HPuc9eci0muuvW2yS/J5/2kwIb
86aUb9tf2c+/7MF/pCMutOsxNW2x5bjj+wL/0pTzbjaIPRNQI736HfOZwMrXhKNG
SmO3OLcWfQYBZn1UiqG3p3GAu6/qA85AyO3ZYuB5y/eoHU360tA2i8PdJDPZhaf7
LhE3MKks3dpIx8aJccu5PWAdYHLhA2RyBA3gqCYCjTY9Dfi8PVuRY4h/inK5sqdh
db/plyXrHM7lHeSckyrdy4m76/W2MTsjfWJQf+mSDnilcS0wdX6C3wKIV1qbZOO8
uv+y/K8jHHzHyN3yJ2i3PRUZLbZUTKSqqQGamAyv1R9FU9fqd1vX98GDY10tK2lC
MEqKG4ECGdHxwutiWdaFbIhEc+yvd97KD6C1RZqF7bCOnbLtAX/AwhaVEpPsqsGR
ppmEykqqYWbORVZQfQ9lD9CEjEuHyeVOIRinFsxsl1LrPV+AhCGbPl0PUe5BjwEy
VPNaJhqKtSLb5zcHONHjn3MdMTacEcPeSjESkWvso/MV4Wz0GyOTPpefYQyVK1qi
bW5ufOscrIAeoZIwnz7MDHtMs0P54L/YU2g77wHU3xPFZcFLzSa7tdMlaGpJDOGv
h3Oj+JvCJDl2kTCgAj6H2T2RsUDuINMv66OHTdDDzImnhYd8VvDUlgL1eZUpAalg
XFuIOP8v86g7lYg3CcZffyU5jkLrBK/eabBnFbcnhdomOV6U3VNw2rAghAEIgA7Q
HVkBKCrC2JQU+Bm8UQX99dv7BD3/cUfJdTKjPgRyan44yDgypnIJkCUjYZhBq8x6
GkshMxT4EUxE4UAZ7NOdPrpwdU7F+3X8UX4NsbT0hcESXBPrsvJHmJ66it15kbEt
BZaXEB17bZyLjW7youvRZisfZtGi1rrQkMV4sJVsGZotHIDoOVmxfSdmCs9pGPzt
b10i9+wXWzp0VL93WP3SkVEKC3vBBd8gsIUN4J2BLZ+/Em1hkUPGLlJrNlhp6PDz
clfrX6mKo8ta7ATxFvsX2KhX7XmaMkmV0eptgeQuwGfnHJFWVgPxNOsoJE1n9tnM
hhucp7VTp7c1kh53vIggvru7W4z+RGDrdv09K/Ff5IT9U5RuYJIKHA4vM/B05TTV
AiOsdMFi+BKtsSbT2Vuof166sV1ygA/wGfKGHSG6saXAviQjl9+fHqpbVypkSGo1
DqrL10DygHi9NgtxfcOhz/8TMe0JpQ/xnGxGmp/ERtLU1u0IEdIGmIxjqUHXfalj
IwAV/N+Jlu8PWUFPU/VlHU7yxPBIMmAcCA3DzpktfMtc+Tk8Uke2AzPbnsETxAMc
Ahj6TfOzD9I0YKShv9pmXhQduk0dN9y2DDGEBvkqJlu8bymJpd0a979JyNlatL+i
aFlrT0EHeIGF9ZBLuTPj1/gqCDeX1EqdtO9QKgrK2XhVZPMjiuT6v1LYnzk6a7JJ
kLIMT4q94JLk9P5fd+kEmpTdUmpo9zFRmVAloygWe0TBimveIXB6I8XhAlzgIiKC
jlUN2ym8kYLAty7JR7T/gYKiP11W4hm2WrnpOBnD66zlWevu4O5PEx59SbrOUjE6
8jPxvB3mGijqsFxagGT381p71asrBJ4KIdwT3MgZ0KFy5U2upsZUAuKT5cs1jT4f
K894Kv0ODzXtEHvjH9xKYhtwM73s7En2pYVDx7PqdNewb29Pt9XV6ByiMK6rCs86
mugApDTPhGlAJFqAir993yTI4FlLSjJ4f5S6Bu1K1+lRK2aPEdezNgD5SOj76/is
PaFPeUQHk4yYVR4uz93/Oh3bInhxIPqGTxTa8jimVrHDQXH8Haep7RaqIIl5e9aW
hjHmJIjo2G2MUq5dBC8oO8qEyEzN31JMeWLnAevw8JnKERWUn7KuVseY5oa3WYEQ
nDj/Y8oTo+3KMK5KvjAi7VO6yKkC1AQykcoQ9/dJTri9aJMafpNaHhv05AI7riZ1
jC2D88+p011tU2QJtGD5FhxUEUvtDJFiVk9ncVvklW+0qnoMWlSFMTuT5NVQ5I2/
BRcFn9R5r8cMF+k9Z4xzA0Q5KNqIuWIpPE5AvbG55PK3pjPiZMqk1C0mmwie+8YH
4BNtXu/F65jlJYXq/FYbKg5cQXT81RrJBWRvueNVKXqO9a+J12dZTGFkOOKXulko
bVY0XpeYbEdAmu80JAasCL/gBEec2Qy7vJ/vKbeH9HBud562egQcdg1TPK6c5TdK
oCZjPyR67PlLu98n4UZ1rqE8UknHjtZQObhaF85RnDMWTCVCF0M0uZ7RZ8UxAB3i
ossJM+Ed/DgbwdiHXEYipvofqNgnH3Fuw5QfhJRU8ELigzc/fNe7DFqF3FcGhAX2
Ob43CVhOYabOBZodxga5X9ePhYUuGs5YHlbwpes0XclTDbh8WZeEyfUXbZTAnqeT
Yv3vUFNL/wvvZ8snzi0g7Lze90zgHhY+g8EGkRDlFF2O9Gg8PFnVUcmQViy7DSfs
Xz0WcYxccvWwvV5FLDbkhShrXZek/8RUQ8CcP5nsJkSvHNDd6gEzQqUhM/1ZVI7q
mBELR33gQZh6bMntV4b7iL4Tftz7PA+ig5jYrvKBSgEa/MuObSIRxezOK4V9SxyP
l4O7i19EPyvkrCSv21O67A1hN3hwUnuQdafPHBegxJC1KGpOmWiEnsHIzoRgu3mH
NlDbFwPNVty6d0gbSrOX6XnMx3hdMWW+TFt1r9UTTMEqyqQl2/vGMTNqY+wHPOSB
lRG8apVI0Ci9qCMZxEBJluemN837vDTXzQRxlxPCTiDFZhL9KPrH9XA4XxB50CTR
h8XiGhcsWXYiR0VsWfC1iXhgII9EcY7TYpDBz4m2J3PX0DfxpbhA9rI70DJ1H4sA
eZEl6Lc+ebFwS9NONtwtNhxueH06JcTb5n9p1BPUO7bmLNX2ubbWFq5xRSQoBI4J
EeRja3/sIyhz19ssSyIUkMNLtR2wC1g7BYRGQUgiLg2Tgp465ATJnWfkLiHpWNf2
vCkYAU5c6ceTGQwB318zbi/xRddKZbSZaRDu0XpMHWAEuePcP9ZuCziHGgokQddK
nR/YQJEm514eHH73uPTMmANebtmaHHFMEtHdur0WUne6yGKG38V+EiQBkkYTBIoB
PI1KAKBa86oMYJ+tgx1hZnWNeyQpIRxVnn2RFO/JihjBFE98HDHvVVSiuEWXxoIl
fKQDVFhnR3F4HCCplkbn48K2BXN1phMKeoDmXL25xNMYQ18BbOHl1dWhYP151Cyj
8WqYfdJf1v6YBB5ISws5KZh7ILj4iFLgTl63IuaxES6V+GH+Jarc0URj6DEuDygY
GhlvzJX95SqYOd/CpXtws5U2MfAXz6YdelcEvU3LWuX7Ykaq7lR9iq7vITwK3nOs
OVLJr89Vcfsg97Xvx6gST/K36a2Hc50mhoplPFivznEKCIZTUoghEEVUGGjuygGD
85AnRr7CCRF/4OeoPKPPlumjpCNSyyxl1FzAY99hlwyhAHepjtcEwAy7CQjHwwN8
UbSa/6Ot5P0FbeAXgLLvu7fBlgeDpCPjdjyo4Zk8swX1t/ozN1iEyQEnhIYvPAYL
ys+ULP7AO0pkQuZjGXx2PCSgd8t/c13tIRio7XhYGVJWHSr21TFlQvRDAtAKVDJO
4JHwYgG0WRc8jVGvD4G5dl6Wiu0qVwIUVAqBfxuvsLw+cj5rB81nArFfvKWKLDS/
ECNeuXhJ5P1EAfV1cySzoZul+bm0zv4ZtxlXfbPZDlic54cnDu94H5iP1/CDHI6Q
xKhTNMPhO52KmqEDefCftLuINfvoBTsqVRDqPlxTFJ49Ex+RWjmcAci312Zaha8B
D3MK+7JY3TkDO7TXwbZZ4UISaTx8I1ZQmgZwbF01b3duKikzOK51vYrFxPT3s9nx
rljZI12DkoE0ZPWCYWQGltL98CTVZ9MZw0piTVLfaI/IeWrhE2Tc3JzujyEmW4yX
eZNOJeYXfDH8bJ315mihCF3XK4YGCBYjeZEsFW7gb8nEEQfbTJNvyF9DhCQOL4NX
5t4Xev9JVtlL7Y0pR1bmZ8R19UjugBm3oVmNZqYfnTI9yGJnv5CW8hvIH/IZNbhZ
wh2xcn63yOEtzUXuX0Pwwx3XND8iIX+oqZ3g3xZ6LTD1Qz6iXa1PJzBsOqT7PLj7
kLQc9bNj29UoBYPwOVz0W8SKpxN5w3bcolZpIdhUU+I3+ujq75tIRV/SIZQD3nAe
GESr8ENwfMyW80kgahsRdFn238aNr6QitAlnI8wxC6pomNxWDqGeYKvoQ3lOW2lA
KaHDf/O2z7N2KiP/e7eNv90rlOfAg7jzx1afwQBxM1PEi76dDKk/Ny32JMFAjL6O
61Z+cMId80FcZsAPLsWWCc6esFFFqfqSkWOtIurwMonEdJgxZwvPRpWWr1Csr/1d
vlRGtQmWIMP5vOVbWHs64XzNXy317iXzKSE6DwyWHVXxVIaUCJIth4TCwBOVL/Bt
vWzQdcUThZj2V9R66ANWVlX47+ITbQ4gaWm7VPtdpPqWSoBFSJnUIUdKg4G03jqi
kKXVaF7yI0n447VztJU0/NPWqnVSwD3niJEELnwQ2xt/ScbNKJUwv2rdeIZoRg2n
QFOEXl409MU4WtZZyMfw34MJbjbuuTDlJfVI0VCVSbNLkK/SbOzBOrGNxPpkOxlH
IH7EK3a9Wr0hHog7Dp8AroVJsX4Ya+WQu9TeN1iZiz65qnTYiX18ZlxYZYxh5VW8
ci98QF9hMlzHkHvYVTiM4E7GI4fagx3aHPgSxMQdXHS+CTwaaS6kzTYoH10f0rLg
qs91jd5w50M86Ls5qAlt8EFAx3Q+iydpQ7FaT8kE0IXVgHS593LE+nnpIDhOISn4
rq/pyBiHgf7Dagr4z/YqtT8zYFerea4jRdivl6wjzAO8ZifsrI3RQsYxqIskJO/b
iMAqT6G4Omw65DiNH5I4uyCkXNldOPP44XQSXTR6qgJf6wpUahnk1i4rU9hM449b
kMJqShI8KPdqGltRGfCFh86gFf6T3FDrhGXt6NmLHEhP4kvXxtXwrT9WFePYEZ5L
dD+qW8JqAW9V6AgO3NtMMbf9GyRLLj1khq8mqGxJXMeOpv6UQvV89wjq3A02+7iB
UrpoLvqkQP/Ce/hb7b9CKdXjWUe+T1gmj7UnSQrmzXllHTOJ/bwgBiT87D3pCrNf
SAgng2ZsCb0A2SgywgTRs4MWmRpTCPzVjvo57Ct9lUJkUoqOFwtY3OKp7fDX6wVC
Llir6sMVtL97m65gPDJyhQg/F3phDk2M6/e1Xqa8BkPkKbYc4kAQWrhN6BPTZqI8
9x/IePpLB/aoAFzdrkhOUVx7t/MejpzFTZUmKfLymfAur45jTk8r/RDMV0G0iEiN
dY+qOZLlsqsMN/QOJUWkigLVDZwYZmEiWpSNzyuTDZX+GMr+SBFVeno9JrxGuXoy
LnzGwDsA+KNrbIMnE96N5ptbct0q5b7eo2y+Ab3YBCxD81YoLnI6jkIve+LijFHI
8Zhk+6dmvI9Qo2aVh2OGNeQWbsOKAqau4Q6WGw3m41XM+IUn6dZHc/G7lX95TOXd
3S8/ES+8nKmLIH+fgK3Q16rmVU6HZ+z5PRhro1XQVTmQB6hnz4JR+aOmp2RSfm90
bv8yyAf8Zs4Sgv+RNDtNnJodwrensgBbr4yXEMPGL/wprtx5p6Ezr7QxN2NWo0aF
XV3NgbxLdZFIR2yV1V0heHc5vQR1xUeUHxCzoQfvwCgB2SGAfbglLnp3z98l9YEe
ivvMmCcL8mqfMBbervhw/cE6qyKxL11+vupEi1lpZGRdxeDMvtorhGEmLb5vbwk0
DTeUWBGPumbPIYiGTEc5UkwBlq27LX8MochP0jry+xHfqUaSNBjjqsbxcDy6k+UY
GDr2Iant8eCgTXm4PGym1MOEf1zmd/SfCHQgPatK4xGHaMjfZXgTFtk82D42pYvY
iDCLEHZKWYbCXS14Tl7oTcdquw/iff/Wx/hyQOgsaykN9ZEvKfAEwB84laP/mW7l
FjW7X5648IhSdP10FOM47ZjAle7icxh3F8tMhGRP6rbSDkrpwcw5bXXlKvU44xHg
WIgkmdRajmnR1TzZZ2QHJcFscLATx6CSmDDWMUAx0YDDHBkNMH+maSeMqfD2m5oF
qc470QeONzRWOKazeQYYV4u+KRCRkjOd/IZBIy+zF8mfv/YQ/15VXFz+0oMjxWrv
y4/3cjzNJAdjDvAmDHwlQLkLSoWPLknvXzYVNcqDXw9OC3NFrTPobnO+a7skUk/S
dntEJLYLIEG/Q5mjwG4XNsd2stdHvQyy9HWP9OkkOeVGC66HXdnXnMLL+SB31djZ
mE6O0iSg/iBjTZ2nCmfVyd7o9T5/0Kry3H8Of6GTXSY/P/AwHNB9H+AsFOmCcH8s
5EV+OJrehyl/PaoMAT0E2Iw01gx7J4E36f1gHqWIxJykkBRUQSwTe6TCQZ0ISJTY
91RPjY2SKhTKQ/0tm5oJe9NvUuIMC/ii0YkVoEVXfwm6WhXABTY4A+umwfHnQaoQ
aEz20VtMO0ONOJyeEZvAVCpI7NsdnLLwP0B412ghe2KI9q3PAi6bGoqNTdnaA6rY
ua9Tp1f1K36/aY4dR0/g29PctSBWah9A0KvqEh1cT8ebfwxrO7MThbtBRXaBfqZ3
JSTMxzcwzaQhdakfU6sSWxiJz7Pdl5wYgLcw6jAtTLCoUDMPSm8dCbz/odx7G4Yn
QBshVblfQvSZELqjmuzu2ASn7ltT6uHzfY/uK5Cz0Mhw6mR+imrVUakmmcxXOw02
qSz6CqVOGdirIinBuynmflXpdVBd+UFLOHsZHlGoB0s1czquH24fDIZhFzjVMHq9
mk6vUNPCRQVn53EHeDoCQyxua7CMmFuzvO0opkJcQ9OP4cPxsL1C4PbBTfjgRMOB
p0ufFHjoBXvCXSS9wonqo44vrdLjVCfE+o991fN2nTUWDa2Cp12t0g7XkbO+kb/U
72zIidJ8kVBD/EsPPz9xioFyAKyQ0JiLQuST9NTPkamAVBwTAk+eKwNwFSDXQL7e
Eh71PdctkMkSm0/mzWqgw/rknorkdtApuEgNJPRKcEqS/6ymhyEQO9dbnyb45pln
YOF6H6qPYvcvqMCB5P8pE/rLpyTyUgT/MHVPLzps8xZx+y5Sb1kWbtP7mcYk7E5C
rD41bbtw9CSH5MO/IgO6JYDPks+zGywcFiOOa0ZF2vte39lDXOA/zxNQbfx9Oazn
Yh/7uSJZoBwdzwYU2mAZUNjMacTSREzsmSGxImYC7+eCurB/wuh6Q8T8t9SYREnA
AogQ1Ana3lEEAi5rW3pxHWmAlx7V9pNIqna/5qYOegGI+8QQ4E+FsAGYXI02EQ9a
3znuSfSN5w9HxGh+3JJmsmR7i6lZ9GBb4QgYASKbL/6tU6zIOJjIbHCgEqWRss+M
05sL2yZsayCSDg9/zAwGUw0YZ5UgPNysDTrA4ScJAW4pIQ+XXHteObad2sBTJdDJ
lFUMj126dcDZcCRbLvgTp/Z6nFPS/AWLtvSLk14Q/KcEWpV8K9sW4ohENwijOeo9
edN6XwgGLfdVmHGuSJOQXz8lV5dF6qde/YNRppwYAN0=
`protect END_PROTECTED
