`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vmJAbxPFQTBUiyqMYWTN3tVPifjcJDv6G9tDow1kaJt7Gx/FSBaQyqdABbd01E/8
CSwgtHDf9MEIC/EIyGK7QGydzAZXg/r/l4tKJLULh9hMVdOc1KmcrN/w4ePe+Vu+
QYYD20atwgYREWSfMz/yD5DntAw5ofeV23WD7ybYplRiEcmslRCAjSi4VnJvu+aa
8uLnHmo3nlIPlZSXQV/5zCrQEaXoMGO+M8mcMcEjhJIPUAECkTogMcqAyQJ8DR8Y
vKI8Km8ncO1GOWCLGRI5Ro5KvK0Ewt8nNFwDmTDnTXpMV6zc9tvFbPY0FFz8QFL+
H+CaofZ447dgB6Aw0srEbdbgUyZtSaoq2APW8jd8NmZLOqMw9/STQusBis5BuKrr
BJUcaxGzfmKzaAV0r5F9ngRYh2OF6mAvt5nmUCjJHA9C52Jn9x8bFoIDiZmJETKY
oGWX+Kp7Mjfao9j4po+twmzpCu4pU12sHjnio12S4c6Af1NOhSMfPMmOrYQWqtXn
5VxVMVkqXPz6aez81KCJJKCAL9YMJuwhq3IhCtsCumd+gezfLU1oGdumyfYZZ4nK
7hFN3ELmYB3KRQcbVTLPv/OZsiyVkKxPeQXfy5JvSfoI6JMjnufz2hdqJWdNTEjw
44laNM3wfHerSz7xOIshOx7H+MvEWBbsf8/40ASI4fgYaLTR/E4RAA6hgx+M3/wV
ur3quzPhMQIgzqEYCNg7zO0sieJCv+fK5hQ9QRmLn1AOIP9soEZg6BNBPMdeCaC8
GFCJaDlEV2ttSmCQTjV2JqtONPJrIgMmWgxmBnPr0RhtjlLSfelUnylrBxkLST+o
TZVL5toM6VuuXZ5SQUDJ5NURlTh77f5fdwn3xN1u0ytlewZ9zRB5Z+8LCy/QDQ4L
PGGa3mKmY59mq32lxn7MyxRcqm5O2ZnvDzyXagu21BbWHDDqBbQDregWAD708ah+
/DMa/0E9PxeqVR8dDIRa5GHYQHASo6ELsagrdxU/0gqMpePHLDGmiHFPJTDyQXr8
19w9r1F8E58nKVIbRcp9dC/65CXbyda4x9A+NOYJkfEcW+bl/4RHwwKjvdv1zWHy
OXOQUxTGAfpaXN9uCfqMf3KsikrKRK0ONvCpIFAvwC0QdWhA7JG7m0C5TBQcfxJp
jO5mOToskRUmshceNXeZGTBPC02/y6pkwvUSJu2Czx8/2GtfUwGwu3/efoqv2xRn
1J2ULyfUDWHGfT1UaJuMSm81mCVCw7ahlvPOqeMUkgQLi0o+YKgwnTe6za+/9vi7
RMDwPmfmrBmtGJ7+U7STr4ehqfZGwEeHGDPQuiFgLcWxQoh0gRodNYaRyYCV+NeU
3hjOa6MZuYEzOZPKB3DeCy3wUnllwhlLrN9oGKRDo7pERm/OOgEc6TgniPcjviuE
6HgjO6A+EgEkpFiXWRjpueqCpbIRo33Fwxy9+JviI2+Y2K+Evh0Adup0mhkDdQKy
FMne3AcPtmeMrBF3pKyuTqIIpAZjGB6N3E3h0MRDI19GyOWtDf3/HP1gl94+32vZ
xyRuBVfeslqrkRSU4zjVbKH4k4B4NAtRSX6OtwXhrLOGUh6V+YkukzaO8T9Skvy8
aGYkRJ28S71tsJn4jT53q1Pxnur134Pnw02rL3ljVpqnwU7/YYCtf3XIy0lzgb/X
NydSfXHeLmycPP8MsLh/G1DIyBbfx+HzF0GiBrKoz5egTL13c9o83Ete7/nQKV+4
c8cC6rhfnt1RhSD8n4cUtjrAAW1ahpnDwmXmS8KXYJ5BuJmh4FtLUqTenXRsJlj3
KRWgUiaoL86fwm7oNRZp44RwJsX0dnsBgdICLHDowiNN5mTcAfD8rrtqHbJOL06B
PFyyJ1AATj5RSvuJKGhYYzXHDEXLHArl6x5vum1b0Kk9iyyLy7W2Q1/Owl4cu99I
ISjNdxrPvzLGBMR/Pr/mn97UAurqTuYiP68AfZErZtufqYZY4AW3KxYqpVTYkkl1
fskNyK9A4oSb4MQI2gskdBe3qNZEWwBSsVczisxK7YAMST6omQNIoyag2Q3pdqvn
8suV4ZhkB7YYiaLnUfkaNsbcQ0T9/uanrZJviBz32A2Hhu6l2aZrTLSBv3draiVx
+AeEdet8NkSM7V6X2iDSCb8/aoV61NgjHEMfi1oWWpLgWiGa515x9xlnsEY6xUNE
klFzJnrjACcY0AQWaoUCRDVsVEjWx2BCA+f//PkJFRU/N/cLUmEcEQIc2nVcdZQ4
tvfBTWfhEnhQ7UadrYnS3On+S3X+4VD3vaJChOBzVTMDjYzgue21TsMREnTUCmYk
dszWU9JwR5AZAFhExH19lnDXHS2BnGFWCDQcNkyxBWIko0s7nMPC+xk1zC+TzJZa
KzPQ++JoU4WcMZvqLuXuHwZEjjGEGg5VOJnQge+c16yba7wMwvtecgQG828ux0/4
bnTkI47qkOTQrtlOynAH2bnBaBjo09NWn4qYYji8JoH0aldaqnwFU4vjjUrPIwWq
KlN+z4KiJYfYK9VfGyONhNIDucHkpnmJp3pjm/GKq7gXCEN9kyqqoFcd6D2lEF7L
/9yT4HafNqMtr1CPypKuIYVWmkkte1NhfvMVlT6OC0BYMT2u5og1GrltYfZnF8tp
urzGmuXzoSmEtm0JihL61PbJy4FAFWWjrweiDbwvzEbY4WqVYEEWJTbObK8HUWdT
IWarBKl8Z5nqD/rsGTGxcDUxny41QmQpksVuP7xnmFWPs+7r0FikL5R9lHgGAozp
VvQDWa8oLHBgLbbfgO2+YQCup/rSypmtdROnHvk3dtXK7buCkXqK72Zn3FK9N7SQ
eogsKf3Yg+3+cSlIOU+JUgxRj4Gxv7d/xhbwuUpV+xiIEQfFWYEJlf8r5TV5K6Jt
+IhZ15KHjXaammnV0uUda+VH1i5OIpV+AJAgiT2NWzfpDU1iIDsBxlZVPq33QQSv
rGHUm4/NqE1aBWSLVdeOkkGNafS4B+b7tzIC5YjQCFc3KoUjG+gXIztnOk5TPprT
6AHRo+bhY03DGuHEwgqv9CTk7BHH1Q7qoAsuLuwqZ69ForisCFEWoh/eVt6ccihf
I8vBS5YOJ0DgCstvSGZIlBN/nbxayGRRhKCcO/ebcnvwCx66rZBnktVhbeeBZi5L
pjOBpHSYJHoEEGGyXUtPUVoMspJRYvqopN6nOkM3xn97m/gVXdg0EUzAKwVYFz70
5b5DBWkFlWnCVBBfflIYkMb645CO6KXVZQQTrmgaaxqRIIiRNrhj8JP+cBnSt5yp
wJvPVQcS6wgkENR6PpzCNcY/Moj3873GzMogqxjE9QLUMsEC1Ivla0lk+ppgbQXm
1/t8OlGhySR4gUNeDUP+ms864I860n+nQYdcjyByHiDLhvBDqk7nesgHNc1PEEjJ
VfGCZ7kuh/fdHogmiwZTMkTvsJlaP1xbIxzOWUqPVN9DCLkXOktG+a24lo22j38F
X/58fRPdAh9y4PYfjw4JXNc7vl7DbceeCtrZLDWbYBcSq2fDE71FOrtKmMST/1mv
OxOoUzZ8ZDZO6spvWV3sDln65autXTCSrnolJ/Pc3pnAU09G2FoKIHyDAzM7g7rQ
xLXdb7uQBcmridxLMziIN6PUvsldSEYt3/6v+hE/hn0Ya55pjqUiTPn85TIQx2UB
oEq7DNBCr0gBP2ZG0qNRtzTHUM4zaO9o11JRNS40hEmSa7vBC2F/oD+Ls6jv8tDB
W/ylU3djTKcebEfBUlEsP82jiBs35saYHrmObpDf/y9vyA9WfYyDDaHMfG8rThBU
erryjxU0cTk602tNOBvheiaHUICCUjstCSmiSnRXPLXGw0IxSZD63QlhcCNgXXc6
4kr+BlKISBmzLTgtJGV9DmPxpdjKlfNiMIm75aCnXkt/ArRd/HtFW0BNNThTt/ys
jlU/kPptBLPUHefRoJkneEGVe4N+LvyRF4XwRmPXXVXEiAi9f0xYuUSTzNuNAXGc
sXFn1hYGX1Edb4bKeQAe1dal59lUAn4+d8tOhwTZ/pF4hXLQOFHnQw6WJdq5s82V
GZXSgzbRDcRX70TiC9nbdw+LD1bJKJdCtbASc82ezaweQbk11DOaJ4wDDhG6htA+
ApC8rJbkP+UsNVpn7sSjdhdBzAT9PXrRSpdnyIp/F31pQRtwlaQ0XrhLWbXOPIVq
7f+W4s6j6o0kX1jjYxHAUVQBLRDZCBkyVTLdBsFuCPCB+tKvpFfxTNtEB4j+RmSE
P3kMNEs4wQPUlj5Fm1Tnj4wIfaBY+oRHV9oBMf7C3GQjSuulGWbWZeHUBG/+D6Lt
LhJCVflI/sAUeVXlFBnr2vKkQd8zglSdfRRHYbZCIIlni1rz2yVLQ1uVfIREv7/x
5YVboccMwPqIWukFxxNLy9a20DuITWG3aJcMXcBlIpMbJlqsBGkOVqRV3I4anD2O
RB1xqaeD/R3AYGA9HDMzzeotMZ2hBBVuIZ6Thb4O/M1moDaoKalhoSY4cewyFcJ3
4qKD44E7hnGMkaKTqNy8olTMBfgaAQDnXMRqy4g4Hx78nWDPnnGLp7Jhn5QxYNAB
8sO8PLptsNDySiboyegz8PtFpb/IZNixDROPOqV+iP3Hk880l4s2TA339cq+rIao
7nImEQFnhplCJ4INbZzfp5F1CSoO0847xP02RzmB0XoWw+sf+oP1QNxisroKfjQv
IEwhJkzoZjfgtLmhoLuIU9m0WhZA35jUnWX7xIleBkF/KF33yxnYHfI6JSyDmkYU
6qWnSoRq+zq6//OLlQVgOx4CzH94aBRZnyF2Hbw6w5zpHBfrbN4DaoqnmSP1KOSn
HLhSq/388peTFseTHysK7mbJUeaY2zQwCmcoPsk15YpSuor8BKfiBZZpNKvSqRHF
qOXIC7542m2lu8I4NS8ZcYFYSW1/qcXT2PbmACM3BbJuHuMsRW0QqXC84PSH3LdH
VA0vbtjmzIi+FHwW/bsvdMm3xhY7qJyLJJ0l2af8dLNZ/K0SNp3bFvMS1Q0uaXfI
DVkZjEJVTqReBFgKyLuFYAchlGUKF7k3Uvyzrpt4eOK2dgZvVMV4VdcrWRa5MZs6
TOQ1T0+ebWSe9nFNPYgaaX/hu5FsTgncPmIqDuw0HvPJ5PGuIOXhKIK0oEUfcRMI
C1JCS/lyhnnxxiFJmujWeiy1faVCSzih/eKhl9PRf6dzz7LTHIBxQCWKUdDxBH45
fKplcy8F9Gd6Nsfue2aLz1AJilkTgNwOoNH3uGgWqqg7dtcim+CtPsbHNqT9Ggos
kyKHM7ZN06AwQlDcNu4yJ8oggORFCWEiuW4DSD8v2JzBkoXEByTfHR7/+5Qk2sw0
KuQy0wGRQV8ezfl3rBOClXC3B+UAkJazHhgBTtyNAuGpOqZAeCC/5vL476a3vq7n
5JrFp03by8AtqiHnarvKEAqHqRqp3/4/Rn/xdGhijueLVBOmINRqFyeJV3OAz6/3
IDe3Ny4g4dYmynMC6rDeagkRpXU0mR5hzZLKGw+w64DoLDJOkyT1apZmd6150qY8
42E84/i9Y6dal1irU43ZVSSrELnZKG5DHWiR/CGSQOKKd7AdnfB08nD77LLiUmqt
BNbp0KH0FTOE57d/BCMTlKsuA+SooV7BYX5eaYTWv1OOYFoRoVq37LiM9/A5etb7
S/Aiwd7KBGpBGmX5aUKir3PZ9Mf2DY6XQIa0LvEwNGxszLdJL1bsvG2x1TvCq14d
DthxW2aOogJzKptICzGxz0AvbAzrh1LE1k1LradRGaX/6qQlD8cAnBC8j0l6kMzt
qideVDANrzKG+Otvqm33tmG208XzSOyjMqiSZC+njd1IaPWSltNyaTafxUBnhhWg
SVwb4ry4Epjja2YuUuTlkM7tomlNXJnJeQ8746ZPFcmW5qeRRNe3uMAJj4j+w6Lh
80L8PvpNsO/XKEAKsw5aAiqiMlqqOQJEBf4YIx3ViUjqdcZ7gvPm0y88LKB94Ql0
u55TFYiaz+7kwgXDzYnTXn3JxtDHamU5Da+harZo8ZGwESF6pMTDU5OzNslJOB/B
0JVcfeKJoxFkC5LUF8oldzAiIWpFUtHYo1GvvPwjTxQOgsvTsptNKkK4FbHcMSD5
ECXuTR6XQWLcoG0lproQAUD/0qL8TCj8FMRROMHE4ieoAMZg0S46/qUfEippgJ8k
iZYYvgs/zKiLSYo7lVN7gmg5oYbmLceMWzaLaWP+1cVsLkT4pm17dFZiZOS1R/ty
tUCYg9gNIe1t44avfLStkVNtXJDy/w5XYpBT9+h8Mzvr/88v2hiU9iMU6fsZZ+53
wLTU+KJBZ762gm0+MBD49BOanpyPcTVV8QbEqA3BHuEFvSC4qO8nXKvzAGbYkiHU
v5kizPgtNnh2UycCIyNZIOJS1dTanOzeGoW8vPfP7C7PrHPFipoSpFrFeKJcVtJ7
wAer2sRSP6d/dlzlVk05IaeqmSmg7qsf7VnmIeEdN/Ok73Uhk4U5qYWYzRjI/f0h
yV6e5dEzQd7X7HqaalcRcdR7p416gEvp5G4Dbgtv7GAnZXuavig2QFxfLDmo35KY
ZSHwzcIy0hc+VYqTDzMmqcU0wyhmkRQ1qPJwelHzmcPGPq50QioyAT6o0QpU30jZ
v0E5t/EdezNoVpqh2tikV96NEuppTTaM1VbIwPGAWKtUeCMX8bwcw8QGw5KbyegD
8bJWaXhMQqK8IGAXlzlauh04ya8OESs0CDoKTEoGJzmsVwabmPj2QnDDbRrkk0oo
S/k4UC8YndujH8Q0roJ57C5RE9s9H+t45rFY3J7Cu6iuZUZeer51rpr9ygqrQkAI
IPbtSQDRdcUVFa4U09suFVgccfzPqBQ9nG6WDwjlmWJ+p118neQFpE3exwEnJKzl
+kK7p9Cewrr9jMqusxdisH5YIxD2XIw3EYW9NHVf/GtOb2uMEPn0m+MF6uoEJVGE
yUsO2i9wDfpTQZDqROmsVCvQJBQK66CSlyqv0qipmb90EF26U1D2H31nor08jhBF
UOGNeR11IKgGc8QVWt0TajvCMljGn6YD7Wjc4ICvifTxnplmPpK8piWB3HybOXBI
hvaXbM5ThKLaKKwuw8xgfOkHRaOq0sr8uYpxyScb8pvFr0jS1q4rMQGdt5MckLUf
zbX8Ck6R4Kw7TMKSsIx8J+k2inOfZk6dnggkjUwu9UOtUPkiQg/OyQGD65x7BcrP
cJKGuYf5RMj50X/uv76XTCHRa7klCsy+m6fFfAKGWt5wYqUUrFpOh4sKsuBuZuo5
SWFjA/GMHdzFYfPo+WM2JWM6yCviNGnvZ8++WxLNlcVYFwENPmKe2VVvhLxE3p9I
Lk2tIQTPsxP5fv+m1Ctastwv+jDV2IJ50IWf1+weX6s0kPJdTK2nH02vaPicMOx7
Ywgmm/xHvwAiEHWvfOFoN3Q074kd1csafKueYX5zP7UF6TymGB9aq/lFijdcq27X
I910TOEBaiw1ko1yhZlbfdSEZet9LGvZBpkriwpSpQJsYT4rqCMJNvpN7qME7KwI
6Q/EJ1ccOgPkjfdFqP92sTzwaVe+AGxF7kLb8iqRrFEDACQIq4RWubIaY/6iritv
tBLKtz9/fD20itivXCJkb4HKm2G5zmcbjkl7z2Y4f8aDjZoCKpBtIhBMGacVauGF
b0wWmQcxF6y4MK899mLO/PzM5tP6rKC7IpYwnjkRv2r+QIWoLyuXsdffe69fFDPv
FPsitqEvhsY1AIgjv86cBlKPjcwCUMAq0hQGNx2xRGHxZ5+0Atlu0VkrQNVePqvW
iF+b+Q0MpFQpSP5w0bTSBScGDMRnJ2q5NMLo99B1nmIEF4G0qWSNsKk7UenQ4uHt
QFDkOwYHpj+emgzhEae7mycsNHagF66gXKouGR+ZKPOwLp68H/zE6kKHJx5EIG7u
t7/nl8+UbpYzLVewvBaQ/yor2TnYq/zX2uEU7SyfK6NQi1XxoSTWYFkJWPHhxAuX
aFS05YDuYADhtKY/YBxlhtW2jsVGj/c9kviG2Es982VtXpulHdcUbMRKU9eUbRW2
QpK8nxkOegzFQzpl1MsDJuUgI3gHgaEFvOnSGhc9LzLS2H91MK1LOdfHPvl9MSnp
Zy+KAjGlRG2KK01HKycHTKQK2jy8ahd1dgMQa599AJNabFvQP/bTrDpuhD5JHPJI
oTLRkFq83A8C8ZI5+9+PDI9zl6hifrQVqNhOjN+YEGAQaiFIncqNouPJn07JFpMS
mzfAvLxY/mzg1PZvFTv3gYozXPFAgy3p7oaWndstD7E/Qtubv07uKAolJB0dF5Ay
BCZzvwYj3RY6fPBOv9dEKmlnOLvJWidJgJvMqYZdvfkQIMVlZIN6I8YmTRw94h8Z
n19+YQjCVIKOocfPyiPFqYDAtm7L2wNkUETnhSo5DTdcSoGWJpUQw5E96s5g3m/5
HQByOKlct1P1tRmmaWKFgldUNVykT0yg/fSAmXG8kls5sz0sJltnqv2K2fd1E6E6
HWQykkZizucAQWpZJZuLIZYS1lxuXhc2WOCYe80N39v8gNRiWK+pjYgwl2EAL7RM
mY/++Xyu/o1e61JPvKGitGqzyorIGvUIraoDRe9IQwIfzAny7+zQMPbJTGGRtX2x
UGagiOMezcYpYw41nBYqywv2fmjTF5IYMoupVjHn44oizXfyzAHEU/tFPwojH0kc
O6pAOhzdVOva+a3WiRCoubbp4QDjKySW16+9ItJbQ4YaTHCcShwiffQX8xvrW2I5
9fFuXyOKaaoUnHImhlN0bKTkZFoW6HJsFOIW9ENbPwfZHZSFQmuWGU0/4O/u3A1C
4PdsGHBMlw2CZUVLhMvKZyOf6oOh2bt5NRniyWRFO+06/6i4u2DXR1IJ/x26oZpW
Wi/SEQl2TFoRIP9Myi6zIwlRKIODTRgZYPUe0FRT38BDM8OIm5r0rFqw6WdXDOmI
23iJddBchg/CUDPxMNRMnleOhlxqlcYcoqq2Hbt4HBYkeNkviXcqn0M1q5hYX6bk
v2uARSsldF9kmhLTSe4dqS6Gycz3CnwEghpwJEPS/s2sdiYHZH1iwbbh6VgxuDEV
zrVBBlhubTe3cnl0NfFUkSgVR0IgDrNIrziTIeamG4gJvc2RZlCwAHFciddjZf5s
yvk1z1DkMFQxGBRXDWuPDDwu0GvzXftzohdFIZBH/e32+DB1zh/dAZ4US2Fu6Uck
F59zMJAm4SDiD0cMGAJvv5ls2mV32nfD+3cGnmHPLBWvVTbRS8KWsBfEhvHdvOC6
HXaBjeByg3h1/UL4Vy1D6bPhsb/0/4FmofqYs9C9qadbjf0oHXHaLLGeJwzpzkuh
1TocwyLvFE/PR9HDwmwtkLdlORrkKL70AbdfJ0DYiNc72HBMHKvcoOnOZNEyisHH
/N7GC7yqqKZAyTUp4LwDUJ7Di/840FuANkOFD5v2c8X7IOXm/yBH9FTcByGSywla
4hE/1+1PmseVZpccyQ96oa0sV8r9ZZGobT3nLeTg0TbTXcHKUqao6apBk+JHqr/+
VFLe7+x3wUgad0cI9lWySzzXqFyvXWdZMQgLO97YA+sAdtW4JE0HAkSpRTuByg8k
xnNvPA99ULKcHRvxDKdYA57XRMI4L1GD4e1uGKHbH1GrN6Q278EdB8lvEOtj89zL
1OBf65+iIpoX6DcYRCbBr/cBNz8sFSzNHkC+mifLJU7sgYCawGZHqW4NU7TJ25bS
WYKoURS8n3PHMuZE1jEeHfo42adq9Rlrtx8CMY6B4T8WvfvcICfG88/Yu1e0dfB1
jwcokD60Dw7x7sedaHPFDKnIKr3SDeW1kYiW+Hz9XCwwrGu8eNx/hZ+xH6s4sGct
rQ15v6mAc+dP2Q81t3P8eD/KmJvkbIZqaW53lJmS7wJ5WzZ9BQXGZWsgyjH7ao0v
/Ov2QyTIXQ7H90XUD3SSwbVRACfFwYAsdvCSIxypQri9U08OSoHkZz3Kc2a2bsSZ
iH54LQHWmD7ej2PLizYf0GL/wCTBg4KEJqEfZ1ZfO6gI/glUj7TwLvolOyVBNDO+
T3nXRb9/hnoAGEhtadIuRm+YE6AmacKFj+xYVPX4jeYinThkGpg+yXmIuh/5VTrF
gL3JR5XImJEbux4vc7ZCqvOkWDNgytmIigBO6EK9BnuE35Fc2a5b5TnMIHBKnJkX
EeM/ki3O0aotHiOpkKaYnm1KRC4Cvs5FFCDiv3gUNRngXGfbErk1fttnDuGikiTa
RgmCnnpNQHG1GVNak/SrH8HO4WhFETyOtJaxNQF61ktY5cFgkc/Vtul2QQyoXStU
ZbZF6gUBzPiw4AO+NzVS6nCEnlzyIhCyJtZb1nhZ1f07R3W+qjrSPVD/4bAxKA5N
Xq5Kfov2MAsC3c5hO/MXsrOE1BLYsBGIcFrARNQtXAHQIU2GmqQrIH4H/dbaGpn1
sbdGXtEFNdESSvhqtwLGftZWjh4iYVcaJxnIJ7f4XP2zzFLPtvhpDg0J1NdkTOSO
7dTBGam8tljy3JzPUgZy7gG++YIEjc+22AvGfm0CwTZLm2FHR0HCKY9GzFtlh9kN
oSqjemIS98aNYIwNiLWWSI9Z572HFrSkDHNIKhiTliOkg4KIwDBHrOxo1QSmKhOL
RuTzxJ9l+y0jOU/nXT+cQ7W0Au8n5OnG6UAAS7ixM1TSmJ7Y5K+PhWsCTuEgbtFg
OirTJ5X99fKQ3/H0241HuRjo5sO+ec3hHmCTmg6uTDSX6l9tC94gGT0DY4xgikN5
uAeO26AqYVJuSYZPIfSJxT42HiwREiMIppb2n1d5Y5VGHvqh8vvD35jHch+K5j4L
bhRR4DyIzmPv5RhM39TqtrxJtUjmFN9YDN79ZfE6iESOVXhISSfj8u8H0XSUBm9s
TCyMFm1YtlnC/gZpd901ow1S/7f1eF+QvhjtLYKqyIw6HSLcx605vQcWFlmHFore
SD4pIjlz6Kvqo40tngG5PvKvsM4Y9OE1OWLYW8sKXv0USfJ2zri7izM8IyKkbaqi
6YBp3NujXlSnca5OQ4JWOJajuOMMpQYoRMo/KVsR2kkLYoxDt3RRNTFaTxP0o27s
4la7o6eDMMa4i+Y9z8LkC3HwoJUTQ7ugWHwzD7jRwQKY/VSoIi4ad5KR7xVild9w
f0e5gxPSa+baYeSNeYqvS0QRPLQQkkNH0rkwYuFGndh+mKKtqTY1hAgTznJanTO+
bUvZG7qx9siu3uPjdTcNpdXTHMq2fKTXsfmucL5v/PH8Icp8+bi+0aTTSbLGVMR+
32O+zLIOGTzC1LINHlZkiX2UPAAvCUy0TGSTm1vj/BeiHjUbsJ8AE86CbIeE2KOo
EDafZszKkEnARk6EzVgLRM5wRgBrAnyYwZFTiaOA1RJbAvZ+SAOzNTzxG+Kr01gw
cXK+auiTdutGZqQCdc5li0y1IY2ZrRGrLy/UBaC+JZdkYesdhlki1vEm+0NvGmI1
2TFzi+bqII6ZZrkwjYAbiHiOTZV59lLfCk+4VAMVB64/KQk/sz37DnNl1Reso0pc
KtGUhyBXHZnRsCj5PH7+hyWsEvwG6iEzJKtQJTcdECCuSekk/0ebK5sXLUyxXvGp
jObxF07AsN/QL/CMHoZSxNV1W6d4IGvv/fJbbBV7VwUPL0jyVSBWBi3bN9GqpSXB
SxWz7+W2YY9ykJxb3qNaF6hKdrrhA0YwkmMwd1Fxdl5sCbHJ//51A7s9d6bJwLrO
0OaLUUjWkhw53jRkcZT7cZeKQMLCTEF/ojPwhlj5NIQWGQDMcH/eYAlYwUGa4XRN
k+J45EWrZ9dRMTsnFP/NXrukhpyYytGyL970O7TeTah8/9GEag3HLD7TsxwBJPah
pMO9rn7wVqLH+VcM7BL5N+dkDZAjzBU7uDB5R9ilr4f7AJzcupu6olvF8V+7itqj
psGa32iJX0VjW5c3uIRbp0QeTIzoeasgLOMB53nCropU7sdUUxU/2nClW6ctCY2Y
suN2HRPt+v98ZR/7LRLsvKAtl5kK5xZrdYcaQuL2qcFtNyrw+1ZzI2v1Wug4ED1w
gElCY0I9xUZOiw3wdWB5XCImoUP/F4mf9dHV5PtwjTNb9UOtY+Ay/eBFMCNXgo8c
eBmORGmsDK6TGYLMKqHM9uSGs4mTIQX3g5o8cDPuZuvKx77lNci+vjKZjt7QCFn2
7b47pBWT9vgOJlC31trX2swNA6UHMBFSYIoJfmQIKB1hViHk2RQKqLla7ALSk7Ft
/bwQOwYDxcjTudSutgCy+jutkKEAUvfZNrRaoXCpGrwBP+ZZhIn5G7SOFter1LLE
nOJu8f82naZJRtkfH7rKSJDeh67YZs9GSwEDTs8LVsXETg9m2SOT7zDnkmPxnxxW
1r01G8PVMbuTHCn/DLEx5YxqWzZwou+45f4CZVcbQtgtaTXKghmwsKDRwmfKxgMi
KxNup2aKRm3VtOU9AKZWx40plcG+hkzZcgJzXgtQMhHDEMXLwvVaimP9AWELLIR4
Ff+gVRCFdHMzPSd0Cf57cTCwdrl4bWUVp6A8T2X9D41UOFenSLjMJWkCn+T78oB4
yqq2A+8Ers+u9h7F6gNGKlTIUL8SLVj/MSR6uDUqVhIVKQx76RLLti60VHBD23uU
eVWXo45KVfOb4wyoHk+0hMV/3gkpv/CPp+68MKBFMNERQ74uqBHwIp1UQo6uV5eM
s94sc5AQ95bzk3Bsxrrzq5jLAcVzqxuXsXW9/HTC+ZtOjHhFYUnAhoXsNvfS6gza
fBmiyj39BQFZ7/wXw7DVV4M0s0WezZYsipjYAfjHqZnnb/kgZarxzC7Giom2SKuE
hXHF19Q4u1qHldrZTZVNys/ripimwiGioVscKZNXiiXceiuGwNTogOHve6LiLREf
ku4a6gEo4bS4YxEqnNO5BBXNm8K9RtKiiat8x3kJvIHWInJI3T0XzfmlmxXqQGI9
DW7pt1wjfo+PshiXimo1faNk36UWmBxcnL0oA6t9TiPHQ1K+rzskajeQfTVya126
wD5kJNiVQUBC3J+XtxX7pnsaIDLcceeWdYol+TScPzJNAbKQgAE7Q7xDERKvU/Tv
wQVJb9XLZyOEEOhv9Iyfmkol1FSXFjCb4/w8vSiHNDPjvzjtOTc3uSxRLqY3Z+vy
CbeXH63jOFesj3TmusFEKFqwyoFIOUkb3lpPcBWwE6aM0GpTGb9+ffhsgz97LQc7
ol4ybPExLPE4w+3oYw1W96laeL2uK4G/6H3K7M9oh4SjnQf6aU1pfbG4DmBPzDte
62um0OR32HvuR/XYrCoxPYohzMllwVUgy1LhhT83G+fwRb4j9D1JmLMbciTvSDuD
glEtjbYYJDg95Dn2CLsokgDTqOt+ZgLX1XaiqoYaH+IX9V7RMYjyS0AfFpqwhM3h
5Og+FLi792gmbxMtbzUb6+9oS++cO/trc3K8evCOydbF6GOUwH6+BxGIMPT027rZ
2kyXNWi4gxhsoNUNHqkwiEvNtKQSxskF1vm9JyvV+CWw9I+Tycve7OazE+n+JT3A
uThPaLU1f8hBmpenUR9lEhFic7lhzJVOXNKfyx7j0ZlNH9gHFgO6JzjbXzVKBwGH
+qayvDNoIV0Wg5e8j1NbkC5AIvHCxL1SUXnQhqnJKcIriBAIhbW0jQtc907a4vfZ
Lc+IcWzJYqvvOg5LhdgSDTOf6Xh7skAJtBcnuVMN37TXnFBmPUzNH/pD1NlLkby3
2YYy/egq20hJNFEQyRWrYh11UpGs12+9X0YXrLXW8YgLumAKoLK9NuTvoEqaLKj8
2HMNrXaAARThtq42wXVMdHjZy3oMl7esUuAsRPU/oqk+TFeVNdB9+cyKGsLRlbpy
M8nMVBssZEwLAXhRUiKn76aaF6XEYI/bmDOs5UJ5ls2kWbIxbi5NF4eLCtd9IwaH
HJbMzdxR/p06hHAUy9YkRqTj6Jn/oz2KYvDk3zxQeT1JLrQI8ao31yTpzvHEBqGP
wC9T9f0ZE1nLVJUOSOoTpo2eHiBkEdqtbBmJOnbt2bsypPYMBVjkETOWAjlgsk63
N2U475JKZtS8Mh5h2nn3O9jgVCpBpoahbwcZyuPDq92FynBrQf38rawT0WGjhG62
GAenB4BXDz60adFXqXAbUwcyWRmaU0f6L3yQPq1jx1a4C38SpsUwg4PAnD6FMRoH
VuHAUl6bi8F7pM/SEXCE1+SjEBpHjA45/HR0DRFEMFfFQSCOh0fKy3gJxRhtl2wh
DbTwhqb8pRODNXkjhexO0BKVICrLnHGMsvmm5JSvYiOwGWUDw7nTnI5XvbWZM44M
4oq9sR5xLWHJgy3WgTVoJeTHwlz5wAgy+heauXMUO+b84sFBuIevWBiJrq9K26L8
nANiIdR02TqBrn8meJJhQNm1TVQkuwUmgpLP+osWRMUrpw6EpZNy/uvGS1naipgc
3xiLjYJqlySrvIbruakHiEus8zavhQ2RKQxZmcRKcLNo953hCihpKtF1R4sSOKEi
OX1QjB6exAOpEqs4AMgVChkFI8dqra8jYhLYW6TGiy8lOVuxKF8mdV4qgVg61+Mz
o7LNjxYSYmKOxSl2wk74xN02nfMyOHJy1pCiVP9L6QFSETrwt2HK49uH0x4JtCLS
U3fJPZOUPZFIIRnUIp1m5qPrK35J8jpu84hHWr0cZaO0HHCUc+GyK1xMPAZBcEgD
+UaO1TX/QqgFTfAQ4zz7FuADnIcF2ygk4sXUIJbsTo/sStm/s5nlX/LiFlxHizuA
lbqlaKPFqYK9MNE76lIiCdCHHcTaXCoKt4k31+h9E/sLdMiONdrqGXO8y+zqgAXe
E2Rm2fppCGOIGD0WJCKQiG4mLRY1jdJjVg7h887Y9KwcyZbefbMPJbo3jq/5MhWA
bidmv75MShAE5ll0glMymO+GRMVJhG4jXE6ZFhOGSNbkDr/tohn0jvhgC5urjCbf
83QVyapScqaQcCJz5KbeNGWt8B/RnKxczDWYRJVZHT7vFCETTmOodWFRtmXdfWOu
67BzgLN8K3Ngnc8uHNiJKG4avU4wIUz76NDBz00N1U2RCntaI8GfZrmslV5C5xV7
G20pl641iZs1dxodpyRTFz3093o3V8FlbqF8294Qf74kdD6wdslMA4zNnlGyBxsU
LElDPjx9zref6dFUDu36/PDijGSndhbe3wN22DBuMn9uhge7oMk7Gc2Sfjvn/ebR
9CySkhlOfiETGaNkQMasqnYB5ceL7wpPSITqt0ES+fkpDOszQhlrR1yV8dN+IkI9
fjcvSQ0q6VONmZZysVPVM+LdXO1MWn96l5z5oufOXn0wnAYA1Omhp/Wp07EEsqED
zh/L0B0RvTU86MDRmGMlzeMUaAIProR2+uPon/mDpeyZaAh7su3pD3HN8wOtbWe1
yn1mqUqZEMiF6nqAP8XKIb3/rbmW4mrmwYZViHkn4Q3WwvgXf8St4nwAr7HXqPib
5x6uOtZnxfEtwwlOeBkAf2/63UPzYPc1/UP38d1HUyOTdT62yLGnow03KeMoey0T
jq0vgIJLVC2Pim/f1cjoewvat6dH2N4Q7K6Djq41Bi2+/1dU9uoHtYkBP8PiOa+R
8zzM3k/i1d+Zp7P+AqNCOT9SxjWzGYZ3bvW2gOUyYFyMKyW+8PHwAGRSR0qm2wba
ApEkiWOFXYgLbYcnO4nPkUqzGzksojVLJqwzp7y61a7TSR6Oj3hBUv20IYlfGZN+
v0tyJlPry8OGmalO4Vz8m4D/f78Zyx4W2g0rpj7OsHe9t358XpiO3FDnbCCRmszJ
7s693+jPUEuHJA/AbopDZZ7dAoGyKqjxGTmSg4KS1r7fi9tR04pQAZxYfBTJGVmi
BtA1vnkFeDlGioh5Z6njkRKlWOX/UmDzwYGwawMqV22JbnCZDpDO4tviMYz5A0hK
MNTTqfhCbFrkGHByUecm1RQln0OTUQGCTJ2RNOvALJbe7kQPFEDFOEPXP4WOJGZs
Eysc3+ZR7vlvjrp2Z2trgsd9+PBwQkH7JWUCCZgYFs4RVsjlmXOarhorskFGF4QV
09dGrPZ3wpFt8eG1D5TWH+6vh43MXqUJwBH52I3la4pS4Wi6jz8zO0VWzQ9FW9wc
SKDtKZrFrWc0Y/kqblMifVBiS9GPv64CIV4sA9OXxa/66ELpTX0jOiJht3O8GnoJ
SbdTj2GPENlK8sVxmx3A2USh6LaIUBIuxSV9KWb2DFlUJ+NI7jXd2d7bAe0QGkcB
LLaISHwFgxJW7pHj1ueXBzyOvB9KCJtKPPLX3ExaQuPl1mhatirL5BL+RavEA9vL
5Pumr0+8OtWF4DPO0ekb19xLVZP9ICwOnkr+ia8hT48OjUPUgP8ZKeIOwa1FQsvw
i1dDRPl3GkJjXUzzCmItgKhEk9m0ftfZLk6uf4Q0kYu6axfNdw7tgG4wPmfRWxdS
NF1OJsaIG1m9ut1QaiYKm89hpLAFBXXartc/dJSs9zz9CYiI6Y2UGK5CLdjdnNop
5x/hiJmE5NCZ5V0nxf4/leUAE51z7DT8gpWzSrfML5gMsiD+tbnVguxYA5l+uZsj
W1lgwmot/uxSjFbMRMNuWZcz/ltKJzPIwvOF9DErmWKEtAPjrTvAoGQ8nGThClg9
5IGJKMYjloOumWB44vW7Ffvc9QIt0cfGEWs3cGVFbg+QqheblSgFEQMVRjfxRRfc
PJg/G8uU5GDjdJzYWHll/vjcZMnV7DSJ/KD8iKYCw3VdfmSTJ00E2y8MaM0B5x57
gwsRnRNwTPhQaz96x60eSBMbCOs04kBszoFbmo+F/lCUl8lPenFgMrfsA6fU3RfY
64SNTO/3/tp5OWU7Q9H203ESgB2VQEoWj+WeFSN6jPLdNfX9oktR7fazNB25DjUw
jrcNbYHXYldkjqbSvz2Xt9xepObO5CHPvYEuekbVMaNkO9jhkUdOZisxBLDSRq6a
UkfyIzO2asjb4cGrhCRWMwI9ibDDqeLSSP5S6knZXe8D0k2k7keykKZqBAAfx2US
OhITw3jUodfOs7qKRpf2rleyClJMLqCOaEzVqgjIEV+KfOZWIyMaKAvOE9MaKHCx
D2ftlKd/7F1F4Iw2A5vrTA2ReiYt6O5DvMJCaj4QeOvMp88x2AjqCCilH1PjVchl
Xy0lsMOuzpQ1KJh1O0gG+26G8+WN9KBdbSzAZev5sXQuwapZgRXh6jrShSP+r4hN
3dQkvJP/v29iEWEOkxNn6DjQTATlD4GTQwDWwgG57OqHXrURipNLYqyyjhlLBxMq
xCnUpdhCQWC8OxwElnopw6R167T1c7B7v61c9xOwZR4jPLKPbEduZ9NPrV+tv2X/
4/hyKJ5RjrBonMpTdUBIxY+18JlhA85+YZ1BJzrsOuBmQ9tg1xxQ+c+Am12rBnfY
m+TyOcM9Dk2xMJo+qIKhjUGrFnyxpe3ZRpTD610+ZL4x+YkCnpcSmkuSI33bycBB
m9O34lTMOe5KCPar33mjh49EjWdjKx3DtA15tpyX9jnq09o7j/udP6beuB4Gyjvc
OtQF2Ut8ydaIdyuMDTpjG/0FzSGVqAXloDrzHAcVMoLA92u3e3gs6ozx5sHFq2q2
nbHJxosz2IzX/NjM3lZM49r5GH4rM4g9Cf5Gzm2RUEEB6bPQAoN/MhyhBZsa1OD6
pp7eNlai51qWu/9sFwCwAzYxS8QOPvbcm9mSmh3GHgw8CLSlexp5eWQgqAWPJ6/j
XUGUr1WSxaGc9DvG7Qq3uM/34uZrydUOVBfWUG4GRTGxz2gcoD92SLszEoOemFZY
pOxilZoDCuJwtbMVI0NnRwr9RTGXfjerd8tFUcZu3PTXtVdLSv/NRUo6dMCoMKAb
Cir2iOwMZ4VMFWbL166E3xGU6F7Gm48HPvq2fgho3Ne7Meks4qbabhLIiTmX76Ac
ltvKjaAZWR7e1ktayZ9jseSqKVeCKPZLt0luOHZZRHVyEQFQ+dP5Noa43+FpEdOc
0hig1A52wT6I/k2AOOg0+4gGjFLUjzTb1Prma0gyaeyN2Js+syJTE5JoSGaXvl+O
iy8lWK8CU+2NqYwfI5+NHCE+AxbgWqDgfBCKBwDOcFQqNlzCY0b2y3ZjRqqVyXvb
fV8GRZuf2pnUiRSXHnc/VEtxpkOBhxe7VbL0tBDArP93r9NfUgyZKoaE/9+LeQwV
n2B3uf4XWkQE2d02VmhZ4pIuR5yMP2Qie8do5oB8cs/ADexhpqUF6D7PntUgTwVk
7WD8uMypTZLO/RAr4dBdYRY0/4Hd+gsYx0FNjbJCESDdI6wlQfvk4JbNmDCNZAeN
gof4yCvBoWTDg7h1xK/hAF33+OFEPFO+73oMsyJNtdEVZ8Gqm9mzbHpIiqGNuHWE
OQVXESK4XOwK/WYgXphwnO9MalqbTIsXFDcHuDsH3xgzcrNPkT9D/StaMGot3ES7
8mFoR2uX7PgHRE255yt04/pcRlA9GZ8dTFZ+V2pg/DNe5Jer09b/1Zj0J430a50c
zFze/5S0N/fb2vRPbEvFY0nXpVF2pIQGZc1r8mQypUhro/tgRZ1txfddKB6oCBMB
90jwAbTikT/d6Vrynmbe0a0QHBMfddOxDdft0mhpJZ5H+Fr19UA575rMwQBgBkhH
TdkNIJHIO+1C4Zsy4E3zPlYNX2l3hTeod7zF60y6bgii9K1ImcBG30jrErmt4nA5
dRVzcX/+m74Hep3ysxJkVuQTVrAMKznTv4StiIOU1yiZDD1JcPWNWM3hHirvgy1z
El8z2+nToftKZBRadsNzfFdHyp6+YNtFT0qmeaYYG23mFeLYLcS14PEvBKrZfqmU
t8Gh1MDaaOfLedCRK7qhjxnUgQEBDA8bvbqeKz8+qi7R0f5mMz8lKTted/7P9e4k
h1DwEfd+ux0q3iRyy65/AlOi36UTcep2UeCIJeKO7fAIMByUN+DwxEWlRK+38Ht8
SUzygFt/O+dn7RjJ75wJ/JX1Zq7dk00Ug+2q5tNykExlV+lPWL4RCPq2OxbNG+3z
JcFd2xg/CHpgoPAjrqa3jgIQOxOStY/vy/XDK8966D3QGe+5d51FSP3i7To61LNG
kGGttTG2+Two6Gb30hzoPiGAQoXrJTsQissBzH/D2vT5PJj7uIHf07VYkrsNbM3S
ENcXDWY/ZgDcKyS8VakxTzw72uDn8796KEoKWWBAMY/3Br4stErIr7YaRGpLU9CC
Moya+tmHMUf+rfoylp6gkSSviuedTCSNHkeZDYRDwovuSWEX90YuyL4KUZ7NRSrV
+duYQpKtFwKJtNGZstg/+ZiTVDnhy8RPwrpOadRQEqRWCuWmbnskAciXr9wX+xcZ
daLurBEzjC2ht7+B2Wuybu84c3AwlptUljbBbRyj2mjBcnr+2zpiGBqHXsCOMYLB
CesftSVv+GErkK9i2UP0CjirvhH8943AG2KFeuEItVutjLLZDiEncWOsX48eytZh
06U6ucH3ztuEiDRsBeX5vXt90yhukl1NbSZDbVMc2+UYNNWUX/X6UnCsWWbO4R9c
Ah1r1AMGP0JuymSBKM1n0UuhUEU4n9DgFpT9ETAt0cBb7XhvFXus2U304RH7L7qZ
HogJXCvUPwnhaTpBhJf1igT/NqtY/nXyUi1eCRxUf32KfXjMkZjaIVHT875BhShA
kKIYhaoFGMBKZJSXPp5iCmj2LfuS1d+PPubKNsR0YlpazAST6qZGpNWKov+C0HW3
mfnYe+9DGC/i6DBIEG0T/NTJqPEOXw76sTQsnilEc1uKI/VDvyjGHdWEuB4c3F6T
ig31IvIkO48SQa1X04KMWeng/6G55UiwOBZ4xS9HU3DZrT4qJfVZ2ZkU1mRFe8n2
xSIguiXI4oXczJUJZE+IF7nx23SJ9ZoYdSKc4A1thXlFCN2/dmD00LsvCle8VToR
QpZP3hN2aVJ7Ws1PnkzOR10o13YzK+KbvlItBU/X2COiyCuXYTtx3TxmgC//59T8
YvOk2pkwNGRNK5XeuemeP9eFuEnz5YUJYdTar+OHLOs1WuIjV07gbxNPutzBFOL7
yCEdMwAkVW9EtCN1ZOl0l4rCLZEcVEZjIVWnKvLaEJ8Y40VjtZ8fPIAxzr1oLHjL
SyBOKLfU3bCQT8wavNORWWZEyqzA/f1+dN8KG0yc9dbv+ieTLBZXiFNVz+p9y5Kk
VInhGwycvew71llUtqL0lB87Scfb6wcctMW/ymY52HG9UiylH6kIlMw2rs2kcvIu
DxNT1x9PjDDtQCS5i40PlFh3+oCaDYfvhqYYHM1Dn3A4suOirbHXlVIUI3l8b1cg
oaP1u05a3NTYVmP7CdnnFzLZGbyLoUezayu3y8yKa9QKp+vjPXwZdw4A8qp6cwVC
NEQWsk5ikkYRE3fKBruB0+Qm9oxi9x5R73NYdaSOcK5GdgKN4jSY2+zQirBgfOWP
9uOzU3Gm/aodlJQfKPz7gxiMpzbiAtZVjsgvEVa6Y5Xe0d45EKwGH+WicEubtZv8
9fPCAXKm9y/FJ4036w5vl2y64ky3cmagpd86oYZyNXOGMrXHH414nZGJfb/7TCzB
QhF/TOeAEPDpDWQyWwPn3yAG+v7coFWQlT8W4GgV9z836TsyuIVx5QrmPJhHTWFm
Bw8madsxszLiOqVe/ogPfmJJQluu8f2mmhuXBNtdhYos+IhAKfS4yVAlDXhmZNeG
R2UOiI4A5PJIzw2UucoY9aQnm5JBE1CLKgAOKDBOYkJXa7G6I8vXUJLz6wpDU6Uh
+nXgPAQKF/Jhn09E3kSHlizV71Bi21j6v73A3d3GDle/7wYDe5PZDz47Bxt8L5L7
Hg+39/+POAh/NdAHe4rR1RmbyhEsGacCfC2rUjU3jtH6GHAb+GyYcOrFMaOvJ1LT
somPWk4o39rdOR4WcOxLqdkXafeR1PysgnTfaRI2eOxOQmdTc5l2nE2R2gLGNp7N
uAWXpaN1f6sD3F+mT0UnBRzXAd+KKkX60iwcBtSxeP6gymFZaMqOy48bT4QajcF/
n23VuC8aKW41gdY9pDVbp51A03Dn4N0DmC7EDHge7IsHB+t+cS1b4Dc1zICBP046
B4xCKuvCQuMcBa6D68LE2yiQdzOj+4AS7Fs+0J3vMLpAg0kGyzVYHwfTvKP4KjuS
Pm63Oi9LNM+AmGEcUeU9MJxppwRpITz+9W9RfhoA0dlZT4ouycpy7EBB0REbaF+l
J2Bz5BS3YchB4nHv9XrrwwxFI60is5LvKsi5ld09c58BR0RBGk9kKp9pBdJ7t8+Y
NHXbVymieRWn8hT7D5YZd3tylxy1kodDdvLW0OQcc4g8Jv0tUScyy+nbrJnExibM
Nc0rsjIv+REtZZPXUlqmyDkOGJdkY/kdwbOabFQ/62tkyEqKY0HSiDYtU/nEPZGK
Kxt9/oT6w6ir+ZpYR2pPkupaT6S6dT+jQ/Lf6/oS3ZmOHSgs2J8XDKfLd6kIo8FN
0jfdIkGTxxdBOMFukGqqb4bKFuSzU2VF3f/rH/5sJLwaecN5Frx7J6TaTzeAcVja
EjwjngPNlc5rfyPxS8o+Xa5DZQimLQLsUCOG0Hldx1KCg245MLog2nCaA/F/eXLL
5hzSPRy6JW19gOpH4ybgW+SaD6nd1sc9/gnf5pYrMHxF9y3oLKEcnzYfikxpkkWw
TUcDmzeniW/PkQ9b/Jp7pp47cDOw7JRzxf0s/IU0mifdwnkcZarGBgSeqs63z/dJ
6e82pJWaCtf01BAnxLWxXuTkfNqthanYjIVNuvrzjqerEgdDMSWBAReWbQHTUivB
/vRRYMWR/aiKxVQWnJXYaWry+HpjyaZNHJuWLQplFbEAsmY/OQacVhQjhyb4laQT
WsC6lgLxuOpMFh7Exd9dS+7oqklg7brmV4cGUs4ZFEK+uw9xGFPD+hbWhDMuuXTi
e83hS6LWNANJFNLsLq0ScShlvDLqKof81u37PZfPRpNB3X8M5ZJuYjPmvqu+0N1r
uwBBnHSkFJWTBElzzFXS+pdXCJYzPGixFiLZbWhu4QPPln5G5ptxTCLmzWQMWbO5
cDuxlyMzx2Hgq5VC/r+e7hqHtjIHRypr4kS3Q+67S8chZ0QETJjbvQrApkcReqd0
NA9frpksWiVkgPSA6zil5aDphowrNv/r5nKISvWA2cNlx4na1BEl/8gPUpMr6C+6
JosEiH4NrJi0RTK8URmW//5u27NGbzbXvPg1BuqsRm2tqY9gwtTvTe8JfOTQLBeZ
gepIvtbBayUJ1m9jVOLiKd+5QYVxKypGMOyzFM4TFP8IDKXgs0lhRAhX3bCC6WOT
XmgBhIhxn9jY5Wcf1LuE/pbqObLyzULc+1VkxUpGgYxhb83R5gI05Em7wowrtYow
0KGtpgApMgmk3V6vR/bxz98klJMmYvphmN0LQ/58TBzqz39qrOG+a7DXVEmJrdR4
JI1OQPY4L1ZeN+2WO81YxlYIkwLkNAlsJxjONL9OqGaPgkm7lVGoSTtnQGq1coBK
04gwBdoXyZ+p+8kUxPFCsTQSC3SAesALkOg3lTD7Ejvx4LRZJdJR+9TCPxcN7lYm
MxjCWcQ1nDJArYJoU+HsQSVUTS5XpcujQrNK0anCVaPhJoj0uQGlCSwW6do+u7uj
wmCZ9MVSK0aRk0eiyh39QCfDDZeQVd9BWEAbYftT+0/MefqKHe3GGAqlG4dBGBqp
hbZODhUAG794efLDJEbo4yobELt2gD5DaXsvOJoXYia4EYaMdBw/3UUY2w/hedaF
9O+rPHcYU3M53D9zfBlaxA7UBBF5PWEOhSp2apB0Qggi3r/Tty92qHaX/LtUbHWc
qzPSCeSvAwfXwnod+b+r6WEZnv9FLdRTs3yA1PG98qw7mJTy+fx0AdG0SO1++2AX
k5K4xayDquivToGCZY4GOY0DteDsHXf5zyShuI26lFy3v4jHM+fIirMglmMtWlh4
fvzSw0atemhZWZy6tLX/5c5T6/jabtc6AbmObuAE32BoiIZ0fooFw1o1fzMgXd7N
Sjci/ntUbS0IOdKsma3auXZWOM2Ly6kZx9Ipv7JxunxB3nAagP6fEtvceRZwBf6z
Atbt/Borfpfi8lotCW5fUrm6Op8qIJfVsvRt/zW5c46Ij0mjg2la3yboZywX2MmI
mNwJz45KEQTybCfA3a+9PbuXUGCNV581V2t9DKmoVdj4o9ICQEMptF5ygy+ICIo7
H6Tl5oanM2DUHIKhaKlESKzYRXSNkhhXKn5XK03kQTs7PUaA5yl+aTtCy3ZS74Ku
WNtVgIQRwphTwG1FYNgFcIUb0w7PcFzwsCtK9YABP5w9WkZJ3l0eeirw6hO3yoIS
CtFDO80G3SmXqH/I6X/z9Wb4Uio909Ft4Vlb5a1c2iAZ5HSin5EYcQ9+oj3vKrQV
DOoHCNKhsSFu70a4rKogN68/BD3LaX9+Nhtrd0A7xYA+FykY0u3352Kbmf621K/p
PD1i6raVxm7g4YeXNKxitQeyfMKi9HqyzRPw+3hVNmHNUEi5JtlsJrS/PRdIi8sy
xztfZSqXdU4sNgSLXDsLZtQcQ9wCHVIxF0WZop0ho1UKuNx2L6n12SpfM7hofZkv
QIDNNyPRvYqwVGrDvHyU/0XP1Zbbx/gvMBdK6JyLFvIiZ6SXUyxFbUx7Rc3YK0AP
FafZ1P3G57mp/twHCzsHnfQV/NmoVig49sLq7PbPrhBJiJeZiPWQq4ZYGrrdA8ER
L3Czy5X95hdOdnn0iC64UtW2mZMjTpvpqQq4NCLuaoUc+14PraTuZeHDj1Eq+WwT
nd7DclB+m0zPySA9Iqcg5NvPnbArH/iY+mWiGrSaxc/mGRUkXBPfMtJef/Apt0ui
mNhK+W0ZRDwlCoQGTg09VUHW3/UBGToYCq9y0Nklby5iEHyaBXRuGFzokssFNzuV
uCmROCm67nALcR4VPKNTrv6pBpiLn9UK5HMwh1D/VC4Y5+a6JSqtM4I413PHtGg6
Z+ElcPIolGGULDjedzqXdMp0aGyCkoeO0+rYMCPnbX3FcTAG48VoZk4oK5BECyv4
63nglecy08sE47EevZfxfKP6te13Lpodl4u9hkGq8tVIfsTYoeQEFeu2yKaGk0Lz
jowylthJfATt0oHQrTPS75vkhLAsKCAueUENDW8FtCAfHlTSKqjS3f8YfDSV/Nah
hl3Fk8hAoBZgCDTLU8nQFD2JVJjwpUI5BaxXcBAMJtPwwkuPHw+2UWrykDvKyGCA
O/ithJjK4tL/2kZGkGJomvSTJoE/QSMdkB4alVkSRCNvZIf9TC/klIeH2JzBinoV
EgOgQt0CHDgrEQXZGgc718xWRweMVJHKmSdZixI6NEWYLvy7AjD0l4xIqX6G68yd
q6c1OPY21iUBBsBcE1UsgR+AaX4dhL+IN31UNa7DaD5WXkgjhE07AD5VrCGvSzxl
dKmSB28+INMI6Rba/RQANZ6nMgrUaH5d2kXz1KfRtHxzIbxUMIIOlwFoMdUZt2TA
rEgHGqD/CsNH3io7KgLXjBbHdBhnQp7ON8b+cY29dPrlmQyFj9MQ7319NBInc8hz
TbooQCl5C+LrYwwAjPZh54kWKagL+njdjnjHCUYPqDqeAeDQ83YEtnY3FjNz0e6u
DwfOHnLBKEtrYzsZVS9U6t1nrs25uQkRCxmREkGvhJFYKu6ReI+wePd8+DGmJCpF
kHR5M0+yZdaEKaoSZkAAJbPps0+mnE3ZzzQfvPu+mUooUzGIX0WDThhv0Qz9pJND
TaVUWIDEtllNxogz8U6oQhgV354hIMsTEh97s6IF290i7sclqkvKltZr5cf6Vis6
jhaEDZCtb3BAJlI/MnFoGL4lX3WBSV9QsI+R74EKXhBMmdsMkLbDANlixl/eLGrk
nXekj93+AekFLx2HDMzVCVBbSo3djDgl8kafFLagEqI/X50wWKLQIooOwt7lKLY5
WFwznzEMNEADUi8oC60dllDW2MvsaLi3/wYxL9SBMtiqevGvNnKhQxK8leqinz5A
QVeJ6lw03hjoTsBEHo/UlJuz/gTFH2DDkVbfZ3Q8NIVFuOXokV8RpjxB/6E4s+Gb
JcO7n4BT6jaa3vO/dvTOHKh8XwaFQ4cyS9dDMGMmyFfGJqbdiqpB0LCXJiex2iwC
mD3jRiF+E9FyLNTSySAkcuMv/Yztf9mZ42UphB1u/li7Zf/eYkHMwID5hlVs+NHl
F071tDS9JjbHKDNFiZ21PMI4OZBR6Ct+MFBDuDM0K0bO7zteoMLymKQ7Ilhz9BWs
dOKBlOA4Qe/OEE+5Fa5/lRjIl0uRv9pzLxMQuyMc6mObw3Yn6Rdn/PQgyHLGBgiA
FCL2Lu9Plw2J+GlvRj3FRNI3FDm48s8iBf1XAgLyS4ib8CEou8L2k8Gn8jmYmZGq
Gw5uNmZ/odoypn3fbKiFz6BJmw3OFrOJHkJIWLTVdtwV/m88lWLuHz9PUeUUVsma
L93KrcGzHENkapyc5RPlufZive1FZHB2ybrY/FXQ75mNtK1N1SGp3BKa/hYhgtnb
EjvIbUTC5GgqvKShSuWqHEdFm/cQp1vzM3j46g2mHpiyhbAm7+TV2I2znYmeZjL7
MIXN1RM8ynblP3NJehQNBUbcImZeaKshsWIJox9GmhhIKm0Lq5rqdiP7WA5N6P1L
M6kmgARmbsE2onQOw8mZquxc7m4hHFfjXYzla2mpLNjAgH0dzxjHUvqvSjGUPZSM
6pfch54/tsf5GkldBlCOQ6qSW/p8TyCpCA6kW4aWDxolSHJsUlxysl+znw98zzEs
VfxrxlGdy9HRK7kMyz+UF+KN6KNS8IwzMgI18oFImj/Zx9q3a9mB9gI8BZOftFRe
FbAm9XarnqhtNmvc3kQ4n/eHjLfBQ+80+Q+2RFUTugCLLOsAxsWBR5QHs/mUT102
kK7NQHUTbCLNwCd4R7SE07PzGJ5o7A0NubANIK1s/qjT9UxQSz0qThjlUa4GeSIj
z6fWo6Lwe+Y8F3YigD1sVTHzqEBbPpDlfzooBUJf121KJ8QOueLBRvX8jFDUmdvB
4TyckD1oxJSoaaeQMfexTqPLdHXw0iA/aVUXzqnpVPnm7/VYRqaxf33D0ZedVbid
IHuZAv8g1bPbX3DrJfef4CDId4hkDShW2uxzMwh+PLgBqz2D581WJxxVLbsztyq3
Fpa6VOaMEyEtW68cx8qTdjB83P25Mizx6vAahBjaWPT/3YbMsx88nT+q0Ew8cYL9
nJU6mCDOaXHXkKovPhWuAQA4AVRaupix2cpLRF5MicTjUo8NTjkjyt8qyRMRp4s1
vrp+Z4X6Jm6tXzCnNoanuipiem29or6loH6sgCshPUjx2kneIFNIMFxO/l+7Hnph
5P0w0jIo1ip1aOzm4QayL1FowpxHDtWa7imulgrAwP/pMrufAjEvQKIERORPiT91
/GQ87v3rCGRBxx8WkBnoBSYGkFaW4UktcoVbnwTjEX9WFaKXcJwkja0onYCqXIDD
7BeoG7MPjDeunnFUjAgztYA/nTNImZjtVju5+8ejto39o+V8LptlI9xbzIbKqAYt
uhJQkr1vB2o4S+0GtskZJRVF6TUxoj6sxWZyVfh+Hu5ialI0dkDGOawBrUNGLVWL
78IxDoGcqGEUT7+QP+mT35EnzKatV00deD1KxyS5e/CimW1kgXA87gL9eIaASTR8
uj1KmWfpCl5YLNfqoS5u7vQQp+svKUURQKm8Lrm8eY17Znddb3yA9pV+0tLKFp1X
4oz9W5+1TG8Gl1AoA7Hl0GC3iSuT1mwHLS5Egwo+u+B9gMAD1L+BMZXHqzAvg31T
JeaxSyTjsm/ef82+sTkZVoRt81YzhL+jEc3AbmDBWX1NeK2CVoEBJU68pD/w4r6a
5UMaYCZttleDC9kJ4zrVqB7AByWmOlzV/i2CLSYMbhxvNIStag0Rjs+Ajj/LXoxZ
6uyvfvSihIsDH3dufGjxuFW7Ry5VrdTTwPu82nwqVF9wZLbOROaYmS7yORB7ZcWb
kz3VN79gTGLD3gdQGFaoNLbIvEY9J6MCCcFW0J+4M5cQEyW/xtZZNLkKop5OtHD/
wPm6NYekZ0GEh6B0OMO1citj/s/bIcfyV7NPSdxXdYM35ySPAmwWqhk49iwqQhDw
w7wF+enbfi5tfFhnWJ4sCdB3gPDLmn8d64k/imgdUaloHDByN213KaUOAgWRfFkI
A4/Az0WscLIMU8sBamHBYiJcgb6gzgW3/zFSgXkVTA4qQ91VXsi/n8L0JxrDIppm
9gRnB8uDdoUgLWhtBQEXv7kIWWbwLxaoM4Wy5d71AGjAJJaNuae4qIMVEylbmjCl
Ex8lANCgbEgq2TuZ0kRfsMNtc1tG8gmkrsN36sxrDSuAvf1X+P1ELgXOIYYsLIy8
j2EW0NcI47b2GiJ79NhPehfQytgLWiC5XSxAnTc/cISAsxaYRBYyMVKH6LJOdrHW
ZshMRJtZLHjM7Tvq7M2j/AgLIvp9+x0NsfzhGM29tz0QgjB/5qUKETd1CxXp/3u9
ewoeahzj6+a8RtqfUP1MRjv3Tu6GHGUWzpuA9JbpSndSUA/Kz5y4jFfNjv6ToLcF
RS3RhSol/HDij6X49hdNCflmlY+K/QwS1+dfNLHzSiaVOMGmP0dqW1kWLSpgiwFB
omi1NCdY2j/O5055YTLQ1t6utc0PfcjhJJuCJYkgqKqgvQwP91MqiUIvmLLjCjps
1tHYuCabjAmpPb1uEYw7d7tdsD4utWgFxVKiFN9E17P7SwHsFvQV637YaPpo/CnL
ee7QpcGe92lW9kQXyUP4dZ+orKbqSVSlirNtt/bQgk66dn3s2aUyvlJyNCHgbfpG
xrA5U/lREMeQDaMTrqR3FSv+ofU1NtM/v0WjZ59CVhs2TmQ1Ang4wqSGmynQRK3Q
ct1UKUhFCqPXN+35z5Z5omvq9LtADVRqUvTEQSVird0jvnywMJgfgo32+xxWTChA
Sikd98cMGEcAtm8i7kzfwU7Y+/WyUfMiFMjy1n7uPTBVDj4t8Jd+wHMAbIFDK5eH
3RF84YGFZ0WKyehsOBQYK+jetjXuXMWbcfjAUNQ7rlGDek3OwQ6aNzr+ynbYPhB7
QGXgFXScgHpzOJqKfzyQ/1XZWACV2M6l6NkNtkcLPtmW+iRi9GfFCJZdEQ28JsIX
MCYFl+WTx8ZOxufgxO1rqz9M1Hb9QInw6YKFXIBF7c6er7EqImY1zsSPydgHowls
4xDxbqLGbO/v3NRq99wyvzFAa7a1jme1mK7OBJgXMo2POIvgvtQhyUcT2G6jdtjH
uRuYPBM4qhVyvsETZqLU9ybSOvJtJibuLuXVMHMJyDPSmL+Ki604aYJ2XXPR6lcH
inG0Gb0IgHJvcbg/yRZ38VuMMbxqQwJUURTOi9PvZGhG8yVn4EGDlqvv3K3igg3v
2O0bC3w9o2iZbtZhR8sAItiT39lq++NN77+w1C6iy6y1Fh+jZNJbUYaGjI114oKw
jSI6TAQgur/y7Ep5tOruJiVJKCwrL9s/ZBcB/6jm7vGsxIWlRjrmv7TM6bnGgVy1
FcfSFieD1jjK4Ez0oJG9w8WppGD5nkBzZiZJzEzJMhgNkDwgyoewrD8XwHMZV1n+
bpQHPfD66QPkGiwM4qvGyW/E/iBvvD8zuPt9uigwajrAxgDAYeHxt9w6IgNtNad5
2aDa05k78bNBB6lJZlhIOB0zVxG/qfPjf2Gjdh/VPV2uzEoZPG+bL6SLGKiaPo+I
bgTEpopc+NlgzGrCH8bTz0Ttz2R7Em2LVZLRasKUkRde7uNYIfPixuSc+T8UZ8Mt
dpUSmGc0RsIIl7sqFewo/biRcaDi6Ce9Q8debEZ+n96Bg1I37VtHS72WrSWEOXyH
nsO7+w7FAHt3Q3dCyI7rwBYwzeNu2lHew5fER/XhgiOEao9T0y6Dqh1/KpvsvkwY
lycdmyQ5YrhvnGBcdB9CoUt7uz/0Xp2twqheD2WEovZKOKYfgZNgUcjqa/hqvRRR
QlSYXbI/h5/43v41cmvEKhVcNkaXcs44qro9B29yej7N6FaW7e0/WNxJN20yEFIR
O4dm7FajxeIRokRfYagArKNkbcBxy1a/eNAdrde9jfJUyNfeUMrYDtMZvS7MvAkO
aBS4/ddeAE8xmb2T7hCFS1FXxsk8dSLtA3Zg04kzMRn/6NX0UGyEQmRIyFK4wGFF
RgILJenNLdrfw52U7Y7R+Nr7rQI/T87XkzYl+AviDqCIQRIWaOsVRoflHW7ihkHQ
N11raiyxqq4kTHdHEP+6DJCqID0N45sEuYNhMSyHTn2f8981dhMadSYOPwXlwSEW
t6RkOsCOV3d0qhRwFQPlaluvdSMOQiF69H9JHWtZFfNPXhbRrzxbF+My+/f7uk40
iYfXljCM3zroZengUR/EnIQ3pxPiN+YpJVn8coT/V9NNs7tcXewfpUh8EDcsiiKk
BRB4W0N1/jq4RRwYXA/byXgI47cM6hSdJ1aPjNGxE2FyUfcVjMJgWSOUnTODI1bc
MC3M8PRlJzyPwmp+OcvloCsTeiirY73vqsFEEgfzDinsEcF9EVJ0WYWi9xpTND/K
3x27CfnBeg57y53V6auRjYRdG/JMX2uR9PuGKC0LF8JJt3+BO3rR13aXIa/FN67x
eX7GuExzYonAsBaNkJXV0ILYOf3di1n2Dn8WqV+mIawZ7k11vvMV31qpJC3gx0Ul
Tg/R0IMWp7hzPOCUpg+bluh2wPDwGadlvtrd+VxPU3SuViB7Z+FakQJ9m1eCWbA1
eJ4U66wWsnruFHmH1SghKs5ioA8DEbBGNsF4Bu2x0XZ+ffyE2Ve5ZOgvtSr7Mv2I
x//He3jRv+jDsE7wUOde7EhMfRmVVFqkpqfI8JKzWP9WRI166LptvOGLUo3QK939
tuOif9mo3pgilx3tGO1V0xvA+R54jckPyMg9z4tFlggW81Kt612qI2EaWuth/FfN
9mw6UFVdccdduNMa2S+FQDVQJFqH0C4fdnQu2XNzCefU6FsTFbt4N+TjLRN5XcIX
7zv5HhlPcDBfYia6pC/B63Aywf3BmACRKjpfSc0YslDJhQz2ofY67n6mBat7fYvu
AU4gRSaFt5OGa86CdTL0FCIfFARMBBPZ7K+TcN+5zBVUDA5g1WI9NwCBmVYuOazy
1ZXzOk9dkX1GRFpPjgg3hx6pzMh344jJmvMHa81VYxI4BYwkJk7rjnFpR58IpOVW
3x4I9hgkWhpz4T6uYPtZmqyBlyI7Y/NMW9hf4EXIpz2n1JCms+iroPfQuuVxwZ/1
7jU/IPBwkzZFIw3bfX8hlEI3vDzQUJzV33mroY6AlYCLZEoejB4AMB30MRoAkNDa
hFy6ffhIMOxy8PUHG9QKSahPSxohJrDSt9GR7tQlpsQFt8RQvRFnY06NmSIiDVFH
sZVlRNgmAH3xM4duR6kKuLBs/ZhkxuGSGTJvejY6BP1K2S7jbVZiuHLB/LIawjOA
Sxsh3fKZdhlzBJvW+XXdpF2aUqkBpDx544qw+j7/UPpH8/hJm7W/XKq6JoezcSo0
TFcroi6Ar182L3vHdsihqZ9aIzD6FRuPJE8vFvWkIyvAjWsDJJTXKqKQSr3kjZNM
Ak9L8gYmmlL0SwuoRSTQBzxVDKzweFo6HvmaEB+QpHCbYFvbf/GqObie+tUSLG0R
C4h3rPswtRlfdoy3qhFjPPAwUb9pGyzQY3OmYie3kjZRauaeYt/aWajOTr+nENwA
7iaGRSSz74CivQPTorvXQmYg+sbsz+s8pKnrhDjyVJ3y7ssT1TCUj7Eb4MS+rjKf
avvWZ92e7BGZPULycHdm8hGu8trCA+7jCVbSGf0IRDRpLO2J1NpBDInzTCg0hS98
3vk/vCVNe/gCJ1UBGu0Tf1mR3saSoEK169uSof33cgBJgcZV0n3JC7Ajg21rNMh/
3DDkd6lwuBvKvoRZB7eLx7YqKBozniw3pLD6NnK8el6XpjY0AGY54Piz+VjzE/FY
9mfj7hT6lTP+jkOh0AeRwyPNTONNHzU1AhXRTRWzbaae/IPuN2x2v/sgKYPrwJab
xBY/adzw9UJlzzWzo0xfocO32kyQTYOCZEcM+uzXmEzPPhid1OwHjmr6lL8O1R4z
ftnj2UbhoOyiy1pEY/HlT2CP4Q9ToHuiKfWJkFOJnPzQn7xHJHbxb4JtnxUcYito
iKXMmM/7PcG30qLN2Mhp/fGkFcBvAch5bqmQnD4LrpU38E1GGAhdOL0gBp6xXQLr
vQl3Bh9M//rwaKDEjggZmGpNYKod+7sztb3t5yGBctDkkTmqmYNci0xse4aL1Vyd
t6+Yi5ikbz1mL3u+Tb0D/GBtqdn90aQ08k7qTrbRSdbY0RYoCW393ggNwVZXTD/z
6RUWNC5zE5JElX78Bbop9wnjWYXe9kVnnhEEFhT9X/TfmJ68V4ZxLeNRTFNy9FXT
q5ppZwOPJG1LnzvxtNkGdeIYCBctPc5tzVueBveWPjycrUbhIWoeKkfVifs5VvtR
/e9RA1pxJMM48d70/9arjRsxs9DW2z5kb9V45t7HxF5JiXmgyCl+tZ6+FlrOuWBf
S9qlNNvFjge4E3vdhIal5CHYw38iuRmdjJSPhNeAlnfR6ZUPI4UNLL6I9hsouRLu
xICX+Y4fkgWnM/XBk9YjiXSToh47QUMVhPeb5LBNZPDHF/Pt2hiaUmBsCA4ZeobL
fJluafWURmUUTp1jduRUlJAq1sApzc8cICF3se+5xYvP/UPGsNW99Q7SZ0Nx/NjX
H0pYTzh6oAWmXGi3GvOT+mFeUaTdSSe+D/BbbJYsE+77Hr+LmZcgdU84fc6AbSAU
JphxVo/S39iEa2FgTKJVrwpoNtHNczt4CYwYuqjRlkbgEazQRYR4pQdjZ3IRFPi0
A7CigfMUQoZ9lVSBiTxydRsbnr34BYmYdHHlzFsiOeJ19dJOMOuz0GZ/dTFfolaU
rkzQco8NWIIpJPWQSL+HCAqQGxPISgOAlMAMvOwmb9VyTRO+duVQv9NT5xwyr683
QsqTc5DXRV8BVcze3cm8CSrgDO9kgI+fiA0/MJhj5JaZbYBytY4WOyYRXHIDbZlP
idhwmuuEqkZ5eEYB50r+rJds/+2e5nDUXjSy6RZ1idrNp5+jtGpV4T3dGrBlnihr
s+tNLWYDYZw4+Tm8dwj+0zhA1Zzm8w53mRukl0Q5zICkcqyJx8PGKo59ULJ5Lbfw
cQqfoH7othZiK0yX6HKPp6uhhMhs+VqRPq/JQtRCkZMk5dzZDGQqrCsAb21Q1qUS
34I6ukytG5OHiSrsVQioQ0rFP4/j/L+E4MryKU/trJOsr5jcv/lPdJpWGQEyYoFL
BY2yfFWUdt02R5MxfVHO7rrI3HTp+uZL5lIRDtkgi+rEk0C9XYT2Dk9XGK/4tuo+
jpSzNUR4jeAHC7KgtPdL11dIjonUGXbHGj+3co9tu90Yb32pxaBSqHp/A772E+A5
xjsR2WfaOhgNgC0V6wXavqiQ6fgsXF61g2E9UBxWX/qhOqnDGYcUjNdxWsMxXmJX
upb0Ff4hm5jEHCnpxtpLY0JxIg0fItEE7WrEwmAkjRk0/TFrsV7uxyL4ccKM798S
RJ7TSFW8HggePbqYF4Q8gtXaTqS0ftbgR2k08MvF9zBEjBLnp5Rlx4YmLKFJCxzX
QRAv8ssFwP4e+5ar4ECXOC/io+P2by+0DQGnb1Nn4365FqC+zY/sIRy/nkhtiQxo
PXPcaIuDxkz+fSkGIsFGIuQseNOBDMB8IS9g86s89DQF5It64X3TRu02OZX8LYza
TqC7u4seQJCnF1Ls0moGRhox1EqgfbGtA9YL6lWPIzQtKqDKdfhsJzXWN01SMhwc
txtdz9FAfVyIAvi5rNmHC9QY+8CygCVUJFzoAFuJn0yQLlWzs/hHY4i2W6Ns55Hh
yTNyU12xWBBQGGLIHapUdQQB0Up7AZuKnoYVSrK9MHG8JTr1iT5zZuZyiCUXjYYm
+5fA1Mja0ZXDmP/fbjj44LxUJWXh8u24VVnTQXJ4IwpZagEDoqBKVitpF+HEjLfB
XKz82fY20jUDMkUzghirqGNfBFwrvYISGCOtXHeiZjlWLGcYa+NjJ+1aTfXUJRqW
sOYKkYE55EZqc8tadRq+E4lrzsUSCp15gmEIyWBL2gxUAM1raAq/2XP+lfSH6YGj
hg8naNz18WFF2B6YN3mMXdqHVeiHAhCbSqhYa2q+8Cp9JTZqNMp/Ud78nCmRAKQp
gD2CWyjyA4906OknPRLrrwJ+sNtcPM8+lzutkq3SMLhovgNFFB1NYJ0m3V4AsZGs
g8CHvejkwCXWR71pM5EErNbps7mfbVDMgV3acHUTBVDTDkuvCg5lERzZmj6nRB4m
LZb7S1sxQLeS12pRszA+p64It8UeD7l00P63GEoIARWYVw7LOQxe5Ae/TJKArHgC
VzyNu+F4PmNpNNGxkg3g+QKSYVeuDae2eThN0Vh4KgejlNukGzBs4p9vPGO6qOja
y2Xf30sJKyI3K9EjfIJHDKrdG+vsVPlrk6ccx9klI1D1HB6MS4+DoiG8rCXZBlu8
TTOfuUryTbAFfbcyJYTeQgGqBSX6TedEpGKHhpaqC7LwMT5+NWITqUB6vgH3vnBx
NWEDMphsnYJooumYi7yjsC8l3GXY0B7QGFO8f31Wz6Ee5WtVu4RKxZ1CvaO/ohdB
yld4TiHAKO4tv7nNUfqE6GsKcXfgWmRVtnQDJMiWvcyuCdHAK5LmbNiiNcGCal69
1nO+a/rl7O4EZcXShM78HHMYXL8TOqEwnwyXS5nWusqDN3baCcj5xCGuBJmQYzOQ
LzTgtC2xFq8X19XnjxGI0HjvbOVcbTX+Tly4XtPBdiea8Pwl9jmAyQSv4xTpqTUc
BB2rlWepST22JCmOEG07cXxho0EsGfMQdqXOM/Xqh3EdlnO3UVWa95bLLr28q7NW
pIT69pu+sNaAOCsOM2CYimpY8f40WrXT3ctHOuZQlLktMQMq5wyMMQKqiDZ1gqig
CYChnjJ/SrwHX/urDIFrvDBV56rzR3M3q+D+Ev51Wq+TajRd/+qepD9ZKX4hms/W
4tw7WfOlCo1C6DgjS1hF+M8WGZkSQzgnGL2gsTbM42EqbrBibPXfJZyQERMkLL+3
lepc109U6OQDBxP+fOC9zv5cXhj7pX2FWCtFDJHQ+hHsiEbIWSqm8ukh0wFlPi1k
Zo5Xp66o3YMb9qwERw52XJkUPB1qJMznyrSC2ZuTqe4cy7YWMvR8Is8KqNho/rUL
rIeSyNUQrwWnzdtpTeV3LkCP2dJn276ngF8Pao1CY4c6I9RodGq647dUzT2JUS21
1sdZeHRzAEQ6Z7XRPDhuIHHVXheNq5xWDbXu7PaGf2vxGF+YC9Aid3vBOXUmb1E7
ex5w2kRMks412sRRhOZgQ/eYHsoYyBaY+gGcgvcvJOEDTLl6XrjoSV4X7xSflsEp
uY3p6ph4k4RKxnbLgu/T20U1K8oq++wf+sHk7NUDo5T/i0KIUIgF4IVkXYulxTiZ
HfON8V9AsIGpO0H8kAlZ9QG1lWcCCGlLqFHPV58JoXL/stkaCjuvRxjegIQRaafl
NJ58C/xs7WQpmk6ueDhlVdrj/QoFPAKOchE+e+jSu43Kc1JZ3JM+Gd30kFuXKsxs
EyvhRVycf+WXgId3l1fLiXrI071pbybW2+Uy24nTc+4SNzqd5CvMsEuavc4dTYZX
5APrANiDNQ77gStbyDWWv9CEcXDkS2Z2RuTtI9wqQgFsyL/lm3OiiSz0bfkFBv1A
vly0JJFfALNmdJx7Y0DqboXHKrmb/sYBOplLlce9k8gcccEvE5Z9Y4ZkoutJLqzH
VNznyrvMFukf1byAknNeXqmplwBYrj1r4yjcBydptJRqalp+708QKKQN6F7ODuqt
oPD6rhAdr2UXARo7I5YurYkW6GO4q9UdJr3Nzn5ZxOlj0EbDHzCi2/5Jwr2Salz9
l+Em75NOpovDtCpN1AFAr4k5MtCe5bopDv8GKc7gwQWBG8xAC71ZdxdM6f1cEiFf
H8VKgDY0/CCu3EeUvMfhPc7L5RL/88/8aJjAuGEgBUV4DcqrHPfyNiyNtEs94wcB
/XR9B4+bXivYY5mC+iUdeuUHC7vNCWk5ZCJsuYRyngvx4+nEFVk430mvCN5V+Zp4
fajhD0UAYH6JECi3MkDOF5ltjo7oUqpIfWnONtORZCv3GiSBXUCA/ZAlrf4lGlUP
3oGM1kWlNq9XXx3ssdlPYxZgv+DkbwaWSSyW6kj//urjM9yxCl0TnIvTzRnOPGba
kzBsrAPpgi1pq27WJ9fAu4G4JD1t0uDUNTcwnqwcLJVHdNSZH6/x8OPHUhGBzyfz
LUOTymN8glTEycUbeHGpnzNbb+TsSSN0IhpF/OlaYGaIr9330lvVpcJvqL4QymnO
ti+Ule21a8TVXRfY3I5AuBsRwH1McmOc8e2RzgbXGtSYtruEl2ZRAOpBbYJmvnUY
ELeFX5xtesWHHkRyuwUbQXq4eRvpyRkgjyVn48p94Mdwu7XMxlrwYqv0v45H6IQy
isZEoap0t782FsktM9LZo6SOSB4el5XPbCi79dyQvfjwWvsQVTLra/dzb9vL7Bwi
fNaGq5uG/XhB/ewosZP6TqSa8A4mknSmaZxTY6bVtz6PBVyH9TD6Ik74iWzUa3j8
6XGt+twJoyl2PmowbrVCLAjaXBSGmITd9GFbWNCbe0lXgvsFLhSg1htyKvYMtePH
WPvpd343HhLHzrID/ZPmMt0ZLAuMA3WBG02NnMBxLX/NJxAMz2DJdEHi8xyEvmz6
qRW8EoSBke2YouvqiEDYaeZZ9sWVLi9nSRVszx5gyv3DdUDdyCSn2mukiWIJQPT5
fztMw1tN8mCCQxQzzoyRW03RMChmh/gbwSlkZ6XpQDH3Lxfa5zbWdriXjIEOTxlI
dgyK26gu5NoTa6S3/FvSrCo63u8tkICpdeWhPDJCXzkYkM3QhdXxf+e5DjnyQYJ6
9W/iErRhSn5rzAQWpSNjVA27u16tg4QydHNCq/6JTpiQk1i8XYGVXkuw7sGYdOds
XciTZGLIE+5bKZVC7Zq/pRdqF1uNEOvm13/PM0CTV2f9kk8E7OWWxxmvw9tKMgRJ
nRTunK1U8bggR9URYQ2k6jHqusF/xbAN833RTgH5u4SmO3av8fayicEzgOlQLyiR
5BFNKTHetydf6B2m6iu4em0+gB6dW8KFm0wz5eazB4DW8uc0N9RE36VSMR3ACzbX
cxY0Km41R9aDeL7r/BkQlHzVKXBAekpktZMGJlDWuiuK7uFCmJlXwl27KfHfLwj6
dNoPbDkx8c0ETSzWGVYwg5+HCXgzAC8/VhFCi/MAVqZOOYMgav0DtpYujnHZrlh8
Sv2Wc9r1EiykxsOIWc24gVgS4Jj+1sNw9vu+ONElzyMSv6+F+3zYFWHde18qxzrs
JP0zZ1TMc876nHOrJrtJDeLwafBsPsMc0OgTybCwhE2Qhyr8MD+Xon0PGE/90uZ6
+j8aexA/3T2S45j9GqDKB4Pwos7DzwI5PCQI8wLwlQw70vLwZG+4lsI3NszeCUF5
8v8ZptCoGgXxGgAnDvZ74EylLkiAh/CwCuoRLHmi9ppWKA7FrYG4SBpF1xjCcwRf
T9hPCDZXDDIyUl88Xu1dOgmK2JJZcBEsehZAroSvD6G9mMPCBzHra7zwUSD/RI9S
1Sha25xf9RkAcQNWeI4jXBtdXnNH+Q2Udtb+HRs+OLzasn/Z141lpPX5FUnSfPY1
C1P+MTowqEkttEWcdSvj9dIGRuqLOR8OcY6EPw+zxV2JZNeZ73Iog5CXIC7a7Khc
ljtsZaCqZfIo6gClFJ5aJ4ehNB3orqvBAA1f5E3wvkx2DXf3IPZdmk1bmTsuLhTX
dMzeFdd2y/c0GtNYNxspnyUX6iWR4Gj2sYAPBqJyeNE2bjDuj7b890JYEECyYcMt
1djVyTepmtmWLpE1zNSZIwSGekyzJpqIlHgFwNEHKXNSUSAZf4wsgaEBSkBwmuMN
yHg9upGThuXN8Lar5RC8yycPt4u78MDclhcL/CrKlhodVFsPHv61yCy9ayT6mpfL
K10Y6O2uCdBcpagA4gTh3UbE9QUwWL8AUbOBY0Y/KVqBCyNfFnq2EQLpzYuE8Ryf
H8Z8iwA/iPsNIrKr6LjSR904+FTXEsexpf+61LhzYTJsV/Iul1lXnEBaoNZIRCHm
LeWNNzaiKP1FfNnff4RnS39oXTzgluIL9Via0pLBmezxycJMy5wHSlz31FyKhoGT
8QlRyWmDKLSOlUrqCpyuMuyszTFd+IZY3eprtaWWUOpLB6gxctp5hCo6wP6Ke6dA
MXtezPqZ3hGXSmOdqamx8rhnRItncLykiEU8C5yzmBDIX4tIQOkt4EANdXVu7TRd
qTzH0FVXZeAfyM2IiVYiO5bYK34/gJu2nigk2MvfgPQwDqJR9cLXib0Qi7N9kTWp
8tI8QNP9AQm7sxs4rerHOy2ytU/oTaQeUxR41TEPvjBlrmBOT7Y5PNKQIBBESOWO
Zv2XsacspWBr7YkXzPKn/hsKMsVVs8msWG7zdPoCOV22KBZp1IYjL62Et6I2a89t
8iCd5iSR7AwuLHM68Uz1dhsxrBB8ngJoP4Aiv0wDAuBC4ihD9EmObYmAA5KhLW2n
3wABNDXJmb3Abt1+EqGdYHeAcTGurf56f7SiPoVIiDUGfxb/XJtD0d3ve7Mu4iu3
+t1Aan8GEARzZRZVM/npYkEZrsWpIJRaqy7zh8oTBBC4jVOJeMbDrxVt6X4luf6U
tY73XHfYJPrGUXq9Tcdj2FOD2f/weGgoFYTbraXy+sg2q7FBU2vUR8hOoL5+qiXU
8GMKXY1v3FPoP4Dtg4tK7/KJNI7zqA8IMS+3ktZvGcFQtt6AD1Hfnw4CL3CmFrzP
xYpXRUCbO1URLObs/SceXTF4rzro+qaqM0A+LaAb9kS/WXw4Y7xpO8p85DjOtOO5
JF9SIH9fwBuf1CkQTsPfLueHsdFiBtKpED+8YDwAjzhtPHRLQf7c64TaVYD9y/BZ
ip/td4GoDZwvO26xU1kIG+oSK+VTh7kGZnlB8aMToz2URKymm3YMGeiN/ou+8YJA
Y4aKV0FEQWMLFxLVhNbtF01kRFsQx4KI/wkGrtSqKTy7Ka+3gZVXj+kXI7oA+WK/
pOJ/FKT3Lw1ww+sHuI5Dmqjf9PE6xhNsf4dZdh6f0pmTTwrjh86BDbLGT3EZO2ga
6bSIbp29vXroqYcuNpd+zOaqQ6jeoRnJb7cLcVYw7YT4+HP4P5mEPWK/bnBChb0I
Rm78xFes7n1JRUOPkHXgHGnOzRJT1juTjUAeKkdNO7vDvWClUfkkFsPWE8nR2F0w
+nCoRuta+41Q+TNU7BjrXgFiU8LnD9lg2mgWG3Cr6U2PE8bNp5S+ae+CvIF/g3o4
hJMsiX2VUhGtn85oICuVVQRS7A7xv+P7H8PkfhpLkofxB0qXOzkgn9aQITR57JFz
hCr3a2kxNC6U+dlkr2Rfvgw2bS2vle8twiK64A2r37snw+GVloGW6xxMM3DSXI1/
hAPw0eCP9Y8g7Yj4LZVzNFajupRTKAubKg3MVlSeC4soBkmg30zBIvh9ChWl+oXj
/GvJjfWr9jyZpo8JkD5GMqVnNzCbDFgxfniXxJdhcUNCZ9Sa1j17khr5O1rby3YO
bhBabBLbrjYa1DEWrcp9Tz8DUNO8uht0Y5EFaq4HzaTUeBe4YlfeYQN15jpJ/F6O
wJM+6eLICKQGqil+Be+W9wiYSvqPUIWD4JAHZ+M9Muh7qt5WEl3hw5lfJOJMF/mB
rlK+TVz06J6U65NKPtlEYumZH02lieDMsY2ecHKLD14TsySAulcy+PeOwrLirrUT
qm+99+z8jQ3nF/ijaHG02UQIdq50+xWdv8rqTtYxd4eA2gHnYDV0D3QVWNlkmuDH
PYT1xkjR6dI+nfE2GYsravMrviV4F6yQ42XXzLWHuYoi84O4TahE5FexLvyUDORz
p0wS7AQnMXz2OOL8bef4PWbAbcVsp+RRfZmpcogLrfmuMsiBWFiafZPmM88e/hdB
5rKAP1gPWo8Ce/Ev5Ae4NBePZl1sgt/yiw0+77/rYfK4tx6E+qoSlRKdrp4CcLeO
Bzl9rKJ6OjwDuQGJ4t1p4xXaUii2TGIfIXMcB+sYZujFkROw0m08OCtFFCRMFobZ
3p0nQxIfWpSOJRfCdu3cUBXzv4bYrzUnu7EpAY63A+P4q3uQ1wfG5jvtFzwEP/Dm
XEp5bpncWdt6rs5hAxxuoe+Z+WMqyYISnEjkfEqM11lU0eDbvEnviO6ssCYFKP18
amAc9YCB2t8ZZSL8w4iw6pMlKcPIx7HK3bbWPLvJPZWEnG4u2q72O6gqAH3J7sr6
/VUzvbbKIiEA5b9XDG1LA5kE9kwd0nNTHgFwd5UxpjsBuA1ic9wBwitJscUsyXgh
dhZE4m4aOci8BQP1snxnmFSh6lhhvnBDa7bVzaX64adq7LG8gK2j9lI7PjgxW30/
8dey9xtmHP9VoWsTo1lhVlk/X1Eaa3zUEY85hZID7LzG+BtKQEla2Y0l9HyLyo/z
NSao/iDv8XPHAHXod7hVHZFunxJ/cqYRqw3OxfQaTtxgDpF4iNTzAj86cPe5LNAs
r9CtwsBczKXp09l6iAnj6CbAu9lCBThYEfOQPyGyI8ePpEFJNXGqFAvIfisc1i2d
yXB2lBncrihYxRvBQZgXZnXhiLyJKNh3eqGpUqVGeD0sOOJD+KvqdddHZFC10PST
+cUqii+VvfoKGA8rhKewpEbYjmVhKEoGKANvLOQxjRxPodDZS7DHDioJiPcZ2E89
3FPbIpktCgvrw+DBrvAgdgJcMCCePEv9JDgAirf2JzZh6CkzUjix7S6kAXSEKW4j
hDSviLmqjcc/WP3hGyoAy6sK9TLD9rdGK+cdXPcG0Xwb+EMg4whao6ixV0BdjFgC
XVW+AwtN+NcbHw8UzKZWZBcg49e7NuIhdLbWgDR2aGpPev4MeI7IOhnYl+oL//fu
ByeaMIPRFY9d4PqAvsh4zBswf4IpqbTmEPrZcNIEAtW5Rcqd8tY5Wn+1mvb0fdSI
Wmg+iK0dLgKxkpiErN97ZwVp65zl1wvADuCR/cWrKMDGf335cA6+MIbuzq6v9Sbv
nF+uxq5JlvLNOuk0TQc0Q9GO0n2rxYwG9P7NyHYdDat6Xv7hSmFlt4+g6cqo1l8F
9qwEeRZyGuYPl3dWhLFKxx2/xs67hd6nFXbhXA26o3RIqf7I/09AYBQrNgTbbAOC
MdgCs+Ac+rrqAxhiWag17hPOQxiRDiwbeRVgeHZ8KmTf+zE1/UF+fNZohOkQDfhk
00o8GZ0eVbiG3Ihh+ykD099KNHe0LT0tPLM7GJ9RECftFfgcS0psanUlrU4F694J
IYRL88rrNLWwdDxyPWFN4NdY196IuuYfO1DKPaIm3TEG63qXzzviUpL+rZMDWlGB
brv4d8pxUK+hn/1UVozLRi5etaGluiPcvafNVMReSXP1y3rnc3aKq4LZ/fs5OQi8
DPnmP8mmSjbRu4Mv+qJfErSTKXNqPB4+X8lFOG5bJ5DZd2SYr7ZpGaHx0dB+DCt8
ZUFpQxTh9ELdv1cqieCohZSMVDsVIAu0XTdocFYSUMY1XxB1SkJQQAF1U2nM6K5P
73Bpj4p13/SMSFCe42am3WCQL4m5AIpQX28GPViGV4Y63V6gUUFH9L7/72lg9a9R
a76hzfZ4hIYbuQpWZ4CmLJNEYEByT37jJu1xM+eW0mqgl55TzuCjXwXACwcfB/xY
zSWcSJozN3AZ2ZeKX7EHLqdLoxZGKxmwuXZ7suECRiZAv2Xg+dlaZfyCksSmLn7T
QTF2usTrdAPbZfcFKwzUGcW4s+NqFBBfWv/dXw2yetal5A93iuXBWMpJwFzM6fNW
jUcSSRYeVyqVrELtC88ohy4agE3w9V1FgWNmylMRfQg5skrTASOvIxrbfIlCfp4D
475ZTW+M7EuAbrsYvSainjtn1NkOJXgW5YF5O/uPpIcUA6aq++a6lCpyHiZkv1Yo
NoUvU3sm9GeXIwFhl6KD0Lq1oasQlSMIrpeMG9pgsDjDL2x7e2NMGKleDdCIiM6b
ks4DhY269EWnDpnrekeqyjcLVx0++FL7cCXkU4dui9z7gYqNmiFJGzC53nLueSjg
W9T32DYTOQAc1gbO/zCl+ornXkVHTfKUdHKhifAbb8NwphBLO9cgqTgqKuEezO9J
K4j1RJ6M3lG4BnB5zp/561lGHubs0hqGNXWIi8nsh8wije8upecXqNt4VY2T8uU5
TVJwnYLq1HjtGu4J+p7e5/LzZPhoLPMK1Fh2dYPNHzk+sxLsZFvLpMMRBsoTl3ez
2bqX9K4X9SjqByEy7LZMy+hcs3uePlnjYFsUSXEfkTfZHfnGiUCaaHe9usJusB3X
t5yZWKVvR79Dwai7VAuEWWLPlrzejJEvPUo4BxdRVh+9k+3JKINHnpD8JLgLlg4N
TxmvpT0LrvFevtl0fV/MsqIAFpbxWZTZwc0z9TqyFvewDONsNah/jZ38C1q7cLwI
Jh71z5nX7YUtNZi67M9A5REzATLRsLc4OUKx3JmvzrbjDhi4kbzFJ8yToJ2CZtPk
fM1sTFqDviojUBV2rAAgPN99zlw3jpd2PtMeLLBrWvgT/PE4L85bc6f1ukAsmJre
nR27ABA7cNGchZIB4VIBgL2piw4hLjAVr/ptF/d5C2crdSq2Fc3e8EOZtGCLQW6R
AzWLVfc/qsCFUvCRVfJWSJ7//doAo+rsbac5fiAT2S58o6vSfPw9v3Z9fzCxLe6+
bPuCgrKFbBNxZNB1waOQhbCutnvMUM6MEgdPzoRujXwHp2ICas82/bT9686bw+uW
RJFFW4bXMIpiUkMoZucAhWUQriqjxUUBTRmE+EtTsPRAj3VrOJ/BH8Xt2quCoQ/d
rj1N2VU5FGvrZurORD+EeZm3yUuHb/J6C6u4M8Jux+a3+3OV+IrBephYXbHNHn2P
R6eb0nVYqTQ1m6mnFFterB9avY60OxbrcK9PQRFCAQJ6oU0VsxjdAfx9t4XiTAs8
8a6+diPKETfuOMakx9DslF9lNDRAwFOJuOAsILludVSUH8QLNbap60h8x/JUpe1X
PVtclhmKdKX2bsMN4TJ/F22bswUPkMt969DO6d4eYTRdxOwl1666w2fiazFcKxGH
JO8k4REcKKr7qpy9zfYYYXv/ySpeiGmCtff8F1usJMfQeAapl6VlsZ3F9bGPfwcr
tbTwaKANPa3eFtNB5LUgAb4aDqaHjeotuM9hcOXltOIrnl1jThtvLgstIVUAluNP
UQ6ONqHlPsawO3fAGKuPoqk5JyR5EcMByVwvY/L0EPQk5/OT2wL0iaW7H0pDyKCZ
bNr9gMlnEeuS7+ia7C5MHLW0q3tJ6ArA/mc2mm0bATJqhssq/iRyQdo96MkEU8mq
Oh5/8zVfrPJ3w0g43w1G857XXB12clMmVDFEZfOPDm4EREq7bPucsxlctxeU172O
RJq4S/3k1+Ur6mdyiOFdSCMe6n/ayegvVV4cRcK8qWAaXPs8ZXuZ5FOPPLjR60Su
nlPmt9MQ68EPRBebmxkorC3fR9pJ3c4dKl+oMLx6qVVWpSM6Y1m7cnDG87OOcELW
Wkd9TGcg+6hLCASr7QtarjleuxOzGa6m7pPrOsQIgwlLQYDywmYZX+SwPCMx0kgi
d96SOkCdg35IrsOPzQH/aVxjhGd0Srj05BGbJmVLrLzATcbg3qeGkFfRbMsXqNoa
IfMoTfBb+O88sTzMuSBpmhYcjui9OXuiTdA3Dupnd6Hr5yu88fo9Xc6VvWd7sPup
bsZ72zAP/L6Rvw8PEkKgNREStUon0dQ1L+aZ4ajL1jzCCRR3jzZX4DXgfYuf9irP
49+CNlDnF0u7Us+HXVvtnyjou3G7LpXyF+3EwizmsxrO0RTJhnB5g9SHISj+nNpk
qZDFaHiIG5T1drpFUtn3v0m5fQFlgKT9fwD9CekmjsxgCU04sZKbc1TN4OGM1yqw
fUYMB9/Hd7Ct+yCgVLxoPZP0KnZHrknygax+7tdd/KhEP5nzCq0kOT+oOZc4v5HB
8PM7RTf08j95eKI813Co0L9poLS29KZnxkCMplh6MQxCQsTsSiHK1c/UPG0TqfBe
EaPONoyGq6eHm4nDfj93wTplabqnS8pozHUuwx2DibV/75ky9YAvQUODcfdCML3p
raZkMZDbrQJQEDoGElTJubN9dAQCgzFjklw0IETGgQrX7jRCH3vcRWcPR2fMigM9
lJJhRWh6Q76z7ltt4lS7s9eGl92bTx3CneLaU4dnq9akgDbqe8EuQ3+H+bpXfjy2
c6aOw2HWWjK/LT8EW7Tr3sTAeCYYOQfDH4WbRQPuu8dyO6E/uUicQA6gtYogGv6h
Dcf8pjUf9PidbnBsheQFAVvMy7/BOce8gJU/wBpFtPzgkvAEepq3CTrtuRHCxF1v
BBcR7CvKAS96iN9zVEtLOkmHlt/n2/iw+Vuf6Njw2mRh7R2s9//Um88EDcpp8rTm
ak/HL3Rw2qWiF6mCJuesbuouzJA7efIyciVZUJ+Ps4oNqhSQ6d3Lx9dsT4U+tn4d
UCDJtVR/KuHkNqveKhagWVLZrGACylxDd5nKud72v38+mJ5hGH+b4sJkVrrr3sn7
ve/8ZgyL7z+vK5pWhyOVoUSAh65qmkyO5t6FfBrossusq5uzlueyJGHqZjalQLYY
VM26tAhe9Ajk1XevfQcjGSeNT3dQquCxA5SmZjBu/LgDNuXElqrGcTHck9t9i5hS
x/MsvCbuck5F9UucrQUoMpj48BYv5E+UBP6EVt67Lh5p7tf1BMEKA6qglsbUAFlQ
gsTcf9Iop7d2cMi8ESO7MFugEDlOGRd3ZH6gbR1JnJCDOUuWlZmiYVuI5pJTMXRS
+zFak1yYEXevjfsTI0FY1b48TW6AXlTiGei8HJmddplcwHXPcBY0Vub0i2TxUoKa
W1j1dYZZnRLYRLGKavN9SJmQj6E7DoqmwAdxz6rHbvGe3oUtcXqkHJDMUCc8accs
zPV7vKSECLYaEGZgu2CRxaCS5tP1RWl1XsF1UDI5FSVDGWu+TQ1QmDW1tURzkpGG
AxspbSG0Oyn9FcZXx6TiThoYFAZkRdZGpQxc6NVUMdyz1if9CN/kkrigFX8TGzZg
lj9AY+WcoTtyDmcdsduSIVnd65aaq9zcrbnt7xftqYG7tdwZSvDu71UE1h3+uhdE
W8dqEki+CvyzfBrwmwJotoqvwILGbtpmZ2TIl5n0Rw6gxT9NoD1TMZ1f6u16xQ0E
jnS8M03PnZcJFeQRlJBm4nRQ2Q8pQtKYgaDlXRvz1vJnY1ecDnRhlq0gK5678oGs
VOXsc2LN5MJe6ToQdDbg4oRheAhIs1bHwPVCJrenJU/hVJ1RrkI+USaQ92LxX52e
lN0Fq7/ideqZVTDGbu+R3z58NXejG9vi4WQUpiM0NZLHkkrHXiOq8Ou2TDUbqCTr
l49K2OR8ZlC/jCl1kZ4gcZUGQ/4bBNtqmQYAtdOPLJ5jsoj8DyBn/vzjcpuvaTtt
8UgVaohQbhHHFeQw29OrAmPIfdzdBj/B5EfDHBMFI+RN+dOxlFjibtg2BdH/iFJJ
9E/CRk+QJVaKvta9Tc2ZT6Xdki1fXb+RJGnltUOpER8d9OQYkuJ/ih8Yy0kJ3dO+
jAT9c1Pb7u35Kz0ATuCsv1vqkpiJ3q0wxXv7UUHS4uma8D4jbP+LBRM6ieAcTmPe
GICEdeA10vblhLRty+ukEBh4YVBY3ScDffUF63kyu7y3FhyPhyiFE5ON1wxxKwnV
sxn8jSy+bdpyRalJfGh32xbp2LpfE4QVhSPqZpKd161WO9mtl4eQyH30bgyq4r0d
foF6rYOiXKCQzazoGPnbjwcCDUBPz9gIU0Vqa1io9tbTT8UnNH8ag1L/qSuBD8F0
G5KJkUouA+SmH+moFDnbhuNW2EELPYK6TCDiiPlXo5HCEWK9FJIKKWr1ABZOO1aL
tqro/c2n8xGUcjQse10uPRn6gCrj0HQgF9Mg774QhV/fOcLz9DJpVC7W3r5zXCzW
0vAo5MXBz56GEIDbXftcVuUQBvf+x1peyea9FOD4goML7Wyd8zohEP+PUJwfCaMO
X7A77yr6RjfKHoeNRfPetGSPVqzPjAuNA+wlAxuj8vc4c7H2su6/lpUU+4rzYbHZ
oufpWeVQ2RVGsGBy3CXznJG70u2gnznjeaLGfdczbGG/3XQgNZuDRG7Rxvfh3CeI
RJHSpfw13xDiiKB1zpq1G6KkJWZ3Ejsm3Xi58wd+/mF79SX5DNbMrM7qeT0kLyQV
Cer+2rw3TydiFKqVycb/21HoT3CSGH0mK2zrFnTHp3VDU/3QwNsKbVihVzsBtGFi
cceLeVtyDA0seuthfpI9uYTC5J2B5J3nYKLB0dOt02LcNy9SmIMtpWnVyC2ooCgY
9mHBWIlVNZrG6XAWueof8T51zwF7k3Q6Oik/3IpaLuC7VLQb17v2NyAgrraxLpy0
wgYCRaHNClfbBj6zVIamONOl0aR1l7z9W8V2Hjpc+xhBEdK12f4gAgJ9VSAPzOI8
8dhKk6kln/eVqonwIBv7rqw3WOH3zntMUXlISzAzD1T9j1E5M78DJw33cUjFO2OI
WfGQzvj1nnB7zYz5BmAwM1m4juVVFBogomNjDlV5kljwanLQRFKyl76N2JcgqC1v
js28xW0PGtKgP64Q1rEVLA4sZQVqNaCTf6UgW2rss4H0MyJK6VVjXfA61yaalqXu
LOj+nVIm1GSU/aa9wVVdf3W189Udc3Vlx0eu8MJKHK6OvbiNvZ8n3XLdUvW8ebDu
QmcRXIhURE0iNzzpkyUbmQZU1nW00QkAr3GdByxh8ZfgvJaN29G0CcOpGO0/7vQE
dC+sDOWQ086GQfexBQibz5xFpJiQcdPNsq9yGTnhJTsidBeApJkSgRL7qEewfHw0
iNdPmXIK2IbypsTbg1M8RrCkTMvglzRo1kx6iTpuN1IULY78pvXlJjeV6sb2hdQa
wIflzybChufEpILm7WWTH5ND8sSB95hhVarlUDmT90/Tv1ETKQx+mqcjR3TV+4rX
l5BJjpG6+cBGf0BeIYTmxv18rpeohIlCU5vcgTMODI0PLEBBsNLZUn4aXGbrrQdj
j+kwnjFo0vSaTBkg+Jdw8Jw4QAM0asqAjsoSf9h7b3x3FbZxI0wLiTpqtzAXisCt
g+aIk0ZSedPApNiSeAUcrlWIsJ0uPmX+qTweYPG82mKEUgSIgCy8j6VUC7ncLZmZ
gp834eXdixIiNVvUI8zcEppOEcFBQP4S+bSlNP7RYezaQBVV+L1L8fu15eCT8sHP
SujCSZbUPPyIXInXstM3FRjTNdajNkqDLBi76xuInzIt7jD/PrYD3B73SpLW0qFy
bFoklZ2TJnxrnkEeAxK9IObRkMzxuvedvwTHrR8HSIpIi6PK8qYrI9HFGfaFw4aM
DCiHN92yJYznKO94CXUHDC1CvHHbQIML6fU5sO+835yiSyT5Zeuzsstb8pjNJj/G
7nujvhsT+ZjBGw+GIdLUOKVgK8lzfJeRKGdKpxt03V6SJOccTu+1YGy5PZuDwquo
1HeRmJzL7lSISdp7WE0tKDXFzcddmHh2cAmeQvEAyhTvkBlptu5XUNLstEqsqyhw
fGaF2uIbl4ukCoF/YIOUzNnbnv+Tb7RGIogTQWx2aarjKkBe/GN9kH466Va8gtpD
XznOHDSZ2LahWQbpN2u2taYXfYb0qRcIpTWzKVB0BGIpP4w8KbHXSusJikPz2stk
Egp5+xhTVXOohh/oGsfVGW/xfPwfaFNsVztSEJRWIHA9/8OEowo6bQBKNAURMEvB
+Gl2xx9864GlvvBkeK1g5SjJLFWVYlsMH5H6q8ctTHC1mJZkes5FapM7GAmEzgau
EMUALEw1pPGKeVm1NFsABuMs7aYjWSE3JdjAuz1hivk2uPsGs76cVbIDOW4zwtEd
ceEUvaQz/KQKoUHT4diyOE4AGkuQUP511Pfc4WYraTPB4GNDfNX/VYIBvvwMACSo
WhMkvOzorcX7hDSJBvB42Acq5E+OzypzynEzUw3UHJmXX3QSCBVFcT+29J3I5/oz
zn/DKDa4mq5RSkxZ8A8Qmg4w14UvJ7Xlnyitln9j/ef/AAz5nD151ETZ0TGrvCuf
FMHOPARcQbAHHjK4FWOYZtqQxYTrgEnics/ZsQh5cEeVUeoWcyXa60jfn7GVC28J
ijBKltk7anmUlgOMEHa79pvU0oq+DVu4ORi/gPd9Fti2O51s9ogsshOl0t2YEZ/a
f35AY77S7OBS8GobVS3J4M5HbaRk0hV7cZfGXI/dn7GJg6ykv9fe0pmQkFuEWi8z
zatkhyQlxQdGAXkT5dsmJbnO0iib27EAuRON0eNUckPpQCAcEZcCtkmhROqp5lGb
1xzsG++Cga0dh7WgKkMv0UhF3rVkgMzFg9iSVLjqpzrDwT0u3yqqfLq9suzCoY17
DcXH6Kii2U16ynYZkaF+aCQrwZcSsIy4NyevAGIQpcFW7i9QB6zbsNu9VTY6BVE/
fINni8gHau9YMx2qx23tr9CPSSS3CxlY/HxoKRmSGW3oQgapeTW2J7yMqI6OGQLj
CQLTRPrbEegOc1y5C/kdPfxkJj/hAcwSUa1lJYc/FTyR2oAoSkti/xKcdZVktCV9
U4n3JPhSGnNszbgGuMAVjtYpY2N0kF2WLN9UvNo2YZCPcjKTPmOoh6QihkWja9uk
RFZwHAbFA+L6k16mVJsFKLavHMlzq4Ry619rTUggXcsEbQsQyyc7TUtfcU3+hjNr
Bwck8YNNc8tG8mLabh5ozORNI3wt5nKBzgqvgIZMGrQ5NaLrHxFJl4ASQAuLlDrQ
gVPgz8QO/zulRAc2ACDNeGdjxhwvQMqEfSQmeZfe9byu0MfCiclouWtVuK6YLUzW
h4sMeNNJEGUj0wm0OYOfMhnrHTn/TYWPZyT/9rosVHg1Xot3jON+Mf8wGfTDG0OC
PCyCDckHOhs8f0CZC3ojUBziLgXe3qzdIwfHVuOKecM5Mg20RV3H0bJxh4s3HuEH
WnLYjPoVEsXTJXxOwNrOLun2Zhe32pP1jUZpH3XJ2jU+csoawGqkGJ8NCPKWdR1I
lIPDOpINLISu2qxAtsUOT437CABdMaVUizJo6yUBrpsIGL5A3bsCtKuPzSAenJTq
gu0t6LiujwgmNkC71TMwoMt8vxZQqhyEgMRExEWnPGvF3yyhgebLG1RDKgurHToK
Rzf5CbQg1//KcR31icRjXnOb4skbmx/iQhrfHXQto4cYUn447AIIqIA7262GP7ae
wOI3d38gpzaU7TsfCQHPLY7xiNPsDgGuZZV8jQrVyVPJEKKhEHhu5EqG8AMRCR6b
bpLNsQ6FSn8Z0imvTLl0f44vEF0m1Ug8kvPp/WF2aAQTTOYAH5HjZbuf5cUze5yI
bViT+qp14JyBDfe1+DA+v5slh0PQMy7amKoP2KfgpXOimwj0DWd01AmX74woMP63
9MnXqQ0twL1TkLvw3px0vIaTGJ0ST0Ay6oa6X5PZmr3slxH0gAvDOYnq6N6nzwhg
yso4xFHDVlJBPfmPgewosJx/BAhNNJLSqZ0L0K5taLAdvjnRKYctUSbdE0sS5myo
s0zD2p91oxm094fww3h8RkHAi8mDnc7euz+wFKKd1jIUyqxBxbZ5jo6uQ8QncKYu
M5i1NAA3pFt72rxNk0HzJUrlBVhrwtj9fRlVYrnLdBIony3z9wM6WSBaGATPrfUH
r3wv73A0dDt+ey0GU7EeJ+0cQbMzzuWINLiqEWG6pJ1nVuDBJNyvH6mKOGejPAg/
QZlWLrrSdbV7jS/IG/Ka4Ngyqqbj4jsiqLBjtYbTYrMTK6CX4KuIB8+BYHURfjCS
4tmp+aadE56hGEs8P2i0zPXDwecNUEuQLgWltfdTWFxpiLXtpmg3K9ahxclQuoew
QmTfvOWFju4eHJf2t4dSDkJXp8mleb3o3vu5hbUfLxaGFsMIPMxZag/TzzyR68+z
Z2VzdwdhoNaNN4TvDG+CeGWQaVCdknojm48k0oNeRgs46AP3SSHe4RF4pnulBUdX
BLuiqZcYYHJMgaG8DjgG9wj3abkB7/+Mptq+w6nfB8lwvSZXuSFtQqZNIDB2krCe
gN3OsXAtjbeWTw18mVsBEEiUEgoVkG5WrKP2exBUes6ww/RHMW8pbu1dXIkkHrE6
JK7Hc/5ZHwgPlUiNXH0N10V4wD5GH20McaYH/e3n+s7Ua7SQ8BMhNHgaSkhsocKO
/zSep5BWta0mo9mhIMcqYEoCfSOJ77vku8WYwH01GZ/Ua+5ZxvcmHb9Fk+C9fwLP
wkCSp6oqCfudIdAWRobCEPOr1Y3OyEfugnAqeohTmMlKlZFRvkLt2bivJG0S7Ee9
HMcny1xRwGpeloOunwrDRzJv8WzQR1l0Rq53JKCZXZWvxjLeIzKBFDWT96Bl332P
Pd2i6qSAIDnDDxx5SdPnV6Ae1z9DpH1gCQXG7WIHIdJq30k7P+MXQglgpjEse+n7
K1xTMq7bVhZXOVIeaq1Jv71cp2BCPVePwEh6YR6ZgsgWTXTMnSqLyD5hKvjALNQ+
viVz7Tu3gbKBduq0dbb7fIjmkXGC3qj0McTBHhXTKGCzOfqjCuJWYgMkv7rP0A+V
AXMUBrsplpzVQI4rQMYtclqmShrJnXodF87z3VV42dc2Zs9XrmbikDp+RDBlbD34
93E0W54DdXTQpjzu6is9yQ+JKNDWLEH3Ys0yYElf1UCH9X2MJjdTwp3J5s8drsxu
Yom+Gqq4W1mMSa8TMClrC29KE0u5ttz4GBZeZNerOd8cVKPbmwJdT9+s8lDA+X0D
V1KrOkuCJI9H3zGA8GUzi6fzfg7BGfWtiD+tAiqpVtnvFPjAMqPPSkcUWEfuJ4Qt
Tj8B4+XOoj0S+8qRPZBJk/NRFO+6O18orGJrRbhFTEl6+JNyGeqSAAoga4u8v8JE
sjUfcgVaiK/EUpdTvT2bmQYwm7gwrAXdp6fZBhA6IabVJYGLkX5MFn92wDARWA80
K9cqazYU0iDHIhyHvVVQ+I1le4M+2kQT6UveBwlZWu/oQwowHHEpqShsc9mOTnB/
Gw8ff63btUUUNqw2y1fInH/hrIq5PW1nUH0ba3SlkCZ+V7U7ZTLIyVoZWE8QnBZL
2ehxGxTExnnKXaALAmwVONVB52zieDOPt9jmr2c04RgSU+LuIR4JWfdkYxvRkU2H
JH0seMDdhmc96mrYrWH0ws3SE5TAb2Cu16q3YinK61pbFHpzqqsEezsQTD72MzHj
YdAHpWXzFJ6PdvnpXxtqUi2fGRDidzMaUSSv+c2fdvMyDvqefULieIvwoYTU2mOH
z/cQ1E7NjZy3rHnnNMPzZpVxaGmc7HSoBxj/5FW2//2tvDTHX3h9/yJjY5S01Hab
t4Kpqp95x+NmS56p2xF688f5JRHBx2opyviKuN2+xAlIx+ZBya8MzFQ7i91vHy3K
KS3eD/sVXkGb8Jcr36272Mnp7dblieAm+lQuKCQLBaSnRmiLOiX1QKujmKbE9luh
yN++HphsP0SG405oSpq6eUrMN3jQ7ma/yZK7AhE8zX7Ik1zEKXFaeh900EDOzUv3
1ZayQEHJ/nuJ4Mh2an1tO0OQYmbgCvvjkGhHRACDNrZRLnn6DvpENkcxBkRK13Lj
FRlOL82rhIH/Xhw1ATU0kyr4ukhKDoRCfebd2eIADtKRy6OBzxwbyaZmXaHuIwVv
YCuHXMVZ/76kh2P651DPOJAkEcSGPVuSChCHZJq1sQeFJx7XzxI/c79bLkNtBJEt
xPRJnuWE6yKunSXTKJuUmtXn8Zsbh4Cw90oSLd7kqwOEgTqSsSPsUKnLJt1iG1Mk
H2lNP6FaZu3bZF7ESl6W9WDNXbw8dh0WN/gxCaHPgEhaHiLXcpBOeVYE/PcL6MvP
TGGHEP1NcO9PC4SMYCl8h4+lm7roMj3Am2SsjFuYZyG0r8Y2ofPYUlgyjwRkF5fq
SX/lN610aVeDl5X9zjH8gAYyKnOP5cZ4FJ9ixy+e2Eb0nSxNHJA2SFSBccanGUpr
sxJu1yZELQV1zwCIrmJtrZJiDyh/jL89o5p3BLrCO7xoAza/yJ8+VGF5w1ZlsCvm
4kF5X6paKnkbGyqjMMozn0UtwYUPoMelTg+uViGuCfgaUaMk0T0V11zVHgBpt/4+
HLqzirwfythP7YqhA0n6Ihl6/J0VfKc27lQxKcXT9Ggl1T7cUIc0DDlgJzJgJwto
2AL8qn9D4p7kDGEUIktQfdSMRw2Nsk+CdgCJBvp01tacTMFBVW3TNsLjRoxmN275
RM3smb+01gJk6pvdl09MMPliW8dTZz7Vrvp29ycq8YBztcORFPkzlAbb24TyFdLg
FJU3zOBUToPG8rvqUCyzz21nFRi69XHNYVcMKpfHdGUxx0GLxi9ASNjpkkxJs4jr
rWIwCbbH6DZKV8hZE0jk3ngGnrqHzlYXnk9+pLLH2O4uUteADDqXN8AmJdCvdBV0
q6QsmtOiVw7oDIGEQx6xe5VhXddmyV+j3q2zrGBhvGqsTExQX/iUBLHgWR5/eUzT
o0pcH6tZjTDZnRYwYVUP9YoePWLaR4ZmYPJ2PQdy0tEYsdHYLlSmmTlnXfU/FUrX
yfslTDfdssW9Gt7Dgm6/BtMN1PKveUAUm6Fl3VINePpzwIqP6EC6T2QrUROdlh32
TAkxDBYYstZeYft7e2zoHjOyff27hjycIHg4KafO62glJVghfqHdW7p0mu/TJoYB
OSpR9xwGTw87kjFyTRo5ptRqtOX/pXeQ6kbXfl3Ex8bpvaFFHIbpgZfj8vijutHa
T8wW9//1Us9G6QOc2S3/Kcr4nlh1SmOHozcXJHL8XM/ErE7ehs25xxOHPAgudC4M
uXzayntYpvVoQDosgWEN4B3OsYKaUSz7LYtiLoEagzkn7pRLeLnJeifqE3IOf6lI
O4aBfz07pG8WeUlmhvHWawZLgzKGrZeUHiFvyz66/8ZRRz+lfWhuj/YUFQk1Ntr7
M3lTOOs+JXK4gdSj3B36F0I0VSZiQ0lSWWE6QEvmCtELekPm5mCuhj2R9JmeK2+e
jKTgeWcC9TbAycP7mmd+/ptdkk+UbK8zsU5P05sB/SDq1jD9QJRVOFh8whVhB2/t
J5+cF9iqnVJ0HypwbqJogO/Esy93YFLIv+5m0OZbfV7/LtYJK/5SFUja2tF1QJ4K
Ksq7uBG2oSJQmdG8q4NFiwy2AYNiQEsMzrwNPz/9O4oTbf/VaHRrC7Kl6CBj/fnn
SBhjPtkiDMdfbiAxOAx3nnlQ5/IDrYUqQTARqcLp0pbMtvj/Xw6hXDQPbcfB6Fwf
XqXq60NTuRBLEl70YOQSJLy+u5/bQZw7nvw6WvgO6sHFHTrxuBnyBREOh3b5QepL
CdDo6+rE/kpkZQJWyLnc10k8haw2PjVg+EFELyLjDFXeG3THPVvfOxxBfHEwzOn4
GvP/nH8DQTppqTpxzg7+W+XESmp4lmxZIsFrZ+F0jwS99l1rEyynvFD4j2SM1WSn
6gsYF4ZZ/HmLRf9Kktj6LvsJxMaqE18XBBwin53rnYQCXS+3i4tTnlCp7827u2Bk
JogVoOVU7Vv/UquK9fjvEJKlostkzSNdLlSibYwZreaWrjskCuod4hQf54P5Zv6o
UJjf1VH0nv7Ib0Pu19PnxRortOq618iIrevbf13Q+D+TRKl7M/u1jlMisXcyzLQ5
k1R3kbKqj96nkSAuAtb7JXiLMQ0nW3vFcRDm4F8jKPotqR3t1jTUcfLBTV60ZbZI
7QUMegog9z2R63AQT863t8nDkIDd/aFzPyAnEOCnbgmw+n1BkjNwFkCooyPE8AjI
ba2Er1hKsrSkcntZEOuTz/Lf95DlaoeMc3iMEIH8BsfABDsL3ZK1hyYIrSO9iwlx
gN8nVsHfyGB93Ek+skeV6hUUpK1A4nMhcgtr7zYbjvSntkg55VPEv3b+cAVy40YR
IUz/8z3tiVSzaJYggoibi3FDT/38w+SrLpjeru9RpSKWU1YooRqvwfrQAWZ3gQqj
9/bebK20/8TnCMTTFfjYajtiRDxXAxOWS4RH63xfRUPVjBhLfRlEMWdKjsm/aR5J
nkUNvsWtopBe5ABz1kAOmQQ4DS0MVR0JxU7zx9h9ksiMyrQQbeUqfUAGcqvCp6o5
WCZwlHdJ+ZG0Ez+ylebLtC5Z6tDqR2BFDWAnzzxWvPnNovWzXyU1DG/ktPjVTABW
lan4wMV6TuipYS1nBIMe0C1L1KfEmVRL84wOkTglw3G+9GvldhRRnAwxojXnBJ03
Clorx74TXZi6g1xkIP5/sCFx0D+ZpmY0GM+tF7fbtRbCwAykMaXQubgEFKcaktkX
j14fXem1Q2QHacPXQHDGho8EpEQaNuFv4phWoHZhiLNQZsx302hLMRutWq6ehZgl
4/rsAFBtdexIbkuQOa1XzzW37uEqJJLmhHUo9XP0pSkt8ReNvvgLTIxEqx16i4i5
PBsR2I/rabLOTVaoFCOEvmPlw3D2KPZ82wSucuNWj7gRui2KyJZvLRn6D82EuxWo
hoSKvdvll0bieKzjdWX89oXluIEjjsEGGDjT5Pd40JM1yPP4aRGg+fOMUjxhi7UL
EEYCzhk2K3rf5qDyYE+yX4gF7wRmA+eXgarshXRr+hMc/8RqyWlZKlsPeMstF0rC
ftjk7b4NLunwGCoCY0JpwtB0RZ7g9yupiUFqNgp3r7hWQhpQb5Wl5gBEqqEevhxJ
9AlgV0IASFuyzPmfSYE/+yuem35+OLpp8RxTj+3PWgpGZFasg9nShM9zmlXJWru/
ah4Lrliu22RiGGHlgHL+c0CSGyjiY2Qx9JgGmWIWnBW563AvxOH7NfHVc+r3Uw/g
FVqtUKvbaPirx9oFG1w5qnrmmfBH8W5/oVbcsrJZZCVFc9A2GyfEdLIDxBPtblL3
bcxie+9bpSxReJNwLlQ/Oo+Zxhzn1f2FXr34Fn0R1M58/12+GBdX6H3PLJX01J9g
38s5VCoziPNILDJiQdEF/NVkZkySGSyOo57D9Skf+cZox8j3tpJspsXLy83C8zCU
0/wYtoxIQOTWhrP2xQzSKhG2XWptJ6IxLUhd0CqYpn35hAbld1Ejz4pJz8kqE0GO
Iq8Ir7ZVQUnj/1nraR9IQme4appDUgraMZZ348O6fGcczU/Q5DmdunJUQEAJJL17
vYZ8bOSBntBeF7fm4Z1TYzdrI8jAWaA9Z7hmfo1zIuM4um72juUJ+/RAAu0SguZz
2L+XRfUN4gE4wqJTBWpN6wFbjU1KlTZHgCsYOINhmnfNiSAcbOAOKrAtBxkbwURn
Yoqb8IJgTA6hV4QSQdh16FyN9nJVDtLsoQa8pIQ+WfaLEhhDjDnn9qpmn3WBCuhw
x61JUALApZYkbe3yVbztaeD3nqLqFqtWiwWOFbnDu/nE6yTC8lkuG2K5Pc6GPVDm
R6vbGX4MU+PflzE09TlwWsGDU/wxTE7SduCL4CzzB4uELSMSv3PA/VUip58aHzNC
rfHux67X62gazqPOmag2Y+ieambXbirCWGfFYjb/9ok4bGaXtfY9NpQrC7k9HcWa
YK8UxVlVqdDiZkJsK3kvqY0UoId8aymBYM00+hEZE9A5KJdYsMJUSs3Kff4wnNW8
ouNoQ2XgIHRWh2Kh5LtIkoL7tyLsQWpx23K1DR8ymJuOzclclAOkhlxZzNCWfDl8
ML/apyms1L+Bo/x9d7pongjdSB0kZwFUFRmb2HfKYFA6YLgq/Y4DocSiXCOqFs/F
x2qC9FB/1t8xR6Cxn18iG54bWAMa0/niieVAhtAEVBtRviN/rqjeaDXfWjZuSb7C
JQvHdN6GmRfsFjY16tmJb8QrpJEtCuBBFLUmXiFXiUrM062b1PtXNxP0RVXWDfC3
OxCkpd/EMCmljHHPgudRZ+Cnq9U1FlLOCY8U7RqgfvwIWcBkIKi4byNfm2qeATVt
/zP2Ia+5rEDCuRWNUSuKZb649AFXVMsDmGD3UpQxfDhaX48qmNWRTiUjZlw+gfjZ
3oKRd00f7oTKnp/9a+TS8Iv5GW3lfEo7u9D26D5KwLOtQ/y7+S9if5LYGxudF2j3
PPWiB3HoLP3EOAlPm7qzUFrsCuNeT3eIIbCMrvTxbu2zvgqcJubR27+HgUGR0in0
IndgsvWlnYuEXtLJlUTFI6ACtxB1x+P5Ffch1Ksg8ysufJAd/uZI3CgD3hPlr26g
yuiq3YrLljjYPnmE/jXEnxh+msSe6CMhSUfkPSl4Hpg1EzTHOK5Zplen33qRb410
ICl5M8dNKU+ryMS0UDEWdSwdSLv7ju3rEjzJ7ba0vLGcIg9ooGcoxUyDihsg8jgo
2u0ldNlEd9EFMdv+uqdl6jUYd7HkAXxCB3yb10H6LQmzZxZ+TXtncg2/M9u534H/
eRPaUSFqpOC8FTjggu32tOjfc03ENNkXuD4L9tE5iBA6VQR/Fty6a79b8QG9ZYqg
IK6lvvTbJXqV9NZDA1Gqus5D4SQ5wZj0CPnkRNhbTbjr2HPCQodlu8n8PxLIslCW
1azEll/zKitNPFTZXDVehXsuiGl+OfJzH40h3G16fFt1BQ5pP/gde0UcdJ8E9QRG
jlEsHA2CHwim+5vlGHYfjwGvixRtLWOy2MfbFhErTx8dUZPp72VQd6YXRHVkOrtz
+/2YqZh18YD1J8KSAV1gaOQVf8Ddx9Xfe2B6yRFIJOw05DJ/jUZyDOaxyG4ccafb
r6yyuAWCvv6iAcGXFxOX6WY7s8OSwA6YuwGONCD2V3ZhE7ZPlQDla3D5+woKOcXa
9dnOKBu8orb3uwT1LZM3nFqbpATOYL0tTKyDGE0fbBKTAvyG7Dhr+6FxS9Ha8LZq
muJ9ptjMZZNCWdRS1oKOHUD3n+pZfnXXwm+CN0ZXF+PrMYF18dtjOsyyoAGZ+REg
6ecFr9pjY+drmDyK3DhYeUcBFWJvosl0tUzN+KWGlnr71vr21mIw//TDCSrrV7od
Oo0Y0qCaxxbL1u7S4K+8Tfvp4PEgJTfVgg9qWT8p2ZivzndJ37c3PUqwtvHdzf4t
6ExroS/+8P3k92bM2L6rEAUcSUGQej2XpvedCXuhtUFVnVMBEMblV/MQ+RhFtZCG
yegUcRFkSatp/WRU7cMLYlmhGkFmaicazFiZi9KRnTveitbkyPlLQ371pPvJduzt
N0CDTj48UTZBRPvreuYZQW6kNxoplVYGr6BsFLg0f6Xq/9JHwNPQddSgVrWgp5LE
hh52MzHMHcthGN0d278eYSNj6ZYxuGUusLy5izrnHVNUz2sgfFIIdrpYCxzVoZ8v
eTg8z2GdQ2P5wqd1TRBLlW6FZBB+p1Maubox2Cjy4+bMFoMTsf25Y2BCv6N4EAtK
Gi3PU0KprdTMY3/VJ46aYfGlpIy3GDBJlr8KsfXI4MIdTyM5XyDdjj8N4d6jCyhK
q0NN/r+XPDnenSiEqVyV7srgQE0qsWTssAiXV60IvGby1Z4Wl/+VA574nOuSvGuh
rnRwUNUHSsjBoLyCanKOkR8kzUFRStxuKMu0n1vSmhH2BribAGZex4r/zS958Sm6
VTbMpJX2laGjn+n54r8O+34MJcJMsf9SWfPXTKDHeCnDJSuF4EGHwBLgc3+CKaul
PalGvhXOKwZJNkj36KwH4TD+gz/3GGrT+6B0DQcoudS38NYgB0Uj1WXmcd7WHpMi
eZLJo5sAjU7cjEUnhkoHVBYSYyYxYbCMjpXcDJ7nD9j4WmA45zIfBz7rAXFEefTW
l3zTjIYyO/vpcrjBWNKHoyhgRUTAbXC+PuLZMmeB59M=
`protect END_PROTECTED
