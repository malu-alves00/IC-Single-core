`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ee0/5I6aoP/UeFUpcavxDZLXI5kgxLfQMjPRl9HxRaxKF0yq7WOhUxp8xs25by0p
kCsGYCVEBjcseDkkjEI/d9naZ2Yb70wXonUXXlx5dYJZLbqMjTrWpFstDBiqkFr0
6AgNVZDI9LlfUnqVUQj6xd0eqSNZ8vDPP8+r8yrQ2u/2PeF9xeKTjPXSJkCksd2R
F9zppCg47O6Zpvr+SKFceKt+uhej5HL3TlT4B5t0/0cGubT8JhP6jsneVNdElRpV
ZvipsykEaycC6GE+XUSLK4qx5NDq9rnCmcj9IQfWLnISWGJIq4HURF6dRsZQvwbg
fgD0pIJoC+ARbTtl6gHu/rQVKBAwWyCPoBzNwk5D2sJ9tEVLd7y6hGYfwWbeJ5Hz
UcbfesIwFxYad2mPy3DJrpHokmjQAoRmd+04oeBh7cRb4+XsIeXPMSv65IRpVit4
GOyP9lvbtHErHhUTE/+MO2dKNy3VpDTuUIhogGyXB1gF9rnxYYqWOIgkDy/70AMx
bjsOAUmW085AisIXkIQpGyHoJoLLO/sIh2jN4QF7boqyZNBjiOyqg3G1xyO6fqz6
O+we4kG02uI6AKXl29w2HiWVcFMPEPBmHBQ5D5JI2yelNQXjLDlN069W+4if+tby
KbYYWKYuFZSC9X/hlooIeJDrOjtlb5cYxsadA+r5vMO5boUEWDv/+NYjbiG0LJrY
pxf9YD37esDY/FEhgnyBF1LL0jIIxULWIlaYnWQxTOTZxeShSRtbNPGbOD/ia7BC
wfsuMY83xxpd2j55vr+2CFxu9PQKgjsfgErKrqALILvmOOeMfO2Ah99Z0jFSY+Kk
`protect END_PROTECTED
