`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XEw/W6hUgWzyFUca+xQ0m3k0rN2Q7sT9Oehmjcp65CPZFqCTMnjaHg1QYOfHqHQG
djc7eLlRlD2heQEJe5NVJpA7nve99ZZrxFBgFbNenwunXEN+zfHIpots8mKHc9DZ
ewvv7sT8gQkg2m9ZIMT0fMw0CYh8CcMKR8U4Q2tvGDnnzW55R2jc3M5+PLKsCVsY
wyvizqh363uoCp7EZBmT7u4WKYOyudoZ4RRgid8qhs04KSZjuuaFutaViu4nNJcT
ytKL4TeqhvQEQnbnNFVhb1WK5fcUCXeNDGncjCLcgMPGZXaWJ7Rh5ScaZy4/ktG2
dwJD0v0Wq/3yC2srRj7hk88D4dn81AA1Rm3Jo24FXnl6KgLv5BTwkdDzpS8jDbCH
a1HaMrMhsupWhxB3T47uzKal1cJ3tHmd4+wSAd/dd2iCxuZRtfuFiKmeQEHFbaMT
yewJsk6kvbT5lWkGq1k3tDN/kzuAQTVIFcSBM9r4pGxAbAzT0avj+aqvVURVW+Q2
jo+4sao2JRKlZnbjOF0bbwNMf7/LwJM3S/BUbpFsG/+KSGPrDNzc2MFb9NzDHgRU
TZTTtX4J4ObNtZGf8K1Xf51cAQSDptmsFXJBXUX1d31NDS/c/RYD1jCLwy33FZf5
3tyWOYyhk5MTpoReIzU8XGLJa5ynNkwF6DgPlQzhXKa+5stzF66d52Z8U15umItA
WqveDeGQy1ItUWtPdt7zfN2nNe5X7h8He632PRdiA+0QkNBTpoNs55JYGenc4b1y
2T1UU4wQCUxr6KWIUYzL/HdKzgmmbtDBHmXsCNPrpee5FWhhwory64J4yfAb2vvX
gVUWNcNWpXU/2fQGQC1TdyR6BvvG6+vo6Sg8ImBVZG/56K2ZTErMmAaH6jxS2Htd
UIAdDIPFvb66F9VPbpqgsqD1SCso6AGemVZ1rIUpPc9rrFYIG7krXEa4FF08l72+
K+F0dUGYn6s1tnZGaxiPSX91cl9s1i1PNTHUmQqaFsNeVS/dRvUrenp3fqnfDxdt
gNs17Tlxh8t1QQHXRPoYgWYM1vq54xprrYQ+XAA8hzQzRo2y9xmid4PYhPb1QvHr
sxE8e59447h3Rpaf6BRSjkevmJxBU2BdpGDu3JC2QUdElpNASt3Mf2ZOvWFrHAH0
cMSlGT4V+jI051TUxukXWCM6Q8A8MbXbTwFfAXR2dAIoNSHIUhqu5TMfR2SDoNMW
/ZDfHdGY1Y7F6J9UDiAHt7bJVH55aRXrwMlTwvWTe86i5C6Ds8K0MKBMn+P+4ywE
SND9L2vHUlY3rGJ2YiSkIktopDo/n99dN1vTo87bItP7gx5oBzymJG3fjzDy/CKH
+eBI0NvcdgJtpyO8YVF/dxdQH+U11+V5GO/65DhvsV8udZTarL6hgyZfR+lwZx1Q
Ir/ngNDvvTRQ8OBjjfKCfrkY850vZra7bryFM95INX2hsZ2jkAJwGV0OkWHsFY5S
zsvVzNZyaApN22DsMag75C/HVA4h7UKS0bCSeXcS9Rg=
`protect END_PROTECTED
