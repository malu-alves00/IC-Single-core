`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FpqMj3mqNjgIeQ82yAUAwIgehBpZz+uYLMJPkB8R0aiDjrFCJMcxIl8+27VNg+xb
7bbvoRX6bJj+XpQy6EzrWy062KMnT854Bp7CokKp9Rf3HWTMwKGzW/Mna6sjr6DO
4NoLZ0cexFe6v6O1ZRoadqNn0c1IO/WsRcWKDoiOLMnHmWV+dbSxeluZqSP2x2xM
UgBqeRo0yz03NO/tsVESGAR8aIu6T0l9sZRraIMCQ1CFnjoU0mVfblM+mGNtz9es
RfotD4SfucaLRnToXCKjl4z4ULBpPu3guT+LFRo90DBx8oGGMrBtsNDBuoZOciqm
Ly77SrADgtlK7xuENIKMriYK1WivJZwZ8V6FzQ4hEYNEgEB8g1w3eTEI0/JQpviY
O3tBpsIw3aisZp0iwZo8LQhKB54Ju5RXO6ah5Mnkx7VAT++dvWqFIZa8hYTFMOV4
Yl6hb2EOtnl6o8UkySUdNyGveimk3ScsOH9NYVMLS7L9XW6uKqHFley98sDR+ba9
tRS2IpqcNAAl7Ws7WTMVqNPOeXPRbNeCgEs/OotbaxCzBgrosWw8k5Dvfti0jxRI
BWTL8D83YqG3Cfx7iz5DCvHMf3YZOLxM7INmafQrEFZ3TTQSzaxfZ5olcoSMNuy2
pmqffN315damQjivSMCQZSAllCb06oQYtahwSA2wZHO236LGsRDSKtNuedicotPl
9mAb0L4H5TvyvAe/k9EfV3W+kW1poci5jNIxPxDtIDIWcYdzyx37EwhOthsGuns9
olF4XWWU0zWW7mud7HgsRqthHChvYSTIeoNCjfC6IFPplfDOZnthFpbsXf6zXtbq
9VGyqeGG18vk5zwkUv1MUs8hTN0R8ojitC+OB6nTWah+FAfdG216bv9AoDg8xoJm
jb6XHDxAD6uZvLHAPJhw7knul8SL8tHDPwnRKD4Ma1XL2Pj+iWC48YHGERGZx1b9
aNnDD7vlb+GZcjos4nJDnuIESxfjZsdFbY0jC6XKWvaRtxHl04PSOqY+P2vwnw8W
iFY598Qich47qDeEULkmuHgDcIDz66k8+mmdY2riiIZ/zDdccFxNYobEkg1r3KGZ
oU6r1dYJTlkPhRBk1k4yb0hH7vRgfOiQVk4+ElR9SnNNcUH1vZ92rlT1tYyh3qF5
nGLl6GFOIBBnIqZRA3jZ9gJBU94e/1PybS7ASS7S4n5r7PBxML392kUiifOBhD1L
DOJ6uMnUy6xvUG1rMiTeggsUxRI47uCWiCqi7HwVGKwxSvBPcAkhzL8WoPjNj1Yf
oyx+skicPaP8bQPwRji47XP3WrhgUmXnWk+Qn7PeTpPItYXFWOHZ4DpLUv7DwFY1
DA80D2VXJ/RpjM4LVkY4xkUoLCPS7DziU4gmvnqr3or1OeT7iWndKeTVaq6AJtRZ
n1jRItIuSJcTZocZvAqYvATo2SABE8d2eZyxs4dNban9odDjbuiCgAvEInzQyTi1
Xp9TX0sjompKCbfrJjCKxQ0tqmlu8wsaYel0BFwhryk9RB64dMhRAP66pdPbPvfR
ZglzKcSrmfvDmojaNbjF/lPFLSbtu+n7QA8w45xQ7JfKIromRkqW8C2ayt+ZVpUd
9aHq4M+yUy7+EsczrmxvcsbO4i2jWleL4PEqrEHzBnyYdLZRUclj1TZ/kjXqTvDp
GFCHusKDY+N27FLeZIoFJa1lzf8Dau4e/Spm2n82jNB3igtSVq3PcbgifB5iN9ij
VpZdz/QEBTbf+D2Kxx95H/enf7ZGiz1upaMInsxgPvHrtG5dXBdntzcGiOzC1tPy
E1nt4bqpmCF9Bsx3UybNDcaRKyvc7pKkAzuvcUUSRIaX0dr1rquwrdxkV41e3rVK
n4GqO/5Yv9zuO1Jl8IYevwRTbQBfRN586+YTbWRD9X2NsysSYNy+8C8FKPBipod2
NkwGp+3TyfoNk/wMkxB+7Q4hnTIFVxV3OTw62BdjP6np8Dauf+gaFeAfvy6utlme
sgSamb3LUri9erwubz2qE4oYjdT8FVe/9zWtlq3Du5QIBsnLB2P8pTppZ/9IAWE6
NtraZJncefEQsixJNwbMbPB5NaRlaOn2LU6fByNnwyRoUq4N2jODad0Z6+XcaVo0
InuTnm+SZ2X6ZHY5Pdw8cuQ8jXJEQo0EUbW6f/V2C/tyoJIwAI6/YIvGCgPqGdZu
w2RQqL6vPyTZ3Xge/97XKUXzfk0DYRnQlKYWUsPyvgTObYnob48clPt6odWZtswN
5UuUYAmzK6M2gi+mmmRKwPxa/mjW9rs3FFP8YsasLp4mM/y5ASCe68JGGNXINuoe
33uus8BOpm2lQgmnSWa1ActnbPFo5b+sKYfnbahKGrb+4wAgwyN8CIPR+2fkCbut
Dwn/FwSjRckqBCafplNGAd/nq8YiHzvMOe6rreZ7v2oMuOXqKDlvxfkuYIc2wpVH
Y0b9CpFeudMmkP1GXVaITrDhlEDKtUqeATvtnhi8RWLoJ4p0fsyQlheIdv9ei49n
C6ItNKGETqrBGGq/xFRkAt7Y4XnNZ8tw0OPBtE+h2pBb7yBzH2QonSO1yVi1pMmF
yyiDDehT+mGbGIFEuQ55mZrBk+FYZWRAUsAmKoiPQck6Aklpdk7lmqy6rDpUxhyF
UPbWo+NVOq0qoUZaD6k9i0zYIFuw+EbcRbdJfl9f9kfImGFSUfSC2cgSn2XymoSu
78BL2AEX/XX9aTUz+S2AG7AHZQitHMGG/stg9yppw5hFNKmwIP0pmJhDsIMjV0Kr
eue8Q/xN55CkRh23PsJUNm4MFu/sWopFGeuV0RnYX5Wp9xqypiMCk5lzGJdgPuWO
Gb831605OUu2thDsdWTi5ETZKXivH56WXu24cSRwYArYBQhmBW2lG0ECUfOWnAEx
daFRB/2XlMeQinjjnPG6r86MkBbu9cEGxl9MX9D97ri5pSGodrfED7NG844bRh1z
CVimr3v/OQJW7rrqE9cdwxJ6UI0eDIhm0pUERlw3n7HQC1dkQ20laTE18QGOysgr
OtTigV4v1eCgwtiE64KVgFffgKedIN6exDOjDF/5VG0l8/Sg+K6LY0tqpOLQd+iU
ChvGhbr//dCGNWbjPMNYxOYcVjBkRQkeajGvzzZq3og8jA9e8ZRQ4AtG0Al9w2g5
4qaGmoKTDdGTHl1oIMpl4LhoFZN8qwPTjGUdxIdlmwiShJs1chiNx7x9BEpe0iyM
ofsvRQzJd89TquDLh+gAFk8NBNMaUncdPbRUMTDu2i217B3/8vPG8zlkzodB3Pjr
aFhF1eGkF1ChbXthcwaqDYzGBPLOLtXsk1ocHj+ttJNS+Lugqmzv7b5W6CCVH/6P
PzJolaVg1YjxfzoOxcl0uyGGrb7HBFtv0YucHyLL75HbhQIhbZuTnsKPo2oQm30g
3fc8jCfl1SSVq+9OBTwofFPS/3hQl+A6FT4gE+nWG8/Ml7kBxCbOuy3mUaXvtv+S
qMjcHL5N+UrJUz9ZLOw9cjOt6+HzzBEwBMT4MUm9GDMt5COeJqGetPg0zGQDg9P6
3CtSi/aYZmKqThIau2qzLWTdcC8t1Ug+jJbY7h47lDdBExAWmyrCjL4y7PCIyYK3
4u9T6AKKY6/wC424uta2RSdW8y7jm7T4NelbUpH/YogYiKPmC4XRFOqrc3C+Lv9J
IDeB4bEDzn7Lxl2WpqA6aO//Q+fUHTy3zZxRpK8FFdp13XIH17cPoP2cQRyexj6J
ThXyVju9SP6nxFxNlzcXxQWckaGHJvZJzySqpiZ6A6MCHaOpwzDqoyo8kmZJA6Q/
h08xEnZntm4sKgTpEL0Wn8vmA9hhirS8EmWO1PS21IdSAyfq4koMIswjk3xPbzaR
JgDjk+4Ydy4YS77zfivYSci5Wcis8t7fbBHkd4Exr5O1PlYiyHLmV7crwL+Wbe0H
RtFq7WCc8wnj7WtQQRGR6OJUbrZ0f6CgmSsigg8W8L8lfnxmHV533NM50F9kbq+9
Jn6pYic9mlxk+ncMifbS/H7zRuPAWUogVx8Tfqq0ac7uMYUSfRKBlwrIVBjcCWWz
n3PSoirjgjCeTAID/a4hi1NHgA8AkHKGb57CrZ0+rWtW+BeEoX2RxXegwFBjEQew
j9npxOALj/k57BXM5OHhUlBdI25mRIjI04VEDZ90pf5YEiXWSOd0Yp157cwObHlD
LwBfIrKp9I8rz1U/sFhHCVse1HtAJRRR2XOkmZvrAZxtYKTQKw7xQtdBZXLkTZCN
JIK3EXjF/u+9estnNSiPAjAgujs5EyZJ2PFkvL4sPxIVH9IkNkeRUoYpyq+yL5/+
aINtMAwa89R7edKonkJX50QTrAPP0SIY5L2iKHAO1rEcnEHgP8SzbTlwGatOG6lq
7BcRXV2YCMzmJip31p4roBDu5xCJXKmtgEr6SFSBeJeI1QiZlYSa7EQWbltfpjN7
Bq83Envi4INZs8zNy8hnkOCYKHF2V4oVa8GODvAc9WX3Q38i2vK94+ICo6Zoas5i
59LWeJngr/MRAg0c0PFXW93418CpnmIh2vqIdIjhAjOAH6dbKdkz/GcZAXgr6WjS
Gd8ghNe1cha8QVBQ5dFlWwio6QrfQ8loaDxzUlXg2mY230V1mwYhvGARpHkDbBhB
sOBrdYnFnQ6CoJM9TuwTmMFNQFu2BUN5nu27PjeZ7a/iWs/QUHuUl73rE/RSDkZw
16op1OTCNrMb3BCcnFq/SPyqauKXmkgi1ircEg7MJBoaIEukMPEye/CY3mhZsQnE
NR7XhEX2fHq+iXE57lakY43OAxFKdROeteA3+v9lm5foroduuUuGfFgBrWtB/AIz
EBcwKyXO5C1Qox/E3jU4x91EktEd/8Vj3qOtRnrxpGC5Nrd70ksQru6jr+GotANT
AhW5yh7WJwR5VUmhAFyZYNerzT/0Rdif9jXswKu+wKIvSLqQBZRDmtUFOrJQKJ9T
yf0PnTvxKitE7R+61nntIRN4w/Fk5G4JGs6MMVgqaHGOYbF7momnXFzDcFA+yhI5
VR+xAMbaN7g3nV+L4LeUheXEuHzy55UZPQ4NVYVa/GMcgp9oNESx1nVK4x5v3TH3
nzEGXElqM9UdShv9lFgA7zKWzyr+Hk9lH86ubyuYr+aIOCqXhNQUCQn3MAMdQgfb
HQSi30udVZ2T/KH+Ujli5hfNDNi4WoKHxJa8YavQHJwCsrXvN+9PnoeIZs385SL1
k9TCrzHK7non8WW3lftfeL77F5WIO0TQdzUOSS+2As219O9G2P+pyRzQJWeBcChH
+QB7wRIwQ/j6q4H5v+amfTIUfg4qbRTVjNTYSxbYO2x8VathGcGgcs5xIQNc/EY0
UcIjjRFc5tA3wXKn1AXPUIRYDT6x3t23hltRmMemjIdwPBmqcg4vv/cQUY1/h61a
mQ9dJrYFgFcGEVcf1X5rKP0QSXuNmi1QpMrVGBf43b6vZ1QgjkxSRmrvlQavSPPO
vE291ZEEwDneaRGt2UFwTKS0bOfyI/WP9RWW4FKkMEYcdhF3JRr8JxuC3SKdqtcq
NssXsjglNdusbwagEzww8sUzTETFKqp0oaqQ6ZxEbo2iM7s4oL+LELtpOt1gqbt9
UgD6IT3SysgHKiGKTRUiKdDNEINt2O2qcXdg785k7DRKyIq985TumH8dM3Q3xihy
jzuprQsldjkA1/0d9WIXYkUo3+YAJO5anj0s/csVBqKXiS5/5M7CKicjtXpn80mE
ywXd1eQGk/rORRiTzc2oMhho6hZtDbeG1TQiZXs5Lh2SQALU1Pw2i7SN6bPQXN0B
lEeHrM8QKoWuu0dlIFk2CuI5ejeJDQ8ucZ+eFlrZHrebvO9LkvbDpapRbv3qDjLf
W1STnJnJpOqUEpQR1EgOrpi4nkjze4waUX6GtpkZacM5Ouodry5xpTMO95JIiDPB
blyKan7JX+wHrpuCwxMLRHdp2xBqj17R5LsagrsSx0VgLD7fMeITgp1wMYRHxqYB
cfZrU188s5eOEkygX+ByqVWxAUvQXscysMYXmIBgN+G4Z5eI2yCItaq14LeZbiI1
/HRegP0SlI6O1uWhCCckylCnQ3q3on75UKBpEdQUWNli8EQYSvrkjchb74dzSgng
kCNFe4twSHKZhq1OabF4ptWQq9mwqNzFnj8GtCRDeP9b5DuK72OMYAOW4nNdPUUR
SMQU5mJWWfY6CDCTa2CwNwPBotV/5tyxWERVwZAgeksQOYzjCF2WRkpsZ0tlf4Q+
G5jl3m9wG2lPzPLc1ilb5UhMak8TWC/Ft6u0e2klDWUEAW2qn0Jom/3kjBgtBaGs
OC2sfNHxsfgStUIxkHE3g5ngw8mkVuX3w2NDMwvaycO/OpvICIbKklfxKWhV0Z3/
6Hy5Jadc1ZGPF7fqwmxh0EgVtSU890Lv46VkYbmeQBfFoDnXgv4Ys/OE4CV8CPVG
o1R0FwI7pND1MlvTV5dpIgceoh/1dgcY27HjdzZ/5dl5dXXFQ8v1nKIFCbk8K32T
u5Mb5cwQVXgiENiJZVvmrF+02KlZS1czllyJjsJZiCWYlVHni6FlXVeX99051E8H
03JQdMuCWgvRyZ8qhqXnVaCAHgdrejoQOkHCMr8bphCRKgw70HJBJr916A+oSaIM
p0LUnLWNMnsq+0R1fMOsZLVr5/+iaI5D6dp8ReDSMqnOwesekPCko4qEesecGamS
rrncH9PKd6Nx8q6r9AdJQGcpWHODw7qr65C/wBzhmra5TuV57L5rM4a8ZKm2JWHl
TzpkZpbfaQ25Pn8n3/tJpkeiWPHYx52NNvNvb/Uq+xiDRYS1bLWZGcz336wFOYuC
nWEVXDcgAFRAE8hFm80lzsfagtSbvuE1D9kkzXVVQlfOc0nvX0nzs+NOrz1U4bts
6w6644u+PZS1Hgjc7LshHsTb6eTOHRlkVgcsg7F1hsu3fygGQDAHYznX8TLMAOno
Tl0CK5Lk6FvoaQ1K3zo530Bp8XA+z3lk8pK4+SlHgAFXfoUHw3qnchai3EtdAgzf
pRJtKtqVxPJ1S1I0CU7Mu+cIaRW7DsdnAP9Wfpv5vBElsKm1sdLNNGNJqiaLKrPU
U32l++xuMAsPt2CgtHYuEDOR359uT+6hbiflLkztWpe32jofuHHZzP+OWvTufSnS
JQjNk31yhuHBrSUiYF7x1sJNnSrC0Ov7OBxSSRczPkLwla62GzUPiCgW+r3YwTIw
6BzEdKdlBFX1WrojI4J7vFcX7d5fuFpL45XQgtYHNyOHkDNUfP4vexVQItMcnA+1
Ri0+Rl5gQiCoG6w5lFe9G/cay5+MdCPgPTqiCOuyIXsu6u/AgKwu9b6tT88F0s9e
THbA7VZTxbtTFTaDWA6y6zI7hZKTG+mwPvwM3sNs2rUEeg7t7/r9gss80xb36M3Y
mzJcGaQsKBm3pMBX3xjnvu5y3RD9960lQJTskOhpXmLlcuqDwevB3ioDN7jnwits
tary7YbLxJ7vQAWjSvJeqBGVZZSUySzo0grz39P+yFfm4SnJgiQwZECUubwSa+Fg
G+KFbrxJAJrvb9Nd+6qHBnsbKqj1B4HHGWxGvXOVyQU4kquaZzDeTiYTiBOrcbfJ
e2yx9rldVC7yWYTJ2eJKBqU62yzFPmtDwKjXCpy3q3KBgn6tY5uPiGwu2tVilRVk
jtnKCemqw8NzpBVCRt1nXVI4m824o6Nd8mAxKoQj7VNxRjgImvluEjA6Ozddz/0M
XJxRuiJYbk+E5j3cpaFDBYzx5FvzzKTGVIWICjTe7U4z/mt9Aj2idkkfAScrSyJh
MWPm0D6AoWbwEmtoa2mDNsT/3bS4vgB8cJ56tcEJrIDaTgrd1zxGGnjkRIp0gueR
KMCg9hBJThmoNByuFCAczUJpvbxX+pgdoc39msB3JideE8mOpmSQu+tzpRCX02qT
NdErwqy9m5h/+ywTCqR8OOPqLrFa3GFVnbTbNyodoQ0OvRrkhLiOheOjIND2fkCh
zF47GSw1WqZqxV+Banq/CSplUdOmLAiZ9yH0c0faxNRB1HrK2uwJVkkGwabtuMNE
F+2L3bYIqbBwax91RcPijkwOVaXC0fMW0SjDdtJ9OPEc5Xr7/a7jm8gVEv/1kboj
0ObbCyaRUwKwi+u1PnG3spUSpQAlvs1xpmf47Iq8ZTxKRi94Z4XQCp2jyd8ZaSAI
1bB1Y25MhpfiIAuMR7QPHfbAJwpPsEe9NtRsc6G7sGU/NXQVHoGg0+YyiflJvR87
I7zxqRP1lFEPGAOtE1NzLvoN2AF1oKqKVMk5M760Z4aSRYV0yXfBpiWH+sZ+vwqG
uhQ+ab3GgQK99ClLZpj7gVwVKMPkweVlbtpIxIBuanQBxiVrm7XybMPX8CyG5O1y
zsg//5+fEsFGa8Ji4iINbfkBzWDEdJGXoZUD479c7EMhjVeYNBNpf2RKcoCHjwKR
qcf2ioBBQlqP3lccOqIDnIgt1jFtx0xBkOL6EJ8wsLPDCmQ7j4kZKuDtBB4MwPSF
wVhsdhsbKj7LIgaG4nKv6t87MXgqKObDzRPrGdHfcD88eYYDAUKz5dZ3c+bUtxfz
pA7+GJc7hMelzsJkrEVUxAu8y6eRYvw6loEhU01TDj49vD0DNl4+WlnzdTMIPZPm
hWtrfjAWf4H5XsLErB2psKnL6mwLMWgkYp1r3VwXu9is/Ur/CyUkWbZdjGWqOjpS
56TCRMD1pPG6zYQb1DZy/nnSgyIp7NfM9BRIcYAcN3NCtZPzdrh0cx0sKRDYRhge
Wy1Lqzf7J0ep7WBHRxslkP/1ObiWNSdb98/zsM+gQWPLpCVGNtQZv/9k4EUQtMOv
k3FU2sWPt/+OPLYxvaDjnbSMLgh6Cbo/Ql8086DM3RhJlwC37ELGX8L9ZQNJAky6
S14elUquLHOZ02N8OuZshVgCIeYx/gRFTnpKOLcUgxSjYyz0f7Drg6Qv0aFrM2tl
6GV/TSiRtQT5MLMlHQlX2YucpZ15ywptAqYDjtdcHM33RUUVWAF55WVC4xkkxVnj
5WurgKLoJ80hHCSuqkTVxEKB6hKQaE0ZI6rFAr9HLSI38p58r0BbqFVs0PKH+gr0
NXJzUZizj3pQcdGu14jOpkjPvriVRgBERenbW8s9Fcahfg/OHgNhNwwLapXgz4p8
wgJxo/KOADqd2DCG1oQPIaGYjCEMuqG2yefWSKhjh7SLjUMnC1YqyacLamnmAPUI
MgX+n3S7HYII5R4pUWusL4ZRv8yxT9/NJCemzd5JnWPT6s9balUQDdzo/bgghNdI
qNpH62EYaIN1gVv5IdaAyFYaGyYxvXL4qISlZlYUveJTiiOR6FhVrEwO+sSoAgq2
7sEa1IiUaLMdoSgJovM+3OU9SsEDaec6VdBPYMxEIheh7SLZQM2HzVT9owFg0L4j
6rey8yLUdEoILxtlrCEkd5+cou/t9jjYlmvKFmC60YC5NbZ/dSKVQTy95Q6R+t4j
n+Hq2UavIbRKiNKxJVLwHodFoacqUBFRaEgdnnvVj56+sQ5h+vZyc7yrkplp3JLP
gwnI8Vawsz5WVkmS4NJmVzNia190p5KPZt4SJsUDOXhsxueCE9asUlaPCiM5LInA
9sdb3yrWW0xR8sbEXdjXd1cup/wlM2gUeyEBPT7Va7MU8DeijQh7wmxuPLTPUE4x
0TKQdh7Upb/LH2dOgbH0th24KlQ8TMwtBIbvtse5k1v5mu8W3ri4fmSxcfKkuPEL
6Pz8iKodGT4e1pvZXVnztrzjWb3LEoYIlDf6jxOWi4XsCmc7ReHADTtY4CH7QNno
ZkZItoD7+bxjSmlZKWeNCMrMbVihgWkhgWAdT7wIv/JLg8xDWwlh3TDHTs4nJP67
8GDRnrJcZvNeAiNqLB9hUOIpbkPi23Nc5QaafqMQELaKWiyc24/XMGj53E7//Nev
Ed5CY8rf37uOrQf+IH5CI15VzGPClzqbWaFzOdNElLgRw2WRhHpprI87IE4znn93
hfmCS3sY8OrLNOxvRMNdpkFwTsy1OB/E5Vd7K17s5jjHtgFNuhJNGqjvd1YAYUKA
vznlu0C45k9vfNVNkcyEyEGDMi/39rREDPe/qTZOesFuxfC52zmRfQVqiMCDoqww
ZBMBtzZK4Md0t4KQQSDxICvDeU+oiSvidMUIfo05bZIPaLQEzkRvWASg3BB7DRpV
T6n1ZE6GFC2AO0Nn20fsXYkbQgsWYLe2xmnrwrY5n9QPX2HGR44nuSouQc0jXScP
Rwp4MvfZ8dTWbAJokNaVXksGVf+yeMUpzg8Qx17elVmT+G0wcKZO6qC15yYlbWxE
OM5Cr8r4VkrpEIuNsrHeK/JMN8BYnlg7kHqMay0OYvUF47ujUsI1n8ZJYenaK6KK
xvVsr+jOC8p4HIa4yO5RIXProyKm0p4e7tKpW7DrStIZSCSMh6yvrrRB/QDf+mjU
d1pnuPeEkXgSgBx6SJiHFi4E83Yvt9HNQ8hfitNjkR9w1PhBjrVjUFDnuXW88/Sq
8CqRnbQjXrCJTMrGG7BRrxFygmC32+UhSPScprB8Ru5X4k4jJ/Vu0f7tsaim5/n8
I3UrCN4oWXnnUeHYRJwaQtEOsEy814xqZrMoSUK0dwkwyOE/6jLkmFbTEdaI1xZI
C8F4+FguSRAl0e93vx/ZlbTBHnedxrvqWhIdwB8jG45nknaigQ++uv36St71vf3H
IolxKuRcBunqptaeWVGkeFpfkOE26IFEh/tuUDXpC4d2nNaXESzwpjIN08lfBxoI
PHrfQoxIsljeGkKgRVdPWqpmReD6FePnNC37FtZDde2nZ0LCG7XUMg37bxmml7+M
VVuy4SaA5KY0Bi4Jl+R2knWXQ43Egy7AmrlaYQs3bFTq7TkRIqaIxnbkpCgufJmD
XPD796lOdeFgUz2v1tvUqINwN6Bgb4H0aJsT42VTFXmQVjfDxyFnjoMVnrwuWv8+
fIIiFf3dJKrt2JLaXVp1tHiFVIaEBwILGDu0F0+5zV2LmwuFQcQ9g7twYq2p1vVe
pNL75G3t5MMkEGc77OL0KL3ytxg3Ln4s99GUEkn5D8bGwlz5v0qCb18T9X4Y3dZM
UCxTlkKGPngQKLUZ3/5qOmLeKP9XPIb+t0z9iC2OEX7soKtYfuaMh9FHy/2+Qdj8
KdH0OtubuGQosLSPbPcbFiuQMvVj6OWslKaBqIE5/TN0VQ1b6rm+LVqmkLY+iUB3
4BtQL51rzNa+hQPmoweBay8FArFNW9LomMEsEFoDzA34cdHLlU9OSnx78WN93Jdu
xR+OLbJc/BLByH15Lv5elxJ8095dekYKL7XXeRhM0Px3cLXK45zjKVAUu91COCFG
ly7u8eJIbqj45rmeTV4KyoGd4pGLl630OU/NQb228lPKCB/F5yTKSCh3VvKLfgic
iMOX8j0Xc72XMI7VyD6KuFu11sjYXuIpZZlTdUnYi08xHXt5rg3GEhXLfLrQbw+o
8IpB7nERCiTPxSzmeD50s+Ega5vukzU1kycdSvzMl4McmxfLXnvAQOMSIalVipGl
LPaX0Mpyw1Hyjw3Dy8aB+PqcB3/wvocl8/VRZJrfKa0pS9adniJONrlIx2vaMUfb
fHsnVLWlnGemGYaD50bAPn90J7uUpwpArzFAGSop9qN7CYoDbmEpBo11ZcgimC0i
uqrrfXjL2upYv7hF8aaluIkDvG04V6BvSAdEqC8sXgNSP4+VkhSmjKiy/kkRmtws
Md8u2cbu9KsNhgW7PvHXrLjyG9vaeusjHgejSnbolqS1dM998vq+yHe6O3bXWIyB
pBmW3HxcfcjBofslXbCbFRde8pl5d/IxtdE5Cd6JYJBU4gTebmxDZeANmOdLqDur
/eJdKouOTZWqXu9YsEImhxD95Wef4xa322lOvqBAlCpOk2TDCR3HFMzRADS5+oj5
dnqBC8GMMYBSNba/Rdvkg/+3R+HQw+lq8TAhIbGBQZDZ3J1U6NAODiucMCFrnTpJ
rOWyQIh65rlYnfN1m/pVNtLrtNqjcKbVdhix52gGHlG0JeJI+AsrA2B+/f5ig1as
MuRL+GTc0YTmfhnZ4R3Sfo+uN+v6wnllWTbGOG5GdJQF6qHo1GBdd6/qJgunDKmB
HhvrpdLrr4Q8BA85pPd6cI23Iu6QdNYw/sBd5BhiLaEtTq4/GBACTjLukQWnr860
H5afLVsIgNhrp3jT8joHn68RHJZwqg2JHDYypY/7qKnB84fwGmtHJh3dMceduPAs
TpxwLoRG2y6DD8v5O4n50Sf12KbqrbVjL02MecfuYNl33SuwOc5vik8WKAwR2GRe
adB0vaqIUYYOo9VTQSnOr3LxwdjMq52RYS2Q6Gl0agXrBf5UwyB6VkKjbLMQPL1O
LoBfdGF2tnNGcuS/cSB2yK7zz18LXzV5TwZQz2IG161wqhsHL9KVCK6ftAYvn4Cm
pGTyGocwuDJEDI/FMsXZRy5kbEjA1reAZE5A7Qmo53VKm3qW0FXybyIhgfiZPfkM
x0jeTuI/XxxmeIyo7KpnUAI/f/twScHdBMJi/CmVKoC5xuQeOjMl8hl74IvK9cIx
xtNxoXgh/n4DN56mLzpg7x0vObGvsGlBkdD+igkId1U1sHPNFDRa5JLPlhpdhmyH
x7vC1cdI9CyiXXjQOcM4FJn2K1v7SZwU2XJhMInPkio7a6TK3nS1e0Qb4nHjHW55
AIvyEPu7MN9sXNvZ582bLmnRlc1SVZCz/46UUdRxiyNvl1yt4KJEoezRtlJa9ZLE
vHRARsN6iIdkSKGwp0yF42JMzXdv/N/MwNciFOAganJcefmzoA/ijPQsGiPKCanM
MRgDY3bwRQ3fZ/WrDzvk6U5saq0RpxwDEFGBi8Gr9s7rGCY7CuxRpF6lx8ky9gBL
hYyX2e35yyKrAuLct0QghkXVf1tJslq5i04K+JLW3MxOoT8bLv+QUkZL2jGiyeJ4
CQqHGjn3Khg6wa5diMXHD8QMQS9jxVf6yllsYAjCpLx0whzq6v1sgKLvAeqaavEj
LELFLBSfB7iedCJplmag9ihgYzax5gefSEtwJL+6UJrN7Apcg7FrnCryA17T+IRf
p8yWLzh5tidfbqJ0G9sX7NRdDj/RfKcaP4slKsfnut5j9SAsU9dr3l19SZlB0lTd
S54sENLrTsXarg1FT1SJZ2UzuzWeIPGyE7iUQtIzPoIMTsOKQ5TR1OadojDTPNYM
HK14y0PJF9UjtuDgpSOSuXgd/SSlGony5LDNJeUK2m/8DdJT/JaO6Gm7wxgRa8Y2
`protect END_PROTECTED
