`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BuUgcJM07z8q1C5+GdUeoXPYPpPfwgFmAm7HYkQb3PYRcTNS4svAjHW9y4WYEsNE
ys54XNEhUZAnFMGXgP9HLCJWVOewVSqMjNnBvTtk6yAnA0rvBkyvVjX1xDFOJQKm
HenhUicjRADxwq7ZSABbrsX+VG5tB0wMKcWPzWx01MFARW7XvF9x+YveJw3nK5jN
EjWyVyJH5nfx79gOZyPl0RXikZ8JbFXRNe0/km5YG+DvR1mE4LfVuvJ8PMsQtChZ
EjyamxJxaHu9UI/1SRE29NRNwmNjggCuMptvWBlxpatFg7xIdi913Rxk8yCKqYaO
J7NJJXfnmk3cP2DBT7NeO3oio/oCCz1xavym/BFTncSNdJjUoVRiuiC2AAnlAh+u
4fqvf2/yyVUUwlOIJ4Nak0VMrHLQnGBEjqv77Rapo9UkUBM4IVrTbd1iBakM4MkI
+EC4TCb1ui7aQyAldI6IcopjGOz62SxNtma6jKzw+N0WfMNqsY/ReBQ8Rmx6mJnh
uo+WUe5oobah7P5IrZ+xO54V0SidsiPEUgj4bW9O2B72Zs6RPF8lSbI/tDsRjFX4
wHMMTRtfiAavJU4eUzuHN3tE+35RW/XM9oS5bBiEqseh03oZmPRNMXLw8oE8lgt7
pEECzHdLjWEoWfNwEfIXM+GZIUqM6TH/T2uqhurB1ro=
`protect END_PROTECTED
