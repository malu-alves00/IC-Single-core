`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
K/JtS1L38UZkk47BXpCS5x023JldYgeOOtMj179cWKD8DzqbG/eiN0Nb39xN3yVG
vOa0eR91FSrR5hxyG2TLieKqu6SS+bT5AuD/e9BeWlUUHnN+LHvAaWPl8g/n2BHV
ASOVtb47fVhUbPp4XKVkb7hRACXAX9ZWuNjuwydVf20hmFyCkutL59xpggFzOEEg
JcyLMTIznCdICjNNGDBuClx9M5PdepHeQmUrGDWe4GsVsj0y24NOR0uz7vZVsbLv
AoRYmTeTfT8GaAJ2JiVhgN7/1LemfDUudUSBiESQJOjL0CJraKHaijQeufN0SO0J
ar8XTEwiPDw/SiLgg1yNitsjy+sQKLuVkUAB29svEhgjDxQhNEKievd+wqEdvoN5
fk1iBbpbov6e1tpheZaJ9qkd1O7eGknbyrMjl96Jv+A0ZIZQiUj3FE7fztN7uJ5t
sxJEOjS8PNVoc0pn7tFI66X8gSdgwT7g5U+9TDdIp+OanouVdXcfw8kmU6DBsPmY
W/fTxdgTFIK4C+W1izhHdOPBBgvgH/k5jcjRvTobB0L3UANBRMsVDuj0cE/znkX3
HuoWFIMY0nUb0Kl/azvrJCI6ef34CJXNjwwFvwFCrwjVH8eWGKKau/rnxIIXh5Kr
vmRWNWtoRg3MNntdTmKOdtSGrnjJikz8VonfajUq8rFOosphJ8o0DcAX/lEVOh5G
bT1f57LK4i5DfnpDXGgkvsZyJQuPvBszSYqlcVb4DMDVEkExh8jVsbR+casAgs8s
mq/tTgm7ksYcuGevahTQx/ayL00TrxqIVBXRe1+VK2zde5Dq3c5AcISVq0mI36nU
SsjhCBQjogshDrYhq+753OtIa1VfXQPH643maIgYJNI6OLvdbTFGz/d+bYjYxM32
6hOxsEkjfQ0dopJpkkbUZHsDY7/uXs2wISfrPBlIpsC1LTiyUfT2303MQ/qoAeRN
S6hoplDZzumpsaW8pzIcLTl4PlOCv7aiD1+JVOwnTVrWnqqjmX445ZpMghyC0EsM
2uwh+s89aQAYSxQCsUMIliKxWXHydnxJk0MURofdx6WUsYraRjWCBH5MPgYybOKV
bcXPQifZQdzjtaAWNCFiFbEOtZpWt9UlvIp2WBFOLugGUnY/ScgUnpc356+bNZgx
aPlL+7vxFHp776/IBH9wpKYKhRwi16kEhODariTeknrUYDAWx61MyT/q6EMCUZFJ
bC86XyExgm8d+UZCIWpDPGmfVeX1pe08a9S80QgcuN6z/1L+0hB51/3NObz2kvbl
IWcegW80MssZg2X9opFWvZ49UXIxQpzMb+IydruUFbES06Af5CZbuhGcjRYmD3l/
yICoOUHgSOXUBhArOHN0KMMFFy3dAvyhfyd5LHuEqbBOMBDBkUTJKcvmzCmh0SuJ
lsJk2CibRUHrES1yWnlLrIVGPSgG3vyj8qVlTqxTW2bbfi2avhKXjssb6Zi0PdSp
uu9gp9a9MeCGoUYIoOkb30j8RPgA+AN7lH0Z0fQWqRMdcDQ9SXfiYYJb+r4G8l2w
2a2Yz8fdck0vGUHfFR8Zz2lKQNlp+yMVcCd7957IbP4R2qRh+D3cBPqbTRgc9AKg
zkGs+Qs5DjM0CK2fIoMZjzxU80vjB+6UzraNno9utWC22prbS/bkSKHReMCK4GXV
opAzRDZlL6VytCdQK9E+A4zjPEIMgx75LFX7nsAqIW5eGptJl9lLWOSlqlQhc5aR
+5sEiumaJe2WOcSoavaDeadwciX5Y0LMRwlH1A0RKm+SY43ZB9eIoSDzXy2x+96a
UeeIupNEc0zZ+MNz2DiPqj2tV3j89xLJsi319IATeGgmeM6QrRU4IyDOt2+KFdm4
cj5u9LAKl27cSB/oKO5EQk1QpLKUgNrud41qJEdK/vf+L9FK1bzzG6LIzDBpqaLV
6OjUFfv5k2mXC+6GNdFNAYzGUVIkfqUf0bLcnhEwsGo4mjbMahseuRjKHyJRdKXv
6HQoeh/p+/VNHVAHk/f79cC/VoWqv7y7wVzURf6tY2Q+Pl0ngDs90Y3gAVzm83FI
NVjTn6ZSHoq0DMl8cU4zU8qElcVx0jTmmmklsv8+hFSMFP7vSHdfiZB7U6l3ENUh
6rjN2OZY2/alNYAo13fnr5qCsVt7V3sB+QZ0wWn+Ig2gwQCREv25TaNXpEqGrcoi
jDSZfASvziFft3ZhvCpkBvPWG6XnPBWr9QUAHZX86DVxblEmm2U3Efr6tkwJQL9D
V3jhhG9+rrRtmPwj1/k5z7C/7BdzJUpofyQgmDu9qdo0BRoCDAQadGplm5T3AiVh
4M/jJ5/2nPawui9D66qjZY+YYpVfb4V4n55/nHro79TuUtWcOCXM8EUb+oMNh11m
Mmbkw79OxRcpTpu5aTcS4k4kCeB1hhWdoOWJOIBKj/TLzQbmjjAFyYwJZZgLfU4F
tkIEiLL7XSnoZGx/J6cPEedr+GO3WPQfKoaxBNhM57K3eCXHXA4H2bRNhPELHf75
1qdsifQ1+f7f8sgmSRe/iWvzlgB19Mtweg8nFT5kO//NxNyJBRi2wdCSY9UUvulb
SHhlgmVB4hxhIAclICgwwLBq3CCI46Of7l8ZF3wMjjX6PSuqTLnlaCwzPJsTngWW
a2AGF8C4BxYyxqFHCoNPTprSVikRw/eMUMWGczgFMAg4m/Troj9QftJf/AoLteSt
++sNAtqhlr3vExyuK5C8rKACeDJyGfyIG7mHJCpaTf6F6ZnDaHzDP2K3GlswPZeE
Mcb6F04OnzQ5Bx7la9nDXDPG1ukDKnKLQ0Fvk/9Wc93OQGOqhA34+2HCE2suOzax
1HLAe6QBKZKdzxwz8Q1FPdF/Go/haADEaIzPFx9I4OMA7FVtQhw1WzANyIBncV8G
0nF1yK1pL3o7IvKcATP+imDDm41/u7svRXw614/MQrCzDaacbRIH6f2284eRe6AX
wFm3cG/rh/QsalXaA0utuTZ+NipVZlMdKU28/SlzX8PTHZHta5DNn4BR4Ulh6oxH
MFrxCvHRFDElwb2TGSi57gzd5N40ZTzv6FRj3v2Kds5ZxT/0W+OpUo0iF6aCFgUg
Iot+8dneFiuN3Stu8IOp5peMpZPCQrg+jXz8Qa2ST90y88uvxxA4MnojeL8TJpjo
rPEAgIOZGqRhOx4iezOJcRfWnhEOeEptiPRV0Fd96awXeNJNqhVmyKkORGVD9s4Z
SaK1xbGcYpyykOtUhMMeXPOA/zLwLniY5syV/M/VczELekWs2agjAyn2nht+ODux
HpgezGJ1OtU47DWVN1msDD4iIFLEeT0RQ3znC9Q1yYTKkk1xStWxToyWCatnSrVb
vib3dWmvDLkh0la1Fv/bcqO3h5+pBITJ/GfDeaDdNTo+u2pnrVHDyV84M2hOFI+R
r306uN9CTGZR9XjAeyzhfrEjqJXKc8MyVIt50YTueFV/AYjQ1AoRYDrkZfjMpGlx
fj0oSELtG/T8RN2lQgiDO9AXe0xS8PhIPaSyzw+oOvQ7uwBm5UaRCID7n9Xpwc9N
O7AZ1RymOkul4WYtDx9UMuuPbgRnxZA3yr9mptUDwsAXBNiZMJkeRj2DPsoe37tW
jfytJKtxsVImvfSsokR+IRq3h/QRRqGdTHZJo+vb/tKBkQQ39GSe56LkZqZ7xtOP
8TTqFeDN8sDq3yz9+KO8IHtcycGEF5Gaj9ex/xQQ3Xs8q4xIGajfGmtn1nIBS2rL
qJ4ITkxfEM7YoiwasC17kdlxybwi4MA4SdQse3MxHY+Aa85ZW8mTh06ztlDyIgGk
8eBo3LtoX1khY+ooLK8tsRrJyFL3HBiI1DmyoTxEVLRnt1ylBbkkt23/Pk/CFB6K
xccjm+MJS2H84vm+eapy6Re8qLDJBgb7TQU6FmctTkZVKc1lrfe1O6z0cO48t6E5
/4hzDdZorsnTLWDnfrwONWp1xVOTMgh4Dmue0acwoo6A+twBRUPAZ+Ey0aPcaqpS
3/+nTH9rhjhxHBH1cde7P6jffF2dHTXi5np8x/3qqE/TaOyduz+7xVnd3MhhDN2D
CadvQ9XtkDStAdOKyi95zntdLAqNTW2y+9cL4LDECSWLEkANyyeWNELU1G9UHg2u
5b0D5lcB2x9EG1zrIQcCefcu3/Q2Gf7t06LgSQMk2QLTglMt17il+rx6TmxFfZtk
942UgD3tpsp4QP3hwy6/DlwDF1ic+ycm/T4asawmjwh+G9o3D5m7lGqZbC7fxR/v
gQ1cXpOUoBrI1pqoUuAbfWwajJ9QtigeNOmaIpR2n3HhvJx3DH9NaJGdcqnQbU2d
7+H6MjpcUlJOSHydsVRAvhy10LwFTO8QYnxrr7mPOjw8/W+7FCS0/hAme/6O6ELR
bjaiEDMvlzaUpI/SzmjX6qzGNNosNSsC22O75WeC8LHtSJCYhKltZeLZVsIRpQLo
HQdhi3gloNO0VRrs4Kx6NWtGU6mFgbr7wD5TtXa6+8afwCetg9pv/3AWBJ7Rb4pa
Z6ZKg0iqA5iin+HOhpUrZbtmI8JeKw0ZBzw/dbaahyY693xMJiyhPN+SX8L+AGbD
4QJ+P5cwB2OvkyK5Qi8iCrXm+0b383QlINhKmQjgxFl2bm7Wy72445TiLG+v3zGU
/n67+drKwOvRGlmsxdWuqnhHLIh8up41uALD2q+9YvKeeHpPi8V0fVgQFmij9+nu
fPs2GMmjwKirLrxlwHemhaGEpUfYFBhs/9Q61ugnrNqamMTWJDO2okOirqesd2K2
L3mmvHeuAY4hFvffNiTAxL0esAgyuUbGPYOSRiUMcTO2oyX4FbyHylOr6XXHuJ5+
smYqaflZo484hZcN4BdwN9vamrVU820facDAu52a01ZAXIcvA5Uy2ZY7wwJdXMte
4CwDzPEW5Xs8+yTcvsQCPMDUr1dLQLMZ6nlY7Mat9cfkk56vNC3Ei5qYP1SDBRZw
rjO4LsL4ECMuJHn8Zjpt6sZsfsIves8IO+zRo8l75l59b/NMY/FiPITmuxD00cHA
xbUfOyJjsWrsLpLL7+jUJANrj0oG618b0DEH6y7DD+jm6+rbAhvPWC3Ap/FyQqj9
SZZc+NNCSPY2eFiE6l35uHvicwcz9rgW9aYsNctMyKpI7Klf5uIsdR7EWwaL9iC8
cQUrc7C4nvweAhqlt0jkxblEPER8f/vbSbiyATU1BgGx/W49t+iaNFiHd7GRFXdp
/fm1v7TDLm671rur9sySKbSwhzXoMuT8jNtiZPUZETfcrHmgJAR/B7pG3ntjbmU+
ZJGeYP7S5EHpVRYecvkLN9hY+s+AeLNO+6swdbqqzNIowk0whX4kkATid1irtGgX
r4IQegUgk7EFXfmVVx6CmlVEKEyEn0DzOrdilQR/se2WnKKL5wu6j7L6umBH9Lkt
SuEthbsLkhIaDMLxvB1WO7Wh1xVj5MjRbmeB7qziZHhdK6DRnZrIHTqtOsd778HZ
eoQFD+UwP7cwudB4N7s+u4vcyEddO4d+1ircEBWpkXj71TMzGnoxjAh+AJUwhmuK
HsOb2TvOLKyFfMpQFaYIXtPncxO6UzEVLJ+6xa/On4cMT5Jv+JWQThm/tSD/H8oH
jJIRQIzttJnURyKGvqmF3F7b4gjaqxjOrD4Vgdh7I9OTc55MINWZVmNpIFHAFSOk
emOO8of1MLlry4yn3cNrXvY4TUHOHkzH+/kDn48qplVnkuLPI9JtMq95JfHsuQJY
61PWLkXvBfZI9/8N3dxf1ULrGq8askw6OysD56Wsk0Qo585Bd/vROdqhYSEjfiXZ
6LuMMRLFhfvBcyhu9qEjG10OV5eLFkz6alE0lSred4DMPGpBkHxi9rorgGJWR3tA
kfSy9N5HCqgbcNTK0zbbaFPRuHEeFbsBCVaXBk0qmO0=
`protect END_PROTECTED
