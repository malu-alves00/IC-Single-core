`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3RS15eM2HrHSz+BGSc0kiIrqigG1XIh7xR5JtJex8Cv/pCgSzcEYX3OL+AD67NRZ
Drcnnwm7e1tkIaosWV72uD8rmGkSGOcL6gzADq5pGyRQBdEn0aGN+bOILFqFfAc/
xfOMCfUKNS8wXfZcz5E67EuNyBKLjFm+3biZj4PtxgGKYeYznAO9x0ad8Ci4KwHE
ZzeWu57HQofQ9r4xtifm0qLanJU+uYu6dmJ055u2xRkkgln++BE7TkbSJSzskUMj
QTgSOxNwn3atzt2Obn24FBZbgUAWvbiwZ2C5GspVBOUIlaE3u1Zm7SHvNW7Jaiea
kyqaUmaJnST+ph2MF/1+tHW3wIQ7jINgbyYhw0huxZsBKF4t0osN8fu6gFoZVlZ6
yCdaQyzjBl+1+tvLsBChliCpxUhLGBjO4fLz18tx1D0tcMbN5sbXy1gXe32ejaqT
jH/O8rah6vv4lDGI8R35DD4nfmsiXWdftd5/dEZFhsnE6wMdB45QF4XyGnh7CrPj
+5aOSBxnxmjgK1hP6uZoKOLQ+O7mVjyKi0s6C9GBec/VcVjgalqWWH4WNWuVgB8u
2ojGeXKh8wNmDFZoxxKzFXw1uBg/ybP0s/MwB4Vb+apTqNsYndav+EvAhLBzO74L
bYOXcoy5S9Y6j67tyIFdTi+ghIXGly1Ob8Vj38X/HpHlGhY5uLyI44XgjGnPsrHU
Khqqwm8L2tMIXmezTo9UVohDL7Zpb+/zg1C1grKtXXlT7eTvfkOppbdQKrGIOC5h
r0IJ263ALhqUjEruljB+mU6rP0pOLEZMVESqK0yrAzFe3WhZuwX8lDr2u+ncOhtJ
nQiRmmwMNz740w7wh6XHVoOPCt486+Nn2OVdlvrW1x4WqNSRptJg8DoNSYclqu/d
IlEh/JZOhPC63knPVECtEKlNS0Pv00jxnfBer2kBBvqUjrdlX4lZZ5EcfJMRTEkm
QzTHeNHZCjqMzik9esy4ZKLCPxoeYjHBpf4cDO9AiVTSF3ul4mMrLS033d+r/kJw
P2n4vMMOr7Egjm+HN1luQMfdQXF2jpva8x9l6fCeKMEtlLjlKsUsxL0F5GHP+Stm
Nhj0T5PcemYderwO2dMqKh0YIdfi6F1ErckcJpfdgNnu79J4QqnueFvJheZuCZyX
dQCCSSmtC2Yv44sLXxO1fgxeF6HmxxcM7wyNYLwrAgVoRtrjfR5/R4CWAOhAPJfX
1RMlgabe9GqS/8/yne8/EwV3OX1Lw7oM+SNO4kVu/NfwgCFdVXt60d4pwYqvf6XP
mV+5pYFT1AnwDLaOS464XPVX/QLXwDFmpmOTGieC2cqRXaClApD+GxxeJuGaMeOl
R5NbjizVA4Vv3G3Ol/iEYp3HzbmTrju/AbpelHpAMf5GHyljL5OIy8kOKdLHpUk7
`protect END_PROTECTED
