`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Rj794v2/3oEnIzo5p+cZhcQVItAHsHyg9YQrDhfyLju6LcOKzBvnIjN6qaiJ7oV6
fh9nQ2SfPt2BA2OQNEO/bip0AaH6p7fgy+VzK1xWQ+VAT7M8Ldl0Lcjpj+0JiMAH
9pmbCkSarxH2SgmmLPP2sBB7NWPWNiW5u02FQr9hGIgAoQnsDFU2BIMrGYPj0JLA
88cAbcnJ3TZdcgNGLnFa+hp+/OmtEdW5tvrYU+Mf8XvFueY7Lh3PJdYJlpYA7dTd
baci92z+xSOGWSboaA9GRjtoUHj/Xh4UtF5fxLYtkB4RogDPKrhn5hO1bbL60kuD
SetdDPJNqkD8h1AG5nZz9Qo6mpdVjeJ2pvABC1Xx+vv8AcP/WgbgsK1bTjY2KIXF
8B++jMnmBh4lgGPcB046rx56ON5PBu82hPyMYi/XDUqxyAR/jTlVKWjqz9OoQtfS
WJzSI8ClOP3zM7BlU0ohaWaPJgF68MEOZ01VCxA6LSlxrAZnBIBR0sNMMbT+W7iY
janXuGFeNTC3Tf7WADz0jIDlouhgv1XUS7GRIXqxDZjTW1ZkHDOJsjSvDYvjAodv
8CBrxhXRG4TMDh1R3d3N9bsxM2a+TqjO3Rkh5YU6xSKKsLae13YVA45Ma0nTORC/
HEJFZMxHfnLqB/m1kDn77M8F/MBugXo4j619ISAphyAEUzeewbo8CmfDGGx4YusU
9nwU62BJc/WJK91y2oSmltgtQM32HYhxFaEPdPzpkDc3v+87WYA0DfXU4GSfMnB7
fCoixy0bZj6cJvJq0syESde7KGybcpyfYtTA5afJd0u9NCQTXk7OcuvplgAn2HZm
vJ03YPx2wco8Bp1YRaUpee+EqCzSU0RAD3Qz/lOQO1tzghFStANR2rq2lkJogEhj
940kMC8ob9ZcUT1HOZdzETLeBf51ZIRRygeXx/tqBM7hQwM5I4wMnEj9+iWMPcqh
rQmwKk2f2uO/qtva+PPznDHALgRq5+8aFSrLNiF82/fwADq0XYCuNVUQ0b1kyzOL
WL/GjUj8fC4MhBb0Hgrc/gdHu9NZqYiZkoQVyMwu5NSFucVc5Qw3CYSAcUMrThvF
J1GyKe20WcQ78ygE/a69916nFjMbGtw17tdS+sPAJeFZh+6uVIrxuJWKxwroiwbp
XZOIJ03uw4URLI6PD9bWn/j3f4KuFZkT7QPWW/SvrLtHd1nVpstk5Z7cAjMoUzJc
zwBOVILezbJCLvHuQVYr0ORXwK6yHGlWMYBrw0/MfDBFg3N+PUFL5QIDnKGJKSb1
6n0hqSrblrNagfgDteTfhBct2gWgEUOtv7irzFu0PWWXyF5Q8RHdoeS0DAwNN32Z
3Mk8kuNZmEu0epJhqtJSABEEgVWwBx5gVv5sqBS25vAhsrgvRqtsoM/rKPMnKFlp
TzivWgmXx2ePC3MpShCb3Ox4kK3/OOzfeusEEWMyansIDuSy9z4joUfmEI+jzuSh
ZTCk1bYVQAS1Cc4aVIwYJ1bAPZS6peFrG4jRRfg5vXWweUblc1dS07mQQX8rGt67
wCWq+xCxPvFcGL9mMig7nKpz84TCeDdYinnkOolb7iz6ZJR6Teqyld5Fzl+5DmhL
Dn8mqyMBlPodLVoq/dAykOsSsQ5G5vl3UNKznPO9sjmLU+UsBntdnE05ZZNdCfU4
o+KNsil9A55dDCEZyRJS5J9ZFEkiy4faJrJz02M65tY3vTY3FElxJ4H3VyPVkZJF
btsiDW2MHS2P9Y2mBN0w4GvKHBd2Tk3mw+MsVlNeabRT52AhQ7AAm0YweZw0dnrX
LeMDVjHe0bqGhn+b177+GdiVnPyBWfaP/fpmP7ERUKiC5mDLh81LeaelgVul2JLL
wfx3tV9zSro5l5rHNpM7Obv2H8HmbgYSH94fbpMOcgr1tUQdTSZubbYeIavekO4q
kLrzsC3sw3kJbCY3CYpjc2QyP8Q3Ul7oh1PVVkOF9yf1t7Hyfsc5LZV+GJfcLu/j
vL+ogLrM8S2hwsgQtKvFXFdLcWwzvKPKbsUKma6WHWR4/z1ehO0e4TyEEDZBAHrQ
lBekRsSlLkjTvkEIhcycoXMdhnAkgER4HY8MlOLLXVpJA8bxt4nnvgm8CRTp0bOh
WOfN2VVSWkS9M/TtKkKqBw==
`protect END_PROTECTED
