`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bgQqDDAqTL6O3WPGk+lZeY4U8jXnHRvYM2ZXApOGr+CeTZLul2DUb3ZV7MKqcxNj
/3xfGRz60km2YpVlvRbS5HkDJjkOlSKYWyt7eH14/RjRCU2sJhj2QgMWkSeD8Qdd
oG1AvwskNY3jynypGW2tsAbW0ACKHAjdgcTfebKECaD6Ke3+Y98JHD4AHPrJ0rjx
U/r7HWM5JLiKebL8JF9EyJhg+6tNQUcO18Ut8MpdzHvPD4p1yOdbMcHdcBIXxlXb
5mRI03bpivESflISqA/PVURCNICG9fKQ10Bm9kbbx7ElREHX9SnVe4qWUGa4eGv9
QV+UuKPHnzjSRD5oG7/c5aV4mw7szy23C7nGJsZGEqwUC1Aw+trZa5CZ27fJ3ODi
4C9316HYzLvssocnCRvcC92/LwPIfrrj270mZt0zI3OgV+3GK943x59qqEm3zSMp
eToMxRx159r+k7vub2FeIyvYJeVbPuVadhgmldHA7BZS98PkfDtIOj7hY5+lgzRU
L21k9/+smG4KVokQfSH1bO6mAK1RGgw5O6aYVudYWaiYJB93jfqag2OfmkD33ZeT
YOM3ohOO8XFubX8xvlRB0XA5qe5vcunNTomZUAF/urX+aa9T7vwWRyMVlG/pSsEU
wK3d8VoE7MjWj7GfCcFz0aa/2P5uxPT2kz3T5J2L9SEjrnN2+IoS5oSm4YwIjCCM
wbjVUyjh5/P/+OgN+s2wnSyoDVF9ST3QcIuNw/npXigAyw9wqeJNRsiaeWINZ16J
C38GfKdDvZhlM9fJ2P3lcUDSbdKuLZuku94496PFiCrRrDbvk5Ukur7b057jPi+g
8cAo/BgRF1UhQxyACILzuKGEIXRcaoSN3Fekq0xsqgfsTUgUQXx8E7bgcTUom5Uf
fiDlMa0AU2N3XxDXj0wmLsR0IFHVo/26AA9/aS4sxPdbRa/6jjZMHFKnwOTItR9S
BCfONKMeAwtkFInf9WlKZLqg8Gmj0h+KTC+enxkoEce7WC0OQUnYKRZPD44hTFJk
K9Ym9RGh/FBXjKS6Qw0zQa3XlmV7eK5lloozd8tBP7WGdB2tGCV98juZDch36DId
JPUhEH0VC/58x067L+J+bvFdFJbtmiBSAXGs7n/IzkXnhB4qZiB6aubhNSCHwQJk
pu/jd7lXDq7C0rJKNS82QZOfdLvEjQTlfyaWO2vA1nqc/UxSTLe5OJAQ3prxLWGH
xNjwJW+WYLIU0C0n0ic5IUBjg2/paYAj71OQi6/uN2zdbmEDteHkHyaalZwG69vr
gLl+flxIq3sXmd6lslZ2acBmSxzJuvoTXDqkgIIqdkwVbi/28N6qFQfmWn2nIdZd
mPHFfxViA1fACo9ZEgMtrADhN1hiEE5KZbdqugtX9FTUNXQLljOmd6KLFlQa17CD
kPT8QLJj+ASTKrOWOgDaEs9Tt9dGRYUOp++aIQZk9HQDszjuW+nxtfg/lbUQUFRt
GDbTWwAukAsyPVa4YAoV7XmZH5mZ8XBgAr00fsA93ogAJha1BbFoM9U8vDDd34rl
hBOEHPd/t0HP7eP+2wF3e3UnfPp5A6JEouGW3ok3I/6VzPmQcFfGyr/883FBcRoz
4unCEXFZgdlUpo/3fGTsmMzOG+sRLazV46qjWBvxFeNimOX0sQYhqRVRlD6nYoHJ
GzMV0bztMdpBEp3Eefg+Ay09nMHbVubEvtMqWbFnfK37aH8Sfs3q/jQ0gj53/qKl
VZifTmawmkCvgZbKr3N/uEARGTlc0/+Rj3WCJzVWp2xpRKyxHZIqiV7F6NFTHMjQ
ILNzqU355HApR26ZLzHqfTEbns2rqOEFRCrbo5Y7Gt3fF1rDGM55FQl113gJ/X3h
`protect END_PROTECTED
