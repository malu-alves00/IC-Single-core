`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
l9esXbhglzT57A+ak0ifxPrqslECXRMFrMUXyEPNBegAMdPAh8YbcOHRT8gywwhA
G9Ou7nHl3eNPe3+OT3TrRPx0dnaF0B7kCKLLfiao68DcnsWLjZzZjHVUARLYcaWN
gJXm7JB6fYxO9GUFumIScUqKrq6mQI7zDEur8dPYLrL5IMz+rT+jU021t3pzqGht
R02hJK10uWbpe8noCGGiyonBJep7YjLSNOSVPFGEgkr3XwvU4ltZ4bN1QCsN24Un
gYiCw5v21HiYxaXAw//LX0pQY2HNrja6mtJGryWZoG3eKRPa0KfoBeYXpqPhO8Fw
9IZhRunb6Ys6A4ua48Us/XTj2N+f4rKnpzIFpYPIDUY2YV22oERwNNfViJoPRcWc
R9MCqutiPvuw1w+jWDq6zMc4HD0KnzQFyQlSsYpcpssGm6uaxOqny6kVJaqP4vFD
PH6OWUCLpHibbCQlEwg1D4urCWbc6MnBEQEnPrKGjA/sIW2WwDP+vbMDVLldyhHR
y12DbCMMjv1/OQTabaV2YJcZSHrvoHFiNfvD1BxYVayD3agbs/ZhJP299s+/pDsc
q6LehALsmDq0vTaWAnRzIG8SyFQ6T80HHqh5Msqa2GgPoA2CJBn5xK3xzYBMJdAb
MWEtuPp4PzH6bzFyF+tPlHKUiqE0Y2BhkcjgqYo4dn7Ys2Ozq2RCz25sdqBj7O8L
6MuUGVYeY3DNN2vhb+U6EnetvyMsWjM17K/h0/ag39wG7G+4YQ7JtDLTV3TFpd6A
Cte3l7RVDzNUaFUyZ8NEF0khNxj4iAb5Jfc2nbUXaRS18G2OloNzw08mJ1GPg18V
UvnurFOGTIITvzXuQY3+uRnIXgXL25tb7Sg9NoCIVKU3vvtwbSNgpvWcwraVUXfG
LOT10dB35viguGGsOsxX0tIUuGzyg7tWvmLnT6g9xwBSRqPg5vG6uo/S9v2zeC7W
HY/6R/67KOLwOOboSzM9nLu5/uT69x7BFaJ64TP4TXM0U+wP/zksloCJPIXWPSwW
p2GCD5cnhN28KgvyBlV8D3fAB6uUpQgQ1GwFwG81BI3+1zvZwaQ3LFIIjlKKTBAt
fRp7rQRFXEt7xZv+0bJPThHWbP08hjYviPx8mkuOOCRdMpl/DMEeswEXye/2VVsz
sZ6plSRZPTdwKxCv7qXq5Q1nbl8JkrfpxodnRynpkVm7GFe2jkUORSRr+9Fv/dbb
9000fwLQZxBcLMaaNB7/ZGJbb2bD/8en+bG/l7U64jMu5otTr1xwK3TVeIl5vfH0
nEVGgLklOVzYWd8NkC7PG3RjgmUUEt5Klgvq3x1cjwS6N2Q6CiSuOlheoTKruTMN
JrfaRw9JdJJTKAF9RyXv41Va0tEVEr1AnkNGVysVSXzSIfbA0GbL3htiHbB9t7U+
TuQVl73vJzMBu6wkBKGzi5Jd6XxHT9HOOmhxiAJmAjvQrPJClvMwf8NnBebxhWq9
Y8+I9UDlXmIMVNjOVPlGo487Uzqsr7VV7YbDoYeoCMWKKBsBhAqffSuU06wJSEwi
h61xELPuAa0i2lRmJAw4VRnRA+CbUgIrsCwQEydERfZ1ZI9HPoo9GWj8txbthg3s
xX/0bB9Di6AGxDpjgoUUjitqCSREGTieALTvKwCNGiLJeyNwPAEJXhBK/JJ4RDPF
NAOpkOr1gkT+E7jurblHXBxVutIh988tTs/WYgljCuU2PLD0goQZHXmwFiEnZklL
k/rKeJGd3LBC8QfvNS5iVlP8z51lv8aNsD3lwMLWf9QGXgQyiF4piudTAnnZtsn2
4/RSF040aS8SbQjBByQ1nE3fqhmDmcgsm4VzwCB27CDmKWam4IJSy1TN4UpVKvr6
PyP9uHxaplUfo6h654aI8KTL+PO9rURpd2GXfff5iF4NAs677kHpeSpUwi+yVPcG
GXrVp+Nuf3vvnO+l5pi49FG4Z7IDqPtVWPJI8wcxrmvOPPidQwT7KHXFcyTAY/id
+dIY1TvnWFLtONxUCHVn9jcwy/xAtOLIV3Ugr9qmAEqtZj+Zw1Ou8CNymX2Ej8kJ
fN+mcUodXhk/c/NrkEYt+KMcZbLXFZZSfRzU2FWUNCr0aQU6YLh7b1aQ4fU9eA/T
Mt0lfIwRpCVbkfqXFmcaJ1cMTj33zhvnaPo4GUURV7C6ipWVCWie6DTv5JTDxvJA
WgOogPVnivecbJVn+Roe1ZHf8xhlgrZGKDTGVp6iGd33qgS3GCK285Thc5AZTzsY
YTMHcaEW6Czaojcv1cbrs/VWOr3O3zjAfJJUg1TECWyVG5I39tn3C2AU+NC76Xns
cGdJjcJq//h8Z70HCSzt2KT4anUMpaoa5IGb80PUrnUB2oqGN0hlTXxqoR4XBs28
nnAO8cNMALN9mDBcy9mP0EIeVrGW1gL0/ViPtH33r/YI4GWQEJIFepTKV3AUm2j5
eNABT6//tboBSZxKpYp/vS8bT5KRl61tu/hpmRjmQ2mlxOfdwXav8zwHOeXfGkoY
x3KYL9JNffA8qGqRcdmcNbkW10WS6iiDAiMT95qS6G4itDti5rKJ9L3IU07kz7fY
xorGTNlmADCNCY0cIdn2W9aP75Zt3cXGJJCfWoS0trQ1upLnj8iHpNs2mmoFNJGJ
WSMRBFZ6bFuiqWyNbcaqfRp3HKE5uEq2i47jOa6lzaExnzsOu9TGv0kT8hbWG/Zm
urg0mATNGPD1Ro4kRZ/Je7lYrPyZQm2lzdPfTpIJnY1hRA9hr5hAXkc12NcQ/1wc
N4SNl6sAGV+KecAj5cYQAGTF2ZH0ZUUeW7nUMNDw0QGNXDUObuW4TnADljsAgt6u
E1EWI+/0bz2AtPScZv5Kb5ckqc8MdG+nZxeqWO94f4Klnn9Hj+sVYWjI5PdarO9Z
1QoHGpOivvuMq/XUsU5+qOKxarzZg7CvOlicJUEMbj/xOKrPiY+ShWBDX6dzqRvR
4vpilXzp68uswZgIBKPQkULpJXgFA6HDZYjRKZ6B0Tm89FCBVHogkQFoQZvbhipX
kMaLSI2xJ++9JINt9QdGI1x6sNODUEVNrgtUgo3Gwv9JGFFxG258X7SCR28PYMlh
UcxNyf1v06ckWeML55zUfF6XrQ8tTio7dsplFGMKj1fM2Aj/TY9B55AUM4xwDWrX
JenHXgAeigKbHBogvenevhQf0Ew3xA3+idOZiz6rmJjRK0S2WW81Xdoa816j2c9E
DZv7VSYBn4eYBV4l+cj/S2fURuSSJu8gho7LFvUSqQ6p0OMC+o3UZvkRXo2G0O6X
rMB1ik8z44cOqWQjBajpHih938TEdvRloSPd7XAQPf+3C4l6HU5PKb+TbvVos8Sp
HvbEncmecDhH7lGjU5CRbJ+Z41C3X4CSostlS3UwokvE8KaysL5xUW5Y+FW97mtC
s2UGS9gUrbxMYWHLbDMjUkWx+/GMFiBwjXypi76txyZbIGFAQDrGDhecVxQj7qoN
3VucIBj20t8zjf69OLIB2b1I8HWXx0CgARfzCJxYSQpxifTt4hZRZl+R7Sk2GiR0
pCtwU5e/HplQ3FhkWLEFh2HrVrL7WSjexg8MRU2Bx3gPvsGxfED2i0AzCi9MR7kZ
e6dFg5SWiFBTVD/prwjC9CRpasZ2lYVp2XmsGFWifAXs0W1Uc67sSL10Fyu9f4kP
zTWtNukX5y34LWDtCx5z464+U0Wzu/gcIRvCMBkVoq/Ls5/qu4maX4ysX3tU+8Bg
T0+L5UsuKs6m8ei28A6nv98LgcOcJHpdOOETnqEwA8V97HlxsNx/lX4LdXaxafvR
CoDTZmzFKeR0FDWNF7VXTIjxOfxedINEfK2ebGqRm0dE8PeVCfiJofn/8zhfVM9Y
ucpJZu93jdF5e1dLY0fTiCIk51hXS7gSYO+koCeyhKjpLSDexnmL0EU+OAyGZS55
iq/MbfUDZnY+PCWd+3Y360ZrKySFhPxFh0vh37LRen81dUWvmu3F869QzuF5hSJ8
kcQhpfUyrTEwcb15016EJuOY/seSb0rW4jWCdGaK8x+aYwKCb77ghZsd83p9jXPp
ttL0y4i5Uhry1cFGPQ6/NxufP869663QDaCWY+YdO9Pio40cIGy1mE/kJ7cKW3Rj
P26FXCYuLgFCDO1B3Ft+Mry34kye/DNOKuXXY1nCOuRJdVcwrXSl8i7bqVzLs9es
/Aob/9GKcxxJjzRmntDnny5dnBMXgmWYvNwOmLp4IZ/tz9lC5VN/w0uY3CAYKUVW
KIm9FsLGNLlMmGJfBaz9D+iYnH5/P56ZXub+MCRmaMS32NEqG9EZ6+to8FcdwK9J
DOAjlOPDS3hczwBeDmuwZDMkVVTJ3IbHpTwrdZsspNdq4Vo9HtBUKre8isw7rWl1
P0t1VLNgIgMdpbvtgxTsJoLhZnYC/v2wU4DNdTCZ7xeXAhg78hIPNvC9pclop1yH
sKUQSrRtI6TwjZQBYx1B7P1Duo0kEVgC4/06+JsXOmQDHuxsEYUlNJyPcst7C0h+
JyLqiQzLZ/CEjyhQvD7NUNFjKZ9IobLU+fm+QvdsA2sM9Ryrt/4ywyKMDsV9q1sa
BxQUaYsvrGP0Z0ydC7oPnXB7H+J1cObp5tIMQ9r9TVg7a2wKhM9g+Zxu5sSpKJJD
Gj7KVqdcAiJ5Bj6EjsoEBoLPd9P8tlqHsHpLZbfkch6DKciNWiCyPbUqmWyCpr6N
iZ6rfNDd+buDPiENIsfjG4qkurXCCtq9fnj3f1TGRfOLX6VnizqYHPl1jzXvgfHa
KBK4EOjqkqQSKkpGEC2Fxks9e3guLEWNhk2QsJO44stbVRl9pkAUTky1mUkPeoS6
xD5Y+vl4XewYCf9gI5kZ+tg89T1uo1cDizfz/9V5m/g+lulC0idy65C9vU4LRut9
jqDKJpC0iFrY+s6YOVgYjmgTNaUcRoysJI+lfIXr43PnJUf6AwMHFPLqfZP1dY8e
LS5FrnPkK5Gpg7t6rbjroDE5EgZ1fkcI9V3NPt3h1OBeVU+Mz4TgN47U0p2djkKd
ZVF8/TLi6ohszv4rFdOUj+rz1L97Oy4EXkWtOkin8OjCN5qdwBDqS0g/aSHkH4g5
Sws2zH6R+kI9L+iYNI5EJA==
`protect END_PROTECTED
