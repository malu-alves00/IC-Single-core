`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QDc89Omc53ZuM6sl9I5iSym6YgNcmxiLHRJJ41HL2TRJS3JcAdG64nhUKnGKl+B9
0gcda/YAo1CbrPiME8j+wllHC7zJJsRDrL4t8p4MSTtQjlduBdYRf0Cwj38UAxkt
whJ6SGjKOp9s4reJp00epBEUxOhGyjuz1ImZl+wlWJTX45jdAIOXI/kHIgdT/WtC
uVcZe3EkVEs7RAqSQANuI8G3ljV0NBWaIqFRxAVA55rEkvJd1VVH8uLiMFcg8Zrc
APD/TZeW5WVeF783co6WemUrUR+Mb3C5qZ7xr7E9qktCNSwhtIRnNDeBBWkK0vbP
dwPfK1ZDcegdjiZaBxQucYZqqOKfNmsBteIN/yx6CTeVO17gwpS0SjxBOwixVzdh
nE/zAnNnq0DnthQeleoOV548OLSpy3ufqVVeB06z0QAttuMceisHM5oodfIwpWQ2
WdV1HMIQI4j4t33yyej9lwtpv4ZQk9a0mVz/slAg302jujMnKtMYZNsF4lVy9rKO
h/cg4DL/r6IqMZs1DcYkvk54R96UXYGXMvCHC9GJyf2el0hrSufpZM/HOIZSEIYs
/X1MsKv9x0hfywbh/TaEv56+Ad3WJtqDJEz8NGLmyGyC02AFS+aUzstNsXuhhTDo
QY8UPRBJA10zhlivYe5KRAODfwsmOZuxOC8VPQzF6U6gDOjpp4ZCq0YNKO5Jrx79
n1VcsCY1Xao7LxhLVOYohLcDJmizkt3pyMmq24zR1PmarhjPZrAs2Ybt6BqTPFw0
3/gDfAuCNbQKyZ1q25NjIcCIHPNP2DQUgDDOwNARcjH/C9q9E6nTtIWNMSSBuvXt
KY5o1gkTx/4Oad65tKZFHI+nzbjAkWCRDyXxXj2Onw39HACjs425pNeoWOQ7jKrf
MbjutOAyp3FqmTfmGYbVYSik1YzaR3Azkxv16QjQ4WeImRsRB564aijvM5odiWzk
jmgn7+hinK9ALdJyzJ+zD69L6T5ILOFrFGHLjkBF7XUkJf7uqQFBiBgPa1k+ApDY
UbasuXi+S/9IAWiff8zEYs7xgpORb2OTawRQucpvPcbshtutaXDLLKf4rJ/vO2hj
diGQvPhpKhxCIQBapp6Un+B3kfXX5uysQlsQ8wdPOao5VCCilzDszPJpqAPvuFPU
BT0Zzez/RgpbGhNpfpknHvzG40P/DyKPlU3gMbRsvfGPtGdct5h6PS6l+GuteZRD
l8oKBq1h+6jr0DEewEKs0Mr48H60jffg1glRjtRVBjNHMEkKyh16juampTf+KBX3
LNwuXhignl8v/fSHKQFQnTAthLeQRk7qc391kawyAhiz26zPQ9Kr1jJNdW/Fjdo5
A2i5rd7iCDOQqxGhV15U5JER1cWoYRReMHMsS+nTkelsOoFGsFkDQw8ftlcVtB9v
4PhzDbxAJBqysa2PZnUCZ88bwhzkDsHAIarx5PU8hwFWrZWGARK//TpO0Wy8WHiN
`protect END_PROTECTED
