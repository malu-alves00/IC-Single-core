`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
T3vSTzeYghTwRQKsXsfEKW/WAUmApZkZkl8ZiGfi4LN5ea/+FJCqmrbe6GLgVhIY
CGTBwzE66ZNqsO6QFUlk2H3R57zfLk98keDNnQwpGOXPzD/rxvBXlByxA4yHlfSD
4sOxdpRV0DoyhlWJ40d3JwyrFeMkbk4fcjl0RI4iFT3aJKnh8bXv8bHNc9uDLXNz
6NpkHgrUkQiIB2xW3JGAQBbnxdXUExVXHkksPQ7C+5s6h3ChC2UxhrNbqJqcFXNi
5PW4SEl5H6lnJlDbCLiJayRFh2OBIku8EbUAXyoYNirBZem6I2yEReIe+V2Jy2md
OSDYuousOir27WRKi3kdxeTNmF4BAG8YXqjM8stj0EDEoegEjzR1txA6BDmAmv+s
pWYnqTlghzi51JVcZh3f8TB2hrIU/E6RVkQ0NqJ/JIIcjGQKHzP/3IQ0fPjsA+Ni
v3e9CHOmiQ0rjxjrkEIlcjZk/ZA7pvSRxG4C4D/qJIsqYCBajcqS4A61MzL4x70D
MWu6Fth6uUnplYOUivlol1/ZqFuImZqKxCyAmeMxGyMrVOYlBU4o9EqJonn1bgWk
N0NU5zwRpoGiaUWqeGodUisayAPyWNPaUI2InNxqk3+esNlWGTqXc7YfwxX9eyjd
pzxP6YdNSDd9QgCYCflmOEk92ZMqkU7d/49xuJPQA6+BQiLQNOD/JxgrICOzPi26
TQTGjx+ijYPoZdXsuLSppFA1REMyGD7Z+K1fa84+89jWivdhL6AnSdtTNxg4/DPZ
BTJB6dpPq6EvT8OZXP1W3Eae0H5t6KInWvRapMV2xuBtb3MAwAaTKG3lgwENrGwN
cLtKhcs0AO79XpniohdmwAlZApMlemT7ttbn+gtwagwqshloIsWXzVqLfKQ+dMtu
O6jnp9pCCKACwvo1naKmQsFwXDYnUDdMsN0EXlgxkP51Lemxon7Xm5iL9o6ZxyRx
dxWoKEi6QvGH0h9RfYyj2KuWGfMXxhardsSpAzwmx9A7J2I8bTcZLHAs2meOuBfF
nGIRxgC/DL3rwgysNF2YVMtAjucx70/ImW5wqQIFFbkl+cnsEzBI9utNGs5w0MHm
OQ7DErjilwSf+HPnrTqt5H1hp1ndG5uAnCRNYbHEzw8wHVCFujhUXFGkUHGfpOfV
+VGqTJ8/8SCFT+2HciwrPGZpgPScCjqN94U8eE5ZuOVcdh5N43kB/n3axDfk44WD
`protect END_PROTECTED
