`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jLwUIE0IgonSSHpPCI7wzZAOiF6aBJ08YKjx4Zdb+kupUluDXpkb8qg3M34o+qvc
FDAMvwA7GyqRUSK6fm4VTHg8p6xmDnoGnvpzxZ2LstLqUsGZZ3PMDK5u4iEhL4t2
398GiL2sEycGm3Ul6mnJhj7le5KV7/FiX/f9QU854unW1egL96AA6blLENnnSOQY
B6ryizksiXEHagPwE8iZMc/otyVknpf41fQF4ZHs01LtfB95fxSFUar9w3GeTeo0
KqUmcjZ/e6TpFtHPMlFySMzFrbjN7a1uFAmkj1Wue9gdpmURjOY1vSbv440F5DKW
tZIFfGHjOiJGZ4JdufLRcbA0tP7FNl5OOudx8Y7AjCVt/2t3fz5YmlxSTe7L6qsj
n5Mkas8XYe65rQkkcn0soFBeYCCP4qe3n/GRte6L6HLSaj8h4C6ftzHbrl4Vsmzh
kNG+X3+gGzk8DRAJ9qa1RQ==
`protect END_PROTECTED
