`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AuMiw22OBKmbxbxvqxhuJmgZfrSVnnbv/vfuo7FdgvuIeg4BFkgbyowKadsrfTnx
VOnnIirdFCjtLQoUdt4MOgdFAT8cvjeWdSXzKaiZy/7nUEEriglws0bcCdaOrUrR
hV/Q9def4wUR2GLEH3ObSKnWiDAT5giYgvDlYTvL1298OQncliTgIgl+eWS5kIHb
vh449jshHO6bDCB+KlWOVUCOF+QdGrDcPp6ERQvn1/hCTK9VQhseJ0fK1/Q3ZHqw
fexzLtxnGj1u52snOQQVAmDXAAfDF1LxismjX2NjMZyYtIKQniZryoTRetLBCuuH
K7gKDUI+NjHFypdKhNF8UW4NqWheizIf0uPZIMMDg0KLmOTV1wqk4ATHP5XwWa+U
wuHCgZIaDDI66baJvp77zC7x1RNsa3Jqw3dYEP20K4O1RuCVJbApx9fYMk/aN60m
FIWqXFvusjRJF2UPT0+g6lKIZcWBUFv2BL6M9gtlEYnI+cmOodW+8WH8amifImRV
bnK/HC8DxCCD1gCBHv3z3j752EF4z+dm6R4g/DkNZbP2oKa4pjn7JXXWmXEAWdp6
bjiV5DZwR0GLs7yamHIL22ibeN14PoBovnFsg0Kdo8UAFnSxuOR8uo/e4WWIwpgN
vxjIVeoF9+AuL4BiMUof0g1iO+nV5/Cm0eac62H92wx+5xaKGFWctvv92YSN+SWU
TN7ji19kPB2VZ2mYxyEx5IsmNVNRXJ4tqJzZ4nAg2i/Ip/ZHiEPSbJSQYbfJzRkr
13J5DGAF8aTR22YD0jy0ScEFU2FJXiNPRnQ7Qd+rEebzdcqlzXyb4xtBJpVWgbys
JjgivZLowHiVCLy31n8gCNo6iDqdyy6K54KeBcY0M99HIyYUUpCyp1q1xeEu0snY
GgJAiG9cg9wyM1hfxafx/HdaqN3LA9uFInbgNqeL3erFmUFAGcZJvsczIWHBv6cg
YKNSsmUZJQZx5RcrMet7kzYT/fPg92zQR9emlrDZkmB9iUfF8H6/9w+8aetfEMvn
xqwbWjF3YZFrviIOCx4+3si1Sva7eVUOF9sDoTBVXRPre3/6JFk55V5qgyD+L+T0
vyoV35cfTLE/UUPisTrUpnD8WRj8mkx0/sU7wpcPfT8zmhw04c2Bz30Cc8klP6p2
RIwN7k4sOKYtfl3BWOXyC4mNjZVUp5r3MrRianfCQTxwjrruTSrebjwLEUbst4Kh
BDH5Mw9556hDLtRubRdYelIy3L4gYXqL0F0j5aku4A7FSHHqJSZk0qgkGeWkAfL/
iMeDfMm9XEi4WlWQeU+nJz9lRoFVT5JRpWGuoiUnXoqr+sZOO+LcWt7D2Zkvpg7z
KZdT3P+tDfwG5v8nxOg606K1SJMjrFaSeYOlAMQUQeRadR7Bz9A6hlnlYhGUtiJl
H0Cho1AHQZvCQ3gWdeej/YHJDZseIw6x9F4wlm+KJ37bYgbKEb/skcFRBCd75Mfz
C9+GebRUVnjNFqGNcQca6JfJ/euZxx2rr+/2K55+qj9qQ+mXVs7MP0d9etX6ilcQ
vLw/o6v47p/4e7fote+Y+P/Fwkddg5Lkp8T+Txmnh8vlpwA5EcPQO+H55q+OJ16n
LgYYXUHLRZ/aL7eP6rfaMYkPl58+DW8e9/htJDJktP13U6jf3MEIhtdWGLdY1ZNz
jyIiFK49mKTvfHapqqxVO9UYmXgcLz2BT2lryC/UWFbmm2VV4lF1sTusScobUa88
EgLORWkR+23PNzvnGm/cYD962cqB3NEbb1iOPg+z/YZluSQfCuDGDry1BE1gYWFY
Mwadt/rO69AhjLv6IApiL0oq/2Hkx4Jme5becHis/GB5Q+rQLEKOpbPAO0v653Wj
+MeQnGOgbLr0zSXGlXeD4DBhZ7T8OytA42kvqs2VXruD8LhzkRIkYIUBMpCg8CTF
Fuoes8FKkuINY5m6bL/N9eJcfYwl3gxS2rNR9E9ZIKaZzXrLcuC6Z7W/1FOs40NR
U3qkyXgDNk92DbAbHP52f08mfH+/x8Tvdgxp/rrHYkgde8JnJWLm3OWQx8mH8+Pg
iD/mKzbphU1Y7bUzIdRc4n3/ZaX1C6jQpG4yG2OSME/uwpBvqvpQIVdK1EV2Exvx
PlBPxBc0zA5oEXIzowMTKNxVixi08M9oE5f2/LmDK78t+f9AIRE85m7WGHYzvg3j
GwvDI0VF/pnfPMbh2Pj7VZqs9hmC+VmUckJhX6xD5b7SHPR2HG8I4XybmkLhXSP/
4ZFEJcX+8+PDVfX49bfoyybzOUjGIgCCwur1RtMuGq7kcJjC/aXbvOfwnQJ3P5Wv
4T5OucHR5vShP2qbtoI9Y7YwGAOlmfZz9ZxGi6nIaD12OMtEkLMzavFCzd2ohIee
bxx6htD3dzlOlgKqGBWb8sh09vMYBT5qFkd8XEdxuCQtaZnB/GJu8r4/kRu+WE1o
DVYoqUEx3C9hFjPteM80UVFP7Ne0eq9ZOFNP4RAEQeuUWVo6zAt1U8q4ZDaKG7XG
Qx5R+RVWcM4K3y5tYpWDcwnN8CVrzN/wzy9sHPFQNPKRn8TcuUZdWaUQwTGw6n+1
jScNUXGK1gSJp1Lg+YJI9zkMK1+4i+ECPpfav12TadAk+pdRYWG/wl0hNISZYgjL
yR/Ujk8MwXdYqVXrBRX3I0og/I3sHuhlMESzLNgy4YSkpIGGUCuwpCSQioeNrqjH
wSei0pJoJrJ0sno8sOPOUUq2ZHwF1Q/ImF39chlKZO072x+/5fMBEHdw/ERK0xgc
jtIHBHSOZKugXcdIF2fOuFz6gQ+74uyvMRIB/TUZse1n0+EDKuupeEPqMTcP8Y4h
H1benfwflbqMQFhZrsfjSfsk6g0cBIGEM37+zl5bzhiMaV1WWIOYR98/AVAILgE8
se9AnoRQyt6++qxlEXMbOeKCm5rHW3lewew2UcjI3//1c0k5ODqWxtacOGY1bk1C
y7olIX7QZYgNMUez+AGZPT+6z/EoiKLsiVfEbeKZC4x7niWGLHIyhu0xAsbBZj+W
KQMTTiy1Xixh6uzbQxtG/IJCEIK7HT/7uCetU4YgkYR5WCzVJUykhOEwPSeaBdD1
cQ7nQ5PByUSX1FRldKhBycYBe29Pe54ukkj+61oVIbOJN9cyEdc1dt2mL6Fd4uod
a6gP5l13adohOmvjzdFLiqimt71Q1LUQJxVj8TEAemquIjNVe2FOTEq8Lj6/kcvZ
XSHekd2QnNtJc88dSO5rXwhnVWc+CRur8G57Ll63R89kRuzXCQZu7pR42G4VEgg2
n1ggoYUrWhBp7EGytHU8eSm1lV5O4N1zQIB4U6XQOMDXb2hjGYpCGl4RI00k5fxb
nCxqFgpECs2v8ndMtPirmhibPRkL11QYCniHs03J2BAusUQYnVkfh9wVLArIlPjZ
AdQuDD66W3PyfdKa/6Ku7aLzDu9jMrb+y/0ysukLLocIM9N70ZXHU6FgbFSEoeky
ZC89OFzHHfPAEWxVmULpVFV2Xbk2wP4PTlaZdhUvrkpIBbGWZbyN6+0jfz3mhYN/
Q6FjG6wJ1k0ZCyhUk6nu2vHd07ApX5gN+viLGjc/hVTfuypU3YhVzpNTyUN0PANz
1Cz97HHgL5JNMtNm645k03M5ogmx/uvISjwcsZR4wuVODD8cu1DveE/FrgyHms9X
xQJ3UHwqznCAj2QAHmecvApeLRrxUG71xYoVxuQP6rAArjrDJ3omuodT/PQCLi+9
FQTb3p+nA9Z8wicMjC+wJK1kMeHFcddHBzNXp4N14SC2BaqCLxpMJEYYT6gwswzj
3SHNkWTnDEhlGNPRdff6eaH1qWQCGMSl1vsA00sDPYWzc6yR/TvmgZhd07xPFWsh
rMFjDU1nCOMPhGjHThInWQ40J+e/Ty43S6ukLCtGO53FhJKkmCC72vcgOYHXG1G6
JZ/hP12qCKj0E8wlKRTApzBdo6qushJE24qcLj+DEd45BdFFL+44gInNSoBj3wyQ
FNuUG4F66IxlSLmsCC/OfyFIh2MmspK8OHEVERJ6ENzQ6lRhsXRiznxmXoxIBwMq
Z/CEFTG4PIP2+jsoIr6GaIIuy3475WnBWhlhjM6uxI0Sre0l0CNLKXGvbRZJAyCX
SOCzPykZxU6wvzl4wFWT7UKJMzGWpcKbzzIk8ZtcT9kcVKIH/oSRpPu3V3IKIg11
/2+26dGlPj5yukLMNLc8Wy7vNQAvvKnsSM1JsRvWSmjbduGmxYO6VsvTbDvMJ91G
zNYm+glXi21pBFlruSzeWRLVN60aQbFNR+Qwa+sXLyLK3ssD/qx6pzr0HGVIiX/F
hkpU9lvZSgLKWCa2tO1/F7zW6mQ7ACf4DTlLhwDuhVlK6Lut77DoDIe8FRPviAoJ
v23I1cHu+UVSMBW4yFhPkg32+kBGIORPL/fW+kR9kzktDbojFUEI0tu+wJWf9y9T
Nc7YzM5BIn0Q5YJ5iHQEgpzkCSylRX3ZJ8nc6HzDI0CzVOUbtkIRu9DeI4oOfUEu
YQFPQ1lmXOKSJnLiMtKwyd3u//oTjPlIe7AerZYCl+tR/tNomHoSWb/r+PhmvEoY
KFPEZYRHBDM5GhPcTi+csnlz6kUfcroo2b4hT7o+m9dPZiOiJvRxBKjo8Uzhllpx
dspxyuCONEH70b9ji7HaZ+DSV0+TvkLum+II2xoGPvxr6kc0m1qOBisAr1V/5B2S
u0kD2ihCjqZbPhxE2nHRtcrxrSeA1S6Y83v0mHzc9jNuP+KL/HNiS+CJtXjkmKcX
fulOMOwZCl9gQjmMGPWa3dMSuCjL21h3XOcZhCoGx3yGhrMhjanml0tGC30Yo+Ft
amt8zcswX4tHxYaroA88FlRUo79Lnj4HCyNYc1tm9JTdZmCS6yOahO3ExeH3sVBr
QHsHG3p1Q+7Ip2I5e01G803vkEmS5lna5XTFXztWbz0ZP/wPszf1In2iDIU4Eire
XHmgPQ+23pevrI0xuqs21PHcHi5acdBGCNbq3sC8Htkftq6kr0/GEhsibbCmwcq9
Bu+Sn3uIFr72snIBOPSZ31yHofhEenKoVXev07OvZA1rtFxxYYms5RwynuiT01uC
FhgEPSqdr/0TaDv3+6EdMyqOh6iaFpriNN/wQkRXEdDH10W7gM6pGCEpU/9ANbxj
lPonZ7+gZdUOY7Ih0P1avh045oZiY71gDragjaB+rDPjnHpwxT4Po+rQ9FP8DTSw
2qwJJf5TXOfZjkp7BcIt4tbAKdhLx5JNry4W9qU+Nr184Jyx+0G4MY0Oa6DWe0nS
IX7xDUTPR6XCobCmMBYXOk+BAbexEqghbjwGfSl8qbs7PRTLuKoOkIwvUwfWKBed
OKIjYZfQ4BnJMil6jieNsFxWXMdOAR0yIDHARRA/tMcOH15zzbAsoFdp333u0wEE
PcGclf/RaW45/tOEJ2AgDf6zgv6zc+1xtk2XfbFH7/MaGEhScigGd7FJgGbqhcvL
VS8FTQ6Lem8SWRcCB8j8cYQu9Q4rUKafcIFnVq6zrS/tVbW8mSFiLkdip4YiIXX3
SiqvtFsWUNnJEzjqB+T9BFS2BNpFJc13HawCCp52ZQ6MEMXbduia/hBkgLdZK6d2
clw/wDgrFb3KMc8JeJB/lFcrBXgKHMvVLzpo1dsWf6Rdrn8BugFEmrCd5pKdiWQ8
La/PB/xOT75cpwG2uut3Sc/qlwfQCf2NRf7wHEovI0zZRE0wfx2kRCZVTmz1x9zF
YBVPb3p1SDNRA1eWKHu72x+F+Cyn79MPbhDyWAXHE882DuPpAmo+xg8oweuFbOHJ
V2a1PKbk/4bKQ9MUi4HP/cTfUvwD2DBduLdZ3dlYzN+eKDqPfH2XH2X7GvvyEwf2
MsSIxn7F3hXmxDXBE+ZqnSPFihU5BAvbSoVYrVsZ+FuASAho59M9x7/S24pn60ha
Ub0NeJclBOCn6CWPW0+4fSJYbhNM1Ei8zBex/vZw8F8lQ3wqa5imadNc8e3vZ3C7
1VEDvQXbJAxP8typTAzbbSI2zyls+W+xUL5SE69pynYOaNy7U8B7xc6/QDTgEGVf
+D8a+g95f4J1k4boyDuBCvofYALgOUr2L+FuNMavkn72nJBWueSLtlvFqT3vqaUY
cWrWRmjaVAqFbP0UVEhKjK1IsrTrVLyOMZiarNffPfHTFLy49ekLDBYMbD4WAUX0
nlQ7JjdbdDa7UNjOpEAxFvc39Du0OI3JTOCFZVO5KCEVcizceGUarOFTr25HcsIM
Cb76AmVp5zCUBUNlRUvaVh8qGmAO/bkofCY9PfDtp3e70NlQrixdCKhK01p49rzb
xW83zSYecqBhdzHuKRz+bpFCtSBB+JnUgLegoA6chMTdONPONKV06cTF6spuEx6o
5kPdW2NHl9VRwlO+RuQZawXcdacWvlXxP25UkdV+Fiv5LmDjfaitb5ETHVpJwTu0
d6CSf58DiC35DvTPdYhxQDNShh4MFvp0gSimQD9EBkMykAe8HWgQwOwmTIcZfsgm
jYt0wxTSaglCTtwna6fZFlIOYbBv826DmkI+gQCTSkVDcC5BuMUJkdz9sNEfTV8K
ZSXYxYyyvahtRECQLyegSlWbg2fnahvzO4PU/weZEBZIBILLyUXzp7dKBMQhWxQH
HtQ4yugnbmzEOFBk6wIp+8Jn5ncb6aIWYdHfpAoEF6g5ytyr7/nXbBFvPoLfV8KF
iW8qIR+gt4fW236RNNnULsnmHjJ30or6UfKJ1p8qC9DK6fnrIH/KmtkEhaKb5g4E
1+aiwM08NIDW7xaGj7EtD6cwK9sIhWp+iUjHkPf0jHghZ0/yLztO+xr27yXddk/o
/0Nbft30cXwhfTYq5jYANPyS/FieGMEX9qaRLtWH9UxxZfFeHb7tkiwQhMfeeiP3
k3nwaX6/U4wQQ2m6aYlVfqxwz92aVb6Hpa9bK+lSJYZYuU+n/UBjRAP8l194NLqs
hyrT/CijIjqvVMC2trrdOq6OzoVETvDhv+f3JFs0UKXxpSKU+OPZr0PlXUYatPyc
FYckrgi3fxpHaE9EACR0IMgaOgxmOZOxJr5VTlZy8XGD9+N9STI6SxMku05GOE4t
IefSaj6nG2jc4qdS10pzLWF0hv9iTwulkHhMSSP4kVMAoM5OHIpPNUqEGTXOk0M8
6xqoGuJZP9miyVFXiFxY9+uGFrvy0S4062bBWRjn4kvxHoQMi60+wX+vLImmGSkc
EQl0liL9dOSwDMdfSeM3eciyq+yvDTfagNKKNixGlHHxoLaPx1PFHVun7Go1La9h
dV31DkFCiG4OCjP4cC3ksUZs4GZWseaBmjCB851DlO+ikQUyYbU/mHCfhD4hqfB6
Rrj2LE+XoDXuObjKhWiQTPg8c4AgP7+ZV/QYf8ubPg0GPz2abovyoOI7/X93vZ1v
TB2OknB1BwrmJC6PppQNFGftgUZz1Pu52h3Wex5netpAOx2S+aLdZHBepX86DbwP
6f3wI5Ar5JO4t/pH79zPOrp2n+LBCL5ehS2wtYs230/GFqxd8XJNGI9mGwPEvkFn
ZC+WOG1qXZEIYFAQBZ2DxtgRh6bpgxJbZNWT6mf8m/vsba7sxq3DSdhdMH/maHuU
e2XtMtW0mieKDV6yuq6v7te8+LBXUY+vH8SPz7WELMHM0Sp07gB2+T3EcpsXMhZT
NI/kgdKwH0f4uVrdY0nNGgDSS5mBXl2Gzjf30Cu5Lx2inap+dZUczTjjvcQt5zkV
jMgtNbVzpQu8+YXLbReic0gXmL1C7alG65Tv8i1DFGfws03LuyCsEKB7X/EAK1GW
5nhzhEzftEn+xqicxmaEdo8B8YAbEB631+llURDKx36ySk8cEa57r77X8xOEHaln
UrKOjsLQjPdUA8vc/7wwoBjcZZ6WoAr13vEd/JBp+DM=
`protect END_PROTECTED
