`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
r9xXvEnmjtWczKLZtRJSd8QnsLfGydFtLkP9fFDAM3pSkvRfUjPNQDCKk0939ikE
h1pvCEuS0iiJmoQGVr9/H3PxHkjpuf9isgbWasXweknpg6CYv/+d01T1sCujMC3F
jwdOa9RUTqzDUitFXiCoKkhjnIu1zmOOxc+5tssRISwoisSv4cF1j2h06acXiyEF
4d/clZR7AyGjw6AuxX3xBmSFKKDSo0hpsavUhGohfV2moSEZoht808CypD77ZvdR
J+4JWMSnNKino60GP0r7IajH8tD/Z3Wcl8telDVxIlu4ruLS1yMl0UeBSpneXCc+
TEhLKL5yOsNpW9pME15FnUMoSLfUZN7FI6B6uOczD29cVstJ63PO4w6y5tFS5jHg
z3LWUBHv7sYHTA4MWmSZOiwkIOwzFXx70Zc23x0Bs8kJTPFPs29UJi8Bpb7wxa4D
1PZ+YpmNfVWMChJAP9wn+0CMzjhv7O3GrrEvw1UOC8GhPNrojLe7oq+5Gld/41sd
cu7ZO12RKdbaK7okYSVI+e4s2FP8eTLmuKL8h32z27BAvgENNq3K+bkzzFF+E3C7
ZXwrIDybvdsT93rBZAqdFfV6HhJI7biFwdUjq8B6pA0ZcnfvZf2ElDbNX62p77wq
7gt2Wy5zSK5j4UiaG6uLKaA7vA7+iTAbsO1586wkmMVX302JeH23//h6h/J30Xn8
wtYN+3ZhHWgsqFqgzlC/ZEhM8EQTNe/5epZgKD50SAxj6QPjuhCEN1JSwuJGRX/h
UdsaPUIFdPTIUpYaStZnw5Uz6oAbzjjSLHjTLnLZKFA5AZLb589mEJDq3D/mn1Go
ViIGAS+5sy7coxKZecJ8ljwn6WlehKRJPN0ReNdjTwHlkxPyF1jYXsYk46sMTW2c
rn/qEgHoKZDrSgHDUXTCr+zDxy0G3lKdvreRRPHaTzeEieQaoNFeWoA0gGgKYDFH
fAuCjDo7Mc3G8AYQvV71/Eg3SavggZv5zzSyyMffWW3zFQVFO65afmdxmqtqFj3y
tdqz0BZYOC1ijOzemswH0L4fuu/+tmMTctzeVrnc4FtVM9O4CfW7cMcgV2xtYZTD
XQLHO2w/0YRKGM7hGQPZoFhZbyOt3vWOLXiyxG7jA4pcchajMCqqX+N6HRvDdMQp
FfNvX6oTfvfmLgtmp/vrjGXN7kz9n62qSsexcEJbMzyoi1sV+ilLZenJx/kJHGi0
O70TgacSaue6BDHDpieVUIRPThuqBPd6vey8GMIZNce0ckc+VgJffowdC2jpSl4r
5N5GdMwtOSM6oS8XDQTs3X6HLnws+h8iMMCMEgT+cWzcwap9tw1P0qoLGtlFbUqY
nltmfeoFD2mPYGM1NV5lIti/a7fBjH21FgeDwuB+utE7m+PK+7uDHBOAbxKkeWJp
1I5DWK9eaqPynu1tSOhn+LBaB00RIe4BBfQ4Jj/ZYD5TvhfyA8m/Jllpng9N6t3H
I3HgryotQrbq+QiwrNqMjmZZbShO4CKPccnn3UfS6t0ffYjELMSd9UHQURHN7UAL
95jyedUkCFwqmYVNjBIl/4vaWlCkOX/vCr4T9EGFqFRYGi9Ba5DOa/2+YyiN7QYk
fgHu5le0oYt5/nYGHp8plD77tpnle9DkNHwL4kFk8QvgfHQUluZdv7j64SaUJsBw
RFJWF1kOsSfvzoBeFSmSMN/TlXuK+zVuA4aJ78AONTEZNMvracordLSi8eG8/a81
tj4Oi2nSv5t3rU5A+cYbWbcjj2Gb/nkJccbmcZnqHUD+RwFR9iYdCES6aFi1l2Kh
A3Qps3AacLS6Y2YDsqf70uBMrrjw0wjSdPmVR8cJDZk4b2sjtk5Sfe9ndRDUUQxC
j2aNFZP/ZT3fmLHKrtAH+Kcc9aeUlwtsnSLlenudWNZoH112zLoTzzcaDQXP9DXe
uqwM9ptOmV9rKiS55LQwL8v/71ucW01H1IkdshrlxGjoNPLWPM29/sLxdKqgWVNe
Kd1ekI5tfYLXHZUp+pkyhW4r1cMYWymJ38TVwMk+bdpxIcGXMaQCYhdWTTdM4Yc7
zJjyRKfIvBGNe+SyF8tuL6ms4QHx9xhdj1itKicGiXSeilxR+pZ/fp4D2udTtU1o
/01L1nCExqULdK+tRmu/11XbXaX9OIZKrZ/l4tMJOh8ABQ5Z1NAXi7/Usc6Wydkj
ujz0POh9iROxPoqU6ku5852DENLNqbQn3vtd/lwg/TjgR37iNy3IV05G6huLNjpr
oziAiCuQZ88YEk7dMxhj3GYeynvXk/RoYdYnHYW3WK+yx8KZvH71mt4RGj/X0NzB
HrUI18s1IAO0hNyNir8mx6fucqfdAmlboi0TfFoie4m0AOUhyuU9HNVejr8Szy8c
1XnyPhYuDcLLUqtkPEWQonpWF503ikKda39nqJOKDG53WBAYo5XWyhXk/6oIo1kh
9SeBohhINAQnLm/FI7pg/284narjHpAthPgHe0AD+Nc3wx5nHo43GGwDNxolwvdr
vHsjDF4yFXUW0ZettHchDGEAFp9mrofshN+IUzwqxC/617qP0JkAVF0KSj7/+gKW
BeuSs4v8WtTujTo7nAHD2oTS6wmg4VuCrg5FuMektkNZnrEppB515rG/YTsCNwPd
mkvFNLU4KVLq1ARNBx2GUKX/yAH61LOfI9V0R1SmsfDKiIhNaR34WfJ4VjyTaQkw
QFqghURtj4SEgJpW9ZNFIPwLwTgXBOtVHcJbJ3JSc1jag0n7W8ZGwkGBV7zlM4XV
YPKgtc+5SzAiTbyK9jhlWq2ewlNSNxh1/3H8vMUnYhwV1NXcVeFU18zbOHYnvs1i
j1BsynpXsfbcsYbgPx93CBBBmCyOsyQoZmjCoJ1uSQt5giBBYyUZ0Hn681ld9pqC
mqVmcOCVeOQ7DLMA21Z8SPhGqvWMv8QUCBJjWWiQ7dB/k7X9EqgVdyFtMagYI3T9
EBYae+5/bGxpTwj0LjDrSU9p+XPsUTjdnRK0x+wsth3OlhjkJxlNgDcFj80XJWhC
k7zA/3+egJNIr+GKgs4Y79hmDNE3n7bSXZxpOesuZ/S7naCyc6nxS2psfm7Cd9Dv
XgdPpRUi8crRNA6iBs2ArcAmxAxPXDellGvD5HdxICvY4v5FrkBgamzeIiFXbGlA
SDnAaAO8tkaDTEJts9pH6j5qLvaFOSOPn3LINEAzigDbgmSR6bPZZcgLkKkkWEND
OorK3By3o1FOKiQt041srii8WMTz5T5Rmoc+PqwkSSOj8Xj2qnmDMYZm+XouaXYS
9B6239y0ns9j/tulf3jwlcq+8aRtePzyw2OCSomdoLfQLb3+GfhgL7eyEsZe6EdL
1vDbVfn0c4JYhLKkViV/fNGEwKIQf9yECcOdYXHglp7KhNdNwnr0jvK95v0/fY8z
bb0YoDsokQ+Jo3ULmEyiV7Xjbmkeps603O5bZyYszBGLxGZSzrvER8vxFUBjRJOS
VFyRAd+huXMEnWSLbKqArlXqFBvtP5ugFiU4rNXHHVYglm7nVMrmdD7EyQDm3Beu
FVP5eaeWGlFu56c/NI10DQrIL8HOWgonMAPx8TVvTl4IP5BByXKiln4GS8JZtkvH
GcRljJ9otWYOXUW8Nb+gTn1v3xKXW+YZ8hFsuhytHAQyLSMRPoZ0BpDyr+FMJzTI
b0N5vxjUQc5EGoVnXBGNfC8oHnSSQxvTn3RJ7zlDA+gbo9wxu2Dsfvd2hihP6FvP
TmmeIfCMjZTbBIEAsjmSu+M982BXY5eQkIMlY1Leb3mIouNDV2Ml7L6TsXYVLLnZ
LcfC94XhzVCuTnJYmMY8RX3WirXDfopKrzFSd0voTNdYMtr8VwXlxlMMDfWLPGDT
dKJOUH6uZAdtVlEF1Y55qcMuwNV/m0INW6iuSP3Hbv4SkoF4kqGbITLi4x7hf8Fo
HJf/8DcmBGS7rm5SujyiLzghrq1iY2jezi89sYNvEHJw/LtqeBK210e/B8vtw8Is
`protect END_PROTECTED
