`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
C9MWxrti9qNSaA/Fho62hx6e34A+KfbpNm1oWmr+qLxA74pH3pCk6f56D7GEgpZn
AhAU+d/tX9LOYtTiODKLmH7KJDerIgdUSrrCl5zEAjJz03Jda56LBJEW3iCPqT2S
DvbUVQ4vDG+lm8cKwlSPxBU2IHExqSXr/U2swHzWtlUxukPYhdaxT8pdng/WZpYc
3OKYk46UtWw1nqexGTxQt+8hRhugYUewsHZQptowTdGijmPHqtTk6XXV1GpWXDmS
TPfZI8L2z1DHxSpiPdq1nu9OewJU6BG3XSBQTQ4qZp3xt3HD87kVkzLK0rhBhgB6
xdYPG6GdFp/smEV0YwiraVfx8xTQdooXQxoK4lkN84mqyPqrOr1iUgnZnY04GjU+
nuv5oqo6K6X186ld6NMIcBlnXQp+W8i656mooTi2FQe6HppwVp2lZkeeb1GkFWDk
wmgMZIdKKMJ3hq+5AfaJnYbpeH15GpggIQ5+PmbXCl1r8oRrTV9CM/ud55bF9WBe
sIHTO8sAgg9u261IsaeppEStyS/PUjejLLZ+9M6e6cdRSMiY7Tt8SlxVfqJXkcxT
BvozLGf16kO4kocgzZMexpTsbMgl+aIr7slprdzF/y04U98KUppMOgF9pNozExqI
dBoG5tKHZ717uQLokoyRZhB3sYKugR8AqURABmrdWC0c4uUNdYOoGb8CeOb6JOtu
cTIkcFTaotmY6IwsiZX4kqQa+4iP/l2SNerciCfXRLL83j6cxoVjfeBkr59o1mkX
wDb9ENMGs/65fWIaZXQTchV+KmPi6mkWdVhQkGVLdJBpVmQbKlBJOqFy2W0COOpT
WG0ExDlkhFmUfJedbxEl4CDzBxKoW3S9eR8RhapYtgufkuYKZ4YRwgmmm/OtixhG
iwW4QXj/2Ljvu0k5WVDrUnJHresm7USrKkkJfn053/BHdbbzo9OAObygP9+Sxt36
b4h7SnktlhxJr7KNRyzth0kVVq2zKOV58WgqxwAZfgMOKvWLYiyfV8zhq/jQWU6u
5W+K+CFTD2BNsZHB2uHCH0NGKdtLN3BUR/rSB1XSQvG8pJctF+bYjAdEuLGnNiia
bZoXs0FXSwDuT321pD5nxthBjOlAg2WgtPsODxTOdEzi8AdnjzdpcKHl6e7tuqDc
GYJSpWJuNu6Jp4KuvNExKY4xGhAHOhFD4w7O1q0Nu3HF4b6J1EYZBVn7Pgad2d0P
mJ1avqWkrYNA4O1G9N2mlSOExGXifFBLou+/307uZYFSrZIaqToEPbFs0IjRgpIy
W5opp5gOv9JR5XbBhRd/GsNisjNXZuZWqG201WttP44CKL9u6IBQfTT6WPor8PZP
N17ODTiAJBzMgUv7GI514P+8Ah6KZmxyzO7STfJPLMeMxtoXSQ0zU1uKwvt/2EsL
Qu7Yd5x94IAECcd6NF1uSlRZ3DXpL1LC3har7zoEqKFaSfJDxfeaqEFDjoyO92VL
W5GxM1ETA0LbaXl9/pAx4XunJwQ+FYQslfqA8GEQWb5f+FXRhoZXPiJ70J/fQHcH
tqQPeR75x1t2e+ac4l/foYCLv8Ibf0qJ6ltz1wXc1UwwSf2tHxBCuARTGgiRybVj
4RLa4ndduY5pAUVtdposUVDJu84dj78JlOcug8YUDc/yTkQZKP8wIvS0ZXAtT2+B
Wn6kv93wgNx+j2OFdIAgCvIPn/r3h5W2WpgiO4E81E5qL4iKs4fnqNxx4e4m/ved
7huUOeN7yp6PSCejTkym813PA8zGUxHM3mS0FdCu5YWG3hlfQj+2oL7UB3r06eqM
jU7OwszHlDUEc69pzItbL0nyd7Rp/mC89xzOR0U3Zhh7az0ym39MS/z12eaIss8o
g9qxJJz5dvFZ0uz+xG6Y05BI2pTUUJNbfYInD8tRmSz/zfSyOVk1gUCvsmtHDema
mINQ85VC1n4nDKxWb7sxZR9TOEe1+sAy5e9zHOjZUjQjCzcLeER5JZHvWlfIoAzH
5CVQqVLsNa9phPwudem3YM5W2OX7cpkUg6l7uQwPIqq5nZRrHlrBJ3Z3GEQiauGC
MFxQQ+zoiJk05hIwwulMGM1EtVf2sLkOdg3BS3wHoqrNb/GKFUzXJT6UroqA9lqs
qvhUEIKtk6EnUfl/RvYzt5JzEOKzE8Swn8UIQEk4859W+PFjyI7UOy4yL2bgq8y5
zZUAKFMzaY4TR2cTKNPATGSfWL7Odhb/qo4Tb4k8RHv1gmbuWW0gzVaSY4Zbi0LX
+cHNDXYINE3k6k2w+m6bT0R7jyzH1Tgr+LLYwM5weI3D3bdoPNnt4eD+dwK17a31
lKuFLEtdWaBnPqogvrsakZP1nkWQMDFN12/bpgyzEYQ0DhXfkLcB4nmIEsofI7e/
LxDvIdvVnFuS2QZnldFV7XF1GZrY6TlwDsEGvdPxHuQvny3c1LIJNbhlXKw9r4Ow
Wn62GP0ojVxTZjvqHpnNxk+O6bIyVQ/eIsFedzlhm6u55Fl+SbhHhJjD2uT8zeen
ZOOpFZbr317+uKGn9zb+Psav9XNbOOjhRHAzeT9M2pc=
`protect END_PROTECTED
