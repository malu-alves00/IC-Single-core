`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1jc1xto53WHlRxPFhejVLrju+t9ZFjgFHv2wMkqyvfBuvlf9hUGLauWJlTCahky/
5/apvTL1+KvNuXFvK/Ci4fNLt57wEK1XWmO1lJOaIW41h+MZdgIuMeEm4eYakuUr
EUTNpnEFyPcMdejjpuqtoAgMsKZZV2eRhAN0Cxt+dCLVYs+l8EVgqp+6s7tC3QKm
nt/Gdy9KjM/c+LVtM5+hna1lxD5QeHoi3amVrUVg+x+jThdyBPbNQ7guWLktxyEx
ztmpkXU8us/vjagUvh6UgRdaDJcyY5LWltJ19/5Gy5YY2TGMt1oGiNN3SubwxZzh
7jW+UFu36dRO+vfY1e2t5G+dA1QeLnuWusrvKItNQzI43L24TJEGTvz/auNnGBPU
uVVJIyedFod2AkzZ+MiLwcphpNu5BaxlLJvs2wUWaJjTlzmTTRG9+NdEFICZPEI6
JZMu/aY5L7RmhOxkrlVEV/L/VpDcLmiEpqg1I5wzlmd4+pn2XoOg+zr72zde7GGw
iyELCNsCJBlQcl0EenvOL+lyrlH9q2hZCCN+ZOVd9v+PysjSedo9AQgFMWVIBnZh
vmgZiv9JgL7xUNd9dhfhAShJmjHo0t80lAaMnnGDOPz2W7F5TUQeNjdt99uFQBwq
j+YFRx61ENW6hfNCwL2uYCuG6xaMkkpk6mV1AxjfIsrbiAdcrZRmHcicXuxy8Ifj
PDVq18tB0BJ89MFaUf+1SDofUqfyfZVVhIoHJ9X+D5+jzj0jy4Dz/YfaG1PuFdhe
X/djJrVEqEY5+pYslVi3DJPu9/hpXzTs9mQ6smW8vhU0qRRjtdbX8k9lPGVweZ/A
E58SVdLhkVeUyfn7dTHo4g3hIvyAlB7gM1GjkL6BvC02VXLAxG+dMMKdcPZwvmM9
7CA0SfgkbuvOUwXkD7STAOb33HqlxX0ilGIiHnq0Dhtg3ehtUd55brw58aQZW7DB
Ghot162AvBzPxCmWAlF4v71K8aRhzQgAmssX8+6QOWIcEEm/a5O91/sUjKGZx3kJ
tXkKPQx17TeCP6bD3RKve6Aqv9kXoJsRHCrtZZY6bS/1f7FrVj2yvQYIDrBf0uow
6hLRR98eDkU31lDGao/+sXxqDBSvsrdon9OIaTniX4vCcISQDkjSeuN8QhIHC8vC
bniEUbcJbvlHvCkFtUILn7rMHiPtf7jYZ/DWvOlq6XHDbyOQlcDr3NDwbEV3g915
zmRTTHqrvBDt5C6mct+obF7MLuFCEO8U2TaUMxK1Z0c=
`protect END_PROTECTED
