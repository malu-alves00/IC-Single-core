`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Q0EaLQNVlLIOR+luDSlUQbwfOF35zk3HWg6ymMypNXWuWMazYDBs2TqZ9128S2BE
Z6i9W9+a0S63cl6qhi7YioH3Bb+Gcye8/Bdfyppmi8VfsUFF1zrc6XBmA6ZTWakS
d8NNot5IApDj36Tl8eOozvedNbWVRoTGjMQQGTSutz8zjBGWXFDyqIQP1YQI0/t/
k1kE9g5Y++0GlWIfT5CJav1MHG2ZTSkrWdrGRL7mYf7yAFt3N3flCwjIvLZ/AxMf
Y96L79LCrf5y+/4eXWfZ3/pF0iFyKM8WL7gQc4PzEnK33dST1PgVEmNNTnT6e/DO
JwcT38EhjSQ5hRWqi8NTtHuqXuWwR99emyCCj+EzOW3/B1OEN0daZo/d4wBbmQhi
UVLPM38007+LkY2zbEiG1naYUuIHwNERH9KgNKAzcpRNyTZmD6G9xdI1SqKa9FDX
LTmwIdUx9sMHGAVjHKVwvqRGmpeO2BHFJmNedcPLAUNCF5b8DmZQqXGFr9clP/Tm
WYF+PBCwYoWBOBmHqblCcaYHjmjR8JBD1+Htp7XSAMc=
`protect END_PROTECTED
