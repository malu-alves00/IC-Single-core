`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2/U+OLL3p5lF5UegPsMUZw8738/r7TtJKKQc/QcsgVfUedFwCowBynreqZ1+4Zlf
fAkBslMCB0bQ/FVUn1dRp8v6W1oU8k6eG4GRwTbEgBuAjW55qVmwm/hyWr3eOnw3
cn3Tzg2qdMnqt/XwmkcFrMV5QZD8z3FRhnYHNQ/5KslgU9yb7ANkOBanTFwXIwfR
`protect END_PROTECTED
