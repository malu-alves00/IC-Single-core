`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
W+JwAyOwrJ2+8CAHRzxbcYS564KpMMGV9QciP0GyS7b1uZiPy8jfh0jv1Gruqf+X
GmwiL1k6XKEg9Oe5LGjxztCMMDCG5OAs/ddjF+OYIhKz1P2NdxZQdFtB3nl/3kYU
cw2lBDYM0Ebq8owTB9l/tibvWzapCz/I8KRrbl5Qf8r9KZnXasVkvtWCPKw8tHVO
dfugMedi9k16cMgg6SuKkPwbH7QM4c6cYE1xNE+sYKV3ldteShwOqUlXgLxXmTjt
45+znEp04H1q66bweICw7LUeM0l1bK+2lk9mqqd/cIy5vXt1GGTz5TVDb6MxlFT8
lxq8YdaLAThpwjRhUUtToepI4J6Nt5TAuFKQDw8UHKkGUYhqiWuHKdXvXm5lWDjt
RpN0JynNBpJivE7WUe4H3543ySSz76m+/N5Ca8uzUzrloHXixpeUI8QspCevNoeh
GIqgET6uH8OufbRGi8RxsjLODW1zyv6gnUgN+VYz3fS36MzlSZLdUusr4rP9Hltt
IgkBwTTUqOc8UPyhMyUFwhNSHl/SwvH07MpyCRL/KTcgFLzXhT5Cz4o5BNaUMa/C
Rkwf1uFi94LKtoAW9rR1tjtDQ0ZYMOuvuTbbGKLM4Ws6XxLLrPdf7ADS1yRA1w5x
`protect END_PROTECTED
