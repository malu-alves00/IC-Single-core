`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cjFWPNjACq35nkFqln/23p/Ucl6y8ODUOMgsckSrWl5UIq0Bzt/uMcQzTdqEOslo
ufpC+yIxvI9DOZN/UVXEnKPsN9kfV7l5LbfQ0yezettub308GWeDQzVB08SvAGph
Tdzkfg10UxLIr4wmA6IeLA6OvjTSUQNsQi2DWW+E9IUKtDxFFErguGa/K3FBeWCB
FNqDL7xXFCPNjWUMvVaQMaGkgjFWeaD+pDrl6IuRT6arYja1tzs/VRaKsQ3kj7dr
M4zfcyCE3eH8EC67NT1HTwLfKehy9xzOmgTzAhEvNKwRBYGjGUEI/3vJtWzIqubs
V5TDncGJD/4RZ3cA0pyCgU26E7zqN0SwOcMg97AEmzLAwoVyuDGWhfHRLDMzOX2Q
qkhB+YlSQUDwkCOC7T0YSA==
`protect END_PROTECTED
