`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PlgTeMdaWTmB1uYOm2h32bvPS487cxGG7aZ9xqp3Bo83JdEFdp52dINMDrQ6vPj2
SJQhktk7SVuwV/WJm4Vw9ZWEl1xqJnJAGJ8nVCQs553JZHQjGJz53T0W5yz2kpyu
63H0YuJh7X0ROp8Xh5Srs/OwqRsATYkln/iG1qhMzLYikO7I1xwkbDX32rBwmfuM
opfXFHDb8Pxd4P33cJUGi2wcOCCtYmGyvu2jfAdn1aS2zAWGtGoqrROvr8tlWY31
+AfvgBqDUirqQtB4CheiXAjBCFgUZ83yV0YxdMwz4D4JhC5xAm+yIj1zJexhTdqx
jIzXwfJaRMDSlhozURTxizaIstHz2dKe6HYfl7yarubIVn4HtaGMNM/y6Z31xmms
tQCD3AbV/540I9PO5o+jLDk9y57gwbGYZsrXSj2dze/h7x285+u+rfrPfMLvj2g9
Gy+3mH0D1/CIHw3Hq1IQgNXpWQnxuAsuBFBuMrzVV/4=
`protect END_PROTECTED
