`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jyjmV7dMlH2wRCeTe98dAcNLqfHFwKkvRUh5pYGimR1KJV9JrN4vs93jAE5R1JKg
9zjG1hjg4qb9qub41wx3Rdgss3oiMutzIv1EJPCRKejizZu6tOSEmmXea5EBu425
vb8Gt2p12BmYd2/VhvgTyHpH2Y3V7R5IDfJmeucOegqwJMWkzvCNshAOPYs0+obg
OJosW0a08u4eX/p21Hm/TWJh1CgZERE9PP6rP9oZRFxR3TCSiNFd0MHfbAM+tquN
zdR1tiQwtXspQJlR9sq5vS4POcDjooX5zm30dM+7ibhhs/z7ajVde0ZpzU7jo0GY
+HKZY1booEcIfiVrC6lmfxjIwOT2co02uGtK0pp4LRhy6a1RwFJvuDOHdi3l8eKJ
cdI6qmarQI2AzBw13xH1DQ8IjGNUX+H4/u+6i5sk+2AUlp89JjjBl54Q2ZsN6i2N
t4u0P6clTRw0TqsnGwflKd8zbn9JRfnWV0cYa1I25u38vtzH1/+F8IEpplvZ1KlX
Nt8yf6hni9rF2KNPmqsXAvMfMde4899+Xrpo9mxmysmdRFS7VepZXqrguaDDuFZE
V/2Pi5blVCfj0TXCm4Kq87J2e/uDYpl6xPQq5KVrtRAXpj6OsOD3nMOoE3I2+dKn
tatFuQQgtq/jxvHVlQbB5IbWfLNeA9b78IG71X/YZxii9vphjp0q28yLW2WPa0SP
NN1dKIKGxyQ40vThSNkUPPELykjrfxU8vYXFq7NFRm1FnvVOwkKZbH3nHIt0HQg1
5dk8CH5ileqzD4U0AEAfx/NCTw9E7g5DAHXXO0N8TX122X0yucu2/Gd6fYMYwBBL
Xb13aHChj9jAeL8LWkmBHz+HMheeSkKdJQqiYcHwK087o/SwGCH1C+e/dmFMbVHV
fg4AND/Cr/nCnb71bE1+CXpkbbiESSK6f2J6NqjhW0xh/K+YzVLIbqSOHkzhnhbW
SDwhqzABXlkOqv8KdC+7VjMR9d8irQc86f+9qwuyI5BPsQYg8rDdg0L2J1k/u8IC
pt0MjOWb3NKfIC1z5CUwjEfY9YL6iVYMr9GN8tFLG9bOPwP1IDXqpldIM0wU7c8R
PsRkGT8Vg14RUSPmN9ZwWSfspPoHpzO2/Mekf8qr+P9eIVA7v2tMtJI8+Cv1HOaI
44Q3+XchQF72P4W2w2Qc+Gi0hcgvs64CHsQdcECvx3Fp0K3ftc9wSNVTSM3TzukL
eXvcGtayzJLg7CFuR/t/EJXdxdr0edAZ90+crGpl37WMk3dYIQd2tQHJOV2nwkce
ClXgsNMsqJpj2URX3H27KVycZf90/BcX0yP50/sn9PnFqyn1LhJ5HYcVB3QjqSUJ
ty2gvGbjNOQC5KiMx+Y9vFCP7kI4yHiTZvG+cfzsTpiAK8N+TMM0LoAcTtQSqV+2
ysEb7yj77OwhgCkFRhKg8Rzg2GdAPXEpDraYyqP+P13guOn+gE9gV8VmHUN2zO90
10c/GvJpyeIcVyTJwg0Yb0KCi0xmQpBToTcZge4XCSnYF6hp9PswYnO3WBBUNPn9
Ky0CYFQetrzyxYwbADRM7fH6vj/ZCn6Z5DX1QRjdyZAv+cPePccvJN93oPXB57qd
vWH+k3TXmbmIjsh//CyECJSciAb9fB4IK2OlvuC2j/umrMLTnd12bFkeob1WK1RH
QclFGnHIg+/9zBUDVTAx+n1RQK30AmGWEr63ErDWajwSuI1W5Gr8f+LH36xBkD45
hV7A+tHtaHb1PY8HHDrrTUkxtV8gptnWYIwQqBoQyAzwKMCgfPH3yKHVMJmzXAu4
g67+3/V53xXFUP0sIEzK1pjrAWd435V8m7FjHjn7gqYMxfkzbNlAoqdJI8TM17X3
AfgV6xYLn/YyVtrW244qQj1xFpfJA3Ma8Cy4HirR7LefKgUdQR6gE9Y5YCbS6iJM
xLxU6qkRhOcWgsE879twiDQ7y84Bd/UpVCBjSLKYlJD3+gEJQklRWrLAR7WQM35N
R6aIZlwBXjOWCIo1+SDJmgAi94FZ9FI84rRKm90Ac5zlvm0A8jOlSLVc5Kqr0DCb
sw5atq9ozpuAv9t6Y1ETM6CHCj+Q2GPBe6RWqlkTx4Is7GmSu7beZNBXJx6mV0NN
bxWVmniWWi7ANzCI5p9Te9DO/l5USUapOH38Y9TiWaYfZYNQf//2rdSFWeCuv1SA
sAaU8aZaC3XbRkQNOB88rvsTSCQl01++CusCME8fdfYNLJ+UmG/49ud1mVDXMpvt
5uvxSpl2BVvUeaPfDr30GrY1R5sCpGkOhaEDfhH/yOCehCIdBIT+IPW5hpxQLYPg
Fwe59rrdqL6BMCwPHsdnrEDqxZo52Pvbs4sKqlfjCrVbZVeUSOXQRonguTFdc7Eb
cWmLfhTz9NXx7jb6OjggJam0c0Rk+zPZKBeaWqv9E+x/x3vy20VXlnIYDW5lSpOQ
CmglKf1GyVKXOcYMgrj4PdrkTn+7sDsBECICBHnMn524n8EL28ktCEsu7ukZxPpV
Owc6MEv+uWLO/zMancqlZmJJ9F3MZgN4KtjXhe1IVQjfehos9rBWgiU90L31ogX0
sMiMOMlBieeyGhKN+kWWFdvkBzg50nnSI27CEvNfjank1B0UkioVtJaMTVittHgu
zI5RuuMh5ZXWl4ekP6vKSaWZ/sYGR+O8rJwFtb1dCAHuCh1Hz7edC4DLAdd8t7D3
fRkhCCuYDIw8ZLJjGfoohAdTEswnRbRPmkxjQZi20v4NqliTpzCyZ2RtfVMiw+SM
FDlpVKnoJp3IcAB3E6M49lPqWv+MG8UW3pwHFu2LX42iZwX0YxxG+u7n+WzT5Ko0
puLQUmG6bsyyW6QEqu5TtIKUl7V4KhmYW70zQAKgcn8frJTIZg61rl5pkvQPF4sw
2KyG4nvjvHI52eGn40VtNsTetyYDqMLoOuMgnYtd7NeBZauBDSQT4tyxtkxFg7Kg
QF8aDz7HfthzSLdITWPq1d1g9X81h/FMFN9QPePnaDZe4qU4h6HgyYA5CLNM4d90
DCNw/m7nrngCOVxBCNPFBgHipOGbSx1lpvd5StMNOiEuUSFkSODaKbnoh0ecl+MS
eay2tERs1zKbd7vnFJYttmqPMY5QKW/UuftC3xLIQDbmzYVRwDhYt/kxpkxUSMxF
+obDFiCSpROLTGxrcvkwqxbL4M9jGS9pxCMMFMCSDtLZ6ax5ZcvpxCGqNmWOdeK7
FJmhRXD1Ur29OWu9BhqIQWELfYfkmKk7rcC6DB+hoSVRnRteJC3r4yJaldb7Y+Kx
uoQOlRIrnG3WbNgT0wOIxfFd5zyzsts+P6E1DQW4zXbpQFtt/qXRbXd/rNqz5LTj
cpA9o2F3jRgvehNKieDF0JpN14NpJszN6cYbuKr0RDDczIyiN9ClWzbFkMFlVV4c
igZ8hk3Vn1W/N9q5+YSU83Bj7wOf8jnmH0myoFeQ4X/s7grBjdaZWRq+SQKEe0d0
snSodGszlZZo0Upk8Jj6c1n1K4uScsL+TbWkE3PFSQ9rtcRciYE9dn4ZEM08scnf
rCsuAok13njvf4BeyFZig4w3t4a6rxkaje9dr1vqmgrdRGfkzoPmhPNT3G/ijtbA
sk4KSrIy3W9Kcw5P2zuTQNMAXQ4XVgby8G2WGqAv1//Ux52wooNQye0VRE+sWVCB
nQ7cUtsTLhqk8eopdmhxJO+I8hzaKyS6k6CEp1BFcZDhrF/OUX7nLzB3XbtqvUPV
L25gcpGxiFUohTXxgBV57dxkfxgS3LV5IKholJwRhirVPxKfRLPkpo/m3qSL0L7n
oJC2o5YNXI0DMVCPJrVtwtbkSKZhw0boo9NJgK/Ead3nEHjYo+sc1cFGMYaEFMbC
Jh1oPl/GIWSJo/B6bT/8qZSHmtqE9oPJapYl1BywkUsIln3KNARgZACnxotNK2kc
N/Hxv+LweKenBDPAshWEDcKxMhrUQu2GM7GZ61rx9z553UBDn6evMH+7NalHXoGO
dGB+VgLjuS1MpOpXmCnkUxpPqMtJW8oBkVXc3QEy9rg3Ly0ljq8s47zGBE9t6GSI
F7Fqho1jVRS7alW/pVcvyeos/Whib30DOY18brL6Neisbq39VZW+3RPQURPCPoT1
HgjqfX/cUt2amoCctpD+bXGS2pOlvVB/MwtU8t4So0CQpQQK9MSXcWxELKY5BoaA
0ItWfYSCiu1o556GOtpZJnAchXwScEvnLNEBR7JgzwARKA6Jl79AwV7BQtXaEbbX
`protect END_PROTECTED
