`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
doE8X/u9aflxSVHgH5/CdWCy9vO/X/taICbRMpxrKFyKHruBo6zySpBpfWQDPQ2i
u6AXYbM3NU1QlERg3yYZQ2auWKiGyEV4xsLykzw0Ywp2GjHy9CXsBHqAVMR+WFnm
EZbgPlotxl/N1/JOi/Z2Z+VFhtTLu8jNd6d5bghPDDghh6zFD1L4LNF5qjt0Gyrz
0LHuYs/qL7LqO30F05kqCO4gokv7Acv8Jve9S3G3il7ymxqPc5lSKpGE1rN+HRM7
qL6RBah5y0z/oMBhex2Rn66Jug/bsKBzvkatLMjsm0T98TGR94HmHeKIu4wLBgw/
K37+Ap0cLKlVQsgufKD5fsCoe8t3SnZbYnrilHQAh4pqdAlhPOT9+PHpRO2Qlu5P
V+W7aiccRNmE834lgDUSosOFsgR6FZ0jKBOWfMVMwynb9kD7WU91gB9fmTJb6ORN
WVS1Lbe8xbTy0KH9H90az6qL2sXg9KSTAEokRi9YZNUg38N1Lf3HZQZpWjk1ETYb
DYe9HiltOovuwE+QQxO6zHcRw6UpOnEFjv/i2rBnVD5rXKRxYs7QCx4xbUv07Aim
5V2J9fslKuC+rtsZaKjH16jPqN4S/H3GS8ufEKoNtgnA4xoBrHFFKipCjPXP/rKg
vrK+hOW0Ho+dR77T4cTCLkf8iCED/ZE/H4i5daLv4HI2ilDakgBxcHqc98tdgMxv
JFOiXh9diyzpCJWAnHZkQnX1qVkId32FsX55B5HYKZIQXX0RNrw7lUR72dqFkwdn
w7cwRE8SFx3+XmEyOkTlfVZr03L7wzex2lip5jqZvP2eHr5mZGoewa9d8DORo+P6
yHxOLZEb5V6Jfl7G41y+8BhIhG92Dxj0oXavXIJPT7cGHAXcQKhvESsu8hcvkaCL
9mFATSdZNbpgIuiDUfiy7+NoqhTS7n8jqAg4oRzucWmJhCnT2WzMqo4wK3KLNgSU
NNebb8w7CuuHF2IhRZIUI5cQN4SgHkbvDgVyPXn34zN3bICxyim1BW1jXWlBm4q7
fOWmOG7JalfytyKFQwjP9PC7gZhH31TlhVcOaThFCw6dzKm9KA0CL7oMdMuwyz7v
ZvpvqChbWiVe6W4z4MWzZDaJNUsbjTsxqw/eryY2B6EZLaqdHFZZGxc221u2jiar
IY9tfp2KUWVJkTaJMYD9DP84yRdiA5CbqnYyyHpAlQPYvroD3hhs0ukV/uycX+v4
BeTiUdGo+vW7nMddBiXBTHcHvLY5esuQn3heb8ZlVol78sm6kxYBsNTYuKiDuC12
8EYsTlEH0sBz8ITq2BU+ruPeusI74eLJINaWggXUcFsbeQNv49ONaKFOB0kpyfuD
DUAHPDgQjsD2cmCXaUTF8d2EonUT2RUTLeAeHyB9jcUQmwu50B0U41b8qAsJDP8L
jdq/E5b0q5JHXOmvghzHD+UVdKgHdExEo4MqBwLXygdxBQqIUGU1GyWRs921FgFO
Ph5rEEuW88o+yRtmEY2JO3qQFLIXJwEIKQgV9puzsKfYsdz7luS/r6kxMR9LGuaQ
PIYRD4jk2jHi3SkXg+s9YU33+acKcm356JmLHfTT2B4xo5x0Z4Uf77THcq+0KXE7
H5yZhPY5rTymhwuWhhVk4B8K0wEdbGz2i2PBw/8kRhWvDiX3TaXlbMSkkriOyPu4
qFzVz990El+xbEnWcSR8oaPHFfWcKM5BhE2Q5nvCe/s+j3f9+/DBuIB6s6S/A6iR
LBdEd6Gk+lbHv842a+K2YlXOXrdHIVe/UjHreX7RU0nr18IuAG2mrpXagnoSOnDA
OKeyq0THVRtcrwCdMuBhUW/ss3GA2yUacTzVgnsQJ4BfpsqCRDhWrf2xqQxPMxWo
TE7IN+6ayUzzVA/eBBc5mzeYI5FfQ0t3Wj6FXMurOA04+wlcYJd7Lsy8aG6VxBSP
EJqlVoJIKsM2k/g2hit1HJgZIIyEiWqIz8ypf+SFrG2+EvfMTITFpq3vElNB1HvI
Pp+bFRBeTEOVCXlJgrpUD13f8nazUHQE7vq+vH3kzxnFZqwW52ChjC2ftV0KivuE
t8ztXkOzYATcps+4bNcbEeKmQI8riPV6Zg+Dr2T0fa5GJGf5SEzNs9ikkTfASpJQ
mbL7ubnvAbt6ezxvW9HtcwsY6SMmDDdB7lYBdGvG2n4PKO6N2DqmltYs1kGuJmQB
74OiI9TuK7ivQGszUn7tj1shRPw/1eJCt7MbmrfXJPj2WrPfET+08Gw/+3C1+8EY
OZHHbtEg2Vf+PMnOBVaAWS9kv7x211yYYOoROk6KCFWlV7Iu4RNmnAgFIgFLLYcN
la/91PWcYiNLittE35J4StFCP3lQSeTllGq4izMGa6RqGqlkB+cu4x6fAzyoGSMX
481H/Jn1wLUGY+tVMxnh2DDpt+W9k9twRW+IZw05KQ8ZIgYdqpsCbeHXyLZRsmoB
wNdg+0oHSRIGGrgaYvXHezh5V1nnrCR2B6u47B+PGl6I9j3yvAplhweFw2PHz7Kl
skIn+viu9DGhy4OBYK6zsUTud0N70V8Zkc8PAbATw2hqr4mdcfRZ0ozCJe7868Je
wIkzxg7QVYRd5sl9D62hGGVsKU/kcYWvcZfECxEECCxO1Bx1T17h7KSuUqF22z46
UtiAQ1O2rrc+YPGltTCO8LIui5YWi2bkJYXZJbQLyizjdMwaDzKB3K7O93pQXgDI
2lAsCyPFQsCXbWvI9NURp+GNduFSx8apohfH0MeTtqiZtrYyO37SyybZrWKp/GDv
F6IILANlrAhZw+U3ZTjRfDjEF24l6iIKNzcsd04qjnU1VY17XciMGyoDm1RXAiNV
Gdq1nsywnQC2uD5Fj2pIkp22fdh02NixTUm4FHPOzNa9j4QBV3Vsesvp/DpTI3I5
P3Nii4TtWMYTqrqAgTZPlY6BdrtPWBKsuXoQvdlz3LTI6raiJ79PMPIdNcvRTpFx
n/lVzR9BTmBvepRgy9ZxQUtN2GHq+G1wUX54kB5FOGm5jbMB8WWIR5HOT1uNc4vl
Clns7847IMNWCmy2iejpF6m4gSPr/hUt7DDGkV8W3EeV3j9sex+iZBCAISSz1LPJ
M4fn4EPhQCVVAWukVkffurqybRtvJkT/EZJCcSrDkjXWVQUN1XLEKGfE3cL8jeC5
eR7odCdxrr2Hozhe29QVBxDkIIs7Zz+/JzlBdBOc/oFtmxUcxP5gGxKTGHkilNEk
VnJT1EdImtGPucMmHv0pYwd0iozXE32oHfPHyKYXYxd5AovVOHyNHvfYae2VmufF
ogGfjm4e2nop3WzcDCoLpne/dG9VePS23XMiBnmf4MSTjSkjnjsVNACelH5UdBMt
JaEwfAocDEqkA5MPfqmovR5X/Cj7MTHnT3T98yK0E00L965LanAJoXiqOpDt2AMc
d0mfcyyYm2WtNSvnMZm2FciQ+yivV3TnWid//n9spTE103KQ22IJTT1kj/xASaFZ
nzrK4sGOjKfWpHK+XFqT9Dk7p/gLOnvS6GXwldoor/L9MNj4tbH/51Gt7g3bIfkn
5JlqdrkxjAqbAQyzj7EbTIbf3CGK2ZMnOE6YHrUdnkDFti+uzAZr5dSdq6fRhtt7
eQXS5YIbWUgwhruUjh3W3KrrJrERaHVF00rrFXB53QmUXsMP3xi4kEy1hGOBLqZv
O3qL9W9vlprxrclxKkWIPafOrPeDrC+X5BgjXoIV5UC7Pu+L5g7W2J4GXvGhNiPg
uqePDMN5BsiFPWBRqhztNqoVdNPtU1KFLeCYCx9wJWUaXUj7mGEcQWWJbSVOqcTX
5h2Ve+VWXnBy2TA3ZEFr0mhsrUw+heat5EbiyeXt9E03f3gH0enybztCFfZFTLZD
pbG2P8bLZBZiQa1ETpjFfsia5bUk4Fpz0a4ibBdLKvBWMRnYhkfw2fkhowHWlvqs
ZN/w2atl6rLJDG45khDubsRVsIFvoqQB9ZmT9tHn1CLCDRYR3psMLaiz0KNEEopM
3o+kMvgBDEyXYQbNpgtkY0J57zvdfaME9qxoniYwYpgTmBUWhEOLW1fCOtuWZJof
TWOOIfHkRChjBSV9styO/XErC9DnFUgC1mSRwGrTY7TLUmzBN5MLmtQcEjur3z5K
hrZ9tjrilDlbRgDrEQR5Cfngsa8HdOdDeveXhMfpFHcvw/NlvuXxCfvPAAnOZzjs
kFgqd/+rxCtnjstQ7UrWvHbZkLQj3jJCaIRKd0X466dGoMVXeFwYUk4XzHp8HF9a
CJf4/fAgZJt+ioWsIo0kzV376ELNBL1RwlG1T+MTl2eqZsCkZ75FAfoKiT9YPSiQ
lOPzH2Xs0KF8uIxE2WY/rJ+OqyTQwKCjQbf1GLc7Wcgtgl7fvbybitggJEJA/Y2r
mSa6VxaXHoy3m5udmjNidBCSZSIPDWvufMV7eyqVdiNi1qaOnsxJEb7+/M4THTxO
SMfj4kVSuOg/+kA7ZlqaAlVaBjVJuh71faX5qa0Ca57LPyRD13ggFoISddK1AKzY
S87q2qBV5GeHGkDK6Tot9xEFRvM78WqW4aK4wLoXsA9LgvxDNT763jnGlKxiXrJx
t5M9/K2dHkmrUmlcl2kPbWd4+OWsehbG9rm3iBFdFRbei8ffcPj1+SDaFV/eFcdT
uuDNXSLfiaGx/LBbGWtgl3pBJdaVC+h9UX87fLrIGxZWh4VAa0vtXbX7dxGwbWD4
FnXaNDJNFshT2I4l0PM25FFtqz8dkYswZuv6LeQggBY+FrGQSasufVg0VppgPT2q
mOw/IyPJklN94SmisqAJkF/2JR8dnxouCMP3gtUfhBICahKw0hoCLLyTMJUE04BQ
JBmAB7C+xUyANgVGOQMCHOwfjEsBLmzGCnVx7tQDLOSl4FNi2RIFZOWoON8Bk6uL
csG1VrLclIOd9Pos4j5MQXFEnVj7DaQXRuhxVksKScOAVXaifGR/q0vahV0WUT/h
P1fuWr0YSVbI2SVXBRaicLCqWwdElfufiDUIS4onZxFeWcfNm6phNZ6EBvPzoFvB
HuImq7euxYfxtXCVc38mp27Ot3sWTEr9D5ZVRTssjNugXDs++UGzau68eoAxfK1d
gp/qgj+mQAW/jKob045/fUVAMlOckA1POghsgo4UUg/xSnWoKlO5ST4dR7iXVmPa
EA9k2LUVaBlJQJ8fX2CJelaMg7EmuYYsF7QsofJowNNTNQtazo0Xudmw7IrewNJO
PQoXIHMY6F/yjXR6dACdox6UEnM/Y/7jU2aivIGJUB4rfXAGdj+waopRzAy/P99E
6+/kzuS0F1rXeBvWm0bLeqkAs4OWDwp4FcL6f6PRY/TT4ZQN8culc57wE5RjiZH8
O7Oolf9tWrsENzva5BmpTj8kKLm8zGEPA1bB95C+zgzxpHwNx+DGwXrDO/tlkxRM
ipg67aSt8bQNN0MTaNxKND4yqwOGXGMToePXEpBinTcnLmKKj76z6lgouEJwOcft
qytMJhMh/ADekyyqYC8sdoitYPWt6dyj6UndcX14fjRQP1NoVMjleZ3S0qizJ/nz
vgomnTSLbwVFR41AmxY3+zV08hhgc+wlwmC9mWXoLlnFZvSNiYNtbOfZmc208/ec
DEZtIaYv/OUk9bW8SIfjLjZB8vUkD4///pq1PoUCpkpksNv3S9wpnZGuOBYPORHm
4T/90QJGMcfhlu3xudUPc9wXUXIRh6wWttlzKojprPr92UiV489K8l+2RZOSaRJc
QS2bqdq9bEeF+77Dmrag2wSXvOD69kuQniqyuJFdnxe8eU5z6Dy6buwbBJAsHxrH
tMG8371xVNxq50Z8Lbjh1w4mhD4giTAdrhTfWS7lLvG5e9m42uGAUbe8wsVwENEh
45mngYjao0vNlD7GCEc25DPWANahi0xsI7YbbmF0FUUwqtT53f40IGimZWmUBQuY
Oi9N+j5dxfoCMjORYqgYqCQcFQxBXtSKuQmVh37PS0WA6L0aVhfJb+rdsCMGNTsr
b0gjn5Q6JcYh1p5RkX9IozuS0LFwxikzO2j1hInkOTI8xbntVvCKTCKqusXKmDhP
J9CIVrb8/ybMvuHrLim85WJ0P/V5So4BkG3wVY12sBer9FE0P7jPH/ZG5Fi7zdIH
/fQp+AgfofTcwLMdBfqPnJubhvUhjVxav959UxEIckaUzQvMQESiauZEMVm5Ax31
l+DaV5Un0CWng89Fjic3e1JcnIZ/JfJQqoJ2TRp6mEOk0QbQkfkkEFcDMzxCrA6+
zesuePYPX0H1e8kWXddQn5g8Lxg323s1FSM2Qxkv3/NxZxuPdTaY7SYMFcmsu4cV
mpwaYUPioypnOR/R2nhszoB7UbcSpGC8qO349EQs+6UxdrOacS+gtvWCbaLMXXXM
kWTAvDfH4db/vVESeeiuVMz1RMyg9D7x0lf+w6DPlCdwakTjyzHyppIWmTlhCjhx
dYpJ9iqkIwiKkWYcO4CGJBUZYXFTju8+818/TAeXjPVl19YI1Lbn3QB40AqdQcT7
dMpfNvHs9cNSsL5wwXqksL40noW8uM0SrAI8x7sQVPxsl6cLZgoYCnxFU2nuCgI7
NTJTaH6wNkjZPV4p8WCqeAzcRh+TDgLtaAaMSKn7LYpXa2WSw5Pcn6b9VvCLOLUL
SUiRLUmm3dt5ldKb6nCAKhBhn+sYnsBsPFguycVLhbIj0GfsRIqDnRgYncrXPbfr
cN7S4f+OdHB8UWf8XZcYFn9LpjC+R9cSaoSkYqGA7287LYXk6WhK1SvgphbfnApp
eb8hTKKbeSLz8MJApSdXjeXctK3mYU/2C0ey45B8xr91s/62/jhh3s8B2+eu3600
/RipH/7WA0TQC/jwNynUipQ7MHOH0ByBILHpJ4kr3eW7x7QZqmGiAhGx1z0z9M2T
6tyk+iAYJ0NQqSyGLjz+NcRGB2g/mv6PlhpA/YU8A0hObjtkhgbSHQmIgUGb8JFA
2isOhlSAF3zqN3x6E8IkvXBQIo1kt6KUBH4WQaUyuG9+H7cSLPv/nsrAjBUj0rV4
gC+ZmPzHGiEWABNmgwit22lqU4bSNpXgAbROMMBPoxCIuAbrb90+PPXylmbVYwpE
MRuBWpmgufGY0qweV8BtVa1hVzEIWzj5Mf/R+F7UBe2ovo+DYukthkmhrCA3JKe+
DjV3Y/oQChSB3sbI6hKhOaEp3DKNDVqoVgn4SGZq4JAlnZAn8rIWy12pmNwR4F6z
rBZyquw4wvUkUmPo1hUbFPLnnRIAGyRKmO03W1Xo5aqaLniJ+15iJPediRvLp7EE
Ud8NtLeiFbZlY1VQ6yFH9KVGGDYPVx9tXhUtuc2m5PxN42T8QEbVB5U9WdKxFV4T
vI2FDnVYXuhGWYEWU2I9VlZnUrLfwBM5tVaPRVOAD+oHab2qDd59BX6uVZ6wzd94
fsvq937ImObo030kdg43q2ETiOpaf5yJKWMK7pQrTwndKAv6jgNh3DSYbfI995kd
eZIcYpY9YedGne2hkqaLbgxlL+kfuwCiPE4o4K/tGBfu56fj0PnI6qvCdNa2gc+R
6Ee8aCPFJeIa02UWN2TwmwSPb+eRS8QE22vcDO5xrulflnYiCLCb2JqG75j3rYva
8lRvBcwMWrt2Ho0+KRdMcG7FrPwwdnM4p1PNaYUq/qqHJHL0dOWSdEBsh02Fv5Yw
oszZd4X9kleCxxuNqkl/o+pcjf0paQ+mGb/UlZ2/Cc1rR9hWJfxQ2rVIkRbAistP
Y1IL2cL4MdxL/crOpsZaksdBFK6ko8mlVgTbfP8xkgExZj419ICNkkXMR3BHqt6N
1qYYFBz9cVqBpei/1Z5+L5Xv1FSqdmIiGVrQrgrPPq2SJLUfU5erbRaXmPz9fECg
KGO9Ql2459UMbN79qZFFKLFjhxLSCSjIbbuUBCQmkTuCeH1AvS4g/jwSoFlk6Nkg
nA61ns6Sc2YZuY/Cz3rq5O40t5OdebKNvz+blGWNecNvkkS69Qlf2H4e6CbpIyL8
AL2pzpEbTPHE2t/xzeTWXDoy2yIN2JwzHZtyj8+C5NOFiWoin0u6dXSrPwoN6irp
XKE22l13Cg24Zoba/Ruk1A8fb+aOyb3mCDJk1WoMNCzpDk3pAt9gfVjT9f9528Ex
TdCSD+4XS2MQYwXUbBex/6Gqw0jVFXb5lC9waFyKkdG+LgvQ/3GW2Hpjh7AmYi9o
OjGPw7hiN+biV+qVnme1nu4l0YKBSFDQhQA2mA+LXziUaU4XF8Iz/OPyNbSwGj7b
ODgHxumtG8xfmQEMqsGj22Nms1fGA6aYCxqU84UP0xLfW0DAp/Yr3w41Od9EAo6N
BaQ3UeGy76XU4qVGO5hlrUptUDYQPVYrTRasHRFL+aURcxL9s90bGvtwQtwCp5g0
G8BcxV7bzYT6ilXEJJXDDpWH9MbopPpS13MqiLCQRXkV7TG3bC0kfu6VPcxpnt+w
DI1kOclSRKJnCBIe+wgsnEnnjjMLCfFkY6mdk25HW/X+qQht41yvgND4TnzyvkDn
ZhuPIhmL0Da8PzL3Omp4S7KfifVei4o5R1zyZH0SwAWKzVLQfjAJieqw8sazzwtq
gWK4VuOgc/n/V0YWSsL1w2OBJt0iN2YibWoIy4YgjW3MQGwi+hB/oZYuR9K8g9Q7
c+wD/UfSYD1py9rNY0tzYw==
`protect END_PROTECTED
