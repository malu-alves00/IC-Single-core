`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
he/Pbp6VUdTQYBTqHZgPSIaFAX+ge7NNi9qj8e5HZscV+hX5oLWamXELAWLiX7Ff
H08DxHRbMlzEG731/+neBHUUwzzpjj3ELjuXXtK5tsgx7EyKPrFbgQvKZwD4M7Cx
XwGHnPCxLc8IFNbzEXrE66kz7ZBh/2pC7IoED2jhhXEIKwfyPLUNSe2ueteUJ0mQ
BA+Gc5gfPtyt+pZWjqxg52N3ajQVxqczQmhGYicmfxpAmvX6DxaltOqeenfXmgJo
ppQ/Zy8wajLHpXxzNUzrQVzdmBribRYZyhjh9ypjJnpzSlgTmhLP6q4JXIKdWRE4
Ysrci95XLMJi53Irm/URzH/YW21EShKeQ5+Pp5Zda3wiXQy77z32bKSOFXvgfqs0
rqpGXQn2tlpVK6tzAKQaLW2Pj5E8zAiNIPnQsZqEhYmFn6tMqblbLxQZ2DpTaXEc
iB0rXCGoaa1iWvT/HSVXjB0mbCDi8ZJbOsi+ID5I8GoG+4i66gkt6eybrIMZpc4H
O1PyIR/cMvbKi4sNNOmO0+eu9YyIjAu61d5FLqChv7XMhzTvC/DQNUylYD+NQOBd
yEwOwPGl2NDaVKq2JL5Ib6KG0kPpzym10sNeMVbJsBXzjlVQ0p2E461prbLweN/O
rMI5IGO1RjamCXW3C0HGe19pIfeLlF69Do3sdPeSL8W1bMNo0vizNWoJmvuPsPxC
5R5/vaDwYYuIbIy6y1PRgX1GbvdyDNvqs11mJYSO+jG9elfpQvFb7OaifTLECF/L
wZlE9dgacuDpa81XJk9TpGSwZDzecWh1qEyCPG4Jr7DzgtCqFq5lVaQ+Ox9LLYFZ
+9I+21c78Zkp9aX9f7YP8/GPaFWiDjZDvzIhxOUZ0bwip+zZT6s6WGAitvcFcckI
uUce4c+Pm+vk2Oo2bKES8nzXi54iWKEFK04unhl9+idfFG9P266R1I7A5KM9Juzs
wuO7Bj04NqoZOOdO6KeLjfjy9wUKLJYDPwd9zJ6k8+CIrYzvijkLEFcOvQhJ6n65
9nCwbrDwwsy8zcsqNCFNhQfTq25j0Rztylt4SlPmG3T6cvJzCr3sBCJfF/mytav8
CR23jtssuX0koTU+D1Zv32eDf2eJLF/WYNvHm5guYC5bP9m1dMilKn310Y0RV2zY
ZBZwgOhQq3FudZPCLtr5pZ5FEXQcN4hYhdT2Q/OdyVtbb7mwxVOdkCXdMzOzet59
LVe/6s94kJF9k6Ro7qHLIdYTUZZ8BwMzkpAwwC+/jCmSxoiSvLiLSWvjIN5gS39m
J5iTnQwq8blrQHMq/ytF3qwzIk5zgWtTVdiQG4X5GZxvRlzHPh7g8AlFbywtp316
/ogwxicrXkzC3ew0JvIRyRdcTKvF/BjduVWeBoyhLOdgQ7gRbZwtr4pWxM8swGuY
IICwCcVsvohG87gw6ZDeQy1fvqA/1H5Z9HE9BGC05eCEOMSRrbwXoYqbDQ7VXNKf
2vqyCOUKC0R55RPhxSlCjHcR/cQo0aKgADvgSDPx8TxxasR4utXFx4VO7CUWs9Ul
0R4I4d+kYAMc74gDTIW3ko0pJ0uQGuunOuJrgSR2rKCJ+wU2K71t8BWMLTUIi5zJ
2SdVdfxlo56ouPVAgVmzsutuLaD3XUSkSvoSNWIU/Vj8nj5b8KWmT+SpLLLIIJ8k
32W6B2QkwKWqkwKylwtr8m8d7XPOWkumgkph+nbwqaHTej5h0lWtmfdT96e7+Z57
o//qKjRsGKXn3WVjvWT5Ia7vwijhg8NiwOZvLETw96TVZRnngGgUb14fVr/LD6D8
6FEU+i3/2aqV7xxFycLB0wDngAcCU5Cuz5rI2srhuLhb98HDPasl6FASv0StY+cc
5yo6EzHTwAQFg7TYqu+n70WYwvegu726uI0Z2afxHvOWec7LqMWL/HW6tGEeNPba
kFlqq3FSR+l+3FPk2R9HX9vUSzl8DRPaRH6w/Ur+thOtBeVsM8MPe8CPpfTzBi1n
JCMCC5XkMaXkE7TSXm4zm7RyAUL8x25dD/8wW3unlSVkhOq3Ghe61PeYAnaKXxy7
kU+knlIQ3b/G3NfpdqgjRuYUPF+he0F6efoZmuP/G4UpSr6q7DWY6H1rAd9xXjsM
YRPKS8++gp+yplhVltCju5jtAQqBp/7MlARN704qfdMyGuDE9Oe9rcqBAvWY7zjP
5ii+4Ok+iyn3HLqK+/G6FYkdN33vcTJACEzEUsEGFiELUolz9R/+I6QGVK2VYnwr
XOGOBzNPysNOWYfE+K9ZVMC4tQcTCf4Bmij77n/O62DPSlL/PnP2zo+kum0eEZqR
f4A+PqS22tPMKOVV8JprB54BbQkpaLVlkOgJPm2TD2cgWnfSlp/iaRmfggRw1Y54
LlcrWY0BzoY42iHhHlvKdSzV5zBuK9S5lNE8ls4cCMGk+1gZZ26bpL8guzuUqLGK
VCLC47qgeHTbcU/V3+TQOMUgBt0VydHGFEw4ip7KWLOnCc6FRjHw+UvGVs/7kRyx
U5K0IgSGu1Bhb4Jz24tDA/wzBASOK3skWonzut94ghseSIRJDF0SVZ9Q6jo7pH1q
DSFgjx8UcvwJXCZ8PhgEHX2/nF5HaE2kqlySzL9IM7/6YaOV1h9BRvSLnc21ENjH
/77K2YD8/UYK5cYDky1BFkS1dDRsr0eq/Uw0FV2UQ+c+knUXjevajX60CS2ucLg9
W+R0pbdjr9P7MD9zUmJyUfYiJ/xNEotH3m3WwB8pBYc8aI7mutvzCtBQWgMMA96o
83fwuXf7NHH+5Q0G2sRE40X11uukITwrR/lZjZY7z+r4ieYmN9QDTMz2mTUUbp/w
0bVR07BaySYozJKbyyq4r06r3OBPGSyCW6kXwGYT54t+JCYDFlOq+b/LAZoqhC7o
+Hab/4UT9i69LWo0HnmNUpvGaAPKAEjjtaoyjb0qVixogFnvq8HI4HXnhFyVfTdt
6NWkiXSvUjSYLC6fHbVImcjziZt4HRiWLyU3zvQol2Zh3KPAKJRkpQQEOX8BNHEI
bHl7UcHRuWcLf7iqInaDpp6LSiW3l1lLoL4q7ycw15Q3MgnDJQ2mTgDTlHJEYnOC
Nbrq4XlRejGPcbSW0+IVfxsK2Zoh2eniFPNQq2/w2w7WxxgorXIzcjsV8tUe4rBh
raQoJhsaoF9C9bZhEgzdyuaNw3S9t1LggEydv7SAfQxy7TcRopuQ2Pc12VJhkVoE
kY4HJt4TtKyIaNuA+i1VHcHUSMCDI+gg7XVEs+TUtFKm6E99c494ESENQ7/NO+5A
tF5YziriWkWn1naNJ5PeljWlAslpVzYLNPSFzF1oRhVo9AUQ68Egdmiv2c+PgVQM
alg12TL8uP6zvu4bKlAfp8JVXSvL98iH02N2y+ajgCTw1GUsF2my9D0qfViTlvqw
b3uQma4Rr0BoOOGdPp4nf+khK+CaCB1ZyPys4HtZ5vtNe/l8FfTVu5okl/fW8nkh
EHHWCgnFWKu0HKr2/W6ta0gW5uQSbuOXJymVyLJM0cvcW0vnxVIKSvewqG3PFcyl
ZYk+7thXIRJ7OAj0o28xuEts14bcI+CYILdJmsXO1j/6dufb9XnPVoG2Ok+T4tTy
YG2B4GqeUjHwLzSTwL7+o6AQoEGeCivjoYWZ0WnLWi/EavAU26AVJdd1dPqjiXwK
X30WUuEu1gQ+vWyDPb6DZ+na6hhEzvgtt+vODcIvEpav7RJkqKVDvGIgzW0thLC8
nfVf4L23IhaTV2Cq0vIeLAz40wOY/yA+qPe+lMzhbAKcL/TDDJbJ/qJHM29v1XZZ
5oL6DybkCGn7QIm4U/OWYjJHVOY1CcnPVTf0csw9aPr88AgPcfNelnMHb35rAL5h
LeZBEckq9L8wE9oSGHNJ72/+kYpQx0exaIjrxL8M4fvAxVe160c46hQ8ikd811td
isRarn06iBpsSzcwFYGDfAZ9HxHH4laijYi8uXotv5z3QuWDPTBNy2Cd4o4B1dhK
Y5ulAzyz6QmY7vGyZoffge/LVERhAM83qiLAiQgled0BflwnrDIdgVbkMxGnDRW+
KWDWa1XViiJU9PcdYsy4Gr1jVmWXE7ATWPH9v2UFLDRAg0UyU8nvhdh9RXMoWNLa
VWIwzNdlDS8PAQe0/qgCXr7l6etLfAqe26cAVP16JOrnW/U/w+qqvu93igZ7HUvQ
q4gSU2HkBtrdS/otRtX0Bg6MKGd971AD2EspxAOECDm5DkdMzd5/5/wBFaWfgHov
FnawFAwBbGNZB+TXCsqw9CEftDHnBr3A/6d2EhUUv6BNGWOzuXrVpiJpd61R9ACB
wiOpK/wHM9SBfBgqylq8iDnqhdr6tDTE3/0/ShEMjwypwOjI9jQYSzE+dIezuZjz
O/iWCrrW3pjUigHjiJqh6ngew3iqCZ5PsBGk21ZnlRxqoSI/n80oecEWm10pGHLc
qHAkNHcBd5hA39YNBQ3SviREisKdGqkA3XSzVXoDlE9+UpoYH8XQ+cgCe+/Qfp1K
kEzBzFBPJLS0bpPZZp/iQScQ9h+yrIBLkJd6Jno24mbRY/snbPhojHrFUW+0BsDt
QOtu5RV1N/p16l2lYwqf/hmQRl9Qr7YVe38LfHuIuqsXk62YlK2rscgxOH3OTktw
iSKFccwB1TLS4ixcgmJrfkB6nBmZaxOVjuOAyIYpoi+AjmqX0OTe0rG/VGM4GXNl
UkeNLhhCIL/CchCKio1+sfc1GUKmZb5jdwdx4ddkpZb6H2cG+UJZ89Z+eUM+SSOp
h3YtfP+nKVraZrC8RV0sFVA9mdYScxsBCyC74nFZuaPQ7/2hDo9T/78pT1I9MeI/
yq+Tk3ypToNbEQgRmZv3mYDCNGPBBgiD0gSzFs6oi5k/0k116+WjhYjQTuFAzOSs
Ko05HY2vGFse67AlArbWmzIwriME3TLJLOUSvnSsPtwPX/jyxEZXTp9V+WlcGJvn
fZrsp5h5lyYEH/rGFEpxWVcFfnvwuhw5ZkVlzeGBu9kVkuoDAhsqcEp6r9tWXUzP
NQ7b8M53O0riGnNajrTvYtpzrRcVtQc4WeaneGBBWDl/+Cx3LPF9QJDXwhygUaqj
aWEaCgG7K4o+LE2/v2FvDG7W6xYcZWNedtmKcvOj3EOgwLSCH+I6GjAI9fy6muyB
D1UOL7Gnc6YdQD6WF/moT8lWfIomH8dGlMIzDEolQJlKJSxrAVC4+gMah6NxJO/n
ZQk43n2nLvHNmGEH5CXVynLSP0be26dHUP2nJ23iwrTD1XZcSXJfD16NdCnGJNNk
rkKUVNW6Z1s2W8Bfb2efXEzkDleCoheQ85A+5K6hDAxUypPStCri6cGXidC6RFzm
2OpJqbPO5Oq4DK6mbZjaudsfrSxHn0ZSUMG+xRoeg17cZ7FqFXb8PrmxJNXGzogo
o9dyddenrVr6j8+Jnts6GKM8DqJWYnLENNhHkBXBsuy9+q5SqJaddMvpOOaiWOXK
jDn8uEEYhH1HiHKCwo3B01AUmUG+KHl/2PjFPEVjP/p+mCTaPclwNXYZ3QpyOtKg
rnrrfC0DlY20ifgIAgamvKEdCg3iGXQE04aAlarRqg8hr7fBubhL6oNVsdHZkwH4
YEZWheXtmaYuJSp5DKFbGXunj8qybNW6EEXqa3v/xyN7dx4YByly2LQAb24alXbw
nDQ0hCJ+CW6mSArIc2FU1i1DwR/B3GEzWkA4EKNxuR67PBlP1guDlehAYnL3Mn8G
e2z2rP0vNFDPTiFexmUI31PFhTEcuu4uQfWy6PJ8o+XKR8lZzaQjA0p2PJVqoJ5C
PlvgJsDEcJt4eO3i2h6+UvtsG0zL1hf10dQ8G35rpo301PreDQZrRWQ8pf+8EmJv
FkaLCy9C5/2cNuLgQUKRaXHDXqBDVSNSH+Di1vaQgmAO1UpqIgmk5cGJAnhhqYq2
xwjpalcwzN1t5l3fHI3ShuEe9O9Cusm7SF//EIdpfUMV5GlWKKB1ySBfb4vS9mF1
GqesABQyL7aUTQNVSUpM+2bOL6/1S5MJB3GbVcwQYt1AVtItl4KRhuItU4yhP6rg
q+GG+GZeP0F2DAbte2eqorzNZHThmnwzQYTg6W/5DGS8qaFLZy/l1aj1dldYuz7B
Mqku/NiRfcYetvzdnVoHu477IvVMZat3PuFrcPQgjwoExESVD8ZYGcCZURyNYRCZ
YdmBrqAP8FGXlYcDBH3vp6LwnQGTz6YD8K3zH4OW0AFP//utR+To25BxLmnia0qT
4BuZ4ERXyDHhvotsJqOXaMe2zATE27eSPlxIBe3RqFbSKFaVCV5BGo1wHKteP+tU
r00cYFV4my5fYGZsz3pUbvNdAx9fbj/FcrUO64OSNpXE7Pfx8ObxsCUXmRcuNjpd
WwOPPOJiwWLOb5d7ya14FXtJVDn/2aRXhS8vAq0HIPkz+H0KQeTn3kYMHTxlXq51
3ordiOBYS5H3PEXAxnp6xOrFIdSCIu0HyoXzdJdvKHS/2omY5NHwmRxyDZXHWxmT
KrVq6W1A9xY6kOKkbb8MxeFF+DRPcSknLvEH9mzW4hNiHV3JAC7LhoAWFBf9AMTf
BGlE2pb482LiXfuMAaVu0gUxWJDO9Z1lG7llsaB6rlAs/gVvhKrG7vqekK6VS1gt
TENLEMXYYIvzPMG8tp2vbESc4fzjbjf2sciawtNy9dRU2Kv6SV9xxUYgYDAeGjG0
LkqVl8Cup0+n8V7kMJmZpb/nAjxnLbCtT3VNuKqvx6Si2Sq1k0z/spyzyTud+Q6E
LO5lSyGSomdnU0MAoQZCqBgRAKU7U8s4RFEDmPYB80kfxW6+2RnqveBxTMd01Hyd
pcRzzgA0Nn+Tw8Ia4EnhpLSbj05RMUsRuY6gjVegnLtkG7CWdXme5/uLEOXh01XF
uCpCecbpyKKORHCcEsjUhvm0wg57tNkk6MydUs6QjSGXz8Hf9dNF69JBhn1Zkxu9
90Q75b8Imh6IzGG3PzIXLLHYtYQEKW+/CRMPhwYGkfdWCz9M8rzd2mwIDM9kRVeo
hNfXtbXCr5+U29IVR9wZhI6rgA2RetEhwbM/uXBO2WwqXjtM2g4kRT+sxFFZjFqO
zUjzL8kutun6SXqChvYPXkE4K+6Pq/p1EdqWm1Tu5MijpxWGM8OJ49J/mgxhYr8f
GjomFRpiO1L2XoHLcPbfQp4CBzx4bPgSQC5J2M/wCEOH0vOE0q0iNP0Nr0ZshyId
32vRXa0nF9LQcrbznn875DJDzme+MjwPWcUb6WUldnty8xLIiEOST264trMIuKNv
3p2nqXg7YpD4t5p4PWikdU8HkfJhx9Gka1zgxIpICqhNvMMw80I2B4vOY1rw5/8y
n5b7uvmQ8hGEOElJPiAlqw5zEWCorJHnj/ndshpkH+g+k8C1vfsTS2BCGa6n6oZd
Q+1Gp169wpIPw+9j5oVBgbWd90VN9q/+ouNSkOv0TAo1t42T2Q9ks8yb1nG5tuyx
26n3/6g2pncWxs5FGv72lh9UUakC84gUULJEYSDrZjvJiZblIPBUZRiLM8LYL1vg
j1WXUkt8TpGYq2IpQkcb+ctytc2kqRTII5X4JK17Y3hu9oaC/scTJaFgFRuS5vlY
GfbOH/6BqYeu8tOZiWMdX+M9XZOIl0EBDAxk4Ue2w/LBpzq8re8rZkyRttHuNvk+
8abRDfJpVNmfNZ9ATeYSVF5pnWJ9KZsi8fyWSSe1+qNPqygcRrOPDUNHNABOuXXv
v3ZGABYh35xyFrFrSXEWQN5sffinSTMrmqV0yKj8s0tSQ1Mk2p431jGpk23ZB+m9
tbMUVz0pRFGQSvBZy12cA0YA8R5i8IfROZvX+oBiokR9+o/+BugDS/JAAwzDk//7
IejztmhDKOlWdybLtkVbrfUV+fQV6/rzCzOZmqFYAKFRsghTHtnDGpuzbxsFdRb8
8b1DZFAk8iO4OiMWBBsyYDMsfEzUT3KRo3R5lnPXimBp9YKlOamjOPLTV4VnS6m2
2nFP9a3xoM92BembynLu7qCNon1KH0Qv3TaLLZsoEFfN/5uIaSAtp7rUODEnv1DI
BWEWjFY9o8J1LKOVHaalg55TMmgXsBnm7JV2i3FnR52R8WqAz25DrfQYZ0Nzz+NK
cZiXAvznhVKEIrvHTzEBPFhlu3D0uhCvaeo3W2D9hBbVLcDoUa2P4DW4VTGO4Bmi
HPT+wIkZYO1HaAewq8JcFvQX7upw59vrOhoVOav7KEPE2SPzfMQ9WbRjg+dMhD/O
JJ7dvUm7CQ9P1ZZWuLqZf3YMaCpFY87mZqQNVXuhLz8qRW1fi/yAgvk+U0pntgOQ
mFoV6xzP/zuw9ycTunkXfHg7rmr/X0vI4M1K6HgrRV7qYtBjJqDWTY/tac00xtoI
FsasKUCXnGkdGlKLbkXkWkp+vWBrwYc9/d4x97wRJ5cDRGSd+vuG2bWGFOmjnPxv
w0i1vIc/llFr/vbACHOm40nXIavprOPTStm+H4ULWYxsRclgI5GVHkUALYM3D8sL
zwahsCXmCpZOgep5NEMkUnHmbh27MOOYl+XNuhUrHN4Nt5yEsHVsD2WukfVEWCAY
hbhnEAJi9fMthzBbk1RAEJ6LHr2MV3kA9aGeTZalK5iTlxMbjFi+Hf9u9pLhVeKa
WBXhAKjaY5wfJwiCuvcrFWec1+mZPKCs+zdMNyjU4ujLH6J1LtC0PNGwamW8wZZO
BH51Vs8ekYkDpXjNQm2miJkSXiakbYaqbJ2PVrsBiFRK0vswp73EpEQPe7sitHPF
5CVQpN/p9tCVnJdmQmRv2iWMVZWuHgpHCPrAfn1ZgWLEcmnpZevcsGdRkH2KaNrI
iQE31N22wz8YpxQvheaGTl1/c+/4GlTAhyZpV7CldphDKlwrI/2lIlaC3M1A/dPT
3uIzBEnKDCzGPjAXhoZrdYbGnfSiSUo0ycdsrVWAj2GuobhmqntFK2/4PNcn6vKj
b+8YUjSAo048riK6L00hHVzGfoXEsQ7zLSUZjW402rvAsQiHQbzky4/zefabl5mh
DzJqFE7N9NMBCNGuliuTIKHme7sNJbi6jFT/CYgv9Tg1E3XGTQ0LzF9dy4LKGYZr
I29P/ZBZR+RRERyOcDxydBuo5AtT2MwRbz3OKM38aSWqkDZ3wQ0K8XCh27R9yLo1
ZeJ2w0yOYs4cuTG3gtYtN+vgwlnzrSetzEImFfxZ0TEDpj4ZyFm+hohDpsFQv6Lj
RPCwxcgzmOD6c7dnaHg3YhSG4G3wd/bUrh1ORKopaeZneZN1rrBceyTlN13WqCAl
yuDIE8DDDuiBTI84ZywtOAYrEDID+xrmYpmwSMp7tHaYuqvAMwkl0+MJhukoWpL3
6CFnN+RWDSCzOFxAXfMaAzBymbyRBg4TP+y3jq3WDwt1VYRhGFF5cwB6bo9Zy0ox
VZUWWOK06cKEmORcIzHGjYK1k3gskowyBNKydI2POnEMoc21CMriGZNGF76b2XKr
qucoV9yaHYoNdX1LspjodwOFvmYk2ZJR/14Zzoyij4HAKqkKbhhb5prtnymlCv78
Uu8kKnVj6tZrtKucyzIR6APHmGA4NzbR4hn6w4V4PMwTivWzdcoBE3+mu2TkhaSf
jDc0tWtyrzn/wXygcS5VmGBfgI1ccWuyzfwkdx5jkfFcPc8+IQ4WE9WNYd2NET10
4kUH+pGRk0SE0QYj1IhZr+m9eohwmNNvubTTiUDE2gGHbKozMDkWCg05eqF/Tyov
3Raev5LwDoK8kBgHaoes5B8JrxqClt1kzdiuBiWPjZ4BecdD4motPbILQ1t/rlHL
nzoKleGmJEH5b2fLaeqfhudUahlwDXS+KQy6dFmEh5GLltJerb13d2eFGKpfApkM
Oj/5W4GLIBBEkU5QhlZjj4rXZvUa5kG1MIh0/7grQsLyJhkQdJygP3iSr2h1Owzt
kFtjUryfWwT8IchgVuyT81GJaVzPoMrB1CxEn5bIRVZsGSINekC6Y07nv0np+6Rq
k3P4UxBByo5ENLTc/b9zgCFtm3z9TEQtkYdAq+qFEY9HpQk35yXPSVGw4sLjDMGx
xBXcVPC3o/M9pYxgYdnXQwWtwlw+iQfyPA7H9bNqqUq3TYNxi/bgeE2GTWt1XXBY
4Qb3RDRRV3PPkiav2BJckjKdJ8znQEhEWIyyaU1KHWYst+su17znAWDqFwQE+0bM
JZaSD1eAzW0pyAgr7OBVnQqPMUxFzNd4NdZtYtWlv3OseBqk+p7xRrns1hKcFBej
BPv+I+wsQcj5R+OTocuIsBzQ1nfLfkoRAxVX+HiaTAf3sVgtj+Yw3ssJv8j0TAs4
KYiJSgKVkxnTiZlb2ytfLhrMP7aNDJMa9OFv7mCT5K41t09EL3JURpsSG9vQXaUd
SGUep/ZRM/KoKNB45+29632ZIvouQwi8Chc03syT76C/Rrb4AWbEj45xM1dJIu3c
9UBiixOooDMm+80cMTVNi0AtSCSI+cGraqHE7Q5CF6DR6fXTabZLRVV2gE0Tingl
Uv6W1C7dBc8KJWjJ3q5jO8AXKG9hpANfC7SB3BDlhA43Ly94eJ5G4cUkScLzWSAZ
rvCPzI34Xm9DT3TMeKji4pgo+koSI+dDOyWROtvT5PMaCwkD11T1MSaQrQXlQUQ4
v8pM2uxeH1rAw95UnP4vg3JbiuiCPc3yVdXhbe8XSdySVWhZOBPr0ReudGHFUnzF
rGGfuDEg7yvc7dAl3PFmw2E6rRd1o/39etqvdzoqc0pCEUaMtc71qn6yB4V07lIT
6atgMa/gtZdsV3Oa3Ny/nA/hh3BX5RBmCIvpWwiqhhvs9mifJtG+M6LQT9//SaJb
FFSlU33N3rizvgSP+RNEYteh9qbjdFEjgjRGhBq/lR/K2WV8pxLuDW94ROn0/G0N
sIhYO1kBTJxnVjhOJYwTstTRUD+zxwJ5wnSxnFjVTjQjlYoTu8BLTtqvQiWO9vyj
ilHzC/pArUeejDR+SbYXMhdSjg/s2Dboe+k7Qls4QTYOqSWxT7pDDvo35HZ11KsA
Q3toQcGWVindbA22/C9ZXNzcDWNOttfylWaesh9RJGqmUkwO1VeCyPVcArHcTZch
T4J7p/y5JQxOIyCD9H0sRZXScV/RMvTO0Y6ceZauCj3u6wclEwegtsj9h1mSDdSE
9euuO8A9SjTKWg6wgX+e4KSoYhxVz/pJFQxP76gbzwVxqICGe+7w6SDMHKw6q507
BW+P3mmKhIq/Gs3RoncYOh8sGBUGOXayEDJtHjC3FYcJFGRlPrLpvNd4mcjKC2a1
bpAHfjifxWmR1LZuFYgOGGTWVNqfDderGJidMxHYPgXUZmTQZ9hjt/WeKkbKPj8w
qgAljNbuEfFBtvXu57jXVr3rEGCeXmGRaqpsiltkOm5+2h8JGk3Vs3cz/NS1bYTk
vy99NPjUUDeGr8GWvg713ybb/HIyxHLV7R911v6ZDB2pX7UjjAy9dVNtCEEiqroT
WqnZdU+a3emw6rWO/srcXOiat4mYboSWAFviq0qtdfVT0lGxrbpJn/OHMRtengZl
3RZbuCBkQWKLAmQzsjA+7QB7jZljaiuM4kqeGjHajnQ6Zd5H7cRrr6T3C4bYAfZO
xOOaKzqNZMvVY9JU7wyG014ByacLtG9g0l2fM47WwWK1jS4/Rc15A/arBAUlvAAY
cFrj0UF8uLDp3FjOHcm6JppBaKeJY6KBo5xUcnmh2/+nYsKV+va06Xqmf+g3py7a
YV8IaMmFKcYFzG6ki3DuhA3+v+3R+CvigP+U3IIJMmCAyICNs2/AFKTv5pCwgnKk
Y35JejJ9EbSXc2y7YIIyrASXCJmSfnn4DDKj0QKKMO9g69+Z9S4f1wM+ipqjJuB3
YNAyQhY1x0QosdfXyL/y0fORXXEtdKoRU3UAcMkiNnt/bcj2PxWgOycSt49TodHU
gS58xr+lneDvWyXUg7aSC29wP5EIdWxvg3yvk0qveFLsfsW4ZdWW2Q1cxms9NdvC
s/Ay+YqHZNxGloMsoCfeqRPt37eUzcR7M+Rwl/6len6WsUfDZ71ow1lDtRxTUnyx
tN0F/EB1SVaJsQF+tQvK6FqyR9hCCa8gLQnMyoGrm4UUusE1nLoGggDoC9mkk9hF
AIhMezmKG7vWznQWtg2j3b8zJiyv5Dzuy+DFbQa6sjTApf+m5OwLu/p+dEjv3Ixo
Oye41QZP/Fx7fNkjW78gZ0JNO/CVriAGn8LRKNl55p3sjMjdf6GIxqV78lEwqBN2
k3mCNmOpTvef8nsMeb4fvGB7G3o8GEtzyQ2rCi7PTpZO1473Gf2gQm2//Yg7LYvG
1kUM8weNbWurLpcb7UlTrkC2AYD3/3OSuZ1+m/rSYkXBvjvDfjIeWUP/w6o/ScSZ
BenMPZxABY9SH12bgNtUqdUMqxCrqRtYqPXxiwyqPwPGZdQMmlQYJoiCYK+x6GA+
lAWNHR1uto48+jIqdfE6vQJqjTQCThS5Uxi/0taqj/OSwa48qRdbIFpduClE4ehH
GcNM+hyEJMOF1uZV0YiIdGysSlQ8puIlcxPPWpdhat5qOAM8YDMEowOAD3rmbaX9
9Ej+4YInsTwkfZgOj8P5Ocd7aa8AImveDMabtHEH2twzg5zaK/ESu4rtZKQHdKRu
12PUosh7hPY4mDrM90s9IQAGZyKdPMc+ANKDWirE/oXzdRhHxeIMG1cyvvoMfGGT
a+IPX3Fj8FW/f5pf/c13iWyTPi005G+ST8IFX2JxMYPQsovnZBlgkwi02wI0oQ1E
teG4l7q8DWipsJkZO5HDazokt0mpshkAMhY+f2nS0qihq7ZIZ6kdg9pFBEEDDObq
QVfaP4mxBvdo3CgO9MwzuaLSP0dKLG0JBGaT+kRY5iWLf20dHCPn3518NJz51p/y
Yp60CiLeDTWWdJM8CIJHMXW2mzXnXctEo1DAsxytl2zGnuSQioEU6cGaegch+hDc
wuclBWd/XV+a4gX1pnu+r5zf75kUYt/uW0CXPz5IJ+Sc3kxg6Hi182Hps74X+OPx
f78UHqIj+XDOy3hoDY8FZTJTUSHDZujLGh5lmQoKPn2x6LYZGGB1Zrx9UJaOQEeG
EZtRfjweJnEO8NPVjqmirKPtHBX9n2+bYGCaUhgZco6arD1esgl3A0gnE5ka4ebe
acMZEmgEuiaYPA/1k+ZFGFc7H11N9XFYIAW9G9Z0hqUsO+V7uZD004ky2x1xX9gP
abp2yDM/kVyjuP+AnBIG1C4fsTnFMFePcLibQrrv3N1G6nmBAhCuXVW41BA3Nmph
ERb/m1IfUSMSdrH++pfeqKN8ch1WESGlvrHZTBuiq068rZGCoxPIFWYBdMut0OcS
1RTRLwb7k0MSTY9L52pogZDFIiDw94D0sANCa5KYrPkeDiMmq7S+++Yl1eD2os4N
kWwxJ44jZKqvfOAgSCMUAQscakT/eTJunPUW6QiHjmJYYlauYEqtYSw+/qrpnp7W
mrBXZ/UCxhrNG67iQpnJWknLTXAdRQPILZxOQ1fDrziQDYPpt7kOqrnCedh9dpSD
451NTY1fYljvHI+NgWBIYpVSWwIAu7WfO/BF4spNoPLdJa6Lm43onIILfZDwjHMp
jMeUPcZQel87sZ8Y7QOkJjgC1OG3E/YYJle8AbULZPeVz9mGdxdTFpv/flQeWm65
OlBsi25aQ0n5ORWBLzCsea52x6gl5X2la5/3k9nHciCUosxFdmvPCjZXkaKyn+Rk
82Pc6ZySZV4vnO+ViuKLcEqd0M4JpnVGAs8BiqTW7ST6XaAfdZzsauJ6vEqsgYt/
SUHzpwF2M9xGh0ea2w3+8p72jqyw6l8tOG3wvqfnwkmC4aU1QbvdCNyDRsPW9KjV
7q35HjanO0ZjjrhYoT9RX5VDPXahZrhTcqSpzPy71MNTSCqVZ71RlX/LauL8u72M
kj33GqNMdYI5gIPXhMQ/hjj62lOwMgcMQNEQT8YwCv8m2PzDOepeeD6Vt0sOWGNZ
9H/YjfbCc6/iAyeHrM0yDU7cJ1lyZgMikyaRu1P7AoAsX07Bh8VAkivT1nhUjAzi
RjMaCj5fba4JwCO+dqUziiGOLUZhqOuiCWt7Ho9NQN8x1RU7AUyHmY7NNcwqCIMi
7fFnoz0PQfL1ZHE5yJq8fynPAKQqYk7XqgVZzYwKKcd21elkqae7Xz0XAyxCMJvq
Gdm3gYWS2jh0nnT62PKMm9SVJDK2cmu+/JxLB4oC7r2F0Q0TkFr6uZ2d5XcSSBnW
CXWDYdqRKNlwGAkULouOXYKDRx/bf5543vRBskrP5jPVbfJikq+Um5QQU6mObunp
z71FQ7Lao5mYDtMdpUssVea4vO9Kt1zpPIUKXPGirteq0VUPxBlSxyhT9NHkDADY
ki57h+FA0EJ23zF3hhR+Xi2QKU+n9W8j1knH7LP89NMTtAKo9KktMxkG9RvshDwt
p4PPvw/B8DkPa6hie5JzU6j2OkX7bJ2zly05e/OFDRkIoIiZKE34ClaUnks3xE5z
qTrA24hYsAaUtFwKnRjsUv6Ecp8Xd5cwTSpqlaCTi9lppfN6oQx77JRZQIePG8o1
4kDrBDdiND6Vx85LWr7zxVBG3p3NzGQvEdvCwfqhNDHgvFXpbBvhynHkkJzgKSKv
BDWJclLzpv/dK1QjZc3kQtV+fyh+Zwqn0QvVIcdlxENOuvZFJS++LWuuWi2UXxOV
AW/JC0FciPV5mJkLis++64NEV6BYlhvPOaG0HM43MOAkytcOpRM6vqJK+Nrv4yrG
b5bUuZxo8ItSXtfdq+NWGbUeVdT+hOxJaxZIUZTYBUhArOOstSPujLwQFV4qTHOZ
ZboU5L+MivSxUV3BXvkI2fygWzpIkUAI3BuoA0Lui5zSYh2MsK32T8wHCfwQE+nt
k1i+cGb4tR+WxhlJRt+s6IzNS08m9eIwr4LKv1fhBxI0zZ+e76//HEgbL71cy6W8
/TNk2BUEn/J6mUYhE4spgdO/m1kPjZ9HPYDlk/oItVxk4mExMZBJc87LXf7NFPuz
Zq8MobGG4yqaFU2x/LOGqPTanY+6I3ttTaD09o4jSPzgVUY7A3M5IsFIkKDTmCgG
1goiP8gbrZa/Z9CpEpLKRHsnpPN0byxdPjkQ+dQe9hMoOaPuifrsaOZG/NjnJhTX
U86YHmfYn9KXq/acxodcfkTqcqTkxjNUdufI/4wSaD479FkWci7txkN46q6WD60V
/Gyw2iN+fEtF6NbgWZOb6pc/dtzTdJsQ0NRcfO8Jl6mH86pdGP5o9SHLYD1ykgp5
Hm7bsD7F953TXLbQngmAXLyvtGrtJRnDemLGjF3os+3u+ycm/zQNXvOgbiTIWfQU
qSt/xQMNGVFzoWUxLQiC0CD/ALzrAJlN+Bq7TJ6iZOK4crOhWXh+uLV8lC0I4FLN
uSc+nSDWRf1cMeMsxqXH88tep7ZPnmDZH1Cu8IPXTB1o4kCFamk0FZSw38BBy24I
XgbpjUfQD3m8ZdeP/GH4LR85FUBaebmCsfwTk358MgXvs5m4I/kTd5Ky0CQOZ0JQ
wXQzkY46QeMkOYkizIWXragzjXYjYUXNMxi2c7w2Q5Fe5icIT5e5LZXSB/3a0HOo
1uXDBF8QX8zGo6sE0nXvQ7MsLJy4cnGsGbJGX8dVYYwJRwMJB47oJiuJxKbub/nV
hDqlNifuPpqfggmoEauYoKWAdgZpfxwfowrOWc01Qjju0bktcWIXtrH9EQ96ovfM
fXA8C48CXVsNjZ3pe7QslpS6CLcFmE1F1uSaldASIK36qiX38MAmCzlSDlAyyokv
cm+be0mf2Jl04TFacTTfE1jU4xjgR2I/ZS3JY5DW5R6fZpr+MNutVMV5VxvP5fv/
CkOQj1lUnd0849pfkS8r0Ro5D5Rsn9zv302O5bn+WPP3XbWm/sXtW7mudOad8AAl
3ytRjJbSfy4bUiQMhVcCsOPyyiA6STJYi2yCxmpSexlZoaK0r+eyovGJ/MJLS6cN
IOJ4cCvi2SMiKMWRDwReYd8QjG+ff8rKlB0f5RRKxZw27HoNcrNUSsZWBsyIA/E5
OT2SdGhMPPrQfpIugOKgEPWY2vhTpNbvZDut2QkBgWVQBfju9jCWGTtq6n8uu6bc
G/dIQvUZQ9L7CtZ6iDXLw5WTIiHNGcjFo2IGaG27zj7AI0ZR5pui8QcaOrySu7CF
naeI2FSk2lEQz3iHJz13qs13zhqmRACyLXvamBUuHvsjQny6+qBcnKYCSXPPdNGs
bJvdA9G478wTM5EfpyuhSGjvWuDd6TY7seHzfj4kCPaNuJaFm9LkKAUfUoomGMpR
hn8X+m1xKIaAKsDRuNG0Q05q24Pdfhv240/w903a1Knv4gfm1r8JFb8iW3RIkMXT
TU2YE7CLpgr7EaN4ytolM34H9ctjXcJJNeQLYVVwxzZYD3UqimZZ8L6QCkxN6jlE
RYEfudr0p8d5uKSKam4U5CWIt2onDda+6i4hHr5yxIwI0e+m5b3fpIbX6pOTVV/N
S9v4TDZjaioHBebenHtMufHSXgQRztmZlBQoijzguuNYF6gff+NCDi9fHc45PGc0
1rWjTc87JlVl6AEopT3Th0nQVGCnzLU0OeCOjH1G+ujCiM7Sbsqoe6VFtd8N9bR5
8barC/7TIpFFrQdcsVyBXFYntNmDgSACXEsFC0O8/BCE9MkyUO+nsBbz5srvCxJ/
qSjWQ5z6Bvp05ZJC5uk6WN2hEBLWd6ohpxpRV+e18Pl3QLRClcvjCRxR+OE/6w3s
+w6NjCnisLRwb9E03qasEj9CVCErtWEbSwPepzGHBRgC23YwFrtJhGImsBrH045k
goutUD8Eiy5I3K5SWaSBSMCK8nrRnxyBBWpmZCLQDxRilfY8X7Hd6fJuZq/40VjK
FJYZcE6gAFVf0c/HRW9AnuCf49RO7sRnFBpjN3MyQZWOxNGlXxJIqnEflO6U0fCN
f0mbqgjOU8Z+lt+NG0EgFtamCar0VficPsW9EcEMdeIUDybKMjneaN3iFaHDmbQ3
tAjyj1IM4qY5AeGeK3bQs41LndqmOcKzDMA1DAWdxsG0YGdAtP7V9DrIQzAqU0SA
BJ0YWnoBT7+Sh8S4MRaIJhxed1xyFEmi8HtfEKvyxVgrXeLEHsOl7tq4tUToADTo
YTEt8ke7qi90/xMpxmPBuAoyzmN/fVzOOnuASA1Z0cO7gB9Lv4nlbtPKeoM6aJAU
YnztY8G0Kym5H2kvoLpiO8Y80vAp2yUjSylkS060QNpOzbfcPeEDMSOOKT42YLgG
jllqT+wGVfy+t/qa0+/L/y4JmaEDGrKqWnmG9X0BShQSrdnEL6Wh0+8+m4GiidgM
31mCrXoeQh5YKdUDZLnDHkPUzjSrpUQGx5V6CmzYCo/Wpa8dNUlRBRy8GQKTTcTr
H5TEEnuZtTHKPW4Uah1BSWg+e0tmVuj4k+CVZ2Adi7DGskyS4dLgrUErgt8Iq6vw
DEshghZZvE5TbJXTzfsNiwZSa3hPXSaqkwrZSsPmFB9V5nz75Br7COS5KJS11UN9
+F2bevsNxcJ8KjLPTLoyWSi5FJRd06aW6gTOFHIrQpKGNoghJMdbyEeZvOQt8hH8
0M+V2EHez3ghPAev/py7wur+aAFHVZNVOhYwmcI5dkkJfAwIfw14Q1s1+TnaMEF1
r/4fTQbRJKaPva5pBxN/6NkXHZLmR4lIuc65qWfZWzhnH5IjnbPEK3HheL5Qe0oP
keVqL5GtiSOZqPJNLVAQOONqJOelauZvydTSNwQu4Y5w9HEH+wyqIhXOaHhfvXae
xu4htImGu3sZGndxcmW6+xfItKohKq7yvg0f9QHO/eTQVL+vanIJi+F5wNdOzwm8
DKh6suhRKORUhQArIVWZ3yRWvA72DhX3XN4Op24s7tSd22M1E1EMZQgrSQDOkWRA
DgGL9n0l+kg74zrkDrIFNz6JRENCfIvmY3iHL2Rd8VhFm5E9puI4/WTosSOq++am
tew+VGQObljugQvsbmArhT1OtKelPRuq+XlS9llBc2HC/5H7a3R3xJr/yae6Cf3T
Hce2Oe7spw8Ly5KsL5CMI4Nql2FrMoMU1+wANT6F4arsnry1VLMXrCi5riWKqf+S
ne/2qp+91aUePo1qLDjwLpyh5DPMvo/tFoTNbpN+OnIReqb74QjMkK1X377vLIps
iVbdMSWjO0ElOq4DALwqBxVnt/yBC8fXdlOZuUFgJ4lnlW8qwzEPkVNgMpbqhRoI
/kQWAZC+f3jcQpn5ne/LpU/WGoVry8tHPZtq4Nx+5dNDTFZrnRg9gz/S7AHWg0sC
2CQ3lktKziT0W7aafETQJHCGGXGCSOBoxXemBJ3I4USjciSkAWM1vct60b+R7y1+
tdx18AzDoGMM3bUzKTjgAaRfI6od5hX01QcZasFB+ksdIIdoUrv31Zv8gjK6gmrG
I7LxyQQ7510Ogr5mwi8BI69ZRcSGm4SkRTnpQb/B4c0ir/DA40I0oexd+M/b/OeF
ggccsumFJR/o1jmp/BKfE+FgMPdOUjZBJ3antA5dbg8esUo/LdF7C+3n5bfC2E0k
JGFeDWAMl90E9RNF5On7LgL5UzhgD2kBiJ9j7AZtehaVlvA/Bp345kCjBXwpeas+
xLLSUB9GvXL+KpmURDJSnEXAnH5WU79GwcC/v1vnoRXqRvgybkj+5xnHLFWaE1dL
0e2sYUg0d0TJvZziNo1WiJCDAfUitL0N4+smXp08p90sQWXlAF74PCm8CjCqJLBS
AJVU4+d+tXlqsK8Y4X9iQToT9qsLDNNYIms+WelvvvsSwLsjKaYEleofq2qNlJm2
pO3Sb8bMrS99dz1GgWrrrviCSxle7RIxrTajnWakA4rR27lTSolvopRwsuVgEGt2
uimq630gvQNXHpMX76rPVxO5DKLvXqdZGbphcRV0BA0nn1zUhDCFvjlJ6tzlXJ/b
rm+IxliQHyJzKmguCqsCyHOjrpQZNtTlcK/6UdC3KVyyHwkM5IsU229qZ+khioPx
h+9no5otzUH1/luja5eEMVIs7QPYsnevrEKIveG4YsZcPWsdvZccfwMCzTJ8IZid
yJ1ktfkeF5Nonv5TbPVU1MSUbxPNL+RkBW7uCoJ6huLjdmGsWCKVpEre4nrdL8EH
mJUTHRSpDxMIHWkI7Paqyh4IqVrWmVTXcWCjdsAKut9bMjClFnGw5z/HbRaXBNTc
E89TK+G/4pdavuoaflqnNPxxQSfg0jHHSybqGiFdDlh4hRgk2Z1Q4yFewk8IR1sv
RaoPjSq8e7lyW2s5+jv3WsDDt3G7TQCqhaPXabSAg65+O1TLmg7WaVDEAJrUB+Cm
bY2v9ntmRWN7aq2AbPo5caiukVGzkfo/bVk+J4xTrDnPptTr7DCvCZJjMYj+Fwdv
Oth3CrxE05S00eeEvhZSxhCndg/AIKC/JwdGiA9xzxqg2fGEkTQspENGei8v3jtX
0SwHWizMa1TCFJmyYwMUL/Aj7JpLUE+ldp4xJ14/ymS7lQfPhNZrsPZLL9OnQkvK
zGwoKTP9KPLfCrLm3+HtEWBcZZPRUVJC8XWp1Q0GIpRmyQVWRClmyjjF1aeiXUlN
XefgAu2rDgo9383F7e9aLPbq0lCiP2cPX9P6FZP9kkYALzg2axlw4dKUvOSlWJhR
2eo5bYqldidmaa95HSeAc3wqd+R25yAKlKDSr7OED1ASfJqS5s777Zmg85rgmDJg
yggVUAa7+sLVt8Udyh3jD8AZCU3sXkIHTJVAaxcsD1yLI4Q+EgVi+tOsrTHgCjqX
Zr3UGWEn9yGavrtj3609b4nOhvmnlV4+nCDceybnqSp4XXnwgmLD7tz2DpZUWe1w
MSCMDiMssA74uDElgLLdo/IWYZGdzFqkjQ67SwyIkZLTIHXoRRE8hx4ZhV2Uv1b0
9j7zhyH0ddbjqipX13PC6JetiZWMVrXb71BZ5Vb6HHHPdn1f4wy3jAi0xmEkwe57
cJWrdkzWAmqVB26FIqs4pVgc3+6za4DvN9Oc8y6Yec7nWvXcV/I0uOdeXVidr0eF
elVBwQSa9+g8WJSO/pe9B/J5MJt4WxJWzYSmkfCf2P8y/t8F3O5IsF3hTbOvh/dY
Z9tg08wOYb792qOphHhhowwlwqxUhubcnf3zzPjbe9HBX56TFsxWv0Mi3EM+Clrm
7WmRwuRMat7YcIXoLTkWkA1zPl0bGYWIgzyD7f0k8bgVjvUlxpKQIwAszT2yT3On
pvJFIQaLGOUl9e6AfEOQH0g8/J+51NaP2j88sTzHVDaSYon07tlNohMsyfj20qhe
ab9BTrWduz/y5GLctjWWFEubpyfc/urgBhJdswZJpnnQGuLWC/wGlooPW3ItaN9i
wkafFu5ABOVW3hkqiJUzAHrLGLgwGjjgCIJoYZmrzFO3ud4g5sh6tVki0Cr8p52w
Rs0RsGtkwchiiyPxOH0x4c5OxRC/klwr/bOLj416UNNtRQufAdVeqq7dmc9krMZh
DS9GYHXzJKFw/2cdzxVxlRNlXhjpQ5ZeMmGfygj8A26aXI/hYtoFVsex4ouxWR1A
Ra6CgZVp2CT9XyuBWFTQwicV3b1dh7xscy62SFGTEpgi1a7MHyydYQlByc+URZUQ
7gBZCaGrIe5a9SXcitZsEc5il5McMXnluYJBwEa6XX4gftWJ/dg3Y7Oq/bl2+Sfx
QpMxT5gXf/YQM2tzxLDM0OS4brhQ7WHera6t18HK2/gOHxzd9QklJ9+62pmflGHc
quH7Cu8+O6F8vMb7U6DCJrfKk9WW7AAdfTMnD02qJx8X1/2agy+YkTQkxVUfYyGH
rNmDkTMj7dZ4lVuQ0QXy2aImqWIckrzFnC5lRy9yLr0pEOzCQsS/iB+fxT62JJdf
Sx5Mb4Ei0N5GXeyRP8/XNaub7gwZsW9hBD+V0r4/j3SFvpd5Wjf+9P2zyi5r/gM1
a0J/qgEl1fwYjSjvWtJO9LMf1Vzh1jTW95/HjocK8c+sazmvYLPNRUU6+joYa+qi
ecxKMvtjK4eJOdgFidHRZd0MvIWLct/yN9QahyIEweOC/4OE9kgDtvleRUE/EVhX
33f/SpnCXOYedcFbUm9UaRPklOSIhYV5HDL1cLoyWsWN3yZysqhMoedaIVTOWjGy
f2eFrjCt2JlXFHiO104QxWW2FG21u9yDNzTfsxIfnHiwQd51sey6tdClVj5qYvhr
qhElDz170qGM5S5ubcThYgB5bUR3D+bKtpvlUPRKykKiuSswZDzleOL/cn7we3kS
Xq2y7epNkh83r3a0D73bkpshi7lb+qU9UpwOkYCgEGDy51oB1/Fu85KjG2E9JIaQ
7Hp53t/DEu2nEeLepMuR36q4SU7Oez3n56kBirRnYCJmxL28PbD7D/8io3nHADI9
rL7aQy1ldAX5WxAiWKyjebADa/jAORV0qng2TRFvg/1EhTNm3yr6OGiFYQGiF9Hy
xSLkfn2tdtaYdTzH1z9xhJ8v7r649jS4IlUPM2YDBnxslK24ThWnGJ/i+1eFRxq5
dn71voHuJ4luumO/b9SMrWkH15guqvfTXhJAwfFh2EcZqMP80NUrEBtzG83D6gyZ
E+VP6hcDxTC7jItUXH+Ke+Txw6odloEgy/Qgz2NQYJ0TML0ICTbRsqfsZJX5qcqc
yw0LOPvmnbplPV9Wr8va5wfHr86wWPNmDzsjkpUuvQYX8CutunbzfVYsCIr9vSx/
SQ7w6cP0EIunzVHLbdYx+8tNpXpHKPi5DHN0qCQWXn8Jff1jtjR+Y1Rnx/5/jjDp
QhGOWiCsVvVpLXWchOE2ClSUNuJ0yGHucCn5zYw7r9GG5n+Y/h820jIUDGqiYdv5
G4F9pEzFUihpqzXuDiEcRdOkc7ea/oooamDUBVKV4Ud65II6XgX/2w5ImV6Br9Fw
WF4f8AMiuy2UiJ22GP2cCuaaNsRvOXSOM4xMyiVbITNY5kgl9/xKQZ6dPbIbA9jP
NjutgdfF+YYzUCu6b8iIxftzNxBh3dSsvky2EXgwCn6fFtKPH9KoziMTbZmB+0hu
tQjX2n3ZIfzInUlL8RRHla1GIae8GMT5CN0Z55uLutFitYOxgEWzKYxzJXLt2JcA
NEIRbQYtKX2taferZU1Zm8PMeauhnBkOVvSSx/mrYWOoeygyFH5Z9UpRiHFAqhl7
nKpqRjSmlfCwRW6klCaAeqIiPnZqbO0evqDTiTxAcvD0hVFTIwU9ZcIOuzTlEkuF
D3k7p2XcooxxyjrluvMQuWlMISFfVWVRfQcUrJ9UHmHN+/dIuN0YVIyoLA4Bx5Am
QN7DqW3zOA8/Srri5L2oQHy2PZSW5bVZiQgNqlEkC7Uiibq8NHgRwzsw2MNU8j/V
+rC11EM0Ew62KCgSwlbu2GPNfEX2GKgAvRPcci4GtFRAzNOSTlKn0Bd7FWvSKxQs
6Is+skuU0Msek3if7/FwpA==
`protect END_PROTECTED
