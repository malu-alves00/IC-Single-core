`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nj7xkpqsQE5zHpuDYuFdSBODqV4ACWMtX1rE1+AYcRk0212ri4bt30sRMwXHibDc
A0HzaxS2yzLXpzvOJfDDSfsrm9XRJ/SJLF8PHjdnLvISvopsuZPr/kp6dB6W47SK
Ep1QwTD+OhnElG5pUu/m0U194++DhCvwNheWs8VZ/MQqSaXCM2I9SqTWR4Y/XBcr
Y4y8x+ymqO5vJnPqLK/x/f3RIo9srNo9ktxubbJTywLKmDmhoYMf+8ERWon9Sw2r
5G4WWfrBndFDYsoHFuq3muhMXdOklC3+BSxmyRngQ5xUvKkKBu5ezJit2+ENQHQS
/9BkXBXM0HPTmRADePfa+N7SEri3cNQFE0nB3lKyy9/VOzQp6GLVeFe7ffEZMa0d
gFKUPZzh7hf7gjwDtVplbStl2t2nqHDNFoxEasFCulOPKX9prKxqNmTGsZ6GggJu
9DAGDwsvCaSd8GoOC3oqvTb8l4NLRmx1/LtbeeUODvxCKBJuQdVZeGmjUW+ZlSci
CjwQjunctFrMTskjx1RvXZKNAh08+ryHLxMFPU5b1k1BfivYorgAM3jm+Y1cloNM
TckY2R93JWt0MI+jAnt4NcVPx2a0YKIXmJXzzRz74kty7OMnqPDVZOthuFOJXE5S
07aw1/zQ1K4BtXrujGq7UmiUXpF+bxn05OjSywS0flgdktrS4t/CUlPEFjPmc921
/KvGztbtjUvsZIh9oks/9/OmFZcWcBYZFagHuu4t9ONoRNWySIUMAByZ50tvC3oy
hbNFaJ+9YIq4JgjHd8Hy3Ghk1equJzGe0OvbQose58jqpboVUzV5zLuo9qiIP5Us
RnpBWKxNgAlQHh7RsrI71J/w2n/v/sHWuQLSi1lssPNih7B8hFjWoUvtcR6aa653
l8U2czBXsOJvUwvkLrUZTJ2QVS+LufQ59LOYxwD1ysfZqBBCjhBEYUe6n+GNjeJz
9M4Pr+JT83jRt4gIU6qCTNZ/OnJmXsJEl7ecyaMK0CH1cZdVZmbzTHGsTr+0NoRq
C4yUisq78hLUS3bB2deQD6Spbp+gYgzIqi5Crk6cY1EAl/sIiGugdVUir7ZuDmZv
vr2PmVum4IiQbOnO11lV6MzahgY++71RN7AdISHEqTR1y+1n3HmO31H4zPIk3PEL
3Ou1LM/Wq1sEV/qzDU8jT2lOjtcKnvSBHhGjQ14BTtNPC/jZXHigHGrpKpT8fa47
VxkkOptDADFLnMJ3bLJw/h8uzLD0JBZoxq5AVstHWhR09agFe/RYcLbOqDXhNAs2
v/L1oaXpSfMYczrXbjoRpXX/8M2I0WxeXdqRzz9wYMlu8I+OPE16QM90SffmWdMf
aYU8WfPuH2HQfYgJTU8ew/FGM/FepeKnYd/Ps5DKlUF5ndl+xxhfFh78tSyeXhTM
uk3w9tGvvRb9zBq4hzN8aPTCBxM896C2TUfForOQ3hD6R/IgohKKwsjTZ+JmwhF3
lt2H9E+tookkLE4evWuHrG9VzZw6xrPrGE2E/m3hJutHBnMG/NY2yT5zFB7Hb3Lb
gyeVEN7elb506l+zQ2rAngDDq9P7rUUPV/7UaBIUjWEZdr5HW8+jsPiyig/OIvyi
4iQRfpp9gk2VD+Y5qXNBKcRijEHQHdSELTm9eXdmVBjoDjasqpuZGb/OkkSXEYqB
RSkkooaG2RAj/9zCuP1AnWFOz6ExhYER9+5uDViq/4AP6QN2dHwMrqJV/IgEeJDv
53MCk5gvD+2t17v+EbPieF4CRMqLJ6IYrSY3r887lg4mnD0npF2APxQynbaYstu+
p8PkVl9Oh6KcT2hy9k6LuQIQeCmEPh/SMxQufPhtk0IxyL4Nio8IB2shkmxezgiC
JwUsHk91MYgTbM/XHD8pleqjgjpqY0uZcDJDqkSEKcxQZXhh/sHSCyFoUem0yHY5
gLnwsl72S7qbDXs3lGTAArQ3Hfkn12q/ZXZFj+ULuKg86jyxrKXLnxxHiAoyRFSl
r5XjfOxHoZ343HKIh596shFUdYrYfGrQRMYxSQksU93KkQin+gCPJk1/2gdmAYur
fPu+FI/nBqGdr9aBc6Neuxic9aYEeqiQ/nu6ADY9AeenR7ZU3Vi4Jz35V9497B3h
Wg3D0cDt/11QA/9ekYlgPkrLe0W7hAy3vZ6ySRn0wH8FIxZwHISLdpBWaVnWnQK9
aw61KPTdmVVs7nH2IizYSNkzwggldh1T0KvHd0A3HZpcvKmo5KNWbSGJU1J6UgAe
goxVHLJVWA337LLj1h9bawsoHt/L7VVj+Tujilbs4jroth6D1cZ+xeT+Ii0GgbHT
o5dHDOc1J/imvBFQCejs/Mf9vGHvj4rsDzQCpwawap1wFi8YYTPyZNglBEiz6WdY
Bn3emseiXnFYux4O1dL2nGyjLDNyy2SB3yIH87cCFcON9C8105hVaUJeWQJrv8A8
syBojBu+g8hSlcHQS053DPJYFmcYMp3faXjG0KD4cT+hyRGnZkMYkAvOU7XGwY+j
eUZQ1DBLkhOtXe3/vzoXBXfRjlb3yE8bf1c2b08HgVfzhhAjuEyB9hgXShGEdKLC
mK+5NIaUjHkVP0C8tboGeh1lUos2gNK5yXIlRuWZyCwnpaqRV39JuVbXREhdqDS5
jAzeLcei9Tv9H0L3Jn8d+Q6LfzywRqEkZmeJxUX15gMqKXx3DuC4AAKSNou3dklr
EKcNTp35VT/04wte1HJ+LwtUQpLOztLADFy2ERIJh90yklFoWlWhkUdFVfAryHTU
5Pxx0Y0K4kl65x3dPlJfPh7bhhYVEmWlriFTBrFdR2TBpfEB3ww+mP1iCulGv/Fn
uyOQRuJWsBMBpjDuikix1XdKzAYHL7J7bz1Q2eyr7sPj1H6RyWnA2O1jcdr6Jh8A
I0hrGzCyx1PdiPFmNPveUmtRRR+PoMliov3/vyIteUoEmqCA12Kou3QLUxcNAlfl
e/x1nUdMxJUMrVZ7uSH620FDD3kHbWbgJqp9rKn/6NW5+9MCAe4waIOGDgrMyOAr
BeQndApYqfgBpNz/Y7TVgw8SDh615VLVdye6PT4yg+q0pwHRa/ubXOXX9MIIKxAw
E8ZXFYyDIE69eUKVn+l8I/d6OTjoXJ4RImIr6mAQHqWRhdR08HBH6SDasoGuP9I2
43HmFuDtyu8VnOBZaSO8a1jL03o+A4vhsgM8iYVv0QXbStDxrjR7mGoZTbyc5ygn
a71d7R78S/dwfYOZqgpgfb/xzJqSggCGCYfaqkx4X5ZWhYdoJrGUIqHD5YOHvjfQ
kNKmY+Wkw8gkLdIODiqOklhu8oe80GmCryDq1/72Nyhl/bkW31s065Okqu1Ns/Xw
E8MWBnHyI4swk/cq7CTT6gIVk99opFrKBdH4QLiVrTQJLK8tSRGWmoH1+v8QTDKN
OChIGs0kUt5+v5UD9qjuNzUOHD4sEQR4p6uR9byGJKCSUW5l2eB089Tehcj238kU
7l9q70A97QEsrbnUNU5qhQqPGF+18nClMDoFqxxeGmakiX2Sa3NNbg2BdkW4wsp8
EqARnrPBx9XAdT0yRzEWJvtMi6hmf8uqdwwduh95ZB69zoi/gr4zzle7A2h3+0Sj
mAwnI9I0MHeHL7ywvtkKhQMtRsoiU0GDt1tJ/N/lqb9MqmTXDBMWO7Lgd0aEp4Lc
80/BNrlcRwsTVCyY+zRCqpmr6/b35R+sD0k1W5DEyW1PNYfe0OziSLt78lXn7I7h
xSu0EWOFYKYXQmomw1CYZlbrNA+Wts0mF7AjBOPq95nJpFzxvj76LI161HP7QfVW
MfgcaeKVEX/6nGEU8OWTMwVxvVGh87GLC+soeO8e14I9RZceTHUtM+0emTBe+1tu
oCjpVSy8Pa7B3NHnPWMt4ZuH66hCU99wpO9PigyGBsLkxOkOR7ymh0t9YD8O/hgt
CCrh3vfSLbqNH7+IN2wugRdZT1MF9SABu84vsVKNXv4tHLRBDClnaodf0bjrJ8WI
uNVEepgyIBTQAYFQE5H++9Ml2mKMmljh+DK4xsq+w0+5ovvm0C5gSM3sea71gnS7
vzjTe8CGrkESLrH249gUsWAK3ngDBfq56E0D4sJkfTI3ukVmp6CNx6Hl888/ICrW
0ZdMrqwFZjbuo8wVNVUpFT18P+Ugw+hEGZeSFvT3GibvlJE9b7wNrf0fQVLHbfC4
RW3Bsanj59R2vc8P/gOj56mcE3ZzX3tpPrKpMftbyUeldm6gCgmaq9WSLSiihRxV
UELzteXcYrQwZQHqZFsJ2xnx6Aj/wAXVljR7IwAhVp/H5ANM9VRxAbq1ZvsLVKgI
cCTNAh06ADPtuwaXdu3st6B0Na+oxPwaN+/ICnPEWQ0I0+ChPNZmLB4hAVKhNA5U
b5pwVhNsZDn8WXBwhjQTAudW5v09FpVu3k8kaJ9KD1Q5VpcQNI/rNCLKj/dTfjku
u9xsq93l8bvAl3DoNsV4eyWurV5Slm/wuXxI3Tt3PkC1pbKDLMNq8U0n53SIJbC/
zfzwUj6eXXOza+240FZ16W61rI9lJRUaVBLTGnRJyH8Bm9lL0un+udKRUqWUj5wb
4ND7O3DyzgFP1EKWalThTeKaS+jviAvRs3ZOOxkj0YXWNTEWW0U1jSDMqU+dcs1T
KSm63NYlWx1DuQb/T+3olrBZAKopJuoU80p3E4WewNWQgXN07UMkvM3giVHoSYzW
EIGDobXM7d8WaDfr4mj0js/6PrQ2O9OuxAjQ8lPRRkXwhWcCGiKqUMLmr1TjaM2Y
1j8GbhScYgED0Hry0FvI6eHmB+MwCDskE4fLp/767Rxl9Iskt7iV6nXM0zJ/yE41
rrLy4zeKnjB0xnZ19oAO3lOPOiGRzziysTJrz03FeMNU4BkqNhoJJOCFMS3wvZy4
gT/zzBYfPDNzdsFRzP1S7z8bYtwNknz1DZcGsrciwQfav7Tdc07zTSAI1GURmHAe
1jmRBBm5l/N/kFV3e4ZvKeczgFHc5IzXKiA1FWlm87Fh0D6BvL0hFkhJcDo27DVW
7PYGnm573V4JifiFJuDrh0tHTC2CEqYAkCGhETYrrNOZy20sjs5qZxMNq3EbVpDA
+3QxlTHvq55BpJN5Z9DkgPLfDHZsEoTQgVgqHgwPDo19P7+pbOEIm3AG3ITkGLhN
0X0QD+N21KMPD5NfeMstDGLBO5ZyPZi5aTo6Yiyer0clVqqHHy+Pc99d5y5W8cEz
a20fTg7fAi8pwobDjYvHZed/45hdof4lHs53zIPRMJ5F6TZWbUFi3BBwKwMRSUEU
mRfUNqfQOwcBXCl24cImqlL+6Lgzbx5B1HuWOpwIlqmlhrDHoYGoAsOYaRS9WgRr
xcb51mKOfmsr7vUhOEEceauIvRxp7CV0Gqc8tfaTBK4AIvx1ZsmBRacAfogBzlSG
nn6/4ZawDk2OJpZ/jPPtj0dJlJgHrIsfyR9LeKs1hx9h40QkseXnNKK7zGty6g+Z
VnAK4iCn0F3FwvkFoZqAA0gDxO/dBVEY6Pp5pY/V1BFSvS6HdxTtNdRWmM513oRw
sqqpdjrC+M8tX2QYdRfSWyRZ1OCgbD2rlm2d7rsIOkNDLZXBTu8Rob0iovQYZGfv
Rq3sJpCfZZw3et2JIEq9s2umah59AGEk4alcGIBJBHsXlJAz+NshZigxzZY82aSz
KgJdvq48/QlRGRqczc00zPGUzNuDyRlxuxPgNxGnH1NEWi7b0eJloGMyDO3Biz5u
wG0PpCdsoofxK2+oRVj/YeztEfONneaIAz2SiF8ym42uAgTnoEOW+MrfVRq8gGNH
cPYy4M6qOq4ewlWwXGBQ9aYK74yxVA6bCOVdEckI9wGuEdZzO+pep1/HEx2Xt0w7
vl4+9h1MqLsdKWgonzcdPjZuWvSMb8mrlb2JEwFXs261XPVPneqasqgebSa32StE
Vhq7jM3EhRbcdEBtebhAmZCdRBzmJ/JuiCRTO4luGizXGbLxZYCkhdMnuMjme2LH
BwsUE8QdSIp9KefoglNtoY7zbsWDE7G4iPgf29kS85sWdYFixLU7RINK+vPPRVJX
iisp+7oDuJS+rM0RkdlJc7ZAZWpDVDWDqwJkGOsErSilDTViwQsJKBpAhPI0RReF
8FXjwPzcSjo/gtVjJLSxCVlWyLfiva2noUxPs2SzBwEDk+nPAmNGdrrAlFKCRmtv
xGpxnhxVt1sjpiwey+FRb6voO4HWtnk4+mgiSmJXcczTYg9BiGJYyy+edyzF90b8
P7l3KdJ0vjnUvWGuJjVCTTfpeB4OP2Lo/5EMTYFEH2AseiStz1AtcNFlIJOm2MK7
dMSQvNj9yEEzl4HRT5x0o6cMVv00oiz7+d+VHE7XUStaT3fZnatbpzCnPyC6kcTq
lE7+9+lfvDGiB5fHbf82fTig/8p1z7ZWlB3C4nCM++Tn72ebCaEN9dqnDMxLPGyS
vuoo4O93U4naOx0Ogsx9opXQihpHPwuSSE3ZkWTAp7asKHvqPFudRbVWLHMJPhBQ
xznaPF4gPLRNY5l3GZAEioUTYz+an7g7yR3WhzMkkOD4bO3H1DThyTdVryB0tsra
Mp381F9Z4zPLG5VRfsV6e6Y7QqkBhjHDXOwQ4ny9fy8PcBc+rOOiSRR5++EpmWIs
5dbjEgdE7KLHZvGMUibCZxDWKwpzD4kqdDlP27lfJOXuXenjEkRBw/XrUdQVrtob
Ddph4bxdIbfAmxQMcWLVAjIoGbesdtkLSUcBmjbawe5WY5MRz6Mx16hKAp+Jx/ow
8VV+fMpDlHlYLgLffm8s3X7Aanm6meL+kVZOWQMpIbUMjoOvYdJ1BAD6pGTMX8eT
bfybaQ5dfWsR4Lf4vZ903dTiFUIdbUQ9184GDkWgfae//PBAzuY2bBsD50qGLFMu
kWEWQFkhREPq6G/oRVpOUteEFiPQjs9rpVc7oQ4QvHTIo29/2fqHiNMCN5fOKjTd
gvoPaZ5upeVQt8gCWUBbzA1L9TLFjqkQ+7aWCrtsY3Z6/yjXABQoekPNz09FiLVW
UiRjsouOtaHurYFlKODLAV962fO5R2d0Xj9TgMOup9MaMV9Ael57iiUVRKijAxdh
o9U4TBfhjEdSvvn8ZtWJB8ren2LCvhdbEaYrELXNu2Y2jNrXw6sTXJr4WsrfI7TE
QCDkXYdPx6WVRyvdpHrkufaoda6BTD4Xjvrzr6XNyFEsIGxLX+xp4iwbV3q7p6Pk
G6GWmDi2fjZjZtVUhZtoM4LD1TNgo0ThkmDk457/n8/DWSWqXWNHrYb8CynHCvbd
Zz/1csM8u944F4iGzFrM+TsQPSfNmakE4Acbu7UI4yF9NI/yk5HM+I/RDD2dDLTY
x5va40QNju0LJTAwULohPfNXOhZdZi1QgWfoZCXgTaAiUX/YC3PIcOb6gRPdwtq5
SNVeQZM5ONnrfZEiV+uAVpnMY3MU0nRCdVIr9TFij9pRz3Ri0xCN+1/BlmchwpOm
FB70y2vv6OlFji72B1cXTVCFmHc94jSqsburQL5LGT6aQE9FwiJ4tzX6ji32KhL/
tZGGaGokI0oQkZtKXY/gxvX63Y1+D0pP3KG45dcSpbGb/GsS5AOIEzlvui7lk/Ve
B+EC7IIOjnMeWUwFhOk1Hmg1zC8whmNFw2Z8C8eco9DxX+evO4I/eM4k+UCKcA4I
OhUBsNMtAqVf2tsuzTgUAkfioNmAZy/ZvECdUsNJl7/y3veCbzlT0AkhH+hBgenY
lhv6KzeX+V3qSIvUCbQ871aVAYtbTKw2LPWDduanFRFFDQ80t5nGUUBcB88vPT6V
0t+HEtPV0dQGqSbW229tpqVjJACHchid0kC8z7SulXclEMPFzRFB1bIclXXXjjbb
bOVv1qiZ+UwIHSOpCps8vNse5riQ9EhYAFEO3lK7eZoFptrIXuMGa6vnMxrgSLPD
fZVHTvYPWwa0ALeWetT+tG3rlFncOCBMY5R1QSMB5F8g68eI2zzAQc4a/JgDsyWE
DxwLhZ/mLleW7m+sF/5E/3rtUV1a/5NyEUMgVPzm19f1KALDm/sFvwwfSorRzTxx
J8ZJgCRS0mOxyGwnrKzBOcDl+w2YeppJZdvGzLTcLAWotGnroYAfUvbudKqxADag
ghVn9owI6EElTsQ6DZy9hmcAzUTf1fIagnbCfxQ5QTVxW8Vp+gmQmohIYnSeiKBv
DZ460a6Jbr6kmWxgiEAo0WlNVu+EiJApi/kssxyIfXo=
`protect END_PROTECTED
