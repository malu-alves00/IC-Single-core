`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ghNNngyaAfysHOlmr4fW7TpIy2yZpYhbeoOHj3xzWn+hOCgw+lpJZWUlJ4e6dIKC
dV6eGeHa6GNV8i9zTRg7oHM8nZ6TfJlZHvTvJtuJ1ecUJk0mD2xSuVihcopaIDsY
gBNBw9XtvuxDBUm2GJG24L2eInVzhwHq6Z7MBblOBfbCDWuRSihiapHJZKOn6DSD
XTTdC+PVt8tm+B0nV1bjOBIlxLiHWjkJFS3Wq1GnCiKgJOGrDLk5Q10muF73tjLO
R+rEpwxem0nDFSRip80FnABaUmKlTFVoPtQEP8f0s2qFyDCzQ93dpzLUIIkkUhH9
7D0TXFHMjgEgnGComNzfp3z10/f1LNjLldAIFPJ6Fd+rvAEkyWYwQLZ+DUerdanp
3QSzMey/88KjPTbrBoQ9eoo6+J7lAT9CxslclT54lkX+zzH/qFowgIO/aTAG/F6A
J/s+btXr1UvLfo3I0YY5h1HYyiyiK48wFdzS4NlW8lmjpbDHUVakTyoDdX5TA9Xi
tMqfu4x6krUSMVEsnIzu/nqaTjkHIG/N6FPJyeRWh8UuQ57Q2JLNRounzPLfOsBg
zrPJ7QOS56WpZ7xM0ou4gSaAVtHyZBb/UsxVhC4fj0d4o6KsxUmUzd3Lm+vVHVJx
ogsIXXrfIOw/HdG19i06ElSayKXmGGlPxVanVVDOBYRydkmnPNMuMZ7L+X71JHBd
INmOYmB/Rkahf92sClA/2E/2c7bvI3FliNLePvZV4XhkHiSAQ+L6+PBJLz0r2B3+
rYK1t622pNlhTe+GX2yAZaMpShV9xhpA4AfeM1Mea57wkbEEc34fqvQ31dRIxj7t
BEcDBxAKLLRFOm26ke3Que9S1mEl7hFhcdy+x4rFP3bjNvLpCFurZhnlOjJgGSx1
M09gJOBYElv4BV8u0WLwAmNiZqVAfddiFfT5G4XPrxlMgvIdypM0NoYWMsxq3GqA
H4QuG7heOZqC4lHCw3VKGxvgn7iE34qW1oWsYh0QNKY13Q9y/YbP8Pf80xyq1jE6
WEXuEaajTqwgW2PdodhZ0W4V1gSEFcNk33Ta5DNndowZHQkNfQ/nOV1aeZB834G2
50Oey8hl7emYnJsHpZMdf66IBmvShnS/cWClGIdEYVQRgW3unucLwNHbdcMIk8qt
6oAr+zJzRkl7yvYFlumHjefcZBpw2EaTbyz4Qe8PuQBw2tAMoMnfClMnTDs7eCNA
1p2xlZrbzCmSQmGUzkViJ3LNV6FFERqSRSwCzDphC/61t/t88DsyvRWyc1Mg/O0T
xW2c/9Xozty9EES5QXHoSI0nr71eCmgEBFoTfWYPMTFMUr9+mD5tOJxnnt7fXS71
iyzqw8zYZHS1KPMEx8WwdlKPLWoGin5XHDl1w2c0sWxW0p7BsprZja+hBfEgixjO
`protect END_PROTECTED
