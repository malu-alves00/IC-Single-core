`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
naJ90WuDDTxIapu3cu18P8M4rb8S2fWxc0OzmoXoAErIGoWIDW9S0i0UXYHkzcEz
9cd867DjoGTL+a3uKzkXR/tQmoZ/RZwiC01ru1aKjVzcZnEadyHtuoihqvBsUkwM
F7ajq13IXhbCkFVsxZBj4y6FGu8beM9sOhm2b4idg7W3k4/gO9Tp5Kux5IMGjvQ5
FbWMhvmrY7zHHtDKvixiwYq8G7RMgJOuyX1NKmnavEmhJrQYRvhCmkTJ+YKnc/Sw
V1LdD34h5m5gNLomlzn3cywGIcw27zbyAKqbwqEd/b1wJbNnabWx+h8pBZ7vLiOm
9GF7xDuCEbXG2ehBY+E7uj2+HATRlx3jBFDe0xJodIIcHK4+fU0BYOZnOrcUN4H1
tjKUtbSHvZDYWzIDkdRCxycL1YzOc2qa3z8N8Oxnn3i4Gx8SsSrK7xt6GI4LVfwz
MbhC3RYjWwLybDYa2kjo93qcwQot1WpFubwU6kNZ6ecA9zhXARtirCGvoGk5hOFd
ujO+ILojcPLBeZ2/SuGFlNgnUdj5sqhXEp0fjgd3lCMJM0GDzIkk2widO9S/VERW
a0xrk+unnKsZ4QoQVFyUqrr0XlHpy+dgUMdb6q55KAAWrtTAJEAInz8CcqXw3S7O
A/WrerW6MiRCakl6HIh8cIWr1N1e7elJfmrCUI6bXSIyjib6a9dn04IS4JL6uuiZ
J5AGx1V5Uf6OrkZmPFkKjVoM14h0n16nAqvhSHiZoSo4mN8Wi8Jaupq/3lvmPx06
OnUhRh/CiU1eOrw90kASEwViKMJHdcdPAqYc4mKhmW1Obluz5JaU94BtC371hsWF
G9atWH+czSKCbmR0SQSBJD9Qi/N90UXkCF9DykVgv33zQX/Em0lJ2GHI1AqDcFbR
Qk2zB5LjhNElQ03nfPnXzCYwcX4d4wTH75J8Uu/VWlsWHzp9HALTNI1MzZBrMGga
8UiQD1sIJM2xu2Il8SujFe/A20nZ0OmF8DeWpGuHf+FjU0Dcm2gR5rKEtpKb7WJH
IfXUeyc78VsPNhF9zByNDrs9gSFRNofJk2bMJzTk/9AT/HYqbYQM2oeeqDYt0gqB
qCJ2GNnRLhnUNGYv9T3K7I144+WTByHgIsAfih39iVPONtZUdPM3SkyMitYlY5bE
2l6fz7B4XGdcatjPnzfUcTl+x/cSQrTCvolHPiTuTfP3ZFxRgcKSkzuW2CHna1w8
kXwgpRAdxNiZxDlr46b+w/MOmU6o0pDsTjFTPEYuxuufqe7guNF70MWHqFhMa42d
0UCaNpmYo4Zh97AakS9DegtLHRurLD6CfKMiTYMdP+OGF3hqbNjVSXqWMjJLV4be
45a2m6j5AuP2+nG1tH9/vn/wNqqrcusRVcLTS1JJn2bXcpYTIhptOZLBRWJ3GJz5
UMElmwZ121NcXvbkcsOqXdhDEbgMdH8FZWhyt7Tk8ZsJdmIhTrDTe9yz7v0OxkfH
FqI7IV2MWmwIdPixvcWyWy2/f6LexBkHwVTduSBqC0ThWQD/rQ6tAF1YOdN7QNFt
1MlSvFHVID3G3NMjkPdDlEIqM5p/eXy9D4u/lI6QNdVk7rke0apqlejlq9KN8ez4
lGNTGXnQGZ81YB35Va4PrCuJLdahU1DbeSNQzhWUfRJWnHJwyVmTTM2EnwYUXCoc
zhuThYXG4Vs05Wn4f8pbQWlL0bAlgBiLbae8DqFEkbRQBIqauPsEbcuf8gPQMpw/
30NZGeXEx0Lql8/7uY/bc8lM72rufz+BsgbBzHGjiJ6jta6C1LKC6lSD4ElHb0Ng
c431dUjyQtaxW0dTbEZbA/MfN3R+vnt2PmnSeWE5Ciud3/RjHDBTGPPRmZq1MeK9
rpyg+2gnS1jzJsyHDd6aXw0h65R4vdk5vjVAI7UVCDrOoAYFBKFipu9UUQeYXRAF
wx2Wa9rkRR0QralS5o7u/pTaETP/Uuq+X2eteFZK2kCPlEQAKqbstAOHFIqCrwnO
Zc2U0kFGZopBVxFKZr1w9O/v9g/AEBlC/62tnxfk/qcIy4gp6NQ8ypHF2fuUsKMJ
hqsPGNs9TgsOXgXeInaFyKUzVRjY2nT9Ah/VnjiVuJoqMGX7wnZTxHBzriMTLrsW
x3odGTe91A/0+Q5HEBEe6qNw0FtdUzeeEkG1oNZ+ZR2lXaUzFAlmVfB2uaM7BZK4
NgkFghfxj6BzViq299owN+6Itfm4O2200L8Md16uBiC4zuPAPS5oTT3ixja/PzL4
87iLQGwAb/HKcw5yGWMfdl1iKXrzET4eHzOouio7G0v2kW39F2gLHqi2QZYH2Z39
A31sSQjbTOc71mRFfbzoa5Sxr7pla+4vF3jHRxgFMcdk1isVe8Dx3ycWtI0siRPV
nZIuovne7T6fRxMAHC0ZcFGc6KEnRsU/J2fieROrzV/213cxmaR2dYFBhT0Mic2p
GMO6cSwknLUN8Gl7z/kei/iSeTuIl6ik6SVUqh/vTZN1ObMF8OlYQ9NbvpsHbSio
oid1/J0MR1X3OtVAD84YvHE71YuNZRfHMQiRT5rHTQiwN6kR167Omd3aucnjYpp4
gxlbZOsQvgDTb5iOtWGK7en+hfT7Yzf5gWug5lCYw/uQTUXTZ/il8XsiCfNpNsId
ubmd+B3xOAdUtY6HUwWwp3gfvF2gx5sdRRffsAmR1yLo6TX5t/xubFBn6ejS/VaS
YZmQtqpNw6ExnlEaKoAbgoY6CQC3fHglfGFET7gqYOCdpn8jeFQRhjt+d/hOXM7C
CJ1mFCv9bx4No9iE5ByIFPghnlpNH7JdR1TpuADmyqKs8eFFj0NHn4E3W8I9e7ka
ewNmiF2wqp/uFplnG35Z4HfrbkuuJSBAbXDdWO+4SQ06Byj7EVRgSKlSK0L8lMnX
u0PnHWiJP9wtg8F+vM4BZQM3580VaQ3lMD3BO0nNxDd0M0cDdtAsgY3oliRjjwXo
pXdxmZA421EHgW0BnI8Id9h22HruylafG9eHv/klQH4Hvr7O2HT79MCChZqa6Vrd
AVVK/I8X/7WavGJpPS1/Wz2jLrXQbJcQPAiLL/J+b2Lz/tU40nOcIjCHxPf1b4LY
TaDOePo3gmnZEbcFXwC4KSyxh6T2PkWtbHi9to/GYnagOTLGH3AkmccwNRmmjO5j
dOo0bGZHqjaxznX9QQOaBSpvLXuXrmm/n/OJ1UzNI6CCpLzN4vmmjRg8i8f42S9o
JaAbnue7NyMg8KF01H+eYBK///ahqgTcfCI1wiD1IIIQIlAZZNtq2j1mb35b+/0w
fIvqe6fVBOv70NejPq1fWxW8uJSdqHxisMSBB5BSCyVbRWPhclTUruta4o7Twd/b
lcLZqPX4BBcuTfMO58IUaMpjsCmvIymVuaane5AYfku5oklg/hTE5saTFmbPrgsz
pwv43iTQ2ef3Rj5aJA9aVbDGoN95/C6FvsK80hAu57ad8zB4yQ/pm2mjNhuaB78a
sy26i2KmzTRbjI7fcJ4PLsiHGkHYiG8b5t/ngg9LPYnihoni7flXy11unwS9kx3o
AvsntbaL22nHpOUZkaNt0LWvHyxObz/JLYn5ZM6EOICBUcwrDC2geKkm7KEhgac0
lmSbw8uGjGm3CinVOGUj+zmiS41AImni9O3RILX0CVAWQ0uC5sLrJDw4cNXOkZyi
v18Wv2WwMOtTqCS/jDsHg2J+12vx8YEpfJ/XzCKgljJf2gowJwMUAiuusegeOWn1
0yxi4v2nuBy+nacKicgrl/TFNPQ9hyLe8feEI/eP4SWgs+q9G0s7ElEje2y8g+Lh
VMEt58VC+J+mKpAu1sSwVa7C/wzodUQvmLcqlsX+pYeCLyP6cnNFl8OkzchuvVLW
VQPF6U6hzbk7h/yrtAYrceaynA1ICIUkLKcR270g0sFjg3t4w95ZWlRcoX8HjLd6
IaqxD8wB/5s7+9uR6q7NLiIV0Sn0CsMNqkyTZElTwULG2bFDpeargABThMVLIz7A
NYsKMVrvCvNz79M3lUrwyDMMHsb+erwW4Cy4oE8JJzMb9zTmklxQv6SHoaCkdxnP
3rKyVBbWhhOMrlpZr/XgAZzw+sSLCiUoJt4p1lSK9PCnjKVtliLKedkOKJIwQAEI
xJBexvyp/dNCBDX3VB+mzdvffeyi6FPaQ735S+QVYGtvDuRjUW9tCKrjZysSgQBT
BXz/IMLFnLpDJJlxNoBCIac3PYitYh4kZg1wH3z3qkeHgzf8Un/TjkCfmfNOLcxv
ZZA1lJ8qLLktyUtJP3dSMMUA1BGit4jknP9xVIHmBsDMayGzUiQM2hl8mr0kfWw5
HasetpzsK6MyRluwFycjJvq107v/uvsaacJ96KA5DOZlRNM7mqfXO57xP6hjjfho
3pBPAOLNbljpmpI2hbBmQBx2ZoHtLhXzWozLd1V9CVR42zY0H3WbPBHmRN/XyCF6
mYxGBLMAEC3Qvt4+I91Sovw2rEtJ3qGPGAlcN6oqB6dUzIIMDLz7p0xniXgJy88A
EZH9jPDVFCbbOpXI8BYru0O+q3VUF6rVpJRL7Q+9k5lQ/qK45Q4xPUUfVVx9KTk5
hCwQ5/OyvzMpeYTCdHXzFTythe//M82ZeuOQbnY+Mf4/FnRrVtDcZoHqBw9DmYeo
hSis68l7kzcvqpzwVgt2CFo05DMvK4QZmEyPbyo25E3Ix+m4ZQ3tqA2KnaZG4lzd
2YtOSMyGM2ItgpJoOAbddoYAR5p+2HeMplB0yxVJsuMgq0x+xYB2nvVlaPGgBjBz
tvzW5K8VmadrXDRLUFZynTdqmyxPfTwLJpOX9/6L4be12ve5slDssL3iu1kxznOl
2wx32bkGMIdHjxm4iFTUI6Lx20ztzvTUxbD5MM3xMEwzzwvzifAX8wJIVrkf8WFK
r41PqU2mquA6qvMn6lzbl9jlFv0vjR4WJI480KMt4YwwX6Jx8sBOh43Gbjw7N3d2
TDc1d2Yw9aSwZzZJd7YVEzrp7sP3Zs7rtFGK81Y4WJXUNWaZ1hI2HwuOiHU9Pb69
+Ilt7HMqiuRjQ7FLXjaNuFDUzo864nEQ0nGXfG/3g6peROMZAG2l2mjclhr7k0JU
U6Q4RXZb9WwDSJ7ejMen7Q==
`protect END_PROTECTED
