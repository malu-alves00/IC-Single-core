`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2u9Rqw++RDMEc/4TNbXY6npUsRgC/ybEdxemP69jaEcMgY7E05Q94CHB++K3mYlf
4K5SPajP76NVX/mjMdU1/PNPYkHXJXSmq7IkCw2niDryntY1zcqE9xMh9memi5QI
oGF7HXSCz2tUwcIXWIvnN1WIFjiE0t9eU2rGOp+u5EK2zkS7MsxQsOpRmclyVq7D
74D8DZ+1aF+66D6VfK9Wm4UjJq2XzhB0mur6UG9rKSokzRS9t7mfq8z9O32N/PSW
c9eSdlpFl+VmKGO0ZdXMMYvdraUNmIjzImmFCsiG7BgDTgJ8v6M2DpDVZ72x7dua
l8tG2D8irwFTpiLtOQrHLmZkaAe7nbzbZyio9mhIVdT1oV6d8LT22l3Xh1t+ilK/
1PoTr1gm5iBbgWgd/xwq6eigJF7In3OPllePUSiPkaZ7dNVtjYwuvXV+qdX4EwpN
XKzqePnRPRMt6fltCGi+yWV/sPuFXeEZkeIgNHzkRNRMerZXEsSBmThgnzvqqZFI
5KJWY08st5ZnC/3/NkAv+p16nutdJScsrcGJuZ/CWjBsOURI7qzV2pIKmMjEcJAo
b3zr08PxnoX2ueuiEbGDNYasp/YQMt71Vl4D2meU080zOSBTN5af9KXUeDIskQ5V
SapbQeEQM/8HTR1qgb6JfC4XputjWtJZqU2ixj8fIbTXwjCnKiHU7xf+H4JD/m4L
c7dhDV7bdO9gJ+45arvM+4aYWXVgK4tkEqYMblnsloHUtlm2CK7AAwhcUZ8JwivV
Kjg+xDjZeNKApYxUyS/z1cpD9gsWQnmCsUPwZzo9lPeKT05OZAyej0NtpqfrcWXN
7Dal2pHJPmkpKjoL57Fdm7p21PaUPRyb6eNp7p62of1zQj0UWCyJwrrDOWX0unsC
4FxYMCtOGcxzMLkUMeNvglEGXHND6xmctH04EZV/d1cEiNrVbxyC8YA5Xc4FMQZ6
aWIbN0NbXY9tZeR8tdXPuxvX618jmVIDrUlHDnbaQTEfyOrNXCHFjpMXhkCeVLsY
rVlBbHnR+X0ulS/KIS/ZlOa2xIEH8Pm3zQq1maTBv91/c3sMderZaivMVyzynXcj
IcAex7qQCf9DZ3ImJbE7y/S+8e1hc5z9UFwyIq+ZD9rEM/1ZAkjXUzc6Iyj2FiDn
xjeXwggSs6X2aOiFFUxjFSpgofuWrbGCKZdptt/K0HFZBL2vGQWpaoRp0IX17yhI
QT79/K0NLsHrDiH9l3dXeogtyIzhF+WfR49fOCg1p8S56yZaCl0HtrcktmdICqgv
w9xwZt6ARau/6Q3yfg15ag4rIFyAbs7poQr/0Dr9VtZmZSp1bdze+jw+/XQfjNJ7
kc6MR58QGbRbvsQoZ1zljQ==
`protect END_PROTECTED
