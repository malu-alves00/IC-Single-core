`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8zM50zlWRX35R6D8XEi2y79IkMEFqr8BXrl055HW+0NlaZ09Mo3X66pljKtff3IH
96Mg/tNqsgzuNzI7vCt0g7C05dkUEstmc6L/fJMgSbowfYPYbxnZNquyvhmPHPVn
jWBidEgNXFOXwlkCoXcSO7MT+quZdods12I3Wq3GPQjz3MJ73ZitbuUSWNGWhT7/
D7JYAZNK4kCjL63aEQgu9RH29EjHF9EndVROMG/WZeM4VWpcQrIbSnEKzKZGTFzX
mL+7R380UU0gwIbspParHl1CxhTX8PtYB7qbyF/QkoJd4N4dg7DgHTDQzUHg1tln
BVstRKA3LGxlo+/aP4wsYcJ19XiSsWEMxZv1zz2ixHwSpHiq2/sCiQ5SvsfN8bZO
7CXaBJ8z/kuSRcjpuVrxgvI9uDbKkabIm0HoJKUvlJ6gMaRb8JYY1D7dEgRecRDs
aB41PM5Ei4IS6tTFu0eHrLBnSk3IN+mdDiI9EJ6hLZUtF3DYFPa6n3FCNxJHJTSP
FTOQyOWBJVmszBHWiuls8DpoMEq7pcT6nuxe+4lnuGmYEGy4V5YzSK486Ef8lwy8
/giHamxF2xiYM36EoiiXMwg/HlPPdrIeIsBJmGhrx3Pxa7XO5H1/RrkokOk1Y5uf
k9o/p2aH23dcrnoIOB5t1QyIVwifnbE8FqHvEBmLDXCMAHZFMHkwwVpYHoUTaTn+
SuVlYDUl4cTSYJOk99eUL9dUyFBqTKLmTN6W9bwRMsX5QmihsdjZ+KZYM3QzQ6iv
ktp8+pqGRiDKOOsVmDklmnNxIBNYcOIrgFI6MSlzOdtw0+QevKg57xUqVbGlEbpe
xO90UUoRpC5WX9b8O4V06RzknIAESWm0PRfUMqRXP5ELOsqBUL3edi6wP54IMULz
T8P2qEn8fiVCywwLwOeifehFi2X1tomBqQnC/b9fQMlHpNTZxMk45MUkaxlMiN6w
Y5VyxJ+x8ACd3B94JdKRpBmrFP7SF5ScxNA7RChQniI1s+Ihvu+F9+A5Wi75owiV
Xv/DQrs9WWCzVnw6nD46JJNjrtGECfTiZ/P/3SgGP1L1UX5NDCegUNTVRl424eWs
M63OHJZHLOjD/udnPnbkVFv0VBfM4NW+gsPqZCQ344FIRlQ1PEM5baX9CvSOZhqR
6C2dttjtqM1miowtOlkd98g16rIWydP01DCdkeWv6i7rIeiYxoAVIi7b3M8BE6wJ
gpEuJdBHKJHzP6iBWKus2JTdYuOn0o2IXVes2gT9zRnPqGQzwAqEKZq6lGcHrwO7
U3SrZLMS33KCZJe06IpKhFmVB9vILB64IGAc0vuPOgHOBcZG8SDYrLLG2x5r40cS
Y20pbOqzy+mzGAjhwZVmWQsDuJSV1RC+ezeKJQyolLQBptHcPVBwIF50+ZHrGWTT
nSb+qf0LPR909VC8+BUUUJx7snRekYywgicfPPVD5R9/c2lMjCnchP8GIqkNUOTy
Ub4liGo+fLfofEtUvHIsnMLPL52zGt7Jo6TIMtJF5uG+6vIBkDwNIBi1jXGSeTuJ
4Aq9u22GeA0A4x+jM8NjH2wcwT/8hZIX0unbSVVXuGwWLl5OKP8DQ2iknWEd5APT
XNFI9b6RyTv4aGJl9/QAX8S0GoCI+zXgJe/kX8YILMdyG+2hQUC8XyvNQduNWCUX
57jNS/L8pLFGjWG30AMXrzQzrDkizHVn6Z/6KtUhaAj32Pvb5Nd5GOsOFCuUME7p
PLKG8N7s64bK9qe9cJckj7HvIE9VWi750RWGI6rEpAp13+NjPdBDU7uzKFEJKDsT
4bfijCebuho0HetXvk3t83ISsQnEQVmNDIodtpL4wdnuwd8j6vZri3esIEoQkbQQ
VYT7MZwsuL15/VAr/Zk7yOFKB/abNxOI/OgPgmCh2kFGMNkTUgguoB/oo621PkXy
2/eUIyNb7q6yDWulN48TuQ==
`protect END_PROTECTED
