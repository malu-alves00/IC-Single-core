`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Y73t1WnUzVd0HShymjiTqdSr1w/WzhJibMlN3x3WAOoPzE+3MXgVRuyImA+t3reu
cRXCj5UlKg9CKnjIb4MsY/sYETlcaTU5M0/AfDrnAP5NlDCz1CZL0ySo9vEfnq/D
JxXOGVUDtYlLsBVxlmaThFftb/NrXoqd07QrkaRvSeLNfA1XBs7R/prmGx1OlvQ/
9HpupqqP1trUZ//V8V8JRho0DJtmzMuBd0g64S2vylHZQ0V0S/4mumfkpXc1hlsX
qELdVj40YhGGJG+eS1CGGYOTc1dmKaYu0T5wl5aCYQPPrUG8XAiT6qeUtoIRyhTB
rNTZWoc9dcthwMw+Gq5FQtNAkXeWjJteGIqq1u3/V7JKBM2tI1Rcs/GVsIAqGTN8
ChZhFdctkygokGB6HrzQiEbAHRre046lH0mRXfZDZZIxPi1D1qiPRFyFXdqSv1ky
yTp5w998r1rx2om1M+TrBVL7dcSCoyGRu2lnreZ35XfhNb6nhGzt6kg8LnNsd38N
YdintEfBqYYnAjbNJ4jiHQ9fQTfNcEdnFOsjnxry8eIuy23HXjvaro13N+Pa5iej
J7Yf/z/T9HvbEK04q7JFMRjLZZad7UQlyH50yPm5Fs8xoFb/bg/gLlpiFjcxTw8U
EK+aRSLMDJCm66R8NQmpudH1DZoqt5IXrRD6vbwgE1+AsV0DYhaV9XmAmtw4I5cx
duMpleCUHcUwFs24eBxGH8FletXQaeud3r7ONq2aVk2+v+vlXSXaBzOZSZLMldx+
c7ROX9Etp9oavPk/7ZOONmry+fYzgmsSyAKA8J72HbD79s+brK8pByGAiLr+0vvx
dDr5OIgvHzCfvHDdBo77t2T3U0iPFzndH63tUHwxChrfjU6O8xpjvwvFvJRfCUCU
isfcicyeesibUq7OjVhaDX+0jGbJio9HzcmwtGXb+QYsIK8chQ140kwrY2B5bN25
rlTMe8MnbnyuJOGJ9907l5Q4fia1caBhv/utQ0uxDtj2enPNbuBAA4GtgbnJ7DgM
x+CbFnl7yyhjj03BxIy3XZdLk6q+4pWJAFo6gZJvDOTW06dqjgB6HVIPu2F/hwj5
ht5FwPx2+MPtEVydUFkZdgY3PZrxc/iwXcYMw5sOx9RVP+WCLUCopjV4tnsAPmJM
DkAWttbE/SGg7lfmwWwKJinc00QuBCWL+bB3OocJgo4I2dIRJ+JdU8XX56s6aXt0
SzKzyBWlYLoWAWflFfMdY9mCRN519I4AgfnygouPIpZMdvLngXJFuONwmIWDCg5p
p70eNj5koZ2cT3T2XY34Z35Mc+L3N393WJiqh5HP9XyX1ktJfI6ejkqBLkcBzuqp
mPl8OK7Nqso3NRPJIPd527t0rfCgRqfxVG3462Rtw7LoP6XxCNkRNs+9DIDpK75G
vBjGbmiDkh5OPyuako305QjO/OplLQOab+M7JYaj/QiEUKOpMdBZMMrGdxInEXk4
PunjNTgxT8vX8saNdurLsWmyeRab15m6+TFnvMwIHEmGdSbByT8kSK6lcVFPDW77
w41GuQCKAGLdXPbkS1/DrOyqjtC6ou/RJXilOU4tmun6oUzEJEVnPhXNi6XpzZ9+
9RQyvmZvvWklzqcbxhLDTyW521mbmGLNx4UIZUBIIqnMU/qul8Gg8UybU8o2DJpy
grNvAHLQW/XYH7KiGroRqSPowgbUmcH4xGQbSFm5+OhYno+2LT67LFee2yr1VWJP
lnXq0+W78QjyfScJjGk/HOnnG8iINm2OWoWGRYPPhkule77hArciiuhPB1OuqcdH
ljRbBZK5bRdjc/6BxaNaw2GQ5tKsr3hWWyfX6o4JJp95Cx0sNWn8MJo3PoKM5Xev
A1UV/IBz7nPU/9wL0whKwEVnAKsnTazF3Al56TwKvqRSIEL75nEc/I+7zTTfwvTl
ceUriNcn3TKY9GqUYlaGCEqUHbN16G/6X91LaghycR+yLGeV9sTfM8aXZiD7/69c
0GPbduHKHB7snlYOzMZ9U6CfC0SvLJ70JSjAnoJm6r7/4ubJzWsNB8SgCiBoHhc8
d+04cTzuWfmUvKq3zNmri1srb/gEe+tSQJlanLMQItnIcIdHFENy9o+b9rp+eB1p
XVHs5SWh5JG1i3a2OXczH/g5RU7p1Hs5Q9k0bSe/3CKFZIk73kHx2Izqx9o1Zogu
rROoro2154IKu0/P6iMZLtM3L535byQ5i+fjQHtElZ3xvYne4MmUaGb63746mdv8
HKGAWLzIszr2gAHT2yVljsphH0HVe2WUbavBRBP5Rhna4Sk9qcdQh792dGN956Fa
nhFwcHOIUQG10rK3X9s0lsQxA78COUOTu4gDenFig2YpA0/pQwjnl4KNeKflTqNq
6A1/oJ/tlD3G3B3D6zS0Iss0UkzNt5IsiYAXRmM0iTC1fefezk8P0cpLGJczig/5
mOKfl2kJ+NhOevJt9N+WrvTJY4gTIVDnrBOIERdYVK+ccul6f9dozfaWx7BlRUZ7
g6rv9w40W/L2nCVlCGfwjOYTKvUxYzJ5OzaKs0D2GPRuCcBhJtss/tjhBJkgMS1m
rji27DAccZ6ks+g5uX1VguX2Q8TCJB+LMbVYRWp093D30ykp/cBQOwQdV3bE6n4g
i9lpLsNhYM8LThYK4Kh1gLPRt65kUamHThA3es9kRPtl6JF4NjPbYfD2Ys6tRLxR
/X+Foa1pv+hYKTxe5tjILmdF7afpI2jriQ7QHQeyWSsRMfp4bR//JQcFrE9hOmaq
FW8QjwySzYog3hXds/6ZsKL9+5jza81yrwPq2bzyc7fXKIf5ODf4NFVQo0EfXaFX
WBlbh3/46NbY4HhpabvkYAa0nU2h/yRpGhulEdudb1mz0peAEMvnPC/F+JhjF54F
Uta6UzOb6GkgvpWDq23BEkJfOFgVrPnN22kfZp+NY1LNPRawUrFxs8lz5y+3BOxY
TkAddBfRuFy6O75ZkVZ4EK94lU93KTz5aWYB9IC2XCbB0kZ2jspG1NJKKORxBh+R
q2yHUz/v9NFESOp73fCYYCo30zkgqV9l2RH/SBeLRk84mAWFLIzCwvUJX46oyJPk
s1Oj5U3CdNxSkfV/etW9pyqlcBToLsa73fWOHXua9O8ruNylOpAotZf6TJA5O8Fx
ePKHkdX4JiLEO+/UDKTk75IVpBOD3oezlF65ZMLHpuy76VH4WmtgZZss12kKfrSQ
FV7h3ZFPbr/EE9i/KGtAUNV1DlA3werATfxvi9GdIEGd2JXcNYbk74xel/St5szi
+riD/SBDgj1RjW7s20ldkTNqyT9uUiZpGexCrR4iBaRIb0PrQSUfvoM3NL8sZF1b
kUsRDL6YroZZMP5ePjgNT0kw0axbktm7S3UpETYOMJYMuxa/jKowizoWB0Prwgb2
XTUYbzB4/1zB21UfN4XyLgB12ItLXOoAiKK3Xehnh8u7BeE8t6Yh0WT5BQrlqj3y
5XI1XkQn5lL4EOWbDI5VLA==
`protect END_PROTECTED
