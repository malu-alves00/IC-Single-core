`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jTgHPEOxB8+PKczL2Tb9vSYm8hOPw4UjOiufJA+ZqnWl5HrjCkfiW9+rgUO89KgF
W5qgSS8HnQ5FrNb6dNa8V8lBSf9vwO+zRiWmwFrFo1JWVJUPGWvIPq1KWXkP7Bla
MyQh2or+lDOg0f9p63UnksSNQwv/EBNsCv62TvMPrbbDWC6dI6ZNR2Ft+TB1Ymor
AzuBY/im1LQE7B1j42bUYAjKEL8Evt3GTbjXmsEtdIcnLCsCrns3zgYnq86rtTvc
vFb+cTUy5Om2rKye8cJVdQku2EgfKtlZoxrhpu3JhEdhQ/CoXc3kogv08JZSU+Q7
vXifYYtLqHTP/Op18XsA3p0dt00kwwmQjHMOUnGCHW2BCi4HhlrEUnXuMtfTBBBx
/t8CW0WZB+efFK/nXgLF5tRKic8lbdKkqGQyKb2vDfuFf7XGYtKw4WKscyb6MYfC
waU1YI3W8WLd6h44HkKz9VxcURsqiZrweNoafczYkfuc8NyU5HEDwgVm24YtHU72
+xcDuFG+WDENuJFmhjUmf0OJu3QgRMfFKAmNH4O/K3XRI9lYtst1YThsDKaRInhd
jWWqEc39ms+CUjTPXccMWXAgrtb5ywYaNCBovaIqJEA0mKaWU7Fw2LDZKqiUV6jt
+tegyvANHL349gIf3GW8hdxXe+z+aXDh6q/bX/VAZLvb1n8hokNKz8AJ440Nucds
Cr1CDS2nBiZ04di/wjhcrmYXrn5nHu7kpzR+k0Uw4Ugser0gKGbwzpAqL6gjHLhp
gHaxYKDnPFza8x3YJYVAY/Y4p2Pxls/5Qm+IijTfLIHMq35Rg9Tfxgl85fTSKpct
zS31bdUTMuGkFMZhtEopv3uXNaa1LgIkprDy1XT+DA9+I+2L0T1ABXia3yOjJqmQ
vjhwFhqE/xeFU6zL5xXAlw3Dx7Q06/VWEnrdRAY9UxQaFx8rQhZSihZx2KG0T+YD
/CN1f7IhowljatRr2a8Jgb/qq4S/WogC4QCVUABKUdTFvZLXON/IJh1V9jzFHWzG
RuPkRB9ai5EEvlrAzRWb43RgARdPbXKkYEuUOYtsVKjowzIzZqhiomrKu8kFT0dr
dtbLT/n26N4GV46wqVtKcnz4W+cikphUEXikCEP1ytlv+cIJs7rbj1lQqwZl5i22
Al2Dd2kFA6g71htvOr7TTqH7Afn9TSFk+7wd8fvpRwPUvFXU6kDv7SfC727E9fgB
Nk4BYdXpgICmvbCaehDKwv3Em3UnOK/xdozS/9oiDfQCMo8ToCeGVMBnMnoEgLBx
ElwPuI8GNf/uuvWQeeTYMhT1ugvYRnqr2nNyYj4yjR9oZlzUrhgqjTG3OaIipF4w
p0rxWwmy4n99nuCm91Xo7y6zBqzYqsFEdRFDME6yHLMBvJmDqO+MlkpD0KlKiixS
n/hHsW+xvo5bpuQ6ojaU+1LVnrQQgS95j4Sj2XrawYkeQjQEkrtL5cEm0XG4pNQL
zXTDh7y3mBE+irmQ40cqSPMyifY0yuSxLe3L7PEh2pp02eZsyU/0b64alX+7DZbH
kM/28JYfugQOpMV1Y+oBhrK9u8hqQRklpcFrAYoYMKdEiuR3oQ95FtvrulnvN+WZ
hv9SQmo2BW5EigY1yN7b+qFghF4wbVvGmAExcRZAn1Ajb1UlWgcVtfzd4TvnpYpP
`protect END_PROTECTED
