`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
khRlJqksK3UU7lKQQk+OaQeOGDAxejFOXc75DJPoEuUO0ijUFYGDbnaONlSKiKCM
tXM3MaPMotBNMLbQyRnfFyAcvzGKVXClhBy4bVqjsLljZXYurM/q8oIgkVf/EsK4
n8zlmgOiP2AqMKx7jo/d4VfYLcwog/QQV5/x2MgmtnRgJpGEBPpGYuic603Tt2qe
xhN+GeoE45bj0O3ywm4IuNb1jrth35t3i27IshmBl7RGWE9WoWnItei1mcSLjM1w
38iTJ4HYrpOCxQcjyF8xC9bHgM5Aejm0oGdzXifj8/Om4x2HN0ZVxeeQFUDLepA2
UHjinOA0+5T0PcbXjo0TBGGQZ0js07+5Sl2w+uC8cuWxLxK+KotRkrHpIoal1ApS
oPxx7tcvpaAns8lJ6KCDL292KAJbR9+MTX3rogUh7CCnJus/kmmiU90/0n2tpH1c
9ygTzTxlUgddLHQUfUNwK4zVk5aF1DYM+bc2F8ZahhNDpc+A96U2j5v/OrlhTmiH
xNJujeUNhJJm5RAtI+BZ5A6SghdczkBhmQ4/+fJixiqjTHqSxW5p9gEYGzoTyb1S
EodouuiqjTi8SgDKyD5n3Pg1M6+uHGHHJW87NsePRPWqNWlMd0PQ2D9e/s5AZljE
GZuoH2zPFgazg6n18bpW043EwzcknxdCDHCsRIy2NYaI7k5XFLSovbM25FnIWxu/
1e2rMnH2btZeFwPRBP9/YNRUDFfpRoa7nfIHAWcKA8teeh87dWGqwMNuBHeeBgFr
F8s4qW91uvc6mbNL/DK8YlH9KsqSPIO96ReWAKnDRjqtho4c47/GrJK+H3PfBtpe
Co3lF8LFQ8dEmYqzyY1nqqlE0uBVxqyKkp2NCYgqvglnH9wmxi1PdMy5lGsYUdNz
lBW/7+NrdXcGokMGK8PrvNunRuptVvmXa/tvDYkx83yOPsSw/RBye1ymC84ZhCUR
jlKxZuNahSld1rNvhYaoTJPl2ViHzKmo37tenhUvkCuLazlXRp5N1YRYrufTNBTL
UrwiGMGwcBgU1zPNKntv9jQZ6dtWxZmZa3STNt3j3LCoMzFJY9F/tWj9DDQUhbSK
nz37dzz3MPw1q+zQPNPVFHZ+R836Hqx1wmGP8wWlFTY4GpaZSdSixzx5spAmbJ/1
HGloD5lAqhIBCVteSwUTR/4JNhVEKTCnYeVmEvxjfwBlhvY1/Qb8VICzoyrvHs2U
/CHxMLBbQFzHg855nK4HKXRPCcwvJHcEN5BKx38XIvJh9Numk6EEG5UXeKPstenZ
mcYCtmK1EqEJzY2E0vICBgdasyRFM+w/+dhjPTKFS3AgmyEHT5vg29u+8TOyoEz1
w2336Fllirx7jBtu3ginBe0YjbTcSicNpsdYY7QZDq0=
`protect END_PROTECTED
