`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mE+Ftr8eoH/Oe1k2m05XaA5Kmf9HGoYQnw0pV6LN8C9JGpJ0g2QoPhPiRwutlr8T
vd/P52u5/HrQkfhC7vML9Sp0fHo7/bZvoLWFX3wnph1Z+TMsFCfnW7gJDcki2Ice
8PZubxgaYmorG1ZfWt/tKnAV+u2h120H47KGoIIQOK2f8qMz13hgdRVXVtOV4gdI
yh9FrHvwKuY0ElVGX/UrERl4IY1CsAjU5qhWH6dxUwnjtWvlsdQXc6+f1uD4t24Y
GzXh9vMlFgvWKdiJ63AmBhkXc0sHj+NqXwLLuxcVcbGGgMAftTSVS9D6bgShewX9
o7gyaRIwTqNG8FeGEzmFeY029OgwzOVeYQ2S3zous3WYZF3EymdBncfUtB0hsiqg
XkziH8Uoy9quS/qaaVyfyIoDvb5FWIZwg5ywwKMqlhqF+qVfJickorKSGl41Y+4e
ge6j/Bet9JxL4XzMmmc+Pbm9Jo0Q+iQPA4xJ3iY6aP7KkKDBKd/3eAkMTE+rl634
Y86m4EUJJCI60UUN0ZwZJYzHFwsprPUpGxcUTxwhb4U2VC4rSDB+cztBfP+5YhPK
Gxwiva6ez7texJBJTAvLBsuvJf5u8c/iljCzXBpFtPy+j6X2DYGM6TrKn/k1p3Qz
7UPHxEhND1fgUG4q54BVaCBzjtUfS+gDKhnX5LZQoZ/oBU/U4mDeKLS7LSSjM9LL
viY7wcsJ0wJOfYkhWvi/tW9hx+bB5OjOXGZcbRstPSlWBHfZYNEOML4SnH+0mUP+
qJwauNH17swZvINkBqEwXQ==
`protect END_PROTECTED
