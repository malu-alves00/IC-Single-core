`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FQBJ+kfAobi0ZUM3IBV50wEfjkrjCuUUZkkXhsEWDgHta0VuRiHSnl8pRl/6Ggmj
ARSzwK8v9FMXidy8VKL1j4ZogOVMEs1PxXkM9bR5yuCrR58+8o5UtMtAizuJYGiF
QOJgJaL4bE64eqpf+aoQTycF/bbrOu1GSvNDUfcBQKkR7NK1n4Nk3b+T/CoqlbxZ
qB0HoxUBXtxSGKYDqkbCSh+egub9/k6KB3qfy0/9HqCpcTWH5uEXoVwdeRW6EiEP
lD1r673/RaRYjXD/gSxb5rQeEd+JWkBaRQ11LfN5EoPoLJH+B5ujfwCTFo6NWQpD
XId5P4PTNHdGGjxEk3TRyQPL/2EoJVaX8uUP55v7HlDqCVBxZLuPhjFZJmDug9/a
PkVfvjxt7S/hkqC2FdOYPJ2UsH4LEJdHatAQ0dopiNNuaZodjaqxERdTpTSnkgmc
neOLMUcHq9xV4RdVT+C1CFHVR88U0T1g70xu0uBZgu73z6hIIRFKgqbnihshSvbQ
ok6uTrZDT7NkZ64rVVy+chr0NoLNHRYiKlDPYpfn986YQliQYiq+OyiqhnjVpOgB
0RSiMcAgQ1kAwdjg3QGtBTiPH229J0/eE4H6fCerApqkbX4UyB/+yeEEhdx8VM8D
7RPA46rLf8tKHWCx8PnBGcyWvaQBljck/9qXWog4MLsdXw1C14HHVcPtYEbKL25B
q74Vcw5htcQL9sBoedUhHyuTBfoleUtoufsoGR5rm9lYNtLsgPESL9yMDJQ8/reI
1RUyDUZdLCEEqbXLQrEVhI6TU/cN/CojSXoNw4JNzFE4nQYMFA4FreXTAhdUWlNj
rz7LJTG6WtFOj1eswTRveySdxoPJ3nmkDrrTRkQ2cC1/bFNGaWjRIMXFvOob5X+h
JXymnk8uAfdqwB5l++zfb/GMfL/0+9FLkAKtKfPLAoP1zDPnyNzazJRAq2cQjp5d
oBcuebCZBbbC3Zuakh+HcqmW5PJz8qL2xncCV1tzRB2l/la9uMj6NmfvWY36QNf3
FJVrsCUJGrTvPvpfrJy4wKQJNB8Nz1Ka1Yz2USX/pRc8GMO37w6LgrZ3/t4Li0nj
sKKlO7ZhZhal13DH2uoXZkkRDx1I3CUocsETH1d/S+6FqOYzFF1qQlDwzB8gEvg1
ulKL+oId0Z1Ie7nU2nkCPvBlqeUtRaF7s2kz9zboYxnOxmRSlQuyN92+3kOj2ghf
eO1rBPHBtctEIo5fIOWl5tY/ReHrFkgkx49QtSL7WjMyf5ZpoyoxAgs4knI1lok/
su2YJHJkFXn3r/8gNG2uMgmiKGzNkCAAWtVGr2QJfe2QiAdd+21rPVo+mmBYLX/r
Zlb9XTFFp0ze7mC8TZkikbIdvC1hip/2gHRJ4HgsN0iVwgTbAh5oMDrYySNJnngD
xWyqAAZhj1MSlQ5SiwBH/hU1UaZLNVPk/F/PPiMJJSg9YMS2Q06Wx2Fgwupl4LgZ
08/7KSSnP1dH99p2NKbuliFzYTEYYmRJ3yQKvXZ/p/kpDD+XODfSvCQa2RCgzbxZ
u2wJi00TOLkjrhOxHkzpfY5Vi1bvKJOBy1AwMJWefYZuuTu5pdh40OMEBXODkWia
CPrMD4OONNERTEEYyKFAKOizN1+Nml/4VKHCRB5Gy4uZz72P4d4+ZujOT++Q9fZa
Nsfhj8FsuQEiKeQt1YFdMqaD257lBS9ghtLqWIEg0s9HVgPoPR/ngb1JgeSB74LN
57x35rhk16EAgbFq7gZgeSFZFxr9/v2RSIOhvWsLGcGZK56bp7GajWH2Gn7OrQzU
SBhyBzvL5AimvOJ/rrjhzktCYiuc9GwwEy2D0f3nhErpCQJOJHgFcJ53keUvMdb3
jltoH1t1OVNg/Pb4YkSnsuBQ+bQUp6uAAP8lqLekmoFZEy6pyYI24LQMXdDswM28
BtvJldASeKvlFX+SIWGCdZZ+1fnVNMsOhh1mQQuaigKmeXX/sKcSxx5A83dYnfnn
3UZl4gJx0mS+efjoM00VE3vvjudtpgKFFKkzf6sMgSXmvbKiwlCPPKDCLkQ3ffjG
CyKnYhOOlf4AXVII89mdq7eTNGNJlom8ZuZ2Wrq2nABBjU6JV3WeDYnMHmMVWKyw
7TRXwFPJMdflXsMqrGYv+wg4gsWSEobX/uZXlWRPmjlms/TWFapC26bl/KJFLu+u
Sbc46cdMCQt0Ssatv94EYpJdICdOXe4MrG13k2xRz/ikzKn7yHTiCDcC9WRQYbkf
xE7NmuI26fe4oQSxSN+zcYdFUCE77ClCknRFMGfXjQ7v1qBVxNreRFG1b+dsqEN2
4qw8CBZijtQBR+seXFu1XaRO0iO1qiggwx7mSCGnQWl6+6DqXm3kHgKrRFrwt3As
GOimCqnmp2SS2QIUdftcyWa0CNMz4q65gdFNVsO31sVM5NlGt0ZPjkruZhLFyECX
rc44xkAmt3t6xK2pr2gkjbmT908suvIk8OWepK5+HfymiOLnT3nukMbC9mGUjQ3y
WiYcs86rG1XZeEN5pUbXbXaSBAtuYqTWgjVxHgauUjkBdzOhScQPdYuW26k7q2lC
hJKANdqUAmiRN4jlTVoR/RBZpRpBN37kvEEJTHaYDM8bmxDaKKwcn+S93c3SAF3b
xXK8j2sRULz9WxPhWoMl4WpQDoLSQLLxGVNqAO4Qwwk7QJ2Lstd64d7DwMe2u5Mp
Kse3Ffr4jukRFUCDwYS7Ab3elDRBFO9aL2uNE8p6+haKyKAMAzCO3fjYGl19QzXb
8lq7zEeHZQ50cxgvjUU6C4VP1oxZirIQo37625S5CcKFB+r0cOp0D5xvJDuHSqH1
0AzTd3g4lsBjotsYz5mwh7FxuYgo0D6v2DPn7TI9bJdhwjVB5PHTy3/8SFxmmjDO
MJfnbZKPfEeqV2+/zeNlqyNTqIyCTvp1oK0/Tbc5F9xadAl3dO7LiYudsFP9o+wd
c2OoPmCTdBU+OnJr81g5Rd0qgU3JqpjXQLd6hT3NQs1TgNazPqLREwbq6d4ZyrJg
eK3QUgAEaCEcFElUhOj7Gbs3gnsRmkIdKjqaYSzewv0esUUHgPmBFVhj4xilnIZN
WV5WhTMyhsPTSH+L7QK6KyPVKor+MVo03GIxvTJNWaVQ1yWsIwHxYZU1J4BtNWA4
yRlti2TBbx/xNEPYXZAnVyKpVMWdFZBHN4z0gXxMIwbiclGb3twrqqHlGc+Ns05P
hDnTrUZQe8flpFSVSCheBr8kky1N2fDoCz7fKJvL3wxTCCChkQAGIoZsfdga6/UP
e+ac++YtSxFRUAzxpWjGBa3LYagDAeX3Sy1t68GMAeB6bDPIP7c1Uf7O0iZSHIVa
UfX1WRNttzdngsQxAI4y7q+gsIhb7RWgl6FbBsdOooU=
`protect END_PROTECTED
