`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nULilZjZtQyCLLEO+Af4uKC17b+/1MO5GHYwrt6bnOJUgIddeOFFMoMCmTQkdNUB
2C23E3U78mxWhnzUMRg3XjrPs1UwS1BJDxn64iQDpp8GTylidtf+pJufSXV/NQOp
Vqy0+5wPCu8UbWbIwbU9I0HOMoU6ZrLpP2J770jld8wr233mWOeelLzOElDR4wb0
cqnl54+8d7hTAUJULelUgQ4skJt9yipSGuWCEzuRytKVxx4l7Q6PTQgdNyW3uBoY
GVPO46qpCdJieVx5kydCPu6i9Y2XBv/W2nWWcWNK8IfUwhUQqIXDv9LdlIHSvY9b
enmxnpQKQK+pmAlSjRWe1Q3Q34KNzK1Wc2dANbp9aaxaxOfx7rXDc0uJXkHpZDEc
Y2uws9epCgtf26wobCHmxAeaybgYU4fE3mYEFQmANmUWrtqKChZzrvpkZZdQuyE6
Kfw1VLZJ/QVpFRJ8dFwD5m+bvcQGdUqih/AJNacagwkbGEaS1rZSFIT3WBjR4pFG
hSU6EaUF1LCRNnmoPC0ItgdsKGoqQ0eaoRKdmxd5RJaxZm2oStC5uTB/IReKy6ty
+UudqREYXaak/z+jX7E89Vs536wbyfwP0kwcTuEL98KQSoA+XMpODRhvAXALOZDc
nANMl/Yjtfj3HGttr6raerXUbmiCTK8CyV8K8Z39GWoIEXIRQtMCEGH54sxewnSW
CAijnlWICG9hksO4Bzx+J5RCg23OfL063zSMTTm89IhS/ENmFej+onnycFvE6GbY
M2Zjn/iuZHfsScptYw0i3w==
`protect END_PROTECTED
