`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HbeY0rk+ukv9PUGSF9+hJyNnXNG6nnfmPBV+E2TQ6+6PaoFFI36ctVvxsEw+BFtP
zwdOb+PvS4terf1ZkLBaY1ajLYUwzpQS38j5OZvx14/gpRaS4Aw9B3+NGTO0MqmN
M/BfAoX2qP7phvewvErFNvUa5lpVKkqXdzgItUXYHQUv9RGaFk7ERJerZj5wzqSF
V5+lL4PCbBoyrW/CAKb0xxpTMpDn9bpO5v9VAeCOHSsf2XWCX2YQJTnQZOs89EB3
XTNB9IvafqCfOTKdY+Mtef4twI1CrVzwB2i6ks0X2UtN29Usc389h3CKxP1+gRFc
CB00eZZGYPXunEQciu1G6miWHgnWya6v0od4BeFQa9oOJ6d28NXc9Dl8CSJsvkoa
h4uf1qMnyE2khnIaySvDe62MLy85VozVu5Fgl4AYvCyT1GmmnqZRjvBRzvFobAGN
X9sbxuszASMFGaJY6oE667t0s45C/ocUnql8nPmavj4rzCTL2qvJCxKDWaR+a9T3
KeunzlaukipJBUSCEE7ei72OBojtyJIyLpITnRXSKdDg2vPqfGanYP6nesMyThQy
1zKa+/NV68kVQlfJP6sKN+n/br8r3Is45e3NwDgdvfxAJlACvM3EFjkOnmcO+NHm
mihN9SryLKmjCmPGOKPT2EggEYUMhbv644JGmSulTJljGeVpS1zKFhbKjIYqCPix
hwqzNdTh2gq5p2Rn3Z9i6ebD7XfO6Z+WuTh0eSuCtyYseGyCCi5nbeiWkz1DBNds
ofZ711beWyrc6LK2O0L+1ECEMzOzitM9eJVdzBbAuLfPSQyCKlz3pQgz66aBDE/K
bSs5+iQM1eWKGu0gaE78d+mo4dploOoYwBk9LDXzsU7eXZM692KwrLuAdjv0Tznf
freAsFjVbN/tnBP46Xzx/l6mkIq6O85/Csbp+Y9dClRoWL5dvKZiqUpgP/DmoJFV
djaVnLgELjUNa8M6OVawxR1APASZh9Z6TRAGwk0c8gTCzd+i4LT0eDjxD/KBIMDS
RUCO7qquPGpj/L0jhJkyGdB4L78SQwIm53Da6EMjxyxbr4shUaCJMofxK3AvJhI7
4Dc/M6qm1jHQOv1DXOl2OKbpWwnOAR670c+QzrkyQ5RCO8hq+doM3CWOk9HAEE3y
8z+CWixm0cK9drQ6o4Fttb2U3U5yrOOElAMk5NLEnUf5A4LQ8Axcpi2D92AAf8Mv
7CKI6rUiHMSD1lEjH6M+N4F+4j54VBBHIGn/G5b3PiOydOnG4YbHJLneyW1IX333
9x1bGfKe21fzc7v1IYJWq9ijs0OrUN5/rPMCdFoi2hzaqSsaEmHOFY0pgh7bw+dx
v5VrDz/kgpRsahcdKun65daKFbNBiS/fQlvY6qD4px8o1tWMybNsEDdJSLsAf8SY
o67ILQoWYcIM6HfBZUe82jrGdsuXMCqFkSG1jtdUVCPW6RYn625Gs8uL5ILmyFKX
G2ULyOl/s16gixUz+vnv91Jwl2/BLbrBmbZL/w8y3F3sIYSPyOyk2ZKBhFXzzobd
91KREOC4kaB/gcI1OgPbssdNO/Pdep0XHP5zR8/upgFA0F9HQeD28ajS4Mf3OZje
xsSFq/IRiFksefJkMcA9fkXZGXA4DElxK8kgzT6z6/gF19C1QHkCiH4AhMHTAkF8
Fp/xLhqAsWN1WAfZpKcHle5NNzjhJhL+US4oFU1V9RD75QqETNcod+5MvhZa16qk
GjwcHOX4/42C4iQ6YNeXEDa+DMGhCSPaKWMQQS/PzAMotlZ+DviMfBPMHRVd/IJX
K6NADCSxzhoUja41YtojbHzQEzeV+ZIO+PRktJlL6EFd1jf/+TgjPT3dnn6QmQ+C
nDdBlIptzOKJ0pbjB8OfNAg/fLBGvyMU/XHOQ9DSb6/mRWBIumm9b571G7Uaq8Yp
zzpfTEPzKab5zNNjoTBRSGmO9OnBGb7OwfNSji5pCne2I4lqHKFbJIiME8qxvmLX
jgYENevsMD7Y+9ZZcyqqoDthCQy+P8DCeyCAYI3RmvhKNnUx3NAh4hyzxhDX5WaW
rliJjOU8kgILNYDq0fhUF4DUHZJjPm810acvne1U/3jk6KEpR2sVXNo2vDShkdvb
eRXM50dyY4sE9xxEzIkJol78O2mwrP1WJVuJGDSsMdMuqH239x1HU82WRYl9NFTe
9BieYDdww3bFAQnWZ0EMzr+0lv21flVNRpgk4XRB/TjHgAcKCqSQIbMOCSmcVxVz
IMJ2tqoxLPcujxet3xMAcAu90KNJOpJ6DnlX7EKcd1QQsM+DmCQE5mxscGamtR8D
KKsTIFgzb0aDnyxUaGTfX4wgsNF228uJirRycazcrQunExWEAi5ccosbaKC2ByiR
tayn8kFK8IejjCEg2QgNDDSqHRGvtxAm3+8xY11/iXyemTws7X+3wO4Xp3/0ul/h
SEDeNZUo+fGa/L87o4ZkAxdJv+L6cZv2Qoy9ri6ThdstNdbzytZWf6fXYK2Zlk7C
Ux21PXJio7GkrHjfUf1xSMS1dFimeeo+dXIcCdWt8RSNaNFixGifpO2GjX7Mk4WU
jyfs+Yk+IZn5iAoh0hekQzsOG0ObbYnJcvQBSmiOy63cwAK+zbE/FfQjtiP3PICH
JWPTwi398rftVKDITSI6YrXICse/U5QNi3Ky9rsRmI+FiyaxuYn/xvc9WE+ioCtT
xzXQGJzMRyKyZ4WbjeevUmL3KxqsGNgWoJTrjS4iuSKf3L+CvqE+zeW0B8iVBTQm
BM50EqzT7LDI1WUCPLqCQ/R1nAGt0sQ+Q7dmeBap4hg1khGj0MFTs3ZdWXXuGo3K
AuBfHgXJ8QCT/TLadpyf+HxgiFgeGLL0TFWByWfZChMYgGMEBKn40s4kZ/+gmtQe
yjT0r3r0p6Yz0sWze4/GsjFXUTIyW+I4i42pnKM137lLBTenKrJrhsurJqB8z430
qjHyGdVqTKF3inlLyOZCC+oK7YlIzLvRWMaBPZQMVDjBCrCO6+gFdG+FxidP44eE
YtG698rJo7miO/OnIGXRpg/HOpvIbAazWg4H6zP4Xck4YDkmnugAo32hYeduT/ty
W2FoxFOgJh84D6l3XBTNm/RE92/GOlQJmzkmUrBwL1Fv4pLbzhrZqwguoLo8FWql
eO4VQTlpEStnBwGdhvF8n0ysdDWzVaFLTAwz+uETZawj37otAeV1JaftflE263k+
W/lnCBZWm25aZudl3rn/v9JAq2HdAY5PZo2mDAcg0mDiu7kTgacjhYQ+MrZGN2CA
hE4xGhnxZheZ/DGZORn4ZzrKinJieKnAoMvdOmL8fnP8ap7kwgA6Plg9xLG5YZoJ
fRYdT3AmjfEEf5yzq4NPDs44EGv+d9p/AxvxHV891XecuZZm0/pKCWjSMS34GW53
qW0jMBP5KEzvFHqBVG17dk1c+RMJp5KLJw2U06lOAxRnak8gWDMYmPMEZF6kBPMC
cJ6WQEl77QwVQGUJTiJti56rHfFNWeyRVYiQy3GshkfP/pXLgWgF3g0i7R9Hhktj
JAg4QVjlOz4yndeG7RpZsvUFpFOX22OvN12MnMMIQTtYegoYkP+kNhxPGz2kZwSe
+XxsKLsHkeWrMVySTy51FWZIC3WIUmUtDEn02krowhVvfwZ91o6BNReo7H2SgxJV
B4rM7dbiDxTP14kePPbn3JL4KAFFa9FGhkLwrYohAATgtn/bv4VoKumZc6bBfcD8
HgIwHp++0NLMSMoZPNh3agqt2TiQLw+CS0MwL6dwAm9w0psUU0Z5C4W81yJCvmZK
Zl0PY3Lqqs0/bcYA8GScgK+1pL97VNmz5DmI7an9GMtnlJIw/DzCL0swz/ICTX8l
sgnVjApE2LETBhj55uNDRf+SDgFQ5rw5V1nWLH1EK9KXwHvuso4f0P9NCI3njrRf
ZiM5GlXOdhADzOSQF2jWFeslZl6J6AuP/oRS8pgxEXtt5UVmOQWYnwk/F32s5t9f
QeQCZzgiXZKnAIf8Hm+YRlfifUpqi3/JbcuE0KwqizwwmYiUhU1T3B2RWejYLX8u
5zw/RqVE/oHVwrGWjW8AlIrzShFrumj+vTDw1PHX8Ut3t5S/4Sdp1ZxQQmxhy3RV
vts2/ntVX2seFVxaZ4NR0vzJBCVNPKO/Mv7pBrq++MOjcCN59d0+jkUGgXWe/aVK
P7FAvGEbfYkotx79/VNOLyulovsDYZGBy9faIIkaz99Z1sgjYAZWrxz1YlqANfFq
XMSPtWP4Jq4ONweAUt2X02vdOsYdO8/SMYJrjPEH2cHd78HoW1z+SWma0th/lsXU
F3wS0Yaki8cHKSWt///zAsIigIMzOm7bGrsbuvJyUaT6E8azA73fkiRQbx9zHiWd
hs3306WZdhgh97oO/7W0zSvLGfYuOJA0D5/ovydwUHv6S+dq2N974e/u+5kxAU56
3zZY/70/vbdoipVrdIDYtMeeIP/57IJhCOO87uwwu8S2++Xw2HwpGgtkHNJxMN3l
HH2dtFEz22WTOaqI/83pokBlmQis2FxdpRpxDTDlH3uunKYPeDJsEADN4OZaPQdF
uTsNjLANuYjnv/6YdGPgw0QX2gId6a9E0citsldi00JeyuKJH43i25BNJiJO2/tG
Hr485AzobK8Ou6uSt/YLzdJFhW+RDJv0+pVIsS2dYEIqykUD56oU8i7Y30nVk0K/
57Bf3e/i1ZaeBcYhq5AXbH8Wn4nO9cnK8dyLvnCkazvk3axy6QyMATqWRFHX7+Fj
kytONkyo3dzsyPBWf6uY7zaU9c7QDwMNWswf2M1sMd/Ndyak3CLxeH/15E6FhMis
oL1mOTptI+xSIYdQReO+oIYs67iuaSy8h8fcG1GLBatkeKM1rWEzuUdxxpR5Xo8f
vLFQcawiUC7YEqCnKvrwWd3kZWzL3Fd70iH1H8m6pvMxg5fZJYPsO22OJpG32udU
ZPJbi5omxW75oGPgU1Y8ZCVt1bGqWfJgTJvqvOSAOgXswuv9lidyWF8BP+bMnubf
9ypmd3kWCfspW57SMxxrG5SAM3S8Od+Bi7k7QkSDmn56mLcNw7JMkkLJuHswMfsa
13oCRzNpl+PCrnkvuzKhRbnhtnlvbIXna3GCk4EjYPf2Gg5yc2yP+ZewOSbz4ccy
KjdrvzjchR85Mp8sEnb3IvtWxGoIqhUSiOzXopzJg1vUKGk7HQGq24wJP3XQvFZ4
32G4ZcTbjmryTcMojURNX2mNHkfwAbB6RSkbweQYBe0VzY7yWQbNqzt0dr0ohOd1
NHe3/JaBcGVQjDa9E0Z8yrepP0RB1JyDrmGM02QHPmGWl/2uPyogpHMcIdTbJhUS
M/nowDnCiB5CW4NaQM7pgz7e8MPo9wMYYNHElf4x4hzjIdX6pWLc8WFTSziocqWz
mgrSxM+sL0EF22IQjs3u1QFh+6Y80QsWWMzaqGUfLgpJ98skauYAEjbGZf4H/ffb
wt0GqawfSmQh1M/KSE2BlWAsWCQF+Hz7zPni3XVFJdqHZM2cui++N5Iz1MdG6eEe
v4tQ67P6WRkJL891v9XlE9/Cwuc+0Osl/C7tc+gx56QlSDZ109vNhjzRPYr5LmGo
f5yI9P9vcdZbIC2zbpK1bMU0ebi4cilrhk9YruvkJ9v7DvN/QjNDmoELPJK5Ab6n
tnikM8iXqncl4IcGrjaz/Of7TwtJY9oA+maElrDh+FADVhTJowvhLITeVMmLO9JW
/Iike2Iif4lWLH3uzB+ollc+7puP4eiVBtdbnG3uRMGo86urn+s6jjaCgIHvwthW
6Ye5DsGUQtkia8f8yx3Z1y+3KI6Yp/6n1s755vvPcbJvOemFbhfNhTkDzWR6s3k4
1AjyuEsYDjNrbzpjnuxF9b2nh2DZ4IjPmX4V8YSR9TZ99mAOxHpUXnZv13kfSSxl
HpPFlFQ/zA9v9LK+fuILqw2ymWPiG+HlqnaiA/RQqrl5MnkbONXoKhFH09HqS4rA
81l7mObj3ap3h6W8mamav+DtTYmUEBcMfab84IjfZQzfBzg58LYFKKAPCzL1Hfkm
74wG6Su9YNWCuuK/OP03YS0C703U+qpVlPCljfhNui4mRVuxAosaN7XJ6qVcgoww
6hHluWvHAY2+WvMHJFjUYvXPSDBPhDflnNvoRMy6H6RdNbpBOlDtl+o0Qo8uqKXJ
Rt4YG+C2gglREPS7+w/T4368eLvW0J0NUJI6ly2pb1C2Vvbr2bbFjAqnhoU8LFoA
J8TGT9h3pvr4YaJ/49x7KSKEOta6ZFXImpYkYdOaYJ/WIVGg96ldAFE3T/vTwubf
2OO9m0XXLMo+1Plqx+hFgTt1HW1Gtkn+9xKoD7w229Ps/WHV15rFMz/jXTsNiZj+
Fin2vOltSDG+WSwOcgnWskLHGlJ93XDpnMm7eqa68WSl+v7nuY6ZAyCNSstBwMxf
+ANzRAnH1R4yfFoFWJbUA19u/duanZx99gS445KmeEZ+A+AtTTQ66iiwAaKFzqft
okI2K1cDK3zXSNVdUq62dOA9wBzebaUxLNqWn6XhfMPmhonwqqUlTwymQXLsfnL5
7GlOTU4gATpX8AklH7t/qVu3svmt9WEus0SqWSDW5BGOkf4pLNvsfxaK7yltncPS
aDoFJf85QZpkivL/CoZWEDlZw0MUmHIjMByObhYQ2ezw4g+M+XQKMluhuJWDTj3v
nxXD7OZ9zQqdlk46RHutigEEDbiNqXC65R07Yj7a2C7as9HNjGWZeCYtFYQ4Ep/P
ZBD+c4Xbcf6PIdx5cttQi6+hzaTuVPY9nLhUqufvEWVYXfs+YcWcOam1u9YYUWZx
DYXpU9Fj+PhaxEBQFHwrrcHjB66BR4lyFvPcpV432pV1VteLeCn8NklEb9uGLAKW
heWbmAksdEYuLvAOM6jv6kaDHTguiS/wcogx9IYxiofKc8gTJUARDqMrwrC+tS4n
6kMagNTLNS9juJhZbIDPOHb7JZWoiE/5lI4/Yyu/tO1bFAoPym7to93hLMOxbhTf
hLDkVDrcSIKps6180sm3MSHo0sKfjURpdlMTh2FQeAeCoyjrcKeCFgwm5cE8PpMY
RvNLmwId0dcbnzrgU7bFlD8udHNVOewRP6CQu/3HpIYRpWFM7ynYMRhbjb7mLSTZ
AK++snrM5dkqwdWjYXX0zYjpmwyO32jv6IOW7QVcUi+ivtlbDmrFU7vkwfSKtlQH
+iDqneg627heVYnfGzijofX4y60spKXobMwdeHyLQziO3IIFQaLSaxX9rF0iZgxO
rSsNRsXM5RjVXXjqb6VS67Af/6CGldSVkSGWgAPmbYnAQzU5EvQG/kLYq8vjsV0T
035ol2h565nZ3YfSiyXhjgfrFg7CLSroG17XVUoDbAQOXF+hbaVYOfEA0WBAcf0y
EenbRzIuY3FIbaKx4nTEFzsoTQeM4SIARZYCkzjOYlk3PNeWVVBzn8UeXZSbj0Z0
XuKB+czO8Yf3+iR1MUoYgPGwM7PSlpBzFuUMBs8nucCuIBXxkfm8bpcTEQrEGxlC
e9nUM8NHOlfvfDMUt+vWw4q7wyKEpNPrnicXZfI8ZMwyzXBbtDKSsRL9qppFhSOZ
nf0TGcIwbXHVdrrqHQ5P1Z2kUX8wdEXZxtO++Zj2cOMSEj2EYsNKccL2kO0b6+Ym
1NG1OHAmizImkicBz2tlZgua2+RSMsOZTMmFS4HWSk1qZomu8Bfj3ZgXXnFECkWf
LdEyT7kjgfpU1Nnlo2nm1NXJ/3gh6E+U0cnNoV187/L6wvpc5BpJ7SFI18wnp9ro
Cyv0FvEukgUgp6YxjAV99ZTUfMNWKJWzzdoaRDauJ/NdT2yZDgWQiWXKwER1tDuf
QH2bBOwHJIDVFwxwFFjtOUTqc8/eKEnZL0RmMdizMZ+VCj00ICsaMCk2sDGZojx5
WVz4uXxqiYpyN7FxqVvMqtDplPwUq9EOy+/wUug1Q9yEoV5FosrBKs+648xLxEPN
DncWGWmCUjJMZa+Lj6m+74oP8t79R6c5k9b6WOFVvzJY82qTgVXbuPQuuau6w6mt
kDwIpxx3hWygd5eYYW7NrQyRzZqoO34x9V+N93ChVVPkkMRVTDJQXCWvZWue0/TM
jl+GgqHAEEpfdg2U8pr16aWcEZnRwgGKOcvb8NwLrCcMmjT3WsD8FaWQY995l998
XCkCw05dNSPhSqZn3Ho4WS4TQ0mBBTu+y6DETabg1sA0uWHPdis00vTvBc9876jN
OUXcv765i3ppsxpsKgYV2jb0hFIOB5etSYbiNdONLOlOd6pYmPBUQCdQXSPOzUTI
i2Ji0x8i5DYb5cKRADOKOs4LZcYc9AbxdHz70b3sohpwTynBsv7X5PtIzsjgo2X0
LkXvtM4UaCid7KQ3d9Wg5tGVLQcE3nYRFUJbpAXprYibhrVmsHaI7UXLNL4EsEP6
o3VWfFF/8k0MSl2GBq2c5q9AeyjPE9xl95DRuyHq7rnFn8iL0smPhVMZ4QdRYOPs
0C33sHEZzJe9gHU1ppdaxN9J/40twWqXdQ33ocnZ9V6mMo13w6hYg6a0vTa3w9HS
1TNzSZtlf4c4NSzUwpRhEZots9P5JZ+SzS0AqQ8B7S8lKUHDTA5ryMQ375NDdkYI
Xun0sXbe7DOyBZaF1IcTVGbjjV9E432+HZEwNAGkb1RumaL5MN4637VKLYfTy2up
7S8UYGuWdCVhODixuOsHjYGISnLQFMaBK80GTw5Yda7NdMzQMHy7XbkF3mroE8H0
2BP5dySvv0IN0YrfgsXCwZSSIWdGT+De7c/24BjZJ9+8Hb1g9mw4QRXqijHDp2Ba
veCubc21SQOGCaXyrwpyQzETuEARDsLj5gd0MSKCUFaZHA0EtXYj6pMHUaRLoejA
a5BLmh96xQw5LItEMVGuPZ74sSI4H4u/Q7YN5fIf2ABnt4/1V/q4NIylIxunn2Vf
+kb03guNNsD8t1EGbXNtkmdn/tLDhiJ8g7wl51Iet5Q9KJU959XwFY5xfs9fWQFg
47o2LgXnzCMdnmzt2a6OJLvbI17mREPHaYF3yZy5vUC7i6wq6lGbiUweQvLG71iX
PPyWWs9E89rMi5U9B6nvK9WoYakyctMnfjxyFgx9fT0T2shwiQYJCryRem6ZL/eG
SD83D4a586iVD/Wxg2XmUZIIAfIERCadvG1Sc6V/F3Mg73QW3MSNSMQhlDvLoGSY
B/VlXcT8450NAp9/IO52ii+ZwONvbSJtalob1VSNEcnSjkjGettQZW0k0m7VWfpG
QQ9cehG7a3U/hPiZ4Nugz5xC6tUvz2SJKhdt0YoYS95uQmVEtY27vaNA4zmFaFDG
GcYPt0d50ri8nnitH1lmaHvP+jDa17aZ2oNS/r2Mfwxegut/WAC0OIxlrWT9yIdA
X4huOVVTtzACBMyHWNm4PwDIhdHWrH45Vu/E5EsW2GO2MflXhAZ3tOonMa2cE03C
ksUVX52kTDeaVFiEhTKMa/JngjXvdiNlM6FwM6/f3c9wBUuy70FdYQFtsB/2g0VD
NaqzdxIB9iSlDY6DUa9FqtZ6s7wXN3uTd2OFE9ewWUBuTu1ToFdjoQyCGkgBx7uz
Soilgfb5RRbE6pc3HZTZf8VyzsxJht2khPtAo6DB5Dwk+42FXJ2G9t78kffJivEd
DNRhdTrpbUDI25I51C0tf4QzXKuA40Y0OtfAypnkXf8OXWrCFN+KZ388iFIl3cgI
HHBYE+FH0mE62XoW3Rj2CWkRdH5y6ZzZiBHTBLWfAqKDgMIVf8F2ch++mWdBRWrz
+UW4PCZ2ZDMVUm+9p1mN9L2X2QhtGomPPor8PeCi87m0eeMpq33VOi+hSKZo+6ue
DM+8B+iqQElryHzb27cycqu/L9Fb1SvYaU7rGmvlxm7Oq4Hjl8Zkb/0J5CEbX/vO
7pSZpbv6sMQ4cYMCis5rhd4Wci5W2W/wZ7QY6isQHY2VjTpvf7ilCTx6T8yIgEuZ
Dcb6GJmW43GHbfcN6Sn8qJ0gG+x+2rMQtdqWJ2WgnBHsjK2JObjqZAruSJbqx7j3
XqDLAbOzuh/4NDA3TmIMN23saDy/TACt1FmXuhM0O099RrqpOHpk+wZ500k6wmbO
fLwrJ1Lkrq5T3vpGwHqsvqv0vzoefgP+gNFvw1MRSj0Cz+b1TW44o/bmRN5gtbf/
/S0LCDzAUK/VWDtPxFAQ1ZOWMTTWxxEt/k83qG8hIOP/SW1ql5HB/pDRsluY475a
HFls61a3XlOIDtrKItKfpQ+Oxhi1rx3Esl1nMx51L4JqLmmJlfz+TeVysDOTGIQr
6aFXnOdXUoRaZ07WOc9ma4YyeKg5BG9Wj/vatukKTMlDmtHgqiemjNjsR718dH9j
6Y8t8vVcaxBqo57Ci3EUCw/7vE0wqZ0Gv6fbKVkchkuBZ2WYg5QpSkrmuF7FIcVn
Z3wgWOtjckEAzs9zdykGRDufcb8OZt0QPzVH80pPVci1ggUN6wMXRME2SOq0x3YK
ycknPMfJEa5tVqKqUhkztQ711HNWRoyJH9K5gC0f5R9NHbtAGt8jNpGDp2cpgv6m
xL9Yv/MmBZo7Ra+XcnbNtQ==
`protect END_PROTECTED
