`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CmNifKsrogP/apI9NTFHlzbxbS2IwE4HeAWZqAtW+AXFWBJ5vUyl0B+TNznSQJ7b
s+a27HAetPie/AJ8s8R97gBmdk6PeK+Z+C60oBvoBeBooan1HqgiF3GbRyU8HRwM
owiHnESMG7iMHLxq+O58ZX2Myj15m0x71K3jOxy8KS73Q/SOi6+C37t3CCJLQDdC
lzy3tW8AyXy10/a/+2GIX0mCGAGrLR+z8UDQwdxb0misp9WiW61bDCWRhNKJ7i8p
a01inE/NJ8hSoedIMrt0t87syM3yE2arCofk81hCy4eUAHYj6x/P2zBsHmyMSiA4
SFE4npdrQ6e7zeHNNQboyqE56BhUy3HTeOnGobeNevgUjtYXAqMqFpMFhrVSjbyG
6YZSPXPAcCYu7owr/naFcJ/PTMyOaILeu7UDcQKVwy8UVW77ony2sTJG6fM+tQXK
Ce3pejyff+iqndrtkGkY+QqHCamweMQh76hzLORpNUXEyipOqzsOhkZ8oPp9bVv8
+sXfRzp+r7kajMFsLkwwshtXuJgIqOKyBE4e7xiUBM75XpCzl4/cSIwKe2DrNg3Z
O28YJnSvCv8Q05qjEn2FCWigY1KnsKd7UHNMg80w5hJda25vs/ZZp60KRUtT2d95
WvBXjNc+71Zpq8QOtFcxuHk6kuqXKXRdcbrY93ZkUTgXcz+11heDc6hSpxlZpqmc
gcCz9/Bsbh7sQtYUeE/bsEiNx98q4VUfMwf/uHU7UENpWOokjNL8YxT+JnnbH1+B
93ujrrkpPi2ZO+rloz6vdh4SpvsvHeM0bmsOhcUE2wUTv7w/NNV4WtO44eeXeMWt
YQYm/n2/sv3thLAhYpM3f+jcVMTG2eoRy8gKAouzAZKZVgwa2TXdMRK6j2WNKo8V
dXO4boGdEVRXTr4tqubSn+MB16QIT/iLDzSxWPKisHoaZGZ7mSyDHfi12UmYiNg8
75UcBTn5wfcjSavx9l7y6CpSjIeBcysU9ZZzpNFzZTwSc2y9mH4UPCgD43spPqnv
/fgUgFzA0pL94NzqRovBJiOWUUtW9SOt/n5k8Fxwsio7tEzO17/Y6O7sAeqqCQ32
N3FXl17l2QU3DAQGTM5PWL1vxwfh9oupb+JGd9vkQ0vYrwS6O7sdguJGoTccIuOP
5jkdig3Pseub3VWF5xwriRKmIKlpT1JmCTpbelCw5VVJfGkV6D2M+jjvx1/hBX+Y
XB+gd3Vp2ERiPALl2AImNNmqj8zqoGiM4LxRlOuUOU5GxGt4YaUDL5tdFbL0E27K
l7kAHq3COsrEF9L94Pyf8NY+ayII/TnkFq3kOPFxbOjuq9dnumqG15fPI2nUtewS
DTkmiCsSjeVxc4VCWZvbGms7SYd/dqybjeGxNlgOP1tSiXTLKwncnibiiENCoEnU
jdRu3E1QdRUV3LdzK6Er3T34iyl0C9ytjEmS8TQ/1PPZvYRytCNlsIeWWn0k6Mt+
BYEHcNzPL8rzg3anKvfAl2ENDBdu0Si9QfjFuVpTgHeVla+JWP63eOq6jRJdsjLv
4whfBKasnrV+mEJJbQ526AcyKj+vEsNcImUTvtNSC6vbdctzXxaZ3erppdYRkpmn
dXmHr13+f6/WsYo8YAtQMXBwtXgSRyjPgyX3hJfk3j7dSYCT413am1Nt+fHqPf9r
RjT2iivx1eudBWTnRKZ4CntDWl8dtzPcZ8i+245/uq5/e8LY+uyR3DKDWKp1lzRO
0aKvzE8G3L/mpoDWwg2ctmHow1lDofdTZ6QV1l7lxup8FjL3PxMA1gkT9FzTTbKx
xNUCRb2FRBGWqdogDcDy95K179L7P3hZ9YumX02zIBSLzn/C/qXc/+FUhF0uk+Dh
WyqYx8AsmMudMyAc5IbRSSbipv0/LpUsoBhuppfo5g7dyahtiTZA2WuYMPcymWT3
sCjNGuNwAw+orbbAQIWxczJC5tQ/GVh0kL1bkYzmJK9Sl1idSJm608++qfPTunk/
YbJ7tbhl7rTqGvfjc9kMy4rNP7ITb0QLXeZ1hK+43tGpJQ2Qf62sfVIXhycWM5OD
75KvYMcYMJb+Ru8DHOiKzECo+KmjDNN+HAxstxMk/vibgochoS9SRZGE4LaE4Nrx
DQAJmZj5J7W3Am5CVJJpWKh852qmalSVKJWRJydFTTI=
`protect END_PROTECTED
