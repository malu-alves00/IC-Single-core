`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nWlEWNNX4avnwn/gC4y+jud+XgNpqbuC6pxCMMV9aKaNVAjXRJ+IYI0UM6sh5Zdu
Ze5w/9+dGzRnJwSt/aoj/5De9VLWwxOiMvXBAFAYO3H53n8f6YEnHo7pspDM6ktu
1c7//IIce+TY/lIoamZM2m0ncSgeVMM89NE1pe9ay7Gk6lqG2NfGcti2pi8KOX7W
UiI0xPwSEWiVZT/21AIdfRqsCZNUga31J13YdRxsSv1GizPbhz5PiBLSKOlV/2+G
h4+BgYc2K+a1TD/0eAYiAdL5ppBFFixqE8S8qp+lKSsLLGL7SajUvTeVMH1B+dZe
IV6FY/zI3UJuYPA+2Ynpy92xe/XA0aFGiIIjvINnN1sf4nXitH+SPz34QjM48P/A
Qq9uh+x7biIRhtpeL4eol2ph+pWHuv1t0jB7VHeDmEIwpsAcWuoXx+sBu3MXcZbS
krmXdATnUenESaS9EXPbZXrkGcxQJjG6Ly0K5dpevnS37EEzC4CBu+vBZtVgfxxL
mnLzk2TgZWEwr53C3LWK6cH+N94jrGcq5gTDIMnMYKn4VG/T4es2nrfXQEJKFiXJ
MBH2g2nqONQYvIzOujKwPsfsSoERTcGWwyRQYXZpsjFZixM35Jh3DPdrVFwy4ibi
wDmznd7tW5PGuqze5BH9fvQNsutEYuH6k0KeAdfIMpg0YtWsL0bOi5iAEEMd7X1u
Fi9QOc/I7bEmfQIeteSRm2fiwg/5XxJMqn3MCZUbkYU0TFxjMdsZABW9O/f23kX0
4tY6lkGhVYzyHDOxmryOuO1ZKLgc4Pv6Yym1yRS3kzNokr34wsv6ArsTwSvIn6qz
I0GSTO3i57QGLsC3iIgzGS7Tt1aRgbyfic4oaCjCMBcqh5WGKfDNJB+ql+z49JhJ
/SHhXoHmq4Spr+o4reyP2/GMoJb34LxMelyIAAvdk/7WjX16d2DmZAdZXEHE7rKx
LSrd4oVH4/pLP1STpEwzU56d5F35CljfdKUbCz4w/n55cWX2HQ4kgXo02UEd8lsh
0XyMjpHj2oSzjiJjQVLtfihQwB9LXnpq62a4Dg2fhDlOa4Xfq9eZQHQh+JswhGXd
snGonBdA/SLajP7aWQD7Wj+Ncz7x2I+GlFFcv/bOP08VWoEh8qdeEYuYb27rwYVM
AQktcz/DzOTxaXMzvHZr+ngBUZwWA7kCrEfn6OV3lKaesu71XyIFUE2EgLOoyCc+
adzD7E8fcZTmbszjiQu/EJP7GF84GWQk0sx1g+/BYDxibskAMADppZksB1AiXKVp
hrSZtNnaTEXXqihxBQOLIes94CPxY08tB0o12mztjFJ+pqYilmSGBdAaGge4ZT+d
w6BKCphNYzP3XcX5e5w7V5kDcCpaS8PbvNmSioGpAN1InW/VYRHoRWfXYrA+RIoO
EF+MkqoA5khZOqMWEhUWHqMi9Q0/olNHla9dunv9kDvYLeDlZDD/bTtBOnBSvtVY
m9G3EIW979tm3PdHY9ej0HauRYyo7OyyqUl08JPhwOyHh72EIhD9vs2CchkMNLvV
I4ZwKt9Z3FwZ8MPYiR0DiMQwc0myjW2iKj3ocSRfn+LE/vLNxzp1pasQhI5RzOer
r9mQhvgwrlYXtyylG0hOChmAS4vnxMEXNUbjrFgKFERZGDHglMSHqKtNh70UwaRk
glqsN3678IPjHY5za9swWqeFf1FPQdsIJhqMhvwqfDZR7gH631/hbS51432QLGmW
ewOGlxq0PYzf9hiKTc6j1/kMjAS4VaamFudlO/Krq44Q6NnxjTnOuct1dN4fV9Jn
7gi96IPcArtgJqWuE2tLKcx7x58H+b2A+69kAaEo1RicPpPeJpQH1nmfwF1l27kw
`protect END_PROTECTED
