`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BFN96z/egvPH9TyUmxnpnPva6+2aAGX/VE4EP/Q7QKW+5o8xckDEbj+TU4fjdVLu
f3NPyecszr+57/sVo2D3SXnJFGebmfsV+KvK7oFYleuiOoKCVpze/ZPHGQo+DQXf
CNvuxAti47sAl8k2nPHJMdUgvUe2xdGQ3s1O6mvpArf2ylf1FpGCjTyFdANOHvW1
csQTpZ4ypMiTW7B02wpk9Jz5dLAO8512phLK4zKgG1CkloyOz7+qX9muef9nrYVO
lMzKiGsF/f6BJejjj6nKMH+qvQF/X7aUbIFENuwUz2EVp2pfmsY/guKCJgLBw9+v
SCNswcCzg5gdIaDyGtbDwDeZMWCumaLVYQgj2LcJs2srvfY3zpinfpwRCOTpt3zr
N2AQaDuEkG3zL3Ww8H1Sfqd/X8wnaY7/bUwGNrcz1F9HWq1luNXWTs98BT7Wb/2X
UvQJvUGPbOvvPx+kWMSAIbJi7eEKT3BdXR6rwesGymMLniTOhjmDsqXMclolEwDZ
HZzJk6x0tq2vqAqvTVzw+Mw4z0bRqLrmTwHmQhqXgOkOR+F/TT34YFzRXEbTMfac
Q+97g0uCIp3fKFxnI8NTXMD2yDKsR5AQjUX3nUuhqd6DkcQwe0c5b4Ml1NXir1Gf
3CwX/kWU3jJE9hXVf1bSe+d/IlD9Ij2fKQ1onuYo0751olMhiz0HVqS2hE+At+Sy
VL49UimNv8bBmkMUW3Mah9dRBwGxIVbAAijIf0FWDPK/5bc3uDJP7aPrNblg3CHN
dst/iORISMgzFPKAIO66YIBmw4JyF3sXcspHvEx0V4IXioPQxZmRodVMutN20r+Z
1zuFspXcxc9ATqd40G1Mpz9OAXp3Gm5T2FnZmVDBYvE=
`protect END_PROTECTED
