`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eItwNzr/iJamD4H4y+SbsYqfjf/hhisnvtZLAx/qPjatZcBwWeQS60KwaZdAnQ33
TAJ6z9gB3wanjLqBqRObN8BBVr32GR4+OVG3MgqVx362skNsy1zN32K3EFOcqgcd
omsn4kAr57EuiY7mDsjMHriNGIOdbCX0b0zgBVO9NVHibPRlWFIKGhVvoOfAwKtT
2D9dZiWAhoS9Ae9ONjXe3DJH6Ibh/Ft3RPIDGTBsbUHAcXzHku49SkdCuOqi/S3k
FOv4xJtanJxeCKoculeC304k65e/FNR+f8ZaeIWNhniSi34hldUui8Y1mXo8AYDg
BMqog1ohefWKnX51Yl0EwtUO5ix0J7DLZ10RHEyMTwcbomAvi5Rs32WxTM1S30Rq
DU/iu7Q/TVzTENRO+YIQfmBsqutEajHQ14jgrTDTZdoZXJL5MjlYUdUDbhV62/GR
u55VvgriTxhj7YPHT5Hb9lVFO94opv6dKAujKWh04TP5BSRHd7nzetS02wb2GWCU
+8NT3tmkZGdaMMI5BCE5fJJ2qY2QsvergOt5JkjzughS5Hl+kfa0/fUXe6BYEMPN
RVIfRr5OZd/Qc84EmQ7qJGNdMT31yaW+mEhBqsrAROgkpuohSEeb+k3BcYkRc4YQ
9BRB/qLm76cKF4yT5tk8z5pBgv2DstbPVMbyqB4yCrmY0ZwAeMj/nTwvjUz5Vcdn
keJ9j6eunDOZnqfCHEZri+TZUVvEzQou8ogJaTfnKU8bh4WtMT864gKtN5EhkFyY
k7bOE7aBeZUwgHXy4UlmAxFbQiAVAVbsKqJLlaazPGphaLSiTSVvpeBfsyz7/UC6
jWtUTjwC6m1nCWhc00rfG8o08zd0TyQBw2Uuu1U6taJzX9l5Hm5pXKV1QKvsMLEo
B2oRiOqUATNb5nSQSiOqUG73A9IpIW0epW1OhvgvWsI=
`protect END_PROTECTED
