`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9Qg8E4TCuKYFdfGxgKjG4EroJER+CZu7aIUY53kzqEFbu0oAWtrF0SNvjYtVQofs
6R4WX9C8PtgVFaDP6QHxHR+GCACcotFgQvKKEWsLtix6msKdZSPGrmf5Jo2PFi2v
TAxke6b1bINeo1g59WiE0A4DqIZfViXfRO3X6InD80rbNEH0y+OvICIdAbzL66Df
7Zn40cT0zWhA+wql+OHutYLRAhK+5iD0zC4oZOuoZjntkn+sSSPgTTWyxf04lPFW
Du6F9THw1vjU9uTPJrNzA07Yp8KACjLnRYR6DrPcRIA4lgniNgDgXIQHIDOkj+G9
wfglTIJcP10Cy4pn4DJmHxV8LOjvKmqFsjVXZ/dsqRJvgP2Xq9+KBLMwcpIQS2aP
FQCzBR/+W1Ujz58r+0wYOyjEuo0Mp4n6AN0sPAellP9P+cs8wv8rP0oQe9/H6gOG
22v+/lnSoe4CRIuYvwhpE4aGPs42qBN2BnwHOwImDHQPrCcql36EVfhBGJ4gjxUx
swFPRiLFY6E8z2R2zPiRuwRla/aIMbiBtMIgvmW0ExPUMwfqO0+YFLUTwEpIr0Xb
Tu8GnN21prouuT+wzcKoO+uDuRehBJ0SMCNOxIEp0Bw4NtX+Jyu0htdeMjRb2QyZ
B+ig6jdnRiBmtORj8s8YlP/lqKvt2tM05oq8e6KCGXkcnq7tDGInQtrPgR9Bq343
hI091x2sZEKFm5pj3jJySm2ofmZxEsVZer/DAzwkJ2N033jxRpmbRzLX4KeDFj6U
bitNc2MEYN3ETzdjWm4pZ6sy9Yf0s8hWF+8+rJVEv0u7seNVJ6p70BwofD+NcsDs
XVnibsUjwyrFAdy+bLVwwQZyMqb9efMdmKLsWQ/OJRChp7Y8ZhgdvCt9kPw/mt6Q
LhqUjr9VuSHOMZd0Vv3Pec2I2bGLED714RZv0blqkYmyMN9jaeTv5N+wHJZMEUXJ
fXr1fNc64UoQBElVsY6FaJPQA+6PupgN51nIgcXRUn69Q2RD+n7gRv6bserfVNxN
zK0G/x6/z+zH0tBBCPrBfjWJy/ItFBDdzYKhKS1iUIq59SvDAM8OFDFWqn2fJ8XJ
XR+DzpTNHrNrHuSTrt8ZzV7K8s8zz7i7/SGRJR+WgK30GTEoSTdisP4gX2HJfKSu
dHFRxO9WO9kDyplfqiQjGtDF2sKciYKxf52YzWOP6a45gu2jSF3qa6ZgW3MBzjuy
wWNEWfMN8havvsjkA2oaOe3ttTPWrHFininpLHsEdgTR9lC0ABJbUWy/A6L9HPYM
a4fJdKM2N5Q6JuxiVG+9t0TwbwC5pYS16JPEWQ+IcRQfhvshki+NlYZgtzGATDSj
f3tnNWwkZga9eWYfxjCUQBSo7jBNNnGcM/+sOi3Nc3OOWYh2pV0IlGSvyaCG02nG
IQriSZ/+0DPOx/8C+H2NUb7qGlu9tud/f8z2lFYa0i8MIct3p9e2Icso/ZW7ZKlU
OEQKdV7HRQ+UkRK3O7HsUjHgIcwzMVkLACaorY9lGRgqiANpLPk38SRaf445NXgn
IiXo0otRYILrHKdf8WvK4L+8bmdb4xZJBjLFfcG17sDBIbZ7C86LjWa45zKbLarQ
IvlBChhvnNyzryFrTgKNsk6Z7rjgxl/uWRL9uk/rgONjPTenjJ8yU4Mif8Xs1YrL
0f7DyJViKvyzgKOi9P67ifqsU38senucufl31HFC3R/NlX8ZKiefPW8xF4ye55Rr
z4cj1nMJD9Jw996daDjDhg==
`protect END_PROTECTED
