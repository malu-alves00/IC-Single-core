`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
E5VRnmLPH2nrJsK4SZkf+GFjevlW3i28jDwfhqItEuIdmFYviYIVbO4DvAV/+UkG
kEHy9z40dJzhrDcGKBG4kSj1H/Twdc3rkh373MShT0rzt5v4CFBRdBuWRWbEWmKG
qyoN+GLOogoUUKXZaG3AvRuU6R35TRYeaXNIpAMvEmRfpXgAzUwAwxaL57WeKYfc
Q81m7HztHKl9S6kTLSVTHWsH0EKQUCRdWfSZqVX5iTnX0mMC8JR7gIgc8pjiTEjD
2iE8S4S/Qo9KWt289f6Xqe5GHr8rMpBo4EE3XGwT3iBUkGk2I8P4yiW9zrAnhshK
c9EDbWM/jwIgk+7xPvU00jna5uqY4trMFGcW3ED7JA+2NyB2FWHNzewGtSW8sCnj
AZVoUTPuNBqdE4k74+aRQgNmPw29qEaDEQPhdEX9+nK0gX52pbb8n8uuoiX0n+eM
rdQ+uUGM3wuYjsdpiBrqtTgPNeyk9T9+67G+HtiuaIYV51gSdSIslDi3UzIICE49
SNFoXw+7Q2SuYiUumrQFxIM5k66VRv8YtaH1pgXWmvPKFAVqDih6Fhv4Xs+FI9//
c+xHjOSmNuWNlD5rMsZYjM7rOwzvrKLLL/yfbQ8oVKmuib4dt4RiDZgo6Of4o5+H
Ep8hDDrak6dmRGgodNMFuoHDvA71FtOAABbDFAN/NzX/YQudedhzm0fj/zoXMyLR
wopKve1BBB5SKL8NPIyvldJWdGiGNzfngojbSqVa5lgpaNuMTR0fBinvNGI9iyEr
fCkjnqhE8d5iP98PaEVvYdjcinIflSyhzcAv87BSqKJ8gEDjZUNra1pBL31Athge
P34G6KeOOMPe4B+4dGCl8LUV6J96ekczBF7z/WD8MKzt8pSPSbyDJttGPW4rRQFl
HgbsywviyLF4OquqvBkB/mobg+NjERTg70lg5aRSZAM1E2gQsfm1huAoDnvQugOn
JXNnB9n5R5nKXvJ3OvFIBia9KfdZd7JA+lXM2yd1pfgqtHR8P6L4EJsEMJUcvmTG
wRVzQZmRh9KEnfYC5UQWHIgCIf5oLqgOxhZh43MogE37307gaxqYnm62/oEwzhqW
LAv+HkDxWLbXa5IAHD5d2k1HMscekRLMXNKoz5y+62rED1/XkIQY6Nwe3NR7j+y9
f81xIN643V01hq9vuDtm2fewQpQiuI/89qXZBVXr3/bl+U9NF3EIBPj60PXHnsz8
v3+NlnQuxv6Ek00Enj1Q0WfHNtX2B38kbFBQ+KgevzL+tSZyJKiPlaiEK/6sC174
Tn4WN2E+CdVDrvEDwHKh5VvphBDG17ZOtRouxrEJo1nwcz5kyhUtNjdxnP0Av60/
f6qvEuiqUu5+4Ai1mbwdaNV5rgj36zfEluPnBjfg4tF6uE/9Pht8CRBRqXlP4sJ2
PuNsSzqwPF5jldoh61OOOVeE+sQWOjYWrujdMT7Vt9YYdTu0JxX4Rq+QbuWvIbMX
hAZZrFQPNGsvP9UjIg31zPmLmsjY5dObBGEfmXOubjbUFbLgZcKJMtS+QwXZpddn
ugvYZknl5ug2TUK6GkqHnzJaFBfYfPxeCr318CPhwH704Pi4YBcJpDXgbVVIHUvx
F3sTP5+yk7wRsS0uk+MaXWxXC3EWy5NbLqA3hvJ3eN4gwTrygwgBJO8udljdpEbW
Lc+k3HRPdX+ezeffcOD1Mv7r10nq2wNYzxUCGR93R9ZmeyQ52IK44J7Rvi7pyUPl
WfZoExQ8SAEFryaPwE+mG51bNgukxKNDo1vIzWhqlS+Iam9xcXSmkgaAX6SEUwDd
qjmWdIGHGTPiXzcyevj7XUAJUgbmr3ph3X+95CaHRv85TYZ5CF72/1CsZZx8plSC
jEuS+3J71N8Iw+5DomHl0/sBeInmASF8USJ8FSShyJw+oXN0pwIILvLNTtIqxOMR
yi52TNlXG0NzEal0mRILpk1ZopZAB6vLIa67tojrSSJtc8EbleIy/TTYK56/khVb
8slPT8YqpMMs1C9AgVCsOVtFhOcyjXxQEaSG/M6uZNveCJGCAZzD9T2LiMFmRnpq
obu1ezgQ9EBYgoYZZ6UMI/ejVj1T8GAooNXP7hV8NjvX7bkO8PmO/Pj3uind6i55
IA7Hx/ge15QnK1twBdr4GEVoVzmrtb+K13F2ea4EdGYzBpn/HjsQ2uee83gZnFcA
yHUf913LIWwVjVlR9mcw3iyURQpMqIqLN9FrP4R1KW9oppLBhJfMbPe9UIy3cwEi
nz2VX9WaP2TLeTWb0KX5gYQldnSlX1uv6dh2w/XoNmF6FGPEjnmCRcW9773szCqQ
nDYThFIroBVmwQsEc7Wfsn9gPqw9tUG+TjGsyEFvVVMA4775HvWNFrymKnQTE76q
cX4oF2TsoqzHUqwvcM9lp1UzgcxGt+3c/ApGAtlLa2f2abRA9z4W3H3KgT61qS8o
bW7T84xWaZh9lED8SIQDtJjCTUJGIQjKkWHW6de87j3SvKPHcqEwtfJ3Jsgqn1c5
dO7gqkzGLjYXVZCw1FUpg1amCwwobGZYP90Km89PD44NYxjKXcV1YFzsk7Worpgi
cPBGdv+7PPWxkIrMguMJz3rXIfpdEk945TyH7dhoq1qyIeJHQrZxoQ5VQoeA7DsD
pdY9L2F5m6jWXZsJudJm1H5A1wpzrp7BnnXrvA6Js/YXJnAzTbEhhs7bg52nttIS
131GnttjGt/wQwZfIy/+0INTkE0nefM0SvIhW2MtTEYioPkN1737SWVsN8BG3nN2
aGhlAUZ05cOKF+VZSTMgjIAaibDMVpc+JhXJL5KriRoala6uhFO/FUrt6m4/a8Sb
j8N24DSunPHD0TlbwSaf5hNcEaoTqB9r6bsOAykwe8ZNgDs+VAoEs68go/QxDoqE
PemxFtzrDBO0hCKuOshYljsqNYv2mUZIDCK1KEPvzvM89FHPXd3dBQszl3oXq9d4
p8AXPUbL0qJYMQrbc0zM2QeXgU2tubRN/XRR9ANPZup3WHFw0eIkcv3XBJwQXxkT
NbEVPAZfm1oNXjheWSrUCuyGZNanxdrsYImrR6/L2kXV12RAE5F4VWDxeIXiTUmW
u1rA21V+O4rBtiowNszR4nZWaFStx6fh9xIgYb7P/09Mpjbu4z9xOJ6IgX2Fri5J
Cb5/PODNntyz7XgpCrb1o1S4/DR6xlXBRZKVv3ICnBroEBGsz1MRTjpY3CLfJhYm
NC51WMCCTUbkvyuYAKAX0nRQOS6YFdCeOJ98UnfsYxMrtcw7sp2M0I0xSxBn04X/
CF6rmQ28vfQ+k0pSQT6cHQRylZ3o3AwkXZaM8PJpUrRXvjud+waD2BHxMECCNTE4
qzusjw6lg/thqcIDj28nDAzQzOr3zm7919rre8yo4n5FnOf4HGgb07/w87niushw
eYUQBECJYdf5/0ah4n2ZgOuZ0LPWhxnFKmSotUBX17SHttr0+echIL5jW4+ae6XI
nW4YV7I4LHERPwUyCusY1kNFJXbXKWV/Bb/GeiXHSxKQOsNKsy8W8AfsRbOl6M9E
lFioUZ5kup+UdrcsvhgzIkWx8vNjQGNkOJj6joWpz807gAqSZysG3IojzjT8MTp5
IZogxVxL07i/G3dyCJKSQMBfryzqn6LWWsfpCw2TXrFycnZWH4fVznJW5+uQPoHG
LxhExSH9XKRhgYDDdxQwnjpMJzPKKAA9YYnRAUR6POW2XNvdWGYc7nrICPdcmC/f
xjU6Su/oiMpZjPk7srCZEChkC2Fc952xvLWnLB1pDo7v3d5IPkH4/Sopdxfl3C+n
+fNKgOH302oLUsN28eZ9Yukxrny4VDpdXpNOR5xo3FPsALSrOkEgWTDc8cysGNuj
BZ7hACHNnJaA1Scg7cAqy/GezCxgQlUpl0o0aZLv2xFGltPc5KaB+fQaWymWgwEz
vmRDVKgVXN4DLX85lcJ6HjSIog8+n86L3j+uTgRAue7CBH9/QMraFNJL1AmIuFAA
EJUxL0A+Duxuqmfb+qqAKX2BJtkBxzp0GttLVj1hlVDQ35X6QeSLG2BFJyW/ALDu
cqImQgPe5JIWUX7XKOD7xfhDm1z9r02u5sbf4fvo3bxP1LGhp4WWzhLcl8C1useB
p6CqRc2yvYH4IgmrtzXpTdlnHGvltucCPWyXoDbZf4IIwnzGgt7krtK3JYwPFEm/
sYLQDTf5TiZgVcTZEaAuWY7WRddMCuUs0kAzFBdaW0KNyvZhTmItkspyUBQossUt
X4/kk8JLmZI5wT054bZ6SF/SJlVR9ukPK8mvwnxB2NlqVqc0RRq0VDdIx3r2nYZA
Mep77lQsz+wXk6iOhRoIadg6HDgGW1BEl1nhEy5WJU3AlC9YxQCTVdZ/yxuY23SK
3CdhD0ZkEEPwgCe1LIc2IYX+t7YZjWla2gerCV+OwUQ+QStjgDYuz6YYyQXmf5W5
Kyp8r6U0MUV8owu5wlQapNJyWDYau50rKxJ8tIbp8oUF1Xc72Nqg9EbJ6VuLNcQU
UE6f4c/bqLo3CmqUgwTUfkpEVtm75THbUcmZe09+gJQqTZtFVTb0FddMv2XUDN4h
DUfjdYHASBKAdqH+KlBtx0nNgKI57th7fabbfQ/J8SLzF9InzjjC6f5BJgcmLmUX
YP/5Q62r6gLMJn/LxDPqKC5Bopa/2H9KkOJqbSqfR711qLl8rTetMTijJK7K6PmU
0xnEttu/8xBMi8mS2CH56RiRGsDf51KWO3EhJlbSunlo9mANw2fBAfQ+j2y8uihG
mPAwokmi0sKvK0zlKzHAxDzC5FLm1Xm15aIzEjMn3l9xykcEEFmtWNPA4i2n82e7
6DWTpC9WwENp/prFuL/Pg0mfzzSKJClafSs2Nu4nl2TRU3l9PhyNceVAYOteiWP3
cuWSX7yqykMaqkMlG6wAp3lm7y1rJbfDlBS7dh5kfso+GBsXGj59s3QIUlp8bbif
aYtY+twIQm05l53FDqFc6/zvD0CUptVeLm85QWHueZUyjyT7DF4XSufGubdZ3Cud
rXFmblaNRBiILHZiSihAHzkHR4ebJaAxLlzub0AxJw5BWH6QH4fr15Dxx7XwHFQC
t2MNyQ/rrP5VY/W11y0N5QyJzwgvIdp/IPSdMhQUHwGnevYMKhX3OuWW19MWa/Uo
peh+5qwqLhfq63NhgrCyNHVy5AssHLszXYrzRQ1hLW1Dd69ugAldbv4o7lgjdGSk
C2rmGf8CadGjvdguGLBIPf482jojOa3847LwRWQtbNIVzECmocP9uocs9tCoKO7p
3x7c3ThaoRccfuqhXSXB2+3IpRRfWAKWc07P6YsacjewrFrTuLPHzbSOX7ztrSe/
lq9yOw16ZgKIzcowA8bwKbe3Hna37v3nOFnPtsKE3Ytj87N7xJK7ayywUdpZK9q0
bTeKI0YKXmXo9eO0wZb4py4hkcV4MLc+YJ0rJMm3XKjZahXnCdVUDYYxW/KqN3/2
e+zyFbbvXws9c3CjPomOdQVXvr/74ATxUfRRUiNfXBWEQMsPppEyrLzPqSjV7WT3
GqUrCw3T7C6V7TSCQ1qG9Wt3YTrbgdaafXGdjgLh4L2rwjmIPH0p65R7Fj2TPbYJ
iNIJ8OPdWhH11fiYcyNisvt4trTJ5qu1JR0sGrpO1qDcNKZJkwkPlCCs2KgvHXFr
4pzV5NhLLEUIcgUJ5jgutHq59XFh+gH/7NFesT3jE5hCqJY7zYrPgk78A8dxWoBf
By2aFqvfpJtnnHjdDT/dJjFOuAftaBt0hDM3paDOs5OoCquzTmD0ENM9LN3xnEsl
kmr7bvkD5317oWI9z5g1STbcUVQ/b3ABJEXrmg724005+YvKFybfX0BaZ315I+UK
3ta275i5+LYVUJkiSr1yGYme+PIoVwQWWvM4XFX0fLLR6jxAQtsRpxtvdvTYlVh5
RTBYl/9lpmjW2kU4BJ6znYiVzsvQykJNwAtyykr5tZhrxln5nGGg+rkGRrlJMHlh
Rq7u7JeQxF39N6t9vNU+0u8zSKQwDY+R0aRvLXsf9isS4xF147g/xbNJjsiXmWqX
Da5JarcLt4x29S57wHZywx2cOKi4hK3NACGogI23bFvpc+DliOt4C90WH9JJInJ3
jWTjb0B+5wGTFjnPAo73iyMFk4XVHjiFzeDblwVWSE3f9IPRnTi3vDkAAiJnJIZU
fH5lNWmiprnR/PSFyhZRnQ0TkfoJaLSjmGnE+YmYvOEDIVrO75b3EijSL63iMsBL
0tQ1TcVusoGbR9j+PiTmHSwU89fbSv4tbst2vnVRtd1wQgx5tPdZUZBj3b4OMk7y
6tmopMHm1ydydqqKKunE3bQ1BX7nPQWdX1dxFa6Eu391PB1zCOUFsXdtzLW+DXP5
roo9Ejv5NhIzpW/4wgBngraZ/mFo7pDLhZLlLm/O2OaQTU6qiYesweoIkyp3cK4U
qi1kFjU9G+R+4UuIvqyElDCYQopFk/hVtPZPeFYwjZad3nZ00u/G3G23oxrLt/sY
q6Ftz4hMRAW9GchQpWc5DAOawJc3ayvmf3cliTYoD1eaLTufNYl8Zq9Yh6EBddIq
VVeU3iGmhxSX109554rEfVV8KQQVhMRRFErmst6Xp7wDQgyM189dry3loAulXGGv
v4N+TzO9ZTdN4pXhKeedjX7WY5ubKWUBx4OcseBbUy/6Outa/azlKWUxSvPYCX02
jyYb3cSjiDrdHr9ZvnbY7WTvW2urRKNBuHQmnNY2oM3vGdBJSzgGhtgjCcEJMyfs
miGnLA3dzfPTwcRViWqLw4alJ1RUOiEWjXv6Mdhh1H2nGhMtuEZuL8D3yQtY/dIM
KIilp+Q9nUFgW8hMQXpaH7AXdULd9wiGieHc+qoSwO5QIE+tZcvUVCZSSLlQGL/b
WAyNLsnqc/Sop/pF4zzz+3X7f7MnB6/O2B9nXNU9eB6qBUOX77YInuY+Q8rkrk1V
HGVcV+Jw46dVxQYn4C26MB1icEl9wLwHczi02sVxBjBcsVWKh1xJERAnpsJYGjN4
YnoI9h799zQcCfxTDa80/4CLwJTFLWlhQa7z5NhpNl+IElapRkCG0AT3hVuhRtSw
dL2ueQyMooqgpz2y108t6w6oylU6gkXQgpee48IzQw5JaziuqEiXWk/ayew09NH3
10joXfjaUN6KJ1/S1QiADy7GsWSWY2VDFTaYObxnJ6ZShykXq1eHK61H2kO71P/s
mhdmEcPUqoEs6syG4u7Wo8Cl6rLfGvQVGfu3GTe/Ed2Nn3Xa+F0xPgQ3ZPZCTvYR
8X51Rak2mrQAu9A+TZ0GWa8aq8XO9LKPvMiN9rSQmOx+0HSuF22reY5Abp7vWeDG
ldOJU8cpF9x91kM7ykTUj4QePiucIo/VmbQnkfUm5VJ5njXj9Xl83A28Ev07W6F7
9t6RL79F8ePGris75V3koIA8P7U1MTn9b+nJ+aLi3O1DQ1I8g5eIYC3QSvs8a28b
RwnHFcw5dVwDkFIx2Xj+1xMUGehQsALjxLnFDEpxTb68IV2m6288+H626N59Dd4l
Tk1iVf8nctmYNeAf/Wv7eLpaDdDF/b2MnmdTY5Prsba7oQiFwgzFgc1WmWInqG0+
Jv4L9LJESqLqa4IEUkt4oLjH+oAIMUY0vYFm1VPqZaSafPMBnTU6JH70/vbhA+9W
TaOadddrMqpOg+tqIrw9YZpiBZPXrs3bar4ndYxO13fT4gM2PMmqK5o3r3f7xkOj
dk6hqM3J430wqg4BJ0iYZT3neGaqrBikf1dPcq/Q+degu3ZO9HgVae93DM+20I1x
bsgjyb8DXed0UfF4FCo9esHB2UYPExV8UkqB689cGKNT+9FFNhxsSRnKwnZcH+e4
ovt6cSnIZ8WPSyyJ+DB+bAugD8Iy1LUw8/eOwze6vdZ51y9PmQ/zhF3EdSZXB+yf
KSEAqVghUEZ8Fn+MMLkYPofuk6mbNclKEOWd+f184OO3r8FNkVJktp3Rk3PQ797y
0VMoxLJdLp4Z/rn+vL606s/ucAqpcewXKTx6OzgoHekHGBIHq+MtLNVUuy3WvN+Z
Z4kAortP02+ik+tM3yVNnCRgdrzMiCsqV8JinVkBC/xLtTsp+9Vwbylcy6VzfiNH
WxbNmixYKXfuxKaIl95TskWah0njK4GL9r752h+IJjzCG9MGkoO6c+YslMJV1FYZ
g4ma+L/3VgusCWwel6JBM9mzARygx/2Xbmd2Gi2QR2ZrBmCDRtYdm7rLCmorBsn+
8N/KSGKnbkEP15yQVc1tSDTJkjYjfanZCWJfQ+wVf5Krl7Z77PJDJimJUA5qn546
rvS7Jw5RSVCesIowN5/GEmOsI2yfpUwmtUsForCw11l/FrMhza1lhwhdjmo8P+LJ
P2T8BIB/fCWzZfxT+tP98Bdm3ONqYmBOD7J+MTfJVeD3aQeYQPTy8duy1FtfjsBo
35zN8/4v8UWe2ZoUna90vylGfIIJM9Sl8FWEGLY/1pfq17aa9gF+36hjSA20OZ8y
UOZI1MKnCy+B0n6YYfqWPObqwBjkOegO7dDuzYLSvHGa1PQRxJOKNizvsdPRMKQe
0q565SK+bVC0TMAXavvGuJ/RVDZgegFXa/UEfFiNChlNpjr1coEMd17xYhtdzdzQ
naGIvvR6zP6t57aBnNtX8Z8dRTgF4x/RCviecv+ZZh6pFaG9YotxdX1DcNWMLPXA
h+nFRvqau+9Ca2hr5DLCr2cO3G44ows1YGQUOv127vXSn3/+J6my1DqBR2Xw7QnA
kevviXZdlja4cP+JoFV2ULyK887y/JEjEeWqDLFjgs5hRAbZHYc8VxQt9MQ7MzhJ
D/z4cbvDBbZGMj19MgPYEgSYb/Fiou6AIkPBw5O25K2fMW/9MKJ/mGnj/Sfxs9Mp
adP0GKKxfsgsemqNWYGFQDxiuR1kq+6c+wwVKZSJa8sYYNtrVbOhyVXOZyx5h5Om
+wPmOXsiNFrSPmvk2XkiHx7bsbaKcyupNCxrjOcHhlWExYFPdfhgvse0TsBtmWuO
Z8fdRVvJb9peFNBhaH2RYey3h07FvTP1bzlTGsq3l8njoOQaM7X27zw0ZYtrnGou
9OwlvyiejoZ45N42CFBu4USd3Dctyow+k00zMXERZO6XFamwGImRRsPX5FL3NhCg
o01pqYSzty10zIiFyamNFTJXFd8eOp5X5UdbTOWj3AilrkZtq9RGmwBAN7DwiAj/
yIslSqvf334MMY8kCU3bLr0NESySjaN4XRtGuqwHyvJNFUN5azXlGs11I/oY/pYC
XXNKXRAx5az0+6Oj0Kv/alkp7TTgUeRUAaUYRibLvIqsjv9YPdL7JAhf5LEusR6l
ViHQ8NTmzrwGaWu9STaGo8Mj3d2uJuOXWMJhjU77h1/yaAjDTMuaSbmvof4U1wtW
5DaLzuW1m9QEYSGLdlo2Idwshareq4zrQ/yHgxI4z/IKFjFcernQ9VKAkdT9OuX4
OfrQ3Zp4XU1jr8MI8zxSsahWvUJtXCdidGSG7uICFTHRNjQ8zTysE6J9lyKRVLk5
Phirwzet0Yc3di/PrkY8CCvTVtbVvfbP/cmKwweq3QMFC7Goal6tQWSXEqUcEnvg
cg3paIJID1Samenj6xlgnCVVLr0k3TDX5JxrFZTaHcAP7nYDCF/yO1LMgxAE/H34
h3n8NQ1gtRbJm3qvkxJ3RYU+ObCiBjx86KX2O/SCCeFQCdj5ocyElCp8WOEXfLuY
Sh8aVMlLJju5MGXPHH2G0KPH1JanYCGorIjIs1bp2ssCmu36g9EO46I0Wc0SEjkR
jQ3cWmHtG6pSjEGI1i6BjENyfNOk7xT97nhT07wEdL1zYctW2nPs/w3jykkKSAL9
/HMGPzLF1N/CqRtyWmGETR0mdA7+tdPoZkDWwoXc8TWVcqCkmzswXLJurD3of4ap
TzMByqdNbYLSB9bI+JZl3Ot9IxamVPmOrZobEyLhFzlELq6ONmE3a7Vztf5qYZVo
CFvc/wSiQTzwEhAw1sFPiCi2tP/3CJqTUCZxok7k6KHT5l59vixujHob1YbBkWoc
jTvYuAMdm7hhrow56K5yLj14qdaWWKDCerklViZBROZGRMAdvZoBEpEP5hWZ7WYd
6zl+2/BKnGKsassweHRzmTjYQB8AoYObisZC2XN8sC+t0P0/6A3vFxQYNFuAIqBQ
R/Ll69gbkpGpvLS1DnpUsj+ZNyHFyQaJvnqjZmaWPqKoXMm+usEeEGEzuVIT1P3s
NKJ1Q+sU99uj2av6e1kgSmElvmaFN4/oHPtgbUwLvKgCd5uy+HdnroMjyl8PHn0V
saqstZ4J2O/vRujTlsvuk3D73xedNF773L1oMoJ0yxoGGuA7cqhGIRmjU3ks0YVp
IVPzWEZDpViCd5PF7rmS+zlwo4Po5/G3yHoTf5tAlnbPFcP5eamQNiIv8EwOeJ9f
SI78me6dqOIdcTaWw1SbZnzl1+Klya1ZeH3W+wOpR+4YGCwSxjEic64aPOJrN4hV
ZbGfT8RYqvBIqA6hwFK3gcNGiSPQBJKvTgXV/wgcF0mhG501BGdf4gQNZ1g70/dk
vwqLfLyPzlFndqdbIZikaKz9F/nJH/6ZdTBrPXHSuPRL2+/326PqzO3d0ZukqYoU
cyN+UwCQSgK2FM9O4BUfsQ8LUzgHICuHhO3Tq/CVyIw5ml6OJRmlL4b+8x7BS6D+
jbr4Rbrh/Kg11WDvzoKTIgDdaEAHkPGwtDmMK/2x87Xi+CW547uqQ+tRYqH16xYE
xWJ4G2u8Xe2vjiuCDo7EJ8sKo1PqLum/5Xf9NqYpfufHjTdiLmji4BbZa6mAN8bN
/QCKer29H+nWiR2BFbo75zIj4VEJFt2wbR7EYYW9aFnXzeFrd8QjDHmy9C9fgkRg
1DLV80n+g/9s6O41Cqcx+R0OhvcEGeti9H+tETB+9A/O1qLKbJEgVy7vRsd6Uy3a
vZSdXaQc+E9ETErvhZwV3TTABpJ1HzA786VEKZXJxw7GHY76g/IuOWirQlLKlVhP
pk/V4Po13B0ll37LQiQFTMzEg6pjiDaCaz+Ztjcfc9nqn0hecfSsWUdW2WcESN8c
bh3fSYdDG8c6vRVhMR07SFgaJLR7Ul3Y1YhJKrrzrMXE3yZ7vMGtL01ikspWMM+k
v9RB4p5v9p0vF7ffcxya6TYvunk6PEY5kBtfOXD/2kFDGDtfk73Ezl68TdnxIXhT
HA+ER25kIMDTQrlpixp9PhK3zvun7C9FkM/IkbQGJWqFMRwCQoltrM/ub91cHRg1
sHf26sj9XL8sY0OLEBuVGk69YQBifZqH8GdXnLX+0sY0MUc4D9Jr5sU12bCkgA4M
B9ihUMwRb4LIFwO0dA3td77NEIGjx4492BntlOtSVU1htr2ocMtrKFNZQD1sSiuk
hJcHom0jnfKbpY5vhOnxlRGoPRdB34EO3OAY6UCunMj1CKIq2m3Xc4MrC+7gHxqY
9Knd3956yEvTFPFmrPxhMbSwLGCEGchxxxhieqmofig0zaEuKgN5gZD3UDhjRHpt
M2DNE73OJiLB81DqZjYWlzgw9+eCOMxqM4UDM0fcDmpgswtWy+kgxbfIuRteRoN6
J/ssA3eNlPcj+wsAIkHZUj0CbSZQxnndebIzt23KB/8+TTosbGjHlW7wi8SdJcyK
3dIW7MnJrdGnJyptT9/hQG7bXqaPnc1zJLk0JoUFeYdalMXJq0KqKF09AD3MV+hy
XBO8tXKBQ2YmLC9QWgVfP8Ju4GC0KvLoahvTWHCu4jTD5LPTx1kOw1HkXfzs2ca1
Y5yg12Hluh3wQZVOtEtbc1Mu4Tu3BH+jv3iQJ6jUdS9rUHrpg2xB3mqPT4acPXYp
FEaQ12gmfGL7WD4iuWA58TxCXj+liWOO/hfUHIwNU87ssGUcM7xusnnwSrSCUFom
wd+W8vj7UcsHpPefyZ1C7k1dUF66mb9K3eq5VFLsAisXa4J5Eelr0A5KmNnBt2vT
SRFMSDhWf/LP6WcHd8fuxTYJ8HEOkDNzgrFbBOfrbgr4UP211qN3oxppZiUL5hIk
9gg2p5+JDc5KmcWFzlTsHcJ6uPxzd+tKI+JFRwMMBhyCcT1q6sIDjeFDuuzee68v
WjFrdrHODLYs/GcXkEPnRl3g6D0bYovqhXN2GrwyUf+9brEfAtarO4RpEZpdJiAe
E74FD1JUmpbhyUGaaiSVM5mQI5+AIoYoqFmnFsPzv276ZODjhSBeOMS2EWnwWCXf
iRUR8cuUZvn6ep7WICt/mGHD2/h99BOC+AiqWXiAPCG/wsFQpnGbfaeIEh6tPsNY
Zae/stqARIb+nmoZVXZ2hEZuc0ZMfJwQ2A29Sjoa09+WIdMTrAFlrSnLKRMsoebx
x+CHpLACT3hG8Z7yH/CgDR/k37QWIWRZhy23N87jQAeS6BFMtpmX7sx5DJRyJr6w
IWyUuybCCQqIHejc3FKUnYbpYbBuH49adu06nnNo+X0zeNr1CMZrlz5PsM4wkpZl
CHWAotzVrHdqvIYhmtWEHwtwtSGJaBzgo6OS8gkOETdOXSmdMZdMind3TbUBuf8W
MBWI1fnfGXTpgZX8eomILHqaHsw2/z9T8fZqQHTWDG3+AVQYmjylFu/fV59/rUPO
yS0QcGCRWL2cCIKP1ow0Ry4ZnlF+nmLgjd7c8EjiMIeMcN2f3W3phxNFcXTN/Sx8
s7r3M64BaX7nCL3kjVWAMa9EHN147hRm58FGUuQSZO9aVUBCOHiQYpYji5+oACdu
EPsbz7BXjGdTAvih6STETmzUVm/twp6neL6cM+jk4KEWRdb7kxWO3/xzCyplULOm
iIYOGbcu0v9clziKW18hbn0XO91mIgCFfb/ST/P0LWosUc245Hg7II20wr7GbFBP
ypx7LCkpm4FCP1cTUiCa538Yhu1ZEOFm2wOaEl+o1NhDDaMAx0H6VddNvIQeQuaJ
doPecAXAf0GMDpiXIhuXvK4pBT8vIc/rENiJpNX9Hgu5lIooLJ9lT1QFM+2Se/xo
M55xJPp4oj+Q2hr+0vxBBJFO6MGEsPtYXXk/9XAAyQvTyWL4HY8TaSCkK56VmgGl
lI6+XZqx+474pGlc1PqASrPN93XQeVm8Ck5t7kHCBjHnyHklKMeXE4douFzMHDz3
Jq5JhIuy31M2oVrVG6cbhiwZy1TYxJV7rLE68BvQJjPkwZniqHs2zVc2x00DDOdD
EfdaTy2HWRn+fD6KwHmNF/Wg12u4qight5ebBlsOhxcPgA6hCsSTQZ1zYKkfGVQ5
tmxNP2hS1HrNIXHGdAeZ4obNKUHaJgs4bfDfo9aoBlA/W830Fx9GWincfbNDHzha
F5oqRL7PsuPJAf4yQIisQvwxMpwyrZMGpgxWHW0BdKRYApSfVlWvDIZlpXxLi8VG
1oXUqIDwo9T77AWll75SWmeCBXeYRwDsjFszXMEgojvgE+mGF+MS9wZ+4PF++xsR
IZrijzOdr1jNaaP5oGVtTOBTlBBp4e4sq5o8GHzMjiqUY3a1kaa8XHIZLqlm6nil
0uBscGOew+Mj0r43b+DZpxQKaUdBbp1M4TBl9QCCaiHL8QQ5zbRyZJ5KHR/w2af3
uc6fkfZp5MmBfq6i4aVtV5/VvLvg2rRfOcIrIYCsCsAkJJvP3pw6eMwKkOTMWqSc
cXkT+Q5LEabYM1szUIuDnp5ad9KaGGJ4flIIZcga+OyDy/UUuUbZPEcIHO5A8OXj
OiToPFSCvK8b3JWK0cN49AB7U/SIjPQFCXyu1sK3KRg3XTYinnJeNXq7jrix5bgO
58E+XwzXxNurAKjiIxVXms1J93zryV1E0nmk+dRxsFYFUXgaQLp59lBIF1NmOlPe
6idBMqMg1teRrfwp5tgBdX1lT63bVBOBLR6pQ97Gyuy84h67A3iHVwTdla54e7Pz
Khx60Y3k/sfvAoaQhPcs6o/U2O80UbQ5F+BKdF+RTfTXco40EAeF/XWcRIvKRjyb
P1/mhZr0jYORSjQwHg3QsOaV7lWhYnr6ggBxqL2p+aX5NaSAr0Br2QN5spL9RQcE
HolTFdGmCDogQ3LOc+W7f5lAvOof/xu6zlpnTRzjJK/CyE8wg3/wsvbwsOn42QAZ
NYAr5qk1qoTytKBzx8WxpC2FekIA3BLv4RLUJUXDAeh/V0anGbndf05mODaSj0wr
FSTBjCyvzs3RDe52dDC8W+egxZRiaDVaz5ved587dnGc4L2jBvYrXV7pIarMydAA
or1HcNPYQi6vD6Fe6YW8r4UiNd/HBETeNQn4PNGfI356suXOgtDF3+sb4WGQCq3h
8SR++yv6mpyIyrqi035rIMgWe28mSsDJqC+jqTKlMuDn5IirAEU2KAzBIjr66jsf
sNDfcbn4kNvX9IbvaXsYLUo/M9yuKdkg/TxDp1iFJvAzDVBpcVm1b2VjT13lzQwg
QvZ+cDv8D476JUjAraIkVeXfZMJToAxw8r425eov/cjgB2Mt8UjYyyoixxKzO0ZB
SrDHigSQy2MKTwCIjsL3ISbjVOXSUCdC9tga6Wm0n0bnWcUs3ZMd5VV9m5wQzXm5
S/+zrVCctTuYX8MKNxazuP31fxovpzNXXxC211eE5n8kwdiNP9smkFu8mpZvv6t8
p8Xnm8BXvrKp0MwILIqMmZi1dMnRdpteS91vRsW/kRsmqs2i0uTwn4RopGNmCrRj
Phaijli2f0q57QCAS0+AwsMJkdGWkYpAHIOH4ktPrpJcKH9yN4xTnU16Q+RoyPUb
R3EteM7heFvCE3QcwqFaNuZGRot1E+9+wfe27XubZAoJSivE/WTbWPGAJzVUu9fc
7ssoHPUZL3j62VeEQ9415h0eGfxZElOAZs1pUSOnuWE5JDoQxbKm/oDql1otNFDJ
8B3H5FMt4Ab47wiW23XedSNKmykX+x6SYyOuWvohf647nDXOBEW3NqoRmIVamNib
XzODdCKgieBjbVsfMK1JcuQh8/rCdYLR9NMfmBuKUM66+bpw0bpqI3HlzTok4u9g
nSUrT3RRFJWOLfwRU3CUSlXXCGgLtEwNUghww34s3N7EwT5im04dSbT78IPuUEHz
yCUW7y6Z46G6vYyOSTpkctCsyf8OQ8MzHmhVG2j+34OxsIZ8mw6QNERG3c5zyQqN
jJD9lHbYYn+i/9kvHqOEw+HE0ZlkrzfvouIt2DRbfSE3Q7YfGDml/6NgmCo0hHLI
8jkY+RHt/Op01nzBxoI2wKxr5zmbuesv4hdgvqPisjN+LsqZVlPG3x4+RKDz6C29
1bojStC6nnUxDer7kOAO0jCf345Nu9PlIsgdUdWy7EryH6LsizJNhDd7hfrOlPhq
VzXNspIcZs/02g06FB/TI7cZpxkYqPGnmd9ya/eHs0rcb9I++aOW7XXbOZD8fPAC
1R+GxOPEPcM5KgHOSBgKd5eB+GLp2GfAyXbpd2aPAw6+KpF0i8U4pBBkjZTA8Xqj
cPBvsKM3y6Gfk4GYaBhBjXy/svdAQIrMltCUXCFXHR+sAwfEyRTU+DJjcQZ8/ysY
unJH4Os6PBumNhP0i53XXKhahW1DaVeh5v2ypM+uhNNyx1JCBHv3AFl3U5ZFEAfl
K6HU7OkJ2b9v0pvg0/Fas5r8rq/wqatuSUOP9JGzi7k=
`protect END_PROTECTED
