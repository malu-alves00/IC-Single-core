`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4irTUO0AfpdQghLQ7zAJTvkroM+SWJSDCs3/CnNn5Y5Wb8SUfa0KjoB6vCUkkC0S
guvnIx70i90vMj5fybf3QM507rbDx0dkcXO+f/6entpbJTepeeR4LkhfwIgQ87/W
VWCT7IVEw7p/UJcKRvdSm7i4V8xOSChay8mYCoW3Y4G1otqMUAKbG38V/5/JkkWB
szzyzzSljZFhRf1dsHIU3W4a6c4LnH7LLJOqbFOMk1KZZ9Z2mQsKrLnJlYe7wcVk
bsPSHkWFZAJT3hvElVxMKrZUOlC0eOBEyB85fEthSUc3tc6kxLmdxDovAGdJBBOr
5HGYczIlOnJY6H87BEeuCm9y/CEbGLHF6Guh2hWw2EOv3G6qlG9cReHu22MRcuK0
dcCk4zuvkAQgZ1q6oAu6Ls67ecRlbBzz02cy86YO+Z314vnlm7Lm5GOaxdND1sAP
4x3l0u7arfo3lS7dGkTzM9cuZBqnJwLkSVPkp4hjgzSmFmalGqmdNJZJLbrMR8PB
Ru7ggRo/zoIlBjg77XdJz923L7h4Mzivp2zphT0Uga3qUkdV1G8Upzh8MXbIvj84
oOUCiCun5c2U4Siq3YNyHeYO1ye1Ss7zyeZWRMlGWFQgLlag7gD/CCc5p8LuV3gc
f45lM3oKguRllr6p4SGcXpA7yvGw+kSoiLGsfyFCsrjBoWGLyebi40US9yexgwvg
YvjeqVNqQYLgZUk/CnoQnlhTBAZpXtJJlTuiCsIwcnyXs7XTR+XrgNYoOO/ulTz+
clQNFsbqd4y9x09eALPJwom7geZqguktXASGpp4QU/t+2oZMOhxtwETp41sXky/J
1GESAxJLkhR2Aut90ryzTU6JqKuqz5X2ipDkFj7rt7ndih/UjJ4wI/y61oLAb30H
jelJUU+P+WzZLY+f54bN2qwL6ynjs2YzDX8vQZVnfeq9dXdcrWTwwriK8TyVqjy7
GSxgFRGlrO3tvfzj3Duagsx/abNNPKdsGrGNrFJ24bRa7TPZkCYoklXUpGRhQzhh
6xdY4muxEfud+2sXHVeJwwweTFH9/gzvFcj//+Y+2G0K2NFkip5iaYJlQkDrr8JB
iJ3gXkc3TbystSk+xYthrLaf3B97x3p8eKeJ/UMrK0ySPzJ9Ee8gkABv7b33WBui
mkhghxiXVqu09Wi0CJdyNn8Qr1wFBPczqPJSWcXTtxl7ZVuKeAefFBFynDi27BUP
spSOIoZ5o8WOeEznvhuQSTveaPkC5/QgUhRNZKE8pzAlbJ/hl+wKeqkrgoFFl0bq
EVBpbFS1fkZWDmj8iOIv8RmDk82J7H2wZbNO6ErSuePuahnWU6wlnJx3pvMQHnY4
dc/cJVznv9SHSCWjdqbr2hjCwkNZgZ7PsMzn8uDb6F0LC30mmkEFmPXoRsX/W+BR
yIM0qFmmsNr6VZOTm1N8GUEFAw3VbuCCZTeDCNoWXxp5eBGqivm51skWrZER0U9U
+FmfBInm5H2Es/9km80ele7geWjJDI7TH6I93PYDO08CgEQMksnBSeTI0Dw1dt6m
0c1vz0Ljl1Xp9JulPNi4RiIwLkpKY3IQJEGhpfkidnzyKMuNYXeXS2Se/Ml8mOGH
wfMnrhsiTYDjWGhFhxb4ZuUMNG0Vhl791HmHfYq5weTUBaAIQhlxTWcLsNVbxBSY
K0k8UXxdiwXGrlet1WiZVcHFvhDp1wvZqwGsDR7P9hO1OVzFlIzTxea1rZzSLICT
iJxCK4kkn0HWuK6krBXIcyP9WLs4MiQEB/ohj2yTIWM6Yh5IQ2+SCUppe7OhOGcw
oRy9pRrAu9/N5CF+aWOWjRwqk0Xsv5eCvwvu79nBVIInzy5bv5om+aPzXV5PaL9g
NpDmqt4fDzw+H3dRFd7NwTFtyjRfDyE7tfX2wmX5KVfQq3k2pymXCTzMGed5dFsT
MlYH8u9fgN2mb8If+3QMljVXxQD7ispmFT++wlAjuVzEmkMe/ppSZYI0Zl8klhZL
5QCrSSBxDFLtgiSKgD1HE2D+GYDPZAzu4TVhz1KoJ4SLqIaaMJX4HHf4EYQLEpJW
jQ0pjcfIijPUjkoPGQR1abBFHxgDYxIlWsp/vJ9wwAgwJ7DcASDe1NIsZ+yHhF0E
u11LdBUPMDGih2KEODHcrg/1/kyvz2k3vj+9DlRYRaP3j82KOvX8njm/Q07kJFdc
K3yZhtwaRoRwEYSjtc4FA4+YWG/eexnSocmOvgM/sA3yudQflSskInsZwCAfjq1a
EfQL8D6PFlW8ccA9LUSVDkQ0yNaxLWC6zec76DdolmOk/vAVpkqJ4ZfY9eT1UgL5
fm4iNmv7Cpqd+sunzCejS8Qe9TyQDJUXLAM7/CVBGuBGNdu+V/WVQfLVpaKCi2oF
EbQ+PQA9Qjr7ocMf0mxxb9SdOY4AZCxy7weN66iXKQpyiX8yUDZb2KrLQRpm4kpL
2FCQQ1UfUaOaeCVBm2sXIOZUc9Mt1UoK1927j0KeYBMFQ+R+SKXvQggJJds3DfaZ
t1hQoQWTjwrhj4z3Ry+rMAnIY/3zQ6+SUZNSs6buod+crWzevnnsT8efl8nCOR52
OmHyFvvHrG14UeadF9GKIsHjFXvOXv9EbYyxeIPP8XmoYP63/ydHgj5/RRHjARt4
m92X8mHJUZhBLD2Yfg5LlDNAXA9OODukClB1k2kOviCA2O3T2qcPXjZeLDwQLoG4
scrLtKaqaLlWqcgyDazkBHSm154oAjyeGgqryu+OQE8IES3wNPh70JHtlws+urv6
jyMoi9piAM3GYZv7i0DM4PykosFL7g1e1KbE0pA5VUNDr+MIClMSPgeVPh9UBqEL
qBjV6l1rNE14H+xfs4ZJ2d098YWnS8xwSKyDjncUZQ41VWBaFOvNc+f2aSIz0N2a
y04BIfJLIaOFZqf8+hP5Hg2/91BXGovFAMcZPBPELol1pRInqoH3zkqV7iILcv8h
htwvZqFsIdgk37X4LR29qdY4KUWxh09UntsEp5OXlTFI9pjM4UQM+rdwojFCdFQD
8IXbgpw/4V1ku9S24OvtYgnKgAfcYTKYw3B60bdaTuzk3Q4l+6Wekw2S+wh2xyOY
QRJTUfaksO36AC8TV4vTK720e4et/UwWr51SC39JdamWUI7LfrqXh4n2jkza32Eq
H9yHrCb9KYJH64i8ZyGItS/dSSMSs0oPHQyhJAZOtlB1pQHpJoBAoMwxS46Gdy/z
r7PvnmwwNOufKYkIdnRuqIDe/2Q6CeBia19RyEbsnmvw3S3MyWcpDMSYIf9xuYa4
rKKvhr7eKfdxM6VOKBdQ54u6yrm5s0f8m1gh8WpDhG44SdchgoEoh7EKkdbft3Gs
UBJWRqo7ZywfQh+1LreujzY8Qy5DhruE4nypldy+yFei/32saoE7MpLbSKNeff4O
oD4eqbELcb7lqbBmF0Ht6dH9c10KdOm4oO11Dxv0zxtBsSHpiRLc3F+BoUy+XoWl
BS6/mu7e3x+h0naREAwfpUjmDPFBZTzoAiNloZEK3PQWoM+xr3oLoVerG5ecJP/H
hBLio6phN1hZIsl0tds8/ueYZMXtLu6iJVLIFh1XnZx8A/O9IM9dZF39X/P9pNAx
vRiYo36IsIFKjmObzp9GybCKf9nKpZz0HnFECCmpNGA5UZL7q2SzG9as8/KS73NU
BVmcSEEgRzdFz1PYrDNW41pe/++Af2jyN8rzL6H1r/3uCiqBBkQ1qq+UevWlz3yZ
7cA4GHSQQlFjYOcAZ08QQA1+gqnmrGUQqaGpFe4OQTyTpHBongpci5Nd+J9UB8n/
5Eks+WA7cw2wNuAT7E6E2Hex/KKvs+fYJ+dUNcnoWpI6rOeGqPtikXIVUYOcJg3D
ePio5F5LU4ks0sBah3+rtNXQfaOBMw06eXgIAjUy48P0pJ193wqvWfjNdxpTFAbK
Bzs9wswsqJAMr/UBzt50qLwatp5aokoJhWSSfuRfBqYUZrAFfe/LfYTpuB36XRWC
L+IYheiWKYDs2AEiO1VUHB0kHLjXmxF7wZoUuF4Supy34mgiPZQ5841qgf3ZMXuh
tkVpZHdmE+zLn2tPz2aJt1f8GAjq+qjEgITT8jBKyuNcVyzK7We2qMUF7FNbTBS6
wPOJw1FivzQbCGtJQuKzoIgr4hKp0QRDhq14FE6f8rR0c8s++RCnFjlsRAuD4489
ekF4o/1DXiWTVl997VTN4dZ5PA7BPekeXoKjJXz81CZhbLxFdnE66D9OC3uR8AWs
xdFlGGtFhkjXBqvV38uHE9xnSMZX/6RIEovG9Cp6iLk7aU19BSNDoqEmdD97nOt7
KoUz6jl9UAeHxeB0hRmju3OHlFWskZOK5dTHfpBsFvTE12D20OIb1J4fRu20dPgV
itiqnyyz0r1THoKwieHXjAeREtx7lShe9xobJCWM8uALA1PDOSGto22MJxC3vS9g
nbak3+SI/SbldyjCXOF1LQ7oJFlTbCMPZbQkbMXCyn2f2QTU+9iyrTIgfjxnL62p
Fxrap6oMYgu/1AltI1tB2/X84MjQjr/y6TEYHGA2ry+94mfI+Opq63rJwPdZo2qi
8DPY2IEAcEx8E2OB06weFnDyzZrDKK0geE0bEt9KA3xHRz5VCf8Kk9Zr1VQJMCZ1
PEjQVWM2L0eLo+dXXtJcSHS7jhAPn4HAxsFHpeSlyZsl1FX5eDqj9VHbPmsxdStk
ao1H+ouGKGaT60uV7bxv0b4JIhETl424Z3INeaprogiCP9kOwI0Dihu7w7Zq/jsp
3Pz24MyJIdtSgwZyD3MWE1GhAlX7Ex8FQrxv5IeqobgS3YjnBGdiJ/L5D19Z6MzO
oW5m1qUZO67GBIzsP+rTsw/lmTDN2V+uxoFksLQFpibXrVm3OyPIBnhbooDU7G9G
E9bn6FP+SjCkxrHNDhhDdt0XCXrOrMwEkLxCyo5gop9C2t4rAz8EVqvsALqxhHMR
Mh3J6W/2tgGhXZx1pYyzmMvo2Ai9UqBq0z8h7KKTVg5ExQokOryGqw9bSM9+l3Up
xYCVorORes0EEy9KP6HD669nFKCZ8c0pk91nGEpZhgs6fAIS/ENsPVlq4/BF0Xs2
nQjom9niieVeSp6g93QLYFjf9sgWaAPGldZ7PED9xR6Iwb+fgZUtEEGjkrt8gF4Z
syL6BNmlZBHVYCQUQ+14I1DjOX0ah1rhcRpwRjyTff4GEQpe5W1Dwf8sQEZy0KgK
6NKsRsM81WkKD9yHfFvHV+ITJTc0syREmN4FiCVKu6RduZFeSkxGMiSmO/KAxfvF
sVZQT+z72i2lh+vmSQHwGtgnQ+TPHWDArLUxR4L8fZplRGWEQeCbIfbKhYgqgJp/
qQOvOuoZX98xf0JICLucboI67qdNdJJ60/IIoqvXfFxD8SXMJcLYMQCKXlILJYh/
gz+TDVtpkcNtKC39bCNKbuk9BNrwOJvXwL+4Hk/Io7a7Y2e7/g8WM2Kj3B8Q8Lmg
BwR3QXiPJ7eJDTCqA2bxcqj0tCwCugx7+54Hpu3Pxd7EDNzhZSEu+fycLCe+akXE
yK3mO20Y1r/gjf4SytDsz6B65ZTkias7RZS+tl/Vc2E=
`protect END_PROTECTED
