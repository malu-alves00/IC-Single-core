`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YmBEVb4w0SK/ec2FMbix2cOC4y0HNihozYFvBgaVOWpnS5z1r7ZUGTR89aRpJ90d
rZ32V8tsVBv8SOX33noOeOrUwVhG3AGUiH1kSiA9k1cyiFtUHzXIcDSS5kV0h+bC
IlhrrYdS+sJBaGHqzOhEwBtAdv++vMbWbX77rU269RQzXcTMMN7PVb4bLmSBbaMP
PiHsU/cHl2BCuTIGPH4341/ghUPKxYx48b6FU8ZthFOI+BdcHrznTwaZffOzdTDB
LhurwT8SPSPuuCoXkz/PgjZBchROdy4hfayxMYvI79tnhY4B0U5MkHMDtTdxEYpR
k6z9RkKYzvdt+j3EU3wG+uapT/1TDcYpGNQaX6g26dwd9kXOx2IHoebZ59+pKowM
IWoguEhdU7oIe/Ey4Fd68SeDgF0Y+rgaal1PNSGcyBnpwtY3da52glvhBjc6icxP
xzNjcjzuxIhZ2+yD+1kryKsa+j7PKMvD41hR1iejUIiqARtzmD4vH1GDFHg3pvy0
FEpwSkL6bFI46QnUGW7224WOtioI7ulHDXGn8A5Sc/M=
`protect END_PROTECTED
