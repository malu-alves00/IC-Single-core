`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
imOpljF6NlDfqeBsA62hAZjCOSyl2tczglsS92B1bDJD7zFbGCm0z6cQJWAFpqij
N0pEs2+NqUZp0YRlyHrAsJqH8oCiOIsImGbA/3DNhomeSHJ/A/QP/m/sfGmjSJxI
xb6KCUDc/tYChwgch01lVoiMD7zQ24fOa7TD77i6pC403Qubui0bQWII3ufHU2qS
uznNyBbZgZrOZWRYthsay/vBM0dhMTc8BSt6W4ug1LsS0uJDsDOWxlnNXQaPjQiD
Uk9qUcrZ5N9Fy1rBMAdAp9OiqL5x31uaGRyitP9wDTAnuHlVSNIiiQnTuoektXBN
elzC1PocDe39mDNxujKVXhPUpElUHSaXkkWs6ORJKMshjckhfP4QmbI6KW7Wh0Uy
jyabQWw1L6FTpUrEijhkQXk7iDfTEau0qs8GaPBVAg81i6MianT4/nmptdjcU8J1
3jmR9TIzMeEZsYZ3lb7jrljg4sPfv0m0efUvk4Ipim/UrrX/+afMAPPns28y/yBr
SiiWaiMHQgZt3HSlY68WpbkjnXErq8kDk5kcuUxlPSzxJreCKjsXyQu4nZA2qxwV
gkvhO4agOaflU715lFt1RsMs896VYg9VzcUVYJQvdffrNdtJlv/ukeXtsxEMaA3j
+AV7y3LKPs9Ma265Z4rf8Ee/8FkXR+49Dn+BgUsRXCScaEhiYo1+DhMvEMBicvBp
GnIKv+H2Gs9LBYt9KXEAp7Cc76awkjPZuvJrjoyTX5QboEmgRj+LRBRDkljuxfsO
Rq0c9a48NBmRmWdJgshhaW2RrsMLNY3IDhuqNvjEjfg4jD1Om+5JuULc8UE6zq8a
NNRJ2/7LWF6G8VqrNLv4nSpwJXXQpnRAf5lcFTTGc/IRKWAbGk0F/1kFB6CHUK4d
w3xlJ0HxRK8Yj7I4Hs91SasknRIJEQCpe6YZkG4Hs/7Z/LH2nGee1UM090qZNTpY
`protect END_PROTECTED
