`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+9iP63eGA6qXethffwJEowdipSxOkxgHVZH/azS2jqRX5xyOnYBVFzsj4A4YuAwd
aRWA3qrZbl8I9tTlOKsloaFyLoFhJV02XezlJuxE+youQsTIGYu0o4RRn/GjXogO
Rl4/sqXia33QPvsTHJcvEHff3XNfiD7HFg0K56WgrW2Rz/BRHMRIPaN5X5jjjGhd
zc6kp+fhhRe+AOuk37X7L1SvQ0WqElZfmcszhjNAhzGX/buZb6aDcUUswmjmBohA
8iQ/jONZiJComsfXRyYU8UkCgVfXs5Txk29BIowDom3wccAjcIa7hi0jTVpvTD5M
7q4LINiq3YgfbZvmBhFK1LGoodqLVgpGwdbZnFaofvWYdCQxUeB3WPlDNUGFeMz7
QNvaQPTKRpudceCqaD8s/nVazk0+JdP1KEcTUgduaU6BGYio/6AwjTcH/+mJq3HT
CxY5D2PJ4YXkLV+wOd5/e1NmXhGZjiq+bsdVUWb0v9A3OmoNi0HzTJBFqPU5o1px
l13p1fWl4Wp/h0Z7AVJmqvlsEXhxw4vtdL0aH9RcL1Pykq5E8YB2LrGs/p3R7qCX
VbK2c2FXnM/V+N/FhlxLaztUr1DmQjKVNgk1Afbg8R5rKdALMybFHrtRB+g1Yffl
Y+bp6IrkEmG2vH/G2JctZpEOAIdIDcz3mTYjA/pUH6cTPKJmDFV8PgnRGufGgMKG
IcCl0kBJdndE0krZcph8LIOPB/V4s5mYHfKUzMGLIKLVgIL/piSriB0N2svyHEn+
DUfW+hLhcqC/nzEi3/4GfPPlpJbwuU+xktQq+K2GQjR1bZmMeZ8QyPOv7IWzlaKz
edfFsM1H+tmMyzVCoeXdAQb7ZqrO56GFo6J/onA1cpfkr2FmQ9p2wVBaxar/D1+l
5CprOC3/sGyNunMsE//krfvarAjBkz72tVhkXhjWu6IU3VF1O+qHVx4vUgrEQ+KZ
ekK8237Tf1ZUqOoNSjKF1b3snxzW6VUFoBmgq4PBiEj/yJWbtAcHIK1UJq+l+knu
ZQ3sjcDalkWL3yvPwBpCFyt1tUZId3H9wtztRUKjsu+VBpY8y6Rd6VAfY1kdTSt2
Wauqr8jDhzyfF/gjgZ3sU2j9v17spTa9P0GA95TMfMZKQg7GbC49lCFbcYaEBaY+
AyzZzB8wWAuv36OpLxWNdDzBiauOMxVZTcAEX4hh7JT7u34FFasYafn7sXp1fIlI
i92wLTtassXeCgYsS6dFeK675mNkoimkJdCsyjn9voY06TNi+snubhMDw8HKIiVQ
e3mYQycUQqC86u72c4/k8xXdAQVnBHYCxDWwLpd3QemTxgcVF+FrFFqsBxGgS1Wh
BdZ7TJHHWBa4JvK7Lo/SXg1Y57bSU9pMHtpyq1H7GqKL2oRdzBFy19uvM9g3yoXM
jyDs7wTV/CDAES8QNZcS372GBXo6NZCxB1PR+YVY/rIdUtihdafP3a1qY2tyeGQV
RIVFmv76avh1172SfhpohkjdXk6iSD6UXdkIUnqqtL+kh/5NUeZUcKu0WvvE8EIu
+j9iJuVqp5uifiq6bttDJGdqCg8O9GdzdH0ueJH3p7p9QeIIVtqA8TgcanNLTdft
DitrpDFyytIM3P2UZX7r2MTB2wo67KRagyoijcQcrxtTiOjOOnDz2ocQUfg1kzPj
PzpR5CUGcJJBiLQGACdZfNoNV06d2LGI7DKLoALQtPWdHCCFnXQOjebArPOLzqFF
lF7s/WVW5L3pcxusx9VtSUFCm7XYvcH6ZRDixZfQE6A9WkijkT6NH2YMW5KMnnOd
vad3nMohRUAtss8A4A0J7mXZF7DOF06WAfI7jI3CDSDmC7W2wym6z48Jo5b25veP
DtTWL3BUbF0eHM8+C0hbjwv95sdOKslNcItigEjHxmacHt3wcOFpwl38xLZwz/+R
La8tQqo/nFkCCigB7ZHBYllStf7J/OVH9yJuDk1H2B4=
`protect END_PROTECTED
