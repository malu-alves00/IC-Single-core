`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lbkubWCHsAwbKBg3+wIECoR8SdVxKQJ7oSjJdduVsjK9Y+bheSGtjl9giLjTfFT7
w6mZ/+JpjI9SEymKXzSTAFF6pJABDnDYbjpq7O1BG/a1LPhqZfmIjw1bBWCUv/r4
Ywewjx1E0J32wRD+PcoefSRsMlfC7GUOqQjHLhggTN1drTCwqoFK4aTQo0FN3jC3
X5wrbhH78zvYbYfK659t5qAJQNMWfsxrsxDboR2F0d2jx8Hic5wGFQ0NQjWqwBzf
Ls/SLn/SogT9aPwDtoYHCZ8+FrsmrsXUC+1X4bmDbYmAhqOYJbmdBmoMLuUzFRPJ
ltQOtlW4Un4BbDt1Qokb44wRSRCJylgNB3ySSsMpox8jhpcLN+Ul5mIOCKaem1xV
b4NfD4NGIiJ3p/vLEZiqDqgxQXLQSVlmsDUeBZbm5gXi7NSrkmQUXsHqooPFqI8N
GAhfliHTFM5u04YfqNYm3EXKzfH1AM1xL6YXCt8MvqCYuBA8Z1FQd0UrwkSfso6n
McgOFjIgp0rrWKPTD7G62p5q7rV6bh7+/DkSbnFWCRDG8W8fSZGEwNnzfCIbqY9U
eAHMF3YJqSWCuIN16IZ11Hnh9H+1UArJIhepvGcJSB42hEk6HtdY/O9ZhklJMarI
YwIkhC2MXmyFl4u1yN+V8Lzqa8nU+ln0/LCWHOyl5rSI/sDVLKdHsvBIkgBCdrs7
vy1DxUINgyiSM/ADrvAAafeEjNPILAsfL6laKK5sYQTBRo3YSPYlRHXPZRnZznC/
eUzhoP/AXOYPkO7pTPcv3bsjsu6qqGOHsuU7FxGvIK1ICBGUn54OieeTliMEcwvQ
HCqEQ6Q2ftkfAULt8LQjlC9GFSBpH5IqQs7ZNYi/lO3ta1JRi5kyjKV2ZTU1+9M8
aOSIXkAiGusa7ywJqjwVfA+TiedpSpWK7kYpuu3H6FX77Yq3V1QrzfUKzJDzkb4k
SPNbjhKL3zto/uQETNQvlyl+0NJ6voFwW2fOPhuPkATNhMW/thEjTyMh/YN56fDi
kv9b4COnGcw/IqtVd4t8bQyfwZNYYGywpMDENWP8LqmH2XqFlXknJsic33yaSdty
a0nUzXADAwS+VjbMdSkGpq8Jp1Pt3HO/m9LWAF9FF1JcxbsNKx26Yq8zyqGUlHeO
fCPJjX9dM+dFjnnF7NEXzPGGRRw2xlCcuKGrZi2OW91BqtVdpQoIAOnEjZux6w9c
sCqpftDfcQkLOpbTP7O3ahpyLEGWtwlE8xzMAbFLUaxxAQtg2zJx3ZWiTWmDbBtC
wCMET4mEz2xg+7kcgEEhaJDq6e/ZhuiJ9HZ3aDxNfiy9opZhb648LYHX3aWB0mPp
duq8Jzn65IPFxHHOqKkLP8QG+39fA+XYQBef9O21XgEC5gujcIObQtJ4FeSAwq8p
1RfmzwnZYoOcY5iew8uBx6iQilvYRqrB5s/KwJNkpeY6oiSJ6H4tXVAQjQbKd/n1
ToXSxW2KoOKr8ygRj6/kAsOVVI1l3hzu0P+3XlQeIdMNInvf2COZg7IprIsjk85W
9OZmPPanWLlWbZ8GvWav8nqqPfYL+3ylFWFNat8hxUE/+dYuJGYaG5EjRzdt2uk7
ImdtFxpithqYsozi2D/0os8g3qgsXbFHhY2p1j5KbIq6qRXZu8ArU35ENOhJjuY8
jLpgh46niWZnjZeQnezPQM2CLlFHn41FYxzLJL80GFt/cWVqU8NovoqgwfKujbMh
kUBaLO+3jhnlVHSQe18DHcfaRac1ZKl736vucBuJfb5i0jmxWpPWKuthlJf30WQ5
a0kr28RCx+9lS8c2Wlt5ycHSyjJIHMB//+KwmDbVcFuvNuLFytViaQUKlRhIGTTq
WQPTroMhkSHmCltv6kBbZjetWR0CdzWEq6eLY5cuo1rgCP7bp/3DdfMmOUq3YyIx
cuAPt+/Zyx2aSo3zPx5AwBYsU7mTat2VQ7QIxrOH1qPfZJdnhmrf2mhoiUr6yYwI
3a6y5O5xoiE6Dg3wDlgpb9EqP0tYKU0Qk+KnESAcWVrZN8XYb8FXIeNPwbstkfqL
`protect END_PROTECTED
