`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/8dW2PYUckJvIGdbXV1F5woA2Ait2dBDZRLPhyGd6HoBE6J9bz9pSsfNiZohbsEr
XFRk/A5gYcKSDJwQy3HkcOwDL++wPsvYZM+KSaPpwtBcuZBV3kqmaEpxldS02p0q
TfUcDP0bPe1Dwx6RSkWBVc+qITfh7VdAL/zXe4niJT6TbS2+3xWQWACnY9vFkVsH
fCSKqzoB3g1h0AncBIcRus6PHxu4TAcQFvDiFdTCN48crHhYLafpt5E/iZx9Mz5/
S+fu0Jyp8XC3EyiLS8QrHfkF0viqU4OP8pWUhFdmW/0sMm3lKbbU+NTGn769iDCa
fvVbN2xKLPlP5MCbAnYrmoPULMSXDTdw3XtPXoM0i+yY7c0kjMT89jUmkDI7c4o7
Tp6i1/rQfbJQXenbdwdisV/nKK9zQWxPYBp9+fAS3xuwTdwMGWRcINb4/hR0wPEH
s921V2pWN8+DYnuJpfvndoo7ikGocPFQp+ot8wMh/yFFLDrM6TSaCXDJvOLzevAQ
sZ5ZNXoUMd5J1d/H1e+JSY+zjOntAwpzMrUSn5LFxaoIwx0xuEZJv3IZu25Wlsqb
h+hPwd1pR3xqBBG0dRu+8BqVXi9NLK/QrCNFUAtr/0Lvv/Uz75Z3jzNs7G9N6N9d
E9bQyWQVfPbWQa6Q9ctWInlaFFnfBf1Fkv7i7qVeSGZiacoZ/ExcBzk/fsDbZ89O
VI4Qf56bDWyUvKkF2515AyysC72o4lwv7SqW38l/PeM/KqDZ1o2UOm98ujrlR9Sf
S4VgSSc1aNB7qndkoznM0MOusBIkU0N6R+lUxco08WVQISCUMYrUNTYPzn5xf8Wa
IVIyr4iGO30uYfjYedtXdoMCHVzghIyIyHzFKCzfLb7kWNx3Y2pmEqHPzcAFXFd/
aSgzlTk+7P+P8grdRiuFSq9CUWv7C5gNeaiOY+jom1JgscFRfzekQaGopHaUOUz8
XB/wJBuRPrcvBTpTiV4RMzw2FQnqYskfJ4LZo/WYbwnYlWnSemHbupjuYkADZFXK
rLjkH9vY4bp+CbBy/qaIvqx07G0JVcR9RGNXDmSKrbfsztalMFLdrPKSEmJDsf0M
hJdHv7B9CFw31F5tp1CfGhLGV6OOEmqzZZz5pHZzNmNVU73EXNnP1BOjZuvPYqs4
vIS9GlEz2JtmsY+rE/3LyxlCPmhiBMtydiN6z9Jts5oXwBTlQ5DI4/MrDngsyc7t
sz4j4DSBu3NRafF04636O+54Exg/dVN77dQiNCBODbIFbO/ZVUiLCYIYhaHASBK7
+L8ZQMPBnlSPNZKtyWiYNLy7BUuZp3lFofWC1fr9JrrkUvnHuTx48wokS9RwMyvE
hOlUEYgpQ1Mp/fRVxy93VJazJcMT/5qEG9Kyo/cMPHeQsSk3jHNUUr+pK360tuZE
CS5kfXQf6j8ikYQ5AYPE5A+6QKEfVmv2M/1LWBJWUB781b9+ilCgfKB2yDrOR+6F
0wPOxdWPrgtpKR33OIzM9NfHFu/ZJi4EvD6LpPJR/3i+1dBl08TO+354fQzOqJxR
cEvzjx0m2on/q3NR0rCkoyztBJ2BNb61HL+3Da+rf+wyGYCSl1d5ODhT1/NxqXk4
iqDVO7ol7swW2m2CyFJhNATIqd/09xkII3DFZVx0TEpSz4nvP4LlsEwa6HiTUGMw
WtNrfiS6+akEMRHr/vCK9/lZumpRcfplwbN+I0n8Mf9Al4HuBujOG3BdomoeJMPU
EIY+b/hoLpgGtz3Zkb16q8cVIARABnhpS3+q9A9wwWvlUhGrYKRmFHFHDsrf46Ht
5WmV4sqDvmJNSy6hDoYFhxSt0VPCCrK+SkqZhAUqrkJ+Q/k7wApQhTHjFhKUAvTD
Lt6bTqxmUPNBEikLQZBswXhxWxAofGsb2D+yw2UWrrWYPX41BR8waU2zhGUnyV27
OKWNgjLwMAevj1WgGB+xlWhoC3foHtR5oPSRvHM+Rdj0UmBY57dKoMFvwCrtXWXO
6nlmoblsJ4w+cA4e+jR3wsCqI1zZB4qfxxQEFTEEEOMuWXcworutc/AHqTmWbr6f
d15pOp8ik3YErXUA2uEve75btAKRgt2juwhKeA9pldbmx0sinMTiAm1vRpkMleS+
AqlDeiDoysc1X4QpHXYKLslXxQ77OOQEImpRy+tOpgBlBB66OW0+wHpU9FgHpvMW
BD+K2nEHNPUfI30ql86W+NcO8gDuRKlH1eZoxMnAb8zmkupGIsDNWYxWBKva861w
lgljPlXGX2rfro+DDlFlm93aBZrIdYUJNsCsIYKwwOhgka3AZh83HnNPYr0//CSC
aJw/sOBLtDVdP34WM/+/t24zQOJuWDAQfK9OKc3S/fkM3I+dJNUwdS+J5xndvOMv
P0jU7GmsUT1njN6i3b+JuUDhBa3jTZQoBvkg3DbW2wSZwokPwe1MZ5kZtPB2+sn5
x/0WQzHQqG/wk5sljWRXTsqzO+dlcNet6JPhC+vNI5UlIA+t0VJuCF2M2rz7B6Zr
OaN4u49uk13tly0ZoEQ79nQbGTQxRAc1hLWDOHggqfnXk9hQBPJpHkE7oDQbZopa
PCWmbodzphye8AA47DYB3xyzf9/WdTdaAllUUPRI3sq5Gb2WaTNf3Laen5gOmxj1
jxK8WTfGZpHqVrg3c4ZxDxT6YzLKZfFTClu4rZDWiCRlW6wAwT5AbbUK7JiUJHi+
9sUhmmOxYHGbYggJE2iPPdnJDGlt88+KtnZzEi6DzCLhZL57WC1HNBkxYJgkahlD
my5leClIycIvGeimuAx34hiznJ9vndNpNtJ+z/OFXIXph1DVxvkdjmZL5/P1mbTf
h9FnLdCpeWPw+LtXxksKmJqqJywRisSEtDGZ43FUEAAmEOcVN+d03t5n+gVCY3I+
s2+nAq7WuYKDgSMM2qiL7xP5SinlnIPjhfI3dFWA9PdATTZCjGD0GzJanMDyzx7/
vBS16pHmfyerWyIckjM+rlucOFh/WnOyh8VSnQfpxqr3kJwhiP2DZcOasw77aM7e
mi6ZtjTLBFPCDl5cpE+5QHTaIag0O71UTIiamodzA0cTBlcE/WSS7GPtWrAR2hKI
oVdIHlm72O0qwcJJN8QOVHCrqLHPNnpVcnn4S/qxhPLzCPZQEpMPKBlgiAbEW+BL
Lf4ocM6yXSA2Zjm7aoCOo+n7iONVLiAktZDwHlqo5l/4AswdgmY7QJs2N7d2OIPy
ohNB+sS5CFAg+mad1/ncOYxfzePC03dgQTatoR7tvpURk7uCnS7ZjzpiSdE+eBMd
6aR/MANIb6ptVdxX+nbjoDni0h6F9xeapLQ1F4Gomw7LvI/8/1V6QWnUF0FtKWK6
lDLmblDhEw4m/uIC7xH7e9Uq1Mooh70RQoNX/6VsSOXB9pFdaa0s5B4+2+J+R7sY
F1fyu22b90FftjESpv6IY+qXbP1CvAlxaXLMmhiaOM7dXxp5nIErN1zhM3Sx+brE
XCjZotJPNUxcwSH+BSvAg/MJytXVNTPWEeBG9gYCAT5pT1RkBHFcJ5k1gEdHI9/A
f8+15ZT82vsLjnq+1UBgH3+TgcMfgvpglX3f6LaRVerfitrNiFBd6raIyQ+7pyTG
fhGwT7LyH3PziPTmI8XMAJhXAUAEXS1Xvw5t4ZhOn6/ePgtFHRDDMrBLzj+HizNc
GcoUv0O1R+jg0Q79o5oSMJZXFzW7xv0vy9eYQueS+GEtWln4ZqpCQnNbq3FiWunb
ACsS2gozbFgHvAvN9ydMxACr5S+nSodrwNcRjnuoqsr+nhOYZe5ZcSk8XuGdXmMO
3NkYx7n2kRC6DLrrkQDCl4rnDfw1IyLZec67ZfTCoXWzg6oGASpApQnVaijeC1dN
J+MmAhcfk2brlIs4UrEOkvdMpi1Uq0rFoq2vgizBPa6jIZ8ZrRuSjk2Sdz4e1loM
tPBGVdIKbyzsBxShS1sHkKSX5j/kD+x4MdgZq+lKsc2np5y9WsuAwZaw9bM1PrX6
TdF641WIUCp2u2d7TNk+qJwTWENzwGGUX+UXoM7n5IPnbpdBzEe/0em3CHPr833E
vH3a/Fd72EFWr/J7XqDlTd5oBC7EXBJrE30KlSqEbHHNl3VTajUVstJN7SOEk6gp
xyF+dVP9lHvakVCPekWG08Uzc3HQIAVaLGwYqlnmuHKaRXjapmnnNVXp5dIvIe1t
GeJpcdtVPZ9Rn/aSZu0jIJM4GWtkewrBHepCKBj5uYxf9N2brk9vmRVSeGh+br1+
/34Xig6B93uZ0s31b0/ymbgQhDKSGGv7pOevRIQ+p92t/tRtiQDezOjisqBu2Mg6
jd8YEgF0zdhKjiEvyOWRPopxgWczg8uVYxgoYOSmoUDLjHno5Mag6fKjMh8Tt8JT
yj5UKurw01QrJATYTK+UPz253LV4Ub51FaHjTPrh9l6D2/+3q1/OnCnVVUUIE2AE
9rAJY6JyfPhih8cwUfM3Daz10Ba1mCNgGu7U88FYvKrc28P+7tt0JUcMD9MJew4d
`protect END_PROTECTED
