`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CSH7ya7Pl6xdUtMgFsmtadiIKGPAXBbaAxJyHqozzubY1I2nQ32+Af/XN/LJ5Ole
/uCTiP+PLSYwFpzU3f+fDqdg8RzZo+uB9WaHarr8mvPEJJpb2Hw2XPPAVyL8PgNU
7uMw00+XzmrLz7yKV+th/Wd5h008XlDc/+I2lA8DIdzc+9GqS9L5AtNwvegkrKrq
4AqmTMTo7nkWJhHQe7KMFCKCNwRy+9K5nDPkPV1PHrsSi6KFZ2z6OuwqWQaa2jTJ
ZQFYCmNLJeytWJyz0ntUQG6Ku/C1nrAFCibK52ib0uEO90FlGoAe6bPEMcDGPoaf
cbugmJJN21uLo7RSIpkPRTpAx1S0wZ+jzWD4K8Iuo8n5SIqg46+g18v9VHwRMQt+
2bBziP414m4o9uo/c2JqYrG9BXM7irWsMqRWFyb/U0B3uG+bdwSzamGSiuL4ywXH
GH3bbOXCGmifQWC4k68HlULDdBShMOZLYJ6Ehg+6XooNQUagB85zvFcVNCZ7VEO+
sAhe7/XowkC0PWILibXApaExOgiv0BqiHxBb1i/pSmb5WlSfmvrj1h1GfKXYnf3z
zku5/QwrCr3L+r1sAGAlFhTI8sIorofS93V9stAxbnF+CDox1yiH9hILbeTicr1a
TRy/HLN2qJsyf+VVdQmriTrp5SPGk2sJG9mol39T0C5PmBKrl9Kbokfx4l9ymYID
77gnHibZsLbs78I0L4Rz9kfOaDzgzxrwW9BLgkUfJhmENQOisHIB1ks6kiTCQE08
xHIE18GUr+l5cwqm8GGuxb5WADQ1tUTNJ3IB8pRjj8l+vzf/hwSS+a7NnzZxhE1s
LeN/bnMV+t9pAz0Kt+zN0XpP3luYEKh9drNzQ/QYHpw9iCgmVCn7iSj+WhzfcTwl
HeL5iai/wE84vuZHOXxo0y0amsCCJh+RHCeqEHaW2ZcFVjWuqHSUjIiNt2wTQm0w
`protect END_PROTECTED
