`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fIDgg1o5OKiUzvVgeRnKHDOysVGPhPr6fMG1j2UMKu2X0wUhJSRJL3ZQUzVWkYxn
ABERlm3npfQiXhevhfyaYegmyAJah7jz0VA0kub2P1FMLg/n+QhfqSZj6+1WuLTv
IcGNFuQanZ11r90vZ42PRdkbWaTYC3JS85C9RFBpCY3eU3wtEvTM7k09kX9dN1e5
OgkufinwFbRMCyoUTOVQ52k+z1mzPKyQL9T8EQif5O0QzIHaTOFrt4Ix6HUs3WeZ
4BNECEjdKBI/8hybA2dEipD5nISF8TChtEkKhcneNMEkAbQ9krwzL1Kdr97ceosd
Upv1aEh1Xsh52aStyFowVT+P6RwLZ3QvFNCGX8VEH7NopR8OXSmRkAvLIemM9nyE
PuYOyEoE8914aQyvqqcNxpBDK55RcW4t5fL6gAl6VkL4GS7nhd3PPBQxdnAMFh0I
kIQwNmwNU3LMY1khDm7/9crO1UowHs65PcRjCeGX6KLDhktHrT4nIZLxHplThFKd
XcQm9purUE6ooY2OAbUSL2skLYK4ZN0K2W80GvVdeUSQh9bRD9P26XYBB+Y1xupu
LIZkxVLHDWT0cWfZuyQ2PcxJ6LNe3R2WPNS/BsAvl9FJ/oVc3dzAq1tpZX0f9mDi
BSc0Lj6zK3Ywcz/hC3ZExOm+y4QjW72TRDCdU9yJ0ZkPO95mUq5GVeTgA5EFUMeS
9F56UXjBtOJDafPTchy+wc7If+5uwMP9HcqFwA2nt7JcJyEr67ydwy8JEKgihzU1
haE5i4C3nIAJan+MjBJ4TaJwvxOe0QaYXStrKInAtgZMfEqQp99lDsrRxIIFk+zz
jr+hG8ywADRQlOAGbeDK0+vqBNBKxtOhHyjtwPy3zYG1rgKOCb4ATG2yQn33wCpG
Adf9K0yUlALf3xVQtIsnwnR3qzlLOCR7X/eOkY80j0ouE56XizL8eT8ZYswW9J2h
Wt3p70xH2AfJympa4ZK1i25DbrY3Z7ezHYFmZYiivz6r+SUYO8ZyQA7mzCrbP/7s
HyFzOAOi52JaaPesctsZLigAyJ1aSenSl6KRA0duIYrXUAHat2Hz+WMmHiVgFESk
Ql08Rzb0tsq6USn+LmACNdjlZ/vzZXQdypWRUTUj8LUsc6PtFV0IvXc5yjG91GT6
CzjtuQRBUecPmbOUtZ0eHmiUXUK6lYa/gm/rOMOMQRRHorDnQqeAqPIYmxG5B16G
nbLt4RK0AN63ZCt16hrfAkEw4KAt+f1GuDEGyS4nZbKSYWj4/sZOopAXy+Z8pqTS
eqcQh5gyKWGTYp3F3znh0V0vjHiGDcz6S7fwQy1x7LT/qDLPKip6HjryEOXXW/9K
8GZZbScHaD8TziV1O3VwXcHaqK1WnvMXoUHMW/OvzaiIbIvetGKNo/Ie0+p1IluA
JOH4K0HebEiHqXVieRIGYTnP2kZQ1zhCnW9ughRg7TOAAHszRO4uet80UzJ136XB
EiXSSEK73YfJqa3Y7Oq/oRwKwCqgqYLYjyF/poCx7qf+vPxX6QGVL5dmQVSHvhpN
stIFI846UlJhQo/XjnPUHd6+GBFSJJB4F1TwEQ6Topdc4Eck29mMuTb0sihgjkLv
BJ50FuaxEmiUIKwBiTDdLdYJQevtaoGmE53Q0xQ5VR46LT+4v/Hi19BOZRe4/hyZ
LWfc4TbwxXM1qarp6cH5D+fM0WX1T2mJyaubfSBWbdO+ylEu2q4tXtwBJXQmML7z
cFHb70rdJ8cLcyFA+H/xEdMMmsZru/dk0BA41uN2iDIrIxnMryTjlF9+43aOrF6R
iXZ6bbp4+8Y7tl6ET54o6Mu/l1nZYUYaar05TOe+xPEGTtu7160VJntYcaiKGOHK
tKZTNWabCRB2KPhi5cASbAgjtzXqvFrmkcWRIGMedJ8hVt0SoOGKLTq5QidNSdL/
v+u+QM4c7CXiJeuKgl6Ls/KVrcd0mNGerXk3wYS4IM/VVSS/ANpaTlg0aDjrH1Jv
HdNnkJkp1+WL7OwToe3iN9rB3jpQ2gqARI+bQIb2HwGqqNcU7QdySU1mj2pE6wn2
K9C5TocN/or9Pw6JllNoO5qDtpNfLdk++th0GNIjaD0AbXa7eIkopjLmdWF3/jfO
9CPuCvMdidby+NsA9KO9ZvXTs6+qpsPa+n5Hw34QVFWFRfWsh9lr5b0nlxEt9BsJ
pJm6HAiWDAWzkDVbNl571kh/iaOz+LsdTSR2+ZYWV0ijWBYGtia1FZBV3u+eTuKy
jEWbm2JCrWBvRSoiAxEl7eGpBwc1bb31eCZng4IZWK+WEW/P0L8khJ0YPFcWPHLr
2pEsdIEM72EMzYxOo/zNUwuqxQE0+dzGQ2+dO16GZCrO4VbbZYDStbB6zvutuF1T
SuY6EZkw66TvtEnaXQIKK+CnmUQYALf2X4XlF92RO+mY89skKkHvw295W40a9Hkk
w5Xd/KQDimHfZM/aWUXwMwYHk7ZdoARM1DSVukCa18c9ZlhPuGk5a0BmwljKVD8x
SAuMKqgmH+erLici8SLHj6vGbS77x/vxU6Yra5xUND1p88AuR8Bu0YMDR1y3jZkG
BGPKG5vv1PmygSQol05S4eXP7OTs5GbNxVYyM9cjWcFQ/rD9zRH3NdDw7a1CarZ+
LwQRK1v9QvUDbg5necX0/23xj1J86uZaq22xK4nd4Du6KCgE6l/WWjNtx0CliOiF
l1jn0Efe2cHjw+h+otz78vIPWXc0Kk8bid9IUr9le69ougz77G75FwiwgDfGLaxX
dyJYHAwZLCKHW/A4wjoqBpRbo8GPtx/5WGlC4oI3Ro0u7a75rOfaSZcGK/YuvACp
KzqNyajkMAntRqXQc5DgfRy33nLNzFtMFI+08KZmcuH+wib7sGb9aqZnhh0+Wzac
1W+6AtGi6vWZQLrj6HXGzsINZ1ZIbXmN9a1KlIcpNcyhBqAP3D0DZhL0DCq5HP9R
Q3eD1/1sJGH7jktLVpF41M3MVItQJnHaRmNldukqT5+ucbaRsCF0a0oVdGLIyTFR
K6RNpmNxjlVAghEdzRpocwHJ3xXDPDyGHoQbw43okgPFWD9HP6t8TZBDuCM2q0oM
j9y5Bar8rNdmLPEdD8CVuY6Jwr+lDKBvfjIS+V3MAWIDg4M1ieXVXwX3Ux/xw9MM
DMhnHg9myfBwKG9BiG9f1jpWSjanG1DSkpACdP9kLaRm/V1fED/69qGMfnVpG9Rw
QoTB+qZ6Elk2EIG69TyfQTk56I61Y+sOlx7yUnXVr/5CVEaC5UfPkPsH8sgP4EgM
eZmjnskZ0JQwLs11Zo9lxwe6jONBugCE0gBIdiul/cHkDfmt4eu+yXSD6KeJ+vxK
Y126jWT+DjfKehVN4CiTia8XXyumRsPP3rUGCbK3C4O3ZytLr3mRZjiXueEavupK
8/bgSeLnJcUYgmLwft/86281YmI+NtvuBbwI1HP/oelGxg4Jd+RFqyBLSGPhPXJY
bQw6x19wI4l6t9iub3eDx3uZtttn61K1Lk5stVo5GPAexbIjy80D3kGBvmlARhRq
S1IU71A/UYDZ6ncCvCcLfm6t1l5RolvndQ5Zq5g0n0enkIWZ2BtB2pxbTDzLy4B0
1NaMSUU3oiMHtMz2IYdmIaeEb0AuC5vfr6saNwTOKfCkLWfgYokQMMtOYpRNiPh6
DdImIPYg4PXwX1waaLqxZ1XgnB14rXVoeJpAt1Si2TROC6QzKByybpaVSBfekMjR
zn3Xr6Eqtv1cRcty/4WI8apGNaJ5NIKpwyqLthuwm4iyFyazDJ3k40JAxdbhXFcT
MLs2FWBB+4U+u2NIhBCkQmMMGfGt6bDLgForeeRPrhCGi63aWyUsw8iJFOSwy4e1
VQkpmf+HakcHQ3pElMefWxSUI0x3muyNBIstza5SjojoKGF0An2ArP5RT1zy2B7n
lj0sgzxtK4vB757H3B1BABstLvdvwDmo2JgsqvxZJQeGdaPbUmN/5cS0zJgjWhI4
9yRefycM4NgQ+uOADyUL1f82sXP8x6upxPh4s5NxnQ7uk2n36Lh2XavYfgfPShPd
Fyx7OV69ruaCLUK6DmV7+4JRlHyc/fa244bGu3pXMcKkOe1BVOj9fjGzGqQ8nhGr
M/SGRzZerNmQFCK7gaxvOPij3T0veAsIyyY5aig8MkbVBaiMpcawJRUXRmWmg2Ow
SaMYS/ldwbO+IZPZqXBMMQM6G8gCBCycUCgBnsfpikIhZEOoSXout3N8rrgXhRTd
G71Q+ziiGbpVuGWEdcmafIxRXL+geg9DEaHhtU3Mp2MyjC4VVgzn4WDhc5Sj6QGB
u8Ra/u6T/n0h7jCyh/yYFo0L1oUgzgnasbKfPRb+pJZQGeCNvmvJ2mHfhdAo1bKO
qvwb5k3wxJCtR7wR4uPH1Se/gE4kTAuEF29uac8KBYTZPukFcp9wGoK6x+F/RQhr
cOAu7Edn9TUTK/Zv/OrHb3vGFg5tAaHqWT4ZQkDHAq0iRkp6Cq4pPB0SRbtQWHG9
RT6LIBujDa+tx7eqQpxOhf7iuDBRPn3Rt0g36RkMvVOxup1HJStvYsgXPGS7lt8F
BMsfVbmdx2UaL+HcuUbDBJfmtIkTmGVQYPkjvjq/o8ZdKDmjMDwimsF7CWBzQjB8
9i2aB7vZySANL2AepPRSEqx5OMsA3V87qeBhSBhYO7jxFwvd2gTUk8CZlr2RXrgO
TM3CFtBtjE/qc1aRzm+CqkrRFJdQrGNEEKTAbxAfdFDCbc2hVbA/ZNPveYp8MJCf
lWKqIBe6LfadJOR9HvHmxL3pb1py12TkDAeHSUpT9uw0tMUhd3gbSq0uPnFYfv6U
4BEiETP2/v1OkWrvIS7HopSg9t+mL8vamGoQlis7w3L+MGWCgeCxFjBtPULB6iFS
dN8Tya+NGe/7mus97wGZYfLvceL0+m+1YcS9pHS/jSa/5xQBxwJ5anPHDtbMGOqW
Dhax6vBPmFpKYi/DyfoTKlzZvxgTlYbZJkFDi3VFffJAop6pV25n9ReXaaZ76btU
bfIWLwlyshr3dUEZ+HSadWzDRUHrBqWvzkOwu+R5z5qaKhf0YuYTRXZFl3uhkxwA
6m6bgqS2j13pLDzDqaUp4a4q+zSpEAy69SyGl3XwKwZMk1ZSGzN3f+spvXlcOHox
dwgQXYHs+nNNDeo1QqABPCQgs61pTUZZ1TU0w+XsZSBew5jGT3HvkQXgyuo1X/0E
o97nSiqSm5bUITv/QEyphhw5gkkRdDsOGF9Cv9Mizp9jy9vpiN3UXIWFDn8SucL4
CRuHjLXY5Ex+ahgWj+64OmhKuBeMT3wqgR57m6Jk0ctAjVg8A+abC2Pq2Vnr3lLE
b7eGkc1APQojSsU3oIuatT/3u6QpHccoeJRGdgyu7gP2/YCLHujorvB1L9Swlpbp
4pWL4olQBj1VPVg2yPqdANYl7q5YMl4ZMHvoqBTDymk6R1hWfkzplCWG52n/ZQNp
FEh0l8F9LCu+4/OmnR5rOVBZdz+Ecuf1t34jyAqZ0eMbUi1JpdN0Yx+QNG5MG389
upWoRRuTTbHGRp6cCM/m7LLiRkRo4nSKNiYHJudt0Mi8nuw6glgMi/SErkRjjHvp
XdmW96+XnnOQppK6TA1Mu41asEvr+BDNXRYiFku+OLMG3ZZJuBT4kZM4M5kQrUpD
HZayYrFMeFRclpRn1yaR0hmd9/zO1xTc9QfBcbpHyETFZyPnOOh6TAodJXJWdWDy
uFjt1edCeCLs5MIfb2o7x06y/NOkiO/JlkpNZfmEqqhbqzBMUYfYWoERUH07nfT1
fcojNwUrd+FGEyvk7PUjO3Oeos2vkNSQTsK+1y72jJ8LeyjaP03Fz/ZouPPx6jov
imLuA01hUxEcl89p7F+eXYMiBtSuPn6RPbdmypH70Gu1a2mswHpS+qsWSR5JMlG3
6qa6ht4VCt00urO6fnxHcD20lLpZrKPgX0UioeD7yDQuVj8pvFEp1le51Yfn2w7B
G7XZcuSWrKZKJfmukh+W3qbnRnGumhd/qx9pZD30leKCkheoPdjQynaTNFGLrh5y
fYagM2zRxOZWAFPQfdIbT++xsAfGr+VuzhLiry/Oc5HJRzUzBzKcnUqmAqWXbMzy
ddapcuO7E+CF30Ub7nbIuCg/rzza4JmsbM61MTkvW65bpktpRENz0ay9zeZNs9lc
QagEOWEKHVJH0dhaoFOsdDT53bxLhUyzhSzewzc1a2ELUjVJ1FFjFJyfBGNAIPoC
mD2rtyEbQ7iiok++h69m9j6iHuqDYuULpttuU6ZDn6dYPBJDTXpNH6Rwg33baTZc
mx1Wp7vpMU45dLRVmw7mC6payMCjhnEucJ2yeO6yvDC0PodVWWL/vVXb2GXNdiOg
nX+ckXp9iTRW1/h7qnKPp/AYgbSJck3s12Uyq8dadMJO8UAzauW1E3mg1GJva18E
LXmLsbfKyHgiggPhpWmMg98BskJWq30ZdcUh/qO0Fh86o+hr6WIXsPVs4guxIt9I
C616pPupIL6P4PoonKxSXR5C8cRZgwwFhy+P2iC9hYt2ay81VJV/3BY1nAdHyOGu
rVR6IWLhYbm46qIufeDN30lXo2Aqe6QYPPLRO0uty3K8GyqU3MYuzbp3fsTe1AT/
76qctXOokB36/mJ85SQ+Ka2JAZuImKqS2+zRdzyxD3wvqgv3JJOQDw3/zQgXYRI5
roZ1sYed9lCEdj0V5FumyoVnIHLs4HUzBg4dkgdDTw3bxQFMbx8RPkk1F7WIFBAB
ax2lvW8vZ+MZMx912e+Kd+3opYXKk+Uk9TaWrDZtzN0oYvu2fYhfTejfaMr/eOqj
Razp10EZLuQnEyGshOY/YeRzVnsOrrMJCSXMJJ4U1Dd8IB1nF755ceab1uMvB21f
16vzul2Zi5iizEvElvQBr1XAuUhxVr9toIwtZwSn/zaAyE4UliU9AryQVShEQX23
4pqCwT/OM1r+cR1nJNObOYVTz15cp0H40rBMhEw94zKPUnu0OdE8A6wnrMbpqZWt
H31ra+PrGLetG5C1zPrsBrsfa1OTs2KQHYx+IujREBUQRl5GzpOT/cginxVfibNR
Lo5GLJzlNtrjYV4RgbxHQLak7C3hXwyaMzbmyBlFQcb7Wkvvq38HXctYpepVLM6+
EHEApzIClC38mWmu9XwufqgtH3qJ/P2XuMmCzO4CIyzamXNpqbM9Ar22CgOdrEMB
4nRoDRd6tXX2KA8wdGpNWRnGqVlJHnuHDwXTFPhuXQI8/POMrSCZxfcoYvIO7RxR
KpNXV/bniBBlYSwNeDhwXES0y6qSTScRWIlAmRu1cG1qWuM23LFV8+cnNwmvfDNF
j9BcjPzKECkJZ7YkOzDJinAnczE/oQJ1j+JEfaGEGSkoCRGk/Z0r1S889V7shWZl
ZBjXKEf9AEoqG8YGseYaCYt24Y568nRbJ8XV8kU6+bHCemqAZuA3ELb+TDuLxoin
C4062bIRmqujyvi4qgrYzDx47x6ahN9XRPEg9IkinYFcqWFyOGH6/+M/WXd5yAwg
WS9x2U8g10sNkUFhIeVa6fLySTHnIcUqpsgM+ruIpkRq4C8LilfgURQrcUUSRUCo
Ro7eY1tp6YtYrpgtesgOU80PSv2dYLfEOsFzqtBSIqYsBiiFZGyITe41/DKFDniU
x0sYW6ZRsm79fCjkYj/w0bkp7hZrhCBAYogiicEkfJgLj2fzaoPLo1C8trhaQbPx
AoHGJCuvlxcBdsFfuZohfuRJyjmly6i86r/aV8LISBQTSeB6QjJTwYKU42iXQbS6
O2bqdn+AId5566kGplsFHo3PI8EuEm95uO5bjZp2PiUaAUd3jDE0zcMrsfhOk5mu
HLrQIoIEUHgRcoJ347ySKAoy6/oWAaY03Nr9RRG9U1PeI69e/gSaSGaoG4xVOi5w
yphf+AGY1JhEYS/Aqz+75z032IZuvZLFRbtdVKEiKJqAi8Qnt04LDQs+8/E8oFT1
WMLznDVqETT9YIvihg7+dxA1Z83cV8Hh510Y7YvIhn8DGuEClSHucQU3YRYzU9qg
yzv8oSj6sVM1KmVjm0GkC3xy+xuIgsPfpugSKF/rltTGNJH1eujejjAvj0Uvx0Wk
OqNy8HAIqI2xCMMjY7QUY4OSMfiX+GlyzWsY3WjM17uPlMUaSTh19sczjcfeuIgt
McLKS8AwRq9wYLr2wnHd+CrR8w8Vx24VsCaynBhGzhZGInMoIInyfOm3tTXfo+IR
/Ze2HZbuffOAieGjcafiSx0hIkzPonVXXMOyPm0/w7lziy7V2PpRhg361cpjxnmj
iwc/GnUB3il5XFE+0Z5GnNuNGOj7o8xzhkJuC0DFOGqet3LAFu9tSdKdVLE6yQQc
oghUdnfwBIatHLqg7Q62xML/daxU9NWkek3w2Irrh4qIJDSItYm3WHkjAPxq6WJ2
FHFlfPnppa6elkmBIC/FxuH71kXZEHH9mp+znBvqglociUft9bo6/fjulee93Tj+
u5tGdDCTikNyziGHSeuHRw2RsZq0mCEJejLvxykZOZkW+i8jFigI5mVXztmVL9Fr
UZ8+yAtQ459gqBX1Y7tXMWgDANMKdTWfHZT87hi7DDWZ4L8QJsOCQb+hv8q5Vwic
xLnd/X5rH7wfGr64x9Qdzo9fCJfV/tDi68CCIpzq+9H1r13j7q2EHWSdTxX2jNWn
WmoolsRYW0Dh+IJd4kzSr14jZ3WhPH4Zbw44vVD1PdFVmmHknKVXLBr3vOXECeCy
23QZ7QopeW90796fnL9eQM5HridqTYWatWDOA1bZkwlovCIKB+Pt/pX6XH4H0XQy
ZOC3ZjaMx8g1pnUPmntKOY2+NWNC0URt6dmCO11CO8uGpnJVTyap8VpFVFKNSPhN
eRGyyczyzjFTqJcEYshRc7aALqB4MhmZXQWMky6MeAPaNR6ol46HneG7TRgaYZkp
UNRpcrdNKyHtgxCe2Y5fdiVgIJn/PH4kH3R5WxWQGfYBJTOrcbMeLLXpcshGydg7
EOxVk80MrmtlrvbL9lVVQet5Qrnb2UYB9Rbwz8f0eiO/CldrpoeD5CnJzoBxYAYz
ckkWjsrcGYGa4hl1VS7aoiSDzbP+WBoPX4PCcj8Wxkbjm5ieSJ7VqRWjz7uniPN/
G1mX3wP9sxxdsSQ4s6jLAjarhjJ4A0zaH6bCLUjWbP9ydmPgzuEv8tB1pgKoPCy1
zL5Bg6gJGK8K3/YKPEJplEX7Y7dX4w4nXAPlEDPrS8jDmwDJAp8NX2hbbOhhyXP0
Y+4AUhRYUOYh64o2un2jHPz34lFmkeEezMdCDp7F+jeOkKRnUejOsA7E8dugFo22
a8opJJfXZ+UM5VK0WtDCuQOANMgWYgIemo1dFXFw76J4BMWq6yKLfKQDUwKxtN8Q
NVFYpeIXSjGMOovV3Iw7IBpR6R85q+QZuGwiqqYYi3qF1Gq9WqvE5LCmW5kUfjIz
EMlwCA6dpa6ML4I4Xg+eT3jyOJkRk0Kwq23tRrxZP9eTe7SpyyWYuUgALkJv/giR
wGu65k3ncS6Q6KLzeL4G/z6esXKjeENGdoiMxW0iRxGHQ0Mkrj2dxobpHmnbQLv3
YK0wyPTWMzlduaR8ESHtyt0Ck+hYyQHtDQ1EpDG9k0srG5szADv1FtzTxaECNGNr
mIFyl4kyXcmxLC0ndXPnUbqnmT0ynE7K6iaFzQ7RWh5S1ogtkjIInekampwZC2bH
HmJ4+ox8xBr1hEnK9+1xw4uA/b9ZMeQ0HFKaSN/Yg5e+as5AmZ3i4Q0YkBfu9Wot
jIHwbMdCDNnUZii9C5/p96SorCQ2JSzMAogvgbDoJI/zkcVUIQky8lP8WrMWutCQ
+V+XWf8cuukVjj3drDn29ti5Ock6GBS0U5BOEA36LZRSXNBLWNn42NPwW1SofS/1
Dj6WnjY1P2F88mui1qX6hcoHenvPNIoSMuMImJzWZq8X/gRMGt5Vb5B81fPTzUcL
S7NBoKSYmOIxKfY5ijyQdzI3CIaecZlrdKNiDl5mrSWgZP07G0xoEROnhAv4HJxI
y1jdMUC8eeWPsyPhnMDZewmljurFGfZu32rq8J9d+CS+EcHU+mPEvxIIXqukEPlw
CQ0ccKpHjq2ZwidBZoYYR8DPjforJOMXKnNkafTz0/aAqczT57FJjE/IFZw7xGtS
AnckyfliU3tZ1u1WG/jD+q7nCO8e06qR/36Ur6/OYs885EMcpbHyFVX+5lrTqeK/
O9JfThQ919vd4l4LuIHOKvx06IF2nTY7Uc27RXd7H6Ir37H4co0ySW6qTGGvXwE3
aZO5X+eKRORH174l9xPf9xIG6FCCK8V73H1QDMGsg/pu4vd9dM8/faUkWuFPIZ0O
V3A7JRkAAjfUiKLUYc3+o03mjJT6mQhN5aZffmwRT2ly9tM9y+PVn4H1M/rClmt5
YeoqFoPF4ZNCeUgtfuRKjNDZQumK/zJVslVzmZt/Uogmv6h6MSknm6SUXM3ZznEH
5seD9plpn1bUuiK6/q32qBPUDRJAXH47ZBH1Rc2fNIfJGZZvvzyj0ILYVVPHXnU+
+u3cFHuLi3TiyqTohIsCSLXv7OunaAxxE4OzgrAFadC8dpRUiMLHWjY9OU8dgJ84
lQWp+mdu/ULQ5mTSxDdXhklO69UdRP5PxdZQkmzujCS73wCzxhsaAVa1kexydavn
BL2o0BRoUMRDan4tYosjgSEzHRa6wB7UTJxSWrGdetwahUJKJ4Mp1sd2VkDvVaFR
4cnWVWtjFHSc0C2OFsv9dqb6CesCYEbmcLejaxjrc0QXxcPmgOq/HdXp7dDM6dco
AjV4UczCq6OVL3ZNuNiAypcL5rAZzAkwsV3yTIZ6rIgKB4DIwua6hGP9dv8WViVD
LXf88pNmtCN78QWl+xgWKKddiA6aXdMcGFPjI/G0nRTc2OLC6WeBWW5+Aw7Ex6dm
Uyh41g5AqPPADe9Vpt/n/xPxZByQFOEPJErkK5ojSh9YreUIQ3suQFhNqlbp2e/1
J8KxeRv+3iNtVIgR4qO4dNKpSbhQHX+TFC8HI74AZFQxMk1ZgLxl4TaqY2hoikn9
hxe/YW/Dp/xJhLUcP6csp18LFL7cFPO1QLPqSzdv/qcYLA4UrPJkzZWClkVNPIcw
OWBjENbGL3JxWiRFrPeXd4n4x4yYVZi1jc1RoQ+2UAZH0IkewwWhzWdup7AoLj47
HGdrsQfNdCWbzc33N5i4vvDfXEjKrFQBx17tXnoLROypwAnKANmBVn/hpOcdWhAI
k3t8sxeaINvhnZlr4y99rEqW5LiuXRkCoBiJnJlvltP4WOTuMLWWoTEyetJ7+C7i
pG52HsvkOhCLaIE48zJ5u0Ympn6A2EnK5VDezlWufG3IwSawC609nmWvgJFgAR1x
N0gNTO2nISwlK7QW1SADAiv5Kovov1BCjjW0uaVMKjFLY2VLIt5Ji6spMi2tz4NX
p47UnJ/9Aa37Dt0Anaz/uRxOTYIt0vdubWRRv/eN+TRmo9Lpa+GfOvYZ8cv6sTJI
l6CdoPGGk+Ks8niU8vHvIhA/yK0dTrSe7F119FpR3AXp7e3x1vj8mlyGCDy7sR4b
0e8zeFRPSgnKY16gnDhTmK+ztgNJN3SxZbQpRtwCo04PE1cvbMhLZHE8pOvgV9Ov
+oFoSOCnJcQAU9tdg3tCN92BbGeUFaeLrmI8IQLfFMYvi3bRXP6iKY4hJGwbjVcI
ZPKAUG685n9iHBcHklf4RCqhkJ9oOMkZsHCpoRhsB47PJsxoxFq2QnQPxn2tWyoj
f83ZPDIrBwamDfHIcV+D53Xn+cySqyprgKp4i/7BCE8JW18Zoo8bKtv4DWhS0owQ
oHeAE2fbapa/nb/PFWKJxiBUWgJZTnj4kxTR2AaGJjteDlCORGdBRTUwVfwe47y4
ZZ+HRvu5NvZu1TI8ELARnIq3bbig+EkMK6KW61mVrCIQIst/dPC6EYPk94OqLtPx
F02aZD2ASqVRJZGIuXaA4S7Em58m8nUwL6XF0YYVz8rJzq2t/CpjKdSIbD+dq+43
urqSgBml+OoTWve3MPrek6Gzv9EYp35efKSq6m/ohxw+xJYxXXrBjTs+5BHfB4iE
0RxZifWhEzJH1nIj19k7tmIeVvYDft6AcyECyq9RIutWs8kvcQJlJZwGkiTjK3zu
EJ8nybf0VJVPa5Zvj5bqjFv7AkGKN6OraLx84VzGsaHYXfnUu89e5DPET9ZkZxSg
tro9zLcItZzKnPAHddocz+wjGLf85vc/VozYTIT9wkwuhL/TQwXWvvPn+N6BM+mk
TlRMhPRQCqRFnaSC1j2osq2pxXBB6gIQ1dprNqDSmZb/y4IaK1VAwRTvJYt8QmqE
41IPXN1GbJxuguHorT8gjWLQza9Lz3zeOc8Vj3guflR5foGFSC9cNEQJjKD0Y4/X
buqXZtGSAeFpw8hoP/EtYisfnTuIXzpXxdnst80DRdTLwhSAxMiDyp9WfmUjhtKC
rs2bpHN1/2tsFIXc8+dDtlf5oTSuYiIXWEW6CUnrs8HRr1xl6WonvSWxlbmeEP1a
rSAXa8tctYYfFDvuS4Sh+A==
`protect END_PROTECTED
