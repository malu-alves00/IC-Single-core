`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qbqjOqeM+f8uOlHLYUpDrRGAq3rvBWkpmfWWVo4jqTE218s6aKyNlcCPpxoZ3H/7
CZD2dNSMeeofdQ5fYEP84ccaZnOj/QNrwHhcl0OfadvXuFnR+urEK+osjBKtY+AL
m8o5+kezSpEfpGl6Fi94bLwjDY/kKP3HIdX4QLCvLlnRzu0OwyUqGy5DL8rYJzRq
qKg0gn8WZGMybEh8uoWvpw==
`protect END_PROTECTED
