`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vE5BRspuJu9gaVZaq8iJAHvH5OvLDTMHyuA9nb5k7oULqGnGkATJWbrcjL9sN4Ei
2KRFWA9cqQcUzEdWH0Wt+A10TRVCyAVuGlk3VwZ+FVE94fmckIFkkc0uCMKNcGc1
pxkpFuGIv5JRAyUUoFWcftCrSxuR81IXYCibpO4KdSqsLm+ykRWieyJMfNWIfxz+
vUuHgDOa7Y1QuTjeG+yf4Q/Y+wfFOeq6225fRf4HvGVtu28x9iMcxi6Gg5ALDlMS
IM/0/fxP7f3mQeuMOK3YLAb02/gvBKONkAUzZR7hAqyaPi6jxmuW5UxxwX71D9iZ
hGUrRHVDDnmy0hOeMfYjllGbYWH2EZoH6iKlSdF3lA32GWhM8B/uX70+MmhvAIJK
RmrXCVbPnK0B7m1WUC5Ty3M2gvxQLjGmUZF+FvF8+5rJDwM2MWgp2cuawwc+HAyK
CwwltIPW5733WP+kUYUsN4E9HbJOh7SSuQQ0slY7JqyeMUclFgRWnuFaXOQI+WzN
l0ZB5Emu5WN4ZrWTHALlCHskvm1zfV90vsJYUjmDf/lZLZuIuw9m5cAzApSZkS9D
c+u232K2sZSN7bTlDhw65VfTMbBkYrCgJrRz49637HyxraIPmqlcYCnTBD1A1BHP
lgUSXJKM6s1choKMgHue2NLEGQtMoFL7esADfCq9DuhIs3OHZYDanZj7gKLfcqjq
binQAD48J/fN7kJQokp6wPRGKzyi3cl5GIu1os58uqmaoI1SbzvmrUGQyrZD7Rzx
/9wDg5nSAmOiMd7xyizwOOllqJvDuIVD06KjOz2821iGjHmfykk/uJ0HQmbjfI+9
sbRXSKvoHXXr5vOWuI19SG6w581o90Tfx5rHrTA+OWm0p3dfEwrUFmpQ2sab+XsU
jBN162+/20I0Ys81ZIZ/UD3FNcufoEdgwCwPmMSV/ydykvHu4SaJMkxRAc3GW0/X
holqdzcTMVpfQnfYBBCUkeRhuCJs8kNZDxZ/ffCsxsN8qjWcPeVM/wI398RssKZ5
JWI1jGoCi7zXyq7764Jg+JLRBy+nVgt1T2XCiDfl855xe5b50AtD2UVRpXsRsT0D
aoahDRQ4+wmnHWSmv8QZ9tPijJ/dgmlg9Jcf8yM97noXxo+93WDcG6gq/Vs8ZlOo
VJbfAqanmCx62XFImVEQm2Wh/gRGZ+XdfU5WT4lc9cIk6Hc8BDNyJbVMQM0EfbZ7
QiV78ac4vNw/T/0a91kUbh6RcVtFCA7Il74mZ2I2GhTr7hoGsMYHtRevh/WTTsln
QDuMBR0qenu2yrMskGV0GGIIbr05sffdjv7YZAjLKInK3hRG2vDANUeK7WVS4OEB
CQxEJuLhLZ/7ATxcUI8+qc441DfskQ1IHxUFq+Aty+EwHSWbV8ZEExRRNbcGuPTf
4kwVjJtmJlzOxhV5fuba7eIs5NThkJyZ1wbyhjLLmwxZVdmOsLMRgxOhbBQ5q0Rr
UnSBqbuHzqBAh32oxtenKmJYvw7T0AQIBlF7LusVrFV261NXO3pqRthSiEiIcw3o
3AsfaREkS6fwAs0YVoIz3sVkAGWe4REV/YvIRQyYEaQctsvGxoUOYeqnQHBKmM4n
ue3Nf3703fOSO3DgVlcZyj4sM90BqwYvZQ5xxgIXr6Q8nRMYyXE1SDc0dbe7PkK8
/gp/LawlXtzqLFvvqA0NTfm1lAR7Z7UC5Xd7lxRSsB1b5D3kDlAAwW+GfcnnPWLI
y8zobwnmaPfUebrUAd/5gkDMjBRbP67CSmiA1nC2TZM2iHXNhEEs8Z6jS/RMbwf/
lbx9T/nbxN3WFLlGXg3zzTG6uy0dGRILhsMhclPN05xCiiaNmbHKDVaSyQLJ0Xrb
DeHA1V+VG2YBCG3vm8ceS9vphySccW6OSPTooY9vD8aemUf1ktrz3dzBI3D65edH
Jv0gz2tQw/gI3JXnh1JrF2Mqcn3VSHL0QO83g+vaHk2flckNUZ9bRmPl9ot6xovT
7v/nypgjIKpj1rcoGU2cH/ahdui5DaHxtD6RvQ83ICCsBo8sYtMPqcrfJ9cgPTDO
JCVSUvMB4Tz4RPG3WYmPMQGCdOgFBS91ekAg4H5krNJ7G/k/iBnHWcQmTGpbv3+z
8Mm7lFblot5n1507PgUlCPYNp1iVl/1zQRJfJwUIBwEjAjgTl+1opciKy8eNMXTq
u3lbqAVD8U3zpZO8EacGZ/ygckHEcdRh4Vm0/Jyr+D3xRRk0n1IrO3cQLH3X2Wc9
ykBFBfwiN4f2UZWZ6qjDcDl6w9t1mMH/sCzdYJb0JZEwLD3FZOOl6LRnIy706fZ/
pg892J/Zj7pCh187r3yxmIxRSiif+yufPh7kG+DF1hJ9ulvu+0+ZBXBE/HYVmQgX
GSfTcjae7As4kf3b0zLkzQbYj0mBM1RIRBoO8GtdfpaQCblT5RafvEJuhFRpBP7B
4bqNX+VYAepvqUq+CkL3ahDPXSpKnIyR8u/nfCrFxSxT29FRuewXxpmH5qR4kAAo
PEhV78U+c+3dJb1QHlUib2AZ0uXcZB1veasB76y3WPTfR//EQlbWR1Ur4ZtN+4uI
lPCiZ/BPqKkBzZz5j8zMdw6Jq7FAeZJx8nD+4mPDBx7TF15MkcJLl0Ad2PSsaztt
2U3894nFnQKsnt0onV4nJOtAI0KbIp9N+KEhDzGzNEqs9ptEfo+UEykAYhn374RZ
x1PZFdpBKBijopSmCoJE1mhIYMkGRoRUkV6/5d77PowVN7yzjoaofgw5RWSD8IKC
XfXexzX2QOzcvklmRaS/GDUP/IGTA7nvofUZ5XxWwg5m6ASnqnDLqQCQ6o1eRTic
ExrhLbI10MxQj9CxvZtmWkp+2tklhl5Off97fRKgAANP/au96SDw5sEepdZV5XNY
Y3AuKWkIjqKGN9zwgfwwJph5SI+cbDdj2D2CASX6YrDisUBL4DY9e0nNCg+ZgpIW
cGgP36Xr9ANhV2s9ufqMQY1xVutD98ewENE05BknktSIQHuzoQo4ti6Wuvg1jeT7
dJ+C6PqIeDcgumUZW5I+eZM55rWKVH5P0v+Vp2uRheFsgzjrIpIjq1BDB+LUpsso
tPaKQC8Qqc7EzwNIHxpATcbclm7kSgCYQKdZt/SwQKHBeLRi+KS2yPrk3qOSU6zA
tFp3sJnz/LyJe2ByxZGh+ad/MDJArDNnCa0w6XqssW7NF0DMxEYUUIQekonBOMEd
GYVbFP3ufnAwV1GQd80N34p8bmiPAJ2u/wggWSh43MyAHbpiCPwHePLQye/qI0LF
uW5/NTkaPgN4JcIarOf0pvvvXqCOM5o9DX//zKCkYrnyBm6O0dgyXJvOziyqzLDk
XQupA0jqIAZPGCutrIdD+RAGwUgmrK6ZYZc7lpJL45DCFV6/FCI0ImxmOediagAc
ZbkwXbwlCeWnF67p2IUr0Tjhd4Vo01TbfhM+cEl3pO9422M2XRTW+6UgAcm379G4
ehD+Q4tfuGIHr7uOnty8fNmFo5HItpLO7cyMOFIhGf944Pnoic2F39+rvMJ3YI66
`protect END_PROTECTED
