`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
73UPcsVs60p9C+jApdx/nna5J8fqbLpRTUdQEorMjgWXxZueELWXGH7u00Qlq94o
7LWVB/STWKGMTycSQns6YdeWa6KDFGkLEfywd9yqjdSsqf2d8J8G7EBKBz7G0VH/
eTJyl8rrH2ctjdPMZVDY3pEDEuhZ/fag2d0lyrFG0WP+5P1ciq0qO7wNN23stnoW
JAceRYl0MchNWA7vbSg8zaD8cv2e6twLWcVuwuivau9YT7KZd63gt3w1RpsKlUJK
u64F82x4qVeeN74+UNVb+qHV4+fC69TdA2TtTXWgxoMyeDLMDl0PqJg2fo8T7sJA
u6Iu4UpyjMCjjH0W5+FrLWVaOp/gBEerfxOGKY9sSTkV3OgF50WNDJgVt1bcoB0i
yLif/Y/sX0qxdIUsNngUnAjf0optSoJKGc20HrRYuzUUX5OeTNadPgg+ZRqYXv2K
5jPfwS8crK21+lIJ7gPV0s3tSDcik22TXRcvNsbfOPy1bR57TZ6d90nH+SV9AKTD
QDuPyuOyZSIG0j1mmPfjPxz/gsvpRkP3Ha3jFN8AJIo4oOi/I+NGFtgJo7gOyUkP
OgSNVl0PdrJLv/1jR4BZAN7gWgEDlciTvg18+sKzl7MjyITKjvM68MM5Zl7hnZ+L
6967VrMBhznxFhGv90kaGUZrpiHC6jMJb74pz9VrraqG+kd9XPW/NcLaB2Wu99ER
3mWnrvDtc5eIkVtmpYD/JwCgtKglWm770rwD3PbEc5bQzkjYkKRrYIEbbrtlY2Os
kalRC8EPPtc5xpQPgvGAZFlkgpOqF1nrErVhQItZV5UrJLBEWFOpbg97gba/fL8C
KH7RKz6E5BmY3p+kwQBcXnaqCW5x3VYpaOBTJykZDdoAu6rRuCVs4RIBu+IZoOIt
0LsJ2TYq7lvqtRsan+JGwChjBP6nyGOEK+SqyCM15WisdLcijRA9ymYrINVrCPJT
9FTMsWkr6gHVaB46cVKgNbOIilIsJhBgdZZqX0yINTxtAy/zCST9G6sHdv+OR2L1
jhCo8w1rCEbk2husskxGCFcIQ5ZmkEfIDyzw0oEL7BnlH/6T1ZbqWp54NTqBMQxH
vMBqlcHEEVfCeadyiQSNq6rivyK7F9vcwhZorebI069Qvg27ihdTqwz02snhxtlQ
bGpwvGbgYRG6QXsqIYBwJUwAKZpM3s+CY7n+jjbqKvyexIbqiM3KFjRhTfwIvj3K
MGUdCBT31qlyTuCgTZdxeqBcIEjemHq3OSSleJL4bLOdEau+T/rPjLviEejVLKHX
IoytKr0k3ye8naxoKLdeVkMPTMWHmbfA2O4KY+vfTrWTB4qOfWOR/xg72XU7TFLs
9M2Dq++W97YSl+zZXSCPSM1QmfVi4xHDKVCtUum8+Tx21IrnFptWY5I8u6rWq/wY
RJjLQ9BBtN3zX+TOh3bIcW+1xeInTsZTIXz3FjU+FX1pG5U2Xt6pjruB3dxQlFDT
bPInc3EqrLzzr61++RU5RPyElC7J5z+Uf98Oiz9Po0MvS6IL0IKzxU1GrZr8Nybj
+PK45XwH7+an6mTtKOf8+mmdoOF+ATZo9Gs8c1BBt3T0m/5C3HnzL7coOIvRp9zO
X9mt0al5n633pQCRDaHbvkgJ1GZEG0APh6M83ALvVSPGbYvLL1+8nGC57WT3dRyh
ntCvBy+3/5oCRsOV7SURTAca3cpsYqubLuF8e3rklksABkoBhXm45Lqu+jdxyc+F
E7m/On2IsOutVQ2MJssp9ZYBN8jK6otCe3ejISYklUeM1Abrpb67n+EOf0fYS/tL
vE6+EO4tLAX/sJiZfsMGKtViclXgCy8Itrvm51ypFuOpAVspJOuZa0s/m1ZhXWEd
AMElG9K3FhtKeRVT5lNCMms7D6Y3Y90D7TYiXAff1QrPd/KkBBCi9ISs/cFGFHUA
kXa+3hUwyrpftPjv2wDol9ZNxm9Ba2T+XVHWRKTr0tYra3hMjt4BLJMOjEkKwKuj
Lbr05i5citc+Zu9Gn+A7zOjPskiFDfjK35qfUKKT4/a93B4JvCgi+0u4MvnaOW41
wKiLfAfL1qhLOFwMmK1gaqGDFy1lFtp/GCPimmeULkQnwkLCJgXfg6pivBSY1bYf
w4+QRHWUSkf5U9TcmOSU7R7HzeMabA0zI5E7eis0c9dSTizWcL27vxdi8XZ8uU8r
9B4Go37+kOaQ6pU1AlpfJxSxZ2l2bPKaSSRH5W7iB7qQJGUZsC+OBzfEctrs6k4i
tgw7sdsRQKufkPOwAW4rgTMpXDyklF2+lGJ/r+UJVmGfJIEDH+jXltXiAlL44VlI
uNIVhDyHuI04xzcE31piZmojTSymV4PK/sNVMfpArxukJUVN6I8HxTcrAVhHwWZh
27yEo7sUi8UsimhW7kgKtsfWOdZjcXYEam8pl5OAdgaoPHQwp4JUcRu6cLOqgSt+
IB4eTSeTFPbaLQcXBY49MkDhHdNM0f0YHRdaV08ITBWtHPyOjYJV0Re//DQsNa+y
8qTBwMF09DSmUKoKOlKtPQO7Q/LvIwiZUDwNzPBKc+lXehDnLUBMz9haPe5ohlzU
KOjxqyIShz4Dqfwbb52wxFqZ8HSCZ7dh12pYIFejHNomDYfs+zFtq/whrQ/+7J0g
fzd7d7pQjtvv7p4sVAU5oP52taDZugv98afTLu/jNU9/3pSEnkZofrh9l7OMRUbB
9QJWVAqPA146WFObV1NE9vTa87nu3ADaJL0Fmu1wpDe9DutJprY2Rn71vs9JjcUS
mv1kpbzUvyeHvymakGD1Ibw0fmZHkfFWzBdoJSUdK7vDacPwOqb2qzNU0vuEyFpV
XD2kGqO0uqCtZeaGhKTwdGaZxCtGIgSnujxjqtFsKpWjugEzVcBbShjPt7dS8SnQ
Pjfu7sIsYuQ+Y5/jgiI08wRe8BZjFvHL+O0LTW1c2u9DgM0UIbQiiF4/Umrc9giJ
1ld+o/Hqvt+EUdI1wT4NHk78Z0TJ29gWuDJQzmCg7etZLO0cceJOghjS6A6q1WkS
1y8pKYnCTimAygEodnE5h6nEzuTw3PxVazWKcj4x/gazKYhVdTzZKXGBrSzzUKV/
pJGhO0RLk06v2xpZ+ShN4unoAcPbrmxMZkwSq8A6sBdxUb+rBu55R/Nm5tnbgvuj
Mlw+OE3sGXtZ2F93StUyYxMNED7CmlSOlT8F7zVFyWEXEVGXrjD7If5wvDeECJrm
hZexaPScqqtuSnCwu1tOPRKnZRCJ8lAfZ4VrgYpe+DzzUv3gFU3IHIf1Zr7Q9eKk
vQvWLm1fTQSgMSn6BjaeG61CmKpmwPodVyFdo/XCIf0=
`protect END_PROTECTED
