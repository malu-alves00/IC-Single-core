`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AANvK2Pff1X/R3MWcU1X0blwI+FBWZucuk9RKPYsLJhcnddE6kjW1TMG+hbUK9R1
cOHqasEyOSUXX3EPQRNcvD6jSRphX/rBIvKmbAEAllLVlKNQsXHe04+5dCqwCH0a
qhvWe9oowwHJwKOLU9O3SlmXSSCb+F/ccfNvqPEwrqQ7iLjQhHXj7ciKCUh5uCz8
q2mwzhTFTCpNpKaqH+baebGOCgnwHwvgLqVyccACswQWLKsA4L0cvFYqJS2yWise
2oYMHm3MqjMZ9rzERWgIVA6kvYR4YNbEphj8wKuWQYgBTPBhH82CBoedvJEazuMa
e2JOYNJj8cw03qBnhtznhwlHvwwAr/mjfX/oYyb2QdBbGJ+YYEWJRpbE2Z4hIHP1
T+Kxp+9KdH12dZGVSPjzHvM4RUveD9B7G4bVad6qMLHrVyV9rGMuRYmVugdBIIHl
Z3MC0yP6wXq7CDPFiXQ4Cel0mm2F9V1Y+Scz0jdtDP1TAjNzgei0GE45v9jku/hl
tnLMU4balFLB7tJcqFM/Mg==
`protect END_PROTECTED
