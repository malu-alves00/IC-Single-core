`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IOzQI0kG3LyjReWc3rd10vA47eCtMq8Z/8maPhWHMwzpbTsyZof/8vF//CYRp6nm
Mg7OW2xPqcQ9CNO0fBAPmAkarzEDtoZrDdqlGyrD5lerQxOz8LVi1QuvMEZo0OHV
cw50NYe7ZeNiZucrjYHNh2t90vGNmMi9I039k30GJ90ylkbIsWef+vlD3bHmARfX
pzdiuUj7XhjCzfDnc24P0SNTPwvnOjZinlNafdLSF9cQRRIAl1/VIfumKnqfLEa8
9CLBsSx+/QAHCKV5xlyUWWZ7AuLS6wPIEc3PIBB3wizo7TphvfuSTp2vzecKIqiD
+neJ+Atr5AnScZrpvl03voXf1NX1/CCrq36uB0Lr6YS9bmQS6qNBzZ1FS/t+mRp7
6IBCtsDTGbrQ44D41ZV/Xo57d/WPOq5dFwS2WYzGgX/8LtREA9YSe9gMSe3U98PG
likSQg+yZTELFgkVPWw1sIrDYiq5lyYBEhpvU5gQSj6nOSRELls6B7yUPYPRzkjn
989F6CnohDTZGYf11Jkcnf/2JtgVoQxGg95xrTBJLB2giF/Ifxs/RppBgajQcKGo
Iz8ij0XOHLK4zN6G+pKARU4vM0WgozrlbFHayU7MZrbhylFVBv2OYhzlv2oFPTQT
cuf1jgq/wIVQ0dXkZ26tfExStYpmKmI6L6SlRM9xKfp/VfvGKek5XG1l9bKYHu8Y
nqRlO2I9tsuRYd1PvcEjzlSu0LJV5hWD039fy4Eost1qKQvxd8vZLGcaleAhzTAn
uWQSOUBu393rEVUNsmoKdymlP6A/GC6jBc0tIWsjWzl0csQpo6qwlcB5fLPVISV+
t5Sf/Xk+DMwmBXBS27bBMuKgXXqj0a5RAqypzVSVP2IlpO2objYz3OrE1hOpx7Ml
OiN3K7ZBvyF9i1CQxs23kzIdP4uOA3nSvHgriwIdKXukBcid+H2PkQQCLxUHgYdJ
bD3X39MZmShAHBkM78ze4a6aTj9esMcxj4B9PAHJniXhpuaQetUotq77fgSrJtbQ
OVYxMR5mQvhTWOhQjuaJgYo4Zwm+i0zzRDhMrUuKIc6Xo3Rt6xikMgKFKtSQaLa+
jck3blgYM5ap1UHR9wXlVn1jFdzCfNyDRkaG1jk6t7m6JLSh7t3K7lQqOCauFYqO
EapLvBN3/mXO4OSg767rp3yqVFWfX2Cryj3muixTBqkqjBNasS72eRvct5nueIF0
kU94OP2ycfj79HluFoT0VGKuR9r2pF/1nszyrZo2IJUsUD/Xt9bsJ22RE/rmSKpy
aWUZGtv8RCzZ+XhghG23/OpwUo6VbfrRtyUvL/YubJ2R3srZISkFCU8s9AGUriBU
NXA9DYDh/z6k8xZKDsESqo94hXu+5DYx9PUEOKIkK32ziZ4XGUFck4xWcdUUzEEt
KWEH2aq+X4EVkRKXiXRhfVDg67vM0W75uVsemaIJEuDiv1vovHwx/p/y15VkLX5f
of517mrcbEVFCQrIOOjil9D0G0+tX7BouP+oMVFBzXpvr6jw7UctXKuw5niP9N1e
8P4USm50MS05DxbJKrkXvV7P2I/hL2hqnVKp9H2vn1CS2oJNlu0BU8xUIV7LfxQj
uXAaFhSCwrBImsi8lqT5EL43aAHZFlGBTmF1R0VSdOuYwFu6yygVm6nCecfiqqAP
RLE960yjD0sF9tnA8oIhC64pOH5OLXur28u083KayX2Oain/85v7mVr47aKpWnwL
dFQzuwEu6wCwslz8Xkz+RPrCrWIfzk2HtVmHwS/s6Nz7uIPTMx1IBRuvmX248qex
Vf+buj4dF58UDhoP0gHHLvKO7UL7aBbkNur2Ju0b3yyPcYk3I5n/6O/bTN0rZd4o
YmYkGw0RFN3SGS3jbZaoTd1gBwCyUALrzu/XyCLOvPtes7ecXqBn2E/y4UTPajZs
MYg4l8YnujD0x6xkZHrrsuRHYuvsnbuXBV9OezSMVcKGh1tFQB4J7VDt0JQrApP5
BiOHgBx5vavUO1kE3uji/PuGqFQ3hG0jVoI0jmBISMPeEIHQB8swbcckn8M6dVcO
FUBQSaMTlNUyhynRTd4Ogun2/M1/sMSTQCOhGt5EKzLfgorAt7IxtX66XEk0exsY
OwqIpVEF3bjY8QmUewN0RNLdZYKkDGljjoUbgdP2QFZdS+Cxx/ROdZjNYdHh9JJG
ud4ixe0C5R09mrhQ4eWJc+MExcsdi8CZz30c00l7COetebBalNWpZNQx5HqjVHg+
IplyO+8yneoV9weVzkpIl2h8QDix01EDeynZViQtICUPrGlZa6hd4Zw1w6XOzYDE
Pxojd/PaBLKXfVsoOO2z1cu2/t68flnltP9UDkKT3HtadPKsJewCINOGDuPkiatM
zUyerhqH+Zwp0dz537hGpn2/pjcQmErIK0dJFoDvJhYGYY/woorQP11zI+thcE3r
`protect END_PROTECTED
