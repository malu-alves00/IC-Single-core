`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GTn7Lr6Kbza8jI5e2Wl9tSGHFjoqaLUgaGkHBIFSlI1PbqNxDBZL2LabsxlYH/jk
M2fm4mZ+3novsL1LttFNKKJSLtM3aEXo86si+GqGENru3Wbc93NfFmh2jUIyXM16
F1BjdRNEF45W+IB2yrMSyg6tdFGQkMeLlHyMOsJevfp+f2yar06Dpfyjx4kdnjss
IPH70VvBuc7saXE1DBP0B31vXl/K1LAdWdgCz2h8WkL4cvCxJYUVWP4tn3nRekvT
U30PX4kcN8nu9hoGzhwvgbFBGFpNcZYgHL44Xw7fk9c5xC3RU4zS5NXwiQFOuwxS
DJi2CoAD/SuDaGY2Wh5wuy5QEz4cGA9CYDcFl1jFrBuE636C0E7+qC3balYOjtc+
SznQhbKw2HI9Bk9xJXfYsizNKt+OuGM4oAvMtzNb4hH89vnW6pkXk3IIHL0wr/DH
uM0kKFQtc5AFmUpAEfWApI3X1hMBnSzFRA91aS9TrzcKqbxb3YctNcMr8iemIYrB
coyhHlbetoiH7HU9S1TZWaBuOvxoIG8NyRIYg7B2zRjNq+n5vSr2sIHOQzAqOOmv
LcB8G2o7Gp99A0LTTMY68UzGavH2KllzaQ7K5hT8enCwYQB3nXDC3DWiCb9sDctd
+xAmTrOUcD+h1TAsPmCRl7oM7rOPNdrwFGAN1nSplpk5CirPO1pHihp9jB0vhbXJ
vW8RuR5WLqk8yOaPspEWCLkmeEqojNob97x3aokpAdS7ESX3ilWxo4R8NnXQiqPY
vTsmvDzGKjwVXL9jUXUHzO7JBizUQndreSEu8gJayacXXSCr7Z0r7hAx0Bm+Y12u
MINNOQu5k2dt9fk0L7XSdSJEwosnIESfvT0yPBf+/pfZfDsztmo1YSlu5kQ3dvJt
O1D4OCUUj4Gtksa+Lkmwp1wevjqx+MNrJLH/DybHw//+VScqZQCYfMOamkN8M6Hi
FuQkD2WufcNqkXLdzJBKfPA8qKeVxxMMxs2KDIsmzdEhO49tIbyuZDOy2yVfCjsg
Ve3rHWKv/mGSjVOv9I5X7uAXlJwBKuib/6KCr2wYJnlHpPvzEvtjBoeiPtlJhVu5
cJbBUAjO6st8RTyT3OYwFGHbAigAtT2zWNne7Jk7CyE5V2n29S/kew18wuyeb8LE
yPq6EMx9p1OsjWVvvcknWPpk7qBigipD7QuZbavmXiR2oTVbYuEimsJMgdAAiQlo
ZFImsNLrfikIgL0qu5JxdCe5HGVgwIcVu96AzPGL8hplkQRM/BRZr17gKSZRaOag
8AZ/bJ83wb1zmvhTxJuehcZbdm/LKqI4Lrj5aRcqsqFIUNU7gv8OA8jsa+EoOITu
xt8MK2UO+MnKpucTknS6wfcSPneLFmiEQ1QUUu2p3+F9a+1FnLv8/pM8nZXvdkgO
u0RX58WDVnn6rXGsC9xgClqRLocuBcjeDe/5mG2Uo0dBsqEZqssKV2AaktAAx+eT
Wkr7Y2baKprvYw0uh4pgr9Pw8jad9NhyYdK82N8xEEeBWQxalJqYLk3KCu1Dm7UH
r+yNsB3tLiNSJQhQ8Qy2S/sCMq3h7x2+t3b4vrMfUU3BYtMRlKcKE89hNPXexwtN
oFn3m9zQaLISXI11k+tod2TMEIlR/bzeb0u0No+uqIFtPqAvvaZACVvQ28R+DGwR
V43HxVyKIzklfGOqYb1Oimw3woFwIFXVDuUpXukWniEtYjEPD3rr1uuJz4hBIm+V
PPQZPYhwd5pmqDQ8Oc+DM7mgUm7A9sPvlMAYrPv7VDXOJI5fiXksIGp+4Cf8eKYt
B2duHPzDOTETh9MDjT3dKF6gmhRAmM/QtWzpBSGsSUoDnEKOITYWDA8VmujtpjYp
/cwPcafH+WJWPL8XziUJTC3QNxwnq8WQWCnaEVXqBZkxs3hKqozkEcLfKL37OykI
uaSZlWW8Z0WfxfuDar0c4FWxysNbURzPeWlk2D9DI9Q0kcV8Tx528zAbDN56/NX6
pvU3lSeyAACQ/v0Uamj3VSkm9Zfb/hK/5CmGaFb/zzZFE8bMbMXewlcU1MPb3lF6
nPQaXWyC/1iwq7QL04NFOtyvNxJjrWxk+l7ZqFyjAWSBp8m6IH5PbICHTom0r4zD
F7mFVmQNO+89kdiVupJCQEE5f5V6PjsQLXSa9HXfVAhRhpYRMKhVwBx5kxiz0huO
w9rdnr4UGqx9iab6hnrwVbqsKr4olrt23mNugUSgi0rNryTXhajYeKKcLNViPwgX
eJqR8yBTuCmOES7RcpIiehgK7LM+UPCC05AtGrOjKuZSD/IpRAMjNnL0LKCXw3dR
OjzCbMGlweokR9AtiGO98CJnlq4HPZqRBGjdW9zdftPoMcV9EDUxx/wWK8avoLfT
rJa4cLPi7Uv9yxNqJImEACqkqFgxidPLBATxodjz+sxFqY8GnN79lV1h/0AYDkqH
jxIrXom8I+AyJ19cxAIQsriMcGX5Cu3pe8m1Ex3BQ9Db2PwpfXNtG695nwGXpfVJ
excinnOudHg40FecHt04ysK7MrV8CKbv2SH1WK5X6/Y1VssefIPhfrONOgePdD9V
N7uMKuWG74ipHBKN0Yf59JmvFM1Y0kKJIgySUMB/njIIB4vHdXD0ijNk++R9/KXx
jowhX9ZGKBBJudQ1Fsgy8Xk5tvbYuHmxI6eDnG8q6cjZcJ57wbBiJxXS91H7sAdf
j7Qw397yqsRGtpe6YUIofODmsxo2s1dXYj21UMxaAGNCBQAoU6IrQVlyms+8s6cL
QWRjNBFko2qgnwH9kOt8B6nmuhijAdv/NmXHOQRa5jTLUPcOq3KXRUsJ2lipDfI1
pwJFnDMpyBpI4OZgLv0fx9Q8Yov3KFoUG6P0Mh0CYql6MvevapxguPSp+vE0oMZg
eJgWhJ4LVCM+pn+iE9JER0c2RhamUdDepH1GVak17WBL+mHg+8zAh20/naQLvRgG
Ot1o92ByVKyO1fe/Bqqa7M3LIZ7KpkxatQwINvErxBQDfJSBXl1rNMNlkThZcEns
cAz19Zu64EfqKJJUBnbH2jNRDKzcHExMN+dtLkYJ+pIxhUznh3jugqMoB4Y1D6bQ
2zTWEconiKjb/oQbBbSzXNtxUM1LJgfVQrulouA9TlfJyJidNsfn989l1EHiF8Wn
g/NO6McP+H3sqXnf9W6pscAIz5nohhR/M08nNgaNdy/adkUKmJUJouvWcgd9j+bP
oEoub2gNE6BhuWF9z9B/AYu0Y38Lr4eGLiI5tY4fF9sCE2jJFxQnbrHrFekiMTlo
1Apagkwwl431sJ+ytDn6wGVuB/hZm/toJgeY9GWhCMeMhLVbTuc5wOqVwY2SKqGP
0JeezHMgkfdR/WZJgoUnkaAO7x9fEDIyw6W/uyaxEy1uKGkrV9Gj3SFUIU4IPQUr
NCW30pVBNcrvY9Hg6zjme3Do+9wT2ppVugdyO2ei+bYHxZYhZYcWvfkNnIBuHNpT
2nAMSwO1hgronWajIBoXO9PArNguAeYvvxrBMTBzA5QAuk8k4aRSzBEMPt/6OAp/
HbIJXWyVsJ8nkDa9OnE+wKmI4ldNl9Ifbh7bJUyuPQvuEb52MSoYYsXTAfzf6dfu
eneWH2LTmWb4Zp3Gu6to5QlXUhuZBLVZd3Dy+3dHemrofazgeali3Uamy93zbcDb
GXqMIXwzenLWpHSb4qJquMEQ08gFfzjMNCIXLosSRbMT1Ivb7gUsiNsDyhAT3GxQ
funClqL7ga2uo6YChpuuawdP/bic/mUIy10sslJ2fokgdYZUGf0lcs+E4vMAV6V7
XP2OHK/t0eNT0PfGYEHnP+1CI9kvAMzpjlZt1qoiAi35oGsOj0HcrTiBO1EDqj7c
xMPylP7yGEWuNed/Aqn3/aG/GHa1v4Q5mj7CROpaYReC70onzWAxp/pZea5miWRY
iXel1auDkIIzZER9RlDNLV96GHPYfpZxnDtUrE78ZCTnIfCGvoXGEXSMw1THoN5I
BMaApSDJwU11aK7culdo7JhFs97UBpi82utZ/+XXmkcqEFZdJLU0kVZp2pz2DLbJ
F/IHvch/k+8vUoZUKjMRaufpMYH8VZVa0EYT7BpK3gSWBh19EXiMDN5hFGQf1Sp9
fLt9OlglPq8hYh1gMO8XIT6EUcijCmhZeY5Nm77Eoarf3FHlOY1v6TTPqz52AnYW
XNg/gQdsrkIC2w52pzRcpf8UZyzA8qXnl1+DbW827ILKUvb6EibHBWqZi0GoUpPP
jdgZRhvTymQDBMWJ4jdi3W8PuouuRg7xLVh0DQJaPGQqOp2hB22trB6MDVk1WWWN
B1y6K/f3gE0Z99+zh2YPIM9146qJ7OZHEhhZ8FBqkhuZmpNpY0EUTz9abUDR+i9s
EMRZIo6RLPS8zGCmb/TJbelcVEG8ydHjQz77YU6aGfrwK/HSHoFOrZB8KNocOh2L
ELK53mPT2cH/CnuLmEHnkQykBITq9dEbfBOhh7nXrzwaga30tzMtnTo5/M49RCqU
HHTByN+B4O5KZUsSTYfZsnW+J4yJb3ErO1w7vz8wcijrbkQjreIZJzHCWbgDkLhn
KUnlp9LDTmaHsUrFEEvOpqj38QzJoiGTF0EnbCcuICmlntRDyr/DFOkOnxHTMcwa
3GG7l2Bx/0NlCSQRKiM4LzFTSUhsTYyPPEeLIlPVnwZHqnA4LwkTPWCiJ1YaxxnD
2j7man18smscVUWKxijQG5MWhTDNHDDq35TsG1dKZ5gUg3AI7mih6beXpL/CDQl1
tWQP8UCuzWHlJTZtv+o3UTkwow8KjbiEv9bJyudJRVAOYZ4Gus8YvSYq9tTnz3uh
WafZRGVVr04gmCtRQj88B9OzBU4oLIMMG7/zMzAaSroI3X7awy5ZIC4TxhclnCoD
/UGZZK9lMHdSL4UakYuTVQJGjpHB/4JP2yfZnTe/5/VfmKFhUIXXJDvN2WqESGvi
BHPCFh9SYbWJCLp/UTgLL5dEdqalxZVwluj1efbH5pc0jACrEQ1xBGvgS1KfEzqe
y/Sjo8MgZc5sy78VrLz2KZssb4czavKpUGICo/yqt91kqwOkOlXxQp/N6RjfdgL7
OxaOqryBrfqXkGG/DsC2D/oT60+rHnAkAbdSUcrQdipvo8LFy5E+2dubvzi9u2hR
fk/c7xCwh+CFHPVnkq2XzDO0hTt/ZluxLpTTHLUXYG7XKGPE+x6Wfzycncn7E556
TXB1usXB94SDGqMeRz9WGJb9lgyVgM7rgdDJmy4gzgQ7lP1yYlE5VGd7WLQyVHxR
p4IJ1y7EnGb1VzyB/X4+D5vYkGPBlQoiw93y5ooGddUN2n5phW1of0bF/jWILCpF
gKmRE1wQ97kReRL/uV/KzZDP9Tc2DlltgGyY5FoG6ER6VSx0CwTBigHKVNPXoOeA
WEULocfRh5dnfFoJNjh1W6NpF8/+GEZAwYRxg8/Ym7gsXXY3zPQNS+/22vhd7ChT
U1k+FmVRHODIatgfYG1TnGerhMr7hBLQdXL/M7+dP0EM/xINqAAamZz3pNmLi4Zu
uMHmhKWNL00Gq0kvjIiN9ghvwSsKJpaU6Zq+R5806DEOwK+vr/3jDKggevIUxG9k
enFDMsfCTBKv3BTcWdHtq53Pz5wxzmog76+S1jC6OJ/VA9b+ifmps75mU8w+PKcV
3hP7n5uEn5qAD0vaiN2jnjp1Ufkkkyi9EoMqjR8xrTniJudKDBcyp8J4chsxoR+s
Q3emKy3Xhy94goArxZh7Osw+qi3Qwx+wUYmWpw0ankeQp2e6YrpwvV0lS9mFoeoM
7fzTTlmSkD4SKYhG62FMKj4umIKbT9iwpFex7GggiHxNYYEaiACwshNtUuKfT6TS
A6wVCeJaOfjd3fZy/OuK6t70IaHk1UqvoHFEeEX2dwgKYygOL3IDqeL8j9mVXlN1
a5l67TEotcvZ8njfoKK+sUEuGTUdeBxHZXY7GyzGyc46kT/mtBA5MDyPTQHtIRfr
`protect END_PROTECTED
