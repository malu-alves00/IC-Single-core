`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
K3WLiCuPWIAbIHfVswm4KVDOOzxcNQ4U4G4gr9EvSUlzdfwN4MpwFyYLYfLQfnwS
mXKTQIqov7g3g1+dsJJXTfNaJ7/fuFva6omPG7xfsqkwaguqW5AeLt7H/KueW3Og
hvbgQB/2azC0+oDZl6ZcUirmICPmBQrF59//uGX6eLdMTYYqW7n4HT/vxyvunOig
jcc9Utqs4w8Q55Svi9bX/yjscXsM/iCL837M3kqz0RCqaKKP+D1SBMOPgNBkFp1H
WFTUoDVi4bGv9VFDWaB2i8QP7vbfNqcy29rFw4eVwAjJnRInsHG6sDDgcAk4+9mF
HPZ+h57yF08TE/iEMHa/epwaQH8SIHKLXFQb9v01Y3vdBeeDXiXS9WPAQUOokrEG
YynvZRWpW4KBqG3vWove3luV3J3yhKEbFM+Ln8keMM7DWxz/FnDNBk+0B46yHRce
tJznjqLtveXERPso89oyRtrKy0bP8WnuX8rxOZQnK5W7IgFBW/GdWvqdNeMqji4n
TPTPJ9sY7bY6pAzk/Dofp0Z3klyKIBzR9/R+tYRfzYhPVk4ZPHeAQZ555NDJK5FG
BenwzIXbSKLHzR44Bf0ItME7xLbQJiJ1cpPC0IbxZ120swD+yVjad4E1V34F6/oW
eZVL10O0Y48eTdYubiqHqw8TeQ/zw4t5XEclYmK6SMm0wn19va6e1vv3ZqDP5a2v
TJCoyVr1Dhj7dT4bvSKmRkK2vjxsHmeX/mB+rcWbrRwnrX+BEFwWQBAzaZT57v8l
spY0ljXlYPEQMl08W7eEsA==
`protect END_PROTECTED
