`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0IUN6t6gzUaI/biK1hfa6EBlm0uX3kF1ZQMRILhAI0IleN6sIK3Qc254+eDrttjL
qe0fwd9alHJpdbwAl9+hEpMzi6/8suxf6RRTP6XnNvhAs2bmPDV2njYQ/5wRCcpG
a5Xd43m3HYZjArTFvA6VyBCE5Zzc5UfLziK0mq+up3aNMBfgKvpXbgF9ov93Vjzn
MytAPulqK+sWEkABWwvohjwhx5QbwjN1sv2o831NW6edwU12b0aCM09Lx18Ru+Qc
lyKR1OXt/7DcAP2A2lf2bmm6Nlqby4HcHPfs/jUae0HLuXQ/gVwfrTmQogOnbJw+
COCuTX6WcqRUHIea8uLzpLkydjYJIiC4DHPDNA53OrLDdIS8JMefGrS+qlfYthH4
KgvmbRvW4PRIf42MpgVm1+uemzqXgxP6ujHxZCfXo03bk5/mu/JYSDmoR6kVNlJc
pCSAhXhJetrUpqVNj0enJWPB0QnpurRuVjcbOhsFDPPihSDAgh67R/X3t8mjcGLg
tzpQ3oHQCLrJV+WFJC42MxSI7gDyAsE8s5Au/Ocy8IHfI06UOyNfhhtr6GnHpOad
R70Q9w2XLgdIItZ4dFM3Dfvo5R15o5v+r11w8y2i6W5aqo6OpMY/Yoot3qth5BRI
RtgtIb5yQm8vRBc1jzjzfKAO572p79rVR6ykz0yZ6ZFSONgTsUfsyxLnEwg8H0EJ
BmdtDhi4+B4zKgFkkfaK6kJGy6nHCyEOl8o9tn5ZoHS1GkDGiD/zI4Yjrx9XPB3c
6DR5v7pQldJdNyTKu+pFQS+gcjgIRI1ay7ddkJAwDeS1OiXHM0uMQKajEcCCZaHl
ZzVP5uCuMiogF0LrtD/2N8QWO0xzvjKKXqONWYm/fj+bfKWIaZMTZ+A6US7DyMVJ
I4dL7JfCsSf8kugXblgbbSrnV/E5qIS91JqV+L4EV4RY0LYqZ1qhnTwLJ4vCrEmH
rMNTf8qMbGXe82Rde3NIZQlTeehzgqtQqVNMsm6Brj3+EgOVuK1b9a70/Zo3zQBm
jwsPmyhzNmq9jPWhP57EsGTuNKh4oNkH0CZpunSDXGRagH935QQFDzLIiFiCKIlj
7qqWMcC7o7GOkuALhVLuUoabI3+IlnwTQpUbyPAIAYFVaIwmdQB2cK5ERAUPYMN6
5aKJyKR8cdkIWvjpYmP9/jk0hzZOh/ktbwjt3BTxEXPY9sc291EpptUuqN+tmBNG
az2M2qbHFdWmQfVJi9XrNVomSUX/hpBYcoA/BZQn7iZ/MxK9l1LetYo3ga/MSPYZ
M/HEslKzD5zc/4PnZv7Ru+KS0lS78ZzzuwrxVqVGKSJIWAaQBRIpWq48PZKnpC1Z
qmPE046/dYxaOy6gH08/NB1Z/OqcCvTC1iZL40dacgan1tE7BNrkkxoY1HSoa9h7
7loZ6o7cSJiv2Ek1xX5k00yIOey/9d7ujOH/wzdEwpfI3rvjismR0ISkD8MW4ANy
rYxJyhd/eFiu0Bn90ZTfCbWc9UQxx1zc4Lrp0aQtO4Jf6LnJn8o8qDqp+ifk+tv2
JLoIoBwLppirUvqByrYjwauB/9p3AIsmr1V+KEuqKD7CS8tRn+opz0SsOItq4Wge
sC1HCiDOn7OFHjt+kLLAJPvUg4wUkA/iw130ddjQieWPGR4vbGte56+ZTgSegjsM
2VU0/W4jpvsVoust9RUCkfkIWueC4o+TMgOL/uUb48IM6PYlAhTu8Tzweydy+HMG
aYUdkK3FY0T00xplVQKCkML9v0EupqAA9+MhPyy4t8feZireRNt4PzESzHsRmIT/
y0aTaf07AHuj4RST7VJ3lVrc+xRpp7O9foRQf9GKcftKy0aDMUQ2ekXV0Xva66jJ
p6aJsvjpJnVmJsgG2/+g5jn5w3PXPQxzj5a7vrsfNLr4A8YxvAlftPj3N/+sej/I
ziHIhjgyRDzCmLKOBnnag1yr6VofN7P0iakIRb0NTVNAJPutFLVu01+ISaH7333d
fShzaEw3aWAzg2sQrnv/XW3vjtPVI7/sGLhS258H9nMzegoXDq+sSJj5S/opcrY/
FXlixL5jtB/8VcdG5cFpcrEdi2AhO7hFEszwhgLHhsAxhbE1ruzHm37nlg8sZcOt
7+m//0ZGcVrrOHvD0VYvcfmrSX2Cn3cRL4+MPlA0ZbWie4kQSYgCC/O7nBIgA+Dy
WAxkCExhCbmN4Qw0ouF4MH5HScEGeDKb+6vCiwCo3bLWEhYZ9PIJyEkUxAUVU3J/
Wu461fiN4n/yp09ZpHvYdNMMTxFh2eBtLsXj0Tir/2ngUmT4FMYfwbO8Jio3S5JV
0khXnqrNj2tnYBxv9JOdDKQkuzDkd3vVmfSpZp3+W+4qxUQWBrN6Jkw8fP5NqLQO
tVHTr8qUKCUi8T+8jj6n1m2lys3y+fP3xSOupXMsGj9r6M7GuGkakAcIgIGyVbhf
dACjQEW34WhWyCO9rC98qGZ472w30cBUq4ERDV66OHCTKmYhvu0uHDbnHRgfT+qV
g/bS03Af2Oh+wq3lIj0ehRLGr09WFNDS1kVPI2p5rWtj4jqp8HFoO/f4pUjJU5VY
fayJBK5g3RdZt+16UTuvO3Yno5/cX8J8MuXD3WL4lNRAbkrdUz6XM0pMAiKuS9qn
suO+OThXBgr63BgJ7ENohxFBZR0P0u0GO6lO3VrHHhaMnusI5Ho3DV6Ef5B+YBus
M9o+sIkIlHWAQSa44FknV7FjIiGD8TRc5n3uEMoKfZOE8P/dRfPxzVMViXpPSXiM
eoycovjfn6BB3D4pQF1ur8F4tHvN+6rYfum25yw2Dg/3jyRH/h7jnyRLZ1x5ZrLn
Up4zMBQ3/ElerrtWuDpKau1VqVegNX0IUHa9T91d3cSnxtIlB/U0Ys/1/ZNKnTEg
3XT9ZgmsACf4mv4Xr053j6ZyK8dA/HtaOt+hnyhKiCAm1Dr/Tc0+QqZhyHU+2Nhg
wv0fEMPb3UtKL/Bi/HGjytGQCZW2ZC92CofMqAprisiooMRQ3TeKlp1QQ2xfULFN
FgIRJkDcrt3aMUPwUdwuoTTAo5g1lw+FW63A38LbbrEqqq1RB+3wIybteuIJQ91O
IIOGNxXrE2zgR0QQIvRa3Vutl3ol5ieUU4Zgzq2j1wipPapOKxIBfJUi9p+wi4lU
vj2rtH4dqkTa02UZ7FGE+V/BikZns5Gj5EWJJWbR/cGMtkau2AIuLrLBRe0LTrZL
RH76ueSstBkT59h/oEJfkhsp9wEe0I+yeYsq/9PV8XvLKFXob1VqZIthoi0XBVfw
vniynJXPHRfq4bDksMj61d8+DEMV3/ltUVyrQshg7c3xv6XCGMPTbtojzx1kHss1
G0X7wRJObqwFYlb0akSgTMV70JE2NG/cSb/9NttKXPnqgeReNwUduYB/BfeFvnxn
kYv0iF1JTop4f05Jr9V/V7utA3ZlR6JbHc4Z0SEDGj/Rhhu7bJCq0hKs7h+ajijR
d8e5qPyEmDjEig9QYipft/lCjuL8MjuLNJSmM0j78wo9cQvmze0lBT/St+qq/1th
AEJJm7a6VJbZfV+MiDmid/p5VM01InTGny+cJjbeY3HM9f7YG0ks86eAbgQ14MQX
e7y0YpKXXv0/jX+M0qA1cDY+UY2rnJH+SeJPSQFl4d4nD5vyMRb/kotbirqNJ6UL
NUML+0F5IrA4XsDLvd94QKAr0ktx85O5spcC/fceD4nSCSAzn12xVFcNUZzPHEdD
CXcTqXNlaISXrYa+yqqlX4aZR+m0WAdq2H+ysW8GWoHZLYVvfkmj7PPu7jcH4mhq
ZNwscH/7U4RncwKDzPgb1e/I1/RyG7eajz+vdZw32oxdgCgyTDGzhKvw76h3KCq5
J6RRgXI8Ls2L7Tp//JOfxOa75an7IvJeoY36oDi3Jybl0kQSjdUJtzzcTCVcBy+g
5iIRlj/0Ameuya37WRgpzCXtAeEMdfg+6bBI7CXyMQs1YxS7xsQQLGAP/HXWtPkV
641n4d5Nc0JB5VYx1BnUo8RffghsJ6tE3I3lDjIgxvCXf5Gi5AeVS3R81Oq1ZkgJ
dF2r+opcwklsRh9w3MeKBfo99a1D+mbNEAVOOdfMBHwQ9wMLY6BTdJ/PT1E6bPps
fiBELhCqOWyvIjS6mS9m59X8aNhhoRyndv0TiArH9U+w/6cvZ2ptamEAoMRDJTrV
7t2hOG1YAmU0QVJc79VujeypbORpGwYIj8LS3TVSpN7hFf9wSPjUtnetvJ+JkbB1
M9eGR0b7iLv789prNvlWGG4sJbb4F3xL52Ukzje+pAXz87Ui8LUFkBFpo12EtKvC
VeA+HJnjUcwp+XRMEe9WDyD3gh+TZlE3V/Ui9kN658KwSnLQQQM8NDGy0E+7ZkdQ
f0VdF4JXtgK8HOLUiKk+mdfpK/qEa9U0ePgW8km2TADbdsS1luMAAdhswH7TOcuw
xouRNnb7Bzt4kzGJa1WjFVAvGnszO3Tx3LRHbLk7hxWjt7zdw2pL90riohC7ovAC
qndkWT8K4V612WMYuhrAglbCdyeWyLmg/z8WvycZYeKf/xKaHn7GopUOGyEE/dHC
R6nJE3AY8B2g3fq8/ebR59mgLWmRY1R3UHHGJXriEtJilMQN8CFTXfOv61OR5S0L
bFRg6pLuGHMUA8ycQBI4sfs4aCj4FD9CXzumBMK5r9CGUzYyHcSlcpeAeVsBKS4B
bI508rdB0I3YBasVq3/zE2GAbJRFV5iyrZjLRGuar7MYVZO+LDHEpUybk9y7kbPo
W36yfiylfzEqwAqiIMSifc6PV/I5zKZryaojY7cFRLtQcFjHF0PlyN3dMkmStp3e
wi30Y8SFK6n+x7MWEN6EvT3oHPGWQR+J9rHRrQWt/IVKKgwLHI9SLoVZJD2QJAvI
V5k2+A28mB/I+2UF0vKyV5CQxFVBl2n2PB5IXxSxZNbosdeJ8dF9InP57GbNRVHk
OmXhpDjJc4yEKY/CbxA4aOQNGjtZ41c5+tNMKWTJvjBk5l8+XXsIFrBpqLfrcNx3
Cp54kU95P9v6e5EsjIXuFTLTsoogpZd2ApZDdDKO86jAsghZXC6fz5nWOOLfsRaa
iqh7LL+lBTSgYxbLJElmylpcNBm1bumqyr5NtYcb4nN4DbmLS2Ju2sBX6+b5eIPD
kWkTSOpLRTjqMNi54Ftam/JtrLPg+HVP7hvBjog/abDmIK6G3z3qspnDA2Xw6cbe
21YOSy8GGk0x9oIwAcAJ84KyOLEqGccEJrp5ZgDdHeQFWSXiVQNPFMSkZpqggC2n
Pje9xtufKCz1LQfoiGfh+MgeUq6org9kDcNJirpkZ8KL8vGYKaPjELjs2NNNJdDn
XSW80XejWsVR+zG+sXsngsmrDfoy2+6z2K+AEPpG1prNcyKbV9SEKnEhOUWtWE5M
sAau+VeaNj5VTCKZ06uKEDfowgQ1c/5fcnvCdOcb7pUVLYvou3C8s2AfbKxyfYDq
wAyHD/NSq9/YGrWhlyMYtLG1cgJIwcQ/0aSBagctUf8yRs8iEZRmItYi4SiqrJ8F
XyvWkHh0YapFUOSC/iyPVC9puAN7w9OR+sHDqlk5K2hJGgiMZrlBRyb1uapQRbsu
sbaE3n7m7szpAT+0Y2hKsmJvkGftNXPhTU7l1Zd9ZOnzxv49cd27nLTeB0T4KaxJ
/n80mGrVmg9Gpgh8dPCqogQtEgVrdhNN3PcytPsywlk/SHJANlhlVJ3vpSexs+ot
jD0oOuSdfpxRUtpe2CWhFfqsT5miFZKVOQnDOyYR4axzbA91zNY9/eY6A6KM1peE
3VRGsAO85wF60fFQx7j3GHsLMlG/5mH6pdGaJPCHSwAh1OlAouOwaDIufCDcKnm+
2ug/FDyIAMSGzcsSe7oqIKfw+2uT04Olr5FZOjyWK3phR+SmacgSl+vdQbqvH1nS
zc6bVZrvaLC1qYD9xQV5ReTWsX1MDelKVMwz4+7tuCmJWYTT9N8uE36nf6Hi5t68
J6ozpCDswKyfMX2t1ADflnYFTEwUQL9dhNBJr0O6Q65AsXKfAqKLVlq6KhFOiJxV
0zFxXGyapP1gNWUyk9E/m+ksZkafm1zYYk/OissPQszn3rRrkIi02Dx9sfUaC0lW
ZTXhZkVhIyTNeOg4XsDF2unztD2DdsOMAMWkKYarDNEzAh2zxTieOMLqOWY2HHS1
2bcPvgH43CVJJGX+2y0fLxzrvLlUc91BWjeBMx6XgXBcGmgyDqCBt7J2QndkNsan
PIaFGGDZp4weyoNjaPaqi3EgByknsP4oVX65mbn1gK80CRhigXuXldoE658jnu0I
a86HefHdkbKZbNPFOURcZtX1rPHCVn5DQ7evPj9NKq5Wz0rzJQvllK4nVCsibdMi
RpOlYeql+hiKxLl3VgzUY42CaiAFYc+XCqbdhTy8BUfIPV8LHqTpscLYuXbOrpwV
sJ4g1konveKZA5LZAXYOyVKpDCEhYAe4vZQU2dQlMJ3cA9ZLFLVX2oXyFM+DAg5C
zYx8bIPCvEMBvf3kC8cH9AxraN6DrCVCVxEaNuwld2NV2K9Zri0BrUfgn/wYdjU7
9vnayIc2n2xxpY3lqDkyCTJZm1+7hZZvvX4z+yODifoMQGDccnLabelaToVuXWf0
Q+OPLX7dwRPFRJ5y/C4DFSziGsEdUTciaInMloHRHs34oQn0oG0xvXBRlajHfnVQ
3PfKe5krexRPqmnv45ZYSgK4Lnfm89u/nENlMy/6uIW8LnDDYZwDZhdj7itRaxc2
LHQKK38Y/H0JzM82yCzfLPy2jVTDs0YAV+uniayzhYXVjQmEF5iMGa7SJh/j0O3T
zV9jnx+a7qkE+BuxdUrNBbkpvWUH8ghYNQabsZ3tiMGEhGNXJU8Z6awuHhTg3emW
8s7tX7rpJsdP8IO74dhPeSOOrvimTEKN7PN42A3BggKpD1ipld4vqr30x0ceyOB0
DoIljCTpOeazpKyzjZdSCShoqHAX3KEzyXMfPHR4LukoOuK7t+UjueICJQ/tj7AR
8zZFF6saaTKrquCvs1rp4FqP83WFHvU+XGbIz++OPETARRsxU4bu3eEza2H6LFLS
wSP2TvJs7axGoEz6BZAUydwAybRRATRTUCwwAE84q5Q13mCNP0rMUgdRtrFH5GVK
I2UG7G2L8uTNI7tif6YjgnxQy3GMlpTf26Hqo5Wg8lFdqmDsATy0V/oezFQtlcNn
KwNPCR6oCgFOXZU5jbaRkHcbV1EsTMebDe1ZcHFLXCTyqE0dEINWc/wgV+z3+GkM
YK0DQHpQPuGWKYhWZGziH2wXuhMx2n5X16ZU0AMVsyzALqXOO9q6d6h3iIh3ZVF0
chCTAJJrJfbiVEG03nsLjRP91ieBqT3GTR5ndXwRmKT9bLrcsltNhbF5AUi4x5xL
NoLg+tWZDIR0mc+AlYJrnmS79m84LYAZKb93WO/R2fWtXMPkDdnCwZIZgnnuCJOD
fEzfL6W94PyOS5PAZKUK45QwZnZc7H15Zk6aDhKPgwkDDg9QbibbFIx5eOhdYsH1
D7j75oJFY1xdZESin1jSRCJ0ExVs3fIV+Nb40TOrbrImL0HDUaz0yoPioN9yeMLK
5Hue1tGa/ec8yWT3PwVVRQ==
`protect END_PROTECTED
