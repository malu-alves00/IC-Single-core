`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iphkOcExkp3YV8IJDNMF8IL7oxGve88BhxuKcB0EG1L0Bl+DqEDEhki+BcoN4x6o
Fl6bYnxKTwBt1iawJN+CrgOCw2vGhMvTqn03KeG//V9ZydQEl8onM4LUhRan4FlA
khwBN2ZcLp9yS6yzwIhzabVtPAmFXNO01EalogrIl3qAZdwXT83SM85C7pLknU7R
zcjU35Glq7xyNfPN+Z0lZADudaE4bfdaXFI/QubVrIL0FnaI05xAjIpQjVaN6tkK
RZ2w0CEV/QhlrpEbEmUJ7dhGU6KSvYOoiwXJIxA9lZdpLWfmBWLrGE/Fd4YFwAnU
j1a4wpFnlr5SxsA2EOxLP7zHDWHKEFPqvb88/y21VqoNfXTxc3IwF0x6f/BmkBvv
KpVMoETV7a+73/MniOczW4jfRMu4hhLVYRYr/IRiLR770KTK8SI+3iSGZtOzxd15
eKuy+2gtHwd7Szev57C3oH+ulJ0kV3JJYNZtoOBreM0aCAvag6rE0MP+Oz45HeNb
C31KKldj+oJl7XomN2okrTqSrGQQeHwTEp7/YHEBu7JE5BnqXnCJLhuhPs8Jj0AB
NHqMTjOnn3qnMIgnjxJ38ps2AjWjQmR4VRBs3tL+UThz9wyz7g5HvQo2k3MpbvAj
kRUSrkbWjRSse2TmJL31bSKdZBZbbv596t2OPe7IeV2TtIpsYppIxXNWhye8J/g8
T4yBDU0Un9OAUrpjW9d9n37lNURvTlME9+7fpwg4vR8Xy5IcBPw7pkGhk6rQZiuU
w2FEaby8U8euLq9L/f3qNHtgVp5aJHfzFA4CqHLJ1K/2CL3qSa4LPqOBFrQiBWVJ
fT7KSuOJXfru609cZleWbw2NO6E+SoQJm2gDdcp8gR3WfsK3VownHeo9Xw4M4wDr
ev9RxUusB/dIrLilUMzh8IboyHatgyEx1bqOz8/eTOgOw1iJDigS0m/idnWRKVeK
/ZTJdVIJJZ44WgHBB/X/SnpmFGf6io3PwXQ3RZ2CG5we5/omzOr46P7DLmfNi3iC
+XZBvozDup/b1so99/ocsPA2XZQQGVMkBpkf/eQWAaOoe2mPthhzIMYLGUl9hBo0
YYYWsgzx9T2k2w/ZA7jIDgB2oMr1xhzVvYJ3KxexscnYLYfo47y1lFL48JT7gTYT
WnZmL1E6eMq+pct29DBVi/CqUDoITzMOdpg67d7oCXw+tXztVgRkusfQ6LYbG3i+
ux4K/PsFk1zDNSYbejoforqSU1WS2XzzTaAATUZP98Uuf/fZ4BQxFxDzStCAMgZF
wJICPaWRrnAL7Jmh2KbwJoPSNQITM3MaqlA9DaG4V2Q/tJfP+o2NhfU41soGWkTH
bbZehwIp++tO+ka1BHKNIeDbJCCK//Xp7/7B14+BD1a1cLav0eSJRTW1pLEU5EFP
xaS8Vy9i1flwyQB+7nBeIBlQfzzZ9hi9FwK2QwIC2KvlsxKMjuw9ojERY5TTGlUO
lBLtLowXh9GgKf6NUiU0PYHkKYYqeG0BrELWo4CMrJkTAX/UP1OnFPXebfWodJ9k
4CoxJoPGmnxLRlyPEGt2siSWDkDuaIu1eZiVuGmFXF7ivaPqpQ6pFxQ7mm4gTZmc
xm8qAVwXVL+snJQVqZTO9dboK3lyuErE5zGZIlLrC6gkJNwTn3EHSjtgj+XThzy+
VlncdAqhTyQR+GhXgyFlgzcE9hlSuHX2K5kwqPra9slvb3E6Ec9l3nEL3RNlPUf4
lp8JRMB2UbgLn2SSwMuaQ5usD7HL24Uc98jU4qjnKiQls1LyubXW0u90saL4jQmx
TVmPHV4g7tDU9cTYmkphItAOwiwGl6S/hl6sOzvm8C+9N57uDIfOyS9hmzNeLAku
Enr5SJZIPzylj7DMQcT+plrK831kfY/Ilnel4Pyp2x5qiGC7IpfR8Axe+5ypxeXW
L+yp52FIyYU7VAT8bU7BaKLSPPmyFLu6849camyVU7up/zgsY3W6BwWcBkAd5IRy
h+SjDL+bj5nt+ApPz41w133KNbqh1kNv5iGdNw/t/8/M6HzebS1tnFwG+pcp3wOV
`protect END_PROTECTED
