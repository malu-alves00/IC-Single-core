`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TM7cxSXUVWZL7wttwy+xAn9X1jrWL5UwfIcLc5DsXYsznnWONI/mldGDidDLxzRK
q+QnoJSVv5bwDiC0SUbXzPgr+QV2Vddz72TooZQ3Mr4M5Q45+40OHEj0/gYDSmmE
soz9F+206E4o44zjBxG/SHeZruhAEuYsjwyAKnkyLvlpjmp+KdfMecZcXWqkANdi
BSWiQ03Bx+V87/Q0JGR/lG3GLGg/Ymxl5IcwKT/G0opqJxkh7j3ru3mTSLI9RwX/
jPK+b/3khF/1mRCk1aroFTZtsjyA6zdo+rSaZORnejgQRHt+A9F70rTcfVnjTCA7
UNMRkA/8WdjIhq74zM4R7Fjy7TYxMc1SPg8gHZPxpO1o9U1wLr7ACDaoMJJkLUtF
8dv5YL3VdSqWcTDyClWnu3XJ6utEewt1udlwLwa6cjTbKKQ70lOw/VN9Pgq/xttg
T18zUT9hORDQmoirg080j0QaZYtbBopqKun+LA1U59GyFkjXjSqzf7l2nwFLWUYY
kxSVn4GhCDMD3IYo2aaEwSqjF8vM5V1s2bP926kwGiToYDV1O0EQ4ayMVibumfXR
zBszc+UPZuvdzR1SUYw4HFLfDRw19U/CKl4mwfnB6TsP5TXFD/nZXmMozZzrXpB6
3bWzmmkO/zW4yLz3OQ/GYAXPZfIK2dEQjsT4UvBkHbEIu5g6E0iRIMX8wAGJWQPb
9aMD6B1DZ+gExHU7/oUapxWPj/RS8MWBiz30+rxDcBo7oE+TQqS0NoJJB4Imsckk
+dDLca6y8vcPsEZfMI5vwE2GxIMKLV2v6mQcMpASWJfmhM/Mw2Pe7aZBlV2/u+6R
gBvuYm5kn/dWYQADwRHH7LEf4vkYhtNfttHtXnCuEavRn09xXM2qMji5URTqKYJW
BWX4nxOCmUXKAOhA2lovSmYK+IamiMZ66PVuE4fxlCVOlqzaEh86eBefVvjkpcip
JogxxVoX32IMgtkE97zg/XhuG0BOSqYWtWMUzn97BtPiUyzDXN8RHxk4jT7KiMU7
Ft99Ax8O54e814d4p75UoHIPnikeyKhO4VYlOOGzohKB/jnXj3Adzo0Tg9RfwwCZ
FljuM095IYAjT9n/TtkJsrZJD+FZC2jRBuY7cp5eSHWTFyWmC3523P2J7CPLgaoV
bOkWw9UgfbWw8zsACgexwddwVY9E44CE8BBTl2Lk5F0CeBFZhzTKpIVQHyifNL/n
6Eo9fsKy8KCegKS9q/m2tFckQTKOKXEZQ6Nl/38q/vKksjh2dlhcISXpA5DrBGxJ
ycsu0au+h6vGJugiIkyZU/t7y1UmCyMIXhmPWuM7NSrSXWKotCb1DhZT8GNe2JgL
xVewBgr4iIQ3K4R8bxiQFtNHYA0iqe12BkAfZu2vKFkfW9oI9qtT7aANl6tttAui
MgEAq4sQqNqgC2i1L5A1lergdZJhqNJAu+5RN7pwafOHmz7bMoN48v9dzkqc+fBh
7RzX33o+D9qQWVKIoTZInQRrAMQQpdZ0wMo3A6O6RtgvCnTLIm/waV9vTYKUIfg3
oEyNnbmvA+ky4GE107467wloj8ZPqiBV98EWImycFNnyR9ehOPhf/RqTwJmPYbq7
PHx31dTdvMXa6lCtvX79Mmr21Vu4+i56hbCI8MT9/UvsX7EwlUBXwIKS9UfscQEb
A5sZCyzNh7BcUUxn6WyFURU8FteUCvGoYotTy6HpHbYxKUgSZSF3yVjs8w0UHUH2
jXMnYMOA8uXb9+KoGXVx4u7kCwpecFW279FeONPM0lbJxkWoshbI2n0yWLJW4oIx
Lw1ShNG32AJMucvqew6EUwwmsREJps9W0MG/ax61vv64H+TBPsBUkGEIAXsYuDtN
h6J5IbgmlrFuLYlisgMEluwdZf+PL+aGwETaj7X5MEmqPOHsxEQSSEH0QgOFvcR3
VeV77To0tjVlKDkvcMm/t2yPrfq4j/ZCzRUtrFD7m6mPXf6B74JrIu1HmyZwK62y
vmHAvOXBQFhghgrLLZHdOactDo7cAEksSVUiuOKYBaH9t0WcGjDdXZMkeTNITPbR
XOH42FKCk87qnFXITUw4aw==
`protect END_PROTECTED
