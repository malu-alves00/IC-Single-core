`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ANAZ8E9QeIvA0+8EGQCdiFK6dn/viRQFC4x9sqk3A2Lj/TCK9qt8P9qDgy4HMUxN
A7gINqHesa5XeAk43ZHaJRvMiKufnqCd2hy6qzzG6id8o/JI7HrQCZXz0r6g63Mp
SGA/h1loPwFSoYiDzZHDz3fn020hYjBufVyotD6yHVYUrHjpIT8tcyM9V3ITnRkw
tfGnttaMaVyr83fghl9ww/rPdsMGh7z9Go0W3vC9HyGnFw+VpCYwUSC23PJTBZ84
MS1nmKNZWebAYWFXUs9TZX9F3AIYNRe7OEsiHjUQdbVyLI/AQrwaAso7dm62dryk
v1BAkTs9j5UWFfuETnxTlwthuJHFX9RLLR9yXYhlGUiArzslBRy2dmoGHwFGox7c
6OAe71I+BfFlE41X+hRGmrSvYWnThILV9ye6jd72HC/zn6HbgB2wsBSEx/iZ3leo
Ot1GuppY5DMa4LBUnqXenscMBKo07j7MykPB5/BMMTWLC+YerE+OCYUnKPj6Q/iX
EdW6w62aojZQyATsPm2ofrFiO1kmPqgLxGvutow013K97a/VQSrXmJZRXcSZ5EK3
1YCWm980/dNGsZnmUCZzZg8RPAqTMgc/GQPInphMMdwNxIjUP8QceQLRWqSp22pV
odh11wWNVtD/2mnek0Vif7b30qNVom4xj7ejnuq4f15bsW/HZmLZmhACrOcG2v6N
vqEdYQ+J8f4WGuVF/aDcbBQ10nY53fG4rjmy+viuDPhHpzxm5c98cxFS4bbJpiN+
0msaQM4UqmMBMR84+NpISdpXdhtNDyqZKYKUYN8iaLMeRbNiKsU5b9dXN/flnnDb
spYamOIAkbkoq7+BnIscn2z5bA9jQU/LA3KrZnnhC0Zd7y4aYVQ01oYzFcaJBUOW
p1AVgV/d8Chi2z78UFTCoGiypffs8snMHMty54lQKrOJevLTax9Sv+e/9lsObzHL
G2Xf9B12O33y4QYTS/y6VFelAnTp4BaNgWuY3Nl8Yc+Issngd2TdHMyaVJrtSnsl
UDuoLZU8YJw9aYWh8aDpRt1qMuPdL+cywtAGJdeyeA94U53l2arw6SqUFefmojZe
DjXKcDzZHaoLvf3eV5CC/oM7ijhkU+qkQdZnOUylW2vAcPERg3wXmbVit6Dj/joQ
PE9xorlfqgUpDY0RNb1C8kNoo/t+wIedo6VwZaaY/vWJ3fpQtvL3twIiWwUKxf4Y
DG4f8D78npsnD74/msPHIMegyfnCCr2fKf1nggNmFDdKGDcYbxSrYvzAZmbhd0of
L3BxZt7MEDhbJhl3ZkVU2HsLScXZXpfYPBn9Hl7y6fC9sHm5rEsYkKCcKwu5GOOe
+KvJxSksQRlV1e3RVYymoXXEhMiLjl552Aatd+lVHljbcUsIAQlG+G/4RZIZTzFo
7fH+IhZMVIFpu3ywTBV5f7N4w3qLGf1p4W5ipJSTRDIMKciH7XZrm6imNx+uwA14
wOyKldxXr0YasKXqzmVRdEsJlcq+CELHrri32aDrmym6nlWj2XmWD2P0Z6ye2IN/
WvViOR8CpELzP2sCUjYENMx7AcswDmI/pT0W69eUJzoaOIWFsCGUQzAXUTMk8xCA
Z11hBmVlYCT2QmCr78bSzaND7tMqF1vHW11m6UwqWMky4t7EbstkjCevw2qpG7Te
QcG3venvX9hrKpWEbJKjpvtJlJVsK+85ruRJcz4ebYZ58T41BkJi6b+NybemrW3S
E70zcxi4LV5CvTwtTorDjQy5E+9j9EA4DFvCNULscteYJ6MZOk0Z4bWRhrLsAIkV
IJmInstN3WYQtBI3Lc6vXbgSP9h0Q48UqgGuuOZQkBtJDUu2EGEK6pGP+Zn5azQY
JJ/4wQQkBuKSjxM6TxDloJhXtdVjMrDv69kUBxHsFNUlhHrdQAHKRqE1FH2pW4oH
+e8Pa3Y6CTOoQPDy+PVxFHGM0OMG4M3B3bF2nGMETrzUAry/8qpRu+AUcJGqbpVP
UncPYTWn0wJeQ9FEztA4o20t0FSntpiuw72v6RBpgw2JXBxmPNwvNPLploj0kty7
ApehBeygkXzAUWfmaUbFo+ImTddbaH16gNr/O/Vl44LioMoI3fTzU/QD/vY2PGbH
wMMvyw6kBpmmlZK3GmS/0n66IxQ0Vr67qn99SFCQYU2eulpOnlL0TRtoswP8NMR4
a1SQnLy/Nd/GrwtXsdcoZbuphO9xMHuCgqgOrWwaGT+5KdZsvWGacIKaoqVSItwD
Apf9pWl2XJfIGG1c7YjEEqwtUWDGCttvHMIa/GKAqWOdt6c+T9SSWajOI4k4YisY
ccacKQcUwRpVuYZNZBNnYZ9l5nMveWWi/0MDZ2iHzATDbAcPKr6c7SAPeA4BlKgb
kz1jVpdFsbQLzXXXOSUXfAh8dWHf43D2K+2mEXD3/GgcctlQemXUF2iottC5VgCn
Kn1pwY0hTBuiZriJ4yweSW3Yx/0MTEFjwdgpTsz3mU/OgmKQ11rVm3yGhLM+cL1I
aWS6HhQW2ASjUNsvKbFj5flnKk25iRzmNcBHsnU4wEP6ISkIuFmI6m8MIG4b8bHk
MEbeDQzCttiLjXfk4PWL1bkTDNFLAcOepyllSDzOdswoZGuoY1WScDLMyAymJTY9
0AjPWOJ/EHxiAnUiqPp8abfDSRHZGLQbUFHM6DEaeC9gh1j0ZA0j53XJVQWJeCCt
CKBfrG5LARpqqZ+Ok5wPdMJW0vVvewJQ+dSh64Bze6ngmINjScnUysR9hvrhOqQA
PxWbP1HdQjFR+SNilmLRvmKZpxQu6jhcclxE7bPoKtq/Q8caaw+0D6H5xtXRHVGk
VkoXf9byxewrWAJNUPKm/Ef8jkf+/LXa9hNotoPqtqskwjOHrDOX7Qw56nQsTips
M2gMsfmyAWPD1Lq3J+d5jEoMsVdU73JUe6bJoJ4YpMgqO08p1xOrNUzM6pKrlm3D
OVuwIv61/DW3mOcIbhbYUqWAwba6ww0DcbWXf6M8B5BuPLsFZIiOuUU8bcGWMU3d
B5GSPkbuE7iYTD8Pwgr8pB1gSxEwOvUMdWTuEAkwX8MfFm/igqezmRcnVclzGYHp
8VGN5ic4EDQNppMkAKC54gCP50pnEDjinBvLg0l9dGHoFrrUpm96esFdDN2SqZCr
0Vl0iAsh1siGVTGp3p+DCY69sCFpZzFZ9eF4vhtgbA9W77IFzmnNGKCsbUQ1B0xR
19I6ESmfhH7Gp0z1WqtXCtUiAX04ovrS3u2yBUiCR5yjcsAJ/IgBebDag2ECGqaA
nyUSUoTHA/EkpMubFaJnLyCNzVZ2V8fvM2+8/mfo3Z5MvpYXy5ZjqQHheNPF1Dod
dgc8YEl8BSWwrgBnSTN0eTxfrHG6AJ0Ye5GWx0GyeHe4Saqws7PyKxyPIyzob9ZT
RgTZKXEeo6TUdpOZxLdm5YwGrc4RkCIZaX9ugDmjxEYAAwVDJFX4O6uj6l2CoEyF
d32umEPSkUjvkG7yMRuHem5s5MAAGf0CLD1JHiFjqLllEG/l4s8B5lE5olxjCwPG
gexqZdTwqxWt+RGWKbw3Rv1j66zxDJQPjyNyQfSE/BeBDDWc69OKhWrqTimFxi3K
031v75TmOnq5CpXbEU+t9d7UtKxVvEvO3fvstld69+Uwx9fk7nXC8d0aWvliI1w/
PZN5DJJOLY6ilZTAmXBUmaQGNSJrEt4FABOsDRwDPEBNGfS8thJ9tpyZOiR1e0HW
xcdq9LTW3kYaxcwTOoSRSiRCAGx6o7uKK6GCyblO4WvDxXv9e8XWB1fRYqJv/cOT
JjYu7EGfdKTJ2Eg4bKeTNgLe+l7ORmWXJ7T+eqJ+3cr3Tl2n4ydszqKgBpmhqf+n
JTEb9PtbS/WJ1TukaVQ77KIaNuuN/l/hWNuolNB8qN1hj7FmpYSv/nBCsmd02lWT
aDOsJgEuhFbrFZq2iFL1/7Pik2fBvfAu8q+X4fb6Vb1Sqo3l7boolqtxRIqdGGGi
kNLdLgPqvySx7eqwR6eplq5JfdojK+bg5eh1voJNiyx4yIkWw+Y2lVJWRj4NY+DZ
FEymQ31yvzArwoEZUUKcPMCQDlfZBthZUqeAahDpkK7af2Vky1rCLSsiVwqPLheX
rLF8aRUqGZkTFBQ3KFUt1oZjAsOQ9AQo5JnJK/a2FygxsmIC4EdYIEjltjryD77Q
VxgSH+UP78Zqyy9Zj6RlQ+UJD8OY8VramX95ot3VmgC12Bhj+9mLq/hKsuDQbuc9
GkNO9ek4sGOlhUX6DI0KTHSXPaQGSPz0mMJ4So31coqTQI2c+R+A3oKaS11iyZpT
tZ7OlQtB9YnUxtwJ9EXCj7CdrPIHtExFLDzzngENmkN/A8L17vC2pUgyCAsuxu/s
DOp1Tv5rVBO2DaYowHhnS8JzaCinCEpFnqF+A4QlfqJpz763l/gZ5BIqfh4amEu7
S1GQQRdLbxB2/waMDVELlmsSZlt9wdrAvWsYWqYlPao=
`protect END_PROTECTED
