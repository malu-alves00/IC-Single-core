`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VHd+9ByeAta+Z7LdDC3ahCKSyyKW8e34BdkNbbEwd46zcGWkRFaDQIovMWZSN3Sf
/JL7Suyk9ioCwLXM/JwpxLN4WBZUXNY+htViPEZ66l+8o1wL/5V8DyZB/MmOtMk0
hjCn0yFuXNIWupoFsvPXBsd0RrIpCJz6XswFdmR357/5XEyE8QTWOVXRVxisQTnl
lU/p5lAcQhy1oaLDPe9U+LLpywxyZ/G6nAyaPm9UNe20XjGHJNbTAHROPTP7rfHN
piW/qfSCZSgTMWW2x0xwwKuSo8tYZqmPlfPkWo+30r4MQYbqpbcbcdnaaTvJvApn
efIcPCCWJYjr5VAwyNHF7H6gQs6MYuTFXHdDwxv3bCSBi2fK8PtbyFxT/VNPzwoO
UKoOiuDT3Q+gtvVbQp0+jacgPlikc29FOkgDW0rkC7fS5E8UY+IphxIVwi7YAuQN
NleeqONAqkBU94ElVpHRhqSsM6Zt2DjO7akFX59NApP4iFd+LhMR73tu2XtPrGB0
LmWBPU7jF3nFZGyEvmW7dPAtmOOh9Rv2aN9hgmlvvOQAIh572vobBV8noJ0MEtOZ
GW/DjM5PDbVWLB9cT+6X8W+xy86Lgy4e4kT0GEw/cbPxIV8C8akmsHwSwGi+neqJ
950B9wtzfcTxJfkY37GF6GOKmytvg8vIzoqvVJaZWCoP+zBBk8XnD7ozhLoLiL6X
f9zVYqvMfXgTd3DnZqWKz99zNOTqJgFx+Wt81qcya/rPKy2z8Eq4/dVidlC0jCIe
aHnpE88fjOmxvE8Fpuj//dWWU/Y0pu7GwYB5jN0SGIKotgaaxkH0/IljOsO0hf3j
eXOVN2glJWNsHxOf0/BeTNYXZecgHjzjsgdZvEK/npPsjoUqYmF5ZYmbix4Smt5t
tSxxXcmt0XELAtkBnXzpgOVgICTLvko3y0Whj4tqk5IS8XBNjxZP+8MXPm7qiw4V
1JamrWdmg7hipYuc7Z+sToGIf2AbWCHMb3buwNFEVTn3QwI8Dj1yOw40BdsXplgE
Pved11wrlRRpC8k3o2ExDIGo5DAo8uBmJ6gvhMuZiY54SiRdrZax65c7akEYh9dn
MYH/rW+/FtFirny3nteChwU5P+0nW3SM8WsykAnOSTjQfhV6ckMRhN7OnNg9F06B
doUP2JTS8npPsY7O5Oe9ohiyGjm+/evQZeko5PzkeKxVBeLrkLbZvIi5W+WaxgZf
u0uSlSQHJLV3LATGnD6z8N1Vvjkii4ArrLI/S8E7CqkFBuSm2ssiwn5/BbvTZ893
9ZaCPiPkUBN9mvwpgQlMTA==
`protect END_PROTECTED
