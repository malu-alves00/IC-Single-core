`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
P/JVY6mE5tB78g48bVdqtw/T9DxOdr3QNUD0lm7R/sXrnRksBleVy34zIfZ4B/eS
2jRoMzEoXLylPjrv8k08bZ/eOMevX5oogpPV4Fl1j68WibeAkUBpSaWwQj5A8cGS
csIWj4nuOs10UXss+7BaaPkvyaE4SlL9+mq2oh35NVeauL8hW1RsjPKaq8dWgiai
Yb9pe04sSK9ipf7dJ9dlMACVK0mh59rqrT51OFpNHAFyuhMTFSUhl3tidFWigbr2
5RchEMWU5hIei2GPRkdXDfzkVvd9Ob/TsvuBDqYT2aXuUcjlX3N4kQgSJSbj5cif
wLOIbB0sC9BrH4gyTg1JyYcysOyLh8R8e2gIE5vuQRTo6wpN5nmcQnE5z7QjddwF
zPmk1OYPoaajfsatPPEcQcwdIfJWELm2AZ4DdmAIkUyfCxFDY26p1KqTZMs330my
EkrE1Hz/zj3wKAv4R74gpJjqB30nakjFcIMmYuxO2t3ais7frEAvRkK0O+rdSHXr
S1vFRJdfLvkH4QoKkOsRummkik7MHyY1d33rCtG6+4pO4BTFQGj5TVl5GintfEf+
ZVtBMXuRK9LIh4sDYx/Wzw==
`protect END_PROTECTED
