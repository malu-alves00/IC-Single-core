`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
s7LEUepZbkI3WU1A/veAS61PdHwagJxb3SrtMYAqnRhNJ2nhhPUX0XwqDCE/M81e
uFoOAlt2JZQ/pveLZ2BdhLgzBn76Gk0w81pprjqUbdkFM8r3Bt8w4+eXDfxIz8YM
HMtL3aww1w4svoxQZ5xLJHrhKx/C3o36XGevODcLDx7u1qXYm2EaY8YwYf6fk/Hp
YzPtHruLNiEHmAgSomRMBBsLTITC+rACdJkFlJC/W9xV1qEY71qMWbM8s5/CKc5d
2badzAphnvRJU0Ra8sZT3H4hpC58irMWNyfLlYcIJOi1rb5OxDkbYXewBCfVyC5+
Q8IU+P0bdwsf7cYuGB8Hgqd8eIGJMBwjDOvBDsllh91dFrCnBVWyY89r9pYc+UVE
W/qDTw41qs6/63GNWSue//1LyXtLTxrS+/WU07d6eH2eX4C71Ze+H9u7jaRclqcG
7/QEVIDJvxiu9TfBWoCqvF3f6hUxU2dFWTb4BGXZLH3gCsNRjVvW1Bq0MzHbFwU4
tS2pKFD62oa0ucPthFjrZfBRS6IuNbR6nfBcTSDZARth2zznMHwBYXkgugm3adRm
X04RYBSK7Dhg7rvAH/+BzGCxiG8y+sV1UmLEyJuyBlRsyFQC+4oncwCRYA7E+qoy
2XB3Ol2uyPIpbcz2Nk861I5jhsVHu8Wkx2Qpf7dORnXtGzSyKlD6gJ2oaIymFEXY
472ochihZK+kcBCH01/ua+x7VHSrfDVvk+Ac3o2CSBKEK34um47Vl3P+3xTXB+41
VhOKv4rreY98Holu+jOsF4Mtu9XQmlbubY/brbNEmSrR46+PtL7pm21wXbRjiidd
V6UTqFPJtctMRz8q0I428wQwywG1J0RTlRUuiy7BdNufzTPkmjDhe57kFAntc5AW
rbhwhhznx2+y2HbRRdV8eT0xzX2tlPv1TFzPwgWQIWVwf1S27uFMN67nUR/5JMV3
bnpGIMGpEeqBFzUrT9GY8uNN32Cdz398yBWIcsFH6FNLaV7p+LVvHNOO/JYOzGtk
IsqycgxRTa6hhht+CXbpWpwJKxPUx7Hm8v0o5cPK/PjMZOQzN9/xfGofKdoFLqtr
jsuNj4pSD3mkLv3/cxj9HOcwEP3pwwkYmqRKTRqiHPruzccneHzeXBfO1tIkSQx8
88NtUCZ0Rh3cLL5Id72nfRCHY4LwLjHRuf+t6FFt4Bg09kr8zenDQEUFDyYk+bzD
pYa4Ty8ZkqevIuw6wb///I06XS5wvbtp3+rbDYqA2mbdTD2vrkQt78ABZbxIVqMi
ZI4Cu5ZRLw1LKWaS5sYwhOqnIaAJZxtIt6R8+c/sHO14/3V/jmUslJvW/NK1oTJy
MMB2L7gHw1hdOGtQNjdNfKaftlt7zaGcJYnWuwk5OhhfpG3lrXQuGlk7hdcXBIff
rYAdQm2EXwkJtYn/YRmZNvIMjlPiMgZ7RRCOpfE5dI3tLvh1qxx6jjQSuZFiLEOC
JFegV+3mfh4UzQG3N3ysrWSuoiMQ2h/GT0M2QZDTCclJW1nwtzWdmpkbm4eavvOo
rXwzqeJfGWcfgZVnfaYMI8DKkaZOH3uDIdqQRXEFlA8dIsqrxiWzDv2krt1K34mm
kzpBpcZQILAM1mJOmYLlFAkM+/9LIJC5EcF2CswrfOlY7dGeQE+bdi8iE9PkLpG2
g0x2hibmV0nThMvIkKF5qdf9rvuPi4VaJy1uonofqRVFwhV/8KLaua55La7AakVn
OGCULbZSugbNh2q0atoLFQ==
`protect END_PROTECTED
