`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
x2Tus5dudb1XbhXelX9X6Xup+aulWerPsqaQpxTvFkmikaQnmfvG2eGiRBBJA9ma
WAWhocs0fcGy5SsvKTHsWLvwE1BvcQZIra3RDxp+ZfqZSVsJH4tfbNvLkwaWZHBm
JyUnq3NflHw+N4m4/V0viqTia5IBVwfpq8kantYj2rWKrqyqFvPRmcBwbuVyYDOq
WL7kUa3YsEXp6qrPnZaTVGrSlBBlChXQV5NUdCHPpSNYePU7Nsje8FWS3yRx5KSa
hxVzCC1bkZMKdkcP+hFdT5u9fvRumgU9qSO1p6KDkC9wIAlFrrdk/SlwQ43S425m
Icxj5Bg0bcHkogyUVjPpJ/dBCpFhgoV14ZLSXArYYcDiYjof4Sct7tFLHqOT4SJY
M0q4cFmgUZKNN4pZZYAayZ1Mcd1nTaT2X/ALqE/b8p8JuQLf7K/ziBm9tHhIlTMD
iUb0iE2O2vzYr/nVE0lhy+PnPv8jeqnpb/IUg2YOGsabuPX/lqr3kTL1tTkpPj+G
EoFz5sbTv67SOpy3MpGOQKTGmrdweFn2OUnEfFfyqpodR9lbZgqNOlerZ9/Ucyjo
g7gGg9q8bmFj3jjoQ61CUrJGyORE3zt8ETxrZ5li7OcbzV25qFwYqQHEhn+j7Ywg
P84F9pweb0ns2x9AWsHpSyZkqeg817OKWDyXN4hWVkuH5sHrwyp7nPK2xWPZ7jKo
opba1Hh+jPoxbWBGFVUiQgJn63PWnZPBdl1/RIN+qyA+Rq8uy7hA/wBf0vQ7hSsn
OXZbKAYD1QI+rc+0e7DCbECzWL4BNeL6l1kpl7ud+eLZboUBsepey6FVcAc9FHMP
REaZkD6dBgliTfRzgDZR06xVA5GVEodnQ15l6KjXEPrpx+XwcFCaM+KuOmlqW5U0
V+ssGGKTHn9FjTJCnZrwa0jCAZsvwC0DvN3310yjcbw92QAaQCRhKQjij+Z03SHi
cgv2t8A4qIQnQwFRhUdsu/0/mJ6gh4yNqJC329W8ujjAGMoiXGVnxZXiTPqy5tfD
5NvKlf6FMSHUpKPvRU2Sqwa/fhtq25GnIV3qb+xdj8a+Wrf/vNsPzBwxoWwsQJgu
EZ2fzEYq9Eot2I0Yfw0oGh//sFqAfmzHuSw5+bKeLyEkOBp0idzd3B7Oe9N8Mo5O
t029xpUwbZP/VJvtyhi/HoR5k2AmA4TPlMUXgm+K/5ChUMCVegUB5TjrOtUD+fQM
Zv0pZFgYa0N3pftjlQXBOBh1srBvvfPVdpEk2YtERwx74ZJrFLDlm6aAlpG/xBXk
mOnpw0ZkrtNQBdxYU7BclNEuD7btSK0DC9RUMq8huBycMUXV4quNJZYEhv/iN0o2
9GXeCm96SCyLJMqt2GsMNSpvfIQW4w+ObrEukL8Lgc8G+7YaIGQCElji9upX1mpG
/xgtZGv0Zp23xVqodxd+vmqhhKLahIAHrdmdiO3MIwwAu+EXweGEYfaxFf9IRskd
Uzg49buVkEudQhtpUPDzRvxAnfy+DEaEvCpY4vE37eBNKmqlcgW1h2MGMvIMx2br
jOOCF++zF7RlHeGRwqZJt5+yi79sXYQ7vB0+A4CwsMInLWm6QBtWAJhqJa3Pfb5B
VPvADk8Yby9/Sm3EE6oA8Un3r/p9cVtE0ArEmlGXP+WZqAF9VpO8LOX/LLa0Lu9R
LeOEHJPrA3IPSfQNHiQa3Y2BOb46dAFwegHfTeQFHFmuHu6hILsqsz2C9iOpUM46
FRUwLWlsg3UA6bcPSIhjKDg7936U5fH9Ao0uYEU3SFE6Ra59jcgvUZXs97RJio0x
1QcZQJ9eiRvhNq5baNvNA7H6UlDyruZFUOwh9texg+2epziDZr11NjvCan0Jj9OQ
3MFqbJj/pZJIDvvfZAiTbpph72UGlNExan23pGjbzxmlguGy4lgcs5UntqNXXbGK
BPSAdsDpfVIGr2DJCLWkELacZ75oArZaKxP69J3mQUmF7pI42kq2pYvCOQI5nrWJ
LlAcD4jWzPOBbxnPufpsmuvjpcZHmHszwkZTnpltkHxn+KlbLzxUG1dta9WYlMp+
ce9hK9yV7CjEdcD7Wgq0gPdLZMH9ULCmT+JX4I2gi4T1CVE2talXnK9Y5Hsb/DNR
5IoXepiwYXdch5Tlz92auuKVL/44Al0t0hcPfjXd4sr1b24++G7tJlZEjXTB9cTa
4AuXy8mPpkaA4F23b0gUCOFwXjz4mKoM3SMmSCFCRT07B6LeMmmfc0DrPPpdo7FX
fVTemDigmaHy3eo/phuwbehmR8xZcNU0tshMuO8LAriPHexRIa92jAd2/eZDRY26
Mte3d4gH+5EoVdB4ASv7STzirnN+OzqcTRBkN1fip1vcNYAtTi1WPM+b6cy/9rzE
rbbP1i7wbdb/SmQtOVX7VfIQlbou011Ei9kgk20tDP3/ClyQljd8d3jmmod8wt4P
xbuSfzRFMLkQ1nyhrEjDWSoi91MdQGqdLdvgRa/UANE7gi09/4f7q1kuQFvHgysP
aGY/9ZRXLfVcPYWvoiUYBdFOB4/jiQNpYnEEtigh4uspoNF2DVVRSks4lmbSCmsR
JV0KPn309yRTiXqN1FmeqfIAV6e93j7ESb1unaTgdG3WodHt41hoczEw4BfExVI4
XDoJOb1FUDDgQX+2eAq0Vuhd2R2pwaM0eA2hY74aGnBrmqn+a8xqO7h5vssqOuhd
bqciTXvrT37QLhFIT/XN/Gh35Kyz8FFyayzBXI5ygbXgOR/bFsUjODRGeg6bulw1
3jhmDHh1njV1VH+yQh/R1yVnrRgNRRrRyGDfn5ucVp9yMt+Lh+qx1/mqdJTtxFs9
RVoZTI5OGoyW+2OcVdXnzmr3yZMzlUxCRIhXHk2JJrmsT7iW8E5kwQ+oWU0WgWXi
yG8hLrDOztZ5VBGEo5CSgv60vvqk0sm8jWNmXFNmUaNaZPQrfM8X2ojCMjrpzL+V
JUQ9JjNpDh+w3ITCJ7fMP4pO1mSDUrB9J2z4MjqUozeNN3KLHNRPCVFM/gjszPvl
M60NHhGxf24rbUYLSfrkrUmrDb0+AMebNu4jtWqzt/zGZaF3z64YpJHWp1pjwm0P
F5Q3jvoFIRE1ySjZxMhlORfRhqNrYc5GbxQDqd0RtppQk/ia71dVO04+abnaC0YS
fON1t5sqvfzbbIdrhoBmzQfqL3Pv/iaeRP0WnFlknbE8C/fE9npa8jIIlKH7mbWK
g1NArD1Aqq5iQ1Hq9q0OkJEmJUwo/LCU5Bm1PhndCFHa2dE+R0VFZCWvhoRq4jQk
Lf+N3J8KEqQimJBGZyrfoUO3hPEbrCNkG+IGwYCQbgdCfPJXILTLf/qsNHLxlr/d
Ri4P9eTPURyZSzKbGZgHr7px9dThKle5qW1my+gNblQ7yLVslCotyi6TNIfBtsfP
VHgj/Brzjc59HtibLQJy/Jb/va0cxjdW+DiLTb58APkQ0SaFcsoe4vxkvOdegO7J
ULoP8yWq0cXA3k5km+nXAWEZOK60XX+zghp1bonFAeCqeF41L5INwknlxGmh98f4
smmP3Vh//h06bzTFSY2k9XNwmwpPT6er8LRG3YmMNA/sd/YOa3MRYmEE1Qr11Gbh
X+yHVySgXfFKUR43FJES0kpq4rYhcTC9h2N8ZNpWkGaazFP8qNMi/ntnM3KIbl6Q
10CebD11JFoGlrxJtIHPknh0nqpGGKxBVZeKehjLCAX66McFGRTuGuDVjF2Ns5pE
2TQN+uU4MYJlFZRwisi0ZqIYb4IcU717vhOO9hpXi1OUhhc/FNcCBOOmzKxHtifp
K8mKf2xvh3SkQGrUs5N9E9wKvG2ONK6tVL3wDdVZ0eMrfTqNjAHcOSHgTT5GZU+I
NgfOn0lSOCP4cW5JloWtk+yLqElIK16I9WRsq+MGXbtZTRlyGl8RZ8wAl3Mme1DQ
MeiyxR9RZ2VKwhkpq/cZzPb9ITe6Bx2PAZWJm4LtbQVFdAckLcqytvZj/Yn+tcgW
z4ds0Sv59dYbPgjmij9dJ5M1q31QLLSSKeqAZlm/mH5rkBVDT/DTSYdQDuyKvybB
uWceWEieaL/ZyHQpBWF4LS8XM8O8kzARP5GCkvGDT7lUmkME7Y68Q3N/8nUxt4Gh
KAJ21PKUEP4/2BAWVgS338uPbJD76YDgBsbhT9WbiSHjXuLfUWpAXXm/PZ+lLsfQ
Lo4Iu2j3BA8+iU1/Xq4YQqJSjKurvuPYKe+A5gjGHRRtO6ISFblLHTgAxFiFNaVT
OYrsA10K4FEJ6D6/kF/2CfvoWvJUT93hPkWh6iK6Sq5+hbNHW79h+US2ORqskQ0f
xLr0nbp8XmjfKicQ4aJ232CCSogOj5Ps6Iu9U+Ji7HWM1BvFE9Tb1Xg58rtdZ5w8
zmDb+9NJd9NcioK5RCoe+ymWPWIEEebOynkbX5Y3LvRcyGBBWs+CzqCaQ2krP3/C
nhtq8hhWn0bzc4w92SetxTkAEH7dsRDXm7IGecdqlNaNsBuNVJbn0Kz8GcTQsz1s
mdy7sguTs3p31aNLOOzwqW3yKGlHTM+lCC4Ux7VAVyVA7loHq+svnoLUhB3LHGH5
jlOtLFrEIEC9E5U9wWbR0ieVeNQhbEwgWnrT0We1UEIyd9wyn/5i5kF0TlwH+arA
eP7okwhzLUKY5DRL5G3iuYgJc3kh72yEsSapoNWWpYtZL1zVe8kM0aEFmPgX8og9
Q65Gn1ecsTOJ3fF1bVR7ciOPhrtQfEu2Bce6UW3MyjPDKt5HCPvl7VbSPgPirSxp
slsllNMQTmd993X8RyQgvnB2s+CigXSLkZAZq971C7Cu2e4PpBy0P3rJsA5P+EKu
i8iWl/Rdkg1xC7VzbLZuQblzOZ2ES99pNyuHqUxIUa4CvkW5OuKJ85K3xhiGWOdY
7qEun80gBj+T1Ucvvqwjg7+dhfRR9FUkagyZU5DLkn2D7oGuEi7SvgYTrus9lHB3
hc4ddEL00mhiK8XTEkQD+BYlw1RPmBPhD2/8ZE7G96iUM+lurUmWaTV7f2pXJuQk
JSVRnE1NSK+Ymo+keaE+jHGKLxD8VBMYbPzTPetH6BtmI0xEtCY1lDix7CUAMrTe
D+4Zm19yhVuZ2Q9h4Vqy1KfxD/i1gbMNCDTBX05Wcmg/BF/GRcE9lqoswW6P83j0
XmzIq8LTo/n/LcsVmcNsKPXbjPzQdjCVDihOAaweSCgasVnrn4N49PimTIWP3fJm
WD6VUxaueKfij/t+N6Vz1RchKrMus25gHxCYPQceYUPjP1A97VFyvLgWzc9YCmq5
WwCFv5F8w8OGjQmqwBgJpMxqt3SH4yToFqeBPsZThWqw3N7bMw7XNEELtlDVx8vu
lYPKeyYl5vF0lTihtBZoVWeHu78z+QD0tVr5PugQuICQiacEhE0Zu2UTZL9rTE6k
2tWab6bxXOJxIONtNS3JOzpt3oPlH0WMP5oT+wGPGp7/2FVU5UjIaOJkZ+GzMK06
dx2TcvhupyKxYdDsuwPqCQ==
`protect END_PROTECTED
