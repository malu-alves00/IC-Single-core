`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
r7D4/RLaI8Nn9M0VDriXDzZivIZGGlv4ZQTjJOkjMs9YZO9EDPuiin3bvjwUcVrP
4Rzxt5j1ePg2uzE1UE4vvOjiJm9RZuzX6jR8OLtTrw3/FZL7c+mUL+LzwXd0a6bc
SiL8q9bfcQD3xczY8yMH/HPjZzEF3lF5kY11BGTlZRAtEkM5rN37UGu08XVavv+8
ioeSY53eW9lNo7X1loqttc7iwBy5nSG5M53HA513d300k9M1N2s8ZGLpQwX5bQ7K
iL0mdFe9HZUrfoXTIDmKHF9z8drpYs/b9W+FvbkfDjYdImwD0P6GYmXsXgY/5Tg2
E7mey8WpGXrNV5qJX8Pr5JPXyeSkYJTyG4vI933a1JJUFctR3gOrlu4SOUhNMMbl
CJaDUHaDf1eTLAmYZsHqiulB3/WLQcvSOEPDz9WvkYyaFAx+LNAFQCrKjuBZi/0T
Aau56a5WqhFSaCQCB2P5EhT4WdVytvPf3PZPHcSTd+Mfhdn4eQfrxyL9pMEFzQa1
U0eHJDrC7dKLarLM1bRPD8qbokLVYZFg0rkjMAyOnYgzmOLLInaFjhaZhsyBSiHh
3RvFJKQwkiMY6WhY4NfVGA1uWx+ZPrgTwd3wib+s6Gpr/BbOEEpJ8ZdhVTgJwkL3
dDRlO2UNhNhZnIZt5Oj4b7ijzgPHtHIlUYWUPgRK6GSZNFKFz/Sjc5VJL9AydAzK
`protect END_PROTECTED
