`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IZEy5NrHKxJ6F7+dAe25mc7yirUeQxgclYe56V3Vzmx448EFSlFYvC3jpXaqfCVg
2+JHRqY9k7IVDg9JnHodBP50MaPtmtEdt8hmtWOLfef/UrKox4lgaKwaHaLVS2VU
3GFrz68HY6YDPzGGepw2+VBcev+kxxYxVAWAMLCP3sPjx6wvWHUsSVwY2RT29NxD
RJV78git0zc/8ivhO4wpP7C+ya77UtsqNXaW4a5gSI0YmCG4bnAuf09ni/f2ihhx
3WKxzA+ieaoToSs+h/qGdrxg50ErAhaZ2nRPyNkH8/n/e0QMjtELiENSiStEaf7g
IDlmYx1sIT9zehhoUx/QJKkDcnzUzct7pXF4PeR7iTwPViee9tmSayBpgCf2hZTF
SaSnit05DW/T1WSJUxMhbxzCWoJHezpmXNEMqMPiWC2TJnfCRSvUhNq6SjW9CzG8
jQnElno9P0lZEvz7aGnQC29JloHT7dC65em+E8dsDYvp5AFyGQKgmFhLi4D7oyA8
cTrlYk0b+VcxVYf3kDH6fNy7a8aq/te35d2OMpn2UEnHAfaYHmHenvDbjaBGxLTl
tzU0mx6Tz+OjuW23Ac21KkVfYZ8SWILennnmritOkd1mJlG4EDOhraNe2I792vRW
FltJhc5LneFEmeFoAyXlwEnetGeXgt1ZnSIsEal5ctx5YvG5sahO4n7XwbVh47UV
RAhidCVsW3+0Xgo3H5LGW2uKMOrTKPX7TYoCeMjH9mNWwJFwzVl8c5qSrPeB47Gt
oiSGq6YjpI1kUEIiKZXkuShYU6l7ny9lFL+1BoF4O1OQ03pmiD9LxYUpy8TxUool
K5FbWbKrE7/wpWd46PMIDtPxOcvtXVGz+12cXiPTfT8UBKzzvSdC8FkpfI4RG127
XBWPqOPWQebIqVf94y+i0hjJqEeaguIjNHtgTPsob1nAW8oZoFLWclu+AQjf6KPJ
c29Z8DRQWqQPKsohpIzphCy9bL1WHsYaPZmLElU9RhujU/9C+Fnjonx/k2D1IZqS
cioIRPl4X6LekB4Q5dljxFuI6giuSaWP3CruYWik99Ag9x0phEOtU9OFbhUGUB4F
QpeUoc28Oq/cLDxA5Z7AfOfmrP2AkWhp0LAW41rsTRtW3xRghwpDoE+jeLJ6d+mm
GOrZaR08kkoSBpbAWpjq9SYLav2UtjYp9McTobV7T+0R4ZN3z7to9NXYJbwdr1mX
EURLMvX9mRBfkfEx12dh/B3G/gXbPLvTkKB8aWbYbrSZoDaBtGLOdZ7R+8Qltmgw
ODJZOCsodoE/hcouTTnXsDcyeULSlAWrQIs98reVzyAU3vFudouRXyagjHttXJdW
Nd344QeeEFkFf+t70hji7mb6MsO4gQ/8QZUa9ICuPqkzhbE56gkGHm4fxiuKZliO
LI/5VmjKaKTQomhKq1Zo90T/Ic9uB+ZcvQ5evlNSWzAUfZKHiXSEItL1XQJdhvhe
kn9rlhtQgirMWjgImkoLcpILFuGJScqEvN01ehI4ZNlenGBi4ptl2Yg+LKkKFdvl
QBxSSeLx2msJcfhuqeRmV/p4e3yI6c/ILlNubIm7dFYa+z/qU6aRUpYYVV5lmYVG
FWZDRKUijnKrk37z4wEIIKE3gWmEYykg0p0qK5zg8Jv3bXxkzxnZS2eaOHNiJrcv
jvz/lFa8KhxagByaqUInvTlKtiaUKWtKvTn9fEhVluLuBkoKWKJxz04HNROJPVa3
`protect END_PROTECTED
