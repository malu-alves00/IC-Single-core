`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
p18s0GeKISv+kI9jWpwsMI64xFOwrH1XaBlv212dx6T55HKQXYBZ4I35YJCk+stb
poLQkXj+RH6GVhnb7edJcpCWzi5xCFBoDavsP3kuueltCatH2JJD+Fj0dVZ7JRnM
a31gz2nLr7O9se4yZKawp62p1Wt2qJLTcHxu3JNsSnGZ3ojrBIbnkwqt/TmbTMfl
WBOUcl+NAZba4Dl0ihMg4K4SKcAhEB/gbIcHnzfsRK3rlneGO7SicR4LCZnXfkDw
0/iu8jxDsfz/NY32KJBX8qKctOlShDP2pPXMkyZIjxULWOShqG78UCSGRTaSaZ0e
rDLs5nYmmchxiSQLQcv9H/VSEzHj3IInuGt4ibsZbtAOLtEHHuNrVdjMH1Ch3PMY
Kk5x02WW9BTpk66ct3LvSoPtS0ThJf2I3jp7tWYGtwQS6J1pdiKu43qQFaOxrOSr
/spj8J19N7MU2u7QqoFtl8W/V2hym71Ee67tiXZKiyDxzRCjNcRd/5EjqJNOBUb0
11ABNjJHag8hvYLQKifZvLYq95U3LVEE6DGc/IC98O6KKDiajuR6v8NMHeuVgCDn
0HxPoGpJLF2gqj9NAbXJ69VceIlAVvdJCL9LkSypFkg=
`protect END_PROTECTED
