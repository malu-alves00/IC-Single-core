`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9CoKPImRVji1TwidLaeAmonyZqbXmLcY3W8mk5uzHTgluY+9/mT1sCkfSAGt0uBw
bV43PWP8SY1907Cem+P/6zvH2uYJi/+P7fXwkR8IxPhNAwa9962hCbB6W4vBWFkF
T9CEoeZKBpvJGSx2daWOuXqzKbYVYNMGmUAstjv483JiU35pYNDcmav/Ry5ZZ5Uu
wDkHJnNJzb6De7MGAzImd0bZeD8o4jZJW3unWZHUocPjy1WBiHMbcdBfG8HZunF8
+v+PESgAJX6iDR7YgJCR1Df9m5zpRJhpeT52So/hjhvqbu9UBfgaTlGY7+dytjjG
RJ+5cxc5bsJ7l2S6foJ9Ym6JOV/873milPFi0XwBhc27EYVMt9D+W7Z16oc5IuCJ
VBXm20ZNDPDoIw9tBpOX+0q8jEPfMrDp8rnEvrXTGwwo4YOh2+JqLtd/hIXK5wWv
IvE+RtZyWr++/lF3z105eh2pSmGvkKv3It/Vn7vD+3pYo977uWm2rGNWWF2zcNRR
fryvPk5k1nlMBemZjVMDl0XSJCxkd7sZ/DfxcOCUHGKCcdT8u+LgcdAxlzxxYSL6
uG0EoXvz5hUtJvIUkR3vKg==
`protect END_PROTECTED
