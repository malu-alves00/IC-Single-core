`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8qRKUNJNCtfiFETJvrQyzGJE9hRQIaPJARWd7mjHeCfmS5LkgEw+v7sCKHhFiYH6
Gb/52tHobtFz3Xcqr0FZCOCKi8HxEB1M3AcpVXPSlXQqdrTEqNOGJWpGVJohYUmd
nPDytBmPkftGCE1H3c5d8K1b4jO6aMrzDwNEVbp+qdV7HZ8iWMmIXWXWsfHxTCCO
0kocaCu+yY5fVKJpWgvx9L/wXZ1j0b7RyUxuTMmdXZtyDy7Rzoeo0H13u+rFZzWJ
hFldFPfrREOUl4/3bXw3aXYsxop/p28UWAAhAZYPzBkgghyKw0wodKlMgRHdnCRv
KpvGr4+x1aquBl1FY5kUVq2A7E7UYVBBrETcclcA43uDPKEI5ImkAhbPfqB/eL8V
E+DWc2G8n9PAvVpeVv7DrGWPPVP6I4XT50lDPDxKoLs=
`protect END_PROTECTED
