`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Wkz47kKdN0NUWurwmfkm7pxdJcUqFj9f9qsO0IvChS9dhAB+1kblDUa/C2T5y0Y5
d6z8uCeBbk1reTc6JXvsrr0sKjFSM0cmFh5BM6xrKVqKRx/AzLdz3u9Io5qjSQQI
ai7o4PpEl0tJOozpLOPuBtLh/Wrg8KwriH+QYMugRwpHlGC86Ng2Tk/9Fiyx1WTW
jcIp5IYR4TMKoXqtMIzTyuSz24PsYxPRMWqG0goEiXTW3I7MDxiDpEjoIJPwxxgw
K8em/eJTSO1dDoQ6ydM46Vk0pPmRzB1Vn090a4wHdTBZWVOsYoSNzfcZ2LJ1OAYL
CvGD26GNWLVWq+L8HErjtw5GQrOQwpJbz7SiJTzgjbvRxmpduSrrFOT5liUGd2bd
xMpUjzo4EmNuBOQ3hxBMt7tV4WNPtEwUQ0OwHly8kncwW+hoYK4ASs2EDZd+B+01
RHeV8twU9iiPru5tSDNZ6x2LZLeD/DCx0v+HiQmoCKMi2TVgTzstDy7r6jo0OLmH
wEOqFqnIWpTMHk/WyhrI8t+SNL1OOJ1tCK/EZQAsTF95d1WdqoaBOPlCcdRkVnae
D0LNbH4VFgg7eIboRuFXPZwnaNXJdFzCKoyZQrBgSpEOLX5/CUkaE0NbIYCppa7b
nOv2GCfhVhVpwNIh1Y/D2ggMA4g+nC0yQ/6OFHBHUHaVHhLmgxBlbcsiagUhu4D/
+mD0gPEGGHn9LTJa9ZwgY+WVmVC7ANSFFIAx2tWn9kuR0JNmnYFjeKyW2dkep0Lb
+fv2glfIjgaxku4VH0dOsBk7LbPf/C3vNuQj/SXbfnbmgFhRm/yIRv5P+5lmEn+Q
wQxspfiwpMM93I5zUL4NsUvvcGH0zZ/6saeVPBT87fan3bLc2vpdf7kSqi1gYKmq
ZWbUm/YF9xZ2ymOtPuLcsW1Oks/Gdy8Zj6cXi7QGgfP2Soc12mNH8f6UH8pAaeIc
TdGezzTMg/FrJcDxA6UStuCYxbbhqo5UkB4xQ9Wal6JaPQsKzUSffd9xw3Tepr6b
wNYn60JctejXgXVds0+FefRcQSqSkU0deWco5nHD2PlbbHF9WJjB2FT4B1g67WlD
9WrE+HZNKTolJqIqURJiLHa0E9p9qXhNRSaj5M97at1gac8e2vDMQiid6qUMD3cd
f2lTwOIio038dzkcPmj3KNL2c7Bi1IY09yNxTq8EGWk2kUarCOvzNBHHNOxzTC/6
8735d3SxUiup4POn8uhWGfTgTw3YcgTYixoABCdQY1OrIV0hC4UNClLqz68uGc7t
om3eoc66mvdKb/LSf/bPhl3tQ03xp+3Qn86ivPFXnnqXJNrDtAgI2jUhfXIZL9Io
oYjc3ZhWRgMdvEN7BkSa4APIqs4UWKZAN0H2mHXTFbFGH6mj+pskC1cqFUPQk6Di
jKS3zn4BHlxF4IzAODet+uPySVH0jiF8aTBopup1A5VeYjSf2bKdUayPGBm72N3a
sGmK1pzr03/iJHUpTlcBYZ24sCR6RHMUmjmtUT06JFKNECNh9Y0YRnMnGlMUicZJ
EVQkv8Xr3sS1E825XeSIF2kQq/H2WMw/DYNE58vm0hRTGBllc/HxXeVA+4HuUuhi
AuB4pdF895bX98weeysVOwtv/Mt1E0hnxKAEnxPfKLKngZlAIz5fCYCxVaavx0Ke
qxiKAFCzVdtoqlgNo3JRUySnNBBcINoZSQkB0kfx7CfxkHqg68DsX7brxiCNeHmJ
saM1Re4oECYmsS/SMESPVox2W5gxJ4vwTwx3TQiAaTigGNN6MiTDHUs6wNKJGkZo
E+KOAyOYYCcCblzRcy94zHvxsiIrawY/USKwWe5ZW9ALTTjDT3PhKa8rTcAn5NYB
ys6Fyy5QtCXERAvjvRylajThWyHVRCZMaFPKmftzUjILvOF4R5j8h1xF3xINuOWM
HUwy7nz6C6QggEETLRuqB3IGrHnh8qEVIaRNKpcWE55Gx41W+Y84F8FQVnbeyUc9
m9EfcgK41GJfRKthUcNgoZ4PXKwBneF6PLpsaCqMQzsCk6xlwfLvTcaDPoUnFtRX
ffbO+Netd/kPghsLYtCqzJKrsBywy0/HDpquY3+1G/ZaKfq7r57VnlvxBxlLfIsT
kIRSA7nfo7VRThjmDOcdaHdjgmH1du04rNs/tAvDB3mjnYR90IKmm+oGzeZPj7C5
HLXdcEYRKtUtuvtkBtWRxg7on9Xq3Dc0kcjcNoZvBLPx0JutzOWyzNF28rjeHhwP
Sf1RfS8TTm+mLfJzmINAaEaLfVdec5kDeMJIzK1oE/8JPqSRwpi6wjlJJVQumweU
vLfs2oKc0E+VeFgzWehAloIuSbzvtSmNi/Eyp2gkxsuZ36b9sB/vRQLGc5Y/yWDn
UDfc/wlF0yJRKzFbpM7hUTFJZ7485mMgtruTupEQ5V4s6ib7AVGNd8oI0V2//68w
ykBx7vd0FjBmmZOgMHyH7wWwdrz40bh1z1UwqvlBM7Aj2IwHXEO7gLViBExRvjkg
BxxaDxKq0r7/tstSJuhnLaP63hieuBU17511SgcPuROjzEKxRWKtqa0CMu6gpLJ9
P2oxMNTKXjipg5T4i822F2tkO7zC2j3baW6pWPW0PmcTlnIaxYw0tnkNHtZCku91
deUmqg9bsLu5RkfUVpu4FRYybyLh3b68NEI1juJVVbzfeda6qnTWOo5uhizWjE2+
Bs0XT0jNEz3NX7SMzUbPQlt/TtgZYJCFYFKIVvY4Z2kL5AWub6Qg3qNFdbuMxX6E
NzwFxhjaev66UIvZ35LD6wA0zAib6Sgids/ln368zTRsDn5zsFH3MkBsMUEYeb4a
Nt8sFO+ihM9AYlbpm4ifHjUbUEdTmLbF04SJOzCWIcH6R9xqhPgprja0CiX68z2T
lUoN4KuFEm3M005YERBUDwuzXONwg1YL2FyW0A5fDB1lgzKb0fW9nE09G9PVkmcE
6qBE+iFEBZVzL7+ZlS0jHYqjHpLEg4m+4dPByMYvOWD9t0gjb5EmC9V3r/1T27Ob
5QaThIl0GxdFPLfqWh5ZnqAoR+IwRC1ephv8FTJi9COLTJfILHkdwuzzSnOVrhi3
b6rcD5AnBa9Xdgw1apM/7hJCDpzE/yA4tXzAAiLnfn1zNDi9J+CvUZEhOKWidLQl
ugyMVMHPVDej29CXCFIWm8YmrtypFRnwiTYjhXVvUxOzk3P1ylVYud8YloTfDOOq
qcqpeOrtajqDw9IumXFdLyWhwiZBBuhDlAh8B7dhPGIbpeC07o3vd4r2qlXhphym
K/TFtf4lsRJhL7MIh1kEHXgrVS+qBYMY/Ga8FyDV+12qYEfVMU8e+QxBjgiE1Myi
PURK1aOOomxUnJUcHTGLtyUQZEAPrUlfxnofg27BVAug2R9MztdtclYftZWrt/T7
BEUUSM9bunQnNR2eQk5nRz4/cF7mBspN/eTmugcOaFjGVv+eD6iuGhnCCJu9OUIG
qHBVpF3j8WAB838HY3dNiBl2ZtFWcnnCN3ybD7aHYhwwqKmqFMvXSmshfZyGLon1
niKffqVYDGK5cPde7UugcSjgm3h6fCx86v/r3Duzc22OaUxkFqK700N4RV7cjrwC
arpAnSIZ2NCv/34zQazd5qCIRBOFtA95IzZR1Ypr00InlsjqPk8D9BOtium2qhMI
jr7VW/zvWl8XGoYifHfsUz2V2IGWjc2oQawnehfca2VFzgKZeZOfgTOb69XhDySp
`protect END_PROTECTED
