`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FA0m67NyEpfioe5D5BHxLks57wvm2qLuRoBhh4mYLa7vWdZU4H0/o7IVYvIU8bfC
9eOCarkZhp3hlidzLgucc9cwoesjqphLUfPi3ad6rc8bpVktAI6UEyWjOVRw1Xtc
9u8Z4myMfurHqGYID21ZtDf/MlFvVlLqmD0rTd0IQysg6TRGha3ymU0TBgdxyN1R
BjsQQk+9ug0W3SG6bRwge0vpueE+XqI6XhhPo4AsLWRTfYuHe6ueWFLlKc3Ypwx9
IIAyvD1nW7elDMXba1VU4/FpRLw6dOdCwbzjz6dvdipJMk21vY2mf2iKg+DOVmse
sfalRJEcQcAbAJaYWHXqW/Y2X6QtN5pv4gT2j6vfMfvme/UiPg/xniL5ZmQ05Ki1
zbdS63QbiD7s1vd/fM2k6jpQrf/4+jm1gl31+K7G4zAG0uUt+ql+pIn+lI5kYTES
v+NHs/KtD1CeBkygZpAcH1DiDJkJdYB+fzytvZCLlW/jO2QXvVMFCwJc2Voaa4T3
Qwb4cfdLzXrksEDxpbMb8d7iEVwlT7htVhPGk46HJzw48hb0IWw3CbEzfLtoQdAb
cFZQozmFpo80VjtgWHI9tLXA4anlgDPhILEaEc7+ixm4AjLwr3dtV3Q6LQQdIF4M
t+w5E+P3LWtHrr4se6YOpNTGYY53TpEj163Xaftzrjst5/3y5PhuLbKul/0TzX9H
ljrhmIjDWiLaiiBrCmdDqpUMzNYjJiX1pYufu9+xzHRxJI/exKYoFdfr7sR/QR+Z
bEiHK708VHTxPrCYV0buvloFhYCmR9TlERBjtfq7GLz0F9BCLp7jhWe3A3dVms9I
TZyhGnMhPXv3GassRe3VnK+wrhZiMJYFpyTDfbxWLYGMxjtsThYOX1P2gPcXWmFC
dH/clcIIQMKJF1NupfbE6anyFrb8h5zrAcwj3xC/B2GPOA3WSrgt1ss84XgUS1tB
t8bikSphBbrwbTU2zd2npvm4fSQfvctDSdfIfvi8xqNFmPfBKRAoRMDlwmkWbNpI
RMYhprctxHsry9ouvNNZTZTN5AkHBskz7UNtErQUe3cVfs1OuSGaPRlpYrt6PWY+
3W8TTDdUeXdYaco4oxazdbD8W7xK+7odHEEB+GwF/5s=
`protect END_PROTECTED
