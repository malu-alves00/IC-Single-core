`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vDAw1XXH/gp3H4UyzNCa6nG/mKkLEf1rYWxZudTE5PiglFeyQTCPTnSTDV3CjToX
lb0emCj3pokoqXo4Cd/Jx7mqn8lX1Vnu1kFNiJ8X1oIfU1z7qfhDVPHaqc9wjFis
8uQTgs9ielsBHcfD3nEajWlOe7428PwF360+VexJdUyjYeUusGdN4ORWh3wu5zBI
SEo7rOnHZB1SmlD/Qu9mbRCIwLWMPDETazAUO3vwV3yMoNgzxW81iFqjgg7X3PVf
kjFUY+xdjuWW0Tbs3VnYOXHrkSi5uLXraXbhFclgAvL+ea6Al0DwDPNVrI7NB57t
oBgk0AbepfnqbdTuVh0Ua15jFy9q4ESp35hrPyDllVFi5tSI44yj+/+MusUAktNA
l2MIUIqCM+fIN+GeFaQhNJ6Ma9uDBJg4vzwvfj8HeEA/FIdBJ7c2A/kvas0ih2uJ
l6ok2s22rnZ+YwkQtJQwLuJSHnNwWjrEQIX06JtTBcrEE1+lwBTSKs8uNDoqRNoJ
8EOnnDYjfyS5a/9pbnTJNAh5bavl4ZJaUOvuFl50yUvtV1B09t5MsWfU7WXvl9an
15l+Bn0E4CuR0jnRoM36PPd+TzthDSQuk0T7lvDGGm2++UefFpwrGWw783I6gGXH
RS6p3CAHDbmKaUjTALFtY9Vea37tZgSTpar/IGAbFNlDQnT388X6Ss1VX8XyS4rL
ImKdF0Knr4cu1VOOHnmN3JO9ZnBageGjMIBhlhWvi0mBWAKmaSU9psQH4XQst1ls
51h7snNyMBGPRQ0eunpwkELqkah5R8LbaJxopeT+Wdaa58A2DqAaEBkWS2X6L+WE
MP/6/zifhzH0U0hoN6vHJQ040Wju8RL3etnUr5sSwEJ7NNWkm39pwvgBpILofV7G
QN4MNrr/lXOW2i6NiE0xSZ9/tuqO9O+SkksFWKqj3Y5FsBdNBhc5Xfw7/WnCYacO
tpihxjO8VXXpfgEzXh1FQOUXct1bu7Oip10VHmvcj3eDdiUSAtZ0zObbRE9RJ4ok
/z97jPSTgVJEMAtCaFuZFNKOp1ZJ3/SecsmX1JU/NMKiIxYvonVAOoiR+/s4fdEb
`protect END_PROTECTED
