`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lRetx2nsSNyFv69TzgYgM1ks2jSyOWMDmitFhN2tF/Y/32C8P7racfM+C30XqxRT
VredDJdUdjtfp5DGC0U8WAmyWiYh8u7n7YWD0cdrqVd3EwKLYtAn2+1Az4DqU/w9
r9WQsccSbcMY5rqHpcwyIe028Ynv7nQ9/Iq6SVbqs5yf9N477vN6EjxnPuBKrGAV
901SkSZ1IGHm0LXL3bf9cQ/mvZfOh32kxoWTC90fG5sqrEHNvVnkYWsUBbe5jUai
qfyiHwLRfq1mOwvSSQXvEY+1gi1uaBG7ovj9fTLVuUrSk8QiiYcxGDTlkzWoHv9b
pcdWHOpM/2gnimz9qdPd3O/dhQhqa1henD86Tbv8hIyrTkkNzBZM/obx+a4M1t4a
xFfVa9gMSdjQvem4PfG6wfC3xMBn3dSFB9Lg4gil4fMnsmoL975CuGWSpUi4G6Fr
c1D+spy606UfhVWz+1zhySIS/6PUFrh+J3IZ/LGDGecgsJz05QGbVDc7VD/h2OSj
mI05unW9Jr407r7492t6g122vCa6c3Oe/FmLrY4CNR1qz9Gt6eIij+4+AGDB7OO4
KkzEY/ky3JrcJjxIDZGsh6eAZ6QQKNrE1V5BCJ4blO/J4YF4reavYXAUrSlipHAZ
g0nmgyWjSAcrHB1QTRqKDK90jhTa0g1W6HWr173mZehdP9Hm0MUxm5piLi1Zp6RX
S57Lc/6ukQAwVPtxno/ZRJW9gMKxLvL9IqC+nEBtRLomucwADpf7EFCWPRiBn4G9
MDY+3tu6ST3a0Zh+VG++1m27qP1LLLyqbhAMBM9LrQo+sLPo2061gOXgaOJr0U+O
ICZd2udrHPvlqAkDKt8SsA==
`protect END_PROTECTED
