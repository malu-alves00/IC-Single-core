`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cRAFJCDvlAPF6IlB0wEPE3tJbwS05D2zQ3PE25wetSo1WqqgULnDJ7L/llG0gLk6
LpREpxzU7AK/oKER7emoQOsJtPNRQVBC33sSeIGEtG35OeSdYo4aAavOlwwdpFC4
E2vWUS9sNa87ax5tu9EQT8bWlJ3bA4pjfMFAP9tGlHYblZDHL1I/TdWSLeoeHHLp
wSLt8earXdjiVDjNwcBeGE47PgwD6uVba1/3N6+QELyIrot1sR81D+/08D9IYAHb
E4JWtjiLo8QzC/LJkrllvVX0T1E/05q29oCD//8pJNlNgNybD/yAVeQ9fNwnRsqX
xrG1pQNGopfmOgQ562BX1hymk66u8fn8ijKLSt9wNMIr7CfjZsvNraU0W40loGNf
BQbT7QwN0hnnl4BxbFr8jXgKfsIiExWCMCEMCPfyL+6trV4SDkLGDTsnspUnuOvC
6amCsBuvQjGb1DkJcCM6yxFcR4HxmCyoQQfvzGX/+NFbZgOtBotvdIjWyM3Pro6G
zCfr21991bAm6A4rtgCxCF9mmFmZYx+dMznHqj7D7IOrJLubiH02XdnL4Nu2V9y3
NgohLji7fo3W37vgB3rjVqoCuK7HMMUk9/766R4P3c+u6i20lzF43Kon+JP6TEYe
kXqaSqVHAxMIV6l1UOgdYjlWElJP2LIrNRFWGllMYUz42W3QFhWeabY0YTavkdAQ
k8mCYkvigntftxvyIhTdVReg6lN+6fAekEcoXOZAJf2dt+ois21kRetzhxY8pEUE
oqI5CYe9a9wfYfekbyC3WA+1+clzgxwwIUtIYWw37oFQKrIfp8tPsGZ85ubO3orO
no1W1mjcqVijHeitrqCdGkGr+mr48sci3yFdZl8d+hvN3sYklmlixkYRtClfpmlp
VlIIqdkGdveKSrhuxGzwAozjJ0veRImvzeu2ESY7A28CERJxjdDXz2fd+RA5M/W1
15bdp5OskxIP7lDtEiRAsXUrPVALry723mve2N4ySFb2o2Eyo3khOgWJ5HhktNYV
psGG2ZL7lWdVqCOgn0DIvNFFslCmOLwlMukWhCGVzVtnopc5gFjx2UfK1ueCDbWf
5jEUy4erJzvh2HbQC3Y6p3pidNr2J7deUSYOFFkrhfR5rar6QKyfphOUMNc9WRWX
jkvX/hrE/gpnwM/AXO+edA39ENWRiGcM4C3MoeMzl2mTwYmci0QmkvJe3cx/qb4O
tl11flNAJsnnncIkvC3JHYi2IQZQDYumWwC5KTiD1GcY/VuZAZkbNBG2E7ad/hYQ
GHNKdFExiiyVDPvm4LnhfT5J/yPvO0Bkod/ZU8rydWicVnFrYcgwC2iFsTj3387L
y96RLlUnc8vxSySJejqPvpOWjiq9PYwXuohCMWTUIb9PywXUNBYJDnYmQBagOAVM
r9Za5aRzhJZYGcT+qvxOYgiYm6zWsourJpqmJJ+eOrDwg8xG9IhUdWMh9pobo4sx
5qCx5GJXLM3myy2eBE6AEpbsst8E06KueARrZk2oxcv8LIoiYj+vK2ZhjWC9rUpS
lHi8L+c88BIMIL8f76riFQ0aUPb0TW0F7Q0Yw4oE6813gB/mROxFD7pkDU1hASXz
y7NuFio5WmxdpZdYlaTgM7PaCCDWqUDcNEFQ2WAJWvAtHxtW5etap5DalC9Kq/IF
HDlP8UslYLP/eP5a+dEGYjKmFw6PwKklgxT1XEA8QsMnXgShPDZbriXf5ShuUWmc
lu8Y4LVaF5jf3OVf3ZKIafyD7+xl+H27qxgb8lNRtLDoF0ayuGKBzz+sq8Y3NRfQ
MWH3Nbd/+lXL2z4HYHBRLvtkDvvNQi/VWSwuOhPeTzT1NRJNllU9M03JFOwVztin
E2M6s1XzF2HBOx/3zF/BgJibv08HUTsYizwzN/XtA8ka4pBLg6W3mv+AhjZeIhbU
0QT38nKIlo7J51O6yKn1nry/ZwVWeNGHMWpQMaqr4OfHyMsefeBIJLRNoKLOFwSU
+F3PUefaMd1CpldvuVctciy+PaRap+rzVOTZOkxYef2AwLao2PYx2JTc+2EcKU8v
P6VMJXz89Y7FHiVGndjQnToRhSkYqdB7bc0CeNz79I0EfiCzDcF3aNIUJx6LEUgP
IN8J2rnWenWbgc4S+pAyT8nnorIWoJX1hT82sdChgiF7orvLLmaxcNKcFqyEG/CP
njk/EKzcgtvpxoKXXcQ8ZC0RCSqbmsT24AZ6QMGWBQcIdQ14lRF5hRDrcRLIpj3/
gTQoZjNZCBeYWLVNhqX3ZfDQ+j9j34MvlnP7EM3rxhy4wVtG6LXbwz779NpU8mvu
3gEEYNHviTAv6yJTZH+Gjx4S26bFM4l6M5M/Z9XWNDzEaxmycrPuE7VMPKXgCsQR
qYoTymgvgErkWImb1EPBdxDsLajs4LhO8tUdN8C5D1EwuIiq5hs2ZYfJlsxkoeRz
5NGHCllxtMMy2b0L4re7EOtDjQRk3wyib458c21aX6HiZ/y1TbbJJcJQt1PHjb/E
vx2iwL1fKVjkwra4OJR3L+hSVyzjSvlMtqTj2C56oRAeS5nI6hyZSzdVOeYIdbem
yqFQZaX/BzCQy6OQR1NOZLUwsB9oRyRv1l/rxb9orZyDQLlmALekPkCKzcy2WF6g
PqPtZfwfPg15qsGSnemPRSEb8Ars31EMBuXTVbHcXJu1eT/ffly04BG7ELnucuxQ
ddNW2/kxgfOpnvBhVZV8zQBna69z2uS1xlRFgEcelMp8BF+ze58oQ9F59J2bM/AL
ng5q1OKLG0xnY1hSoADS/XSGjmMV2HuLDXQYGApr1EvC8jmtITz/7KE3gcSoakGR
7+k3YNf/D0KYOqlUjZijhc5rfBTtTIgxyL/rIXt4Em5uy0FA4xWGJGHp8CLYvAJI
6TlkFWdUY2fSvscchMoj9XksNNvHg9aZMTF7vndA8RKYqC3zOyPcMW2f6a6KeK30
9eUTxi9/cyviRtQqLQd8P0/+8bUf8rjhRyu51K2hIJTxamc574323wAGUHAeyJNY
05j5xa95MRxfl3JDUJmfp2M4adKRcvnrnQLzwcspg3BG7aF8eCEp7rcugX5z+BNC
tEynIiYV+t22q7W3U7ttsxQvH2QdUjP985VX+MT7rIxUMmnxjKqtkMyYFkrnuMWe
6KuRuBzae/8WqiFBHmkfUIpbWxq5wsqVqTQtjmzYNM7DbqqhZ6ckcWlZc07KZpsq
hxvtTcf0yFsRcmmodc3XOSo3K7IH7WiGUOH8UIbv0nZx3SCrVy4WQCS7FgBrhS/f
nElMAv4xMw67oggGPOeWTVG1JiN6tvR/rGpLYPjlyVqDqK7RxpQTu62R4wY8jV4R
s68iRo90EXKVG0O3VemCVvd+EowOLahK9O5oj2W93EAUQlNTtiFdURFm5tsDoGM8
jTQ6a9XtL5FuINc9vGwnRDjxrAuUcX3GUxeLcHIHNYMtPzyhzGIYlQ+vA2yUYRp8
VYF0A/jIt4AVOydcU+NAWzhS0MTd0AFSI5ut+QPdLjkk62B3F9mcMr1+mupokc0Z
DoDS0wtLs6aHI9J75A5GDLygeAkHxd0HnVPWnORsy+m44jbc343l70qmHkhr/2So
Pswj6mLSVDPxeWlCFrHESRSAf1wA45Hksh/Ut1c99wjOCiYA4He9uRAeaX00ow0f
zWkgwuVZ+OptBGtwFbdy5J65ZtBHLnWxFSZeYUSr30toMvze2+Hip7CZ5GhnVH4j
BgK5ST7oFH1385q6p+paj8WnEsPuuNIXCzXtLX0P/ctvKzFQqltW6Jz7KQO+YsaS
WSHsFUN59FXmfVlKt71tCpzxQMRqimFUt+NpNCf7KedoOM36pNTR48+Tw+R2Gjim
/9ScU6I/0z/kfUsifaXZig==
`protect END_PROTECTED
