`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3dWgKPiBz2nX8tZx/TW9SdowaAe366HPiMPLDMsT/tEKrOtpA019I0uLIBivRf71
SHKVtwLMshYDoJbo/G9yl6kNepMzaAvqwJ4E34iYvOqNfOwptXLvwtnpmVg2qJaj
7Db7Q6CLDoROtYG7J8WKeUaQlVdrTckDUpAymPqaZPIpjU90u5imwGkWQuroDNMC
V1dDeQsiZG0CQcZLQF4Ir5LjEV6JF2HVuG48QDBQ0Bihy3+lU23SWveda2MK1FpS
aQifaQqkoz4MJvYB+2V2SGBElp0LtmtMnlkSO467huXZdVf52dNrmrk9ak6oVQJx
ghqOfhS73b51EIPOWsrPXvIdbRagdl3sqFf3f3j2wop6O9inV/Pk6YkL3NaIQsel
KtdynOqOD/OMmGl2reepkVWiJkNE+riCfbUSm3s2E7YjwJ6ZL0D8lNYPjfh2hg4e
1easqlfHqwbLjiV1D9K1kgB6bTbUrKXMO0u3O/X9L3DngD0+KS3WSQpghauUYlTg
YUJqe/+3OPn/N4sXKLPeNuaBubQ8pxdK5cZgZCeO69i6NwvBRrDrcn+tHb+Q4QR6
VGQVDocwxH0/3wD2IeJ1tyBlP+AZYWdoEp75r/tJeNxHkfIoHrr0RJR4Uc6AtQtN
3zSVLY9EEo/kTQPe0yvTbAPlrje6BrWR6oUSRtDWldo5w3Cskv6aJTJyBYOjMx99
cRf4QTREskpJjYO7o9iiBC5LKIWrISSYVDdV2BGyXc0VzhhpxbuDPmIhtm43xKx/
UldVHB0tJ3NARUa3NG+Ao5aSfSO68WpSUgElGY6XsAe+2/krt1XMlvohr48GsHQ+
AU+GjVKZbhDGqmLha9Tkpdz9h5T/BgrydWZVPQWTxWfsZQDTmC7UQysS3EW3Uc4M
fv+wMdm2Ag5JX0osBxVz0KagARV9dchWKR9deAdJoKoobB+AoK4NAtuGSdavsrAt
iwlQwqAe9IqfUIBITvqpxDEhG2f33N/a9wgYWGFlhAyZVV14a7cwmYwT7YW9uA6D
Otx56hrMiQkCVEf1WCovLZtJwV8pHCcO4LEi0PC5stxbfEhQ8la39Lf10wMPnBKu
rpTg/I3g2k4WHD5LWVCEMKXO+Lak68Lh6dlzr8xAKex5TUbSbvf3oslTMh45J8Nc
lXomFqdTlk7gaXyOyVwEk5GlMwJSxG9TFsmHOn+Xl1x6B5Rmz9IZaGDxQJMPRYve
kB5ZOMxJsh1h8U1mhJ6EMjr70z1U3cloC1e/IZ8UhFZwnky87UkUWVahGCaQXNSi
C1kSQsLue7Z/jQwd9eGXkqkvwmEufuAu3SWkg5+99CvJSjBYPjOoLgVa04FOIcn5
6NIKddTh0Z9nQP4vwNPTmMhMLlV85QhcQ+jX2W3n1/GtWfdfzSFPl9qVjzV346A3
Ei6EaZDYdRIh25jgQ5IDwCxuJ0W1eVkZj7UFBpEr7KVM/3bz0lsJYgfts/gWYA1E
3p2ozEnovxLpQYYFrmxBiT3qlXIdF8IvTQYKlNcLIxc2NFrbtVVP2/1h0N9ud2+4
na5eL7qIssBpvZgBtyaLvsQNa1avpiWxHDAEGVGg8NuAnBAFQFBQ/G/mChqGx770
FXBymLJ6WUU+AwAh+vqb6a3OsfhkfKCb5tjbMfijOjA/t/+sWdg2Rx3FLaU23G09
Pa3wVjee/f9WmC333LldRoAU3vnuSEMTi0cQlkj/vv2RX2XiZfnQhlosxaool72p
l+6GFt0jh2aX/C9GzD9jO7vJRGK+Jc3TxPTsveev3O8cRh/oEcO9jE1m0neGNjFF
P6ryp6xfGz2CGCmJVwbeJ8Sh9XMH8nmxHJpMY/ZSN4VuWT2I+3ghtGKjzpb0jql6
xJEpmgdWeGOjuB3CLflqIZ5HTKW7jmjmSnsfydTjzzf+7LGhjeRSWx4It0wAH8jb
rLN7oz8aYIK+eGWrEE2dM/QCAyPebWAJRJ8RTszB8es5MSaRJwecjS3WFYQjv45o
uRg2XLjYEVerCGtFDS9ee8BvZwFCxypcb0MEv+FL/WKIK+lPJsPC8FjVkh12bGOA
DCHhz+4IenmO4q37YyJzm1uux9ak/c6qSIJlCtXrnCj23mwfUxj5/OwY9dyWWRXB
T7/2ZK9wrzjbTPiiCF1RBdUDsOC4iFZrz7bKIOwM3PULyQCaFf9F1Cjie1yF4lD7
479hi80FrhKjHnIiOEx54BpwCkdaTTJNxrQ3WBJPIcBE9Ju5mhvITy+39P/fb80i
JzzXApySC170DBrpXmfTyN7WRZ8tGT3IeMTPFvtauge/vRzCK1gJl6DHcIoiiIQa
NWhUuH0EfY8szOX4FXkhodMsKYy3N4Fjb1Q4CnvPNduV5kH56J3+FfzDqMLG1HFK
62xXOhDErtrXJcS27X46iYUNWUSi1DB3E0p7pjlxzHYXeYa+VlwhKwncos/xwjf5
hjAyRczIAwGniqz7UzlvCeroJisdLESA35sFICvAiS+rpZ++UxShQpIXo5ofgJ+m
yZzQZW+lARtAFxuFzCrlKrbXh9FoW7sSRxtIyQlgYFmwnZ+woXQqX7itSWH4QzbE
EkpfiOkTanAW2XXJvIJchsZlT6RgHDbNxAIxvz7GxlAkbAyqkqDwB7VpHdlCbsQt
ZM/TVV7IRB0mpeRFSwpvDxGxKPlIaBwnGNNi9yCFhyb2apXTyk/MYgcx4mSBsifV
NKHrphb2qOGrtRx+Q2+KL/Mw3P4UGoCg/P2nd471oHnv2dxcM45XNY87OFTnjGyJ
YFtKW6wJmhPc+sUT1DwwfTFBWiNAMx5wOXeOd+DVIxZHQNK+2VZPBjhcpEXpsLYw
CMeou3hHkK1okXX450PECzKfhsyqtvb/3FBpcNVrHwapi89mulzv1C1S3jfV5AoF
ASW1c1RS3QSBZ67I0J2+1pmVkWpHKXLSsJhLzKHr1bKr7SLGbhH23OpSIsQfh9HO
7I8zbXq1MJG6SmyWVi9j1LumnfQZBEQ8WwI1fqt5JxpF8uwC795puo/+xYjj1eCV
n1mCDKuqB91xQAeUvwlGvNOtzcUUoqIw8nHtJ3GL1x7lGGMjWU1agaxEE72utA0g
j455TE5A9VAEeknFX52xvdcNn6/xP9pySzmq0D7w08xNGjpZ7/GsB0U89cRd8083
EYWNr4PCs2SZquztUIGy52YvIRw9M4ZE6rqGgZqmPQ7JaK7cGpZRw2Kp4PZVsxqi
/9EYC52mFJOvuhvGp9WF0gJ0Ubs0pTyx8+rRpVxr0zFj7xrgSphTs7L15OZZrsmi
esvw0IJeDLNygQQ8Al01iageoCwQdEO/gWbrVARMx2ma3wP+4fVViU+yArKwrcHP
kKp8tYrHUANZTVy7Z1gPrnlnT5Kase9uYh9phE4W3JoSUz+wtRUkaMhjQrG33ygF
OAm+IDtnMqQd/bpl6VGP0+/7SfdPIRj3+G40JGnLB6WI5n750FE1JBEd9JQsnm8w
doe2t+0c7NP+mrlUhcsUVbX4fsVDcmQHjQlVO+Y5xisHpsMZzo9ZXm10GzUaHQV5
GfH3q740+IfDoOHOpztEcRUoGsxWYUG/a84KESPLK2rgbiY7zX153CiKNW/EziCQ
ypaBfjd3PNtio5A+Ttx+oeTPnq8OA78bJkCTwi0cZ1JpIHDh+ZUp1BA8deR55KY7
fd1upOnofQNcrw9X7lwCUQbcWiEw3ohfy9Wst+0i3dRJnsdktdgLE25XvfurOQld
/9zFRgsZ/48XKorTQCK2F0bLTnsg+A0dHZSMfMrYLyXURBgu+uz152hp7bpFfkLq
2jiVZd1aLKY70GufvSvZw5MIalJJBxr/mA7DaJ9ixR3FRhSZW8Jqp3bWXsRlyOjn
lHel1JMKQ4fXE36u6wA2rxF2rkHqYfOWJa9oFuQlfh/9vOnOAg0mYKbVTyWjFSMJ
C2ecqkp8S1hAwjQEgZnE9iTeYq0wI4w9btq/hTgCbDesNpXFdmVcEoVQ2Z3P8/yS
7sRX2pE/W29iOHa9A4IB9aQdpYBwfHSG/Ks3SI71N826GCJ6VwvSRII2HkfE1Qxj
C4UMZeCkMN1inlNC+/o9eQsraD8jUOavqkU0JEy9PAnP1cJEA9rxvcVGhGCaQEBP
TJHXVUgL6/5Eczu+59OiLJTmjXJtSYShGWEqBj3xligNjDYOmRH0GsfNeryafCgu
xiw/5QlzjfmA8ALsB87ayo7leBigz3gJLuf3rVxfZp8D3zqBF8dz6Rnrc0x2Cube
sTXsdFAi1PHEMC/uD49L0nJcQZboBlX53T5cOOuAjoA+J77+uIYK6yj99aprbBfX
2gPnxTWW+wSQDIKPJO2lW0XrVpaf1eXC/neIRPwPUZtTB2V8IRawWkR4ub6gewit
q62KrLUmp4lYBtt/pH3oHDkCOLN36hyeIkkB7lPqNyZiQqpZQbvYfhsaS9wr/qmr
foEt6ohNlBEdd1AtYUwyWjX9DQG7SjmHBF81yblrjV8hs/Ra3vgx86jH7yanXRRM
xSHr6VfOZKyJFhYdtgMAFUwMBr36votEJAjs3wD9cNHSX0O0pD6Ju/l7pqFnG2FR
6gMzpfsNL++spyJB15PlvuKVBvLYwQcOmkIKCbdJmxvK6KhTObXOmIbWZrQ3XRX/
JtGHgSf4b1RfaPOkvdzCUU0KOUV/gss+AwQ4IXje78s56tkx5UfSEkPucUTJlKi6
XVZQbGIiIZP5fUdLIK3vfvpLu1esyk651T9+XHFo9Ebk1BJrulJFbHI8p57fcOnq
lpYEmWTNK/QkRlfr6oC8jb0Upt6RUd3hTerOS2UumbfFAuWKTnHqgVZ6ydBJMBSh
rrDffoV1ffQIGv49QhNfkWsiWbLL3wHgdW4ku4CqDIu/GjYCErcwTEc7TH5Y9g0G
JNA31qTlhD+oa4SClC/AZRl9OZ1WkErOZYEnQOCcc1BKJ1jTX500Ael9kDH8s9VA
6/JfFRzcOIbZp8nZ3ZcRLe/mJ+Kv3HOwQw1Q0XQNZ0KUdMl6MYcM3KmNsS1MCmdA
fuusgyvvvbNGUa1P2iBH1EP7OkdJK/iPV7VdSNiuls9tbF78KXBYEktIj4TGmyBD
t/tZ5YIhxxm38hwZVbNWMVrX5Ea8aH2+SUIUOuliF99uKBMJg9hUD+VyzCAvaBBw
95mQ9ibdHG+cfYz5LC7VJi6wm6raU/0KqSOVpejfF9I8gunENBwBqXsZk5zxxrBC
GaBDtQ+ZpM7qPrLR2GNCW9WjQX4IPwEQxVqIoBZiycItwJqqFGDSkfY6TsLsv2tv
x2zIjb9g/9OC000ByzX8Xi6ssCYFSc5PvPchtQIHf/ylLFW0yTzMIrExp9w/bhSH
7bip1qleLKglgCVRVYCbiBgTeqbQ3vdPhHLcG+VZidKdW8pUx6YMnz8a/Rugu5Be
9AZ9ohpqdCfuZrIH6zmKcq1EHzFRzXf1NF1JUibq01Hl1I5Zo1MsbRl09bBDSdCR
t2jif881jg+8h4B79paNdurOVDAlUMKFGxHfTPqeWIRfkZuyWbnZnes+jAfQd0FY
ky42LZTQj2QOJEAh06RnGkHw/20eSf0HGR3AqCuZAtFLR7hrZ5Mvk+xJPo4blgQg
QNJReuS483qNOZYTwUSrrF3tdQ+kHBa1RXoX8F5eZP0HcrcWQSyud0qN9t46f7dD
lWSeHB0t/N8oL+kRgwMaQGEKZXgdjcX+zzyS3nFQe61AiPv+8tZvzaQyJIkitD8t
DeyZ5jKJR2QEmDtSRQhhoh9mH+WqR+BG4Ix3JHglcVjx4aETnscv6zbC1PSsXzbH
tBfrI1D9ZqZrJ398ty1S4cVaNjycGxipWwXcvk5xr8xqy00LABl2vbUfCJrFW9V0
1VXOa0sIzpEO1ftlVKGkmtnHDvalE3wXk5GGI7FGyVWB3u5so9o1uGupk9wjW8ZY
w+B36CiX2+5wJJXE2WY+V1IXYNw+/vbTwP/wGQDkEr4NGmdHFyzlalfPTdJXAw0n
Sfht4TfBO6qPsbwgGfTVNDjLU6me1jv3ESwQ/RQWWc2ca2syFCKGav+gRp7CXmXI
sXkkNpVEbMQsQ4kUsB8s/OM29TJ441rpXmXKJXifHf2R5cyy6P1IsZGjQh9jLo8o
zii8bOzrfjdjmyMXxkgyrWiXAOHdlD7wfwbiR6I5dumfu+U+lWg59wsTcSdG4cz7
ObLIcetB7uJTrFT01wkqRkFaXIL8gR4HmIyk0cqtnYZPbxHlKpfw/ojTCgFyu3eN
Wewz3/otFR/d+wQFExPnBpszzMdwBFX4bam9Hx/Ep8u0+zGZSOuM9Og9Dry/OQQ+
PV9q/BHEiywqzjNTqhSzpx/5oBw2v2v6xVWegMK1XIN7CeIx1cq1Lq/IsPzFk8Cr
52UaVKHA5LUXxRgKz+fOgqw4V8fhrSJBgYXCbzd+P0KvUjpaJXKw2eZjPJHafHSW
+zfm+0YJSRIYis4EZOzZxApjYZ622sQplPd9syGb9CWOP4ymHqabO+0xyjK90UI6
hwBVQkfNUERy4bd/rbtvH4D33QbCWbcIZ85VLTHuwVlf7cPEM0HjGCvASiDhT+jR
zl994UBZ8IF0ZrOzEvQVdO49sgejmYXX/+DOoNH7Dh4dSpX74DUHY5M7WkTOX3/i
8/ZuISEsZuszsTfGrfebDmIk7b3pRf8JhFZGDeMBVjM/NvZQwtMtrF48ju43PcZb
g1gwRAogJ5uN22DVfSvUxnAKTp9NhNB/37zzaETCD1WkOfgQmwq2AZorG8uqvpEy
nzfsFgIdFeFr9HRNva3drp1D/XY4jvo1xC5Ga5g1TnM4gYdFq4r0FSQDJTI2BDJJ
9jCfmt3gv+OYJrQUUgSlU0QpmY/L6JU/GuRge83lcfiiSSA2lDYC6MbFocoamZ2Z
BzyH3jmM6gHYtDjipa6Ve9/14WDGY5ksanz+Ox5DuPSnRvB9t9WqNQjmbSjw7/2/
p9jOGuSW52NMlCLQgnbF/F2zF8QE9CGoD3YOI7ZqVNlVzwWmgjnIxHrF1MbYhBtN
`protect END_PROTECTED
