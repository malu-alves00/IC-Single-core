`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kjXtpAFfGiGGgJwvuSuY9rSgQxEbw5JBbucBkEwnD4r2hXZ1t9sszmFR4JhGGxH/
Cvhyau/PKBqWEWqk9vwAPDarNqhNlPrAguEwBKdeuOfCsV6N54Zln4cC17jUlUOR
aznHctGjMR9krtSkdInb4aYBr5fBpodGqgBqAYU2SKNkAZJ2jnt8wkc5s44J6ZGi
BLkme7KYCERGmqXRgYj5+sJUkmkDPmXmlmNyatMXGxiSceQL7brol5dB6AsWVfi7
GwYo1S0+XN7MOlkAARY315TcyLV1DHDe6J7Fu0N9x80IWXPgiWH3b0HqcbDpc2eU
kjiLWbFv7c1UC84eVLNl1+6mTzkUaJSucMUzlWz3liJvsftqH9vKnZRSgr/cAdcl
r17q4jEP+E0xROvELjZsh4VQYJuFFILum33ch/o52Y9m/Hjm32c04WQNhxfDZWbs
QaKpxUmWy1Qa6s8fAvFky9j0liC3ACt1uYfyiIOgV/+kUin76smigLR6bmHTvQ9o
ynyfB8RZYjAjuWtHZOfCbRML5wxIhquA4NyLXb0MiSIx+AhB5H1z32aU2ggLcrwe
FiP66aVdw+kX9u8IcHq23aXi5DmtFsEJFhgdF2FYv6tM7HklGQjfuPOXQLulAgvP
Ixhxl2SCXI8mFSBJ9b4IW6PRjPUTAoSSFqFqsaMCAJh8LALZIP0XIH+XlZhpYwQK
Aky7rLJ5hPLXl08tPsbO82R5TTNeerF4SG8fUTvVQ1c8D1rUC1V8ujsgigM6pphn
9RHQDeETSr2eelFVFxZQIa3QYW1lsLknB1qvOnVYzHry7WSWDZ3cm/yUuRJoZeMP
`protect END_PROTECTED
