`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uyqALG4i6ibsNRCAXBt3oggG7Xp2DPGOI8Jc1o3A1C4TIrEdm5bYpOCZG/n6WSN+
aUAFnt5ZEDGf0ndX3wQm8Z0dbpagANVVC+RJks5I+RQf+c2jQD4vborDZgz7vNIu
OemIAy1OtbbhrQCi8CtjmqmWzVUwzXq0NaH1D3n15FqXks1tKt1SwHb1OtmHTR+g
RGXR/z1KKUqCTyL22nbsCIuVsE8cVHY/Il/LfJEHVAwQvNmrU2gZwxWteiHQNN8P
jAMVICmnSaSsFgZrUPweeNgjM3CU++BdU72AFfSQHGVq0Liso2HtbzvJlJ5z0Fij
dokcwmcVmw+qvhMvo/I4KDbMluwqHipN6kaFPTqBpgPG1x58sjpyNraRKbD2Zvnn
5kA4HUIf/YR53Y1g6hCPesM2V7TPsRFQpvAb31b4OCy0Uj7/kBzzuuHaV4He/CGs
t+L5AMJ4ServzVd1S1cwbAg7zqFnMFUDDo+ABEFqzF++hACRPwXIbaALu4apdQXS
dAJ1S7ii/ka/wyMUCMucVP13DyfxMlp3xX1KI2aggYVzCO+HSBJ5kHLERxNchSok
genH/77wWqJL6/3aNojHVIaKzxlAd0NynfwT2BhUkz0ZTYv47H3dGN6BIrmaAdBH
V6uOcbNccRt55Kv7n0ikBG2nM39TuWXCwIfeeTJUaT5NahnYBcLseCWrSv+nnlzb
/Uj9aghJ7EBNgDd1Oj3sCJXKDmi3r4j7zMCXPXhvX6VmI9yDP7/H16lwGdBW501h
Wt3OfF0gz243muy9PzES9qVMe7/Vx9prXifWdNGH7SHZR/e6Yv17tcEgX0sEjb7W
I8+8mZF4qY2kyaQjMQ4PXomoK8O0h+gakdcLEPbduvE96Ww2YP0tgnHUOoOYipC9
u2WsjTiiB6WR9HSB1XOaYyr+ksyAo9mMZB0DLWtBI3gNFtHxn0W0sRFRJf3bL3tY
poT0Ig423pu8OiJvCNQarU52cZWi9SAVsuwO5EdJnweDXIR0s5vx4gLJxJeA5dNQ
ou6cl/4YMOwUQba5zQVVdP+1PVGs2QABFzEW35V1pk4KDjuK+nYEHUtmpDeFtPxk
S4hyff0/byvLl2Uy+Gyspnj8E9JrkN7nPtALqKMQ7g3WUgoOV1aMPHCNr8rZm9wh
DFZd+W9FgYbTqYbXyWZJMKy5VMnduc8IMmI6Hvp8zmsqaZpVwgAQ9nZ1ltQp7q+p
JSywz2IDUkx/k02tblBrFqERf5aqNGELUTTbadTcpfoekSCP/eqzxbfxPDbcgBtw
DP8L6E5WiK32Wb42tQD3OUxGw6C6C1o+a4RDdjWmPJP8B9z8HlpdCvGv7f5W0srq
SPH+ELzquyBV1mmu7ZELml2KAPEbFDwnRYnnsJ2RtTBkiAlwFFIpJrOBxq/GFTFN
v3vvXN7WlVTYKquKutLIj8d9gTg8RIKw0CLvuqXczBbYYLI+f9I2OVd6HWpEUs0W
5TdRLR4QZ8dgAoJsEYRmk/Iqtmn4C/EmGA1q6iBBIxN9hDH0dF4QXXnDsbOzjxNe
8xypwl+ss978mb+neUeKu6j+zKNMGdlYk4+uZEQXfJq05PYbyF9U6BcWRXM7Kch2
2fbLr8EaD1xhAfyv31f9U415TFta263S16kdHAjixTKrSyDV2rLfQOuXdGz+OitA
0dRv58orG899piDVzaNDam/9HWIhruyMj3gSuwQuT3cs3PjkqR6gbYUg8OFRPkg7
OQb5yQDlr2hYU+zgZscPnA==
`protect END_PROTECTED
