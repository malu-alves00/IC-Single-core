`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mcaTsncxib/wr0wD1nfC60nSvdvd5sFGfGilJkFJ+JekYVkESeyeWPS0NkDz/sbL
prOIaXLyTQDdTl/SdacxZsvKrpHmpg5GiKx053kSdjYXvgP8Su58LQIbOAM8bfDI
07fQbQ2PbXz6vVvXazGAt7hIfqtUSMuQ/2l6N6xDC368OoDVhRgWULNQR10WHgaH
1fvzH4m9ycGh7SDeEgWoja8YQcaDnuquh4mXHG2KD5wydORO3RH3+wg3ORu+Km9o
ETNZicsyXUthu9RUcDg/CbSjyWi7s7pbpFAwKvW/rF6UF4JOqYk4AQjci4SRyo7g
VoytuGRF3T4INHyBfD8IpE4OYneueol6StEnL6F+Edho7zasA81evB1htvQwfKbL
Nd+F7ydyVLIaqw7Usbn6+284hXqTbtpWYx23AJt0srxl0tMxZK7ZOILWujZZ5nmi
Mc/C+UnuUzl4elb79zOu4o9t0tW1C+vTtMnxOL5UEh9nATvILRwixXBk255UurpJ
xeKBXyVfpatc9GbYvTm+grItTr2FIGzyVzDjIQ+mcXqYUeFv6CTFLIJF7ONJgf30
SXhrUP9MHlltVEYLGpUcoQNi2AWhxrIPZGELCdL8kNNhNWkjEkssLTK3/vpRcrHn
6+UM1zVNcFIF4EpP8axkhGcLcbv7EoEE39jqpGXNaoy0hPJ7a9mIanOsZBBsJGon
fA2fxUO1HkRM435R2lL6pP81mCx6ozUX0zwKVjmfhzL8a425/XgNiJv1h/9UAQ0y
S2QOLVpoXWfRsqiSqshTzNUDQorNla0N5cVbyagQ+jF8F1dYh2t0Kzfw2PeLwnNz
b/0iIR2CKIb25p8CUmDwQx+O/rE2h7aSijVxEV9Wm2nfYuQrKlwhSQlOTKNFabR3
V2dm3Qa5EhovIb1RQvClDk5E7jY4PrzPHIqgwAFr9BJUwi5s0QFeUPXcULtDorzn
s0furAKS5X+d/oSp+rofVsWcIMqDqE5hSTxSFoUkuJMQ8wpF3LyQhUA4J/aV69bW
qKFYVKU8auGSOeN9z0EUS88slKNCfX8Gx3k6CELjyjuieFfA77dafToSJrfe7Rmr
G7UvsDI8EmR+GBaCi0FmOQGO5qQ9N8bYas6RazQo9eWeB5gWGzMoRXrXtTN9My6B
0RL/MgJHM/7UlpqJrdbY+QOHKJPBjMRtB083DGaykvGMq0+ofsCQbRHrRX3zFNH0
llzowzQl4wRH9picSHKnSf4noNfgokaJT4FfL08LiwbTMHGKSMi9KpDn7GKv9e2j
HqCas8nMVjqGfoypt5pRJFP/J/Q3NMe6Ky4Q8y/QS7oeEwsfVEURrphz4QrCNDuS
Bv64gtiszMVouGEP/LUpPpCkP3/o9zDFBNUidfIsKIEiHf9fhl0YqmQ3jl1n3Ger
SycjzHytm3keyONkUGu8gld4uehXCiBUvxJhSeiZIsYM05q50v5dymCygWQgDupP
le5wqxIiDm6ZnTxuWcuQTSk2MszUeZ3UdTf2hDLsJzscu9WEI8cT1kEX6owWO1Sm
yE4WQiQUoM1tM1DNI4dTV4dCdPWkTBRSwA9eBrs+NCdjAfQCD+bxoMz8gSDuNnt6
szuNPZa3CGjj56F3s4nXWei9plV/5j5UGIxaOWmIHfc4ViLKW7PSlQmb5vBXgvFh
SvWJdeaf7QX5970zbMVk5wpRHTXtNaIoycH9/tYUdncS0uGSnA6tu1NMzPjdR/XK
vr+vuI4n30cE0iCaYWyejtUd/ywmNJZjUSKDjZjT4EtNE7DpbLZVaZRwyBB7VVl9
eq11P6yHZ8aTuocmajmGLaxfcQjMp6xPAoxoMD2d6oQ3e+xF5okEAVy2hgR6rVPC
ZLgnkJRZXivAfNpV3QkxcaBdmRzUaSK7ocT3CS+Qq63E3ZZ7g+MHyGPJ/pS2heap
K5Y0K5iXxu4YjX9/aFa4zasD8GMVtpU3YusURowmAawzg/Ck7ySbKVzRaAwn3IFQ
duiCXfkoNEGXLIJxxEG0fiDkKbAMQs89FXl0iw61wnd7UZxXEBxpdMeGITWx+LLL
6ztTHL3YWIdiUkGLs2NjpFLGzf+SPeLW+YXFhQ6+Y0GIsH5f6Q8R/Ibd9dW3Gnvz
umKxyEROuoMd/mOCKKdvrnaXlduuLirps832y8fO+O5Yy8Fckrem3hifq3ttrVl6
PpMpYGax3mqB/tNGETvTbvUQFhnT/cgRUcWCidnIhUIM3HW2Vq0+Fy4B3Bz+eti6
7cQ3aAWv5+K9u8yp9XKl0bhX01TpZlfdXoyYeDoJnw/BNlEccolwPbec/UcEYKbC
AdY+keGQGUbCw1ZKpAViqjYjItU1X89pya99E5L7jbEu9zeQt3ovRGkJMbz4HgMU
nms662ehKdy5QinJIpRyiJhVD2np9yaxsBc/LJaGWT953+l7iczslFBCE6mZ7j2d
OIJ9UDAG48Uy1OMZgtUtsX4Vb13vIsGE7dLf3envBBKphY3c0TYJhqnS6mznh77i
XevgeqhZrGZMA7t2jh3Qzd0h9dkB/0W2/yGIqxZ3ubbuQgNtl1aNBVhkCzTUUqkc
NQghr9THvyN1i4NZY2NHG4Ku0gnvE3W1cWEFNMFC90tugpZ7JPk7uvqB6YhTdwCS
mvUJYBAHjmTHQ5XXl1VL88ZmDeT+gqwHyEC+N8yA2FHNLKxme4bbrNUyHf9madlD
aVm6tI6aU/nj969UgMZslPjk8VvPD6MOkBWbshvfRYvu9ZRb2VbTv/CzDn8dAwKm
O4+b32lB5NyY/6MltxIWGPzPlR2GbJivhtYcixrYLIozLBpt88hNOQ9m0chHc1Tv
QaJM62xvSfClLyQdHGM79SdIxsispQ2wAp4Tvk3WvU3wneamuDUKtbH3aU9cJQ7l
ruXXsmh/9vxsCNfupSIKclTdXo9GfpPzVhHbvG7dfNY3FoSsoYS4Fm9EWqKRSrC0
frwHSE8chUTb+XUQMKIE54aV73WHk5iA9jZ1FYf//i0CEoxvRjdIW+SpM0Z5PGG7
S5DS9XnvKq70nOyHr148QENFWRPmSSnKg9LuOu2UcjDrRnxR1UaujIbMHGRul9jk
0kWNQrDiNPt1QHEUAo1ozgO8xUUrGDLgIj3/qs0yrd386L8STj5KnDsPaomSjkkc
NDoEOFPv8BCJzSw1VUGGYlnIMcoHvpIY3JbTYvGs0QyS8ujGxPPwDkNAudFUB+Np
8blYmCEmYn2XiTeTYffj6uI6fZI3Cfa8K+Ghh6N7NiNjKqkroz96ztk+CNocKkKk
YA+v98gL10ktxtYhy4BU5xiavwL7q6PmM1Keaet+/9cckAyg+OVmIt01hrdw6hzz
dmFiYHRrPq/D8bci7rUUQ+lW7xhflBnim5Sl+MPR5YRKnqv59ogr2JqMmstLUsuz
iSqxJh+bK3Fjs9ZgJzGw7RD20gCATltaThJSGIIeTrNrqBngKo2/gAEWObZkUGiP
4U5Q9wGO+MqDFQou+ohr+kTolzM/iYXhIq3rLT39HujMR86vNs+ZdzlWnMkZkNKa
in6ijw76TA8ML1HbZ1A9OmU7doxvCjaFsfyCTWZIzqRuMxQvBjeY7jZlJWgGQj56
S3OfW8GhnY+mmM7l9MlEDg7CTGmWRgpOmG4fsRutBQFQUKAX/k+9SIiDUCcCxWqu
ZFZYocQx44j06wbEBEKkCckGOUdVo+jQhhObM3ibBpEdP+588vkYtuCZ3PdZTY2k
Cz6bKin+YWEdsqUIZVHOeZoA1zgokaKRMgU1otKLUERdNrn2AJHCNHt0eCi9rKNa
4mcazurWTHc7x/tr77FJIORSAaS8BmrkAA036CeHzqe3QyALleDsy/nwaRq6VcQb
TKgzOv4LM6m+0GCpouyiHY3VlsrLo+4/pKGhLqPo59O3PtYrKM3a8FsEpXIJHxrx
MepxaptbvicY8URkUOeZ6M5hQeI/OGbMvAU5pmKWV2CAPIZJp/8LJQGT9WY4SW29
k3B8v7JQhDWkbjO3RSxliNyu2DXYITYoYaexCBom4juHJfaGr2qrOc7Gt9GQvnnC
oTEraPb6giAJn/ghmJ+j1NhTQ2Hsr3eVTU5IJ3qHPdoIDUjlppJdfIqf1Nk7DUfZ
Vo4xoMVVehJOn5mpgvgKUYI1EbD8myjbi0C1EM6uW5xcp9MAYc1pYXDFTIeGT9gF
L2rkgcHAIfrndVR5qUmGx1QowroFQhqZY9ZCwVNsg+P8VFtlIzEuUvyl1vFsANal
dRPgRHwCxgkXP/mMYnQOykc8vM3UidmI6C87kyQbwAJHm9+o0KReLCqGet+mSlfX
mu8LXo3hRc16Gjjrwk2p03It88qQK2tlRvOkNO4vFNYFx3ZZ9TygJQuV80+yaB7e
XtcrrEl9AF9dOREY3aiMOBhvn50iMgNxfHSKcNrvjqov5RKPnsGQHwc/Atoic/cT
2EYa47CbK1stiJKXBbBfpqQ4/lReIzYXPFZGqRwjBZj2zP53dwDdx5WeoJmjEA9x
7wBW9qxfRnhKbR9j+GGTlyfH0A2mILxnasA2aX/+0mCTRnPZmM7gY3xBJjskJnfz
CH1u0jpro4OdXKsu9LHuAHwDRAeLWUlIYmro8jdpnRPVJ/s/yBgwNE5zhyEFRJ3n
Y8eVSSRC0h9F7/Mq+kY4I7mNk75KD22pgmJnYg9oGLzl4Il35oVP/Na/5+qIPrlA
HituKq3tW4tDbd+29tv9fL+MZ3DDJcatDmm5MMU4S4pToNZzFWvGFdGwaQytaD/l
I4Mwm5NB/pnlPA6NggQIl07GF5hY55bCLb8Ej7YP0RvzSll0qdhFtoIvWsbpZf2Y
e8YorojCNtUEvz5qBOQiHfO9f9QDbSKdj7TX4lUOGTEJ7eanB+3AyrUaOxST/2SR
uuYLoa6ci2cD2Q8eIyY+vyqvNGWEB1WjvdUpY+8wjWYcR6ZM2Q0MbG9LfyYUvI3d
zqIXAxhvciZhLTDZvQToXbufq7Ll362E7NK2Op2Iy8Dl0dngFteQ38tJLQP9Ijra
V0gmcC8behsgkhBBCad2lKZs4pmZ4mj8O5SH5KTSZd2OVT+Rghx4AIFP5k3mM6bY
dRHdJg0+USAafKeTCyEG2OVTNae9PKkKk7h5qlhg3WGgJKxb16V5gvCBpYpQ8aYt
LHJrrCvehaAP+r/xBVxkUlKnCunHjjzScrFThFjbiaSpKtDLv+RMkgihP/LEAPTm
Wi6342G/HdWmEhnPriGecWhg6PaI9x4eCgeHcc+YaRqLnsF5pTkAR7wFQnOwN9iL
5IYnRPYfTSJyIxb6JDR96RI2X1tdmfmKRa6v4/Pvlm2ah8+0rr6lBNIRpKcj/ils
nwJMaDIsTijHwZB2DeYw61WT5NVzMoigX0n7mw70KMtd8C4wk8Mwof/QuSSO0BAQ
5/zQZY207t0KwjDTlkniCNTCUiP5kd3PEAP/eRV9qg+D9UdNhqDh03Dgn+Fc/4Po
U9hr7udsJHR/wDrBPqszNOwqGke62s+7yglr4ZioEFZQGXzv7drtdL60bb6ad5Jm
s7NEajLxf1jsEuX3Mc/A9sWn48jJiave410eboQO6qkwloGfZ747NtW6irwKTAtl
YqKRO6xdUhesVxuIGWjzP3MGHTaH4Zq4hJYGuZ2efgCA26JMizKA1d7D2B+0adFE
83UrqEV92wZ8KoL2PZ+rY71cPUwwM/7ryhupOFmFyfxlKXfZ2V2/cWUXrkk67nwN
TevXgvCzPK6nA50i+49rs8a2Krt7DGSBmRaSdhF/Y3nBTQ+kk3Y/H9tlYbPQaXh7
AZmFGYJTTfvq8dyEb5dD/M7Ck1n6su2RFXAzWnocGq3Dxy92hdFTWeFqafjgG3y6
tFKGIrqUqmxF89sJOdxUC6Uw18Et0/dGklwivzKRPk1FaH0G2F5xKVYW9ucMtHD/
GT/kLRCSPAO5FT8FA76RZ4Db61U4fAWgFzK/2OD/bmUOruO0/wMvOI83Uj/2bbwz
VaDsGVMX7yh1/kwRpT7I6QM2IrLs1KOeKqGZHhYNmqF8A3cfnZ0G85TROKmzkg3K
dCxtkiGdb71vfoF3YwYDH7LNc3rXgGDTv12tplvqMg6edjzrqMcTHnnxBxboIwsM
mYZ7CTa6LjBArKStxoy1lkXD/ZL/FlWV3je4MaDA+9qomp3PzC2HA8pNcqMYhJoL
jaqrQq64JbwoEtA6SOYMlFaNr/pj78FqfSiI96/9uft84P94nMAYXNBXcGXtCCF6
Q4bpDIax5FUkj8ntHR9YYiXS7cqyRX+OOm8lmHrzONNBga9yF+MAGgpGWeeH+wng
amCN2EwAR5iiZm5MD8iVDyc32zYmxey4ZthdrS4SInDn3oXNbHXDlItCPWHb6ti9
OMZgnMC1YpqkDErhOp4V1feJ0GU7El76JE/An/ChCZoiu1f68IqO9MG7HiHYdfx7
oSzMFwt7NKn5T5LZ2DR/pQ==
`protect END_PROTECTED
