`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bQvoT7V2fcOO/NxBXWokdZSkPZaHBqrUDLF4yaqPp4l5ugE5Fsi6uaFxeLNOnWBD
rR+uk3/pyKmElq4DTkcaXqxtkgFamr46dtyVLLxefHfnYATBRQDE97upKZlEjBme
+diozm9fLBb3007lKz0iu+HhPIDVV+3BDzePuxW6vwc8Iw24Jj82DqjtQL4ACOHy
E2Ji+fQIQr0AYH8eEcTUDi1GD7bL5iE/mxEIze/1HrzP3jefUadDfbdOV1zLGRTr
lwtNNENfsSoL9KKdB96xMoKEHk07cufCdYKdiGCFjLw5lFVFqYk7tRSX7P4FhHJm
GZxNunvVkLj8mFxdUUwwhrL0P5+DMB5vlH31XOgxrfUSp4sMH5e6qcPmtAHk3f5I
7lCrKgKLuY4qj9W0uT31oled2IjnsKgcA8pvWf8DE+T3qKEzijXotqHCTzGEur+k
u67z14uvNdPzmkJ4ijJqk1eP6uqLCmB4GyG4Y4487D0FA1wmM9vHuhcJb2n52wTc
2Ez/+hA486omoYTX2d4ElWbFBfMhWY02ZIG6euFBQO0=
`protect END_PROTECTED
