`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jYJLxV0m7V6D+Ire6X2Sz312KLUxM3mxfPNCLgg5EjOztD2gPzN8VfRChslGE3aS
uSoYKaf4meLf7bkCOUP7+exgt1TBNCYQolC3WPsC4rqqsUWLDK9rtW2Y9U7W9/KG
V6vD4badZr3+KTkfZmC2PXDIi16BzWRhbQS5jin0ZGORRWKoM1GBg/Ip4StQtwJv
91zssSeIm/VKIBKmMdHYMgkokK1ZgBvVWpXy+A5txsBQmSiXV0b6E6AfCUQ+ZUW6
2Spvtngtzp/nxWYxXrubS03NKVhp4L9bqLGZ4ZpI28TT5pGWP8vaiWPsYSJyckX0
3whg9taGidaxig4+6N8+ZVqlMLocHEQTfHcwD9pvjv9F7a7R/ykIeqsAHCVnFvp5
5tq0CZO2nBiEwIorTgU9BIBTMnPVXQAJp1sbwSdfoanveUbwuNkdxpGKt77ITwJR
43yKhHwK8tqOjb7BzBcQEL3qF13hqKpoAuEUMGeo+GSsEpBns+AkSun3YI8gFNBy
ofcWI6Tgybx/bYDjQ2WKZwPt0KuZ0LtNcl0ZpAlllxsGRqP4F85/QR0yPsCjEZQj
OtbU8WYJmKaQQd3XIv+MYCMOH9fYnXMGuK5pdTI9DH/1EmdRX3nfTRT0eUEpayxJ
DOHLDTC5FcktTbpPSwjNbpZNS6m50EHjN6Bz7L5lQ3Oj2rrCVW7gTakMaZi3GKjD
B0ZLOjElUkC0d4TXMgZt4XShn/zgP3JoqVumyKh7gPvV0AodUB2jOLNFpxLY24PZ
dYqmEXT998mQdWRjRE3z0uZCJLtJX/HipeTQ9/PwtGrZaJBdxoI4cBiCMzs5+07V
5yYebZ3k/EsYBXTubt54QNnsQWFlSR9fOOWKigDTMhQEIFhgBUypvykQ0biXS+Th
zVlVt6nAkQRsALJfZ65OsvR/IRNCF2cX6B25+giMnOwtvwnc+U9CjID+JwQGrnnu
wKWbT6n6o1YPfoSfrR/QGFw7YYdLuaJ/zoFUNgupriJsmaE3I8OuwJx6BOC9aif4
XT0eHL7GsAUGUo1WuE0N5VQxszQLh35Qn8vq+uXeAxfFt0wa1zx9IhC7BbDkgFNA
vtTSegMSHKZFEwhQ5kO0hcDswUxnM+Dn9Lz/glEAgV4ry5HlPfNGdc5DQhDkulaw
0GXcI4AW3VNMnc0ohCGhakny5gq3G0nTohmHm/xX3LtMiGqiV3RTLeT9xuLLoKgF
wA3QPUDPfre8iUeHJQEIs5kHvfWkvnya4DdHbpbqx4UlcULfKMNclOkvwmGy183V
UZQjhsUxwqPtmdSKI8KZe+p5Ab21r8hdqRSrj8Udg2KWM4Z/Pq73cDiGvt6PqJnT
ROvk11YqlMfG4JghwV8H8adaHpnxDpJ+BubTpLpDQ+NTBvRAA3W4Tfzs3OfEjGSD
3nGABDo0JI3OUOr9UbIG5ky73hIoGy7bsFPaH+iBdp2IlkKTEhp5zn9Or1ZxzUZq
zKu1ogxIAjm1wxk1b5LWSMptTlHCegX8tjd2woBTE3PSZbipCsAkrnawneKMSZ1m
EsnYH5ytBJP3lR2ZRb86zRoK/MY+VCguaXrzrcaTaL69YDdVwpMee3vPkFiVJH6w
Mf7wapjWD3i7WIvSugabrO+sslIpjSNcGMCqsWVNnzJdTdtWGEOcGJXfW9XQtxTI
6BlsPtK6ek24zCetwBB+2CyBeco3DSHb474BRa6M0fanPkmpLFSbNSoLH+/qfLi7
5vEzLB/Zr06DI5CyebxLgIQW7KiOtxIQ7NcyXcj/sp654KRTZkHDHFNPYUdlKQNV
M6kHPB5F26u8qPCrFsje4XnCxJZEbT2VtR//3XBIhb0YE+ICoMe6NEo8+EOVph3K
UT8w210YpNZ3dn2+BSRtI3nkWX8jSuTSH6/FMdtPnrmx8SPu0R7UKZKBP21C83mp
h52urEzGZFlA9ZxX40hVKGZUtBw9Jq0L7Ds25wvkWN39iRxiRmZlPklnBXcWKthR
G09t8POEfJVXFxiZO/v7SxJVI1DX9HWnxWdpFZ7Jx8hkw6HiTmNnUGhlc3Ip77zV
8ErizIykNU17Kh9LZyZTD7vQb3AcyRhDICdSKK/Ch+eAPqso59WySWcBl0UvDHVr
yR33OWSya3ZSqOn0BJZ/1HE2Vw9tswQJz+OoU8eeQcKSP3yb1mv8mmE3H5bTelT4
qW9ra4LsFljL01TcqPbHMiwKOuM7JFK6/UDw98Dp1Jvgj0V+sCF3Lr13hDhS9vA8
eqtJ/VG68IQPSqxDHyFZYRcgGS7dEQd8fE/CxuKJ39TVGl2QwNLwQ1xv8fBLfWNs
KlWqoZUcqmmf3D0hLzQgKYLHUrWOdm1P3a9oXkcqr0YdYuZBWlX3Xn7XHTKAPTDR
raMvgx9Xp5E4QTMrjLodC/3DduyWNbaeCjJk+wvI+Xe+yV5VkMjPnEFYyVaaLkpE
xCW2yq5B99GXJCSJFSB2+mziPGJ+BYRFdnSYSYA5f3B118RrKQPcB9cUgCszZuXM
65UAA1KYFtSJk+F/0b4gbk9yQMi+1XO08dsNC3DL2YWOhNZFtf23B4SOK78O3yaA
I+IXISGumlEUIto6NZM/Gw==
`protect END_PROTECTED
