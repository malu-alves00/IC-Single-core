`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yUBimHZ90irBaPbR5BFwXhjim/GZ4+DDe6WGzeHJdCNDOXSmWaz5YMOKlIwGPaUa
8xtikkkyycgi+3H3EmrH1bWwZQl/qSKA6oIf96jBc1SxWR4ieSOxaMlvUf9ZpJyb
kUZBZH5nyptJv1T8cuIlyJBeHHrVFUEcOTSij7uCGnhUZdIjehtYQK6hHMVCXjki
qAartl+EhTFaJEsSOC0K1aoG94eEGkgh0VnOOh3QMryxVJpyUWCSSv8WX1zlVSUN
ZJLseDqG95haaj0YIQtBkMVQq446Gd9+Nx/cxFbNW2x0ghs+CbQG91I/taGSXq2Z
MnsPKA98JSb8n5ZhkM7oz9MhliGTsFtYaD1y6EuRp5tzgr9pUGGcj7Arn28nm7DE
mjK7uJn5zjGGCBqKeMKH7TVfOUDRMJRMoTDOi6abW/1QRddrEZvi8RzEYuVLRI3f
/laRbDBbBAQayW8gUuN+QouFcYHuxggLxAIEDzo1mdaUjobFh0nWQgmXWtUe+kvp
nBTKJCcp0W3w8qkSJuATElTYFVCo4XXeIJdWMwiQDoUXgYd8A2i2+dSmGtp0Psd0
B++99afyNvRsYib4KBWALd2YR1kNjdqwfWZXJ+nTh6iGw/23X8SKpN+pZD+isOet
YMPhcU/vthDlh4IALl1Sp6blaEot84+lAnrjfFX1QOQs0sh4jUNCgCUBhO++khBR
fx68JjppsgNCJDGd5Wg9ZHlVwJjtnhsLxkeY34a2n6CAoicDHITRB4QnK1MZYRSF
vypG1/DLJ77+LW+ibhXiTSgW2fibihDunMJWcnNWs3O5/o5Sr+qyn34IhyGTq8MM
ysWR/WmMcxQvoP/kSK+7eY6oisy1au6dIn36ZWq7Wg2WE9vw5HZwKPqGjzAmrJar
iMDEbefzjE2zox/hSNwGv/h7Jz0/rAT7XOsMSVI+WlgLd3sWdHgyomKflDovSIZq
YzfHQBKk0mSbcapfeAVZCwVsN2uyzGAC7CiISH07htOac7XUiu7ml0hK96j8Taop
idV2WZ01z0LHitrOiadn6t+PE8/zzAnpsR/PgnEXvBXtghhTrGJX08YcFCOyBpyU
sp2Unygus+LXS4Wq8XsayV5tn38L9CnrKCiimZ4KpjpNfMd7f1OImgbso0Gb4jPt
wXkOgnoZ8lktoFkC+kdMhkCVxLLbudzAv05blihb63AWNroUjFQ3JwFcV4jsoWz9
3LVCmqyD/lvuXfYk2EGaSYYz42gLLwYW4QNbLT/sTQv8IGFxx82VeugKvfcY7ylF
`protect END_PROTECTED
