`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5DiYb+D0NuHanmlJvppr28D7+K7/JkRQkboT2HHOyTc9/QLVw9ShWcHdaGSkfu+q
duGCflkj6kHTxh06fO2j/i/GmZvWULcw7IQcajEHw6/bQTnfT86No3KI3tEpBhEG
n2Wr8ox/5v5dNN6Mt62GM3HbErouRhCaqLyX9YY/Qt3WfI0yTQUxohEwrRNnvZQo
OFHjv5E6O66wlWuZy5jtERUdq68xqDnvFAjOkj/5BXZvHNAMGO/DbrbUIfX5YGYF
Anu0QYQhMQ5yl1SvH17TYSuPYwgCV+lpk9Q/G0MBWv0YOJQ8xviL8+b3k5l4Gc3w
uQWB7UNKcP4ZGm+1Qs9rZAjreYmQB+WrVkX61g0LtKUEr/cQLgqWv4Hu4iqeqhA5
WMhUALDoQn7dD/dkCAsHLK5LZjRFFNqaa3VNmopRT+4GaXdGJ6u3P7Pee1Gjs3Cj
/LIZ2SKKa25LaRBGUgsfZFk8T8dnnXRaKKR8C9cCUAHo5c/szP/K/LNxLfUJLpb1
S+5WXWXCWwYJJUpugHH9YJxYaPa62gyygV/wMvbFlui7YOY0fjR+0hTfAgSks+pi
aoWE5bCt0uOaHc2DohltxAWWmXgVvxiT/2/UrN3GmrKAk3puyn73zLzigg/6bCyJ
FhbzeLwli9ZMC9Sp2MYPR7hjr7uyUWTavdLHb0JGXVz1rIaYt2tmfEKCjb5CSuVr
ywsIlGrfioCTvby87iC5WMUf0xFDbAvJx1WCKMrh8iJEW7eEYj3xMNv2KW4r3U3s
VzfHHDhYV9jfKEROscKwVa7Sj7L1Hs+nidVDmvGa6oq2kLCiRfn839QSEs47eo2T
tIIPEEnL1u8sKSA7dsy85MdfjbJenVQVCswV4kJYCwyHDetOWEnja2P9aadRenn1
/zTHqi9rnKYRW2QNk3orkwIDWddK8f0BoXaUthuR9mFp1b1Sa7AphN2SatRQI3BA
T4UlfwllCbiQk6bhrrAzFUSDh438yR579YqDWXS8pTpPBSQelEWuWHKFbXBHNTdr
5dmfiruqUeHaATc4ojmQbevcEJVZ4i90Jbzbb0ndnWehO8wsZ+Ipzo/moYsgdubo
FiHBwHsglPD7SmGmqa2LNXCBSNHF5K+85BduJCDhD3r1DPciHpVyk4D1tMoJMr1y
Q8xFfJO6vk8HOt/Bt5pGbw==
`protect END_PROTECTED
