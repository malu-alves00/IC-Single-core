`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2mWTOd3ZsoNlBUe/XgrLrImsjpYeLuCGdwL3gN2B6nJLC34ahhwmW5CrTgVgMypk
6NKIGSHc+TIz1qzl3lbqImzwIpW8VEmGYr9vN2nH7rEb4IzxVjk8gjS64oD5mpu6
GZ9ytOyoHbai4EHQS3wG+YX3YK+NxwoBJnvJw55PCVvP/AxDmePItPW5ReMypFzH
r+ERxxZes+Z4iSUe1D7raUaWiCe2MgGOo7jXrtHct07UBAhlsbfm934+VIvz50Lb
TX76z7WMrkyH+e/k4G4IdDqphkrDb2BqhqU4g+4iE4mDMIsgHT4dcZF4NGRKsI2f
m3yKMrf1GiMP5bFBZ3s8SD/1YS5ia9rHAJB8i1liZzUQYGLWv3fkl9w+mU+HxKgA
SLEbccOaIvsgUbJwd1Ckl9JKCIXqypGPaK4QOqHdqZG6CVApa541EgKDT10TWMxr
oQkXSPXYXLBUIUfAUJXXyLwFipbY0yNwR16saySMEjQfYZBoWYW8zZJzMiCG5XDM
if2/yc0FGdOJlo6UGf3atBkBKxXdWU3/6UQNF8OcxjXZE1LMRSo1HL3sZxMLWKk2
pAQiW7REsyCZUk9VNLEWtCWzq5Azepec/CbE/BQIkQg6UpX2Ghj8BWlDHW8AlWcL
N4UcbxjPwgI6cj0PFUSGzWkUpPZGyIaIAJCh6V/U7GeXfhJC2W2OCOg6KoL8TYrG
FxSKcnocc5nnlnrFGdy9LzVtySeYVkKAE8V3mBYcKg6LlWOcsTaTXH3ZqRnnSIeb
bDeCr9tC0s+B1wAvP83EvGXYswvoVIqM8gkOj9+PmP7Ho3vuNTO9HqG6m6FqkIfy
N/uFdncifUCqlv+2AwnJBRRYv/27IIqIn7DDFlLR1hWQTwQTwykhE5Z+c4TPZ2MX
Bool2qXOJ8cfEzIVul9veDVhE+m4iYQtgjJis4yla5ihWlIndpSURVInbgfvJsNb
UW8+kpwV3eeLDImEp4ElrYsKR2cn5rKpDMgpQYsqPBlPbfJt4Ky+FPE9NK/F9w4s
fINhmJs110JnROcMtEAcnHsQ7w0T3uMNirO8DltKzwYlcOsX4g05eN77my02J7R2
pr6IzZ4PaGgt3j1zCAOeGFLgHbPBKLuXEGGfJ8OgSLT3xGx8weBHmDxVlvXWy4GM
uwqdJcxKi5mDQOQVjOww/UTdNjklAB0dINyjG/fT5H9d+eqfTONXwFIjrRIJOEuL
lSS4QyfslnTeQiXAFP4chVrPETcmsP7TU7tqZLJXjd0EGy63sNMIJoYan0MjVUUF
wBtZRu37ppqfKi5/mt+K9la8yziS8oeCEc6xpEgL1CYEYQVwOH574n1/new5NFm1
XBLMFmhJJyXrLfRTV8UIkv3t5zFlkIQ3MhObtXnskGR/ozBxBSSpAgHry5vy2JPK
bGuffQ1XoDdHQ6L1wsznuU/WdNLynYQPIuT2bkYp5sLCjeyvd5LnAmvHRqZX3+Yu
AyLTCJfttA/QUwwUZTYJTnIwZSgD0SHniYljmlgqc3CUZl+RSTCTqowRxmxD8yZk
T1Kl6o+KMQC7hvivbOink1UU6AlefYo9LLSxV+KJOWxyYQd2sEoYJsD2fOMOOmL9
38shEOMdC6U+zQXU2D0oCsJReIVHjbc5LIWRzGvXFD0ElC9c97QTxt0U/ThjXIBu
4Dvi61ZdKbXxWL8OMnvjfh+qFoAU5EFnxqknovGl1ZWzWBALpRXuksNGmmLBpTYv
XGTD1+L02/y8fmGLeter8CKjzrrTt5c6k5O/rja+BUbGPJAEoqkzyB2W/kCuAeDV
lEbmu6/cua98wRkGkOuW1pUjl2Y0MIcmfvaHnK6vJENHoBu+ffoowpLmfeHci0MI
e+7gUTGsKAZY/w6xJRAJDd1Kx/8ICay4FU3im8CvOMjk4wFEMahrTIi/RhBIBMsb
v4ozSeaNRAIZn0j4WVELZMG1HqvN4aIAcZvloSq7JvPuNGkIdV24xBUfP1j6Eq04
VAEd1hdxZjmXfIyPH19eaKHcirrugDruragLoEi9Q6E+kiiHKGVzgQ7Sa+lMcjKR
wVoGFSMSMnahuxzVq7+79EREp1ZcqVRk60EEz99hmS+T3LFVxqhhW4GNAxW/UMai
Bq1jhovRnY8HPZ2dl0hKu40dfJIEe9twjOm3wo1XZqDRYxSsUazeFPTi7FV3+YIy
Wn5qHSQa5wxl25Mik3ESohvuOGqIcZkepGbHZtZfUsnnF+pqn+vUJ98U1LKsCNvT
A6uH6FuaUYADW1xziIuspTPlu+2TgTSFjJi66/rWvFbKMAljvCK5/w7wQWLedZTB
PII0pT6WhZNSf5hNRELVtzOu0yp/xJJTnWByjE5nTleHN2+CLbMYyZNc2wrdiMYt
XMrPRZFxYV9R+/bcSsj9Fo0Oovniat3qJKqwOOdnGHcOJVQf9BD5kL2wWOYL8h+a
5l9PrDocdaHfN/wYE05FwdAScgugC6GqPLWJMvsU1vSrlfTRefC/YvwHX09K796F
B3W4uX3U00XgpCbNj55zX3CqpWtRNVbA25CZlLnK30XHORPYD8W/kLnBaSYqY3CR
skCx5wevGil6WK7vN4URTHIwl33T2O29s82PrurcizSVeFHDGz6wAQMsu/6OKO05
tvgor766Q0IHoEyVWP4y/w8mPnJTVZWNGYgWN2OEuQ4DNCdS6K2jRs0f0hh83Os4
FTw0WnbCpvF6Mc7S1XdOKR3ysNwWzA74JaxG4HSj/SiEljGhXmzhcl/Gcr1dvJjh
ZiOl+JCoVcWxcVYl5puD/9VtPdUmihV1qa9BQ/br3MIFyyfniJSrvXO+HYOPVRAR
3wtqr5HHJwQKRS5YgkJmsJ2RgjfqYq3V/LEKu7wsvLs9vgC/t9smDE/MYv556Ozb
Bz71RQBd6sIqAJ4LSU5CEAXj0me2RfMY35hkVyZsLO03xHxQq2imykCRlm8qn0kL
JgjeJulWGGy3tc+9xbHu/G3zJcN1IStNmLmi6y0amTWevp7fA/SQs9I9MosoEnaC
87fg2ZxbV0jtfRkqmK5BFUbR1UnZxLpAOLTvk0SV6YfZnMri89DEvXF+TEPEn+8f
C02wVCfGYe9yuNK/a9c+yWIwvxCL52bEp8FAje/p+PSKYp00V5IrtiVgmubWhEu4
XWZ8IQcYwVA5MVcMjynvOlEm7SixAUI3SMf7eWAURGAakbXWLGL4QtOn7BK+u2F/
qWIgqNnfnnYFF6aOZK0A8fY1EwdQQE2ExK3fSBejA/8dqEtG0VMbBRFHWVE5U1j8
uz28La5lMlsW9iAIEBAoerwqoZztjm+h9slRjjJJVmlWWk4aCvchU0bxkj7h/p2R
NhUikrFXsENMvWv4pRgV3uCSn3nSNdo4sm9arHTJhb9+LPzEZenqarBbwKXsLMPS
PzCYDwmK0FX/BATLON9TOZop0KeXsIzsizi4/ZRlcPYETFCTt2KxXJfZBRzdDpHN
Xt0Uje0qrya9UIeupfpk2irUzBDb7u0QfJBfWn+VIaMB9zJpZzt27rwusGdfOI6U
bCXj3mbg0De4pCfC7w1aEw6oTrBTrczwORNhajJ2QRoOQau2Pup3ek7dtCOaBdfg
T4K4vl+a9ypdeXPThtyFbqUwJpjmrF5v3abG+85QvnIes9vHiENIYzAdd9qgeWB2
6iQ4U8Ns+6GpNBsTMRQH4GO0dCXs8IzXLoo0yC04LieVvwSZI8ssNtMolz9JXSmB
GaR/wpoIlBrhbko1lZrrjs+KL2laYswzAkKMVFHuuvgmQtlPAhwlC2cAlg1FRcqY
sXfOuIUYnkRiJVAM0jRQLsLdBXSYvQBCRFmGovGXAofsS8JoBQz658XbuSHRkG3i
KMOyOASqROVvgZO+s/GUP9b/kH9LEc4UEIN0lrq/6fe/+yffS3SZf9t0BURexn5F
pmCFCVIyh2FxZZDLbigWakywb7pRb4CKIsR75j2Cl+Wgmb737yOd+XDTudhUwS5r
4Lkz8U1j6qan2AUgp7gDWvURVRafAkFsFQLeKEqbQdY=
`protect END_PROTECTED
