`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ovRVGaVveHESztVrocnXgVBT+sSFkwgcOWORXum4GaKJEBvKBqqIIkDHY3If+UKe
yd7NLY7fF9xyJmLyvcQn42814ToVUeaHSauXIF8yQOTFGoPide7tbEg224hKx83r
tkioH2DrL3/LNRRkVqDKl0qwZCoYGNDlyZD36Kr8faD0mngN1gOlLInOqpWN33vO
A8H5R+xT2bBTYrRjAhgpaqvgsxzmtXKxdUV0DYpKwnATl6l3rrhrSnM+tVWAfoX+
CkLtbMPDP8c5SS8hwNTe73H8lPzUSf5on2YG3MPS+QUhZaIJtN+jvh21ACXxnKhm
n50hlGL/lDE0U+TN33hi+sm57nNOwhSTeNaN28xc5D1GOyaWLPSpW35n3m94PIaZ
ZosMaVjKoede2VzaSrnuydGAZLYvt482L98pdjZIe56gxXKr2+ReutNQo+9anHRy
pVFu2MxJs7pLkfv0ENy5I1wW3lLH1OKGdsYKgduXuPZxS3MKx4t5KXTM1v72nsEy
2YCz1IBfw2Z5bnhq+YCjNYKQ2MGeRpa3KjPls2q7IJk=
`protect END_PROTECTED
