`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HFpheEYJFHikDMty0pWV81R8o2dSodKPpcXBBss4+pTHKv1TIFW+3a8i0f+3Bhgq
jw/Z4xaFsBw5oKSsNk/OAw7MmHzKyLsGpQvvt3I5mWDWIEpvBdA7erPhc3UEdRYp
x5nAefQ8rED48OiZvXhE18k/BFZeau6LOWRPoFli5DsnnGdvHWfR2tu9seR3NPQk
xt6dI1JyWv7Xt/ZDBC5BWk2YrQGZtqtNM6wcONLZg89F3JI0nIs2CUwyrJs1d41x
3OFwRbCn2+Fo27cLLLDJbR8aUmFNCfzGFq0SjT0D+C37/xObnf2aPsk4zIqi+eUH
Qen5r+wVWnwPOwn7z7d25+QHs6aUPPXOSLV2S7HXk6TGF6QJTCvHzpjfBlbFK3xc
eDw897V1cxpXwpZAurMpu8B5YLhz02W+a2pprmlorpjU5F6ja8qOMUs30eU5zQ4K
LUsEPSazQ0Cq0TKbbD+ZGFrsyp8aHNTO+/oxpEOpYO5mbTfBBLu2l3GZcZciFwQH
UjqRnriAV9BlR4VK11pEed7ZZi7So/BQgH2reI5wwFKZMedbn8MagJb8PAnsJ9Yr
jLBpf2zAoCjVdsAPQPMBKht+T630n03hIcr7nCiO5eMRXxkO9vJKqg35dMn25+XN
K/qbUJ+0FIrQU4bOfDc78ZrBxOjd7mL9NctB/KHc1xIeRZwjCw9e7w61NQ4ipJjv
pc+rCh43Cg4IsMEPhCl4yQ5vj84v6mJwpoprbPQE3Z5UQPCUu1uwZ82JcsXzDIN6
rdPSGZxD+RJ0rkU2sSBruZD06hmWdIcviPb6D0tuYN/B9Grw3f0qiya3e/dBU2Il
4xgxGuneLw0RTXyZ7nRY3SWl/Jmh5z0Oi6JhHhFx/sACvigGmHpTxobI9wkv/XTo
GIy1ICLQUtfzLJfqZgJmbmQH8ZX/OvTx7/aUzadcT3sBgTn+1o+Gmjkcd70L1HQK
LwLTJTLoeMKBzOPfIu1kVW9BktxjTu4ZUVrmuK1HfdewJvAUGvZmodLsus33+xpc
riCxsM3btRNhD6wqHARQueyH7uG3x+tY8pmyD1pCj8PXa0RmTMjywB2Ddsh15gLm
KruDygvoceHqz5USZOXYyi+6D6iCoZHN21owCMb8phY14HjC9ziOzOmvMuXl1KIg
BPDmyWQVPE4PAyDNhxf1g9f1pyqD324uIoTVEWyLZF6YpmbJTQt3nsM66fd2KHXg
Nf6A0oipXG5XSjy0FgOXR94V4pYHueQOGsdsF9k+Wcq7wLuXTdk43g/qgsCCY7Jo
OryGg8n8coThTMDCTcpRe2QXt8rAWnrEJP1hlxy6wxOXIH2snDOpRJQIeJwc/+RI
47yqYwm+LdEe/gLdn0/An93xjZi/t3foJ1eUjZ+mO4pGFhos8Q/8uiXmRvMUT+io
1Z4L1B58314lvmDpJh3rJ9VpzlYQNU9f6uvjtnqEMnVvz4dpRYO/rdzFgJL55NEZ
FuVZ6Mjh0FC3503IEfzZLyDqLO/bguBG6qcZHWcajfkGSYjxypA5WEaAPqEKSlei
7VHcoVgA8RTLkkas7YwmW87S5gVqS5uXmATGuzlinoJj4g+52fDOSAWTevfLzRCj
iRVJNNwGnNMrsRAuJx9Kvkr0+OWDtEY7JNrHGUb58nEBf486Ni6Pw166qz8EKNcW
0vaJumoRaLkv+u9UcqygjC0m45sILl/Clm/OlFs6JfNk8HS+UcyQvqvbSniIdoTZ
lxRGsI+37vkbR67hFQAS18taj+G9F/qPGzOYBqdKmnvuaJMw5ZT/kTa+okjVrP0q
I6QQATUETmAfrBPEu+e7hSyvogWonxtI09zo6HHHc5awDs5C++Ewh+YEsQiejpgH
sz22AruP6RHw/W9Ryw42uBSqP/oj5Xn3IFgXUVlNkBqnST9+yPRYy+7wWDR5E2tW
/PrDI03reiziyZY4vKYoDQ==
`protect END_PROTECTED
