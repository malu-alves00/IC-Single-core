`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bl8S6/Rx3BuyDWRgStS/ZoN1crnsZrP1z8Wen+WvBzJjAp6X8Wl8XysiptcaDyS0
NEli7lkQKJ1aGtz+IAb66vY+0wEHve4XofAU4zu8ZS822MGRsNbRuHPjlE2oQMYi
Sfo/la6FTUabMHOKc8I31+w1289QCOiqKLYRu1qIjac/OQ+IcqPiDXX5gsNo2nEA
RWFHxQGeGB9hxeNcFdOxNVQ9sltM2h2AxD3kZTsIjX8Mvrbyz0A/fQYBTWy/EiK9
pjh7dndpleOHuRB1NA1ruONXM/pw6S30WPu2CyFFqVOuPyPW7y8anFDTbSTPlt85
DHyYbEhCyYsC51p3MF9Wj8Th33Pa+hncC8QW3EKGjCtab/wH7pjZPFTuo3oF69Il
H87IrRSLAV4jglfwJLUobbKBGszAuZOuILQouHmHw0AiS/+xMnfX9We5kq/6hIvp
iB4a7t40kndAaD/eI82oyLQoxp46zav4taiuu6vbvmamPasucVwb+99N1oqlT0h3
XyhQRX9BitE4L9k6ibqgP7ZiZr1pm5iA5X+J1JPeRuasb/UkoSWw1MVHkDQrE8TD
wBk84Ubib85LVWLKgbqa4BkA4dBAbMGHXLd3Wlw4qZez1Ckk3yUw4KE7VTl/U8XK
AZwc8Lbohp2Ra7tJSadFQxoqSbcwILikymndb/svR9ci1WkCBXqHs8soK5TZiCCD
8O6kxX7sx8/gYJy2qBCR0H6U5pQWJy5U0UWvNxbnzz033K3fP/MQfOTBItx50m04
66t8c9mGvJibN/qZNLVi/8L9H08Mf/4XGkTCRVwsbNDHHj94OoDDqVx4KbubrRYD
p9zrxbJmPeST11pTztUG4+E1pi6JeHrxT4E94CXyTmGMS4RGsvQk8CX8KYZfhxZP
x7MVLkvo6h/7StsOeYVxxGodyGfw8guOq5zSQX4OAbX+zVq/SNfrZ3Ohnq9O87l/
NH5/D0vXHeoEIDoPQwoF/CAH7urP3qYqHXbQvTizZSfNnJX7vrMj1EInqNv6SThh
zW+8Kr4Dqfg+KtR69A5gdQy50zUFkHs+2bRQakFH/+0TKLEh/7mP0xT3JQkCBlU4
mT/WzN+237G7yjEKJ91N+Z4SzPne3vYsuXEfDne+Dokaa8A/l8MUIfjdtfOaghaX
bbBVNMcqoLX7fc8ot4Rt98lrA2krwmIT1RB3258Umcq+/jhR7mqzHA+VFnwcbUcG
ii7pgJ+i8llzAyP5nETK3cyPssODiDeQj24Dx+8riR5Sp63W53OzdEH5+rbvpb7t
/xi3FTzmEMnV2QhWgQRHEeNtmc4WUTXdZ22fluo+FEcJya+wz12r6/86vuO9mJvB
8biUeodLNoefKlPivhRsbRAR1InKUEFl7gB7LNrVYeR6LCH/BXob6olbTFOP4x0E
C9ZBrGom/+l1LfWF69w9nD2d1lLHQIi/JgyfMoDR5Btbd/kU7qTi94ORuVr0+Upz
J4Z+N24wtt3ddtV9FbgFCsLJTx4r8KMMNcZV8v6Yf/ACInM5rtgaQfrVG3kz6AW4
VFP5VdUW2HnmM/zqALHYgUeAauQwHLbvn4xke1lPz1PpjgqVfJISZQ4UBOx0eEB4
yksltW7dJ608P09TYvBmQR7q1YtIpVytDtvPm2xbzfbrifydXkAzj9eD1x0J3qrG
YfrxygwYhS3i4AWFktGpLxvxhG4RwSmsuX6/jLjQXReE7ejyrMWbCszUCnDHZadu
EMDYrIRi/hsccnP+usb6cmSztvaPVtNB3gPE2ELnS6FXk0UOuOzXvGO41JrD3Ble
zpx/svpPkmsGkZhFMVNjTlzMiNv+buuS9AdNGAUd+BHQHfJo4k7uIkiZflKPIQjy
RRG9v+iz61WJy1dB+2cRHvaHp5Oi/JK1feFdlXey7f6LSUBMKF/5H/SY3eDHiz7x
wZiA1giznN1r+HIgKY6TB48WHZd9QZ9JQx2FcHA6f6OHaqSDUUbm0mBrqRHYjlCd
1ZN5FOtZfaIn/ccl1vsGOwLFN29qBA2O+vQ3sjFUEG8zfL+T943NwvvrTnR3Nc7E
jkSKtfm6U4Fp5hChKN2DM7scmJ5+Bv5diMbDrkmBDIc1IhrHI/RDkkUH3knuzbHb
Zjs05rWDm9oybwD6jXDedVKq8KQswbpej+EsVgtKM2xsngCP5OBnSE4fYb0/SiX1
68IznScK8nooVUuDSFA/Uu61pEBbacMY4cIaSozcuch2tVRJockCGwteUaLHIHb6
tMHRwHSC4Ql0ENg756fMC5gC3+WzJbA9hw/U75wJACRZ07AhymeuRjs/USXO5LJQ
j4wmAH1fgEoDtXa8UlaD1DOXqsjI17c+FPWlrOndPltiYDgVdKMl/7jGF/H2af4i
vGvdfN1uf2T1Dxw8TZnb0cOBKDaGuwJbmsFLKtLlztQrChBsPcTmIvnFKJpC2RYY
NH0FmOVD08y7S0G8sms5EcAEUhw4XJpzeg1/v4+v04B4Zu/gN238NrF/2PuCQuaZ
b0uRh38PaNqgfC5MWh1Qy2tm0eGLZ1TrmpwYhjNOOP1fDYtxmuO6C8C7qv7JXbwp
LOJeJ9VMzWnfwfxUJJRo7xABePTYMiOl8f0909j07/J8+r5efQycAleFuo1QWGqa
x2LwYdyUmLDQoP+fUofztmUfNVAxpzNufxDQq68r8hy6JYAimeruL7eJhn6EOyYO
6zxvNA1IljcBnds/hxvB69Y+DYq4lFVOXkueQlPNmA5J9d1Y5+EKrsfiqS4E8/Kh
g0IgQFcJs8svNID7QPofYBDPoiEUi+5Dl+7uR6MBy9djWOJ/HqRufoXQK8dWwoTz
BbXue+O+bnQt9/Ygg6Ty7NKCvQ0BnTNFWUcIJ+/zn3jZFPMYluFWeK+zBf6YxiE+
+A7LXzDYHHRfSPXxQacFjpLQx/7+I6ulq09IzgKKL2Da8R892gYc1m61P3jX/wSB
CH93fmwEwR4eoroi6YbGf/D4CJUlW/cdZD5CJ+JAl754lAU4jzazT1EJcklKquqv
w+/3WzQcYcE0v171CmbDbpU8t8QZhiBj1d0vqC2WATNFuKwWbK5PrPjIRLp4BLW6
eWhpU71pUwdKlTTL/VGcf5Up3SE+Z5HpDZt7fK0Krql19+No0kec/Ddffzjb+zLC
0PKhf6us5MDxF/N92c1fa3XlgZUwYNsipmmKSpJfk23ZDHW0n/x+Y5Yi6DKNIlgB
i9JOeTWHZYAKLpHCfnCmHn69PaZpULqEMnXUpFAwxbuB+/IN/2yJTxjOWZBA/sWg
flwZJeim7pxcZIzy3j8+QwnBYnZwnxTzANDCh8JQZ2AChNgh6lYAYtaYtaw/ObGC
KjkzjUWqyktTveDMLrz4zBt5zAoXsnvLTMEwGSfwZA7URM/4+5dhw4Ghu6pa1qOA
0EUJj/KTX6M56OFTBVmFr+em+GUgF51v6aPese/IqwqtL6mxd2ssQ5d1IRCzI85t
M3U0YjMe0hcOvYxuSAVdIJWsqgeGHrFixQAFvg2wDjO+kq4jVpP0QCP0SqLhh6vI
dlcWRsHr/GHojPJB4pX9a9dMvfspwPXTjrzrkSGP2zqeN/Awf7bcGUaNaL9KXcZC
u6kB9v+RlLsVReMl4N4BWPumoVDFBvSG7dLNUJHDAYOMWe6p3o6Tz4mbVBH6T2eq
ZvDMivrJt9m0CRKtOuVOS/nHDOoEdPNxM6fgRbg1HWf3GNhfHlO+F0A1uKy8t32k
C71Pz5OLoPYVl9gnqI9I96ujgeWzMatHinDhlesT78NTDUJCgpBlN2ySSJBqlPlJ
njf/zXgBFwuwy/1HA0DHh2mO/VhpMzdQPIcydhSyv3I/ebIw5VQ7W00r+W/55Lxh
i7dU8uDZIOs7Jd2L43U2oywWAOGJw25oOqeqKwwoEIl2eHn9Z5SYPsG3dnqFKRYD
0aJbL1G3NVNfHtALrnKIWEw/NgJ473gcximbQgSbisCu3Kn5AztiiBdHyFrloDYE
0C0jSTimIw2LocdDwgiOj8oldcLwYrIa/0zon9u+MsLPrV6k8LbbQ66ZXZNBN8SW
BtUGQ8HgZCDdKsLnq3GtdRkT6dIzhPy+ENqovZpWEphaKcNXqvTyijjCk+kHCJ3z
OkIDfqzQIqFkEPgXkhqbZobR/ZvON7nZ+i5KVcffjswU+TV/8i0AZrTwRgH9g1KW
vTH5sgEmlVil23DZ9W9/rREEP5T4DL0eRHW5csLWhULaHtbHhqx3ugu30aaYilm0
OlN3/EYm7SKmJMOCjwDVQfc3ubFE5vkeYuWAY/m1ziijsFzK12GLuFEVjEsAAODQ
xLM9jn4Yhi+Fau/Xy+IACbbimM4kscc6cXdqL/9mZ1DcEpWxTfJ8ZTdZS6n3Z5H3
nY5zXly3fuYbMjOkb219+Sv7O54TNMgFUiiPdTPRLTmd2qJhtueiQDt0YZbwIBFE
izaiPbiAdUcPjWkcYIIgBxZPTtnHDZO1Ex4SuuIzcboVWMC/Xe+2ie7p9wA32h4r
K8SFl71u89M2jrXIAZP2VkKJLlwl6iN7CqThBW+Yjzu/Oof52Ld77wQFdEacKvfT
hiJVnfRItssYZuPKNZuxvrZ8UxUCJmJILlytfXehU8Pe0uDKTZgheHzvRJXJqza/
Sekl4iAjphIaDGNpGctD1xiOluhmNBh5qNrEE/+QsinQZDGSu3eciDctEUI50MMA
cmRH0g0rg4MmlytL3pRR2+5dIxgQq9jYDumk0aq6w3HyNt6m0kd0V8LNQDFmhE66
FnF2oCixmTttxiHFHJzMnYnbIcyUVWuU0y7vxvPuUzVf3Xoggly7RYCXE7VxGfmt
qTx9A4sO+E0XKFzdr+njJNARwzHGQbQZYAMJbHHrZ6sVrf2Wjj52Elaww4wW0+8U
vRu8Hhsp6TlnTT3Btf52V7cq6yWCptMrr56XQUhNWcTNRl/knpiDJGGOvJkKQQkM
LXCb3JfyQWMvj9v9kdBAkOn4vp9apGRikTfzm8zwEwoEd6mUvoCF33apKT6Fdipp
rOUyy4PpC18kWY1fo2qyxbs0p5Lb8uxVTyDcY/jbEiNKNBTF/woztY32sSq6sT+2
5GtC4UX7BtUlEvWT3GQQD/YGXLIwkdSRt1truyC4SDepJuOq1kh5Lw84MzgFX/hk
6ZtjhGuTy3I9KYK6NjCmxrD1K+OJoWl0a+e8PVyCfZVpEOPZb/Mp2x1b/9h2weLi
3mY5wriYS4C9EoKTizf37ErgXdD05xRk6Rx4WphxrpgdyeW14RiH9utCOLxI/OVm
hsKMoV4BtA1EtFS20/1x4AE8iunSVbsTUZubedc3tfwH+1Gw21tHn713FT6+eV+J
In6yIwiynsfUxq431QidLQfmRuL7CSBK7jaegVQZXi9Xu7J1kUUAxOsAN0JMcS3P
C8PMVWKn1W29FI6vGRJeeoS180jc2f1gxsUxeZWLIrK9313LxfcC1vNIGhvlra/J
C6YqUfsqFr1ccUs7NhymOkX1XZq9RGa2UP6qH+U7S8vaDgKri07IQ42/fWSNcwJy
vcQmRdLN3nM5X907dzHki0gtyPiikW+h+UUs2+1Bh6jtUb+B0+JY/9gbAfZaWfrY
awRwlUNqWRU3D7Tzf8f9xw97FGnzh/oHN+Smk1OJQf5eEy4cLJV0VvzQOhoPlXCv
QsVt0ESboVW15jcTRx4bx2ITXS5hoD3nD8iiv3A9NIvyGTmF+wjyuWPjINqW3xWB
AMz+nNTgcrAy3h6SUJbLIfk+4g+M3rrzkLu6xstT8zW1bF8lnix3TApxXoFajuLH
qVeO2ynXoiEYHcxfL+Cz47PkBtIvBh49pIlanZTetVN1WK9YefsRUNtay+604KTq
IORS1Pja5fjDImShlyzf8wZ9Ye8EV8/rFxZGDDRrEreleQxBht4wf6afk8zG2B1o
TqjHcbPY/ZWDI+8Bf0JVdDwuJHt9L6W2HN7BpxDbD7GciStZlbSN5Xd2onY+wgzT
zjMKBuSQSFp84R47MraCmL7xAqm/rA4ey6CGEP9LedE1S40vvGk4jFFxJmgbODl5
i/j1eI1dkj43PGAQt5XZ9t/hk5zf6yF6WvtUveZHhg4=
`protect END_PROTECTED
