`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
e9k3HRTTg+KKDwyMXGqXqXvewnZrdW2RtVFO+Bmps4q8NcrWmtPdFuDrZzkXlbK8
DCKxdlhch9CsFCroK5EVpga0rx/1Z1BaWBMFgf50nrPYXeGUZL6dEQZrgGzD3Z7q
XYXDCBnIyRIcisBa7HFSFhuafA4Q6P8ufMW+prwhaA80dFVLFpZijTapIRnp29iY
mi4z+yQOvnM9T/YPsJO5nzFxqkFA3uZcsA8UfeUo8iTHz0shgQju8rjjlEzCSP2J
1PuMoe1XO2sQ9vC7kleuwzzR+uk+E2VYivdBPxFqrKehuhx1yoV6hUwps5yEUSna
OK20cv+oTlSexnvO9cGPwmFXEImsWng/Smkqf8VfHodD7pH6JJkMQ3V5y8MHsN4z
VBGZg3Ru7WJOsUOYddZ+sCuY6BCNI7ezv4dU3gd4L1iHybqzyAWSbtk50YkhX8xa
KodY8Vn159vh3OBVkIj/DdBukaEFS7LAx6+jNzpKHQ6wdQq5aaPTRaE+a+VnF+aZ
eblJ67vGOHCifQUEtAB9lkmGJvjJ/W4tOCbsFhjcL/bCl7EaLuUcBhPeqQaDYE/0
JYABMJP86imieprbOe8ftWJn+J8j/A6LujOuJCRg/YFW2y6S/p3kcQOZdnxaN/Az
gF/q2Ns1mQYmEb1j9pjEho4bsyuVieLCgauy57tG3ajEILqH+poP3PEWBmfBvjU8
is7uFhkKoDFy3GSYSgTHYZlNNEEU0fFjH7/PbddiA5V7BhzqD5He6b+fiCpmjj75
ya7FDdhJJ9A6UBBu7nnXDLhouhKRvgE01tLczduOJtxUA5oahzfMnkADuWF4LKBd
Tz60XeSq+nBD+0OVNdVL3yhVDguiiJVAC2fXugrba5OgkVqAZ/QKlyqvyb1Kbzob
s+b7GbIsbjT123MdpiGhGPYFJuQkvuI/KwyVSs1dG7flmfENSAZ1RQMfvRzndKE8
ByfoGOoEb418Q9RNzl2jgXxjPJTHr1l8E03cqiV9sDc/cO+fIpgT3KvG9ynGHN5X
sTNi1SN9MSBMkP1hAchcQzzNfAJpgMK9EHyklsx1Fc9pxiW3NlyFOytcZSSQGIhi
Gm14a6EWJOapS5k6F77cjt7G94InOr3E04mkjAx7wPMyr0i+fKjzczCB9pXWikQg
J8DC6OhDLou+u3n6Y5LQ3+EFwyvAAumTDfW+LrrAURlFif0KLxG+1qVi2OV8Z0nt
IjE1YykuO1ce5HA/hEtGCO6K3SKvMyQ3mCPJ0U3HZYBONowB+tvGhtmR9zTlxkou
N8ENLLdQuwhStpL8sk3Tg1bs03JRl4xepPrE9KJRwymShdXby/rRAPHdBTgAGMI8
mLppuzCqW96neu64n99NYeKpVQnDE8CAGPXLgM3VbAdocKNa2pPBRqqQb6lCEVkt
w91Xs04WhQdvw3vEWXXX7ZOuR+Qb4QfAcmFJ1Xi3ctmeUEG6izDl7fIEXE3sOegW
SoYwop0sJYCZ76YvUq7kpKyNByZzP4PKcTYkzvfUKw/zo50/AM3tKEZuSltcJqvT
WoaxxUb/CFqV628j3JvdK+wVyxD704OaB9NrzFsUAUubRW3qWmNrnQeHvyThuQPg
`protect END_PROTECTED
