`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
n1ewOv+rzppiVx/u8JG8Jy949gJcGAcGwW66xr5SCKHhgPgCxCDGVMqkrzhnMeIk
8yjA34IcRdcz0iSZiy5+UOa/8zjmjlfnxdLUaUXws4cS3yOz0GDZcFQPcmJDCn6o
1m7N7697b4oiWtL/pezI6axEpB48euy4y0eZfjvizzUFzujg3zM8q/ktQG0kwOPC
HQuTShaVQuDIgTr1vL7LjtPp7FUaQhA5wXFfdCdz2l733jQ7vOaGVyiYnUZM9zvX
bTA6yxigxvZ7ANsm6WnslADyoeJM76ERtK3CfokXqV7pJYkve+hcM6HJIFswePuF
NmSq4zrwiUjjxcTiosttzZ72Mma+mbRjU2J86UyYQcsNs0AQDjgA/PCDZ2vFzAGp
QSLy1hbaQHpQXUhXZRuJbrSSTxbW23ADce8+TAUawnfHi7L7ANoTg+7oTBIurfva
i9FhoGer49bh3RjmMH/fEKwwhWwgHRL46xn6F7VapkkEJJOjprAP23z27zhkfP+S
6B+jEpMuKAYKKNzvxphXMA==
`protect END_PROTECTED
