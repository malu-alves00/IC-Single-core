`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rf5udWBccJcA2rJQ1ZPS2lsLMYr8ar1bFair5bvnSfhkWPLXlWQ7v38sfcduFdYJ
PSTVmgJhURMpLbFIytcM2HEO1TC3aMBSN3S9SkTBAzznOvs9mkCzkDhoXYkojIZ9
eqBBZABea8dSAswguxmE2ro60q89C7x6dl/UKTZ9L+4nDMAMMdG5t2udydfgVUca
OwjvgssT98A3NKjo2Q3Yt1v2UbWZqffSAp0+3SEuRliOlAsRiR7OuvwnhSiWgEGY
WBrznBnzQLcIArhU+FA/acrzjUueDc6uSNNrFvOXoWEvaQeAfMoHQvPQcS98arlc
y0/7XmeKrekqTpWzEcd3G2eKvTjUr9rYomTOF6QXLqrppoU0kohBzeNdueIpL56U
WOmND2QEPjr+OoAxAtBrv6xdl6WnC/XsWhRkPR/PmOVhDhpQZOF16K5iCQ6Uceny
U4VC/CrMr6FeXGC1mZEfn2SYyptqA8CTaHTmiutKLBxVSQJcVLrdqcrQhcRkzF4u
n6B8TwC1sgQc/58B2Cf9QQDlks013c+TSQ1od/hN8nqofEWo6Kj4orS3hQP211JA
VQRuhcvm1EAHcD9r50vJd3iYcEEUFdHXJPKPu8s8Fjgg4yil308vnXb2ma/ALbAh
KmIEzTypBsyRPduXeZuJrytv/gAkyVLlsZdMJDRXEXtuSBYsimeCCZ5HQEkZABQ3
xMQr3zXebgkZqo00dvyAl2mANfZLdhGq7/vwmwf8GRgICrHDf7kFQTJxjkDs3bbA
gd4FyuLaxeSZoU5P3HsE58rB5IHmN23cxp4dQ6FDccI=
`protect END_PROTECTED
