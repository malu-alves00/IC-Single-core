`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2MhKkijb0SD8EnW8cYTvOAKBvXLxZ96/jVFeXPsFUkx+3mJnAQyZMUMuRBcjrvL2
P9SBVavxkhTGzx1XUHpOrzrKAtSTtBjtYF/512MVy3gdF4F4VTvHlD2jFparJfqn
NYJhaQjiCWGA3zD3bDUtGJ3vW1+rfa9Jp04dHdS+arQYj4y452NFuoFijtp2ArXf
EKztbdyvX25ngnCnLR2nFwqi1HB8gFtwD01xO1rESGaxy2rdvdfYZC+3ocjd4O/1
l9EO11O2t7c6EM3oKCOuLd+gnp9yKZfAbcCdygZW0CkouHRfBCABKrRozw1kUPs1
KO9F1CXDZiCt25BsHzY7zfH1KrUvDZZrv2KXjn7JAh04QJBJdeB7S6tIiBO15lix
pZQLSsTde8xm3WuyQzTpASxGg0YdAdTtvz21rrXWb97LYBNs8Mkcd0mBAONbKJNM
geKccRp/nByCy6rtnYC7ATOp6NmITUfCESgDvc3xJ5bPSJnkwgkMVc6xdgaiJdWe
X+Ihu7DfWou2T3kiBjAQUBT6uzF6bqac8zpEiW7kIYi1IRB29Ai/l1yi94BbvQGr
iVwkIQ7Kg3U1hf8PWZLSkPgDR4gb9ygOFl52Z3tV+HhCfIG3QEEZ82Y8hlzYJRia
NwwIXfvF/gi0v5Y1FLM5B8BfB4dlNNC4zVzCDyPTfVPahtVgA/JS/pFS80fF8Ya1
i6fHuifUhlWD5ARHLECSr1UW7v+3PTN8JLrsHjRf/95VPoIfCP6yuzJzV3nmjULD
7wf3l+iTjae61k8L9RZeFpYMQK2SKjQKCdsjtFIYYx+DurLnCMd8qibDDwanFU5R
daMbkeJJP20p07p4A0zaPQ==
`protect END_PROTECTED
