`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mLLH3piZQU8weCG/sUkY3houW0z26qZ5KqUh0Lxa4YqVl0jC0OMqCBKTIGlKhzpK
dkh0KSAgeCBarmvrSOJxpcTiJyyLL7+t0JGqRUopGWZMKywVgt9mIOET0U8FGZ20
wKLrdQ1bWLwQNYwETFX6QIsCjJb3evGMdSmLlWEHtE3bF+vgyj4HLpN59L7jFA1+
90IbM6W/NRwsOv29qmDzm1fusowspL0+cHb1n3orA0YvIKd6Lu4TcBQfQEi0apk7
F2L3t3GkrBo5IG1R9Ojc0vM9N7C4+w3w+OJMtbfPiuvxnDfK+Bc+/Qy3trUfdCkM
YcXxiD8j8GfnBrsBaj3ut6ScgNeNoFs+ri/8iYI4nwsusZP/ar5M8rS9bzxuKluf
llNGpdGG9PauhOHl9IOScF+6CFMZD2kRK+qbQqf9qQ0pVauxqYTDAR5IDwqA7xDh
DVVyqkt7e+hmBW8aOxUxJrk++Z5HlqAjOTYNZM9sD7Y8av9Tc05r43rgzJzFcNGH
DcL9smQnyDW+RIJu7ZMsLLKn2Mu/moej3oIMeV0gRzMnaiN9l4R0MLgmofpfGpjo
jvgW6sfkuwfw4PClgRNJyCvYwmnXuJ96cw2AWOHMvNFAgmOoe+na/+/JjTvnxNyQ
O2EgYug+2f85jpe2D+o4DzoqSy0H2ChLBSYRp8Tu+SDqu3mTrLO78AeY0z8OPQvq
a8XDW7OTMJA+pf1VAh9jGEluBUqgdKyG1Jp7TZ72aFL4aWyOCyUbdMXXgnWd7fM1
WMkxtdsCyto9umOdVgsymyF18Z0SyFdxYLuZXku+Mc3/cfXX9Cfnpjkx2RsnFxuc
luscWur9G29rftVfp/V51NMV1C13NJ14QD42sMSdkspAd1ONfru/GlZ+h4uGM+lZ
U4iJRn03X+2XHRjydt6HhEPaoqPaI6eTeWV1WkisrEYOKj4aqSmGUSAn2X/NHFMG
yvkY1zJhPme4LBrlEk8lyNvoyiQART12ADJ/A7IjWyHueHe0cR2VbeZHP/z0cIYR
XdscO50S+uf7Pf3b03HMyQmtLgNEHqfvAx86A5RwTdnW2tR08lPHqx6ICxv966Wn
ZQ3cY5cNpOqyYm1nuVGnQDLAz6A1OXhcyb0VH5/YtmDpid53ii2yYotwsRGomi1e
adWFm0WG1oqG4nNBTd3Gz2T9Xhvi5CHudqVndadvnpih8NwPLkw8xbJItmFmW+fm
lARF3uayeXxEckdKKNSUrA==
`protect END_PROTECTED
