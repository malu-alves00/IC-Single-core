`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vvvLFMNLEf+/xq00Kh4fI28RDj05gvKsYSCyXhYK6i8IHlmurtaNtwGZYZo/uTMB
yJ1K2IvJZvTkTl94nCH3Tg/ZK+B1DDc42rbQXsCMaswVvYaaE9NdtA3yJ7GuO6vS
+HuFrFNruZu9+jnkmgkgDw+FTe9eWASA+2aTSiRXTsG5uriQQk4zNUgPILjuoO9G
ZdDxNW3LxLT28kBXYbvi+Er9HwU0OLFB55QTug96K8Mn4I/wUNCSRnW7XzmSK4Ni
ywgx8utgTLw56PGigpNjdAYUS1ehF+Da+YV5ixZWbW+5+24PM9VRpQJOBEDJUNcQ
hRPKjAgnGI/GQylXaGXbJ6ksnDmEd04EBJ5Yrbr9TIky3kEG6j7GZ0m9JejDKtjx
HCaPsiwOuc4dfMKR6cLPh7nDKg+Sib34MLO2QVFFEg45cgFXxBQpRzTZ3xi9SYi+
7A+Y+aKmdHREoXmrZn1gui6fXF779XcQEgygl4uFQJqgjzrXquTuk1XN7F4CJrRK
LLNhB8DPUNyqYsn+Ddie964lfe48cyQVIpg1Qp/ltp34vpMjoBChYV4XR/dEQW8f
Tl/WbDLSeG07h4bMjuF2grAQzyCsSZnkfXxyWb2hg8MEsGhsjLA+4l2lBfP3psif
2OXaPGOuPK9d6vrqY+mBy8aWw20lQ6DNZIinpwmFWmIlxCpLeXAaCOA4NCv0TNG3
CxFX+rNwroy+trGqcpipjRBaVlyBqDev57kpfpxvJ/WRdR2jyopYMqbfp7zI1tfK
NP0GJexD2cy+9L3BgHP0H0MswrWB90X8U5Xl0oH0tEUv/kHeVwg5zVrRqSMrP9x+
pj1nbD4D+feWlyvYoqqUyZIKnKUchTeAhVrxla0orwJlwnPeflipD6PiWnbo3Okb
ePZyznztZFahBJAc6ikC7l0oMFCC03VtHmJWqMdcgmKj/DboRxvK3+0GES7Z02J2
ar/hoxFTclzESsjw28mikePQDX1psBVgaVAXML177tRxCWqm5oPwvzQtCgt6kPr0
IOwpsYpTVQsr69tqiZRsNImDYRBv52fdHTFRFcHQsizqqO95bKFcghW1kV/HA5Jq
ABemfzS3mOdSQwsisHloKbZ1XHkxpmiW+BIpn+zp3wcNemQz07qEvccTRwF2f7Wu
6CnrkQi3EwaL1fCcWp7tl8WfpsHgwyXIl5lpaNfidCq2Jz6PMFESeaJdgWtLc70H
l6+rEUeRrArIlh/EiCraJdlX6DmU5/G5svPZA5OJfEVDBT21kjO+dWymKLocnsgu
38dLbn6xIHDEH3dGv5bJD37KyWYa6LoohMRNC3Fg1Xn+qZFi6fkqzPOeZlH4Ohah
q2LNEwxPi1B699kstgimEXc2X7K+nHKTfSkydQGpdAmQWlcXI/SDzvF+K3U2u0GE
nCTqaifjKCJbrW3ga9B4B68ihfxS/Z83t8aH/MUFlPdhMRMLO10YnEIRpMxA79q6
6xfSWkYRE/xVbMjKI15dM3tf02o9beCWI5SNm5Z1ZklT6bVwzXiBvXF75yZZ2oMm
hlET9goyFsKWfyTlrTTvtsLukEJS+McHNTU2/H+8g+RwdJE+mWBu22DTMZgzOZzJ
Ul8eVUoRIG3DsD1hykzJYrB1mDWq7ZFNjPtU42vMhAZ7t0QhQLr0jEF6/nhkKrsD
bHLozGWtJz0XTaIhkv+mIkuqQZMIOiM7pznRV0qRonM=
`protect END_PROTECTED
