`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
p210o2cp3PNadm8RZiEl+dq9SUtrylu89KGSzrHo3tvWDzMKO89QVScZTp4XDXu7
WTId60giBg3maGC4NW0AwjNIRpKwvyDiYSppALgyvWxdQ1DERvqDRT/6teZPj2LY
VQH5bbXtzrS2Umf8NGeM4kO/eB/hJ+ZFTVKTUEQY8d83rr5xDSSKJZn/KKBdlZkX
o0qad4g8cJPKeMYeQDXqomhsrjYNjJ4c3ctDaYHY+HnhNNc/krPbMu1g0xA2Cntu
PzvK5l5SlPqwxqDgH33L9UnXilRiW0lo5Q24fe6cqQDO5BNBpmwcWKTq20x6Oex3
KqBvcM/mud9kNDKvr0eJ65e/CYIpV1ijuRlRvWTvRaXa6LOJYztE4P5M5gX5Kpjm
cuVKnrSm07IqNEfSFNXcvac18iv1wmpt3isya5VVw9ChcJbr376SYNphi2Q4Ae4P
Xbg/qEGHjqXBS0zCKxnisaYmBqNSDP/pdLuT6zCuTr0ZNSZnrOuavqWwlEQA5QIe
nBLa/0fgC5JxeQNh8Fo4Q3GDJ0lKDbdrZ8Fy9BrF6pnJj6dN4NAE/wRRALCNGQot
qOCwYD5EM/mew8dqdY1qCMr76UkDLDg8Rj4+EuKFkduAVEkDbXLjU9omcSCJapQV
6ssxgGiVVtG63nZGmxJP4AQHZG2950RtIowRUYY8H5CoLlOyoqUizGudTO2MEfRK
TimKr438EEe5NM6ZyvTwf+Qw0gd+tO1z9rb1wj7GDd5t+EgMjOZ4Lo5CyOeq4Vq4
5OSpX9FWT6Ds+gY3Be/PmQK9wPEbrJrMXfIkkrL7Dcc52v7PHrljOmYjTpWJYcR3
gkNerIbx52VtirDLH+w2E0li4wOEvOJPNFKd8zRdKCHWd93rmuVfX6uMYwB7z/+7
hAv/sEz5AQPDatj/4cPWilWuW4sHGHtI7q40LS7rkSGwv1OuHZynBaDItxR3xQlu
H8dyMkJpuE76JbtP/xsgXqGr/KHqygSbVFY0Fi2gLQDzQ7xINlLct5vStgcOl30E
xEDIQWwfOlgJfDjGUESAYtJjCTThbddpUI7XV1qJU6yU3ooIP8co4AHzbp4wF343
fCYZThqFAYLRA1wGKKTwwx1CJOyuVs4ND5oN4CFfPBMgtg25s3xCZeLQznj5b6WI
/Kc2QfFMnp37ha9c+wFNKNiaVPjhKol6J3bmITpvvIBC7T+8rEA92rH5z60sCj1r
Nv5+IqSPEFjQrMSOgQOOhX4743k6ihoK+WpChgD0CLkuYMSarEgB4VYD6os9ugDd
qpT3nZrjOpSc7J0z1QmsQbVfrrqSCiQ0dI9e+0RP8XybIme/pKb4VQNsXxs+H+wC
ioPdo/Z2upSkOyxzVFAHtvnGwt8QPqNeGA15MX1tGgWAx0MAqpR4lHLpKFA5mfQn
QA6kuM2hXtgg4SeA/FzxCHuljzl61k0Kaiam+9wwtLU=
`protect END_PROTECTED
