`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nbLh12F7f35mjLS0OSc8ChP2zgCJrPjF9szrl0Yrim24Z16pW5JnmC5e3zSj0/ZE
C/6Y5NqOyUQLxDTbf94aFuX+m6owLNoZAsoXzXO/O15xqMckOHOKZh8VH0LdH0Lu
X6qxeAII6aDv2rzHOkjGciVIopu7bg43PLlZUrKslHe3o4te/BkrhTXbsyeLY0PX
ZRDsMUkLqWmdzCKw5wVvIlFi1eERGXfCRwY0FdSMXJqQuAtXl3PscGRa/Qp88hP9
u46VYkulC8i4loHxEkf6WYxbcJT4Y6uOiNmoqo5UQX1AlTjXId7qN3kY/F8bsRBT
TFQQSUBkBM+kQ4QY7EZ7C6WcfCjF22F+rK/6EAvfTQI94Lx/Ok4p/3MI3Svtv/2k
d9whA3n2Udk5QT7vJ1SG8h6ua7mb3iawj0L74tjySEKUjM2S2e7aygvoMNdojj2a
D5ty1QHcYPnHE3578ZzDVKzaR5C6Uv6W+4iZIS0AUY9PVP2oLv1hKmxgz7aWpm0L
A4MFce/VzEObX3RXhUuOFSAlKcvhNsAUd8vw9mYGzzTChN45CxJquOhxqQ5YrR3C
/xbbyx7XSFM1/n5Dlt0aXjN2GNTU8UM+lbDLX1rJRgOgwkv66u2Nmje0RNvjfN8e
Ri+F05EC88QOznKSCxArWIX8S73JA0Hy04hhh1kiQ8/Xn2jE6rUTaflmxPLZI5jD
0Ydvwk2jfEXevFj8QrhOqbsrTAlcsMNlmapVjaarlis2PfSoyCdRr8PjGNj7vJMc
6DeqC6P92pntFTqszBSMDySYpGZy0XB3RIsJIvo10aOn5KB00qhQ9mZc+olwYjND
xXj2fMCahG57ZgGT3Nn7aTS/+42j4PJ1TJ9EpQ4Twt9Jysh7YzJy4Og8so08FJzS
dQ+AbsnmerEnX8Fyb2JrTIg2AfkINdGYT92xShf8YokYywTmWxQJnAFSUoMm3LUW
JlZwSV+IRlBv5uHqsujqPJJXzpBcVFjxJbZRPQp0LMwIYcMRZz2qswrzJ2TpJyBB
mwsOeXBHXU5hpST6fHDxZmNcyWWzep6xALUqilwMMVCbY0tvwXGUUCEGGshPLGBm
XP1FJTUui4ED0ENUXUnYQFIGiezcFHdFcaLDCAkyopuKSIuD1w2m2wKOZJcBkrxU
0qZNNvyNi0fQYCDRO1Vh2cBfva2cuITaY4h6IilSdaQJA+ou2nKEp5+ebZsJKyEh
mI5l/F1RmyKjqLWdQ0aRGugk2u4nkxm2bT+mjiyrVHt3E/Y2hfOZrAGZ3/nQz4L0
sfhpcyrB8OuctnnQZyhMUYnQUQwfLi/zMLRpAwMbVtOxDnqOKmVVFVI3xMJLhbJL
oW29JHY59f4RVGRFQ+oGtlVxuvE3RA4mhxKSAJ82wjyjI+WkbP1M6pW+wTI6xm1b
eIrNJKIPQhujb6XXWUlTAfrSDKGw63NQoBx2Pt+0ccuODpXUsWRpi3EUPgwqXf7r
`protect END_PROTECTED
