`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vjAPWKsYcZDOHbNMzH81u+5loG2TTbmu00Z5Q6eWatJ9156QwlU2Psp5TVxY+U66
GMG1UQD3hkEAp+4bYWA/cbS2czokLw5AHgh7RkMZ0bibP2b51bxlTBHJGg6e075J
OsCpl4XjxiAHQiM+GSpV6HYR1Nm7AZEg4P1VDgJi0yitCwbKYYtxQOzSYah1dXm3
S2OuVV9hmi0PXmoZukYgf8/9X2j7MDlnE19EigujGpQUlIAOK8haGC3Qgs6V65Og
+lYu+lczxVf0kLEzL4yJQYNRhzGMd2bF/Z9LOQwAL+yBW1Cp5rcgtb3GIGhGpYl1
jYnTe0TjVR6oJO+ddhiv/NIIiBek+NI0lJofjv0iIleqWbylEGw4NYCMNdj24vKh
aJTaiSOJPkkFVcz0rDfQVFofu7SCeLCKSYWMR6dc2ZVQVGtq/071Hz5x971AS0g2
8XKfnkmY6m1DoPtm9EcrIxxnRRiix5TKIeRe4BvbWensfOYb4juxsfbBx7BUum+5
crRbtEPns7nG2N/o2I8NNsJdQpKC0sUWs92tnBnjOeGmpVo1OeBy4YyXOdcKtgEJ
eLAaeu8p0aGlke6HOvszCUutUfZsSPe+2MRvRwIjmFgJ5pmBdvn8q8rfgr+vjFks
n0wkeKV9VPhrGqFqGZj4aCf77F4id8R8AgtpKHPBlP7MpDHbus473lUqJLdDrWQO
MYL6U+qbMg5guUQ20kAwMx/FApn858agU0lFm1Q1huohF9aw3U99eaSg5eyQB+yN
Zy/JFH+dTaiSsEUDKGFkqCzUVh7k8AAOQCvPshUg+0WsoeWsm2bW3ln3ViuWIIKE
Rn53PAuWn+qtgaKVsspWYHs7cGZmCNZ8u1GiqzR8d+FxiHcg0RAGxgmBTVmn/hS1
ZSiFg7Q5Eg8G+gYf4Ez6wCCRPx67HMJ2mezvGqVeLeAfrA3fWkmYoraqbcFBjrLx
UBAB91bGq/3jl12KXpHrzvzEkzaAEDbHzTHe+B9I5AVucNcMeeEZxXOH9RvLiDSG
lq+FeUJF3DUz3f+u4oPfOoJ1aWYsVxw/kjvioxqj/90H4W4TXNsME//+j5tQO2Px
Qv0ZoM9hYiiQsfEUdU8HT3nLbhxVCBOBSnkhRySVA3ASGxVY54W4jmmpM1N3/SLQ
0FiXzB2EPcDmuoZ9Byy5xvs3puG+ZEN9HqwnnOT6S+DxGIE8w9oGrTcbFVmK5HOz
gSDxmAGW5ZGpwh0ZSAnblcT504cY1QFpeqbAONVP2qrGyrRFeBAmUgKG73iBN8kP
HWEdIO+LLN7snLyP98J9odq46zLWAz2DQYvkjrN/daNDbFoscbros7VJ7gh1O14l
zEXvew9H9/i7AyWPENoMaEWPmGiGiFl+al3VUMCqvSU+16F/L8thoj8e231RJdYL
0BsPl182EkBVW+08N6Hq+3CFC7/XPix4wwYOu9JAXGzTEx40yhqAobd1uRm9Vswg
l7b3ioxWJ+wKS/SUjRZGzqRenNB5YoNh0rUdhm4isDjfBxuKImF2zXPTXLdH8KdX
8vSuQPz+ia2sdP4G7gD+oUPARQ/TON2EHxeiYVPEQhgaL7rupE4hR45qEJWjO+VZ
yN43lGAQ/ulCO5xptY0VRAt2wLTRspICZizmLLsw164=
`protect END_PROTECTED
