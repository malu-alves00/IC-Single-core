`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
i9jqQNwnQ/6+5glfKsNOA1n/whpl0QR8wcbTWWTV9oMUXLA4yajtZYmkAZMXttVt
xKwdobzeKwBJXWFJjLz9E+eLDI3L2ojTvgQAFuNy1QUzmFxx6P/w0WuxA2DJ/hGp
rVi2L5GfYWvap44uRldMnJQDZp0nsALYQMcxRrBq7hBn/Hv+cLGDegf2V5ORbwoF
AB6dV79i3G1CWQ4CfCrx05vL4mNpFUVQ1Rxy+mJe56jJ++pV9nwilSln9gKg0LEY
SA8+H9VtqKBMa+lPxTAlaYWcOJpFyLtiraenJaf5fWZZA+G9SATciIvAJflQkH8f
74M/V56DCKjXB7vhR++zfAWod1i+jhywMZ+KmSIdkJI1zUq7Dg4fzqx+M7Na4w9G
coiGeSrGF8aKse9mrbtjV6wBFpw+DaGU4oPqSVvtpJMxzX2ttz5KqUBiU73OJM4d
z6gxJmSKggOWdV648M/eKxdXJ/zjn6bpD7ITJANSlGk7EmcwFvay0NqsUdGYYNhv
KIBLv1c71u/G89Odw0DN03HnbPUIuEL+6TWuipFbuY8E3iLggostzumPwz4RE1Hp
Cw5csDeoyC6NjpCPeOTikozC7qiJzyR6uGvpBn4gLGSwxlDJOTk8A07x79F8zuj+
aGDg0/Q0Gy7/4oUSKtZwEf45gB1rZNonUzf2dTNaYXN0puqYPaWSsuTq1JP5VEWF
/WcW83Eqb120FVGi4Ik5FMpn5xNfnyrJk8o8fQTDwNcVSLE7qebV4pqoKx9BfWrO
vV9JVj3sLSAsK98YUT1z8rcesDPT/0vySnrSzGrZMsbtG+Ym27c6fJa2DuS4/Z2L
z+XTSm5v/9P2nfX6g09PuOrXSIWpgEufM0kFA3kP+EGA5ae2CPssj6aUNetiUDra
bJby6DCASBXIJnWnbyDLXhnlISMSz/sJXEeLarzb2yW6806Ua52OD6qT+LfXdEHZ
ArGMkREJOxDwkvB5+CrdbGj3jB96GPcCfJlG3ReuEGerpBW9HqteGRquxZ3ct1Y/
Iozj2hP6s3o1hRU4B9tOlbn0IPyiiYKNzSJnJmUXlqGaNNPfr7wTSMHmvEkVZeo1
MurNHkyYkcrcbVoAVRpL3wqSGMaGI1eB2ihAafrptnzBIkBnKGUb0w8oPCgYw96T
aEB/Q+gTSKn3u6aAWQw1hR34ACna/vYpyl+VcHv17Yn7nTPmXiBe7Me6HAKp6QTm
V1xPLyfAr9BCrsVuI9grh4YLLb8OfpP0kufTGAE+7zu3sO2GFH6yZV/rwmcsy/Zh
66Y8AHLj1A1I8gUlxndUgBV0xtBi/hjGghcIBHYMIlmxvjWhsewPvcWq0/73g2M3
XIp7OBVJ3EJozBz3GxWkP4DBzo7uoe3W8vT9fHr2ylD+cgcecp3iExL3wGw7S9L8
411AiCiw//hnCcGWsszVpv3bGnzAfmyXbGGvsZg2c0l4JoBCuHdjsM+CggWk/YCS
UA3es5ir5p934Q6LWF/jSarJet9WcO7Wi1nr4mmM44nbf8AUZEbiGga7B+TCQ0Wk
Z1q4DYii7b/jaBgkyPnDbRCo+y91cb2lco+j6PRp67fZSfPcEcUFVQa75m1/KjM3
wbvD/rElIeceLXrsORGJWGxkYU2xXH04huBvxCzKEFBso+lPx3T0q1o+KC9q6EPy
OM54ZF3UnQgF+VXTR63+zlNKblHH7YHM8vS594L4lN1ZWd8c+Bgb5CFBQAOlRLTv
oZikDAVaeocncMCOYbONSBYcWof+AJWZlTtAKliQP8q6wRRlntRS0+jt42Sspb3y
dCRHM/t83kXylaYW0Gr49EX8loV3Vv41TRBGNpSwi9aTiZUqjKhrCatsZX3CpNZo
zZBId7bOw/L9eLV9D5XV+NRD2QTcI9KlHq+JkNLqxK2LZZVG7vTWHWdFBhnt6SZ+
F7AB1efIRzt5Jv1KEsHKqymzWsQasllQ3QqJSx7pwmIn/gv05DWBL0omHt0/dC0Y
K+9oJOgNcVO54RBUSC57nyl47Zo9jpDljvOtbUx6FMvEko6gbFZnkW6kUJaYz9Qk
KJGT6Hetlls+ANrVUuezuUCNcrHkr9+1KyOOSBzbiCMnCj1vdyRyUI88PrBnDKCI
FINSjd6uw9BrRc/u4kDNIzaGU/Dg50ISA4dz80N1YgFPeU7wg8J5APp77HZw5wjc
T28FaIhCN7ymsV3/W/l7Ivh8bCwgffmzRwXnodkl4xumej//yzem4Sh7jcDlBWC2
70YFrnfh2/6ZYQf1pdcpqfCJjE0AVfdGWHJIQbI52EgHYdLhrmmVDGYlh/uIIZw5
QNNPgVhITAQv/0aT+wKtrZLv29RAp6jWg8QEwlLSztyW6n3mIERK8z4EnTf6+Ck1
7BSpkjWQB7xDtfo1r6PwsZPpFU0Rbe32UR/yXKHqYiqpgN/xD3nyt2HgU+1ez0kv
6y2JOWqRRq4GaFv1vhSaHWF4owedD5Q161KjbQITfn+5wHkGPnfwHoF0+z6TnGtj
ZMhbLkefcRpgbMixWVzXQTcIpCw90b3tVYhn0QO2u+L/gSbsBVxYENB3WwBE36tV
kVKTK8Vw8GCOQgpk595iP5g3wigGat4oTni+1mp1Po2C5Ee003IdH9Rs3MDfxCGf
GMDG6vcKdDqzorw8ToRQtsrpPGwFnnFK/0sN0uvLqCHE9aZs/BHwbztFvtoFrZw1
E2DucOUnHWvhge+8BcjypXBV8G+aCOfOXZDvD90KBntOQ7dEwkez/tUrOYuKSRyG
f6+lbjt0HeAsTVOef6bRtH3FmmAn0y0p6WMY14OZigsoOKt4FxYdiRpxjwLx/KMH
Sdoi5i65JSAMzEsvsdJ2JZy6Wyhxk1LArZqwvecPo9U/cMSg5TvCc7eRX2wGfBRQ
k51SuOPMxlH3EjXqAhMDD5m3+wOMoDeyxXXjvOx2CpE8drBrBNFxFty5se5z6S07
eheyqydnJYncnETZkoIfO9nSy710xSUCzumgptM4Iibu2Zz5m8lsdXKhJImdqLtD
I7q/zWd0R37EeQizRceDYyfCZvk4/b1ntnOr0NessXJSx8D5TfwUQPWmZhOnsJLn
pVjU2iYgaowOvpUG/v0zoWwWWp3NrrMxocaB9zxD4J8h/xRFWrkOirBwWvKHUtyg
RxevMpgL1+J+WlrQI8YuY01K2N+6HaHCR0Bupjcjw+At6ViAvTk7XQ8qOEzc3dz0
XLu7/8A0l0jWbBhVzcqa5g24tJfICWJtGs/6yDJTcik+D0w/5WZ9Ld4k4Ibkd86a
8Z9GhnQotJCp+0UrgTbdetGSYVkdhOXFLszhVW1Mic5oMeFtl9fxFLeJmUF2250S
fFiN9tms22DgLJlOui2TeoD1o2XoM+IOkgQJloUQp2naePqweh1sBhuB+u6wgMVx
Xrm9Phv5yx04n1su0iO4uQwtGDEBSfRviRDJrL9YU8qMg72C5+jWBXR7RaPU+xi1
`protect END_PROTECTED
