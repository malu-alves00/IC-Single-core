`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8afXhMykMSQnFbd0c/REJBg1MDNCth5ZReTgpA2VE+gqDKp0BaRk46bcWLbsxCBx
ewkXhV4sLXNbT2evGTY/9PTpKN612m1YkJWJ/4D7WipyCM6o/SOOj8Zaqg3Weaqw
dXKYz7WuKujfVuOIfXr1eiJqIYR4f/XXAcMcswiKe8BzA5iCTYMGFLdvawd4a1g8
FiwwsmOG3rk/01OlVOnnWNFPxKAiENrWydbQ9VvnOTnoyLLquFwyKGqgtf4XRg18
DGFWdPVG9lhHCf8gcHcTOEWKD+z620yt6DeE+wzeVHwz2lsmRIvApOBnMi9hAhqX
/rDKubecIMS1ncDrUHH1f+6MIgAFqA7A4H40pS9hVE/+9SfgbWm5bSsPu6BP3CSg
8O5wQn4oYs8K1xxuUh6fHejykVtWJKL1CWTz6//Jmxcy2krl9JDpTIFmDYlvI821
LDA7U6xtiWhXVx1ZTZ+EzLEsX+a9R9K+K1M/dSOUeANnClbm6xvF5ctNpYYnaIo2
xBBnvRcOBvM4e17WpP4ZeqlasOAFDUKKawVHUmCbFcCn3EC3tVlaB0ckW+e1E8sq
+LRFzmD+dSvCSA82nsBNOg==
`protect END_PROTECTED
