`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uv87Ig8df5NIYIYwu/VGBhKVSGRK4xUcW4kV9DVmZ40DIX8e5aKuwPtHS6WdrrmQ
yUfc0z3qhhpVFzeKVrDPq1JGDLEfStYW9sLc7pq184uOC7Muwdf77Qt4eeYtPxL5
trhn4oP0QBqt4h1flAGSYPDcQDwzARynngvcMbgc4qb/KW/AFfBYO0/bqOuBT9u+
WlbRZONBWC15GiTAH4Pgj49bYZT+rPs7W/oAODJWSz6a5ChgXp18OLVGSJ3amEPp
QbHO7eOsbaFGqa+lza03dy0kePn8th9Vx5bvSk1iMBWs5MLgUICZ7JgjvcPMZ6zV
aBxV2ObELaGXdsQ6xjVKAmRHulio4Vvlx8U0S/aleYF2n+axImN7SXvP6SL3QbuU
RPNkteHOFR0UQAJCdPFiwiPdDHf7a/ez9uCVL1BY7IO6ej89RjeZT5k8vfoIRcgp
o+AcoMK+7/SjPtSbSaRt6WZNLszHSOWdwIUYVrkk+K3RvDrkPOc8YgQwlzq0E0R4
OdckvGESsgn27tlh0YpWOf8uTsOlBCO6kI2Jwmkt1aGeBwcdCgiotn08uzRHaWKE
/wgiE52VsSqP3sic+i0CCaTjYreNkaXYA4OQTi6bA25Fooh2WzbXEE6397nJ7EZb
x5D+uMk9b9cqSYjsbr6RSashWkWm2yHY6g8oC0Dp3Ap3/Iscs859B7So8UAp6j3Q
Q9ZfJeaYnV2uSTg51eC4QeAvdvz7TzuKh9f8g76uT1LdVzQWZB9jDv1JenumnzBX
yw53CDRnn08wGqKVYAK1XPCHwswiZnIT9/S3B1NDGVptcvgaUjeQc7VaGBGAa6AY
vkAgo3HaOFOzKqoMi3hJG+4gz611xKywBQOhqdUlsALyuoBOp/VfTFDWD4X9QabS
1YUvFIq1FIu33JmYDBPFdRK8DRdvrik/DAPgPjfO3aDPiTMnUOo6rJghEjM2Iukr
`protect END_PROTECTED
