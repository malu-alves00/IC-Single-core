`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7yHy89zVWMv4IBemmEpOEQhUlmIPfvWCkRxMH94bDSAJ0Z6e8dVyHuIwwiBOCCHn
DjedXKI1qSXApKBTlzVYAFHlBQrygbZIiLneXGxKLC7PeC6xO7+JnfTTj5fnTyTt
wfdn5QSHjUJDMoD5eMBKvoVjPa7T7CpmUaqxOzpvgwexgLCczNvb9x2XRmhhAFUF
gcx+zrP30LJdl7bIoPeIyyMff74BuYiGy/RabXBnlHZGhTo/u2ZwrTNVyQ3pOZj/
VdhqJgMz6KCibaVKm93CubenDtk+y3sG4QcL1vg4IDw3qvlFbrcUqsjEoJLXfrwX
KmBb6avQJ8VioKl2c7cWkItua3OQPgeWkhC3PZ2eXgI1qpbb9uGDDy579HXA6hn1
nabP0sQ72YfPLH31DhtRuC9pmExFiJ4TY4YPmncVaplx1JL7PG/jlTFj/8f8Vciw
on8U6+uKTR4rPqh7FQ2OhS7ZouufQOtEx437IIFaTRl2Uduyp9dYHVlU9Snf0wHZ
dHzFjGxfkXgoVqPekUGhJyXEruF7ENmFbscrw25GoJwYieCbFfyWkrrUdPfnAEBk
Avm9xexQ+dnUAmSNR20rBHKVBKEAl4naWV2fLAZ8wDJHOO5xdMjjWaYSUe+UAN9b
Yyhlvl178cew2sMlAfH6emaAYnP4XRSz8gxdvufqhoz+h5C7TX13dtGqq7pRcvmp
NdtJ51fS1289fKyZdKts0TXYkLjibF3kB/WanbBHwfWjLwed7EcuXk7ZRn9N0I01
bLVvyTmq7xO4KHGA9nk8uUsGonOpeEqEL9IzcY4/eQ9RytU8vtcAyu0+RhyEacpN
IYyMhcfKE3FPhnhhVsc6/7TO61XriRcMi9T0dcwkCIv9FYV6lBww97T5Dsq1CnDg
NHk1wYxOTKOzfa4HyHsbJT1UVB5DU2ZYiv1PGkVmxjFRt6MWMNKLWh0M40h5Eu8N
alptSnnBFblIwkITA7YA78xKNUB1JKQyFI6X3ki31DR5HnUAFCNetiEwWHTR2GVm
uujKFdz2Z0zUEGB1kfrlVJm+3lr9FZDh7p7YZNKZaKNOgAgR7u5mksdYvJqtp7LB
URswqt11OKpDsMynLsQ1D/BZcztrQJovssOcpP1sjr9yyK6cA5M/tkp7z5oGCfDc
liRVR6DBJ026/Frb6N09jph8IHhuJxtG02wi7w6s570IzugdG5miXTCOI7YxywP+
7TmgZ8hd4zaP8SpQxaTfnBO1e50nIgprw6R1DdhDS3+s9yeYEIK7C1lKqd3g9lRd
xvaiG/PTS6j4ThUOfTW88Y59zJzlTxFfpUpSjMh70SBXL6iYtho62iimQY/tVJHC
NZmCKqzdsC7n7zYQZlX+DD6rg1JrJxtZkBg6DFy+2ER1Ejjt6YxUuLUMOURjOZdD
Nm6/WH9J3QXsRhUmp8A85GP7UApN8aoDQsotw8gd4a6fddwLL+b4ZNFT+7x4Uqtc
d9/a+tflpMwbmSUCkvElvUjZ65dOwQeCu8kOkZz6CMUkzd2DPHb+Oi//AL4xB/6b
GoG6dfp2mU/3QDpm1tDmdl3os4zwxAvR0+7x9kv/gLP8m/IbnesZgAx5Yjaqr+Sb
USHzgEepl+TjkU5ZOGLWz0b9peVOQ+2Zss+Fh8t+orrfde+lhOhW/Llv8DI6rjA/
Q0LXOzG0coxTIpv+mG3kr5NvmABySAMifrjJgTiIkI6xQiZZMfIyGjwbOcVaPh9A
XL5qf9JwNLFIiFVQaZnuqj4JQGhYT065kR7t4MESpR5crTM64BnpcNW3ZcPnBCEn
0MivaboXPsItnxbQrXfMik6m7is0fq4Ky6XUeF+lGJ/va8ae+QNs6EiW7oUqGIX9
bvFXVwMPEmJjwq5lQPPriXXAEp3c6w06dtGsDJWFOR+1Qdv5Dr19dt0PowAN2KzZ
jyFB3KbuRUgm3ihHQVF7NGbeEnooG3nXq0epPiXAHZF7Qw/MABCjYRutR+n9I0S6
PmKCXtFqQ2WhKFczNQeJGLcJb9Sgat96YlS1IVp+w1ED75ls7jCcIRLLBGTQaNoC
Rt+2dICO6tiijBG9bGuC8fGBnKLTBbUubS6/7zEcpNfEK/nGaZ59xZf10UAvfnlG
FAvivBQKvLkVEA0b7lWnoOxUJHYUngdYm894cIG+L8tK6ner/nL6nyObXGvQQsNO
0TvRWZkn5s8OKZsVhoqOvomlEuaskliL6JvMu01eyA9vbFJmvZr39TNBZy6QwiM1
Y6j0YAU6ZVfRvDmk3ScB1zg0RD/osSsU2h24DJltKqLZWUHQOji2CfWbov8/LmT0
WDcbvIpJiuEcoOt/ZsnVyKiYUiTz42vNn/CTiyXy8oxSsRZmM3KplR2X2rJ6Jkrx
bF1rWMqZO4XmKkZlEH+MkzSCgfaGYxycmv2418CvXx741VBozeLv3BCK9l1SXj90
uTZ2FJ8PwgUWvF/IxEFeccBs0fGsfV/xFvFus3i6aBRVmystk2d0Leqs9ZaiZ3iK
RPi2J2DC7lDFwsvWqcdc511mk6oKlsuxbwAv3EBedOYLF5tNLmFUkP5lvOaIfCCi
/EL2iRtOjJcQrdk7VqO8FlTpz7ODo80/mWbNJzVXuQvldesaZto1ZXXMtwNXb6gh
SfgtcMI+FbMMB0lqhpw8iDZ3D0oQmtfmoEakx8qsVa9SlZDHeEgKmbVha4KuwWXh
ZIJ6p/s0CWe01FPLr6UxGVCfxCXVrFlmyWsd/yfSmPfca0gUGrEjvtZBgUDG44lz
47mTqDZAWyuNfdSUJ03fb2oW5HZLel7wEGLBZnEH6i5VfK2Kgc7WmLdGJYu5KbsP
2cF/wNOxeX7UVKIhjt0+kZED+ySt5PA5oyzkCWmtPB9xkaTugBJS5dFe/ZRPGv8E
+OPIFvTxPZjsc2q/GwlRJnX47ETNTe0e9HGJQDPUvdIa/aHhYate02N6LhAqNKcY
aULF1At593emVFmTpe0mkB7ByKrfK7HvQBm29JH0gsYQortzQnvaXVkJnNPd1hxc
d8/N112H0pGpogt1NjjdVcV3etNhUAxFhdtZjCWevzJHz24THJM4OzYUGL46HAxQ
u9z3XKt6WtqgI0n91Kf23U7viN7ieCjcPZ9dp6mYGPutM4yOmUaCsFdN4iTLgp1J
GACQn6jDL4p4vMMH1tgVVBcfdLILX0m9M+sVIdkqB7fHFd1oL9OBDVQw0rLQN3KZ
w1AjTAXxjvLOWJ6zyEmF6daw1S7fDO4QrIpZq+9ieMFjQpoyw9gXrmAP4rnBkGUy
Xea7W6bx5D56Q7RZqofo7qhkLP+T0Kkb2zo/8amhItIIJ2OWnWMQTA6N8jCaJaiP
+F2x6fCEHKg5BGCsNLyLNbKNIdPzJnaXUXUdpPE+FSnasTbTBfVzs19M2EklJ+Lj
EY+bFTikbr2Y2AeXjW7aocoDQvGf4wiL8f2AK9tl8wxka4I2zXy7qjH/PeocKeLB
kAx4nonGuZNJEAP9Fis/IJbYi4sffsdOhQKu5aDShTkor9N5aDV1ah222SHRhIuO
6UJ3cvHLKiQH4lvrZqDdUasc81XbtYUgWlOZzjBwAyZyJO97biqzbqOt7IM3nnCT
1x9VVPuMGR6WJSHTtH/tKS3Xe9c8BL8zFZ4cmr7EkI27RXdY9/fi3bxohG5Mr3DB
K3/WyrSrgWN6YdX84SQK3fkY8NemAMu2TWeTYBsj3/qYPm82S3MRs5b8Szu02CHR
l3vTOe6PXUmGtP+rxOB8GJtaSAc+fWKGlHkvsqo5QxwIxI2YD+7ntVmd9UH4/+AS
QL6GUCW59Vx0hb+FY8y2xdHQzhk0btQBLPxfIrN0B1JyDvwyFMTLgoo9NTEnNOqm
Fj1seSolTanL/Ex2zz+dtg==
`protect END_PROTECTED
