`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
T3FfzPxpvuQRU/ZzMvXfXRl6dfEukEdNbw+ZlMjafHsCzjccVkGDIiM/TIlFQ5Hm
bj2eQNyMT7aLVTjsxmmLxsJ8Wk3TnDUEUarEY50t6CiDv/OqJm32XQ7z6IGy8bxs
VY8yZcYNt2FXIhKM5hEY2HwN7Jyfj6rxXk05FsrsvepPcR+gt55kBXQo0AoCEXKK
FcufRAxvaQ4n9s7nEl5RHu0pN+afBVvsokfgps4WbAW9ZVyW5JWmwVEYRp2/k6ds
zR69niEL9MDTYZ9/uvWeS1AYzMh1L0UaNf1qufnpa5mYSKGDL9Xrv9uP8HSN+724
nGH3gHguMkrUxNGl3jlUqSwXYrIpeJn9CSLRM2ATcFixZ6U1f1Il35qzNIVY1BTm
XuQgJe5cCpNks0GXbT2ej+m8lOjfbSYKeYarfjoJCTHn9jORXutsy5Z6EXbqKFms
yeLtiKuSW3KDQOnAyqiaABls828yHvvnYWGpsXl41rDahAJpcFFmThJQAehKQQ9C
+Ft1508j/HTccmVcEH/b+HYHNRsyj6/jcRZ16NO22zwPqlKOE/RrqLvyVf2oj5cx
S7Hy99Kl62VdLVqrEuD/8l0ISotG+nyk9NoyO5iOyEM4btFC/R1ij75ORreQUkrl
gvNXYQp89wd4Rr2HKwM+NqVFMTPcxZzpqaBwlkTBs/QP58xEomfheghU1Gbpf+FU
x999RM8oVStceCjGZE5PPJcSu6Z5mXkcZxbsBb/EuAYPTFF4/W3pSKahr1V0/+go
szCMm3mRtJZ/m1N79NwXeaV1oR96AATRX9+4eJcpHeNYGfr45WQIDqnklk/WmGyQ
8KJo0DaBLegYy/xaUopWTDwxwiWnmr0YdWv78+4bFmlZz3Nng/OJjYe3aL9QSxO5
eKhNOR7uLjw3EBMlKTCqV4MEQGcesDoSHkkSsqJGVD8OdDnujyIBDiA7cHrIWNt7
BY3QIKegVwjUxe/LZwcMdNG+OcJ2bY8SrtgElj4mdEHuMARpEm7bc7X0/8yxZPeY
8arU3WMDTLvjkJME0tz6bCXTbJQTF8QJb1wmVa88u2wwl+HsraeX/3HAM7h78Xv9
i4epv/nbyRROSF8rUbCIL0HjQM9izWP5k1rK2ivTmKT4J5EWlZtxLwwcJqjYum8N
4uxwn+EPv08STet9a1J1+weTotDna+B6pqQX98kLg7mKkGfbCVrdpdtQr6SMBfaR
FIzgwvomhUooh6GALTDQRTRNJwtsNuT1BvkmDNXVrxSP4HNMWQy7Q/KUb9IvtyQj
81/Kwc//YYKio+P2qu4GeCzijbjFEGSOHFt6xqNxhyG60jr0S6yDMP8rxWPxvkHI
XEff1874keupI81wqLA5pBoNwrDCi67oO9z9DY1IuM9+fO5H2GDPxzllBX8tT+hl
YXgupL+TSIqZzhCFKt23A3oYE91lN0MY2Lo0aTc7g7KnFx7SKUscwm8+i3TWsZXG
V2cLsWwtzVil5AxRSxHx3BwzKmlOccd5CA+c03p8ZiRtmgSXaGBg2grMev5VPlBe
GTa9aC9z0bmBDMeHduVIoQ3m3JmtA09fOL6jGfr5RHoM7Leix5jZa4k9qmpttV/P
Lj/01cPxysWQ3KkUlAfUPthcYpN8xsMQoP0OGOpcGonSdAoqqt1S5HWe4wrDT5tX
BsVzW+jomW5p8vdjG5DgYkSiWCtdVooq84qUsHLZvu1fsGM76oTzwM3bgw223xW/
FAX4r08bvc5jC3vQmEswrBnzsD9YlUJVU2lD2bV/zl+y0kb6IVuYNeIScdfxmq9k
5+QAFhDVaxiUeyC4AP3CnvS3BaEQE8e0I3oN09d7DZW/cQBHDPWfNBu6jXfof9c8
5sVQfCaCIbYTAlwiPFvKED9mniT/p0++c7o4MiZWzyjBAVCVjIjlpjdMKT3JErHU
XCueSJ+rh50Jz5o5H5wsw5ZTbJReIE+v0LgHf7mNauZoCcUIlmZI0RDjut7VUW3b
lVwt+OBf9WZqwRw3OggmGIFjYX0+U5r9no94TdP2ww6FncuM9AF3NgVLMM3fGU2P
pTmitblb0+xfHLNL5Jeo2e1m4s0l77eym5oNLX/Pbon0u4A2JpyhJRtTZKhb7KHd
nUO5mfABbZhzTj16d4g8TZnqvWLb1jHZe0G8IbfmZGZ8J3C0pHH+RIEBbuIpINFg
nMiIR3S1UdxUY3jN3XRcPZWV0CAzgulyZs8HdWq9843GNVEsvy5NCb8GjuPRQnd2
ZTByc5H7xoA3Wz4M2zlEVSYZFZg+WtYA+ZyLtZ4Ln0p/dAeI4shfhX3HXQmKFt21
wesAlO9HjYigv6XkWGR87HjjROJTN+4H58ZFlzBAY5WeLIybEzbfz5UxKxKKfhNt
eh+ETX4UNunPa2Elnaq+JYvX2IXcFEtrTtSexRFAU9r8uIc9vb8uWU07YA+20l5K
nkT9H1bf5V8mtXihwriqpAZLFThuht4DxHMuNLQs0qgmCUbnrroJL6vQ5triWZHP
HyRWontOVEp/VpNBmCj9r30pWqZk73fn8hhpn1hmBwZWClXaFPM0XYuVDJ9zrW9A
YsO5EQdImf19oL/lBsE5r5Vbg0xOfP1vyxtirM3/PadB/yLzBlUxV2HlBhbnGpQI
DsosqCpJh5YGbbQ9bbCKF5WXcx/5vYrqnPPS3jHabEXHM1xpglU2XL99xMhqC7bB
XfG9ii4yfu8zsA6sIw6PCI7I4bHX1m9ZrnkF7rQiX/K3iFyfYRg9f05Il/LU0u4f
Jz6T1HzvP0pKYCjVk5WXpsMbN5nOlwAI4Kd4/rvTLEvivoffP6Axnd6r5msrT10v
r1MSCN+9BHAUK+F47ty/BbX/IhWH/uGdGuTXOBIAo59kPJvUCAWoX5dnkckL9Dap
VRy8+8jmftRhbt1UyDWWRGFoBeMWox8RxMYXfF5e0Qwu7kLKaqqlMEbLVTvfLp4e
1+VqFz9kVVB4RkjViLovXCeaUUG8sj5ENL0WBD/DyBZW1yNW+A4fpn4mJLsdD2bw
j6ik26phFspaGD/1W8SN0keloFjfbjZq4iTCXhhGVGUn9x8NqBw5WV36cQmgljgc
0QLa2U4GZ+GTy6fCv4wQ3/PUAAk6TOf20uvdcxMIIvmN6IJSZuRZbHZgBW9mt7jl
kvxK/t4iCx1ExsHmgQUgx0b6PAUEeYBpymXA2VS0fzzUO4GItAGd0ptl2EdGVOGO
DiNiCu7NGC6u5mo9CV2B8yjSR3WvWqjLjQ2BF0D8ShHZBSNKGXIlVaK5nuS8tUWQ
ao5jyxLESaSXUwLt+uu8smr6w7O96FuT/pVDxFnWCbF3PEsyPAHUwm78CccGgwA8
MQtlbp/HEPr5UDQbvYRJx88ZoVM9DHuWa8j+Pv3OIl0LJ+bkSGCSbEvlLVb/4mQQ
RVXF8X3GFnFAxnKton1TW45hpZuQ7tHmR5Ala/eMbBmjTVUzw3Bk9jsrhs/+njZe
RyHdqvnjNh1CwH6xbBLYUki/dfvc/lP0doSdOSPttjHTM5H5LT7Tpk15NRXu+oJm
fr7JzCI6Bs9rZT8LBeYRWDwDrjTIw1B2IcKWnLXvZ436be7xNQbBi3I23MfQq5PJ
Ganr/o4lnwVxU0LYmNeIuR3mu2bIetyOOMaB3snwI+CYTNLfBKbZ39q29IW5Dnbd
Cvpt00d40S162rjE91yJYmkrCFGvj4O+xEJDrm4sFe8lIUdJ45oTAz3WE/GnrbhN
ez5/+0q+0i7fhZTK1MXnLYL7jQ9Mx7WFdXZ7HLihYnhHNLXrxl5PWak1dUiCmMcv
1TmX9g77vTXcgkgw9GsTh0ZbEZ1xCr1nq7hCJ502DgKFScdoCiffvg0+wCMCjw4Q
Dmkf5ycixh1l7ewqDWSAo6yYdu1tyBH/HvxpjfGIChFKakDJbEJOtmFyjsBKBZpe
cDkRM/aHfX6DjVrWqjPrJiTVZuKiyLR/8Dn3nu8/2ee0ETqRJMz4ZGzGnw28UqsS
ADkh1RGrSA1CkDJGpij3Wf3epxFXDN7SxRtLVKt3YBBtkyTm9Vx4KmeDaQYfjPfy
XGkTZ7DYql8uJfmvr4Qw/YdRgzci8XX8xobzHpjStvMlbGqM2Vong+ABzTr4OKMd
veu45ouljbHwluDhlA7JeJ1g2/Bpb0r4287CXaboIojBdfVPz4Lk/Fiz7OUzsaTY
vxvLbkJ+r+FAWcHs6T3CexCi17rMMWsFnE3rGw9DeWlyFavwfw2+fbzfFPK4zH7B
y5YD1bJrmq+P6N4rZWTq/CM/eyaRUUVqX+uW5mlFwk6fI43LFaFIABFEVKVDk2mD
qBaB1AJK+26t5De2zpQkrycSiS2yAN7kmUTqPYfsI2LSGnEB6A/DQGGtej5DguXc
3KPoBZJ5z9rJdDngd8uSbKrLYbxaJ7venfK+S8ifdBpbp71NJ7ReouCuwm6ehPZy
5PDfreT1AGtuhu9nxavnI4NYk/lmGODrK2t8hhhZSUvhjZ7vv3My3iccHZSViQ+w
d3Kgd/jCI+zc9XKXQQcN+gbME35McHSHHe18fuuJTHhbWgrCEhulL5iT4qOTbnzW
AuV+pbwLzCCFiyHkzkw/9VVvCeX+RO1x+lPMf8yuClZFkWqKdb7lMPTWHiQZAH7R
Xh2J8UwLx3NCKfIEmOjogTqlE+6k8yDUsOIguWmw/rT4pazhX92zSyBArGZwCQjW
Btkfrfa9ziJ9poM4tGeEpVah+G0qdNydT6sn6qnfNK9IX2E/TMApr0Jaj47jZh7F
hreQtQ/vySLsBcC2K+KwEtulL77Cmsjr0oLew0XV7J32syKKgYUIhtdkhmm0VwbD
4XXtcVHgHFcSzLUbU3gyJI4BquEl7FctgmrUCHz+GcjcR5Sl7ppnU6hS5guklSdj
HbAWaxifYdbcsNId2Fl0mt6c9bbO8hT53nug9fluzA1GYyzcJkUFNtySsp3+FM++
oedQymKnAZ/AegSFyUIRE2VA1hNidU8YLZyv5G4az68heSoOvfTIb81jH/1AaRTK
2qqciqcntIVDhEOIQudvr02JbU9WZOu3WQSe+IoR7eIVAKuNzOa7QkW8NV9Yn8H1
3Kun8yj5RZyqKhyiH6TQYQ==
`protect END_PROTECTED
