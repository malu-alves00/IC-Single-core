`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JqCd0rGoL6vBlsbOuy+Pgl9JVkEc7WIKnvzI5TPkWULmj5b+ngiqykTVFEPBYxp6
msZgA547/Z4GdRGnofWRACcUnPpv+z8qLDf5Ridh3r6cq1633lTypU2ARlUe077C
oSiMRfnvBP1CLfxBZk0gvAhayIwpDAJ7sVT3lGIEyjbElceLCq7YWIqoiGrkZ+3i
TBqP5uQSf21xY2c5heVcE3Oo7zwBXA3swprGh8fzQFhg7H+uOSoZVhTqcHRqcDst
PaphDXIWdao7uN2K2PIT4C9woKcTT7KcyKs+HqhHtOeUIYJyjtjCiJuVw9H73Ih+
B8/ScpqbHEcohu5wteGaO7pppTAyGmcBQriqBBw0w0jSfyJRQw+eyqk1AQ/srOOr
LbtKdv/4YNAUbb9aeZBKUCFDPs/Ogbh/aI+1eTh44YdSFIeKbP5WknCgXGyAdG6y
ybYryCgQMvYqEIw3BoF+x96UUuRhnXBxhT5uxbXPWxgAJtjOsLVVAjbvZWLntyLP
8mynDztWv39l8RtHDqJjBvzK8XzUwzzeDvxbDVSdIRGC2K9IPdusbFul8VDInIsn
i2/cZcFQqjCXAdQpsBGrSaD0r81dzYYZkcf5BxSA5cuvA8wbkQ8Qtl2l0map8gZ+
kn9jKxsm5/EIrAzWGDKM5fqV50/H9S0GvN2QH0hJ5K3M8SH76wtlwyliwyZUsQ1B
zGyb6Pqg7s59k8VIEdCmeeVPiVNm5BVE/8BgG8+q34EMhqYrzfhyxLajRDnCsUG6
UfVxuxzL9kBlNSDSRootjdBazn9vaoWp9896c8UJ+OyjdgRakh+TX/iy5AflX4Ss
A6bYOeVbToCyMdePgg7pD9odO7qcLCX3c73SRw0W5J9c7VFOHUiAfI27NHB2/Ekk
KXJCDopj12Tcfk7WnVHd+5MrYQvD3mY4tGpYxSV5DrUVu5lN4hMq9K4k/qx3xaku
0qWn7vvoQQHjjTMA+grxTWjy6UuD8opMY5xwRdQs6vUgeExAgy0jsJcFikqO5xF5
h+zoOeN1HKwQbROyWderWLwSl6rwY5ZrgQeLbQZm3uGEz7QxWsRb9wpuDzjE68WR
MfFHzFhU2Xw4UkugZnqipR8C/e4XImqBZaXoAG/xvJCtZ7Vh2hhrna8tLPuZcGdy
hT/+i7581aXx5OhQoLr0/+2+2z/4AHo/ROW7p8hxdwdlG3lSbjckfgQPWKtK7xWH
or0sUmmfICxB/kG+QfpcdB5VItnbL0ogQRhQoZUVzbbzEKzm5zH6ie58a1kvSbU6
JAiJ/N3z3PUKoHwf9t+zaR/sfl3A/RtU5oia6K8d69P9IRQKyAj5g9gkZIiF+sFw
WBJ7QjlXwNEYbCNimSNVHE+hRasrd/wW4jTSVAr8luU2XWhTFSpORzo0R9eRYy/L
y6Kt+II0rysGijGRl4bqAlDWy9Cd4IFsxZ3/dpYlouCSzl3gITgilT0j4Ns83Y+X
xDqXAgcMVJAFyTgQkSlUygsp8tn3F17A7/jfKelGof3YEs4nk47mO8yh9F49swN/
5UxO7vZqqvYbFtk0P1k4IVUguZ9h69tQUezvrJYoigujZz1R7dEuIut9kamCSLa1
hZz4lOlCpqQYvKk8h5oluU3VLuDn1yGwwQOQVySBH5zr+EEGQcpKRkD3QpiGm4XA
XZM67WBbvdd4QSVZIS4H0ALTZH559K9ny+uwDKY+k3cTQlTx9cNmFFmeQHdwKKi4
ZmLqzK5/BLIrKsOpuA3nI6IWe6FCLO5lCQ8om+Q5C0FWJhiRsTylOBTN+Lfxvw2h
i2zRxMhrZvFL52+iilMJ9pKI+zkoDgUxLnuiqDdKPAAXWr2LAVmVYeUCflyW6qQJ
bIgPVn2hp7GgBBp4nAmokURJoYAQ+yzwcyRS2z6CVMcD0/wv2C1loEv8WcwlKT+x
LZRMtwNNQw86iW4PQKpVOhA8bnnjUS3AtzLlnoGBTt9kukdeCESuIMv6WETOWYwy
7tb5IVVj/aPBIaqRJ/0MWXdVHwqb9GdwoG50eA7KnpVB9ic81AV9jb/s5sipqSe2
Q1/9etzAhUosX7SgMaI3HTCQS7ZFxwfTGaqUkAidP6I8NmoZpUQ65HvEYlFhEodi
4A59ALD0OtDFyIKJwKtu1oehIBdYOPw5HotPv+kIgBUokhhj6y36IksXU9N07kM6
n6DqkzCQWCGASJgGKh58VQQdrbnDppPcr3zn1Uw+qLbgy/c5f1a9DJmZKGoXMGGd
hvXQcQdoEMYwPLGHjC7KhXOGXKb+35g90s3zc6BRccBFkCqz+osXYn4bnr6/iAJq
fSCU32O3j3/N8O7yqFAQPlXBtYdlrTGmthWHdxlKhK7DULRif15fz0HaBamOJjPy
JdRHAgou3hbcwCsKPRl9NINRoPU6jjJh9P6wyD+TgCZSiCxAg8woMeO7pxxipEVL
4IwbtdCT04XRZVaOhJNgo6Cn1VepmU2BB3i6XCDRgU/UBZ/KFh4CF+H0wqhQty76
+Ham/9Dazqldn2SyLlwv4rPKFvwphG8vcIouLMDLlnuon0jKp1Tm47v3oA9QcPzo
473lMIgTUJ3zh7clzO6D+vcNDh+EyAS5vlNshEwz4K52KqVkla5VfBzXwGjVtLLG
FyVHcsqUJWtmog4/h/ko4L1/8M6JFDp3lkKx9JwxwoQZf3bcGttnjKVpV0+/XlZz
z5Pbfu8aVDHc/esCvxXwVKn4PqjSEC3yMmTZgIt046tEYtqp3ApF8fl3KovQcnF0
1GrONpU5pflH8NCJZNtOQJ66JA22uS6LHPLbAE9qEhTxOSHEOZH1gMoyqTFUZXh2
W73Z8G455JngWPpwZyKqtGUxGEv9Smf09HQgGVe8wCM5kiOf1rhSp/XYXwjOP+Gn
rp1+6+K9rmldovEbDzkj1rrYlM9mAyHF6Ge73xC2hIIM8/2C0d/1BpItk+CU9Pnf
uV+i1IBvmZwQjgs3Q7KzqbZgQwQ6gVU8I+ZMTgrbHtHfHWFtu5yGMP9IcFpnPtls
9H9GjeMRsN6Z02L5O3tjSNHBBuKdRBwP9xWUxMNnOpmTDrcf2kzpgZ7TMx0eCPTx
wlgkbmBoP4FT1bb7ZESjDUhnAGSKCp3CctXnXnuoTW70viYVERL8yuv962xbZ2Bo
hUUpL2v61ZeepIyVCGSlncWYF7IyEg0wk8kRZd5rd5i+u7ZM3GTXqoWfdN63Nfdf
KLBAzQSEc7luQB0xnqKMRcF3gLiBcx1NnVeA8qDY8eVRRPT2fXuu9L7oe9Th9uVL
Z1qYGdxK1c3BsYJAbMM/t3aWJtwuNvocBLOolmXJseDMbURiD3F+rl34glXmbAib
g/BVHBFU8z7Qb43lQHOKTjHFpAWw99MrBOlOpNEzcPei3xVpSbnSfaf/lPMaaaZl
WpUoNgfmkqgQnKELyCd35glkDyICoTePJK11MwMn4lSgtA7K+VN30aNuq43nq2QC
g7ghVVi4Hob8Ht3KfDTD/4zJ6YE366IpXqwFlAllDy0ZWiv4EKVihulK65pZj4kP
HIXD+s56Wnl9HnlEiKd/GgbcV6FWNzVYYvB9n+ETAg03RzsYb/Yg87keKdbdxGVU
45K3Hq+zChLg5gpZzxT+FUUUoGE4oXszOCtQ5QP+c67eyzL22f1zNnXw+4OSPsmo
8SeAIdxr0No+g+GACfoD1jxfTU6b/R4Q6XCptMSHDjN9J308ZCzsS56hYhQBz8wC
IoiO5SFLfwJvu5yO03GEmjQ3iEn+r2hMJR/Cc3bVk9qlh3sjGwvMYeQ5/qUt2EXn
bDoeiN0hxW3SJNB2EdV05wvM6KFDDQtiI9QyFKvDP5YGF4ju5rndOZoyxR0QugXg
NmmX6yQ1jjPLOKKhuFzmDIKKpbgKktlnsj9eIS3A4HyzeHPdJJK0GW9beOJO03Fd
EgGPiVNhgRJDpKAyhU0jRv/CgqYpnzFrORaXyhjFemH5GRQPLh2kHp6yDa7cy+GE
2sgw9rrzHoBbeeuYs2NVSR7kkOGCb5wsYZ7ngR61iK8I8lafxXmRLHI6bSmGPTN6
qsRudJjSEVO9ZQ3cajaSoAp0BdNUUq8CozKK+/7JNuQjzox+SFm4yGqeCF5wEsTo
HIDsdpKcChELHwAvrqfMIadY6IQhjmgFhkNaQwOMgoaZ1DFC72TF8GgcqUsxWXv7
K974h+fQsz7iP4mIU6NTKuZzbk7gaz8yKLKIxgXHSXoz+hKxQ/KvBHdR0P0Dp8C3
JG7owJYb3knuS3MLU6uQnnZDPMLF3RuraHTy1QWNcQw5VY88ZaCqqsH+Mzktqxjw
iPzjtkbg4zT1u2t2L9F+BaWOKOlnlXwPrMgGPC4mVqSqqZHZZNqrpEpYPfVPHDFx
bq9CeWaKTqkm6Pk5/4QPciFA4yCAmF1XLvTHVbgCazWjy1X5Nu4DObk35UNHUxN1
CXjfDRUlRgxsJ6QEn4wkqDRhI1ktK5CwN+AKEJ+Z7EPmf4agW1GKNint3CoJeOAC
O6LF9M5eCG63q1zOi52xES8YqYKabnzBsT0We+uMj3j+LDHYfJL6GPWFRduKikLK
VrnciK2glaZwKKoF6cYBvEksDCr6ChCjK7zUfiqikoF4UKTQpARVpejU+N6t4n+I
RvthjhZf0nrE52Li3tRpaR9RgYAvuBvtfRiG/LF94m6JS/Bf4QMR7X9t7AZ7bmbC
YNarrB/+utfgYr5BaLKjAk4+tXhqse0g5B3bPM+NOYzghAmH0M+p64tlV9AF8Nl1
w3GGQfkAd7ByWPcBcKcoVO4RSwS4TJ1mr8NZSLj/VOeT9P92XJZCRM2axMhVIXjy
aZj1s4V77ltWj7Cz7qprNBW7KZP738dTXpy8+V7Oxppvx4HIBt1ObU1cecCR3Z+s
RH4d9Z1DcuYQxClDpNL+3edNaQ0l0lgrBvyB6grDUa5DXCdrsR6FctxrlElNDa2v
TohMsv3zSfMOiBSoKqsYOEdKp/OnmBjd5CHev0KO1wV1BP9eudWmbm+MxFrMlgi6
DP9EclSrEnoe5+PlTb2JCKKs+AonTEqf3KPYZKZpAjAYzH7Q6xhlvedqWce5jzjz
wjiuioIg3F5UAnGydNaK7K8WkBNNWC94fRrOAiKvrbE5K/Zje7nlrOB2Z5yEBu4u
It2ltrgfYoo91yPT0dWYCHkSgkgN7vdP43dd+82ptCV3noYATBTT1L8UIPSxLk+P
nLn0HtfOmT/IC9XHq65RuzdRQ+LtRdjIEpVba7y7/disOFC4DEhAYaYj53asqD7x
W6vFtxiwmvOOEtBn4Va5xwfnMTb6pGDA0Zhm27FJX/yEDuAEb5Ai/IiQK711YmWC
Nck1i159WGNDbT61s2ycofYUIOWUAPG5WOEMhmak80P3miZTjGngGyH7yMqn/QYL
zF4iibcsWF7C4LMF/AJ0vKJz+FbVgztpOadrOd2gE8iGZ+68Xiw1a17vQBTqKjLJ
LEgMeQPNnCu/D3Fxz8AdMWfG2s3+5x0EUZfjADtv100mWu2YZekXT/WdI0CJ9VNt
oqS349yY0nTPIVWc6QoELk0w2K6mUBIo2/1jDTlxMNMyIyAP3IY1dOeLrPjlPWh3
aZvoMhfVdVSrKmOCFjH7/w+6kyva21ySSYuZc8ilzI8BuZKADQGyy8r+JESiwscV
fdeCE7DuER8Ygte1D8ItCylqn6+VkgEryg8TZnqPlOPMo04sqaB7ow2PBf1YsSLR
7mdXw5gxTsUfFlOTnocCEQlb6ZR0ukPQ6Oi48qe0amrRbvE4UhJnhpERLAsYCmfk
siGOOP/Cmdi1GtJziQ8ZFIU34DynS8nupUpnNz0BepOHsqN3zY/Rkh1ZXg/ImWYx
6GloZFjiGoq7f/BMxEwldvdN5ltbJ8d9hEqYOCbxiZLFA18auEW6Vt/B/HPfoONg
Wu9KHwxs5cz7W0DI2osLXxbAR6DuqQpxrrBUsIKTk/N1Gxe7w+1BjEx8JB49YW5l
Tg3BLYc9dGqI7LxHzUkdJHfQAFuL342N+UVMCsjAgMcH//cbvzdtLR58N4Go6m0d
ctE/lcI3Y6Evkapae0sStKixf9Jtrtz/4okBC/l955kj6LV6hoz5XRLrmah716Yo
+cgMthHEghGG+qMFGGdAz04PvzXYYVCNP7e2oFWZYffvZ0EUAmodYJcfk5RbPMXW
xmgJoHkX1qcyT6jl/ewropIWJIBizCBnSaa40JbJKKcF8nwKNBVf5cVXxrtf6SJH
fN+lNOaq56aur6oqbP0ysCgnmYEH+mdZqB9y5fywha9aIo7CBtMH4YTT9XmqCIMs
DQc7Crzgmr/W3092eym+aC6NBAIMnS5nAONHyjgxZnI5coou2+bq6d2mnk3JvWoG
lJJEEt17Y+gz/FPYKw7zolNav/C5VVQ+hVMc7dyu27Xgu9Vyeqn0cjzWPTCciiWf
48tZFhfNe/j5QuLsoxKoPK7WvfTWEUGuP6AOHICvkp2FwNehmITdU0pVhHrNQ2GW
2bs7dyszv/wsOdKDEsbVNG2Da6rbR4AEpmPiRx4vmzT6XqQoCIguH6grI5Gf2i09
9z+lgmpwsucVQaRmssitBFmWOeag/D/1v4lZwzvrFEQTkRIhEz7fb5FjoXGsgFlh
2plFpXfh8SlD/RGUjcQw0WUyLePNuVitGj5+qRtDR7oOuOSpDZmQbzLnp/CqlRl/
f5mauEOxbPpZjpd/UxbW3smIJevkmBOYtpG5omyOmivZsQKrzCOO05XsFTOMh+Ml
fclbitiPNaPoGCVKjx7BKsFMikYjJP1Npf8+jbwLBq0Euazj702gAOFDxBgdz5v5
LexkPh/t/zQIDM6Hxhtb3bbHhtz8YAtn1uxEWw0sjKVD1DOde3Ad2nXvbgelGt40
BYwCaCB9f6i2pHbxSwG1eLMmN7ifVA8urZtqZ+r35MCiG2LO5k62Z7YMVMEoEW9I
FCmKhFVAQGvGcnzB6LqQ+jy2WZUYyNdw/NPfGYtaH4UYLmRlmJK910cj3yMtCW0+
cGI2/G23NmfiAAXlv53ugZQcRqmLHKsQj1Nt9QZcaeBQ10byrCrORglVeT4oZm6T
dCBDfMXdpfIicNCFfpYAOL3UyP2nqzGNIDdNtTV5dwoAzOulX0nveca57v04SoqX
wis7D946IyUi3m72Wot/W31/8PA29N6J3lqkiB9HRorKZa2sax2D8oAD/HmNdLb0
heh+JSyzqhVwNJ8GxO4rlq+oVpfqNir4n1kPcgvAYra9YY9r5xJzS3I+VHfUtbaG
0JyGIIhLE11w21ebuou4Nqwf8x7wGbKBK0bq7OlEUWl+AERQ2tT0U4f1HjZr5VR7
SAWdGAJkLU2Fjzt6+A8hqbiB9kqX4sZaw1Nyn8pXxbUZ3b0WquQJJqb1kTxpqbY1
Oryoxv9RseBLfaj+OERmWbLJ16fEnvGAr7hQxO6nmHdAd2moNB1xmh9C2NtUQF2+
F4cEi6HwRBAnuG0aubSNNak9s9ghfy6hoGHho2Us+HIvL6s4txY9Cymetsv6dw9R
WkpdTQ8PUZrPX5ZqDJxazPRIttrOp/vBhM5Kq5JCgqbLrdHriIH5dvmqasxgQUDh
ZcLb7v37DJNOBXYTFITv2dbfj5ILn477PMd0VRERTtMfPltSQIjkoJ9cz9j1drYA
xb0H/hpEWlq8M+UZyM3hBr8epTVBTMxK53ra3yUeu4C+0MCej4Gr3JGYmyGA8zBG
TCWoqTKH1Xiw7z01SW0J3ULTLZ5zzhL0zEzl5XTaWHoB+G4IVXIMya1jGlXQNEZT
XVyLaZPxp289Bc2W6Jv3niyF0L9E3K5U60B7/dFVEyHqoPNzIcz+92c3TbBhPfmj
Y5UdxhWMatHn6O/MTKyqOOrHEE4WGkN3db3jDiaYaXOQN14x/VICuA+d+eSC3gef
cOKXLN5sDKFhp6kE87q7DmmDpuXCM8pFUMHwXg7KpOZahc2rAbXgNQjmdCGm22Z3
406oYi3VPZANL/S4mZe1jkTPns1gyp4/QhQcQR8TJn/7BY5zHwR0D8A258DvBwP+
BU2B6xKe9O1J+BKGp4aFfcNPsDV9vLcuUcquQhwkfaNmX0OvQLNioeq2t0VrfAJX
UBPu9iBbgrCwVotICss2UUwBmw3kYXD0qn2thvoeasFqWT2IHaeeNy3qaXBsuAG1
JCpBVQ6t1udoyYnGhrqbR2SH4gK48UKe52oT2RQLUB5sU0wVPLNSYmwLRjlT4giJ
zYaG5bI4y/he8aClwQq7mQMsikjY3nD0tGQbh8H+/w3ws9U1vk1isTtfl4r1zmHC
t43swYMsghYuL/ADFhvq8akt8Laf18mOdDpW2ZrjH/zQ/Vnsp9JWDcGRs0dwKOQk
FqXkLkc2WzihEnBZJQeSSlirmmdRRtyn3QbSMT4QhywrqnH+TAiaOBoZxZb9S2vm
v5N2718y+k+8YWtpnO78tIBGHfI2JwvOSFKGid1/5Hf5eKMguzls84j9xE+a+jdd
MJwpNTwP7wlNBkpCS8TIsP/yTRGu7V5ifWOdk2TCXgAs01exUAkuGGA6mQxu0ae/
bKb7tmHW2nF52kDdbJkqZmKaU11LRsp3rivb8DnweugBfBM3ptaB7bp6KOaL6KLw
9H09r4JTag289z7XjsRtJ+oR7w7LGWkbBNH//ZdFLqj1xxf99bpbzCileXOxdrFx
rBYQ9c+63WEVwl0kVAm201ydMHpE188m6TFk0afUyoSqbJQmPwj7E3axdNlI3ImO
zOsc1/9hfjn3FTw36AithUWW6fRnNDqpoW1V/HwDjdvhi0HBUHJ68LqHhrxkDgF1
9z2Gvv9ba1qDpmS7ZA5k+Nz3iDHGIl9sWY2MRLYnRboLBYqgicYuMWCObEnp226F
Z1+mZsyWnGZR5WLtWfQQ9fSxBO2OHBsB6z8mnESBfHyAmFzWDKf8jkUiZN3EW3ZL
K7PDG2lLwwNr28cNkvJO7tnDSgYcLG0NTRvEhmFG3WMaRwVQX80VQezZmvLfXquX
X9LMmznLBJ10hZL9+4hWBdlCaTpHEDrnpp+qFhZHrWpJUqN7Az/66MPThlRsQhqk
xEMvDQ2m/AsJ2viVPedBtX7kt06565eyEhRbvTqylX/z0DMsQweAn9pshJ3138m9
Xm/TwVFilKkP4MbfiWJ5u6i4yuHp6a/VZYoIGaOGMpRFSaa6pEdnAvtj+3T6C8Hx
H/MwBLKcaeSu+3GqwwPv314iDtrddj6dju6sKJ+v6MFtJKH4MI3Dur7byd6dWS6p
ZZtS3wCUjrX0+uYj/1DSdAXcP92nXDpEwxtuTy4iEx3d1glXORo1TNTjuMk/aGPO
Ap2P8DeUJPxEJlm6Zp9+H/J19BeKdyFsTQeWjb1ZFdjL8vcbHAXGZL8fI0Jzzapn
IMrPL6zp7mMHpMQksg4a4GfTm60x6/01mDP6VG2dWQ2DJvUZJWqtZ5ZvkInfVeKr
`protect END_PROTECTED
