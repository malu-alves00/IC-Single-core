`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TiApwcZWGeqmzk6mMeGUiAw12u7CqTGiWa2ofm3lXcg8gAcpI/i6bSbPeYccKKN1
eu3TaTDv9L4isFK1edCD28/fuNBx2YV3XZWAYNsoNub+qRHm8oIjcWHyPV4L2C/h
HpaH5W4iATMi8UI6NjbLXYg4G5ZjqPeLKDqCCcXOUYhZ0XghBh205jQ1HjIMKa1f
catMUxHjSfKRb9ovVEULAWILKdUf7l96gASzg1VWjNEhWDqLMQv8o9chSyBPcoJd
sQUQ1WU6aObEy0HAz/gagCOHiY4zfHjx9m+NPH1b/CzAipwZHYc80ytCLPC2D/rM
Gu6XLjpgTBGEp6u2PuA4LKQwf2/jaF4PD64EwcvuFRNBJgOom91E0PLNL6Mt8qKE
rbRj9YdU5qfFRofJo5vMKv8Ala0UqrTFo4O59S6lGIRPXYeknsF2SHJbXj7xu8/C
XNBIpb8lgSQlpsk0Rg6idbOCOqgKZwm3CHAxY3UXHnWG4ERJ1wTq/f3BMYqUluvt
YiDrrGCgmb3Gui618qEEBtleJd7r9AIms8o1LnbYuuL0eJFBJWrh2HW8d1uVCTmH
wZcC9zmi2bd8dXkIF74xHjFhB8DV6kX8QWhZUtx7mjbUu7RL21WXbCa9VxtQH8wN
yVrezeSGmxvtFTe20XbPeIJyvOJczZ++lw4B4oAy9HW7TWV97LCZaN0Qcy0yLcue
Cc9nhkkd5EsSb8DEMRCPgfbX9aHGLRpAFjvEi3fJciMN/XwI57/9HVT49iQAbYbT
5jzPyfpORF9Yt/YLfL6yDVFb1aJhotaPJKjUJ9ojqSZFhuyRSIk4lLMJCEezzIEp
CGs96S2i0ZHHLc+N23wJ/s2c2T2nF8xeUenUlCZt7qh/ukemEWRXTbEv/uuUgw9X
a6HjqERDfqoZNp6HWnkVtkkU2KMQVOxFQbWdvJyqB4w3I3U9tl2UabqQl8rSVXpJ
IAPC0PSkt8qbu5qQpxyYbdSJeQA1r3Bmia5jki32fTFx09Ghtn3hQydXtQy6EwhB
+0kssNOCWGShBAmEZd6JUuAcrKPkGXd+d2urGZAdFNpqlZ0cPAnipkfI86PmXYb4
kfhTTPbl6wf0x2LphIWS/g1uuImdZJN8y5PAljw2NdLcoSW0bKdVffNvPLxm4amR
uuH1N9W8sZuMwGAiWf4v1jU0lxzGQcCASrGi3MYp6LnrJL6l97GCmUZrxsIGtBnM
uB86q3IT8XW9AhbnQYXEI4c/gGsm6X5bwOZGkVMeDwLVyrQirX4EnF7fvy16j9Je
wdLX/EWKqljzv36Z/u6bOz5ayOjlgV569KpD/iK0qlbq4a8DA53jbfTBYquCPi6d
v5KUlqVBdxxiJ1U1n2uCpQNA3g1o7vSoqhQoPmYu0cqdIrL1xer08F0Ruch/vvPC
S88xZE/gXqx7azsIioMazK/vgkS5PwZ0MOuFo9weCz/8BzM7xxWEssfocNgG4Y5D
0cyfz3hV0BRm2BB96gAl3FUZZiVPEwCNwrvX5qit2mnGvqQ6n31t1sTQV+ZZiT8c
ij4acB4KD3oHRTeKmjHX6gYlsnL/QyKsdJYvyDggPrqosKIjVpQjaUqwOHW5IPt+
CFMO+fLfP6k3uRpbC+Ya33r6UrQ2kaMD8Bo8CAkUR1FjndhagFjhgPV48slsMBah
/4Wmv/tmsScvPt2YtJ4xWvYQdQMYPRxOd3eA5ZP79U6Ne/PUo36Gu4BDP/A8SZwM
dRVWGUzb6CMlSv4wKd5FZOCd9md2nwwcIsVkf36luDmXYx8TbmZjxXtUpZvf19I/
wQjx5k5YBHdbBMWkhvXOifMVSOwzzLIHGF2DDg3S6fcBJzpPUaNKq5nPkfwB83b8
tCrntKbRZd5s0LshPPBLx/a/vNxmASrxfCHVvmWtn40qNSIZAhgS5d0Pf8VwLxk2
NcBZntIePGfcMWbk2O9BYri3kO4Q734T4YQsBRD1BSAFTuZU2n90v8ESPZl0QrOo
02R5eneiyfBFTAQLGGc2aloyj8Xfi52ilJJJKykPSu+DSd4xO/K5uRQgIPqyfa6X
3l8EiZigxvcCPGKsvzsbHy8khc/o/2/T9Km96EYthVq7gLWMLoxpuSZeYxmgDSgO
bDO/z3xXbV0dQmpebu4MAgoBuTxXxX52xXoT8ayGuCRBPx73yBwfWkmygj8El9PJ
JF8/R3OrBVbgGjSgqKpDMUqJK4+svqd1bW4GnPydZZRbUdxyH08vPOlVn+opymsd
qFznALVd9yk3RPfG3tLauj1SJuq2mt+D/oPw40U+cS1SdyH71x75oZ16Z/3uviWv
KWGFKDw63nYBBA5uvs1hl2lvew04TpzRwDLah1BzgtWhRPJeeT5puXV9QjEHMnqS
dKOO2vpcHKE3YupIBkD2sTpMPcVwYjVaoMPJeb7v7LZzTP0LynGbvgGkFxDoaJ4X
22lsMKkibHI0oz+tUelqk8gl9E91cVsZHjN9YVzTFop+JRreZVe3a0QVafjyj8G8
ffYUanC5UwnfDr6gFGsssqWwSJ8Wvh3+vkHXR/+Xe5TFaRtDIRWoqxI5ZUFANTeJ
9ebBgOU4nCZDCyuPr3zmzz5y4Sji7vlzpCjfLHT0HJ/ZpMFYauIzuztzgFL90qJ7
WjRvW4LG2xJDqrH0NYcMcsjzByum/LknLvWYYGtUTZsYW1R1n3a+C9Nb5R9KGMAg
fe8+GWRpa2MnYzUGkT+cmUDgYkBTCg37FYFRkTMwK9L2UuuYMJJcXFgrgd3BLDc4
ANyqo9FrL6aQB+7jcPwrs/KzPAqJGChmbDnpZ+uex9aUqHRbuBbUy1wiiLiTBe0f
vyEnRq9re1gJ1MuUduvH6OpfueoY+FaNiiqTIGdxDBzsV89asLyb/h/4Kp9p9OPc
A1DzQMEVnYYC64jfJYwXu49MKy9SrDoR8Dbl2sph/UDCSzqGeNuPvS9bTvOCXhvF
t98uy9jKvTtut5q0734vD2RrUobzWXKZZSSTOJ3N/MeSA5cMNlf5cQoaN2wKmJNF
cVG7TusA57d9DiHfoFgNf1w6kxP92bHtOKICOBaK+tMiVHG6j/RZuSWSxEIGxzmd
Yzg2LKA7i2xHtkqJotmYXZ6AnsAAPd8T+VB1p3lkJJenHX2BHWofPCXiw1qqLlAq
YEZvx9dDw5ZEUWiqceS43YImKyPa6reBUha4aORzbRjF94Zln5Govq1fs11ZZTxc
dx3mTXPh3vx9DTskp0l7U5+kuRdvq1gGuuZRLFicTP/yKDetzvfFiX/sVkeTFuIF
vnWC1IcxcbTOo+CutoJCCaYnjT+FYcDSzSziz91BaR+HO7C7mvCveGVJkGGVgByE
RGJBcchN7/mMZbxz2o8TsHqvvMWK0Ajry0y97scEuEh7w0vxWy8L4O6sfCO7vlVZ
3iYYPXcqw52hGc8OvHf0rYRA9yarOrjeI+FRe/r9hlNCHXqGLF78gpf5YbeaqL/r
wshY2VXBmVvsjFt3FROmkKDEBs6CcJJahrdUGfyeBU/otupjBEISsHEa3X6lISya
vw7ltQK0aC5JsUhUyTYN0eoT8GIOSQaX9HR5glLzUWhPtVOvBkMrN5/veovV/UQk
UcUwdp3ZxBjp479Y6RhvxtuVR1uMN8V6u7PZCJ7DhZhWjTU79lDRsb8nC6/nUlN4
DE0vNqp7zhaJIhgsoqF0AF/H6mM4ty8s0uoU1bNBUQLg8Ar1T+jr7SuSszCcp8Ki
U8tfFBtZ+yytxFm2DmnUHtymcDUidKHkELU/+bZSdXLJaTdsk4rZuMNN9Pns8tdg
qrQt+LS7yXNOk0orEXmF2AczdvrZwVFTgJ5+SfoSx9vKqHQh/KEE/PwU+nzPYH0Z
eGryfXV0sU3b6pQL+5FsPtACMBFfG/OO+bV+gx9AUP6NHZnO3tHSCgGnq9/dy1cv
NAu+y869L43QvBOfQV4KebSbWa71iJ/TujfHUbNKlYKuloeYG+JRXZIC2mkAipSd
c1KnC3VyY0P89DOpYcKK8GfhrKa+7C0pFO+8ep5Ykxcjxsnj4MxXgGAHwtBlthoS
pkuUdl83R6st2q0VtDrk7YzNKFAg9UnOoEw7KRjEbjKIXBLRQF7U93TNA9kg3uEa
YhWtxPXeBmpOqOos7gPoOWngLgPRF/rgUUkf+bRQfQJxQ5Ktpgz2a7xnIUlLRxQb
couKti09s1Potw5VPsYT8Emwxl5i/lq4R2wxqF5pbg434WXNtcDfU66DwhCFuLAW
j3RpTJ1BU9Q1TBbbO5cc+fNJfeDaKfcTjo7RfJrONW6A9WHxMF3LOya/p+IkQChd
xFDWVhuBhy84uK9L+B4ZNJtaxohGb+TkNaOSRBRoo9VwimQvsJEUCfOK0kQkW51d
GiYc6nCwf6GSfkyEPo433qeIjU+dVtQDcOVEYBnkZtXtN1cm/n0SkxIHl4srNy5e
CU/X5fX7d0UVZUZrqKzsfIbsNiFT944W5FYbK71dOKgJonCroU1J65HKoXjaEkXQ
JsyjbquI9TRwax4Y7x2X6XSNJxpRbAawvdwwf0VOWd1yCH/7z4RHdt2FauyMB0aP
UcnSu2fiPDEuEfaJ7R7KnHFA/AMgaQRX54Kk39HNu6JQyXxCTpimS1KmqPIErgAN
X2irwZoZA5lERmkHRuaK2Bc6nxx8602z1U+24gcQwZuOCPWrG+id0MVmHB+V5uP4
sGQnUC2fRlSm1fObkDdg+BrD2pBSaEvHKmzVIMZUVFs=
`protect END_PROTECTED
