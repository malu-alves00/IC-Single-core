`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zgKaSPjQNePdbd66wd5qzdb50vHSC1B9NcFj9+MLZFqorz5wntstWAi/yak67IP5
v+P0JpE3lNghbnLUwFu5EBlLj4FMb70LwRYCWd6O+Jmw2Sveik/UxjLQCU5TmMDs
v1lszA/SC3hzillSLbFO6jsubzpVoQlVrQ0rHRWtkw2o4Yi5piZXMCTiDkZ3nmz1
CHPTQP9G33FmBTimV+S8s124wHGt7A7fTeJOXKFxouXznH23PvSKUZnFNwvylm5M
8y0yp7/AVuX7sRxX36XaUYaxAlE+jgke98FrUFpMz/WHQ2wHLjJuHhGJgsadhITq
EWsc/peu6F+5DCiEV43aPETKrpnxUxSvmC62B1PdEp343NPGTYrrtGhH30h3qanj
5IK8n3ZgsNqPNwnWVVBFTHgM9BOeDc0/eQ9uctVOC6x1DwZ/l6br/6NugGX+NmuV
9T1wVm9DR9Div3/eHol0fd2OVND6Gf2wb5lqDoa7zHE9kr+QAGwCDcRl6LIFta3K
`protect END_PROTECTED
