`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
o0AybZkf4bpdYFmWbBq59MWNGsDBujNTD1ExItOjPT9X59SFviD5leDcyzKc8rW4
+89Jqrux8pAROWd7394053uUQanRaL5BuJR1RXB6C+EPGxTOwCcUk1nbxd2DyKzF
AjDtqFVriRz0n1ffRYGuBd4rpQZwrh9NQTEn2qbEthXjBWC8IFUOa7JQ8CDtJCB1
HR2n4zLQVpqR2tmSFJBVL7Eiqb9YAeBOlo7bOxo8O35jJ6bqAv69YVY9pRAKc0Vr
3w/hyK7+r/mJC6S2L13ulmhWIGsqAsBKMYK8PqWfi+81jD42kUwwmRXEj0m9KG47
O1rezaVDKtbtkDDl4xWkS3MRRGHTc12HVTX8abrkZKQPGbH7A8AzaoxJPxecbwDV
5+kwHpC4uz0hqtPBKvp+C8/f6iju8ohoZjDa0VW0qfsZoBZ6aOsYA2LXaOj6agU0
N9ErfNoVEd/46lfLKUjoQ4+iJA0Ak2pnl2c23JP2pm8edOpsOcMrI6Fsx/13GZVa
WqGLFyfuw8hscJdad5VSmfFh7iGp36cz881rtWx1oVj0zPzY0pxdquba7g2GJts+
OBjm6vMfANca/Eh1XaHdf6pKJqE8d2+2PpiyYSCU8tF55C/jTlIWjA841zpFDRp/
zU2AaXLeJFEWZ4RVDKw03yOVSCpzBktORqBWdgQnOtssxJSNKckcRoC3FiCrnCee
ZMQz5zoyqr2srZze/TckzlsbKH1SaJeQ0s52Ps21QLQ8JYqo/j2FPTCQnTdIg+/o
2j2/YGI+snGUAousi0HEQY+/qOTX51tOTaVEPIFfgXpKvzw8xO23oHizxiUrudjP
9sCwBKjJc0Tiz9CJX5S4AlAz5iPlu1UZPkI02IESHk+aye9KqswfsXhqSb4Ymf77
uHMgIPMy25niyatLR1vLNziebwnO+Q3zH3paB4Fazf5StdMhuLS0XL8Z1AaCI7lN
WB3jalHdPwHdC20wuf0kDmPAUIiwezvoT7nNUyXK+5QiiaYCIZ8gpmLNsCM3s3OW
YItNNnsjjoXg+w2fm3AHX93X/ZdQla1y+LhTj/J/0pWiPi05zS4a6s44ryJ5Dr0n
+1oNZS0MYdKC9PDTx4ZAhm22CyvLq8fTG/rrFhtx9vpblNQqiGgdTDPJjlI5TUtq
wBOytwmAZk0AeujRLCiaByr7t1YOgPTVDlVsTd/xfec/YbI/GVlAoQ8K+HqTDQGZ
AGpL35m0NLD0+F7JcDqUsw06jO/pA6nJ7JnungQgLYAOwvY5sAvJ0FFdZwkfPmlq
tyF2eURKgHjZD8iSFeBmEp427dNQyJ7eC73am1cmVqkzMo9OmkMuAtXXfWP9a60h
fu6nVNVgrMwkiTCAqaRRqJ5L+dxVVWEihEdkrvmAvlkldLBGrH6seWQ1Sv90G6Rd
/PfgWA0zDfS6N5xrKnCu+UaBPJy9tuSgoah3FSwoWyUXP4C6so1bZQ2NVBvMSAHb
Q2IVN5U5nmDj5Tm2+kEMze6Bl711zOspYbfReJ8vJskjWruf03Toqd+i3dMjBMPr
Mbq8Dzfjoae7wlGHKRPIIn3vIf2YAjgVjq1PM5bpXoF9qRQUt323Ghf7irPpDZcY
QfM/m2+EIGi5HElzhhsgL+kPzGXx+cd/p62ao9e+x3qDAsKpws5U3b2gQVMQL0lT
KN+1EUpcAr4zmadQdXbQQAMMZs6c2UtVuMbx8pcJjHBz/hQsNzfeYyqwEExT2TWD
BGA/vrlAhLIVWnt4AdQhA5xKZdtJACAoIckV4tRS2OxYq6hwjOy77sC0BLheBhoS
1SqcGV4aCzP1wNx/JYMyWDkFp0luKYqcZfro2YLUPL9jyh8aU9NLVVZrTNkMfJqF
ouCTHvKts92d9xfIWPiNVK1XFQzVFlx2qw44MDm0Eubzn8CU+kVE+8fYM4A6H9hL
aze+hZ0uQbNxNymJlG2w6Xrip2gpVpQLBa4Dc0gX4w9dTR6NYVbZSsFBjSrqi5Ns
Kfu6Z5OOxiSYQdM+JpTtKoc9PvlUYo3V+iV7VctqeuijjDYr77LqShDfikJYszfc
XAjljdkAorM8pv/6FCTDCRS2TNDp3YxXJmVargetOKjAR1GF8gX1501kZKOHH/HG
1zE5elAiHHxvLBjgpoMm/rSQuJvsqzofzmYAd43hjv4LkslgZ5H8zfbE31bHMHaA
wPEbVVH77geWRdtm5K3UdY5pBcDSsRIBxBXZuO2PzDEONHgNnNWXged6NMbieavy
z2uFlvv4DhgrD9cBlPjbueSoN+vjbSFKWVTmjfdDU67WqRyq5IYqrannW+vI2hc9
pXGyof48MtJ3ob2hv53+7cFAdGWEd0AoDIY9RCm2qaELUQ84EtAMKfKSyKJDREyG
JvEetsOWcnPUX1e9/8gt/SjYN+nVyL7dycKhDTsenu0xG9IuJ+G3/lHSdpSVNAIA
lKXNNq0KHsAexJThZog785Keae25dXzbj0kxfDaoBmAPwEGGTjH5qMFrMurtr1Tt
vLiEQ1Q7NT7AF1RBIyAUAewkjBQ9TfZ0PIlmN6TdAnYCLfm8Bh0PuqkW/ou9PxvG
eG6UJ9FD5JkYp5oQoVFV8ZZmgqdzbSVZ3z/enRUdYKNHAz21gsD8L2Zw+zcQoxn3
kaQXVjJ5T865RAdXi4nIYzPeCUZ7bQwJrhaNRhMVRXcGHJzIwnkuMRRR7PO2bz9M
itfMUH71aTS2k6EIn7N9svDrzJVnO9PlUfHJ1YVluV6qbrxPp0AVZRBd3Ff9GZdg
6cYNtcs+MFRB6vsw1wIeXou/ic4dI899gRlbFqdoofB3ldbliWtk6GmD85i50IvC
7wtn/8rELOlbjjrc8cKPBB8S2kTALnpg7MnlA8kjm21Su2IjNtS8lCwEBevp1QOg
vkCkVCPs8be0H2Ut47D/REq218nHCvww9KRNRIsw2FMF1MiN0hrNLLo9FAg493bt
glUpo8wgCZ8I2cLLJngvGEtZDufZb0XnU2C/OdeBaEs37OxGda2D/uXxQ68biD+4
01+J9LVof4JglnOKbt3L4+rgL2F9u3T3rZnNYmiYE8sONzmmyWDIf0AWOGcebAPC
qwuvWUdW/BjN/jvNVobCvqCCAYg2p0P6hJrmgUSGeV0vdq6E+UbWOzBE9KoqOoj4
wFIjov166CEflEetu498uV95T7jrt71qeHSryH1BslJxesbxHZ09YwK0hB4bkjhN
wF+R6dJHBVz9Mh5utQZY7lg5Nh0/bLdrstJZt/l0D8lxbKfv6hxbC+2l5lHw3AdQ
cJjDGnn8dEviyN1Cvm9PF7q6vVBXGqB9OyG1BjVzM11FaKsBmpGik3uo7kN7Ri9B
GO/DNdDOuOeCxB1lRmZFsbnZClvF/LyRzh2M3LXWp6qX6vQEtyJXai/wigVS7osC
QOp9/dYRKilztfx+ePIyDHvc2aa3XVcl0Vo6wOfcqzaqEsPTh2wubX3rGlBwonkB
eBgmaF6WG1gEOxbCfuLqAdXVWdlCM+oZmdXvWlPOlpRL+BXAgE/URZNerMJQxfw5
JM+QXk08rBZ9eNaEaPMmTkKuDDuAIG6r8CLJ4UrNusjRML+BT9Bg3NMluoapr0ec
F/ZQfLV0xmDygAcXyCWhtsqzAdJrt1yCmmArf2Ipdt73chwVqRVpV1aIMMu808Xa
w1LN7NN6Yl+3iZBFskjiXQWfQhCGrJhP803mYrQYwQfIokwY4m0luw0jAkI82hCi
45JDrhcxOWbpo+aW9PmZXMqUenOQ0z+FkOl2RhAsE9oKmGF0/TTeZXmCwsoNUGOI
nBR+aVxkMVdotS86AGLOWGv5jYtHYh+GkLkAmlQvTyeJ6oSzImafyYrcMvA509pn
LnSykF2owq2fcb9cJhMzw5Q5t/fOJs1+ucAqxErpG9ub7S6bUfFdMqdBUpgX37Et
ci9VZDFyA77Xj8PNc7AEQq/+xEkaLUGfbjW3XsW61ORWnf0jbwojFShwQl8PIcQI
Fh3v76KP4qMwQQCDT72uqjsVv5Gzl84Unpsp0+u9tLPF/b0xNsRcLNqH18vmjHC9
ovGsp8PdJYecu4FR+6Ld/3zUllUIGQ7CANGqGylmqKnJpZHR+espmh+9A1OowDOn
8cp/GlZnhScv1gu/79fazyxcPbwdrBp6ZZITN1CHSZYHIx93Ok6K2ehyck7m63MT
5MtxvlSIz/ob2W6FjqEDl/4bKUSD7PCKplgrITwtmpifcXbwuunEfynX3gzGOl3+
75H4AK30FmRuCsXHz9JAKiXNIHYXT8et0AM8Kzr+J2xg+AWgf4XKQWv9q5Q+iLcw
Ye8zGgsvUD+R+dGA78jS5hXp1nu8SXSd6rsupRU0ZN88g5p00BTRSkx5MfOZ+gUX
FCFIhXi3tZseUrQByRB1Jctd7AVs0NXca02wSqCXKffuz3ZiV3e09aj5rypfYyEk
jvdO1psR1Kz83JEUiHTeehPulzQUdGIGCuSCCZxzAjVwtM6GBNNt97a/1ug2OsDe
BVsXMs+4hLBN7VYM/l839osJC5/ZcOJFRG3VHBMkx/M4SVpRlFIgHf7asvLTMdjT
RWVoAj2EKKSRwUNJqXTEVa6/9Po36Yd24VXXWRdqxciNpVMOHGC0CYM0OEXfT+N8
NUJEPEfDTPfzJANSvKZbXZHr06ghw1G1lbIjzdpgI4bW6Gb4+O4wyJVckMZkdoiD
d4kfQURwwvb30PAiC+KyapY2GcypaNMvm6AMgLH+WnPsdP90N1lMtR1+TQqFY+tT
Rt4mK0GAY3IN+6wqZa//dXeJHZiuuMmbhlOVkc5VHxz3PU4fgMiVxf+AiWD9iCGJ
FCNX6sKjeT9V7QSjmAocnLfEZzU/IstCOAkOIel5UzyO2k8geSD15Cn7nabqu4RA
escWAr7qsfHk57cZ2nFKU/36OGXFUIj6VF7o5H5XlD6nhfgJsIpVLLdlIOtD+F9Q
MXM12zZuQkaU2+MeVQ7TIMcmhCOrhMdlgyZ50GtMf0iqLlxZdGRqWro48sMsvv9x
tjEFWXq/8SG8j9b4kbGXSa2SeHcYi6Ai8Em7rx3rgbNEqQTtNObfqrzhasXWym7o
ZQvvesV+zRP7xqjG6vCKXsc0cGv+SiGL2CItTJVqsB2pJ2NLcMNQqrMO4gvmOAm+
1ucsTH4QKrFoWCW9PdeCf6hcQUyMRwt+B0LfzcyYY4ToOEqmv1oe+0bdlmg3vk0i
RBLW1QVDT5tNc+0kYuMyU7b7ymj3tpMeXrLRcnb2GBW0ZR944xj0+XisotabLnvA
eI1TCjC2nFmDQOZcsqshQehr88A4gW/K/8EvbhMHFnVtXdHkXKHJvi9al0Yel3mF
rIgFc4psIupPkOe3+0ou1N4Dqd+Ghx94PQkV9mOq4PPg9B0RlNbWKGIx+lf5nnC1
ER4LU2bNwlSXT/dM8LFbRHGKJpYFnJNdvpmuliW3+/ddt2hodbt2hrm1Pu2Qc/zD
9rJ++YSARiroSHZ8NOTS+1Gu9V81/YTa/aU66/D94JyiWa+L7mDVsSB7sB9OK8zJ
KWp3ewz5hhGj8aklMGnT3uZ3sVc1p/hocyGak0BLaRZg6RVcPuNh80tR87QdO5SD
yT9681KfrrKHRMCUtb55CXnczOipPjdvkcBj0nOvSmozse5BRaeYT8hM9VrGCHda
AKTNZqi7nIMqozqma4ov0dEuQQRk5XX3ScUDVIfMwQl+STAHH9+sVE6uipKVlJ7K
N9OwBVWUvb1O5MJIi54TwWKdUQ3PLBxQa35goA/2e3xmzXQupp77XHiAgy4Bjjta
8hdT5hd/1dXaACCTWJ1qByUaVPOQ1iHP9gl9WJfn8J8V0mO8dd8fwJ7mX0RiS/UT
xeLbVE2K0rPYyoIonOCpVBP7NC6azE5/o29xkOHfrOD1FSZA+BPeN9TkrJY3fTAj
Bt82GGSWius4z75p9T5t7rUW3Ve48NuGdBz80q27uXuDiAyx3WKUxMlFo/bjdPjv
JG1woFo04qJNQlWON02ZLWprkClyLMy3DB8cFYj5TMUIH3QHLfx8Uzlu9dZIgH0w
CIdGgl+57h80GnU+qn0SXZSXPnDPbUI4AELiTxeif4DKoBsM7+Y5I557pdNfpCIT
IdvQ+LojmPhjPDy2lAbd8rrud6YP9XlET8wjnP85A+/02BYpCzgj0uZ47/YA1eYT
jYVUavbXZ0EyXr+juGRIVtIdge0n+feb2PT9pIkXusvYFZEp0q9ew0CRQVbQ+L65
2qzrONiCq34xpuw8SbC/H3+ehzOLJNOlZ/XhvirhRS8sGxdMtkJV53qyzhDvvANx
UD/9A68zJzF8U/jAUJ3KBau+Fet1E0SejV7jAcXx4qIO5LSsLaSn9oYc2YZt0aQ7
z6sc3c6/m687BvsbFb3hBdUkFeg0qhFO/YzQTWnnTcH//0w+15kAXCXFruqg5x7O
L48z+ZBWUbFWf1Jn9wun/NnXmvsOssv7TyWvFU+yUKQhyiE+9Vdi3ZIqlOahib+J
G/VaZ+niDSMB2S5Lxo+UcZBHe8x1onUcy9ehuPv1OsqGV5UD1I2hcmvLhqmC/0a1
rFsUaNlxCb5x1X3CtJeauzSf466snn5aoGK205XngWZZA22+CnMA0lZS4BrA5rok
FzzxQRa9iWs11p2VL+Y++6RIHS+Yim6v1lpi0sinUGRqgpeBv8vHuuNZoYtH0Ltx
xn+p4WXUhNaaBf3dT3VmAqBMpSNvdxBu4NpsVpDPOmUZtoVffqZtjo91kT5bwBb7
qV5dRPMmeiQyP0kaFOoF3ipPN5YgMqGu2FlnoRtTyW6sbrhwvHCJ4ycGlLJkFPYk
L23yI3+nkXmJcvYKA6HL628exAUF8SzxXaDNYuPz0rghcEoRpx1gj4mx6f9Y1pbD
/D8AzV8Dui6GGh7HsOxgWZgdYho5b0soVeFz8fxW5DeJCcS1NeTJsR6tq41+tD5Y
brYJ5aEhwEch4XEeP8tDxtljrPgWNgCh3tm0lhLfbjE3eAEgrKqNZOckFVJDCDeE
a0Ns8rajL4An12HdPF6MGjgAKNkOuPIadHo4i8jrkuZRuS9EtIduq3mzOCnhDDfk
vxACLkn9gPOBcYlAV/L5yCet0qIchjSzCMQldpLjsTmvaIy5c11DBTm8WYl+aDjo
XAKv9bMVSDZxrQuHIC0H9aVS66dKd4tlRVjQuPpam/KQTm7mXaq+Mw42I8cTUM9A
uA9Ibmqmz0zobmCgkUapOQJMglo1Ee3LwWGvN/5O+7jYzbf/Y+2Ivns3+NWYRRAz
MZ3En7g52hi/5xmUEjYRXHiz9Z8nrXxjdELJeqPxZrwGcfuoEERa1nV5PVM9jC15
oqqAkmsHlWHi+q2UGjUuGXKQ2eQDISh6uTQKFN0wIqkngttFVXFI68FZqyWY68Lu
bkQZ5/3lPZZ1XNxu/vFtXItB5Qz5JOL8jIobY4STlILwOCIoFLizwh+ey07EISlV
7Yl0W574OcbAucQpR4HDr779k7szew9K9SlMfX+56K315+gubansKtcrsJEDz0ZS
m3xpMWdASyuulMFUFEY1sfUPOjDYqHMnCFhRQWCfOZTzw5uk/wjQlqjWl/Zv1zTX
MudmxXB9qtJdvtXB51WH+b55wJGsWbj/c4MykQotGVmaGoQ3Gv+N+MlatGJYZgFM
kxYETs4/PxsRgugvaHA3iWqiKycLfO6hXtorReGrQ2lh7Vz3dGufN4glkbk2Wyd9
9xtasQLL/09A7LWSgtP0BM1wdnGLT57n/Bc/bZFkWOmFvYKBSLEe6M+SrT5ZV5+6
OoM5aH28JNG7zLJevcbPHdsZ9it0X37fbhGlYlBDITsLASp/VthbhjWk7r/DQqNs
a2dyP5v0PrvZx2Hrh5OhJZThfUnTckVAZWr0HAMCSn89fBs5Dab7Olv0FNUUdnvF
xBrzegP6qPZh78bzSnQKI9NLjqVMm81UGqHgeO/LO/5qn7eDtsFLHzJKTpqIM7IY
S3uJRstJ9tZrEaLX3jyrASVLAY5/jJhuWfHXFkYUmvXlXJXKbzJss0mV69YXBG0N
ii43k9mACy0NsApAPc+0PrLkQLK4czTltN1bpb8DYpryV0iP2hvfc5SjycW+XNRG
Nc3KbQ3gWw0Ui2eR1yaXVGafXfbN3eHdo2wHM6pWE9qZkLaejH609LmML6Gxv+E0
na96nvAYd2Q8G2Es00XEYkyxZiARukCPX3KE3Qio4LjNmKHTAu8wHwUmE80pDmSy
BaIJIf/bGWRNWEElF9chRHOkbLcOg3mgRTEqMUgGA6CpHnbbyu53zzz1KC4WD8/o
8zokRLoPDruNM2MDFJOPz01VMeNjiYHljJFW+sGUBaymAtOcrMf+pSBEkmiiOtDq
xRG/WNN+CIHAgIbzMzx06UNaewJj+AUVkdMpIVm9iNmlg6xZ3yKwfwWLZr3yPyyV
yZ0tqDrQtgABBIhDIBKaZadsNVz1ysJWVKBthAfjYPkr6Clg0vYPEe48WfrE1n0a
AHQxvxKisSVIkaNAS/ghWB35a/C9Mw6Q0egysHKyiPaUN4zk4jHJ/+T/rmClA348
YABiJ41yYM7rLfHdnrZYLUbQEaRPcVgBjYj9xoJAXfl+wtzjbTNWv7nYMfNThATk
Nz8tAYDTtzX8s7cJDEr1SI89FPrk8tFzbnHF61K3KxmO9YEXXAEuJEwzhjs5E69s
gdAy2+Qyb6aQjESWfNGrgGjY4hwH3m3BK0xfBZTO4+bwttMQ0izEO8JH+O7TqVsd
KeSdE+HMuoKIJgJpIMePxvFpb1FBTlfZZ0viiJi69xFtC8lwI1vrRfeLHNz9JDs8
J0IAnE4CXZvsfHjOQoW6aGdaHDjFT7LoKPBx4mj1T6o2nzEwlrpCOys6AOqFopqK
KNdgo6UYGW8/MHAzrkFSZAoOkMO8TZMzbggl4vEKYQIuaNH8NSusKE+Z6h1fHlRi
1sqivNivhu6jANeJBKJBZaThJ0/mAmTLmRkMkOI2D/Wt3mLRJR0VZvpfdKdfQDKU
SE8DZAAQleWyk1pf9NHyFHNlIDeiHbqyj15c2dxmdRHo6rmoFvMcNTWq2dl1PnhX
PJqN/YYlrg5e5o1Os/1CWEs6LMHcJFtlh0DqEw003cl+5Dl3pXddlDaGHtaKe/ut
V9914pqEXIVJLB/+N2A+mPS+fGbdYfjT7ueZzzorhcsWV7s2fDgrmH/RaiFCVsww
dScyqydtFp+dkJcpYFY/i4yxqIgzRN4pCICqydHDG332EgToJFC8y6PRoYJz4pMk
7gt8B0OLuar1ZkudlqSQ4GnmrbB4Xebvf+t0B2hNNQGV23tSuiU3k+UiuJ4x+m/l
7y9rrkSkrmKg46JmtnrbQoQiOFliqbeZKZA+7FxtlpUrNArWFdRtT+I32BAKCDaD
k7luBv70N4Lwr0RseBWAfbdFZR5M03VI1tABFEVrOdK73sev/nD6ea+cFXJ6LfbV
sw9CLrkMdAL/Q0ZElEDHvZu5T/medwjwGOZlJUEetLZ6eeIdFyho+pZWbXpapH1t
cpUULdcmamk+SQvvj17ql96fb6nmFXPN+FqMvLpO3E05JYLtaN0aGBERZKIxCCZa
yMCVfqLExBWWpdEqwXDpNSPozhtdmgiuZMSOjk430KJsO3/xk+svft1yZUNHg/AS
B+iui6vb8HQL4GS9LvoZHCfZsTEbrEIr1f2kV6vpXMZxOU6S5sf/s0FSrdvGfjT5
Gnpov4lQbs7A4tS9Kxyxrorie2Dd6c0bT2kcwGYM7HYcj13IFnRIgQq7dgFbkw8q
x3oP4lQpeA5RTEIYQQJgIAItwo0MzyJ1TaotKttHrcIst6JS1WsFwGU8WrrPcL6J
ZVnmgJBK2oFc1ZVDDT7ETQYOehtjEKGn3FO7hQ5ho4G24tJ32VgXyhwuHlBp2iOz
JlpopTJaEX8X4iGz1aO9YV/FVmKdZpCycVYluXrQhSgyOQZ7aORcL4LGQdXyfxUp
8aUBHZetECAa2I+Np8f1NqGxeGRhu3Zha7+YA6JbVcPq5nDVF+ltPlFaivzHum1Q
cN4iXJbJyIAB0pGeNdU7hbVPTrKISQkVynC3hmOh1qG9hzmN1GMW/qwOpBqMHHSs
Vza1KtN4lP2isL/+Q70AIZGIAHip0w0WZdTIFg16a2B88ib0j3EsozxFxK/sZQ5Z
IIf0FgFemwKIVJzd7cHgV3Fj0Y6YPPS1HeRBZTOw8Ipla+CDHzQxoX3vho9FJ4FF
1WKdlMPhttFGG3Evn7nuX+/50uLWNl32+araUdqS04MiACcdsc6NDjZaPE65QXgp
BSJv04dx5+RhwDRqiq9hKgTB3cvcm9wXNWWzKgxDNkP/IdDYXeTf+gYzSGEShd+z
jeWXv4hsoHOVLOycnjhCatrhHXJGmJDmXpOhB1eITtWtWirJkqWkhXCaglrMwn3C
WEtKvFyyGypXoN34c70abNAK5ixDha9L8O3tp1JurxPJOCBG7t6lC+SGK1FEb3Hq
yCqIkP14aR5yEEoLm6cF7yoETdSVfHxKjHbkaR2ss5q2OfyFBkDCxGqXUjTuBKE/
QLA2+q5CJhX4p+Umsw4X5jM99yzTQKBx+qjqq2DVghTXQQvQBsMstZ8alclNxkyx
6XNEhwmDu546qP8MD+C81dGgl/As/7lhgLjFOKCDKAFmjpb+pJVAZ6e2daFA691y
sRL57z5NXwSJ75LRhuSiQkZxs6PLssE5A57jpPhQVC3TfTVNUmuKucWTaP/wEJIi
3ZUkm3nJneZxhXfcR0rB6pvxTZAFewt/pSwn7quzJZk9LOtFDopwTIqWY2ZJIBKz
+ICK9cDzEX62jVf94asoSzY+lgcnozwCHR0n3e2kXR5OgcxIpJYMrorQMuJ65KCO
8QyM/ixAMJ6SQFygogL4QxJcj62feb/QBEOhpoTrQIaBS06KSCTYXHBL8bul55HY
BcGGvtyQzHYcdEiaJ+WWQ+iNQjZyFt8qx5Pxg6w02rip9uMWoM8IoNZKflwjBlfm
oLuJAnsu1F3VVMXs+07Vmtsn2X/3basG1qry1DdtnRKWXlOb0yG6zbXxmPFF7Zpz
fg/yy4X5TSqOSGnQkfwagDmsqBmY+lQggkrARWAL6OksfyJF7QKfZfMI3y3Lm28e
zXWUYlMacZI78n7+1M7LZOZBNmjTcyCFsy/lP9uGkjN7AwNLP/MTQVmzv9/OvXr/
TiqTZZFfvcslmyzgKKxDxTNf6kgV65pwrl4v7aubQH37j0lWUBOmhOyonY8tn+JV
sfsCJfc6Jlotyao56c1Tb/BPYVIYeBJA6MZ6hg3XI8Ar5Y0HRdB0RSpXDBr4W3pH
jYheXl8kydWTG7cCbzQNkNnc+QnXyDN0WUTZCTRitk8dBZnaNrdyhxLsdhauCkmt
+gMjGaDpulu1xr/TLezl66ZUU20cpEROLBVSV4/lTmdmCCCRhVAVGOwxuqz1z5D4
W8dZv8gYf5FW0sYLyYMlP6k6dotVkFo1eneV+5CZXLV8Ii+VTIMww4JO7OW8hnlW
rSj5pvXetVV8MifHkYNWb6vfPmpOsCcIqo0SNKD/iqLu/8n9LHhjeL/UM/WRprnL
G+P+V/N8byeB0OuCCqJqH5z8NP7eq0G5jmOg3RUB/YbFBFrGlG41kNrv5Zevdy42
YUnhHh8i+P+ktvsuI4jO+4E2Ibr+Vkz4eN+9H+uOTQqhR8HNUO1IOQ2319bE00Ug
+/nigNPD3AUmq59zHdwxmVM1w8WfnMNmnNgU6ySxZexF0nYG60Jq31gg7Sz+fpyW
bYZ1pEksG+JZzA3SlHjQUFDeLSy11fYxc7BXhaPgfebi7oSvXn9lGRwF3pA0BU1v
jOSIWBdUoXY4jI3yRw+H2clI1GfCYbrbuMr12dT6CFQeWFbKCgcyG1nQcKcdCT8F
uXf7K1ZQ774LEKtO5OQyJuOWcm00xMrLkEKkcWQaXQtH77z7zlKgAgwkGoSkVbCP
lSq28dMbKWeFuuGjWD4RE+Kw/1ZDqXMi8sKiP/J4rMjLKOZCWbXunvxDnJykji0r
QDjYoxPMKN2SCW2qVynwRI0wn6D0kXt2fgWIIcvmvZL9tWlE9heopOP0Rh+6vCBb
F79yJmPK+/XQfjW3Z0ac2eMfipYyocZDbzaPCjXayPuiqMSveORE9nlmjZy6ZzX7
5iVxfekmt6BDrVCjert81judE0P++BdbGnMwfP3JwN+73URg104D1u3mi9JFpYLl
yzVdo6j1D8pn4WVC1+x1GeyJ1MwuTNgC6Z2dtKJrHKJxcmGtkzE7X8N8+OS097w8
JAzUFv7FFCugpQrKPefBTvBfFbenVejPBBsfCtyilV9/u8wnRZsUeA46A1ghLapy
+pp/zC4SGuawurG1R/uv18qx+/q2KX+nNkQoTTsGTPz4PRkNlm4U6jp3QZzFS7Y4
81/SPiUsK56uarkL+t2eRIS3yKh7Vly28JmtyN0QvTr21URu6mlzNOYT2pg2TwYa
Ew4K5y6yRExa3A3BjhOcetkzHKJgg6aBh53WNcrqiE1mpQ4Ys94rtZa1I7mHfJTp
HFkYIfsrbOAjxWRU6DEcDbpg3KoTnjOTY1TDWtQNJf1giBJRw/8VcyeKppo57gMU
cDUmxqsQf25AOYUpTVVvNIzRV5p9pmpswM6rznpodXOCdPZPDpv3rI66wOipkSUH
9v6pZRInWRVTyrVPXIYZNmeBHxtoiIIXyOBikcffkoOxd/RmHwQTzeYli4kOKVOh
2HIb5/uHIFt8Wk1x915JLQ==
`protect END_PROTECTED
