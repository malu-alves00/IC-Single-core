`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NuPciji5VB4W4YMD2PKZUm3NAludk4jiEo+CgJdGhaq8vnzmzmbYHGbjyhnluEEp
g5i1Iznw1ORa9a39PPCxszlXT1u5Sxrlqd+Q3JnJN1dmrrmPeEjPjf6kaxhsHbyu
AqapvJKlL3m4RlIvSe3BDqg6ptMWEdUHJmjoeb+dqOPvfTHmZwncuins5phuKjnv
8JM9UPqQzPu3i8VdBGTYhVo1blTeD7DSm22KyD89j7TRf5zgzxddEeZYaLIZTgyn
w6NrEar7CDeb/Fs/5DKm9yZrhoIgpAKX7YV2V3r/HBUvUlZsbZA1T8SWviB/KlJX
5E3RQpUHl7AMr+TeJHDhu5B32pvmkjrEuOhIOinaNX5be9F5ALarNumxDanf093F
w38+Doms41bWDUmatuzbJFd9/WKme1h5rO/cwZ/M5PC6C13mlwX+oRCHr4H7Rtu3
IfUqLSMSbprx68NCKtZ4DooHPo2kls/K3bqe2Bqj975xWwBaooDS9s43j5LYTW8+
mKlDKNCRbMoFLip+/fU9KOCbtmUXjXo15zaYwEetLrPJpX/NbO2SBTMzVqjpvtJT
hNU2eYT8BWv2onuZp1D+BjpUQsnOms0f9Lzr3ScJVaftHkiIFw3QGgd42I2E0wBj
FSDzWGuraMND1/Bkm/lgD3ONHyes1/EBtiN/MVu8k1ga+3hgmUPt9mnDPnXC9Ypn
++CyYw48M++9w/3U2ayx0W3WS3uYEIiHph4Vhkgv1fXkgblJttcEGNQdCn1XSsBI
V6x1TyffYr4NCoOmV80uDx7U6ze6Y3EPx/o1wdBrj0K/RYQNzmzh6WrXf1DNrRD3
Cd80GOa9uPRATxZCuM04iUKDuhgKAxoa+gdCeht3Wln6kZxAevAaUnTYwPYITo5x
3ykkO852u4jL/3O9jQmo4xVFvrvia34hf/ijuQtufCs4sRux+5Nxrb1YikDJd08/
+2tS0mcw+zizYrv+GDAJSRdi5Sax2RyR5i1lZp/Iv/6qJcCzSl9SIMi0SvO0vcFu
hmgHpKaP2gsk6nq+3poawTrxTYo0X+lsrZA8l1u/FrRZpnhbb4SNImjadbmgyn4C
ivxDEy+4uPiYECm7ywRw3sCR2zC0EhGwbGbJ/zg0jOApETAipkfGjDaYFOfFSMrB
3KQC2P4T0UusLFdE3v9YakJmaKpqeIjWPNwrsGhd2/Mjtu57yPbUDsjtk7/ArAbP
40XrVeBi459blfAJKrS8MNeEfIGx2XfYkU5AGkYttQxJkuqiwOr9xk4JxKIAmaC0
cm8esDkjAvHMCfcPgL8QIi9/QLeHBMRZcg4dJ1t745Kbrh7gjZP753Rbqf9yhW1f
tKp9GgcNuv0Ohu0SH5XqQuUjzSnlltW9IQV8RcXjF1A49/w1P3dewa+Y7NuMZ+NB
expv6crr73ySn9iBhielgo6CNTQUjo0oCJtFoWlyaILAoxN2iOfh8KglQ1oXTXLI
eb2qh88fcGdKkg0HKSLt6wVTipLqGfMkKbGlwAxW8Ze++siggge4SD6Z2cvKSWNz
dmoNUVsDegc0G6HKJ2T23hw955g/EaC50EvNzOafWQQ7fGNER1bqjlQM+9shwu8C
NkNGdpseDIZzc1zgqPvxpfdAYeDWwIewV3BIBGZ1Kl6NHYk0idoY196ZMNLl0lRT
jShlOhVJcdK+Ex+0YikUqlJehQQsqB44QTPCfB5cos54Sh26zQd2vXVg7IHF9AwT
ORhbf7pB3duu6uhYotsB90AHAVUXiR8OQ40H4dYHazWJimgHwNnXrnyBmVRlpR1G
TutxEMu5m1YsvSX+76PUG1i/O4ZRhXz1pyW10GlLhEEbmP2sq2Ix3YEpC+mQ1vCS
ZKDzcHUrhenRc6K83TPRW1xm98e0S/cXmbmqe0T+IL151h8obNVHzTioYl1aWfhK
qvw81BCvmXlbed1m5HlaAxcsFW89RKWS5NGvVlK5wIFFDUAh/p9bwzfHCK/eTs2d
DCeBl2Aw1/5qH3IHctA2C91+xnJW+PXSLnUlqM6GS0Hi8vVh/sbPgSbBUjo9FYot
OYwYPKWuY/uiIEG53paProcsefOGXOm9xI3Oez/6PjEQOZRMQbRVAFg9UipaRXDr
IpUxaeGgNDM6VBTFW+yN8GOBOGQKzAb2/0Xua9dmmOrfZqQY3wcX2WzAqfLn1y+k
2dkYExvM7NJmUBqw1OPRfvhCjoxEImQDBM/NTP4aWnRxEl/rstFVbq83XCaZzRBT
TBiWhenxPCjLRajcfKhHsr5eRCXx1u2+VCf9oyLGU4G2WyGXlItfd6TAQpIyTz4U
ev+WcLb6Sa2cPH4t6FnUFwGHZi4lu30D7vB3AdbeW7CNU64El8bpTHBKvOlXvmDT
U373lbVlHO+0ChlNqiK/UXSU3PJzmRNEF52cRxWJqNLpFVYQfZragczbwvDcv4Mh
lqdniCS4TxpfnChSahTXP2UBo16O4rpox4aBs6qwpT7W7lHIpleonBISr2fOV+Bv
+dOrqNTtBdhAD6raoHBz/4AiYBuZS/74Z2s+F7V6ZZZF/7UVYerrHQkdshaBwmCi
FaJnM9x1QmfeVyZPaM8qPvLfX7WYarz8jrPdy6ic43A7Po63j2L7F3bBgECdby7V
TxJcHuO2k9q51G43KhcqRrGhnjYsEQKiQ/oOET7VEnyC54BTCQWPdJFdqMRrHpjU
n1WNYdU3J+Pvb+PbMEdUZ0a0t5WshPcEng9SkPLdrII7jC2irvNsgK2cNSDIEZWV
cDIwDvjNW6AP6tgBDgNsSw5+1YtX/vuJndjJCXCnN5IcMxca2uKaa1mCvgFwd5PP
95tKrgGSWdiJ6pm62hbo099ilVV7TCBOUlMEGMxmF8WLCS75SmUHC2C2Qv1LmkLi
tQdUh7grOytRuvWAT6l5mcLuXurkvxfuDB8DdDbbisTSNlF3VzFDIMq1/KH6CUoz
Q1ywTI27ZDtTY+Si9E1Q2b4yvI4GtXNJeAwHAbKCitx9B2qJdGxBuCt2+Uqmh4mD
JZihFbpuuw5HDT7kMKC50r25YUmzc8+ERzRYxmJEch9Apo70M02LsvuzNgUn23kX
qLkwtA3UGJWTIy+x+kQFB1NZpzuguobIcUX2Z5ThpQKYAfxmmss2FO99/QU8tXcl
zxyyiiOudWWTCiJ60j3rMOL9oV459eUGjqOTUCuczgoaxDLLV873NylnOOiFfir4
/swVzA43JnaHFZy7b3NzqClC9UQoD0hiQOKwPdsQNgH5te8MwuZJEsCcjlzmd6S5
VBEReHRJCA3B1Oc2jgpHu6MqcvXc7afaRkWmPqnUYlZRpCcIKi2QRbNLXoXECSkN
Wb+rs77YclL08Ylh1Rn3mYBgIiGMrENSKa91WRtkG3FQw2Wm0cS17PaXZkb6HpNe
UNQ2tWsU/A+sJaI3lvMIXLmin9OtPYC5UR6Glo8tLkGvNAyR84KRbLcTVdZKMK61
C+dcZhOfZDU1/r7WV2BiKrwtuKbwg4f90GV7jICFiEYDnqXorpmKISwE7/ckuaMc
`protect END_PROTECTED
