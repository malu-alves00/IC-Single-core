`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Gx+94qLsdRDp77RVgcWzxuOf2Mk/l3dL/TFw4deeyPjcM8X6THnHkEpwXTpz9zji
kC8Z4CR07mRm0IpD1I4LE6x1+yaUgqXcBN6QjD24PLKxHcrDnE7qdIQwzy4pB+DW
sEzoctVMuRehMrw14lXqd3t/58fhFIbG403GcfEcL12ZXvAOnDWdQ1N8S2PA3bSl
damq/YgupWOGO57OjYzRMCzTS+3rCN9KDDMZP0FeDhd67TI9lJLrJ7NGxA/qx3L9
nUa0sjytPfYtrwSORfpC7iodDPep//PHwtLB2gNVznPNyh5SEzDy+c4XiVZsuiY2
k5Aihgq7oxic8uM6t0uXhbL6hxtiTuD6VN/HMH5isvn6KIC73Y65ExOo1vBDNegF
8xrcYL8E9vGYsVOiR5p/SEDHdzJQzxvVHCteNmsWvlE0tHtyrxo0bexnO5kBf2RE
uEMYp/26fjdd/nQ9qnBHmF27MJ9ymw0Ch1de9aOPvmUWfsU6rbP+dMT/mdapxgDm
z8RQECdGjzAtyMgJmQFORQHQ6F/LfiarpzMv3ILW+pA4i9z34XzU0m7P7jA9jC6f
RQSmIiOubxeiklnJQqLo2ddQENV9IS2ObOLkgd7EXxi/+L6ZUfvLZbRmU5J8WSQb
3CO2KF5cJlXwy8sLq/9USk2s9ZwxjjTfQl1w7SDozqz0oDky7xfNlV6kjms8nVDF
pTccvYqgLi2GCFqdVhFq8hfWw4HWkIAj2rqBJnLDw3z7VPU+Vfq1UEKiqhRufawn
ojTk2FY3B5DmG7PfRZ2Qh7k7p0EjuBgqDG18qlaHgfv1IVPtQeVBxQ2lEVWnOftV
buLUBtgIoQWbr1u+pJko/0xjuiwSJRKJt1nhph1hvcHcW4n+POO8Ldv849RXxO1Y
5hIG/lsjuPR1+9APC2O5WnuXutOdJE7/8VIvMU6wrY8rs2YLJ3s+EjtzqethYejl
onH375521EU0cTaX7G7TmZ2UvNmEex2GxDN88y3asR8JWzEYo3Z96fZkJwjIA855
E7n7wm5eAhd8sbRx75EHtjZen4bSR9BhRTIm9XfB7mbzhnkBEOWqhm2BMm+x6NhN
tfgfmcjEJLPKoa2MXvAQD9kaB7+vJQnSy1iSfooOnxSbogdi/ZVSv5C4oef0KzTn
3svZOR0PP6trWgWY+m1atjHVBgaeXY83U7XCb+OqogTJbbCgLE1lcWhpkuvP6o+d
ah+HxO88Sy7i+2V/SSP96K1a+oXX+JWh6x8pWyqOjhQrMdALuo5vpRSIZ5J4BiVF
/l5N1cBkGcZ1kn+SMzyCFcaXo8Dq4u9xY452ruLlLleqryqWarTmd3mhO0uQGF/5
djYwPo4H+wlPMlMoCvi5t9PE4FWoSWcu3GEuzUrMb30K/yALh93IEyWbOf1BnCxP
JxEk+O8JcuKFdcUJluUXWvpgz/+iJFETI4koIwcr29ub0iovhHcVe0GJpHK60ZPQ
gcDFLUd3i8pqBD+NwupXzmJrbTYLQN0BDdlEWjzqigtPRLVctff7MkG7tZ9XpU89
2D+KPR0Ov3l6yafIf8MOm9OOmri/TkMoX3my3qzge2JYnUjke2qV89l74LsAZ+pf
A/6Grzd/FIAgHSgm8i55LNmHBEnNrxDg34PDYmJC3ZreG82FqbaLCTcFALjGwSx5
ld8OCIZdPriE+EG0Hhbj/xavMu3ewfsJZpx4VtRLkgTfQt3asTFwA3OKmtVuWS46
NpbhwuyLyB5hWMQjVBWOiR5vuD/vWhWG2I5dT7E4k70e+c7rpgNZW3t4bS7sYJY1
cTsz9Db3NdK+BF5bOc4bLkjdcJuhyCAwJHKOv+YvReyQ4zvpWuKTCLhXZ9sG/j9j
2My0rlsBSBEoQWo9qiRAf8tK2Xf6pzmu2ZP0d89SXWcdJCiIIp9rV2JGgR921Hhv
NhfWXT9YTXP11s4GpEgUZOBYbWM3lSHySFwYKffzGvXlZoJf4H+tbmXyi90GExb5
qzrt7xOY7+riVxsz/mI8/ZShUuS2b29oTeAY+YUKdfS8tVgjvT/vRoF6vyrQR9fI
3ZRbcmgvB1G6Ng44yW3FAdjK9xUW3IQzFDvIvPDZio9b4HJPIBdWAxvkV0a84HtU
MKVG23DfqJmTQjiit0PYXLjM0jFIneDX15spobOr3sYQb99M+5UhM9tgjpNZ9awZ
qBPVzzG9ST+zJ3DJ2VPIOBgQ2EUh6p/kQ9kHgaFH+FRoQ/Fgse3DbnGJngEGWLQ1
V82bJABwdcm4vmOvEA0AYGxI9lr5Z8einx79gEeoPbzmXtvE8OaFbhH1HOy0THa7
e8RIsXXGd9WaSq+dvcjo3LdI9M2OWThkGuy5eYUm0x0Tmtx9kO+tgZLbo8kcoMSz
oO616rQgQZlMpPURZAed5Rg6WkyJpChPB0JIau7FEkEJr2yZULcri2rp/xKgDJQx
ufNXA2rf4sh7wfPZ97DfYS5fk4E1qwjJtPbl39TzpkUMYy+BOxkERtYbpHAk38Vq
toz02I+83mnA2XuytSwXlaR3Gkc3Sb6zSbhv/fe+MUoGz6YR6k7IcxcBH+GmLBCV
/x6Tiz0P6mqSDsXcldI9MVmoVWmT8uAonYbC/b2DidsMeRQ7iKeJxIrYkjsWtfHO
0HYqzi74mh0k1bokiSWZNZyb8VV0H7yKMLcecqD+Ul8IW3OvSeAqm2Kz4nos9E4Z
9yITBrSRJ3LGuvk6dLK4+yyEuCzLFoJHdQki/pc1QUa59pVLL0IVpycIRCaFoOKr
Q1kyXG0lRuvVfABRZ26kgEJM3kIyPI9VGP+7NKi+x7tGwfzq8jAj8oPp98JhfsYn
HpKCbX0MWGAHMJyn3e07URxNFxW6N6dZgctdxMp0L8i6GMlFTgHTM9C9SqlAz5oV
1ja+ke4jaywFxtRv/G36fkpwN7Nf1lydQPqDT+h5cB4rfhZ4JeS9BAC/0dxGyaum
P+OX4QV+LmbjZ7iK1rHZ3yv35a9MEar97zJzJ4dz/BIHQdGKlqwVMpybIKLQCZVb
JbmaCdCtH/PaAGI+FdfYGUzr9RFjvs1BfHrDF8Q1VWPSyPbXb11Fvui084PKCP2r
AVgjUsKExeIDgp850iWN5kO0fe1mhPIU1p8sBYbtJdeN3S1DTKIBIWULaQDes0+C
r6x7rRhKX96m3VFS0Aje40THnpee1D/OyRHCrCbBYR6THfDCCmhMdwRDQomfFhY8
oo7khs2+b4Mw9IpbSVNkG5eOk0Fhazad0VgpHWg0RCCYgdeSqC2ahQRansAXWuox
9jrz0uwz8iVHFkA9glvHe3aT4OQgGJuRjQlCGf/5BCgoWo8GlWlJ1OvwdPnUwveh
sGQDeDZn7b6sgQgc4LeodQLuV9Lt6y1XXM/SlCn0QDe6yP8UfnbX+5m1m61K7C3k
38kmi8wyweOyDBr9kvRN1fygusfsXDXnx88rQXQi3wVRKMQe/LMxte6UpyRxyKQR
yDr4QKnqCxV9XXy1E2ssz6Nm1/VRc5Y+kRvhnkKlnup+KBFkf3SHGJE+DyL/bj5C
SxdAit8cfr1Luvsp29E0LnhWwj1Ikv+nRxQdC49gdZQTgNmoR5Rt4LR0mdzzhb8G
GQ8N1kUXPgrph4SMamA4MHp4q11fb+WOsC7KeQtOINto+NqBvxJsAhuLXveCwuL+
tdfHK2Sgq3rFaZYvbra3I9R5bjMP29e+z448vNkIxtAqjrx/fema492D1Ouy07w6
Yhty+Mj1Ebpv1K51eaRyrU+qgXw2Hx+nCOySzgVGLCHC+u53ooyaKHfTlq72xxN2
PLgqPCqqh24JaE0NH9OdIFPxPEaAnLuFFyt6ND89ngJ4/pEmEn1ncK3VeCle2+xb
FYtQVOUqCS2MW05991a9P6GQhYZ/f8eNf8odu2w1U2W9DedqzlRBK2BymA+v3kJI
PO0+ff7Tjklm5rfi7MPHzieu9tqIsZzgZk790YccL2XphZxINnh1jU2epkexAacK
d60L3bO42IYiRshqO+oUpm3A3zdfdOraG4H4W2wUiJtfEqpvGtBlgBAYW29tKFdx
DPnvsXQ0HSj7mlq32h6+SluH4m5ZHLU7LHOOUOe1RA+hurBLeSg3Ycqfa5bJdtp7
n85izMbrwNYx/1QEhdTP0tA6iQ7xrforfHQw3IjTxA9GpWCP14pNCvjd4vyTid3V
Adm0Nk4sMSTVZB2/kkTnz5GiLAsZggrvTdQ2A7Ph3fU73tNl1BLTqtzk4AwUfRwU
oe+pWRi+DX473xRgkkkXTMisbhnQObBw6WWWu7uXJsmpGCYSmZ2yOw4QtGAQZmGm
SJ750U1Q+nHEyx2BfXM0FnAqtpQ/vH0qG0JxW9HzRiGxhCxQAxs8SEiKjUy1iTHm
KQyHWA/Nt36dfWCXJ0b7uc0AfapIY07bqglQS9GxmElA5WSHRNiI1zWFO2f1CD+u
/pFBygzEYQ9jXShBDNqYIFqd0cCFrOS26AUNUpVPoutk363QZU0B2kiaaje+Bj7b
jQ2lNilhb8jy2fdvpEdkvzMqs/dwmuTHbbCgOP+9i8BffgHBapijb8RoyKdZ2qT4
l7ppR5UZfyl67xz+Z4Pm0igdNijxTEauSL6sqs7Puf/97GE3KooyVGAcqy0NziCf
GUyNcPCFbAIfd+eLYHrvr8sZqqF/4YQhZWcUit5Z3cVCJykeDiHP/3NovIJwCXgo
0BsiZwcr1sH1eu1/YJSuRglCnwmG4Pwxa/BYxYdlpLw+sRV7Vhgn8oV7xM6s8p5b
ri50eAvKRcRVsKB3RHkZFGRmPuUzprbjs7k77JstUkas7/hta3MFzurQPCYVmdIj
PQTP266IwV+C6T1vJBK/SMbDLOVnqGZCkvFw/UoCNOisrmA+DD3Nk/KVlkKxAVi4
SRfClO3R2lJlU1MFAfd7pyiMtnq4lNBd7H+E9heEVXJ/IEAZWqvUaYQ6ubEUCuZd
ogEDdcIs5gcIQMj1KRqWcs+29CHeG6Q7/MWuhsliQDwrm7sV9mx6zKLuoYGPD+oh
DL85nDqsjf5ps+qRYIuFmI0AU97fvlX8kIC5Hc5w+7oIKsbTwBp23jF+a4iaK3CW
BjWAdE91HsimATtMaXZK/ISl9/63D3Cx7jZ0bfAUjHHNE/w6oinfjt8RbBfWHApr
Vwd77yxYNLUZYFYzGuspTGjFkrqNw2vdcxuWqvSfnt6LXc/ILGhEiGxaxYEGMtJ1
tBbNONtoxPM/fxJLnthi3gY5dxD8WrNEkMGnuXikufrhLqx83VcPnkNbyaFxn4m2
GYMia59D+eQ69gpM3yIMgV8y3KRfKB9sndZGTHbD3fJaWvOKX1EioUYBa0VwYcPd
74u8hz8SCD5Q0r+FNBYu/CaI74X46GyQUTsVWUQZyhrOcRS9suTkBkhaP5aF4tfG
2dG6HmX49FJ4yhu8lqd3+o9Sf/DWRSG0b5YEbDT/ClZSADXlkwBi0lRIUOTFxr/+
sb04JrBIM8X6ZtcYAUHAvEILnoyU5N6XlM50c210/+sGHB2A2naTEzIRsxAQGQ/I
8bbYsCIyhREs4bXsDmTVXZtaXNBQJvqEoZ5YcM33s8/2bfo6+meMGVFcgJjVBhQn
S9jypRsU6pVhv9ePH1DRRV/aScPscTAH7WOapusaM1GGKoLOY6gN73EFOPb2mVye
jEi4mozi+MoaivF4K+TyQeFrF6ubQRO6ajFY3rgWz915OZdVDxR3zYfKvKJetdwN
lt/pSwFhVBbhnxmGNGE3cZUqu7JDK3ANXOnQVVyaqJNGGr4KZU+k6juep++SnVMn
mj8BSE1ywhwQdBt2yYRc8VJfzwKqyHQHgCE5wBQuDbbhlVWTqZ/H0tb1wAiAKmdy
PnmuoBdTJkxrkpmTkdHN5HKje4w5vEJGYsbJVLGw3ONUc2z25ZIvmzx75LymDT4d
LtYuetVjX4Dw4n14Osre70KwhtHqwCRh/VoN2yZq7Kb00QFadhopLSzx3Jhzdx1P
OcPDsTCmWZw4Ss1PBT4mWCHPkCrRLDKiYX66KEir6C0RcAs3J4xNqLrJgbq1l+75
L33pKtTS7s5PqaT5zc7NMPe9QQy7Z+lk+Fq8eDaSyY/nSYq/0/02c2jRgvm/BTGI
r2pwDTRhv9ffY5n55zbeOCaREb8A4SduhbxVLhvldZWmM2RXmACXu/JyxFAimXkp
7t2ieAYPWIFdm5SIoJme1ftKFoP5ZDwg1JUKFg9LZBjS+izVD53NjptLhg1neefB
n3LgB+S5ZJ14tcOUMEtgBSXZJD3WKp1/WR7B32ibaeImFbm6lay6IntJXW2djFUW
GGX5yNDU0NUQKH7REO6YzWCawZGIzhDI+/LB0oHhI6yMo7EyjlrTJiH8SXuComVx
wVHbIW9w1ELqS3ZcqZgYB+i1/ans9Jpbcnv71z9UBd9h08ksKbS2NtbtywHxwmhm
31estJmlztGIbYpJEFYK79Dr5806xoibRUUZf5f2XMBNN89Dz79wdCb0TPSfst/w
ugZs3YWanSulx4z9zn+okA==
`protect END_PROTECTED
