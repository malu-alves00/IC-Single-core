`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
L0nqW2ykOgZUHvs71t6dBaxQ5RZToa/sRi9pIbS1vfQReImHwnAT00TVR3EE2Y73
VAXmCyzc9ini/YZ2bg4oiNdUkD+I8YWPiyyIgBmLpHiMhZKa3XF0+NRu5En4yFm8
bw72QQrWPtjkgsPgOcZ2tfd+P/Urj6gNRJLZW6vDLwF9KZ0i78G58Z+6h5mjkly4
hHpVUl6MS7oO8EcfjJGBVZJc9HtKrFBBjTWrW8J+sfuX2ZEstm0r6Na0O1EePU42
TE8296jWCd7rOOFq0Cwk4EimBCE4It/4X0CIv4pYMyYV2clJ1Hy074QP+m9MJNFn
nubdZ1tEcBKjwsg7zuQt/m1Y8igX5jyY2Vf/gnrQ7CGnsMRzyFcLQkeatP9ljakf
cCLEYaQqv3Hhpl7LrAp/b1xhONuRKpxIHuh5tCJZtSrHzXBIaMmVFnMwNkS7FT5h
U/y+NCvEQVuTqqnFgJKGf9kxm9meSXTSBIvewr6SHvapAq6ZsLVPhsJLpjBhjBNM
4bUCwdx4MtLIJ9TlraURLiKpr4Cwou+VJny7y28b8ZU+LWHEhQVmkGft5kXBUE31
xIhnhunYEBHgEE+ed6eDqRId4DN17hORBGgxe0LcqxdiYVeWzMJVy4i2OxYKc+sp
ZKVmF39angzXRARnllllHCejn5pq36x4K3mb1GuSFvtoP3Qy2bY9o7Vlb5RnAXc5
okxCm56O9DEPEQfuwGdzv0FquMcvb+0YSc1yPA5RMue87r3fgpNetC69dx9QzfJm
IdP9S52iNOCuz/b2S+p7Dh35SoeWHeZ/1/z+4SRNDeg8GbBXrKGln1DihACmgepR
jeux8J6xA9l/2GNfWLBM9OBPxG0M22Vn86KAlN+iR7I=
`protect END_PROTECTED
