`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
D0qwi6ATxbkirH88QLwVuxu8uFZ73bpvGzBqci26qOLQyKKVsGTaf+pd3AaIghnH
FJujkQpyBl2iy4mYg6vqJzJcOZUm55wGqUjLdCpEr33lUnYrIfhlIdUXdi7Ju5yf
1fGO7Jsazy3tpthvNXctBqizt8kh7aVpZFVyXozvKssoh4YRJFvMZo9xMQRX/NHU
Wjv+Gta51GEkWmgKHIFuLG7+qi/rZvnbdIETbqkiXBW/9zS19uh2QtWROflp6PcY
JP41fwRjFGg7zuQPydYDo0SR8V5LV2K2x1mr9ng2piy6o68/5JLFD4ie2/iub359
FM1M9SEwvmzphIkq72lYtufPgLEfMbhEFxOqjJIFo7uyHFHctVSBvtipi7bYYIua
j957OIshP/eF3NKGU8vNOnSmlGx70YAlUCzcRPR4szzvfyPLpWu3aqZqyJBfeQz9
VqUPyxRxhcghSMyAW5B0hBAMf7DrdtJfY8Uc9sl7yQXZQdZLatDiQ2p/CjJKUHQ6
ScmoIhj9E3SQ2KMrXjIndhGtMtzULtrZ3PpoVBJaR0O0s8rj7j5GWH8LX3dkrE0a
y/XlkI6i+7hUNbbEncMnn3wqIp+bytj/6y66aHF67t9VFoRwMeOwcP6jwpsDrhmZ
iNowFTeUOnve9ZHL+hDWA+5Tc9rfB945F0TWBsq5eid/Iv5qKl83MoyofFSkHvhs
JoR/Aq1k/B3uJTwr0MzVpGChhNSQmJ8Y7HLXR/je22ZfsatWWZLIp8bgW7M7GiU8
Qdsx8htG21d2UxFrp6LsqngSnOYBsy/fYgWSK0I3fNjUEmgoEeaErChLdtj+Ogrn
3ca3ZzQrZaI9rf+x4yVVufg7TuPQIzZxH8NBjC42+sq5csMIS4lPyVykh9rD5uJa
SVCALItgxG3pZiiyrbzB460eiQaDiEWbgHhBv+uVaBhHQ69Df4AWGeEaLajaHKc7
1Nh5VjuN7ev/NswCj1l0U8KsJ//i8ES7WNKgeQ77qh9NnsgH5X/khl3633C8RFei
sR1JbS8GEqobkLMWHDV+1owIJgc0V6/j3WIdysGC5C5DgMUi9NkuPdYUawUbgZhX
badsa+d+wA9YJQa4BXmJXJ/D1tcJAZcmenvMXQKkC1tzqOSNisU+aNotYtXD3kg/
I68TSP1pbrMOZKYA5PM8b5U0Snjgnno6kOshjGrTCQleX3DWk/rIlbmLhFR5AlIo
+oHo229sejFjmij5vouiVtUfDOvBp1XIRbNvRBgjwJGhf/rbGfnhc5qYJRaRPGRn
rtxBpwiSs+ujoI381yZDRr6Qdf6hRl9mIRD54nCcWFRMLZpd0TGzfxPR7IXW5TDE
N17OIbk4jpR03Tv8+3GlGeGlECFcNQTO+U7mPGkyib23PunNyeBAqnb7uxyWC7B9
V5U3T0vecRorvgNxq27YLHI4qYR2e0TuXweWx6Z2i5Szt9vmhJ+h+/zk2qYhdSBg
oPyoYQUNTFkmKru3GTXWx6JyLQyB1NHCsdTzGzva7AoCIcK4exVOWwT1a3b8+TgO
sXQ/HYMVADhtC0EOfMvWREIirl6bQFFly3oSwWaZ6Wl3ZqveVLQ+wGMgMrP4bF2W
CQcDoXYPATWLCFX6kI5FJyJFsW7sAVTuAbPORg9FdR+70oA8dRSCwG45LZJkkmqb
zC4gJC+vvJ16jRCLAHW47CfdSTHMXA71bi++4QZ+iyVLZLqwDKT3byVO0rN/Hti9
GFXnWYc8tW1weMAqi46QLM/KIsz8cMjuKNE0djR2H36tPBl105SdUN2PVyabQC2A
g0EwZYktBM69CbraH/2mQkVoCc6WpYW4tn6Rf0aGvPpkLliJFsYyRF+oDhKFGAzC
SiElQh0OCbJ1yYRYH/TDw6Bh9LKXUT4XSqeanXbU/ws9E5/DvIeLnDCXffK/cPz6
WBZef/PGaLzfyDk2PU47cMzVODcKr4JbOSP9ZYoR1WuoTAt6Asyc1uMzMxejVurV
`protect END_PROTECTED
