`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jyRorf0ZieBHvKIEAe2rQ32+UXYAJUjAcXYUEPqU49+AYRukbxkSXupXyXwBaiJT
vdf9spPiB6RjxHkZk03/nlO7XAwUXJG8fn/CKVM4LPd0l0/oZ/1miYtDxEtkVsZB
q0MxESwkneM/KCM/yVdL8HzeST/OHSUtgthG/+uE8ahH9RKfCCfrdbbWlX/1RTFI
d5rtHuLSr1rTR/uWfttbPMXKGI4ksNaMtM9I9zz0plxl/LOZSieOOHsTooHcwyyS
ZlWj9S9F3kSSc86cxkvV3vWnZnTbc/j0wiw98PU4MoP5AaNJKA6rHskemW532fxy
j01LMlEIWTSuR69Ul3W+9DsojH/GwTPqDBiwbL5+5sibU6ZEnTFdHdaAWrwZEXZ9
8JyeVpf908QrDPXe8Wt07aYZkPIZjYIjZBuc+9x+PcR+yNodZk6aUL/czmqyZ7Pd
eymG58PBpWklUFtBbNGJlW7VALeTbzMjXKE0fqKY1H/Q5V5wLPb16xx+bhr5j+UO
QR3OXZh7XLZopaE0TOyOmOn0Q0bcM5w+7AMX4l8ys8y1Nyc/89vP/sFsZ4TZCWxz
M1n0OhIGJDGqvAGHcFByKa+saoxh9JF4RVNLZPN2kAl/tMTP/queDOSydiCTM4OE
x7dbZ0LpCBi5frEnNAaDZF6Dd5ZykH7Cd9IaGcIWYP7FkPC4at4D/SaDRqD4ykh7
/mHvyLH8Pjinkf3dXuOetstGaJaX79F1Jq3/P158hSpMDLyMHUuf8AmJBr2jJzFA
1z6aBfVHPsOTEY/F1gWMA/RD1pO1hvpKDwXsXIOlrcXL302/kZDXsPJn5v7keE67
r12epB54AaPBIfN2qpr0Dzovmj/3VwyoCY7wXe7Gn4Dk5CCNdY/8TfVt+D1r/P+o
bX1ib3HZNLFuIKa1+s5gqI55/agDmR7SZ20xLg06nlUCnu+aoVFRerNlZ55La0OG
RjHIuPsLQqDahrIoaHEgeQb2fF18KDpbxmardu64Qq/Rq+afezRR4eO+g7Le89M6
EVNPyotccxZ6sTeimhKzSGYiRK1sOgzbjEJuAdAoMH17OxMrYBHfFwCQ+YWyFQhq
rr4aTd6wv5HANtFQie1poHxhF0gdbx0rx2sili2qFc43+iB1Ffxm77Qu3xWm5BRC
N7c0vW/Uor1rR8njJWCjFPzAGVlMV8LmJjhEJ9ki8wBUSW3PvKXa+W/nwXtZyIFd
ZeesKCzrYkuxpY5uYXAdJdwAOriDBBMCQxbifsLR2jeEJhqNFOp90WR9h3S/pWFL
8i3mgWHl7ssRvd6o9hKo7n/7kx5UD6AQAIVpxqm3vWdR6OEqM+E4RlElOwFgmLoN
c4QYf7OyPHo3w3BRI+q0EETLcJfswoF7qLHy5ozfi8HqKXt2ej+p5Lp7N6J/4eyf
G2z9rZBkpvNWV2jFRWdnh5CHdBRsu6P0spjs+Xu564rC3RxToB1kxr8LI0kXMR2G
+tdT2ISPUZ6AFxYstWI9duBut31iOYFcGebLsGTNY+rPJBcXsct93lGLudSAll1D
nXC94f4jTbV3JEjYU3uPhVXD0XaQVwUIdPqFC/ZgaDIesd6YX0PCDeyZLr091wzx
Slik+4n3swN1KOStuaHfJYdI6/zkjdL+z33O41lffymwSprJvJlFmwP4GJApVKnm
JMVHIfUfRwqxuA7CvtNB4Ej8q1jA/j1NjKFwsfe9V7DY9AkjoJBcrL3+ZWyqIdSg
H63M+7zn8TvLDTo34D1LrBuWKEioBDgLHxI/2K4YJfPf5oUJMO9lmURKdLQOgGr3
vO65yygl3a/Yh7YL7vmFLhsRF/sntTMBgmYzHb2uIA4AN/QyHkHvlM9iZXOlu0xY
zm+XEV4nbg83zrufIs2KrigY5JWQfjIQwkGxeU2O1Q60Q4VKjcIMvcr5Yl2QvWWd
3CW3qksP3OmdvgSK49vT5X3DcNv1pTvOoRxLAoDcwQau7PsuxgOia7EsIb+v601x
hDA6HWwRVNlzrnFAcCvFuUsvUYF5M+CJ2pgFdptIxaBMlRBbAeZdRFiqRxpE5Efb
u/mFdxGAjHudi7l2+/TQUGesv9+u22R+FvA99NepGoPPjwqxMA09cJmKiAHQtrxw
EoMYX5w4tXharY+9Z3AJltQVx7kn1qAy1r+Gh1e53cNb1FfDFYngtmK9/kIxs2lS
Yuop5mz1kjLE2YLT75XChBRbssdX/n7rTs0bdhmYuAOKRr+D2j+0G0vKt5DYxRLW
wmXHWSwC3sQ4VsJuy9qQ2+wdurUqI0mpmcBeVXAYtDnl2KPjfrqXw0tRc9i5Tv3I
7i+kQ3HfpxBjRt3dsBndCH8N3i+Y1kJCPhRKNGfafeLXouV2xX4JnKKesqk9BeDV
m1BrWwFpjJrH9Ahhx8cRzPs/leuVDTO2ldnR6IOJuZnzwgFAboe3z0DXyAnsKFUQ
TtoZizh1SpKw9KtxUDFokzVesLD6KQlPweAoyqK3HNixH+6RF+tmkgx46PL/JBQV
Ewub4rrz0bX79ryfuoe/MEsqN5Dr64GOhBFMcvFrsOs7WpMYRV68+DQ8iGFStYuH
aywHQEH2CcsPYIdH8YSEaj7e4rQPAecq6cqhK/Zew2RPvR6vQ/ecOVxiUvN0SQDV
aerywBiRDBP92EfMzKHMIvBsAosrMFg4V66dm5TvQASFjQ5Rig4KAyPiV3Nl6q9o
RhOZbSgBzKUGPxwmTEYc8/0Q7gbE3XDu1L8RlRvQDq3Yv/iSaMMhIy3s8GgYaORE
dcbVZEvnP60i/sFpqCy7RGmZs1PcmXOTuJpiGdc061ToUeoJMurbLTdgRV9BrVH4
zuRt4shwiGzS7LRxZ03Ky74vNY+CUmGLmtFYKkM4kDWh6451LLW5JZGE0xipYOBk
+nqnuUUzT4ruV7jxoBpyLA==
`protect END_PROTECTED
