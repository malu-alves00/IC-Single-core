`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
K+O4qm5Xy0fhlnvEsxZi/LEzSZt7Vd2gbdeeV4oqeGYPOTUT4fQbokWTZdqKD8Pc
JGF85Rdi0lTlS6LtRzCiAZFt3rID2ktJtC90aFsIRGLoJEJcWD94eKX6Xj1vOCcB
LEs5FLOdVs6KQVJ40RofDKNaiEyckUT+SRputp3wrBX9aIbAK02hIhaiNZCW/yz1
zWR5BrErQo2jwb3UIUmrbSwy6sAfevS9r/TAclHGDmqv5uEuckNHKA2I/lZ+Uv/Y
Y+41NjHm5pGK5WRzh7Pj+zi3VU7W7NG7DZPWdBSC5YPOJCcgmTGVdwwppzZlGgZi
es3wu7TtGWHAaverbNwMo8gP1jF26brK8Dcaz8vHJshECd1Jgl9OHaEVSsVOX8cJ
g57ez6Vj48mZx/+kWM0WL8Q4oFMYBtEfQQbogZI1HdM3KKL+6Cf4OI8nLQQ4QGWE
ScSTjADNTp5Fle7h7eK+nC9EDdPxxWhT0mcw2NUPlm8jGCM0StQuQRFfKptlQktS
6WHtdlixmfqVqmmwImuxJQW4jOTfHGaPHKDbT5V0MkQQh/x/mkBVzHuxiBVer/mu
6DjKoM9jbwvkJ5uQGn6mK66S2creG4EKsf01c4YxcZ3owQ9Ppb3CnE1g2GKz2gYK
dv94RmO7E9TPxRQFAGawSpRYflQKN9rpIuz3tmTQa5eYxo35VbAGUVIkMJ+HsRPN
uZ3fBjZsWzQxm3OLci5MJen6Afp+P4AHMn2jUrBpE9ijK/9NlXahwSDLI8tDNIHn
qPu4kldKX3gTFTe4u3oRARkuNaSgT6JEltrxDtQxo0cQqYv52IztEH3P2xxyIh4s
nBdsJ5Ng1UUj/iW/tDxC5VTMsks9Qkdf4XjcoUonAsxqnJsxbYFay7MbQsJd+MWm
VcwauCgZS2/YQNv9I4koSaJnruMDBvU9HUe6gOXbFTk5Qvg9d5XV6onHoSKfUQWg
DDnUDXPNw1URUc3hBLTFt7H2agnXEvpJLyshMocxYK7sUovNvJ4QYThR6JB7DVc9
W0gfgbRe4lB4lZJvsMspeExh1TEpS+Lag9fGsdpDLBh97ZmFBX2dN8LOGRqhH8Qu
KtcQRqhGy0w0IYfTJq5lMiYDcQBBSVWlZhnqWzRu974=
`protect END_PROTECTED
