`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yg5EJqc5g5P1Vuhz09+jq9NKGOy47ufbNkkve0AEhd7nFPZPYQzT3qKLMQ6YE6pb
rteGP1cIyB4qeQw5GcG3ZsYwBdsYapzIIPAllFUt8g1Y7ZihYj6Yii6uKVcdyzj7
ebt85EA//PJ5vvYa83S0POw/PmcNYESNU/REaHbUIZ41MXhMzgP/0FaW23ZA4AQi
gpqKJNpatQPSjSqieBqWOUecE8IzaXW8Y1gLAlImwHdm5etep/6OfreKQ0CbiYYr
XdbA7eSoDxepVOb7Yw4IV5d9wr4D9LPTxZvGHoJF0Qv9qK4Y7R9/tiKnikaSe1L0
oknzLLdkCPjJ+rF3fiAgiqtvyyw/BnSts7DHbmJgttM9NpWe5PWzEdjN4pR+8JAH
QJLYiNoRtl4Kq+JJ/9doGsu4t1KatXSi2ztFjghAk51BaAx8F+uVJJdOpUNWlFf4
v4zP2yS8L3VXoR8ihVtTaC/n+8A3VLSdRoaRDPQ7j8RGm4eInwnwYzT0Ugo3h9UZ
Mw7dozkzhmCLJCuQDKLBmrOqFsmLmU0T24prDKlsTr3s2iymIOHsZhE9s97fXxsi
czzGClHfykpNQ8LHocJVT2WdtuAoR5jInDSW9/ekAJfSdVJDkGJng+enA9ZhyZcz
vf2IurDrpj4DEij1AV6OmA==
`protect END_PROTECTED
