`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/Q2EeF7tcQLpi8a298EzOoSq+3bBT6n2le/VBfpgF17ySa+pUI1onSqkeBrvy6nz
IpT2ytfnqJaNrXNDI4R0W/lLLdQY3Qkcm1TgpW1OuT5QnDCOOP+o1rn1cc7znt8u
jPlZQA3qmDXkLphNXBL4Rb3oPvfA5+TxgIUK6gKVAzSvxe+mGJrzjKzulkXb3hlW
v8hspcb8ttNAB96BZVmIoTcYUMySkoucDoS0ZYQUZWzhVmFndWnMhydCTxQ3dmcG
W0Yh9cbxGIQUIPJ1O5cCZspEtA0953mEnQHqvkpnAaI/zZzngBbtushDSds1qFDn
B+opZBmCwRZ5Lji7UJs5xqL01dj/mZMhIEy9JVUSIvan7aH3MM1w2tPf8prGQxUV
7i0KZZ9sbZJUqllbCr9sEOxtygS/zZA/Zg3koF1otwN+4Jie+qTvq+/iiEcp5iCA
sgOXTmM487EK4yqAPxJnCm4AXJYcuj49coEZKxq8n2KvIdrX/NiAJCFddilHZwNH
2Zmbi9sDS9bDO8bWDQ7K9J8e638bBF4OKV3IA+EuOF/2LbrZ+0q0WJ1urj7OCbFr
MrTboz2c6N+UyCYYEBuQl6/y0BSVItMDg7YxEjtAk/tQ6OPXZKiDnprckIA2NSrd
amIUAJ6IjsKgjCRXjjSOD2XHTN8Qj/4fMRj45YXi5pFLPfxcFB2k4n9gFIuxkmwa
qdc9e+hZkTnhwP1qb8tCMwioqxqdxSePHedRu66cGVywRPMQGrLsWU01YVvmMUO9
TVj6/gkXGgvWXdYF/cm1FvoLQ4Yy7nIBV+IrjyJLUj0XesMciUJFf+Epb8dxnWMR
ThMYRMWuRQuLDVA5Lmvgy5yp5OpQDI205gqUCfKcitjKbxnuIMBTfYxUsKofEC16
kqdnIkU77wqdklNZuyNdi1r0sX9GGZjLTr3b423Nzdf3xBdtZO+2+szG7tScf//w
QLvzd/rOxafSchQkIFshz5yWBWUlOGOV1tpsGwE0oadD/+1gAU+UxwnpNoNoWUSg
pODB0g3Nn6Sa7/Xzbi0Lbyx/LwFnxQSg/UD2IxgG7FHUDzctTYwWGpvGukqpxOUd
MptzBpjVoxNEuZiN7dXeE5OjWw0F4MKgKxZF3G5dC8P/gsZ4OYhT3964ZCOaJc/4
F76NZmgc5VTI4o/L7LU8lXOnm5Ca4btG1z5037LQV9ElGzdUiy7G4ZvvVikT1szs
Pr2bfmfSdxywfTFn2W8TOFaPxxn5tscvAtGu98fy6ohp8vB0loaZgVNCghXdRzRt
dDWecBSuJsz11Iyt353J1NQsGXIn+VNUhL/XhlFmqV1/R4kBjX8LwOd4TaoDNkTL
4xV1w0JToDiO4H5pSq/WcVCsJKs8mbqZSwSiy47KLXBxWrbsmizEV9d10VgGzsiQ
WNkzKyzKGEYCswJH1a3vV/VWPo+Mqi7Ey+zjzrezA3fU0JbWeYsgb2LBfJXT0B96
xOOJtT6g5iH5tY9Mey3SrPunUEePZdaQhvLC1tgE96D7WWijYHBGxM5UtBeXT21y
tab46gqk4hsqp0zoahNQuobI+obqB/MSGH+VzndFGxu8tV2nNuyhvQ/WzHZdzcPm
GEz1glWZQBEKaZzEoIGXwHyE7AIU+OzD2UsWnNXFA80fyOKF7RGvE5cn45XasIcT
Hpr5AqrNm4Sjca3EEPDT2H4bxl4/XKZYgG0jtnuQ3CIrUIbY3+PWMDmHT1mkvGwT
d1JLNjAiof41g4RCpT7vtOElPvfcV/UGvK6mIW0uKwG8Q6I7bAQylViMW2xlzT9z
kWXv8pbufief3ebRJRb8J0vIw2IyhOQ+1Q0T1FQomk155cH0O6dr6IeDL3yVGfGB
L2QbqT2vuemjKdYsfSOIoJdW++JT2jyDH/H8g65nBqRkPj9Nx7q3mlUhdSf8Y7UG
istYsvUdFAcYQNzh9YV5kU70HUxlZuBh9c55WigJKGNxV05bWiS75Xyfkc148CI2
5iHtETtsoG7MbwxczMl7LtMC+7mES6Kf9834n2icoNU6iEriON+RSwSvSPyj0xEw
oQgatJimJyga7clUvMO2YtxSw5eF/QJ1sunHEW2dNXBnQVN6XHzwT0ZqIvZoapoV
wvvErTw6xwpX7i4skLGFS24oZ4lFa+Aczrwj+GpLALIJ5mco4xs/N2OGdQZa5mi+
25hP/u6cYp0riCa75nzsQc9yk8UL8hkmeI4lj5NUj9tNXd5nLIsVzDiKmZ5SBSO/
pQqhvEdVX7vTokNbcxyM/f8adHaUszfZase5FCdlTMbKalJYP/tJlhfBh/p7JJ61
JYGnayfFe4UWvLRwg1HZV9SwMKPBNG5s0ZLTjc+z8VISEHwCbk+Idlwh3+JdqnTz
WaI4qZhvCJN5s3fwNYBwlxJZ9BcWZR+9FLcrRzGxA9DtVTXmXFrcuYZn9nlHrOVS
O6v7E862/a7b0rN/aLDtmp8/m8dJCBKatVC1E9BXxXSX2HVU1lj2oe++hVmG/I0j
QUUhb+9I0+cPwtl+E4NRvE+IHDPNRLyGJEbLE4EMzIl895VF4umBN0lz2E8nHeqN
cUmshHpe4cHVbehMVWfQg2g+NZYxyfFK51UChHJ4spzE5J1PJmQcDO0L/+A8cA3w
i0yqss1te8M2PHE91ausQP0tTGjk16X6Ecks911YW7eflcUDc/AN07DIAFUgu6+7
PMY5keKqRQdxGhe/70eQARq86TNA2du/4DbiV+69eLjpZJlXeOR72wMPdtwSFLfQ
tw9lXja91AkAgiC88mUDT6URSE8Bxdb+nK1aei/lDZkHwDlzW842t8LVxZlWnxW5
O/6HWtck7K2R/pkF426hmdwEt1cCWXFRRUaGTw/tNBrvlukzy8xW1L5p9mcGm/zG
2L4rDwmrfG3vimIVj4Xw9VQR3v9a0I9HuTuaQqRpEaEictXptGYq6kOOvyNCVtsZ
gplx/J9uuf2u9LeruknJdL07AqLBAROhd8AsEHoWVepU/7YWeh8F4SWUz3gbFqVj
FZZ4FXJUl9A6uyUzMh42lXBFBAgrCqaZEPH6XaOLueEm+UyKmAALxWrAe2+8bUJ3
FbU75ZioY32b1lIkNSbKsYCkQD312v02bPabPQ0me7A+8ALCFmu87AhXbZvyAUGF
iu/AYsWjuT35WDW54Qdy/uiOmz+dHe7mCbPxraIDMS98A4DON4He50ti+E/HklXh
lJCAeOTDqkDgqEKfvyq+TrUrUrt2pqFF4rFtFZos+mByyJMzahAW8bHqWFurnT52
pwLnFK8TgZPuKnxFDVOpzanC3HwSDFdiWoP/vkSQA3LfsVUDPurA2lzKA3voSJNx
nedCVVI6yyjjWBT3wOzrDdF1SUWRm0lc2Gk3Xlah8ohBq2vE3PiURGuVcVKXpy+J
y9R9ny8MwQGq/BUAPIelOqb/MWrV12fsXARb3Q8/R1rvDA37Y3w1e3KhZg7Ez40J
y8qHNMyuoBDrQVDzTjyfIO9TBMQ2HUaVYMeFmQGHjGDJzYBxrPo5HK08R7OYVCnh
VHC4/59GxmoHKSMAxTWkVoRPdy0UiQUJVaLUyukF9nyz4U36BndSIOqnFdZBt3mq
nTecfKW3+kphkYb6o9Qp1i91rSSuzQ9JElW86dYodPuOTj89vG81x0/uAtFxI2Ox
5cmpkVY2NfL02yh2vbnC4Kod0eycVdwxjBMLoHrYgfs3yQDLSODEuGVaEDgamRE7
Mtxs/I5Rk6sogjBnw94IYdsX4BILndwnH60NyQTaNvoln4tnyL/bjysjooAdC+wV
FjaDF1OEfX4roVNhA0/Ffo6enGRLQ0e5E0wxCVj32jMuWrKSGtjzTmfPVgBFFT9N
IdOAuP1mlw2R0JLfzMJQBpMrsQ61pWGJDB6fGPHgrYxuMHrtnmDvnWcfcLLy983M
zuJbIUWqbU1bnLjnPDBKaPiAKUXqMxhvxokndElWmvtPA1WmWPMbl5UO6Vr9uQu6
v1ATOAMCgh6l0o7jNkft5LNsh1lEUbzZJaFfBuDyTldTAO4yFrFs14i/ipwpc6RR
Be1uVbI699W4YrnR7eMDFllOjeEl3wSrK/MN+W+oo4H0XWl/+zDNeJtmZpVZa/d2
ypHq4x1SXERp9be9f3zyKJfhi01waH3Xp2mW1IJlcAuR1piCo+xAWr/cS9xGvXSz
keb0kcLfxyRYajPPhbwBlFMmke3H+EFuX95gZG03dwr3G5fc3MZtf0xY9vmX/cjc
zsDfE8ryE3gNOQ/jEywIJWx0xAPmKHYU0yfsvAWsKC5kJyv8axoxQlVPO1XddAaE
dZRG6w1HyYE56oxKkO5lBTkedTF4LMDeOt6OpjV080ptQWjfz+aZlT+NoCkyLOqj
37ox6ENvbuu2K86VQBLgrEU7jjTUESF94LoItHtMbOZNn1AimhipMDFK9JF8e6M7
5byl+DhIvvwz9fMme0XPjKtqawAHc5C803RL1iNliPLSJxWI/e5OnQJpLpWzgdMD
kOcyATaMTjoj19A7rvXmuTUUNuRF5FE8849qnte20VN/SEbRxONvv1DwQxMzldnK
EELLpGT+RWE3zgAGnublqclDM/RLhhE6H6028Aj1Ljl6DLsLGDWeau/W9jPccOit
8KeONQxrgbCbuSwkZvKsUQJQWWP6UflkAzr1JkB40h+CMzPSQ29IvLHBnZNdalg2
beLYGAgaW1BkWpuAq2Zk4n+Ypxpc0Fi3RfmysSMy1QPBeOgS/Xwj5+GXetdtn0k6
wkD7SXohNHcckf8IO8AU3hoB45jc5WCEqgL3NQw4nrQpTtJ8GY17quLLAQpqyzZq
Qyips4vJWs9STppVk6PAgt3EbajbRttRgWk3zxhTYbabAp2p7ctP862gt8VsYWFq
t8joBywTv1YlerU70dkJCnvaJnDySP9pd9dkspWVC2JY+gHO75tJPbNzrF3ZBva9
B7gUqkDP0Xs1mYvRborDuBie+WtCdJnkeUIo50xbkcEcZzaON/Sk8TB0gwhpBlsG
uGls9DHdCVKSLnXMsBVN4KZGcyYnMjSUxyEQ6yfF4NCtfXPhLPs3G2qjxzThnujd
J7eO+tTo85zLVEV5HlFdVbuB5CklH2C1DuZDyyikgmXOmCr6C5kfmmJ3vC9OwY9+
EDyeUsyvK0sy4iSofLEO7VZchFY8UQIEpucSbjoYbNUaGFzMgh4Ta3bSn0f5q6rY
Pde/Dt9oPWJuEqDPT+uQkIKIXhhkjZhG7e+6v2Ir/Agd6EVUyF0Ql+Xg9fRlyThg
mhcXNgTqy/xTTXB2FuetW5MaNSYD4gZ+fNfxocQ205YI6pdqTrdZcRR73sPX9Bjv
tazyIxhepIrIzgyUPTYkTbESh5xEiLvnyusisYLD7ATUiEoeIlPq/feeIsVdnVVg
omufEIkGjuNtXZTceytWUHqyFqZb8Y4gnQzChoaZUjbhwFK5P2y9+O23vtjgnoQ1
J9u0AUSfbhNZOePtcGtzLk7ytmgmC4sl2En0uGCay+jFQ/mUKsMOrXrdj9IYcKE+
icLaCnbOVXr34WtzUkmE46mFYApeOpPU56Q+U0TOU3eeL0FljmhlTrikk1nAPoGW
q4qBLyHkF2Mg2K+flOa7C6/LKNXAzE+59x2ijbVgslza/lGxLCz/hJBsQvOUpKwq
b11UoFjZI1qZAVdJKhiehiZW/IL6En4WdfS8JOxsQI3VO7FNDa/iL4ptBMFUxq/d
SfFDGy8vqtQR1Mc10/GAvgpq1G/C3XgaFQsaP9j0TDNvMJX+3idha33KgFriyMnz
EM18JQFsbpNl2sQll127MDhqeDCHDrbqoQnadppaARY/Iqp9EwGemmjZ9m8VkbYO
HFR1AN250fl+FI/waheQV5f1CuRXyUF35/ZNw8kfQOLziXCIZ4vK4mELaMULKFK8
racwviWpoSXqGh2KGyraE3i0y95Wo661De8MgNXSa0USN6Zl4+a2fX0kK0EHpo/z
IcQyt2cQvAaj8l/tWNRKFkvlUWJG1t0lr5A6rNYlH0zhGbS6EqsUPV1z8wFJ9xMV
UJHf4MwCdiEp60mddI5n6Mj9EkEuawhuKLVOkKpsvoy3m6OAbniMCsIityP1ltCM
sufekzVqJCR6tYWmXq4grAg26cLikUwXDUYB7vVXh8j60g+c7mkEMFE9XvDrDPCs
AC062FMTkOzEob7yxbL+/Eq3R4wY6elqdW5Dxf9KFPwH2NjN5ELhvq4EgYaBylg8
X9m/Y34LbyorMGagB0Ij3C58lkGvcYNu7qKkeWAPlBZGhnkutvh2Lh5ET8g2H6fl
uOG0W26lnZLMQYuX4z2J5hA9UuznoZd0DLQs5faYmTPqXuF0UD1J4+WwSDQlB6PN
06qE51oLsr8D9km4j8gam1vm9j7bS36d8y+cEV1svYw4QLub3WmJ1R+UZKOdoZSC
y4Jjw/YWa9ImPIvORvUs5TY+33tzQcFC3D+cg4NGC8juwiQbwQuIvTSwIsmIGIJH
vuvn1hsJekFEhuS/XLD/oojV/hZgPpnV3AbgZgigG1O81OjbYkBRogF5TA0EKwE5
OH+igzbVUoJxWPg63udhw15uLytDjN/RoZtBDu67i1a3/eiwstg4QvLRKx/AQdGa
aawzDuKX9AJAr/omGNJM/xEAbbWtNRkK9AZIyulh4CDKLIEqD0PAPG1+PaFzzjkV
wZMeZsH2JcVxJLjayHbbT5nER01oDb/3TM85Lb7Nvi+DpMxTqUuxc3S+fMEN6Bzo
N3FAzB/870ZvmkUDJpin+5H9qZvXAh53huIBwkbbPP6NPpxp6WulMYPE3i1WrklR
zYR/F7h2dBqhFXnFKxT/S8zLNA/TiiYK+7IBqZrsFK/oEyuQftpKIFwGJHUye3h0
mNdQLODFYYdJertJO+oKjBB3qMeGiXFanagPmAS+eRkhCzZLkeeDo/fVlSHAqIh2
7Qz5mZgeuuhtqnal6IvavnoqZYn0euDAe+6eM1rQYp4RnOcStTCXU63eMMrh6UZM
zq02KweU5OAqPztFV+TxaLHLt82IDMKKkwGj2UY+bYSHhrlBnn1RSeNtu4jh29NW
IcfC/hUYRX2sAyHDyDSv65wkyaNVAsa7A0fIj79xnYNWIEkeLwcsyB1LvQ13cCVv
vSEycqKuXOjdtxOCKfWA2trCs2j35wvTd2/cztYavZDte7RYTOgT2bKZcU7Buwc8
EG11oykBxL9TqyRsEa9yvo85YKsD+OsU8eYaweI8zB0NjjnIY5Dq9nK8Ao8drYHg
6KBgN+qf59kNaUkW+CZXsJoGvNdzjaUvEVa2BzGzgeS4RAs4h/jeI9d5Yq4vnXcU
dGVe6YpyoE943bBtgEaygBKawQ4kLkAGvHgMdaxH0A8Vm/YU7HAA6xgj3lgdmKFG
WCWV8HdzW6YwVgSAjA9AZNAIwCFaiUzu8Mi5VPj7FVP9ml/POmbUen2kcOG/qN8C
NlQ5WMA1YmZkHarvmrryMRo6fxwPAlMZCdNvjpRra2D8/3uwk2sKswAzlgDNkjoz
89+1oxLarMX71FzeygQPTloOF7g8RQgW7xx01BZPkk6XnYb88J9XekYe6N4cjITe
RrxmZHzwgh9htPPySKTbywZ7z+fD5LWsYAqMhNIIAEEaqkzqjruSExCmHGQPA45o
1t3DaWWUsOh9yikC3JH3XWN2/1WdCqCXqUP0DZMVzi4O4zwpAVog9v588sJt79gJ
4wDkhPZkIJ2HFBctbdalBtC98yQGWNeNCUxV5mmxgqI/6dGzWMH3doB4+/rZeZ9O
Sjq/Pzk4kFGL5LqdrnhMnk7JTfddeFi7JnueJitE+tbaMqonGswwTBPUvWBUbpbC
FsPecJlnoFYfJTulmaKfDyfo6PDdzuq+pxjm1TTNZKRVPP4EmVAxwnPx0L4sW/48
X4zwt6k1qcR5BK0zkLSbMNynihUscTNJKOfs2719M9WEw+xNzFgRB53Ag6/Vph9L
ipxJOv0NP2BhiTzKVrQUaATXprCsIpiSb2DjikQNn9I/lXuPGTqQmKiRLpmgy+/x
DPSiVI5qBS9oD2WPtzjiQs8O3J+E+64Ort/xTBpVDdeSiTvG+qmTfPtD720N6Rut
/KWhTD6/s6y5vXmyxTS/RO+BEV63n3nEg1/CXU4G37ncR31bQwOnwIwtuOyMaF23
6aChdD49KOWu3rl8nPFEk3f5TdFTf8hId5l0Fk0F0yHduS4L6ttrRvkfs4BxMf4R
s/DQ0Eeqnlw43lQZ8OGJ9BvLRatJA2+C9UDZedA3XXXBlAY1dwkKqu9Yl5Lh3t4E
Oe5ufE9A6hePdxINcN8MQPkIyYzF8HaQTAyRbgpn+sdGvhdr7V3EjWC/3eEnxLQ8
A35kI1KVLuPJvbXWKbxJD7jI/0gX5f3dvPPkC89MvQMA4+HlaKEiVFj56hi+XuRe
NZtzmDwXHfdF3o+W4ByyDDeTcByrERDsdIAo2vihKep7COSfg+z1tIAUfy463/8O
11iF/u3bF136vsSGI/k9NDdEFgK0UougHtaj7KAQnuHf7gMJcko0BBNbF9u3m/Rp
mWtIMWu99mr3Z6vUIpE1B3cOdt9qSAxPPmJVcE0mqGbOkxckmYaxMhck3tP6H25T
luE+FpstEB3p6gg1j+VGYcMFzDQiTvafpRKixfNH3s9/+JBxVgQLPBU1Nc6946Ux
A/m8KISL2eOotaC9A38pAXOZBE7B/E3c/mPZ+2nWejoJrJVzH23HLy6b/FnrVYpo
gHwwJF2vZaCMoCUnFXtswKQn/nHhwGufb9nZSHWRRXahP/8Xsu2pLol0mFqLK3AR
zz27sas2Yx6+TmqpjcSj6YqHCATzhXxQbx0pwlj2tuX2Wbq8pdxsVGIYEOx6HeyW
WPvg28aMcR9dXYTbdmn8tIWpCAt8Nzmv2BbHoMOJw/QdAcd02wLbw28f5IjeIg7a
noo6RQsDKnO6BUNJOlLi8iNDYhl02RNHcqmzpYda9JL2Rp02oGNjs59cJwjWfFZH
yqPcf4lGQXI2e+GAEO6u/hjciAp99SdmUNsY+hdgEfe9UjprlU3dN3n6vHPmg1nU
GXQouhwlw1dBHj2FOvyfja+fL5Gfrx7lGMQowkhBIWfEQgOpaF8RND3XCT2ZIcmp
eEZV8TEzACUTb+6CUcoLCMWpqmPL4IhGuER3VK25sqDKG+rT6gAIMJWgLxwAscje
PQBi5gyCoA/0fpMY3lFv+h+BbHxPVcPJS12UnhPuhcDKwTp5YP5AJn6BHEUlfxwD
n72fUeLuM/vWg7X4BU+Jpb8DPGqvAOJmWW+6493QldqPmv4trBA4s+164hIRFpdm
FvThA6sBNcRMXOIvCLHQmoxQB4W1yCP3YaxPv7DoErrEahcUaQKJ02DVWdQzVQ2c
mhrQ9rzW85txM8iPx4GtTYprpzWIGlrK8Pq7ee2uyLkUJc6niPPdCTF1LhQJ3cKY
A7l9OV5zvtlszkpd/yoeO8lPt6mvk9I3A2uOnSS/G1psB2oEVYNFxZPg4rtXCjal
WGC+gYnFN3Vr1HOVUkSmmVlM6iszFsIrBv7LVQA4e4tV6H7JGYyVPPCF1zr0/cT8
X60tpnTLs0m6dIcnW4GrMHoG6daccR0t5IaaHe94MMLqGFvzNxb2JNos27FbkS20
2THT9ziJaD2mhP9InWE67wNzHSnLZOasjWcM6YuBc39asTFKuxzw9rbhA7BXxjL6
cKhZYvegzjllzwY89PVxly6Lnqe+mxgwv0ee91fI3KW+vuTRNB7M67ZEw8u6VM36
1jKEZGz/jbwwD702XRQWnYBfroro2wDzWiT9PNB3HDc5DBCrsLtCORrH2vWe3WWx
eaZPcmYeG475NF3/sG1V0IzAQ8iS5dzxSe3y253lbos3+9qgyHvR99EtPh5M2sLL
LWXXtzQjgbyaMGcVzVddDYbziCVRDnwfloNKN7EBSiZ8wiCZtkbSvSuKKvdC0RWB
pR5/ME63R7dz+JLzdUpP1Qy50u7EGxZ0IWHqNmXwjbN/LWx6VI0yxoeWE8cd+KCd
7pJ4/FXgHMm6FXeagETXkZ4KH+fZWn/ZS/xompnzgl5LAx9WvQ7obOYuhbiv1vf1
OP2UywRmoRocJmFtGRrREXxzovSq6QOMoyK/48nGXcYUfOMNEDEan25jyRbVTYF7
z3S/UnSJowBZ7O9tsSbrEk2mvECa2OskXsR2LcrYGt4awGbKi7U/ViprU12TxLrv
9A9fAT7lMuRjH3Zqho7p8hlTnUn7WAaKVF6OVU3hw2Aw5I6oOqSWjZQ377NR8BJG
tu0z3r/eeVJpTHR1tu5rzx4Jmzx074nu0uMjir3YiGOsyZkrmCCAltKvSSPANCZq
PSdX/IVBBUGxsvOgX4vo+ibV7Rd66C2siyk17xameyOAj9C7mpqsKuuXAYGhlSHi
KnuFOS6FSyz94p2pWzArh/ve3mm8YCpgeMXGD/AsxjeGNJpMcK2/fYJEraFC0Tt8
jxP/4Jg9daMzxclqxI0y/XU9FIDS4p+Wh6zOfgAbV2Ph65yzK0JGiaRkryxVygYR
9eER1+/ueZ4yPJkndrxqvCB6g2fjwNMvkqIob4NV3ReG1PmDKiCh3Gzc496OV4sa
bVPJEWphLNMLbUmGrsWU2cL5Mdq8g0R/WZwi/eZmQ6bmxKIqmf7+tOq42pQxSUMO
8A+t3VacGbI7NnOSfeWmkj+QbERM3ciLgBoEA3Cw6VSdbC7cd8bvHU+WoOPe3Rf7
PeIrQ+9VGrU0igMd+iOtDEexoGVudcErD8JUHMFBuLD9HJhkCKq1JgfPs0aE0Oy2
YtK+Znr7T75XgHHs01zc7xywKzGPg6SsaQ9rf32ofdpDKJJGtmYSpMAXyENxfXZ3
HCZHRC9Th6NSUdAPwLh3JasqcCBfbR6FFmyQMl8BUkDY0UK57cCJh8Gt96ssgFAy
BNhUj+/XhhHq165nGSbSp91FuJh97yzmFG7ewa53bVqPcCpz5Oi1nzKsSrQhIf8f
ubbFrRKzR0jU3M06M2Te5UNEzMOd5UTes2iC0qNK0iiTWhuxVJeY51Tlgtf9xLeu
15m6TCKPyRp2QuDJpb3toyAmtGDET4opx3Tnc4GDbaTR6q7bceg8Ao3srZEPTyOA
QW2oKQIHKrl8kRB2zJombg+mObX/W3RAUOFgY/JtA+37eMA8iGzrKucZcq4/9YRs
B1j3LDEvWBfvxfFeL0ldDL4i6t3WM24U2DaA7VQcmIS1Hlxt0JNEQ7otPuy84+8Z
2sgLYdN9YoBxGoy+r+lf1waAa5iPmSTnGdFHLndbUnw2NOvZRS7prwbAqQun+7xd
ykea/PDtmGXMvOQqc5fo7rszvZa46b04RidevVrF5ImpWI0zCXVQxtvBpo6WAJtA
wfI2pfpXHcC6ni5qyFiDeflcxjwqDCE/naQuRTf9QyfsngIn1jxAsYfg62rFlTOH
qt7taKTdOHcrwUgEhQjSw3e1bhF8kGgkxmXeQSfZ2Di8s0WCXLxjX1MXSe0u/X2u
GyFq/gP/LmPXdbl9x/azglpGmvF2rzh1tENZ7Kc/1tUN/MjbmE2G2Fk6s7bT+hq7
MKGo/7OYeGCRHlJJXR1VSM/1Df7u33G2L5EALja+0BbGKk+Mvk/xMwiBkxRXOiE1
tHbamfm/l1goK61d0n9F1Jov67fFyCtAYAWkDqTFA0m/4Ewuo5MXwxHPNToVdEDd
eF67YM5g0lfT00ICzGonzBEk+0TageELB5YB19NZgTxMck1Rpvw5rjdUJl0h9g0z
uXi2GcAKchzXI1iKC5feBeFT2Hr8DBP3/jZ+eyLWMZ44hB33IEz8MMu1ndQ/mwiS
0IYz+ILSKGS2ccqolJgHIj9YpGLLdM2Mw0FBecG9YyEH9kV8rIy1/SprheXPgxGV
+jY3qdwNNFAsfXptYKQPv5cLwjKoPAlR687pvtfohmidm3Ksp0mACOxWCU0xwLcJ
M/28x/I1DNroNV6k1Xc2yo4oZMNJ1+VTiEQhAFaWm4dG4xOYeOOiyyIacNUmeqZk
gcquczBVvKiB5sAo5lvPBH1CcyJgGbhSsvybGAmNA5QwrCwwrSGwi1EmNrwSTmaG
vQjYKJV2p5gFc2MoeZvC3t5mbOdRajpQUpAdn8Qz9EXZiNZ8tai0XNDrwreFn/3B
EbVGoJ2O0FpURXvThICefj4MhxmSa7Eks1pyDkbqvH72fJC1PI9Toa2M5CE97LPK
X5uuKc3sGKLJf3+yoF4T6o/3YMacBZnThZAGMnKEH+x8Ar7iMi3QZVH3tXmV8yeT
dZSkO8sJME3rV5n2Wa6dpoQhC1sOLosi2fqyRJQUMkdeXAVAY5xwiLKjJ4uf03J7
lXz+pOMy5tCaHOExkOWnQRJG7B4GmcpAD2z/1iFqKcGMpFczpKpA3Zn3fVbPQUnD
hNChQYtaTja8AUycvEwvcZoocZPEJ8X8A5W2MS4vcMR9v12gaWmlfbdWKbEjLKYH
/RKEmlBgKHhWlpV5qUB8G58AYyIGK5rF2Vs6OnOkcZR6xlyJ89/Aj6Cfb2Yt6E1V
+hzCVC/k61xrc4z+Mnh4o6qdqNfLHEwO8tKnD/Cbe+JgT/vxcyeJwWkUDL2dCA4H
HcDPRopJX4LF7xwITDy0z4ET8Z6eve3Zl3c97Q7Q7Wf6SootKNeDfqyEDwhXTk65
QK/TdeoI0eSU7yiSkHbD4kWl3toqDH9hKoOZ3olmMQu/u4LYQCp1PQ+XMPsV5mz2
BCk4VCggttOLdMz5Bc2mXcu5jKFN6Uhd7b/l2tfodEFl5l7NrsmHTgT1mpgrTQNc
XZO0mTxcBZYv0CCVEwvbnb2NbbdtZIQqFOC55mkom6GbdW+optQ1+zyjeq2webWa
cNNMH0ATLOSl/ozuL7YIt8u6FAIPmYNTyry6+/XaJAA3N86xfBD7BKdhh5/72NF3
BHIm05Z3rkNq45/S3uqDPBNBj59b+98sRcVo7ZCXlECEXyQwTBxZ6vWYe5r5nxfC
WrZwvT9h/3vRVV2jWGFZuzWBFgy5hg66RnC1V6FfY6KsMTpM9OmmzSxtTVX+wHpX
4FFwfIZRGkbU+i7RO5OkYXWFKdKQmyS6DOZv0Z8kM1hGk2X5VtE09bXRFD66Ao8l
1+ia1i4/uN6hT67s+Q44RbuDxtKljsh6UvcXTcIxSvswELGl0bD/cEmwwRSbOUCi
8ZF5YCehjjz/gfedA0utR1StEi0XvQZuTbPNPRemHz8Pa26bgiz0z0bLSsAuTBu8
`protect END_PROTECTED
