`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8BEY65GVmrxc+cpEiWR9y192d09d16+rvdutmaC5xXWB5qOM3ZOthD6FilKCDHmV
lJ0ypcLBP00ckBJYiLXgOUp5kOdX653qPow3iIFi04Upqzf9aa8SgaAuuy3pebaR
c1Zuy8S9nn6LJtTrm/NsvixS02kYCpKTybtmwxr4iCNPgwAfgLBisj8JyuSN71S5
SeyWj+Kc2dhRws599B9dbWcymHXwMaJitSY8ptaj7mgyEY1TerSxHh2jR6b1dn/K
+fKqicLXmsPo9pLZs/vo0piwLnTHd9rXb0LGAYE8IrHO32LBdHdHuRQ+sHn/d/b0
iSXMmQJ1hmAMvi8taLN8HlQRoe75WOREgySs/dQFthLcSsFosSGRpxXuF+xok27W
kTcvIXZ9lTyqsVuHAAonryGY/hk1VPdgi+bLNM78/25gdK+2LPkr69ILosSSOoHT
dO8YUj+TvGtPrdLP2pFRo77poVabh1r/2cT3XOyhRTh+XSUFS/mw+qBxvUM055qn
7GoXq8nJgDsB2O/ZF2ZNKHNMMBFpO3N7QF3MYO7B4jnuaIm6YyQRSh6MP/pJku7f
4yCkvAS0DG7ll4LFAp2Wl/w3hkvpCK6AoVPeI+4ATNK/meLK/ZSJyjCLxho01QgC
RiHK4UiyjYIKgpoBptNcn1lb4VwN1NlsGQ6McV4BhTS1SmPUqpynXcRy0Cpz0CY6
JLMDEBinkAXzd2cYGR1XEUWzNnw0cZrKMrR6feHeZ5909a2O5BL1myy5vJywjfXA
vSDS6+KCiIlh+FDEO4WUvDLIy5nklcxbZn9jMpSv1z6TR6KRtyVjNG4shJ1B2QG7
XcBkza7LwqHnoZ/AtOsRNZbS9Ghbq2cI/2TFw9dbd1juAukxEyGmGh4lbwA0Ef0g
4x0KiUKboRTKPj4nTRILoBm4OJhWCF9XrAqIs0PenODyOk6lzH5XhGwGOr65yTIF
SQxmdbVMjQWVXFi9sMRKVAjCPXT3Ww0ztEN6olKr7RIQ3HjAQBNCq2FeQIA9goX+
M92qD4OTaOruyaUyEe707Vst8pN8DggxjnajbYOG12cqzNXQfyeKpdbRxAbw1F/t
EN7Tzo8W5+YDzCdeJS1A1sGTosCTANL/bJ+dE5MnSg3AK6DsgJPidnAWHvnuSSwk
g5TL+KHTP0CAm5VpKsls21+PqdAvX75ZEmEA/2McuNPGdIqP5yJK4JIEJpef8gym
cu/9qpizz5dELB7bE1ACHkyI0VOZAB3iJSP5pxkfbr1NBXc+z+UH21KarGP7yCGN
OTcU3oVWeH/JkcporqyavP+AigxAwnElbKGgWYxsKpLMvUYqlAWgs2P+2nhkSJqD
byBr3P2tPYozDT2nHyi+t/1IYu9UtOnewk32hB/TX2YgljLI2NDxbO2N04tozJqr
7L99YwBmQBZN3H9jNDa3bBhsllnAYuGDtRe+gmCekG4/4ICZYPWCDIJtXL6nooOR
qTHGmgvNeT57F5TLCYYw34KojVkV6yt2AYypnq2aEZy/b85Fh/JTGHFRI2CYXhDE
a/jwHQl/ROsUbYw1iC8hDfzyqBm/powD7zwB+nhmV4Pve8VWnyHIDRfPsoq4R66R
RMWs2LAkgW7FxQhLxOmfMiSqPg6gtdjdQh500jHQM8Eq4nqmZapj9Lp0nopPImmD
cdvadK6JEWZkd8/9ITJjeWsGU1eK95s815ODQs0vhCpU3cf5Mb1iLDS7An3pRwhM
mCNjWHgCi68JiASzQhUbAmzJbgkVSRN3hnmyYQ/TBtyluXSGK6E/JgMO4TneLgJD
lAlK8NgZzJ1Z5+yS6NDNuLyhhx4iKHHTHCO/alrRKlV04rKu/wji7IsFC0oZWuB4
ZmN1KUD6eAv98LoBocrI+TzqtJvZES0Bg6Asi86FZ9XVSkv9xX9rpJOIHdk301AA
CI2/1Kjx8igIryxVPt8UOgJfAMTJaBOAtjy2hXbii8fu/+SEuS/ahw7QTYX1cZaB
aHnLpSv0z1ZwRijrnFiVqTLLI/UbOimNJ78PUQvJg7r8Ls0oEV3eF9HelabZGGeg
+72CJiODPtbsJRc9j4BqA8YsuotbqyWW3Ja2BiAORemUJUFmM1Uavy0bgjukbkPE
zwWlCuNDym4cmLgDe47g9QxSa8DGwmTSVmUeJKx1iVmpDmFsQmcmPlQg0f6BgLPo
5rDf4VjJ1oy/Xtg6EsauxkGSV6ejUjx6Cnr5cCW0s/5mo9fVrAvk5bh5Ydrh9u35
q0ofijZiTeLR0UPasKtGgOETpXxMc5NjEOp4Cjs5MOpGt4Y2kxiBpEPLzwcEodnD
Qi3zNnqGQUlD7LlpICjx1/vgjBQwh/O3645QBqLzrwBX4Z+CfsAVVgLz6ja9Itpg
CfBk0bndsPE5sAxRF+JujhHQG1XgxyyjZItAOMhAj9ndB2QM7frLLuzr+ERHJ7Zj
+NEQNOtYcxPN3xk3PcEAULkTz+fX0Lb7cHCarGtHkUAN9IfOgH0MCWZwbOmj/WiN
z24So+3+kAWdrVIhg8zhxasZHaMBtVp/RwsUWoxZWXHH/a4E3UV8W4vPiazB5KaJ
mIq3V0wn0Xc+xlKYMfisi4AMDBwgmQ1onrZuJEZC9MuOWIh4n2PqJoqPFUTpNxnK
9kDSZ8kCHyxSaCcpMrkxFqaxRgqkNcZPInNQdGkrWggd5U8O6NOmhMIfFkVVV4a7
R2K1+1Ab6XoN1vcOMoZY01q+PRLQZWUapEBZpKsGfkfb69t/gDW7a53g0d+aIUFv
/noczoJJoR9gAtN/63bOSOMvkNoW/XeiUPGqWMpiLHZNGTYKzyPyXlhiNK1FV8UK
PfqsZIYgMZCdlFsXVOLWojZ7biucBhsARkFKjiHilcMbOuPR43j6zo55QogE50sg
jgj740kpi1IRlU3XEsoPiMzlkCx+b/Ahq/zMqhkwgY09cnPWz/GQI0CltMfY9/fW
NVsySqStrWG4SMclW340uQhubywLEqzwpXJkj9sE3WWY7zCAJSJm8Pw4d27FMAG+
sxqhj+uRTAKn8D1sx4MvHGwIsxFUNDc3WANQ2c4u4hXCOhKi8jpMHWSIV1T7q7Qi
fnadmR1GGp66CYu/3bXuqefIMRjIkFXk2UrzZa1OgXbt1U/ZfHJxeJ82swv+5x9L
9AZHl52KroGKBuujatMCco9BiQjSMW3gWSXkxFADw16ZroaolN6zDwUQyruzZQzs
cKvBfFOBd6aitztj/USASqJZsvuJb+rN9PQ+LEbiYg8tNQ7aNECn/nMp2NDDGy7y
i/HDDWxSEZWgVBBHb8Q9SuoK96OQne2SmNfGGitWViv+JndG9Z6hNeEbT3wjQDfG
hyIz7d7PbZwMJzC7M99UlOJeYeZ+IzdyQ/4yJPABDNuoo3Y9Yl4xbd2nL5bPdc2Q
MXCXpNfbePscaSI0rLXYW+JM7jkYlFsUGazw2MskZSOMAxpy3SfcCnuG4IYfHZKa
NMp+S5GWqeRFwdmYugjLOGkTdxfkk1sRm1PlFTWgt0+c2ppWaeui1fbShA1T2eAL
CorNjv4UwBDfbXeBZOPSP4Ie51BHCzopRrcosfYb/iutRuyAghAgvFlY4jhbCELL
j5ZuMChbz6cqOR/NjZR8J7ebr6Rr+4aIZ00zwFnziFQKBDvdiwbvVJTP02uR4j3K
MiyoW8pUNuU4k7fdmZ8zyp0aFoLhGLYUNcswZ0me4Ycsnkk87rrmPYygnoSB/lDL
Df7kDE6RrDEnMBC4skh20YPWuIV9k/r/PI2iU7Do630wdWtbi0KUYr9aD+Qv2BEe
pHDRrV4QPZNGeBuNloiD9MBxNYAs3FsUzOcaiZZgadkKYPRncKdY1IeB7ZNoydvQ
qW/Vw/03wPDek4MDINvZr2xO+lDee+aK1IqBcmbCJlT7bCfDFB5BUkOwBLGrtAXu
QvlqX9QHXgKSrJqiVg+V6trarCLsBQWUgpyEMz4qo3RYl3cNCXDswd7MQrbCdeU/
jrd/Khmlm+O/K4SmZK+30/s2vgVVOrO5Aiiqbh1HcV3ejMZtr9czhPS39P7rAN+0
GdS23zAIreDeNH+ct9rFyqIdBjMi7NLO3UwINTa51t399tsYSHRtw9uu1drPIDhQ
4Jl/DWBoHs5614lX1+rYmg2CPn2QN0OxJBZOi7sPduAddydrI29FArk/LQPjoJlg
jIK7iVDmcLOmTU0mpLPL6OJHakNC3VfNmutxxBwkVZOCeN2WG9MlyfshEK+1clQ9
oNq8sQ0XjW8h+sG8IBmc6MO9Bpt7k6jXwGXSh8eN7fbEb92f4dUx73AHb/VfOoOg
WXmCxeBcObedDKTZqV1nRGF3H/BS7f+BCXli7APVgNWwuISzabqQmDzsyAERZV3t
oaQ3/j6ZuP+AhOq1B2GmXP4sicJu6abdqRgvedcMn/5jDhoO7uoh0DDmK3eHq94n
dtoqOnk0OmRDj6QAyrKs4l4OzwPM59YY0dntQ2W71XxXmTOX0voCfIr2QBTX8juh
WZzITkkTjFUYvLvKj3YKdZQADntv+KSmNF46pKjDYIT0brXJdrkj5zA06CubPL6K
4OEIWHfP8/p5AaHaM58a5s7OPoHnp5F3of1wCVvPozw9OVvA4VzCcbNt1DQvBHpd
KG+MDGNEdY60XG70xVZ9BESmFgvfe6YpZi7XKMorbjbGVfMjDUlMXLqDmdEzlUN3
DhUU08IIJ3XJFB1JTTNuMvXB6a10bMIW4hAHyBjLS98dbYlbRDpJdseq6s3oVJIc
nNI7l+0epYuwE8z33rRcM3fqQJGJZm91dLnPgk58j+Q0/GhZU5W6B2JjZeubG83S
pzX8BumMwsOukniz7EK6MtUfHYDy5Kr2t3k/nMfGa1zpSAov972/tTopA6r1ZBop
XvAGzxgbijttBBxCJlsaqyPM6/ye+koHGXOcRknbe70XbiKowly+o2SZEbCbJXYL
H7PEIDvTh5Qf/LGy8R1BHVMSGnFiaimkXJPhPVTzeTdEVdGzkii8gwGV1aqawYcV
0RM77CGRJydzJAA9FyCWgJ5Vslw24qIDN6/qO7w2arqigrEvNYBz4TBsXj4aWihZ
m1I6mSvTgvdJOzjgKblX+9eFG90pN2l8P9NgBMpW9pohxSsoJHJpRu4SMaBfrTRD
R1onQ6hXnzYjxYMbAbZ4I6xxRiixcr84qnaq1D2ztdnYlPdK6yT7Q9+2yzC+ZQBk
O4IvcTWVr13wvJNsxhvPsGq+JEJppHEvEZvzK8nTIog0fJyfTay27U/OGcC3Z9kx
Av2K7haeCQw5pveyNLSw5rVsFKEnJxWEdHgqV0eNjN8Fmh/p3iqrhrTwk8bfVUhl
GIDf4KSrs8Xfr5DB0n6rXDbTtvlaFch16gEmqj2uytlPxl7XjDsF7aWul00cgONv
h0pGI7OKmx5+Os60jnF1JsyIogxo3eO8B5wJfqZc+8gRZZT6IVK9279VWYCbzfSw
0YLVd3vIDvvLkaTdEcTzTH/LZLZpSZDsRgTB8IFmnLfiHdhw2RxlzF89Xuy76z2r
ef2tXGtSfj989eUxwA/82+D011dIccxHICEQSvMzkTMLv/J43JWnaZKt+b59qao/
Mz0Ko9eAwOeBg7dq/bQ7DZueM5AYuoYuv4iOd3k5+b0K6EmGJn70/0TatjKjMmAb
8IEJ3qkRaBVHLwsYBIlneRO/TrwMLpeX8eg78S13MLh1bgZNsqTBAaYCyJP8iswL
na4XGye2iLKP1Fxgufj/68JRhkS6PG5t0+X7maK6riDtmkO/M7IT72TJrJdNmQsW
SAo4S33Tk4WjoZKiKofShrknQrGLTmhUVkfUFDIZHgZg9IZeWmm/nRDFqivReO6o
ncwSWn/7JNrEKNm57HFzMAR34Ror6dvfK/ir4ptWgNAJ8T52Tu8M65ShB9jgTHwA
SpX443YGnbp8+7XLKNqYtOpKyY44c3+SOT3JLeQsA7jhVWmoPk9KgwWvvHp1tuTs
+FOchSubA3+mc6j6t8nrc4Nc+EagjOsqBAy+Qd9bZTeZ48NFkELFHPgwyNp+gphY
ZVY2s/M0mie0xdnHqgsL4uYzk8/os5k7pygAiV7UJzbN1+de2HCwc0dJ/Umw+TFX
kVHQOF8ioRMfj6H0r4RAEgnyG4KwH+6hxRkfkIb8Q+i6q0GFJGJ4SgQyRWIWTtqy
wsQwDKwDrF6gmy3JwfHHz4WBbyC5L3akpo/NvyqP0bgbh5NGm5TeLDyTBThr/UoW
hj2lmXEKGsuE4H37PuRCMnTGycX88g0PD5/MSuOIT5VzKmO+8XLhHyHsUyQel2ah
1/0bF8BP05gxV/g9WRbI9lgr4nNUBLfYv930cv5exWFpc2PMJug5/CjJYDvQ90li
h0DZnIQMXeZItmhgSblswFpAGqS85QnCMbG3M0ivZHs8QwKJ/uHE/jNOLKiqckXS
1SRU1U63eywwiyuSDLQCBQLz/CnLbgm3+KV/3UfAf1nNAKSPVj8+26mg5Tj/UZCy
EvJjahlWDXkQ/ATLbeTjIA==
`protect END_PROTECTED
