`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LZRlD98d1756bkU474xEV6HQ60M0DqxLMAtsN71OHAREhCsIVE5mM9joD5M/mP7w
v3OLAK3Dw0UTf71IE/dXZT8QyE9hFWXYxkJSQqDrmOJdEKjaEQFtBiJhEZP4pjOz
0Mr2VQ5gwuFMMJ6vWixyN19rXNcqd3D5wivQePfZ0Te/a2s5gAaeBqbAqQOm7V1H
j+F+sKKQkMMvvpwm77RxUUFVG3uVsCvQ5jUNgJPORs4h830W/nU2goaPbPPfrmx/
nYkZZ/wrZLW6d1eB6Vwh1/HfSO5ZNha3WVKQaT1VyYbk7iveO4rSxq3FWQRUycfm
IeiJFZD4IHTTJm5jbYTePtqIM95Vnavac4y4fxhbNUtgySKX5L4UhFA/K3UtO2us
OVM6lf75PeTKCGkeA/o6kODW7EhGNnYL5sHvELXWjtF6v3J+OaT6JEMQwA+y4W2g
HrpsHEvsvsNw32bzGGLQSGdDobMbe6E9NgONCc6QDhu7DBoJuSNaSJr2u+qXyQRi
Z/qaFnTT8FOiOMcmn6w08yAMM+no27aDxINAAjaX4O1unp6gqdW//8xMJ0DG9utU
TQQvkLErtEu2wMVCDJZulwQBoiHeGNmL7EESwIiJxlyykbrjmZ7yTI/9NNTofCwI
9QPC8b+PpUnji53FFPuqPUF4xgJTqTcFty4ojstAYo/1Oq69YkchfM3Ww+w6Dn3F
sodOXaHN9uF165ZURn6Q2N9zhONIsJ7Emu3sj1T0gX8n3DGfGbIA3BVG/HRSJPq7
I68aDqW/e6WkpgK2Tqyizb4puWeLxsS7Pr7kv0Ap6iJVD/co2RLIwKGwhzmCS5zn
1ADA2+xES7JMXP9Ip/yruJbGk9hbnu4O5bGSWTtvZ6O3JqR2PCJjsztiOD1KFKej
KUO4HhJnE3AA0itOJ+Fkk7ct8abU5mNgDWo3GXfL7vpXMCX5af5XhiDvO3VFqF+4
4FoSn6EtRKrvr+F7FjLmXPB3JIoY4NHNiyse83zYz1X5Ub57wUdZfDnSLVXv22IN
ENvOQ+vp35h0NupDoR7jVpSvXnkrEsJ9y6CxrHY1oMuAn+K9MX8S8VtKMMb10TTz
v/RmwTcq9Xubv5/v8dncOmg7A6C+ZV6QHNsRAtJ7RdGPhKZVUQV1TVkDUxc3ZTCk
jxqdBXbmycS4ERXxwM4oUFNQHc26ZGjw3qmJ6kUBOwQkKltpVSZTRjN3LNZErC4u
ZAy3AMqMebdq72xoFtQnVy5HHKbz1fcuEBol39UvyK5J5q4e1RhQqUwKrmD2A/s8
cK0EwdIr6RAPBA3WjL37h5EkCAljWL+t6ieWa/kjy1eA+fgyQO8IO22x3YrwGK4F
lOtdwfjAAsg7f0UEBCHQ/ufbVERicpqVbeDn1BWBOfdoxBMSkMp1QO2o5IBcCdMh
P//9vFximTb6Br4ZOs8HlRDo4tN430ckp016tjpxV5xo9m3FATYhdTijs/7WZF/A
fatFLPZeHLC/fhkQW8jlAEcvgLZBMo0LjkLg/Qh+oTlIkc8qhj+p2A+Fqd5e6GgE
hjGnEXey02yRQ7XAIJk8Cs0Yan6xikL3yUp+C2wq3WnEPcySHOq8MsRl8+k3HzZW
x8k0cmrbe5R9YhOTk0CtcSw3QrNVvDeRG7vq2ylxb4CQowrgvl0A3ibxGKqE2ZXh
p/WHqqlAqw1Oe4j5OWMlPgCv7L6jw+fBHj14crBlQQtxDIKDd+gNbmzD+LJc0D3W
/AqKcOhZW6GtZGmHIcDZ/cLcvtF/oNrQpSd2tD0pU8MQRuhtynIBjulQMJeAPpSs
mzvUL1Md6RVkufaCRitBC1Dc9nlssb5KLOz4esRBRNaPUb4tYUnZY/E84JRy77rs
hlq+k6MeMr1rYxqOh+HppUvlgakq6KYKYFKSNmEiFU/SLuRXQL8igEyEcOqEpMpd
/I6v5AUgK9pMTCq4piAf+CVEdGxpjJeN/HNcfutFk+I269DaqIbfyeYHb43bka3l
Y7iqLrFVMDoc1P4q+RWeRuHXFNXSAs9ZlcLFmt8dG7WA0OZvXRXq/W+RdA8ck7Vq
Ipu0KVaJQ5kbvUWWS9BWGlAweOZQDiH+SVE21kINHJZ/1Cie/nzouu4NabyPuH2o
IlskTH8kvMDbdGV4UWJDTMLsbtoVsOL+K65X0s9IROxnbd7I57VfyU40V7MwMLMA
1Mt+ZRt1eNW+Gm0gjZOvbODXpo7x2ft3CMKKiD0wDP5vd9y2oiLZtgLIibPcOpE4
yoeYELUQBZrph1k4Heg/2gppVV2Am0t4pmJlqxeIJWZKNE9CF1slhrveEdYZsZ3k
dAGvWeisioC+2rPrJfzSUQIWhzZMTG7+6YX+Tfk/H4vJG7cToCYInpAsCNGImD74
1AMiGdcQ0PKLW5fBFHUbLx/luw8/xG83vmUwZhzmo0W3SJnxAEOPt6JQl2shjpbU
HR+L1cJDh3dpGnhDUSu9rJNwX3wVBrb777pSc27CR8OyqI1WkfuLJUveHA7FX++1
BSFPHvV/wX+GRreJK3c6oD5uEkQ65j+1bU/Bgz4BL1DlH2nb6JJUP53uWw75F12B
uD6++YqnhF50rpCN1bAk5Q4RL7D9H8cP6lc9C7+KN36JCFAJFR3gfiDNQrjZWsKf
yEAq8MnroD5Y2e9/WHCRf+jV37dFE1eBgbxViy+EwP9duQTwHs4tO5TvazeQ6MjJ
kWioVXEsm495CPTZbGSWbMkMBjjVpCIOl39IkBUYweYb4NwzekJv1+7yhLwCasWY
9i6OGBupsKKlfZAMw4pe81Wos9PcbDKDzaGoJmju6veh9K+opY6NN3uUwTiIMdsc
U62GRNv7dBsmeCyiLyNgK7bnVkkSlR8Ak/RO6cgva+u7hsvJlbhxoDautvzTUlOM
jY1hvlB1KuFAxbb6SdFxMf1Y7+2LvdflKSSyODdmI0b6bajN5Coj8pfUWN7DLtXL
m831/b6SKJo9wIWEGt+//hWZeFoturH3suteoRdFp9iawyu7Oy/Gttf+Q8pdg+P4
X/VkIewYDgmGakS8dR4+41J8GkQykTnOQGaRLTU8Lk/IeSGev7JzFWfm1hCsRg/J
+sSt2lhI3kThjndB/XWycILO9Q1Dfa/uQgh8Avrb8PqkUEZwuPWLdTAlGpZAYtO4
ElJkheJjBKGqepquZV1hBxDELwCCGdEINK26UlDZpFDygR3ZTfdmlD7BIn3ISKzO
kyFCfPWPqDi4z2aD1xahkm3L+eO/LNlZINiGt3EmjXTaFZaCD6s+8P8A4JNW9KpD
Amq74FutexnR9yaD2tLdDc/Rq1bTrmDnEPyvBGOUBC96ksnPoeZ3QuLEOpVV4ArX
iCX/ycqDwQ3mPAEjcykmQHNAsyW2j84PrGiGIkyDAv0hV0CCViBCr+l4P7KhANfU
N38X8yrSiRxKwEjfklDZNEgxAOu1lJTySjfSTI/f3wh3tUSxEgxlFsoMwlhQbqAN
yp6Tbb8XfHG9fBsPuqxQRZLxCQ2iZRKQE9q1J5FmCL6fGwDknTkjv+56lgm9SFTv
HFXwcJ6ekAHOPIpI8WgOy8i7BBu9yS/ALq5QampQ+k3Obj4bb0H6sp2bO1urc8gd
An4+OFhGl9wunjkQqcPo9m7phjUZBtTPMeodWSmZVwW/OU760UPejkVf8TdeOLwq
93RaRxNX2GjxPun3CH7HDAEZlXw8IRYLE89s0z5BwzxfymOYsiRlJDPJiqqdSXki
/wmBenw+7LZ3jJvAmyyObXOkAJflKx1iFcltA8BTEUWCWtfXr1BryVtSxJD75kYj
0mjGEIxbJLrUTbX4u12WeExarJpkfg319cevdchb3EVF4vYujK9OKj31AcabXuvu
Xs+4H2+yGROfsz62XTyWGXYAg4UsWyJIvAO2sIErildkgz5Rdl42fSHe5wm93ILq
9D/kRdy9bPszvNTd5tGd368fNY7euPNPLpqHIEnXwqD4273kS/TzPfgI++EYGIsa
0FqWneIltu+q54Mhirsc2AyOdoYZw9XPrqwWw/8nSu+xyi2EzXl8m6SbTpypN9Dq
2WpXv64cqqM5jNBIVkmX4YRobk4hZThsMr7U6P9SUjjXAgs6+EV0goouq0ChruYU
FvQmY2hbGdiFovGCSMS8boGR4zNsL4QSOlR+hXlREY7hpMp+nJ1N8u3vjlJJdY1y
EgqAOsaUiHedhuM1/dAOoVieBfSU+zFcDFlfuVJTZ0jQJfSp5H4KNFaEIWNceEXb
`protect END_PROTECTED
