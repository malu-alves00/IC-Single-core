`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lDMVKcLjebH79V/YafEtVOaeqMPtSJYW7ctdqIh4H8HwXgLccD3fqpFR8vEPjYs9
6c2MrPY4+w8QHtw7/qMCnhgL9Wh+8myHDd67hXzSSVpMqSG+rWg11VptC+K6Y9cY
7BoEc951KagwDu/ajj+IHJDJGiNTG96ssY+pHslbS4GnKLwcEGutdAzBKVb/NDDz
kcyvSBqVvDB01equoPl6zoEZZvbnsGPxUHjX2aVEWqsTM1W0LY1At5KGEYr0/cLs
b13k5b0Juy2DVEjhf2A6H3IpmdIBwhz0lk0dQHupWz9PaPS4v9kzYdHRsUs7fptp
OVbqsrEpbG1YlKkNcrWqGGJbEufqt2Kt3ndQo5sWsq1OBi9xecTAh0hzNJmHyhik
BblPf3AeaHlc4dqC5bwGxYTcjn6Pu8wmyuOTRZh5c0hcsJ7r4CV8URVbiBnvQX35
6FZuZGF+GYbdnVSime0etgRzSvdcIckzjzLxn6dE8vfjJA/OzmN7EWWR8Jz/TkIg
J2eGmfqt5lVasdXb5Mw2XBSJyBwinIMj8FhT+m3aSxZW5i/mQX+m5TzsWE2Q4Y5p
ydupcrZl7bJdC/D1VaQZ7YCOWnHWK26DENm/q57mv3mmNi0ZuE2Z6WTeIlbQ/4/u
RUUbUpLPvrCMjT5JdwxyytvTsiVWs2t71Fj3zbJxCiPxwjcylVQlqcbYSoJBK1Ly
A72IhLGn44jvVdWflhtx5Qz+zFizgjl6j/7XWerXSwAqiZKrW/Vng+lWW58QYp54
KxRgza4JEd9ktr54OWoJOj55dVvxKzJx29/onlWs2YN8waY4ILMNkwwmFvfWzgo2
+e8SsC/lBL1az1CyGn+80zpiGUhrpzMOOd3NGvl/XxwqIZS5T3JzSRtY6ZgYkUiJ
n8VmvhSo+V6Ao4Tmffg835jTR660sxRytgSGg2YXH42YfYyh++34XqXzGRYbHULM
l/csCWK/C9fKPbywHvjTlXuCyZMWjJiHPzfdgOcLbs0PSSQrz5sNo3IfA7Gk9ali
qdFx112QMuwM5GE1QHE+o5bMGDuHnippwy1GaBPoBRo1P91PWLo23g+Fy7hU9nEc
J782Zf9JzPnynn3iJFA6w1+WeEvdCGptZDZPa03FuhFVYVbfozvZ1ulFjsIxR+f2
65x/+4jTPicaVMwWPizpQsFPwM9+FjFO6cTYG5JajzXrOlbwc5iDBZg/UyAuK7/2
xnSr/fWWiOfGMGIzSW09G1q+7sarKkhgKdvcfQzdC5AVTXdLnTJSKebLqYZuQD6a
+mwFjNIVpRGT6Eh1wtHgJFglH/MWDWM+a8A1/xLcGss7LIWTMXSkQROcSyBqCnZF
KrhKS3mt+/YlTLto6ojQ87MQwbE3aAxQjXLw8rX42aGMtdm+pkPUXH9Vn9ZmS1/v
WuC3renXBPJMQp7ZPiaKi6/IVdxHRSmOimc4LoDXJNZbOcu9MfdNiAxmVLySwkF+
4fh5tAWqssSBsvifpOvd/GA3UtIkCaf8f9g7KzWVX0uIUR93808U6jE3sYMbiWui
xARMIbBiJPdxMqVZvlLXUwzVoI2JNLseQ5QOCpLrXWk5J6iJ28MDuo9o08vr4nwA
ZuzonC8FAJhSu+T+LC3yQErgbFad2Tgrg5GzkPF6V0Wl5BSfeQBXVLIvOFsoQl/o
Gq8/TQXCaTdb2EqNYiO9tyIUjXxAsOmTmFv9jYAiDtRdx7RjG/W6h/0rBzqoOj2r
GpifbY6XM9J1Y4UZ3Mc0DNAIkWslpVv2pofY92/I76TWnKqt9RvAg3Hx7IlE8c5G
gZbPlwSjhn2eie+JuUuXDNyUUT6MrQRhjyygVyFD0Q6DuiZ0Dh39BO4V2r/J9qY/
1AL2CSMqNwzF2tXGJkkaSqyo70xxwvQ72vxvVj7Ff7Lmd0FzQtgkO1wfCXInNLgM
pO3vQSCxaCpE66vNyt+J6GWaoAJJWVPGhSBQUVtOgBLL4j56Gh14liXCsX61yv2v
YPD7ejArj29r7+QVyTJlwMadhBMrnBIFr2zpi5oVTxFhnHXmA5BqZuDmZKrQF1s3
m/qd54/paRRdWyAL9RgGrkyPxo3VATANH5N3JriBtZ1dUxvRWCKXhX69Jz2AedkL
YUWVIvwvb7YqP3DOyoMzfh6tEe9MepcmIGDJemlNjgYho38pOZOGU2n8UCQwhIbx
xcwlHiiulfQMNRMypcHaQ6b2KSRILVEHHouRHQYqIIJYFS19UnewV9PCZXLxw1Tv
iPFdwrAlMllCW4P9qCmepg==
`protect END_PROTECTED
