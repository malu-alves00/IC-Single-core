`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AV7u0NdFWzIz8nUk9qQAZtinDUhKS9AVrYbr5MYH5AaoBdxhoHYQa/92+n5boRPg
CGMSrNEQZ+0kTFgXErSTZf8kphzoYbKEaq65ItfdZfblhselB6HPKdvRoGOao7E2
6rsNBljPOqK6Uwx/xSyE6O605OpKVOWaI/Y5oybzkW8VnJQkbyfzzvSlKsbAw6c+
B/2jHAboni+JhCwlL/XcCUbqCHvxS9DF3Ry7BLz8u6zakMR0sqOPlzrday3KOO+N
7AL/HH6STN0NgMEBtQstgHgDdfesgwooztt8bviCxg3C2hFzhFoWK+dgty6PfgPR
W9YRMHVPWMjnJrxPIHT/gr3B+Lg3App2ayZQA8fgMzs0BTmLV6A5IVxmcRm3x8Dq
GGU19ZxLUYjT1b9qowCgJMMGjQXpm0aUfwrCSs2EWDeRLWpxOFN9WZ3KzyKzXx5h
UydiBq4BU4bP5IjI72/zuMhMpgNu5gyJyNUoUuSmuulhEOvgOAKexP6bnREjWSCc
`protect END_PROTECTED
