`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IaSJSHDl+uh8SAHBboFBTibhEziE2p6d7xIvblsbgtgnv0SPNjZKzuAZtumhbMps
dIGWziWyoTnboTJA1wd/+/9kf38OopdZqETffBZMvSlOI2dwu6vsUKpz1g9CB3c7
XsCa+92RQ1C8zGo4lvWPL0IUnc+EAlQXJ3hL+Bzwe2pHmtbsxhM9wHUrEMuiBt7t
Ots7pu1i1uQwSKV0g4nMgUL1yLfbWePORkENfJWiqmzPJGV4CZOw50henwY4Anc2
Wr6sV7o9srlrG8s45iiv9sFT+tcZLAu5VKQqMap/wJaWnDaZTU1KvTX+AtPPnKGn
FaC12u25YujpItM+z3ENXXa2ziErB7eBh6HFMP87zmmpRb5toMV46i0MZqwd21ZI
1uFSEROojWpUCbH17ffN4F7BgXQmvH1E22wTyawT9xXSVEtxfcHaRYlfgnPmiFgW
i8j5MidkAOnIjNo8I11XaacuThslgK8g8nFPJ761Ha8EVo0ndU9RUrVicoLeeT3d
UnRBrnA87McxTOXbBkj26qvg86coyEve4at/uydZcZdlNqSJnSns94nNXa7yRD4E
KQEwk43iC3aXbGsB/2VYQBRN/6tgmGqXQIdiFpJIBWks7KyFNJHzN8qA933LcbN/
Pb/+woiqmNG0SaGeI93ncXoQYZ8Q2cCGrzRQ/H1tqaY8bjpS62FRMEoIFIBVL4TA
cgn7vmpd5jz4F61ADYqTtWlXfsOxy6lJ+wpkMyjfjhPqUVWFhneZcCzyDSPhpDgS
ySoK2IjuBmA2BGtOA7W6Gdk0cfngLUoUgVKJ3g/rnxCNRC7aIFvUz+czFzn5kH25
Ce7+LabUzNDwbzADTFGq5h5KrRWaN9GfhoEwXKYyokveNQpYxmjvy381e6EbK1LA
VwcSrcyc2A6AkQiWcwQAv/n1d3ZgWMCRd9BbxubJNGgRy8AsXWbAuAB/cKXnseuS
m0br4OatO5qydqegHCkDj4lomdPn+baZbsnJa/yvb/TF117DfDc1UDJrstJ6awUD
hR00DjFecBrMgjLAHh21MKvfd+/mZjv38og7EnrQjmCgrdj1Nbd7NwE7jcHccXLf
HMC6vTHRKx1MQDFr4ofMknjMqm5zeW2H3d83wh5l49bBOuN3SMRq7v5WeP5u57zO
JYJjlHvvZo907Xa/Rzg0xYPpJ33Wa3gUpdQH3nH5LNNq+ymaIo1ULvrfgPoxt17i
0HSgNS9cljsX9cPdmh23N8SHqUeHJl0UYEEAnohRcAN++rSjVcvSLJJZdXXKYNNy
`protect END_PROTECTED
