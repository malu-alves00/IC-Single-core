`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
58Y7Ba+g/FeWGKbDshC+VAXFyXd0kxRd+RQAizesFcjiEW/H1sddFcGqOyPbi1k0
FYZRp2yYRDqLsxJN7HGPkwDiCdf00CRlmiL5oCFn418Bk74BrSTHa21HJwwTO8N9
/E7PFYp3llXa3Js4N7XPGODkwlt5ZXvnTY6asFatvLI9DIVthEstS62AeFxPRLTv
zPrqFn9SEl+XF9MC1SX4eHAiNaGWQJFULOcSyyxd12v5/h33gQyDsTRBvXaxW83h
OxLXt4zEKaSVGaqd22LXucUEZnKlmDsq0ryfnomKPuf5j2cJjSquyWaaONU37a/1
QOOokIeW5hHiY32AovSX2b1fAEkX5wOvvdkb9Uedud3Le9UxX/X8N66Bcty+i2Ny
zcrPkSUAYMoc8hleF/1aXg==
`protect END_PROTECTED
