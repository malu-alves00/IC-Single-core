`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pAEIaxw4PqBjaQ8hLB7G2k85Sc4+UKeuWHRrwLTB5RiG0pR3xNo79BZfYyJLeHvR
PBXtqO2POsIYY45QIf6yFax4pFC8iEeM4QmaUfsaGq5rBfuMKckbtp6WsrT8PXvh
hmr87D9BV3JzamV341ZHuqKzZFA0Y0MB3a7UQvpyEzanprGZqol5Mxy4gW93fbiM
9GmcO7P54LsrHFB3PLzzXmBKD+qB+UkpMdubdFadDhSKHe1Ncy71HrAibEKp7tLg
xHuoc3n8a5KGYxeXxAa9QrLpj+4muZMpREKtg9p/a9D7iFuyfSIUT05G3VMFXPiG
xj8Nae7DvsErHAlGlwqPVc6Nw7vxE6b2qSfdVEPp+MGWnBQGddPZA65qyTvuq8+G
N4qPbmr/9BwYNJo1T4H8/QUjDdawwsxnCSSrV3Y0svfBfhRyfZOiV88nHd1X35xi
CK8UsT85tSKond4pYryT+7adr62BNMLUZN1a7a+6s2clruPSMSmHEI6ADDGstdHM
o0HvvVOn/m7LjJcis5ufh9/G3m6hwMkAgApAzwAMPKUzgVWQFfIcFDfhNdQp6zn7
Ks0Gpr4N/Pbf9b7Onh9DuStvl+rTAr6qY85q0NL9hQ+L4tc/gCtbbkXzlww4xE0O
DXlKXiMlAiMqsd6oFa5CI05mVuAJ0R2+3NFXmOW2B1UZHGpardaeUtvAGLhlsLXv
t+9YwNHIpafShMJZ8BqgxnZz714kgvlGv8TDnkCxdNK78y/o4aylA0JSulusNxym
0XKLUe7zZhsDvN0p5p6XJvkov2UdhOOz7qMJCmSA36KpmWnO0ecy1Cv3gG8oNbkd
hQw7dr6jkGwYf3Br4oL/MLOBeVRRrcuqbypji56IAXjIoJZ8QsQCicWJMCmTZWgu
`protect END_PROTECTED
