`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
44EDWSsDa96dWeoQCWPXuq0aQWbR2L9GujEgmp6LRJWv9jgBq32F+2iDvbWWwAsM
/8CQ/xblw2ZK6wHiYAXz9AyCkfBNa4sMpEYaZU/ma39aOn7EPEgoxodmTLcBo5nH
mbmyH8bLxB2Gnvqr/40UIPcp6PjDROwWPf2netS0pWnSXgEz3Kp5uLBN0J3DMTvO
ItEn568D1ftmchp0DXBmPz2PzBtwgvADMC7CEekR0Ev5gJKWk5udnQRFtRuDRWyz
GuKPGxzKJ/MPr9PFmqDGVTmD1ruQOM3LI+CkI5KlWlxZ4b3tB4O7XPVgcBcVEKih
MysFJBvqhuxzI18tzsXH4pVQS0YkPs5T3AG7JcUvBVrM3tVL4t43wsMcpsKKXjL2
HJNXs5HcMXOcslsBoicTSuI8LctSV/SAfPxtBaZiLSuiMqsSiERd6Aaia/x1NwNy
kHYxtj96aLRzuH4jzNsUH5TWPtN1Dy87r2no3vtRTOFoU0YppiOvu8RC9qQTGsYK
Qh/zfHSdmB77p2KIGyEiLZ45TRX26kWa7KUDCid1r/fEuixEON5i5HcUduVnEr1d
4rSFhfso43pJLBh4NZqFbICvBtaGAqA6sbtX1hj8H3q4C29EpN3Y5KQka/vvLz8J
YTQLr+VMiuG2ZD7N7zb5su2SEcka1Yx7ALTv8Zgdmb372NqtxpRYAj+5JK6i4BDr
qE8hjH7qA5HnpKb7595NusTexVs7tHTa8m/w8jiysa19/M4HGep8HcpZkgPjWfRJ
o3uTYgA2vLzQ/BdOjkG2FkhpWNQ7SZdjU8WZczIGraakr2mE6YefTrYhHpNDmr5i
7j4o0oh3yV2Frpsg6QjlaucS/IEiIhPmVJlnj37VUCyEDEdaqfdtWUYpLYfkFXMS
WLAbs9trnK2Mup74xc7dovkkGwRS0qavbnd/A1CeMbW7sPxSjU4BHBbXaYxt7x8E
5HQwDug3+D4/klzQSg7+oK/Lb0o7BhhHphmvniUBK4pTzp8/Sq56o1H9xB+AVYDY
DsvfYVcXtlXeVJ4qRW8rLD1f3JyuY3yESspeTDrO1NC90UeZUfYBCJCHj+y2u/IL
j1BvUsp8mv0MgHK/lIVySfWuKSXixb4ysYJM5KIMGjzS6lkzRvn7UduDeB+rmlf4
Vxv9FtOlQF4ykaZzKhf5eyniaO96HdxQsiQnl1LPZQOQSl57NAQU7z4pa6ukDH2w
OMDJj5GKfbdQJ2J7dRPT/HkZV7BQ3oJf3/+thbONzOpG3+hc9C4cJkbQk6tP5+GQ
7P9Ny3SCw0Lf9ns8TB8kl2YURVBL5/Fa/UneQVrCsD3BRZOAfBRNnSl4CfwSc81B
D54oxnBiOVJzOt229lgnt/f/aIyhtvrYm1WpxzxPc7tI47kGTrUZ74Eu+h3R6S9s
0QLsKC81QOV6iTIh+bt8mV2/KJxDA63rKBjhLxNiThIkdeGl0s1KzJ5AYWrqA2Sz
FCC2ULGugmo2EFbRhI0DoO2alRyfpmvSvSETAHc0oVt/e9qrhrQVB9TgHIxLzh2S
GXp9Nc41AsPdJbFijO70nOgM4LqRSr81CiN2/tHohQ+mTczjecXVEQTKPGHQdnlX
ix5WRxzLVb9G1I7wAgbZ1scsym9+XRtSQGpbHRuPtjBI3IA8mrqR1QqDS+75ELaj
NGAWF/slqACeaIvJ3D3gg7FILnh7Ua+pgN/+Lc9jj81egZnxSSnnwYfsvNfMGRvI
90L5X/d89Mg0Cw0z0AOPkl2b2B5RwWBapanRrXdtvW1YewjUyDkXGYKTEDEg3X2N
fDHi/ahfy+SyM7SHhmpWUYme9QiT3LLaJfKsRd74aois0UQn9rZEuu9KznBUaefL
KB7lYFU+N6O1X5rfYei7efFNDsPchwWarb5qEXd6vdgQZ5/1Y4EgSRU9L7CeChNo
Ck+F4AW5LKHkLtUfuA6mARPq7hdRBa5U2VAyuX0ZVJYssuTauSzRhfb8gGhWnUda
33KvE56kBOdlVqGROjYcbhAZEPYJnbZTsZLSDjcpNRXF2VZBzaIooIBOZ4RTtC8f
wMPZXePiFlk1WkkRWjSN5DFQd5ORImtwYa60HfYhatZnsgiHcxg22YFhi/L6+TAs
h6GOKGuhezknSOUsxs7hFs1Twb5DdhBuln3pauSn3RQvc9qLiarCk+MmdcCxWjxd
uyXL2dAH9cvtPQcdjy0jhdD1FrggxHXkfpqSxxrdT9OgO5NhFSUbBOhv15AkpV56
o8s19CNTGQVeP3QcfXdUsoKoImq7tmeEVH6hVCUhJ2joPAAtccj/sF7cR8oVyNbU
YKPSe9ihZK/+QOM5GvuxVWTy/Cib5uMvB4ECX39s89Vfj6/lbdmaFNnSStBY3lDj
5FsXwmIF7SSo8aPFYIbD9Yuy5ioX1+czr3U46MY6/vpi+nEJe3p+4qYPeplEvxkC
tMtMvo38QzkaTbjLBlfdJA/ucSRgOlthIUL6V13l8DnwYpsCAu0DNZcMoGVH4Ack
YVdTOitfXBYfgRX4Woot7i/W8RLMYE3mF+PP8FTcGDegKS1+nJc1RQ+HpZkeoJVI
H1nPFgbQsGVwtreSyKhtudtQCKb21igdWc5Fz+UJM+/d5YjSLP10x0ihZbjTXrlD
AGuNx9xAPWUzwebwHnXSjqqQkRLyGMJzR+mgmpIaALJYGMuueUkmvwj64FrrmxS/
1ADnslMDKCGl5B/6oBEv87dWkzxBzuXJM1CY41kL1AWXetAuJvJiclTSN0ZH20ig
SC2RXux6UJmS1V3dpqio7sYuOSELp/zCnoRBglDEG+mnR74LWv6VvWlapJeagvuY
Q6Otm9fsV+5zYDJhKFy56lAXx8Iga2vhqe4raN+us6l4A08Agvoy1cBD88m2EFUe
4RknFh5crafUm35eF+2AhvcwIhQeVIURs9vRuKAVa8cDcBcTqyInbRY3C/GBjK3t
H1L8qMlUgKbJHp3x+A+7haHQK/5QpHrfCzNR6+2vbvwF2RJd0zSR9UgMGy6UynR4
KOclN9kWBj0uAs5RfzUyT1WbaQqeErhD8xEo8Pyyk71AlaqKSqqPVe+nLNw+0y5p
QrpFvWPxJ7Qmf3gQw4eDmwmZPAwVU2qhVdBioSNPyOAzoYvb6DIVGoKYv5Q+Z8l+
6SRpBSqs4ZzMY1ZsoIm4qZtoE2+TIR7zJenXnU44P2ENGlqItsxjCZy3ujehxGXi
b36ZyHn/vK37x2eITCQ6NnF+H1xrLn2B7YC2Yt1vRYp0hPG25rW3P1OaS5jsM8bq
mBKDqgLr/NgpDE6Cb+I7dvSzK87ppJIGFgQbHjt+dvkWh+ISeSkEL0LvYItBzEE6
TLOO1nXkEMb6pLE8aRfkq8WalWh/gLQXHr0g5zTA+DwqpZAQH0SRcXneuda6jf//
/y0f2R+r7n/CuBVgs3HjoZihuEyVPgwef2h3s6lxHyoBzWpRyP1oW0qfSBH+6eB5
XB/wF5pD2Fr0nmKpoBPhXAarCRPbh1Z7owgBqHpvsz3wcd4XaEDFA9Y9GhzSS1bi
eIdXy68dSQYE7MkRrRjgHdSkIhGgeIYWs8rD0H5hGAO3Xfmd8l7bspbkwvS8h2EE
xl7MZj/D83pghw/1w//aMj9+HpxRdx3flbIacOPTMKkQiXiOIJFsqAPeP1of8Pyg
rnTmCqcFiiOjd82WP7ODV5ku8+KkpkCvGlexBN9FQwZCZjMJc3L2MtWqipGm3onC
J0vEF2Y3hi3pcEag7Ke9+4H0kb9Ye31hBi6kpiT9gXjRDHKviPGNa6NM0HRannSF
ihdBjwp+l9uxN+LuLvixfhtfe7wWWePCf94SRyKEH9VKOTBKNc4fJjBQCDdXVHB2
4Sv1I83yxWbVP3LHkVLvc8CX8DeS8u58aq1emQHLLun02iIwUaFLXvunfupkE55d
8MbwGCjCZ1lYrLQyfedwA/JWmIbEq9Nvd+9wDhEJV5psMCzw96vaubnqp7qHgqua
UfSaqgus6wjk5KCcwkmehAaL6Wg0cP0ipnIg15biwUgBHCmV+vdlFj/9yLNi1WR6
C26rtiu1c0aqUv45W/0FZBNxsSBNc/wNoFvxbqRYgw193gRzJieL48VPnItDAFhm
3rZcrz6g78husXJ2rDZbwF6IFG9Ziodd6Rg6wcEQ3qBDF/R8Q3SX6vqM12An5IgB
g8fbfbWsT4Oayu3BHtdYxgNBok8bYzdpsIoV7N+gQYqYrqCD7B/eMhrfH37yBoOc
Ss9vxD160f9Nxrl6B4J34tbdU2+yd1ftWogKHKqY4pOomB82GM2/VmiJFfL/hMoC
UReROl9SUldgI2GS4MjS3cuf0PEBrOZKi78fmBIAuhcouQJA0PM3VgyWOoDmB1TB
mBmRtCBNih12nRoODXFBKBxdi0m0/ER0DKggGsyt5HdHjTwAO9D099u8WRUvpS7v
Zty6PDORYgGPU+g+MtU4okY8lh5WpodHbNAf5gPIQ7jMwr/2VRCF08PCEuN4dGsZ
5UyS/lhdVydjfohU4yARG1H33AlRhOQzz2fiZe7bnlxbGIMbPwecZPZU0xIl/6iW
FEJ89mhTJK+xQGtgpAPBBsyZt0y+BpJ03euELMR9OBw5WEpu/LKmRmoFN3Q/LfFW
z4//ww508P0fMU18kxIDSeehRjRgUESrprp0XqbT17rcAVkStAp3bfItaJ7MzG4I
6Y9MFtwopySaF40S/cfDtaoZWhI7cO1FFAo5Vr3z7amlT2Q4+Nr1XyyfkF1aZhQI
nKLyD6KqB8brrV+V0XLsMrCgFHEGffR6EiVeuFWAQktAW2ndYrXk7rhvsV3a/bUM
b5fPNfUHDJW4OaYP5ibKwoAXqCveOTw8YCbxavIAv2upZIQj6Bvv2FiMtjCqhF8I
B3IkJ/rn4A0And2CDzVT01wusd/jaq/URetmQqo6ZipQM+G86OubNweLIpcY2H2c
ZDZUTV6qYjjlio4SCwob3OVlCg3utRHqzZV6n9hroxMskuo7JHjFo9Ehi8r0onlK
B9Vhi0zA86vdpVYImy/R1W5VncWkqu6OF650iijNV9Uk4P3BbJ4mDb/oNQDkJ40g
LzkZdJb6NAsbdM9HdnvgfpNjZxyNq/5Fhd2bdoTGGa0udxBBamKMj2I9IH+mBJAv
xIveI/xFvryaH/jzCY//mksHHOrlq8fMO0ulrhikUi6NCdPcL1JOKRjtEqknaqBv
1Xur4K/NJXOpdrtkW3FamU7dszxXWH0WXXGWShZExD091odYtcueezWBhRcD4ty1
8L4k4OubzdU6yRja0mR5Hcl3AV321x2DjNmsQnMGSc9tfPVawiQwQGorEuGTtArt
VwuLh/LnfEMFqjO5hAfudk0ALbcQgcGL4lKDFJlQ46VhFe7zZYPGFRW1LKxUEZkK
5q++ONOFl+2Z+BCFCrV4PAKALjvtDBi1nDiHvQX+c3ec9EmRwR/3cch/DllXjy0u
/pXHmDLNXQwmMwff8/Vaia6dRmQ9PFM9RYoL+uklquQ+qa1Dwpnxkcd+NY9pDWEV
mVvknzBSO7KClZ9stIELm1bcNzeyyutufLAsvccWpiuyci8wImdrmPkyl3HqsQOK
Hn1hHYx6Z34Wq3WYA/7t/5XgFFsQcpwlG6TICOUz+7hb7Lo9NuxmorL9JhiOOo4A
967JKLt6474/aI7y8n8YJpoF2Y8Zvt3TNaCJWNBn4MtmQg2B38diRJP5QJEaWNT4
FHa4OJUZ2y7CFofTDHMnc4Zff8e0LN1MFHXyBdA2HJHrMM9QgeRPQRC1lkBhaWp0
rGg4lqCwCmjLpT5jY7Z7Vf3czkteGq5EPOtlmwbhrG3EruVgrS2k9cyrbZp6kbb8
dQNudE01GSLo6xx5SZpaU5O9fIfMPGSLvF/pPMDEE0HxDGIZD7i0WQZ2aptaKrLT
f2bS7uiDTNdBq+mBJXHF9hYcftZX1sPxD7IY/xCfWL7P7ERh8wj+TZE7SOfwE1qm
N/inEARK+dJbAqcLjJ523BP8U1tPanw3M6gRoAcXYgDJcJcSXLFZhPNBK26uG8ES
mLbMhDO/q1/k0y+lbiAqrteCgyPFttOIcL4VbHH2/3QYJL1UO7zf12/HqfrADyNH
l/NRoq3k0J/Tt+Xp/UDDZHMuRezFduYXofdxPXwCBXU8vISTvJ/afcYqlEDKLtB7
H1R1TNJrmd/nFg9pZMdBtJWldXqrTxndQgih3HbR6fvUV9H7WrsEMwebbJo4GlRb
0hHUvmqHd3ujs0IZvHcJJl0qh1GbeGe8s38DvJWuGebOKbMfVPMWZ4anmfBCAd5C
nvOTEra+XOftDIIcoknEd+fo9FKvA2rj5VNPyJZYYq8urvx/ht8XluUcEuuzPMkB
hGP7yMFlrpoRsrDvDUn7cBYXgTk7MBAvD0v14LP9qcBehUitnkd0pOOI3MRiIwKC
UTI3Xs4qeSwcyp2HrU6XKE9NQdc8xItsJlmsssSuU2dj1L8pdtbIMKsD5rgvrA8V
V2+MFdMqp39kIABvVmaRK6QUS7G6uVitSsGb73fwVHyX8xyP9LaIPQNCvtHdtrHk
NJqsaipKwTivwJs/Gh3ua0vxkciTSRbgye7a+5gVsXXJoBu+t8GI+miAcnopYqKx
w1Z2WNGTxPksfBXzlfoDSeYwvg2usDwDbDGSnjS38/DUG19JSV7KSl1zLnFDYbgS
OXTAq1gtuWExtJJmwW/EvEDWxPkyIwyG1RKQDiuKgP8C80VgL4Eg2MpQcaukD3zZ
04F8nUzwo+8Cry9jqUF+q1P8JfP0lwFt9Wnzm9O6vqVJ3MElKAWFUK4LxGa2kFQ5
PlMsFUUh/ohZD+j7qHOpgIqF2dEaGQ1yI63AgTDls0YLkq2px8cr/+480DgSs9VY
nYoqGS/tJP/1O6r4OMAWbUKS9I6pKNnDAK+rkx2mPdz9SH2FVFloOrmzXVHwZqFF
bd0JA7F7rF+D30fDH22p+AUYvbpOIf219Esym5jvOWxp8W+JKxd++Zvabq8aVDye
/UlPOk5blOhkMndq6F0HqCy+FGeakIOutz8T0YIi0XBxzv+gOC+cs7999asss8m8
isa7iL+5KZ2HTJGYg//Hbdkb3a0GWvaXW+xiSoA0rUZRIYLJXTWMa9ONcEadhpS5
n2hP1ZkjLcX1KyJZCJzIKlYvz98hOvzjSTrBPiUKgnC8EiIs9H9VDKD/4XaxJGfI
amzpdDUSiN2NlCuilZ9OSHPDPGZLvVSicOLEaAwn/rQf13JTWi6tbatgY8eNXjVY
g7+C4M5BOq0m1qzTI2AYxquGgK+jgEEYrTstDva3R/4DwTd3YWUPj7WapR0KK5jT
9Ru9AtW5EAZPE8dRZYn+TXt2AYFjgHrQ1+kgLRgqY3sY8brwQkK3yIlsUi86dRSb
1zvgVToqtTErFqyUY682eoo4HjLNSSb6vnZIHoWNxnf1k3xofcXRp1bBcNFQ2Obb
NmkdSMWNI6HYPR42UBboH/hWmoDpVbGUcPjKCcMP4emLlvPCS17YKNpa4p/69MWj
WgQdI0emUmbedoQwzfBai+kKuHYrSzy9vo1Ze7Y65ECF5HmGIjihMnu01BTzdkv5
L2ZgZp4q4qomuJYglIz9cuvOTA2Dy2t8yoOG7w8FOmZ8NGZq4QhyvBJqkVtNHUjD
i7l9gsTS5mp4YEVsK2fVyr6DepB/eIQ8iexZax6xKtHttWijbxfH62+CBYK6mRoA
OFoOQSbI4rQWLM0f3/5QFI8CClTAPBs5lZZS9Wd8W/g5v5EwRbvzS8ZqzUwO67Ox
SsRJkvYMhxI7SbOIQqnl9ARHYW0szcrnKWcBqAUEPqQP0F5TPyZrIhmBj7MnPJlD
wyaVGNQcu4jGK0bOjPmwSmYZ9lqDCjcGjGZYfO2IZNOJ/dvcVf7caf4lstmG3+jw
5xaI+LHss91r+VxgSVu6Zs4rbkTZz77aQDvDVYGNlpbPTy3uKKSJOuEwYuQmF+JZ
7Wxyh9wc+54Dm8FrWT5DTzggJcaDqZytX2s/xFMHeBmMohAjZArGJ++Yj+37n15f
blrSiQQAbZrxAvszZ2/HzUTR5snBxYVP0lOq9vISgjGf+y/kM+9or2nhx+jReHiO
ETPot4gJIbVYgVcdqWTb0JjQOv61FlXftwLLDoEQdH8l8pOreuQPB2j731z2GnVd
NAcnRw7MRZpb/W6u/y3rpxqvCNIzCzsyWFcaRp4bW5LKwBzVhpjygwrUV+ErynIa
BWj3KJ+u6KimD5/TP2jh4JE8JqsFFHySHdEXlzkl7HAtypcpGNU29w+Kjwd9wE9R
T6j9vNGHJHGjWxZ/v5IR8J5j3o9JUYvTBLPgB9zBwgyyBcrzwSGSXZ/LcppmIv+O
V6ISJUKmeiU3VHJUjTPDQeJcbhdvmL7xpm+KxB39X6vieHpC44epWbGLH+TK4oAi
06szVpCK3IFKJ1ubJf7lZ8r1u1eK6Y26cYFi7E9xv0TulyQaJsRZxSBOabV9Dh6S
1q+i8jtlsFXwy12IylW6dkHExWYvgZuMpYjL2/1Z0+QCzl2w28YwRww8lyh5H5uL
Xs9JK9tKBLHMjA4nbj2argH1cSrLS6LfC7MWr8F9aiNsaPfrCE3PLEHlqCzLxzDE
wb5nC5N2kEiS9vAV6POP5FZJfzvuKs2tJOLA+F66gckvlBgKxevuMb2PcxOtFPwQ
cR2R+47J6fS3bOSaOCJ4ZoTwZcfTpk5vO9yCw0mSJXowRGNu1Tnj4xs2LZeDsZIE
X8TSVHJj7zPrWb6hJ8odOjwutiqwYVoz6h8suspJFMh+DNAM9VyOX0MjFJMWc9AB
iKv++zCgOpNNNpt4/xzbJBTbcHU30Hgrf2l4xpTLI0reRlXW5w0cZwdFWVtzZVIS
nkD0PaEBvsBaiZjuQxHLFQ/4F3+ROqLsYjIxQIaUtI+JlrL3XF6DVrCV6BHOvB41
vPGsspXr5nxk8FiyLvKhQmToYkTefwtVo68j38+7F2sNjoQFS08bbFdse1FpxqCx
/Neh9mKkQVu+uukc9Ff3ewU00z5hEmEn553dHv18cOgVX8uESYfTRypjLSvR0189
wDXtYtDGARRnbxiRwd9bKUPQUNOcLAgd+4tfYEZp73g7K/J/rAPPEpWgPyJ9PmKz
YAV/22OIxNgHRrGkHTerY38hhB20uq3/W7+C5jS9T7i+8CMAxweO1Y1IV2WIFs/h
FdM03QY4u4W2K/bHdZ98ObxXssDsLw7Rwxw2LjVPQjQJiMF/N1AJOFpaAZEAJpiW
PGlXHtWxbXzSkZLTC9mJlSCGe/HFtRGwGRHCkyjrleE/3hOmMFElzV96Cb0zfMOz
QGXiuX80HEdKtIAf/PMwbWGqiYqsnwjOGMTh24D+rr5UM7iCNwUt0IBo4PUJCHko
FCnTH72BWrQgB0kTlTBswRtGAhG1tVYPkmSdFtg3ZCBPVcK3/mKXnsyFaLP/ncMb
I9yMKOWlhYvaoIFJPjoyMlKFUVjSMuKUBfcUFg7MEFP5HotNIutTl/CvOATmJn9H
8G2f7jZiAoiRJEjFXztzkCa6V5mGaJ7d6qWsuE9SwBdixOMp4TVbpljh6Mo8eMhE
TORmG+htQoCnn4mf9iMp3HHPXIr5QUSdVN1bf8fP6I1PDgZKPQeeyGRvOKsuKjx3
vwY/ZduCGxU561Mi3Ew/QvjI8Vypsj6B0GjH+q/TtlSvvFtEaKPCIMP6CftzaI1/
ZhvVYQncwkTMmJO1v2REt54srCoDDvUCVIjpXXQlIbeMnKokDxX/ABtyWdVdJd4v
hzQxZJFFSddYEUgO2DIyHnb6f1+AUMdVob++G+ifslt+ijHM1g5l44XKDp5S5Z5P
qsmGbPPu4d6vdLSnvh+hMsc7ZAzlIM0szo5GIu7c4Yw5Q4vIJCBXNxDRwlYvd5GO
S1u1bHMA56RAMJ8NxlYax+vohz8zHXeNZcrXCSOjOnmOtcAGDgsGZVstsjyY/aLf
DiRF8un3P7pPwUWvn2lzE/d9wESSMikvV6zMqATldOPqCVNTZhufQbgcWDXGBWza
LeGhrFJFHV/nB83yoD4x0rK6bIWGPIWuToUrKbFwXa3sg/YChtB5AIEI+LBT5M0Z
/6DPJnIE9G6fMQ4/qXNNqJBDuIrQ7tR//qMFuWYcsiDGO/ROx4E1XczlrRy4AywZ
hxN+EWRn9JtwafuNy/MGsAJ970KdCjWsJCxnGYAMNVqZjVKA8j5b+oOyTlyWI0h6
lSTOwc0dUC3J4CGxCRA5MWdDVhKG42hkTzAw9drSt8B28erIK0/acUobxF9sXd15
KsVoZnVdPJD4KGdPEWNYAZW/3aDbFCIXKjtT0B0FP9HYb3qcz23k1TxhGyLWYgt+
oHxq0G87jXzi2ydMpZSilFg6TgePIlTg8qLIj1EHBM7OIgVniQzbn4NimfS8mQmh
qY3Z6dtx3m0OBTzc54L6ugk/nwY7SGJ95LbIg7JXnRfFh+TXJ2w3Gfq1p0ZiCWFo
vHqGl0Z7lYsSVFN05DoWoZiAvBSyCY6yteAYzVCkAhNmUJcrdP5a+lBs9FxwuOoZ
cGzXAlsBtAQjMf7d0uxyVw/FSx1ZVMLgG0BcZzFFEldQFti1O6sDnN83L2lPh+Dx
wSgAyRMumLkeue8mcql9VP1KW02o9bDkcgt5d5WoLIB4ITZOORC/8sZxXK9HC49b
BUGo12im07XAnsQmzRIXIklaLtdCzqqeeI55zLCC7RChXubvPbU5U9FSKyDSxgv8
6IpVJztvmcIlh4aaAF+z/J8LuXPZVWoQR/Gpm7wRcboBsUbSHo++MGVQuYK+Dj/h
ksReiec25k4IHVfkI33s+5/Qyag+6scFiYzj/nQiUm/rJxDtpZNtVrvP+3ZToOxq
du+T+ehb9e7g9+ji6Ox6qefDt1J7Dy5hsGMT7El/Cv69Orun3TTiqqkH7mGS7Q5t
cyq7KDYYAuz3mOwQkSmh5wJvEQdghh5Sn6n+sCT0m1v+Oi5jSMvZM4kBBoc2ADA7
+V3HBBfihfPj7/sjklV0Mi/fmJn/CDMT9QpWGeYWBaYuVhBBJigEzvV8mS6igJz8
ea3icPpWVc4jDeCsRBGQFiLwKnbBk1OIm2fDteiEc5Qrn/snpde2x9q6GesKi7Ph
9RBIXgxSaJOmOEYEf1XVwbU8ZlvnuUnhEpz2N+ZmhV6qtbOjbDhK5mG3HflWYpcl
Wk9yxB2cyczAcnSwk/jlp5wnNYyMeGJ2a/TO7oWeAz1DoywJBvKaN0J7W56uHBtH
AZ6jU6R1rTg7HCCmlu2XcxR1eIAzdK2y3J83Bk3TN5wx4Rn+i4pBfBtwz07zkmVz
JxT5UCieeODkF89C1YDK1bx4T4iVTnBHIlS+9s5goYqdVm/kDFryKQzMMSko4wZR
gNVlRwuJghjF0JJfA5gH8O6uAADihISgvkGGVBykW5R4MYbvarXK4/be0lXHUFrX
AenqHH+tygeapNk9fE5moEoocvB/nxvTS0O3ozCovF8mN7ux/W/ZTJiKHmf6uIVT
cB1Ii0/WT4Ns7iYm0kvG+M7QV1naT4yGteZPvjLTri+9v7KLJ+fsrOQxkZ3447kV
PafylXv1G59YLRGU9t4l2xXdqId8s1WG+ET5um5DyWx/9ANZWB69PCIYptdwzIkD
5mXbCKQChc41tal8gmP1RMW4LjyETwIv1Nm7QjlSQdZI9PgYDCYTxTHt34tCOwIH
pK3/ViwQz3jz3RjTbpycZBV5eN+Pc7PLDbdRVpE2sRnpP+AgVzVeX9tJxjlgxCUa
8eKL3vEqkA0JbIyoa912ZlWOlDf6GuyHNaLlju3ermIEpXJJoqKNXFKxKcf38DhR
lNFFMuF79ONt+hUI3Q5d0WBLTHzHWp1WoyE2/aJUqFfXzE3eiTJ1miqzY8cnu0Z+
06m75zbD73U6+4roKR8DvH+IgwFr3AhjgT6LwhkMAIqBZmo+7/iGb+2AIqTZpNps
cYREEY24tHjn5tBOopeMdeb9uEw/1KkZMd8RAOV4Aguqr5H21KK2+IFXvGna2cuv
AZ4ap2Io+2+IgaWH4O4b7DQDtFO/7yD43dWvgHHP+uJ5XQV+0iM+4GZc1Re7oeAQ
+wvJstC0hFAAPuND0ulL2feiLU+J1P2uavwIl6jp3Pjv4cx7wM2SuFWSURsRfiAn
u3ufj0Lcy4bzCZ3AbSMgp4tF8CFkqKqlkF2FFa4dbt2qcgpNS1+QK8BR7Eau45qI
ZKTU7rBwN6VOfKOdROSsxZI4EzLyLSGMic4vqcBGEjKVwxHUQge+gPdXrCrL1j45
3tynBmvYPqDERfkyR/x4Xy0V3tbVPlTlLXOuRXhGzplxOliD+DDMAcTUfxshy+LN
blmFjCAMvsLQaU33V6K+/lugEoXncNRrH1m5PAt6b5GhhfG3w5Auo+huCyYdiAn6
d6i1WD+tGQCVLEiCH6Hazk+Wieo6ib/VhKizbUrNMa7icm2F9t40iyZl5cNG0Yqm
0OO2QhtwGaM+/L27rHzHTLSeiFa2/hBt7b2U1/cuzRRze283F6S/2ZiIGZLOAHrz
cX5m1olAPgAwZQxSnMXW0SYlssLVoNXX1ZO6Y8T0MsEWM5Rg7slGKMATUgTGdywC
anrghs5gOWpKM3+IeXdhP2XMlsd/ycVgAF+MKaqjP5KmEcpJZkEVzbeTdY1AjDby
cT5tPp34Xc6hygdBlpOAuJ2H07Zh+sZYFIfBgALb2fwOpSZSzi2m3QNaUCDiF+0f
eWsYNsQigQtnF3tiaQYkoB+DMYcxNJjoAsE0fmujfhOVd9EKCIz69HuFXMwMsTAM
Tmu7Z+DzrLn6WntxeJ/PmgAC0xRQOzXTUbRSQig0W+q+GncWpRjpGZt/pbdNwJRQ
jtYYNFcM6j6hSju1Wr7r6LCEJiA1xzWKUKUYxHzJzRmGIbB+EBG19go1alJuhvBO
4kttg7uigEwiSzEKRX1NYhXtvXsCaawqW1bUxgjAl16YsD0fc2owAj6a7WV8ZBBV
HRAnLJEEUVgUAlSVAy5BQ5O7w4XhiP30l4qd6K3r/rl7q7izPliNI6VGQPwUIFnf
qaGh/9vKq4vFYSlUBX/u9+EXyMNs2PyvCIrTajtvPwQpMFOBkKEE8a7BXiwuEzow
VIHgGS2vzf718eF0+Y2GULGM6qjsM/t2r0LC1olhhxZzEaDSVMXzsb5AhHZu8JZJ
VdPjlc5+DEGi5vipim9Fu7W501PkLjuF0l/ySPJ3QKhjsNtBhmp4AFMqC43Y6jAZ
MWYgHOn1uoYuxAuGQ7GQt9LgabocKidgRDHCs7I32qk=
`protect END_PROTECTED
