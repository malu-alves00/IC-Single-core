`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TCcbV6qlmfLkyQXohNl/o3WwbMNJyw2AerZaxAzvQI1zxne726lB59vokT6aBi8u
58KA4PuaMwaTZaC/JqV0bplKNgx01OGuoqrkanIoF2eripOHEJP9teTLEZ3vtSeh
6+/uk3AuoAKkHXjKu9JL41ZKWPmovAmimZzdzixYl53JShRUyuFSPFbeI2ecGomu
2+5ER2ZKa2F1Z+8S+feT+jB0/UjvMMhOFIn72RyvqH6eL4z0RFpyGdy7YdTlzhTQ
vR/W66r6Ud88JuK8qssquoAQ18m80XuJtQYWDRcT1cIQ+bqGY80YyoCcEdFoUqsq
mAibZFA160Z2NBFYQHv9oFWdaa40K8MknYYzp0Se4ol1ZGv84NWwy236msz5qImk
63XM/GDKj0ACDQwU7hWWj7CYf7QkyzEaBNk/fyia5kB6t4GWKGDzDpO+dE98C7js
uqh6TqR5Pyb1MtwHP0qqoNPBw/oqU9HMR5zWjrBdR7xsmI39+SFfritRtPneUYb0
lyTWw7C6dPIs67HCNrMF1fSnuRNfnm6T2AwdHVLNLCwaPz9UP5qype74Ff/8CncG
rZN8OIVC8iD07v3aPlTl8AuLIrpVNwbjLun49svsipgjsRAoLc1maqMhXS2ZW9QA
+tDSguT1LuzvYhVXy8W+F8N0b904axqXhkJr/Hzt7bAwGuOI3Pwq3M/DD/thZ0y+
wF5tW7wheN1hhXOzVC2RZZNTkRzQSeWH0b19hBKUMFx8OEgsgkPSZ9oosytL0NbP
UIyZAlA6Nqm7Kje+36f2P4YV3urY6GrRiADB9qKCbVSh7sgg5nipGFOChIjJIfVD
9znBWY/iTk002KJx/ityLp9rB3yaPXnqssLRGNMTBq995FhIdYmFouLDjNa+7vsu
63JEtx0aW6rnk7L0L9LUaLD6mySj/x2RxM0jt6BGNKgTltCu5rUrzEUJ6faMtgkW
Lp5v2b753WGefK6uP8LPurECig2rrJaZo0IDcf1Ad3P98Hn8vS3yV9VCrRhdSNlf
hFWEas4HqpSncXElsKgMEPVbccWpMV7PxIuDL4bUjaLhF3NknkgXv9F+ZfkwufAF
Abj/g2gWQA9inu/6ITCHWkni1qvn1JheGojn0xGPnNFU/OHfmhJJtUfC3oQrOa32
7zYa7PFuVHTfZ0/p61LpTUXfhvgWZc8xGZYmjvZJesGJo1glB3spiTN/z3wyRPwg
CsJXUa1YABKISb+ecokXX6PkOHWXxl/cFy/fZwX43PU2qemwXEjrg7/TQ3kU5iOE
vfkwEFhWJ5aUyPVx7EcPJy1VLTBZYQScELojA8dtIyiTF31DxJ4YLaPvGeXjrxf8
NHHuJSYpH1AdQrmvJxOsVj7LPIAx1V3k1OAUFRdGH7s7WKuoc7EsmYKy1HS/sbcK
XteYGoiSszMtpvC3kuyvkuZsYAHFEGuJMTsYX6rv3pJQ1SoTRJkPMr/b+0Rv163H
8x+of6V7+4lQxCCYiGBPq5NcR8nAB9aVUI5fgvN3v46gTI5nsm1Op6XZohETtAFp
ZqKSoaOkm88ou11ch2KYlCwTeESgOhtwNebYYwVsEDTB6VCRB/TL2AdglnSbmcvM
+smliArKfpeI7qfMm/u9c+R2rvQgq4PrY8CkVyCoEibgPXYOIi04Q7k/sJ1SEwne
RdqhO+esNjurD2tCo71uXHbcDVSIjrkj/c518LEkChBvmTMLJh5dNf5pcQogYpcK
IrIgS/5VQaMB+NfWm6d5ewiNCh7iBqVHQ38BCufy05eRp9Q1OZMd8s8utg/cIJo7
0gb7eRm+EXf1+SOZShCD3fzm+LNsdk5hEpLSD7x4Omx6MS8Z8qOr/bWDnXtTRk2f
L0Dbv+sCdBxDi7Fs4znz/2fedWfX6aJbxIkwSp13BoTZC3w5nWlXGot6ZYXELtWW
rSWXzgqCVC+VupKh7bqdNzvSYpI3NMj6vWzXKp8j4hF0ThfPxJCcVQJtCTpMaSUe
cQhIQfDcEIaHDz3tKvszF2urpEHaHTLHDwc4+tSLDyaGF9VXYLFMYZTp5UaQEjiR
uUb+4TYhg7iNqeRQUbIzK5QBqHSZpncGQDfQ6vTa5dRmcGkdlaTnp0H0RXT1yrJ4
k7iBU0u+uqyJtESormzVKV62wNKShpGDjBnHVphjh3EC2/Ej5KW0DlX2vWuafXxW
cLQxp2503ewk5BRV5TpktzHnLzpyBx60fgTLG6QozQ2vR6Iitc3MwE78ktz4Erdx
QOYljEW8pNgLIYMOcJk+UPB+OdFCy1HRbqIhqVBAZJ00LeFeI1XhWZ0WaTXkaM7d
QrxzsO2xyMXMZA6TCqT9wAOeXH36Sbc0fqglzIv1Cr7H33JJQOKbFJpN0f+kCbtH
jAmC9EJ6kyjKw4oi5rowMvvBNQUJXWhfOgQJ/XuntAe2YNNEggIa1b44rjH0kRZg
vskDxVj51/A8s3pBShmEJ9T/GUA7k34JgscNu6Rq1y/AfGmT69f4J8dkSzHjNzh0
869ar6Jdt+sK8az0GeWTt/Iht12Q4/pFtGuAa4vcPBFtLLjtobsZ1joGdy/Fsz64
Iy0/8fPvxK87joqQtf/6WBiLsjKNaRmarqdV1u9s0sMU64JTBoQe6RaF6p5bHgPa
sgw975Skk21xrbf+8nucmIh8PFfyEv5R6dFJmzE+ndPdy2naa7xTN0o3uiHY10hy
NHsRCyetRYCCYEUVYlMAxqqcGCvGuVYOMuqu6GqpGzEMuhFb5ALYW94Lucnwq+/y
WlV4Y3z9ImwrSRq+Nrnw/KP+bADsS34Y74Ap9Wifl0ZyF0Yewf4vpLalgEcv3T3Q
5lybqoDdPAg+xGOmkj8772zMGOUEGBQSLDIpzJwS5F1MJvbkl0IszCKTZb7bCBIn
ImTDgDrObh27ZeIZWnHuEAQju7p9YobPgBTY74vATn9zqCENovLfDUGAWpvmo3I1
wdLzr+jNss31wkndWXkch0kXpq4ltQynyMCvr1prx/p1djolOYqFY2tv7BLHyqAs
3ejg6hJnTB0qKckxuVttkwQX+CnqPiM3yv2oVJxQ3ZtvSadygBme7rxBpKMy1Rf5
+Vj379hH2hv4lGQAYOQSQLrTfBRPq24ymhgPrJY7lk5p5oy44I/2FUUCG2iYLgvD
/naPKEWav4ri/jGadJtrFfPQ8YOvGwBQ9vdsDwJIfKIlPYcKbO4mLDA+sOe7moJM
aIXHAgEE7bLJpQzsaFd/VOqWYQvBX9Nb/5YkcSFQnbUkBCDHAFreOH0KDrWqnAsn
6yiAQ+2PCE/4pXdXoewcBdjNkAegkzu7Vr6Dj6UfoUVaWtc+ElwFouL9ovdN5wSL
BqzpX3iQBGZYGgetzxn9BDh1kpf9Ck1Z04rpfIsXwlQopOLUqQCise9r1YcTxh1h
WYy7QaMAWYZEVwBROItRpI3QK2GYRC8ZC259MdGzkaHM/Ir9h9tK8UXqqXEN/VGO
qXvpUccfVwfjHynJrlCTq9NzebNWvg6Wp749vEP/fXRCkm3VRlYaQr/2tMCqqWlM
jDtGICOfMqnSUIHpyBZ34WmEf9dUC6cKhVRaJFECaEkRACi4+kZcUVisXT5E16/T
6eqoxBQihRxKwr/c1ar3Q1bGyNNhay5omomSyMjnpYI5qPnegAZMEmKEYKR1vrbr
4/D35Z357OmQon0MvgYlKq4N1aV9dUjolMFY6pdaWN0Yt9Qv8mnFm90gpOMF7DDa
DVbRQiJ41QYDzAX3QkaiX9Rd2rxEyUuZ1DBYD9LFRz4AFSYgGvVptYVw38yWfAC2
JxjiYe55zAhkJjNZg5u1/qJgV6lcOBWSfxe+9ctki2yzWqSwIcog5xjD1biVxoxD
zvf7kOceePt/vbjOtvq5LOJOT+gxRx6PtLmkPapzKtA1i1TnEDtrZtR8lCT5plKX
+/0yfIVURt7pY/MDQcQDdJcvmNoT5UmKSLYW7S0pmK195n1WrGEzkeEjWuJx0CwT
8LI8muOqlXmvwosvxygmDnhoeQ5GjeaDh72wQXVmYwN9NvDgdWpcJE2sl3nCR4wW
ESPLILTiF3/Cn8q/sydZwvP4hxt6te182hE8RHL0X9Io5hZiZL5sb6T06ykPA9Xb
T7+Eg1fDcxZu/C2XvZMUfM09yswdb2XOyAdkwfIVl/5y6C0x5N5eKJi0D5SOORi5
NS+S6yk70ew6DAqmyAWvxk2E6O615oqq109mA4Ldpm7VEHXc1G+a2af72FihxWC5
V9SVEA2J6oHZskziiQyczYYrJbvIXWmBjSr3E3mJFDLmDfBICofi/gdMX35rTDME
TsTDsChqp91d9ia9/mtE4B0iCJKqWtcCCaCSZn4qKgwNJiuvtDlHfXU/HeEi8SS7
bfDJIrHyNi2/fLsJ3fN4a36zNlCHcLwAGEjpksY1l8xlNnkS5HowD9oVnuRweA8Z
6KjcpxJcsgDhGon4Q6zPNehvC62BC7Lh0PBHuV4Q5fLxH9A1D833whi88clZA6zj
Pp3dKbyQcWQmpirmKs1Yc70JiDUf+ETGD4C96Jbr5gwL2o2o0yWgl5v2diBpanLp
OpmatZ5WB9873gIKKE76bWmiZzWs+8akOrLvv5mqMzu4e91cB2B81FKk6gJPSbU6
EvNxaFcB0/uRMBLzSG60yx8opJ8FvxSJ53LnTqsfELDocPf4x03qt7F3aIvvHbuT
7y8EVSVnyCsezMmC/9ii67krUEsQQgHSSBR8bAEzxzWROHP0bpCB6d7I+GP00fPj
WRalhb58VJPcZ2+pmom+BwV6sGNNfZlrc++pTqsQTs4+1OqGbXTITPxV2Dn0WyNE
UjARYzrHTH2A2VhQAYWoxD+bbYf9dgemScwz+j6bJupYv76ksCZsGW9FwlDTboUE
kW9IDjQxkh/6bQmOs1AfJl3XJwDOBJsOGA+HWJgMivPkCgIHT5OhfdVtjRpu3Jyf
Fd2hvkI28pA84SaLyKMwmaTUxYXVDl6JDmbECvFrMbLhj2SwE0UfhyHYGdYZ2tsy
oR1ynOUNJuAXuSOfN3CyNlqn8OAw2QPSB85ZPKYb4rDc3uvogH+QOH6W4uFj7Tmi
W/cImP2STzi32iNj8aJXCgrxBpkpYuYFK43GeSPeZzksXZmMsk8POE2bh/8A3qek
+Z6yw6RcDUYLJ5IVKeCeHYZr1fZqVwa4x8DopROeu/nEBPDAvZizRDdyKdA51g/v
3lhD2zV8fSG3nGdzr7nMr5aJGPJyK9JkpD4fGL3C4KhmcnxQnXnTix3T7Y7iuwKG
F37cW4JRu87LHtimumQaTI+mzzvstEz+c7kdnaQq9lZ3Yxge1Xj9zHtfF9z2FVvw
rOv/IFM0xuYzveR+Qufmq99TpxXI45XGLNLgU0xgWReK2UOEFDg28M04GOSceDN7
PS32N/mGi/id8n0ilWuX3VUxDGyWeKWQAlJCgkFznwCf/K6pJXmHXZIQOoTrTdsI
rRACklEVr9xcfgEWpeHNVwVzauv2UfIUAIayPGEXWH5jU+rkmBeGC8Cik4BmpPt3
woJGOy1g9tlH88GCVV8SqYUYCKJtPfTX/3+gKXp0zroBV8MUTHTgqjmUYdjibTgp
VKu2Tj3Yh+ddE7rHvV/IqJjL2T0bXv89UVKThubbYmPxrgVOm2rJuAOF+EF6oJ/V
9Maxi/V04VGhgS1oh1w6PueLigokgEyIK2nMgGoGarD+l6aEvEApM3uZdeJ0XOTa
dhQW1iLkclEN+CyZ6vzuUMDMAbyc22dfuyGUC1mTJYmVFJulNrQLf+OUuGhz//4j
DmCKjwn/uTXE+2VINARYv9+ov+ub17S/JDYUnyIoZUg9rS4Nyup+24+JZXrc4fZ1
hWnNzbUfuEBEbQtJEpRtMmCFDvfIi+sMMf1FW8lrF29Om87u8PxVGaFEYdkF2jo5
v5n8qetYmYEfeJYGpv+DkQ8bbacQJNC4fsFu1V5RX8+PCAqDMWkravpXsdTR7SbG
timDRkgk+7uN+gR89zmL6Ly1PM5me5Hfcxhu0gj9QI4enVHdxHz1H2vx4pkPuopW
0An7HcRolAzamVORMQDuDHpF88rmqKxh8QzW/YDjQaitVjdkCNHNmH7mOx/A+I7D
kY7yvxlXx/WklkPCoy4OqyJCU6tI7xJSiZmm0sVEfCHIWaFAXfD9vcRKP0yH+ufb
k8tFz0WqD0ZkGVyKeRwkRLwxrXbC/F4EC4XGeQoyD/7Dh+4puL7ogI9zt27lTL2R
TnJDPlke5x3RaSG96hFf7CTczLy6/8NaZq8ojODcxkcskNu5DmFtezpHPFz6fQGF
OkyMbqCQE99NZmOtU09xGWurXc/cfFAJN1XIF0fHVh4iWwHvKVEKfAtFsFxqlROa
YV/BrFHJemBl1zWAssfwNYzhDxCNPZ5TErNoC9mkq5f5KqgZ1Z08AC/r327dvAga
lOHyPgffyza4zyMXe5bCZuLrIwxj/E4PiGMS8Dc31qhxPLhjWuta69ppLwMOhPN8
i8uatD4gn8KdU/nrhLrl2MBaGoEGynNhICz63/mbLREs2wsYQodq0i7VMrfUe+jv
hopqE9dfRjSK+d1czlo2/AlcjW+gyK050Pwyr1oiyXK71XFq6qQbpyQMT2CIl6hy
rpolv5R0FQvPodiM6lRThXol31njqfJ1sPSlJ+yDNY2SvXbT9+BEmaDYTPoRTyag
CVgDh9xKcA6+HeOIPmsxpR5LgO9rRUjJ33HuZoZVZAlrHtrtRd7p9d60niITwqrV
L02/N9hCo+G1BSVcz4Uhwe0PvLKfQkARc75ARAkhbtOcXksbfo51Q7cdbziv93fV
kyOxlpSHePT1viFLZyq1/cB9wDwekaXZc05zptTVeZc2eFMt6Y7zD7HgvgFuathc
Jkj9ZR1Xbtgy9k4pihwlmTJqgYM8Agc5WGCBWGkODIAClWqtrVqoPvhcdk0giUYg
hQSq6cRslJIRlRZtofqZER8Li453CAqy78HnXCzZ3JOqHlffoZLdFsEVH5zZ5S7P
iCrim5YHVfJ28wWeDOWmh97juNu8f6RsK5wHlvq0Fdw4j8DSPGjpphbGwnEvnK4M
0E4nRm7fvTs0VJpOjZ7F6ksod8KZzmu5DfiAcHAM+7LKbhrEvRot79/FPhQVreUB
rA3agjocBls7NvzD8I7qPT14jDGgf04GEtdBy2RgPMSa2D1obNlB8LIxPegQLp7F
bPadLDLvPsqsqSeq4Db689hro4VVaKR+3D9YrImkVPnClyh9dhWCejDDXBUh+TCi
BIaYmeai/+rDeBRyHF8Rfvq32t/RegGqsGbOFoD1Kj2y/7p7h1mdhhg8QkDG6P7h
WpWCYw3b+DrZqwA0ZR+XqPfCZXWoqLXKwyWUzoR1j4aa4z0FRylzJ+yEwt06nq9P
RHreBKCK43C9Le18+DWo6h1hU6liKAQgzxNfuTMoGYT0dKGFU1fW/TbF7T4WmI53
N+MwSWBgaBH5CRUDbmX1TvqQzsjg69M96Nro8mKJGbnqx77yGRV5FjLeacVZfHYF
iUUSYllDELPG+VoP2XG/Uq79zuOWQUXz+Y5tbUVoyVYMIwJx8R5NnhiEcLFhBmbo
Jf2BqaQJo1qu8x5pKXb/T0jKdVDpXBaJfd2hQOJ35zrudbzRYuFAJ73tmxy+K58R
bU/kGi+CGRsZu+Awtl0KHqnBCTEaNdgAqutRjAKcuaN60g6CoDYDSQM2h211p01N
r2Tq3ofvQ1DFdtk27a9riQ8EAuxIEBA8B59I9qcWgq4BabZF3BFZbVKqKbWa0eZV
AIGJCBeqMwOQDo/qjYHvq9L7AU1c1IEt7TcHt0j4Fw4ZMxOv25kMlWNSqXJfXsm6
6LOMlKYPxziYgifNYpE8GSQnNXndUAM+qWyunSR+jrvumWUOtozWpEb/rab6mv0k
V4hdMMYiYt/0q7BgmAC1FOJmZK22KXfgosBD/E7iEzy85rfojtTMkXn0IMPak2BY
dlqSVIBQz5Vc56vTOpw4RcyyuANqigl85DZIqHjl5nwgCiDbloGC9YGuEb2pnOpY
Pc0f14Sd8ImboIDwM95XbldY6y/lhSYryJ55/4s14oFjAANjhM88OoB35QQ+F/6X
uKgqBqNQI+/ifo6c1AsPMwODlYcgU8bm15s+hIhYrhd7DMgSyrLwS39xPEpAYQ6G
F3xmMoo3KiuzlyrZMTbe9MJ3L5G70NFsZjeQi2Sohemh+SsMGW+zbYJ2sIH0vajP
IE+DP5TSm1KbMF6knF+pvoN2Do/O/nH52qnrpQ/wCYNi8jRH7T0E2at69LfARlWQ
YDQS7pSGSPZ8wlIFx46rjFNs0utdY8YArA55Uwd2Aj6mwlRlw6yeJRXR4gIZfM1m
5ezGWZonP2PQdQvAo358ybBUmLWTHpI06qN1iUQ4tiZQ7bsLkET0d16doF7icwEl
51EHnK3VmX1s4HFahkO13VeMvjSzR47LadgbKRA2JwhvmEHKKYbbqcdeFnkgFiuy
7dbVBi+uIte4CKa3okeS8LymiiDTU8cmroi9SxSEtwFh1ag4BzsExlBxVRNZPz09
Og/gJFJNbZVwt85DeaRDWJQpgDT1RHNzR0EKRjLXqZrXv7UWXlTTCNh56HgPg64V
o5oATM1KGDR9CoJf/28IMsJeQGaE+Bx9ZIG3zQKG7/1H2dbhpHBpolqO6C+BOQzM
hkZuzGbi1dQZlzvo7wJukiHaRWA6xRaibmZJGcRF4Z8hRaJiste3ThuaNUmqNbqJ
+7siZaIK86BOS5d755I0bt20fWrt7UqjaZNORp5da7KxMW5uuPnHnpqVV5+a3D6g
mkmD/6kbtcbTmofkUysQYg5RhFnMopgD+IZlw4pw96vN6lufMnQzCQl8lylseW/U
WybDsfQB6qRaDsYkawinI7+O0NPPOXTt+75awpo2Fkgi3WNOMdgt2CyxOYj9IGSy
6EO25HoChUmeiDKoayqYPYUszsk6vSiGM+jw+c6srhVz83j84xMpY6xO7jENsggA
98DFGsvs801pECJXTncwxpYDks35Mvm5a2ccbjsP6+x6Fsxlx/zp1Qvzw5tfajK6
gIy7eDDuCb05KTVyLJc5Hzm0BmQElJbIoQUy7W7gZ+kZvJLWcwrGLIXzaiyeK43h
rX9y52vNWFguZUjsRyRSK4LT2XcoF2sLGSF0plsRlJsfOyIpnc84MAW27yQyG9PO
lEEiqUQRrMm52HJp9FvI+M594K+y0b6X/KxbWomWV46lwr+3z5NHvNANAjAJZtAy
Q2Av8bE4rNyDRra3ilLuktzM6vacsid06znOnf1hQ2UKiRFnWF6t5dUdAM/AszLl
YmkbdiJ7knHI0RBuIJ6T07FXDSrGJH6QFJRSIB5dW0WxIDCShtLF4UybdUq+OyRF
Ga2R8QdIDuj9zTdVGnMBQu3vIHEuZAvHlpKTwsTd3kOTtm2tj0Cfd80Zm9P7XSd0
OpVT/taG7bDTFyp+RJsZJ04NDiqvgINQd+kd3ISwz6whxgm7ws7ZsvSvNz2vb+dn
ULKTyQmyvNL18kM28wzrNf5q63e3iqCxR1Ih3szcYv7jc9cOr3Q0usp+DF+wXCLW
nr+8wJUozDKK7MZScttEB1MQTRQQcGABubwgho5CP6p2wVUUNsGqe1YQPE/VQlmS
andHP31hW4aOeEo8ODcd7lUei+ZoheZDO+oocIvXcg4olkPwOpy1qcw0pL/bsFx7
ll3ju/khpmk8PL8h78tMQCvYK4PCDkv/TQSvdPF1uKngvyRJe99Hy5AbSBsrdNkD
wT11EYLs7rMQBsLWI9EtYkQ5OkcubzRISm/I4kwJumfYCaKV1evKZqOPPXUNU5M8
jwISeng/ECrISK/Yq3av7bcJ0r8mUll9rA8oK6K8rc1Nf9BViekem5MV1nw60wWz
oewDO0LjAgaQKg2aGWi0VHBkTVe7ByDAikujb/YWoXkfZzEbJhN2/a3hr4Nx383h
B7mDK5wEobe4zZSGdlydZ1m+/dhYE6ru4Xw9cIBRu2FGW+Oc39L0gqw/QDI0THOo
EeHmu3fdUHkahDBRnWBiml4xfrhTNL6r1dV3viqJHYO159ZXkJE3ghkptjm2IS3g
3ndh1hIFJc1aE/0tdlNgtL+ZHsTZ2elD+EpksVQM4WadjgMq5TbsZAillLgdwZ2S
8CDCvEtwcSAx4a1jn7uahynpdbWqcRjs2qMLHc06VFjmCagJBtA0agG1o2A2rzke
vsUjeNRfpTX0WVu8JguY8JTnxOFLlHgx+u7hL0a1IeGHGStc3T1Mzu7HF/JBwlKx
+nr1Eyyok5us8oekauBpSLBdiAPaOLkba50gxcXcXRPdPiTifIJEIN/zkWvFwpR3
b0m92EraOiMY0TwZa3BYNrgQmE6M12/thx2OfjKiN1H5qn46WuPSopsvDrFK3wAC
YXPfRt7ouk0K1dfSGfJs+ivuNIxL+0O5jCL0Sa06+29kXXxUP+TMzcCs9WzCNoll
qAqmk1Vd63sqghaW4liFr+lgOocMBb7tik9ZvXEj/DTr3DtTPHbab7TrV3LBGdrx
OiQHB2P6zZFA3YJ6OVc25J8m1YGrvXfA08s3EFOco6IwtebuiOAtbn6ySbRLp80Z
8p77TmbFyiZe5gLKu32+Jbxwued7dmxn2kcCMf/QCOTyyAGWSzK+UWVO850JrdCm
ZrM30ralORFo930L83BwnNatd4jgiNBrhVkAGVjwA7uNQiH5vp7hzUF7YWibKcPc
Yxah/bO7V3b1zhb8nkwYkZbkh7jlvtnrLRgOd3HGjdbqHAUCxzJPAyxpPWmUUudh
dvVx9CfzOMd0LnpLQ+zq7nyKVvfSuz0w/I4Tm1CNPgtW0+4r5aDr6ELtvMzs0RRZ
/OMKvrAbCrMrpnvmGcIQZ49FmsK6H/SZVfFi0p6t5pmYwlBy5OJfFbl8I4VxHF6t
o+Pq6ZKgBZXKqRYbHGkc4s+sn4SRxK4FTWmIITIGcSIstvuW1bYLXX0lU0EwLnGx
b4XMcuHmtoxV/hgHXGPAO5KDet7CGXYIFIG/n6X9KzIcAO1GtLn1gPQWd+qMDwza
yDkZIy57IKfXqhh7yMgZ2ecqT2lmszmrfMrPDXpqUQOt0YmwoViGW6cg0G1vG2zD
iDzCgl5NiZzXF7tl4/lGIeLgpwmIcCi468tC5p/sxgll6Taco9b6DUxGfLYt8cnv
SI52ZGWfRKB52LQBp7n3bg4M4AuUWz/lmx25sOQsR1sunojxvl8S7Hxt6XADeEP2
q0Llfmmtw9r3NAfzz5h9lQvWPa9QIvP9g/EJ/bgAIQQMBtJncY16cHde7mJM+Qa/
gxktR8EZj0eJid0nOi6nqeeq7xFlD6STMPkHdK8PEeo2EHS+pwN5WunVd4lxBEFn
9YfPY9o4A51pFL0BkszZ9T3qFjJIkAt6aBctsIlUvskYA5fV4DaLk6BhcgR3Zxc9
aSXmac86JImzYHf7SbEhh4xjYdpw13t0RihKXf+Io/FFkt6nOXJDtQGL0Lecu694
MzoKxHLtSA6D2ME/hYkbP9MvYrGSkUueky8qVwcUvOoMv+knowK/oPrk7sQ+7T7n
vWMNwAgQPs3Ck9MM1e0nuMGbDPeEkQag8sKoijNCkpO4prG5X0pwNomkxDMpI9qf
szWO6230NG75Vy2budIne/YIk96sOLPAmSIVSQjU/f4a9GlwtiPfVQCfAxGcS/Pn
EhHTgrU4JhpSchVxmqezGW3//W685Rkr0iQZ0PwB+ByFc11E5KDqGxP8K1nd9J15
C798ypgQcLSmImmz4VUa0Pgz8YXjBtLlvncUzWuU3P7uXL+Aphu41awjpwewbAWt
sCUMU9ovawQTQAh4FiZdNaJYUUcbO1eFY11Xa62U/IgBulNdqO/AUGCiA7df4cPm
l0PTo+i5kMYnf2aLxF6TfqQFVRhIWHeQiQTtxuP7aqf9FceydqyOnHZ/WFcx1/Yn
EWWgpATR/s8r8ZCLE1ju8HRMSjngM5viU0XBea5y6oL6emdY8abSOHpL/nKWMD9K
ysZXKAdBLd6PvGhi2Pu46CseGiz3nvF7D/2TduiU5MHjmYMcaaEYeBiueaGmpYO2
0RTXhTO2ehT6VQOCHmTF6ZaYpwnc9cS3lrBQjQc6eWpAqmWWLhUrxgwOJNUE+qd9
/S+6nstKs+jGHr/DchpU9L6atW78Ju28wrj+ys5oaVdwBRT+vPgok/Vz7U2LqQu1
xTYui2TibrKPEu56AUxdBMd6HUkdcHkBXWITttP7tVqQvEJyyuvt5SIkz8mDB9FZ
CfKcscz/XyO+C4/Jxx8N4itW8VbIvDX561pBLosAxP9fvUrWD+oXfzT+AVlERNQR
fH7IU8sN6Mrg3c9GW4soDVe4qAefwPWfoWdRSx6rZ9+3kdybXl6pF2lOHp0Y2ugH
x8zBY3Iksa+aQme8oWnbODmeZCsGDJ9WJhjsne9KKDx3edyA+yS2rK/9Pg3jicRj
90mH8LPUBFJMsRpJcbPYZ3mXvYfU4L5CMgPy05QXtnsc6cHKaMzaxChvB/tyBhGA
EhVBwaXVZJnt0uPj5kd5C2+/RAItF6P3V6k2OpbqYSngeooy1B6gPF4tWulx0Dc1
DBbR/R0xUF0/R7+LEs2s195vmxjqCl6fWvkYTSphmNIuJdbIiOa6H78kzQn3xtQk
V8nW7DDC8VbsBmd/xWOfrFBBJHurbld3kRpLh//q29/e7vR4Ox07k0AHGP18mGrI
xLHxeNQkYsY5fx7EusIjUoEbshMBNl08MOG1tD5t+8exo1xABNz8WKp1eMhuVJNY
vIf/DWxnONNeQOkKRuoRSWAh9B1TKe1yx1TT+dHYFVD9KinR1eVh45OjbxVE5PAz
ObWrORbOFNq8BErRG/e7/NrzDDCRSTQC/ghD11dNfIIsCZbTugpP9fDwKeXsGdRQ
FOCGPbYb1KTxrCPDfANY78lxxFujDDLAbgmIWsOvWKJL4UeVhV7Y+BtkS+gWKbD4
0FqyPcOoFeHcp21Lq6JSRAv9LcZnsRzP38SpSOk/aHwr4pNkQ3LwVFdCnIcTF0dJ
SJ4lqQ30+r2OiJwlxZutNQ1XR+GHe7kM9CuU4onWC6kMEvJTFSW9Kk4gbDx4oQ2v
KM+wqlhvWLPd2fpDDHrX7IYTjIf55nt3w1Tln7FkFiTeoLi6MnYbEHLlvXc8OpwW
fLZdhEJCboLLJFQt7cWrh/3LCHlUUf6/THJdvTSutHo8xW9kjSAyanP24xnyyJss
pv2GXMlxV5owJzpBy/1jxC5xrF4pkByW72WNnBAC3vlLyd9nflskewXj0+1t4Cd5
dPejxFlMQU8iYxxJKYCCeYifNR9AV17dvSK2xJwZAFePJPHsAES3eUF8xnBH4S+5
xYJeCH7VEPFmXG4ET7VGKLL+Qi0jQk9BlFdYhbffrcCdbQVwUfGlm1RPpKJEFao5
7kAYbqJrAYDEHIJMuHEQrIK2p4JuCeHMa83XpZy6+k0ARJowf7vsgZfnxPOJAnjX
tQvFUEcfvWcGYriQ4LzZGtKLbVSVkbcouTMLe95CE5YJmKdF9SrXDXV+SnKA8VfQ
WowHvxbXQdu4zZa0jWS44OJ68eJQK8X3ng/uuY61/3gcYC09aC9ZhoqUmRPMWHXU
M3SYfb+r0Q3nDhc2Q5PrlEEmNWbCYtE4E5I1F34IvF8x7+H1oQysWfWB/kePl1Yk
FRRCKYIP/FjLjm6ssef1vP6EqcqAIvqqqKIqzmngbvT4j2EH3AfDlqX05SW2xrJM
0HLl4R7QSCQZ9pOld+Z2zNb+s53XhEri/iiMEEubbFilu1wiBBo9MFLPmwq1hNWr
kJ8pZafGksuyQAQIpI7JEUs227vvmOWRVDrBspfkdUgiTtzlFXjicoZCJ2JYXC3h
PUgh1DAOpPquzVJ8jBTovD8NdaA+zoN2h+EqYq+PXXVIjHp4qzZLM/EcAw1AfmQC
TnMMvQrMLHrJdtPjHCxFi3QN2i6iXxhBlgtzukPHNLBDWbxlLDawjwUfkbtwuaeR
dxBhRa1dVd7bRPNsZHZxqpZs4zJgNJwc8iX5j4p8Mr6CNBdDh088JR15rzFm6qE7
4lJ74JfWtqeK95+ltLrQWrvO7s02FK8kNoRtbHv340m1guru7hjTnBNWc1sJVEXp
Sc20q2VtBKakRBWtc23/KXOrMK1ymZlOo9pqqlCTbVRsDIXcZ97AVQBUsujzLOSr
ERY81Ih3+lPMlAIFJ7waSmDS6xzLksh2JrcTryPF3xYAPxAjDmRE2zuUyyPnD/Vg
72jzs/X2/tse3l0ygs9Kd0iKgIVRz3nqgwyjMfjFTC0eBtz325zzR+jx36RVzuwv
LKTfK2eiKRQH4Ev+EJWyYCv3v5H4SmuvWsOAJBVd/1QksQyomHZwvIgQAvdGJraS
KDtDjoLaDLZWNcyXD4c+Njc8FJAXRGSQrBjQvsTJ0nH+l4G94m+7bSx7Zb98yIAF
kh2HRiN0URC3CK1iZrs1oq0g5M+apDhzj23m3Eu8M99Df1cvcKcci4tHwiTBsx2G
c3WnulWbGtSBXlyIwiBDPyf6yWhzO6c999UjgIhJqaNLZX5+EBw7uUMYQCKMz96T
yrIMfGzQrAI6sNjZ4A2boBcJFRjJF2nVjyHyG7bQqvgG4d3Y6httPUjapNGz+aaB
TVApnivgKsvPXEo4cPevlOnPE0tpwyBDia8U8Hehp8agcE9j1oO1QeSpwd6A014o
rv3UIeMCbeOX1SINGzn6g1nEnkmJMfAE2R6vXf/Kq8j+nmH2PcM4ZjDAA9Ck8Uj8
7KG1PZsD3uMWaFwvX+8K19Y6Kn+xOm62kfA8zhc988Ke38qImTcKu/DKIy+jfSq6
+AlWeFTLn6gn+l1VMKOlI5ju+5MW6BUR/7c3N9jskBpqjEYmo1oh8lSOKdNR/G1t
DKKeu+9B+aNGWSsHsvVPRDEAXe8lVdj0YusCLFk+AVbdhVXSXwe3JMrl2orSN4Fc
WnNR02MRs4G6bOkrjc5y22fep0EmnQze0QlLFT0WmmCYYeqF2gmjvA3kBZAAeeS9
K+ewTTfAmcaGYfaiRgHhtnDqcNm6s4Y9AIKC2qLqS4oeb/XO4hDxKJlL13Io+R3A
ZjgfSiCEu4aUTKSH3mMO7Q+TkLpO1dGXTsyjdUx4LTClub1CGMsUTYqfMycog66E
O1Xfm/o2TINpSVXL1ifL5ksO+PMqFN8PsHFzHXJmVH0jIKRGkAkoP1rpBHWu57eB
YrKs/ywPs5ClxFckk7VwWmXKKAoIB+MQviJ7QGBEJFcvvOKrSSeMPIbJHzTeDNqt
nuBFP5bNpZVozFPEhOULEbDGEWzioh2Te/uwEWTc61yO55XBTH9lQ0kGhSzYEQuc
4QLaIhYhSxEYEWsiFFUA53LscrySNA9/GzMp6zmtnZsAQHh/5HzkBAIpvU2PqINQ
q3PV1n83wDzjGPcGd8/GA7SqLB6h2mK0FS+Mm6qn6N9AhG17OGCe3gMObKfy3Jub
cR1sMgoBRgD/bkOviuW1Jrp2P2aiMMaGkG9qA9kq2xZ81kM98WS8aqPoXrxqA+aG
tjRBDuoBYYya9YnKmhVqvkapycr7fYpP0n8i4ovzJ/lY0sN3rydOpzA5YgeSpefq
VTKy5urjk6sSa6QmaQJ3o1WDc0AdSUaUMHCbj1HD7Pej4oDknZDV04ZSrpla7GwY
ya53Y3j6/WT669imF3rn1ZKzkZU66tIYOG/WgWDdV2JmtIYa1ho7wx1Pxu9GDI48
k+zw0CRosPJpZt6BBhxnnvZvogm3VCwiGczBKB0+AfKXc5rxGmiOQoUuR7S53VDD
Wxk/0FkFMzeggsdVxJBAUGxgX/Nuq5KVm5e7SIuQShF+drd4keJBieZ7hWTrBQBZ
/dhgDK47S/djU1QhGIi4eboQ2/oyx/MUeH2sdt/RAfDnELOIP2c9DN3LkIyH1Uhm
2pMKaGR9dvkwyY0IGzXsTdoJAob6HeY8vQE+MANtWr1VprRroreInH1efcPtzOYG
26tiwwWzsGRHHL7Q0puhOVlVlfpezyC2ply4Px5FsKLzHN9SUSzTd4ivo9N5tJQP
NT5OcQTBlP/wZv8CLSyROjoBh+4hnleQt6zmoU+9pC0SMLG7j0VAf7djGV7iRuQY
CZh1jLALC0Ymk0Oe/zxPf4snzyeRl35z9iixqCzcn3tCBN/MePE6hyvM6K/hXeMf
HfPZi1SWdnjulPc6HIprx51JRIE9x0OUzYMiM1MKmcgPHwtwAntMLz9w1122/v0d
2M6pUB0pP50lGKzL0GnWhVps3ZbLAfVTV8kMo+36rc3HYYsB8qFjgEA6YNj4P2vY
tQDrNE4xe08gCT/F/yEuoMea5SPhIxOzS5pvOo4UgG1vPVZIbj/TqJMhu6zTtdG5
XJz0hLTSdOmpOhLzGX7ORec0bHCznHGDf1RshXo2luU23ieWwRw1UIOLB+t3IU/8
DEhC0HsItplgiCIgJ6sqZl9qyClUynwoi846Lbo5l32CRYQULi7tO4f/kWJhyVET
R+aibzVqjiNXfElvHUUWTg8qtjMCi7iV3vIN5gufetiZKUReSw/1WxriHHfRb9w2
DrCQsMaDwJRww0b+PP7kNm8zeEw/FlIlSvnaEq0KGm6LY4hk6AgONglm9TLPyAxc
2s6SxmcFuOh7w20WVsIOSl8vU04b4hwImRXNQKWSRmI4MHjn2wAuMotr9TlKp0NA
ZEnmLT0+DySvN4UOEWcFuLxE+qrHXdjzDWpseE/nKDya4D1UoMVQ5BX+bQ0b0/k3
PJDURbIyAcVfDhg70loN8JIHnLa2/lj8D3/UN9F2qljbbTOaSXrGqnEMbgWYKQE4
zGNgg0ZTtZR1upWhAXDa51OAton3ddS2mEyYuAwk5lJiKfpJPfpPOjUrWwNi//iE
1VsKfoweAxjm/GVQJTijTHxZBVO+IogEPiOKQyWengnfiQ3oCA+ZS7Ff/UbDeHg8
Z1yqutcNfl88Pow7b5dzJsLG1M3/rWYoloneh92yQkknczIBVoBJOu1k76RgQpi6
JwtvthKhx8Xe7rxRklDNrXgDcaJmue0VHM1+ruZJJPydOe98fml73tB0kH4GBF5R
DoHvAIOJ2x6gs9gVbtUrXczpRhl8nSnQrY7QFjKV4D896NUfR8Vsg1DYenxnH2bG
RfseDsKE9IyU6/9xewUfs6FDxJNOKHey9a5jDSgz6IOOtqkU52qNIR8f18vSViVm
ZJi5rO4nIq/X4SwEJLpPYJ+B3gy0WAz9D2KPFRc8qpn2VGz3piLTsbqnhtsbw0Ph
Rj9TTewK9VdbP5nUjOK0qvjk4OnQJhE2RZslOOaj2tesB99TnFbAZUOSxzrDhY0R
zHMfIys2qY71jZ7ye92kdmY4+eCIe3fm+AFAuCjB6f1vCsx7r1KbS9GPqRb/ab6S
FuKORBHu+bI6rq2qNhVZh5sElUFVPO9EUT6KKkEAVihfGElrry+lakQlxJEOUyKI
V2tufCyYOlpI7lK9i/RpatRmlczD9x+W0E+VKQVGTbjKvdPRzD96VGG7kQtrufjD
6bTV7HMf1rAY6g0xfjtpLjPnA3IYSAYk1oJnVKAbuNRCCNwk81bVcMMbziuQdi0Z
rymuUIIplo/N7tzayyIUhZJy9tZAPunDYLr2El6mI7jA6Pyg4LblK3QqzIJ1pOCW
YG8E2n9n0UFQ4+sWK5i7JlghSSlAEWjHFpw3PgI9fDjSC3CeCTnPP2I8lpg+J1mp
q688TCNpDW+GcmAYhO6qpS+cjT7BXVUd3XbWj6Bas5kO/byVp3m91skdCmB009W2
8wJK2TIDgrZ9xhl+yUawBq6GYZQisxCMkYSwNb32nsW6NkQOtdzV7WhndjFhVSa/
vOWMAjFjHT9CG0Ts1QklOucJ+4rVIrD9WqCMfG0dCeQuvH57/B8gRGsJ4ZMWe20d
TpuyfqX9X5LXirRCUv09ni7AGGC5w615MHsCxZZ507weXs6APKQhyW3euBDOlvH1
wL8P1NY3RpVg3ccznVdO85cMT6uwOJuytQJ3fYLVCIGQ0pfP9w+w3rOWCLA6Xl0F
E4/icPQ4elkV7P3Fqdnb+AOpJtvJ0L6GHGkq3qCyCf11qJ+rCaRPOHHQNbkmBt0c
QddemeyEQo2wf35dEsS11BX+1r2UQHLc1+5d6R8tyJH2C7rAoFpGpRMq7E+HEd72
70gb0SpLGzk/SjN7V3Unpvq+NSgbmd6XIujrCloRvt+iQTFmYjaE1E7ipMk4cocj
unO+Y9fK+LViNtOojNQaVvFahmEiP0rz3Nb5ydjoerqVDZNbrX5eAZh/L+vKRGWt
foJwl4/Wldae/peBmajDkVsTiB3lav/XyAJuDoAzUcoRcC1/7rksTlOBAvCWxPvC
/Y4yFfcVyB1l86cKW8JXbAJg8Nl4zLnRrSbf5I0Ci49Ocz/EUSAWGB+F04ZnYCA/
P9yGZQDzvn9zYMVOxWod4oqFWb0eC/cHhso69/8ZdXEoWXmRI+s984PFJeNF+97f
ujCPeaH+16JG0QNujPkUOVKFy+PedT0z+j/1fcBwRwoSOkiwk1F8eWaGzZ+phGVP
uRrqctG2T46mVmqVr070C7G+5RVnE5XS0YO68xpcbgFewiLjF1Xji2EHELCMF21Q
xdeyDYpyL+ojxoo8tve9gsoL6OUIz6tiqp7aiPBdOm5j7UnDqNda+palsl6aq1n8
Rbpu4BgzHehHP9ba19mX97oer6y9RacTGu7CPVQwKoGVhL2s/DGDLpPNz86iczMD
DMUchInutJ72y4MOX8y+0OeaDTHwOz/qyE762fH8qhQlN4kxNllkgNQn+RBwQVuJ
Si9Ww9DJZ87OkJ89wn4Skyk6jY8KINFQrALTIn9mVgXwAXKCKRM+IFKIh7BsE9a6
57mxl6Nbq8q/F3eSEsqcqpkpBEw7U1lHykAriBoK1HU6D577a6wTv7IbmwKZyFWk
Kg/roRObOK7fbyXw+BkLpR06ode44MIfdbV8OpBdQemYz7j/C/9qQw7aJW/18GaN
94OxrIjSBkKMOwdVEJfVVgR0/iGHebdWsbhZEMnKCWvxPjjf+KITZuaHHv9fUluW
J++9nCDJhaYyl+26OrA1KJw7TcfpMYuuX3KDev2PG5oL37n/0R7qG+dLE8AbV087
IzYn/qGeT3goSgozL9q8oVgS8JLBckPszLKpqA3vcfG2RyBq8rYFYqcK2C59US0w
0XOcJ+aaTbfy2/R7oKANu3wwm/AAFPpGc7mxnWu0R77TkXxUUBDFVaHtw2hdTg5U
dYcNMkDwr2+OHy9DZaa/CS3RPRYeEJsDfKqPNZy1iiV988USOMDyijar4oPSQL3F
LJdlK50N2maGPpzsi8xBwj7pVWxqAYSGtGD4qz58KjfTVrxMQbJQgI/HWjkH1/jG
kbdRDFcg6nJq2bQrfBMN5Qyn3b9Yt1+6Xv/Y7vEqbdZWG37LMiIttVNxUN1NFjLQ
dQjgpiRUK+IO+CMg7v8jWnmf5GPvEZtss2yrqPrBN4JOqEQOMyjtaAX4TXW531cq
UVc2jqY6NstMKRo2R4OaPs8GX+gES+4RzeHSTM/i/h+vcHQm8wm7BrQzInas8Ikx
6p9FDUdL7nymFHvt0G/mpmmfnA2lvyQMC1djkxlae+Re4cLWitoSw1dmzPG3IopQ
0dxQbbIiAk/jUC7/bJ3sBJjoPPVsl2QTG+30ot5/VvAgSfH5XSd17nr84a0snFO2
Tq3ujdlY4/SoqfQsjcEEVBEmdlBnqSwT3w2scOHh0YSVw+QIV50Zyc/RwnS586Lz
ZOnDrqdYHnTsq3usMbZkuOYqFyybgcR4XUqjrnx5+ivl6TTRVTBDid3CKTz+EL+7
Ggz/6h68zsufgnaso1+3YdhNnNQCOy1JiuGZiDSp4P6w2hvHsCojfGhTJVFHBMie
4b2WyGRy6FXpBgLGCzzFnEbgDtO7b/72z/Zmo2cBX2Be17DSceMYCBi3Edqc5ZEd
BmardQSAltUvavomo2CVfgpK1j36Nnn/0RwL/uthyG6fa3h7TIivelYV3qBwUFrN
SEEONhtTuQV1Fp4FMnPrsCT5QyzurOp43gegxwuIQyet+Ki4XFQyYS9hE7orBEpG
ABnyYZEkpPuGHHfSfd1tEZtjgBF2SIQ0OVCGyWKco6QE5q4sJIVyq+U0mNT2KYI8
JRLh4MRYoZtxInCa3KFQW+BMJXBls1JKIlpc1370bG2oGNWttBQdAw9GMXTgGne+
HJAStDKsK3NDgvn6+JstjjvakmnqrHfMJ/oLCrj72CdDMCIhQThQTrJDusMN0PV+
UQWw+HQS0y+MYvmh/HPuDwzdC0jzfSJtC0jXakP47H+IgLUIEwBs0GFHZB6cUKF0
XaZtQZ8B9OqUiPX/5z8Hb61wqO+J3J9dhkr09wpBm3Xw+mLsbDOBLJTy0aE2n/Mh
sVPrexMp3ew9MJDfuz2RFWIUhKPT5pa45Wh2ja6baao7e5A0JPAn5Bc/ITQb81kA
h6u9PJtzGzoRJ0ojb6SCpRU8Eicnzxd/1GMs9qNvCyFDngbwtzmSPs5mu0354d8U
wRLlF3+2DYzTNKT9Tp5ILGWau9j36gMVgFKc7bDSNvbDCaBcCgEqw/eLZ7wfw3RA
pKB16GEo+oREB5ubZZXD1dSLXhvmGUcdcm07U/aOC2leQz3bZYZeFJMWXLPT51Kq
IGLkbG1Yyt85rRmqA64DD0I6QZW8BuHzMSXJ1woqEA89gQXDn1liDwaQDLIyBceR
6p64VcJwdLhFZqthf+ztdjOYkb83Uwha3lCHRyEoFgwfgWFfcbbz6k9J/G84S1rQ
E4lH65OKqqAP+7qdeoGFaZrep45peTsKj8phqYt/GYKM6+uSFpnLz+f9IW2yVSGK
QlUzFZ1Mi+DLORn3EKMmxRRvj/uGLtAeP7Na4+DDfaNPUIOoywhR+O1qhZvFFBEC
ODZonXOSmZL8MNEzBjDp/urp5rAJAesJkvdnXPIJa+yapUfT6ZsKLiXy0FuZ7ubS
2WKzH3t19E5IU3aw22qNizHY6DL+Qai5/fx7CAVa1Y+nqejLammC3JKNqWXOneoU
DyQVi+lHENWjnOsIQycu8iLXZDx0poBZgEyP5kRzFan7Dj/ZE/9v8H2w6IYbVA4q
HILIld+YoGkG/Uj4ptu83cYvaHEp6gcZ0wmqPKXdx4GGOzZMJJF8RLj+ZOlXc8QS
4auuz5AUSGmwCAcR59gZpYKd4SEd48+VX7QYZcU+xoK8Ukuzt6sEdo/9GMDZKXch
EWlOFO1ZkriSmnP9nNM42zSulkYxOyGqX5X+r4qAZZUa+sEjysm6aw5x6OJxE0Yc
2QcZdSOajneGWIWlzvT5Z6esy8izWOMi9eWza7LHFq/EWlmpAcjcSsAdY/0LXkki
xr/+5CTjVpciu1/HTIdDtJLYLw5YgQLnIky4ytDeGYb9RV5aOd0uB7sAYrRTHCrh
1w2fiqFvvnFPlzpM/+sDIUgaJYOw8Fo+Hb3f0DzlKbLH52OoZdhMdWPP9bsCx60z
1bW7H9E0zeqEdD4CIXcxZd5k8/vC3MV5A5kCayyF3EDVAPe4Z81w929UN40p+/2O
l8NjxTpoWPSXyU+06OTBYiPSU+Ntam9pQD7aDfdR0gO9yAWXbr1HFeAglCd3wFDc
xgTTSCJ26/GFMOw6vf6uUwBYY4B1Z2Zv72/u6ech2kQg6QLC2W/beEyzJtwzsdey
N2E4AryYN0P+O6JmST0FynAv/8O5Y9FFwTEK92No6pJWg4+vM0nHW07BrU8Ey2NP
AxqUuOpWlplv3jxihPvoQBjfAC1Ql/G5q1UKkunU/Djmoc2XpHIUShMdlfiKeyWg
Gc7cPvLAruwRYbUf2+S9fs93tgl8txkGSR783qNg6W5uCPJA5Z14KXOe/vTmJ4eJ
Cfec/AEvk8OfF2XOuKztyGqCMz0YXfBN0NTLUA4L/OOQoeuiMI/T78r0+nQulZkx
hlXYIx1zGfnAjgWPj/Bu9c58tnRMFyzK5PgxAXcIrj1+6mIU1a/vfaGdShuepWgl
aKEUxTu2ySqMcjxv+Imh2Pm9JlGzl9PVFS2iZkVyJY0oYbBVSumZ75LM0CmXPFoN
GreBzaxH79YLHIrQB1qF6TyR3VXnm+30EORCtZ22mekXsci2i/yJYj2UfuT0aHP+
7isbJ2QkLMuHbibMxTMpLEnbMI8kfFXGVdrvrd0wJ0hDxzjgK0wDuDhaKgy9gmr/
oGHjGyk1p3t2T53VtHbqXoTGhXE8BzSmQHV9eH0BvgIBsa3YPvWaYflEAo+4N1EW
qc5JKe+YGclpPO4768jyR88TD0Rc6VrBV5KcZILoiWjS3MXGZk1GAiJhvkQiLxYd
QBwd3fXh7zvMGEZbhJHuQ8S+3xcqDFZE6z846BXFEMemzKp1+eirvihs1lnoKNBf
yFxNFiTEouOfVneX1qtJdnK4QF7M/nxncm5fP2rg6tfFbXQf7AETSvGwlMJHYKEs
fL8CuLyDbBWlr4K4WfopE8uSoV4bIrGRYU+Nzi6MFBZefQwx2FUMmMNyo2YxpsnS
xcXSQNkrBZk3qXM2ssP+L+aOeoj6P9tAoZURQULM4PRhI2xV20ReTNO3DLLA+AWD
kS/M8CrSfLUVWQD/m5Zqur+6vG5RTYwdhNkf2m+R/nPyrY3R3kkQ/qZIh9oqVsM/
xSvc+CkS6tDqgp2ilv7UTsN0k73r1Y5Wsv2P4dT725faRB5RIALlxBbfEed3XQbN
XJ1Atr+Ev7Mi6H8gWTK7iXoOXaPuqWgUW5TmXVm/ahDwr0Hyr2jnG6bxBa7UwdXg
4zeomPNOhzWDqgz/UjdBEPSFhprJHFekBPk4py3EBh7E6/mYBoaBOtKkb/nhI8C8
LWlhoj29nX0ylEOYuXjSYGuEnDaru3VWlQJZI4ZNWXqngwGhwYEA874rnTvih/g6
05BCWE0W9t/QOzOUW45LvhJVIUx6qUtQQYe3vUjjsd5Ew9XINFq8f/9I9FJWKl0x
3Zovbq2dG11t/muooSPrrA+lCuyYz1A96fwfWZpIS8rkKWSBbSkoE97v5JXBDjF6
f6jDOuBGlrZH0+2ooalj4cWPTfXy+OfZYzMjJt31NwEDNh41U7XSZfQ1Cg9xWg6K
lT5om9dx4N+uO70m8LzOqQ6kKKa/MVmbECydKiDpQ1GEe7ctM0ejHR2jX4Gs1k5/
i2MSBykHAxCc9z292XMj0W1tU8V6lSLfjxlbMQ0m5D6kIZgDEqpD32xEdFL0E028
soGRKhfAFe5c+5IvBQGemglwOZkA7lCMKY1NLPfr1pPXr26gbvHakcifCYnjf8Uf
T8E7Ct7+Ywp+aMORHA9+9/FRvW6NizKJ9bewxklNaAIBQonUtB3V7GRR5g/M6lVt
I+NHgvG3DBoOOvM2oEgwtjQg03Yajyp2wmLg33txDEt8NWMAFaHO2tOf5tEgh/6A
dimarWN9sa1lAZBXKUsiQTEBwr+OWChzDqBYpYx86AY5/XrOjcFErhf7Cc3pdNvi
dOVyyNERBzP4lBGl8RjrwtqW2FOXckEHhLCqQ0lQWxbiQRXD248SeiJln2G6q90n
1nyOGmiIwaiaBLybo9Ow08ki6Hp1bDXQ5S1dzbLEl8IMSdxlopPc34KBJIOoZl/C
XZgVELXJqlRTTgeC7gEI+IAFc7VonIzvalbS4mOEHTVIJHIAY48qqaV/s6OjwjTq
NwMBaUnmEBIZaywemGqlz21yeOdGOUjOq5s27H5b0hr8pGYk2v+uhBXC3FCtw8iw
S9qc0rCFU3MQ/X+q4LW/ZyIVRIUw0bKg2cE/n6pw8zp4r1T8rLPdZc6+cEZlo654
xPAl1Z47h4k5FkBe5ABAqi/isES/XWHu5cicP/nqHVpsQDHrraPQGBnHg01oSbJ6
po/KZzDHCjV9BRVouxxBS4UwbDkeAnoFmTvZ72m55kapk8zZa7r8xu2YqAVm6V+u
2BcnrSnpX4faqJ90QwL4zt4keHu3p8Ss/JiB3baFtNgVZ1sZ6lz/JH/Wt/Gpd+06
D8rjvin57CEDWhmvKxsb2V3oEU3rZfOlvlBvQDI/yvIYgEMxShPqbzzropifTQlR
78RKtpit9yOkiyIBkmvL9YxUAuP+xjeomVgn0zrDeFd1+erQERRhlXyflr8z513z
PneA3zMPFs7Bmy3KLuBB0j1xX6p3xVpzAp4ynOxZOlM0ICZ6wHd55pn/zjKDS6PQ
/gU5p+eRflsFNuSbNU3ez1mDhLDFeufvE2/aaaJrt1NGuWcs2XmCLMKtXULjdop0
VwxnAoV9avBG7UzacOeIRW2/4Hp5QgwUD3TmDdrCdNO7UmFgJytofrkEFU5rbdym
VoQgf1fH7B9bNiMQ92ONjNCP5mhko3BbCryuyQMQs5lo7QIBwPLtC8gGItA8m0GT
PW/0fE/fmsIXbKJcu924196rfBFU06dloihFu3A/DJpafMPFq9bLHonmcMJ3UcTE
a0OTxnYXNipYqpv3HENvBGxImMcuNpYHIhrfOrYdEt4bJK8c2///AuTu/ixHPuq1
AXA7gqyT3bKMt9tsZkLW5Bxi472FikBJRDYfnmUg2iIFkyTTPrBU69oq7rC1VCZM
8SxTmNtjbdRJZ7B/WIeqxhYk2fB1Uqo52FTiy9zrjGos9m7lrJN5hx8HyHm9Dgvl
jDiddvkj4gjrkXo90GiBvLPF1axAJzSxLuSUyGiNioeCj6gAAfIuv+wd4i3nWZy+
Gl4p+HzSjrL94nhNRKZIKmfHl1Y4NzRLECRjCKzTjRvF4npXC2yhDxR1XwFFBOM+
BAkrwD1Ax4+1YExfc8MvdA2Cw/5oKLvh4zmSQvWsHcjT/UtcTVYBbdHrrIoPikRZ
1JHaydfzFIBMlN44tAX4mzqQZM47cskSMmhJWZoCZZD0wLXjlyWdQXOx6a6stpWy
a9MxPY6g5l9RwGoh60kMvHvoOO7J2qeALsCzNgednZxN4C4UzAvXyYpB+gXzgU/e
xJFJLmEBaQJnQERX/xRrz2q7pOHPPc1SiA8ufVKszkVJmF4VhBIKFyD9ec3wG2dH
Zmzd+jv3fEAY7VnlJru68b8tWDshiVZgH5bnT+h3YyB6nQjOhrwv2+ffB2mintyU
tGJ+W9vkNj+K057KSXig150nTF7aJUzKJVVDxdHZ5JcN2p1uT1eJKYKWQhqH1O4N
zczM7FgRFbk3nVQy9JkHaZPcs5Ef3Hl48HGMO7NUhNoLm0zKzstc2+OEv8LKmfxN
tnuznYP+EaVRvqvpISeCcqhO6/+y23AkRfTFOjNTzcF8vu/eMWY9CR2ZIA6fJCD9
L9nPhiIgDd3YkRXVEdy3oM2CF/gVwLiUQLgnCXuM8KD9V6iSEgA1INnEu5pVThKy
oFNT8Ev5BF6KL35vt+/Anm9sJyXdk4QhAM3p2Tu4XzxqPYOcrSeGX9CaoZBFom9c
7dibrdWapJX9qBMsGJbbI+S5JSeDEceQxqprB5ud43dZhi7pZkZBvwIxAqWvEuNE
mJ54HU9BReq7/D2P+CIhllYuB9ok6BDjzTfEHfPaUwgVmRTcJiR+EBA9m0MxIsXt
Jkdll0iMUcj1jYCnlBJrm0ZeYsww1femYIRmn7vcDB5zOebfAjuU2/herDtV57/y
uQXC0d9+qUygruEJjK0d5mOCpryRa/1dP2QkvNBZsNJqqnwh3yGrYOG/WEAgTQSo
658jAie9heAktaf+V3VNDpLFso86RNScOAlnrbR1Cdc2i3iZe8LFtUpnBuoquaeP
5DR4w2B6OzEAGR0m4osgs8QJJH7uVWKVPebT1wCs/i2LC2sFJxOV32QOiw6EbI1s
zvHD/yLIlDc5I+GIJnXkb02Z6uIJlpNMVuvDF7LCtaceWvbhG/0bsH6uilLquFbN
cqej9ufSndAKmd6ZCAJ5SXRI3DGLvXnyHgEH03YfyG6DAtrlBklxyWIB66qhtkc7
Ivx6uA+dm8h42g5wyQ9d4IMofito7jtBcT2F0MY9VRj0DGzOIKmohVOMy98Md7yT
orT57w8cx5L6ApbS26dxeV4mHMlRsmypttZEhp2wk6CpSsutP61tVrSKAdh4sgYD
mwQZaa5yS6uMSj4DpNW4+IEGOf7vmvilvwmwSnAPuJqvZw70ifAmFwYL+WY1BE0m
1+ztlQ6Ks+19oeXK9BKZVkbGK31zCq6HK6ccRo0E9V8mdll0k9FO70yLTqt5D83C
u/wMdIk9ug1aWKN9yYiac9hE3ZV5zwx4wzDSmbhsjUL7iMBlluXG2Yo8ekL2txP6
XNFIcHyJ0rnYdtpoI4dDVtyWj73eYb0ozyTx9yCke8HG1MQPwMoDNMcti7O+jkqE
LQl5LwBILkIxBSPVIbTppTGZep7VPQZeZ3waQ0dH434OoZVcAynhREwt8TudRYsq
z52rS+lOed1YILMSdeDk1fSQD4Bzs2KR4zdz0wCVJurZV1L3VhWKDiqgXEmcFXUp
9rJxF1uRYji3fQtsq21P/xo79ztSkPMLsmai8BF97sOxsi+zca1nPcBe9CeGkz57
Rlh+A13GjHYx6bLRzXcsfJ+KNq6pA5YVmjJ8E66D1O3XkA2MPv+Ro6OBIPgugF0k
xZ4Bnf19jFyoB28bTChNlJ9loFqVIHreK3LmtAJluTJsSAHPopaoVKF+J119CBo+
P8uG5KxvLFCDaLEUeDNUK+6KcT8TUnhgyHX05KpdeWBSPh+NMaTtQJtaGd/GWclV
pL1Ec1cldC7pydmmfqUP/0Eu3qDbhKhfFFB78xQJBhI8JnnEEg0BJn1pvueDw3zq
9C8vGiDzn+pqRHkUImyY3b2TDiO8KjqWgb9aaN1xna7mr/cteXnRJwy9zQHMZnK6
xDVjq1sdjxH6XyKPO/Tu76W/FmW7v/IPbIERvSpZDDPMGVdkL1yOixl453YX2Mmq
Coq5dukYllOmyKYmw9U5PoWiCE//spG3DQ+QelPDrO72x/09ZMdn3lP8eM8fKutN
3R9as0kKYH6XRlRmxm79SPwXdUY121X478xTXVPU2c3pKdI1W7f2hwhzkQ3i+XPT
9Ttt/ssNmEplS1Yv4RcFX3UZc1dRSvIFImPxJa/mHAszDmrymmeJWmXUNChbne5f
nA/pGgEG58Ke3f8BvKnzpxZWbdR/sSMzXMOjbJyeGv7yPzly0eMwo9q5xICpbXqZ
uvwaQh5Oo2hU+Ih+MqWtZ01rKxXt2BKUxxgFBrZ4ag5Nm7BhyAEj27QN3T5s9i83
OTxAZM7DpH/fniNgpHEvMXA9HFNPFIxqztQRAUN5RudJ3SrjWz0YlwC0hUeC8njB
kWLuBH0kb+2+tpyedP2zHO3Skx2PAaOt4fFB0cMoRbu9XPJATwmLhbwjEFfYSkAf
UGDrxUDt7705CoDRFRxgJgQIjtE/Rqyt4ierv9m1hVdvhdM44bJlAdZtI/KmBlsT
jCUf1hWBIW3A2CSK76YRD5KLnc0ftFkwjJyiawpc+h93s2rr+G1Ji94Twg0GGXVZ
IeNKdDH8r0BfenVcEpLveZMrXg0vcov8+B7tHp681xD7vP5zMdBWrTDmuvz6USnd
jpB626V1IPKEfXxsKX8O8gVfAXJMjJ5QMVTTdmX9PTFpWP0mhUbduPW1PUt8vnTB
vkuc/zSLSKCBMombPNefLdYRibmBnRasM1CWE/+501TG/W1VJD5nj3AzYlLsEXvw
qwK16fIdD409LooYe0SpxLl8+BGVmHw3+UqtZBNplrAUNILhqTPsKNq2tMMJFTXW
loiNFLd1aE2krNzA2mfEd4ormCoc9Bt9SteMPC2ZJEIWYIDtxeO4cj+TLj4KbrTY
DsFqg7a6m49lPjgjDmgvy4MDQVpt+HJktQzUUFiuQaEVXQgqtxdbie14DBlMAuno
lVnooD/w+fU2RwjWcY8rLyvEmS0hrUlxi6QOpY1lb0vQ5HRx43tWQcsrnD10EwnX
blqJBtUJywI45tpCCXg4N8m/pbbXOA+Ry786elFBFAsbPIdzS83lmrxvw0ViC5Gu
qf6u500iN50b3O3QjwaWluBAFFRmGNEvkyj4LFF0P9Ytlk38c6UN2/tCT9JBX3cy
0R/jmiQ3Isl+8D7jRAJOkPmRMwKwzz17nWBP7etq+1f1MjdQJh12xQieX/SXfHrC
TM91leWayXoKKeV4hBys+q3NcJMshTjudWpBnBMoVH2drvw4r+wh3/+o9USBJLFF
CykepkiN/VuGLst8iJYiF06b9fss4W7wiMQ75JeJrBWn60byExl66LHZVSNWUvHv
BT6/uXEB2+hJ9BJpZQQdaDlr3m+ZWZttdW77F2fT9I/iKF3IdvNaUgnI1Q3v8B1l
8HKbCJSrLYXiBSyjxQmg+bADK2JwwpUoB3x4Cxgs97of1PXZgYAYvJ59e5B9dsL+
Be4dGY06m9hYnsgxBqRyFg+iZBr/9HRQPBsmix1zIH6muCDLzJLTzzdIb4O21R72
qRAhsEvF6gbHm26MolaAr81Sn6nOGczp+0Z65HmNLbqaxgeBdAOMfsdQGPM509f9
IuNnzqDsWmdjRHIQRz4lVeIGF39HpCgO+IeEGVOQkPRLJ5blxzYbgfIV5SDBD2Fc
CGR2uNmgX2EfYz2Q5HeMmizmMRIzjGNvCeCRZMFUEdwfdMI0Yusk9wyJ3knAVwtc
k4PjaUgLwhNOvhyqyyR/K1CQjZO3RjiM9b6IemVv1h4me8K1PuxSlkCRQdVLi75L
Xrid1M9Cbr1nZwpp6P4sX1Tg/9KV/j0Ovj+RDen+9yJB03h8BMub9fe3ebx+sjnf
lnRxtJeZP8MeDX+lyeYMgDwbxg6vH2ravwJxeSGS8xrS8I+5z+sCY+xJe3ftptqe
usJDm1+0sIe0HNow4JtmswkMriBQpg2QSbjQqcYSvAj/mMDIjoh/ejGIbMLwzeeF
HmN2nMf5NHMXK93hS47BUqWhDe32M47EAk55AFS5SAm1Qytss/JF4Gvf3C7V0O9u
bsnaqrI2qplbag1FiKdFTXHSz4HsnBPO23UpusHT9WJS/XZVs0i+v8SibnoFUHmA
RmiINcFlsMxAGeCtslaoy+Yg7Z0uKITPA6uhituPWQcDRBPdALxJXpq+HB8vLvHr
oYJ5GeL9NwZJbLubsBpw3n2K8mEFd9w3d0A5aimc5z/jG/H+yoNYrRQOqOff7I6C
YZfAR6ZQZqtm1082pk8176Mu71vTWWif2YX58OJCFJK7MDEFtL7YJzh7d0InaIci
KxfiWCwhEoj4P3T/YgthjzPvEAqCYIf2L0meHN8wIrYyqyHRaUa1fY9txQfbWzO5
XVqygIprhgyOrwJklpxSCHri3R+KVe7RydnEMn+0Z/r1e/Xw6ioqA/S8DoTkpaBm
zlxClQ8zcrvVwO9vukdd7Vj44WJo6SmNC5uzQ4Xr/dysKPL7m27yCX9BrWneptP/
zsUh7p+XR4BITVoBVTGPfK/c8LDiGWFMjcIViOUaW0JCOG6hEhPZhe7EkvyAYp2J
wPJBthj+1Clp/MSV+ugVseIEePTScEc+LhqMYlBIjCAOYODo20PuCcxUcbLqwfI4
+/HrCV6IjHNo+80adZIpivLTGdgzOMEqifAhA52tcO1/Wmxym9y5HOrDi119K/pi
OWL2SzvOLQERdHnYSB+kQMiYyaSEOqFIua8jNTawpt4aPDa6j5YpCAl2MQTct16h
jrnKbX0x7gH2cUfJDGjAy+jM7FJ4UDiodPffY3Koxiod+shs6lc/8xUlEJjvFZYq
NoIBrk6UZThdEUU38H8egYcYWwWSRRQA5hqjmVLLYnNMz8s9sptDngODyJxD5ycQ
p4h+/FenULveIBAMFNH0Fu44JNHqDrfszIXPytaToeDKwJQ+Z6kB9s3dPFjROAqx
sVfOfDSArbDmKsWQ0QKEzvzMxcj70Ry3NAGGkI2eUT9lFdx9reWpVznxWmGTuQBP
9JmKhNTTzYOQruM28vZdIXcM9sTlS+aS83Zpg2FdM8ULdPCH9V3YSRRquvqLhWYe
RtlQYTbv3EvCQJeYqFJ2xNSdgG75Y85niZk/A9fiPj172x227Q6k5wAj9VROf/lt
EcXgUCfsBue9mrRSiKZqaWvtQP/CDiJjmroeVZW6axguanrU0TYAyNpcUqv6fR6j
Ho7jLw3mXRbjfJCG77r98M2ZcngWzcFOAZLjrM8o3tqqCnishFeecuWH/OHPKmHe
pa1hvLsMfqH3J5jW+f2GoslY+bMY1Onw4/+OUqfhV9BlQTW6kGjk0scD7CKG4bMs
TPZtKF37SfNg/ebZJq2Hc8ZmGwVqEJsH5pNVe85JK5IlJDBRsIW4DXcqlQF269NT
Xe08R0TRD1AiKXcChNK0epCCmtyXDzo/CD++frVZYV8ceqyr3+EVut0V9rgbdmqz
LvWjdu9jAtM3/u8WGz/qQC+G37LtFHOOZ3HUX2szD0ySGj4gwlpXlnEYkgYUHnxU
fJXgLucXt7vOdHrK+Ltep7GXn7AvLD6Ndpuu3F9jgX2iAskAvvkSDA+dHBUo8Zjx
FPf4Ted2gvR5gBw9mVSYC04DC2CBw8AF6uKv5vR9HLKwMjQTuuY208lgXZoMZoHn
DGfsvOajyMbYliteA/KCp+Li3TL1KA+mdAvFeqb4JoFteZq3DmdJjPa4fH+Eu7LJ
dcdPi4sfx8FwR+1xr5JINrz+exErLWE9h+cu+MQcECkFX5ZK483bnWRJn4zWcJI7
66bMhDaxMkS0OZr3NZS12xIhf+45GH4CevolZOHGazfFHXLfKyAT9IjtZJNPsWz9
xReu0QMabQohVqyR5GHsGnqN6Onnorp8Lzg+brhQZIcUGSFW9h652HBBPXk6hYei
989mmgQIJoxnDl7zVIwhp+bPvSMxiYTR+iuvJoEYCfm07yfIJF6nzXhAQB2+FeSt
FLueLEu6GVzg9R8wuL7CuiZKyjOQz9izau7bA5oBlBbUGFTxbhpiUeGxoo546DRU
AgUPvRoiOFyPa3QlYSgNtDzLxb8AmvFDeRxU4Y7fIiYXwY6bxD/CwN/ZIFMhKDQv
qC0p1yoaWZdLvStF5+5lfrexbeG39CtoiuzXc6K5+LnyXoe+OEmbm9BQTG9uVGn0
LGm1a6VFuXb7VsAScwZF9jpBeMgYA6H3ij5+CiiLlCanh/p+Iqons/5ODi8BAoXo
AwLVKXEQkf23YGt7F8QfXNAp8aUMHBFehcpZ7zwc7v2hsvex0RCeyJhV0AWyibGY
Q/ywuflDeX88vbprcUPkCzospbUansbUA4zC7YuzrCPXplK7EMzwCgHVW5CnecKZ
n+y6XQgg1QkIRqrXLHTZ4976h0SezLaNPu3n/Vs+/YgvItip2GqqIOlDFqc0uYsU
d5M+fpmYxFhbxcRnQrDwi9RSWV3E4iWT6jLl1HjRPsGJbvzAVFkvJOxsIGWPd1p5
Ba8e1wweuQlyOKTJnj7AvoAhBVEs9zvvJ59JeqeoOGa2IFyts4vG4S7NKAu+n0h6
a976HvlthwShFSBBwaNydLQm3CsnDyUVeqhqFTRF7mvRJaDV7uNptgIppLyE3Zz3
HItJdr2GlDT+X22RPnVK6E08Hn+ZIzWOSLrfvXrBA5OuJn3rWMztqCfiYHZUKQv5
7Ow0smOTlCUF+AzuJWKkvc/Zot0Et9dTbur8tFN5iYTWzOJiiLoytlZpZppJfdw6
QKBtB3gprenLQUpnU0uoG4thuAq5iScbk7KtJPAYSyV1rgBx+hyGaRKHoSp6SDv3
LFRd2RuBs6roinXIC3jr3n8IP4WO1jac+20vU2H5iWklNQpIpinlM0hN5W7fjXKk
Z9NuvrHa1+4iM5eLYSbZdmIri9fcFiSSoHuNBv6VaSLoWs5Y8ix79mZUzu8jbQPD
wvLjDV9y/2TuXTJ/Au8gZcZytJP2bt335aZEcRO/vNjUVDrs/skhL7SaDhCIRDIV
Z8zCd1ij8cY1MyKz2zJTM9DzF3QzAqutBHAlyB3FjPUTs2ugdEO6rc8E4jrtJD7S
TviwphxXwcsiTYPLki9mcfokfMlzFEAKKV8cqKsWcaJQpb4elOGH7beDQKProT6m
4E1pHZoTwuR3cFsvPpektj78md/eMhK9G+y/8WOWcFeDbMNpo9ETYyQMHuLXHs0D
YYhbsbqXSPozg7JgAbSxJtt7kiW72ILGXiAFr7aX8KoIP9+uA2toWJxGFxl71RAb
5yWcUUyjrzRH8mCaDSye/w3DiDzA773TpDkZ5Suvb1hb6d5HYp61QJ8NACqCKGrN
oopfY1P8TyylbO4bGKM3be02V3F3ArVEwmYhu9EjIoNAmyGne7QUVhLohgm6pqXu
GBGFY3hugb1xTSVWWfFmhUCJzLghFU07a9s3oc37NXPkyLwuE5VtElD6uGaIEQzv
PgaXUGFAKnwYHTh3QogvTm5pIMQg2ekoyMdYBt9JDLgU6HlI8qHsFsAbk+ld1hDT
2NlYqwD05ODr5DkUD2Rei3OreP2agWDrxtep+a5QI5GVd/MKNLhKZo8G/z7GlsdL
ImikUxftlTnJ8F7c9y31kZElv615WEcvg8PDVkaTDlLRfQ/5Y3azC2vZRziMLm4Q
w+2TnJ5hxSH8UtqRBlm5jfcRH5vq7MNMEGCOEnQaPo2ckGn5CoW7qALpnKSEZYLt
0it/OnEv7HptF5xHwXMvTqcBXmXhsQfso9xvDivm/kXC/hNHA24AVkrserNTPnrQ
VeQ4Pl7Hu1qcF/dilEkmFM2IuxcOwiz4OJeDvZIVHMMXpPVm1gP0V/z9QtZ+gl5c
Gy6reFvkAvxnEgYO8168ebaxp2HHr0G5uofch1wBL3gODeFf88wPwRhM0NoBYmmN
68Y1z+4egHNbRL6HcqNvrQVL2Z0amwoVv4SRcppIqmAo12TvRgw5VCxqShE/5+fx
eFyDwGSK0hJqdDEMCIEHS6J5M/9/t2mZ/N5wgGjwQKHA155hgeMsPIadFgmpuF1u
/Ftj44v+clvcE81I/f/q8KxinMpi64L0fdNY/fR8hqef9gvi1TO4XyyJy3fCytot
pu4pOZd8LnQZXfyfeRqSy2KNB7L1wQixqAPsIjMVaTGPfiWJsA/NvP/O5smUqZYC
ugU7EYPEIgb5lorScNoiYwgkLZvhO7AJr9PBbzj8M+Ij5HIGRMvbaCz7vN2pfUaG
WFT7wWZLXZJJZDSPPOSixo8jvU3LQsgJdUtfoubEo2WMOG2PmcUDYTlv7u8d/S4Y
t/myYcUjxmxQ5QBa1ZcnC0AhC2odOgHn4toVjMWI34BUFOYKYEh+5mQcFuhUzijm
fwadcH1lWjVgtyiBPPn8PDfieRRyaGacW3MFMxbvWccvdmlOwfiUT1MW0EtNuGyb
PhwTSm7BwTgt1CGU8vKQMv5OX5XZOPYV8ds9QCMbKAZndlsaTD/u7/v4AJqghbnx
gOZtL+WjAt3B+maojn8ZtT42+lbgfqqNv7Fv+yPaxAPTbhk9anhfcurqYx+liYHk
axaDzjBktW1nFtUZcvEJhw07O4A52M5koY8Jk7Ctb96T0G9/85gVTOtlshwkP9Ur
bGjZ6iRIr+Co5746Getae+66+7K/XK7hepUhNYLzgck8XOkMUe3QnNHtusRHEeOO
FT6xetfGd2T6MMEQEq08Lm0e3NahBeo7B+aFYKFy/oEvzWjFTi9kcn5fgL5qI/Bj
21hDGph1RouEkpHKDKDMSNwJSSe2juVvEbtiTpxZRrlhxY9tAGinIkK2Uf6p7LId
183hw5jkjxNpS3uB1rDGtbviOACcbhL//2pHIWo7jn4a1wTI+rkcBdfZy2ahEMfj
9fsMcd7PJIyzsHXqFs+12GfC5DvpzbaFMlDX+PX69iflJHNmtnQHdBH8r8f7mu9Z
V4c/ir5tl2akLVdiRT2DuFmC+Fq2MQOC7+70hnMx/qgf+q2mfpCzlukfcC2/Dgwl
jAXvH5ZNV14iAx3kLFfUmnaj9afd9r11Hldrm31jkUezeBnIigayEUA7NxunXo1o
l4xzJpUYU2M7xQ9rgkGS5ExBUdmDzEy7C/9uBCGT6bs5cFOZGT9SL1700FGkz6ik
ysydBJKaanj7PaZ6vM8/UobFaMQLccpGQqJxlLiMAR45llaRBZzb4pcYKKzW6+3T
vRLD1asvut45Dsqb2S9bzm7V/AEwGR59HtJRTDoCa4VKfYnYoY3wUewGzbk7czlA
EwDWo/4LPv85ugwqOThhwylwE0LbAnkR49L45cNIOeCoopZA0RKRWEQTwxASHmjv
C3licCTvBrsehG48nxLwfWFwddVmub2x8foKTR2SNbFNXw3vmZ75fMaEa3bOIQIR
mvf3zAowV5d5cTSIi8Lxopp9I7yJT1PzMyW5+5OyKy6+cU0mFU01vqzZQKfLq+Nx
3jDF3WinPC4/Se0aO2Vmp6BKxU5UwWVh6uVOTkpYl6Tg1ctLIECUYO+g45s1o9y3
8pCgChUmpYBSqU7oYKEH3pfs0vY9Ga2QA7Ki00j0fqjKUANB8KvTEswVtW8boO3c
lFYjCoUxZRkCcOJdAlNUcOsK0xq0FhanIR6kDB6N3OJStUMaRqBnDvHEuQY0Xcn7
2WZdIxs6i24KG6/fohGm7cMWQ0lgqz9vXIk+CwR4jgOdV3YdFD3oo5lkSQHNnsnR
C44deUlfFcMgeW2rKvyYjKScbi1dwchAF9Pyek+MhTW1ckOPJ59kB46hYTzJvXB9
ad+DL/pWwAXg21YGsS2QsGiZRb91einsV+lzjzO+c9+4Qpy15XBoT712n6yI/8LB
wcZC7LnVKsOg0zEagS+UumKLIAzaUURf8aZWBlKn0x2HVRlVe3dGYQztQ/qLC55N
f0UmZ56rXHUk9noHWYyLxwp2ksW1TB6kSvB+7On4d2r9DEAnzupkGg6rcA2irQEu
sb4LW/dCXw+qM3sW0bZH3hYerVbm9/Rl9sNRPxREPzq0dTcyq6oGwBP6mkHC7J0V
FMrEAaENU6hW/9BuS+nnHfv6SjL4cCizSyG9dRFPf33hg9/zwR/K/IzyZnPPp0pm
HAVxathQ043gtzET+fip13nhJrfEX7Jc28x+ehqDrfdYw0CNrCmh8gHXD5TIoNem
WC7msYiIgDxz60qOOnVDuVqpGBlpbKuC2MAw1R+MkHwy3NhuyzmRxLJUpiRLXht0
KRQacRFy9ScxUi5xf6Jfjh3UUBUBe4x8NFIccvMHp7xJYQhOJslfumVm55RLaXKX
52gTpbBQLADhSC1buVTBDiXjElUaOcpn21BONTOAu3vbyVzx7MU5Ow+GECb4cSYy
ybeNdvofP4umAWRUP66a/NrJHpYq9R/NGcY6i2tj8Ne/uejVgOxzmpMWXI0f7Qzp
5C5wciyU5uaYzIsX3lX2yUkH2pMGe7p/2huBlXhiDXIKQ5b2pZrF4Ohu9XE3BRXn
ZgHx06Shxh3jNlLg+85RxpHWlQaLhKZ7L+1tPCL5ddvtwwXW9scZEH28lAz0YuyB
F0uLvDeTZtqpyPDJ1Bgno7wJp5mFGWTplviGyHey6JcP8678SNk7L5elNgAfFI0+
xOtsoSaBX6PyFbNLWnimDzlQI/xX+n2ZWsvFlOw8W0mmEk5rRSi2Z03QsJsrJ3gE
vMezqPz7dBUkknOUlWrx2GT0nluldDQY5WM01FFE71Q16W0ptRSqmQ/oo9R3LKkq
UlK8Dy2faFtlLR56H9Ss6mgfwiWHTpxqbeznjLC5nqyhjydPJ4IiQ9+o52fo4P71
Y1gt2WAhSNErRaHXU2nRj517Z4Mo55kFXwrtMl/pqUQBACeFQSQdoDVwavIPCefo
z6JpxxtLY7puETODt7cyIG/m5DdEaNs0gTLPEWIWt0yT6bVpr2+pEFDk0g+eulGf
jQ3nVT3xiohoP2viApU52C4lgWZMTjqgWOpV4qO1n3je1T1u/OwtJvrxa4w/W9cG
hYpvy1MB6shLwgnKX4h8q17iFHIfwQuKK5ENwKav55YH6C8Yq5xnWDfMcrR/8e9Y
8zw3CJ1hRptfy9Pm2jTMqOgEVtkJeYZlqiwfE6qWw+9JVLAorDq45zVRtE3C9dHi
XrT7t2bkhddVonb5lqK+ZX3HBa5tVSiBdlTpFTu/agPZn02bIDZgu5TAOSO7F8qq
5SRlLvJJ1PU64I062WiiRgG4MKmfygNSjBZKXcYMl3iC+yg4ic5jv0dEQF/kv68I
06/kzyhJyCNi96HlV/kBoSjwAzRG6KYFc73MYKcFvj6NB5GcqTj715T/iEMBwMHl
XSIkvg+tZ/0MxvFUD6S5XfIiyGdgtaW8H0/qsgBEKFmYo/qVCNqGgN2JxIQB3Qi/
DlZSIwYErxlf1UBAq6m1G6234EJfwbQaNVc/KA+7oFZt6EvaV5BQKN3Z2V0yQDhT
+30qSOePGhDpbbXHw44nhlKG95QGMWeOjwR7TLb5WE3M8v9vPz3J4F17+H607NdR
IjhXO4r5jVixC+b9FW+lNzzTEKaf6KjtVH6s/HosyS9emvQnlA4muI4qkin5KAmy
px9Do3tciJ9YmWE0HdtxD2+kDoRILGbc06cnsR1LWBswa9rt+jSplBXrnz7Yr50d
tn/viqhHabTh34euHl+yCxKW0k8qSFB+6lIaYoxOtHdZrqflyKvu7ey18bNUh2kE
C7qO8NJ0gHldFQA6ruJLcyAJoJL9PFDYqNfp63di5yVhX96UdLluz8vuN5YzAp0K
5QA1p9HIXW3CTQMUC+gckZtBvnllnrX0J13ismv40anww6JeLcFajviKpqVaWrB6
T1GQRAnscKH7CrrXXqnk1xDL3sWb2l+lpvl0IIr7Rs2WQQ0rhDHP3sAuvWnuckp8
SMmu4ExNy5UnS/EaWcrU6HrGOvPztoJbrh1ZOA1QsJTEFUN0pBRmxnScvxSeR/cr
NRd5QnXpUCw2jYffDp/phO7OUlczQM/t/mN0z8sS20tyMH/29Q/3OnCU9hAEThMx
chZbV4ZyYPF19x0ciDkTB8EfFNhEJQaJjZ8Q9HEd/+qbCoofbxWM5lh7xl1p/1Jy
nt/d5Mzq/Vji1UXRBhrirBzuTznESnIs0BO9ZnSIbRc6wsoFPV0z6zUQsjH5b9DR
hocTtYNFM5ZscaUcDMXt/9NhfAwOQfQJFsPico6VKIDhHy0ucctcBRm9i/PoSB/q
8Rq47rtiIZM0w5rhj2Eg5siwScAngjbTFcIDWa1jMpZXyGC2ZLW0yfQZDX3lE2kg
yblh+cQpjI3rKxvHLTfRrf4PRWqvS7fJTSfl7+w7jBEwBybQYKtQRUbkLdHBuXwA
vqU0ZVq9s+3ru18ZJnkg+h35csXNAbTCV35rFhYxOS6VC+2dW61UWgZy+1dXdzHB
60vPM0W0tJ+mqPWv94zI83TA0ecuTWYgUhaMapu56s1WkeiT+w5WUx3u6e6ag3wD
4MgvUgY8SJtvV/V6XjXrfqP8ltI6kxGR+mzUAm8CEUK4ANRuhSKDvZembxt+Ia7K
B7KE309cbVKy8LQxYsLkDY4YaVqxrkrNibq7pD4D1hmn6OBIykWZ18PWu7nacRZd
b6uwheHbUWcDNwITTNcno2GfIqAuNLi9EmsG6VSFrqyxvOKwLg8CmuENZiZlDiX2
rYCKMk+F+9SekVOa2TpshawVE8JTJ8Ol4AMxWXV0uwGL5RtWgXpCGwPaJA8lbfap
SaX4zGwgoOeb1PE7XoljIWCeTKsLzAzFWeWUiXEdujQP3WjHjq5CUMhYsEim/2we
xzIzl/PNYtjYkrS87qlyr6W0xTvDcDRRPfk7bcWqQDQ9TnL2pSyAv+5eFkFDoRb0
9rmFywUE9VVbEculq/5x0pgbHooxJtNHtUvnF+1Zg0BZ7EZdze7xv0J4ULUxCMHt
MJTbRtRhr6RjFZ3gc0qckqDp+zEp/WeWCv9LEtc4fjruFbdoU2MJ9NHCGkJiDw3B
0c8OBf1Uo4c56Jnjk+9+tPVuEKJRxkQyhQUwlRiAkOQt4rOcceLLzOZ+ENmVovCp
8Leb7cIqoOvEgQCcEuu/cM4J/9wokB0Z2RbUoTD7DtRa9RO9dHV9hQ9suEqA02c7
Jujd0kJlEHHL5h0qKvfTPiYjWZxQZLXCswRXjAC49qgjDdRqqHv9UG75bZpvNhcR
/qlDHVlStknA+d9XKixwa2DbDcS2zvw794L4SI4x45mKx1mlkEd2lkAQwKYtEdEf
8ACvRk8n3zPix/cX/5HDBrMfpjlloJ5fxfLkPWvoaFIMnUm3f+p29kKEu7Es/Z4H
j/6bd4ti3PvgjzXuyW3tFZCfkhxMPFXrVLAmmY/rNEUq/9/DcFGmXfr+49KRNHOA
hLjY1lJdAO5stkwNSQz1w321CFGS+g4PIGbcN0pcdhF5JYNRHO8jPB4sL7InN5xP
9+M2eIBf5FdG2UtWNCXFuJYE8kvRInuWEVmVvXM9JEL0km1q2mHxHRwQY1deZ0O+
HuSu1XdzLfGYh58m783afGyF8t9zYDpxvkIsZ4mZfhJUGVN+h4YpItsJZScfkCW0
6Fdv02OqwnndO+buyswW+D8p0dyTPleKTQpnEKUBHcxPoA8rkyqxLLIFrxvC6S7K
TAOL8Hl2gzSdLDXsFCEIeuxfrJfz5q41+C8z7p9/+1Zu8To9w4gwEMu6NGIdz5mc
DmXfi0blHS3VvMMSdFX/wTelj3zJHGhiAHLjM3SZJ56H21HBKAEKpBvqtX+UJz4a
UcNk/3i9zOvJHU6vK0gPCXIhBd3E4IcGTMhoduDmVZBhO0T09xq8B+GXbCg5nDLL
Z36m+1ybR0zaNo5ANSz3QYE6MqPZyXPb6w44QO+SKcDklVYgegIpI4SsqkSTjqnF
AQ6FaFaRgT2LDg/8YMoFYrBJdGKt96dpFp10fxfBx2D0UBuCMuDb122lSM7408cV
e/iEBqooZBUFLLcG1euE7UN6RVfv0bvuT5IbvM3/kDIziHbVmiMCnVo+CPJsalS+
gQi/02VqSk6Hj4nm9i7ovGMem2hTN4KRvxjqWVUJCuu0fiQHp6ACSzOWotfzzQ7Z
4k0fEqYd42McGG8rUDOhwtKFcgM+rFnn/CG19yQFZSrn8mKpY1okkyRa5S2UDRfY
0mMDWnZsAa7U4VpP261CZKu/NvhPtwekj/SAUnArOOBMKZ2PpCl2o/i/TNt7bfNL
8toyNRuPIZwn46enP8sD1g/6LkVow61J8MLrL+BkKQP8/itN55Dlp/REtP+XEb+0
2g12w1dXvlr1huDJBfpzoFmdmVbxdPuR8S0uVP/rFf0ZenyEpi0s5ME2euUxNfAF
EiZNaaSzPkLs8rB5xMTteobdoexkwSNgqXbVM8g5nbjWOvNHSWJSR+GnecAauvJ+
Euo2WHfUz8Imo8Rs9zFdn5frow/lZg+zyT6isZ9w4D/pPQuLEeF5xVDjR85jR6Wj
VxoqSb6DvT7vacX/grlFnsDiUzUR2qaM7nEv0AMaUGnVVCVBtSsOCpS41B6NBVfL
PsYeWU5oXn1SNFuGFFYBSofvjJ6tlFj0clycVSMO4nskEm063xIVDqIgZdMaHvl8
LS6bVAkUqRtkSwyHmcu2V7Q2FsZYL4GfCwr08KWQ/2gdzVEjreOc5ZZzTxLtDFFP
XfgcRbIB/y33DY1p+l7ulLP1V0ZlHHzd+x+xBSdYhoNnzwu0nWGsezHn42pb8rMn
pOdfhsEr+Wknxc3ecXF1z1Z0GzbU8RHBb63JUr9H/CzV/+481Dv1MELV2dFGW8i1
nSca62CvgQGygz4R1zG9uyPZ41pZ+NxigpuJ1p3H8/0YAFf8svggkXVI+S4zaufU
5ZiECkJpayZtzkkYfwJBrmtAgozmO7Bj3AGxehhFZN2gVDUlGl9W7DeGjdcTzT8W
yB5cP0eAPkS/de6RoDh50XflDLhL6zI4ybm/E1npLTB9v1dp4mKSnM0jG5UVw/2E
7+dM1hhit5tT2kYDokSkPs2LTcUM0eOoUX0bN5QgGugO6du+azZKeHrRoCTrmutS
KDoxi286w5cv7VM1NEQJyPh7WD51efOk5xvrMMVQb4nxd5A520eqV2ZCb+4h+9gE
SCUvve2ja89gBhB3OwnEEuprhc8pv9ZztZBm8SvOEdcBM5H93iAuGDci8swC6IyL
sbgcmZwAvKg7cedklVgID6O2sD2IB/SwyZcIrP40OdCuv9oPheivnd95eSVGXI8F
509t84e1dOOJ/4b6kzRaFaCNrz8DIZpVgTVsv1To76IGEShiqPV/Zha1ESGzXSZ3
xdEggf6drk4Ly97z7cacYmGMCN8Itn2U6/jd/Id+fLC5R5t6aRq1PV9oKcL7x6fC
ER5+bgJOAlGXimS9BzR/HbKSUBJZFKo1L3M9dGhmXeIOtLn4K+VC/ovB9NPiTQzz
abojRKeHxqvWhDj0fn41IYnf2ezH0X6SoZnVxOz2QxXGuHzKdad3kczPtMFY4TeG
KccI+Q2WOb2NQp9TJaS3YbHqwNxOjpbdSfYdWWyXAq0PucJXAf8WzfE/qa6gyUK1
/JIYz6m2uWvRnfpIzzeqbjGvOEb+mjpdbQFfbj59fEdiS9n33iW+vtggL8t+2CVe
uNrDwdDB/E23SQeuX73NTFR2jpjQWlbDs6NEiw+RXMMIGijv7FLAcswSued5rBzw
3RAbWXFuoYq64mqXh0XZ3nXj/Nu9x+auCOnAq8yQsmrzeWMcWCOa0OQu87kZ7TOm
SMZNQpYqSTjkc8W3Go3eVbDdmpT6rKwjIAxdaq5iqzyUtvKmAlqQl0DzsnsSNHa0
XA2ruMbzZBawXfWQPPpE7slCsEgak2MOl9bi2J9Jd+uswKUy8paafu7EknPs7XwT
kTBJaWGSgT6z2M8OpTVm2ojpz4bh8ZlHo0+pf2odbU51CNXtG1ecAGw6lNRFnT2E
3pyF9rbYsRis1i6OjMYb7eWeypHQRnbzeasPmG3Q4zp6i8iNZfR5w4oeHBLbho8c
1IEc/UmuU35zkRVLmgzOEvLQAZ8elYw1g6+5VLZuFKDRf2BBBESpJ4okqQbSwhfi
I3V0RDWVYqAryK8IuC0UVAmjR1biP7D2UHWk4JudMXf1D4Jej5TxqEPX+ViRyT/M
FNFa2oU24WDwFeUJb4Db5rZ6VMhjWDLywA4Tt33QWG0qjAaHNialvfm6SrwXjokA
yrSkgI6FgbsdwZdn53FdKqL9GfsNaQHs7N1X+KytoMDepXIkYdthBApTyW53n9hp
1hMvygJ521aOQNBJpz+wU1P6NVZRRypJ0sPtj7mBkxYdd424V5Gwwu0HVso2TAk+
TxUcNOZNwF0yE/hW+b2LIgf03OQSJKoN+Gg1mZxn8bmJvqBcRwxwk5Lh1QN1z5zG
PQsbBY+eEErftJwZAIqdkycCQpXsb3p3/3jPfJadVMMnGMlqozQesfzmF+xwIy7a
LYD/H9WREy3Y//gjKEN+OEDEhEIZG0TduKa0Ku9ttYAwDB/IHxHAG12IxPoxr3GA
2fO5yEE3b6bl33WH3AOXqaUc/0LElwNBA8FZe/YnQhu0/a5abVutIpTYOfE2khmt
FtIO5fNHDvb8Gj+6lPhCbrW+kdu91yEFTtXnQWo7BEl+w2xYDcVQTzmclZI2dmMx
7f5gvcRqY98f7mPahj3mohmsnMRMvQxy5Rmtr6cJKhW5rbAiVR96XC3kfHy+Q09i
8mf01gwqvm4xZpLgkFlXdMNlYoiZzORnB+IViDq2YjS8S9jA8cZEfviOHjg5E8R1
cD8LCslEGIMfzFdd6JS9fKV5koVsQzefU7vMDWdiHyYQB2K4zDTLCCecI2ujCaNu
wKq5itmrzONKJR9wXQGXJsNQ5sbYLbn0ZJdwsJqOdjpJkXscNWjKzJwrf5rnBqND
3scQ0scEn6o1EXSB/Xs/a/3Yvb7BtQT+rjOJbaTQMt7+ojmos03A4BJnIeQ0nANJ
Bac//pTkI3MkrJwA+MGqVvxzTTwQJ8nC7d75HD713gIrGzBHVht/K7oAF1kaXuON
/I/hYfnCpZM+tSUr3iFlmAyHuieEqL56TnUfNPoF99IoDtGtmxEktKWJ/6rqu+IQ
Sk5MrJcFCQTyuRaffIUozL/Yg5MbyVHJBucEpm2Tz5o/cCWBVjV6Y9h0swKaJKZW
m0LxicKQw4gDEVXTE4G07aZwKlRfmDWR5jM56MIOUS3buupIIa8srIIu8vNXWl3f
sgOxGBnZld50pbck/L42W+9gKatBaIIY1sWHFOQdVtfgObHsoncE0MmfbXeP8+xf
3BONUqj5FvtO6dbQD1Gbo8oytC+yaTCwu9kVqEoZraYYiA2gxU167rf/6lbv/4I4
n8gzRC4d4O8JLTNCIiWa17FIQjlKgB7RgsTmneZvdvM8WysjltRX34iBISYaNx7G
Ty5sKAvGBgvD5ncfJD8xCtlzh1sbYQ85TI0ocyS32tpb1blR4KCit58f4kmWqdng
OLh6oOHDK6RziedlRtFo1lX3VWsHGaaS6dwFmh/8HmNNtGaxGrozFJphuQWux6Sf
CgballK0ZCrcYO2Y4HbstwEPb/sodTqSrBhotePFBVGcRzrwh1Jvb+VEYuukDSEZ
fyNnl+X+T6ftfAZcktPuYs+T7r6eyOuxYNHm9hQMNj32As/e0qZUwYlxPeO/wRR5
P+jGNd4Gt0JIInAZh3qV2AiHDBW10DbUkoGiyK65dSS65fHFxA5OYNnzXNdvCICA
wS3iVRqz8yu4tTWJy41FIeyDj44KYceZWLSZl3P2MCyzopZwKU/lH/un/utB3IFy
6jPuv+IsZy6OpeM1g9eokC8NKT69kyjsZCVvAVMczkIa0bivpY/FM9nf8tNfziVJ
n1o4ya+kFOZf/WxprQEqM6ORO5irF5Sbvybvw5j5I4KmUP9rD97TJs1st1oRKRLj
4jO8JLpCJgUOFXbFcFmlXU+L79Y1t9KQH48VLXDYLPz+JEAYyW6iyHzlUQxnMYqA
d6B91sHjWsTH9rXNPluXprRnakHNp3x8M/iuQPduqohpBmp4QDaEnL56DXWrQ7XU
+/06RsgN1OQ+5WcTFrzEtyW3qMNusFyQ/3H6IpkJ1zuKzoPdGYnmnjCwoOCGXZYe
xZSRMRkJaOTJ2nHbcwtgyltWe4pI450uk2gQWhKDCb/qlhQNACWzy6BEp/NWuGcB
ejgCHofjvM+PHN4iwICUO2IV9lGExg27JB7xOeY6r47bni855Vf5t0UMOuY+InXZ
saglDYcgqrjz9oq8wJ/QNv2yEXMG8Amo8E8sdYDvub7J2ci/WuJNNJ+/xOAqW1P/
jrEiVkHOjEqzEjE5mgev96YAVNRQ9O/fQDNInPazTIurch9y1n4TRqP+qyBUDlmp
JzHFyAolYPgeePr7jNF/r+y+41uxLmbYNBmEBBoXGYWAoQ7UiJZt9yub9rOcVZl+
nZ5JXoIw6YJSJK3RWw5OkUJn8iP9I+nHml+cPe4G74QHqU0ftm9vFGQmdK8KFriH
fgTXit8kk9BTXvraxJ0al2fNfmyCugaaCfKYHmiLmgB30trlezBDQHz7NdemCvc2
xNhsHGJiXgQZpq4HFOGhdurfuJvvPZEFHX6MP+/u9i2LMH1BdRS0l9+bzMAIcRbf
HIP6MhZlwvPIzbcDTsP124nNan235qH5cxSwgvuchfkjQWzhujW+P3zT8JLtJBno
gx87fMKnGDFDvpMA5AaEu6mhzgNvKuEURbT6QKgv9QpU900v6ipLTgkkTEqdUfQZ
yUZhxLiywTuuOjHAT2ZO7867f1iQvhXKx/YCHo+iNMbfhdfSW+3mp10C7zLYYCKq
8GFardrqu9+2Ts/zKArlw8D01zEoBH4Y4jdIV9AacXgBkO7Xh8RK7mAJxA3ebp9V
MSSGa44aSr6kLqgWVrriAi/2Y7lgobecqDtMcWWfFzNyl7Iql4Ej3hlpJmaTsNQc
RvD6KyjYf17lToe0rpZ9YxGyOatmF4L3JQV9j203MLVgrYI0LZAaxKSYgzX8If4K
2YaIiHI6U7ipwR/j53fUBzQgtY1/zLd+UU/AW7hdL5gpFvfZVfpPPgsPIq6qYAmv
qR/dO6Pwt+aEdtx8E1sLekudP/tvlnX4WbZV78lu8YlQ/lsWkQUD/gKDdWJyWd9J
nFD9JqMEq/NlCV613+AjheK31fJnipUlLHTHWmFAAQF8egnFBGbn2NQM31D2VuuY
jR7UHdpvfg/rUI7sGIYZWIzs8VttiQVoZta3zhmn+MjlJjBAd/p0dPXaim1cSoIT
dl6bUfhjE0D7Tumr5lKCaVRse4laOSVFFoAzYG6bgCr3uohqm6nufnztohuqxrc7
5JXT/SnMi1Q6Si16wvCMy6UQZ+tzgZbp36jCcVWzssWN8F5S+5sBKzz31DWgmKvu
XAzXhcIrboWwS/hTzC9rdOxC7gh8v6SYk++iCTF0c90HW0H+fO5Jiq8ujmI9smb5
jQqJ1lqMDmOZcvvqcxh4/c00BqfL6/y4jWiwRpXTvybrFkUgQiSJUPBB2MRhqlNs
M5Yl8Xrvmpl7QUjruBQoGX/VliRjyIUT3w9X4ysCsteyiUnNCUCji/V1MFSJe3QK
vZSYhdJuDr4TkfGTG++R34UWu+vidswjDTOp0Ijsilw35dVa97+wp2bg0ji2NZPE
ozJ0nev5Jcn87tEcPJdxqlqW4HvXJeVUFaxKDtI/V0x2J/fxtCent88hLyptlUix
CHPa78iks991qusBGEgavTK4LqRvbvYQdIIiH5MXRv5FJfYL4A5L2VO9tG+p73Cg
ubbghVin1kNQA/eyyao4Oh0YVW5oswsCKGRwmqS8DJjGfbHdXZFpm5Ts/L9hXFl4
gXHZPY+te+tLuCis+WOAClEkk9nwCaH3yk7fwMl28rCH14o4dG+RsR+5aGsCKCRE
Vkfwmsc3lSYuFISKQ4VtJi5MhIDV1N6ramymIcjbhEYXxMtrtWRKA3CeCp4PzrD5
H6MGCX13U4mYRXbAmstiok9ax34xKKH1YVPtkYbNnmIrpyP+rx46tD65MQAZ0/Pi
CGLwYiWv4cghandF+0Kf+kYJF0e43pvRVmoDdR38oBJGL4OaTyn/OP9bSI1gJqj6
ij0cRbBdLZmsCrnbYsWX+jjdoq0wYQUrFWvrkqw3/iGxcoLjD6Dn8GP9/wNLEQLF
ylzLWP7PQFd+YZKUq0ao1e/R/6NYfYOKUktiThguZ0JChaRL+nbjso2TdtFHLbxp
PhJeOhpstpVLxJCdmUYfbrixMXhdo3T5Qe/4nl9RZ+BZvg1OjTSAo7QnyjNFh34a
AvaGqBnDdYswPFETj3IlcXuWlYy8HlNW+8huiqfZ/pJNT8k1iHKnT20Uud9MfDAa
gdpMSyrwiqDN5PbW7a/NYw9EeBWZix5GZ8va8CH06Ksp43qVJmASW+iAoKJJKQw8
6IZnxWszUsVQSpCX0/HEVhYQ4Rxyu0HU1X0ZzS+GApG3/R9hzv6qZVPJ6oDc/7sR
imaRGbanubPHyq91VOlcc4Eba1dr2OHBaLY0fehNtPXa1SGBRl1gDJ/rWSsbsxcq
MkJ8Bo8hcD0TsmtIa3gn3IeOhhspjCX2JWoaKPVV0fXgii4wtTEu4J8ZyTOb6AkU
T25KvX5cgN8qhIeHOvBpKpFgB6k3UbG0L6S/z48L6QEd5T7AVruZu+IQYNCEL7Ck
Io4NYp3imvMqGkq+mOU7NZrE7Cfn0PsPuMIe9bUOWcOMZvQam5GdWf+Ujzt/9vbj
5L3VFUiQuyU3KlY2fM2lrLDmCiOIUE6tw5Slu/Sgp47qyWyefgn6p42l5daLx1de
XZYXrNDlYa5wszXqZIklzOfvskRU9q9/YzZ7B14Oy2Rt1BfBd8HdRvLVRDYUwFve
GXcJhLvSBHNS6es9GxtEmw2odZxY7WDeh6+971hiaQyX0jeQQjwxaIWBNERFIwFc
KEu8le0SVvsj/cQGo5MBqjGA2gHd4HVH0IWDcnTICt1xv8RZBO6lqXx1oVK9YtsT
7r9Jdeg6I88/dRwJiaSizRBYK8Xc1K63ERDEIf4MEhBKoo7CT3kHXRoZRAaZeOOO
10KDrs6GNB4IzhW33DZvekIfdyBuS7J1bOc4I3IDX06lDOhJSdgEtCCulJ6GLu+e
NuGwG9/02H2sOjXYH3KyF8S+6C/SiTM+lEbobRapbW7DQIaLTM3ZDIqnvz4H400b
59dkROyiH80WAWs14hvui1jdvelVft/gAVXKAmNmGXLKkQMcKpwRwTw0izQk2G+2
1PcmHoL5TK3bVj45h59+LentEGGgi+nDNqrKwNU0MMMeUST1j9JkIS92doTDa7xY
1fqqWU7Fg3vF7hgXZvMUUbx1OI2M5b9ZZbsWjW0y+3pRjBnA8Xmev1LyTj0hvSHN
mRj87Q5xzoKrBt+Wm3CdSeUulT6CNGbfCc4km3gkC3Ou+yGleyEBZFNV8EstD/Xn
LCVd7GTGF5NnFhphvuJQnm3gFOmNWshfN3cghWcPU0aE1bBSzebUQ+OQIwtFwWhQ
kHuXHmoYVpwLU0pmR/PjNoDkYB9KuFHra0ZIJHXeR786upVWsl+v5NHW+H6/Vmqo
tuDRZO+U8CjlYiDEkxc8C+C4pAbqF8k55kuCCY695d9RETIpZn2rwNGXkFqga3tK
G0Q25iIqJdalhyJW9zgzYqIbQC1Gu/zUZU9Bn4ig942VyoaecO2n9mj4yrwemSLh
GDBfx4NHLlqmKYVNgcEk6qoBpD6fng2v7NJSCo/vwWnpfKNFXNbuoVoyhtwcWulj
aeWSefZY3xVeDwcr6DE6+kwPtrSRq/6DjTmhq1EiT/AK0IA0Bwg7UoKfsH7b+Kph
Qi4t8zWfoYK856FPcSmxrru7N0hKWIkHTR/gVfwLcZKW+Cjm7TouQ17QJfwbWAl/
08tUFBcHOvvq/XWXQN0rEa4NsYsV0IEtvNT04S7uxWcDN7NQclKstrLgt9K3gaUH
iWJUhTLDt2Cyq321JjEvItnQtQlQ5hhgr4iZSeNagzHBa9tpFTHdTjT8OV6kzPPQ
0C8VW+KTVA+iQONM5gyge0+7R1WI1ku+L+4c/EasL6QJD0moG5lZCOaLiGOQsIwq
+Qlq0R1SqN4PtKRdDgltPlQNZ/wTDHkdKXX8P2iRnTrDvT+48WeAHAQsjFIxIUfO
QUkmrV0MCAzge5sKTl9dt+tg288Un/3TuAgL+2+l4CTnMDvZqoXXIEbdTXL6IfjY
SPgx8Xy/ns8zPEf0B1wUt1GqXMCxYV5E9b7cGZXmzcVoNnvhw0wFzI/3MHDpHmxK
qmNnaf6aOmwTu0/SPJZVZO4UfTCv8L/MZTwi2RypqrOc2wdRpY62mwzpVT3LAYBl
+gttXXQXrRAXk9XU2Xnf1nC1wma/iN9Z2Gf7vsfFaeEYCMvt1YkoJSx2Rs4U3QCM
HzRfr94Pv2faqlb3eLHL5zPVKHdykTIHv1bFDyA6JBKYkonTGktKGoTHs02hFzeW
V8xQXi1hNIR2TIr36OlRUvrU2dafUQ6iuQvbzIgVj5WS3sbNhoDysLNT7bCJOzVW
7qI4IdEhw3RhTd2tFDdyusRChMSzA7JoFEXlGvjKELfZ3FgzJgfmj+nKQwXEr1eV
AX/RissBweuw107+PjW74pj6FKXtaylEfYqfoCfNJaYHvj1+NBuEIYg+z7GpV+cy
Py3b+xcDkDROwJms820A4hkinH6suZ+ZXbofsp2wd+k4obeUdZWeTKCuKxYoABn1
WP9aFG8+LO/IN3SA36pux/1pYUfodEhe+1a2dXaGfIZqugW8d0+jznlMKotKWuC+
KLcIpqhSewqYxYVUsyfHzuHNPPIt96YFYnAfBFpmfbiLLcgL35gEDDuJFw/n3Qgb
tqPmI2JM9M9E2jqEVcLcwXTToOo2+Vw/qdDlF+QBgS1yzxMQdUx0udKaTo3ISf9n
ClMPoZucaPtaDZNKCjhCyvDAYqphNtzhjbAT6ihlAE8GFreThNSjf3DYgEMlkBl4
E+SQQk2ILt6Hmca83ZipmJk5+u/uPDCqMHUcbMSazaDe0hw7dS6JeciNr7zNo0Wj
e0VjgMmZZY6ssABA1mHVZ5x0aC9nE5WJ5Hcrs9xHqflGw5NAHmGaiqWrjq8BbT9G
l3mzMcZih1he6vkp61eYkc8uJmEEgIgvw9LsMzok1C0rckBDxz1jtSn2aQL8JDyZ
PE8ecPnwY2gQWE97xrNO+5qN+8Fb57066p5VSMUC/v4j6MISPrwV1TTqK/pOC9t8
rh/sfYBxeDlR/3TPCwvYoqDcnKq3w7AEmSY9OIMWwhscRR+CUC79FImpFi7lpGrr
7Rx7wrgTlmGdC8Ihwkx8mA8Cy9eGrJJI8v7nSiCI3numdLLoN2gewaGCnG0iZDWq
HDZgGjQ5JdLsCNe+4qWw9UKPOJeR7EGg0jtfFrEwpl+gaO3YWW8MlJyVXz8BUEzT
xAKFTeuaD1K6+SC2+g9kFiyHIZtdtqo5IFt1eEI9oKr/SjiXujD5PADFUTb4p1Ul
Q25fWl968QDV0mnXoHzigaUvGLF9yOJRNrcjgaIp+z42lSR0WeciV5oWi9bgn83n
1AulSsHXPjAa2NovsCXYlRbr/1J+Uu4sJjVaghe20qbj9iKnAVwhfA+ksV1W3pn8
I/kcKyBLenm4yMNh91BHCsqi3eeRJ5YjCvs9DH+n3FaUFuruNs6AI4uZ9Acjxtxf
oVCvvB2BTEtmsIK3t25/kGRS0UZK32vvyIpeB5K14TwlrFR9bo4e8pF7Sk8yMm3H
+G6aXX/Lw5dQHv7Ymg6Z8WA2AhUvmPuc+yfYa4RNDIi+7+h7+AOFJ6SsFrB5PbHx
w8mtZmqfo1ZUhleC6hfoF60v6jLsUtAmeSjkQ8sjTzQinPzAjxDMCmAvvfEWKK/w
qkaFZU1Ois5nGJKkBWP6s+nST6zEABvEtrOn8A2YVPhvCRyYno0giYiPg7SHtWje
R78+un78O0Fx6PAmTL+HYOnGShdDI03FyL2l2jXF5kaLJ+ASKj6mkunkdxwhdtz5
13uMWXnV0TzF0qfVAFPoUxdXL80BMBm/dIRhNwZ7Xb8yS6mNFUYm/AusmKh31s72
XiKtJ2xJXs73bDxe97Yb0OMvQ024vtwEvakLHBQpVu0+2+smaru6vW2syhLzvTF+
tCPFiUUzASGShlCtJAJl1cvALPV7RctMlMkYNh6IiiHxCM3uH60bxIweoqiRxCW9
K89+k83YsF7QOPW9UxyF3NHeQBHwu/rnUmywV9MOanBPgzZLRJVNBMHQin3Xd5GG
S1m/HnPtFxMgajHRZVjWCIf+BprPRpj8ACAL7bLw4qqfnjI8hxcizcMsAJh/zWkW
59s+UPiHdx4l1ejpLI3Grwag4V0YVOO52XPaRRrkmHeL2t8MHmgwEUoIhIPN/OLC
3K4Na5gecAztcI5UruHqt7PA0mVqPtIffHJml7tPAIVZTttMWvXdqFHtMl55pCuE
jrPhmAtyUYEtvzCp/Ny2TFebWuZVJClpaD63nX32SuIYvFcPElwPavNotrilk9Kg
fvBASiE6NZUQ19uxZjvKQUzDf/7Ej7AKK+s6b2MV4wUDq8su/FD3CYMLIgIJDRhl
086k9Ulc92yf2jX0ehmTwswgL5ii0IglX5PqPRwIJ3iAa6u0UyvI2ESiKccHMiQy
ABwtVnC+6mb9I7c/pj4xOS2CSnItMn0ezTy1L9YOcL+zSadVsvCriG+CbpFfDlBG
+QzHlwuVZJgPQjsStVw8zEJKxIWT0ATPWpj3g0t9XCi6hGg7JcR8S7lesRtgJJbW
IBsvjzEVXDwLwWiXOQ5hyGtt13IkhMu2UAMI7iW9hXnfxL0Fo133b73oqzxDYVx/
X5khj0S/pFkq1DlaYWZ9DcOGXsGTu5zwEj5IqWmamNMRZIvdJq2c9LZMvw6hKAuV
g6gyuoPwD+n4ft6M5A6RoTYdxZJSkOeQzBmKipT1neWXtcGdiFxVCpBNMmZEqf+j
9KEL11k+QXWP3C4BLI1nPHyMJ/0XkTGg/ivLrJiax7rD/DQn3ZLJVWKJhTpu9obk
ffyovmvTAiuJrkwXZVrxl6C/pvI9SLM20mddJrWbFIcuuz1NIyxQFDP/y4tdQgUL
xklTmA5FvKFStjrzNSbFx3UkWeI0zL1EReFdXek+iL5UIq8SE+pxyeY2mlgbWDtA
edz8DBycAiZhPu49+ULobmWGe8kX4RPsJVCv3O2YvnrtJ6n1naqKBc/1mrZHep2B
9eGFo1qBStDrhoMBI3qSThYhe/oqJRVSqZ9HKo81y8FJo/sEMmAd6UghArvY0oWx
un/sAtYlRK1d0wZ7Ifjm27WyjzbUrbmTTIHY7CaiZIyIzHiVUsPuRbt1fOu207yF
aB21yQ7qRfmdAD10ksR2pL+u2m1oKwYiw7ZHixl7jXAn6sJDAaAJAKyTtp17T871
rVenq/+ceGH84IyOY8legj7tOA/PoJ6MWT9KH16DplRyoOkn1YnD8+NgTJg3AVHl
jwqKCnqW/VNBuw7SaRcXnJT0W9fLEjt3sSV8fjs2le2gSxEG3MFA0IoW2dzIGFFc
vXuDfyAT/k9whCHS0oH2vSy0tDEguYfWaGqPDjLeQgfW/pTK7bKvCXqvI0IrFqhV
qKpkHHjevfPQM1IdeUeTAb1muSW3FvWH+7jc0o7wwYc1oFAbC5EWZAJ3/SXkltRI
03loWmG8GTxpIZXMx+sHOF0ZMPoWhGc3syj6B8CSvXDmKR+V947eU51XDuzO8QQw
2tyxfp757NLC/ymDXF/kZ9S799lsGzZMmdsyUJ2SNUnCFaVjU+G72otlEfKbV0U+
AHeo2S43Xnb5I7TlvENVKZF9zNagIuaaLZaGeW0YBy/PbqbISZlFrpbT3QUQcasL
8sBSPKaDdI0lXGKlAaiqt6UOlcVw6RzMWjH7qRiJ6lyyiHFoCm1f5O8GBX5k7xQ/
Nfil+0LnvfYpv6KeA5qiQIi3n7ojoaeq97BogwnPdXUU68sUrE6q/CKnffzhGkIZ
HJFnQPb+svwP+w0mAK1RusKeQUsadsR8blFLzmAkZBWsudB3+TATZzBX4VS79Jkl
5fnQp7To2guCaNhABJgsqmHxAxIM8FAspQpPxAl2ZM7Utu0ATkWDqTIHP840IYG/
E2ySGgXRWkcDVxEEa8LscddwdLojrefdDlnxAYTsbN3m78M7rzVSoM46bofnT+pc
rqbrpKgR4e2hwwWYkEnMnMvM43VlOB4S6seBWSbLZIq1RmWGE1V/JWIJoaD2Q8ij
s3O56RE0YLaoTVFAO1zihDiw04CYPQjrWtLusPXbDez0lu2z+XWEigiFaQzG3HYb
ezJC0gqHkpiMSNg/5xxCM3jZ2S7vw4C5qkoysFY9LXzrw7C0KQUOUH+PpIdDmtEi
LJva7CkvuKGVJTtvRHSISHP++9y4WvJiTAI1KtKQmJDYWOxHz7BTHiY8oOtsCfCa
9zV9OJL0MBjMYQC2JAFcOYGg02CvMUWTBq+u+YWSMmgZQto4dD6hOvSF6YjY0fgV
UfFX9cXjaKr2AaBZJKbfcCYXX/7wo46Owlr9bk9ve5Os9E51XI2Wz9RFMTllMItI
d4tkVBdJ2hBEqkNhEOXJYw9+vWC7Jzf2GGKYsM8qgimJipr3FTmDrAs0PAqsednh
eWEE3q6MtLjUXnI7LDfy/S1Od7dZf0iiXM606Ns479kZCJmIqjhuEOU4fD+3HqqR
fITExPltExl2U9PP/NwlT9fvKO503EbPhQ8tJlB4vdYyptarofmKOaM3TfV1vGLF
2q+XgvkYC1+wusyxaOoym+5qawcwnQia/GqS6WjHRRlh+CHQQvB1RwObp5soK8HN
mPDEGdd5bM3zKhXMVn7g6iZ+GVtV50S9MnC9NIHEEoLz28uooJbxlJy54RKuPDxY
+U3rFfBcJYtPNcPRdPDPSCmJzIVVFvUCuRet7l+xj0KLIUnirGrO4nM1e160IYKk
Bib+yPsg422l4XL56ZPSyAi18AzfFibMfzmeaCoofzVdBjvgq2zrPw7sttkt3I8t
5FkdPMpfeZmSiAG/ku/DEjDqcXB1GfiCRm46moEMRaGdRQoR9DZKR5d7m5vPAxde
rtSYwzSNKcXO81CgOuuMELRLlK7vUlf6ZFV+8+pupagvDLMqjWt+6h9BeDxrg9qc
pe1EQKTpnNRFCRrrlY559XLEPPRIPTABTnxevNJBmNqEa7bqb5k9vfnNrVGdq4cZ
tijHzF4gIfkBJl6tUMfSIxAXzKu0b3QssCGdKvE5DeNptbnVZ2bhu1tOIX6zDWFp
+kgIH7UIt0dq43H72cTVfsYKzwzbp4Kggs9igJng2S1h9xJR/f0xWiJqRXw30vbA
tidP0RS8R8TYeHPcsrS0YLt0lhfMufusakvFBWVKX1Cw4DpNjBJi5zgDLJonNh5K
HwS5GKzTEF7Z7TgZI211YRui7Z5FcHnlNoX3Ai6XoNrWv29gBGMH+I5DJBNSPgtJ
ZK96PqZxcpZy6PsIiazRJ0BtmF68g/GygzzXrenNV/2D4HcZKwjwpvkeiMHe+y+t
rLHBN7o8ir9PRc8lZvnlVj/pbNJ6T7v5COCBur8fomDsarXHjTAONhMNI5cwzw46
/ixYPjKxK8TjAUhuTICVkGHDIWkgSzom3ETxfVl4hqSOgOyg1irw90u3cbEeKfkA
kdguBTSQBXevFu8B7k08/JSiW46OkQhj4xnntczMh4giD9MGNbrhPPpTrAhMBqiB
wmi21ASgij8bFTDeCRUoxMPY/AFUWw8ai8IdVHEsSZw1KAk75qoEg7M+fquKkOSe
1b5CBiYxK4b/nzcSrxv4nGcHaGGSgGflmeCUtN7OCYq95EFcPj5u4xCb0ZSQ+ufU
j5eX2tw9HyEcz4H68tkRg0oR5ROmZqmiisX9rlewD59S52j/+edatntf5/cWN52S
1JbhqxW6QrQRexDg9bAOw3WuMwfNjkwvaEqTErMHdEULHw/4a5u7p2qfbDg3vi6k
IEJ9m+4Y5JuT8vHVeReI0OOGdEAvuNy45Vn4+MZcIUss/hUGMifgCIy04fSh6tsk
Fu3m4lPVcoYdoQVfGssv7wyVVZN4SEbqpAjfWZt+kPeIunJBOQ3JcWR9QorxLgWv
ONdq2L63VDDNmORSF/+autXsrmnF2Kaulm2NIMZV+5V54nPhswNxRUQ+EhgZoucu
v8ZmjtX9biNyLTj6kUqNSzuZVjrV6pkasWcBnifk54+ghjQL1jNUOFXbOMy6lN6A
8/Y7fKcaH/8PuJphyOEePeVUu7nrQJfpcK/vFZmmaSZ70QcKn4H+LEOy5QmwZ8r/
4UlEqqXfRMmmhsZUae9de1m69SUTfcFBmYxxDiEIRk2DjO3t7uM88xkFtVQ3vu1V
qtjTHwD5lGZWh5r2eN3T3etFqTlq9Ja4liBcinBmGarFejw9FVWUUqFzICA4XR/Q
5rwnqXpbNvNLnCSOybynPFFrKbk/LnCGwn7RsZjwOLX0nM4K3xqiyXiHI+5N4lz2
FDqMkIqAROmaC5MGlcjHLcxbK6gYqY4D6u6F14/X79ryPZLsXBqgafe+iJDQoUSs
qAAzofytY89vS7IC2KOFcq42wypgGnfSpn7EqfzL+PUezVw7pGJ/z42Xgt/3Vpjj
Sa3QlUZCKvqbZV8xkFEbkQmcI6jHC1VlgO3886mlkGFELMuud5WInTtM2VHrdSFz
2BkB4l8/XucxOevd8wQqP+QXlLK9/b8SyjoXZSre1yIVuEJOOStBMhN5Wzkccnsd
V3WiMw1Iok4HAXy8KFDmkBSA1HX3ZLvexCFYV8MHZEaxmkSD0Hk7BeSATHdchkwU
OEb4b2GeH4KNQCeoPD0pns2GCsUSgifWGEtuUyY2FGB9jVmTxOMPdYRvayNrNAEF
/C4zF1ZqhKyFu1QDa6/Vhj+94MHMwT/lDvApxfww1Kc6WQawkv8AQ/q8rT/EWsHs
lgNXbgIzCCxO6jgSOPt/9qfzbYcnpmlBa3/qmRLebjMGqIBX/ZrUaQYP6NAMzvf+
tCMuJa1yc0sqSUQuD2JaxSRK2T+IrJOuB4ZrgmpBeaNBoQo2VQSaTY86YFLrPvK7
KOmhslkyE4suakCzifqZDSSfU5OW7R6lGUPMeZ7KQzIMWeufpiL00NEZq4u4mkQN
BRy39L0vMuV52qz/n/uwhTOic8iWrk0NxG9AmeYCM5yMdC0upAZS3l8rCu0gXAUC
D8QvxrS1+tpg4uCwG1cSJOxXjJ7eq2B4gnydLaLeSmhJRPtOYQx7KhXcsuUBZq2Q
pBh+7yhB1BXW9o9dcMY3p/2yzrc+UnEHqk44NcoAOSAdMCa+S8aVGpnm3P/t9bjn
/o9dG8nAzlYDTjEOuu9hj0sarZUvxuDfn1dx+pIu3+BB/hluklXcPTVCXdP+TGAE
wbaYkiiIX8f9dcHr+I2rfgk/Dc9Pym6J2ntepmczYtGd69iAFB2iiroTgcE10js5
Gz4xxu7E3UhNC79h5MHBqBjsugxeVfwVMAlGqS648qyn9uezKBadqTRw+HONtAXS
iku7AW/UtK+8AHQqQXCRWd3iqUvWmycIbJOOqBOTTPySzCfOlv1Vs5FegZV86SU+
LtzORTdOcUjsn9g/RAEgfQfss7qNj/0gcHSvc2UsqZ6Kl8wi2DXYcKJHArIU+O9Q
QN3mAL7ZyVRFnEFit3TxiOhNM380KE5EoOe7LgcQuuJfEGTpR+dmUwNHy3VT//e1
x0KbycAiAtlSIUhSkh+HIloA0fUYhLVsv1D6d6RPKfnDEQV1Y7d8fTV//Fdk0BNa
yE+vwlQE4EKCLoR1OXgnBMToLvJwdgd0wgf60w6MKl8A2NQ87GBnUeq871cInb52
n//LKLngF4Y0es43G3LjNTddZrGKXK2XTZB0wv5sCOTnTkn1HVni6nk2+QCSel1A
CtEqYYR17XeZQQIAHvhMIezc+ezWtg3ldfDJ2ILeUYzGyTFxb3HJxBRiEgNgm9bK
O99ES4NQCHB2T0AJgN3kE0dAfU0uupkEa+XuxVOJxxuog8q+mSzHYz5QX9/8yef5
O/oRvKCn53y/rl7WDyYuVqP+pbANMqOr0tlI0ppYVK8Njb2gbw5moljkutN3A5sK
QwHW5qBSyFMQoF6ATkYI8Hdx53jVmPgZCMYiM77yKIwgDQ4jRgSZB19z46dX841r
KSZbmeYFhF2a/Fn2TG4ZOUCyS/Vfpz735jU+8B9Pv2wPzJnbH4wt9N5r4wEUc37s
cgr4Y0/GFsEvumAJZIeJBTtOXSB99EFxpfaxntWcENyRl9wUkS3xWH/xk/F+dj5s
ZzQcLRIMIy3E7+7hxRWA/yFctmyUHx1Wk+Kb+4b5EFD+71NQhVohAsdQV2wyXjev
hRJYb/w8cI8uzbTFo8ilULu7jU4fKoEWoBRCOF6AR/YAdkE6JoGrv1jo+C8o10+6
CiuXkze+bSg15Csbvg/2hnbVkwpjeCOdqBY/0+LZK2wGMXjAq3e7NH0qKM/qgrzZ
KWOB+m6qwn+3b3rAD2hxk4GnXn4YyIqS7WrTdR+xKX3+zo0iLQAc+JyVg/CLJqB9
JhU0tcK7yQFktrr7Eos+Gjp7lsI+pmZX01i5yeB07DncNk9k4Ci1yWDCxRcDx35m
wHqs+IC7eotvtvVOA/NZ3OXYfJE8zryN9J3wu5Kal8oayWBmRvQtd4nG4IJBkG5K
KS/6YvN2P1Kjz2ZNbMxbsBLhxqh4FnBN5ejGbYwKsWjnrvQOkobhcZGmsuXy2Bsy
P+lX7d8OMoC5W/4/k2iW+oiKe7oJE6myS+XlExU96IWaHBCkqakcOJMHufhJQ1VO
hrm1PQMAXp3SJ2WPUiQOuKufcpu4CHzEFfgbajzW9iVEW9mu9lyWrF1JqpygzE0U
UwX51DGugA6n0FUMMq7cp2vhsbuwKPANy3uLuG4Ud9iHZH0/QsdggLQ7d65+eb2/
jrFxWoxEHkOHalCEGLtO7quqQ+h0AbjwaZ7BBEk8zjrof0Oil6Tg7/qqRKCNzg0Y
clEHf8dDEzvtY74caKOIKtgjqBIRkVjRFnMaU90PO6lQ80o9YRtN9nViNDSlLMjU
YfYOuAFU2ba60KREu3BCYMwY/XWS4D9+2YoHFfEY7RYJXCnT4XuHSxlMdiVwQPMc
XsGM4Zh1P8exQLaYLikwA436lU9Mcxf9UrgBgDqff/Cm4Vsl2KTLG8PRzufJGPFN
CMBxQXIEgT0fffSLYWtihVp+wARFHeja035GeSUPxIQUOuM5ROUYjga9twE2pSH/
X1HRIEtyzTcUkCdxUG5PGXfDeatXaxH+YQzKNxP9K+CDxRpAAn5/n9YJDZcFuu2g
ZEzuVJXva54H844KR/HcuFR7oPwjqDvYqboy8tTAq1tlOLUA1fkKU5su1yWwTi5H
UQz9lnBiTNKCDXx6qK8HfKV8w98+mt9GU28Hi9HpmUw+seCNfZCRUpmqHLRW+5DA
5/dxmhm3ec65GAAxo8wBrsgTIr5zCXnJLeimU6vFMfnajpM2FAxjb8ZFrfmGM11a
CNLCd88gfYxMJH7YGCZwFAjcXblEFVHaNUOx9FrKPWSjOdc+EVTQcj0tNsCiaHCz
oeinfwZuNazBV07u+Wtvvi3+bV8cUY0EAgsImpg7vJlsYlih4dl30xVozzO6IoYL
/35Wpb1VJlSldpyX9MZtwuk68AyX8b+bApZK4VXvkaPheIDJwCu+FgRrwnHsfaef
Woxl6S15hX6CZdRlJsC1lrVbO9CrXaTmxEkiTjS+7RoB6fRtYuZS8eKPDr/+EuZ2
2F7U3RH7sH9uKdo228LW4uimlaB4GQV20WBJGQTJfQWcojkVCC6wI53c0XIfnz/U
DF6koyPtopzhXLaDTWW5qaTfX8LWB35r36rt2a8O72pFge6KffwaWs1bon3SFePf
7WD6422Y4SkCF6ZcpN6Mk9w6Zc/bM3Ft1c3biIGizxXyIqIVPPvbGx8TMJtWVdQi
9mfY71PQS2YRv0d2ElnPXGuMj281PFnC5DLbblkOsma7Ckbu6GKyx6ZM30Dr66ju
0soZSPY33sWXyYypjRaRollzma4/qbcYEKBDvSAqu/mQ2v/945capRzFC/Ue2kYT
/hlQnQfoaOZ7EFi63o89iYRErPD7xtvk21gfoWnmoe5qP4L5NU9rD/NSKMGkp2Jn
Qd1i/x3GVToXS4JpzUz2bploQlGN6aN5RXCOAgdS7koohIuHkWWqZ4fGcF2MtIBa
Y2sOU28oDFgNmux4LNTdXJAqL07fgcootO/3O59A5mwYteZHvNE7qgLUCHnc4vTA
wq23it9xV4OzOnpbaJoZJEBXfccRBGVmA94MdwAKPAV9f5ZhAzYGSPhanoxVR+86
SW0/aNT0CkiS7LLhPJKyzXB5nB6iJbmXCa7youaB1Q75nl0J0MnMyxhqFXA+Ke2e
rjszaqwnYr4DprRbXQv8h3vNO041iC3h5Llw3UGy5Qrt9ccnaabs+KVKLzHH/aw/
hoFdMXTgInGdUpgOH9RkWXKqUM3KWQbRCgimBxZgxt5PugLzkfmf9umY0HMp8ley
Ii7+iF6gUCMnDDmlIz6uWsgodn7CDDLfcZAIsUGnUtzXTLgUvT3DM2iSOh2qvJjv
b38RGYwRVqkmDtbjM1w92CQ0763neHo9BOCinJ0p48YTSQckcfUIkY0AmAVGy/2S
nx7p5h/B3R9uDkHgYh20xy5A0q8Y8CdoZKTtB72fxv7PVImMiM9hj1piIVT2/w5Q
yhuIam4/hmbJ0s0GjSFTAE1iT64HfH8sE/tUmXu3R1/VzLYMasDz+scyuZcGUTDV
36rjPadDIVkifG5vPWK/PZDcUdHwa/dXd3N4KM229C6PoWkH7AkR9lgJSzvZA47L
52GA2u9yOojRZW3PMAPeJ0VQFbRB3ySYb+YQ4Os0HXLtsnzzWb82bR3GCVnz8stk
lVTppKpQsMvGyoDF4SpW+wkb0RKS4PShUFo/nWvzLGMeb4nGaf1vci/494zklQs8
y9Y3FSml+okR/MyLDoNqSejcuo9Ycj+fXqpKBdyFcqy/OpZLHxOXSxRaTjyy5gsA
JfhoCGZq2dlivFCNn6oBqTYUdPQ9Xtcrl7quJHxAmu3Awb5sHIhEAjvmhHpdgXhC
snCB6ozjhe2tv4ApNYoInzUwkOExw9YkBppSjT18sTaol5GZrt6aD8uPuu0j1DaE
hI/ll5bVVBosxxPaAl7xF97X1oj1+UZOpTg6Ybv0lFb+WRifU9MJpgk4NU2Tklbm
ON5tcOXV4CdlK74tjuvTn5ilQDI/o+pmZG5xA7bVNDKSPeLvs4bl/SV82oevsGrd
jAyqBCgAWgRBVCcrrX4ndkMlkRl8OhA31ogwRE7g1mOVuitpWAjqIiin6Naf0bcD
7os6AhV8kadSfq2Vh2VlxqGbuykKLm9RANga9FtbCdm4HlshOC8VkeJkmEZEBqeY
306ihUxtsXfH98Jb+uKuv6h25/5JHUvlE9RBICXNyxIB1wRc5nwTVfREYCk0OBax
eGWr6Uxb24IItGObCrVxMVo2MxSRtDCrKFkciUxdPf4yNbB7ti4T+iX2ZXQSwcde
nCL1xBXKWlhK9mIjsYWRMPEoFGDpkYI0LQw3zVmnxQk3NHRuO2ZL50hGzt1hxGsW
fLnCpiYwKCtxA0I/sU6Nf4Q4HND6ViAofcMfC0b9aVy6kLUJiqP4OwxBsnPVl4j6
p1wgC0EzzFl/w+1O+MUrl20ev0OdZyJVlpe7DeJ9Hd80aiwFO13p8QG0+tl5rmiL
lJ9WzErxkESTp9MAo0CIumaYNIZq7zJz+gse4msIL7Wtt1XjzZJhMwRn+UcoEk2R
Apt0peLHE0WGG4Se5Qfrtf/EMZucjQJBQrcNS4hZXdTA5dvZxz7i4jFoJqrCZ51y
FvFmJnXevFXYzZeZNZRBDCEaxJEK4Khgph8Ak0mLBp79lpZ3+vC5IXPStNk6KXrW
FodSUDsWiWJ1s12/D/PZd6uy0PSbQYrH4+lvZ6br9KHVX6MEvEi5RwTs2tihTyqB
Z8rXniHFRQKMARQRE0XxkR67NxRWol3aftfVj7UEHWuVxuyCfpFL8Ne87o3hFr1z
2w5KE2E+maR6ZmET7NBe7Wwnif18BsyfcFg5nCm3I/Um1xnFwjyBXUphqGvV+b5e
7Qii3JiwgL2mylHpp4oWilF4COa7Hh7kUH38gobQM8ChuElB2epJZqLBtsAIiXn8
8XDQbpIx6CC4nNLcqAbw0xZ5HAMDAfj/SM5Fhp6ZedoSoC1AVTkRG/5oa24rJ7w6
skfHS5dGi61ooY6jLZx4N4DFc6q/+mRh9YKh8E3D7T/qYnkR8PaKq3h89xBdRLHY
jTdnjnwzz0COaG2zdmMds5si5n2XxH/bijegLGSDbPFYiv8mpGhpTs88xj3izNrn
FZq6noZK8w2rbiriYpxVVMWDS9giPgAR4QE5WD2VEV4XjrbZXhj9Z8OUHXoFyWBX
YFgG0gVFKGHehla35HYLi2D8634jGLrC80oLXyI0U4dwdfGD1zd+EpX8DKwnHWfe
RDcQV9Md/NvtqHA8GPjI8BK0FD2gj1y+Gc5vhtOI40UxYnXe16rJfTgi1bWnLhj0
8Iq/mK4xtwYZ4fApN9baP6jBK4C19X9tuPO/cAcU9u8jzFBnCItMQJExJBlt3qqO
9MpaRIc2ByzA5Q85P/5CwjDFK4ZDtH+c6LIgComwHNqKDECSWjJCr9y/SekdtI7l
Wkw2+6GtJn73b9tHH88Hf6GuItnIjk3Q3LdQij6taWEbW0DC/FFpakMvBUIadgA8
OcxibkktatqgEEYLkMIBLTLuaMikqGw+oPSj0J7LEKj6r1t/oc6jIEoMr6wICfbO
6w8X65ylu7pnGkFcdqe4sWmREF9EFj9eR4onI4QjmL9OIhl/Mqs0yoSguXpgUm+L
lxABbmtn/5MKnriPjfUe5JmaEb22SvP0LeaqXXP+7bmWN5jeFYBztOhjzjNQmdPv
X/MbLyzXm+/1uOeRsYDbH4WETU2DIHOK4HZEbnkrIAM+qB24DE0D0HJWujlZn1XE
vzKU5wJe2qkjS1dHq83olYDEsADjvBhjYREsaH3lHk7yNqGACu2Y6b7w0eXnE8Nd
mTW+wKwGhYOo2sni+jdw19jlcFFdBkR2ULLZbMl7yHA2GS2thwjzCBlFL1KdsAIy
2xOidHofeGgPX+A6PIGOENR9YFhzoXjLvrKROVxSEyT3A2CiPy5K9h/n1kltXCwc
xb/6sCJL6JZWkxbcXANKTi0H5tmifqBx1aDhJAD3sXX3PBeQfbN2a8TMagsm1Rt5
YOUp7F2ET8E9FNPsiuscP+W3CFQAYv05lfln8YCPJPzSqm7AT42+aIgiABOjrX7F
1fgRDUC7eEZYEaguDXIMY9HAlcLMpm0LQ81lKi7/jc60X/h/hb/fzaCACc+d1ISH
RKcfZurcLq5/ZShvwangdGug5n56VzRo4zOcpalOdc59Z3kanjUa8E38h2/av/my
3gmNOLWxaopjcZoXAU97SjsiwRQ3ctxxCI8O7ke5+ymrhOm1BbQ0If0aocz4nb7s
5+OvMkLBifbRVdN3i0WLq642cAkA9r/JEkvvNJFAG/mDN/xvIEp8wVPzz0YLdCRg
KBJUAiqyAmA5jQomr+SNnfF8P3NoyUev893Ghuy+97owFG39FuN7xwRj9Fk29VDL
zyvAOlu22auwMC1OVIkkz5DdmQbon9T+g9v3wHAaxpZ/TADVwgw04HA0HbWz2eMF
E2UKEmuUXIDxYBf82xXuxvbjMY5BHNlJZp/pJ+RgfNDnywEo0WRimEd7K05L5k/B
29C/RLQZc6IGZarJVy+jDOJnM+7T1Ro7krVi61UQfTBlgIY+shGw2r3hbRjPeW3D
In+ILCy8/0VEE93iSceDfwXW3ee1QCHlQour/OJ6wCEVmqKe7Yd1WI5ouJsT/g5Z
jrrlKSZD+9jX+M69Sl0fvAYBpfcg7r8O4vntKuIUp0gnm/zO6F3CjRywP1RsK2ot
33WKYAXrPN7sUs6qvEwxpnbdWyPC884MKwWM4rmGktMQJmmjObvNx3aMMsDncQhv
ByWTtLpy09dQ4jyoMmmFnLKq6DxLebVX4/EBarJ9ptiHPVLTqUCcoKvTHIQO4bmC
7Ig0fRxqjjTjtw04pR3hvuA7xbsyBw7bHWpboaZLqdpl1Bfv6fxKFVVR537LHtip
/D9LEXELZHIO2AQFFwCFNvnWHrmLh95v/0CQIue1XbCYUfd1xfgEGIfZAuoCJK7w
BKiSNX+F7NTzGkNKGbGwmUSyvVE+r2Avk7oGZyYp27XXCJMNTXrHlyE1e5F5ybkn
K9W5R+Ow1FiEaEV9iHGo7imTg7QPyFp+o8hnJc3jV7guMpiCJVLZDOE0RZ7L+UUJ
ZM+yAAr6DGWjeVs03sqi/N0Xqvf1Ydo2ows9ZbsFWDJys/Jvg42PYL3s/JTAOfZq
QbNrtOMFOug19927lE/YSMIxxyrs0GpEJADkM4w3ePb/R3X9QFK7OQgLqOK+nHI7
UKCXDnqSm9AXAjRHmeUfFHT/VuPgYST0rs+NKOPfqYGj52wU63m+JBfMWMEGDJVs
DVZzTG4Ifg5m4bzgA3PbjVUQZSb9j2RRlU26Kr5AkT+83wFRP8+RxmfcVqJIv2S9
j9AfawRoACPEpYn3If5WV2egzA8gKvPWtbhiwLxZk3zJdqpNVgRkhYMOxRzmdjvF
DS9DPqblf7oUR9yKC6TaSooOqFgpK2tX5B14C3l6W2CIi/gJbtW9lIBC59Bonwca
6gflndezv0mbZGfeRtq4A8tmN1V5DjDzYA2+NSUbuk8yFgp5FNLfcx0t8CWKmwea
Lt5bIos2selUCT4KWdFZ63+WlVyst45oZz5Y0A7fbXXpRFSoSxSQ9Mcp6Rx5fOOB
HaG4gztf2odNx42FqwEdZNQEZJszQcP6NDhJoO47GF/J+yhQy2wg16XrPXc81yAs
SQ3XllzqdjB5z6zOFsfr68/xtlhf3DX1PkhO1pREPwxC6rXuW8Tlp9FOqgNSnliR
3gJer9VR5nm7C2OEXA0c382ZL5r5Mq+/3trfacGtj1q4SXTo+1ANl9XEEa6FKK+E
eTp2QoOp2x6g8B4N9QalTYtkuPIxZBoH7N7n494DSkJebsd2/227rGp+eC3RYkLe
/HOAqmHdJTwa21G2pFwFtTN8MYj7KihG4ub/ok0xF2dCpVtUEJH9J2+IcOe6G/JB
9sID8LGFQZZCi+ZczxEd8WrMup5Zagpbl7pXEicBTX+5DtJNPrc9AnrjNzTwGJqB
d5K7zRSbZ0nA7mtu6l5UVqrFvqIfY08PUBHqEj230ZoN1krdmkwdLAVkrxFi+ie7
SmA8J39UFA6ukiXfFLBCEKlz+ZaK2zIixfbfP3jOe3dIoleZSRorlY3G/fiIQjUH
slwcqahVgSptT7pX7ztqaepveLrQZs3XQzGWbq63vujGUbFX5uvp2iWUoNYEfUaH
1GJDMzlQMPgJQJgsthCcpba0qG3O/oEZMidkmd53fm0vGZECaf+3xl43Ee4Awf7X
pS8SBkkR/xsQJuMz1bCw1I1t3OWttkyhAf4RPYa2pRu1A/ikv2sCIelIxXppX6T+
/HDKTYt6r/ga8ygOygM9SDWBcTEiezMX+kUeqLHRhlH7j2pE2WtncYWUDDq38zVG
tw1OOLAzse4gHuBvsJpfgVjdtNIBB7Yw+r/cORtIaqpej1B51lAUGpJIXVMea+Kf
xipYapMPcHJMadX+d+4HhR0eKFCSsUMtqLNjgICLbcY45EkiIbcwPUjPqyJ/lfTC
JaYPPlczyocqOLHkfuo7WiayBCiT0Pa+22uE0/118P5qVmAZmhp6TXv5429qhgTr
3jJ835xL6oDl2B1nFe5Sf/4En1O+WLJif9GROILEgNxmjbVuXz9RJ326WlQlbB4a
VjasnW/GLPj2cTe3gmYFSM7dQ11AFIA28QDSdmRZwWVkd5uecarHtGH9im5s0ed9
oEmR05ht8W5pCkXGGAej8P2d9Qez8h2zCeK8kC/6lR+xpdn+6NJgPAc4jWAm8J0/
YaVehEzMNma1n1X0x3fbAXlg5Q4dGEVXYkfgdQzr+imt7KNz9VMAPf/+7mFbMOJH
TQ0gYdFpZA2WGtunl03lERmv8Ol64YOew2hKW6CodibUIBp28ZsKbyNsGERdj1E4
lGfSedVgz5dwSkdhIH2ZuJSi9+IXL31lGFtTcQ4RFImvIZQ1lSFrvg5fUjrK1RAX
i8D+2xk/xK8vDbe8p+N8Tj3SQwpF82phsVqdM2sGbvlDJ41/k53LOVhoEGEf/Iqg
4llPm9uLtyTlgvCIqIxCwTwx+soIEwBfN9KpMrDu8vHTAjlISq+Wr4yEkp3LzoDp
OgEbJtFnZio46Ahi2IlYHCB3Wq2nI8PE3Uzkl/rtd3P1IYW+jeGjye5aL2wiCBcp
9ChsTKm0Vmo9+PNtYc1L+Gp3E8G8UDFY3/adUTZXgacy0+U618Ixknpv46SwcGER
U5dXDO7334AyTIi6nonWWrUCs7x39tJvXohtz5URyZL/g8x+OSj49RBlNzceRE8K
Z0rGq7LqSfc2bcp0FCAE1NnE3jHOZqFbO6mSwUFjc+I7mPCKuzgYxX6QwjBVIRyG
Nh6XHWm4sNOlBES0A91pgG0Sveci6z0hDKvJrSZSPq5ev3dh9F5D2+JQCM8ZoIVR
Z2D5Ib+0MsszRYa7TAo+mhXs1Iz8lLbKKP0LbkhLW8TdP6z68gT23qJS6gXjGaSx
JjjH2G4/snlNT8wtkRCzsoY4txaaJEkvcRc2crnP+zfNQakAe9h/OeGHB9KZ7D6y
WLBpNZo9ZRXbN4WD8ET5yPHQOkLjw36kNRS2sp5erHP+rJffFxcd6fnnal9Yfblk
VcBAvB/Ju0D9ihuqMCJgM2ZP9WMbVe4xCjCwkTGODkYE/Npp0rt/AciFCVSY3HTn
EqziKYfmPDfLZyBJh//rT6Xo/dfjw+zwGxvCxuX93LnBd1kYLywSKp1MeEiRJ67W
o4PZ1FJNssA0j323AwNvxc3kQ9b5tnc58XyEoWJCugne3OXTJHjfApF6SXzk9+N4
wz47KVOCNu3Ge4I+KJNsSqc1Ampgy2i3wErzWqnQK7nNR/aNYV9dncaC7sP6Co08
rWdAMx6o/ReYIw4g/W0QZp3RPVZM1RPt4XChtYeiQIiiPxjZSKuwjx1JdfJMf87W
DuVHnwyG2yG96RXuzva437Yigcqe0WRqf++3Ie+v/Yk1h4wxDhlGMyQPgqzpnP2x
attCBiPEVbBHxAElMogX0ifl2PzjUHpVsQZbdBo8gtd4Nafe0jtsBVaerQsxGEDM
MCcOeibFw0k+25ktSfCHaihbZH8QNAD8Q4xbZH+nlQrpoVgPuZcS8//J2E20VLqF
aEVcqydy6vjbRZRKT4bn0AEbb2YYFn1A36F37ygEWHXOJ3ZN2HTNFvV41NI3WR9h
eVB3qjgQlo2aAB3MzKGCzvcwRJT6MmxZP0RKUv/prrMJy/VZC9rB1ol33xPKnJ9X
0IJZG7rGwYG2oHpGUnFXFkQOJEJ641ykI5sK8oaxH7BmL6QMc1T6zvlYjq85z9kl
Gcm2hCc5o0+sHk1mJcG7DlEP3CaNpQ3VwNHrlDDaJmde/GAALP0JI6lG4GXb7PJk
OarXdTeeKolN8fygf0Lf0HzMMEA22oL2ZCmORsYEV8AygXu0pOCdPBUULNmikcb2
YiUkJgarg1zvEXyq46sEAKz3P/AsloQpRTEJ9YuuisyhhnVzenx4CsnVgAlPzC2D
FMDDNqRFfdnGQvtWrc5a7BSNIZhcvHGHutWNUGxMQOZbuu5hybbo5+0lVhU2TKIq
a+lrYFxIXDooPtHgsI7YZGCHZ6DGCCwxV8BFhm3MySSho1lTe/ycYOk5mt0Lt+H9
U/YXwVme+I2EOlOPdpKYgDezezAOeMFqTrOdykGjTsEgHnGUPQmCBvPUF8AId5g2
BZDjfIguetMNcoLBny/WJsr5X8AMxoKEZTH0UTzA9sU3Fzky9SNZJmzSTuREyQ16
VfWrmg75kEeqscg1cbai594LHYlYNFb9L8aApOuiODkDbjwzC8aYQmDJ5SQhn5EI
5A3G7wJex1j+PEuG+UDO6f1u5fsQrV8F85ZBWgfBDISZg70dVXcChhX+t83Yue+X
gYsaN5gQSR0Bs5JCXsjlKsaGw7chAhGljuhYyZwmlSMFpuAsL/JTahGb2Mdb5sO3
cpsc7E3lTEhkAxXWsHGSZHlTq1Uk1UVGEFL//Z5hpUuvWjJ7ry+H2fY64CvIZzMK
ZVFryp9HCIhF8iQG0EI8TO3a6ZhqX42CGyDAJJkkM9mKZMP7RptcwX5V3KQiOrOL
YupaZbcw1G+N8nj/Y9/ie1NaP0E3rC5yi6vOhR6ke/Hm16W9nOS1qEvIeIeTbZ/e
mIGuGr9+JRQFZHvTiUd3Qxlqe1ZMbCWZYyYTJe/hqviVu4ug2hBtxkt7WISlgnwn
O7iIzImBJO3qnzhzEeT9mLzTUMxznTIXwk867HcewIkg3rHEXICmeB+pTU/R6VUn
h6VAJmrxicYy6uHIdzpdO93bnijWKesSqGAXusmWLStzF1CLVAhezI/fqQFKVlCR
CVXjljIYmXSGKx7IPFMCSD5Up4AO17Bi3eq0pxNxKfCEIEjs80PIrQfoLIguZIWY
2NRpaH/n/tQ4iYn2WNpLyXmWVhkz8SDUXlQekkLUNdgkC+KSXpjxtE4AjNSwU42O
gVdbnIpavEejxPirzvjgO1B2AOOpU0xG5MwTySchQDtc0PuZJQmE1tIhrERB9LzU
7x9dRuTBT/2oQWOFOEJPzZ6Nm41ar4h1rPIpLQvRtbLktQNNa1ziMV9tbgi/BXUI
YfBGpq80hZCiKWSW0QK1SvRex95XttKTVuF6rROhqD7cNTFol8vCe4do3qMy8jns
rZ+KqDYEdxEhLa4GEsGDKfmRB8KKQ8BILvA967t27EW7F0LPQvZEAJX9ObLNHLJn
JcV1fK8aX+ldST0BWQQ3R/qwy9Kvi9/2Im2jBwD9hy/4ualnFQqvTPMsfYjsT8Iq
ry9Hccq4F+X8RTMfvyRF1LWDTFNFBIXLpIGvOuThnLQMhvEZqRk0tqPy9X04krfw
5vabJIfroB8nUxxU+NXDJiBXezoOZJDNHEmqVAM5gv8MDP5pWx6BH7BgK6p65eBD
DcXuzfwckDu+THXolCIZdqc8cuKrEHoc56VdzP1BidXRNJfzXfc9R/q9kOO9/MhI
SG4dOsJ0k5xLuhGLvytYUiIoklrzUhsevB65BlVAYap5rZGc/jfTarODXhFhmPuH
hpx6BIfEP+mEsfP/Y4qq00A2iHkALrTNg0WKSf2RPA1ghyoB7Oi8fdWeXiywiPwQ
jmBJeO8mgnX3QKXXyVKC+bJVyEjLtx8wysoR/OqVGPz8nmTIU2rKHlUkVv5qnyEg
60vtFJ/dKG+5zqnuaFfW/e5CzLPHhPBMED9dxRy/8DCohRGGkgWVGQF++APkmBpd
MxRYhyoWvH/K8Hdolpyycsc1aEAcZtDgLfFRGmSE+ZV24si3kgbl715bARXERkza
Gm5rTiU4wpRFftA8NkrShowIEphNbmG/n5BOXT5uog7W2QlJOBNEW37nwBhyfMBu
R4xmrFXdz8jhIEYELoO4TuvTKfl0vHciP2SxDq19y23/579M98ZR++lLF5SUdiqi
DIauxTjF6Xscj5YNWj+/G/mLtk7h0kg2yC4lMxF+lc3dRDfflnwAHgP2jG096TS0
YsyxgehCvfA7FIxjsiwKAbY366yYHj4WSyLx+Dr6j4YbJo/U+qbk6mrQktDxNb5E
e14UzBCAPDMCVSmHQ+Xu0J1mf0C//2zCsYrY7TNYnswkck9sNpXAVd7h6kaCNckl
o7Kijzoh23TEvrQHegHcbhxp/95KgbNk+5QBDwPAFDfPpTXjFih7W63yQpZj3HI+
yB8LyujtwzihzLyWNET0PIh4NL5Vu2fYYF8Ssr4RRQG4SKftK9nNkT1Y8hruKhAl
9/CkvG5T+8ovG+IULamOPnr47AxBkSSuKlwkgZdWnwEe8dTOkcVfU/dukrkpFNXN
l0pFOhnT1HSe3waHi57stgZyEPcoSaXYLm7eUDKsU76zzbv2yrH9KlZMuvRHurVD
Bg+BQmfnIK/CjlSBlzdNmmexnW6BdvYHc4WSfCmY5mrNW9FeZJHl/cNlgkx/ETVb
lQqYOpNm9sh4FLjRNQo/KHdYHLGQ+QEzsnx0/nEVrrmQQMfQADVW3/ljz1mFHodc
UI/lnkkW7dYXQ7icFM4dfcOvkpFzfnl4BGbyv1KlnTxQK3oZsiV4X/91Cef3a7r+
mnEeqBuvS1+zaPT94C7IvyFLJL/0Qpb5z3QDHTlhZFDXBq2vReCHj8qoYccNCCwS
l/uNSrtuubQ9p4kRxBON4bu1ZBqUI6T4xI11ljHQt5wCHJf3VjQdEcW82CQaFm5u
mgEE7x+66x8mmu5pxvXsQAuPg/KOaWGTDZJJRKsx+/nZ+mARTDMJsFvH3G1C6jpp
WIOIEur+ZHYNnlAEfH/m8xUyyANqHS85QBA9WGhCvC6Z/RgVBvd3cjgQMAcyaxy2
Qo1PpohvHvHg6B1/mSs+UXShjJWxRAt8BeF1C777MkQchZg1epENFDUtm7HCNv2C
pFOTKcSjqoHJ7mMV20/7iGKniAG+GJo3WIX1MwKUhLFwD2i/LQzglNKqGh/TaEWJ
fYzlvQV/AHRUfvrLcgD0s3RzwTHUR2Y8EK0bjgEzdPoaxQTXFSXTUlaDBpLrr/Cc
59VeU/mTO8xB2pfY4wrmE1GsWy8NlanbYxUprAQkV+of6NJ1VjcZYCYDs4yJmalK
XwNDmZo6EkmFfIsxnZVpnW92Zwdc2MuoQGAvvKjudJAe5Yk6NOHoaLzIbqsEs3v6
kZtz8IWk2eedGIGwz+ydLt9T7zGgs74keG3PjV5kLVqSP11eBWxHAXUHiCDjkTba
J0zO26I/u2qPxjk7SfV42w9/pt7FpudzNFt4KF7mbFkyeRhnrkpezSbqkZYFej/Z
M9WD9slO8XwpegZUz53CW+MrfTXUPPp8NomRLVEYDAGRIggW3wEJeLesfyXIp1RX
bcGRLscAHzFB8EjYxzVW9o5y3Hor8YI1y6SbvyGjvKguaKeL0+uqiYOyDg3ooKJi
JBAvv78Ir8WnIlo+naYIL1NQdlBSe/zufs8RQAsQpOhdEDixe6y2UePBkx+B+j11
O3uYr0ZjyncTX0iL1kiIFW4fLlIKB3s9xHF7Q+ikqDlu/mh483dFcMcoTIm05nkT
+sQbbafTastPpvUvDWAzjKE6ySUMOUpOqcAFd4vNN2Y5XkqasKhFS8234HXInkTt
6kYBMlY4NPwroEd3CgFhFpFD8Bokc/scLQxjLwCBLzKX6uCYR8QS28PrOgFM2Zye
VpZ4Re7WnebSUPLGwUo+lgZf1/F5Pd322NacgyuDzzhh458lxFD1SvPBMdVEZy5g
FFPyVK+srUIGVPSx4ExOQfNBd1dsgwpfb9uZqbJqM0JFn3AUesRVbnZtUg6Ioqli
2PSKSi9uadtmY8slskz3DieZXZEGvrzBD1R0j71cims5YICvhE0RM8xK8+3e/Dq7
40NnTUpMlrjLO12ENf/PETeA01Vq7H6zglL+Lp3jwU7120h7NSS1Sh+Ht1u5Y5+s
yyKPyRpsZ0sZrpirZljtqPBkAqFgDHhT8gp/biLfpAaY7vjesowEm6iaporcR6bh
Cx+Bny3lr2U4PkrYdLD6O4mpNpLMp78183zNHapvPBqo0ubIyS+WjbqLenM1kpMv
o8PGD/zpgk/S4+GnsiK4Q3HxDzeVoGe8ly+P0SrQRqm2JMMpKQMguWjzwMCbB63s
B2KccgLY99otYlUBsVqKyR7WK5hhAY8e2T4BeEvbOolv/Xc3AX9mjYkdwock1PCB
SIttdJu6IhKkbduga3UlOycbyT3ijCx6GicapNvxtxJT6Z6V0xBs5qsxYlRARaP0
EeXeCUb1c2DFLSYCrHC2Yd8aJWFaD0IlkL2loTjvQ9t8clbMTBRtnxufMzm0td5i
z409pUHpgbL6DLgbN9oPXrIlMR3hfRS8f2qjjTajocs37e748UD8Y8vVy3pVDLID
HiXgz3rgWZQuyGM6NO8jbO2iaxxpINU6bEwB4Uxra7hTvg0yRJqtMymDSSV/AUjJ
mXJXnUejuMhF4tCfn+15/cjSqZn5Aut20wM7ENPPhK8UJRkoGB96khPRdswJv0H+
Sn5cSCgLLPv7LK5IP8tKF2w22KHXidlgdEN+BK8DGEk1VeZV+hGAFb4gloFGQVLi
JexNiHx73SM3VGj8e+oEm2qB8Y1OsymUqoVTb8/r/mfAmg/3gFOsBzvSuyc3vGf9
Orrq10bMgI0Oek61q3pY4UUwYY8e2Y8Tny5DPF7P10Z48XZ1Hr1E3qsnE3zImoLY
rxUDFPlmj0x/ZDbvwR3aSOTRi3fy4ENyrNTm6mBPSsRl9XxVenw59k960nWCcW9q
RqdJmwNWYP9cQTBtY7EiOwqCBB2Q0USg3Xs3RKIjUxKPDGWrY+vQ4Apk7gKz1S28
E/tTo/PfxoDqTNG73UeXYc74WwhCD1j+3LDMWRWP2sXPuBVNAXGt0lM8E/RVFqW1
MOZZDlDQgLAW6ufImHulIeT5aM8MEZW2seCVd6ulThF2Ba3GxaHcR+2LNOIG8r4Z
ai6kkRIf+F3el5Mt5cBBvWEvrS8Qbs2NKqFFTTQxyZVVpyP7xRmmBALYhmY3Asv1
bxSZsIqjRWtJpEC9Q/iHDbUvscgirVHeFbXyrYdpRZNTgsv7wQNOEdOp4xt/+RXx
zlheieLZ4c+82lEv+6pBxN1uQZEWNp7IRnTfoHpvhxhi38wwJUjaNg4KNQYPZXw/
jlhq4Vg9OGzzTb+apqkngDrT/l9cN9OTqyhxtlNepRgD5U2M0Yg8CDqFGPEGTVtS
OKg3SQOs/7ka0oOlLARds/3P2lO/m/qRAFh2TEEWFr09PkjaFAaU50lAopQISl4+
oo8H1f73lAvDa2DSx/O8ZrIEK0c3ngCldke0OK4PgJi9bOKUZOkUZ/YSn8ccLeQV
NljoIeNbvWkFbu0GE9EqF63BKqHyR7a2V+0FRa3soL5c+eFzidrocR+OuuIgH0Yw
q4GPhywmxhlh5DEGGUis7XxvgjCeL/ZW47MriXyUBq2QZ/dlNhHcV2Xl/1RvmUcm
ukYoRtctAjWdM53wXscJ2wqj7WGwHS98uhql9Dxf3/Vd70uR7hpzu9Ci8ph0O25O
wYd8cdTtRPt88PvzbW3/nuK3CpKwltGSEgz56Iw1Sl0Uhh5H/2XgybNjTxu8L7XE
HgLk2zWX0qS+PZ6o/5FQ7o7bvGpRR/4FBbAxHNKiojXownWR4TRWt9Xt/gYcvUHl
iuzRKSnETXzf78Q6LZ2mFpbhxvbwT8T1dlQF9gaOV9QFkMSgTa2b3nEEtkrVuNjt
dmMWOLgNRVK+yKllKBv5mZmbQZoNaztTpnp1ujTri2SFmpSwHfVkHpLQbmClYAbx
57JinJRZVIQAWQVoOTbtpS1mXcOTtrfDGQhibcC45LegAyyHyWf2fcHeu+MckZh/
jAkHZeRZPgOaPibFdWaXZBbfS3+yYtHCiTws8sxY7U0gCoudhQ6gvcFsI+arHa8u
y/CP+U/Yhxv5prRfoyQx7a4FveFJEE/uHHa8ULW91+Wu5Bp6RokWOGFNRiyVUyUf
+euUELO0wqlHYn7giRHTFqHRNzjOwIiFyKt4g+1e2ttfBiSnJYKsHHsWi6eMBFEa
qAL1wbw3Z/3ijYexGdcypU0rwEUE4eLULfKmRe9JOGk97oVHIaixZxrfgEUchX8w
9c0Xm7eBBwNvqa9pkOQoxGQKtq25DERHQ7iLd8bptXLG4q8+Rp7TBtJw8GPsHgt+
Wl6jMZ2c5l5XT+exu1NousOfbtxHTZKM6TZWf4J2Xj5BCsk/YZIAv+DAHgthuNDk
cxaARhtNtwu7+6qer9tI2hOFre4TXHtWiSxg6hMhMS1m0lAb2K1oaGxlgn01NFDp
9L2kR3MPLQZrxOBL45tMRUwq7j0MOixjnGndGSDZgnxAjoViuVsuBS2Au9NJZj2R
UXTITaLA1RjMPPbLHr6ThPetRt3Y/nQFWhsokNBLuwvpYmaFO3aYx+y9MMeLrRWQ
8Eolyf0kmSOqJP2/r77z9iifrV325SL87/TdqsL1SogBBTaOcmN9we5MKZFDjx24
Op+P5kSKmBZmlS23Ftp+PhhrWpobq93ASCJCUMnX15kF5yqXGAlcvKTtzDHgxO0Y
No1AD83JRgR12aUQsOOwdk1WN1XkCkjxGn41RFLd1RLiJ9p3ZzvpjFsIR8gftaY6
qNZ/9oQ+S1uBaCg5xjE/TKjnefq62Ho8lkLBRHCRnjSPCrfun8lSKwdUpQZjQMrp
+t2nCSyjJOX6e8OHLJdevLutMmajcaIvGa3x71gtGi83oum26apYENrKF5s8HVs0
svLqPRjZjbJ0A7dxgYTZR3jb78Gy5bnqP6RTQ/soAN34BBD8dqIdU1rbeYZYCcFR
b0eh1lcO9t03aF1kpdtdZl4FgIy4gqlqfw/PtwATmrjYc1FM9UX6ShYUE/FL6QKe
PakFlW89asg0g69xM9dov0wsWiismQe1lpXEy4bakyjk6ouPVehFSZQ8IhEgafQR
7sUx31ka40J4IfUsA6Ik3E/Lst7yKatRYRXfpYSrIM1w9j7lYhyPbZVPTFIbPCi0
hjEqybLsY7gvlKsuhxGiRABNfYDumnZzgVahez6JWaB/OQrjJ1lfBaSIHk+Sl23P
x6Ebuz400YDO1zdWXuMrj5GMaEb/gWfxGA+d5uwREUTW0cmjnXz/A7o0h4QS4kVJ
1HvE5RKU72e6rIi4ClOEnkjKG5lUBDpPJ2R6RroqMvopQKpoPKa+rEw4S85WTC4O
/NxUeaR4Nb2uFj2u824NnY7Vc+tAz2FMopckIo8oew6+dU9b5uL9NXy4rrcjxXcB
aVplEiA7YQuvdMv130oovLz3yUrHrU1AT8HWyh1CpPV25GIR9jBbF3pFkqUBL4hg
B+euwepZiMyRUWwFq1aKk1P3oV7ZCkvJ2+wkEl3yTIW6DfdogcnrCnUozyvPJYKR
gTUjrFkF0RuOQJMTq5DtVeH3oZBQMy6EaiSpeDYvnzMrIHsG/GS9JheJL0s3VI/x
C26rfo8Gs2IZDE5HuiuD6T0ePOcf+QiJAKjUFCoEujQmNoEboPMkhf9dcyuKqCwI
ZzKWtBWxbJqdn0SJb9d8d4Q47Xb+PP0IMEgUJ0NOl2NEG+pN3eU9dTtCR7kNeQHo
oDp/iKBKs+O00DtiPYrfH1LHEizDPzH2cY8wlASelLHPGvsWNFaHaVUGtbz9ZL9d
u1/qbWwEdE9seYKybVX+PibyQCPDA4aERNK5pW75HnVfBx+VEuIP2jVhmrBlmQP3
9P8y9/Pi3iylYaBjdTsXT43QDX4CD+MvU5ukMHABbq1e8xFky5XpQhV56Al4xZ8B
TFLTpo1OHf30dinpdgFQdsRus3xc0D3NS8Uy/cwkI+RPLAJOalHffYy3rQT+3aGI
l27IC0nhQ3JrumGl+BxZFv2LIAEzTMdT02rD/ldwkiJJENkOOUzOyYQsdg8Mobzc
XRSLfpVWEkIu/69WM0pJn4tPBMcns+W1zi3FiBaM+18SCNK/b1jd+RvbkM3sJ1jy
KrisqoK/hSxk/gVIA3pAg9oKimybVh9NGdydLFZP8BT9nA3268xObdo+Cp2BjE9M
xhkajFeb9sNjySKfDCi4/QhNhav0p7vdMiYzS4poBbap2oYhH/GacP3staKTKsMc
8hEqcYrIXuhPJkB+GPl5Oh9qsyyCduKU4tUvdDmtxVjUvF/gWeXtSBYOgRp705LD
8EkKa2nmi5RI57FjkPWPrgydEu2UMpEwcib27qaOxnJWe5y7uBeCg1aBauB8RkLV
znB/AtExZwXdLIsTAI0TfmYIj5uJzT8dMMfkgR2wp18vlk6pbIIihrd44W7Gq4aq
ArjrAIroansM/uABle19q3xz09uBkNWwdJk4KFSJHdegoQIeBzB0FOHmDFZTO6fP
Pshgg2ypwSNDoKGFoJStB3Qw/MuAvhWbvuKAVQFMGhDCRaYiJSbWQ51WzBOUsQBt
nfbyh725F+rS91/HBH/iz6V+LmSwoz/LstDeS7WKO55pZ01q1Gn1qKR+bRMHacpz
EWuWwvHNAkgFIVboLjU78jFMd4JWmAkYPqLEQIhVq1UnznrbDJyo75WvedD6TIbO
6CroXzFVhr2mLleBe+VUfFyN1ljE2dytYAmna0wLrUTzgukLT1txJ8KMfy+d/18u
SO5suMKzqQqMcL+DvA4DAxNxSP8/Aa33ZWr52slXj00uN5TRHMBNk0v9lXaPTYpS
bFXQah/q/DRgMEGx3bLrc9B/yczcypeLeSIyTuLn6C0xlT2ibekUu8XUeghjauCz
m7kzjx0BFRcGoEuUV4w18Ni7QqQytsIIF0sWBiFmrRA8d7kSZ5KUwDQV6hj3Qmh/
hXNeragnPK/wYiyLlxOSodghwWOguWvaxiN6CZXcVMobHxPv91Cbyn6gokaLAEAj
4qbLKe1AOu80p7DIUDtKt+lXxYx39B37Hv2gAFfI3kxRVOkNDly4CsGBlRyZHHfN
8ISBN9NX6OP3zXEwmJC9OA6nQ8lCbH8cwzUUDUVVSeWOMdot7fk4ITHCWNy7we6g
UoAcAdS8i9aO1BFY1LzmibUoYsYKDue/oqCYw3/uu9gGtcmSbgHdHh4zbOaJQOsH
OzwQbXF0fovpvJQQsaWNlVn1r/rundjsCx6S7y6KIee44mq+pEVTNwy3VsXs8fMa
uzCpLKhvza4t/NUfM6XjMKmYsUBxwlyZzaGJqjMOG6mxgB9bZkehtcLvgROT4E9y
/WNkALh8FCZNL2BmkXe8Ct6p7xWxoY255Q9JYFtHvMgFD2yWSviXTpiJ/B1eSU+u
up4oPyYa1D/Z5t811HOUrpQuA+zT3gD/oXTfjByMj9DhAljoruNmnjTcYejdyPA5
nv4SDtfzFb9v3WVKrXw+7ncncgtb/8d6lxtS1XWdGMHq3BFLICTwbl4D+dwxlEvD
6RCjNB5MjfsKBBbEVeROOWvN/47VSydKhxiV7iubQIjygwIh7ZvpVams8wmzEFtz
qy01sqDfmMJNx1/oUNkZ4PYSNK8MG2FAPrqQJsdKzaB5ONOZm7+QRkIQwKhbqpBz
E4ugsmoUNq1rqNRMFtRprHsYPHwYuSoPacuffnH/Kw29Byj4U+0T1IhOfIpkrLam
2F6pyyCr5BEMz8X5fAhiJ2wFAhM8NK2QyFIVDSvMrI+IJ2AEf+nK6Pi6wcWePTw3
m9ObuogK+fZZekPaLDi3uo8PlFzHL5DqTOY80d1eR6sFEcsAdVpAEo/DGzlmGyRK
h3zC2ST4mZIUAfxRiHr8wJjB7IV2DF0x3KKWMKnK5T1Xbhy7nDlUqYCew0dqZZKt
6aLXJSLDeTo9Cqtoj5JjGYRUo809fldVTMOp5kh+kfc2HNWleAeXeKlkUMcRadjF
CVBwM5te2PfIO/Wx7K9igAP4ravgnAd+wLK5GnZ2Bw00QCFijARp8ydBgMEWzVqc
OztIg0LWh3okEiGdW6HSuCFWoz7I05HDgSHaoBaZxsofUZqMZGHvR2ZHPiEvFzpj
mcB7kPNXwTpcc9k7szZLahYCNZhnJPp+847VvnKlaajSrT+MBHxi2gg91pAltPCy
EjrU5uLdsLB8U1SKbrD+iB5vjoAC0XoiEfpWeKMQ41wfxknV1e6zw1B9y3NRrFse
G4opLshWAPgojGop+9NZ/KwDvcH95bw1NTx3ZTLYAMAlXu9Z7c+JLUhtHjG9hJj9
3SCDR6RlhOiLF9G1YU60zFdnvXzwuQKFRe59lzn0WIwX+9uM1x1IIuguT2zKotL+
g4Ppj9LFCJWzLNVSRcNOhLrZFGZm4E8L1nx5nI0oEB5w2gwLLV+dWU5t0rIYLENB
SPhM6H+OVcYsV+ubXxehoEj415aRerBWUOVIWOyczeY9HJCx6cZ3hc/Re18k6mJO
isobpQSoGbgCa7cuByFNAIpQyEqmIIPUsVDZHL2ZItcJXJwF2QdNPj+CWjhQj/L1
z6+FmAWe0E+9C3ALuynx8fSJF6E0tJRUMvCMJdEFHNKzQv2cYc2RU5cT9r7Ff0Mk
ThtGUs0x03dLvqD60LHKu4uDRfGbT7w9el9sZtfwsOjZcNkREzmPNUQeTniuWUpk
O3WaffGoth4ell0tCKuT3pb7FfOZRx5vs6Z1tr85SO4G+A0oMZlSr+lnoBlYLoH8
K5ZLFJK3kmzqUK+TC23+XmP2dMOXPWmUGNAnmriEZOV76d2wBhF/iJqV4Hrh7HlW
zZ1WwfST/0g88lE0HBALjnOIo5TCzzfD0SGwlXIiBxbrcG0B3B+1prJxi/uA2sii
F0VaOzyUcLzXzU6pHLAeBbmIWb1OGjzHWVYIZaHW0mw1Un5pBunok9DE6HcCGXhV
yWyuLcvQDPgPbh0TwPpSGlREvtT/OREHnZeLxjAHeuAB5gw+Sl25mILYn/cGBGxt
98kKbXz7faZOQ/kTCzRhwGvqLBECDPmZSBFieqCFxO+N7W6IRNsF53nZGjJia1Ye
jtYL1NJbQJLEtc8Xa8Ohg00JUe+TG2t1TzRQIZ226zu87vzela9ME1VAzj7d0ESS
ih4E+xJYhRmurqeNPGtPdwffLAR0DGITnTdsD5ORvmgilQ7AtF+4A7cC+QDKJ4Al
cUMol2+GfNILgOgxKU5aETRvfF6G1HHKHmP2nTH30OzWL0v1/sKmkCNZc+veyO7J
Q1OxU/iS33IGdKGKyVMTWUwZ9SbOys/xA/sk6XzaXHRJny6DHUITjKK6jasRwItr
k1ZrvHbRJuBMKsP8gkRKfUg+p5FFraQzHjPvPgcVL082r7tAZsTDK0/2JoqesHaV
YGL9F2aN7o0bxDES72H2DTo1poccrVA5u5H/D/snVKRKN4sn77OZuVvP5HEgTABU
vfYmqGUspTQ3KbWoEPtzegmt0FeVMjno6hiL6NtqGX36ePC2vHGl2lLNNLHYy/YG
ufyPqI9gKZyYd149icDoG0SiFdrkYJgFQ0MxpyUN8SAGmXftl/J3egz3NlQSi5aZ
uQ8Ln1QvRvoiG2TqZoJ+962COvygANHqgxoMF36Wm/fyVCe2f7S0EY7eA/4WSRZq
r8jlm/ZXnzLSmHI8DksygUtauHcgNWhT1wo1HxF5U4VXiNXGErqYk871Nq67fQ7y
6GZeCo3B4hUQsNp97UlSaZiVmfsYLkAcynmX0K1MxzbMsYLuIGcB+VFZaPq3/4eh
aByMyrNJsmXhFdkuaPodkWGUUlrDy/vdjoFEc+gTIoyvP+s2d9mAg5SG+XwyJKqK
/pgymeecTRq1lochHexvzv8owdGyl23BgMfUdMM7EhEVDJCoWpiMO3I+8nhKEQTw
Mt+36YflHxcbJRJRRFzqFJ5p5iJ4BLWqUlHsBj+CHOm8Y2IBOKohTS9NDlMuW3zs
Z3hxfTbKMZa0+k4mKc0/ERktcxlxynpPZl8KZmL9VDndo9Hg+DHTKRpRCfajh6Yn
qVsn0JuVELCjLCmktrgvgo6xDQvgHmDb/thm3k71PbgpzSXufhnG4o9cuLQ7nGK9
5725kTqAPDqVphMWt7Mq85zx+3N49uq7nQQ037HvPEQq4KAfaLoM7QVFY+7Ej/rd
s/CbwXtKbANxYETe0Gp3u/ss0XnJ5G1h7sWbREQj47LmpTUzOnhT6rQUXDvuvqxN
qyhsX4CGusWCnxtRK2fKg90tfPoarIt2jS7seQKrBbNk3ibT+yglqHeQFSSHL7BJ
3COo1PYY6qr3pCYW7f9P8qALpUmVsxdcJQtd0hVJF1lH61MZGd1312cO545pEXIr
oR4oYm7IKR3wFS4UHmMLzyZGDsL8GnL96b5vzKsx5iD7pWP28oZSBKqiI9dHITqJ
frlPM++pfKnIJO43e/vpaiWV4S2FN7iopjUW/RcMKmnqew5wovfeOdpNI+nENx4P
qtZJEJ2KeQX1K82IslQSqmbzGT00AiobyhC3AiUOlB2GwKxnXnceHx+vEK7Ni4HP
mNNAj40YPsyuhv4MPziBPpyOqrUpgdV1bPGWxzRcgizqG+/5ndTWwODGaBkl2SX6
NqFf9yKPua4ndWwaVLCOe9mFK3kE2ryLwtTxzE6s1BwjCEY9OuZKeSAT8UM8kxRy
F+TzdUpcVqPgi/ec/CEnvq98bxTm9cMTF3rYlG6fC/8lcMaw1KQfljwaQhsXEF5r
vKasWag+eSzLF2A66aCZJz/vY6+YXYedbiQeE6Ej3XdXwjWwJtJS+Uk3qE+l8Rmz
gfMN7WB8hNQBK8zj7nJQpgVT+PImUGDHXfyofN2waoAfSc+peCgKloiehIyzLgM8
YxA+RwfCdmHRe0VF/ewFMDlzbNh9GqmSDJcYJLSlrHw46Es2eJRZ22xjPxE+0q4G
nUE7rGn6EPATg5uZOJ0D+XzUCR3+T3fBZcvj+pr4VocetoIu6PRtRxcPWxo+kq2g
krBeRxahvvO0GDu+In32h1c4+/jlUEvfe3ViM19G4s5jKLCAm1eXSc4HGjk8MqtM
EEHBKtDOW3N+nEvZg9XuGWaKe0W5b19TSnuPpeEIiDBgdfufDW0LKzgdnJWQ5Tyl
i70GSrHkoM0j5FfrDOnr4avYW5948YzKedAyn/8RDUC+Yz74imNdf6WP1vBQ9V0L
CWQ6UzCnrwS33AeH50iQKV5pUY4ds0PvEHyi04WT6bHcDkS6nKp2kadOi9bCrkB5
Rs1YBRbGAz3sAoMqKL2XL+R0SKa/ccl7+jBhBML6ntyF+xGE1uMCPdaLeAwzk7SK
xvOKypPkx+2yeGk5xIjfbzuCOaexTLZP3KSTWL11ftdHoDwk7/FevqcTEyL9pTnD
EN6Uu6J0yW9Rc2+vqQjSFa6i0z2NZjawHssXDE3eLYiAIFpFBrcqv0c9a47Tj88Q
ayBn6ssw4OkiBeLWtPuPOYiuVvfeYUdkNbWgLRlx0SgcszJKt2rdiAoWNg5am2zN
IrC96SBURvgGJBDOQQJqq40rZ2JnYbM3j/8jquKzMukZJnhf09zvyaCvasUbMcWb
HTNJef2/uGhgh6iFPDiWe++MtqoeKjyDRcc7oroZ/8TFDAQpaSLrv2gDZ92oiSyl
XXh0JWmY42aox8Uk2eCYVbzepCKGKXnE9SmDuCZhm3CWBB+HwXZowqoss2jWsu8T
V96IYmkt9F5/RRM8mLZhsf+MXEYaIxEVt7noIMKJVh5JMTskcZclfrL03lF3+VS/
nAl/ppe4mbExZkWawybOzittkM/DV84jmlvK+4qMNmAMD+Aw3dT6/tHZ5VDaImGR
LfLT/FFgD1Qenm4Cp/2Vwz1wVg8ftPxMJioReX8SDJPWNTmaI2YipnRy32ZqFvmp
F2jY1ZCGw+m9BucXg5HCSuFqDUShJgoHLEOvKwb7gT9pla6lpGstW6gDHdFWeZ/9
IicP/jrJmfzmp9rgmi4UI8+PAUUh3f5+IdZN7hcPd/i9OCYvn9RHOC/QebslqbJU
Be7Ts6/pOiElc2Q61S0LGIgPY6Z0Kwdg1t9iroVF1cEeal1aHCPYUCCE8lRL+hlE
sl1H7R3YBgb/HtuiRykEKl5CqjwxmWaCdpH/Wgja9l/53SludaoTiBA/DYso2KMS
nAaALnpLFcPJ6maWP+3thcKa+ioBjZkIghLavFhAd86qUXl/EonvTMCq5TLeGtiK
H8GILCvjC5j6KXU2vw7wmzuN2L4F8iekPeYFO3oZqnOG0nvGx++twJseiG/ncKa+
nM8rADrSoYHTWa9oJqjUrjASjkQ+Zy6zlR6RPWXfsJBAG8mKB3d7HT4Cf7OehXMS
+vgPSfddqPTVOZiKYUbRJtQAcjVhVdXoiZE9cpwYHsen3FSKG08P+JZiS276HL8H
pYKJjSz9hTundDQCSmGqcMjUwhENJOPZKTVyAQDI5FWh0gOa4QkCIHKJbdyoCqDU
FnU5n6g/UhreLGrNDRW12z4Ck3YlsIGriSjI9Hz0ovo/oirauLTSWe51z3dwpw+1
2XfyvaG7YR5qtH2vZdNKWfQx2Ro4Fuosxewz7VNJiOdpn5kYFUYoLq4cL+tPTK7l
mhmevj2RLwBcTl/57N7fo/MGX+PviN0jzs0OEUFqxWvLQugepoUc3SbLrDgbrhN3
1f2ulzVR8OWSrFnEJqQtkI8y82fKK4GyPyXkhFVMvK15A614jCAb7pWsLJur/XUe
Cho29Dd4g5sGComSRBeYU6EQKwvyk/yfQY7XfEF5PFDHu0Ci8P37yiL2XkmxvvvO
IDmU0ZhutaQ0IDbVKQRdJUuDGsVfQHneaWjhrBNmcbW9GwXLeauBFmx2gFExmkMg
h3H/YtCo6eSq5I7ICllepNIvy0Ru3Ns1CascrQsSYmltUA88AYnaSk020XFXwLk3
NXOMCcYLHVATuw1liPbK7+MtGXTBW5h1/MMiDRytBqJ/kWevJmJK0X/A10FRIrdl
06mTzBmh5ZjftcK0k0hehcWN5GumXV3nnbCow/c1/MSYasAhdL5V/w/6YFbz0r6c
fXueW/CjgLsZM9+9fdDYIMOy46H4acVFsmR7AIF/8lTYwy5Wyurp6wE9WL/dZT/t
5ZY9kaawImC4KhqI6vuvI9snzm4Jc3s85g8hyl0uKltbYEl+dFCD2OkT7tAx2wrq
mdS7FzT5ol5F/G/6TXsah/kIy8iBAYztF3Y6VeuPzHTrn62Wqd/FNmumtUY8QP4D
Y0bV+QLmuPMi3pSg3Dum+Ykdx9SMhUiMgBCLu3LR9rJgTzYwYSUiTQJ/11V2tg9N
ovVQEBh+kVgIC4RDHGwtDBmyYfBZ+Vge4mV7x5KpG+Cm+J0koElcJTeu5TgA3Z/P
bMEZ1n62pPY2fgNjcdYFTUTF5CxAp067cqDTktvPp4a46SzOYTqTswtebWgBKlJp
VORoU6cHdcFb9olzNC1hVNrCfVHHk9IrK9B5J76rcKYePzgqO7AZERTUf2/kz1TD
kmrqwe4PDf28mdJZIcO5zrNwqLKUb1/Tqat1t+D8LuBYwjnqI/XW7rj1XDCBQDSW
h6kl0CYAwhfr5A4JAU8mYGl2IcsEUZ60JzVFwbtcbtcBT7XDL20O/L5WAeAW38+S
MRG6FJZe7W2zkXF1/p+Z0B4Yiifi34u1sEFYBvFtfkavXV12mOUaboYQqp3orxjK
pJewtUCHkWiQ+kkb6iSebW+i+zbV+bU7oghLFa1amduo2QkaOh61AKwAzVDT8FE7
PWuoEoSQbdsp1gq8kFUaMX0PhMXIWLc5xy3Szt3Ow/3i4+lM0h44bIgmwEfb7Rlz
js+0tiyrws5n6LS6rRnH7ojQC5vlyzrHkCiTGvpVSdZkt3AppgutTbLT3PGH6qKe
mrzpH1fIJo4SNk/Mam6y23vEPd3PWTzBbtwm+ntXWgLs6pzBGRwGpF50GjH3Yrl2
/T71T+XKCCEQMRtcbLmrcQqUqlkKWsENKuFjCLgKDPPTGIhq43H6n34XFgYXcmjK
azR9vnbJbmXmMIpfRcoeILrUUaADc9IdWgJmJhe3tVIKyAAvzw3lXg4CKLRQiq+R
+qbkdvR0lJCQ03hGjX2fIRVr3Oy3Ph5WGWinmTm+oFi60sx//P8IV7B1RbKa94Li
MDbfO4g/c01Ntc9g9DvmYZvPvuUk/I4ZC14RPZS4ScxWw+UqsLpPkTkTbTuCMKkV
SpekHN6A3weOYMxbm8qwkBwF91z3XB8jJiD7EzPYjuYXrE1RaCkGQt3j5NUnmj9D
rSeOC6eOe2wg59qx23iTYMKlZxNNAkXJ4WXqitbfhbay8BCJ5M5I3PX/TKhf4qXf
gCH2lGVJ4p3GTuEsMCyC8waKKMF87xgXYZekWByfsz2g1NaLgFhdsNoKuLBaT1Zv
tkpYF7okQWRXbuN7oJ09TfGLB3JsWgq6ahS6GtDsNFLgSbL184GKniPC/kTY7rPi
KxE/Q+LVeMZu02U/xwzZthX2RLw3Jo+sqkssGaGpk4uKcEh7x84WyQsmSQxKfQhT
De+ZCgvp+vycl7nW0eYPqmf2PgA5Jab2NjsWAvHYOx+Vc9fUgHRe0Tl7rwob//kK
wJrZJmn8AX41AYHIdW77VVk5T9eA59c3LaORbgSiQnOkJDO1o6W0sm/KDWfqDLTj
TxKV5/MbmRX59jcauYhRQ8LBXx6xLu6j+P5IAl3gG1a9/fH7V9GFj7zV9YgZs99i
5NJtfqIQPwxEZr40BFePdONL6rCqj0WkyNfa2jYYixWYp1cKQjWnhJReptwLtXh0
fljwlQGModlEE4fyAl9XFHWgcEbjtUD5N2rbclPWhoJrZxPMzgzpZUXUbgQcoGbO
8BbojA7/kkX9Clrkg6m3KK5sajy04WPs8lB8QvpXZk6135/oHPxc14HP0j+li3Xv
73pPyc19qUN7C25qB5p8q0lyAzVsnMkqOob3w+fAJGYYOxgOutPJDU4bSb3Lcr3W
dNUv6/46R2VmKqAy6OXSVLhxOLIwVHekeF5VcfdgQLuSowYd84u2tVFETLLoASxC
se0v5a8Rh9Iq/TZGI0k0jvcL2R74mBuOVmr6YRUOHf4Ptka+osHioIHEWnXxEuzQ
MNBc6gtFOCBXXusHIMgPDAYJb6ZWTYs8d+wVtx5wCLgP99SSyb3DxY9J6WRe1crA
KVFRVd0hB2DulxW3d67gOcT8YQCa+gXIPCB42s5qRwSixmhX44BTw6En3HcG6nwo
SKNqUqIdzcUQiONoev1eGJTBUStwDLTTDypeIMFeSqLrUcDRweDDest4lQlECQor
fCnMwBWl4B8eBrBbnguFHfu4osluZ2Xh8Cet72Pf6oQFYYixs5m56T7rZVqGN3vr
cX9PKqRE5rVrnWX0epHq4OCxUEnj4KVrx5pjnbBTsGuv1943Kiva39OyjyEt7fq7
b+5bEjMrDjcjPfcppe6Yh9l3gz8ZJ8X6NifEymQ8XnhUfGyPodwK0z3GP1UJNcVs
cA99dG3UgQi4Ye13sUGJ/bnMDZ8iPokp3rPamaANbMfb/8xZSyH/k0vqpKumwo8P
NSk7c2FUFV8ZnUhF/XKDagwsV2qYZEDzT8tWAQzSkTSrSW9IS3DqvIN94b++PPTk
QQrwUCC30YtbOgAzUHs/dQC6uiKMckwNh5NzNDGKfQIAWE+IPWN7MuUXlNIVI+SA
bWaTWSCsgDmQm5ShTbaCg4+Rs6IHkn1848p1yMF/IeWXfroWxSok4yU/K9Ovlu6j
miDq7NfrSIueQs8u0UprsvV0cOlqaoCdwpVpkwEYT0YzdrhFKwtoB6U34bwLEYrh
6NneDZ1aALS00ikC4z6nUbJJwGgRntSIlAYOu7ReFz7e3judomjMeZyXdjrlNwWl
OQqdKVlk4hQYSBDkerZiScniJsPtnoOTxBECPwk85BH0egmwy3/QctqzlMeG8lWO
R7heSRkY/mfied5v2FcUwXIDQWpnS/GIjL5GkFLVq95WuYQtXjKwiOvTTX/X19ST
brOGxhKl/GWrPwQhE6SLb3Dhhuycvx0oDayYxsKeA2ehAjVJintTd35q45x+pbLE
Y29qMA3eNPUuQyeCjB/diAs6dd6JNS+1vf7E9K1Xsyk0rduR6h+qJrwdGoeDcMAW
7pKBoHzCoIizfv2ZMYwovPIc24g5tD/9pc7+CLlGInHBayEAcqg+PxMxtt6NcjpH
ROf0fGsciQy2/uA6WmVZ4snv7B9w1w7mjmxqfCblRhNJN7q4I0VUVoqCCy2YYQWS
OpxUfwnVoOKw7jHIgEgSzbngX48jtJtN63A4Q8Ex/H9I0UFcVquB7nid2ty1PPDh
/suDP034m8UNtksAidmFDKVtVQwSx29L71zVrFkpyJFRzJGMGuYFoArJUA1SRUJG
r0Xmcx6XBoKMo6ifkLp8b8i2wjR/LIQk8mn/kyo/5PYyLF1MusUDx1K44WsicnPU
ozcyDVmemV2XkXhSRY9GHYT9P7kpQSmq/FYGQtAapxIsae9YASCJo14YGRnIX+hr
l0e6op5BtRYVGwdtuSQH/IhXePNdvuuDzVH7/clDrAIFlr8B3NqPSLc1cK1g/efr
LasMsn18B8rjm7BxBoYkvNKirjqCoim2ZMHgL54NGl/y6EA/ZEjNTMS/RLuJ7+F/
YxRlIBTwVfyy/HRBqPqTBVpY90T57RDp0+OAQ9oNRFrz/YDoOuS5+RJRAWt6Cm1c
OuRsf6Adl+UOeEgl9FrfqA5lgK+H1E5dbs/1PTsDr3zqQ38gOP/nbb946fZLfPcG
KKxIAqsr3sE+7l4bGfw+HStPnQJ0M4WcAyjuR5h9q0xHi9AFY+XiqrInxEMuJXX+
v6DTCipxmPfyYGpVzg6yL7TPgxDdmFufJWcJFXxBm2CV4h8SJejaXA/n36LVbO4K
KYeg1udS+CubDdaeonFG6OHKccrw4Qh1VPTJID73grHhlf7ThtVhoN/etTlnqFTp
/abmgxGs2QfRfE9UDEqqA1qZv2EMzfF5j3xA3TTHCIS+NWd+V8fPLSeDzdLpeaC2
sByquc5DaWTOhn4qpDxCjhstxHX8i+Gy1llG3ClHhYodsVcTOtKH5sQWs2zT+Sib
0/ljcRlwpEah2LrZqfFcXhX5O/yIa78lVc4cWOXjO4VgHS8CUZkb/zjaZsqax+rd
dRYTjedFQi8mTEo+o/as36hNSR82NhBOp5m67ZUkSTxMLBczUW+PuYAQZoO0yGHd
JvoN3nSVBHgHidM/GIosFlI228XGrwZxz712WrtW7ZWOJs2Es7X6oHSP6dwlfSUR
q2IOj0E4rSvuU50GHSW0ZqBvRQMmQTOqrxS+09tWLXIZVkrJG60eJTjQBs1YO35e
6d5O1csx10zDHh5J5vn+uTPDEah9/liSNviD9NPy7D4IUmeFFOBhADDApNuZ4fBM
jiQXnBg8INEk4G8bxEgphosBxQDqKThDKfNxHjhAai3pavD3K37WAw49vDcbceP8
RNasCucD9UcaC3q9eyiGigSiG6lyWeqgdN9AOIaMCm7FS/1HaDaQdh3BJmK5NJ0Q
3BQQtGTWVG+nVPYGQJFi/q3dLwLq9XzRYo4hFBnx2SdPsskScnwhUuF2zMGvgI8+
JFVIkzd41xuRFfUJFzNWUhH+belxCTlBSd1jKTxLbcY1Rbu/cwQGnOJDF2Vey3J1
/VwUp6daai+hPw0lrGBBCZLfTaSxuTRh8s50HTiJY8zt+SFi+p3uvY0QqDd5Qwzw
Ogekt2IZFIfl0S72TNXAfJi27Hsp36b0nRdluES8LJYnE+eFgNjpnOQYGqjq9Wn/
k6R26qK2jU8mC1z/wUEot4JAvdRqJirh2vgoqd4OJDV4Yd2jcbUB9tysD1oIX487
S6QrecYcswwGvoDH1lsd/YEYiVf8UAl64GH72YJlQ6mK+u+Uax0ZpiMZui8WXO/s
ZW+X7pgzLcAKCI+A1EodTKzsw560ngj96y22/TQFKAIyqMLdm1Q9k8NcI1Zjt571
gyhNzOZirmU5rXyX1aXVs/+PBqJKsa+G4Muh8MKJpRafSvn5gZYTNWFPGcYItGO9
FSI1Hv+T5KkIDjY5mA/YM7VP3Jk+nkG/RW2fMIXE00R/SEqeLkxkP2q8AzzGQ1O7
rxSdZnwoN9OU9sPvcjRTc/HNAby4l0VcR63ZKVbQfaGO9KPCZrGlP2+GxHZorVML
NjPJsxfvzhJi7v2OcpBo0c6VLbCgFre4ylFzHO0ZtUGVw1KBQKGqOW5O7+LeUZhO
vb8wb1UDsokpz3gWs5/bbqJob/BKhHKZ85gKcmSHE6w1/CyeMqnEcrfWj6r/zNzs
d7Ua4WfxAqiSNcaAoyhQMWGN8CwVly5mLqonG089jwkJCwvkJ6WakPwju/qkV+7P
FC/fiuXncMSO/lTxvKr9wsSOq6u/myI4VysaKNZiV5ezWnDpzOuAVK6a1EP8Ok6h
P1iDXH7O7IlgT33+Azq3YgZc9MH1gVeZclYHI7OLc+ResK+vnnN4w50/Zc1+rpc8
PD+OslMrGZJw5BilY48nnySjlpDgbxoNRHN1dEIgq92Pc7VsqECJ4eidqh+S7gMc
TP8h/cD2kEEypC+C046Zm0LvhKHZaCJ1pMtwW24THmVA5hWdJ22YVYXXTI34Af03
x0iu6gS4FFzJ8nIOMi/l6qXtPvrzwZm9mBi0mKj0A0nrmJLbQE/ccg6QiHOK2mnd
dLyow3w9xk2hCMrGZPrJ8VCerXVYxsHRoZu3Nuzc1/6TcsUmk62JqNUqhayRktZ2
vcTz8mKkebTlJe9oYSus7UkWhuNUgo0XzWW2W72EsZa934I7a4uo2iTYsoHX7oCa
sjQDX7LVwmygTI/fIH64feLMKprjBSL6lL7QP1fsFz8YJN/rVGXuMLUdnb5hn2vX
K29RpOz6lXcCXwn7N+p0JcOBqlZdqpODxXtWHedU35RHXXcnOJth8GzMaNU7ko5G
LNw/9u3EV1d/+EhhMjWI8MNDLr4hWMBlJVtY9RkEBQ2294gPDIlGWu87FziwWHGg
6vxBjx/K5xqU7kNgzZ5pzwwBmV63jxE1eGOglldGC8fOdpohixauvm5+ltnV2ei4
DyIyiW4JeEKc1PE8jYn0BrtIt2oQoviNr/rzZXTm6tdekiifaK5SRCdwC8Kp8aO9
T5bl3M65IUl8J8lkLkG+RG3fazEn+pLc2/aAhyFAd5b6Qh5sU3M100NCYOb/13Tp
fh8h2j1+iFv42LiJ7P1s538apWtWjZXT7L5RpwYBT+cxf+zeO2iR0kgOiJJyjB5S
9ksG8ga6fKBMN2urN7topwHI5hcS4tjx7txts9dWb+YrsG3HnoJQBoROPzpqhcmT
LZTHLRw83TyT6pXIPhGEimUlP1FMZtuOc5oqKhi0jWSpk9m1vyWjK36yj0GPgYvV
xTyA1LHjYlp0q2aCcMUD3PvR8mejaf8sQbRGcgp+JjdyHw2Guwmt24dcVMtA4Ojz
wmUGbDTpk8Q5HE6QcvZQ8xTs5z8N5P96sajD38fAUhOIDa+xmmeDCtf9jc4XUe9K
t25OMkq1ME6LXvCKrT600gcVq/pLc9Z5t800lUyIbIRMp9InkuuIE5uAzzPbEJ8h
dMHG8cW9eSWsIifxJLOZptf3xNR0KvI59A9eys/7leNV8MX38nWzKTG/v6TJX0Hr
IGvesDHTbBuYLnp1yOYb67QS9Gey2Q1Ihfay09M2oggs9p5hEYk/xB+3YBjZHrMm
JGby+aGK77K9SvwET8LJTO3B6je1RObCSBWaFxDGvUE1aIZX2PGsx4BXrrU8koIO
ZIA9YliHOmmrAJn/UPToufO+BoB9VHpY3OgyVUwC9jyzEsRaKLD7r4IEtNhonBl2
0KkbTDDeyH11I3HdAA91PS2JX0AsFQBs4s7TQ9wklk4vwi1T6UG/1LqWzttabpsu
R4T0k73vtpNiymStogIXzL7SHwSNwoyzTwKdBFisvCqM+gg3j3lLeipqwePJUn4l
jLBZSrpim8DaFgHs4kaZ/wkuDlCX2MERHaYIyYj0qfCVonhRS72U/mTPBbgcmRD4
WnikGvnJgN4xiCrGZ1UsJmJdsBYuDRBfIoQrsLPd8nsyNjAo/yT4NcuToHH13s9+
lG7zq5h/dkFIFj+NgG0x1ZFCSn4MSwy++I6G5OTPMgu3ozhIn0ThjhLR86BW8Rm7
//bKkUjJ2qkq0dQC2tQFp0EwUDBWtLV3jbE7wCb2Tti/WhAQZzsvrEWsajxv76zH
nDJCVjU85zPFnYLe6hLnSpi7/ZAhR3Hvib5qmwF2kiZxHcFhl5/ulJPozVmD6MKx
5V3ee0LrRGvcDVIe6kdXfl9MP+0QgR07t1wJ0LpqYd9L6oHbSsNEDjqk+jVuxCRN
claj4ju/QQaV3g17jTCsgGUfq4eyM6guaQQZB0ber+PsAgjprjHdQipPvrvHaTCS
TbD4jND8SHrA2enQDqx236Cd2+7DvqvOfHDtWcX5XRIS7QFkTpX/qu3MruvvO1jB
tDzs+NYwe0ca9ab2JrMwPwnsQ8yYURqxDbiUInVHXMX5gWwHgjWrsdrY2K5Q7Dxj
ddMkJ6uOqUfWkTw9MP2UKyYaXctvHPlttltgKso9KU8ySpeNOTRhAoGojRJz8u6e
g5fQM0xmvUwZFIUeb6K8IYTaZ0SGb9Q6m53EOQJzUz4SUbmTdW2TJXsMOYHqXhC8
QULlFvNsRc1TotDYzuqsDpHXYv2KdyitJMypMMOKDiNUsrLRc21eTDMSfSuLr9ms
+4qjew7lqXUNbdQGW8TYz53wG4FzF+o/zjQu4C/POMI0Z+ML75xG3tz4W8YJfyVG
+HwrhV0HJu98Y+4dZxxigDLl5WEde0O2M3jTXIeyl5jfYxTWN6bMzIX/euQ7Jix2
ecDWSPcrYTq+VW5ivbutyTxwjvstG0zbWEQyRtCfHFqQa/ra2ywZczEepMaB4a10
w8XlZdyKQ9U+cGzI3tjdDzXO6OuYHCn5lcOClmdL7sRY3QSOT5DfRVLR+A8f/mMn
Zgp2Hg2uiS0XQaLVuBG8PtvL8EHV1iFBv6tDcVyAwLgUFjEJR1FVs7+ew5vX4sBx
GbmVTcTTLcdiFwin2PMTwNQuBxpDSsoMOYglnej7UZ+LXuCgAiSGoXX5bCThrbf4
WvUfhCTsjTyWYLJqQFaM2prJfBW9YjNgyE7p3Q9b4NtYzjDWZb9Dxn2IcxZxXO69
cX5zjt8t0O2ZVFPU2PTLQq9sGWVVV67I+PAxuI9hw+gg+xl3Q809r27g20bUPcfh
egq06/JceAM3uK+KALJqvscgz0eMTU6OJAFvz7Cy7rxkebQMdiHf+nwtnYXIhu5L
vSjWAMP+7sy8TMnJ8tZN3OTa2KjWxYcNpP5JBA2acpEML1IQYipb4NzFOCm8P7PY
/yYNyKsO+z95bDfsR5VyRuUoa6OfpGYc4FJNeBcyYt+vtqYwUZPnoa4pZTFDBOVl
ERLYps87AMXu1bYhZcCyMIGBVqD8oyyb9Hv3dtjRVmb+uewfiAyMVwGxpDLPd6FG
JvqEf0Q4Xh1JjOYVU+zqaUcaFV4bhsZzUZfWyi6Y8H3U3mqV98aa6xpDK2UUTYEB
msh68kfZUHsw4HQs6ar59YwFUsz8yKyzx/Xp7ajV/ilwVxvrwc3bWHXxrva6tKlN
X/TcuiqJXIDP+O0CH9TzOenN/aNjT+l9ua8jNegOb/qDmdkIG4spDqGOS21sNTAv
R4PQ/ZbLRr+BYFNDcUrGVCwDxiQDowZ94MvpfyUp8vwFuVWmdSlPvmHlX7ID3Gc2
mU8GVDYM/4ALpq1DU4ZdSmmKmwfzAvI8CYzk2RXUnRaIQKYTqXTBDFnER6KUg6Mj
sGkZ13UWvwTzyJnCk3J1PNKTHTF2SaYu/paESvK8IOSEzdFJ8IeWSEOx36O8spbd
E83HEgXHx6g8Dw2uXMXcJzC1RazjcE1a/sW04urHqf+7DUpTU7zvQNNie0jtvlTk
olLCluOGYc4AdAhG5rb94cQcrTqBXBGLXi7bTERdRr3Or68UFTOz37y+vCdfma+D
k/AMXnw28/bFr+/93KXiF0rsbjCPoDlDqw3zMxJqw7h3vinxvtDRpXtFSqamPAcu
WoSV+I0jm3P8tl9IxkSphlRWh1YD5AHGW85x736aEj8eWaMSM4Du6sr4hHgzj6/j
KNs85/XKEjssZS0S4J2qwtCdJl8HE+WxqgvbtY1XWEUDR8VLelywf/aImu++n69J
luR6S8N5ziQK2Ca5GCajDJKz81lXULVIDarDVc53kheA5co7oVsvPKb+r4imQ5BD
uv449T09sZEvFFuY6yCCs/0hfFQWGtIxgsUPMfWW4swwCjh1+f2FDdbtY8FM4S9q
txJCiShL5UyCsmWRFhbagz5wEZGonxbO9VDrR3cEqKQ55Hhv9bvSW/bDmmbNB1h7
HUGJMj1/It3cXJbZn0a0e1jVmgMAVkq1MWhK1llId7alMeCkHFnAfY8/kTaHAvF9
+VHbqfNA58A5DMuwa5JG4MqggrlSU/WFQfo0T4yn+6WNTUesPUXL61PJQ9KJh709
RFwSPWXV2ixqnQ72GnWXkUVfh0Q1CsU/91sknmNYvQGIb6zIFxaPX3BWFBmHDUU2
Q4sqWbExO9qso7JhviadTIroFX01K2jghfUbP/p47nKlqGex6n7j+iV7SP2dgRrR
SCL8b3yMQ1g5/800LKEO4Sj6scfk97COeJq+YI1V/JfYWbAa/0sODHlwEo+ijFI1
DDR4vqjj2UfmX3ndtKKSGqCBgzXacOfh6tueVlZnlm6bqasffbfvZpBIFPQ2DHt6
CZETdOftR/Kchyw24ZTFx34e52ya/ZWmGSUzgZbsarnrZoC6+xfdiMhty7GBrEgs
ddJBpja5bGczQEkYRHSYTafuJXwfdyvV4tjpegflaNInIUxg7MazNeg/ERWoWqQF
H3pxu/IMALWRDbCdFKEEO0lQpr1xFXVuUzR+AY20R8BuX9rH39jjjbytAPg1F+WE
JFVAYCavwZnHSMwqHyD/72rRfZdQCJLzP7uenBf01eq8oJASQhaQKF+v2SDkcHLw
YxpkfSi+UreUK/WtoalAULz00+MuI7Rq4a2NQrStAFPNocQvXQSTBoQcHW2nR/wL
O4lzPBosr+1paS+zCBnPn6JlfmZ58Lah1euNjWQya3VxbIALUTJu42lssKWyIZIJ
S+UATc9DLHwVknETaT9Mp/7RtoFANs5gcOU2sK1LbZWCEJ/IxD8eo2OKqdbVIurn
hJjjK7V99qYjcOXOKKQHwi3uOqW10LrxoKWrdvWJd56MbR/Hc+CSDv4kSfgoTsRy
e1EGDS7xZYj2MH397vu7JHBvXN3QQNEChvh3KpAP4bUgUT115G6wxmDO6ng+VLQU
yXwbsQvi3HE4oYuQ4LbQpwg9lTep+j4BXFSKdQd+Qd5iTfk3JWoTPU/IU138fyNG
nEcYj0mS18QYReBkA3wS5Q69wtSLiv/PrmD5UqPg/Yeta4vamvB5uxe2XuS+4poV
4ymczsbZXBZy5ulK7z3hg3op60kd7iMH52ca4e6mQ0r5X5psACjT4EFcVbe7rHUY
8CWHqpKzQT2Uud4yJaaGC/sD38OvOqil+L6u6PbjGQsKHpqj+AYFmD1cAw3ZNWoh
S2cD0qDu+wO7IIpj9Ey42eg7NRaZ3NWqIa4LcggD1qF0pKw/g1bGaO82S6cNpPq/
F3zcuCzdWotZ6wMTojP8F0dPH0xzr4CBBFVXRWqK8dM7Mzp/AhdNSWBXqRkaua/n
a55uemcl8wkHBjhk7RxYY3pltwMgP5uNKAXHZ2ce1K4+IzGzOMRCk1HhpYJa9TOi
xdnDb7wwlOH2mL+QL9Le/wK5B9hoeheZHqTzkkMmbVUhj6emqagCn9v7pJpJ5lBo
x0G6WjWiXgDa21/TBXPNonr59x8IVP0PxrTSLRUe73tTd1mT3Gl/or5Jo/JtPolr
1oLjm2ac2EFGlWq6Wks2vFxQphqX4gWMXOAZTrN5mHgDP4c5VUiGsb5HWyd6xdKV
+dEBQXX6WAjM1pouOqSKqBIOVooQcnLbLfVbuOy+/ssymdIeoXDAUedl7Arw8UIa
V0QqZh7wB8ZwNLY2kc+1zxGQ/qj5H8vzetTwegfvo6tVPjBnk25PrntPu5NHkqz3
wJbxnE1INJ49sNDQRKSUmWlzs5jxyQDCIwcaaQ+q6qPDFycwoIAWljVpBT1OpIGT
3tkkmS/K+4D/D6+swPbmhKnc3Dg+GhqbvNuqTNhazKizoLXmtoaID1+TzdUJDnG/
ezq+DPhA/y176tosIN/ULGqCtaiunADyxbz6idgf4FUo6Lhyqnfjl7FOkf6B1TXT
sqmg03Omy2BWfOmS6JvVw1vnWFjePe/HZO1XPP4/mv1V+UTG3Se7RyA3nxynUOSq
+/MlTS7puJevZF2ctubfAcP7hjQchXw3O4kfpcWRsg5u4RDmK0jQIWKY0UihfzSF
ku5lIXy5FlntKPKThZsD9/JRRvbkEauI7dAe583gNMNz93jk2/R9MQtFO+e976lb
PKeXc/tlh3+OW6OxYls6mBbPlonrv6Fwx/cjG11JOKqRE6DdA2H5gvx//Xu9WUab
PkU9Y75ZvUAtkFv26PYVSPrNR1AHQm8aZzDe7cgaEeLKokpUc+iHjF7+SyU9gE1n
forimNMfVqRm3ijTT+u9EZ/9RG9L35apFM4hjW9NUTt49r/3ED6hMr6rfGE9C63P
eopkJtMLwWV72WRkOPFVTM6l30nOigL7ilxSqXIxkxgIXV8JAQ8+Pp/BN99PThNG
4tPmcPUjPhJAEgEHZ6/iKOhnx5Fcxa9vaKpgqRitW6NQGO+KLUk6lJ/wPkM2kkV1
3Mt+BLdOJqbN7HS4NpgrULibJ/Hb6xE0J8hLRth80yr1oyUIvQ6i7/5btMAtKwBj
igiyeCU5weN4/o3AdXZK5E0y+o3Jk/9nMRaXJBPUOHhO7SgodY/qJoXbx3pdOWAZ
6z0Ug3PgUNWuNFOOKTGLMQo2H2A5/5ZlzTuUvwq0yzF42UMYIbbAMGjB4Rk7wlef
6/KTu4l6O2yXcWhnWVSZBVvw23EMdnDRWRiKY1alxevSmg4YODmHpjRJQ3um+/pd
27RxU6gXQUHnmfuiAFaus5vwcNxzt167LliXqNdjIn5YGe1XzPLr6WtvqwMMTv5S
rFm1vHO5ADnUem85PAFUD8sCQ8t3Y69LrSb3y46D01HECusX10AfKQWC63QMnXeP
rydBgLbbsNSAF2sBa78yKO/TIg0YqnqDHhsWbRYmKlIB3QF1F7AGGLrvL6n3+m8U
ghoqeBz2lr/qnBMDVvcgINidmycbT7Y0xiXbsia8FygsD4h771rD57hgKc0HkJws
gDzmbpS1bCSCj72CfT4Qr80ThYeOWe7oTBK0xj9Vy9Rrb/M9huFwNhHxsHl9d82r
dwvMHxyOGX4Dfy2muDk2X/kySrh0Smsevqwb6ZOKHrmPTkmHAVUqwDmZrKyfFzsU
4ERjm2J7koq/l206GQMECkaaj3vBCkz584btlD3beKb0ry5hObHl26NKM4eXqt/A
5Ug9+AXE35LTfh+xshMIduvXXx8+fUDkM5wi+Vjg8uKBfj2zM+t+lVw1+tMtD14+
ga7D/6v26GxPAmjBoPQBRXHX3bDl9mWYSlhXxfWM7I2n6Rm1CUiywdURfrenLenS
C3miY0XTektXih3z0n+2ACxzVNnwkJV1jxmPm1fzg0OZM4IECOh/J3RQYWAQOVao
wxxnMwzUZrylF3WD2D4jYpNe0wRU029Tgxdj2Qd20LU8x1l9M885mLUbXGCrqLVd
INB2C2nvOuWrJ0+fxsD795TOPYMjer4yMS6kROTzH05/K3oueefeQbmlwPtncBgD
8+PM6aHZ2Qk6J+27b3FrZOoxVg5EgzT4AeHl9swsHNoSo84Rau7bIvXJhQrzHo78
Vt+EWxFUm+DkBroybumHPrcknfyglTSATnHWeZdCVa7//TuiVlgxD5SnnCULR3Xe
WS6X4DzEs1HT7oEaq7bNNq7mONHO9nQ9XcIfF9f0XujHtKsS/bYrNOjmhcU42DMK
+DnLPR8Hb+3qMlQmXCWt31N9CM+au3AklapzsRlMogPYEJt8/jGJFvqgAkbbhHA/
/lVX6qhn9pP84eeUWKZrwa2HHg2rznK/g616xW1I0RniDsgIVij7gXnTiOhA7Vk6
CS8DIp/5biH/68nONjmUbhMq01LyTNkjMESK69qvnUnLiDeu5hvLvvNwyLAP7S6b
YOBuB7aERs7xAvyxQ4PGPLF/iX5awqGIg1ZBEpKD+PZy8aB/aWFNr2Kmqbds2rkF
4RQcRQdsod0T/Yrrh17toYCBDRbffVb1aHSTxcual8eKXki39cNkwFceeMx6+tez
YtT84njjy/erxJlCoPwWJ9a2wS8IS6vTFVb3zfOfR8af5X/1zf6VtC7oAROFwN/6
66fTARc/StZqVoUylomm0dy/KJgCq0AOtX7/fL+OemR15pck8hnlEA/5V4IFwimS
2R17YEqOvRw7pmT392JLsbxeAUiuwNOJWlBdkTtVcf3E8NKd927cIZjwwsuY8Q+O
HNcwnpl6TvVHrMjjLZmkYNhFMF0w9x5tDSxvTT34bWibQg9rSebvWP6sf1sfhawB
Z35y17Nb9w7NMbZdcqJd3yY2CuE9MAzht+ILO0AKyOz3Ou0QisIO5E8c3mpfxZAW
/D/y409h6WTAWvoyfA4G+OFDHagzWlPGnjlqH0phP+6HUWMo788l2n7jVbF1MDnO
dHS1liryG5w0AeZoETyPx5fyam4rOfClrJNsUVZSjv977r/HveACDyRqcb8DBSP0
fMN8nLGJm/wIZzvl9tggYeFwyJHWLO6DAxvWr75k/VJ20egrzuAtWlZBuhXgnlxk
WxGkRdPmZG79ARRwsA+kgwqQsXFoqE/QVCoCOeDQdsYAbpc734oSB8BDij8Sd8c1
D+UBm+W6W3xOP7n42V0tjjq9qEfz1jSMbHAQ+YvPsFqWIfP30VsflJ/uzNILJRpM
VGdmxK8YzNyu1kpDnJn3KkW8rUSs7GS9IDgmqh490H302ckgXhw9Ro6TgTINYZHF
al5QX/v22gmalnUOzTvvo0zDRjhZ/FPT/WlY9/1qdS3aTNl20EPRt5uZbpSOqywn
mqnqOL84asUziWpC9dvCkwE+Lk64Ra7+bPdNVlSL6usDxEaeoHCNmokYAbTSBOPZ
G9ctmopXE9MZrUoto8ooKA2QihNHTm6LQTvIT2NfhVgqVpoWE/yoa35YxPWQBPJp
nZE5QYx7YorXIEMvz1S0qzfle1UoiyDCGn4UcSTXUFcsseOWaIMv0xjqKiz3WgMc
Q2ds01Iq2zzE5sYRn9jepcdpaHFZdd536c716HUoGxJJzdBSO4+Ccb3bflz2zRXf
dZ43cf1bmWoRfddMhpYURtNCexCo/ZNS54/MzSJZdITZLU6A4397z4lgXX21kVSr
8R3iwq4CPAF4M6k/CG9vbCn1EPdK/PIeDdpu6FkO+egVuH7FrnX/D05tP+APsCXv
8rhpzFSHIVGGmmvOlNBBFE+C9wwZbaQIxa4t6sml4V+eQ+0VUCHFgps60cF1DFdR
Q2mPRjMmGhJ2BWad9n/IxvXDydUHbswSQPxQuN/3EnoteTWQiP7uoZRWKxzO0DH1
3N89F2Gh4XeXc4X/qBhz+eCROmpVT3kbuBU6cQL/aUrlLAdykXiC5QaIhroqcG0Y
W/UyY9XKvonYWRjc4HQQVinJObzhkX6GhCG1JXZUmKEe6EspNxwQ40bl3nheevFv
Q5Tyspag3cEAyj1P17RuSbj4Oo9/UPUcDcMY2JSWTO3ad8uYuDrf77P8nMGv0e3y
jUVMA4Su31RiLEWSrpZ31MYUqQaI6/YW51Ohyw54ufpkWTLmJ+XEgbho3IEJCVV/
HyfyQevx3b/nhfXUIufi80ewDhQmUMjePmuJePf1DN21nCobJ875HtiD8nxQdJUf
+D1Pkz8q1BaVEKyGkROnQbzFVrOT3l5VeWWpzUswgM0V3GgfJGPrCqezlQ9wozOJ
bPOPskHlNsuSIOo/SWRoPxFzpxZc1r06qebZyXCxuWCuD1Wd/xj0SYpbVptISFMr
HPD4vBNZsY1dtIn3e5KkcEO5iK21ZcGrZm7FoNjV6oy49sacGoP2UUOQ5NIxKWF/
0QDj30pLl+3685lNQApKf6uHfntAA6+5uanc4PlxlSHaq/0brdXMmp2ZJV5vUjmN
4oSiDnnaZC8VGk/5EXWxWLwKiYzbIMz6IxgtZ4CqpJaKaaNt+CWbDF7xkKkjNspu
eyqGvY5eAqA9WpvkOlNU0Ouaj4DqzSHP5/uEMa3x7inxF2rT463Pyi7mYr7tmxCP
I+NUlO3QBn4tyDMxk4V1CwMTNTJ61I96tcfNl9IBRWmxCLSCpox2Zpq3LVT/QHnM
OvblIIQxzcimFF6zDTW4X7rfLW8MSGsDUIaKThxeRBNGhT/pa3/eLpKD/35WUjiu
9UsvTDTkW603pL8Optwu0YBILGso9jWl7PBU26kgy3Hc13NR4XV1i4MSL5gSRmMu
ztq4zn64LfQcsWwx7fiA+6vSjZ9iR6r9b8Ka/wE1JOl5Wvb+DoSwYUdmmUlRndC7
oGYJ6FTRPt7qug5aCzlJLGqThIhV+lAQmaBkFzDCrNYcsO8EkSdUE4xL5ziRCjW8
NXQzi/47IHcW+5S0D/PhKjZezHo252vdN9oKUJJTI2l06HYijceMi618v2TCH5KG
W5TLkHwYebY+dGu1e/GhNnH2tW8XDCFZj1k/zcvcgee9wyw0bJ50TuHURxqPRvTw
UUAHHn42ftnbQ5WuI1p/2Tq7Hm/4LQRtIASBQ8Ny2cKjOIv6iFboN1HT6BiuT+xq
1TBH6eRgpwOR+UyRUUy2VkPG3uxxDN47bHFuqcj2ZWvYON0RS1lP+nh+jf37Pck5
Y+12avXRpnGxdg/ZGLxMltIhTHOu6XU6VKXH3vsrd3HnC6B/wXIrAyOphAFRtAum
QDIwx534ECzkEJHWzhq8GBvjRlNbFOX1EongxPEGT95n5sCnchZCxyw2HbnspBZs
0v6LkqsFCt+zr2gf1bTmXMknhyKs7qeZ2tfifEVfp2J6QevP/FythJr6PfyH6X+J
o1pHtkyLugBWpghx6vn9pBWM06syJm+0azJfM3mmdlcu4YER2cbd3T7xga8pPeGn
bnLAt0klM2WM9Lsg9UImgBZxnuZcawDr8JMzJZo+wQ/jR7LCyW+TKvj5pVdLUShA
h2xJ8OIzcRHhiq5zsPCBClsXoEfjPeDdPDttBjTaT/GuPQP+dhhnjsnyug3IXZTT
lkBo0lST+9q7/FNdai73Q3d3su8br/mhXaBko8CPk4M83gu9PG2EnM32+p/jIAOO
mTMrtDQmu8eoKyblHMtHpyVzmdzwJ9R5jGF5FCwpqUz4wFuuDfbi5zzRw+RN+pJg
/2qSA7eheLGrLitJzrfj5PS/CTC+NwKD07C5c7PvtPVOIB8/lD9HwxxfWEG4WMQZ
yCCRpzZDpRBLNo/rADNjK/p/xhvpQJBhqBLEyO9s8pKwbjOqCj8dUJaYthTHu+iu
nTuH6304Bslm83jJfOMtkhtBzdxe3dMD03faaPP0TdUYSwRagwldpe3LL69GPDM1
Irjg2rtf/To7Tx7fztKHTfFijERgGvchedaayZOxWTmm4HaQhTB9FfVaUUkf7X59
AY2Hw7QmLd0x0OQsCdg8gw0WMOjnLkPL2T2iLaW9OtNIgnMbsZH2zQOnYJmCKEw5
S/pVAZ7kbBKIZlO7C5MEHHOL1N8LeiAlmeBncnaxIu5CZNzldF1DP9UwvTmTOgIu
DlP3nG8V0yyPliyGHkRCIC4FuGd2SWcEiYpQC8xZTKCWXhXiODvvxFYDS6wwvtxi
b7bU9OhgFQ+PatelGSP1fYCWbc6sHHaku23BexgD/in6XuSN2YxzLIE8oh3w1uOs
FGbiQO+9m1yY8CyZWWZqtFBTBtYsdA02ZKsRfoLXAvTybrkKhSNUKHf2fZO6J4gW
xx5IDL9IDzR3zhUCHhZYhHyoFdAjrfuhFzVB6Sob68BbMFg6dMeMm4gaes6KnGXY
AjLobHPVD3khGXcbEV6WesSLKaxvqyKdqW7RLeMrNrCocSp64Cnzi72D/UlzucHy
pYeFh9pD4+soSKoOd6BmbA45Xpsh2jgynbDoAXULUDtsudcaVEpNVaQ794hvirJb
PsMWGhl+7wwZ6qIpqXxs/ZyYJpOWUaY2xp/tRgq36zDmes9a2soIiRWqpNVRH0pt
o3djPuW4RiWJquj1A2vNqb7W3R9F5todTIEySIYmMPkMdWScnFuLTh2dEVobnhH6
Q128WIw05UNlenbDXPb2CU9CT0lEO+VP08dhx4FRikMMpZbLGUAmvoHNG1eRVyuQ
IlcMTTG+oDBU64rZ6RQ2GHN6NJO/IhxauRlt1rIFGt5fUMEBY4yxGbN/tNLe9G4B
zjodwkFHjf829UFAujzZsiTQilFV9bbzOMSo0xSW1UUnxawv1l8m9R733u3sOv1H
81nKmcmDcM9xdrioN65UYXeHPt3kB6IaR17ZBFjKv3jt0JZRO1VTdJ2Q+l4xGb52
3/YEurvTWegOGEhZ7Gj7CphTX+X9PYMwKkoeyOLG8lK6+QOSmOpEwJj5GpjAeviL
Y11Q+9GA9d5ar7hZsxiW6tedOc/3K/1xmwy9T58X1aHmV8Cu6jaDDkwaYKO1aOe0
6LvSs4y3tuQicd7n+/WzEk8L9Sdyk9uGg4esYc9s21UvXWDwwUncl9EDRrrx/hkL
ExCkCo6363eHiRbsMg/ZKkYfqK0dg1JVMnLpdmNh6xlfH9ltb7lpTADsHxuyh40m
7IQnQqKBeTgHipiX9U5r5snONY9jNRAhZYmJjby1c3426mQr6L2lnhdS2iitP/gA
cis5KGZUHHgXfQiNuYH/q4EXOgHM72akgokklk86fziWP+WwAF0Wwi5lx7cEo9sp
dCCVGU/xDsCGswyCuOQlKfzMvbTzbhi1lBoyxOpFWurQjhacQ+uYu/BUZacSxEVD
IGgzv6ZjUNPmNVJvXdG7LeprJKE4cJaDrPeikbME1X0PclK1l+S94ZUqMuAZ4jK9
QEaPgAKEQ3kOO3IoQdp2VnskCbogm1XKTdW4V1cUk42HMkjOoOS/savgTU+JUUI/
SC6pQWTZ9tmu4zN8wqb1iRnvOrflZKB6csHKjPyzp5BBdDlPVWMTrp0moBerrXVE
8IfeRRDZHJbRt6qf6WwSykJJwd1PBil9V5xCYrA6cAyNkFF+gV7hNpnmczhl2IDd
RjygMKgSluX7FpYLswwWlE+f41uDnjal4tn2+nIcEepOyfBTc+i3+EI8a2bMsr5E
NsLlCY/OdnaLGX3RB18LFxU2Y0WSZ5W+3FqGf66m0liR2ID5R3SHmU8uwPfT2/Gr
Y/stBaTToqwuxGpR+bccgmND0H93lCo3CFEL/Ew6TtXxtpab/upr9jIFmwh+smzJ
WNerWKTBTAzUCYQPuc85/YQZo1fIqw6IhlFgT+stCdVUXeG8R6QT2uvti7A2QVGP
wVD9mBQB2h64bF70btLk9P5XtrfLax0AguNAlV6/cJSit6QD9Eg6TC0TyKu1dUwj
0+GfqOZ2qNpI0Ft3iugNaaSjkP32Ti0SxKQHWNMUcqTjKxTZ7lBW1RcWIMbQo7/6
k1dLs/2Rbs+ESyTsZajkvNhu11ZYjH4FAGOzGpyHtnHf1byCg/MQMGtLo/JK+w7M
sQs/XpQ+dcFELyV8pyZiYR1tH1cenQsPSGhGFe5m3U6V59QPdW433BH6+ggDYFRZ
+7E2LrsrMthui/DsHa99jq9BcLPes+E5x1UPkA88/+TnNLvfpRXEEdL1yF+r5abF
7nM7I9U/eTkeD0Xi7CCE+sjCRzl9jl74z/TG7inWTENLLcVCC4yJ1k4jNYMBCrfH
pPRLO6fNeMFaPAcyDXFUvnSCGcelhJDTGBWQzxUH0sGWOMqCGAeImkmi8aHUETCw
sZrmUn3zyt4ZDHJQB3zxc9dpREQ1geFdzc9Czzu5jTpcs/T9UYh1j87ReOivT6UO
Pes5PwWvfvklSgzE3BwzEv7iJT/1+sOjpdPpqSsnPe+uhelns+H7yXkGohBcDtym
iX/ayet6nfffHwGbggtvSgEHQ2FNRnBPLdtimcWbzVpI/YHrLatXMa3qgYJPFKBp
pGoinlbLGvZVR58zaguiANghPAPzJPQZNLoE2DjLKvucljg3tIeSNAjendaxutpZ
mMgkqdKQibXXV2b05DvDPihOMKAeWQ38HRXvOtd4RT39/DzDmMQI3b1G1Zgdc2E/
C+FXqqR0c9aYFm+6ZxNitJlpjn8et+U8BHjmjmG80bQAoRzTi+tWIY7dXdf/WYwU
O9S9Ljrc1XlKTmIcXSTXRL5vVpcL5caNW/Bh/yKUKYlvyyNoKFkcF1GkmmLLnF4u
CsK4k61OOtFV+0179vJBPA2P1D9TPT/QHNM0ao4cqwNMZXGfgqaaSkEqTvcLYMIJ
F00EW/mFqHyI4UcCE/jxOJTxmKuefAMtZEP6N6fdO4f9cEIiqqldmh2n9j8deQ7r
5S4+2vsuAS7vXc/hG1ETHHYDHYK3CVsBuglLJvu/avlQAoHwVcDjZBwFVNFmkA0p
dodgrLKBitOwfFkgZR0LldFubH2VCJVfSUK7bSWwOh2nuN3tt3GUjIJKxS8+Mv7k
iEsU0FLRmvhnMMtlO/fjcE99ZCSBiafI5ZSIDvRJb+Y0jMzqBYp3s8Tn/OnWkx9H
PqtrZisXo+gmIQHRJ74tXbCkAB7bLKxqBotNc+yCZY88HKJA+uuScRxdohJwSlCO
0Et1PRGVOLMW6bWVk1xu3ab5x7LGByY+ukQaPq0ALB4epOSObVUahbsX5oMtcHx7
sIlSZpY1QnsPxmCYkNk08v5TMh6CvNqHXTLzv4bHcNGnIBZ7WKJ5Dwe7dajOH8fh
iCvhvlK3CT5U5K0agRKTdtsvFWfra4IKALC4sKXMnADP1Ay3KIJErB2w+NjBkcEo
ChyruWfcfLKEtz6KoggZ3uwKQqVRPuwrqKLrmpR7kQn1rzCIj7lmIoeLaldSfLK2
HZhRVexMJ1zbeG9xyAzRDiMMlKH5fqiBhDHoLvdVlBmVbK/pg3zG4OiERCT2Sn2q
j9Sz8T1LvNEPazX43UEQj3X5KEy2C0mZk80sNgAn3jX3x84RK3CMmH1xcq8hN0iG
Z+HY1dB8BbTJYlbvwidvLsf/mxdjFa2kyD2TncFXgFQyihrRJHAQRw96AStLXpLL
2TJKigamswmf1UfLITKPf1ANj7lzS3j6BpX5xTj/fDfLhmqO6Hi2fBzWvqU3dt8Y
ScORjuUhTFwZHf5N4jHjsehnqqfzXW2HobyApyVrjTLY5zCegci/+gjqrcewIbB0
NcZqMPmrhOT3fYhb9Q+ja07PkSvzL6bWa4sjaKDjYUNK9x4WgiHSZMd3Et3Uqm5P
liidCnhp0ZcIHnJ1cRDognlouXeMNF73yVLeo2cmDFhJZPH55lhh431eNd0rSvWQ
vGcxGK984U3YOrlgELaD2hx+moJPLTFjAkJTQEnQemXMbbSaLEHYucxsQhfSZXmu
gg496Unbp1wyQjYucW4PfxY9uIkgXkJg7pTW7GNKq2bUo90AfwSkRxs1HS1hFpod
JSkrtOehxxatT+92Tc/OQOOUxPp2SKIU8ARPPGDutcmNHa0UlMjv8pUjng8SIcx/
QWWBzDdKAcG7jMm+6An+lhjzLGaaPAmT32c6qpeoXPAA7VAZNn8mnuVdDptLsy7+
ClKV7AsuABOHjdtheKjpfIg3y0phyvA/j3EJS1adweGmZ/QmH+v7iWFcP4wNmY9f
9V0WofIeF8etESGxGhMw51fOME818HVZgHGMsiTVwypZ/Tjk10HPEGUWRtRI0i4a
7oO0Z69/Kd+ExS6pMIzQUo6HTELjP8qMa3fpg5PGdyPL/VanK4E8zRvUGMXr057T
OSHGQ0I4/UUGgJSDYs5LmeJjQtfQq70FWuavBBkpQU7yrScZqOtx7RpBCdeFXJ3z
FvaNmu9eoHtQE7PJYWp4J1m17aH0cnyJQiNXY/PquFbFodspEZJYIW0XFBiKTPz2
NpeI7cA9lDTAKN7DIaV2OuiIO505GTOLAVXdJdCl0LrPqQwqwTZMNvQ0S6C3388s
4SzEjEUXsx8dhRvKhmYBXsJ9BMC4a1/AdMI7GystjT3HN6H/YyV7YDyVBay4EnQE
/YBEHO2Y9zyvwk12ZlyPbfKELOKCru9t+51ncS3lysx77/ijJ42azx/5Lg7yEh9V
JI3rs0V1wcCMnHMpZ/Sxb9UhlOVvYaU396GjVPpxHtxHqk/XQeCwc/3juU2jvrN+
4gZ6mrxe5P8UzXOk6obrIXAKEusVRg5Krczl49/SVvoikGhUOt9qpuGoT6WKsU6E
K8pkOT/49FT3yxMcUHraMuCi1MrcqtxRzWfBUM4eVRmGyWRZjPE8NpV2Ybcrk0SW
4Vz/IqnP7Gpcc2IAk8T52j3F0Hgel8ocW8ZEjuNJL39MdQ7EauXN/IpQymK1pjfx
NbCEHUiFDXSWJ3+GEfV33VjJqNy3643MeggVqlULpf7hwgLIROdYFS8VaVOShM7W
uQseBY6c3+ZO5uB0SKUzbs9b/b1hQ3BYgJ2OvrT3Ndq+dZ2uWQMGbuTmUMrWOH6G
4LY/sL3iHqN+/rPdGyQPSM4oUOYv1EtOCAwFyFI2t5X0gPtcR1RuY40sx1bbZgUk
ZLftcj8nOFd1UmCXcyssXrnppRXh3h71PSJQKkLJf7qlsmbj207xCNPlSq07Nwbe
A07BPXXkQPTY2f8yvD8CawN82FC1JGTMpK3ioA0KXG6xZd22/ep+ivn8LN6OYW0S
MxVQQJL0uZ22iIIpOJejmThWSFCT9kXH9XmXtvJGshJKix7K1wz2BWUAtQxyxt/3
24YacQ+tt/UNGo6cTe8lfy+GMvQi5rdzCy4yAKMJ2Iq3rqSEjR6mYmzvcPp66poI
yWpF0REd1FLXnJlOU/s/nJ4Co8QWeFc4cTRNw0A5/6eKf69NQv4/tP0ChtBRN9zZ
dSFC7Mna6wDp0LyS+Cp/R2+KuZKGg/idvySdKaaUWUNH29Gd/gcXK/FvH5ZHMRoZ
KLAH+wYry/dk+4A65kb4D1VhaMxvxLE7qJquvxSO0BHTzUQPTvQwXNbj5WDCa4xr
555IrP4iObOwtLK0KTVlY2YArYyVvO1EEylGcl550kwgR0OSWYJdnWsJHVLI2K/h
XxucqXHAq6A8fqKBixYBg42nKZGrsEl6jbQrz9+iPuNZWgpYz7MptZANFya2xNOY
0Rft2EUDdA1jQKN6u04x2Sicn1BCERrfrAG+0c2KsS3eO7trW+yqnZUhd8ZZ6c+G
w25gmBc8tssRYZqwzlSE07pE2v4xexSecdGsTsJg+y0qKkgB2zglIwcAYh3mYPIW
LRhCilBfbU80SDBreXxiMYNr96LyCvH9EpQoEMQu5nmgo4TyQBUzO9sY6O6P7Egi
BzYWDVYe2a5MXDRJU+fvscbVMhBbrkY58YFNqJWNpNLnELxYIOiL37DWfzDR1csO
oWOQE4nVyNwuSuVr+/xH379CJBZ55u9eSG0qw6W/DISAWU/36XXMTDU1DNvP5l/s
qw1GJ2pjblET7R8N9RNsRrSwcXE6drtY7F6nhrY7fXJeZ/E9fmrHzaASYmC+WgQd
+1lG4enZVPeMzvvMPESncqgSG93aZbuhnnPbz6wrZ2+3XshPXyhWta4rf3+1X6L+
heOfE+52Tn9LuJLr2b/mLZB9HBnZZPsZt+RzgnRuQqGdRlC8CCaQPCPFaBEDTuM1
F5ONwAcTZ9n0zQ14gAEVNRnhPTfyuSnWU0M5wWcMLsJ4J5C7LGyAvXPRBJTYeagZ
5H7aFIdqxi5EU5n/GvTAr3raZ6Fe9YsQEKn9O3rxwHkQXSFxgzp8mC7TAyDQJI6f
ryerWqL6SPwHCdgwiQIATfokI4pRwtV48HynKKpJQ+k+xh/WMKn88dAT3LI3HPXB
ZwEyKvsLojbkhe8p7rKIpqFcKljWtWyUUT1siN7hdM4+Zvzsm7i7rUJ/G4BQafDr
T2exVtmBQVqFLlgDoryc0SkI4aidPTrN/ubATuw/RP4ukFkwSik6Fqcihdyoedwp
gLGsXiSXdi/JRHHfdEP33bawebhHGZLn9UQhlNzHRjBMShniqwrVm83NdDRAnmc5
S+PzE9G1CWTMCV6gHoeaTBqnJZyXyG5LiuI8N1TmO0hUrxWAMazBjJpDXG+pKCSE
msTdyaOT43k86kYh7j/omgyk92HKldTw7QSMS9d301gyxTiN2znOzIj1QF4l+DZi
nJI2peTYmmxKCg7lfj4Mh+BPA7a7XHAPvLZgeCSw5I2eLJLSZhAPT91J1fsb2y4u
hkviwygFDNW4tG0OvbkxHGB2TBEvXAh16uhZ6o1hZEHL4uZ0HvVIFApyUDGcNfqL
ZuhRif810e9iTLh6p+6NCUl4lErDnztEdchFvImNjRh1M2qWhkbDsWhzZVkupuSu
C/4v3H7NbyUz75oFmklxkYFEpjpAQXqcpuXPiPYlNU3vR5SadMq47zB1CgWmdBvn
oa1yQg6Eufy0pTLLZzo51wUchsycOUMl2rCt4lgTc2kzGcRWGeCck7itH7+XCA3V
C0wsSjqVkSmlaYzVLZHO9w9EkFjOxQ87pMjoQsCNK7okfSFU0SGXIuWr3+kCdsa9
K/8TI+R9huwBCEz9t37pvMbJxHjf2LQFfNgd5x+hpT/lbsBJsP9hOT/KjQFk72IY
i2KzI+8QcQ3Voz6jAfktzF9wxm49n/5MyHgOsRpEUudpqHpETxDYXvcRCUSp0ze4
QKETtKvyZpQ/ibvQyUziA4RiwjEwOxX4aLUgF+8Gwuxs+8MopbR1Ba7kyPd0EqM7
/aNdn/ZlTN2kzzsu5G9wz/ZvtovLQakeWhX7O7YAGiyb3Dt83RH40eNMNflbxWPM
lIlycUuOJJ8Q2lkGci7TVCdYCaZr9bcg4RWBtRO4ZVlCy5EI6HZJHEPQu3OkVH3Z
f/eheVcKkU+bYTfBa3NMW2fmj/3pYd+tXcMl7ecIcmhvohoNb0H7ZPdg9/il+ukA
C6/Iu+fHFXVSo1NBNmYT25sZuz7M0zErLfqsavEzdO02VxUO8WDOeGPkEedZfCuy
i4kgXxFYl9fs6cUrHAqullsfWil5tIsBncuwiXqbBUYdxzS8NvLEke30r6V1KRmA
m2X/s2HI7LFdyUsXFXQgoZPFIXmJzzLJ2gk9VkLWrU1bxftfk49cPxxRy/hiEEs+
7L5Rj/n8RkzEVPAHcQsYjEm815TDfXC00PkBtvsHhdldAiEwGq6VP7qM11CdejUq
9U2MC4blP4wHzEqX/JMUQiUQlfs/F18afSvT7FOSXjPm2ItauC0GsSGaX4tVdTb6
Vf9bNEq3UkGoXDD7nRCZaAk01fUPhXWoR/qPglNZOgxO3CsFXkOSnGcROD56dvFd
amwS6YyCnnpFnveIEFsD6ZM1I1Ftcc5y3rcaENlUawAR6Y6iqUj79NM0o/ahQDBU
Ii5FRihbCK0vNWycNWX71dsrwlOt9AXFTyYN6Wd1lKXZpcGq0UJl8suhCeMh3tL5
z/lC9RaP3fRSkl5GPn9fYiw8HO4TuxtBobOPBVbvwMPXij8REOdgwkJ+sZbxoZkY
nuWpToUlz2o6NLK8epfuce4FccAnwgiBkbm4cuYsgWE6XMGFyc+Zf9At4k85D6HP
mA58LG7oCFuCT6staXOkJBDem0So2iYxMd8jA4nW4qfY8pOJ0xBQdpBR5jBI9S47
xRwchukyvomNFiw5LiFpyEHsah3BZbdg6weC7GAGWfNAlB883tpMdDxppamxIb7J
ZtM+rY/eUDPoCWTaG+twIX9597Iq0xooKiicYt6ct+oCGlFQ6DIDGTRKQ2IgrDuD
tHEnrVOVKsnKaBRjKY3C7c2llAWn1riyi4nST3+PboeErJor95Cpi+faDYn/tGp4
xGE9hulqDekKRgU+99zzh8lF7eDNhhpn9wtp1s/u4Dw3LP6nrtWoxyxT8TNb/inQ
mDWPJ10wKsUczBU8ArdYSx6l3G+hfPrbdMGTM2SvIw9Hj3DzUZDY0DAMyRdE4ZTD
hfrLKPKxqppNRcvpI8+EFYdsfhTdGAmFErH12q79St80iGJM/38oQJmft71Zx6Aa
IbyKo35dxkt/vHbpXkKFZVI1hmHcuKOMpoXWjFtY+uW8LhMtF592EKJZwNEaRFT9
jtiKG5bI1vFwt+qZBmUM77SIpUjIJYscXxd6vNUCegIY+TGmuLFf0AWjC69BN9E8
vLp0Lc1AIiDRJE6GpcI7MeX+SsbcjG8Dim4HouxU7IQZ5sw5LZk8mLumALABSA8l
69FMcyTKPzYwUfx7Gd7xsGm/P4aAx0DebOr04AzOwyyESjtqJ/xyWdhN9rgy73ru
fvHBUdotWCXeClYrcheeng4pKZ0pOyRYftnXhFmGLc5aTnTcx0/iBGlIJXH56vNW
n4kTD64srUhVJQ96TKFqvpUR/cH03Wyl9fXcAb+D8NCpOU9FjfQ4Ikk31clymHHP
trA2moxxf825yoz+w1lryrAU/NLl6X/VJfYPVOo22+D4K5ahEFGDVAn/op/1BPGy
QCsfAD3WV6ALPz94oE16n8rNczO6rm/sawQvEqOyuAyyBu7GEZu3gYq3c5hbSe4x
pqPjQcTMQTRZzFmgtR9E7RWq6Pv1g6ap1nBTsYB616h+pmsRl+c+UxrjDB+ps8WU
2tPAZB1USAdFL0154cm+HbUX7LGbG6/XPyBHYzt5rMCO7DhYNVX8x6xpFc1czcak
hL8Nkd2xdAkGV2TxkrVfA3nipI63BfYWvdxd9Fomz25BndEST1XfMuqzYFVZ40WJ
j0TlkE9X74gJwzpLNYn1lJzK4JW1qVm0Op85NT5ACu3wCAub8tL5sBTmakO8ZklQ
J3/ubqeGXP+z9StyZpk6R1yBfyUwZnZBYsI7bjvSW9858KaOmANw1VB8FuvjpE6K
PQqylbu2DNT893X5foVW4oagrLEh36O7L2j220GTfzjS377lPDj9amUlMcxAQvlU
VQC06EgochxjxX0tpo8fAu5aOIXzZv18pYHztSMcilZ3Y7f/26ERqyFr6cyMB7r5
VxjcGVtqbUW40vXbl5v+1hdaKoJuOS1E1Tz6xQNc9PUlQpFj9sIlaokKdJN5MCR0
ft43KHLeZGgGvCcFrq5AbjBNT3wl3RKf8nJo07SGzIo1dAn2DCRQkWMCGE57YOQ7
EwsLn7i9L7Ka2hvLz1BUnpaVd9u0ma6P9vcitJdSE1ojsz0V6Z3NU6DGCNWPVH39
XJyBRt7YhfkOvuT/BfGjgsPGUu1MncaE3SCqyjYb2ZtvpF2B5yS2QkeEclz8Ornq
sr5ndaNDr6s5svtVXgR4xNwtjoDrHl5D7Ijy4NiU78EqI+vLV2HnzRDWfT9w66Xu
MmRGgzfHo/rJMJ2X95DQusny3QjuEQ/l6FFjKFehTZr2jDIEoOu2izhfnzmtGSMu
eDU6tIKCnkdFUdIgtk+ALFZ5SgYyThLgJqEGzaElpQP9em35LPDdg7SejPFc2d3e
NYjK1ROWmZLsqD45cFyiidRCh3p36BpDMDIvIKBxOLBopJDk0kSRbztrCfv+C1u6
94nZUM6Z/1Eab4hnMpmK+TDq7bMKJpIVuQEcc96fP/FtO9Vpk9sU+27LP9MA0tIt
N9Cs6UpjoHWHbdzCwnxyjlW0diwLhc2bsHUoW2EmzKGkpBBZzKvQSTdTnj24iUmQ
eBcxyP+fkhy4FW4lyVKnli98HQlk3FB7qdq39uo/u7u44ZIjeOnyaFpHJYrWlTVN
wOiUkTHOE3mxlZjCZG6skKWf04Ze9GNErEfkbSdRGnIflKkNJDAnk9xyTWF+KnYH
XZrLshXiqCGqBc0sNEQY2RBabrnpQbAvfLyOfFSzsI/s+GTvPhzksxenqT/rqgR6
fsbsijibeNcLjXojSNLtaYA+5xoVrKkMgnpv3FmUK/uYfE0hAmH3wLFyMbAhJsJA
eDDYvOwtxjSvEB0KSxtjRUx4jcFM0Z3uiCIHWPme2iR7lkHJqoEgsT0JzYxXp889
3ArdCLt3WR330G7OqWr4OI+X3QYKCqT1c5yMWjw4he/8rKptcBbimk4otGTPQEGB
KRGvYxSr4IAd5/PFNJb2TmDma5c18Dj9ho3mVz+rblphXcuxnEMQUilxlhWLR3MG
SphW7qAcoVpY6dm0Fr/DjNB4etkWA5jJbKxfDqNKy6VmmjAjLvXEuNt74PH3uLy7
JHZbqKlxDX5pSRYtYkECT5v+1habKLLM4fQ8gsl5RK84jBHrLYSRWj2bFocQv+oA
HjIJnY4mV3a7O1Zvfr0bYBGngIcKWpOvVPNVkWOg/PNo2g3Ja0lpukLwPrCK/uaI
kOmNYYfW9XMYZRQi+xR0jpaRgi6N1YKWWCO1gwINyDrip0O3QZn9xVbgfNJbHHnO
ym8GThJvH3wVIDeHTD8GTk28NODvqqSEszHBbgxDCDvVsvXW12srXc82+4pH3LIu
2CuEKsATLr0OiT7tO1btV+8udXKb4/C3W8vIG6wTm5ohsGxjOkW99xe5eSp6EViQ
eqNMDH99KNZnroDSgpc3ET7XCL2lpFYqpI6qskJN+xtY77OPyv8MOU8MPnlk1eO0
CmuDni+wAGZ1nCsUavVUpj/bQjo7L4weWlFaP9rJH8H7KxMHmQ+QgU6TtsdzY5NL
ZEkew0tZYWHMUmHQILp3OsafSlF9o7SNkj5sUN3YkZZKFyZpmzWSPm9dec+i/Jx5
zce86Z8rsNa0MyMzqhiqvZC/vdUuIAcZ05OzZSoYOXi6FPRNCeMlV5igRGBnFYOB
usY4Wk/sXhkv/ZgIS6Oj7fl3XAQlIJPR28xz/QK/oLZIQ52lP7vtDqcTFX8XTLu2
lXa37bnfJnY5JZuo5gbT5hG/nCnP2WSEvmCpcMelwsV9IuDFSPVbPGxadc1uChKJ
gULzAVn4CcGgsba4knjQkThL3n5SyldMS12pjNZLCrvgHv81uTZDlY2FaqPQKWof
az5NqOR93f/+ioyVwZKRahko0leL8V0PHoJkMfHn0xl5Pfqapzz5ccL978JDeYhm
ks49pKyp+s5VOqyZboWzNYY4ZBsjc32+TptREkNoI4Zi+xw+BbPIFEILfGuDrzKz
HQ8qlSExx9Uaw0j+U0PbXOEajTamcEvCTPYBcKHpGO/i/rcEqkmCh3Nn+jV499Q6
LL/ayg0L1oeq1jXJwbNXXW5PkpxaZ/HPrYAkBz63V9vTCOcJVKReVqC6gq/4mZqw
+/FWDI7RDncCTp+XJJjMp6BsWB4pUaOgCkgs5akJBr5N7LBJKGnAHkN897g8naHy
f/tEEKs2590LtFJ6VXSRUbC/wgtokFP8xM++P99KqYi4Ady4pOQ9qMIzxaEIjDxv
dtqEnhBINqhF9nxWOwf8jXLR3OlT3GoeUJG5hYJmxa+YJoxVpH8oH9z3AXNemlga
oIcCEuP+bEZY5QCfjptIyvJCkcEHjaS5YH0jKgjsk4QKYB9RixX2NxeJFl7J+2sA
MZikTgqmgJv8zA7k8ijahmeOPN1MSubjpl7GTGlbEonFs9cS0DHFXFtkfWBNjSi5
CCfMPDvnOei33TIa0kSYfYDxngGmJFig5FNqCpELcS+TAto42d94JpWyc9qgkcQD
J2Q69uo5JVOQU5vSc+RfyWVJxdBm1U22XVqyh1L0x9pPNu49xBOSuSNDxmwZFmBw
BuakRqYc4GsNKLP8pYpGeG2Eslop+VEfVntgy6wbSjXIj8SXPMUeoVLgILqZpr7Z
iTYnV3IX7jXn2r7nne3G70U+R1jgT667RmPR9pozBWH7HvX9O48MouYhppgo2OqT
eqBe9HH5UCMkUk4J0G4atCxBiaWsL5+Xr93HgGq9YRAs12gqBUUgseOQcZ/Tau/7
2oxodvj+LAc0FZKP3sR47MiYEA3HGe+4THMvfaPXmM4SdUPwzzYlkbBCEtNUVtpB
6pnxFOYOUAnKkN8L9ZKOOYTRJuTi4XKkBx+GB94oxLdiqDEcCYYuz/iPLacohMi8
24f6E+AGkRoExaLd0dWTMjvZuYtfPAjiCJm5tETf5a3OOGoCP0MUxNfc7mWVSDun
qc6liK2lgPkFDBOIo1kBWajd9wCuJo3x8D61tu/hUabAI4RnilDBX2yzvb0t9Ak1
uH9QkliEY7z77WN10kry3hbWCUZZrcpRAWlh9mk9+nvMjPcNcwPEHZceGAAZZYTQ
LXY/wyska8WZCMFAWGbEXxD0YnuVsQUQJBkZ8lP7VXpr49h6Ko7HML/ZUwPtVQuQ
p0qdSc6B+0S0ijAmIdwc99pzLTWzNjPuAfpPDaoYCEsxcbeiBrbS6Z8bzSR+PSf0
Fcq6O/orY1PfXafUY35uJsShDoDEna3FV9ayfGsMbpU3G0BZCtbL4FJHZr553gpP
LzG+h51OoET7gi1NZbzehzszpS2qh6CdxWMbQxogfU9r/7yPqWHotbBra4raDFvC
bFNetNR6Dgp/cLWh8+7zOY6dk5SrbrIT01WhUxDuzxe6lmZfbhgbfJSlJxBSnTBr
lnY9QskauP+daVbQxY5uDPkPpLwWN2B3Miio90UoHKbkFQ+oMAYRfkL/95YP2Z+k
KQCVsYsZF6g7McCix2aRpAQiw560URzKO6q4PKLaSAg0UJeQVvk4mFNx1lMY6+L/
byyx49tpVc/wct8lLEkfgsS9twEyN1J7IU0cNygnlI9Z120SiuCuyXcdKuYtYsBP
soL2EvdnOs6eBTMDydsnZI7JDAyvSxYmGDgvIt9d4cXcGnlI9x+xPmDG3Rl3hebE
snP6PVDZUlT0Fk7eA0mESOj55hOo8AE2IrPGiB+VWBmB6l0bKDkGpUl4KxgWtKLC
z8KFrmoqlK6rf2sgoDeykeQusJfnhF0+v+DJ1+JVhDzGcRcWVDFv7EKRk6uyj4ot
256aPvyW2yL+Vau1LM5BQSMnzLoDM0/ahA4I/cm7IMbkEJ14R+gk2DqjnMDJuu0t
5h7yGTYp/nSQQuyQSjBHkvZJb0sdRR2f3eG/5WAeWnYJAhYy1ZiG4ZLxnlCaEbNO
XhrlFxCGc3Aix47yCVuQfaRg3RTGczI5Pw54aHCCawxi4YAWJKnZp7Vg8opc8U2o
n3JmAQ9oSY2dqVE97rJld/qyNVZV2zdG8uGOr4PgHPqzCrF3y8TgCwN3ZTXOcBYg
l1EYuQU60uQFRL5jfV9L7cP0KuMaZiddhu44brX1cAaR8NZoKB02Tqpbg+oypMCf
58+sMtB9JoKYcHRg8sLKV6bu0LrK6HAJoHcFrmz/xvtI0JoUT66ry6TebAR1pgy7
1QuB5/ojHIm8p/hopqqnYaS622o8CvR2E8nru6er8xlbUHfATDgdhLhuqoS50FO0
YMG+PhX7X1LMSX9gdIOHjDBCVMAhKSsd86IAsB6mJK/iYur0y0/EZJZtTw6e5V7F
nTMX0VPqIe/GlTS5xogWBEVXE634K+CWGxywX2pxM1KQkj9Y38zyFGZJdqky8STe
uvJNYpE8rf91kqoPomsQwpYkgXlopOiChqhsmkk1U0plUZE82r4zkUlv3UuwpT0x
1MuhqFhq91ngvnqMLvCyV0AHxmbndcqgHolt1y+Akt/es/nkKqxX1BfFmwW0fIxa
vURVY2CDhiZ+Tpz20wmQD5heiTxy3z6t6UddEtpAky0udk1AVJ43nnHTPI8FhA/j
Y+gDwWEPqC+F39PIWFizbVvhc9JejQy1TlTNQV4nil3XtRqAIvABORi+LDf42fQI
9j0CXNdrcQJyvSDinUfPAmL5XVRTAtr3ZlJh/S908bTQmq5n3q3yEjZgm2S0Kpvy
8cATjQwcJd5U+JXdiugd0YKnQvB19gCrV1WvqTzJgjOd/7+zZqJJBj+EAGAPTnmS
UA5lcSplGmQDdpRPlh4F86G1ZdLHF9MlMfTnA7jOdajLVrbBqJjaNqWzQJhAKEW5
KqlSpw1JkdFrAtSe/PK9NZ8FCOUd1B4/UOBMzGFfnZ9iP0jmAfZH9E0w4o6pI7qM
7DtTNUeVaWB36BcqwaL1Ua61sKOa8gyPv59dxdzHeSXM/QAXhgExCb65uep4doEw
C1DwLDvuUPgZuAKBJ+2QGshsqWwaTh08qHhZbvUP4OdWLb7WedhWkkN67qWJ85B2
PshdaNoMLpD+XuDOIUmhy9g22B9Tl3XO9B2mNjzsxDXJPse8PZXFUUbjNwQbhfgY
sltI6wbelNVqCU2B1aXy0PTVTRwFRf5hD1VHanRufzPmjI8OGIaC0GFUJKtzyQ1U
ov2Hd4AQ9yf/sK9ZcedC2mREmnrnBvHjYxbmhQ8TG19YSfOWTluKrVgNO6SCE8Bt
0DmcAF108hvZpjZhgWa4X06p3iR3uTM1+hK7VMIvRCy54TdN7Fij2RG0VqeWAH/4
EPnPi3Fm2yqMDP0h2LZgaw34DiAyE529k4akRIzYpNqUwhmSDDHH89GjzBeHOtPC
LWrQ1C0NZz5saWXc1auZ6osFrfwCD/0zIur83GVqLbjYr4UuW6WCmnct6GblA+TJ
qao+9Aqnye62ge7eifvzVVddOMtVhbh4qBG6Jyl9BjgmCf5Aj8s6mgetjdCJhoaf
Ho9FGE5eNJSIjPwnK2kvVpm1lGYF800glaqkb3FYI3mPpcIEeBQ9BVgB49hMIvR0
p7irfFKB44DQoY3JPRDpLk7yufB8Jc6wij8b5RHAQf5lpPR5aCJwopb2kp3+2GrH
QMD4t4tDYUdcr+S2Ket+wzM2yyWOuOuoCI/iWDHkIVFJeWm684vDGd/ysq1nXACB
A8H2+HDmjSmgzHJGcHB7OQ7X+QSW2aT5QlkydPYdvL+3uF14x8PWxlnrbT1q8TQV
BiRKete7ts3Lb9aZwhWgEiPmo6WNPLtnkGyev3GtyhDj4BTJ6vtXz5+mOmvgrYII
wrh24gB3YbfsjIOBJqSys3wDJG4AtOthVpAzqXXUoXtkNPLdz7bAnqHzviNP7KSr
Ii7pVS9Wen++xYmZbeQgOI6oMdzrcUtku7fEq6TpyYciQcNYsSTPlrQEahW2QTxu
wRL7VEf6uY2MmdFGjeZW3yhw16PArqEzsqHg0fjTNs9DXdC4mQ5AamTcYQaNJWbX
eCMRlQ8HliWgSXi5kpdiFPE+GuIzMSRng1cVSih2It6jfCLVTzAd/U1bEzJBQDRs
HyYJQByNPm0Ztfq87Y4ahrEJZR08o2v4z/5oznAWCMdhpyF+qcrpc5NOqYyHL1zG
n6fjhRCzUQjINUzjkRxn0Akic5pqk4Qe2gc9zyiPuZFBI9PqfxsHphvK49rx/Cyu
hn1yTRrlphTVMbHZm27Amuf5kaJLuuj3WocQg9Qj3wxDIgVqmSGpCwrATbfIVcR/
Qg/udlLGAg7pVzm64xes2WXfcOn/nv8Xke4LpaHgg1ssCs6OrFLtM5peHzdMDkUz
6QoUp4HrD8YZbFH6TgykQqivhoUS4WIf74MtqUH6pANpdY36b7ONHs7XyEgxdTB7
xBJbqRu2lFCAjapuWwcAF7csRmTy7SeUgDtcCd1c22bOtBRZAk2YaUO82cn6+fxy
zqC80RujXkUmclMV2Rmk4WHh3BlAOJskGIePbJcCF7JNZPU4GMS2YxpYawBL36L+
nxeBdYZmFVEO6kfPcT9YocKYNYa+cYkGktFggWw080/692fNZAQsUiIF7YbdT+E0
jvmIQh8wGufgBMHDgBFk/fxZkc2IBrYqDhPsPQWeD0Y0ziuPUiAPhiZNUNOfhP+N
5N2nIWHBvv+spp/FLEsLkpEKL+a3qQJ3HZA/nDCvGGim/ra6iPS5ASb0+WEUEhJJ
D3nE11veoEwNkfiH4MbACt0ac25brUL+3Dm/X3Sbq0yiija9Qng5YUtO43YDe29Q
chDwM2pchJ8S0dA3G4+BkxQYuHSvMYOMznc4cmbIySDenP2lGdFCRFu3LM07Mvpp
Mb8N36e1dh+DY1Q6dH7iUAVWyuQgCEoj3SFNyENTLXn8d7I7mBaK7W1HJc83Te/r
Ju4X2FOVS27zcLre1WYl9D6rVVk0NRPnFHPJv+ldzlxrePSW/6wmC7elHQOO/G21
wjg/3k5KLqf9Rlh/EDS4yDNiRldIW2iCjVvotemFW3mK9ecdnuDQwAsEicbkiGvR
VPQsQKSu+5YGIRYzAG22MqSBRR4EjrKE59OcixKm6LX8YytXLDvEXJLhFhkjFftN
bRIOxsBWOg42j29mHkoYiZc8Kg60uO29nWBm+G8a+eJt/nrIN7MbYKna5M54hwCF
ijgLF6R8LqeZwq2yxyTY9kH6huJfcXqkBESk8yJD08HXZUPdp0jhUskQTliJobm3
wutuq5nQIsJl+p58ldq70BsCtT/IS3H7X1Nul2rBr0Jd3wIWtJKEdPhT298gGh7b
pfIl/ifRo8e0v0s9ty3ex4222NC/LO7sYyKK7mgS57JubaP2USrk0V7nliG0dNxN
5TXBPqhdyOC1SkQ/sKWs0Pk2AkyzFeFg3+W3njgFlRaD5JqVikduR6AuXAik97ox
73xA2MxTL0nmVJAVFxteOaKW14XdVucfv+b0x+bluzdwvbSJVEqeG1pcR3EqK/OJ
Ag2De+reUhqsJhc8HCfF0bIYsg1q152N+REW+ds29d2Qc/HerMkr3W4QIr1hYkXJ
O6tF10ESuwrvKX+v1JY/404Bq16j0E7LW9hqRTk3JirgRio7kw4PA3pDRPR8U1fq
PznHCf7VB1fu3QF7XjmREan7txcYkW4/b3YayQKxP0jeWDC9tROOLMPRe6jsP5Ui
DKjhDhBNfCuqKprZUbjFavViRbc1CbFwhGL06Zsv7khGf/K9S9da7L3GBbwlsmLV
N3+tkR8TZ6od7l/Vh5pUdoT7OdEH3ltH7ys+OqNY8zsYd79T7S+ucqZ2E67Ky7mx
MqZtyBd1cifty4DdNznVj28ENPNtt4ZoLj+Y/1ZJZg2ZTV774TCe+pXVOgKSJGLH
Ny8p3ZPBOufXoU6uQLZxNQRr5/ZzPo6RuQM1oXtrWMhYrJnEXmNqhxGpa+cW/pe+
UkF/SYzYFHC1cuFs3Tkm6vqklgixGSBKH+QZudNjNpdVNA5l6eDi2fijUbOOoWQi
ZgHA2MwV6lGLpuN6sDst1gquJwl7y57eUcAPe2BtR0hjTfx0bWy4IRrwfaXahGsh
aj7FhSOIiHC3dV0mkt5P1FMia9AgkoPAaejhPNBv9EJlwOVGl64R5zwoxdDHLDks
WB41uVYqNTZS0aCMBX/rYOVbxeMIUT2ui+ICxleVyjMQBrKovujauK99PKP9caG1
qNn038Pf6Xs5BmAzHYWnVmJ2CEpeQl98mGT217ajb/NJOsRN8EeNwAe/4HCmVseF
IjvJYgypxqxBkL1aIQSd6Q4eNOfjljeo6BNDTxJN4RQx2pt/Cx4znCnlLiovF57T
pr074qvGEmahcz9iQZCyVmJMVhUB9JHIYjbcRKi/M8biMkXkOoVgO/06s71F2bwC
SBlGt5HzbF5sgf0SJoshTCZZ2iocn6M8gfuJaF/K0hpiExfm7XcXDD+gWjIp4Kyx
7SqjyE9BUAQCQJTS7IpWblw57zUzgx74ix8ad5giUUjMO/SlbhVsPC1k/zsqtUwO
lkOlQU+1Nq9kncUTdMXHQTlIXah3jUW11NHYavUwkGuetz1mgr3eFYvioij44bwo
5vxMTKgLIz6OXVd/AIwgB4KE2A5pkGPOMzOYJrd6H2NW4E2VPw1SGrHr6S6UPDOm
uM+v4+8ewh63wlbn89fxAGXQMzkDgjeiVnpdOBbqn4hSOTkhZ9QsAW5ljfSSAyP6
AlbT41ycKN9Nr61g0D3DIeiG+DIxxcLNu6wxrvEe8bFksSLH2Z4TEmU6HfDY99cX
cN0wwi2XZVcJee2FF33OP25/KZFh1KWFPcquBOxhWgdK2anizXWi7+96915wj46d
vAroMMz6GQ3bbjIQtKdY2Ynn7sCU1SFHckENBBbGBU5CiAE4RTSEbI6p7jGzV4OS
oVfWYImjLO+g3DcfF4AMQiEL4N3irYO7hUrTEqju8iBwiFWvfwuRUBiXiqLDcD+A
hUG0yo2Py5CBgGkkyUkCuXSLFCuTlnlQjCGmf3D+9M9D+OS5qjRW51aszoSyZjAx
HLsLnNj9cy1jMOH92fHX03eoqVs5EMdzxOnut8jvoyfTZb/kTRVOVoztFQpRO9Bg
IwMHooIrP40QnGrzBUrC0ndiQCqkztpyapYn15g6gsNLkZ8Ihi8r8Y+IqaHZ7RDJ
bDBulbUzWLfdUzWh0e9BHvii83tqyKd6uRfX9yFuZNsMj5YDM8yK+2+yOoKWndue
8Ly7P16QN9g615y8Hcw1dLSYNchXWI4P7xOgm2hJbBAQp/VYq2NNw3e6BiJK10ww
zZmiPBSXL28kIVozPDKk0WgUg+Yb/Q0TYdVksoeSdT5HGLLY8c5ACmBvhE6gBvBH
GP/tUN9zHBfFBaHJUvjU9tCH7wrQtyfg5bksXuqcc4ogDO+z1knusY989IP2jEZa
mN+pK+AukndTNrqn9KcSz5ERIa/nVN39gzcR0luoXy1dd3J71WswgI0ORM3sG+DY
FY5pX3HL285d3qsWDn9CaMHDAEgfcJUB7Hg/FCNHLG23rwiKz795e3jhKz+8qZDb
nLxiLVLcgvCVvlMnmh96ciWYJcq5L+tLGyXlIsp6HXo3FyYDJDuu/sehuoakEcy4
Sr1hUqwQHgAj5/qHa0Wlz/+wLlMJwauDCnZVjjFyf0KO9mKxV0wf628MfchhJGuo
QI7y7UHvsbzjLgg9Mr4WxjKzMOH7WoJWIMEtHCDRiluCiii1bpRSfxkpcBG8kaaG
Rw0xAQ0cyqsmwfy1/nTHK87jt3hxQH4XTLs9phJ76VUwNNI/vq5FWA8xb2uspOKP
F5PhxJWFvTEamqSguzqVCZuWr6puV4mbjnyQ7rC1O6NVLFXlWv7Wjagd2WBZmhKf
eyPXC7FblGWJOgmIzKVscfG6zPIFDrC7bWAN73HRKTO9QqFEpjPK07Z1jNvbVKLz
3WR/peUuX1y43/ANxYPJPPSD12+0vwCqX8Y655sduh3YN3QhBxoZwmtmz79KdaYM
zAph9dBaUJntOzmeHqqZl8NQuGtPmStgcIdyJJettiJETeXtNo3sN3J1OKiepRjK
FgfrMeAWiWJQFkJIxzp5Vf8XZ8Xf+Gik3fDpP0rnFYqsnn/DPxogLGEh/1w7pXQD
yLAJMANmk79h1SFU6ugzNv8RwnjBnpHnR8ET+RhP2Tt+WVTxhsvdptAKFTulKp4l
kkRmEjWz6LNG5n7OtSYD3sHjaDo0m90eqVTJ3LaJ8yiwjYA752wMzo5araKpYzBp
FPl++NffRILGuJlAQOyyTCPBNltE+byJZ1Nyd2f8f/iioaeC+Kd0yRH38HbukhK9
JzfQofNcUHl/X1M9xmyHGYv4gHJbChR2PRGoCkJ8fCg/VK4yqr+DnMJlsE4a1cyW
Fhe1RtpB9hkkxzhqeNCUZUiWt6PrA7jgpw1YrM5yFO6pnwksuhAtrLLmQKXMBYOG
GqIiKN2eGfbjrdQilpLsWFhhTXNfJd4Xx11koODRJcrmt4ZyYcFVzyYNxf7MRtgW
JEQZRG1Imte9Gw3ln5toTgQ5b8EbtB3K/QeRLC0td6EY7HuZg+s32a1HZxWLK8q+
0/MPFXCTq1tG/fgwtCflZZP1QLxlLSMbrqTuho0ejFO1vJpg9tH6tZDCUHykmEls
n/BqQt2FDdLcAtSZviYOCuKvRE5+DUmclekYBQ53UY1zGaeSlYwZ1e67whujowlr
F6FVJSBHPY/GRZodOWJ0CFraYW4RcZS3KXzJEaePzcIa9e4qVIj+kZt2uVIJXXX0
ZBiyh8ZmhkGPh9oJWJPAupkFZHMqxy1gywJx0GOvMdsmAE8OnaUr6maTa7211qlm
GP7aJrICRzqZl7/qxnhFfk2WxigPOlU1Dvei047expKbbkfXgSvWasL8R43iXnuP
7KlrdsXmoKnecDy9tYLxsT5gVkZKyM2dMnlI68EWwuputqF+NGq+po70VW4/xUkS
746SkMAwLyLgwvwPWsD3e8H5mWi05msMlGIRbjbsBTQwjjiJ6xLcR/4IsRDXyWT3
nWPPMGMT9iS/oSQuVFUe0z2iwShekOWazo9NHhbaqm9rMz1WinAkcZ3rkKHD7B7m
Ks3AuILR/1LRrTTtCPZ67lbDv/Psbi0hWf+BuKpdlInndL5WixYxinBnmjzuATVl
0O8Te5q3v6WS2tac1jriU9ObkiQsmb9fLxCR5rN8xx9O/+z7+GZVgf/O+9mvbJiL
kvVoAB4di2V/XElImea/YogRVW13xPE1dvGDrYN7yQ0TCg8YP5bOD1tYr88kORIW
gYVeVfKGFISatc3kob/ptM+pXG8GzfKcr+4Q6KhUgBA/KHz6PaK/Mk1vGkcViQoU
5V+uoT5iXhmnyuTm8zC2bE349JSgBAj2onowK0GX/tcI61nNMmZtp8m4oa+t9duC
GiwTNtZFSLjud15aSHXvR0YRDfKRCrszriIWMjI47LAKMDjGffwhhWB3miF9qNpt
76nhlX/HWhB0bAK6TUiD07shLL8EnlKKc3lQcWRvd1Q4DooUi4wqmqgRDt90xrPn
55VazsiwDXkYhyq0ElvIg5SkdlGcvVWp32PMrxp8R8ew+wkDRTtF2pgPN36t/FyI
zIMDK3FYbd/QMCV7GWdRnDVRCwoW8xA15GdwD0YOXjFZq0th/x8JjcQttftxgBiH
UbwC9SJSzqnFYiXvAY/VdAoEF43aIm1w9/+FwEXFpJGQUjAqCbVCtxWVTqQuxBEC
mz5jViOtnXl+cyh5iQj5ekaleaI0tdovcZV85xQKjbY/Hx07k4YzwDdziMuAIDXP
tp0IcwW0SFkT+w4IMghkcoe3m6MURwQ66/XwWgZJ/HbeAAzzzWmR0RG0AgKzvA77
48yuExqz/mZ/1Go/sRBmJi87evq3gCz+OjowefPB9m5qbqbJDf9AK0tO5Jod43P3
DSGTOZaZwr/G9LzNkArkZz9Y0pM1DVMspdeNW73296+gIHIDZbKu/O0YkAf3mSrZ
MJtmQ97SZdhMDo3HhTB71gZysjWmZM2mYOLTB4y9yWqIiP/a5O06uV4XE/PwjFaC
fuUN/1JTWMn2i2eDj8GF5O4HmyA5q0AYGj5Tq3Q/vTNEEIRgK2HyrgjnyKIK+9cC
Umj4RzwPZbh2xCmp1GZf0NSNwlBxK/6Q9uQnxpmUOkZnHF4uCuJQn+nRsDgcW0h+
chJB+nitwZoGkzJnGCRZtKG+bHWfwwYxAfMIPx4fJhq0Gy0mk2OHQWyQ/jEOf5HR
X2h5VboGbPQUS1o8oDbakMujloQHrajS6e+PA/99r4iSahkwsPXDqiE7YkdPDX6T
8kVduSCsUoiqisyfa3nz4LOgi8mwuzWLjrVlgwScSb92t9aodsJ878ksaYQRGT8b
rMI49sW5Zml5ZRhl8Y893M+09k9vd/AACBUoo/Z4lvSCbKHr1J9nyNA/Iiz8/zgH
A9Yle2Q3y+7QkQQA8QdgMPr9JUTdO9TRz98jYTriLlKeiUBC0RdF523CHYxuD+gm
ABXwQ6ViWoddpObYW3YvNM2Mnqf16GLYF785m6LLMPRcllbcqMS4Q7e2gfCwk8q2
GAuennmk9hrvdp6SkIkp2rFuKjnzea5r2tG4d57QKB749PlexeNgF+CSqUMCjaRq
hTxP3rhOzW5F3BtEx4SUGUGEVtbdr+fpHaaVDLsSLIjPN7I8JlrEIJWClBD8X4Gh
PAAAnQrSAVvbMnFuNB3hfcL0NZbcPh6U0DaNm1xk/ITN9+figRKr8z1d30n0JlIf
PY5pQbC5F3J06N3tMlWk3yH5GSh1eWIlqDNFaQ6nh9y9oIEPx5EMHTSjiFkMUY3o
xggI6B6QE7D7MPvSsH2BhgvivF1CZDugutfgbnQxaDP6zZjA/IfREXyG0qCceJjL
EJBjHk8EUlcw7wQUOD0c9zs+6KABbo7ZT0qyYZRyj6WkKwqk6bdds3+ImEEvfUma
paowgGg7Ifopsy2PDg9jK1551dED9j6RjrxQyhcLMKrVW+n35tx8dyFEUNIGaSi1
4XuDpjslC+VH1wqDjifWSZewdzN98C5MKFlJ6C9ENcbQMPpyxb+sr9rTxJB3PcHj
lR5W2ket8iIDr3zDT3+2OtMILLh45PWQDHQ+TPVpKErLtbIg9RjpM+xVg6+6e2eF
D3krnpLJ5kpC5DxWNTF/goU29TpmeFEFiZZuw2wWhngE3YW/7tcJRKtGPbG+mRIz
w2AWm5aeVimeSvKlQTykNwENru8ZALdGj9ry1IQYcrxuFwQdWMzENcIENKDA61GI
ySohZdycEPJJDbsSxxW6NU08LdtEcrEZ6dI06XqDVFvq/V9hgKoQaJ0x0CjD8aS4
oy3M7wJNRTLUYeQ70F7mK+THjjGLbrou3Uh0CWWinjWD0j2rTrYBfAQBlkagu8v9
A4MS/dvm1B0dlA346FfBvobGx4EooTxH2v7iMQogm5f8Gq+scessIrtUBXv/hXoy
s5E8FbEKJxVesEiXCEEdV+870a1QfNvSFh5Fj108XJQBe+rQ61MITFhrDAhPQuP+
gVP+BTPp5NpGI/d4WREmVt55lCjPH5SrhWFcP/iVqRzRs9W0pnUQ25cODBsQSKPp
T/Zj92WQ8hZ0razStO78QtbtCukrykFGf7t0iuym0kiHFx+j0QA6TN0HD/3GCreY
suAduK/DUuIAtWkaHI44MFp6Xn9W+XxpPfYWK86ceLyt6ZxoLnSQ793U3DPeZrk7
aqlR3w7YrdJn6niawvAHjrl0pBJ0uUEFgz7iNB+XslfllTfprJVBK0JK2aRJEgLU
x0LHLky86LvWdEV98P6oXW/dOsEjWR2ybRpwGnNfQ/7JVrY0ahKBRTQdFHK73vww
4L/d/RPC6QAymBoS90uyd/KFVIl7SfXQ0Mufks3hukKiJwH9Lh9rcEKGAm4gQ4JI
ys8iZpSK5rUIPkZNpuSYTLrM97YsjkUSsKoNJSXwoDIMKZ8Tz0QRdqV2sNmwpnwa
WKMy4iLHsq9K056kPv+uSL05LWYGXqclr1te3Cu/pw2h14QUsYW5amsnsqOLXzOt
aFzqRFPPGhi7dApv8e82w6pdCAXdy9manQbNO0owhxFA9rcnx4WoLQo3x9hzSXdy
4qkgFPgbRB3R9kPJjLuZ2bkpb34YUcRJk5yY9cV8ZAAvxYtwucNjqSTdtkUd09G2
iJH+sKv7uDJ3tDkSvLH7LZSyfxwdVT4EpDw9ZbnN0IvwFqh2dHPAvrnDIpj2C0aW
23Nn7t9uZVtmrKWGtXVeptcueoc8L/Z5TBnoYFfPDBLt5nExmK/1XcKwBiN11dEt
lN/41CMuWV+eZRYoIBk3bYUGXJaJIoy0Y16Y9zF4pDCgM6p9qYb4X+HKLrUyEMmI
nrLth+IgpuAOCrN0dvP2pdcRN7+oYxG8kl8MP54xBIYGo3uuz3s8IHqe2Svf8fVC
x2AMJEjdWEKZZEdct9rhEmo0wT7Pswy/yBFYZu/t3nxdN0+GCKs9oNej3fc7Ze9h
gJaVi8SAOuM4Is94Zm8bN548Scz5+4TxJVxUY1gI9kvr2jsyZe3i1K+Z6a5XLFm+
XpFSQLvYAoEKQntTccJ6DcInKj0ycqMnFhvYrykELcioe4K6S7gCMd33CJHTM2Yr
nqb18O+elUQHTzK/fLF9wWs1Ci3K/ujhk/SnAZeIKVbF+gUCA1labqpXi29jX7mM
CEkuEGIw3K4fY8igYFDJVR2Shd48FKEOUQp0d1Gt5YEci6JZ7wke9Sg15NpQULZG
JHOfdi/NGAf0AYQ79JKSyQ0a/wNh9htBbKO10CsaqtCmYVyX/b+jQDJ88NxOSo5o
Tup2zqW29dOVWHfdgsE78PW6aT1u3klnYzXNzM6IjjbJP41lcltBJWZHvQBiw/Vj
3XmjxIXU/oh+FSS82mQlheXlDOd4ezLtVgXJxPXUPfoG1A0CaQqfL0c8HpOaiIGd
Y7lynttMGnIn7NcZ762NveyEzXOq79AjbuVUC1OztG/6qgOWCMFpzctZbxgaGFV2
CMtuLLPxpXpC+/vACDlR2sQZaDvAJyDw50vi76NiBnkIBzfTg9DR99MXDUoX9OW2
ggnLYA8lR9ISti6LehCXtFCly0P/iVTgs2/WKBuECXhZIAFMpwA6zAxIOYW+DJmI
R+6hui9YDN+dY4/6UbXKea1f2bkU7exvSP1KtSWx0AwWP0ZW5/z/POWUiqQDrjZd
J9TGit4fTkorotQQgNqqRVRSdOrKmtDzzAno3h1LB9CCkWkW8DLJRd4XJWXLXnIk
f5l/DTcttV0ZS8w88MyxWWthBmPBfDvLDgCiPuyMeeC58cQMU8pGJVqm0N5uElRq
GX3AMN/bbZ0wLQUwFxeeXYGz7vplnCPXcqy+dg+woyTaRtwBoZjhbt6vcvfubjiE
4nvkIaRwwwK/I/mNDCD3696tq44V0az9Vi0LekDdxN2wUDQUJd2rjWJljVdCVWUy
QLYyzYbhttpRPvMY8W/CMHsfHcnT3idIg6dF/+JualgOagjDWjEZOSelK8H9VGgl
E759OHS106VByt3xwZh/IdDsNHlZbwygVkHKm7cidLXGxsi6WTeZ/6OLyiaWg+2u
G+gjyJ58bBbt2swBYOobrvg4IoHgXbI86Ax+MhzgM9Por2DXIiTTUwUXQUDf+rao
1tOp3dwAz7R/5rDS6n1XNahlH+p6DVzBdHKTiz4hhG83MybRfeb0/nHhUccbAkar
C1+WHTlwY49CK7tIwldA25JY863JqMvRWJvxAArXS8CXhAGlRj0kpTg6ZJAbfHT2
vJk4TunUKpAYYkh68L9EpBMb2D+2CN4tqxzuMhmuBfFX1Q85+PDv/guNZ2jKbXuo
9L2j5hD9Gj1092bzlzjZzBx3Z30QyWY/0e2VAvUnoyUdAnPM/T59SCcYKLW7pMsU
SXBWeC8P3dwo9a/WHEGzKOUn4BNmWPHemoo8vvHNsadbotSAzstpLz8zJg49eLsR
S2chvIB22FVfcxsU/jikUflV1PXMmbm9CUGgTr0UrI1KoTu6Z6ouBiUunYt9sb/8
F5KxuXOxCXfj6iIT/kYRejIO9cYLMURew32KCcTh3QjNaDGjxUjVvPBYBqPVXfZV
q6C49dVofOv7L31lLm5N2/Y8/vw36M9bcuh6VQxdEX200ZYMoHJT2RrATnWyo8K+
kXavYTFYoI4T4u1oJEACdTlfpGSdMk8cYjBhvtDk8XNOGmqor7vV5McLTCcgfsn6
kC9y2MfDNwbKq3MWKkLfSgwMH2BdX3BG7IMyJHgJVaYIQ9mRmgHQl99CT++fqjHr
SfEW9Yldk+iEN/97O2aTMPIj4uX1XJdJeEavykCEnTngCrfivRWxtI1kboPqKMta
UrjYcIsD8S1gqa4L0lYZv5qlgSv7PQRaTtDE4M4KmITlIGltDzOZUl5xTq303mbd
G4dZclyZ9taIx8CpZj3hX4frWJbrvNuriUVowLhNxjifT7I3UBYs1DFu4A5XH3m8
XT5wNIpY8EI0tprKbFugTBsNW4UMOtud8e7YRqjahHR/0TgT36ydUazny2LK/jXQ
6foV+pU4mGs1HlY0YAMrnkURIOxU+A+WGcqKCjWiq5f/HwqhxkPmtgPOQ5K+LUyA
/rTXmzH+PxgX/EEuUvobJB8fkw45thZ4uGxgfb4j2nkiqUU8DFD25hOWxRfchX0K
bJLEMA3RAdHezsb3A9ayV3tWqNh3dVsH+a1cT1usoDHpk/GXi+4GUUP8VuySuVi0
vWlPHMSMaqilqOpU3NKDP0dzbrIIZcneoQDPRuQsCwNwoxgxhbcNnBAnislIU1Rg
djoLf+xT/r8gEyDd7Y4LvHWgGC5WObPiGRb3zdnmB8jPFFNvWr4CBndFQYodrRIv
IHHBqZw6tTgBn5jnRzLVGt4xjrVnQcQ3WcEJBL2AP69hHndBNBAfLIhsYrBlzOkp
tDEz4e3Tn0BmYqPfVx4iLOb1WPiUxrlaq8DEblTMsdixc8Ob7/js3jjxfW8VhiLX
jpE3xV+ry2ZnCH122QuH2B40iSE9WmkQYK2VxdsGYcnW50pMAK7VdhVu7EPNJELo
0N4YrhRerFXhg5lb2RZK/1pDuctwrX3JoAJXL1L8vr3mTRhw0GWNBbguGVlDiNRE
mPfnsfyvsh+Xuir6d4XgK/L/gD20+UMayMcZp9U4Ky4ZpNNbJ9qbkqgRiELqeNCA
bVMaWbE5yOjOtHWFObhyvV/OjP1vycwGu5JvrOE5BWu0M14JOlqiKYu+suL6T0k+
axdeHOVj7RHprTWCFcgQkP1bQYWAT9GlLO3Q1GT4ngt/AXGNks6BK/eW6VFFUB0n
eeq2E2QzxayZ4NdVeTbwsWT8proTxMZHJs+Gw8dlfJNfj4vg+04cXOpKRFEXDG+P
SClmRbglCFI+9fXtNq6/5wr6MWrqHWxIG6+bmZsUV3W8++fRismfilgQGEd5Ksgv
QOgXnA6/1v9ViYMvzQxQCeulgl7kX4/HSIWapof3AXQ1b6qpKji9OkwbQUTQ/xzv
kKEQseEXn+fMEP4bfkO9+z6a9IlOqk7u0u59i4T2wD7Vh06m0XNxsffzL6zvhOEb
KllDCy/a9fHjiSfGHz1brkfHHryiBXpYfufXj+pHQJfU97LJsMz28j2HEPVBVe+X
SgjF4TeNS9PQAOtKF6gI08fMIg1ZxPu+n5IMAG6OcCttdVXGrOdg7MHJDJIYwxB7
ZdKipKcWDHD/XQvkjUq0gG0Oj5MDypJPHMdJvrR2jbxv/R8g7Z8xQs0A1Lc66dn5
b1pPtWVMm6NmYmKeDHn02eqnh//7QdjBVVOdvTjNIndayQ3wZkRm1LerlU1J2jiy
aoCiF0ranQD6Q7Sl88EH/5eHSkBD9gHmwyomFAXFsVmJJJc5QaHLdh9VgCyEkulw
6xJnZpm+bgfwS19vftpReAlsd04XF/NmK7QF60QVSM8XWR4YXT7Nfa3vWhvp8Cx1
9Jz6n4kyQaSnstFVhQsmT47qiRoKD+1wMovnxM6+V3fPhNkt4HhFGTmGLvb1R9Y9
cL3mxtIABUUnhtI4Ft1DE2/bruU2abqz8LT2U/6x1pBJmZcpMVqS2AsGj3m4o9XW
XPXRUYTP9NLE2MDACamUf1eVu+RslZrqo0caQuZ+swSsRlXhZIRbV0QxsJ24rBlF
uHtWlxRa6yrULEvoAIjldaapqJ4yIEfD2zP4AnTMEqLGd4Z/h7POupBfVSItsuIm
WTCwVME2X8QC/T/IiEVg5V6MKzKt4aLazZsQ7+X1hHjeEyQ+BjriCfsjxcxXmQH4
QnHUV1E/pSh8J7DsMMaAmLd0+nAAkFZV1euy09RyocLjips6m/oOXYgOXZOFxfiA
ZSGHGVAceegJpcqd+654KUt/W5nZMVWToTUvDoCGTEXr3jnuODy5x8mp0h5RhVK+
hhXQ5mWAz0iS/9ZQLQOYqUByqTAorSi7JynRgiGy7gqaTBVYFsfQ7H2TYcs4At9y
biejk/jK1BvHg8r4ZdQC2Z6ONWShN4zrr2C3uCamOlejK9dAAte5s3MG6p6qmAUF
y+TYm/suUdng+z4dhgW05ItroezU10M2IXvMBtxUPdi3GEY6mCtcw3c2Wjt7xTNK
b6ONC3vqJ1L7Hk8Un5uIvO4iqsU5awzaNuOBsOYvqiqg03y8U5pR7hRov3mR0YlJ
THBkfIQmF8zbb35Ac6dMVXKbdDoOVqaXmzHElhCW6Fuomqw+lZE4V690f3dHY54o
oHl6oNsZwMZtQoLo3vcdPc3p6W9tIqyiBWX/+uJcYuoKigr2JVB3t5bRMqmtC+Je
iO6KzPk868uhe+ZVoy7z1OLqX8N1VmNfglLjM5NpRvllsGrIra6KyrObBHw6eZg9
/rSLfbxq450yq2GVDHuPYeOzaJNJ90aL9d5WtjiPajMUAEAGbIGB/5agZqxbdvfI
HZbqGiKwwTIuOiApvlV3RY6HkJ/gfAEDGg757xoXEaAuto85wkRn8rhUajn6t4bi
ukJwO/ntst9P6ex9JpZ0y3Oks3bpThZ9CHNVJ/bz8TJl6dcZsNLuUE/VON9XXRpU
bJfgcn/nKLBJclDEPXNn0p66Uw1/g0ho1o3XG7TiIItN6G1mn1t/wFReNcqkSsm7
5ZTUHYzIj4tAF11Vx5rjOw3O6tbMx/87cY6DTCzLR48FGNdkYzZJqu+jwvieQ+6U
9XKhS4o2X95FUF/rMO7229YZYoj2oUmv5nJSBda9+npI+D+VUODF52MTs9E09sIr
om2o5cPtzFzotJbFRknt/Y5AkXots1BxTdXXlVo7A3Stvj2GQrDMKYUGv9PckKYj
f8Y5m5FtnL2EqtxUC0XB6uuOwlmNm2DMUkDXKIbwNS6whr8tfC6UlI9mJkNwOaEh
baPFsctUMNI/Q1TxobfV7yBo7jBCkwkosMjmcGlMZrXA77gLEralCevMSNmgyL8s
dNqotoQhAGxOTIVTcy3NoAQXytwzFaqiZMgoz4ev8puAf0M3nydZyPNvD5WSvu5m
R5JW2yz2YOfpyRZJ5cAgjauLbVr8NIgXr4EtuqIWvXs132hxtcWWU3kLip5JLQj9
yvoFlFhPoG2bR01sdeAAkKCErE7+wd65YCSzyzuLQFe3NMxbpTXc2sj+eZl9ZKYp
VzOg2c3OeOkEakHsw6q9XHswbcAurS2o9X8fr8tX3agDiiyF5Qp+JX7tUO3YkqQc
4LV1xqW32GmhEw92JJTZd4y95SKCIGOhsUv6yYYYcU7FQ4xnltmguJSILc3SEHvf
M753u7e1YyLMxTQ4BgBP1GXq8W7WTo1rH7URKeyRMKMXfSOipSGQhf5GCAqB0eFg
XzkdqsdNFWZDJCu20cn3to1NBftMYsxEwAHR4LBk5jVazHcQ19K3OgJBEmhcgfMX
RxlYPaB3cqams8iZkRCfDNikVGF2MsH4nvros0/RP2DAi8xYUoxcoHAco0FptsCx
eBb8A5hKOkeTnKJWvWwsxa4aOK9oQ49kjPHoJ91jeQdaq86ObPdr21Y627efRSaL
JcGUouPyrHV1das0PzGuIUwM9JJ3iUGS6YG3ru/iIONvepD7TEwlF2DO27zOYE4V
XdMjBovg57uCnpsaWrBamJC3q9fHniOjygqn7Zx7+/ykpJuwEdVqCNSIMEZk+Gja
4CV/bveCOJOQv3Tjd7maIYDrafiKqx8bxsNC0xaaEpghNriJp6qfYc3JgGkLNcW+
2cPn8rQoWDtyFrXqTQoiKBcOIRQBzzJpztYQlsCSAUg3fO52SHKlvA9jMYC+EUdh
qQhXpFgvjTv6THUF1Ba9SdLJ61PT+T1R1sxkoXk/oNl3vkOPPX/hN7Pdj4ejAgye
FtKGFX3HPL4r+ooxyssV1jFwol9j6H7MVFe/hUMwXHl1+nqOyoMjgyGxSlh46Xpy
IE9VabkmiGi7c7LIPJ2luuNm3JFdgxbEFfX64pSjL1bFSAnB61c/E/ee/1NrVRP7
CbJ3PbRhnP+joq0FIAWv2e+6llCfAFO9TD9PwwGfSjWaE+FML6V+NPzimX3vMywp
5a8tBT0FqjVXVy1TrfmLCIi69/uODeeCiliHWEKIMngbQ9sHGvGRgI1Dk+U7z4+U
0C4aFzmvklh3GfJzJQACDYzZHbMZNci8uLXwfueL5aovNpsVBtyhpuZisKxSf1uI
++BDQ/8sPgGxPwfyQV8OtOfsxnyTHm9573gDTFbNcu/fOfuAB/vD9FcK+j+vXheG
JSbFpCHbHEOe23VV8WbNTtkDsrM2FiH0CKZL+pdDM/0RIuBJcdAo3oNChupO/box
HBibwIGLJNkQUesTFsziQ+C/LTWEeG9d66f2F3i/U28oICI89kxe2LmjRCZEGpsl
7ZFh6NpcxhWx1esjm9vGW9Own1BQkfQi09m7hePe9enKwzT8h0ccRtGFa6wf5Igr
c0ILFoD7rLRMaUcoey1LupG2lsJPxzoq3s6dqh2kH8KfIkkeBGqUSrbhuiMdcGCK
sVpbc9eyfb9CwGt8mbtt5k+0Ln6qfLRw/9tasheaagIGRc7HHJFV7YSBaG+7jWdV
Jf0Z9qSi6fsU5FVs77hoQiSiG3ckJ6aN8/b5D+gIw+r66qSYvsMEs7pHjfekvPr4
w+SW2Llxnvq4HzW7lNTPNt+cO8+C7e40I3K4V9mRDjosD+OFC15uQKZZjkJqNMGi
/gjbvgIABoKdQP7JCNTNxG6fnZpyrwa1Ukv1kg5dzG50tmI7F7OhSHRdK15DKXYt
fq8NLXrSUfKNiO0uAeR9UmAQbVRsFBkagD7I3cmZEtrvpQEGNkgPr++mFxOMXF16
tELGyurMMAYXOwfxQLk06UCBobYQIBXi3f47H129sQhAHB0bHq2eBRmHPpcVp4p1
8G3g7/uv5RXHaKIF/I3bW7LUVR7xM1NxkiGAVIyJv2t1ZOlTW8Uxy2VisnHX5Rp0
c4uanIieyGx+YVdpE7ssZIMKwSIfHC/ly2YDznVUWSBuySN9tAHHdYqEl2oPQFI+
N32EdIOTShZ3JL+6rZtjxxG7A5fYJF5K3uVB3BNNxsi6iaXu3E6B1WRS3CTkE6Rm
bbU3Uke0so8H/dsdNdrvKXzeEj0qud/VaJzBBJ06EScETXWb7oThDAoHYIy2I3XG
JnleKBOFCFp8QnlITRSYqWvHGUGZwyNsPkh4GtYFYH5lMcL5rMsQ3jXA7lReL3La
P2To0QhIhoN4H/79rJtZbXOfGG+mXAUjbEWLPYEkLALNmsIaoqlCB5i7FNkLPlEm
b73BtR4ATStfTG55Ekqq/PSMtzfWRIFMZ8OcGB5xw8irpDc1KEoyDvgrRZL81JKh
P+zLRStaSdjojHkXt1wj0U3x3LFFpp2TzitdpvjVku6LnKh6g5NvsxxJq+MEjCCD
J3aTTPKW3tss37Lq3iYBA6bmbRXYeq3OWLNB+xuPMUF/+I2e8zwfbpNyi9aHAsR5
891WHBGgJ0NB6WG5flNang9yP6ajQottGqSX5j2xLsIJOBp+xYvW5F90MvxpvOKt
vJWmNXOfPuY1xaDGz4llZS4tiro0vkNt8E4PILZvDqtF5eUQIVW+RaiamtxGKpMF
X1uyRBbc9AWO3u8y5o/MJgc4VqFBfl3sWkKJU7YdJKdh43r7346YUzIOwJXZYgXC
VY3SO4oJ0ZaAXy1ZQPLqOZ1sZxvGXybz+c+gyim4Oqb7PRJ5f4qXhmVNHVrTDGNH
9UM1UMclkrqXQA1WTkTqayDa473PSHfEwQEVt1NJqT8ri/oOHj5n3AsyfNZ9hBLB
WAEIGv/EptXvz2FphERcu96RW7GAijH8T2ArxIYpjQUuqITVz9m8jIow9pkpQXYu
TyjUp4yEcnkLmhoE6emgqZ1YGrPVvEZW1R3wfkC/PVXn4Wic4iQNdEpejb2bcNUu
gqXYV02B0ke7F3JT391uWZDpVg/hy9x6nP3q/WjjTE1bqM/4DJkqaPSr3yHON4gQ
G02SE+1tgfqUwIrpp2rxyZtiQCkhlQc91lXSredRJBCrzX4t8xGq4MetVvxhy7FL
bKgc9F1hvHCTEp9ojwHxe1z/+TmuttuzoUOOCwW6ZeHdiDz4PQZuR/2KQqhvzUs4
oWFguBQBT5HSJhYyZs2+ZmNn4MhQOdpEkHJDeq8jmucKEpYFOgBy1UOV7+pSTjMw
qEap4Pap1Nsp5mkmRacYxCz8EevQWj+RFXYq4vJeCfXreYvrwFqcB1zsIrrekR3P
SAOv8WJaGVXgV/JTq6Ex5oKvyAcOKSR8ZvgxGR8ryznzedhZyrzameKdBR1LxxJp
Iza5CGvXKbDqMXw0EJR2uz1zLveFW7Fm1YOCLW9vWQ4BasOzAEmyItEaz1dp9UB6
Rxtile9x+jWDwbKOm34wy5KYTITdTR0Qc9Ldye+yfHWLNLL6T2VJbvCaKS2uVUFY
FByxd1i4IwAMaQW9oeu9MBLHxmkzjawVXpnoQcwG0enX0YOYwB9ZJHm0ORzMVhWX
aljqEc4VO+Y+m0PfGovof0XeVQvEt9ZzkDAiINAQyY+w1VG9vjcyotCbfbwJslMz
xFkyc46VfLjPzy0JSC2LQvStjBHfJAcsJvg+4Sjx69C6f+LACqnA1CpeZJNk8wtr
KWzt3PGHHhfis+Tsa+aNkiiTVVV4vgx2mFV3r8xTASbZkIYuqgge9sy7g5NEIb64
XIIXLtRjpgRHlZoKoaAUVfiqEmVdt0WFGqHAzSTmyLVoxB2UIobzUxWUb/gI/EDh
k+rcYvOXx5Xd9ajlUe0rVUEqWCw0kdFkkByKxKWaRTHc848mo5Ij/LsVx20nqNOs
2m7b+QB+dnk528l0vmjw1mbkuvliVVxS9htJKGE//Nsr/HQWT1UtT070D6mIxI+r
VwjbZgQsh+64UObwGixUWVcqe2gRI12HsX/at8bPTEWLGEHmwr0XlBg9GUJ9ftHW
y9jUeKnUMvHIQk2eaoUQ7UXzZq+eNIqluTX7M+XVdZMcxwPSkqDwotJneV4ulF6X
6r2E3IMyP3Hqx++4g6hjlftSFIeceGHGgNeY6nJHguL7MdDbD++ZPjdLZCYkqefL
wlRHV6v95eW2e3iFLaYYQzopUw6gthamVskHJYhmwk8yP85sK+lJP+y8Hlv0acHy
a4dn2w9o3AgRDMOKsjTlz6tD63KmQRZacRMmGJPmLxXCLmzfjy3XkFkNzbaFa26k
KbSRp5rxveDZ+VOF1HxqtLGbp5vsfvj04ftmoOd0JDTzD0WYJEcithNWUoj5yTk4
S06HOGhUjyxwKrxvs5vR8Kzf8yKJ3zv6fH6dCM5tcYXZz2uSUHNgCbkmrB5MKB4m
RxMZC8lLoW+LLPw4wGW8gMAp2eeZZY+s9ZFq9H0ZUNScA8msKE5IOMpLoeYrYghi
fbYsOV7TKllr+UEnKu3qZ1IFbLHjf15zdqkNuVFfXTa+FDkaj6m9mrH3VNNfnrXE
FZPezCxSjq1I5V4WtRRuoQp/KOjy8/q3Y4eujpv9wZSrrvQbZWbidxsqhN9T/nBi
aNCGlzP5Fy5djik3+XmzUpKj31I42kbmE9vWO5d3sj9BHjj+I6KBVLewosqPnzhI
RyzqefKGZsOdZSl43gByYKwbXr4/SRdOHYnxtEjYR/IKrh4sTfZupLN4GlwVM0+d
TPcKO0auMcNS75DaqIP/MfkWAVJ85TbaZKVs4FlqBaGA9BBRZIrtiCZ/p561Hts+
GTuPw7A7wWWwv9uMF/PZl6p6fhZ93rkvUiRG4GTRG8YoYEllXmN+AI6JV+IqoBAg
iIfrhwsZj2OPaFzTWnnsm1XR8xglEYBK2TzHNFpZA/2RfOZx8qPuMYuwyICX1lzq
P95a4ZpdTFWvrggI8SM9hndi6rT82Lv7q4lxfkz0aMR9wZ+uysm7Ag6sMWTWa+VO
7F8dB73lG/4rXEN9iwMpn/OWviGI0WaBcQH2WST/+pmFiqDPN6ez7Q4GKivxy6O5
Ypw9X3/AALkRFp6NoR8szAZ64y3yIg2NhSh8X489qoyj7Hg2lJIMo7zc87xPhNFY
fK5545Ms7u+SUq8Bn1gJOHW9QcMPI5QrB0OzZMFXtYKiLNjZufi9+S1JqqIMfBja
l7NaSOz3g0ejVhMkwuUWm/OsxvmORI1m6Ay9IyZ8qyE0HBOl2777OXLhLr4GVnbM
K1jYBThgmu/nYXzGvTIX+tdGCuKpX0r8bHxihkPxLchS7f+lw1lXYHEallghEsO3
c9ly1xJwIn5ewa13kjOiOxVRyNilTmfUrIlKn3aiwR1/c5yRcu9kGCN3qudxY0hO
qw6e7qBI8ZhuskJoRxucL1b1qyYO7hzIEI1MyOk1rEgEoBK5U+NdzcN3KQzI2krg
1ULnCXcQE5Tl8fht/EaPku+tqIphUaKkniKG50VPBglBnCFUUmT/uq/wrLEXiHdT
AHQal4J913Q0IxIeAyiPKawlbcInbX58J7f2hjfxlY2JTDkQERHCovGxz7DBTxj6
ELor4EL/ghfppMfRPZ21xdOB9tnRAzLZscRWhYyPxT+Y3na3/8VfGkCA/2CDBabm
mp8zPGtgR7/6cQfqzWc7+Nwc2m8LFgZrZT/jWqjm1VEanL2ySr4g10hC/8YmrRBo
3uaceerkW+6BAKbH5AHRlHiYcKDrm62zGG/p3WYmt2aabyPOG5PuE/i6rtBRSx8f
USGrt8DYBOPnMO4GoOFb4/KDZjbEvuV1oOTOlKW78IqMbtI7v4SrFjoJCOIPWPui
XxXgf4Ceyl+dOECdqBKBPoS/31xsqj9+GGDLXCi7NdCtnv6Xxrl84xwEPeYYAGsj
WoHqiSY1CVw5NcF1/9ITe9jkEjfd6KqUBgK5T1cGS2Tgu3QUR9zSq4VYqub1sqnT
31c+MG+1hOdsK93O8xD8f3+TLJnRLcz4yE4gdxWZszELOnI/oFI9drO5r/and4mp
P97UtNJZBtD5kCnnIoAn4HrOH0G5Xo0VAfGpxoffxgNk60799aIKdNj7w1GLSbNa
P9ocrz7DgUChwHVCAiRxXnMMR0umNiXu0+PFrTGJ3Bu7IQm26QpU1YiZpIy5OiTO
cQyyU/6S/IPiq+w+n6/mmUWKlImLRvl9x/19IC0xpnG8hLrkD4YxwQZz+tVeSotJ
ivDlhlKyD4Ho75/66BS7002kMHKExe+setnexTOx6hjL5g3SF8/1BV5z3ZmssqlI
H/t956BxN0iZcR9tNw7xQpcNWiaDm5adPlQc8I6O+ZkTuZebKNKQ3qo81SIY93HP
5irxQTjBjZ3UCb0b88gnD5bDB/SuIgMG5ySFclI1/Q8Lvtd0SQON896tplu1+2Zi
rBXa9EiCW0sBbYR6jEra9viuxyxBlSfe2DyPfrqTCa5zP6G7E1IHnup0DC27tvtE
dCFIw7H03hbF9wk/5D5vQdfK7OrVYrezvYt7wd7VBiVStNUVGR6onMfHpl6+aYCS
BOMNytzx8BV9YttWXNNqVVPI0Nc9U+q4N3e79tZT6K7FSylxixrFoWipigtFV/t0
FHS/Ae0IrtCmj8Eq+Ya1XERyTTzpsj2pz+e2r+u2+yVAqxaIgLYB0l7L7ucquNtX
8OBskSTM9MBxwEKzcIL3Ka7liSfhkpktISCKlsvWcTO50+Kgc7xJ5WqpKMxqai9O
u7ueVUt9EM8IU44Xjr2YZS98SpcqGiI1cZfAGdM/HksMmMmiKrOSV8pOoUGu0l86
ZVQn3QphJpy+M0c7LQi3PENxa0yecmDeaewn6YoGAjzxZMZXrlcKMMEM0fkuQa73
gbuYfGSwxW5/RkPJp1JUQ8YVdYtM523vgrviDdwXk+iUIlfOuynYfvN8CR4JywmH
kDIlA5C2nR+YpeX/8EXuV4CCC0ZSKso9NvL+p5rjfhMhZEGGUXfiuddm0eVmtU3G
8jtQKIamw5XNvrPsRbCwNVNYQB7Fr8y4UTzTyrbIPCXg/r6vMzH7ant0rvFQ6ev1
w/ZenK6oBOTZ0WA27SefXSARnZ5ZixyebJHzZHtMBN2U3VGVWPrW2U+Xx1C88y6D
33D69nVkK4KK+Ey3p4V2AJCjGjUBRB3RkcdI1o5oY+ud7dpeDN31ubOwVZFQ+k99
LrmJLwWpi2v3xOsjNqHjB5Jy2zswgkYk2jsXcLUxAn9IMcctLzi9wXIdYVZzZaKH
IUiamcYxxcuEqQlVm+LadYx6klrf+/A212Q3RDWLlb53Fl9OGJZCRh2w2QLvsnhy
UF9cDGjYWahOuz8dX3OF5DraxS2tVmWWLRz1bFWy6X2+21xV15V/2YFqAATZcFV/
xQSEXWWUq7bhq+I8Ac3mY+8iahfCq16AaZaGH3eKzysaw3PfgwfxdnwAR2VJodrg
mu+4/FaCMv7b2J7HW3+v9BtC2sMN1jGjL+igyPAWWbvRXdiTuCr7rbEsJpKuhntE
gQEzXzr3NrmR5s6DlkOJWQee9LmYu1OhIvVJmaCL2KDzbklUFkWg2NAUHb5TzvC3
ZdJjA63PBgwu6uB6buwNFQsr5Bpwr+Ry76Y2+j79lO3XTclLl4i7bMvhgUgOsoBy
iTvJP/txzKJ6fptLhLrRZ5IGSAL8ZNiyUR4lbMWSYKipwkIaN/aCaGta2g1Fk8HP
Ke5wEhIlEhvKP6AgT+ThWdoeGiRwBDt3sXK/pSqTKOySJCZl2jAdJ0fWYR7VTSu/
p/+J4FxxlbMIRLI2bDm60S15HEIPOy34Gzr2xAb9RvrDpZXgn2UQaZtJt0+WAc2C
W4RlmkcR3EOvvHvNmrl9hDdPW0roS213UaYvDKOjQGSHuNzg2MH3FzTkTo9i3pMY
/pyaThn9lY+ReJBtAG0gboTyVEIv1tOep+4tI3iNhIJ7AO3jGrcYj5w8EPY0iLux
fBUXT1s34nS6y6f5pBwXH5aloMM5ObgB1t0mOUrr+Ml43WC8rMDxRWGs9Fn5QvMi
81RjN1J7CjDzf8aC1rsY6VSXZ84zpiH1YJXV4/4jYOLob7VXdOuLdz/Y2vG/VU17
+491HKNy3lUJooOk+HwrxAAVoXoMQJlolGNdzzt7bj6EyqeluANkfV8FwYP00No+
Nkeh/jAaY0q4C2yeGk18oBebIjONsaGcHATXOFS+Rxmzu/HMRA09eaEQk/FJ3DaW
LGP1qSPSH5Y77AQ6W/rpiT7ag2ZX/xPeYkj9yidr6QlKG+Cd7+WOTwxF+jux9xWz
9ed1gvfrnIPpfVJhkRaWZ4Av3fUCGPGlIX7ynY4gFeJ33mZwajAB2PH8eq0OJu0F
rCGUZ/7SD5ce9RkK4r8fyDwQ+vj+kd42+Dh9RQsfDcBmMtU7C8liIqoIqa0gw00a
FWVLQUH3257WX9BF/y/lNOyLohGq9BlXVIIH8BJ15HnLmAk+ZE8F6M2Qcg0yGmyU
J3kuWgZ3LHndXptZKF3ZIH6UB6AHWbHgLCGp1gt2Hoq/iIj/+J/Lk34M89QVvxdI
THXYkkZk5WPywDHVhMQA3S1IOlQyI8+3cwovZjONKykDVoKYvZUerzyZgEZo6UWw
am9MUb8kTE11Jzuj87opKTgrR8lLC+LfOBJB/p5B14LwWL0fQAna9JPfQ87Km9ai
74AlNL+Cy9FIby/S1BZeXuziZIaf9nQjkXyCo7pfw0d+D+PJWdtDmte24Mm0WXOc
grcStYVXC2THronslGX2gV7lXbegvkW6lgif6/mJ4zVW3qAQDwhrOttzQ3o8rOf0
mZCamN/zGdfeJQ5wedhQ2wx61dJGN2n6acKW7K0a4oFQpR1gZk611OpG1ZSv+/mz
NKyzpmzgAMMi1iSyhZ44zSJ71a91gn7KThsgwBuEih5W+mNwdQc9Fkjc9Nx8qIbH
l2kLt7MqRKPkDxoHd5bYKYJw36iS5ntjBBAOKowq+MhalrgxsbWD6lPAO+Z7fqNy
oinoO5nwjWdOCk23+n6VKwvBGPMIyCuih6wSF3hiOJW/BjOr5ReDba7IfTaFnrj6
VIqkqW1MVG7+OFUK1F1Z2p+ZOrIJecL9TebyQMof3mUdpkMiXAmYXZ3Mt+CRBnHN
ju385GoWp1uoHT/u1FeUowM/Qi5Y6957Vw2ewmEVTswRxPhotL1BcHfZHChezPF6
Cn7WI8XehG4xebZy6pRBeAHGiZgwy+8vMiT/DWbQyxtPWDC+9wSEoypVp5vtrV7t
FlhuBb2SfIXeFbBT1vDucVrZpP6Z7gB7mmfZjIDJhSdH5iKqoMaJTCUsLfSCO/GY
yN8w+zdXls0iK1Ecf0ftEY6FpV+NOkh18NFdck1xLIgjF1dFDe0YVSFIhYCNdh0e
L9i+3KLPS+GnoF2nLSUB5OzJ49GmkciVd4XTIorPsJH0WXVLW+kX5Ld2xXGBiO+o
ZxtSgdod9d3KdHg0hWiWvqgqZNrQnO+BlqmGC1ILJU6CMhaLYkXtXAJf4OSz4J/M
V0k/SEe5eNM7DSSF0j7g5jQAgrB2DRzI6Oy+GBQl9n6jx2lYDTASp7vfeVa8ZK0O
YaDWh/XkOJCUDk+TfHEpRGWjRpwKgB2nTiHiawweZelQkQ/DoPo5qANfnmHO10lG
29PKIlLzC/DuHzaPzpMFinb8jdjbqYkIS7cfRwsImSJCoqwG80KhFT0/u3zNXzTM
8wuE6Yhsdj7AUkiULvSnamLSa/mnVfrIVDCyFEq0ZX+zeaH80sChmxhdd5BSxbQn
ylngXYVIeA4oGkkYy+wqy0A531EsEtgjoKoCbt14kco8zOuaGGA0gRVAHM8Uy1pq
AUnhFZ/hE9IDpDsaqD4snLyoYmvzLpy7CyYagbaIXZxG0zxsVXUOnwsxUtZDSzJf
BVl1weoCDORZbob2UJaYWdpZfJ+Z0AGwt5ewIw+pEwsOIR1fB915B/0fL0epApKN
nsLo9wZJu7wlzrHP5fKZwzaCXUiHiefoU70aiSXFnphumlm8uGPKvn8en8WrFSks
Kp53VWeVbcvImrHvEVAV7q9tKe7kLBxH1Ju/vtJbOW5PMNVwhIPOb7gY/L2Hayh8
ZDeaqu1X3bKdrZSUM6kUoSBTVwj3NrvqtKwAYc89Uz1uoyiRDKezqkQHUDPHx664
xXy6ykUW05irRcsHSUetAUBRB80GU2bmc/j+afYaY++rbhIUIvjqGQLeqn8KIDwv
JDiAap6R0f2VJo2MKEmwqf1q8q6qXapinwv7QP7bED2XvE6Yc9kb53EumrILVeUa
xYb770h3uulrKzzEdjPKtrw4w8N8rsgFm04BlatREqm3w4zHodjypEB4n1I7DMdn
8cKlVGAQEAb/7PEUwca/qaqE6Yr7ZbxRYpEKBi60LCk1fkwh3yz6y8Xo2sTQ+qwz
RkHaYFHiodeqKw0Mug/Enj/9cFb0w7iLVFODquRwYS4woJem02kv6kGjptB+OHLa
1SmcbGa8t0r4IZYq9iPQvTl+GENFOLvt65aTZDK3AxGuC4j5vA3Rlh1qkryUB+oS
7HmvBrIiPnqf7TvgcO5KfJg8e89QgtPdwzQIZjt+wxU8i0TDFm630Vl5CWBPZB1p
au2fOI82N4yM4kax6VW0Bj6kgy9NSY+HX5fbVkHLUtAEedA3MWMPCe85zYDcO576
bNQBAKNFZQEg0XmJAQKFXSkKAnKiZM+p3HEJORjP65zggolNE6baxZe09nzX5t9S
DUzY9VZYdbup+MfhGZtc0aHNsxNYh2qvaEL/dwJLEwNibSWnd1UyfRonCk+ZH84a
EP8mQebkMlYQQa+1WfeJHKrFe/Xu5Ksob8wSkt8HDWEUlHqx/D0mI1ejZEiLpw4Z
eAe4xaWeWLJFHg5dwlVWzEreR5drHCR2BN8YyQR1Bd796UGNSlYV8na2Udc+fcDt
q5EnZqEGucpCbJLpj4B4+WkvpfhQ9Ykr9sHHk+SX68Mm8Ur5N6rd3GsDr6+PybcN
FzBec4Hpmh1K+sG1G94aGRl8AYjBVOqcYXYMZUZ6CJ/3J3GWKjD8XtdHlrdEdVop
j0ge97tb+k2xOiC5YAPqNzGr49hA7K2s8RMCE+A/4qm5/+JTXm1g78mAyZxyW7gX
zeiADvisSK7JiLqYCZsWpI/nXHPMAHxO1OwEkGgg069Wo0O9yVWxwSERE/z3lWyE
vg4aL87ebWcPAL4RqZ0QDgfccvqlHRqFIfua/yKUp/RhjUOwfmIcD9ym5kKHman2
4XDOMIOpLiVjigk5jusFE8mKQq/N1QbbKaQGlUmKZJLX7/EB8de0AHbQwMHcFC+a
vST/IsRQ7XwGOxUIP/kZGr3jm87OywO5cjIEoQleyLJRJVZmhninoM+tPK5Fp1yP
JHJdF0X7ftgKfNV9mfItjvm9ZXgIB90rsB8gs7UqNtMRZFvRUUuPiPrS8Y3dXRG1
zsBeptAA4sJeuCoxsJ6JMgWJwkjMzGulv9zIG1J/C4z6L7Jei5FPvZleH3ggWRQ3
+AQlCZCWiWnRpwnLIVkH1D2pmsfQubpqMrahJtugOvmk8RZ70V2YEhAwfWwLVQZH
VJMLhUWVgHNaPajGcw+rAgXhE5Uqk/En5PO3lURKNJZRQMkWGhPnpaHBJL+Kslaf
XeCojoQO5fI5SMWZRzLfpcKlmFpueCKafbpqWuorwXSWjyNbxIUKeThZ5pSg52Xu
Mw+qDxEZ00m2myPLkmLkJb/UOAtpXRy1Sr5i9DOlAq99x3ICwaYvxBjKGVxN4VOX
Zj8/XKjzDGojueYCSZRro2Nf/9Zj+ku7UiH0wAAE8XCoVpVyAv61QwvxJ4a+6XAz
iaf/E0JCUpJTvEpzEmmoVdTZ1Z3kWH6zJKqicWK+t+YtkmHazUGsT01qkFxutMj0
rjZXFv+I3TL4UFCF5UmpHbyNNmjbF5FemKeVVXEjGZqYgP59Mqi2Cc/G1Ak047K6
GcCcUU+xP+1g10JhPHThjykZ9P/diHyC6AtjVcsHbz9COMirIVOztwmjyWIoksHG
9xwUuNvBmqUhou6ZrEGMZinlNEjanpZ5JFhooLaQB66sgYheXaN6JDE57uN3Bap7
XRLVLO5xwvpnF70bLsSFQr1KBGJZ0n/L8k6oZC0evYWKW20zKopQwsl1fLt1l0dv
igTAYpfD00SOaFGao2rfzsjFaH55vYOeFQYm7RWAPnto3xjMCCyzTteqbwH15uPP
afPSolH11pfOXXMINemogwTIM1MPJLfDmC1tobYWzFV4nBuZ6Pz5+9KZdxiAaK43
3Yut5FZdyhakJzTHSk5kZJBx5/35Ta+UHj/tE+C1NGEk+8rc4+mPCV7LTiQfFN56
YAXjaY55pNYT1TwnIgtd99bjVKJU5EFHNAeh15bQncgDQHmtbdgkzMAokTsRMLxn
A47XVytU/1JlRLLY/MpQXw+y7/IND8bicJR9a7atfKiPMMbzMe4ywOydoAUPQu9J
+pCoTMKGsbMgnIux8IW1K9YSASTjJWJiDx83BWuPXKVwkvWQzKEnSyEmyYxoTlXb
ZWVJXRMobBrjl975d0IvcBXx1vau4vLLWaDs1rG83qGoZlygHbjYeVTJ23C6dIsY
OMi+eJ3p9tf8dHDvi8UfXrpzwRFSU0PJUnm4JZmQiv8H6c7PiI2DvIqgJ8PXdRBz
j3wDo8jTC1KMSfDQ3SSBVH2HbhAHaO4iS3tyJ7Tph2v58F7WQyZni2mGe/zyFa4E
Xyb400GNWNiB1ieytZxhxFxOSGmAKxaERpYXKe52v4BBTaWutGwkwSEE2fRDIyuB
MD8idGweJ3wyWT5vT1JABSIKUZrqk1rrhIw6ft9ivwLmBb9+wc+hpH5EBZZj+gXr
t4h/yJ2STbSzwEHbr2iijPG4QY5EltTdMu6KkAhY/izYbTt2UM0HMoiQq8oP5N+t
Qs//IKcsQkSQu6Pi/rrAK12W0Yi0vbdp5mKvPzGxIoJ44dHu3b3QVnAPuA5sV2ag
Pa+rRZFLa2bz3u7bbt3/Z+/L8OFdJt7dQTcXUee36oM9G5pTZa3uaZLnRbLloX9l
Qd1A+wETlek2l4wUfEuJdEo9YwKQExUAmvCkx9h5WFSYRfNyDTBilh2TSUFZdiMs
E+wtJiWw7VUKCDC0HI4Yd6gHzdLqjlhzEL1ErfqBnggx8nGA1M/Sui6BZv2zV3+n
rcuUGoLAfdXSarP7Gxr5K/jR8I+WvCbOCDnFTpnVgdRpK5N41H3i5FAw47p87sGV
7+zDJry56PsvPrxP0yOJlH+QQ8n/aXBTWwMvP6fkfoh7Yr4gGS4oPxnHeKBFlLdz
Sp8m102iHbXzRuE1GD3x4PC/Gxa3gok/0CxGQ/xvalI3BtSfLcg8OgEftlBddeRc
uQ71o0Dg3r6DbDk7E9VwyR48nD9KIIHcLKiR5yxq3Z2R3/NVi385V9uXYYejYKAv
D1YJ6IF/OvbXGeFXOTWV3RCx43vMeBTKJdelo5AVWNUSxYH+5qLJI+ApPqs9Cy0p
WNpikBsc4Xcl7PhP16WZl8ZCdgjlvns35xwo0cBHtyKTj9QPaRwp2Ijbh6yIytg+
g6sPPLQMiedAITMNQhL2sJMSQv1RFcUBBYo8dfTkB8LAYtq0Adzs4eHQGa8H/u/E
cdpw4QXy2H+8AyfhN+qdXv6XPcoGC7bNO7JS06HqZOD8ROvcmanTzbkFWvbet0Is
hxdxncC/Y4SBVCBsaahAs/G6x3kiHWtCf54bd9ZJ3VeOeI8aPQ0CfZKcJY5aapyc
p8t+XKxBP1BqYLqP4UpAGbxL9OgjxfyCSj6QLgZ4PFvZ30hc/yPzUS0r7I0kW6sT
GfmhICKFz/czQ5vK74PkpXtquZhn+8xi67fcg0Gravq9prqoo45RqVThP0tgBKAn
6nBPTOCgd3ELjaGZ2pUue6LJG5VRCc6/jrO4B1T/42Ouw/4LOEEogvhZViVcnwNF
+KHeseW4pZoqvf0VRts5R1oK9V2GkqsqWFbVGaW/7nb4EPAsYdv4h4hiz4XZiY34
5LqemLfLe8VdLJEocAvTIf5GUYzf4kjmxtXjYEv2FsPJ8K4o7H2+MFkv3oX8NeRl
4czesgxfEjjQr56uoabO7eWci0g1IjVaabB1moU3YyuVKj7WCzVEJwcSqrFsVRy2
k/7DtEf7uKBHbsXpEXB2NjzeSsQ/QAv4UL9qXsyFgi5jDU/SZaZO5lvehjT5XOS2
HhpjfwattAHddpG4irpg8VpCUjZJVPrbM4ndyO25i0u1V2OyF5AMuzYdfMClu5Vm
TWPsymDLa3bBJBE32ASRQSSgvQVPBr6uBHT8+3PndzdQs4JQniN2em58oLWYZHfi
oCdMLy5S4EjgTw1dHgmzOuLDYJDLEZwFqGMW36lAeh+0wN3E5xSFh+I0bnPE5Ld3
bL1zZtBrMkDRRvutpgH+08lA4XZl4ZHVK+l9yQl6iWCeIpC/CN1nFYBCTaRmcO9L
oao/e6to9F5NznFwOYwnakQ0/seO15mlsQOrPaIvZ3hNiEkF3TS2XVpPvDAufJUb
DYCuQ03/8KXtjTlVs57+Fkf6b3DBw7jBgu0Tbrw6hwCij8MiTuyCFU0gNMT9jUGh
lF0Fx5rTCZyq40KvBPXMN+nLDrTuq2TDej144deEvjccw66GnoE1FoZppW5mwB2K
K6S3XMN9VhyZqzCDkH+sfFX3gbjZtVCnSjGWeOBsJMWrIMKZ1WjKH6TTVpSjDpPC
m4htm5cvRan09V2fWHJXaUWsueW9LKOmmfbCSkihA3zLR30sH1CtDUVibJcmr+GM
QZXllU0IWHn/Rhn+Qi8/oOG97pLy7j3wcdraTwmtN5iDVoHoemjukMKLswlP2jG9
5hqyuOAo8QhV630BJX/iHwQqJtXNPEhZFq5KLXJKF5URvJd2yQrQVYJVm+C4Omnu
GA97RfDWD8f6VnPQkcj+ow1fUuQEmoMy0V0mz0hcK8g2VfpSOuSmUHasMKcwcesG
gNSaW7sKADyqQqIQA/mTazmP8sYg4PEjgJW2I6Qo7qrEexe0ZeQkhPLaah0BD7eE
inSBwuLFF/fx5pQKt/xnUn63y3yTsRMOvTGKlxXZKVnu4gYmPecKEwPyq7iiNomW
4gYaN5lso7VnWD/caJqJ13Ju8LZBYYIwf16mhaKGBuFBK3BMlnithrDOMp9zrzyb
i/vVVTddRqkG/17lBBqOL9K3KKejadfdOPzn/wW/kLu2vGBzqeHaw3jZru4HrkgB
bN8HLq8CxpkUQoieKzVcQwu+RZnonErzBJOkw4XXnPR8Q8CXBieav0joZAqn65Kz
vWUoFNXqUskWJIPPCuDnl0gAqLGb1Q6zvXdJ5PoIhbLYtP++5xKL+dm5QLFhY6sl
yk7nEzsN+i09G2X/yC1j8rAn1WE2RFSR8ZTBmZUeF2RPdOcL6zxNsHrp1bCjnuHp
MD0PEvjCFyKMn37+7oe2x8NYvNQq239cThRjc7ik7QkuwULfhZSiD8SXbT+pOQZz
EHpCWnVrp1rLPI+bXAevnzp0EVWBpCWvZzWKeM5nz8leO2MYZf4Lz/4iouFPXUT7
IA83CNZHFXlMZIjE4XgOM2/JhS2J3GsVDgXksJwXcQEZMFY6sxpKZP0YPiyc8lB8
Gy/BoGP46MLWLBRhmf5WPoCNI4LxIcU1RKFX988oNGvWSqGI7+ZXMU/KMo++I7o6
gFhuwGk+ecBjfHSwzh3Bx6BmMURAORyymtH4m5zE+zYsp6drHhEMkPFWiiMYQMGE
oiKtmYipHfI9+YdrQ2OmhOWYg+B3QKebBNfq3R5z8dyKUeweCSwer37TRX9+KQ+K
yynFg/kNIv+IKusxFvcUFZ3ZZRoSKpWiRXahufbw6tAOvj87BYXTLRVE4SVxKNyM
qQ3DUdkrFG0Cs60/s2/EGP4vl2Ppzn+eLhzOO/tgjPOISB0SE0ucy+8mD8hlmqCk
HedgrH7eS2j53yI0UuKT6id3dxsC7WmfMrjQXJJCZhbVasKEnfRyzGFb325rwnBV
E7c4GzAaOUpebGBxyPXsni4Yy88afh8s+gi7NM+KBx67N1pOwrewFvYEXSua20wg
Do955Jv/IX2ND+PaWBxB/fnu6wYdQT0/GC9aqbErgjI8BtinUH4wB3k+ABz323Pr
fCvQDbE7A2HuflnuULD0Y5xEJeGSlgO1XtUPx9l/j77fkuFmhkRD/rEFLMtIH0E0
LnQmDKUxqTET6XfBmFKMtYwQwDcnDNHvfzR6CBE6eOnvJeQu3koz6BX0nE8PYM1j
OyDU+6Z6xt2D0Hlz+VTPVKbjLiWGCZnzjgamZ+EimStaPkh4zCeAQUbaALlYf6/d
rrSfutxnlwy5Mnrg4oRMZepbYxusa8CMFP/MMpAyDLO1fMggBWptHYjzh7hYHmm6
IHAfFZcffhPouOmYqiQMxgYbMBN5YjJ7qK6W43I/VgHctWAC33i/Nl1cVlasw3OK
depaWXgyHXWAhorIqFaqGngBhvk93odPHviVdrsfThW+PfrCUVh8teOqJ4AIvcZ8
3zRImzp4S+YyuTIgUx6FRNpF7XgOokIuVeindoEAj/K2oMK9Ny8BYBjo118rlsvh
1RFxxfLAfdtXcWo3RadyQzFoAbIaZJflQbjJ5FzJHq91nS+IEi+wVlThKTpdHBB4
r+rMZ7OZefsvja1rECdS0anjoLWrYRcgBCe/QFjg3wE9udUQahah3SH1SZ8CHy2R
Xwy5clyXMw46CUIuC4EEZWuPy+Ao2VuOJGS3Fi/8b9K2WsJuQeIqPy5EzF4qifKJ
pp4j5dtj1HdRUxrRRxSgTPLSCdcztyDxRa88XmZJnmbEYmO1WeF3KafvDUp29D2K
Xmis/nUPydaYiu8rs1QvOx4L8e0aZj9WNU5heoPc6P8oH9f8MYwaBz0ugOV+5jMB
Z1Lzd/KO22c7WE5tx3U6r7JyHDD5V/Fi5LGR8uONdZZsvKJSVyFHVJRUkMiXpMId
xpniyXAZdprXGZaHZG15ApOgrlDl6xzjDCS+8b3R/qI9DH6YKA8FHriG9SKXwPeA
rDRTeuQ/ENwXtnNinx8mTZfOugpRWchQ2j/k6LRiohuSB00AmeXSmo/X+642DmiJ
AcCMO3rO18h+fkayiCmOGlT1SdFMMDlf0KBeHoUn30EpcBCpBAKGQBLyhMbscOYK
Z1zNm2rF8lzoAjDqbA7gblmf6T2O0LiD+zRZ04EJsr6RSnr8y2U1qkqrYDpWiRMn
i7wCi+GjD+FgbJ4lZdfsOd/cnWapFQc6VwXRg1JpW0mDXuHlPCVsswOAiq/SWMTX
ID/JAdCq9G2KTAwo+rhoO/9nZ3zFqr19661ZJkiXHG4CaogfXSOkPyTTLjC/prjU
R5tWzll/8pggLA6XgvvBtSAeLo75O67zfjcMkk12kKhilPiERQtamh53zN3sr+Ki
HmFhx/9rSLwhenzHvCFRjAE/ouHw599cqb/4m+e60R5tgPWh4YL9xbghsRhPM4X2
4JFa7GdAPRwFbhdvlKq4Yn3hoZK3hpomUgeqWCh6QwhjvlI2mKynz3QT6xLxe6M5
F6EhgGtL/hCh2iuUGz3ZRf49zG7+zBFoDWypfgTBF3FN73bddv6BbK0VQjltNlSx
7Fn4sP5e+NZioZwEgwLGxq6hKzkkUdVec+VSVez7dSEjmk5YNQ9guZ9kn6riJdgC
ukY+BIL6S+MP39COurJCAEun4Pgg3XBACMVG0KWT5EtGlgiVPOyfELtmse8bA8mP
Kjgvwv8VU1XluvvOwO19RNIN2jsFkyo6DHk0Zr7phBY0kgMMs/cIHnhla1gN7U+5
L+m9sKdp1vxUurQv3obG90AH4Cvv9ZNrnoU9sBM1HeMV0V6Rr31iN3njg2VH2Z06
AcLcSjKh2v9+rdZP0NLl4Go29yrGC7Owgye6A+EHz3GduvQnPJznttxZA0WWC6Dq
g/yl6ZL8lo85mYjvl8snmUYb7muIs2Pe/OxBQpg8ibO0fipndInAA6qx4C2RSMqU
ZWbWMLhfuGgeGILAmWW3QWuZ8HX5hESYnKiqdn2+1JvDXCfdhzYAFEuV1KI0VxUG
qsza2tRbmw/jn3Qgi3Gpp19V3ckRyHYyxhEz7YAyOORnVORXIa9HXZMy/CxBHTia
VEeMtsO2biRRH6QoBVutn3SgvvZ+R2zoSMLrww0Z0usejXQQIoeUADKMvVSaIF5G
O3+dzx5+7X4JCmiq3OmrKQe9NQ+pz/Tyizog1yRu5ARRIZxOGSc9dc24RT75gW4B
YatshK+apffhRCia+LWNIJ13EzpIqC6bIF6qhGVEgvRqyz6o3/Z7TX4Wg8GNSNI6
+0qJH5XNvdSSH9gqE28lGHK5a3Fjgor3oPL4gihpJoiQ2DQ29wXqCaB2RNvS9D/t
mcVyzGlW4Kk8ppibdVP6mLHB2ZpspkV3H4oOMu48hnfy7KL3NaYjfklyGlIYbc4B
4c8aSc+76s7CuC4WznTj801b1SF7YsV1vSuUPWvqDCDicT5ztXB+bINe1mg3+JyB
FZ6gccIAlGqOy/GGkDE9DpLpoNtIvfd4c6WyEdxi5tb6AEdUcToXG1/VzyYu/Ryv
CNQHhUY6Xdw5Gaci3gBHGVuxe3w1VvEVGJoYHAxTNeKQtqL6t0FY6gueBA3QeGpf
H/SSedK0el/uo7YOyt14o21otuATLRgAHh2gPJVMJxD5vcWl0NptJ9d+WLMSFgav
NZohgR9sjasZf+vpp9S4tU95StRtPea6ym5h5wiCMBip/aWyKlPcvuRDE3vY7hor
WAOYyiHQsqxKKq2VujZb+D43qqS9HMvTykT+r+sdvNCRhMfo5kIT0KgrrUJ0U6CQ
ysi5WUivSlD5lO98gk9rH6uUTjWPpIoyLSTBlqJUD2SfLrZg82B6TSCUBUotkHc4
dOhDyNDqyF8vG1P3r0cBBiJ9ThHo6n7vvOORv/HW3gbsrLZ2lToe0Uq1f+qUBTLi
V5V4QCv+PK49D0bwVG+8RcA5P0c5Ldg8Em4yM3oyYD1WIvlGHwAZc3usDPnmnVc8
MH4jEaOddHBrJkftRSLWvSmMDFFF0NtjXf3MDJKXjzmC9/PYHUqEu7lSdfngiGuz
pY/KtAT8LmpexvfUwfubY/5rabEOYDEhtbqkLH/NLxHG+SkbVnny32SmOw4vDQRG
vV6trlJSy9pvCvj1qas1YWy2u68lf9PYoq4lE8tFHjnNmV90Mtv8CLtvsBNJjFoS
pZQHAwfCl6dOLtIjQ/orQV924ShZHLztlG3dJsqUvhRqNWfDy0lm1iDWysFkkGdi
Ijqs6oeUKtqfGYzj7ZciupqJ1qKzhJUDsrH5CZBqOvBFfbj50SOG14dz/9CaQdjk
YK9hGVj6pvW0oWNbo5iYr2//ydgmLCRtgnIR7LfieDyXa2FFE1BtJZAIaaipHdUY
7yXSXbQGYtwt1Xvwk7RQAto47y78NXwnUbjhb+ttO2FpX+LL669A/eGkJ+9Hnyb3
VyDe9+NYnmQgDbS7SHFltPV6AhHrB6gkEOw54pivCJqWGG7FMne0CasH8E9szg90
xv7BnnFzM4WfPFgT0v8Lwm3LmCfi6/HylOP0llPIoFT5DrAJWTZOpADcZUIyMQl4
avUcGb6ERRfIQNKus2tQM3b2jB1xNGtSGCRcv8baRRJkqQJFA7NdjWMT75lkDXwl
mwwga764e/U53GkyfqE5KTVKGbGQnsrQzPWzbR4MC4FqLDNbZq/kozQh8BPb1EQl
x6/Bw0JWBxqHoXDycdrOUrAn9VckX6dTcyV9XL79hgMzc0SPCnmHXcn5Tt+hVTfz
SyFnCxdjvB34Za2aCL11dFrDb0KcUYEpxbzolzwgAKpvWe9rxc3jH/NYzx4fckLW
d8FO9WMP2AYa1z2L3KcXByG1FCJfL6j2aYzlklIrr5+cfj+LyCxcG2nYAqGJYHVC
EdLKOZM+33MANCN2Q4sAA4Ti5ZhC6ChAwbQe132I6ytEVpb/3HWsDPKu68eeqknh
bXFJbNrH5WrAVuKjkcaBoV7MxtLeYxByXFGn3oHQkWXVzhyOfLWUXe8J8ASHqOhM
9aD0YeZFVKI1Dk6ZPxPWU5ZOeV28yb8wE6XPqxFPli6NSLtKLVQVMpZGA36pEl2C
1Bdr7X9T0TTUzfGBtKdQj/8pxMlMkkKyYNoIagC+HdstF5G7XzOu3cgRpdqPOjA2
ZA6QWvkCtOVzB4eEeAYF9JB9Bse2V12Y5dRP3fu4ODGAzCJPNVhDFCE4v3tXaDQP
dJSv0xsXT+vARtf6PNY4aBRPPyJuFPe41yBIulHtpaJCV/B58a1+FHQJ311BQ5ph
og6w+9Mjtg+IYAOIaWgkM67QAsKLEk7I4bnJ2BfHvSdsBn9OpF+sCn+fLqkBBrv3
mfUZmmPxxWQ65plP8BROORpoLE0489/9IKq1XPjtCpPRBU3ogj5jEuAp8BS7PrJo
KKNYZ1UFLMqwn5xhdrVRE8BDFeDUxXUvNEldOU07nI2JujmJzdI/LREiwmKJ6yBZ
0SNlUbW9yODYvZjJ537M80aNuEaJsBLCQiOtO03yo5fsUFbzIrT/07jEZpLe88ht
MlY04Prv4oHif0L3e/AGA3TsrmsIDwfVLX+85Pyd9xYg32hU2VpPkTEm7OrSpfD0
sfo0Ld0GIj5vaMoE57C+5T1uOb853u4prs+Aw2xZUu//nXlfMdFttjcaHpEm57YO
4CIHImt8GQsDoWJm+uUyUDDJ4RFHogU8Z+SXNUfgMtnI05giOiAxkxh0rHDD85Md
n/rhmTmD6hAcj6+R31Y35DsjBBn/g8cc2ZAqXLT13eYnfZ2+pdY/nOkGBuNKS1SK
r7ESgtZgQMcdu3Oa4YrJD6y/07FbddxsvONvyRF+YbWYPmRHYH860LLcPk9Mnssc
FdvCSMasW00oQc1vY+a2dFy6jshpVk9eLby77paVyF66iMk/iU/bC7O5uMCOYvDw
Igdbhb7I6iAHwhWSgHKnSmLGm0dq0kzaiA9kP8FLkn7P8Vxg4XVsH3GGf1lZf9ax
tC5pdGFD3eH0jcTEsjlHKGfBAe+65T1IX8VLgszXSDu8UfWEj6Doz7tQ9NUWaSCP
ahGjf5RurD8/BMga/EvoENDlllLAKPiR2X+KBohiVFjcqu2Qtcd2xhHrwIH1WXX+
CcH8K+Dg8kBwTJcG6JoAk7iOCV4Tw8UtNlq34gKGZA642IHkCRjRh2c28Eb2bUwS
bHoS2APh5cBiH6o53MCFMTngBSoWrJ4HRArnkwN875J7l484X5JZ1JIRJdspBe8+
v+iE5Sjcf9u1E6/vG3wl9ePqi7m3g7KM+E/OJiI7+/pQ8N3A+Sb0YmTfZJUJruaD
9pTBXH9FgsXAHaAmzEJXVkUzZPIBwzAvDiG/SMPRNiRNWSs8YiA/Fqf/v415EZ3i
loE/ymUs4Wfr44Bg9DVpl7PV7vmRRONKMbVtvBBLUM23YEI594ci6NYo3Uzv9AZ5
mijuNO4HPdq+hdJaFdHym88cfROeG/fgIBTg1qVBWhiw46VjwEUkcrfZBJkMPSC5
9F1ofzt2k5D4cBuQK6+vtX2CqZuE1K82jrde2cJ+AcQz6PmuAluMjvrkRumrNYeD
tbLUhryXfACR+2ArBAitHzRdoUfzP+GlpSU6nw5w5mTbr8gOgZ5Au5C36SLsATAu
buiVyOzcBQIJ0gn0NyeZc94r93s8vcwwq7WFUudHv6ZfbakG1pNysqkaKJmf1Tyr
Nna+4rIahWK6qFnu3tNdobXaTHdfPTtFvoMk7aNihJkWcTyJs7nu1V2ZdyPLW2Q5
OHRpQ/LEB8Px2qi6jLuQQk5ClaEsaJaMchf2XPF39tdBxG53G4PQ1ctpefCoUFn7
IphOZt5vZqD/j9zkOxm6fgclJpBwJlM9iptMr0iUlOOba/yiof5eItGE4PpM5+Zt
ckmDx4D55Ns/A0kmypGm5kKUXdQ5i2+W8xdOq+riNZalW+WYYkkcJghyGejp19Di
t7dUObKfld86lTfFeKHgVPXV7H2EHOSQygQxqZlnvy27NgWUJaa6jzGZVTK/yrD0
GqZcc5pAamr3ECrpVIh2UpE7/xTXanE9VkfzMt0z+2y3VnIbL9uSrjdX6gz89D4D
2KrvW1vXQ/saPIb94kowJGGD3OurxoqkHNNQqbXBs5prWWgEQ2qAXWeR9bEtxPMD
G1KWsszKHCekbzxg5Pt8902TeedeXKyhTt+q02SgavRabcFZAz5ZF27HwroC6AcE
L5KOtBHPm7ynIpzi/wFMsd0s3hxzTyk2arpKdVA70W/MM0+n1fY7OAkm1dX/5ICU
gq02k4SRYlu73gZ5G8sls0CllT4Dm7CXuIA3hy9fL2TxMO9XWhvNaDR7Z70d8A6X
5X56Taw9UfqdRjV6FqnjCc03fB0HpOxZzkTdIRcYKbiWSvESbFkyWfpFhvsBgjCk
uky6NvWyT45tgsZOxGU+m/jRg4ST6bPWeTm6xdXM/PExnUvDZUxzmVvCJexT4eOQ
/pQnqNYn4lLljSkpf4LGNL78lVt+HEj0mUwUeyP13E+f1cyYEYa85jktanmeZl0p
00x4eYiK7fiayXztZd/KoCCVq7jgKMXgHf1tAdFEhoBg2JpUiImvblmBExmmB6xt
c9Srq/U0jXnO3k6bAVAiEaNspAtDpEU6kLdN2hxKW/zRBFAS3jrhwIvZzRI8dBkX
9DHZRdXjCyhyWlnXGUxK14iier/YVqXjPEIV3niiKy6H+hgLR1xAfU0kHyiRUcWw
gd/k1eR+CNgVI/1ycHWmmZRumEcHKtjzQ9YcyKXVyUuKf10nOOyS6MZk7FQRoPZC
o15zxkWWZHRGHjwdNX/Qi35dtztjF2lBNXl1dkLxpnkJMO/zapG35vpNeFO21BHo
vsULdw9iJ2ns9mjOG2JO7rfIcLh+Eo+ThWzTOlZmxvzyD+kooDX+UlfVfoGMbJUD
/Xs1khOgpgdifZido41WGPw2LJrZ+vb43AeB6TNaYldSA/M8W1lhb5hVWP60ZLXJ
W3qcLIdCMOJCwW2M+Rw4oab2fRZpsayNxMgrLgBEH/jFwjWVkS19JxzjRyt4CDTh
kcMzpDWtHyBN6yfSt+j0jMI//u4KwolGt043/HQrmlSUw/pUWsNBiFOukvPD1FNe
jQ+ej1r0CE658NFb7NACSrvNFxW61jO+Kx+Dj43kBMvVekrLwjlVbg2wB0cUulL1
gh14QOQfmB+XOF2bEMqTvjh4WWMxOwbwNBvKTnNpKlWsS+5RrYjjRA3EP5oOIQ3X
1ORjremYj1e6fGvtN8hSxckesi82ICml+cbPaM67a4hIq1NhTqKNbFl6eFlgiIOe
bQJW+KgxYw1KoZUYr+yXpflwgu6/PdrNQYSJWlp3m5Alkb4yXqq8kjFdytOvsJ/N
3fx8sek6Aa4sOhUSQJZicaKOa8TuzF5JPV0WO6cACHEliN8htBWUaiO/r5xpXM26
aiR1UR5a9VPyxBXMQ3Py6Dv1s+PSJNMlM8DTliQwpMNmOF/XgIRTdhHn/Hko6+HB
nyPisJeUL/J36luibKhVH37SodttUFoVZmexU3j1U/ImlVi960gTFPgLCM4wMcvU
KAxnW2ctiIhGFXu3EcRcEqGDaVwNiQ9TdRIiZRy70IHNmQeYLL6bz2rWdWz+dP7V
MuZJnH6e8w2hjorj3xApGlz/SnxVEGJ2ES0MCtDlnoKlQupHqiXGKW1qTpO2c5fD
pS4CxYY18hYnlLVxOY6y2saTM9+nfNJXyGR4xaVRFhibHBeJCWT0eTkXaguU3HCU
B4SACirS1kDpniyWTgHOklEf1ekkmSpLcOeIkFAl2dfwDpyvCmgytn6YnYDSu//F
jPeu2V65eh8C84byGOWBtheTYBb+bjgbXVlT+gv2fl9VE+sibRg8SffqzqY9sbK6
gW7trGc9OGPCzAtAGhBq18oQmDr5+YuCCdekaGGoiQMw97+vmQXgjIEgZXXFzbGx
c0HJV8V2mspe33+DbiS1YeAiiydkx5Yi88wdS7zNkoLbfoPtiZvTfO7mHxCoCxZ/
B7+6t4wwwOkmWlvDPBGe5JZ1oc0iLE1ssPmGT0b2SmJ2Bi3cG7wigfUfdirLhfnx
NaudkSv6raA/Pggk5YrkXvuq+SRVZrdlXTGdI3CAagj5LOiNObGt3hjucBzs9BQ6
ZYCTLXytw7qtkTGnfnYkNdSRBARHz9piS+Hxr3gmyc0+bXY+f+RbK2BhmSfNQJNV
AyKy2KHb/9WZo4SJufpSetM183UoMUdYtWITBYVQm3HjLVJoWFRJLtYjretXUfqW
wozRRtW6SblkUDguaV1EjQEsvNJoFksQIb9zWmXqwSMHhjGiIU57MUmHqaKw5wnS
PZT/yHy1BR/X0WPMwf6HOSrpmyOCmgi42L4qmsA6YYx5mb3PCgsKwJOwbOUaP778
7HAOyVjF3EJMAcH12fJwJNYWJ4sq28QSi7YxCxJ7tuJ3L6uW9KT3GHl6fTPM1DIn
3dFflIE6beSHYCcu5Czgmzceqfzkv5LzsWGY1umQ5AFKXQGAR6TRdU6pNRHF0x+x
M75JB39Qzhq0vGoXASVlwFLJOls82f5DUZONM2tQUOTdaWz2WsYmC1Fp0ghucjD1
1gAIa2xyAybb0WZbgOYtMNSnn4DO0wQY450Ly66tAHbuPMF7/QhBbGq+dW3DJhSZ
rp5T8+TeZvper/PFTCI1veCJPoB3i30yqaxJKSBZnLC0Ss8uTQtGN5cYWy+Yi5L4
kWIF2siE3DlYESndekxPlnwclvC485V2b4UIEAyK+wA1bZgGwOPJhB29HJhsiy9c
1EZw5NO1/S86Pe0LgPI6jEUnrSFLKuwllRExNzXb7iiXBtZdC0jZ/xl12P6eTG82
EbmGp9vg4bV4zWq3QYq0c+V5saDMi8P7+oH5IdCOXDnUsSpow8JZiIOhYKHr/3G7
cYzyaP24rYyZsuUGxPyceUW/a05pVfD0S4+Cw9KbJlAZy5qD0TnNZGnNvPtpWmFb
PRqUB3ZHaQRLwT5gLfN3Uw4zsKUkZBmIxxGwLp0am4JDAabQAdSqKWDVjWRYBbKi
Vi+lM4i3aRh6WKJYD1YVjTAd/ufWSPpUmkFwJpIJPjI3FfvVp3+XU7LUmJ7e4mc8
XHHd3OMYugOHd1VmwJ9rLIFgzoWIuI1gkhHje5MXIqFltORj6nQ7HEr8in++uIad
qgelggGctW8J0bbSRUUDdXFQ3ZHIWVD6FdlByOY1PJTxb3b0IaVaVs/vSPxD+biT
jiP0UIChStGgeuXKe6DoC/wzeoY9axvYDnRt83slrgl+xZBM19DQ4ZDlGRn+0zmi
Y1qb4y8xz05VlUgLOZebfNE8VlfS/KYwAWw2cttEMou574k2pTyGN70V1plgSK/E
vfR1H/FPEMcibSQ+LQrLuxxt0dkLuwMtEw5ADxrDpjwjQItHDhWn1bJGLH170reU
hkh2ijnPiDWCHjVvEo+V7RKGeaYVuEnlWDiZRUIYO/Qjm7LR1oQwLHUqie78I4VK
yI2zHwUISOLxzHGzsW4dkwzvmal28lFKs+Qa0ofop7AZFam8IMfYQnXTKPeclu0d
aergUc4atjLu+jpQWRfQ8RdBButsrc/9NBugGr4/0r5zCZbvzGfahVOB/hEwk8Fj
o+q71zOGvAiIVEqdaW5+1e1Z26Zl3O+GWIWNIElC75KYp2q4WQGyjpNnBYzZvnyH
Exz9ac4b6BRO6INxdHSUyLQfO3rWbsOEahs2fTtbTBzt2FcgUrCrAxSxzRe41/uG
m0cY2ndHe3Jm0gor8ZTWMM4HP8KACUotCQNKIqbWeX+yX4O4XpHugEuEtvh6QpCL
HnalaZgBFPAN/laE1aFmyGKXHX236e0jK/IWYWNm66cXxPYgyH8ovpaCPBpz60MX
eyW548QyfyyiTp9w/va94tgLzNm9r+RUtYSOysKajFobHsLoE0WDRlpWlzSqmwvf
W/edAbxeU2Qm9YodtgCRNCTlpqHGvXtUlm+/doLmALdni+VvqM6OwhFbbj0wK6Ko
GyWCNnVOJ+2ATY4ZGeqlCiWSMNIu0iWFUBU+SlO7i3DC/27L4nPtM3qcaYFX3GUK
H8A54jpJBDlap+fzx21F0aJy3saDsIqGnBgeGaaODd1kjR3RJjFYud5qbnYDblG4
xBd2zjx4VuItUxnNHonMc34OanZ+RLxAeAd/6F/JEmM1Y//8SZeptcaw8FRZajjY
YJqYrKkdaSh/JMg7ZgYEBRvxRUZiuSDr0nsJj/ARfGiTL6F9rgH7I6hm2yn1K+CV
Dyxn592IhuJTwiM05btAiHPRMRuis5w2xgc8MUEAJDBOUXS1e+fjQux2W/TblI+K
TTkPB5Vl4jZdcZ0vvw/i8JGD4Lwzf84F5X+hU7YnuVEadVP7kTPRLmNLF4YdgQE9
jGAxLFrVbjIG1S1QlC4gUnBYMD/jmp9vgEPtiNLavoK6cGQCmEUzXs5AIoVyZGRu
ujA9OOLpwetKk2UinA3/7qXfpCMr8k0bpUfLQwiHvBAJzb/K5xwdqwXnWTA6CZp/
kiafhm/foIcRATig2GwKLmFgWB2oD7Mws4yP5j3+OzM5nOeAxyrMq/XT9thMP4BB
Vbpewk5gPuNG2AjLzOrayOfaOVZCB9EXX+PSSqD3tHQawfpdyIMLKgoROVnCtNjv
INdY8XAPG2rCzEHY8OZzhE/WrIbkhszQ7yovqHK5kK8YYp6k8u8orwzCSymvfVw/
PZ2E2EwihBkUFRFmpeIAxVl5FT7SMWefn/9CuveL98iYqRuKoyo5sHsCqZx43LcZ
ETNkeM3w9F7sfLNixExfV/wpzrHb2YElqE/Si0OzU7n1dLcj9p2aq0V4hhoBHtTI
dzosXAl583zBaGjD2azgBQCGBxuMqrFhMwzQMHDygHYA/m8+ZhOL8CrZCUWt/i/X
2vztTjQqgz62/pAaghwAVk8Q/oIfvY8MX6xvk8NWkrsZd19isRBF5Yv9lH18MVvL
6qWqFnPx39vkBMBvTF1FiZDR25GmT+b0fRmRrg5TqprYylXcsEGOky8q7cQBSrbm
r+08C0f38pEh4Jgtr9SYo+Mo1FWXCnQKn85+KKUS97ChavZ9LC8n/mRXWwx2n6fU
FBv7nq7dmEw1xnKaFcTmNZ81Dy8SozH/FTmXJkzTGb2/GOBIAZ13DHmsjhz4LTNS
eOrFhysF1cUWpuhEyk+OZ/weroy1hUlP0By6+D8skxvMVX5dssBWBJdk+JmU/w0i
BR0u4fDWQFH+Q9Fq/nmJyUOAkiVBIb5HgZ2do09Gm13lLaoQe3XLxZM6w3FdYptT
n8O6lrhMHc+FlBGHciDFFHQk/ylHaQTHECuE4t04zrJOzVQNe5Nl7/lLRzZdzy8D
CSGC7fx7BVTiTIGC2nd6yQOCeJHOqzNa/iIAM56KkdJE7OkpsLFOPvqx4WhlPcof
oSuwJJ0Q8tc6gF0ZwI5kjVAEyur8X116jDG//jzJANzUrwGcY5Y5jOyu6dPsL2Zh
nK5xDYMuaP97vquWKuhIHEZSXAiM3EvYJIKxMeKpyHiCgXq7KdJUlLX798Ig8E6N
84dBODIffgCnt8MyldhbR1vZGC+wPr8cHRIX8y7bmTqClE7I+nvxz/RKBxsDQOdE
tSs6bwVR7Mc3ot6mMJLzC/PBO08E39lIAvNDytYTKWYhVSo6zCJgivCbDypi8CzP
dLbSvjD977+FV9c8Agnp8QyZa7TM/puKzt/Hu46WzwOn9YZ5vc/+sM9OrJBW2iYX
TWyjepM1m6Wo4NgncYao+qynkP3j+73/mElpIEVCxEeVUxbmjgZbruGMOzsTtyEk
Pp028vZWbzo6n9+oi39qqDm8ste9FBpVpzlYDVC/DuJu9TQd9IWXZgbbn1wSgsJp
ARp8DerqvCUW2jjfMPVVCyhij5GWN2rgwzxh1hQuYMG1Fm3brSmF1NZNfUod+RQM
DPBDluT3eyCfEwpdNIn62NHt4hBcRoRAfe8VFOHzeKSutS14r/Lbk5Kq0+Ieok98
4SE0cBnYNrwHwKViip5/AGRs+HBcoFRT5qmm7rfAyqvlx/0YT025kJltuyEiOIr0
HC+F02nV/YZVTvvUjP2ZeTxeQdOsey6IAQ9RdL8EPwC2gwq3pXvJ85r+bzr2uxOT
QanoZGNO90LEwYrCtZO+WJWjhZjAGezCZ9tcQ3LEtlC8PelBlPOH620kqifqk5wX
wFaa+0UnyVnsmfrchVRf84Wi70dR7+bDH5J0tVnsGBvaEEUaOWwiAoz4Ozpa6CIL
EqfRqJf78wWBWsnhg7T/SAXodeQ8myIyV+erH6rluzxdcav9baF6Dlkj9dl7A/1x
gY6tm0PPZnkBwWrbuySXp1K/137m1eoDnOX6qZEljbvwCZMDt4aEkCgLm75GFR/S
LO4oYvPCM5ETLPKMbNj8lt01wPdcBz2iOaMXe9q56+A71FCzRDcWlWFxsDFspzQg
MUHst7HJBMYUW2TH9ZsXa3kw480H7MPON1lLwnoZw7sE80mGFCRfibQ2VLw87sml
LQi4m//lWbpJsz1uP/8zEHyMnVTFJJ89FH/GAdTFqHk3StgEjB2pHuimVo0kX5Xq
igtOkBOvxqi1uGzMy3kSIu6dUk3ZvrygTsIVPP7Fvq5e4AkILCnEt5m8eFKNcVhP
iReHaBauSMMvvrCrYa5Fmy7y631U2tLPrec7x5qtW9bse9YTg5SwvRaRYNKVHlCF
PJtcLG4ZbtoBs++N0Cwry8XbClm+aFXIwwHqSuv6uh9Sr/Rkus8RAzeoAuxMa89m
TAzxc8BDccz+GxSKHgJSndcJVm4E3chpZWzR6ckWALzlRBFd2hxk6pAM4JbIn5L+
BFYGaONdTYJ2OJChI3GHsZTGcbEdtSTp/Xh8q25y25tkfWea7BOvjYcykF/hObw4
OSlmQnDzMjMoMiwT1jfFmiDaAEWyo6aK7SHOp8HxEzomvTRjHnZMIkrx8S1JWWtL
BF1jrTpOiHBZlzazC1XqPO+dt1rRgkfJzviz1VJpVRvvutvLV9yHxgd/hUlTzmpf
K6X/yopNlXr4AB7u7WniNdl0+HYGEuCzqZVUVbFJuAHKaW4cEkd1H64Hv8tgo2H+
IBDuFhOe0ZMoEmtod1sVcKbRwYgpJm04heoaPFA+G9TWmdJMVGz9ktbR3xp4yjwM
d/emvkLEAeVX/hjRSj381v5ybNoDAgDkAqM5CZDxq8RoGBEL/Ir2kkaIazAgxIV/
07zTGMgHq9AT8uK5unvNreYONbYBU7g8v/H0hfFkzpQm1tRAX/CA3fXl2AVNDHIl
Aq6r+PSDzHXYqIKWoE8r6FhHqTe0EY4EqYowjo3Py21L8G4mXJMsYS0s2j/qJRt1
9gQduX5IbuftiZr+v43JLcMCc+b7LROVfU+XzjhfbP0BDRUYIh5tacKNKGNcdeOr
pK7hmjAmKM8fQc4VU+cpj4PFgszHVpNX1XlxeN43HCQyn/ODuo1IPXRzb4Z83BiA
Boiu4/4XsL0Zq408t8HSd3DJ9WMPlrOyAObGaByWqrUGVR4HHx9X7nb+ZQwudeXG
edFL5FhroowiTQctqUlVg2XLFgsvJZOzDw7JOMDUqe2lQ10jQEgtO3UYrBAdQXw7
4bhjUKfr/k64d9fzBcR+9gmUUnzt7InN8w35nYT66vabDURIRwn6XpGkczNrQ62V
H78J8Ly6LfRq6F/uAcbhDOdZcDjsFiBv1ljURb0ByU2TzLBxkSznGj1jnGlItYo/
VynCjkDWVw7f2ew0sxJVD2TsMcL7eBw67AvUZoUAa13E/GoMhluO1yHFjBJgJhYD
9ritFK3Ej/82SKZfA85EqpWbeuKL6zKkxpUipbKFF7NuXJTS8oImnqe+fB1cAkyh
fv8dfR8IAXf/JM0Jb8cnR8F43vGVNfmKc2e5FQrp1adptAHfw9hhlncATuwMsdhD
hIpUOc8r2sz1qdPzYa1FdXRwxfz+XRNFN16ysYyBaZr8gimjmz8gU2XycuiAfRUk
+B13w5orlEL2XujyTR86j8JeYHzS7mtSrWouKZoWtjOBLfi0aHolgQTxePYYkYJx
3M8CyzbkBVY5HH+emAUwuIgyUAFubjXpyqpfOB1/pCA6ppqgMwM3DLZB+/smm7a1
kc4RgNaBLMDy7S4hoCbrC4i9Qhi80fz+PorIKDFe/x12/l2wS+EWozZJVjqcmh6u
GuI65s+QwK1XKE/KyUqHfPpTuZj+5RzTlNAQzo+VQjSsAG3YVF7QjumYlvIjslEb
M8CkPy3vijRGU8dF3PdxIvtys1bnAXYX6YxRKKBzvlekvAiC0ndMNOiza5q7hkz1
MjB8H1ZUsA9cMFndIFx6LuFnQudGST8XtNnqkBImVO+JhEJcLZb5FpIyJLrKxXn8
KRibhwArQgrQ00IvkZCxnuowwxl5ZBwYlBnG2wpH2P1riWltErBsVeUBHrZQgfn4
ENnC0HkyBtamxN5ucijHXjfcgUUnawWF48FWFmt16UP5Eb9L+OJwsF8hl0kEk+0p
uXt2qm8EY752JQvllbHRiMtWaot4Ue0NuMZ7psAFxXrzBygN8nlGwsyeYmhj+sy1
jo10YY2gU0HDzffsX65D80I/5npdLkPjaKO3mIf5lR1pw6Y1Ex+lIp44j39QFkV6
3VpkqiOFS2tgfoFVUEXiajZojTQ+JNSPEe+j1RoCCXVdNtc0HkOBUJViMD5DO4en
uOqJaJ1TZOFiFnxKjbtTL9ZcaNaqYRGfC7s4GZJX/dFNdDabAZznE1/2TPNrqXaF
VxamD9O4xNumeYA4bkROgdZRB5z4uQlvd/GktxVcEtQxZZ2TfwqM0bZHDuoLNgiU
LiGb0kkb/ZVP9QBYDe8qBvU2s//l0adsskwgo57oiKEUqM7gSNiDLQfKt71zOXwH
IKanTCVAxuglG9MBX97Ea+LCsscdJThZWQ2fWF3VWdWDhL21+qzbr8jfFm8Na+JC
cFUhWBh4noUwiPZAmEx3JElMEYNPkuWVaHPAmsFK57EVns+lsvxJA+8+pbK/TIwj
AdeWgmwdOiqyRy840RKfhU94A9+8UUEcHhAhI/wWbsa+KwPA0aqCckiS+PQkXPD8
mKPtcKNFU6esH3vF+YtjTrqd/fFmzIdHUnd9MdEK68Pvt0BnvMA15dc/9XcuIGhJ
grCKnRt3CHt8x1/R0tMNP734vEDylydE7tDu3R2dvfFqsQZ7vM+CS2hIFaU7Wb/F
ojp8QeHvLR+7/XybZAsaCXp+BODOMFdecAzxFqVwbGz++lRhS+IiO7rl1N4gx1sT
hGeCiLrEsOyPBVUSnvLI97BdbgsgSW+7XAkUS3WsV5YKTefIm3irIVLlX+r8cD12
OGqrFgSC3Zn1lfqnqbq2cF85gHIC6VMTHOVBTn+oIOvGuVyLbnwNRchVfuuIp4UH
086r0BOX7j5cHjbkZ61HaltmZtBmk7uTKK3R5EF6T1opJxYus0uUBHMgCz/nKkDA
ESt/tNcs6Kb/0IPQQM+dbapPtqWmrgJzsmy+ToelIZ1xb8UUv3cCb4HgJPV2J6S6
PLUnP9mU1e0auLZxTpohwge0QVSItxVma/6dYAZ5ibASlpTd29EKMiS4HvDLsVfm
yeNib1g6443uN2VVlfO1vwLOYkjU/5y+EBhtBL8jj1p8PoN2HD8e+dV3pK/bk9i+
lfGH6Z6mJ3F2oC/Sgh25XJCppGRQBoVkTUt4QWxwpFHxqPEt3miMmyCtG2G3b6he
K6ZFHOmGfn9MaFQIyvJvLFwxgLjECKQfbpNbm32+V0rg1EH5J8mPHnDsB2ND+JvS
XTob2BOzNvc305dyiaSvl45VeSDB6qx5m0kHM25nNGveLNjRXi3UK7HaqlNeehfP
9IwBg6J9U4oHRKEBNnIfx40c1AYcBpRtSpKbLlSgYzOTuo65SsdKQVyTpt/jXcyR
UxLhBnFFc3eD330Cg3uNUXkHL/5kqvsbEmIfKKi1MN6NlHXW4JJyIvAqv/tXMoFL
OpQvVGE7rLwpwAlCuPWHN5feaFiUtzvGt820qG6XiemhrcYSRQuI4fqa85schCxV
AY0gIF/Dlfy3v6tyGBslzxIobvpd7CR/Jk/LDwmLoa9y9PDTHSZhekM/SF4nHODs
oLTFBf0LgtwC1fYoyb0EiyRhfG3wLrMr81wLs6OfwqCyh3Qs6BSK4OxkzjDzsdLq
uwx/ZXWzcQZtaQZfr0MFKFnrDv1cEnfknKxV62XPG4hiF9CYt6PK0LsU2OHFVUKE
xNGLHnZxQEEgdRFt+bYEb8+tNEYIW/WUwD+WhnpaGVouN2k+d+OUNw8QNP4WmBSF
npPhjSNCMfoAi0LpGIQBSE2Bm2BtaPixxhpcRMlRREPS9BKG2oFRNzQ8goQxhr77
zwGvpucT1St1FTLNmJvprh39N5wxdmAVcFfE0xRM3tdjtbUhG8ms4gEB/RM5qtUG
PdnHhesX/Hyqbz8C7K/vvtO1suy3fY2OPJyQUA221L+0X3KxlvzHJ+Fa9flaSQCg
hDHGO8ACjE2hkxGOS8opP1NPjPa+pTKGsPAFADX4+SNcp0Fm2yd5hWRWA5zUyrTt
Gi5ML0Ctu2T/9gtc0nZfyee5PL2h04IvEi5Y0T8NdekVMnl6ppYymPyoinZ/O7aE
Ba9spuFrEYmZfxGlocuSlIqUgyNW3pGi7dU38UTr8Rrjhqat1BVJtGbkxeEi65Ch
O17huOiTJfez6upye4mXuXPxvJH0kZwRtoHNSvsiq8Zdb6C398cbJ5xb2z+Oar5X
5wuIqZ/vESmqi+x6Ugj9m3hOL+Y31ZKj0c0SQ8MwjOfNTuXGf0ZK5mfuK8tJLMgB
cnraqnMAwbobY74g1gbe8ZTTz9DDDBRyZ4j4G0gtUmGsYXfIk3/tFkcsncTIRdmZ
3zGEPRpYSrCrKBpm8bSOImrPabNNCqckTkZXLS7wgcfQEha+mrai0c1zZt/8Pml2
O5lDsU7PDqlcfRZbR49Y6LJYBojfCEd2l6JV0Tnjh/VhT/OkfRDd3nzD+5D5luS8
SHMkKS9WyfwcD8lRbhktDBW2vpFAOQu9Rmw8jbJkwpbEInQpLNYHixYePoH4c4cz
LIQ5xucY0DBWgDE2rOQ1t82FxczG1luBk6SGMdxxrhLk5GRTLWY71KTHs9rEU+57
fSIC+EgqRuLRp9tcg74MCrYWrEDvDFn20/yr7ZyBhat9JISfA8ysrwcmgB/AL/A6
Nu8Wiqnq/jSH7JrhBAZ3ws0ceFsKan8oyfZjSi/188Tw83tM2lUKDbjk8uDEneOU
XFRvXLhQlsetUX3XZlrIpzqWn052HmAXRR2eXPMS0T5uIHTwzQMoWExVZgqF7qNz
kDgmuDnZcL6S2Lx9G1WJyn/KjNqSfhR7r6Pi8whhio3L3Uh1lFnZ1ClHRqx9tGky
fdodAbW3wPOKpiwnhpW8gcTyPFD6XqghcO5VM/aMnd3TPHMpArtsUrjq+jGFQGpQ
9UnyKDTFn6bN0n17eFx9ndhCA612Mp1m9aqskFk8lESz+kH7/QVz4mnWWJNzMj8o
oNjljkPehTTjWVjIS6bLJYCmHmHuw7SDk5Un1TDAs3i3G/ye0juPpyIHnSysD48j
/NEVDaPQyukdi1ptzfD9QPgnAq6wm8Bg4HNpVrooioLC/yzQUAyzx638MX5ry0ii
LwedInZdv8oT8HSFJUsMAbplmeC1cPK4Ep1X5dMqNt+ljkHR5brRdheuuxhN+py2
re5yasOHbdEvmZZ6ranzLuTGXENgCyY4j8rkRgENRRyBm4jsf3qDO8ukYIGqAd7a
CJYtRTzzwIXogmhrnRNKyzitHytRb1WT4Iykcq23sdRSjO0g2KXG0sGyQhySQ/Wt
clwXdAEsIFYYGxrMgqnHTgSuN+fZUXAUrj5t3nyEZi8BbSsBYr26I8/XLuvg6NiW
LVHm3aNrucL4I0S4Pmtw+cQa1ifyYe2IvKtfnayGZ6zYPmFPW5FlHgiC9bx8BzNB
xUJ9Vl1wgezEY8mSasULIC1On1G4OAyki9utIhj2adBRRt+uWOqZfEBgfv/SPm+Z
UZdMvxh1ZA3fJEIWrabx5b9w/+yf1hXnLriKvnC4xf4zU0ls/CAo6D/ah6Bym/HO
Tk4Ua8NLBggLE0fKcQVp6YXBIJ87X8JKq2y0Wc2mPYZrYPOuTa9ZlEW2vdggBJOb
RFMQKjBZR2DzfAvjLGylTuyxFyxfB/xqeti7pNt6BU9wpvX8rvhvLz6DSr80Kvvn
tKPfFoPYEVFXi5Bv3Ma2otfM6dipuGSrsa3ahO34M0dFxiLSJKPn6LONSUK767r4
1yHvyS47JFOiT8+I+M4MVQGxlfKqzQWKOzMm0puiQaVsTX+fSLLXgCC6CnoVwTHT
VQhhveBiBT/yRKmvll7uuCxKj1S1ybWwgqQX4IdGd1/tTCeHLegx2GIZ9keWY7PC
5Jgs6D70oi8V4+/Gl/PJeBU6bUVNG3y1wGrGns1MWMjuyvnT/QaK7X9SvzxfDQwO
PV9KQDpxqehx3hjnZi3cvlmIG7MEdu9PFP98MQ/0K/7T3ElwPjanMbjfGBxKHHvp
+01pBzMqzhltY81jdtCNq6oLMwVnfSDYXUR4+cgixY8eewWf/7Cfsj+Zd89vKgaG
a9nuZ1leeZbD3DLlCiJn4KKK2LLPChiGf8e++QaeNHcesy53a81OkujmtX9EVXq9
Q/bWIziMZatX6PPaMNuJv/vQxs2Jw+cGWo1KziGNEbFvkPr5yUQq1FDwZL9jEfmP
gRqS/e2m1RifzHumBscZhxKdWeBRYmMGnjES8twvajmBAeLkMrA9OeBsGlRmiNug
2KhO0B8kjEfTQhVQDXqD18WEO41wwgwH/bc1WvMwjyH/ZZy5q85zbYmVf1DMDqJ6
Aan0qmt+M6/vq3iB70Zf4I6BDtnjNX3AO/ykcxs0JYw0sH7a+C7KYm5Ekwtrqc1b
dmHV+4wYoQVjBc3wPnEnYO5/Q3FsPVDD1Bq2NMMwi/Zl76bCSAfrjN46EmeBjPy+
eD9DJlgmM5KwXD/x7DFbNG/Iik8I8kwLYvgYVsep7adVGo/GvSxBe4mmaRo4WKnQ
84WSxdYo5WEmLPUCWaT0zuGR+AOyCgAdlx4U+GR4HGZrexH0zvNTeOsfkFPt2xJi
GSWQsqKQTflmCZEFUPejo8ts5ySuepRG9y1eW+sBKqIH2RNpwKITbGIH6EBlQOKa
jdMXvaPh/hnU3CIjdyNqJUf9iKCdnEMKJAs3mwI5bPDAyEnT0UMcAKTBbXmfDoNK
SHnR5qsEIRe9/hr5K7hZzL8kucPlCFaPLMfD5XaEYyEL7VagqWEwlPr45Hm/nNxr
yCOAGrXpRf6u9Cg2xI+FjhuSZolAyrNlI6FXVBACytP9yUjAI2XXwSouSgtwgPAF
VNyOkFHugW/9NM6o9O2YbIZFwCxnBG0qy+H2opoPyE4NusFjWneTSzVAknVyWk3J
7QbDuOO7v3/doQmR5lqgiGtM2u29A9uU13PHU+KHsG8ZNHcrYNq9IHSs5q5OzrYw
+Jm7bkhzX6tKbe6NODkvMzyI/FkEP7ytlARvDS9BHgERgylk3FkOAQrw/KIqRbSS
30ePuqIdQwof4NfuHJX82Uk8Tbmvr/0AO6030QF1uKQDMGT0UhJEzL18TfUWWtnW
tvtXlDf0v0wJZi7fh+GihMImdKZxUIRMKtfBEookC/yjOCoACpvG591AEGtRV1Rl
wa+imcDF/nPj8BJyZgCjwnIhnEMbofhP6k2Rq13jyPIzHJutBtwfQ9y8YKcYMzYQ
55698rTHI/UO5T6bwPd3jjn2DhK9zJGWBsbnTLq0xBZAusIiivIVqVLElxth6rcd
kdoY74uKdXqkSXMoFk65bPGjzeFSq0nXdltCeWCGFWVhz7fPyhwXTkyTeO5OqHHe
oJ3efFZaK/Dg2DbDyOlbB6UmeV53SMQAS4B5oB+LMakQ8856ple7msPdQgsFDJgA
2ehej1baF4Ar2jwhQwNFGClkBEsbwqtRRC7gl1ka7KjARYGRMqOyqi8TLeap+cqc
0GandrESdfmsLX/1+D4omW4NlWiDXP7ESir5A/BGWjzuBLFZKxTz3zMG6VJP1UA/
uivR0ffzfeiMQEpj7cXh067navqnEW2A2GMPZ1IcjCyWVe0/C2mlmNOGYo25IHjj
pjc2sHPoIsCXlFvOfvH0r6n0MDFnTfLozZAJ5YZiYu2lJPJpmo5l4MzVcyRJwJG/
I9R3SaBn9T/Qhjnc3oF/KYnDFd7vN37DBX0hBR2hP36vXJgss+mUYwofcJ6phXOn
+m78pubjWnrTHSqXgpVX4j8nVDr0hFflTXsgK9Eo0SFzR5gNz4Z/iirDm8ECicDt
oUUuSUmkwGSwR6hFi0ABZ2LqLeMt7duQiy1ePfKDOtcL83/RwJmftrHnqB59Jm/6
lK7yl/6cfXROhTert297JvvHpr9geLVIbgkPwNf3ZiMlrc4/X/YGMDCHME9Orgoq
VJ7A7dswNyWaHnI8MpWYZp7GO7nSkEqOWsrm8fh8gmKardswDEODP9jAZ8J4H87K
1MtBLZDt5I3Y9JquHzIO2yQANIAPNKVIkJMbgLPKVj/LFRY5UnH/O8QyXkXQYKVl
ZLGZfkXRHXjZgYrpuEMzImTfFgNRxrr5NCaxAVS5GIHtXQr+dC11AsYhr559kuPz
SF00F+K/xeHmRtwG8JKpqfpaPHK2fakTuwMdWLtTcAWW39n98XIixL8X/hCmoHnX
PrvY4AjmlcyOLyHB8U6FUdk2plEVBq6p8mkcgcZEvq7vj/k+YLlXG8FlL70OYNKP
ja1Yl803uSGRGtFPYRfbekZIIAcgMhqyVjoT0TF0pM69P1I7n+M5gzT0JTf262L3
ovyWEaxVuu8yBqr3iIgHUuay1gJ59JfuBbSNgAqKYxyBIzjRrUBjJKmiLUg8K2gE
nYCHpHFyk1QPHcJ42olG/MklUlz6FeqhZwT655zBJ03s0tuH+tHRIrNTT9NK3Xld
a4zplshve8KT6OHhfhyEGKqrvy2sWMP2G6cIgEbgI1xPN2r1PgVxizPTUp6mjESR
4xJWEKk0XhSzTfs3F9KAo6hxCgtUf3lO8qC7KkX5oELLqI06eCNylldYZBSud1z6
/jvpR89rRAlh/LFaMVPcfDY9UrIsaMT63ijch5dbMSzGtTSJPdr5SpDxRbpRk1oU
g6ow+HCUHkRFSw8TvmqF1f4Dg8Gjj65vzUKG0se1w2C+0TnH0qpzq1mkS5jUQCRx
6PNG7bkkZ+1gEZnYnPhA7Rr2k7X/VNYSrs14kEsAAt4YzRinb75qxBjN7m4Dyq9o
EhNVt/W+vbgtXp+tDzF6fliu3od0p7nMumjdIizLle5lcfL8AVmS+fHO38aN6z2L
rBuFDex+7DGGW3jrtlr2nSMW+S+Yes5ermm2mulPxmhYJmzuNpLjJOkx8k2DsXMI
ocYC9t/XIiO5LPnUQVVC/XYS6fYA/sVX0+schtHkI/PzrnIFza9OBf8UNZjMYK+2
ZBgU+7oCR/SfejZZxAeJ0KL8DF6dstQgEWCZyo3ebeT9DFAV1X9sOtD+BrTur3CF
ncO55aYNkSfMI1H3lDpOEqMMy7bysLNdesrFehgHRniqMr+eqiN1grud6r/Ykzoi
k0Lpum0KGPEGB7gw4jnFU1+29WPwyPQHUJz2AcLpz3rCQDEEn6uNZ2x4Oj3zgEGF
0PNgXFmW9kQBLI3YWgT8MtoRTxEnOvFfjSFtU4k662mFBnnGItSaE+8hTZwZ+bDk
WuOZw6CNNrFt0X00Phu7Gxtea+WsyfYEy2JlG/gBweC9Fp820z+p4RK+0XedMbE4
RWScOl6ScqRh14apCK56N5lMDD3MyzQZSqmgtmi2u+gLV65YeqzW67X/O6NfPKUE
Tofs0gkHfY9kN0E5jOF9FXoSx8lPVMh+JflaLQlGQJlPTuxBtiqSJ9K8wsEOyEXi
AbZAN2xLKuavcuolFSrDu2Nc13woF/soHbwAGCa1GNYrcmm5KujxbzUC0Z8cUnMh
Wb39DCIwL3mbkvT+NeiazpmitzVmk8jGW+s/5Q7XQEENdmMCho6gkHZy8NtXL+Ca
ok1cNPktHoWZCWQIqSMMpsODUUB0P2m3Ttjtya5vrxnLnJVy+MUsfl3e2liRRSOR
XQBpbXKQEe+xGDXajP4iSE+lNpNyEDAnH2DkxCZ7fr8VYs0ILCXjGWyR4dS5Yp0U
9TexlmY9PoHhDDKQCFfssb6rnhej2ztWAgnFdayAnl1Eq2kl9yM0b65Y6F76BfYp
MJV0LBJm5ZuqAzv6qk5ZxH9rPpmqKAG1vgGr05sC8ucaRkCz8p7384bEEzdfSXZx
nw8rPNptJnb9P0pdYMUq/SZEPOOprbhYqExKpYiRE6kyj2b1kSwM2jVjpd+Jl+OR
QWZwhHGCVN49oQ2pEX4EfQV4L4/qvprvofFH/Pcgt8VeP1IvWPJFUShGV+4f0tL7
PUPfN5ZmB6wcGGfU34R83/uXIBk05C8auUM7xR8fMqU2I3bB3VSiY5D7cA9z7xEM
f+OzZI4d3yvO8SGGcNqDmHVUbe9CCAU6b7953nXj7C8CwRwdIs7ErYeHks/3wFb8
Csx4fLPAAlJp9Vulbj1jLRhiHkVK52HsvdAJ1di9D58jW2VfhdzYTJqXJni51Dll
azoJ1DDeupTVWL6XYXiVTbbiQrHSu76dXXoJIzWRt+vES3Fsnq8nEkXBuYKntrjS
G4SvN5Uwo9RKQ3ymAZuLW76egsvzisna2vrPLxltx/YO7L2VSi4JR9Edi97scAEK
bZvzu1PWg0Pmd+ZW5zyNxUgX9MF1cCSmCPYRKypOIjum05NZXa4ZV8uej3ifjCGX
aiUSSBLEctYj3Ler6/87cUaSwuc85IMoirZu056LJtbqfmgNj46FX6BAF4hf3YYz
hgWt/vjshX5FzqQa6k1Evm1dx2ByqIRSD292SEZbLlZKhXt/8WOcjlFu7mY4bkYJ
w9sRG2VLfm1VdQy+/0s+lrqnAs5HhOgQFt6cPohiOK7S1QO1rvqMWTR4XDh22Ydc
yjr+e7s18NkgfCRaqbfAD2wfwVBN7GvkvFhRmwLgPfFFu++pCQjxS0FNi0oQHWPe
C2LQaBIW4FKG/k+XSiYpNIg8K8q+nWg8PnYB/6GpiZ/pTUd5p3+M1gHDnCPLalew
Fm7rccyb4g4BrJnUM18iWq/odvEaGHMlWkBxE8AIuefKtOuBe6/EXiUC23NK65nl
bmIoYZYljXc5MGwO29spabbqmy+me1cDdd8OG7w7SZPJ479ooZ6zNi8Uyi8TU8LM
YZNpdyWb0vjWgA5HOXcuXBkfB7AJ7BFZGyJtMolcMALRy9WK6SRgCGJr76mzWtct
dgr1kUycX0oE+seda2StdgHT9cf1wZ3gVpEOouNMLkhjGr0sAvAt08DjlKImYxuG
iCGYIxtbWXp0TOmTipWbvPL1pBwzKdZTmU+DXQwOti7J25NHemvZRBwu1Hvn4zbJ
j7mFpUQW8jIhBQrFPQkDdTfLe764PvOWkTEggA1/C1MPaJXMmf+2omKhskfEiqmp
rCMlr9/tLsANK0hOLhqWws4hdtR1waoH8p1aNqu79fPyuuYeAJ2/TIPl6r7kmA7V
zfmTOotdnDRzYDyYJAdj4Jvp0iBwhRhVbCcXvRPlaG9REk0M8bSiWgteXagdP7i+
z9GEbZcd4FfvOChxXVtD+2Lmhze6lmh896MVT9XNRQVSFMRvT/uDB8j/noScW4t8
y4pLVdWkR15zEB7iGRZbUS2diY2UneGwLOstQ5gQsN5jzaZYzdQUiP7pTM5Zk5Nl
PQOTaRmrfc48NwZ8NyQ8058fomIeAjf7uHQNrsGh9MoQyj41SkHFt3gloMegYhN+
efbMdUKVXpklJx2buintiDzKnMN4Q18r5WmtYpuE4uzwM4zYKvWrjE5O7srn2zLh
v3gDUbflITOe3KqeBBgGsT9HlmzQdqBT0eE607Zc92HPXJcvr3udw3Xwj90o2t2/
GxJafudNMTEU2njXGCCqNkSI+llSqaeFv8jCGOvEclnR5Y2zQfhIqNRsi7Wx9W2x
CfM+6CzJjMR2OP24mRbAWjOM15drdE52LzZN4pysdew+T8b42qfRQWTmigu1z19U
ti4MV2XBtgLzNjn/yerKix+Ve0csgfdDarj4rY8M0DYXHG10q4I6CJ63g5Xu7SHD
2ZPsFK1YKeLjyb+u2DNCBD3h1B5YzA47+av9Shwb1s5+LW9ZpTpCM+XZkHZTi1+3
GclosyTFZs0skXdYs01WFhTvwVjLNzY1+pGRjxI7k5bAkWjn8+btDH+pqRug/azp
9xj6amkLNFxMKpYprTCZZ/WbQhA6M83nv3wF/THSaki/jT8MAutUU9TSNF2iawg7
ArSSidBNdXSpLleYmus/YvM/F9IO5FUygCevMuNcKBfh6NAYEdArnubVfgG7wteK
9p9S80iLKP0h2rXUVBxaJypzhjfIEr+NR5jn7N1EwMWFccx4NV+1pkdRJN+1EXu/
FUPXdWEz11wOJqiQwABC1CHGSOH6yfH7SOdDpxjarStfQ1rIIzIXlQ4HBWP0ybh8
NFSXQjW6hTpSoxWqdEZwU375atnPm2RiaX8HEVkjBeTu9IXenF8wqDgM2txLbo9o
xJ0SPx2MGCyxIvEL4SDCSv7Vpd0Q+3VYFe6X1SWgUixaDB11sEaSM2EqY0BSRs0Z
LcGZUDQ1C050gJ5Tyjkc2Gb9qrGJmEv1wB7r4/3czi3uEHJbeK7VwPfm6L1srkaM
X8QXTI88mIKNRLzqFY86YG3yfBL64ejb2+ff/et32g8e2Z+cAQw7HhK8N2XvKVax
7ncFEA49Nt/N9LHd4AfVg4IVJ6GcnOnlyhkKCgTKDesZ/vp29NouYR5K8x5+CJrZ
ZFTY/MKdAaHoFTLKQA9YBn0ugfF+rqa0sx6VPgfclCd9UnRmsgFzjuLToXCwq0bd
O4G82aEFIPO/CAR1nSl2q4OZuAEXt+9StvWqxovcNjckvW0PS6CdtS5w/77kWpYd
5YJaTVrOrnU6HMFs215/KRvHFB4p9TZb8ddgvgKqvcXbtz8s9kFEh3mGFjhCfM4k
iL5xeqzkms6VMJiEHNQyzJ8DPs87nyjd3GJfLkTNV3Np1jMnxPOk1Z1wwUXjXqXx
H2NJZc07kmM067ida9G46juJ+VQyBCrI8In1kRzmGX8v0u6kg/yy/jySDUp/mWrS
nG7fmlh13QSn8Fj08kMl020P+s78utVqHKcgDBCi6ZNCwV7k0mXpp++6k9dU4Ig9
G1dLJ8EDyjxhfv50wRQOVHd/wND+rsHdDfVhBpe4brGLmkOfsrpAUbKuO1UVR+np
aJ27PCdOCPd4G5IXIaRuY24NUhogK3i8JKt/8sx6l1+wXxOJJJb6zvWEN4/9AiyO
Xan1jPzHvJkNkENuZ/Y4mC3GHQVNCm6huEO6BvVtafuF7wIa+IGLXKF2O/KvdJxo
rEu5jXrMBYOMd2NJ1ePeOdYB+pnicUg2CMlBvtU+rkiWoJpYxkixdhV+C7m/gein
MAi4AA1leHixGedp9MPUcxcCKEXrWFL2vA+T9mWNYie9oDbXBSsursjZFY2Z3rvh
ULC1QFdXShUTk0WYkETiKCGL74rd/JnxFMvNxmH5y+X5gqRM3rLWDQ9MxY8N0U59
4LxGzspod/nvTjhXxbHTf7S3wu98ful1VnSpaljQFST3Xa0O4jTpESm8qaczttfo
4dddorgzcsSlulkfvUaNYGYRDGbeqIJP9ESmvep8hw1rNfCsXW67jbyjGEGcIkWU
N+dAUwpoNe8yqH0F/05hyQBggGRGgtJifqLJb2PV36q40jT5kjcJU3mfQFFwjGYT
g9qVNYEadxgGWEg86OgxIrUhs0qaUhWddjKtr4xN9pOWsCVLjvmQFNWPga8b2q6V
pqiEk3xaAm0FP37RVVNoG5Z4ces/g0QQf2h7Y6b+/tPVJUdgImz1Ln+hpbzktm6O
9wkiMWbTVuxXg3kPYq955DXv3T3fIQ0pARtK2N7+gb1lyA2/HZDnvEhR1jRsnjuu
eshA57wbZRFw4i4L5ovV77Rbl/KPhQQzVWiXZScHrqbukaDfBP7VUpxqw92rd/1+
5wUEfMjI8BoaCdrdGQ0AHp/JbT6x8IlY1nwtqUWlCDkEuKx8XhTjaA1mH9zLyfFP
eFEJVmf+SfC1Hcu8m/skGNmdscK3sUsfNKZOnzGJ7EzntT3+GxpX5x8s8NWbhex+
zQVmgnzhuoM68sVsWUoPiU5v4pRSJLrrgkAy2bBC5bRpKx5erbDIsLtFZGrfPyaz
QB7w0qapkFrDg/u2vVkA0InSNbvUonQxRb4E5RewtpUX4T/ROnY45F0fRHnWRYgc
d4HfT28ljH2535857xxR67KhocAM8M99lc5Yf14Vv24jG8u5W9FOmMWg/y0KW6Sy
aoHiplprYmIqRcStIszSJ2Rg7iOyl1YCQ35UYykL/rOEKypdFUSpN8rwVLr6bTMq
GOY8QAs5Y5Hert5v2D1TdkAYjuCxP0dWfDcLmXj8H2ly0TyT8+liAGY/xUWIWKdX
aITCrbfNd/rD8acTWjBVsyv8qusQ/GW+YMoQSTTsfqsttxAzGGmS6kIn4e9ivIFU
peI+g8Hnumv2PVr8jzwZfMai27eQJ+NodjOkrzCeaQjHH65aSYWiDfcg90pwrbOl
YiHP2QzU8Xk81gyPq/D3oiLRRuuti15zip78nWn0XZA74is6c0tZw9RWPxF0YKOW
fhoOn5I/5coAGE3MU7ko9baEfwILQpX0FZg90ATtwgAvKW7Pag0e1Y7qtNkZRDGn
++uf6O6bYJYMsc/W+vR8vFEFHJo198cWKSGLTeTod52Br0u8sWoBu+P582DSX+66
pf7KuwkaXOt6UYaZoItfXIBsrQfL3a9kwU86P9xyxayE2Ftv7JFtezavuvWJEkHu
PdcEefsZ5nYiis3paP0+8yK0GLfUNtKB201RsyQ+E8GGE48QTQZRYmjWAHxUWUkM
reWNfLirtT5MZ82YMGr4a02knOkR1Qzc9MPDzDnwxIBZVgbL0ThUksYHQW3nUAVD
vSOMxcD9VPGk3mrr9Z18R2LoTmGU7y17kLulrpKO/VwF6AK7kR+x6yDBRSiPuPo9
U1g2ubJ0iYcq2UzVii3Qs1tinn2Rq2S6gm0uDa4ByNqh2xa0NNNv+13km9gv7nn3
NwSouts7J59cKU+6KOJAhtpUCS+2rQTTfZwzcItd54jNT5cHghmMPfEHmL1v9TeB
6RYP58ItXQnjlgHpLvrdFuGAeZOaqT3MRvokbYtbfyXhjhwcbzfQOo9s020mvHSg
RuWnwo1TK4h5AjH7Uvc9Tx/NyRl/uLtRJEC8GTrSqRW3d6ADFdObs78uZwpMxdxL
I98Rb57OsZO1qth6k3ndRn/0WCHo68s03hJjOS2yYwM2xuzgGKodzq4N2zOvxiWw
Uz+dJVoPaUWMSia6lUykRzoyHys50tvIGCBg4BG4lBcdxKhTZ62eIKDW1/m6nIvM
mSOZF23h+L6ggEOC41ls5DSmQykGWH6N1l8nTVJ+6nnrnfmZ3Gqg72mJvacy5T1q
YnR2y8Hw68aI7xYz6MK52Vtz3Djsdnq9uFFPxh03cE+AH7w2wyDx2hDinZKM9p7P
yOxkO47SNK17P3ovdZi31lIxhMymcfBYNaFmGUlZXzvgE8rUHnM5MDpHS1YsGsAK
8k5NFiY1mhW7R5VXErjun4o2FI/F1gB1pywY+/2LggfSGeNZkq784601f1f6iIoN
DqKquXy6W9bLJmD3yaHL1G3+f1TT/ChW5Dzz11pj8f7hYRHDJEJPWvmpUZ/ykAc8
AXO/YcJ/x+ml6dKebaAis4G6nsiRIVTC2UMJsFcdeXWmezxCeeZ7lnUa8CVVnOTr
aTZJbHsETXrU+izvSOYiSBRQ6zk18JTS0mBusZ/XlQrZ3tLGSyC04NVYgjaxkzP8
GSTVoMps/5SaXzwTn9rqK5TTbGF81nxw+GngaTRSX1o38XTCky2OFJnW1mJbUUnZ
aIFy4eg/rQzNHPDktrchzuUMwtZrSQfCFQ6vjkM7q4eb792WvCpTwDjNsn6NvWwV
IkKGXW6togW3DKZMY5ofBoKU5AMkaTXwz6piVE4TV+jxtB0HW1jqFU8OLuVt3A44
0onAQkrVWqMSegsOtJLh03fBAUANu6YH4ZFZNX0FFGsUMPDqILjdQslChbV6uAoP
q57LUC2smJchHOjJMTG0V30BNeKc7C3DGaAf0PcjqEcG10aAeTWab9wuQ4qLTw8R
TTvRAO6jldBDkH8QVw/65GbO3nEDnVUJPkAPc4LrZBk8LPvfkXNEFbO6M/UnWgYA
c5uFmkWlKNlRjTAkv7xI6KXkAw/nKVqaquoHSX5/qJl/8mEjP1otfxNPAGp8ChjO
sBGGnY1OUiAChkLYX9rBb8Nw6cJ7U8lqQre7cl8zDcO2WmVC5WMzGwZhOCH58U4s
OKwG1Bgb8r8bMMn3B/o64hafabBgpc/1r9qqFbfWDDzVUdf+xxAAT1QJnScRttwz
HnLkFJHipf0Xr9Z7PN61wpe5n0BUy+YvKuNHSUTNpFCfEUoqGKUeMUuJWadTRSO5
Zahzq94kaNO5uLERlZ7jYvc1G90RqAomaEZTcO53jDfhHFgc+gwp6vPJTkHmzqMD
ymt2DC5r5B8LXkTjmrMJwtU6vH96E8rqfpeYlP43LMgJ5i/rvAZbLcIuDUThLLag
UHd5Yw2h5nE7cjw6sXU6TiOCJRLXzV5zElB7QDTTR1ZxwHuh1BySk/AqvdNLrPwc
rpaZNWcz1L40TL3TgJjwm9heq2IiCgdA5b4oxdXsyVgVkipRIGaL20OkNPAAJZl7
QovB0u/AfONPVvrqiCPmI/a9Yt2GpwjHRSGhTK17AP0YNIzG372E2/xVRytzhpZ1
rLluSdqxEyF4xpc0Sw1r+FPnWC3ot67J5JsLR42IU1lTPMCRfVFEjUEx5G9ad6M7
fkV1wm+G8wTgAf/89NctxUgOCW7XN2p0aJmjFZ6/rVWprnnRANtJaC7+Vx3JJQXj
EKTIXasGUFOcFwoTwnDCbGtF7HxDPdsw5zf/gAOcnFKkDl80nR2kQvjK5O6yPpw3
90hbnAqcmxE5C6kLOe8CI1Va6JfqhlSRAZseqgajRJ/Qe9gwN98XW27REoXqBBJc
brBGu2ffB7Znw74xv9+8FPXHzLxFzYzhJuDSu20i8+g6whkRLyRy+V0yRV1Qr+TZ
cZGZe8kIj/Hp79S7pOaQLhf0x6MK8S6I3TSru9SLsXg3OjOIUVTNYvcpn/sLsBRP
yk2MQ51O77QIvTItG9Q0oXlxb27W4OvthfUL2dTtlpAnQdumMYyEkqocHvHArvBV
qvJVMoyfL2CrtwvYT1+u3x6LaTFCZjNBD+UJbRk6zybahcmI2Qdy0sYiILa06T+2
H1j+EVJXKRvg4f87hLO0j3l93GKqu9aCX1Wr4xOtfNDQ5srCbb+uNWlmYD3ELicw
lkGU9x69Ifg6g7bTQxUbi8Vxc3YWfuS5Gd2XJiusumn39TutTRc9o7Wq6ZQU3ONJ
dqMxvpm+Ssf84rfl5e97x+UXdBUnZ3urYG9rq9EIw/6Engd2UqsoYmIPeXOiae7Q
gNuQ42CqsQ0F4JkJfGV+zasze69P/l8+f9w2K+jCtWFZjMo9dX4Ty9O3dB0gEwXk
ALrylV7IraarHN52Cj6eSCWhmAcEMfxQ8fDsCCxUkYLCPzUt+zlZa7RsQIYT+MUb
Uihjj248o7zvhPorPX7PuesinZy8HTy2AGopEKMUO1orxFTU346m6X7dHk4TA+SV
dT0tx/PFJX1c6haKj3byhZYpNMVLz4qc4+eYd7ZM0hd1PJEmrCoUGE2IRZUYwI8g
9NUW0TXIv36SeCH6XRtHRh/vlOucAAgLGFQ7au0HeGsdMrHUiUHWvS7qqchkIZCI
zTAC1NDK5uD0kTZ+yuKfy+mvssHa8DpVIFoEHX5PaiP8eRcwPrvLpr+3Rh5exRcX
7Vwx8w8N6FMilQA7bFdLQbFtIuZ1jQUIMc6U/qIbP0pde3Lm1wDs51QdqwAx6dlD
N+/FwLXbsN5VbcMeLPyK+22Jq2+IWW+sNOJQqFZ8V10Ir73OSO4msdBoiOvWtDw6
gl1RutLtPM1/F8A2ecD90uVpG/hgCoqk9vVa2RYVY2imR+S963Cgi6dGu5ZsI5Ji
8i24Ivs51TGaG0wWp+BVb9DTAds5W+k7NBfPWF/1cXoNXoo+MSdWrRk+8OrzPn2F
f0oF0g/RH2FxE2gR2+kTquqMfa1vPSS++3AkX7SGCwMEb8h1AQhKk8TJruuk9kcF
FtgnqJmSIOSJedYr/KKrI35+/9fopf2xthiSN6DDOtDK4DEDGEBXMryeMaqMz6DU
+KkDQLLbFGlElFm3UYAFr0PzxjUOeAiiFsS4rGHvCmaPPCcYjM9RQzhPNKmz3klz
jDPxYdfH+LfEusYF6jsZMcyrk8NNnuM7Jo2m2+k3m371nlVORRyF2VfSY54SrOsR
TBEjgy5ueP4j6xqKmy7XOmdV3RuNRZeK2p2MFYuYaKpv5GF81c5FOfDCPqgJplW7
azIH2LkYyVDXaNcI9WP0gOFV4xJTnK7JKohgeB73zsYxygdgEnL3R/poSsClb0/T
iFtC9o2sDnW0HMBDfGCTLRGcfW82byExb80t01jJotNCNfsi/oWuu7ym3Zy38QbJ
fR+Lpx6ZAIGvgpdy4gRubJZGXF7EO2iBAvEg7TDsh3YabqIAFCN9PtsQEi1Vr3FL
7RJvUMCStEQlQLjqJV8ahQMAQikGWD2wI7ZYhzs+kujnc9grqYMg0azokKrrkrn1
UShH/s7fYDGZIB+P21akPPaGaFIl3DWQLqJ1Oroah5iwhPxwkZOcrFCsFGGf2wlD
Jl6k27+Nm0KyQG0drc7zbCF9I+MUo3DQYnTfg1AEvJ7pvoLmZ8UI3vnV+3oECgkf
LrNfEsaKezYokgxINsD9xZKoig17R/vkP4/2c+z1f9fXWsfKHHGerQlalMN40QOT
VF4D7SBSF4ndEEm7Y9Ebp7Xp1IOnGoaM0WS9G432ohPB2ZZ5/lmNdHXbynyezspq
Ni+x2XNZWvizqrjU4CK0fYXxxtk9QTdca7UDRu5RGgER+gw8bjDDVTzcsTd+f7/s
NAiewcGqXT6vr93uiaf0vAm4LU39SeG7ugVbYXveZwuyYYiTU/PSmMRY6fW0aERT
XuAgENWkK4GcGojHCJ4m1bBiH2Z5zDJp4J0jHcNZRtzNC69onyoV2pAKOxr0kn8u
4g73qwV2dnaGeo+Ejk8aSDaaGPRZlJlaOs2WXjGKZru/TUwL5jtnM6wHTpQfepOZ
QOUsxKhiSTwvRJZqlQws2J7Zv9VZ82QqTZQrnGCI5eF2KAyJPDlksI5vPWx0V4zn
1e5kv+/5XyqpVtOoF1sLnpbZGAcuLn93hIoqJhbWPteK/7B2MHkJyzU/A3v1Nj1K
VEtga0P3rw2EeqbNzQlEqZO9GD7ASVqv04FrqOHxpRZCr4GPKKu0XVgkPrWn1XrG
ZSBfTyvKF2Bqn/r/T8UThS/LoXDL3AhmVdxfjEkJ7PCQ4GJ+mGf0SXXaiFNs+7eT
Ud5pkAOwJQXYj/6XPLCvRoRgNVaMxNoHpf0LQEHRb+UUd8x9aqoMqj3i3fRBvaeV
w9WEHlzOiWU/AkDqg6I08705nLbFLAKJLMIRKX5l15VhcIsGqbho4+2wPF9mQjXy
3p99ow7RQ9jJn9pzmn8beqyg40UEIHgIoC26t76cHSf51hILOyTwuqgx5AXq7mAf
0Iw/MABoKRzHqF+mMmH4dfD1NTQMXbgcJgHtDJiMm3CRg/H5IRbI5cYX2SRfQWuA
WH8/LjWTc8h6eIiFefrxOR+AfzyMftW6lTLUb6aHLlOML/MYOiL0gUOmJ2FhZuaI
h7+t06F/yXAa3U5A2xCGDId+AAGtgeeL129uHZwHR0eMJnF51upAPPZ7T0PUgRPF
YUGHorK7JNo5xD6eF+jiO0r6/R0RCapigX5oLV8dHrHuPoh8WKawYwTZzXkLkk3b
XRWDsJhyr/c58Tx0peY6P7t+prXeu1R1xzmqeyWWLUOvRQVtLq3mD5Y5qh2+/KKc
GHKwH0HCG1/ov5+cIzsG9VDpPJU3K7uj4OB3c6tQ9VS8/XPf//fDN/0Hl//1TuVD
ZPPNxA+ZQPxw+DoRwDSeSK/cV0zby5sgC/7xcVGJZXXZzzUBaqCfotnhsnXWqiEv
zwvETnlHxg4vvsW9imFH4Qav+w5GdBvllG069yCALhUZim8XlO/PcPjEAKZvrNkK
t4VI4dDRdcF9RKsLF62WsraNGPyl7X2qfDPDYWoy1GQ1tqtLudpmpG/4qQ6L9UCq
Hyrm/IZz4HkxgjN2v/I9T2wXR1H1cByGsLZatgmVqqNLb5uBAvqCdEcM+mCCIMXs
7CJ2oOiyH6KJugf/nUSTNyi41V58zNgBc9MEbc00SHL++XTdUO2moVnWp5f4/Fdm
XRSY0lCRVghbrES6xw7cWuCdfNH4m1aLn+3DYYJNfKPIJiPRX/mhQB4mS/BMMaoq
H2s4MT3tMJDa2ZjgJ08k0X5fptdORhdBgsFJrMuGhX59RGVyjgyEOesgtvnlzray
L69rNK2yfJ9oRO+hS0wg3tJ78GwScyyDjXpzIycZLSqs+AbnFX/+2pG5ufUJe9bY
NMD7eTdT1hX//38jjgeKBP1SnYw6fhZK+u715pT9gx62Zcnh1fk5T/MkMZSFHHw5
UvZpuQNrLEjXMjN1zCWCV1H5spzhV6yLyy3eibzjLXgThtiOd1My/3Tp6/t8npMC
aRns7KyhnLYd4XOn0v5UmIIxPzZyOOw7S/X6xWEchHbxi3WFlLM3h23E59ckYlho
+QjhSszYy1RrPZnhiNxqVy59VZrjRl0dRYgI5NahJCj6azfWaggLrAg/hiSG2Dqs
SRflu5SJO4WNrMSttDXWXDPR4kr1JUtznoCTyhfmbeWeIdy/F/cph85r+u6VR2RN
uFxsBnFIOrh0MtEf1stH0B7A9eBW2VGQ061Es4CRlDx7if2eSFZhsV4y6ixCwWZn
ND45wRk2IAZq0Zwm4GvTc9t+fXkx16W1LSdASW3rRSofGszY5ZQ6jnmJcbdWBZN8
70leY5IP3w3yfggoYz8/6l/4rcJkJKe0q3cmxYMGCMovMpeGibCW+DartLJOtVhz
dskfmaaKxP0IusOPYnn3K5EZB7rB+MO8P8rjgnG5D+QiP3xJ8l0Ja/MfzVxOUBDA
aMw1PqAAtNEUVt+Tn2LmSt+w+ktuga/YOhEoW5vX1eC0WHVKEMtFo4GUtmSHofd2
CP1OVUYZRaagLx/PsGhzCthiBvzUk+yjM2vEeb/wqmOQxRm3wseh/CR9S7BGyeVZ
Uwh63a8NWiB5YcS4p9I5sIB/qjGzlQyoTpJNwrADoslc0JXdAIZHt/rO8c3xB9Us
Zcpxd5yuJt0EUbq+YfDiWcJ6amAhZfWaakvL4mnNz319uiasyUuqE68lTdXqeOV7
thYmEMa7z+JVYkO/QrWKD39/Pn6cMlqyRThqQTu/CWF8TIpOI1GYXDKnhLD6RCve
eou3isciQXMPIlAkijXncA4Fjc6HCxIzP4g9Is5r6HpajD9PDGbi84OqV2tk4HKw
Z5NQg3Mu0jX9VSKFzOLWh9qjR6LwuBb/LDBo461ctQWtwyAyOQGI2TeVSHjWpYAO
qdaKIJtnLsxfRjpeBMK9scbkUFqwvJglFRguY6ug301pNHdEdlfxpYfG/fBMuy4H
X90s5fJrZUE4qG8ej+JmC2MT0oHVP6YDOUDyOqfiPRFkODkZTUFaWaTenIb65K9L
OkrsrSpKUoX1vN+2JjxebVcQPWg9HZVaB6Rxub694ZyTAH5M4Y6kTLZmvFxdILhG
F3lNnGXJZqwmDAyVWKbZphws2u4wy/I7WOWD9gDUeNatbVaTu5oKKQUPZL801oUN
TvTSsUJeXvRn+qznZeRq0QWdYAPEp+19HaEI6dTlzPk7F0zc0pjOBPAPYjms9r8+
6l17paQzblEVLkt85jLuxWrClUZdxv8+mTie/zY3hOUxTtMII7UqSFXbIIApQkZd
RkECaAGeR2lqjLyOt1qcNa0vBWGKfCDtliLKed+CrWzT0TuOJ/yIICskOjFMRj2Z
H/JKyOxTPiPuvjzt3edoyUbcYEDXrkiZgYiH6PvJNGsFtSvze+LrYNkRRRSWKXUf
mTvrHYao9fdOh8HL26XCvoMCqjkcWknbEV7mk7pPxDYeI3zu8y/t4DoIt350uACs
vlRoEPOJKY0ooaqnRL1U10h4m6DQOURYTcXhuLuQ7uxpR4W3gBZ68KlNGmAaOV1S
BR8iR/pQC4tPPrwqvhFw2LrEnvR63sQi711BnqYOZTomuJ2fc6OWsJ8Gg78jRBHM
tT05wwDynQSU6WPkWTmrLmCVV1D2DfSEZVcz5K0TPYr3jkcOemzy0RdvT/Jp6EVC
2oL8HyZnP1lfJe9t/K0nBpivsJQq43rOcpS1RVmAscYkZo9dLYRIB+ZNGhZJA+WU
6w6EBJQCi8CzSOxZFirdtBq6HA8l7lvg+41ZMThcsE5kxnoIPGWfheZS1e5Zkzjw
r27BClWnvta7Rm/0eVjl5LCgQ4S6nfcIFES+JpayJL64GTHAH5wgOmOSEHQpVzUW
G8Y0z0/or1So57vqEakAN9+OB576rVUBPbaR/zRQLAaXrz97x9igHEBxQzgBmXyI
PmcoDhPlrWxWGSS780dMar34Kp6piJcopiPS1KxSDPU98fCQDCFQU0Y7SShEyaU9
WxhxiKVcawjTprT/HpHk39yQTCSG15U5kglhpTwMRweH7K7Xf2km6A7AjEHA6NdJ
Xjfq4xFz5Fq6sRbzQ43NrU3oHNIUSuTcaNhgTCc0QEYTqJ67kq8C32XD75+21A/I
Xzp4uZVPBaZHCsaDcu2j9xLr9zIM72YOD0ptGxfLH54EWzj4f/h0e0LREAZFIkU+
ay1J2HzUHQ1FcyeYRh3h/LWZMKDiK8x6qUNSEujD73VwMJZwiSdEg0mw5d4B22yC
c5awwb4QWf/HhzgGIX8AylUIOnU6eX6uhKmAxLbSeS5R16OC0A7A8cfXtA6SS3yM
S5vosGlbkrN8nzARBq2bHm8to24AoXOnerJrQqouaj+o0xeP4k3FGK79Fb+JQUdf
E9cF7VLq4cwA2gPt8AoqysutJBLJv0vWqUG1Y7bHlMOqjY+FBdvJCEbjq/5ecJ8f
KynAX9r75qKhe4bjgMNXmLbbbBJnm59M1QClrVPtvObNmo/n49GXAEEUT/Fh8fX8
way/18b5udhY2cJs8E/Vetr0upYdqOHX2mD7OLrCEKGJOhYqDGTk1oroxI9jbxqm
76XwjJT8IYCvKOIFWCJb40HwP+lH7Lzs4V0EIG0d36kkSds0ZM1yS5Wo3u9chbOS
IO2j0PJyrvFJMkiszVmFHVb/UKOjysQpSi5NFrfI9sIFIASxOVu44eqizpN4J7sy
c2oSXrDWF3PXG1vxUJXZ87QASFaeDwEOhNFx2oPJOUZTrhzUenmq82P992lBUtSh
UYTGQiUdkhfvRoDHGHLtOs8DJIt/IuEi3TusvhlCgrv2MLRrK8hLEi8oYxElBNTJ
YDSPIymljZScAiAYKQWfh/2ozcY3c+iy5ueFvW+kWMLM/33Xyge04+lqI5imdAVH
LFMjHwaHdsCcvXVFCY81fjEcjT5GJsthCKrul/6s/r3+8aTV7mdPDlpa3eV8eYBF
KfLd+R8PbNZ9VW0pTVgw6cY2F2y0giSnI019gUKq+kBPVUoUtg5cNmfqamRh/pxM
2wJOqo7cyVp2mCKkMj8G/phTHLzQZdX76jWwvfnWE8B/AKorim7ENPYdnepm6Xdj
2yNacfo5jqH5B6bBrsP0qHrIvaU4kP+F5mgNBlr/JVt7y345bLY9MhrcWVBthXEW
/0oh43ZF/bt4rWYHLhoehA87ZtMywVCSDElQitGhohLgSDt4IyM7C1ePzd4T/5mU
amz2t5dPcQ4B2gTdfhDoOfsWHEUnEzVQZ/5bwHF26QRxc7Ni6hJRmVchCYTfJVtZ
2P0seApe6mXtu1qMnmr0JhkIndW5d5uaqUkB75HV17LWdxMZh/up8EpPQTOgK8mx
8u69ShufXxk+s/K0WIO6JkayJQk+o2buqXeujCFnmG58X7MAB5aUhbH+UxQ7NbfL
wiauxYMzht+Y84HDBxSTTmTuFS3rxhb2lpbJiS5obmJHAjY13Qnl4VfGx6ym3zSn
JlWkqjwqS+uK0GHY7j6Lr7Fz5AD/yR1W0LCJ7SMu3vq8Jmf/iZ5s1MRipVAz4Twk
59juMsffK9G9TSx1kAsz/R2sowy22loYbFmINIEePZIlWQuXDRqRBQX8amFbo1nI
Ud8FGqI8RqUlFPagA9YYd2ifpNte5W1LTKK48JQXQyG8p2/ASx2oa3BXVf1OskHE
noQa3XD6nFrDeBLotGbu72+m8R+G243rBYT73R9UP89gNdRhxQ9MWLXr8qM9sG5B
JONtKVjsyQr93n1KKc8ufB4IJBmWNlU+3li5lc591NMybcp4qjueX8IMzk7w5Kvp
97iBsyHJ1eQQkCG4AMOHFdCbai53v7zriRpuVFrjqBCVboB3MZisyiTWUnxIPb0f
dazonIMev4JvjsKqbBeXWAKadUWev6ShMrvDYsajeugUo/XZt0fEftwR1yQYAwiD
J7OrkT799PbcqLkXGPfPBafiA6uoCMX5tHVdgyIWs+ig8gi2k2886/ipfXnw9jHR
Km1V/dpg0Bl0fXYnFl9Hbu4DAH+zfRwXc+KIlOu6CTxjXgb5aenCyuzlwkx/r70s
5dF+PSMuo52sr950i7Zfiea5K7KBQ3JCWu7b3Yij2Pbx5/TmVtmDf4MTz3FpOM3h
OhQci1RKOrTtWARBKREdsyumFA+NCC1V+P8tw+zotPrmN3tsPGsyeqaqdCIfAvT9
PUQqxlG6nNyR+gQqJCuLchEsvAimF2h/n8zxd2+/trKsuHNw7MK3NhB52w+q5Ndj
R+20TzxdVMwFs3hlNJU6psSlsvUBltYUVh6974vz80hldbfphFKHYnHDVaxzqz2C
KfQIMwXnhGQjjl3zBS+gMIhbW9MzLONzM4TVEkNiesNSNAFf5cHUpc75aNzbLeng
O54lgTLGkBDZvt+HKAykM0ujzc8krJbxQYpSelNYMnefRETmesTDqdOy2wEBHnDk
4TNhY//+NMPrJqWht2Bel+0GVr5sfVTPzd/Gw+Gn1YYavY0Z3h+kbDx7gzJGODDd
pGTjOkNt3/UknOW0YVDsQCydbqL6BcOmyuESj31XFKxazw0wgWDO9RyA+b6VqCEY
rMlliCK/aUaNdar41yOYBrPTytMS5AwhSHZSCzUmezGe6r2RsQtQ+SPnyGbiuuFZ
NX07W79Yj2kPTQi4Cagf0jCd2Nx/avtdxyNk4nZujEv12WNvz4VdKjootUepmYH2
HwUHWemga9SG5HLlhIoQD3cfFaH8vwTvvtSOwLu++8XGiZLQSnU0rK2btvsWRcRq
iLMLpt11MfVUQlFi1qrxpMPv80hEG/x4mASTfmumaI3uGqTHoMDCIzlezD04fUIs
WkyqH/6YKcVDhbF9ILK7FegmYXJ8mzD6yusIdq626qOjASHYXNWeyvlL+MJK4RLX
kbGFU6HdMkY5byxwWFpW10KAYZofbrkWy3uAWuunbjvASB/Ws1Q9oCNxKSjmASlp
e0KxAxwtczRWgADabXeJmFsD5qnH/Sl0WSenF4viuLddE5zIshJxqGOwYghEWVHn
7Eb/l0zQNdcDg/wxaEfWr+njw0cAwBAH5QVI9zN1H03znNOjJ6Sl5rquHDEzM7hs
K6H71mWN2GkLfOmm3qSvkD911GpJFj058zendoyCZ4I/W+ytEDs9RHuuGDg6/Oqg
5QmGXaquWyCA6SxN0sjti4TElaJBf9yyMqkb19/DDvjTalFSdyJEbd6otlZ9+eFm
ARTcDbRE9/vq4x2o0PTz3iY+Zg6pOUk1v9wpmGpldRaunLtXOo/5poJ129liICHy
uu2afGZdzRU3woIA45N8Qey3TM8RXbLsYEMkf/lkXRChbGIUwZx+nK3TZTgSJkhn
Vo04z+TJW3e1F0s7A613hmyMhfQYa+IIeWZ0ztWZSjwIl86AXG9H25b0t5CxVkn3
ePWdKmCeeCTx+lg7H9pMjNDfmkkI1DAOmTKofALMOXkWh03+tOZa0WqCCDTuvs2o
sdhzDk/viKoPGJbjWHHblsv4OtLBduHCT1uQ6RcU66BMx0CR8ebe9wcnlVvuiM2x
Fn3y5VBksgr+W0JsOqe/iVhmeCMVXNgk8Uyu5lOqenntDMQtdJGkmJsHASWl70RR
IgQchmDjaHHyWjmipYTDIdO9J+3wxqs1gq9MoojDNvED2LaRgnkzyW+UXlHyHp5n
i2loLlP39+V49vHzP4L3DtPPIy6IrC00b/x6PeapEf52zWAwjDnQR0zVjpjkLzk6
2feOGrX5XJkjaYD+7PppLcnr2hsmZ0fb7mfA+4A9Bq3tTvVLq7utad8kLHEfJHiV
PEkpGFh2MG6RvmozzsitHAaFdKYzILRdrgWWLM4FVrrF3y0JdKpj4C/UVYg7SqI3
wtEiOE5K80Fr+a8s4D1qCngHKOMDVzidCKZmq0GXZQTFxpLQe6G/obfZlfGuxaIM
C3CIipL08KYP1acKdqOHUlTjhe1Y/B0E/IZoHOyT+LvnIzLz7FzDGWol9t4+mUDC
yrgQUoIuTXC/Pb1BeS1tS2BQfjI2l2JZMy52xjDq2FtoCivac7mdGI5Y9QO+6+Ha
q+zw/XNaQjmGv+evS2doyE35Noc8cQ03TNHktDuGX1TVYPIkygC1MRBX4BI9bZvT
k0BidK2mc2hgNBAihjV3S+mxVf/Ap4S0FFA0wBvq4tpUWrAjdFz9waCK6c5aDC1+
WL6cK5+EhkV4pouRWC3PjqbXFlQl0lqZnWAUxyCAVx2bANxoiHp22+1mkoncNS1k
r2VB0VAWi92D1qSWGEYybomRMTBwIwwmTS8kN3ZwCkmMYKzrm4H0hfZAoPaBv/31
GoRHC5M8A42Ll1THtID20elpWrT5XCHvAao49Bp/gRMmUSfpUCN+ZAiUiKsKx7XQ
82oKmsT5qyGmLsve3AXOLZjcm+UQKT3CRBjTC9nSvzTal6zZR3m25J9s/i5jGkg1
uE9YI8czZZGT0SmghdY15hVF7cspYeGHRJe2UzDEdwqVvm387SfUJiRaAxPWnd0Z
X5EXYBQuClojfAtx1jcd+TB/k2HOJGvgs91PQf1NIgIdmMtY22xmm5HrFNGZxROz
CmBV6yaXZwqTsmkuNg6sWoueexcfo5JSExSshBgr/SEw3nPww7JV/7jcHPDrlM3h
8KtQz4KElh55AMVf7/4zxkYUo8UELCrnZTiFvtrdLE9ImgiBK0lHnao3bjI8x4F4
7DZzlIZR7zDdNJv24o3AQ4SGMwkjMZ3JuJojL1LuHQ+MjQkq/0r26jl7D2e4m2/H
+HR7JwDGBRVm3vf4tdoncmWebqfcxEL5QXNaag9LpMCTB/uvo74pjL7MogSlcKUc
gKBpkSptOF2WNZosmJRU6A7vx4FoV8ycmua2zpTlftH8XrTPCAwLY9Cg1WaBFnI8
XIAL1W1qMLWsohf/U7trpo51RMiHDtcVkp5y+xTqsP3b2wFKIM4/ZfPcSOHGaFGD
nQnLPZJ2ojIqxXbIHrFZu40qoZHPZsctNReNbqilZGp8nKyJ+gK818MYUTuCl6OI
XNGrRaIuRiQuJOVgohb1co01PbHE5C73emIX/oX3kB8GcSTs1/Qpxz9rnrOlpV1L
9md3kSCxbK2+cjLCvXqPFy0CnzRKKTim7F0moF+qls/FPQAFfRpxwngmv/cFTeam
mPC+t5hCBoHrWaIz8nFj4aofBLHdQuIS+rYaHMj1kHzKYZmhaYhMAOW1jY/jmIjx
zma05C8DRNHAkSn0TuwKL4fLCo5VPC5BPD2njkn9tIIUTcM5V58FuFyLqZZdt/kz
wfecDXCs49aep+pHNZfcBFnMIdieYCQ04YnNjI+4jvTWYGUA2MTVPOybdHmrbGqx
Kack4L3VgPLk9GcqJEEvSXdYH6yVTNvZQQ5GzOL3sOagZ6uDVznIsdPhPe++745r
hymzdMTbaY8T1ant5ukdCXEOuISbC0E0myihePVtm/ePIIt9FfuesQXI+Mh9DJzq
RExw+1WIf8tMZc3GMwEv0siAqwaltiUDKMP4b3PUTx7UTt+eFw3zfskN6d6hj+QY
TlFSOazxRBdz/VOrG3tbWch7xoqkZV1mVwlNeHdvmjf/mrdWr/M1DIyhK4r3LGUX
uhoNvpr/YZYmh59kmJU2G3FKcF5hsxjGKPfTS3F715JGcGK8qzgBjAE/qJrXbgyb
FybFeXu1arlBhmgd8N0FGarNEYuoF6o37SA/0t9VQDAtWk9z457yRqZOKu+rTfHF
e63kWHITPIyImnaZOMd0TKAYlH2+RDUqipyuyTJGDp1vZcsDnpuWMyUfdZvZ4ZmN
sox6P9P7mscE29omUnUPYlZaIko5CgoD8gAzdyUJrdmvQJ0bLkT2VTWQsuomjj5i
Kmdw6CUE6meE4I/zUGWroR+dSOz3ha7BsohjLpxgqBCrR6L+9Geg+ab9DxGhZu7B
2FvVVCv/hWTu+OrHnQkxuUjKe/YV6QohxbECfTv/99Qiu1KOnOGZBgRUeGSoxO6W
UrpcJb9Q35y4rLQPHiznc3dQP2jtigNn/sCkFBOBbPohhxjRT5mVeCP+TOQHAkYK
mplegYxTF8aPdJ9uQE0sIX7LhPTKlnT2RMcLksI0xVENIOltHDroEzWXy51znahy
yAHnuOHs/vbU1cHDzezZTdzslL7v/6a5SU4sSqkm25CqIMP1I1NPfzMfTkhRLGN+
D4n+prruyr/CoKT98ZTiaOQaVX4AZpnVZyuUZqVqsibUF16JDQC6Sa+78zlasA8s
0R1BiYOT4+YvpNZ+5klWG/1BsKpzSlM/tF3BdhwH82CDM0FqFoEF7qVQ8k/PJC0+
BjoLwmS1WiqOmloSLbDP8vYLN2AITGLURZTnIoY+mTElQVYM311rWT4i0ubo5kUz
j13PTvgfTXCEOlELroR8PbXX8oLCCfnKh4SZBDcH90w5wrhiet9cVTDAL4F7eJz/
+lG3iYLl6I3s8JUpYPjZSKp5tma9MuEW6QgZLhjEtKZdb5q1sBBAFBvZlFm+qve6
8AbP/iZzsVdxfY+1smNNEyGcCvQBlmvFi9RYp/w0bOTNCekivRo/2Rmr3XxkNe/y
3bS5o1QHtB5H13dIOBoNvcz+Pq+IU+PYPc/cTFbqH5iW/b3+jzHz8Dnml60mCLHb
crz85JINPsL/KudFCl24uX3KC6+fMa6JcUzt5Kk4HO99S9b/I4EPg1+cITg9xoUH
2a+q3/zjVos44SDosggsWhlkexMZmNHYY6sbsE9+2ihu4dAlrdXtma61gx7v52q2
UsGKlzUwARdrUhMQFg6edMi8yEJJYKt/uShQxECLJB681Yduxa+nZL5cR2TIyMab
+GVkjx/MJZU88KUpGLhbK/7i1gRkIX3DYCui9Gc8N45Yg2IkBZCTRJgJQj03/u4n
76M50+je9DxAsCRYAu+7SFP5b00eqDRwqej2NmrkiabNtZ7TW/YZtSUpgSvQJfo/
9he9qi0hJkY+cfiL5Hs1PFVacYxYKPCq7RmcNBavo8k6eTtXus23lUwZ5oN1nAjm
e5UvWepJf1mHrHUw89XQuyYcF5c6xuTRLtINQeolOdkvlx07Q/npe4j5dqJwZaeu
jAAdepqcRV3IACgLAHZX5rt91ZcY/nb8JrNfb5CnOXa1GqEpgi6jRMUpf7sktpCz
yuyMne/T9e7MMtg1DUi6ODwTXb76eM+snPzR9vWX1FTuy5mVhcbwTrLj/vAKdx5o
uva6NvDEVQJemeJ4P+YjPH2jRnHYfomWAX0eVqiYQz6b2OqMO/vO/V41WfWNiDjr
nsU79drOWOxxIgT4Gv27uC+awOwMBzLft7qtwJuI+euaA1O9iu9hsDzLTQCnRHxU
OgQGPgSOw/4zseRV5AE/DMncq3QRSV89TAdft43C3cTzY26l7pChnWeYqu4yiZeX
ty8rbfKfHXO8Uf+ochmkXFI75/hmdXOCaiZheveeIu2RJztY1J2faZcMSTdi8HfU
HnCZOPAt7wp8MqlkqJzeQ9RlwfyImJq5/cn4gOXD95WPFU8RBs/WAMZO7NRXgbrm
rRf9TXQV7Ghxz+89OrTbm97dGjG1cZViGO4Ml8j2poecmcCbW6u9JnEuwaD3rv8W
dHlaVFjiBjEghfN8gWKMhP0FYQsGko2dWam3y7+RIwEGeI5KNo5wMkzcJYUfFJWI
9FxvxWKcVPHACSftAZ4Cf8hGLg38Q6W+tGtGn2jcUc+j1TtKVlkJXLDyh+xMf0a+
fcCTyFGpaOwkkY5TEmcWzQzIV0MC27yeK0k9ST1HnaclhKRLgBlVeuWj9aC6UVhg
vjD7eysR2YfirHkVjrcA66lGZTw0NiRthnskD9DT7EcSXEDZRoM181JtY+j0IuOQ
8EvpUuj6xwcG13yYMkTM+NgqXSQmBKL4jXuMH4rtG8uu8DUKISdf6IyHO6VR9G05
rd4+0qeYHnO3CYOd9SCnDcoyHpdYWX/YZw3RAWityZyZuURGN5i1JU/W7FnsY4Xp
suPwMo4I6i865Ts6wtrFnmSMRC3LZTMckZyPIdgds132b8ukiqdXb7bTuzLpYtV1
d+aA0sEzaOSFiqB8Ls1iaBQlyddJAhM38TPDwBUMgNTG7XCCDdnFOBrVPlbTuaAF
CJiLtbd2VF+Kso6TT+qKwqsE8tp7w4/lfqgeYNy9GAQBq8aUgzDxot//Cz3UBQ8K
M9y0kN8d661XFqUqqwhPhe6d922/K4D/yOJkkEg2Anfq4leOZl2JSfSgnIIrO6RZ
v8AbMy7GP6jUlsH2oFhLir7R51mVGdY/5LGhxIixaxzSGQyx17GHNi0vQ5yaPtwm
gQjmFp5nM7fLF64Jdu3g5oSXVQDaUszM7HXjpKXoAVukcZ1ajF4H2i/370Zbc589
R1Ml4+N7j6NWOhffCj6hKW48wfp2yKleNcoY1jDO3PrJPW/m1xpBpCENbxloy/GP
DGm1t5tSGogHKan04ZwAfOKaONwZVlXJ+4hD2mGDZysWOIHF2cXO/KBvtZx2tBtd
S2QRTaQPuGY97w9QNS1eFH2xowC+O8sa/+x3P4Lb84sf3JPYKyJOKhvsxOcfMzI5
qhuWVko80/opsvLm7EfAiuhGJKAsr12kw3Bc3r/OCLz1MdTzjj49DuAuamf8vrQZ
Rd0fJ40+1jbTnc1x8+1nYiroTOOSG9/K7MwLCbM3lnV8N6iECXDimapefTEE9eN4
JyxbREmLyRXNm/o+lJsyJAZuBv/HHz1/7qigAT905RbKhBy9vbr15M4igjBY8ZSb
LcrEDLPdYdFg7thZJY+AvlcQkwIrXp47yPLwSx3tFe5d7tLEnBwG6e30Njs94ICx
UbVgohLthexjxJOio2WLaRWIyFhicdTbrZo5rF4fKTXGmsUVyl9RJ51XYr1vQima
P9mu7jRpuezj9gqont7UYLqKcD4IA6idPWUybSwfi0WvOUCkqAmgQiNB6jWnc2qh
J2mfQussu3IAJUJfkiy9nTnx6/IfSiHCmIfX2/zNdWl4bSKHPaaNNFOe0dXBfxn6
+zLdeG0ytjqN6Jj5OpBigsqe9lpI1pk5KzCqrN81Zd/GxeSql5N3+Bh/J7qM7pk9
QB4P3TUlgLbo6V6VrQbRBKNBr/nwWAmE1aHWkL3IF9GDaExiDb1a8MH9S4NBYa1g
ximv9WMnBgBsxAlTKfh80GnkBYK7+9XIm/g/AnXU+pnImTISrxTAiHuBs5Cnq/M1
yTmT4KYD2Lzxfj0db58GK2Sl6RJIZXUy0wjV1BnBnuMZ42hLGKDU8BZycIXzJk8p
WGBSYhLiiZhnxeGA13gEvRRuCSQgNS/ON9pdCRVMjnhVpvSFDx0htLtAJFjWmisu
58ZNxgmMSy2L6NzvtK9uQX2235OhSvqZZVadzoohlTEKhZMeP7syYBxBym56FJpC
OD/IgV40mTT6zWlF8QTTGLD5SAIdyp1ZvGIdx9COKg/rVlSYt+k9iXVs9BEaZydA
+Wlm5XouFBTXgu+su0cdNU3Vd2HjSs9gDvosKOzje6KJigkMB9eX0/4B4iq6N3Yu
RbGEjd6c4ec8M2tQcINSc/N0IYHXsc26IU2R4+ym5NELaSkNelvewq95g61A7YSh
VhMjcPCNzYyTr3EuNtPCx4afY2Ej9qLUBKId35pCh5gWyXRLUY5MW9aEMfrRYrLL
Haf3gefUzHIq3sRLxc/+vDKp7kAAZoBe/CtgPNsOA74SvfFj4Lfx+zlm2Tujtfc9
8IOeDxnlm0HICqVE+LwlJFcM12sCUH/LP5ZuMuwWQLioJwTchn8HxTVQ7TmoaK4L
hOwr57eAhbD++c+ldg5Im5mrQNW9o8HVi57WO9TXmpP0qYustUn6MXRR0sDTfWGi
x08PPOPp14JFvQIaSDCpzSijZXBrshWZJjMiJmKDUTULmU4vAg+FKun3JY1wvySZ
fqyr8vWA264o5eIF/ixXSyP6NJqD1INoeSUlUx++efZdIgpgfBokWT7BjuT2HojC
D6vw4f5vZ1i6ajSQt4fVkE4SzgAX5dPYtdavgWvTTtZY2RxtaK0yKgf3WzuUO5Op
EqP/QxLDe56QYwW5tFf/xGSbaVr825zZ1HkDzw9BZMD64kCSIHywX+5eTrP5KamV
DDCVIk4R+xeWCs6etMHXWPiS+n7RpJYoZaSdetDks3Olfu8CkVTzksIFFSg5uQlB
tebRd5L0fyUeHBOtqQYRFFV5T4xiiyuB3DMSWqnFAqRs3NYeT5yqKyiRxQ0tXZtw
yimUT0KSBy7shx3wHuIdwiwLGTg4F+TJV87rBQJ6dPCiIG+kjVAqaieYUH4f9hB/
vXe/7FkLgZWTPGZTZ5nrUcPEoPIitZb6RnMzB8yRIJkIwqG7erohPPqEjWflMjO5
ZrX+EqfxB7CbyPppF2uZjtWpbS84CyDZvAa6aqQTm99pXR3Ts8ev4YbcxIQuwbA7
n5TE7ftkU/PVq7ttQhyxPN3PGV2Spqhf5vJohA2rfpXe/vvVR/928V2E/hGrRsJC
EScHM/iaWEHSkwpaasUYoA8na8THxBtiCx+HMWyQYiPs4D9CHGgRn4ypz2cTOU6I
qr/3x8PJe3HpUSTsnFYHPplX2xegjsz2WuDL0v/UjwQX8DnxKUHU0hr8G8gDztOg
Q2Q58O55dSjRFN6FvzkPEbaxBf4hHKVCu4Z0m00niS3EgxaQa9EKCAeKOx0iNMdb
SD4WOPiQW1O/ac1ewZ1h2QNlha9yrURAxN7cAGiawWHmzOXzoPqVCoSntArKoW7y
PmdmNiUtWX2fRavnlj8eCdWvP5xoDMJPgoAyAqZMH4/4vUNjOzTK98vyVCayTiaU
q8jXs7Y66yTpvKSmgbzqNE9H2NDXO3ckYr7bVoIM7BhrM7xeSU8YH8OmDnL6NLDN
tckdFhM11opj0m6EkHmRtrBVNvDmYdvQYDP50blsXTOZf4dAV9s668C21eRLHowH
RJofl9gDrEaMzpsz7lrfemf21/OaRStsoChHGoj//9tXhyYg408WFUp9dVxoQr6Y
mc1Y6l2uVgH4WUR8tWdklH+dyLk08i1/x5sn1ukXQSiV7hF+ChygDzJyslW1G6am
7Cv2aO1XOqNWZztDLFIhOCjDllEgjwRyZry7rdMjq90Xw5U0/RDgW6fg29scpzGw
ZBfKjYZZMRfkaO+SN0VrIcuAA65vvoXfH2/VqdsTsqRK0A89Qkr7vNNjSbat5z38
qOTSNe4VBttllqNzeHuvzVJp8DF66P+iXg6LoTdhzFx25RNlh+/f0uvC5XtW6Tpr
rd8NFf72/J+Zd6QiaQiwb7UaHh4y3f3I0jbat0pq3fQZKYnhseCBNGl9V0tAkZSz
QGe1shpxCCxOC+bW0G8td4Cx/eqOKWoT40guNi0vjTeR6FfaTWmrJJJF6c5CdXnE
ZGxLGOl4Nmf1GmJqRpdExOPFPy2VBgNF8BOLiQ95IMDlEbZcMm78vU8CAJLWEIEl
+0Wz11xvXpBJptL37CHnC4CFCsjvJJaKJUxZl1GY/CVa6Zxy5jdaTXZiyeg5AkB2
Jdr3xJAvT7uQSE3NlGS2MLjMxt4pVXtORPcRTTz0mBJAmXFSj0rOr16/ecuypYnQ
VDbMqyf4Vr5YCWg3+pxY8voBgS8NQNIWh1pWYeHQVOzcGAbupOWuqxlBaIdXcFzM
EldcgFvIEMGne2UPccotDVYKCTjzdTgsbe3RKSBl7a8O+ru+pk89GRIo52JooTmN
HSf5UzSB5YU+wGuyYjCnfdvr3nQUKxs0Nhf1TXgwIjoBtp4Lr9vgn0dstSuYsO/x
NISEh9SfoWBsnleBpp26dft0knJVQoo4G1xwUzEPdfX2+n4ae6XDaj7xzboSdlFj
xbezOTZRna9q288/6XyLelGWTsNvVluQ40kN7oylJGLvW5po2IzMKdMYBPuhEut9
faJJUJZ7n7XKy482jpr5EvwiaCHPMvXF+s3cqmMPezY7KtSf7MtiuFPZvwp6pyHa
Qw+r9nHOjheKDyhyBq7Pi6TT4W8KhCZbaka7Wv1bFHNJBEzaigGvHLmepojMgTKB
XyEEv7yK8QlpZEEH9QroiQffxbSAJbeIhY6i2r5WirQTmz8H+V1nzoEAYg4rPKr0
wK0wzwd54nVm1FP9Tcyta1deJxsueqiJa37NrB1xl1Pinym+GayjCdfqrzBBxXNV
q/0Zo20hPm7IKVJmSxoCQhgC7U/xWVknPxpopgZqkiOFO710W772F8TxU0sOFveA
DsAO+CXAtVRbTto/yYxpFCsO33WktAM0Tb11ioZaowWuDJasdfeDcZynrhJhdp9S
pOx5nA1lHZoAc643G47CESS6ypCPDZfOlYem/3Fi5cpA080hkmxzMU6oeRHzXvqD
UCDm8PAaStgzE9lBnHlKgjmjSNimSXVAuQsUS/Ek+H1ASER2cIb8ijMFBN6zswFX
rl8pOpAyciOGbSe1ocJDoyMY6s3Z4kuSA3xcBewNuPGOJVrrn0hJP5Rx+nR6gC3p
QOUP8n7FAwjqw8SGsE+1BnAoINyiLuu9p5YjazuxmSVMNrkaglVb4EdVRlECDFwJ
y6MK5FgebsF48oYdXAfghmSavsKCOlhkq6SIQusBxuZYP5h7Fp3R+xZr04lZoAhy
tYSeTb+Ozjcpwk/7eCUyOkApmfcuNUqKDj17VAHHRbqvNmH2W7hW7kvKAqTbfhJM
JvyLt4DTd6tHzrKj4J3JHahZEb4s9P9uLZFnln/r1jyh49o+lxcrXp/YOBU7PZs9
Pxw2On64IY5mBWoJXLlIICwUMwEoAcrsJHsPHXvrNSGfQVAiqUkCAAhh+6EqQNn4
wRWgEUsmHNgyejVGLocm82QimOUNFaVAYNlYjM7istgK1AScsKvmQLvlsz0D9J0W
+WY0W032SJLmuX4sEzuzSR0sDG8nSZLDDwRprntxZ8TU1PL4BV6dp/gSurP8g6nu
O2oFn0j0EqKl+6aQ9/qiMDtS/0Z7JKIEnZu5TCvnwcvYdNRMdB5fUi5kcBHqjs1w
dM9KYVJfuEkeLkalcRNiWEjaEySvP/hCyFcHrnJOwBGNYBvNYe2jr2Ngf9crZybB
SvMkIBLXsJyMkkTS/pqmy5/oaiKyGjUNys+grTk0QSuWJcCbKDKV7vn2on6SJoOw
CeDS+xpGDjeUQTp9WYiiDmvoA/ZC+dQGEaNc2VGLYEVld8S5ygCDkrKaEbXN9g1s
3K1kkyGQCW7jSArRIH/cqyFTHg05Yghd4Jm5C+msBvsg8q1Nb29VY84DIZXurUUE
wpFFby68E6H4sfiGpcOgzYF4y3MHSxT2NG93AfVa3UdQY2IpwbqkIU4RClbxlg0G
/Jh2ilSY16kkaqOAuAxckdiyezIXpjfP4JXxDf+cFEeLzu2lKleinuMjWrWUBtAB
U78b6k7GPblWUCV/aE00qRnnaPJ+EzFQreDYZ7RcGueFPVYbXtvM9xgQtilG6knG
zzguik5gYaHVnS8xEvmE5S7z8DJDkloT9Hr9SNc1Y1ss+6DVoNGPJozMwBAv8AHH
d0ORYSTfbric+ZlAK9IENvn4jglG2AbeQKkWeLCW5uub7eOSAY2y6Ivatsaa+ULk
ZZxHZEyWevDSfan2kS64G3hM8jfXh5mZbtMLWkN/OtqEFvC/7s8nIl34uTSsub4P
UscIqXST781xqpVsJoi+iPPHxQBaJSI38oWxF8UhfX6Nf1uW92ULfuoOrG2HUXOH
5DNNrrnD6iyMC2ZlnOUfDh77AEQ6vo/AtyyDIZhEf5ww4O/FUPejfJfiDoXfZYkn
URuRsHiGB7LMUDDky/CXSRBkt8gzNk/2Mj5wSH1ViVsyLNKWIgcBD2wIyyqswrM6
PZGqnTe+AU4Is9vgJdlwW3ouGnp49AznRdVXJzkb+f2jUmaGapU36dyPl1ZXaCK6
HmI81hk44oth5zGqdOMDmIV0MIO2a1Z+eLMxZBZ/wRru88e4Tb/K+3vcSxI9KPG8
EGa/7Um5QPmpkXiSGTm05WGOMDjO5StSJniZytjLGsFITwduIna12dw3wBepOPsD
tqP51Etqzu0TwYmq9ABzdPdGssGuVLFTHJRk0vq14jGul5HegXQQ4kf7cs7VjC08
AMkJ3t55kTOfPMiJlR95pOOYd97WpPhI5cBDB6jvahDpDZdWdMaBghKmk4q4KeAg
b9o9aZuow6UTPe9dw43Bc0e/Cf2W6CuaYQIH1wPDGW0Vg59wYNRq7HeiM8MafFXw
xN8ZLpkCA8A3FO06MMZjQvueWsh9SRln9AGmNAH+gAwWVCx0a8ugtsJgwRkj2zs4
vAnniKvcVB0AWjbN3gv6KV09sbcCvfLeAQKPeyRZg/18JfJa67WM4nE76ntBKHcm
CNJa1pXT9B8/uB9iRpNh4/GjSrIS51ImNLusq9CnLa0AOozczQAtym1bl42uV6qR
2zqtq6klt3OvIzO6THBPYIZdIp0L6e+3hQO5uN/4herOBcka5+SdDt9UwB6HSRt2
6TfMB5n1+IV/uTcx84+AsBOkwgjzVWGa355Ll+4xpmAerD1c1XOPTUndSzvtxnMd
GXwho4bqKIgzol6f7dpdwz9WK3wPIk8frugSkIXawByG0BGpQQC00JFsjOO688VT
Yxq9xaDJUGngkor2aMpX/sc94T+0IdVuZR2i38wjHtLNAlmaD1xN11zDeyJK7Qru
t5FYhubJaeOFOjoKYg3y8qjA592VvOSpUyOsTonBUiAeujFdwpe+Fhu66aaLBSM3
jb3bHMIaf/9/UmT8v7iimRcqdfWmP/V6LrfzLAjFXUsogSeKMeBNt+66HMUH2eUI
D3lg+/lrtonutAMYMHYEbVWmIbWhe/tgTmnm4TOYYx5bBxT+wk0kA1ajUjpXD3Pd
Spvpxfpjr9XNwOwUiNzw+BdZZUhDPY0evGSofe6pCbJsacfSkn/iewNiWkYK7loi
zO+rYtl99cFD2RsvfOId6dMpSqxQPPbDH2mfPddyee0wYL+1qMNNo3vrX7p39xoy
48M6KEtpYlScUQ0YmLCTCg/Oub9Q0z6enckP55jVETrTRm/6bsh1Xsi5OwqLdrqO
4N+rCByBywDqgOCY94+M9HAZoiezje3Y43gq81S3NRW9YSFWAFbPKKnq8TuiSRQR
k5dJpYsky+O4tIppGf5tQZx0+xsaZ/awY26zmHmkMy19oXUlSvNePCTo44OPd6hF
2un5wsehA4E7S5Ipa4y/O+ping/g7njDpP6HVX5EF+AbTZogl6dshPTvSs88Sw0V
z116CqR/S4QMyrE1w+KH0OR04j0n9MGToDg1wVfkQUD79YKNW35zYgH9Z2obxWKo
oZqOtVOxDGP/KZaDAqxrUEteztE9wSd9FC7vRyPVcVKbyBsO7HUCLd0pS2tNBylo
NdvizAUGBsXoVCG+lTmOcdMvfa3r8TkX/2FRa3UbLK+oRT+9VB/xVaTUglMzoJLe
ulMH88pcFD64LpagDQpGRvmTEebxvNqb57he6+DYtcbG4cYt+MQ83LbTJ+QIiQYR
v42/xjxyoJ61O+wb2LEH1fy4aw3PoOoN05+SXb30uRyAILXQ3AnISGquI3pn3MDW
tit1xTXGxTJ838IZM4SmXVGPk9Nw6Jtw/WE8z9DtP4SwAHKxGjEL480x5Qpw8/me
IqCyvHULhim1AqgbDi6+BmW+eraBCWGmp9NSIpG8hE9SJTkMb8i9rtCOGtuNGnWT
i21ayCFt8uCarwRdkpFt7FigJ+buiMyj11s/0a76WEBbh+RNuvgCUgK7/axNcXcr
vf7m+4rf0Nbd8UaoHw5ZJp7fGbI6kkavryReHN1umxydpHNyKqAEmoKUo7ye7hvd
pFUS8j64Xb0U3iN5gKlGq+xpBoSEHZD13BFiLV9VelSbCWDGThkullSRJJl3uizw
6LIh0VYRXyW4m0IkYAozpA4zQgD9pGFV4jlBzTD+zVUwjsBv+TmjotjF80qqkd2O
2t5Isd+jrOAMcrA0pzdi/PwrAkSsw4o7kKHhIwT05GucBtsplcX2b19v+vwRwqlQ
wb2JND/A6uhr/lgiltKRWkma35r9O+gCao9wlbfSr+ZuPjcvJ/qCMKPwzOD9+zmu
MJd4wJgWbESXKIATYY+DSAXW/Qtgs29TlizwYGDuyfEXtfWBTaW+Zunj215l78cB
Oc+39qTvsQtMUMXTWxhiPtP6ShH0pBbLQzhxr76mSDhcEIIEHYM0HtS7ZBMroQtT
gA/hup9qhbJO7+nmX7eNJmXCWQtMIkjtYNIqtuyvDmkKis8FRKKac8GmQoFnIWy8
6ptqDXq/ITQ4qrTfBk3uyzjQ7WtIHgWNUhAmDS3Fh6z/SjVqPWP60yiVw3BxKpPt
EYdcGb7VIrcqC7tgW0Qw3z6mYLDrOC19nsNcKZOfgL0rJeRH21tWD9KyVhIAgzKq
kGeAjWvf3zdDiW8nosqUb29SWTW3ttkDuoMYP/rRe+yzKwfJNgtI3O8Ph/YYh3j6
2j43rXaNW0a4zdIxki6O4a3Wh5izWKCMHXi0xfjkSTEVPPXZEUdS2xgKvNNAUM23
yKXpSt3d5F1z8wN0ZMB+k1OI4NNmW3nrVPkrXVJlIOkDCwBVGjeS9NRq1K2ThVOA
ptipQ02DBcnKsnFju65l0aip4jDJydDHRUGLLa+do+C56OcWBxJstecOqPIbDhpr
2IcHStIdHArHj9Lv0U5HY1C5ld1H0IdUuU9Rg5E2OHlSBDVJJcxR3lDjWERTi0mw
k7x04xzeF3v6Vwi/uQ3062+GC+Z+HoXQ8RYgqZMLOcHvumvY/0lwWYbt9W3j6/vB
nv43Hb6u0CTRMe29eYs/Z2vkdZj9EAa4K0MSKzoGD3/b/rc1G2TCcFd6dyo4IjZb
wTEBB9CAm2JkAsykepFjP7vbtc/a169p+a73zAqPuZa0SYnlmnMPsHBY2OqjzuhI
JYrYi3QKBT1cecNWOWyCktn906nGOnKrQ5nxS9BfWiF4skjVLd/FsAkL4uRl3gff
hwu/fDH19E6IgBtxooWkEpmGtpqV8fSOI11uNcJApLoNUWjAu2RJLZxBpsy3V/k5
NMWEgAMqDABhMEYzvX0/zZ9RsWSM/wY43F87eZFAavYwC0Z6Sgg+wogrAfxNFGR5
6X2Rnw6w7uB6JYJa1LiqJsbphqNrlYKOwVYfnQE75vNXE41fnH27W+U+9C2NlYhB
K/xROJE6GG0ZY6Y5jQa534yfBEho5IAPGNucDxhykFSfJg2LFB4Ff6WPsBdLVWYC
CE3tlFHCv5Y/6D3zjkT2CI2Bs1f5SMLDggiQ13oAUpYNP4MU0SBUrDedWQ7AqxH8
A5+y2Tfdwmb9hkG3imYPZMuoJTKSu6mRlFlJMt61iDBweNV9M+zGLNfVry+9V1Xe
i0YJ2/aayrfZE8qUKQ5DUQvMVDxe5Q2X1/uDmXs6hTaZhYEnSCgzocwu4Uh1bZ25
JvyvNmp1InKHe4WVteTLUh6/qCf5yHfcLK8B5iX/KCQTl4PNI8QqII6+IAQG9UqQ
cB2HBaZgLOuvkKyzyZrj+kJmuQ3iMx1rbMP3bdql/TNeWELwfPeVW/LIsYUU2DZi
aD+J6ZRuq6K5//ynomQg6ZBYP0hS6gRVi17CHibAtIippz1CwXuQfadP58CzIb2M
z0xy/LFGCQLWQm73XZJBXUhfdZwww+sMUMFl5ph/+zWeg1r+lvISInrHtKL38S9u
sT8OhAITvFye+73E9O67eZeX7J5nedwGCJKX89hiFlCcLWi6ldp1lZEP7u88l14+
Ru2fFnW2bSA2J5w4JPi39u62yDC0VwsWy8FKpxJXGqFjlpkqgYhCbu+m44xUajNt
vICOIJZ7gZKBQEEei1/N3iD4QPeNs/fYEx9lAcUcD10MY/dvalfsCVFliRt4nsis
vDQMOsmYEewUbQxBmD7t466zMLubTHBaf8YYQQdslAnXNcjxSn2IIczSQ7bdQiUI
b4u9GNiMFqAep35B2CtVG5CTXCxveWl00QAgGPWSoOcZ3xYcYfJe6riuZD8HhBbu
c+XYOp6PVSSc0gyLXTbrDSG3CkJKP9o82nZmSAqiOapHBjpH1xVoCqQQD+iEpKZo
mTA77QUPCv1lk33/4haspwnKiPYh76iyZQv72w8W4V4sYo4NNQ6yBVCdW5mFu6iL
7xnSgrX9j5NGeu2FTtjpFl1UWDCMmE1MySBvwKDZG6H30lLsprtaNTPl7UJ51HgI
5WD1aaR4KqkTOXo8EJHf+/ZjaAiHlpjjMqni+hzQ2MK0LXcTBAFnMgnZ3Q/fIll9
f3x1tegm4U2/irINx642fUPv+KuXz4zQZNtCTZVMF19+0ts2hE3rtNXjm74ZKSRN
drl6Kd3FnuUh3DVoVt5vbPWSzm/9ajHMikUH+YKiHbmF9EySvsG+3aOxfgnLk0Sv
WkRChauBj7akVM3iJmjH4L3XF5duaIgGZrgzhgJ1xVtstBaTskViScGBXOougd+O
//HUuYL94T+gB9RhUyDiTykEV5TjJj2CQU78+QvNqONbNGxrHQs4h6Od/RXo8olS
4tv5MpqH00j+A5MhVUa/xDgP4J3s1ctoIf1S+4YrZvUaeWpx7qyuSdLIt/mKGHXK
41WYhiGzrbTQFMT7CgRijt/cMRKtMoBC1yyZueixIdf31qNvElKPmNVq26xUF/tD
hrO+qAPTRFHEFZLzNMkhSbWvh5g0mRDdJhK/KeoKXPXbatU929ZA3BV10ydsTLxz
VO/cy0K8TgoAG5VRDXABPbfYnfD4vAa9dERWD5aKYpUEzSYM6JwQSYxq1M9JOEIX
8l1A6wNBKIijOx4pP0iLxlcgZL30Np4U1kb4eLzZ/0TNPtYIqHPK2bfznhGxbryi
WLFvAObutElj1Kdbf9wOXV3Jb0x377yap2f3mAm/Q4hdnJaU5vX/l89PV/NFVc8p
eiY9Ff8CuySWvBhRMDX/cPfcEXzik5rhzCN7r1cSVN5mToACQDj3wOLJ0gsYSEzi
XlIUQceXygvtF35U2Pi7c9r60ScA+1uVLMRpvf3rtEUvhekTYF74idqal6gbHI7f
vWv+cXp/hVckfdVly30+dcPQdgHyKXrEpDcFWxirxFlp+7rIG+HFMdaeGrxIHRuA
I8a56htOnb/y1rnzD74GpAPj74KgMO1PFh1l0fFQj1EWmOW0CimGdY5EZ3bpWVp0
N578g/VTi/+SjQZElurr+rjflxZlqxtMWJI8dskMCoAQX/3o9LUW81fIdZ728i8d
/CxKkC+qbvmSIffpxvbhZlJ4SSGNyJSaa/8fnaQB6vXlsTPKKFeHFatYwp+biRs5
mOJ1Ig79Wqp4QNMGSzFQJ4FnX9xllEKlUGuDLpcWzb5AfLmxFJ87tqLF+DZKl0qX
o+mTvNNBWhY49lR5+rPSYgwGRndve/Z8ewGgGenN29e12txUKnvrCK8yiqXR6rlB
6hO8eJupmT/RdfOHR+b98ZGdxw4SY6d9b0OaNR5sXbfCE1f/aHEQ16CS8dkZXVDc
9jxmu5XvZDDRWR57yIVPmt3Y+ZNLWbbzBiDhiwCDfa3i02Wv49ueqDjOFMSEDMy6
xzRi4vet6O1TU779c9fu3rdZY2M2QJtnvrYZ26Wnyak+rDGIpMFmYHycwJOw97S6
z5/ch57hhhVJqE3n2xldLDJmSPgSepOh8a8gI60JROUyp4YuGw+A/krVNmD+4McA
q+2GwZzeJ2VmIcK8scroMTo5XXmvElIdvWwdKHuPZkExGQ+TdTR8uD3gFjG+Du8c
N6kgLTiJuk/zH9fe5FdCduiAXE0V/hJDCKr+KDfxEntli0wPNwbt3rvk4H52kkRQ
vVO0N+mzFNAz8ILIhTnbeJETjq5e4i9lJIrFz70UTXR+vakNi+Olj/yJ4c+AR4kY
rVtzGY1kpLy4XVN1FDDqM8oUXlgjQoDWdk15+z3luPapAeAwI1FK4BXYYxzG03pu
ZWGy3RG3AiT9v/5k+WwTc5bZwiRurDm8ArBAVejI9vldgJ7B/JYVMdKmHijnR/fG
bMh3felU8oO4CX+ViB/17ZU672VJeoa85KE3rSSJgPsrswJbQ1+lHNecZayjJfKV
lJonP/v/QfBle2SMgIBpFCzVbz8MIxzsZ37AnQGzcIRhdDLbT7fRoeu0wR5cy2Qz
M1sGZflTy8q5oGetDD2WUgNIozxVZB/971wBkUZ9L+LOWBJ0b9Eldciup9GJJVMU
SZrT/orVK8+bGI1ou/dQq3lxb6i0GwKSERR2cP564KvRZFWbW4MB3EJHJ3DjlyIV
aMfLuoLE8TAtx4RIeHYEq8SeLFO03flbZ0E4vuV03tBCVrrsowIUU6LXhmoQ/BfI
4Lw7HWDR5JNKDOm3f2qRoJ8rPTsXULifI4A4n7ZC+X19AJoUpsPWERn1obIgIcR5
5iwDUGJffm2twCXGTZL2cb7qM4NP/Z6dDUDZELzE5devJMaKoJoNl313uUfCrmvy
6URUtifFt4xBVmonIKJ1KlcXUTTFu0fj9iPaHneM9hZK4wqTjOUBzdm4HZZMdEzR
02ePSwo5c2DHbyxH0pzqa/0jFjQ6597B2whtq0TpFXUj40pkud1AJE/YkC5LPDmT
n94DvbOJcWOAWx93aei0coKR+cqmbFPyvZzPQTT9ZxyDtVARpejUJySk8VZHUA7g
BET831yvcBW/ergvrrZpsJrbaUkUnL9kUixC4H+5Jc9dLwnaOVNvRI3PFe7kyHQL
isRjidO7M9h+Wo7xulc2soY9PpCmgyZvaRUnoYFhCfF7KSEKZFht6P+IlcwgtOdp
CMeJyQ+fwXLhB8d7a8L6z/D9Jk7RA/8cGM83nAYK/o+Ae68ia7/6KeWZtcl5U3+J
ksxVYeGBB0CWW8jFWQ1MMCfgObKbAanmIVMr7AkhW5IXQJ+99YEhUBMoRj25dMUN
D7iYlGBFtI/GqgPS1C30it8b4W56cfxRjr8hzhUDvViM5YH3BK8jS40IQPeFmNfg
TbDY+2DBGYUapGhcZ+X7CIybK392r/sxfJcgJySroqApz+kqSSmlDRpWB3z4wDQl
67RHX0WzazzHPRHsjV1PyhgAJDANjhVc8K1/+9y2LQQuAvr0NNPwytXxoqSzvPvR
DLqCC2GuIYDK5WlpPJgDDoITAL7VU1Vsc0JayhZnUj28RQUQ2FoXJ98Dg5l54/AE
nTPK5I/voZs4HaywobUMBXbvwunMYysUOg+8YTM6E+bXpzZPcu8eCJHm73nDYhXy
sdC+scMy3UIDOUOEqUMensXGdtAdkq8uHshiLE0jiGaVJBmrCpkDHsGk8lIDEG8O
/CJECZrXQtp0llhENn1AdD9cDqeW4Puqs4kxJGGiAP+h0YCraiyjh/QvXqPgdgtf
78aWgOB4kAtUwnaR98UpkrSONmDP6BWygLZCWHp4t8SgzauIaf7K+0KmT9J4gN7v
2SRp0EmkaQEcHshpFz2XgY1++Zj8IofJfIxbHASHM6CCNaq4c1c7475T8yVdRO8B
4MS19Fc2jAqlZiCd3WfN2juZmJgmjQb/rBj2j8HR9L7EO5+nT3oQHACCpZNDkBUe
9j2ipWYlJ9kt3G6Z+eIzqHhe1tu8Ib1auoRYnevwTWD009cv4f0zx4DDgINTT/Dy
UDh8MUARQdzaOonZbmOqKSvNhUWHmfZe6z7a03NbuuucMvxlEgtZPCTnvArE99vA
09//a/zQis7AVhqpRQ1PE94Aru27Ekw0rKYA98AlN6U4JhJ9ggM8bEwFyXO9jK31
iKIMPb/pd5JnVcAs1IVAY8RwgaeTleAgt1PcIpXCb9MMH+bxC5MnceM6wxOGLIkR
fphbRgMFIrhxetTos+5MCdLhXtCFpcpNDiUhD9s2uthDfuQhCLueAJ2G0WN7L24Q
qqmC0fe8mmAQFdULgnyogaUs84y/sTQSxcsxjBDE0SBpI5fhszZaMRqa4fZXFxno
hGlNdF6W+dTOpqOllslQsM2KLp+v8DTYq4UT8fiecJi4gXPBTAqqSuFNtMhXwat2
GSKnH70/6J4JKhC5TpJZAzKkv5QrT3J1wkctakH/sXKjHqFb8PSsJP4lZbxo6dB1
GChKa9UHudUYd0qX3kVYuUhBloyFNh8fbZRSRXrMGsHK8iWFHmps8CTPgsbArAOy
/d2lSzuKb9nmN6v8okcKlU81dTwKaEARy2Q/05prKpNSusVQ2UrgOJDkEVy+idbF
cp64Zdm9UKjy2oTUrmqfJ5V7uVm48DVLlIXGcgs4jRuAk7mfdH/R3oVFA+6gyXwl
11p0KQoQitd7TuUr0CtvsF51F1RhftBPRn+Nq6t5I5RFLwJUGwSFKASV16oYCK3H
UuYbEqKQYfqp8PIAqCeM8sjhcUTrG491RnYnkHPXhJtY1y3n2waZeoB/vEaRo9TA
KLr4OmRtHhZisX1wI9fao2Xjj1MH/WbULhcR1gYpd1PdTxi6wkjFM7McdipEzkQo
VDG2pxC3y8vvinbOUod9Nv1nOSTFCd9VAOiaghtHhnxgTdRLPa9KAF/sOlsAfWrB
ECrIxtiU8SCAICNDmAnRuU14LkTJxPv07kRJGB/vyUUTqbh1sv2graoW5YxTk5ru
COumn4imRSXbu3b0CTKR66GxXJfBKO7Lwg7dXreXYmrHUa/ZuroNwFxE0wZJd0dN
2jFWxw9O0+si2LN5WhfUX4C8jbjsxwg1a+lxVMZgwgp5sdUB7sWxBHrS3wg2/H7K
zJHekBlyrHHxuwJbFyZQDPyhMG6gb6DXkOuB6wbwYkmncUGP5MFhpGMY5gS5PUe9
GWCU5oloksgswXvDZVAdwdyLIAQaESLUemqhaqGFMCD33JiRkKMEFwm1ke/spXBi
zGctcMy0repe9QVF7AGwxs7gwHuLT0ZQWtbOS32X11dNKqZJnwSVm/LYS1qGTD1c
HoY+K8tNG1yBBGZBvpoWpyWAsHkIUejCE7S094ii2BwL6VAsOAKHriYrPDfU4PfJ
zffi+r5YTaR48d6FcHZwzDgbwWX6cW9fLY3VhyDxB7jEWR5Wxf3vORODNRn7uApj
keF8d3Lcq4baF8QVsE+etKnsiwxGX+nJ2pY7yVHhnBNzVamjZYHCHzim4vrMdvgm
z5TGMywB427DnOuwJqUEs1OxIBGLcyItXfqj7LsrZo2OvGe55trySIBwcfPIRhcr
yLPV5bwCp7r+oeSbIeKrfvgo+VUrT/HiHilPamjSTiLgkEtetCRSVrTcUF3Cx0BJ
rcP6sPzKNq5f+IerU1Kug/JOIXnn1QE3r6KK4ln+bdj1MfmLszacqKTzSanplBVW
YPXIhXAFOnvE4vlVfyWQY59rQlBBeLkFzIY4eL/ACAuQmK1iS4VzJo32XLvQcqfN
T+vw0JpTzPWpFrFUluFIJBHNZy5biYw49pZOjLDEBhIHyexzW88gBhu9cT+6hcOP
YUbuT2yeCDaMJpW04WkyIkkznSKqtZgbs8UhqIsReJDqRSrnQU47zNF0AIMnVoYr
m4g55/duRpMJt34ODuVzQMENFZjr7XZtHrXSZvtY1dZ7TrKCMrtxd1f0wDBUoYYC
YnZy+hIo5ZOxouQ0CxR/2LYwtPGIi2TbWwIrgT8wBzW3Ai5vZN9Cfq0faItQeA/A
TowTp1kZnj05x35e1eLZ73qlPAqa0ozojNDsjR5RH3Na0YwgUtQnHVqyxfbS45rU
HQpdBMe8eUhzgm59AMq6mnvE44hUc1wgCsxAX9gOKUlj9v1J++lZJnBzJbOZMeK6
vPHh0YYrFS/KifC5Jn6q2LK0uB46+1utZsn89lDBuhNvavoDflyMuyN5GMWglmki
5yhKh1ZHPW/MTes7IXAtRn/UXTbboQ3dmibdUm4fmecWYTO5TRTcMFoyPLhhdsn/
dUA1Ca7A4VIGzpUw0jf4Kk+NbGXilx7CYbVLPCL++wooQDm1mWISyQr/WvjzlPot
1yr+a7ImRfPbI0NOBDMg6IpAp+oO4KoeJOlvLRcF0OcGzbIu2Nei3GPpX0uqULvG
k2RhvjRr9BQAE1Jw0x43DIPkN64dUFuHPo4zhyja3eMukidJthtGrk5nv2QJWKx7
1B6hlnjhfvp6AsYFqGmkLbQjb0kHXlChBYVFK/jSMXPttcSMklwYbo71dzDcBgy0
SOyqV9b2dsxWijHuzsBHWlJ2y7PtLWBwrWkk4uWlkZT4+B8sGOgfNd1qdOgecXMc
VD3f3muwQTyYEMbXFp565Hq8Akg4JRppnyNvMee0w3ZFZTVI8/G3Gvhn7RPxbsjy
oBV1KAg57pW3QM1+tm7LmtUoAIddzvjf8zj5R2bYCJAcIqp9ou0cOlAbmV1Mx4cz
KTH4ok+JyKXQsk9Zou3t/ATUtpY5TnhhX82g1Aje+M2vNHITbJhAMMB7nFIWNJGQ
ymql3FehFtAnDp/6tu3j2I9DsF5c4qyiCmvDwbBrtO2EGTLC6evd9DotlgRKuglD
Y+uQjyoYSEaYvinmeb0kLvrxy7HJ4Uym9m9Nxc2BuJT+T7uBJuqFxGdR8ZNKoEqs
3q233LfQoxdvOlhRIwjYZ7Mqt+7rgtou3i0I2cQ7/xCQAVAcxETj9OTgJQB6bJE2
MpwHSQgQoqRSJVqpBoeSJbvx/0TlCpEqEa1+tnoE4cDKgCW7eXeBhjaVjfiYj03z
Fw9oDu2YX03pHXlXgrTdMiAAaIPLObo7tBMPPXoNX6BWQY7XXyj4iPZCB074Pyqu
D/8mTysjasl3hkiNJEDygeRDWCSEbC6iU6W+zJRqScRNjp/3IUH4/SsEfNr6JU77
fL4A79m5yaMYgNfF1kiW+1M6D4Dx2XZGqwCWR3ecWUGvdukAwj54XicirmjqbKV5
DTHMPM7O1Axc3An3Rg8c2n8oK1yYRvabS0/0Mq8Vo5bCn8YJqZbv2XBo+u7zL49d
v9/O/xiR92Mmf3ySvdhU+Y2YkUDR+T5wSTGmkzis9K0to79GYGCARvXKyC0/Efud
ww1V94B7geJr9WV2vrYFi1KISpqHOANZ9vt7rZtucf/QK8ZTe336BCIEa8t42n/U
94O13XVwQkIko5nsCwRvHwVRY7PzCYUvWVvdUaNQ5jXI8HYlbt7bZdLJ7lb7CXFE
zRiZkdULIkbQq6ivosI2GmbrrRpmSHMG35m+FId+qx3urEPvhIuJntA2PVf/zg4B
L9+xRCXhRkjSR7RsI6hRslx2gStj2o0QRY/NpfMT+Rfq4sSPw29Dqnu0+a9jPnhw
eqSxs+fI+eM1o7pdPUG+PhKZEqqqy5wAz7B8bGyNHuCwuS6mENTEcZ6ORZLDzrRT
yQiXmxNAPMvK64HPoBlguL75nKSs6JLecPm9TqMslZsoTv25j/44+MTxcTrubfD0
YYIC2wjMtQWJ6hd4Cjp9qfdNgPbWtCyESo1/tnnZM5MsQOQAR6Plf85F0VNJQa6x
9bNMbzSce0DP4fJlMVx/Kjd0EG0jTIvYl+mST2GNLfCVhkqb41OGmI2w7EelGDUf
P7XciPKUG2RWgDnZi7QuzdSZoCDXoxuBtmGSqlRLD7ZBDuGuOpD1wBZSr5KW+J5C
/sZDtGfm9oJsIrFU/BOzJm/Y4ZBsWON6Yhl25/kJ3v8v3D/+g0y5uvZLg89OlDj2
AZBKMvduwhoEqbMEe57mZk7y7xTbXSHO0/ajV9ldmy2GoWbWbvgSoUSUYD6bKSjK
6F1Dlj1j8RnRO1sx0okGvY62dg2AE98QdRNu6t3Feh2TFdNasmNB1keJzJfAJKDK
Isl6+qy966ylIxC8Y0LhusRHY5Qy8h5AKG0BxxS7HuQnt8mMJdYvM1rMF0ihbGbk
K88xPNs9TW0MXGgvlnRmm1fzKcJxztjS8ytMKapUbwYLv9YLr+W5X7CuAfM4TYtM
OLEcpMXOcpeLOGiwa8c5o1U6jpHCUiWLM/3dbZDVno/NmgVZlAu9AXr1S4ncB604
vpfa+CKY+WxJN95VWHVG9n148GhVk1zGvpHGqedWl/3DYBYL2XJrD1V3ViwYCWrQ
etrT0M07303MuS5rRkPiN6TDdSIStq6Qg0AOn2g1CwM4wCcvSOvgXw0T1heeN/lK
Hz4KPNLS3S9+1kffePqPsGSmz0a+gyRxcVyyk0wLDu7YTTd8wQWp7mGeSUzFNcBO
/7dPfFpSMlJZTLDjc31odknGC8cf3I9x9ec6x1xgYXF0Nvg4y012Ljk5751JvEeN
DGavZHthlAHCVP64gubE4MwDFEIE0ZV/w7stkxbNNMdRf1PFLeCRwCkIeACo1z7p
Fn329R6p+2RI1cyhxc9faFkWDLDp33LrIlrCDK6Ahre5yGUmQkElHMUwSt/i96dO
hwadVEJSyDPc8OY9f3pGxwi2N71D++2Tp9lGdjupeEI1aRjIIScY1mLN4T5S5ybd
bSQWwC9k1HgLMfuJxCeY9FmF5nSTj5TwTbX85sjmYFe++rdjEwOk2JbXvb5GwsPH
rgifEy96XDW1+ErvfsfEm6XJsThC6EmAwyZmZ8OQzojX09k3xXvUP3g8xGl4+VBG
0YrGaUmOpiuWDiTr6/t0jnzZu5PSznV0QJ5MQzUhBW5ZP0EOb07Pq4Ycr7P/Im1a
jOZ7K7OMkRJ2d4zS8jiYiRf0xEv4BI06SgO8umtJmRf1V0o4+ESO8HLKjziS7IBZ
iVEVnrNLg3Fu8D5rGMM+Nt6dsOXd9jbcC97RRsoI2fAlU+enEsVLxB3r09ttYHDi
b4DT5zNe4gdhu3QHcgpNlml9oxBwDdlgIcIE9jG55Hv00YinN8whr+5kqZoAksYb
HM+JZ8pI8ZevUGFRVPPx5wlDTJJp/S+twRUZidjQgqmHosa8Xc/kBKMahnld777o
zmiFya9o7dzwo1FD+TyiiOCjiVRTEHncs7vt0d7fSKJ5C5+pnpJyelJa9WZMNHnI
oPkEmsLWDKIG/eV/bjBMJs4fd0KKHJgWNh345bKVefcPDDTBjTbCrlJuB20eZJhU
mX6QSQS0F6U8KJ80gKmE0HqXZSgIjW+pOroWRN5q7vdwccRjpP7slSF7y66oqTf3
pt6NISqSPnmyVsIE3iGpfaCnsSzRI3aRHM5A+JhrWEarLApVw3RaqNaKSs95if0w
uyoFBkJ2QxuQ8GX1meHQAkEYnel6tQNrcLxZGT0HHjSFTRJ+8DckepvQut4zC9Ul
spC2KrqZAZ8if8rqVu1gL4Qk2vTvGkDwNj672vQCc83jamnKdyc1IMTBwBALFa6d
l2SdATcLVCViMPJclkfu9erSZgxmd/I9zYFq3uog8P8uw0GTRZk931vizNdR/pFQ
+BxJ+lKDVv0//2qYubRV7kK59S3ER/JY8/eBvBPwB+g0yqx1dE4ArMer6BvSqanh
KiWSHp2EKxJDVDDBCeLROcZbhoHxRcOrtXFaoEoIXGM+0m36BQr8QS6yIzPGZAvr
3jtZ/eLBqqp3dnsdPYsH/iLfuS9U+FhAN9SqwLOnHyQBYYRHk+Tx4hldq+LZy88p
tqGPkVwZrZYoFNfPznKmTpbAvKSuYNTSh5/MOl/cxNjgMRq+cNiBx4WcUVUzaMai
suy1tXbyJ//x2T1hv6XJF2oqLb5At5YVtrhmGMiKXZUBD9IJzsoXpBtJAztYBxRP
jbh4WJhYS2Az0uvNssA8pBZNyVjVxkLeisXvTach6dtgnUcFtLRtHmzSoeFMPvyX
ZFhcG3p+5R9Pwa2K5J/T2etP7dpuMmrX9q1GZDEnbmKCLz0IsscIhuPmQKPdTfNe
Y/yllKIFCmS6APf6skUNtrePuyYNNatOFBe+vb1h76TH9q6q6HMboG4WAld+f3jo
D082ZupMS1Y2HqsUYNZIpfnyyndGMHoN7Ffd2K+z5dhCiPMq7hrGU/m/IbcK8k9X
xdeSKgLljmE508iVLAuoebcMeS892QxSQ8TUnum9r9WLQTaBIQii9CzFWdcKFpYW
OXmQvjXcEd94+bK8gG1PpZugytsRJT59i17GrpXbLj79Lkn7Dgy/J+vg3B23PCj6
deCUKNLNZ9nZFb7NHNktpB6/UJfmlkElOwTDVn1oYUfEQR6utH6BfYAGVKUVpafU
suOz6TPJYc0w0mWSc9E9LrvW6QIlXfoTDh+pxisbw0LnFgjptRoiwZ9FGxRDk/Ve
6GHRoQszI3nZJzjDNmpZ4oxWbWEj3mSI6Se8DxzGNXRWc4d0xdzsy/92qtNerW99
S+7YKDHYEm6C9E6ANmMfpNtVkHkCxBRqoWsta7Ng+MmcMT3bdH5YVhJs8x9QYRe8
xdWQ5SGFhWSzVF8YmKUau14jUx3JjgalqiTlTVfYVXPhehpUUqy0hhkB0ABZPqxr
F3O8ckjT8sQHXsuOfmNNKskhRUamp/4MAXovrxqhVvY8qbDXHxFKv4RrpgocGQLJ
X9VO8JMB0cHOmw76A13oBPOo0AlfLkePBeXpm8FmX4tASJV1AtEkjHMiUREaopeH
7E2rElnyq3AqD8hSaj8k0shwkuhHVvqoLCgnpuZm4y8vv01TJZTiYtprygKA5kfM
67TZzC1jTJVgos05S3d/DtkmfRyiHen26Xz3qkzz170OTElOAEwCMai2GdTe22wr
67lJrHAlsB7caf+m5fXdD5CBLYhypNMBzFKdWjFUPjWaJor1ipk0iUqEaL10/FiJ
H8b5v0pD3cFijUR2/NaiZzVB05sfH6Z0s7xdP9wnE/2urm+Hv1XGj297N35oXsDa
7owTy9E+wMfCVqQiKaW/OGjbGeWLI2u0ZBDClaNOrgx7afLgE6R8Icl4igMzDgde
iOURp/qAg/HkKy/fwx0hbvHy87fhGsLqRQ9ggW9PSRMlH5UWJtjX8ZkIpIV0IWXA
VZWtW/5XgEhehDb7e3sAEPNHmAhTfS3M3B3rw8YGBIE2xEuJgNCtYY4E5iilgray
JNs8mdaXvLAt4cmv+4N37PbBMBnjDDTplZJAjhRJ7yjhYErtLLl/ETageRjn76uN
COqhMtxkwmrWvnxAWVO4PL+wj+MuJDf0c/wNviLIj+V1KxtgI8ldKDS4R4wkLOJI
KrZawaVWNvI3s4n5NCKnHd7J55rIfkJF60brkF798NVC1ZnaBCG44FDd051GJoJY
R3Lf04Rck4KrVt2KJK+S2jIGZYH9CAylmNRO1Xj6gbOiZCsr2Nck8N3htmdg4peW
E4PH2ykOWATbJcWECEly5ZLw4x3tgqR7R3XTyAEeoEyLpVs/IGeGs77OoDP7J1Lj
Wg2ld260CJYPesjoDp2uJBGw8nunriYmC19O0ZCe7QkGHfrL/BUKU4+grz0QBWEt
jqpVWrHCViDPf2OY/pw+KUbnSWS6dWpcz2Wz9lkbcMtDHzCOlvz0s1zpvA+r/PnY
bBJy82x9cdg1o3yoIhBwcDXHZHkfIIEmgJgQAIMIwN/rISIhdP+VQHdAm3KGCkbK
HH9k9c9D+yzHYyxEP2mF3JW21VfEE8qTkvUwNMt2Ikms2Xue8uBhCfFF1XSXTP75
EcrZE2u/Fxukakt8B8BzBCRSU7HcJbbJlOUgDRBLngAXXXpFPUx54DIRfaK+mPrm
S8xW6qP0mcEtcBZF/TLIxoSEy8ZxkcG1SDD8qNpddeg6Y1WBm0f6e7ZQvCbjo7Dx
0xAm+f1WYqdm3kjprsb8gGG5EKOp7NNkWHsbqa9FJzIZ7W5HgEE+FoM2FDsLKw8a
DwZdSwfU43M3ND1S49xpoRwJorLTiZ5Iv4FTVvoYyMzlXYM6tpx1KdTMwY1oafz8
zoWr/epm+usL/l1p+OyIQ2PnaqYPX9avCdTbYdeJ52CR5MXBD/q+/vU65dV1FX2C
FIr3Zv/V9KoC3gDPIbMwXAifHvfUh6VjVo4LFWXIXwTTUv3eD/ByMISjDImDTk2+
Cos1X8a+0VwNUmm3mUZ3KlWXxVZ5ZwEQTH5g5xPt6+6NJLWcVNS312b4NWzQyAtp
pyl5M5A5IIOxUZmZ765gjTY7nrx61H8yQqfqOIKOr0OtLtrOcC7L8Ng3RNxgBVTM
vr1NentiMIrUzk0UuCluwUkTStA+160dUrI4+40FOmZRtvGwChJBHuYiHOVRsreG
E5KOxir93MTNOGOYdd1T+XiloBoB5H8ZZbFoArn/QCLP5sIf2TGZO8tyc18UP8FF
ssY13H6Q6jhyYumXig4IwItygQMFQhV37Ucoed/I3yU6HmuUjom2v5ARVQjJf3jM
2oVOO1NWFzbxMr32ey98TFq/rRYYhbLRgfumundyILVSpPjO9ePFXNBnvOOaF6BM
wKT47Nom6VHVkxMhaaT/5f9Vt+EB7CCwrETE/rec31DctLNOr8xNhj6OzNYqVqXW
0DzwwUCWqf3d6KPhzLxOLK95bIMcdX7/AchmBsLhm/I+UL3/RBcuMA7ZKCZVweak
fxXthD6KYJNtOkITZq3mjEWzlz68ccRjuFxWbt0crbAI1ZSTfhny2mXbn98fAHLm
wfoNRpDoKE/U7bVpc/0sNWw9wVpsak8eErHBYauSpOSWn8j1x/8i/V6wE83IR49w
K1ktJGMlGqYEjVY3RQpRODVszN8DkI69f1YFgQpX0/sScr5P+Kjd9UUyz81abFoN
fDdUptypbyGx5j9MIDNRiMM735QqBSWKJMLpy+YNgZXJ+9d74JKboYN/7zUalL8D
8ziwWdcGwCLYprdwbaT6+3qvR9Mvjqo0KFssBPEXh0s9BtaXZaMUS/APta/AHpoW
BmmmPKaP7XO0PIpi/qhuDCGQIkBDvg14vjoYh0rjPIWYhISVXBKa/Nnxy0E+8TyM
+ktzv5n+YFRYEli6SQRlrigtwmk0D46oH/k9wvyaLQASjqSixDgmHLSW1JjCzd53
sFYYpvdu/65xCCtqgICwEIQ6Yig4eckvA1GLyeHmjVvQ7lvfSLOyzrDPMjcypwef
TMqqWewoxqKBPW7pGeGIU3zJgPao32nqxiAjOkIfsmzYWBAHKisgCUUBTKEcT5R4
/r3A4fsd0ALxDOlxs34bdmwJuQYUx4S3DUfg9/WPEakbAkr8Gcce6QI+q2dwUuan
IL8t0BbeWwFwQZXcXO1mSccpMaCw/DujUDjKQzek0Ra7YcJhjOss4rN5SwEXHEgU
lnUV3nOrJK3hTGjRmr6OZ1KIhANdOLhrg38hYP01sQV6Obv0XR5iKsVHV4n9dNMH
3oRbN3Z/hBdXPk9ey0lM5jRpGLXv8gBmRez+C16fqzNiEmV/WUfsr53njbHUBEO0
gJBSXiiafDKbnaLcGDD+tz6FSIUK+ELy5aAt+Qqklx01Rgr5P10ID1MlMG3DeGE8
HdOjt2geylwAraQGQJ0VrsZyobUoc2vB0/GS75Lm2ImFSGUS2Bx8EGrFx38P7kDC
YukKUP/uCL7kpIpShTBpzoiqHjivJkGnBdXhtn3ar22SUMNEMz01L6hzTglGYhCx
p6f4CRnHoD4PMKVLjo6rX+KVIHE33mG/Mf4Eo4hOv8XHxdS9j/X/A68heSmf6uAD
cy1pS9nFRdBAal2rJVcWzNKmQiY7oFYbERSbnNA8XI2YjpdqxdCgjmT9yj8blhnT
PVsTckaQkeXnoBkIKRBhG3BAh3XDUwmJGymT8kybDkj8E4AeoqotXGVmjQAO9Udq
BZ7SM8AAPas9LFXsVeJLU/1+flUlZ2r9iT9q/bA2hwJqsJHSfhiW64sgKNlaEElP
QTCFQrMynhvfBlY+AnQqXMKqKYKpULOEeMQca6qr9Qow4AHFXcpJbsodgprj9J+6
W3Y6db/4aw9IUGJZomv+aPWRYhoKcVQa7WZbYk4OE2983CgrAPMGEpjxaxhMw3m/
+ZmFJR9esVu0ZMVb0KRPbaqxNrfeaGnBENALYwxQ3F+PIV7afN+VlGxABZE5eFEe
ZwBGRFboyrlv1gnChRErWZ76VXFvtjc7XzMS2DdMu2+KdnxhIqNZQBr7I+wUPLC+
G5Z6tBdQeG0oWsjxEveqFNpFFtl0qJxERDOcDwqZRYoUPV3fYhWd5iNhrx1j6Gr2
OEp3Hu0Eh1EMz3u2D14o29msSYEqJKWWIs1m/EGXGh8OzVFGFgkTP/F0+4Pg+2vs
OsGyu0bLS3ZwsofEBfXdhkwMgNIt16yA8Hd6n5mT7MgHdPwJyuG9wc7Sv1qQ86yM
EjwzJzd7GiQwEQpOtf8+SKrWPA+6P0ASbkuTQpIpPRW8yxFGqBf0F3ImfG1zYJlU
Mrq8IJPYoJSWjNAqqTj4+wDxU8pkTvlVkizI3GHM9mEYAozlRA7et74PAEimd97b
1rT2v4fqOGaq887oENxBX7qi9nyt3SUMjHvHk4j01i0fajdRRH3nkNqRwYH5TPjw
S0QQ0bt4jnZ3+CXzYWf0wFdL0So1Y+iJhvIpndFHzbetZ2acCNe4QUQFWFQJ3VcK
NHq3CSevCAO1wXMeBkt4kd/6urDAMYNe6OD5XA+TzueGNQmOfm7ADeaPKNFMD3TU
7pP9LvO7aBklNzkmI4WSnYqz1xEaXlK0N5q3UunVFyjZKHHEJ9ebKEYanAjtcOXH
cvvdWwNJ9AoZ3bEZZtsAshfEVJmB3M8inLolyy3U0kcPXMvkykmUfXkko0o7RCdW
sS1bchcyM7ch0+FX6dwyzRgDCiXEKrKwuu940vj9+81Z8JWZ6N9q6+yRBkAwf6Bb
fOYq9eBwsJZsGEruVGRa/k2LozbCXjFJGS+M9Vzyzq/SjwPvYC/mC8lggn+vFiB2
5S+BgFas0opZEEpsMm5NvCbs7Xmes9YqtqEczJJjAM/21gRZSWypXlRFz51JjHBz
iA735TeHAeyX9ySlx82ee7JJ8/6h5mxVCNgklAv1IidZocqBryfPAZLnokxaBrOJ
4oD80PBs5U6dnDCpPtx7j8DVDXBh7QjzVMp3LHIr3UQ/E/6gg/RRj5eQ7zW94PhK
/U568cVqhQcJ5lMw0+/nk6KnR5clGb0zJe+t631Hs2mAEqpMKYJcDScrMZm+otUR
hcENGRPFyUoFfRa1lxyXqjgLTVTCn6FEEaUL8wp9qDQF4Naba81qXfIkkJOk5tMK
crK8fgYA9e7cqsoCarXb0dcaD4lvYVnaOmS4KT7t6KTDAzbqYCHVWJwnsxuu14sb
1ecTwvqqXKsFIvhQOjkQTEZZWU66qiuLaUQoejdF/4IGMcI1wQuaBhO27AwWSQvV
95AzwmHFOvQfk6kLtIdEtbFX1SK2lJ39UW1xsgDpheUf05XmKpdFPnShJ3EDBAF7
9z6ZD+fE5lK4iVZ1EKdQIt7K1BjnDncteoeeBBw8Nri8udqYSlRwBUR0159J6LWD
CffGdszhX9ymvSS/IoYXVAiI9QqsnKDrBERtF+0s1UIWA/bnASAuumvtgkLUhvvD
zSOitxH64WD0BQ8nRcnH0Igon1Ahn9FVvwsq7rHqGMMI0MItSyH47Dcx2wtYm8zV
/iTyByxLvJdEDtjWD5zg+RIaucYZPSI/Jyr8CibzGrLtd7yhFBXrd8ynueAMk5Bo
1t2yE+cx72IajegUEoCl2rkP2O+voboI7UuOH+r+Ndx+ujd68b6brG7kodcs8fTa
Mriw+Omm6bCf9L2K2RmHjACy4Nghqki/uThtGripAaKp0hD1azAqbSiH3d+TODzN
qnXDC9BFsYR7tKs+uY3O1dLTIuYYsCHoyRef5PwgrX7N4Xb4tWhoz4zSqPfboiyW
TbcqHike+3cr3r6QOsPIdvTCdpyHzQAuCkpWqSUN+uIrXfGaKqJVXifKKix6EC6+
W34flM8mG++0leGTFgJwLMLqFcpmDz3kP4WgUe0eGF+f5/7D+bjPJf3MtRGxkKYl
chKl4OjguP+9mSYnHp6FH/iV5QKf03VgsP9Abko0TXOyRIuCyY3MfxNkYhMh6CWC
/2YHKaDlbamykji70qR9wPolllx5MciSTYP25oyTZZifuTimwiP0nD4F0yBnu5aW
Hi5fgDh5x4wOdBmPEruH9fW9i+rWdZzlNHesv46Jx7r3MeZN2R67rdEU16GAObAt
6d7jx6yqyXB42EiJ5yEZncv/RusrCQbAJzgkFcNDiUPW2BSSGySOlT3pllghuB+m
QIw1ppBHLeZUH29xvP0niJX5g+wK7dvioflEM7/Aid47emD1mInndnhIfSGt2Qq6
itU3ThatJUw5jomj3A6Dew8rrag2x1WxO5Icvx2rUwOfVsfwUMUtKQ+vNhwkONrn
pComEvKmmmdCSYjsgg2VQ6lRMBV89TMioa1HFthueWkuW9RsxxlR5SRW0eZvHI60
D01CRcwW9A0dD6t4faWAnsefIC+l61c8KxbF45hvcujy3cB3ae0CNzeO9uSldAv0
oIxmcUMqAEFIsLl0yH/Dd8fu7/86yzn+MVesKAVFVNDUiJPNviwttXRaD0L5v5rY
9qA7doE0Q2i6iZ/qf5CmgxoXyUaVIy53ukWuA1KcKpn/eSnapioehWC6oHbqOgBg
mqb8tLoswnL635y70PxdtmqUPwxKmGPBeYONpzy5hteRtqwCC5xOBOTVD5NH0ffc
aL/eN1MZAmaJYwrtrlxa5Nfq6LFuBqfZkTMyUOG7/tFO2gDTVQjN7F9ZGQQSOx2v
2pDUTpy41KN9CHiSgNiWTQdi6QkxObf35QmGrmzqKa+5gacl/BAcHTJiuTVErmf0
r2l8huLYzii9lEurnnY9Q1MY8XzV5B9CBxga2GJsnaEeYb4Lxm3aBtKE9jfUFWna
yxBNlzZA98NC4gij+4jw8ahvkOnsvFkpmZzJa8G7IY8yvQwTpSDf1FKpeipk5rjy
+Xx3h4//DF3NrsZy+9RorEOyTfpKRhqRp2gP4pcfz7xMqK65i+oBOvPl1K8hICBy
8hBpLFk9+OIwyTrApjR1++X6NtT4DPxwo5dm5RYrmvvAsjFp2MEDlz7x1B+cEcMx
0I9nMeCXRxQfmpeU3TE7os9Zf2u8OpoF4XJQmxFjFrUI6TzfEX+zJoh910Hh1By+
ACxksyp+E1IMnDOt4AMBhXOFHt2K6pnxy0Fh1K5PBJ2tgmSBYGQ8xsxy4ZhxKOii
We6nlKJEq7QSfxu/pUiHa9V0cK13HEA7/BZTEHrM+IFwZWuL0nlLcp8EEU9QPI+X
34P1Zb1230bRdM4gkYHWXTvP9AOvyKIREk9Af1BcO+sRq59VzNkg7pW1X0alys+j
L16iLJ27m2N4KsnIPHvJh4jYBRFS6s6mb8M1QcuUHQFj5h0ezQEp0jW+7Tnge0r3
r+hnH3Ej8zOE3cYPHMRsb7E36LaQXs5vdQYZI2CWrOWQeFpB0R2oPgN+7vN50g0K
+4U0zlXI36QnVoniKAWdmm6/RnjJDvOlLRzJsV4m5XzkSYEDXdbC01DVnyTZ7G0v
yt5aAWK06Yz9LDW/JHZtfKJAlHu4USyI/wjHTB75so2H8cTD1VAheE0ZcT2ygkp1
erVal6Al7KTosqekMpj4h+lhFafiRuMstzaLq55dpkkSTTgC4Agj/oyqh0fXer/9
KRjzwk/NwhjcWq6en9DabBP4MQbqEAQTr1aTJG5SMa+glVy5ecOa6mm9Z4fbZKpA
EK0gekFuCRQAZOe0C8PrUO5GxkdQuuUG220V/hrFVBuRQzqfJ9XgbxEHpqUxHxr8
EiKAoVmYAReYrZ9FYd4ndC3grQTs6+j5yNdjbFLo+SE36OMaqxgL78NwcK2EzUvK
pRkXtUVNUqUNyfRh7e7w3bkIXtsdecjSGbs1qNENJajrZsH+u2IPAuhkpMaGOI32
BBu8hj6apEGzTCJvv5G1V7kIG7p546lhQvLyFdnkavUhd2LN2h0Xjkm59K6/DMk+
S0PMvcxTM4Mzd9bnAZE63GcUOCmqAibdR3u2j8sJ2jK9C1biovn2Bp6lKE3nMkZ7
DQVbMFLkKGDiE+GY8lZN1/IH1b4j+B2s5uD0CnLvb6JycnaVJs3+wqT/b65SO4XC
+ZlgYPcLx+4sVIA/JYUAHZUh6aiOFfJdYzYTqJGJn6SAl6yx63idvAHYBmx85toj
0Wwz2fErL/F2TmunfNIG7P2WffNc3VxlH5rc8FgE9upmcwBMiHv6hxKWrYkt9ha5
jNWKzKyAitozhChSbBSNBdX/O5jR3MX6DYgoKdFJC8RjE7FuwcJ5pzuL9tiDqW9C
sbG7YdAMG4YnZ+7e45jFNQrfq5ofcvZRczYZ8cLveOkRJux9LBPIq+bkdGVO9Brt
8kYEDGm/nmM8YlY8tW+4PJLKoReEJkbV0ZvIFgBr8RP+apprHjfyWCrlrhVZtR7r
X+wbYCw3+It4lZjEDeHBaiMoxVk247eA1UgO5+vWpaJ2znGDXjhPbyoHaOdjlnDg
WGBTLQMMYSB6DYNlas5yxw6qFpBSOYmUutnZA2BSfPUJWZT82x1jf/IBie7siSl3
HLW1O+7VOlQhoH7CTYUvURSXUWAy7CGyu5FdUrmGFwuAm2MOyRr0pCdJE0xVyUNh
Ezn0pC/OSKZr7Vh8bcQaUzuiXb2qLHduClsQdxVkUfhcls6lS8DQ0A23lKNpPLRw
KKZJOP8CkUVrZGI+NZuVKfWuglzR75hs4mFpS9Z0YDQbqYi99mfnmUwX+SsBSdZI
HtkT64yeKi2JvuAbHDRRiC/NOHUARyxjgm8a0lPre68oA8fOQET0ne9c58nJnbG4
QB4TXT126ACoH1wy4gXz+XBPEpAxyAf2V6F1gXH8n3fj2Xb58ytFy25FJwji0iBU
oxlFmvbLyyVr06fBtCf7/PMjglqo7PyxCt0cuOit1cOJTXp5lCSClqxWhwNWt2bg
J9vznVA0rL/JAuO4B1UuItILomT+bIApiYaZVeXH8gGWuf2aL625FAZzD013RWwz
U8o851Opu9KtmZ/gLxUH0c57KrB0LL+b0UawgxEn4iYj6WYYW0XwiHvT9oStAleU
nhseNX7vfmNGXVmZze0sDRC/dzM4lhaC3+UnYz4YPd2mL/RlOE6iT1RIf98lEJDS
NL4evnmVHkuBB7uNt+ipeA4CcHKVPswWOOxanEuCFK74KmeZkSfKVxAuvVU4pD9A
OIe3on0MO15owsJm5rdKW5JFGf5rh1nlVSaUhJMt4Uzr3Lsb6gT+sT6LUgbG7ZsS
vg9k4lufaHk30yx6QmYR3bbMQXDinsHKc80IFXhSD86q2C9utQ5D0V350PB434Ed
SZLWWX1A5MTpO5CS45Dm3LSC0OJfvFyTO5aCLKcnfYIaZOUbQFyC4ET7WWaKYXSs
pWK6s0+F5+op8mAkvSRjGrzNinvFwtAP4Ib+IAOD1TODwCIjNXJNQjx4hcoyC2xZ
yWBgvz6SXE0/TZEXAoyZ6rIIU4ksAC6LAWKEWBbM1enfihKu9xQyI38O9u97dHxv
lgCoifN4KEVR5CGDtaAYat0/6dqbLOwbW7qcRu7tIq/eqaCZHNTiNL7Jt/HiEyQD
/NaL/Vav5iZVDjJ0kfNHyc4m7SapICbHRWM6OiYOp98DVoe6Yfa1vDpDQhhWCEbG
LLA3/CIZ8AQXy6nnCD6E6CpOm7iK/7GJhtGItDo6MxmZeRpVarXVmS0+I0c+URLu
chW4t6ZYOig4R7XpYxkLkWWyDMxIJQnHou8YtQRyHq6ynNRgEYA18tF3PuEP5REy
1wLta2MBe0JM88mRDepOAlX46U1MdOBWpw0cPvbMRYkeTHxYBj31aMJF49IgBhY/
jIjy5sNPMdbQiiTM8Ba+FwF5wLxl00ibwQHhXRhA/kx0k96vDIuIMaN0Jo66sa7i
XJXRR8Lqf0dt/Q3CQEru4uA+NGvWp1QCRYAliPS9h0gmKFS8hQhnUtXpaDBDZzT/
1vTAz+nicnIh+gfI3qLhiX27SheEP2kAeXymmmgTWm47O9REaI2SP4AyX/jQ0Fdt
r0YOiTHJ6LhUEoPWq+/0yfE9tUcDOQqfK34aWK4WuAnyNcycYw+VmJBPecwyzbD2
2JUjkbGQSKgV3/gAvniBbvXnzMr6mTotMj4lMFnyd6TQyMLg5YS2brweOsy40JJf
Ip2rsUTqaKPtPTYA+RD4cWs2SYiPdZNx9W4uue2ETGKYzF2kYzpEPtl9gNlU/AXm
2DdRwBCc5N7W8dUx54Khntoqzhi7f2p1nKtBPanm0bcqs8wclomlXxkEH1A4fTsS
Qh9ypVmQHA4HB5GDWG4rr6ovBDcBiHgiHCLoVRgwArAnmV1Hl2sTbTM8M96fyI6Z
h9NJsGv0mL4mak4fDD8v52/hLGPiuXfqdPN5rSmSvJK2kQYqc1621lkh0XqgzTG4
MgACnzMn2gwXt+Ugr4pYoEqfCzLoeY//Af2oFPyit/05iccSCI3CaQ7No0q5GWJP
mgSVn1UgAonOFLAV44t2+HZ0sl5wDGiOkwbjJrzvuTlCHQEDdw/ea1dczi4FFstr
MlLZw/YNEUiMh7ogtdROnN0Z9AhtFQjgtqnf4oTIWl3DcfZ6nAiwnsIqQFdegc7x
hKYVzmGujI+tvo7W++SzBDifQn8O8QZTNngAf/8ht7eiljyLvhF94NqGETg704+w
mVfBxDtCbLiUubgJsrFVGIqrmmuO0p/mZ+RU5mSt8TyZCUBh7DLAPlgH8cAw1syN
wlwQW6Jbcs825evnQC6XtL4n84W1J0T8WN0pZkVXhT28Nf11Jq93skGtynNBJOf3
n8AtelDr7BYluRVqPLx+nSZgpsuIXGa4K5PJhOmhExgWql4adP0At03AdiH1iUWZ
5sFTnLh+Dxa16dTaw/mtz17xTgHe9sd8fG4n1S3KMDO93/AKXbpYlqaCNrxvPjqf
l5k8XQIwC2Iw/cTUB/0NbFQNeAzRtCjxfXZnafxlNWZDlpH8GhMAmYFGK4qUvgyH
8UqZDjux8cHwlGJ3F/oypUXNnXDporh969S+tzHt7sZqBug23i9p7nXfurrme2no
fSAzW52XIyj8NM7hg39zDEg8yNIV1mIoq0PQBkge4Etgls/gFVZ9TieCnSSSgXc0
9RhKW9OoK/SnIneAMG0b5G5HwKbfgv1QcLDGsXyZqb/yCtas3g/Ad8NVe6Rzn4f1
5brGWenMFHnqsydpZFYc6q61uUZ4FokJ7QVNfluGMOJc71DOv9NxLJGL5aDvVPg9
9i+LlPgBfKANVjnZkSAa/N72yJvNSpU316cbZsfmhN9Vm/kalFhGq+BqRXFo7EQ6
JxuCySFEyuAmIjW1wiq9GJSefx1XZYKjgDabavIwxEASOrq2jgYjuQ0CDuJiID3r
jbOHj1F/B12r9rCXUpNTWuLNccV4EKxttR0PhteqMvHWNyrLNINHJ7MsYi0LyQaP
jXZYc8/+gyzhVwY9QrzXX0axVlH3UFGIC73IeW4jnrAFESBeE2Bp2Eq5hNZ7Z5u2
+wjtQy9Mzg8M0St0fSb/voHT26ibCZICieUawAGVvCQpDaFbRpLQKEE/+nxaYwp6
uVJnCK3BgiJkcLq25G3UCtxDaEpSPJ3Sln85KNMigYfbaPBgmk7IcmWSnS4PL0fK
3xkV9XwsTXVUOC9BGYnLMy2S427NCZK7PllRzoX8T50SH6enGqkoAH5WxobxX8GB
AJm13B8ZvL+ZCcbA5CGiyhiwPjCmEQWxgOWyilNif+p3U5mX8qM9P3GW0Cef1ggO
Vo6quJInOzHBtxGD8ZfwoucBhiZc5l288ggX3IVCEGSHf+Pv7BELglrVEJJJNdKR
wTIXxHJlTmEigjGgfZqVDqGZy96fVNoXYZCrdRjk5twuYmwG+VahXwvnxhqN30Hu
2ZGoy6D8oAoM1+80TBC0Wo05+QrvnIPx4g+nZZnDYKzb0sTtzuUJ+oXF0qd7tuXw
EWqe43GluRx+nMPPqoaFWcHGzf/7vOby5qxY+7+eVBgrWcL8X4M5EqINGu8p6XUd
VAESohD09W/U2pLg2QwNwMOB5h9GbhUL1x/bst9HmXbElrigieWSgmRIakLIIfpb
durYMq4kzmCi/z+clFVwblEKRZGgSkMRCKYaWBTKgoGFB4Crh5EGuicff2vSsZm7
5h7w2Cxr0xx+lDg7pyg0tOWQvBnb+xNRv+W1sL5RETDGS6pabVzeI4n0ofUBGdkL
oWdS6QXKd2QCX6uc2ont8Trz1PI+7HP2e4hGE3tTujWJtPqt5bS0WQa30HVwSG7K
zmgEZPCy+HkJznLqikQ/740rq+c9Nco6q4A1Dz0p4ftRhKiFhPO/w4efSazSdqVO
LaIkpMIT3lKttlF65dUajoWWglsQBS9k3cd1SoxFe/9aKUSGNP5wJa1IctlgVOmX
BaPzINhxEf2btZQ7EvpbAUrmeoJozXnApu5RGmydV0DJx5gRmwciFAGbvROP6V0h
Vkt5gNp+eKk5nrmD+BzM5y0jHIqXz9DchYDXByMm3kqo0RY8AAHEGv7ryzIZeH5L
JTw+Ebg2OM3S+qr+T9xsZ+7GfuFNWJvDg07kvI4xAOZrb/lx+iygtFs6TvMptibh
/RWp3TBlSPEbJ5Q71c0GPZCyxKuN2D44/PjRokhcSYlOJZft/8WRl2q9EIKFF0Qs
lxXJvKQ8gxsO4L8NH4+BVBo/3V+jE9DSBah1FI2O0zRwbArZRmQN65No+Jjj6K+7
WwZryUuppDzpRFkKtrd6GuexvOE+VZldvdZcCbwZg9teXIydDOkCtUJO4Xo78M60
cophRyvqaexT9oOgXmtv5ye9xU+XfFL0uOvPpquKHKrsM8PBy6nRRaovR3M6MGln
c7B702xPefAsxmq406tIOfeS9ufIKMpEYBf+E8C/SNfkNzlp+4Ng8beDWg7m6yC/
hb92tGPTztTqEml0GeQDu5NsuaKH7eKO6etV4R9lpn+27n9HwHWtF7J68VtFAL2H
ouTP/6ii0bIRtC+SQabVS8S6oBhtFkHUmwXpN+d8awscQ4bziuUrkrId02cLFuwF
E7M3y81qa1kXf9HzWi2uzZudblpz90CkBnK28xnMq1SNE+10A4IsvtC9x/zebRkP
M/o6aPO1ALA2Soh2hizH11gv9gxIByFO+D9T7qYmvqeBvUC41/ZKuyOMEz8mRaLc
k048hNtDvpVeZthIhxmBCuX9bQOlUtZXiLmlPNlhdDI5cjHzYWw8c8gT8F5O9UFs
cZkEwodYHJvBqvIiabx0MokbkHyjKaKmtPAKarVikN7+s0Z5Tdxpeb8FAiWSemjE
lMc7hTK9yf7Ey3nWq2OfLFOlRXg+fkuVwG2wWJxGerk2hDhvEs+TOBiQAVuuhh8z
8OhRQ6a1UoIji4eNXOMGbDieLTkqpcmVseSxb3tfBc2Uf3AyGgFD37lvSAgqdJOz
1C6RZBqtMMAABMsO4GT3bhB86PLfZ7fQKducLiLvjFFNuk0SeSMZ3KQPcPMNf3FT
YDJiPrUXjVQHSxIMf5rZ950iupS/eQrnvf0y0yVjh0aPs2N/vvEI1ZDWCmIvqtZ1
4Ep/UkFDX2wtqv5EpltwL1lUJmAS48UEZX6FXQmqDUdTvMEOwUwIWPf2ErmD6I2L
jvq+zR/BezfrpdBKGnaIwnJdedMFKgpQEA0uC8AksHnbN3kJYSTd9ks1WYAyH0ga
ZJA9+NGJT4ifDGmZsWw+CnMuZ9WEpElmCPesMNkozL4A5msvYqYdNWHR9EA+sq5J
gUSKzFvorsajM5BjLZ9AFLwnuUdq/ZmWC/n8rOShV4gGeOQLTlc/B+TkELwdZI9I
ElzhubTX8pXWUYfaesq3bi44FrwzTeZ9ntZxOeAh/pZSBcmwqC3d36d9YnfErKdC
FArQPWe7tDPD4z/2lk5JUj0hZfdRWnkkPTDSZr6tNxasc06/Lu/nQpDtr79VNvmZ
Mqh9bvB2Jph4AWbdqBXyCYzou5d0EVXHxAoNlajRY4vqRwHhmibWNjMEZdbkTYd3
O8SBgnJrTkE7ec7qQvPonuh7640G8Yu1K9B4EOBQenCFWudocipEUcYwSsqUS3fv
nzpHIuopvRmJk3l4FtabwSVji3tol2/H1vBpkjCmYXQ/dT3WQgjYn69haKIdRRWt
LEb52gVpV/484r8gOGRqyEl/xKolz4XejpwTSgDin0iIfD9HWmvbSO3b8fJbksQG
MzDcFxFsLBzQPZ+hZF/TvIjLcxcxyfexQry+msFdvUOU5zvd22YFB4TxqqWHUfWC
PrOGu+cw6nKYTfXIKqwNTzGdfRrdIQQr191n5DVPxe6jiIoI0dBZX5ps+ZGFlRek
nTzCYih492aj4dc0sNIz3+qCup684Lcp8xeX0YW50cP9bOoRXNex7SfjuWJFmNr7
B0iQ2WUVm3g8WbB5xpMFIgwybxNMp57cvxAD7qCusHLyu/74J43hT0AeYYUPtc/Z
/kiuvN5UbMsrV3RX5KPdTrUfwHby2jD3ydOryw7XEIN6hSiT+cIc1vJ19jvzrbYr
FRTzT2qjzhow9B8jpX0wmExnC0DiblJ7T6jxVzfgNK8tKVK9IoZ2Cg5el9J/tvKI
Up3HCyroc+cXOeZgqTJ3iWwB+akAtypKM7LLjdiWgPdpsSFUcP8OMP0eZzqfq4/0
NoOHILOwHDbELmQ3YMUdi7/IgP3tBlIlc2l/9h9W6qpNdHOtsG01IvbZTTjf/iue
f+bKGUy0tQcsT9poXt3ofi9FdX/xdnHYKhACZI7OURLEpyyZttXGc2Dt1B7Kl5yM
1dZqWovy/MnylPsddazKZ3nxevluDUczUIROjGdP1cDXV4Erny/6XHK1zYH0l7dv
imI1JlrVpWJ+E75E4DK1rYI1SnfqMz3DYq73xanEkdCLdiGV6em7Tpc9/CY8Ahy+
yQc5mHKpZMyUEdwMhXR8eoGwjxrtrRlWXVLu79WVZGGXbyh0d98UhnFyQq0CcFge
tyFsUqtJxEtueOgJb4ked7dqh/BvW/W6XjEdeD08qf7P/icKrKrHh2ll7PjwZRsM
zL7NGtnp6mfrbASD3n2VQ68JFhDAzQDFUbeAxEWYB7cQ5DvnXOIN2jf9JuUEjACb
N7wLCCPTUV0RA3uW1CVplB7jsoikawfh/jd9R6FlbUggRUZ1UbG3+Ndn+7qWzszz
21EnjUjGUsBuiYtxnGZst+LQwrbwzk0nXKtkw6cOuJnNkQDMvTkkiN4lyvLTHeuQ
YKBuRmZfClWjbAi5WdBIC1F8lM8273q+/O4qXjE+kYR8tOjovHZrXicyjVWhHD0V
BkSpemTx8POEz7y97Mz1OX8gsGR6XH4YfToDgPal3s8pmjzYfSwHAofOz+MS7MOP
srzIBVyNwWDzfTubSrBC51CmThL0m234/phuooIifL/dYzkCHU/XmIf7//TdSyEE
LxP3pWxQWBMb2uBpfaRSro+7Ov+uIVomSGzsNW5DGU+hFSx+9zJkXzKXCOA52XrJ
Amb1xQ+8ZV4IqChDsw+39M/AgQ8KJ4IHxygs6pe/z3VNHAwzLhLH31s7YZvbPGEg
hV3LQoO9/KrucI4RS5g/M2UFrllbRTUBzSGQ5+zG7us4zB2NwOxahqVHDbsaY+3b
E9zQP5YQqNxn1RsfQ3tHq3yM1KogeSG3GTDMqPlD/ergFkjrdYtnSX4TgnJOQMtK
0+yuf6sSF1h+8Dc8pm8hdAKRNBjShBGdDn1Rnl0ifmpmHoAjLEUGxSfJtLb17cvg
n9KWrlr6B2yP9yCtSU7DD7iyC0x86SyAki/Es+2+ubsICRf9ikWN6oy+VFXQfbHQ
jcJVPSI04Hajt2PGWG3JVCGErHqHupHjmZ838c0uFogWr+gb5oySOtvXAXyvpFxv
akWjxhdwpJ3oDgfxbGHSdUhQp1xPdFUc0Vdg2M4b2PCWhcvz3J6cATZt3KrK3b++
OEG3179K3SK6xM8WKI92DObHafiZHFvvBPrt6incIOknNBSacqrgnjpxBMUsbG0L
iIZ33fUQBD50RFmzboPPms+ShFivmQngfww+G2xRGmpeqM1zuMLM00ZFk2VBEsFc
AYRcANSrm7y08D1Qv/TQT2oBYIHJpeBBt0MKtU8MZRLce/liyK7vedU5ZOOtvZHV
R0yN/X1aAZ1hrLG51lMeg8xZIygZ3KL3oGgjWPbbxq79WuYevjtLenTAIBcD7dPQ
KToJ+rp0MH5OcJdr8s7CAy5rIHEggIzL1lFTqCVX6FwYZEsLwGgkGGBWCKlWbMHP
zVy1mGrE18SNE3XWpI4bm5ahic9ZpuSqqNXeXSA4ZTnEcavcYqhabc1DK34dvgX2
Vh1/qYzXSHorr0B/NR6OMu1IKKH9kynExjROT+gOT7s7LNUoP50zLUMQcDVQL6d2
+sPD/C+GsiFY9I+bNxDUx5Rd71BsGvaw72tkaCy4gU0OKVI/pAugaTO5JZf95/SS
L2tZR9Eglq6PAoVgyQqjW7ePqbqY5NbgmNEQn6qaRV2mDb7QplclFUjGgOmkASNE
T4u8NJMfpnPQcFjEB1tCA4pNyqoUXs/DOpQDwsgJnYhxnWdGx4UOfSMHQbtfNxbn
lN/kPjTk+XzAR/utUbMDSEyYBVi6BZ6j58QY3MYPYzapR+M0OzOyttSypgRv4OZd
FAr8LcLRQ+xBiSMqpDduASjLXQ+pOaaczUTPjnQ1rJtG8HVtXGVhbiA9325tc2Y5
9NZUI/2SgXxqU8rNx/6kEXMtpaShaKK29fXPteV7XD/8LGByw9CYC6JXpCQagZ1d
iATQxmkCfnC9m5rxqP15aXu6/Kxi1w3rx0lptqrvVG55dVA/IQ8mbhU5i5JKOg81
yIvWUeAu3b3r/zllKMMqtrNRk4gN5/M1XH/mFJpFmqx7m+/yPAQFia1f6THFLAU+
VV7oc8MgwuFlE+fm5gkn/eUZDvkspjiy4Hob3TeM+qH6wvBXdOEBK2WVrHaQVDBa
Y4uDHnSTuEN8kAEKikOPlZdBKoJMkVyJL/Dn1aU6mzXDRaMW0wOic6JdnikUFhnT
M0syy6+KA+KscB4oEyafZAL/zg5OsWE0Nitd+WvLYdM+rmWD3En4NN/qcH32A5j0
U4XhLweueI0OxhquMJEn6CjBdd0xLERglQwBi5LgpyE+r54muG5ixsyF6MKdCDfm
1xJdG2gfboP5uvRPqsFNDBtyIEpfQ30fBBIxDLDJDsV9HYaavs5EY693StAegyVs
n9VeSj8sUpLT882rpc7LP/cC5VTkvFkzVPETEmDAVCkFe6m42sqW/oqp5NEN7G0J
kzofAdKYs8w8i1uBFTDwJf7z/4I/B+I91erKQwvXizokHeJ4eDDh5wcvdnw445zD
mgcK/bs4ADTjo7h8ab7dVELJT4C1jACG4Tp4j3IyCF6NmeEhFTytyvjJ+pmiaiXf
NU/v9n4rblIWvqkGlm2gvLxzrqYrpiXJiZJT9NCLeRRfK5KlvcXN4sRbSVMYa8u5
YFa1vtYCbxIw818I66rnxSIxg4rEqg2Kaaj1XCDXTkyTvA5kBIeGUzmkfk9FLbX+
gKKPMpJtVAjAFdVO/PDAwUv0rW9GvulBpR/UkQnnI/kJQ5BPdE2NVF65dHRDRzrc
lLCl3IkPqv30uSp7/rZL1IbelKtj0v1nFZx/bA4bkhEUzRKBZ1SWGyy5fP+w7RbD
WnFf5Pwtz5GgdtwVKY8pP+QmXQi+gvFfJ5GgpU6KulwcT6ZAaEhbw5pD9jAEA+5w
VYeTenPqeUOHYONf1xgGQWW/gm7UQNCnZocRBewGGNvLpnPPFD1AIQftc73K11Wv
um3AUc5Pi0fOozz4mm7CDe4CiuMsiqX5RyyMEAVC/7d8B+QQm9NmlJltRSOTRPRL
XHkBVTUuQMnBHMZfqXkS0cyZ3eW5jNrjVA6DUgbOZozQf7cqlFlgw0gpd1ZC2xYd
V9KU2JQeuV/aLFNJvL8TEW1nsmDgBDy5WbFUvFOpvasYqan0jCL4nJ9xotH5YAxu
NDeW7LOG6P8mWxgpYqKalofMJ1dDngYhJeQCbM89rEQ2xaZuxWe4hUesrlSh6Cxu
gG+rjZo3y8NE6J+NVjsunTzjeODkvU6Ih9NMlzxG+nldFxpe5bDtd6WWLyS8GlmB
0iFzaWzArG6YEPQPftYBDDDh8iTwRG6lxpKvh85hNUqVIFrREbdk2tSy2vllChD2
Mcn3h8kc0WASwOpqt8YecO9OQV7xvN0RbC4U8sdhjud/ThH4oMsoGWtZx92Wzl6W
o9Y1fL5IzEGRGzrdofWWz4uO+rJDLMTuSOuzUlvlNkSkSos59FOHDoheokiD6UXf
K5Pvfz5kAyBCW4D9gPWEc7oqjl/3SnB6jG8n216yDGVX/6sWQGCjmjcccfz6Cusb
eYePoTzXgbo8NY0Zz/JiBAHjH8rU67OVB+TGnhLYsJ5xgqHDmzkXdMIGq8Ue1K/R
yasJCranBGUrjq4eGIdxHu0M2KgzlN7Zso9PVhQi0u8oZaQGDuWrpuxXWK6C+boM
366X0PW21zP53+VrmrPlf9Ib4EM9RcAaBAXek3m+lJcYgHShajfFdsnmM2/dm1+q
9B63tIQid7KMDoRhnCrjHoAEtBX0S2/nde4T80AzSQ0AJkcj/XN3O93zNGqKsAA4
HtRdBIisbRIev45wmKuCCLRTsvhmT/Pj/QfrAV+SnllBb4XuaTaCEHJLqOUrHJRC
uU1TMhubOssjr+bqzL0MSAgfOQ3BPbiJ1oRjOJr0NIlG1Ot2+l7AGykE9bwYusN3
ftDtF7ZBCMCSyKVDHRGN1vr3D/ELc1PKihV9EdzRZFTTw7fyYB59Av6aVnw4Kh4b
yaPM2LkdEMPwX1nZ54lcjdt9YoWefFnedL7NrpZz0I4FT59Js+tt9DPrQyCtbRP0
JqYSHQMrvtWqZZEtXPP2nIsbY9Kq1TjgyOcYSSREtcoKbrhqpK4aWSkEoyTLREPD
ykTLoJLUTQdtA4dr4DRNpgZhqB9DjsSJ1VjR+rshntWXPTi4wYuS0Vp56yrLt8bU
e01W732FHDZMOb77jAyZ5BFKuOiLS9uAZkU0UIv1CrI1QCMMTOxeNVIO53jOqPp8
0ROZOFBvI8McrlFkzgqXdZAdybYmZEV9W432lRmvubAC6XSc/1TQotpwCDGydaYb
ylO0uNCTdXs+zKmv6mQtPsEsOKOe4tJtdII5FZ+95eOAtQ2TttRuK4T9OdaW/iHc
l1B7FB4F/X+XmrdDva/21GGFtZKC6dEgOWabJAmxye8LRZkNgElnXRpvDyP773C9
aSZqRYjmQ3qr48KZqUrRmO0/RUjUU+97eB19fvVGZh8LMn9TL4ofAk0YGn/nMcP+
tjoFF66fi9vBHYvBB4hkEwFXb9KX6pcLmFtGx99RiXRNZmGrTxnuICqVeu1+nQ4c
39rBbEWi/y3GkX52IZrQK4WhMEv6um57BG8xwOk88tsTNY9bfp7+gpgEetDq91kU
oxUBEl4exXu9KxKzhMWajeFJQK8aPm97cxUsIs0OT0/75e+o8dgtUACqNbBIXyaA
1vYkUwqpE2zFGKR87RzsTUHeZgxuKdkirBkBtu9bvKMBxHilYqOrN3jWrTVjM064
prgnC1W30v5uf9CJnE2gQ8LEq7nVE87WezwS1hka0LQ4xHgDdSt/hEuV2cVxiGtE
vrKeSszDOdNPMbzvdFYjkaRt6ZdIQR8sJsWU3KmXjKoBOjZB5NQYpX40YvmWWtpV
ThDA9miSYnyaEBa1yHZUYaLosTVgtdgRm04Tcb3jjvj0BUuJkTU6UfNlsXLGC4og
ZvibHDoV8XjnndS8CxSaF4uReBgpmH3cUDz75UFUao0f2e7p2GjxiwDRasAI/AwX
uwQBydQEzpE4YVAs3yR+6nt12kYB4/izolNa/BOG/3PqhakuAl/cSlKz9aLu6+bz
DNS1FN99HHrhEwqHMa54YQKWPbSHbQD0hpl1JmVAF7UCkdClFeUy0xcJCYe4sKtX
VRPrhxRrQACgbR7XEO0NTA7xXkl8TBpY0sPLyTbhnFohA+Robltv0yqx+rb//Zhr
pCRKjPWUeEHv7e43bLxyDTsNFm2Rfysyc1H91kutNY/Gu8PVNijTWIbxmms0q9Qg
bx6iUqII3EsC88moU+ACouxYlBRun3SLVLe1M/dCvcAxHzVwhN32jq4nLDkAIFK7
FD8VCFqS7NhNSmpuJGsTXvNfmIALffPvo0iXzhPQZE44sPmQjNX/t123OutxLVFz
ePh13EqZmwjHSF8q00PXOrnOzeFipy2hQ84xrM5tpApap1jV/dQ975YClBva8+WL
im6SPFhDinB6oR++Gesfmx6VOOzgwpAXs3BnpkJC0rj6wCts00T3tNi2ya11esR1
sjflYfCmmCEg1Z8DqWrm+Ase2r20awcyHXeb4MjHNB5yvEVll5qBxsHg35/zSa2R
TzQgqChLKBGS4LckMEA/vevnEo7PIqYk2tqSpVkTAGSHb8Pc2B+zC8M6MVrS71oc
1JqjTUZuBBObQmUDUb7MIEZ5GtqHBck+Ha9k9PUHPx+VHehK3R7yvEFkhldyhpom
zBrufP0JtRZbMyw1D59gWxLvELfHtICqCSTIz2kLlDWqtwVcP2JTfuxD3XvMIHNm
VGDO8S9x+ISryyecy/NqS124zPVtxDqR6a2CqqDBOnYBcT6/wFooAUo3eBzPdZfn
eNihXW+mDNW+WaWZz1TmF+sdTmmrD8yAFzOH+vSGPIgNknak+5NNw16G2GxqM2/+
HNm1sy1Xwu2P9pjgRflhPuenJlvwIRWkRnecg2s0pUPrEs7EtWHP4mIZ/SqV846f
O55QxBqrBIVpWFyi0157Agj3wlaHFRb7bQgGpGrd6v0ZjYmqTQ5vvqMt8f0J3qrK
S6Hgye4IYFdzUDooUpUOJsYc+rgWUJh6CbZYaRTtWpIzvLxEqsREnxaf8jw4EW1T
AKcv3HzVqv+7nSleTrT8uGHz9KTOsvnODOO9/7meBVWsML1LPBGLFeL4GsEU7ZUp
aYsmYkAXmQNtVe1C5H4pAHhNhHkPXWNwAyMDgdzn/L0miwilUECaCGi0yS03gUi1
qBVRdd4agwkxB+ZtjCQbQehsfmRnwpUqBIVgRYdWrci6sEd3Bon1+EutLKyPpuH9
m3Zn6CZtuialDQE1zXpVeG1WuyZkIZiipdMQK6h7KW3zMQF22lQLIzQhJ+htqCKh
PAB6B9R7toemZzzu3IrHLTzjhqF5Jrokl082UQUHL9YcmUhrlogrowwVoHNeNh2b
hjn5gcuQQ+Mb9oQg1U7UQSdWa3Ff8kSzuJYO6QWsvyKG9Rfh4dTV8xm/SxNHw5l7
PrqsRys/R9HVGKcofeTZTGpx1ezLJCyXqOKBceiHSGQQif3SsPgBRdAik2VjaXZx
9HE/C00jGMNdCntJPxL85IS2DYsVIV9xizwGxtPsSr487MvZ5Qhis5YtzGi2IiUz
KqZEFERuHwCt2R++iLjXiVkeqegq18lqRygrnYFphkZeSCbWWHFuOMdyg2mRT3Gf
xLPhWIMs1nIjkn3avhQxnzneLVdXoq2hfRiYgeLrcEPuxKp1eH9Wef3Xc5gSTyWc
vXwOjJSzzGarj/1OqWdcV6l9UHAbPlV7WFfukGW0Is4RIVjuUS3mAIUOzExhX4WF
qKgdzix6NUAYpPbM4orUHhT//TAwgzfBdOkZeLvabZB5R6ubXGVtNrH2yOQu7Okt
kwTpVzdhYSNMVd7i1lAMRo7djEdGq92MRe9oIjdVvePDVbtEuQeYxWwM7RDQoBIO
mB5aTZQSxuWbyYNtZI3PaVfGZdO0mzOa7nWqf31GZSC0nrJkGoq1NNBTuwtlMPvF
IpBd6EYDcpOBMkG8ZRNx04Lninj+pqP43Dpwk8oVTXiuhNONHd8BusAcc6onoWRH
P+t9mcpub262eMr9pQY4YsmZBbyQntfUcFr8/WTHqDWkqKzqyma26R8A/msXxoOu
J4QI2rD+wcvUo8FY2ylEyt2dFSVReaYEe46nz36JRW565w6PZ1i68B7HyRD9fc+m
mWgIsXVlrE/ovhLnS0+47rzSME9I0GIZuMqskDr+bk/vHSoOGobPpTOfoM/EPcO9
hC/mmSQoOSM5BRhyDvxLH3/+zsA0pYIUFZfJb+7ahZ4c5e0Jbi6NRaVbqYLC053g
0duDTi5GVhrjCAT0Q8upX3gSg7/3aiTdWo0+WHt6TjQRAdE2nXIcwEY/6fSRiytA
P11iYWwXU4emWYQrqwZmLlLsXXgE13La/1XY3KOC+cFTJge1QRt5ONbBJxTnE0q1
bUgGIWccXFPnjCrMYCa1f/ygrsben1nI2DakPb2xqanBSAjHraow7AXlLk115NLd
Jp/r+ryULtsyQtZEVY7Z5dUVXBsYUliQTOTXj09z99+0QLsu42Bedap4OrTDB/hz
pxUpTVR7SHmzDEBTxrONFBGwX0xYxZbUBroLzkUR/2ZMDpuq2zhbT/eOLe/jNce/
KjXCNZDWNzjF2aTU1SG4AK/wG63RJG7iTrd7F5R81G+RhvEkWX7UBrx+PyVDVBsz
/0gzGaI/3jfcYdeS0EkCpdIaDH+46LWvcoyJFHsb8nYuo3mcgxYAoF5UWP8XhRa9
Va5LDtHPp7n7/C+0vG2lcZXiEUCA/TyphvJ0QFR0K+b8RF4YgkdZ8gEciAkf7Yrw
C83/UIflpYOqWpN9s/bWC4+GkDHv7z5kkUZsf+EvLOFmh7jL6bQAqMHOa9G352Rk
ASxquqgYOO4MUHgz3ztckBuQt+x4PZi/5l9yAovabnNwmKvYOytO0BIQK/eAle3g
bNHaCn4ENYatZrdvdFoTFkHiJEHFTMV/DxXKytevPjF3w3is+R6Ot70gvDsRamLb
fekPkbc1t9EIM3fqtKU8KG4kkOTo/amWeqJFLBJpYENeQ+TfgtBM92lTtC9DIWad
BwmlDsOFCnxNa6R9UBp+oFjAGB+WTAab0A+oXKL2xgCvIIneIlKn8GP1paIev0Lf
3XwXbnVlkReFHSib22p8/LTt5E2YvvCEw16pm5+N22rDnLN0x6XdlgNVMwFJ6Wkm
zUejJloEKKWk1FpfeHpuVgOo0rwHrrEWDRA195VDjIaBp9TV7id/1rW6LYzrzw7t
6imJlupyL0kjTFxVlZq7xbHT7FfHZ7ixPWdregJGjjRZzjhvtU0cIsWUjMbRyTxc
dBuQE/Ycf1A4JfCXi0WHAagYiCZF3pBfoQEwHy08ql/CJKgMyujnZdWidZO9CWzh
52D/wNwavpsmeq1QJz0xhty+D0nY6f45zswnFp/iXzK3d4M6m5RS0n+RbBCXLwXq
mjC6Zm7e8j1VYdVeyz7ACHJGJB7858XhQd18Aw0VtHUPZCkH5WCfKoGOfazOIgnE
C8ndfkBBvv9Iha2pB3Inrl6jhWoPbbcme9Q4mIe/IKBGdwAGX+Txu40gEl6YsvG4
34pV4r3zrnSpN0VhY424rwD/g1v3uoxsJ8epxc+hKVLzWOaijIRrxudVnxjP0YQ9
xK5IG8t/IbA56Kte/QhRdRONOBAif5Qn7ddy5DtUNJOYc3kcDzM3sOK0FzTaTotM
Xhbu18Lg54YU+Sa4I1uboEBu07CA1AomhA7ACEkZEB22fP0EwEkmINFZ3g6KRSCk
n6HcArjP3tl7o/0wuvT63E66E4/F+zmGJg6cyGAY98rR9G1zXv7sD/Sk+UwcDzdI
XyAdIHYo6Vz+EGUQoElXDn2yzofTLVqfY/HY01x1wFuAX5snTCVk3xz1FhVBsAus
MSZhctYFXIvU+ESwOHqt3xLWLN8/yLx6j/mtLoIQJjNRI6IinM1p2hJSLe6PsFZN
bW3ranpRujC08MBqq2E7udXhYshb6RDZvrMX3TsGL7yuj7I/sH6X42Hx5BUyFoy9
18rVWYUubt+ZM4la/5OjL8EDmNyEEkKiVzRpNNI5fy+uGZ48j1m4uhuWekPWS0lh
2C9p2cH6J4YdUr0chvFUaOAnavbOYmzPHXFX7yiV5KCVX7iTzPl6Wgl10cyW2P4y
4UKuco0GDleiXY8Yc7GnAWd3RXHUOC7Pa02Xfemu/TiLvVCzsLPwKfYfIKvbnCv2
rYN8nBAmxT34nhMgm+m5nZmbi2Bzin+84HF8e0vZSCCZpzP++AvxLp1GtgpJFePd
zBaDUsYExTq2v2gpSebo7pWWcUNufsjMQQp+6NvZrk4/qi/z/zNICjvCGh6eS5AZ
O47MAlQv7pqxTuwhIlqjiQX7r6w8+NQBu4Wl3I2PtCrndSazqSPiMLKGrtai/6tf
ekoABkTAYXvi7d0XLe6qXYMnrSVz+uGwvE8Oma5dPKako/t/1pGP6RG7prCYDTk8
v1NSlsODDRQ6vhM6O6S0KJXyXbiP1nhEn8WNsv1znVrg7pEINi2AvIjnGNyRN2SE
ujbTolTczMBBjvzrsd63lJefU9B8A/GSyPJPLRJy11ci+MBBQxOepV4f89exKKfU
Ij3O6r+I/lFZen8YZVU3TS31z7Ru3Q8rcLC7+9xkqcDCYu4gFGKi5DV2sBCjeG12
DqMO29dmPRjlOJzISaiql/kxU0LvfCh6Dkwb92eaxUEW9wFXhYtj6bi8uL12fGH5
ifaiK6qcPYkreu2t6HGRXUPg3UM4S9uKGtocLcfFdXFWHN6EYr+MpwK7FfeFaLjS
8dRRX6LYKEQYBeYRrhZG50ZVYh9h2cI++i8JZvQ3YWJsICXTJxBq5sWHFkXikes7
fiaWxPPql2IsQ4iccX4DoTg3gbxgnB9wwc+A6qJTGg/Cz+g8J0CSMeP4T1BRtrut
IP/uULVNKI/Oo5rLpf01gbooxfZwSu5UtL1HqHYZVpGjdlwF97P74XuCrygYdOt1
63T9oy40eXJQAsCnUELD13N7NmxpQ9yEvzfz5KqnvFBEndDc479hUCyGZ1NqZq4U
WtPGRKSlhfxEqyRiKVGEC3EpT+25P6wck88nFXhoNILKFrXG2u6/qoLXJeVLcCrT
7daejYKX1BMzEcNcM+wk/b1MUjU9MycHbsSA9n+kSNxBq5bNA8TghB8qKpeo8dYi
x0BE5p+Sr5jXDOgrUZxC37mx/Wjq3ATmBcxDSc/kx0bx2oY9sjlRfpinZF1MmfyS
U2xjKKlm6LmXCMuAitB/IrpQis0oco8uw539ixU2vlFKV9oDaMa55/w+QuS5ghaS
lM2yU7QcuEjAs4V4WU0vrTZKHXySjCBMMknNWViQLR3CfxLFbjy2BkKZiMsXLo4u
18ZFAwwZMXzSyR7Y+3p083xM9bwpXmkwJ9r4P4VvYY6TSGu3PuaLQVBFF2ngoaVk
QEUJYJKNkoT0rNflsvGoRw31TSNYevuWmgbSRWILSpN6kt0/vxr8chyPJCLOao+H
YSF/LXfpOq6LeyRdeS2UYca9tuMsLGdCIqhvcTFcQl+0NdW9OmhZuzkj1P3CNN+g
wvJVs/R2WX61jrwWdlTusXAaWCOw0s+3qWPAtiKX2ga+Rus+SabRj6ki/oP4A/mF
sE8hO8BPh7gzQVzr/WRIydfPRbiFcgtycCEOmD++VMLJ1f3Nc1MCgG3PGKHVM9qQ
NBc6zIuCT/APlFnBrIOdcg8fvgTQhpWjMXP6SWXKdNGcngP0gSxAG+DKNJH654uP
KGIk9p0oWtITwnRKiHs0ieseYEGKvklIMHn9GVsYzRdgM2OW2cFn35rb/RCI92M0
VTff1TYYjZ0mzZkmfK2huxmQSHgh7djh0cACsXLFiaRLPwVv7WUsok0rA/zenl5C
so0oUHaI037u/JsoWU1U70SpnV4sm2MHtO10LJ92wBe7EV378l2duCLDNp+xKRc5
IqC0s5m7D13IqqyuHjkE9oK9F8L6/zNSpUnLR+McaBeMErlCgihsq7lUzzvM2ESz
iEse4RG/Z6w+uCdXss+pC+MKb5jX9CS6+LB4G18tGmQfpFJZ/FFx3m9FUd3XT9mS
soM5hdFJnU4x+3FgagQGJziogmPTPmJVBBhgNpOqeIZImUr11XhrVf5M0agFz0+R
lbhQXI55v6zYuwXsSTXdNEPWXA4LMTPmF9H+3DkysKoFw0PO9ja+mLQ3ffLBOrZc
XQo2/7H3rz8vhUesvz9IKLrRTpnftiBCp7jb/GOhuMLCT4HX8y2vBKeKrX2ovOHa
5fBdwY9I+2TaC/FSdzpHqhRE4vagNBGOr+SNDYoN7zZq9hEzxvAUKVmlPPffZzQf
5Xnzhb+/59t7M8UZKz0nilZSORTe6cODCQnMPojwdglg6XVR5AdMJ0GyeHwIogKl
DmJ8SEZuwBFcr2EzFH5+Qb2t6V14/BkVjDZOhIbgJBo2dx6Q8O96YdNdjY7Xyr5a
No7SbzHBwnjDDBWkLNV/ErVy7M3nNFcQzK6JaXsVgY9OuDoQS3X+d9raKTzz2Hu1
SItjhlvD6XaC0g21AozDrkIe5zV7fU+DYOXvACtPHTBgmulz/uzler0q4V/lW3m0
nHXWmSfHYXVy3WkGDYe7IGML772wsC6n8SRy/ljmuSMmAHDGcZ26t/XIJL0zwhr1
14PiZARwLuEW2um7eQDPXvk0t9hlHbv0b8ZPeEItkeGhPlld1bcRHSUZvgqi0J/O
FrkwLzgf2YRb0IJRYzdtKFvaqkQfna4HRINjwDavCGw1TP+1x5fSkm1LFS2bmAa+
kP+43BD2KGn5iGRbDghmjSmM+JvL3LqjXbQXs3s+G3AeWO422n2a9jaUsSH5UvAr
765fRFjxh+4qWjHtvNX5OGzrN27WLa03z/keGgKzTsV9lSjhxZ0HnQEeOhTlk5Eq
80s+yNEkc3jvJ0pr6dGylb1VWdpi3RXmr7ND+zvs8InOXBQ+sm4u2qy7Ove1SgZe
Fk3yV9xgprH3D/Zb+6i3GwnP0fCyYBAWHHNtUYFr+dUeezZnhBscfDTu4Io2AXQ/
usS5GRafzi0kiZaI2TXTiCV5HMVJXJQrxxleQIF5blQioSK5u/HipKBtr8hjTQkF
9YnLpP8whw8UIaJ52bLy/BfvQdRFIr6Ld+wNealtTVKb9LWASC9V28pi9TwCb8B5
kkvKr9CozxQZ5NDseaX8BDMBYe86QpgOY/6GgqGxK9TPWEwDZVpnH3Yd/YAyeTCi
YOnRdMGiKopcj4UbhMd6PCMDQpgFOAU/ahjWRaXEgPnhm3YZybkOJcyVltosquNR
MlOE2O/MWNuND8udYjtYCEeuv0FaRZO0/wIJeUZ/UCj0F9ph3tYKypkONXcu58mc
N7v69hLb3rgAoSQ4o9ZV9pTknsPsnQxjM14gSD7osDy7jwNL167KtVX1gmCmqqnT
1G+RGkkGsIZ+Qmvbkk9dwT7q5xpiCpol07p2emPqrS4so0l235fFhFTpHcu/w68z
Ts7d44m/cfS+dv4qNy5Fon6F79P586U8PCDidJK0I2tVNl6KwJ+s01Y6AeOOm50p
5SV8g865b+YE4py9hfGej2c1TcS+iI0kexSdfZpAkkT8V9A5FR1i4CE1xvs/stAh
3VTgTXrfCh+4QiFWlkpLvCU+asmbgQ76V8hQwcWEkC/g0gNWr0hkTpVs4PRGGf3t
K/uX215fMIcCg2AnWywpFxjrgTY0oH1VoydigMivtuF7NZKIkRDUIm4Rqayl2eCL
Vh5C84veCh+AmR+fKC2Z+zqLGRK5faHnaiKTc5F4T2UNenizqXQu3M6ixnZw9E8B
PoAPBpZVkghKvXlsRKSOjxMa+wI7UGkiAaUV1bVJ9QJ/G+czyEaC312z3WvEjZVK
3cjGCq1Jeh6KbHNRu5cfcMvcHVnrT4e5UtK8h+9pM/X5aucz6nmMt7aB+W/L2A6K
YECl+93NrHxJaBrIDS3Y9RAIDPJCCzUuoGNKhVKOsNbImsTJnlTUjQ57SZ1uaCtF
Cn66BxqT6skgZrXEcskX8v1MfGa5bO//CAEb256K/6wlsSD3uwGfd9SSSaputWps
GeDJswDEbCnzD52GhW1H1pgVwCVk8WZzMWDPVWCFw+w/0S/XuKeX+Z36A2xREa/I
2TFEmR9ebsbZwGJvWFICrxgMAZWHITmP8VT3NvirGJV1jIzyRjPEaA2lcfkvLhYa
6MRHDJJIfhAIQel8e/zHFDYuy5stXsrV+wjw0kMw227XGeF61LXZwAjvbqommFft
qTFqbnmCRJgKe1IH7HaFwohTmoyzwPkEmb3qxxvAaAeQ7CzRmqOhTaySJU4b3FZ/
tPrEGUwI1KAtjqSYqIVuh9dI/lxwDAxQQwnHCGvZLcYta7vBtq09B/6neFReBj+9
Zo9qBoGVuN35grQNLfeidS0tVvMKXInZ2nZYmHqhf6XMmMHqUnSMfdqYcIXzYGOY
z+oCsLpvu4Fe05tRKAZYXh3CpzYgvpa6CLmcCym/JNoe2zhc51nOyty28OVgMakW
WIFlK4FG930X2a+jJej0DCSGkCXMRpxi9K0ltoeVeO8/GHHCsHizyObjM7zrzVJo
z9vEkCY4rTSSAJi5JTD0Y5d+SesZv7ckTkx1XXCirMgXUeBPgqWWUiP/Ae+Y9/IG
4REQl7FQidtSL4++nSesaMSvW3Z4lUa5UGNmbT8SsHHUw2QXCfWZsDnz+eG7P1I/
2AdCC26n7f3S0epg5Xn+RR1f6ngf3E3w/erK0r85yJQ7bv/hgt6Voz3+nxRNqx+n
+Siaegb+zrRF8R3mYfY2fD6+Go9gKexzqENkaLX0IQDcplYggsk1PF3PRVB1M3w1
ejwu6l4QUzaB0DekM1vRQ/wh04Rw4rvHzSfGTO4NHpKLVtLDAVWoc02Y8WV6SuOz
35USsiRDcZASJ47Qb9PPap/HcJyjca9jaSYQozSIKKW5g9lc8Wfh1+OHMqFmcV1W
Gp0cgDSQMR6smtqRlI14HZ3Lcsb0Hcvaojvp9eeZX8/2S7sVmODh00qa7MKquCPw
5RAfGOGOGMtVyXWNJjkRGgQjd5cPfy6fSiDdlajBJ1oJnVtz0L17i6YopIx45QGd
uexZ1Volnqhzi8ugerjY2Q47GzTfLSl84OlLMHn8IHKL7+gvKQUUYMl1ejsf29Tn
BHAGZ1/byqkbwUM2/6wOp1BPClIj3dbv/rcAoVm3wmbTeA2glQNEDYFjPlr34EP/
MPHL6a+uAiChCBIJRLggZ6QSlB+vg6oL5oE6eZPwrnqiYNsMKETHsY89UqtnRGAA
G4truP7iR3M0T4zPeXlzfprL1VyKEnF5Qz1zpbGcmW0iXQuuLqEPdInuShKNWuQv
YcIJ5IibpxY9mUAjrmmo+pwKJP4pkdUzHGJN7IQdtMYimsFvQy+MHOvkKePjl/ta
UnlXqqYdZtANt41+JPc2F08K6Rcb7/i2U1vF/dVTdOSm3RbISFwh0i2UhgEPqKpC
286L5B1TABP70hd2TLSuwqs47h/2mBN63lntlr5TGbnYjIYyX3Dz7fkGeRs3Dr9c
9waGk5KhayPCrD4fxLOReIN719LbC3hJIU18Ud/5rFvBwWpj7eanMB+A9N/JSd49
MWA8NPCathnxbnH5epB910awAEL/RYdvujN8GfGcQq91CAsh7KiynQkGwVTdkx39
thQtJay2wQvYMGq4wmJbdlttlplKWIwlnq0wJrkOWloFgDs2JKxeSr3uiPYH6wdY
oGNfzO5vrokzFcfIz4Ky5D6/vf953QenRtXl0K/BvCug8VZo9aWeTM8z7SU0rBaT
PsmTVQUjdRZhwj4xCCWOiMrRHfAUPX3grwKdSyCt5IQ7HUJ8KAMtfy9/TCDdtUmJ
2vwQL279krL5E/u4etEkN5FTZzyDuX/nH+0RzOqu05VMuf4HCdgDKQZPTtcfwSQO
M4+0KBa/zN3YkyjM0uAnnoS2fnbS6Exlo1SD1K8K3ucIN10Hw9DwQM49JciJuqOm
mpSkcVYtOUEu3NcV30fmuwQ2DkMJf6m0evwtsbfgoqbeqEByQ2jvIG2dZvMYx3F8
Ise0843Q7zTZ3440a2oa9bGwLlgh25zDwgHJbKJS1WVWRS1g6/Qikqt5Jj9yPGEM
yrxlAYZibU08xNnGS0jatU/A0lwAIl0nYOybdgvTOI+RAs2nHQqrWdtGqABq0cpw
LbvsyIbMcnWcBCtd7exuaCUP2Fj3IztVym18R9LnDRg8alCxDsVkg2qZpoAOfuSy
S9mRMAAL7OfaEgN1E6XLpv0fSHKOLVZAMpbMv+GpI0a8DIuaVRka+mn9rI1e28bV
9Tg5fLka2slSCCclM29RLbFWqpgcN3XZdoOe/76sZMK0fkfJM8vWfM/B0cFACzLz
sxVPCoQAkybzXNRlMoTKVn72l9ng/IDcYuZ5FqFRim6J3XhUFaTeEouq+o6BFrzG
E4tK+2aBDHRVk9K0IoKKJyLTAYoRfylq0k7j2LuYfh5DNfR0l1rX6baV5Foq6DEl
tSmMgoeXEDryZJwaeuxXhsrATbfXqUJ2YjvBzsSiHr4ZK9C/JfuKtVzz90shMUjQ
Sf4AFeLTK4D1TsHhKN5Vp9iohCjBxPNTMpWa/SzO0OhG/L62YXfE0u7JGcNeSrzi
77adMecte2rUX3FYIMRRblxmkbMG9SlerM/GuLZtgqJEVlwWJrC/pBxpGEcgRURo
Ub8geL2clbtGpp7crTUUZLe7gHIMtcZMNTzSHSnPnoTaDVrNuNXOOJll7imHbKF0
K7a5X01+uc6msB1dq8YMZKEpdZPYOX/nT/I4yIMPH6OoFYLGvS8OOtgEqHMp40WE
REDUZMVRac5DWfQchGpTstNL4k7kkIxX3FpXR0bUXWIPBhNqi1osGaUjjNtoHcJn
o58A4f5KBaDitlBBTx0NigwRwdIOkKoYPIMsndMTiDBhiswXU8jmxJYpgua2zUOH
Uo+FR64/5agt70TfvkfGOB0O1mCHsbS08Pn3832aWONSGHKqHz0qWc+Y3W3t/Khq
Rwotm/YBwbahV1PgG3IW9+coy2NQK4fF5Sl2cE5bQthp2o5ZTspgA8/C1HbYvLf4
5AjDvqedgSvAcmiaLgt+cmwSraOuu5+Xw9Frs00eTFubQVRHDGc1Azz04X6SoJYx
Zxr4dxJeDYdeDm0SUa4C2mMtvrh3/ODQrCrTSd+CxH1numPKGSq+oxdMf413mhzj
Ca4wuzvq6D6q/UIevdDmQLBFnPyADfwfcXRE+E1xwo1yv8DGyhI5JiZnaIs7RxcZ
YmCFYFvQBPupN+Nnqyv9wS6JpeQM9oIXaF1JaZktDJtkNq37ohzD5Rek7DFWTOa2
ZvFnsP61txIPR5z181+mtzEb5ZKsKb9auE3DRBiwIsAV62HopuobqzpagWxaLIT7
2alMzzrIwp2YriwUCbgHSzgAooJcN5Z3gqxK/KsDQ+IqY1o5Ub+kZ2LWdVEvnFdi
b/UGOZttSKGNSNmvq4BS31/P3DqTAjRrJdf9fC7fkq4slumNuMk0G2bXRtZSWk8f
I33mRKbGNX8qQU/oHj5g5Yte9BoLf+MH7GDBf6+jqzLBnwPf/7AWUSm+AX957Rh4
PtYqGMfzCu+kqMbWq71wVjQaXGgPkls7IE3dTxq7CgAlB/ZRUmyH+iS6rFPauXrs
euiOnCOlTa7Thd9TqcP8rHn2vJod6IyyQav9OVfDQ0jy4D/i4RbribE2aoopgEhJ
9e2oY/u4MktUPkh6zl17Tg+0F4y712IXTb/DLUdpvaWZuXWRrGHWm5uEbYaAK81N
GMhppupCztNowBkKMD/arK9XUMl42ChHxA0C/9Cym5/NPVw1VI+SI5wsg9C9iU+C
yT75bIWX5yrbqWCxFIbNUzjGTVhTcRtkmZ72MVOOn7UWDvw9KFeiGoRzruZCJr1p
eaw7EfeRVmNQZqZhEotpuGGS++fvSf8fddPqW86p6UhgI2T16ZOjM/PnnXk4Yh/A
xJRvqVvSZJdmfjy8wId98CSw2wlvO7mh9f9ebGoYAinbRB4sQnE1L8/yMRLoQIlc
DCDSlxFzKNEzgajHloOw39WvxpTtWQkc6PuPMIgpUASPBxXrZ1/xHVOe55TuUwkQ
bhUBzia/4osR8M1xCTFd/0VUhaJ7dmPpDMDFjB9MRzH55P/Cu9EAJP+Lvk86yvJP
0i0Is+n1WGyaQR9nLgmu1OeNxYCooy6CP5Gg1mnEcePwDoP4UG+eo8qEIaTuDkld
GIqE4a/yXYjJmcwGxv1+WTpPeHXuCgSHRnDlmg8rvyr4osbyBxC8bn1TP6VZASiH
bcUC8Ox2pnD9yC5E7KsrwN9jO2JxJ4BmkGS1hlTlojUmUNhps7yvob2vkyFnf8dS
7muo4NWEQ61bBS4zen2jE7+Al0YgeXtH/8vgufR5PRkvTaysmnvOPQ++/2qyIw4m
P9eiYY9QZLpJdSK80FQowpnpIBoi4JQUuvuBG928X0Y4liwUZKLnp05x4Xrmpy00
2eG9GNrGYdmTdZY6+Z9f1V2XpTIgb37HfQpa97tTUjkcluY6dzeSfc64pDFNoBTy
/IQkI+E1yOdCUwbV3bF58uUrfxuWXpNCz5IX08SU/DltBoYx0KguY+7u3uLDMwA8
4iXvHaFTKUcXkSnxKYDvwAUixVsQhR8DXka/XWJaGSicyzATcXPY4lh5BugAI+F7
lufPM6OHaEpMUhqGk4tpD/+hmQuuh7EL8noLgDL7Yic6QJx2Biqj1umgizSoCby7
x/aFMDGZxSGeqIWnBy3kGCQNAItwfrTRG9ZXbO2iQNRJRQG5KsjbGHcsBmetLQ3H
X04dnNIaMm8mIPexDpzeZ4XJqlIguX1naLleuy4jeePi6Uzb/CoG9wwo7sXrfEuE
aZ7v9dG4YqeoGqFW9DlkKcR3Qbtwsf4GoCEaqcDRRYkvN+w3vnkhdGnetrYeILCq
UtcBroBdcB5fAffe2PeV68KrsuUMVh0aZn4QEQrfV7PoK942Chdtb7xuZUZU5KQj
8ezkmVautFcYhYoXY+yPyMCv5F3AXyfMoTkD3stOWE/rWyBSbPQRNbvUjUzjHlwk
c2zC563h8wvUnPKuS+Vtb7q1FGGRlgHrE5QzKmuxxitKNUZKFEf2ZVJQXVWXY5lM
uSdS5N/rCz+GVzbW0SbB+WvTLQFRlPnguliwsBkSmXCGrX5zYN0DYUeaGwGPgD+N
ssZg/mhtpLPNawskh8bJYYvi0MOnKdZFE13Q6D810d7zBWdepdsfh30Q9Utg+ZJM
T84pRFaFTDcg64LNoXejCFdpIMNiWK4Er9mzjHrFWJ7I+aGMgmIzTBvayhirDF3g
EH2IN06pWur09Ewmi9CND4L8uBot8jxxM/ZKrOU6qzRIeT3tst249XDjT1DJ6iyK
Towiw2uDOnBAI1VJ1zZ2VuZJcuSM9AXmCrZhk9eMfehjIPQjuWgh9gSjQqsO3Aj1
5VrgVdqoGZh5ipIDCYPjGlEK+drl35UNCm1iA3wPHmRiJUkwkyUxbhRtUG1UuW3f
2YaEuc63R8FoeGV/flmgTC7LbWKekTb7/I42dR3m0jWLZ2CvbljDsLwuHiUYEbJj
i68Rzulp4RUxVooPeh1gxtx8vMZvEb9kCQ6LNUj+QcQM1DoGaZNEv7Gj7W+m42tn
bG7fXPOYAALNRWp+FHShQNkhLrR96xzJ89Jnxrnk9L9rdTewNGp48rXLi3qrbD7K
onSA15RHTNDOuYkBUePJYzFEExvGlCYcC9CV3ktE+fviVnVM70YaB5VKm5JJm4k1
leLxzlHrUg5xx7GwtUW2A7zXXOs+fuQ4ntx+FORLAPOoXNUusojKfb0ejxMgsmOl
xIxnFdWSiTd8t2OAGKj7diyJuhvOHx55K8rRYxRCoKn9e8RspG3Sq+EviJ7HRE4k
Qh1gwzBJPVlQ2z19Pz08korB56xnA/26CKB7MpPNT5ZwraDR22gg/V9xPd2e7M9e
V12bVYJ4R0SXKivryD8UBK36GPJZxGrDPnd8/T97dZdvt05oDjKaJCbO7RWccW8y
oLoq1THBvw3DHzJnly9YD85cjLDt69G278EwrG0vp9NUaDG/BqOneO7pwhUyr4Qi
3zbhEQ3F5iYE3hoceXgd/6vVtW+Rr3NiqBkvgNBLK6fcdNjpbvvQSwvGrzsX01Fo
mcAc0vlVonDbxyK4BKDzwPe/n/zknUFKbhFqgy08+aYbWnFAgAlA418XQ4/oXXzZ
S7p1Qanceuw6quDtV9NjwgkePnfChnvUnb66pNpCKeDqVpmk5n6u6FTpoyU8PCjZ
dCVo+L6ij2mOfYzw2BmWDoSJHJDWRaiZg8zIrVqBuwS5C2hYv1xOxtKJpKW8SRDo
zO3eerubcnDUR9+fTWm6tsXqPPA8HVFD+7l612NSeQ1JKrENc/wkvgQR+EowNOvB
wbyef1LbXGZ3Kv8DQNHGpmQ5juZqx45uVZEG5mOzDtnD2EtArpslvaTAddP27Z1b
jA1BMNr8HFqkMksaIftOoscSw49v9vxXobzAAbSSATTEccGu87ba/x1+Q1slfC+8
b495w6Tr6tS9h/le4HSfbjklxSNdRh5MkKlmS2pCc9N93EKP2jxMFfrVVygzTq1w
qpOibEuPpsVazfTEtpkU4eG2nbvzevABTjJIRt3RhLpHRMZkmofwwjS4Y4/AmCuE
U6dnlj5Z2gPpVRgZ4aQH2mFOsTJbM2Bdt4C9O5B0FLu0OtuAhj831EpqK57YwDJL
AxEQUKXEu6eFe30de5tkcB547lWfQ6W14+Zn2atJe4LwxrSf8eBi/wYudNrWwfSe
6ejuov8AyNEXuFTm2DMsZpd5KItCS3bxa9ky0+9CxvyqiHgo3HiMGepFexo5fSXh
G9qAiEmHbBvhkEoYTi7nU5p479OMlVBaivzcJKJ78tp9b+GSVMkzS0MtlyvbRQmb
ZdKGXr0zOFwiKf4TVOb6ANdahAdd0KmdOfLO4ghL0HrlzZn1LK0baeZFIW90QdB6
/s5TrJ4Z82o7AEsgpVZuOxIOu3lfPuflq+pya6uW0YzImywcM5ss6qf/uE6MVQ6S
qgqx7i3GhXvPpWg6sDJatk4biTVWRUn+8NYQD0KzyHel6vWlJleTaDRjImT4Whow
qZvFhvYbEFPEljEEpfqLA2pkznzIz4Nx28TLeukyhPsBTM2efgjDFWRb7C1tNV4P
odlKbDASuv5HNzO0QzBH4We+dUP0PoI93KVlgzsYUVGpXTkPM62wC9gmVF+qKSic
Vc3JtF2bYqrZSxmkzyIYZOMNqmLldWSDVFif4P5NjKCh+R5LczLG7BOYrTnQbMWm
h0nTZwuDvGJjGgn3Yo7dfbI4DZeF8F/aolxUMLJ1H97FFqpWEz+aEJmXEwx5lQFf
W1yo5AscKRHy36Gv7e1jfVaneU8UAm7GMiiuI6VzDuBroBbEGT5aBxY7C3GqGSWm
yZMsfibHYnBPeAF6zey5qFxBRHxVM4ZeBJ9/ZlSdzS21SMWy6bq2DzuAEI7lwb1H
CBabBkXPvL859foirXddCbc5f87E2latl/0W3OlPWk2UW2kjajZzo2YPl1PXetjS
BShOVldlWjd6p01U8Ji/G7PBV4i6JWGOh1b5kizECqXvvgPfwPOefJmsAKOk14+V
kfgwdkdybqLlGG3/jYZEpWL0QEyIldTPzuddV/gymD3oVYX7KV4FNzx1u9ynE62l
cy6xd+w20fpTFVbNjJZ8hE9qovFvuA8LcjFgpoIbEwcvKgGehVd6KsW2cQUff+0Q
/r7FgoxXPirLYd0a2yOPJtryIrNAp/S1SMd1XzfPuj9hgMUNA2UNL3Up89pchjC/
rfG/32ZXCPZdV1VCx+h4CouNb1yMecWLMR3YAna7wRCCn7KJtfAyx+eSCb2Npy1Q
as3ucCK0Ab2bWGwEBbYQA9N0iVU8P+hTMlvXA3VADDI2M2uu/O51MlJLfm4JK7Zi
URs1y8UrHAGCXDs7jv9SFbdOzTTyiD881dn/3TCnWgDp4vs7dcPKX3wgG4Jqmgiz
b/73kVoyytMreyVFEX7hbXCFnxMw0J5kYuQi70PplcKf1KhcfllOxWmOoSTThskT
CNylXxu3JnNAL3W96f/6bSmnM5aW+TEYHGeC85jUQEirwQsjrTEE7eO8dFAdzaXi
0aKk2y5icr7xrHFPGxx0+UcBI3acwcM3HpTW5cpmkONPCtPo6GSl/5vFbabwEx95
GHpp2GV4Dg7kcQ/U4fW8gcW57k4A5ziBcSLSn2+KPgIkz9Ghqe/JVLqxNAKhdNym
wqW4GUPbi/iFZvFW6LC8UtNHwMJz8scHwvbUCr2r/a2RygGX1DZctU6AKjsiE4ns
Bh4ATo41wUBjIZdUmcQcjvRD5WQ4d24xg/oMTU6Slso2Yd8da3BlGeM0Gm02sEi4
Ubb1QOxbnDvgKwD1vti4yidvWG1dN58aHjNs3qy4PFzhsqBtTbJmRso7JgUv8zQU
XjmJvTNJL+xKCwaIGrmYemsIw9jVXyo6LsYOMNdw0WE37SeFn1o41WWYjafDorHx
r1hG8vL+q4V8XZUFwh4lkce9EUHBoni1iGmZ6u8XDxVde75VUKvsaA+xc/QLXNaj
gBbqxrapDafWJeYHce7EcamgLt0zXNlmFmfU9SNg0adZtEdkCG8wpm7HeAI2LJ72
S05eGCXT+DP7XdeQrijFEWvllRR7dleIT6/4P+cSCjsdplhNgPMLg6DD/8CVlq2I
jKPUU3jrrN/1xkcTGMmYcO6Ni3OXM1tHxa4axGMsyIx8QaxqCU5xLX8RV3Sx+i7k
yF5mWBrtcJob9xkPtVQKWdeQx6duNvntw8JKgNvtP8fWg0XYyHswGoX7Hoz54egg
6oZutI8RlJ1zWvm4lCDGay9MJ0GwExlrnJARriAqs+mA33ihkokFX83UvInmD4GT
8kJZ6ARquQi5uu4dRSVEtcYpLxgN5Va3scEXbARvC8D5Jcgq++b+cC4n7fpMXiTz
JLDVAeALGPeTAJUMVN/Dho575ehOiFxMvmjTKRfEdpVdh+w0t1qD2E2l4zXGtKjF
yfsLnyXx3KnWvpzF+AKrTr+mOi60fN+Yg/UuBDBW+DKpNChmKTGJKlZ467ennABP
2FumVUcaxKJ8GmbcuIei8mt9VROw71zvVk40wp0QH5NklvET9vG/XLjukNRku82y
bbmtfHbAJDKRNRoJCztHaXg6i+EhDopS+SQzdcMAeUcNipySJYZJxb5dSNkHHVyB
UkWJ/I0ia93UF05a3l/zB+YqkFnJmHsoNh6jNGE5WY/lNg9vPfKfW6O20A/IyRQM
8aWQ15B3TAqNpTh6ncrRGW+iTBtLouWKX9DlNNtQ4n3xcDVTpKEc7gkh+HnMQIHP
44ea6yfsqHavzV2GxCIw/94F36AiJ1lROLI6xl6nNGXf21ZNy7ntjB6Am2dfe0OZ
55Iy7KXhWG+xljbp4Km3ypJSz2QdeqsWGNL0Ig//wT0SNHKiaey4SyCXsUT+K9Bo
sFZEIfoOElYUMfs0iXnknblKZa9+n2ByVuEWzpkgw3xooNn0KXKJwjAL1RYBs1HN
IO5I24mpAQt5PzrgJ/zTe1od7eL1Vw9fKzQgQzNZSNSoDk9v0VrSAXQo8Dc3MlJP
nR58aYE+HdOp3nmhKVw1bhmiRhzjpVOD61/fR8SZEg58yAjoCSYzlIrIMERjoGwW
jSYvy/Nkm7Fftz9aTUt3uagDtZ+kWRaLppBS0D4prLIuZvI7aSp4kPnqyyN/fQ18
ovx/kH1aUNusDkG4DwrUoYrY8/kzB96lBO7IP5gOIUk4XwgJjggDKMl3GE6iRVSP
eEicMvaQPGq16ribfxJTi+4MhnMKhxYJWNhZsfAmzr8nO1EMzlL2XkBhgAajtQQu
8bFGCn2Rix36OEtCjazosmi+X7DWAhKekixGJbBgOybzRcZ83AORcmxCT1Fh8MDo
tfx+zlk9LH718/tbmVWAxgC6wsUsovODvl7Aj1qCgLPvNbQ/hNQInbr2T8iJHNON
wQPfLy6YE0Ft+gEU0uPOoTSrwyfUloqbFjWb9vGRKVQpOOufeEvjEG+K6m8YbUxD
ioQSMZJzGw8K1FwYtZDVDLOFwmuTjaMn/ldcz2S5nl89Pp7pxdJk9mdkmHnY7PM3
RXbuIt3hXf/yB8sXqgjbwFIgX/++rMLfc90iMRvl+cbE/Ql+RqyF+XmfSLvYNSMr
REvxEnyGJbtqgSjKlMxPM/7YWR1XAv9ZY5PO33zrzmCdKu10flz/DpcFRhZF1Ddc
9UIGbwtaWOkbFRbbd0+4PpJI74B57jJeBRFAS+hgTeQXZ474zgzz5xKBKnlFMrnk
SDr002gsBxCJLsJqcaDChbEL0TmR2vXK3YD/E97DA9i9IRFUGp3LI4lsqBL19eEX
s34zz0oJ3X6NJTNbRU95CIH95fmkCWjqn2TC22z6WwSY27NZfoLvNYVLjSAOM7oN
D13h63rPBOZV8I5YGE5wfOAZkgilBpyoFlidmkjUvbMVfx2dBFSDPpDzUEtyDUzI
/PleyOMjDRxqw4XVDCUnq/bvwqzObKDbOjVKeYAEVzPhGs1gTNx5Pb/cdVTSGeXB
css95SKJDONJ5jk1WFGRCl8XkHKIc76BHfC4JnJjjmspFBNSk+EQ/HRyYk5BBI90
yYNpGZE7CXvzzH2p3s6KRaiyeDjMF2GyNGUrWD/DF/WxH7i07VaJQmFdFuWzXORI
BRbbI7TjbokCEDiE3c03yiJOp1zIrzS3BOnmzWAue7FH+lrK7gQvoK2nL6W675Zh
SL1vrwjbIWSfs+iX3w0h/3Cx3f3yZfUqvJ8QYr7YRmuB1KwZLqSdxK1pftAp/ik2
vo/67dak3mjoJbrzLhv2gDnDOKsoLQkG52WggqUGMVW+t/Ae2xQTKGg7qDUuwLQ3
sMo9hsKdC7MIGXjRKADB/g2PVYXuORwQ/Grag+VN57nfwhCZ2s5cl7pGyngp9P+w
+7u3Hq9TTRWr4UXNjpP60GJXIbD6QNy7oX3/VvNlWPivGgyu6z/ipjo7ygWWrOGb
1UnLk+TsyVrx8pOuieZW+8Zy3kMlt2zIVqn8iz3RMy2lEs1ZwJtx7B+tpOZOXOP6
YL1lJyx01hRpryZzanOLPPS0SNG0veldT0YcesjupbEd3kbF1Ep5VSbJ/nieaOGW
3h/rqSftQoCeeYmN5hKYqDKYjYMq0LLgmvfiQFW0AkCu4JRozvIIOOE4XeoZh8Et
TwjjzVE5Ug+DHYBDrp/ginULEK3vKYnPwk1dk7XYlmVULQOxZg6XiKuNtpH+iYqH
RG0nHCSwt+nQ0J+sEAeByqA+IXkfGTdTXiMUI/zpRS2jKkIBR8T6XkKxXTRg76h6
QM6+8idEFPJCS3u+i2qR/US8Abd9uG+b9T5A3k2/w1c6R9L/J9JQy0QtE2kVplIq
mtLkgb+ttKpmHweJqBhKGiGtdkVytF9c1uyTn/+NrJXzeceedBKJe2CEE++Txyun
bj0SyeYSMXHIjtXl+OHnJ6EdmE3uU2hTPEkXCMxLkNo998R1DXM+RD5EK9B9Mzae
iyiu4JsZoDMF3CYB7sgAUTsGNWXdlQ4FJG+q1mh46kfOeghHwCpE+i8zHe8zxGJL
elt0anWiKN+Qf1Fqw/qZAarSn/0sOT/miiUSKRgug8CunqDwN+EQGA6ffrtGm0Z0
T85cfeQuyWloIYedWeiAFlB+EIpbgwAtHUHw3VqI+9F22dAvaO5/LmBq7cE30cCh
FEBlU5bTtc2VW65IbvN7Yht4aacaSGnCHUaNzmJbnf9t6atngDtiV8vmjai6Z04f
n7IiUtj+rZai8QAu4Od1pIGDhOM1o+lhqgNgSbTJnaift6eA9/4kQGIGldhluaFY
/52+JqxKOon1T5VRnen49hL0D46BQW5sVxyiLDypp3z/G07STj/qGtH2r3XABhia
/nD2Zux9hEhZTOEMptC3c26sThCE8hCDMv/zr1+TmW5lz/cv3A+MsXpUDX299JNs
PkAwXrndHKY5cTSEBIqdJJHC2kTKvZw4u0u58f/9JBhCZeIum1jd3mJS/0NFYsAt
H67Tu/c19gkHRzjqEObs/QOUZeSF0enTKV+3kV4ObsDyNzj3chKnIEF8X7RjVOMt
MhymUvK+9PfotieaqfrcbYvC4G43M/qO/tT3I5gRXeB5vOJ0BGnYCHNtO5U5Cf+u
8BEiK6nxPEuItOarEzV1jWgqBkoX1XOQaLTr6S+iOWNQNMqQXuyfTHaqp2jcEQW3
pFzQUdFTWxlMdVeH48zSMI8FdYQpLBZc4nSWwTN1ZqLvQDovfU1VAdbHSyVGT7eH
RzGkxVs81IzfHhfMSZogf6EFuFLtEZYt+pH5P8gFsBsiZu0fW8lMe6desMnLY3bV
vZ7RQAoqnJro81SVfEb2W1RCdLoxnjkcvTf90A4FPsWteWsdxgUwMFRyX8zoR34E
5soGjKWjohlzVNyd9m1j4Dbl37et8Umwy+3GTBIzkdhOODC3Jinto7GXgWWcenKz
+T29ZsqWISRIFzUuK92uvKQGP1tt1rohvFNRCoK6s8xz5K5rt5/URt9SiZeqbDA+
ctcdfLzv8bMqqMoLQTsMKGVhya2EQbVUw7JekL2ogxdJ7heQah0zqIWoz2+0mQ2L
Y0YEY4VL6PSEzjeSHoNmrEav5qBnmcDnfvhMSraUxld5Mo9E5d0Nyh39HqluH/D1
pML64i4a+GPgM65T/hhrBAMFqzRvbr4CWBTyPUywphNEkFNy82lXbumZz/5y/H/C
ZyA8IlrSsbpNQ61Prk+NokjSRyyS9I4L92TUotq3eSxKMLl5jys7DfrSK8ex5Gta
6CxOPeQ+M0XJViibQKdmAXpdE3RVHMtCGdAZh53Yf+k/3U0KFAEWc7ktISVp3FR7
uUfOLkEiPeLO5qJ+Z1L0YXi8TIqRMj2fZiGGLaix9NAygg2ZWEXYkE3eEFCTpX49
PmlATIfHxfLnt3msD6mofuTezVex9SlC7R8Z0kOmScMOdpikfbZsYlIipbZPBVal
GZS3Syd1nOY/F9wCMq3GaaMHRWAY4lsEvXxZ5yysQ4wtzj6e/USypyF3Q68NPZ9I
tuAuGZ+trjat4tP2O+bLMGv9WdNqBPxSfqtndKCmYU5l09SASmfs9Zahm5K+hQ5W
dsheeZtP1sFMeuOO7UZZJc8tQcxvJwbJLwdVKG/Iku8PlLqUysaeSm7wchE3IIbd
FIna+13OknvLJsD7v0aZHp3E9IGqAO7pK4TRiNHs5AXIicLp1hORJlnxCzmJs9WU
Bqt+hEP/1T0zKZWDHYVK9h03nLnXY/u+ByeKIhGGjfy0/Oyfho4NAdLENvL3DKOa
4CT+N7E05n3uMT33stgy1ob/fjI/Gu3G530sGs3vEdvbqBeBFCFgDrqFc3tcLXtl
ydbW98+FVU5EbXI0rC9wjY5SQxd17pGFsucwGDdjas4cVGtLxyBUGaeaxnvQn38Q
gzksFh9KLeHnGv6NfMdkkRYYSi7wpmEeEqG8OCYllY41NwDGd5f4eDgCFtKSr5jq
pzv4LXdqBYD3Gzx9lkyWJ/61r4Z2nXoj/0lOFiE3jFqmgGX2gFsXxHXNSb4XFVUl
1KBIeLGhrk1H3SDl64l9Ct3xhuqXy3frdKicwftu7KrXviFDN6HRwPlruxmvRiGy
37kJR8w3PKNnYZYAuPTGQpVARSAlo6UMCfzZH4TX2CAurVpeaVdFmf+tSzGCbE4t
cXp8gUjazeFFXWJP+rgjxpNDm9sqyvgy8DphM8NrRRqAVmYcTBBl6Do+NewHsIU5
3Te6KVkCLJj+NFUGDBDZHTjMVu+rWct+brEuCCB8t/+VTrmFOeS+EM717Wvz1aex
G2rSHIyNJGP5+vEec0z1aouN4B0ESM5cxCoKQlQcHzo8Phc8C76T6Z/CAbkLBniW
V6tdCX+HcUgaYSeZloo4C2oHZF+8FWZlti3iMgvKTegFSjupU2d8dMS+s26r5GKc
osu+NAXpX6C3J4JAfbRp+bU1yqaMfj8JCnWOeVTb1zZhZEvhejk897O8QaRLaj9B
ZVfRLkdoXBMbwPBKN6uDP5zQYhx/sF51efLYxaUlx0C7u7pZ4jYUQBP23XS1g3uJ
sOZh9LKxrG31X840O+RL58w2COUAYYVAED5BMrLA+inS/KKDgPY5ebpQxw4pu0B0
HA6+y4Lq0wt7FfF54Pi9IY1cmKliUtRBFDNTnmym8717/m6GJ25B+Y/CPWK6grIc
lDm+RTzvu6Ozaq66jMNYXREVo40dyCUImJAgCwza9S6dDaijyb6t4bqkiNEZAeiJ
8xF5a7ELNGeeYTjwr1UZWOUfZyISRPsJFYP8HxDjNqaHxLOeA8O3oz38Xj87E7f3
yelnm6FmSR8zCyfgVfQCcQhdxhdnPpkmq3OKDuRR2ZNHGEJZRKzsUXaB3jJclCwJ
9+f3W1OdE0/7rI0mK499/6CZ7xwoCxm7jCVDs5/NUpNs9Jm5zJcyiwLkUboqC2LE
gsTU2Z74f60OosAiEedIIvtinA5ranPZtW2g2B0AaTWu2y0d0TVPJjiR7ETyyVH9
zkkcG/+V5pBMdvGUy7D5uti0T7g3pPUy/Jfqy5Yz5/sH6PNVAweQ5XZbZpRJOtze
nZ7Vj0uuI4EfMSPfInKMhaLSlzVxIt3HskZBAaWbIOYKmPT8nGYTgcGKR9IGeuNH
OVpjj0+Pr2nk0udkAD2jQhQoLAa3WY2oXSvVv6SGQ+oKngymJUXa5B+2vvHdFU3k
LMEd39vBTCfW5YS7jlO9KAz9Ri8r8afU6yBJ6+Ue/fOvI1wjNRX7XSnK6lHxGYJF
ZBxe6n/x1i7wRXfZSFtBkZYd+P0360533WkS/VsF/Vx0vPWDyT2RpCW2wD4fFcud
R5Djld7Rcl2taViIGpGuucolTl9pYLWmMN3GyZVdX0ZdzbQvYZv5MGuRoKSMTSCT
RpuhNqRDr/8OR7KWf4b/47n8loo4rgl+q854ECcxWzpZYW9OCB9Me+5L4yAHU8Gw
Ezhesimq7KQe9aYaLjXjBRW2PyGRtdEluICK9CMmGWuM9eqSf6sBMjGxj1+vpqZb
arE9nUxRdamFA9eRLP7NFsecXmFW6FPjRCria7SwFUCvPeisbM1bJcj/0dDja0to
lqPazwnqKVgt30e0iAxMPowrSX3R17COBfjtm8fLKYtQXm8WEpxtzt/+bfKt85uq
P+E2P34McVOfS0MJsIhoGcRmN3/HSrCLLqnhgux9y5Pul60wMCgiFSZd6moLKRtw
xCGhWXOGoMqTIkAeoH0imppblAdwy8pUIk7tOAZ3XAXFPkj3N5+f0jAGRlXHBfSl
zQMi0zG8Agfo8UI86+S/BUqdYJn0JRDxF9vfiC/2quK4202bRCFzTobrWm2sD6oo
Q/pm3izoYzlGyDheObzDYRaCHLYSDIRnNk6fPg1Nxzw8nUXnmfxeKsHjbzx2ZMr2
Ar1sa9SASEejRLOGNg6EEpPHe2ZMOhQA9kO0e+YUPKLqYz1rRWitfCEH2LhXFM6n
PjxETmx4eHjMsB5FMN8Q2Zr5xqjgKX2I+bz31VdHReeTB7HpkAUWAud5k4YXrrYC
LGgILB3zz43S6ihK40rs/yu6hNfVyAOFH+oAd4c0cMbTMbhee2vEBOPwNUgTY170
YoFzYeFoAXsD3TO1uKne5CE3JqcrZ3G9zhUy6YOn+a3Dnk83Lw42TXQYdIwBfLzN
+1ZtQxtZK8uP426jjaZVjGtOIdf4T+7JTHgAA+Z2uDCLNA5B3uPKZc8CpxWBkR3T
fCmLDECVJFWuA5Au/iX7btagwCsLF4spRz/xBPJlyARqQ6GfQc/K7RLQB+Sqdkdh
woisK7FzyadGghdceY0njsRh6TzZQmLh4BkSCpRMl4e+l0gR7C3w6QSkEl0/+vQ/
dvUIEcvVo685LYWguc3icpnDS/qTdOyH5d4oZPTzkvI5FwEfLAuR1kBkjPw+suGb
UgqdJW1873MPFaB0uSt2Ay9i3hIKfQMRliHpSS1dTZWz3V8RKokg/Rkg4akNpsVU
ff3QGnhjfF1f2BykE63pDi2KFo+KVmI95y4uhT9ZSqe+BTWKZJCGmZIxwLvMCdip
E9GWI3VNmIGd/Gr8dfovxmU06UyXfc/9feqrRMCiUzOIIoMA7snfIKMJGjW7KYa3
abODYdrAL9vy3FZBO9+3PdCwEHGBAe5AYgrTAVGJacIrM1CS2aacIwWK9xsKF7Xc
URYdzdso8l8tmAFCGE40LZpwhOLL/yL6jsVBlSv+2hWFFDhDZlE6Wz5dmLIujLLC
nwhH+xrm2I5Z20BvyafDzvEJZe0P5j3ZPrISYB59tpwMUvdELqZU3NBuIGHsi1mV
7Y7w5zx0bplOco2k5GRPTB8vEFl1Wyg9FXxGs/GbUHP+uNVU0c7pJ3XghJA/tMq/
mWTC9YWhhUwue0JjGl7LjjBaFXpFuAOhlBDIssU3hYxCRlaMstVVbzuFSH938QRe
zKQigWlmJgu+PYcZZM18B4ZKoLgZSuYXt8Bejrtexq7blgDekxkQqLWsUoQVFM4W
pkwxDceBAdUVlI9ClzrU/yegzTm91/nHMCEQw1p8zVj3KuW+4YQ/E5P0fIL3XkVT
qIBX2dhFSmc8HoPJEZRQlJFcCGIgqCN7SPnm/hoKltllSof17LpnGeRislMuyXxJ
+Kj7RlIns8N27QEPODN19lyCuD/d5thRw/xzO/ycNXyxqM3jvOogg7BFzKMbeINC
BY5hNklFsZH4ZiSyFoSQ7xwAjd7wqF20N8C+v6sPNXOtvnr0fG2h6hX/KrPQBCGC
oLBnp5NdG1ruolf1v+0UNOT1wrrIDOpE8+o14REor/ZaV3ruwLsi/pCe9TW2tEnd
TqipAPdcVqdXwrwF3mYT+fybvgDgRLktL1ziu2m90ClXhRbIbjX3sIihm4yfzh3x
79MgzJMYrSERWq0oUkjIn+sGcHKuj/HInaKZIL38b68hEVdotsJpwPHn14MG3iT3
L2AEwjUZ/9a9XGG13zqprabURLS+4JZSnzAancIo/x1peJp5KfpIAfVuk7s0ulnj
qZzvqU7SDIgQMyvmYWjLcyxEg33LqYIu1i2T9lRYz87YsAOPARLYWhjuoOWYuyRp
pZyStGkWbirYimOz7MYv/gIIEuymwK8dnNRdLXteJlk1MEJAj7mJt2+Y6fMT/wyP
4gURxnHo8vOyNMGLmScSmuocJZt3exlUDsEceIyZiu+1qlTqmv5O6svjuYzEnIj4
5CnIQaq0nb1M8adwI3/g7Z5vS1VpaHbGf5T5EWe1VSBHOhR21weT5RbykHpBh99V
hDqTCMiUbNqtxHUivp2g8CfiJMhI4gwGmvWF9hdOefZjcY1slmJDs9OXrsb1UU6D
X8u4i+gztlgbJ8VrieBNnTUkKQ1T53qoIj+TFA4TvsAWFRMF4MepcJMU41WjFyUf
x44VAo80leib9HlWlkkVOK18R7MYy3p8gSUgYB601jhGIQ9P0irZJkNYWUPMAwMo
4UqlokOQNXTOS6VcRzAq6yo6nb2LrCMGu6LrS3Jfui+YwAoiAELVdZknTN5U5hC7
3uT8H9t1PVD2QDTHSMgq1bABGMM4fPZRz+GrM53PAstlmxr7sOq9kC0Koxl6Oxay
71LSlBjJ9sNkSHctAdE0FGEhmbc4LTvmMcDRCj7YNNzcEIdbjD2qERs1cAl8wqG6
3giHb3JH+ywB/CEG6BttZv/e+7TNff4fD0haKNjnU/yCBp+WQqnx3m9KF/XYqlCZ
SZX40URvnU2LMkk6gMWvDgacP9/TaJLzJltA2k5FBmZEN75hKp/k7H1qnuoBNNPB
MXuzvsgv1tcLktbVODWlaj0q5RepAr84DwT5qzhpELXSuOpH00Lp1XFp5xIgzyyh
7SXRcN1KQfE9oWkMWjIBWuh7foWPVWpw0R9qZTTqxhZPIIp2pJIyURN9YS3dkEOX
XZYDQgf6951dq4jxtMajJ0+HuGjw6mOzX9dcOnsUUBTiOvsRLbZjEGLiCuDesXz7
5IQrC+6tyGlR6Q4uIVrcynCd31m/xbcFisIZUbsPNHSiSK+Su4/uy2kvNx4wo2rI
5zefyiRNXoZ1++dPFgBuH67FWTfDtbQHU7IMJnfMufXy9qPa35EHkmF30HH90WjY
0U0U79sY2w+5T2cTdv4NADTqr7DmC1VGc+vRV4wgXtGv6XlnztpdSQtmNbw5wtXr
sd+vrhoUn5Pr2e2amyEegkMgg8pIqqIFVwl9lY4Ntbzj8GxCSRubpld12nVNtizN
+HSIFz/BrVtoy9E+ojMIQsN2tWYhmuYeK7rAjYgtZR7wKhq9m1mkOnm/p16z+/8P
AkOIUSzvyoHFmiafvxvZVyqI0aoc6HYuGFKJLw4CDcW/b9jc3aDNaWcsa0AZfbaD
L5Y0r0fEu/zCN22Sz49y2hKKwT06Spca9ygPOvw21bSfsGSu9PnNu469iQY0YGVs
4Q0sxO8Xds+eUBwA+R4zOPtXCASzmW5fYlZqjEXOU8aYip5XIcw0zJMdrs55shl5
lC/XYfdA8W1czuXTl9bO0YjwKz6XZwUUxk4bpTIuqsy/N4oJBNmlfAVupcpVf1QV
BIenlKBDbNRf38XUOeeGgTpZXDe6JwQd4EbcsKWtAZPN55QjC6lI2EJ87+yd3bp8
/OnkMI46biiRAxXpJfHWUTUZu01kCASVE4YZhW58DGdoIokwCnftLx0hA6DdfZpc
AW5cVj2rq7ZuYZWYP/2KgxvozzRYlV4EkjKYr5CpiC8IDtBfIQahnEzCQ1MSI1po
izGY6quwS0IeWcMOuIJO2/raIkDpuzWbvBlb7L/vcgAdTqfmBixor2O9gNLNowAT
w/Huig4/ECBEXgxiNrYquiTxqc4LxM8PEe4ETBlH6jOhMxRa3pGbvuW/OaAEScfP
GV+iopk5qi8SxetaYjABwQiyRZvNLjfOhfwIsiAxLQUopLjyv0AAKBm3I9dmvpFd
AlMPHGlcSGNK3Zo9AxC4Q/g50iZF4FhzcJgIJKPp45gIAAr3mO6g77b8WYunlM+p
NMjlTnxf+HmA4a4qWfxv4G0T0YlPUm28SHuh0ElfSmOwLHWQNXdOZGenby8GeFbx
eijnkKsfc7MN6YRoAVHsEtsf7gLoyBMpeWDf8oakGIUeXXa+m/IueQsDo6OeSLgO
ThyHvPSX2wxz9TsNbWlWGAIOp7iYPBugQizvNZZhbO3pdLJPuigasVtZQ+WsHtKj
9qPEpKgK3M6cUS8C0W6bOtDm3fh5tNfhRdw/tBKRA2lCRHkbkMoiowF49zxIBiWs
PqvLoh2j6qMCJiGIX2xO00/0S8Gpy65ReS1pAXbqueTRNCpEMmiPw+M6mshNHpON
6InpsLDf1ImboYeuLKwxV7Le+7NUe2Os54jqZGn1pjFT32owFL4VNaW2qtQ/YnHx
4GqgC3aUfWBmLHYwa6N5qFIYyo4eocCMF5L0eb1cz3tzhFOaZtjdUCpDeq8gJ1tP
jGM6NUjJ9NGBjR0btMiOmcc9CHhWsN5deyIF5tD1bqrj6HFINlpYueE6/+iBsR51
ha2t3OTdvBLm2vM6LmqpKoIGMHS8QZE1gAEjGrKua2WJcVbNHeM74xmeAjaB5DdI
6kwvakfXH8EhGW0irjIq/3Phl/LSq3JgbbWUPChZkEm89mTW7RgTWtG8htc8hkwQ
BhMytpo7HiyJF6Zs/N2uhI/9cbDFT2cADgKfrLj1NvWtIACD4xWeeGqfhOoVlq7Y
P/1mswUmYwhI6fqzcCu3Iax2ZNyqytPQpPUrCDkTp+XrSXpW6mr47zwE0sOhjOJh
ztnJ1h+F8eBDBzdHHpgcyIMrxvemCdQCD6qBqXm7eJmjDWJyUJ3FQnscaez+ybBF
MvrWLUuua64d8iUFELVUOWECe/TS0tGKdRrXD/NixZ/DHT2HkkkgASMz7f/aJvbI
N6DBoRgstJD0mnk+eMCOf/bGa9Yq1CpgzQ2SFrzhwPoDmbQGoGIt47ymwNbrUHo1
DpDDQFggjoOYPSDagYaxdm5ldpTH/6QxhEWI/MAmFa+813P816DcYVS3bnSDFBn1
YQb6+/gaTc1g5nwx9FblQRQ3spfbWooniHk/N10y9jrbIBLW5gGHXLgzhpJAsChq
zubYD3NIyqtp9cJHFCM7o1bhKyXYjrr6U3Zf/JRGNUY4wkcLr0+pt1Io9iSlqU/7
3REJobgHBGnqu7huPp6YwFBZdY/QrOkmjZJX5h6erQHfYkv/1b+5PX3/GHJYa8v1
NU2zkhGp3iemwtRPduyIutV2RFekbTLN0n+AvFARWzTSDyqwJFWm+Rs/HOa2+dRv
inLUqELi94dA1VY8ju+4eetvhaJC1RMHXRU+GjYS2sJJcMUFWLZ6yjhyBkFhTrw6
HVHozcMl5uhjyBkYncSH+6B8cOq8IE0+dpmKrXkPRsZK+GgcpPjkppzS9QWTnw88
/E+ZINDvQO9HkP8kAWqJt29YMrYioFF9fAlpxTqJcAmkKt7j+rCk3Cg4/ZQEAWRH
j6ECESMVV0vjVGXqT5ogIM+KBeQ3HMLg+8OcBAKtlwomZGqW1zCw40q2x2E9lhga
3RYVdoccAJemOmIx9TVa7dcF218U9BRMq6tXL32Wh/Hx0LsSpFkKYenF5ENBVbxx
uovcKqFjgySjzZPLFzCXCuZHuDZV71XTN9G0LaL+4iFBu7CekFUlNSUgXl6V+lLo
5vQlG4nRmaWd6bfjbsGP6QS2ZE3WRhDVzO0v4A82et53fX81ZR/hb3myqnm0YQLh
PsGtnDfC3RZ/cSdRFUZKIkHKmXZgEghgXCnOwyBh5sUuIFWYwEGN4cpbcHkmq50l
gsVpwFN2qiWL/STAk0c2gVaPkKs+2NFTSG90B+jAYAV695ypmdUR/qJKuZhoYCt/
uQMga2CmrEuPpmbs1ejHgPbZWOvjImSzRtrWO1BHC+sP5Amcup7rzSobKMD6PZAk
DGJyWEyLBvqhC7gHfo6u7thjRfjQ/gZCWBl9ET1gT7+g3/8XLjzOLFR/N7CvIEqY
NGlqPVVyVlNSIWIQ3R7ZSt9B/HUYV4QiQPs6IFwCb4I5542OEDyzLzdjri9dwi2P
JchYIh7/FsjZS/5NrHPwg0ar3aoOvw7VSVPQBtwRpSDawyDLz/l/+s+rWqmQpF2M
K25AM5mDkiFH8ttkFX/1AKarMjx01OOdltWxyOtCBUGb22ZrgCjiGAM7sQTrIrdj
oJbH3CUxPg8fBrje+/T9P8KgjCe/JnWDHfVTY/p7AE1qKlrdooYMDBe757YNxbdP
8o4iCp9McCqqpcC/HeDFkUPN+2wGMa8Ua2JXTRuKufx24ImqB3RsDx94cj3cA0BF
AWXqP83RpCW5wfUkL3ZJSmM5mKOZOFxdMXvIye+nehutcLNZkneoOQ9oCANmacdW
3IFkFh3Ve+DXZAAw3rNoV7ogLl9kpV8KvbmVBlZu8LkyMlNsVga6AuHQ0fd3OXCz
0PFZoHt6SQkMYmE0uwfdkTB6hH7I6RfBAFj3NUmwUy+/I/IJ1AElH3pgvSpWi1UP
TQOROsZGXlULjls99GQx/QmyCSVmz6hueo8kKIwLypbS953v6uLh2m4xQY0KEPmZ
n4kRGouIgDeNKU87AWU1gvAAGxyUyN7dRcF+cD2w4RuwDnYiN+aa6ruDuYk6dfyU
TaqNYS9frd/VBpwjt9l45+3Gna20IcUNhT/E0XXRMGh6vfyiI/uKIjzBYZJj/3R1
if6ItZOagwd0pjOkgCzHiA8k4pz8z8rCEgf9XdffDDUXTksjHiOcCscOYm6gLoyc
NhJ1KhIvCTp09HZK+HMo6Lndein+Bh31ObEFABLctpyEyJfUbRrEAfLbA0VGWLx/
Y28yC1dOX2OLxOaLYywV/r98DIu0WSAUTuRjuI56v5LOUrCSqneqqs3jHbYyfoEv
Yj6FLWBFeRT+psXyvAIsHYr0HCGF9ZRq0eEnRUutc+pd3K/AaHwp5tDuGpqEHPyY
dhEUEM6C2L+eUx3hzJPI84SmJZDypzF+JqMlPV1xgZ1VMJLxrddohz0DIWWN8zvE
P9NMSuKiaQmlMeZ3BwUvNuoGL7sGDKILcJVWveHKOzC1m0YgWpHDDp2gYgIfFACp
XiQEeeWbCj9HU56FrNV0i2gdbHfVer9DLwfVEG7Ue4woSl0yODC3U9U+4LNzxyDQ
9lNjhn73c4ndsX453IB5O/lLXA7OcNQF/Z2Cc83TCk9u5SGUhgkunSlaVVr6w+Dl
/GUmFcR0+dA6ABrSMfoae5zbdH9yG3cPfTUyn/0Vi83XSOuQAddyUEYI+oIKKRaE
aX1ODiXvemoazxhCBWCe/S9p/QWr2VIxe76ymaqk0dYXbK9YJZMGA9SoJw/5CvEe
1AEu216uUNB+LelDoF1TcgAudxIYxmbVKHha8OVC85vVrFQZTeMNu4zcJAGiu6FD
98OKiKVEPLzw2Hu9IvFjMqHhFDBZ8tUCbX+1i2c/hCFK0whDQ2fTIcjHyUBjLt0J
8axHqlwNlsuj9s1lfVy1omDqrqFk3R634pCYMITBcTsDfMVr+gh9iDMqE0lMlJVs
U5L6jrOlSBlAb40auCiQAOQjqMTgErWVecXmXin1/xupI0o/FwCCKGnWvgQ/486r
HlqbUYUugOkYOFGVvhTkgR03QUVp0pv9Ik0X5XyAEmVUcGaZ5KYglae6cnQ7V6yY
jrr7izZiRmnQ2PF2jyCXkuWyhCocNJHXlsJhSvY85rGyTKGMH+alM/CS6XI7Pvrj
cgZrgjv1f0l5tsEUEW7YUprkQdxtjrPJLWTzYVngA1fxTGhh07mWCzREjepifEvC
B4TdiGIWy0W+6OzHKmq7VSr8tUTk3Ldh/tiprZ+HlGb74RvGJ7aZttsIwwb/uJZb
PUFyxKc8tnK2n89EKtRiQfgqKFVrNBys7spIjtxqJZUwNb2gerV10lrfrQIV8paI
Ym1eiqExdw7Y/GBfSByI72B3g/oP4cTsB1wYstr59L1cVCFAdkDk+4+qOWLWvPDP
tJDyc6jZWZv3I4eru4yO6zq3Mr3ZE5AmviiaJvoZWZb2h2OJ6DHEBA3jvX2ovvsn
CDD0uA1r+8Bv5JX1pE3x6TD7Cxsgt7y3P2K6NEFxy4MEr+NblzM8ZqTN8D8a+I67
X5/0naVAsXgQpIAPvvPldpuWVTlrHw6INLoVk2zCFOp0FKeWhIbfRMFXKr83B6v7
lgT3xh39X/xNXCAK1tBUlTO3JctDFGLrkYcA8Ng5Rp0u/OeHyfjhs0sCeT9LkaGM
cq2vW0vD4jGzIdPv3Tzwy/sUESI6Fta8uUp8lTNfwwjjkLq9RTDpCbrvMtDu7mXt
tIIsNUhTZ0c31MrMn66Aq1T4M0CJHikrx0/Vw2UG+DlhtwRUdlLWWUVo66+Gq9ew
0xta2ARnlSLajoLHZwh/Cq81LzGWIx5ACQAS7T23PeAi2ntcCCA+umekWAyChEjO
MTVfGlrVs2cNyYZoBCTW7NT+SdgNuqn52F+IYN/7WwPfb0x/BK4ZLxxgMw9kDaMV
miaBwufryaKAne9KFMGEfnk3NKyRh6NL8dTiv4IF65dqpp6/WuAE0ukbhciBdTKE
xIFJUJkDvnDwip3AW8DocDFsGLNSJWvTo8mlz/nZCXZVtfI1WKD9XNw9Uh91EBvw
r32iulm1znbzqTTBUfopDw479ISC63iOuTX10RQ4DkgamaNf+JJWIQIqxCi7DqAr
tTCKh+NLDv+SFj/pnViSYBPmuJN4IsxbnSQh6tWNV6EjakaZejredHjATEUhGToO
4ArMYTH1bUdAqbBNZttUcQ3Y3ZdMdhL9/aqurV5w/e2sq41mgtII+p+UbcYgTLAN
GkqLH2e98Xsah2WebuUCSROTKdY3F+fNBLbx2A7ezfrtuPZPyvQJ6lPogNX2Nrjo
51Tgh3mebSyaxn9DkcXVN8+xGeTynaSmhuCSNRlvjiILfMsZE2FhpVOSuSylH4AZ
RidBghZtC+Lzs2Ra0F/IagQhOoiWW3NtlBOzBTic3IxFQl9vH2Wir75bS717i7wl
lWmB/pcpuypvc1qWR+JXFI8hERL3J6/myMbuC1iXrmpiSFtLxU9iCLQP7yRYZf0i
rTbRFUZcWSK3kRoY9Ar7XyONr3GEJFOla5nZ6OCTs9z8xZIHL4P4ttevkSXXPkt+
n6nSAlzuXMR93fJBLD0+7NwfPpBYy4aLhlmks6vdp0piPYuHxPzU+CMWnmNoWB7m
VMZojdqxlqkHhp9GOYp+Aat1iTdj9VHvckL7pv/3uXSfxZqXI4aYMwwX9joNmR0g
7LFdFIWiDYAtgajMWHquiYg3L1Sbx5ikJnk5qsdm5cZCRA9NhQU4a7W8efTYBes0
/vm0yiKEHd/X2/9egvGbq7E/AfCgdPW5nhhuB47aEEgpoPUm5Fe14+F6SVUxZA6f
KPlMTQBGamQcs/z5QKzsvYWxXmcXjRdxhySszYu0HdbtwYNopVBBJnT6ndjuLO9q
+I8xB+zkmEjvkdP5QUVUDe8TkGeRGL1qvnvjbH52y8N2fNbV6t0UUI5SX6MvhF0H
/hlJ9xVTS1vK65LXnxeX/t8TPAMK4BrYa8Kuhi1xOaKEb7CIpQNUFr3eabE6GqVU
0i6a2dAhYEHuuKliYFtscBS9Xgn5R83THNAko1RMJ7iqsJ155gqRfbDjroENldLn
BAPHa8A27XI6MUhQRO9cwBirdqkQ3S6/cD11OK5P9LBBSINy0BlqEDWBR8A/e7bu
lZtvWhfyncJuljHEJprzUnRZPC5bi0bJXCOryQ/IyM//oWjL0Hfb6gsOCX2IPiVW
p/HWTOhTa77zlVkFe08b4WmjTU/8K7vC/ARO23S5fms99OPKKQdCLMafv/nhqn79
OtmC4H7ERbJFa26QN8H1ldL5JWThUHttXMX7thFqeRSOh71lwg6FxY6DIb/RrPF7
pEKGIEFXxgxaJe133aODNywlmjGqKl/u24NpWr7mzUsH3rG7KBTTTcsXfS0ogMtV
TBvlADTvm+73juRa9l4ag4DBFI3EzwYuhtj1j9zMdTUXxjAIcE0EF3tDBV7CNBYt
1OkjY5FMIlyiVyBBEDhtpiu9uNO7e3sXtaad31adBYuz1a1zULVp5Ygx3ynMhpue
B+znuY5NnuPVzXdUzWP6M6IADljwEfyribR/hlHRb8Fc8A9sF16DKDXIrm1Dwdsh
e264g5/I+80j1/4iEopgQZ5pAoKhkMqLzegjz5mOWqcZbD8lx78W/U8Gydgmrrym
yocuyRDBUgatG5lpQV6ei3lT7810Ejfhe1uB8rcVY5LpKIOyKtlJ9q/ivX0Sxjxj
lzlPyeotJTVEsgTwCnIJoCxLxxlRWvdSkTBfFvD1/FjEl1Nee4CbDSv2fOQrHP12
bNroUDqSJgESd9lO1skXYDgewhm+OG+6QcJrs3yFzQC9R07T9zLiJlcw5tLcFWQt
2a4MqHGwi2yyMW4NR9GXlix+BK76XzSqRxspk7AFa564GQsXnDCKTygMCTSe+Oxz
3Y63x7UgtLaJL3JkiXoS5xKFUqSYIQqVAEt+E1vRoamjHr9FmZMAuQuP/U7lhyQS
rHH47kR+8st5vEO+oz2cgKav4aBFjNdGxNB2PvVvHod2tQiNotApTGuWK/g6v6rj
ZKxtAJLbsnVo707J7s160hsWkkmeKJlxpr+MsHxzF61/riNv590zS49nGD4gUFzG
APkBxGi53tORzKGIdADGYdiFuTIY5gdtPy1jbYWYFpyyJxhAkucd/s31/GNrpVN3
zOEBJ/h8093T7tFjwo8cZNqxOQq3vxmKbXKG+LdG27379ghHvx9OEoRyO/u5Lqw+
0D8LthH7vrIS2fnbQeorm605OII15K4e1aIFZgg4P0pvZcGdsOeco6+BkRMAKyFU
/s+Uko0fW2NosizhZ9iWRLMtGf0zz+UmkVPg9Zr8U2IkRboCixi6YG3Iu3qOX0aI
XKs1Iw0gJ6gMFwrjPsVYECe5AW1q+lhROMQMgJmBco6Rw52zhCeq/pAYKsffVIq2
tvY93yTsBzUofO3phXo5dAFIyWEvPBB/9PNVAvbzxdmkCk/d9A/47LHpEVTsdAGt
cSypYcf3O9i2Rckrx/iww61cukbDhn22gxs+Sfw46UnxBToqp1airOmAnib3bytQ
xS4jmpL9TcvFEhKBScX1YIugYxRsLxFl4LMOM7MvanOh3IyARsOYuzxmcSphuVi/
4PLNU1mTRYDXQohSK83tD35vs93fTUWIboKIUG2qmf0O0DMueDoAZoj0TuCJKHX4
lUZBUZfLKOmNHHn9ZuxpteQzH1v4QGXJ0VL/JydcyR1vKFEQcpSAzP88kn8PQqXm
RbUgVXgXpbsWRPQz6VnBuWtWDXNYFnd3Qd8ow6MQ4MY5n6tdydRBmDuGk3RC8gY2
5uH5HXhghZ6ZVIZFmDBO++TRLLRypASPZn9iWT8VsXBJluJ/a6vOqN7oHqroTWKg
Jadd+lmpgnjn0pTEg2ajzdZZJWFtebCqWzai0nLrMbviWgfNTXhiQPOjMH9t83Ag
Onzy+fX2VERP38/NixxpVQvdiKfkJFG6VnHqzTi5HcQoIhWW0rM8zowMGJ56K99S
6YST51SpF6e+9maaYfPIKjYu/CWmdktr/qjbEsZFQTbGMq9a6/Aoup/Lf4vAM7Qo
NkHK0P9Ugr5bICwZHf3FiUSDhIZUPCxPo0IZpEdkudnHIjww/BL6HEQB3GbwEd+F
IPPWYEUMhRffUmJLTHwB+WPDBAK9PsuWZCrvkf6SQxyOqSbjKenGI6tuAZU9yKnK
DHIYJjzmwMXifnKZHH/mdhadU3NDE3gP9cHqsZARxkiZN7oszS0nTwBanNfxy4dh
cnBDpiMGlTbkLrQX94dAhlJOn4PJTtb0o9Pzaeh1HSgkRxC4cjrA1wPfkNwqiumi
KhGlcA60E/sWkfnqzuyK8VYluZo+41qp2y7lDT+RqVp40yy6r7BTDQlosNjzKK5l
aZ+Ee7uqiAN21jcTGDMY2+Kv8KOmF8526haTbtF+DE5JtpoQuTbR6deB+3zGkUzD
aXgVrAsm7dP8o+qGrgbhepsQtSbxZVmMpKMS8BEPrJ4MceHfg+cjXEO9AY/y3GTt
qwif3WejkRmPuME8ur/+2UOorvP0dQHEyYZsqeB/5UrXvuu5IMYVlY0aKtNDkP6Q
Cz/kvFhzXqb5N7WlyLaieoub3+Q0Hr7vM5FfAI1e+/ki2c+DFnzmVy2AnLGGMYD7
mkyN6B/ahNLzzlw5YqLLbYDhaZhuygaRK+ic63uQOvc+MEBD6Qnuu7C564RhQm+T
lwhUMNPp29X+jr1nfqg/JC/o7O/hc5kjmC70JRaRyghKVsdRuOAGC6XYEF9TvG0p
FrdZcxMo1dnFfbdKLsdR1qB2Jd5vO4Hoqwq6gPwztJC2kdJD2++UnEvRfnp7aRyd
k5ssjGmJEaqJstvWSi6GRDXMIltCow42xAegMepxQuynAlPRXyMJ0k2Oy/v7rBwa
upoJ7p8e3wYbpZ7xfrk/l77f7+BKmR6GjM4G5b3Mas3+boLBhgNubfVcN7uLIVOV
tE0V+PAYZ5assFI8P9GeXCQye3NsGnq69Eh76rVAK3RR6klvN2ZrXZlb+jhJxexZ
oG0X+MjhEgHMNjGJljN1YSAvTOZLXcYIazr7ghsOaOgItwS+j7TpwptVRv+Xe7sh
4RiEufg/8iV90r4DcLD50M59qQ6ALJyxlT60pbT/2y6+4/9A+gFNQTbPmc+pBqZP
BHBQ0cp3BKRkJel45KS4g8XP22QF5FM3mHHRf4alf66jhDcQXCMjom9YHi39LI07
a3Dabfms5fA+V6y//5abCex6jN1zB+ZscMiuxwE/Vy90VC9mJXcF79lxNJWGYWT6
bL9Z6uDrQu51cNs1F/c4WCG8N5U3I5pVjoIcDRCpmSftrda4Z07lkp+TnRRZha1S
lpPbZQC1eVx4OGtTahzkVWhaDcObXOSn4w9q6nKiK0vOlof3J58A4HCU4hWG+0Pr
OiHlLdB9QzcEDkLc9WSiBlQWzvN2qzWJS04Gwyr5Dyh4E8Pw9cjTbIKg/Y1j2Ubn
z7tB1XLG1tyN33aau0WmlpXUYDkBe5BAxs+G1UfOn0wtatLgjcSRwOELRUIm23Ry
AWgfgTESsXZyPznHctDvxmRPwIQ5jyuFL7QgvnH5/B1NhD4qLSrmxv12GDgfzgnN
wE4Omiu1/kfO5tFJnB/8Yh5U6apNxav09/N6l4C4cwOMncKk0DnEeTIN5kTs78F7
E+XmDZ6iVRPlvh+k0hAkRjHvcs448Y2WOYdJVM4cdgh7v8Ut8CFpPd3FYI6zZeeH
EDJhpyRBjjp/FqG2NeYvMvzknwBXga5J94X6kSP3f7tzh8LYvUoskIiIQ35olAf/
h9ARHKaJ8lTm8J19EA6wdMN2bK1VQR/95IlxFvV64dtumyHS0g/NJQPA7Lvnuseb
e4286igmdOGsgXNOLBLblIcs5ksEWVRQCv8L01Sw4Geqllug/dqy9OQp+GJNn/32
pi/RvX+mYqqwe9VKuVksL4YTAi5/vbVSf9KfcHaCvDEXTQ6L54nppbUvQ8BBI/4D
bsqy9lA8uGfsg2qkc1DKhz+U4/Z+kxyZFqw+sc1z5UA70D5e3SI8xNWk0GcRHXCt
L57K2hcRMuRsO2WwvjPkK+YISVyXm4w4ISMgZh09PIK9sYE7JJlR0dLhZNBnvwkv
bUPY8r4dJErr2ZXP7kjZUSPRvbxtNDxPoYGi232gflpCGYprospRF73M7DqLkknd
m+pAe2d8SfsNmqgov2an5kDeUbWeJPof1GyZA5Dm++ea+dADEA7QtPbcy538B0aA
YT0FGFyL+2XNy3kYH5NLFmkF4q9cYJo9uZsePG7rnF3UyxxTfCWcKSSclBCBRQDj
9Kbg7pR4Fw+b0381quzArWPlEvbnBuUnj5SHI25aFb2oz6Ez6eRTppbZlFPaOB9+
lhh5cDfOv2gH4qSFpGIFAS9EUqPyuV1rFQisVL6nzw3MCj1kA1YUYSlM7+j9758g
Z26WNbAvy4hsO5VDZzXtggQVfc8qMHve9k1QYddL/9V94J3gqDKjjcW2awVO9b0s
szSJ4etYxX82c6dMdhp8kvyr/HLe3rMrECWgYEBw79rEiWZ3jvracUMgx8NZK7dP
nnDwlL1we5c8Qzb43UJVNm6gFc1CHC14trnMxbqkuyTuLsAQGHkj+yvqBXazXlZF
iEfIW814Akkm9vFw3TY9fjhTRQpDdZNWGr+KexxVRi1TPmQ0OD4sZSNqvRrUOI5Y
rqMn3dKuLqwKJawPk8prnpA30Yc8v1EX4tCz1orrne72bgePirlaTVEFW1H0xJ+G
RWwDLh+FniztFERr4SfAXl8NAgJ/1f44gcIHzUsm6DBEhvgXEXLRHNFX9oKJcqNk
At1BexHLuskzN9Y/JzklS4e5c1eIKREDvNPkVGW2DGOybWmYl0E9sspXGiRZ6wYT
j/1TpEfFKMYv9MGuAWUWyF1VjoViAm9mlxk8H8d9xaYCratSlWZ8TDJLLdlwuZJh
uP+4fA8272jtbQo4SPFpJxt5Q7M8ag6CI1PqfH7667ecnPMGthM7pWkiVGhuT+vb
1KiqR2LCj3yk0tdBQE2JjLps/4iIu9QLxCpsyOxpOO7RKfXIK8j6bS0+HI4UFtsc
IeBWNNn/+jdn92fuA6wWBxWWwQt+QkjR23bGPkzl57jASkcm3pSI54QPy/997jF8
zho9ryweHVFH2ZJ2W7EddwKa9Psfwb6X3WqhPUIJzvXurQTE3XZ4pH3LyUhp0fOJ
DDG9PY8VOJqMNFegI+bQKztoq0Cbdp08KRjCed1Eo64lmKoJJoNETFh+Qg6JReHL
DCIu+GjYEe33JWzcrudsFOt4T3uNo5XJvmJjxm3GRpBfnkKizdafu63k0k5l6z8D
vs/bNgiyQ0g5GQhERp03HPaJTJS4tOse8+z3L2GtKwnoOef3LaiPnhvqVcHAA9bq
L0+a/hiT0bFRXmaXkldmJ0/XqZlUQtTz/WLMTqspAFHV+OnKx2u3UVQ4UgXJwFaP
ybOZj7GgZf2v9UAKK8rDuCF82+mIEzQ9Zx1ud7WAu0ywMB/+YI5azHdfJ/HvMx+O
E7onrvm9k/S6fygqx9A/XqAQYbMNRU2wmTJ8XzMJcGsqq6VVA8tFGEUN4V6RBnz0
+MyQ/MZ+ozekPNBMyIjUHa0D2jeKBDQ4dev6UEnQ3evLDBrHPyauBGoGJEsRISp0
7GSArBQ/jlmMnQgjTnmeA3OMRwWigvohUWBuD4cat0aL3APu4sB5mDmhha51eQ0Z
1o2xtiWOaQBo6PtQnzVAK5qqi7fHhC9mswjSlJ5cTOZ7ViiKWg96tvtk9xG5ZzQS
i+A0q3oXUqnThO8I8K7Y3/taa5v9QcLeyt+kBfeG33HPrTozKXkgKCP8yp5Egik3
y+Gfy+iNcKFUPmgso6cFYjJ/V4nGOGTGGtHxtIUNyzQizEtGqnMWmRo3EnGwuWcy
lL/wzgF076sm+eeI3sh55xSoSGplZrnSN3kbDi1tsa1OuoWnZZg031Q/EGeyU7Hv
dL6f5I615O+4Go0bMksNBqLfRbeOrgMo8gWKqO6v9wyt5nkwos3eMikS0WOu+X2n
5w8NQ4JRM1lp1ziqBrsQgDCs2HXs0FPcIoJIs0AgzTAh0PavNsGPjFZGL/8Hq2i+
Z5s/tXPSWmhDAZrbhNxkwsGufoSh3ovNtjv9GiObXjOelNwJz/XMKn4xLrVRK1Rs
cV9CWjthDcyEi5o9hJ6ccfJgYREjlxGgeuwF8l2/aw6ouNPTtTcb0KS4sqj8W3CX
9vd/Ph83t0FPeJyu/vpjSqJU7oascIc0FzYLmsMSakz3dIwIjE32yFaqbho7oCxI
uqPKr3fy9IxgWWVRNrHirD92u8rOm2AXyoXnW0FptFkdCs/hDuF2yTHXKUbnOZDn
mtrR70BB0vTeS+vYUEtU5VL6tL68X7dHwzxZc6c2tFbePUb14evG1v8IG0z4jQOM
jzNYnM+HGWB4eDBUUBC1tjVKvKrJasPSYaiBzZGXnC+FklX/ZMbPxROfbxZo+n+Y
PD1QjLd89m8juCmh/9bGr4TY9Bfyc5y4zX7F5it8prTN9Bz9ozeFBobPtmN95Ku2
/GP9apMm55axA+QIYCZgUF2UcztZ+qXkdZgFiGqZXShBN6LCeCCoqWoEOAUIo+fL
75kmFn5AVKIMl8t1fRHiroxweRQlLuysSAScCDPoY6ZXO8vd3YsWhdXS4sHqnZSp
Qt1pLtTavqBVO7WSXvipX+GeSbSckRJcrCExr1AjbKFXK0Zd/ayzc321aWfNNJTD
OMk4DsFHlauVxjBdHAsqsM3IWvQ1yHiHtbmIxfT31u24Q/QByS621SqSsDu9zF/O
/dUIVl/AQAaJAN0Xon4cI5fqHv8MjxWMNdaOEbSQQNMNPvoIwRFBvrVeL6jKgvVa
JS1CWGCJMHbP0APpB05XnqEQNf3Ju1AvEoRoLMJJSs5CsSnAqHYDA9glK7f8Yh3k
weUchH2gVL14hXkIsxWicAgBl6BjraqrICb5xTxBzjYKjE2Ip8OctMLyPXtMV1xl
kGbgIRCsds/iWkS0IgqesWB0ca21dBy6fSXUbZz38b+H7NxZaTpzGK46jxlL8NUP
ozu4Dc88vGyTpuAJmhY3jO6BtjJas539f/7BJJOBPxqFrDgeL0B5k8DVxSI1MDbE
X8NbZDv9Rg0X9IHLHOW3pbca8ZQLbBV73adkMXqmJipIGaftx3Qdf5z1jF5P+++9
iwscdxmSnpdh1ThKZGBq4+xrFi8jpPFDO6i8qae4L/8QawUp0GRNfDUoTOG9+Hl1
c1uo61Eqy10ielaHK8BBfwh64NRAQg8D2FJEPBFvJUDgxp2Pr8WPhYkqZCHML7gM
56wiY5eoRgHey3cnNu2H2aRAuwch8q1QkMNKoBaZJyxiXTLAtqu6o4JZ7STe1W7y
67xJaU/q7L/OMLenbBTmDdS0/sl65rhhRIFZSG33Bn/xlfkZAQAUzLFFlrnPzDNd
GqpJF6xxqtFB0Eh4qh6d2k/Vb3oBJbdchovVnEfgGoH+OiVUWiF7QhxVybKsVdLI
5ghmXL+ZCISQ7deO/vULWk++DZjKk6laYFDixTFwEqXbrt3CTjjlK8rPCQtUSoY3
zmQclLMtdrcdYUjmhOr2FdSE2Zmw7faSMuczJAJx7T+e7yyAqFQoqBPXywljRiyg
IFv+tWJBFVYP8IZTgdnU8A98nLtCT+XmWzKg++9wXHH8/gNvlg3+DRmYcov95rTB
nmgSDYQa+ptqUs6rDunXOY23wC1nQEvuIhXXMHpV23WdMjSqPlS0Bp8ygg4TB4S7
XsCCnRJHG5r5kpPGv8MPLGc4h3OPj3BDcBwDtnwmSKIqbwOSdJjFqWsIGmsjLMUO
aX1oHjq6EqG8KGD54V7d9kmlJg0JxgtlH+qrZbWNRjQqf9GsJChIghvPFDD/fn27
JEGG+u5FfSarGy5/KSbJBjMkz5aoGlPvmdw4W/LygEyniNEcxy27VvVpnGFrZ1qe
BPpg1YNExzVo3eZ6/gk5ZtMQibI/IA6tuqr67Pe+2zuvG0Y7WN8LPDCIcyTauQ1r
wUMp65KWT34KrQ4nnQeI+i3KvYNsDz64SCuBooGvErGwgIB/Yl8LyDeEIzzBAFyN
CYZ6K0BSCTgQsZZ8Ny8x9YoYa58fYABk6/5DEGa5dCZpvohD490yaPcA7dJYjcVD
yjRFMXvkcalAjRJS9DfauacTEMN0NAZyeCc0G+CmIbiMH0AX0LEtpHErtyf3Jcqd
djbw/G6FjRyHPnkpue4j8ecR1sXCTJTsF8NrEDJ1Il6SVC8UGGcvd8MPheA2gyR/
9oLQ2LfOBYERl3scfbE7KBwU4SxVTOHFb1t+Naf43WAaqxHEJ/VKYoHQics55rS7
PlRWlChCISj8YCDTgORgKROxmyft8ilkGJKaQr0R6oYP6xieWXNB+7x7IM8rzmbZ
qj/ywz0Nd/PfITedemK613oLY+p//UgmTpC5FbLdrtBVtz6mnCcYn6PNifoWDkex
5GgS2X5XjAlSioATsLXyqK7a3y9YT4KzDHGeFJf/w5ZQa3rgCeXZzAD0xS9wxzwI
0WhoNNJ47etP3TZEL3rAtQr7TaDkTFjWyHJBAMj6PSCHeOH9yrNfV57Gr/wMf1Yc
v320JHj/bB2nSce/k8XVSLkX1fFkh2QaS+UBbCY5ow55DzYJMQsg/Vz9eNldZ8+n
+2iKMRzCAjYhjwzFeLjlyt4sI8L6eTgIoWLpBFE/6m7OGK4xo/EUq3Ezu/jGPYuW
ydA8jaN4G/YCVNkFZbu3rwrPZoPzVCtLLamQOsWSv3rSfXXLpW3h1LOwoG1f3LN0
pMAxBR/5Aq4BGDF1NqRcbw+WPxb5R5JIY+HI5UFKYYZu4r4iBQcXuwTDl+gjjbWZ
ttqROhEnUcQ7XZHdlzlObEG5Py7gg/UExUygGRAXohTnkWpeU96UQBA9EcibXS75
8GgG8eZNkPDclPingLeSF8OjHZJBrrFl+UAoh3W6jO08hU2Ky7g3zTfRNwqq1QV8
AYQao6Mn/vME+NppCSjjbvg6f9DV9uHGJEl0CAdtCyLHPP0JN/XweMlxNiH5q7yR
6+1Zj1zti+Yvx3lCdpgr3vlCHGijgCbrpbfwkjWUo6edUzlt/F4hEyrvIFPm4ZTY
jIGMfiOxWrQKMJrMYk8Q8VAWlrRNDwApW1E30ByM2xh1lfeTp7XhE1DKatbUlqfb
Z6dkvrAa/kbTJz3aJ5wmOfkoR4Cro67Pm7iKb1Nlm9kjPH+/VBeLfeLRJ/yQbS7n
ECH3dFr1AlA3Evk9JOYGK4dkqSjPPSOrf8tKPfIPypWkGC321RZBuU8e6IfGaHuG
mDI3DKaWb46e0Pbf5Nskth1yoKqTY7FrxUEQR4a/AIvzI+QsXOBm1oR3/qpCgrUm
6nCfDF70wBNG2f9voyJ4lZ2ZzGyBoSfrA5fhmH56+rE41paM1UeQfOUHbec63J+N
vH3Bcjs8dX7T+dVpYOXnNrceiUCoC1DpPrarnwSbD10g+FmRkVXD40nljSZzr7Bk
5xFrTOprOM6MSf1on+6VjNHeNRAkoHgIFPZYEOsX5H+Go8tYVYOK/O7fzegrvv3X
gWJxp6GUhVuqoDkRZy1yx7W3kdZlZA44mrodNHAcJTtrCNwRXA0GxGXwjj5h3Bjw
ZW4oRC+8iI+AP5FSObj6RrDJAEIawZvNLciP+uhFVK8bEJqBBFymIas+RWXmx3mH
Z7AITmA1B4DdoicOKukCW5tl+LTIObdXjFHdsdSka9fG6/+PHMsz1BPJBOis7K/n
TEe5lKlFpf76jada7co6VESAOKMpriSogix6eAAisut+T4l1rIsgyXcazxH7vu81
1oJcZfRfH/WsgHtnLHVdOphBYQYUQLSc5rL2PuEJFj17diL0pIGVTFw+xM+pJWly
yz8Ize3dapZNybR5qowX4KsMpS/WrOexMtIg3Wd7VItI3IG+WHjeBxFDfEtxGVE7
I7HYJ4GQnE5WsuSMTrJzyzojY7FsPuS8RShAw4LPWDfpM1F2AutoeKwte46VHntC
IJxaiQAY1/hlE4bxnC21CVU8JvWxNxfLlsA/Xja/UyRGBhrENSc2Vo7EoijhxT1/
SoKQMYCJV/+fBYgpCCoZoz2xU6gMQOD/Muf9/JpGe3fFTMzfM66V9tNQFqBecPT7
mbddLJzQ5TFek2FBADZD4m97/ZLxoSDnAOkSF7/U86a/DPuQ99TiQBp+MPZg8C6h
p3X/FuYNxRulHHU1vOx9M0MG+i0qAiBnDCnji+vYlfttSeiqvMnQmPXMSUzntyLc
9eA7Tx0CSrnIRQTr11Ie/GZhNpiAGV/ZSGPQKHH3qMV34ad9Wn0xV/zqPFjC//Hg
lN3o+XuVn0OWp0+v9HmeZQCYWV0yxy5AoEZ4++EQRs2K67qhTFzpH+hYRFa0FMBw
gEXL2I300BsSxMs37qQbFZuun6fVTocFzrQ842oNC9WNGghLc6uGA10Yz1tdT784
CUhcO1sv+n/F8/mRttbrkI7J7NB1iu6HAcmiL6kyuHOixjvwcoKYp1wU73824shv
TQwybszTT8Yusxu7qingsvZ8abMppAQ7l2dZ/Z+Qy6EDhRtOTnMoTzCpR6mLrYe+
a28o9mi8gCDmZYqAcPRIRAq2MFA+La1DNpbxJu4kAjH5fovJw9BDSG/Qp511f70v
4YEWFTr8GS7mYU7R/xyH7zqNQO23o7L5eEuFqN0dxNRULTGuCDbvLlpcb2yzA4Th
Psn1y2gnlVHv8No3M5uZ6Hj049b1iKOh+lfave6hQDSVHK/nZxAtxe56O/O0CydK
aMdOZrKpN/OKHhy/ckszjK33QvTH2hE4RdSEu81KGx0wIxqXr2NSVh0ATMlziZAj
vhGOnb6g6oQ63LEGiGf7w70nekRrguRmwu+Do+eZ2gRH2pP4QjqSFkukU/r4+Yeb
OjHJPeqWBMFwTHhKNj5wiHMw3idHdFYh0Phwl3gfKwFRQRMnm36vHKhC0EZwNIy5
+Nyw6x51rwSrBbI9G3We49Zx5F7xRnhFrT8la9ls8WW+oztJexVZacRQXMbIH9Kw
MZN4Ysmky9q9H8Cre0DjMDED0f+Z+6WtjC5x3WTBJVJ9DMS9tVZiYLlIgwwKJYUb
V/C2bUhJ+QaI/ReYW1uPjAhtKE31Kp3jo+bEbTMtrYoy8LYKhOC20gNIrQWZrTjt
ZWk6iNEEpuHHohwB7u0mNOOe5gdQEZG3hxTlXIT9/pFklf4CmEE1cDtcwZKbxePy
gHvgf8qPAPkm1fWsKndamrTC9fRTb7De5EqfYalaas57FFzzsUMuRRt2dp+v27TI
7K3ssQno/n6/6aKhfjPso2z0S6xiVS5vZOpbkg17acaFAd2dl6SEh1j/nZv1Zzw3
JdW/kBfjfW2OuvuEjZ8UAr/hr12ZavBrH/eKjI83MyEaQBa5U8tJCvwJlmpfqN3B
1busdo9z8q0ErzKL6xPIaW/DarmLwXF/Aal6kXqnNNb20d6/CaFXsQaoDCaO2lLh
ZUV/SEr1hXZ4+SqkMGYW8vcKerM2SC9oFBxaqNhKYFVzefm5TLFKyWQLTCH3upMX
6WpUM8umI8utl06w4psabYB+6nwTUh2SmQ4CUZeOMZ075os0RKeBCLIysjba5Sjx
ftpbMhYq+ZVS2RlirENL8eFZnABLyl3uMZtjqf9uDUqCg87eWCTCyrBvtRcm+MKg
pioKGj4/j6vQwLmxY3s/ldq3zacmx78GWwe3jdwJIZk3VUAdN0+ylDQ+SYSLHBQ/
JXXWWg3JHYWVcEuTjAIUW2jiYz0TGvYBXTput6cz5rndRosauA7jGRAsULS6L6Bg
BaK2gHaRZDEDTKhDU4ZJ35465jYyoIMxYkH1EA7Cwkex/qs5iyXFAOxqX+9VPTFb
dkOuEaPYHGHQD1x01hIeSTqnjYhDY0gzzfpY6SmtQ182I0uNCdXoUMTfQIiMK8V5
Us907MkR++jH2bgEIOOUumA9/Qk+5kNbIBDCJH8csHJmSwdFOFm3ZAiGRvPNXGfE
TEu20EQIBOttIizGH9y8FfhhlMPyvmVX5OISNfUIcNMxfpcnItzvB+Ipm3pOALQA
pNWXn+DrCiMMQYnhEhYq7W55rJXEmadv0qGljJS2Hhl0dlNn3xFoBY+ceUiUFsRH
NkxrY5OiZC0BMk2sRGHy80tsTiEnwWCAYZsKC6anvycIn9QJXM3izrj/140hrN5O
jRLTnSbqfmxoKgHAMvdfsTEQdTWfdbL89lIL1px+FgbU7EDVvqG6s/cxHRTTj57Y
twD8UEsyyXyWTrBQGzgnfgumfmBRXVMqQzQTO5YF5wcx4o5Nm/TTNssaNlf8wXwI
hI/CzRhu8UBYLAFO+zNoyPrpo3fuBAgiX4gls/eXOigYWDMWxvAnh8+Zfssw6Y9J
MLEcZehe2zuXeE/PV9xwtSBs+9G6avrn7PcQLqob+G30yTW+JBIBuYv6ah857Mda
KFpWxEsZBUgPhT02e3SLrKhoHCyeKDkbw0EtADdPrwnXCW+g3cFTlQN/lTwbL5b+
S/DAFUI/WwEAmWiE2tRv6OiIYJQVrq0fM+j93tipNeknc/NxQj2nblXlzsAqWgMp
XY+E/COJTiMiwuauw7IipXxHtl5rOWHAB8vhxOkKtwBHO4VU+cieyg7BQaBuNTCC
vQFWajquOnS6iJdZjzDETi6byqUUbNwLQWE5y18gy5ijphx3cIUSeLgGur+50dkV
yGJeCzWXhSAxFoF7mN4kz0FtzGQVIKeA3buWhbrOITjuBjZ+i7EyriyZcHA+aNSe
0/5JDHUmNge2VESKxPK5lXIY77mzdYGicOyXjmjQhvY7orv05IVWV17Hr/WeaojP
3gxqJsWTjaz7jidmexApAPas/5nqo+wEMotw1Eg4IvEJIrFx6BfhNXh5gAescmle
n7ZZCGLpoZoQQQI7GVRTXviu5bT5/w8jPtMd+zdBx58hsQOgpkaregQ1yavA8X+r
y4UVnSB2qTjDIjgGyCQdG2YfLL6yw4ug+k3FSs/4UIfuyEu6B36slfqpaX46cpv2
LFkg/4wixvSEgxm5AM3vDiUjYVFgvqs68foy62LUHCeQXF7r2EgWe/UMvPUFIuvM
jjwaUXKVhReGYkVUG1w4EXa6Znf/RBt3np8ggrirIuqa0sWjw4Ussi4KEBmWWuKM
60DpUPM/hYEo81siCiHq+L/s+/COY7nv5f/GwBtNmQOBkn6lS2AUsYCwR18FPr6B
K6MtTaBybeBGIh0aoync9pdOgxOivlTZsexvdNEpAGE7cDfa8SUgROaH4koQkKV1
PYgpBv4C6CK978fXbvV9QnveolVnIAy4PKXrfuRCiZbbA3Em5YWpH25ApjWj6Bu+
dd6tnuFscUbLbift1j2UnRhqwU4MQSWz8k9xvOUJ9HZu2SfQlu7PwIYI7g6hTcJx
104GS/iylAvUTSJ2S8zMKs0fQYlnl6E65vgmZlMR2/aHoeH3G4whfTnCqN9I8q1m
f8MfhOVV4eEO1OCc0P33ExFuH/mlVM1/EX2GpAPSmyggtmxYiYzXOj2hWEeqhhE/
9F8OPjx2pjwt8/XcWfzUd34nEusJAsXjQhNxFKML7h9hLmpQgqh/36iPrKuAtTzh
foKHtcym+NhfOe8cpIDnPwXmZoVTXNzea2aQDj7zP23hIljR3QP6qnZA8sBGO4uP
HmE++wLXaxk3eP7D0h1DFUvEzKbOcNotSpoyornk58cffEU8hTPE6gh8RrF0/72r
PiEpfQsAuqBr9v25XngjJ3Cr3NER3W5oOFTJOCw37Od+mtJBN5XOsYlVm0zUu1zC
swLHQNlGJi2h+FulE26bfNpxLnBZXhowy/70cw/zXL+xS89poggDdoYVwMigcheM
p1zdt8XH5etzGV2LVQhL8D8KLI85LM1y/wL+b7cX7pidbHL5PU9v/5hlZzq4pteN
blxQYtVUtdHbUMACo3AIrrFQNT+XofaJS1K8A27FPHsfY47cvmH4+tEYsdN1c6NF
9w61aQzzhs209Jrcb9fmCFs1P8T0pWPE6+p1u8npVjNQ0MIUBK5da28gf0RZk1PV
NzIk3oyccHVbyNKY5aaC9QhTTBTLCG/Hx8LMVlYeTIzO2EmzT+k9hE70zXA3r6Pm
KAzZHhkskIAafmE71TO6nAAg8V0UDNYhM/vkePSD//HU+Cji/dKU1N0HWslpPHWR
YqRBSLOAtPOh/pzkFD73sTPQu72M+NaHFX4rvVGDfdJEFYqHL312gHJl9/I+htnp
TYKsPAZjmBzpyEKSKEqQpEapqso1Z503UzR5IODoOdcHyZyPcuwQp+YwZad4H2V7
VPXpEQtnzTd6rq9JA+V9RBN8/9mYSZ5h232LYuYTT/vNnoLDgyx2bjhYq8Hj3J8T
tD5pPH1I3HzzjjmggZl9lMwpYz2hAMIFP6AIfpZTzfrThpNYLHjyk7X8MbP7VkQC
wztE8S6qcXUIcJnst3a73cFPMeIZ55pRihDOUzEywiLhwoBasC5h4PRsXYw0/cQ1
Sj/gEgGTzMrXSjzMmRf2VJWeXoyOXFO4yUZLL1rawVt0muFNd1JiRaBjjqUty3w9
mAjUALcXrJCJdmNQ97y5FSDzX5EALsooWBypX0NsIli5POis7KbupAuEUyUIzQ/w
zZoHt7Q0raF3FWz+ZvOaQuZvkKfZIxQ4rlMVyoaJ76W3l6LcBU+m8VXhdH/3BHEC
CZtYxEqbBU57FgXUp3YzlcUch+upPQsBbLz29xJrZvdgNeZZMn4OcQ7Y1+B13Vgl
UNnMvjdcEqe3kB4hJEXX8CPCSN9gB7ooHddgvR6THZ6UCkuoYlyzBJxkptIbIpRz
4FeFQtgBEWKWdhBG1YS0ID/wdlE4HwB8kxobQUjri62hdnO4PU9BLloNg292qTkJ
VDjGdVp19Vw0JE6Fbpxdh9RhZQ2EFw9UXaU1sySj34f94DnUMx6pXowm5oYNvKO6
g1XW6spxJphZtxh2RWXNPYGmfQTPF759IjE5Ps4KIqfBOpFZARfCMmOF7xPFEnxB
KIhZgYE7QKVwxMArDrSzlSkEjCW6KMl74Z0blz4GVllrS92W6bbeXj7bWdZyIaLu
9S3HHtHrwNN0ZNLVz4lSjlTuC546xYpqxB0PtRcvQUMTCAi4kftFOePHTC0FK4Cw
djPTuSB/LpZDmTT0hqWdxpp5Bg98hEOFz6NdantE+xGTQdTopL9C2Quak2um2h6o
HSikq2NEPAvHrZkdLtZ1JHuUHvLJGNJKXV6bSse1cWjdWeX2nV5E90MuFUm1gYBn
4Ts4a2k5Aw3CfSBaiVX5aow2eRhrFkaTiE2gLBCyPg/pt8dY9L+cqNLlOuUhWN2A
oVAOh0oOHdL29/nXjFGF7JlNX0CM/L3x0DomR/CIDeJj21d0G82r86zt+Qa+2Fw4
05TFXVL5IZTu/N6SXIjxJWpdEn8Jszo1+cK/nnmQ5JDiNQKe5FVvz27xbyj5oPbR
nsPE7eATc8AA+CiVqPcCB4tV2iXkPiHBs914AIOZNvjTWcD4xFYrqtMK3W6EbG1D
RqBZjUIbYMdxCi12KQgCoUBM1fgjDWUMps4C/Mvf+Gt78s+4Vc+GHckkJuK9fmNn
VNKjwxmIlwbQyhU5LteY9+ZctFYNRQoAouD5j3Objk7lI1KBaOfDl3sZQtZcWDO+
xlPcvGAzzm0ePxXrLPS7DhVItc/+WdIzwg1OPk5gRj3YGZqUZmf1mA6WGMMyoxAn
wvfR2s6snIGE5PiKCckMDjUozw9RDxI7t9zc12mvdCTqTvTEiavlhvWzoPa06aUm
Jo4tmldL8yzqYW8DA1iYrOd5viKos/0SdFX6E3jqu9bSySwVz0TIRIywQWJtnenI
w40+WNpFKcNJlwfQPkdc4MTtROMQ4KmtQkzQS69uTUsspbc0YWPfla9OF0G6o1G8
m+IpkbqkYnz/4ztJWc32zCKefkTkekDsABgrJvndBJs4L96gQCLOlfb6naA/7LHS
bOcntHK44UQC00WG54032gyZj3L88Q+iWftl7OW6KpSWNl20WH6altcpBRJoED3p
lmwSCxUFv8+F59Sq6k//N5ByolOcsYBclKuHXGERcwRJAJSfP+fDhjDSYF15Iqdf
5kdxfTODZMe7JtU7MKfSrNDVlo2zyASY3hh8r2RLNFn0ymFC2o3JuFr6eCQhCQis
I9T255fdVuJo0YEhS6kBdWJf8T1JtJmAoJnVVrXCIWYCxkKp3k0NEtctuoTrLFdk
4quNZkRPv85TIeho3sd5RJCMNDL1ZOePapPyTURzaSGQoBFQNaXqBAtHvjpD269W
jBRTQ0wcn9JT9aoZ226UQ+MmXVrYzaBWFsul6+nIsy14CcEmCSG0fYL0ZjsownCk
V938bJDUtIAqdlscYO8TZgwcto7anCWW90rBGmI9LroUngBpGJ6aU8w/4c/MQnBi
EpzhPW6JvU4EnsDh7HPPjK+hES/YWdfW7Td0jB34iS0HcyAnEpUtPh/ZTgKZnT9/
TFjgXY4mhC764g26MHhHOAZSH+ZEBvl7XntdaQGEUl0uQKs54oHhODjXxXWbCXK7
q8f8xSpegNST9Iq1a3FEpSdR5mOoTOudkKZ7PupNd7AdGAwiaRs4zYbdP9E4Vvtf
bVLISM4AIlcON9ypOywGK3CedQtH9yXIA6D4ZWh6xe3Ob4UeJ6QK/FsPh9XlzFdj
MtZt4y2AvtFAUOD5ikmxrIkRBRScP+1rIGYa3VXb0hmJuag8muQOHFqm6NefFNOU
6HedOtR9EWvgYhPyVngkj954C0VsAk1hLWtfs5G0EYWpXZPUpL2ZiS4Yp6I9vIjH
+g9px+e3xvqLJ0Vb7TprERskxm+3UzYvfoBpsYhQhTTRJsIIkMCBS0QRJUlZtMH/
+fWLQpgbxJ12hW+H5nXZpAnC9p0lrYDCIwmVn6kQ1o/JJcKIQjtEH20vcmOvytlr
MrC7sp1nDypoop9qfNoaEqXg5wh07zBTD8fujY7IyVs1SghUaHK054wURBJuECzg
CrItX+zdXUXK7xUNrAf+E/Bj8Yy+B5ov/I4OqtoS+Id676Fc3j4uVDEZahfhHR08
CjzAunlz49kSqu/E0jyoLF3nCKMkjwnayiEnqUrv724LIHYqaexhhFOA8nOor4Pz
DOGVZOS8SZ2OO49lwyMx+rcHrwJNyAMShvGG+UzFgkGsXW7Me6lTjpg5actcU8nH
SFFLBCeD/569ecY/a6vZ/bZQBadh11j9yyQQU7pnCglRTNfwKXyqLMJtM/Ob3FRb
4+EfFOfqxTx/SxhpeivT9kHNC++MAnHN1oUz4pguZSWSN/nXDw+NOPbEIsK5mlqt
PcWplmQn3Wab8pOtsIs7u3D6agDee0xUGYiQHUXOpYh03cgpY1+fXGC+PbxWVq/G
e3cF2coXxkZp95IaMqZvI6jIH0bl8TMu6YN69mVCZY5a3NnYlOM6Q4ubhtgqV4Ta
1S3VOnTjhidmlORyo7FcWEyoOjcZz8L27BiSJ/secudaRuxltXR6XvpshvkflExa
2jSSxXh1KrnNJIP+8uLeBjCT6i1fSYuQkJD44iO4We1uroC2CI5x6GdcC2JTVOO/
V+BIQzKmemgrRXtq3Gzkpeq5X28cw1q44brEnFH/DdVCUzWaPJF5i2+Lvq25+/QF
rvjroB7Zp73pULeQ5XU27lyu68OFBh5diX3txN0HunBjm8NGErxjsp+2Q2rYzeCL
etEJI6/LMI5dKMxc7++AVjmqzm86/JmvhU620GRuIkMf56JB9yeDhioe8yk/l9+2
Zqby96UakgrCVakVAaegPgE9AKWAgU2GMfVCMJ5XkG1PJQ4L+Ep4Rdh5/g2UTAT5
n/+6zjv2iAgbAHtZg+xpzOp8Cgr3wAWvl1mPJvavj6Q0VHROjFpffh/+CopKCyki
F0+aIwKKrx6EY8ncwfD4E9t+BjfNUVRzwTHTr0P+4h2sUhB5LmxUSAnkWSRWbP2u
axkJtAQQIxq5ilzQW3X/0liFxTh8g3FEsjiFg0YWBMibj3bYPd04AvGzfoDWYJcP
k56IRnTag2uB3MNmWqnRkvVcAqnng/2n7GH72Pk6BW52hRNVCtjX6/xkQR3VtHu+
Ei2u44Ovdb8Z9FRj1a73oN3lGDVV80k9Cj3VKRlp1c5JJrpvSp3jChKLpawgLSq+
a9mMoHYfK86chOtzVAA8aIlRu6xLRf9TUoY93p4h4yp3UbUKfStfig32AUuieg3/
1f940Ec+pScuQ1j1jXm3Fgxc4jJnS5ZYOl0CiXVw7HHgAHrlvxel6wBR5dz8iLaI
hiA21ntUtibJCcfp3v5DrBei8vqwYwVTA+9GrwnUYpxbm0f7NZ3aarui2J26Fj3U
3YBi2p5OotmiOsp01gwxcO4cKw7wutgT/BKcL3S4d4naJ/Va7DBEyJkjbu6/K03f
8sRzpQr2gJuVszAulYflu2qcoVsga4xpIabuN6iZMbhbta3u8dJJu3taxENQGlJL
RWT08v+JpQhdMul38YqYQ7o2KOzPh4ZNQAprBx5a9lPdK5CfQrs29Iz3LhWiQMxe
uJkIgYv7/7W1lnAzg7IONmdsY23Hv9/dPyGmTYGZQXPc9sRoy+6IcnzQQnSSw6s6
Ljk27dNa40DngN8nLbThK2fd+1azRiVy8cFgkhw569FWfCTyzMF31kpj+CC3Qtkl
KJK7goa0Lhi5cxd2n/pkBcaVEEDVbCR2+uIBV7VMxDDR+3W5WNoBdH/vW5AaaPpg
BfpBCIhA38lsqz3/zZDSv32gj0+v4Lw1/4toqcifS7eme7KRZqqdgw8BlMyWCcen
uyxXfofHqPWcdQlyJCnB/rJegGQf6M5V2ZjKpJx5mNxBECcci+zaMMNjorgX3deO
UlZ5REbVVySKfQY72NslpzOrH94EcGF7GSZdiRYKJoYtFhwTZtmPg+BLcQeZD89/
hwaGwuff+YxPBjZz2NeLLupMF67hY08Y3yE56HxEIudG5d4EuYHAxt3m6Ztf2qzs
QokresoyAUVw0LFoUri1Yc+VYwki3C5OBSgWITCBb7DiWC6XUEoagnnIRhO0q3j4
Ea0IpKHLpkiwVbK8RgBl4B1xL6VLz2JuQokzsW4dGk18ILBbXMxEPbUb36rILU0p
jI94mVVXxMSkDuhZPFGPd/Kdoxc8gx3twv6VECmvqS3vlWkvKACUcIZUf958uW+S
BZE5oKIs5MiDyCRgoM4oIFZg4YrIb2O1BDMbvXFCQ893cU52hH86ziLIBnB8zFPB
dMGXoo5zqpKYu3LUlMUgd5XTBrarYQE6pHCUNyaGctBljMUQw6lUOi/7lGghmRoc
eG3L7nI/yHCO9tFMsKWC7cSS5rFrckZur1ybsxsVD9OuKUcAFLe8up/V9cf/6cll
7I97iAp5iMaRR5FVukZfXXODJ+VxY1X7pRr05B/lnZl+HL/CnXhixJkCDm3JHcLy
AIzUb7VVnN1HfUfrhbPLq633ueBEARm4YaqQEgzTCwoW3vp1XraMF8GUV2vU21tX
zsTqMVKR3q/dbaJE6CsCZw4t/OLI0RLwk+PJaRfwiCJ0hqBhjGKqA4Xwz3xweP3G
piPi2pe1UuDIYaXkZqjYSR2PebyWMvWxFKCHi9CZpKZiKRbmX/FnrkmQ7QA1s8PR
61LKfsz5XRg+zzTAfWkpR0TDaskRs74adNowuQuSgvwlVS5FyP/JXP+wYBrQhikC
T+PNbG0B8Kv1h0Pviei0A8VXiO0X95oEVCHpkFgnsUw0uqtTZQvadeWUkrjxs7w3
qZCzQiXTjcnH4UwYa35fmrOqWJdLubVMxELlYQpUgxeHISyvLmIxXLDlB9sSsK6L
lT1rrdMdOAU/woIdFqkkImirhaRg4eeb0W4U7XDlnWQFVy2aMUCfO/36ENFog5l5
OBac1ohVJ3nbZ/y56x0YBaCJXtnZ6Aq1b6vhdFwTLXJ58PMeBo7YkxeHS1m+ol10
2tezRYl0KINueScVXCorFROkCN7eEvbPIT4jKkib8/JQR7jtOpeW0q96Of204pRX
PXGuxhapX+exGGmWDqwp+U20YDa7UaYtE12mEyJq3JHUNjdHF1+Adwi/1h/wwgeM
XHq95dlz54Ykr20Yt8mgr0l263WzM2DvaJg81G51XqV3OD+RMN/0LyTdCzeDoVWN
ewhb1fqlcBVystAJQQOLjKUYLegDfSi1amnCUSceEsAhV8qInv2cHzsTG+FOxLc0
F4ucGfSlAO5b+47sro/41/7bkhyLKFaqmFWMTkbwcvXMU2AUTngKoQEuQ6lqo9ZC
FtNhKGfntKEaX7/R+G6BEIKGLFUM74TqYcbqizaHpl64nAeKLw+Pxjfs+cHyU9+8
WCDyCbSIpU4L588Uf2441sQNyjIhLFcbTr55ToJv9yPa8jjZZ/VgpUrx5aw+9fED
r6vc1qxPNAJQkpLgiUXKM1fS/1X12WF9N4HQCc6C8wOgChlnG6AL/ci3ovs11agZ
Mi2KUq9WEyc4CtCVtJNjlvBLezg8tLEjcVJgbWlY2XFwE5yZqmqDdQjh8AqpQNfj
fxwBooEg9jVpin1yfbu7r9jXk6EEadsvE4ZPZWE8+aSj16hJf3FDneqeg/U/EPzR
gLPgA2HAixoAC22J77lt8jcGoGPtCMEXuz3+SxQ31jyJRTmp7ildYWRh0tWlvIuS
iAgcf9enZ2lRj9rlYgfemq7VfhIJwSYR1QrSUhGz9sRZNeG2LQQQUAugX/fjrKu5
wzDOU72Xfcl/Mk4221d7Py4lV1oiiWPlAJZowDKSVyfZbJMKOHXb+pd4CEqEWt3Q
2hJfdw3xpqtZWjyjZRjWhtkjJY7YQlaGQvhiWeJu3G3Kx+M5/eiit9GWpR7iZ473
f22Sym00eRHXTsV/eh8hfdLqdE3NNvq9MArqzYcReDhqnNURX52TtE9TMG0Lnc1l
H6YCv6CMfTmfAlDzD+dMffxQEKU+3Fm9UGfKI7nzfd9emfFJ97KejUdh4Sw4Xqfe
JubPdejPYUuQk1dJafexfB6g9kpWZekP1loG/M2L7FYck7CI6erFP1FZpWRp34KR
GdyN91HUAGwXbc+qMmigFCUz+Znp+h4+vQsjrC5HEe2SeaGHzw68kqFyyDOh911Z
+F02DjypbM1J8JdS54X62x6G1Hf27dAYjLeA8tnm5eh/z7ewcf2yscXoGv7iALjU
RJlU7VJjUmrOMbncEw0DG9VuuMBjBphnTH3Y/gzio/p+X5TsKBdUTOJOnYeUKQi7
dcy/mvLHTI1WLQ4mMqztqF6IE+nXCRT5L1QFZ70oxArm72QMdkRrmvQoHApA5OUm
GKaKJXQGWHQiOTyGQzlMVXtd79kq2QNieR1dpkn/IOnHvx2qkiuZdODz8pgWOOkZ
7s/VK5otlVXOCnTmb60+j/c7pnL8kl1VWnOZulyqK7+1Dfz0t6fZfD/wC1f8WPwT
aU9RZCUqcpR9FyN1r8I2FtvHWYcIKJKvQGXsITkWkVK6Psx+QY8b6uznfQWmwW/X
r9ksdGHOxfIes4kV74ZEldC3WhqkJQdrIRleNaneh0KQoxsxBt8o6R9LgUh/dhqY
YkoEIws7EmPse0IYnuZkviTlD3Xa37xJpAxvg9pGCOqggzU4ZFMb/OJGwblx7wVV
CipRlIsOprV3yzraAqvM/TRcAdmW8H6mDaPdGJGu1LeBrI1Dl0evUwdOdBbC8RhL
ml+NZzQan9Tfhpsb78tU3hxJ3/mjtIvdN5gXvgl+yDvrZRhZuRqARt9j1NaZ6eO+
Z9xiXW3E43KmVcGq0PzLE3KoU48yv5zqG8nabQQhnvjv5IJvimBMlBYz41QeHBZE
5PUKMLCwbrfAY/B06j0OqCTsWG6aeth6HI0ZO8eRo8BCiSsMesNYNf/lEItQcUuJ
zvcR15Hc0h9yA0kuWyy4HoCl460konqz8Wn6mkiIgTZ11ouRH2dZxbVniczjWtxJ
fy+vxg5tyV35+d1FnH2o9de62bXVgAvGw/uUOpSAhzdbnvwK2rDVZKBZWLDrK5eX
kcPOyWfpDlyJ7p7M0ZOUH2zjXUBXmtSGZ5vbab1Brk5AaebPzA7dTyolMkRw2miG
k5qldhszakL6XBHBHU5/y+5MCGV//Jue5dZ0LHXm4CluzAtBDdGHv6nGwrf+HbPN
mGs8hbP3wkmQuotnA5bsnSVVQBVSd1oibwHTvoUj/haf/2xVMl6is4/vhya96Tl9
zejFA1jv1ldzCdnHda3RGh8APtPZeNwyJrrWaKfKX7D24luPYwsgUH559ArSWbsd
nJ/D4Rxse3Neysce3R/m4xOfArGnNVZP+jPzne65iRUO4ychbFOoA9wDHjHw4j7p
SQ+IU+AJEdqZTZKx6UgU0tEoeGO8o3YrqHphz4t4bSwnd66NlTWYXFxig5K1h7IV
yYiQEn4Ag28WnJPsnnkJfZmTr1BU//38UuoXaDiRF7kL6Uht7WxB2fO4hRhwUaZu
2zWzVXl4YAtw7B66vwqyhQMgjb5HBd1PoaPFISJZuu2A3eCW6j08LYOAcM1wLaW4
66vFrhkWb1lftnf3DNTNasY80s+8LRoHMh8uHtIEKze5HMEn0fjZZWDn3JWjE/s5
r5rLFOZwt/N/S9xG9MCr433YEODtEZZow74QK/7TWPLknlQY3KQayPKybBoI8En2
RC+lfbb7n7Hl157TBzE6uIqoONmNjAOfP6gpNFJIhkw15OxOiQC5hiNSVjKbYJ0u
vfFCiLdcZpcMdgY8mJhddH3ud0B9XjhYmdjluCVJ1IMHJS9+bBIO/rXdzdthDTbY
F3m+kNiTj9Ft3mVVqhOayS29P8/tKPTczH4zYX9+sQvtDKEeNPPxJNvSH/KcTKxe
NfAgN9ThKTy8+Ir4JdZSF80Hvg+mpQ+qxuny6QzJJc99BH+3zH68/D3ITCk1517P
evRaiK87DTyelodWbvsHRCV3gFPn2KIyyIPebT4jdEgzBh3W1IhKN1TRkTtFRfWM
h5nxBLDO7RNlZSiM00z5TDXb3jp6nh6RcPGwYnHOulVZYYzLk+FMFC4HYiJ5eX/0
hlOHbCN9gCMHWxEvcmtuDDoK4Qm1f8H32NEIKNP4IyAGt66oQ560cVplOoW9LjEv
2wLd5+oi66CNrHZ4kFYQudse+KhTjXt90T1mS5LYDVVos85xPXVcTogoh7cxHELZ
nTHO80OZ63KQg6Df2cVsCAjdKwVO45JNHhkmtQmpqOfSZzcDZkYMZ511sfcDARNg
tp3t6432Pk2oFWpvx28kBCeWeWnFM9TTn0PXCKOp0Kqk5f2Dh3f86xsDRmwUhm+f
BC3xKKWmHj7A55v2Mflp8hLNcToW8/Az34K5ZK5b8BuzDZhILk5N0fXYRR17KHYt
XmD65VvQUbvyLdBBw+EuotS6jTU6Cw7PJ6GfjnDHSOg9KWdACZiAQfWN1CR+O2Cw
wJNp9D6WG27fuyRyFGAX4eN4eT64krWtTH/35QE62mLamVMQUFV3UpI3fRMtN1+Y
dQK3yCYjA9Z/ldnXxfK9PWUncx3/hnpcnjwWhbCnagKKXAhxs7HqCTuFL2XQiVuy
m7lSKqFkmAv0+mFGVkeP5cS7AUpaiZ0oKMbTw2ax/KsBLRGwrEwSF3Q+r+eY1cT7
IKz2r0JBg5sS9DM+08OtwYvZ9sMmmkPYsuadBpMv9PhyPF0dOp6pIWBMtxd2/XeJ
BnOzuUrLzyUaS5AXqsoRnhEX4t3pKOlmIbF6yWJaB2WGsZvht9M1yzbbcpPFdsEv
0n6CNU7jaFbd1M8k0RrzjZ25FC8n+UZigNSUjedUi2JZjKqQ9A6JxC2yPlQvJDd5
PK0G8AjyNStNbIrSYlOghO+5cyEb/K9jVGXJvDAVc2Fss/su5iNxVkBGwzBWFfOl
3ewx85I+Rd/4t3/kVTqRzYh0gdDFxtxZLx5nLFD6SW1YIjXpGm+fq+L0OnvCLeZw
vD9s3Fo7ZbfIKsEfwPi1MJUgJG6sBE1pIz2ak2oVrvy1Qi5pEpbEfzu+BZ76VjP2
FMw33TNY8iwp5nRb6ucbvjizKf3HM3RYRrfDg1s342vH6EaRjDdlcQSWcxq0+oUJ
lDhVT60YxEUgfrIHly4W7rQvDTkAT+ChaeQv8auOGmiPdUM+ZHBKTTS5YTYaFBx9
t0nNaQY28gqu1L0aO0Mvql0mn4+fWMRLZdFgARUUw+nMP0iGj1Br+fakoK/A5Ukr
DiADjNibdOfmy3Qq/espq3DoIsCb+6LI90suPgx2EXz+zgXoOE+9JHW0iDQDXEEL
CnEM1wL6thQEMJTtu60G5fKIi5VLiC7TVMRFlvRNdmERyh09e1eL6s85AdKvC+Jh
QEZE5HzsP9l6otd9twFmfGV+Fjeyeq3U2Tv6TJGOekz1ujI4SJetujt3V/gzUDhH
myb0oigWIYtzV5ekRqBIykNzlRvxm/RNl6zigLdK3Lqpn3AUFClAxJC+hn06fC5x
CtEa+LmbWMJBk4bkqGuMupkJJMdU9d1fBoG+0tRCmVwYUjKscvNhyVEARVsxILRr
XuK+TxZCbwFxzRenzM1GgbjVdmau0RvdhKAw7FsPgTUg2wx+/1Pz4RZ15PLjZNb6
p4NRCYnJ5FtYt/DNjOzYSsYkI9LH7B/g4EN0rt4aBgVKDze8OWMiFI5hY/LtEt7h
0IgaVGinA4d+9fk6TfypiJOSs98qgU6TR3lRYns6qccflO2ZftqJOy04q5KPAcua
9OPr197XqfdDjm9w4gr9jdlCsAyeDKAGzJiBh7H8Yauz/usi9/EMd8XRXKklrfg4
HQM1S8N3FHMsAfhMglXOrDlKifnK7gRS1MFtVwsM43K8blpyuTbQTuu9Xu+2a/fZ
Uou3x2S197BmRmd4iN/shILt39ByUGS5jlcPGhsfg/eL17/iOdBn1MYpzFZodq+X
mgO8YtBRrueJpSETtC6JRHCLORLv+hQ9RZQ7xEYUcndaVBFZHpTZTACiNwN1B+8v
0vn/HaqyC+plswJgdk6CJyV3f1J4aZj0ytxUMsGpec03lobUmHAhj86fvR16V/Om
IBDKm3WgmlvhJtCfQ/925uiS4WcTIbUwmZdcHvAFvffbPkl6ukWHhfyl1tw6WoiH
+QrV/Grz9ySmaeH1VMJbAxborU+lsY4VlW94eCUb5tkYMWrC8ukFPOjqCMqoIcDR
OZgzmQgB3OsuMZMtBFdNeOeDVuTm/StLd0xkWo9E+7hyizNN7g+966JyfyYluB8U
LXgB5sc+W9GxLD/XWfUTo3YTxUJlnXYZdlFImX/tN2MiWheEjsJuEROFYZbls4fK
e5/VbmzRnCtNvcGumFG+9EjGa1iKWp2vcPnm0LHtEKalDNkMHZee6W9gI64d51qS
wBsF/9yWm3YyWi/5uHWEwtZ3lvJiITxfQmdO6Z2LTrecQT43LgM/o7c2A/14Rti1
nv4GI8h+eofQCaNExrFa9xVVcN1zEZKK5Gr3XcfijN3FRSkWcy5/nHCEvyqvJVum
Mvy1N4w0Rr0pR2WUZ5RbomM7DoFNzPEZBjQ73o+hvzmY5w+i2GgxCTnO1Gv1qoyq
ZxDmYDOr2ju3Wonb9HwQcfBLkHWJvh4YGp3asE6cp2tDM8CXI+j6DDUllGU6IASl
oW0VFiCE3hhscAGix0FQ+YZUg4z3hepuzgiVZPzy1pliXHpofh8NbedZGQkFtQqf
deluNZsy0mfd4mbkrU8n3xN6sRJPx/u6m8hpj19/iz0/roKhBfFBXSr86uOQd7D3
dw4lgThTs44YkjcumOTApHwctRT1gy2Xf6nGHr3sLjfeyl/3tZTwq4k/igi1kRyJ
LsJg0V9YlBCTcJsW4+wv/l/0jNSMtklUg+8wS+WRGTDWXN6pTHiGQs0Fjid5lJu2
FN7O3tHLER3rWZF2ICFyyOdAuuZO+e0C+wwHOpu+Ff4J/68P71L7kX9wGzFThdaP
v/ETXCcpQYZOuowvqZMsARYsRwUy46uCn3X9DS0cxwyQXBpL9tM/eMq2iDEv7o+n
AB0N1jNJWT+VITpNnbCdqV2BXkXZwuRS/Lpc+70mZv85D0rw0AUbfmqzp8bgIIGk
fd0XvEV3hXD4xDIfbWV+/2aUicM7b1y1ucBMkvG9R4Zwg3jED+7pyEyKnQ9ybCG/
oDLeUYjc7HQ6ye9A6M1lnJ7p7EyMxILMUE2uLvEK4MnMjCIIY5Uh2ElKf6vIImzg
gfNyqToNDrpoFSIae/6GmR+B1jEBmRToBk6Ikb6l73xKZjp3HkdwbjO9xOqcVqXG
+6jF6r1vs7bpCqOQnuwFVkDrl4Q6zJyP95R4Oqnf9oLv/WIxllIh7D99OwR0OVDX
7fa0aqMq2jQmmN7KfiHJbiLNchN7A2SqqKpBPTr1xxiWSV4rWk90Zd2xSY+f8eEG
ZRCt0WmAUqcsj6d4rI9+AQNpaij0BTjeKVuRc8macBkPWXWfcCKn4FVei511beiI
mqbCzpiFxCyszCTEfiuRWlQIABkrVaLfToBBDyGMLonBpuXhWOLbqKnx6p34AyPS
edJpYGYWMILl9qiDvegnlproZojecc/xdSGbrs00Qr8mIhf9ErF8FVAnxWP3MFaA
8YOjde74I36hp4DvrzxME2IGMMKCAHdCqvUHr6PUuWJwr8vqN1RrHhWLEn8oR3Y3
PX7fmPP5UvtH3gfr8EWOtv8cwIb8VTdJqoU7iefJfwWo9g+7Ud9bWrHAj8oz9LV+
lQ06/1LXkCBsnfrWlIsJHVArZTGoK2AR6Xqmu1hSH/qwo0SWwe/ecZAL6ey2MPyA
37vCsws3Hvqpyh71Jd8xm/9JCqAY589xzarRkakB+kICDuw3+/5POm0viS7VmL+0
kuodzwJseIrvSrsT24domNbQD/kngtMJY9+tN5amBRKuracIG7TDP2ihvPBussDI
YqZUom0FzID5p6W/BCBeWso+PKTIvJjBlRydsXe/K6qcnoQwZqKtztRX3XeL8thc
YCAbxIu3PRMxK9P9SjbgfAJhCFfU0aOxHI7gaJOcqBPWdYFW+5GI6jW8TlVQn/rz
7KZy6RbeO5wX2a+b3w7SAV0mWZYae28LM0j4zEIaFWaa+gmi6N9A6lTUBGaD1hQ9
kKZnJm6kkSDteAv2ifMGQVwDpOmhGiXb7EHt5oPsdh92p/wy2P9hdRmQUgyv7txp
3xAUWmOSoPnHyt0P31bMOUXpBxn+N0Ea6nCyXzeB8ObbsibYHQIajzBbKDnN70Td
mAfrJRd8qZky2Jna9gFffzi64CHeqdYD8VTajylEkt22/1Fr4GU0vhHYY+0CruH5
zaHj2Xu/vps2AM8FbrqjoKKZDG0xzg00uFmYrf1zs2+2oFNvug000ZTIzgZ9L+Pg
JlhRBBa2u/dHnIXxsU6XwLMDnLkkm8bTZUJG/pRkxO8XHT8vdCxaXvYD2PNbQBq9
ykEYyFKLe1Qa6+gu74isnFf+jom0XYP+T9XqFI3zQYX5wJ1IGwMZCpCzS+rIWeW3
C2Q3zI75OMl2O5PHZa2vE6u/Zz5yo6qToSbc++y6mRW6wW7Qrts/rSGYyIqaA57C
7H9rHSlw/4ScHK2Vtrs9iUdf71U7fJwf1/iRtT409xUs+8pxZV0KS/8VPCXg+a8l
ZKlLj1AlyaqqfoapkvqPSkRAz4meh2a1/6XgeyQZEuEGoRwLUtXW9kekbtkBndj4
bxFUDos6MVHn91iUfcR5QPbEEZGYuoqwUn//FoQoGkqx6g6Untk1ayhvRk9thR5b
CpGi8ctoJd+kmTviDZaAqP2gsq1st2dsLBbdq5mXYJ45+5d3/HigtEdceHCWMc0S
8hOO/JqbEEx6XL7EBDUS+ffGF/8r2JSgINcwzKgJMIfrZdulroyYDor0Eyjx66WT
NP7vw+lC/PUU1/Y5C3tty8cxQXrGzmMQKvj2ILxwMhFa07cbTgHH86sR/BxTxusv
o98QXEOT3TlmfDlwiqGHHpRwtsuwWdB4AowBaOcDDxLwW1Gr0sxe+N80bQ93l/sF
yLj0PGm8PgVJhVBFWy9SY3WlOdERi+DhVoaJPvg73Ib2AitHjNUmEgn3ebaiAAUJ
01jtsu65El204b/h/elQ2GzdbWMyw4eUXpoijZS3LKqvILeI94IhSgc/JhTN36SZ
Ye3Vl0YJY01FGM3kdgHt+4DtLXjZZSuQaWPmRZtulbwHEziEwLZEZy+Ojgol6IB/
RSkdih8yz3mEkoK+hjGO9ZcN0xy32A5rtiYX+TehEybykCXnqGvPCMrnN2CJ1C4H
UjPdAxz2GgFmu1geLEEqqA8tC0XHNj2zrwA9RctBmmhQZ0X56v6x2/9yrUEBJLh1
aH0Rb300Flos3t/N/p9oKkL2+rA9q2sknzEK/t56CoGpGtdne6W4HIqrHsteB8ON
GMbQX959H7mkowBNG4bW2yUf6cAtrc08VDsCPU9EXwTUMJyrb+V3hwuco3zGdEW+
RFtbIuHCR4XvEkzLSNNc8HnVnz6LNCMjWbUGYZ+/kO0VhM3bksd+AEtN+viPpgTj
/OFQSP8AuXQWVxDcyMvdx1bAbKHiRuSRm4g+OykDt3/cZ37zmCzxXgxTGICxAZlz
z47dVOlYJKo9SP8QBL93+w7ZznDEc6yCdoWEtxu+4ou1VrQdlWLAgNAzYVTSY/PZ
sM9FnmFtVHkmIcc1ApI0oSH7gZhbrv3+tcR1L8TzowBxCEhzYcvAd+zJfKJRPymU
h97zh1Z/Y934WUqCLbAor6A9rXWSpQd8DgcY/c1ip8x4rMlB3M8hOA7fo72olaj1
uOcgQqxJB3fO3y8ImIS8G0l4lzx0Yr//W3+6tffXU6MjA7NLK++TbIlFS8WVrzCi
T3WxB38yn/zm7lUYAiVcMeHnodwjUzQtaVJs6dglkQ5Jqs/X9kpT28yFSyTlk1+Z
+fTI2LSoMzood47EkH4NiyzjhnZOim/9cUUCbB9Ksi2SvaWV88+g1QCr3/JAq82E
f6WEhwkKkessHegNfa6MhiSb3eD0o/7TVF8xWqwPVeuJ3aDwfJslXaw6U0M/5mME
H1AU5CJZtRQbSlbeg3w4yBm2uSjtZfIGt2/RjSOYfiKf1hiTvJcMG2INxvzEQeTo
mNdqFSgLKnQ/vEfrMJw4vby6/w9kwR5+vlQ+T9Ky3o5DNXwT+ZJaZrP2Rmic71d8
8icw8x7lU6nXuF3mwgMzx61pgpfWJyI/jssbnDHtjSre1+CcdXNyxDGGF3xG2JGF
tILIIUwvP1D0BvMKswN0IB5kpW/j6oXghyJf14cWbfnjk9UyvfJHijk8PahrWUli
ucWkA9MKDPr+47L6EhIzAB/W06N/dP88E1GgypuzXUzO9EKzc0BEF1EwhCuIduWp
fNaFSVa451uyxJF+9ZGpb3nPFmRttkW+KC3dbH0R9l43bppNrUERzlwh7h40IzkU
6HykPquB1bFWAkX1lQrEGuFzwfLi8CV6TpVL7Rs7s5Ma4AkP5qIpu56v0l9BTOj9
+UEjPXoLNlF3aDtSCHkiUZBFEVB3stpkeSgSSC3U8JidmwPxH+hQLmOWEAUuZfJk
6M9MzFEURCI/DVc+asKhWyOaKJRrfE53juJie0mknw719S6tCWJ8M9jxGKqEgY25
2U9WiWozYQNrNumiOgHVTMJshSibBKT+/DlDx2aHGR+u/k+Zi/MtFlXTNG2OLEnW
uiOD79nTPbd95NgXJG/HZk6nzjC23AEWC1yhB4T1rxJfX+dVBsd5fkEJFVXdPeDz
+6Xt274pp1zq5NJhfgkwHRMSuebknR81UiaFhXs2JuQEm1pPAB0NoR428zP7t8MD
95btqKMytuerVKt+bGzV2enuPcwoVbC+XSF7oSEP7kPuWmGB5Qs5b+e0FPIhgGZs
0hu5yzKaQJ0qHim9MakLBJbFh2t5BfOjp0KFFtRdCaTjQpGQwfi8i3CJ3dGjQwba
qM9xs3D3RgWhx/z/io98q+bPalY3N17cM2Z7fI61ooyFLK9oT21k29I1HEfVdcu9
ABK04YfusPvYgK536V/S99MnwOxcUoRGk1fmbz3OsBys0iOr5RVYFjgDNtVTjh7a
A874NGbXZEZEUZRdfzehhb8+u1VvmuDf9cYsMKoa0Yy7MbJ6ToZruB4jQWK5UuPh
GxDnDtKDyDxU0WXKSWldhNlXIJ2ooIZkCQexl6c3uNAd3KStj8pIHtK3aYtqL4nT
+YtIHBD6MqtZIBIZzv93NLFyZ8kLuufQG0JUE8NWgcf3gAlOelMZLSmLgfzRrPPr
O965382UFUfVSUBhKL46WEwH/7TdSqjGFyOIQcgS0+Oj3yoNytmTNdnu5AsV03Wu
AOJ/JdWL1mHSeahPCDEQQmG7BaM5OqBJ20+dLj5h1dkkk69To3IZgUqmthJ1Wgrz
x0OmAZxAqSpN4quGf1SfdrDpSml1RtbacX1ephengKJFIuwQD5oEM2ey3cuuwhCi
GbNj2wsyQzpROl9tXNGbBA==
`protect END_PROTECTED
