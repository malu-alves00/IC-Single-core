`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JV4k9c77PcbIb0jz5idiTbbtVuKNiJI8oHcaZ2mYbZRGV/th4h9x7031hrOxKfhj
s+x6Ghs5XRpe3GSVCMm8MgQWwtNnN94bjsdoFBDIz5t9R5KlIPIUHNQm9v8XLB28
MwEKYlKRoXTDAe33DIHbWi5mVnX/EzIf8d4W1CMe0HxczJ0R+jze8lPkqCASFjiD
1OxG3fnJk/W1TTQcTIvFm0zqAkKfjkRdMOIDG4pGNmms8OFGqSXmg3doLOS78xye
RqBOUbvopvM6p9adGE9P/Y8+GyuhbHa4JaWjURNVfIY7n/lC37HcCyjNHWSm0oiu
5KHI1roTEGdki/8nS5eeksthT4+bWUg/6PlwwabioCOJUhEJJJmMQZtgjjhZvbra
7xTNVYV245P+q5+GgaSXwN0BZ/WGejeWWFbyP9YqF2QswPzMwdNx7V96WDKBS6XA
j+2hgHSl8AseGVuYhP+RO8O7GCsQ8G9C/GdtjQS92w7g+6/CD7uVWviTUe9GyH4m
BZ3evmRBvHNZ1j2ajltzLcKY0QZTsmib4H9dX/EyI3i6gWwP3diDK0yU5bqr3vPo
VUPAGC5fl9KjT7utbPNB+PQbuUMxK9IuehyO0cjEpdsmogCV9uK9RZFb6O1buCoN
3DO/I1RCBzhXEI9+kwusNlltnYHLvhtavfoiVqkbUZnJ9OCHlIUc7bFB6JASDton
4zNz6VIFRB7TYHcPA/vg3AU4z0rJcMZl0dNOCkxKQ5nldFwPsOyA++vpzj7cxZ2Y
n7dPM5iWEEhbgjmmrqunzSVW/2k3bymUU+A/FAFw/BOgvyeMlPmr5ZrO39MbjpEE
9dpbW5/i4Xs22mdgCXF8O5L+JI1HDql6ev2MEqezhatJQhZP53fpxGfYy/5IAc4M
/e8qSqGlad2XYa1R/6VjT875cDIdlN65vWJJlTb0nak0VpSjyGmfGbu/5KWex2s1
eHrS3D+22Beg4vGBWi+a3OTC0fpc6N+vj12fSUm8y8Nf0wB4ZeBr5zAtFET8n0CA
7AggyGbbP9DCiv3esP05Hvvk85SJifSS7FLzpwF4SOxuVgmJ0z4H2JK8F/MffjUd
sG/A6yiBo+bChiO7G/LPaSuvjYvsFOZFQjEaccMU9DlvLiTPtbcWST7aMSFCdfs/
7xEA0NGYGwLSVtEodjaesSaRbK08sSNppxRQPQ+Jesy4P4WEw0CstCPjxEYwMmZX
ZubYAhYjyaQLIPYLWn8yRDybMjHrT00qiHVQ4SNOLEaKxD6Bi9N5OfeXC4+1IT0i
EEhjF1y73ChQ3WLSWdre/jGYgytZz8bvApO44E/Mbtv92GX+fcz2FleYojz8qjSV
boG+lSPr9qGhnCYlPdhr5yJSh5MBY1m6jubCw3jma5Foavz58Q9geFZJZj3x3+kt
nr0i0SrYG4MHXvv62oSmuXsFGsR5XR/mScx1golmvUMGDmRqe8gV3zKC7W28X9iY
BD9QybETuTI5kU+wX0nfdsq+xIGwawfMOghxQuIPsYTzgLw2vAlSCY6vDdDqO0fL
Q6JD133KBO7b2EgOczeO80RbmN4+DfPMaiSN+mO2s+FztZrpx0IrhNtJBur11vnW
bI6gYCIWW4DGXT2jaJapp043OKGTusLYFQ4O+ctonHY5S4xZ70UOM7GQmfNwCPcw
ZGuaXGozcGl/0UP50kE0/AlM6OZ6M9mNmM2XvYzD/RW3H4XTAmAU74u73spfon06
HhIHTlxsoaZ4CthS1WTgZ4avHz6UG2KHAWQYE3fIb2L30pI74iPR+HcbQ9QgYR/m
MH37IAmXizYK2VMZ/vCOBT9fx1HGjpvkCFJ7cgPvG9EfbEOPsP673MKwHgbaefjd
xHjcvDY9wQPLymv9z3P8IQgcihiHGXiB+2I2/I3zNBufjCsL4cDDVgkpS15LT8pt
rl2LAoKwMhlE+vBa/xPWy1xisX61ot68C+cJHmjRwVTk2XyGIBDZDpdq5FSDXdwi
qXY6s2Jnj9bLGUvpdSqnSsINTO8QFNgNWfUaMpjD4frBXokYL2COHVMJGXOq/Kn3
BG6ABRBfd7K4m3IpEJ2gVSgI6S+NZPF8tVgPCMNDD04U1sU9r+c8e3gNtAgK1mbp
JQiknkCAoG/bLUe3LzDq/XpeuTfZ4u7f9MYogk3rl2VxYfxGKQ4bQoWexq2ihSGh
UqducK9OPfUY3yLGZhoStDr6JggPhWmMz+THcMBG3jSOdFMwUNFxxXjX5jauRtU/
WIRoPuKRi+XZhGvz/tyLzFSZvhU2R/TAXFectI9jUu4zTAbNmNRlD2kO09cARIyZ
MeyfQYVzVjSv0L/WVxmTP7ppp8UHYamN+DuHDnNMP3LE8Xb5bvdr6ViS55qs5gRa
1ApO8xXhBjxaQ28+IpUymV/MkmtsEjITXSp4TATGNJ34/6VBnAaM06uUrZe50QCn
d78D5gMTqnXDK/8+RH6TMQ==
`protect END_PROTECTED
