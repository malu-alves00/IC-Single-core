`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+G2nUo05WtHM4HVyGqA6cn2aHQ0s57mIQ/sgQG8h9s/2G6Gc94Sf/OZq8IZ0Rcx+
G5Zk9bhYOnFz/hiNzdjSInrB5Ql5DhDWLTD5CFEKqa0Pq9DWdPp28sDOSuYRwpCV
tCIqgwFtJK4NBRDP74RoujE4DRJf4bdb8EWdPbMObEhXMzq6UoVfwf32Vf/dqtxH
+mDQ8vIB7LRSOqhQ3sbkPeHBOcgRJUHOZcJuDjVAyp/xzIGnzO+1c1k7OoiTgfW4
PtRWL8q8nXW3z/XLU2AToHZOa+eEGVWqXpv2sN+0IIIR35f0KF89jZspoYg2/2pi
OlRKlaMV2O6qxnV8UIl73r0ngXUIJ/VPIRYolXeuk8TT5lCtPXfFuiANd4OX0WGS
WAbvaRmpJp/g1twyKbHgQlyHK0o5Qwtdc1LPXSi4u/++g2OlPaICU55OfDw0V1Ar
T+Ojr8umafnpPCquk4Wx00zMo3aI+Ccl6lGiD/aTCtHjcKcrFetNJOPoh/dFcD/F
TIYMIWlS48tG7X6laqe9EkaWqWanx0zeUxWRLClXSIZ9TWPlsWnbDS2tYFy5zxzk
KJBB7T6aJoV17/flWzMiEZmSyHt3/kDSfVUb8lgqdGH9ji7llzUnJR17vDeBFKIl
kiOZ+K8wW3hXg+5jrPyizNEpGoXXbf8oUAnUStbmHzdsZ7/yJpDujFmHF1wv5h+b
n/d62CNsc4uapYlDzQqspP3VTwnPT6EnZjiT7ND1gQAOe1Wc/e1hQGUyywv0yQHT
KeJsMjiwjCV8pPg4Dye/QUnedfn2TvKgMssOlBlnwcEMjjguhyMofCFIug79vzOM
c9GUyrYE7yvIcnJrwhuQrYwXSUwNH32/OmRyDfxRrVcyMAJhTxkE+eh6R2vnDkD2
fgf3mCe0TNPWAO32BCdjiYm8uLqq2Oa8XFu9MxalyNqXWuNcrfTjK0EYSbigeQNC
X0V57lvxW0EVEFunOjq2u7Py0xF3XhKPwouPMoFVhZqkgFtFMQCOwwKwHSGduveC
CZtx81jWdtZxHb6Jd0vdjNnoh/8LnTYmp5kTmMve2RUCz8XJr1BNjjv30fAyIEPG
K6eLXcFhiUg3ztWgQmiV9rFeMv4R75O7nwj+/c8y5iLKsOZcuiXa/fXtDSJCCmxV
cN/M/9PT6Cz1X4/sx1neEbjHfj2oypJwSCB7Rbigxo5zZXcTF59FO3iN0/XjSnla
D9mxb9hhSOAQo5x2en0ez17rYnt1s6YMiTZYnTHpVlYSWSPAmvbeorBvd9rFfK8z
vkXdH/jQoyQaJjnOMz2mVfqD1kXaYd3tmXBIzdQ2DbWXFVANBYCy4JuxFD3xETqy
JCsGCMrjic0jBpJAwJjgAtBcqXnM72YEJ6obHtAOiYbQm32g2hOG/Pj+OzAJnhln
uAL3PX7of2HEJBLGP9U1SLKq6ewKUn17GjSh8ZOqVjqT/5Q9pDSQ1wYGKoed6lyQ
CSYm3e8x54NQBqRufKh7GUahhI0jxZy678EGdfWaolXcDLVRTZ6lpPJDdGIEiCgz
4mTQngI/8DRN6cR+Lsnwm6QK1uITxI7YFhEEKc5xanZ03DiVA8h0OIO23b1kVrHn
k7CMjhURkNp+yIbgoYCg7uJ5CltjS0uBBiundTksXHmNa5u1T4BpCereWJlXOeVE
Q/RvQtMD0F7o3bBCOuOms0z//Qr4iwBbYvQlvTqEOsXuuR+Fa+lzJtS3b6k3T/cv
/JfsgqIyNrRRgJi/dQ6o4dm1Rib8T4Kld4Z9xYaEyN+REcgHejLx+PWetjGozEv9
jbiTzfsRrFf/9uUbaGQ0clsO330T63/QyeKa9jpussXJ5/t9ZYedQCQF1GyC4+7o
0f4zX/VUHL0PkaKcn4c22nABZrTmNCI3ALAD97nPhBk/MjkyPsc4xJzExklX/6QV
vJ0WJPzcqIMt/5Eh6kszNkWvtejMavFm2WiFtYdiPG3HZx3sdtOVb5+Z6A7mo8NM
a/i9jr8hvEjUMauJTiM8I3gxAlPpRnZSdV1EONsl1Rt+E+VJj06QSrommB63Q0N3
P0pQN8DGpkGWh2GrOhoyGe1oOCDwkK9YwaIiP3gtk5eg/3QibeE9kXMV3o3tcxzR
KbevnOE8+z2HXw0wJ3IyX1zrMJK0YflJT91fB92GrNYlKm9/8hkjI3JiTrfdLY3f
iB1zgCRy3H/s5sk+OE5IxhVqATsT/Pl4Ox3ctKe2Zk4oKGa+WH2e5mH8SBTVRAUm
FxTDYPUVrdRkUauzW2qR3KEipBLpzzD1PikV/olqcbm+J98o8xSx4zgCER8+Crfd
syYcn5AUOcmwjEZOfzh8ZOO4gR1Imy3CqPkjP9Wa9nV3xSoO2riOaCbjklj+MT6v
fgAhhzHzMpwzPdy3TJahkoorzypC5IH7CThEJ+1C9QUCpjHD8P4vIBFL58wfnTRq
GVb/pqCLam1bxDcpPKe7WLlfxpLxv8H8fBirF0DiE7U3Eok4Xj5+SFqWJlNtN91Z
OzlkktYuPZqTU4V1ZBP1+uqgXe+NNYZ9nldVsxBf9i86yFDUrYM6MD21c6vVT2NN
xu0UJKO+k9DAZ6wHF52tTyaYA1uzM254544+IldM/zAL9UMbjQupWV3phsWlWpUS
j7sV/F98rjCLE6ISRR4pq0IHr3SEroFLTqciy3jFt4UmuwSLDYmERZJ596Mkno1e
/xM3jJFOIBGkKYH1mVvsjRmkxya0qiHaF9Z2jBFOefctHFiU1DmV+6aAmGIi3DtC
16NPfpaLxFJdFHOTsdLsfM91dXUZhqpaTnf+GksgK86ekTrNBWYSgw7NJ6FhWqLk
ex5SWBx+soyfuJk14VvYEvQjVPixhYixKzjHiAo9zug/UCBtXZd0O6ufIKbG4c8m
7cg/hhnyNeQFb0bvYe5uotAYe+jMAMLjjcCEySk51xY9XvFiHI42g4LQK9Av4x0Q
9wGMWihOpdoEUYtU0NtYmQ==
`protect END_PROTECTED
