`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4iUuvLAy4YD6VALLr8saCylFWUgutYzdKQEf0yhgPrB9baCpbFpePNBsAEXwiedi
4eETeZVZz19FVXrmYqqODL86bW03rd8dhIFf4kMHwGws755b1QcA1DX8S8jkbDSu
1tpY2oaPmvRKjjxT+nWdirMHjtkYB/C2ECkS9sRbr9fv3+fLxe+bfdF9bvsafGhr
wBe9fdVsr2ZNMbVamWLw3xSxOEa3ptOzaCMg2d7i3MecF7abpj3EBHqZMKNBsbmW
M5agrHM0riWQnqZuOSN5BfK3wXOoDfLsLgGkn1TyWGqGRvrRoH4p6icfBL/ybHg7
Hv8yT661sxULL7ueKWhuWnXI0iPqeg3X5zxAndAl9OERTaXzX5icMrc/fp02hFd9
rESqyDL6q/CfWSG91/Gh/owfWxcr9f/9fcJ2Hdq7oV1bCF0Dx/j2AADtHpv5REgo
qnH5u1q2SWTkHiwfSRobKw1voxJ903Pu3duPtmmAj7EM+gX4UNA977czIaKZAJtT
tSLC2rq673p4gg33fxWckP5wikFoHcC4qRue+BHNDseeUhrn2I52tWUkgRj1p5n+
zjiwPJQH3OMuBk5aZrHPXTLVXWbSzbq3i4SBKZq3g1TOZI18dkC8RUZgYQsJvbj7
`protect END_PROTECTED
