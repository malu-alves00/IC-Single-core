`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sXDAtgzoWk+m8POib2A5Rpu1c4Lm4kHqcs7+J02hxFFgcqSnJUkFBPX0thyCKuwL
8UO62l+82VbLyPL4WWVpMn2JaeyzSv+8jAxFPkea4VkaSKqGV5eDCjlT0nwN7ycL
atheyj/vlvJGfIb1axjzoCkf41BUAMODamRmgQ7aIAjLuesuKQJh5Pdlb6IoxEpG
y3nP393Yh/fzDCT39HmZ2R3qacD52YCEHFasm02C515ZrC7AtSz031CcwVg1UCk8
M7K5KBe+mZMVIWS0qN3kuqyJzkcV8tB+eLGet5+5SlCxpkGuLEInmJLdJ2I0raI/
t8hIrSxflaUxomMG2YQMMgKGmp7ii7zRuK/KLLpiHxMhZhgS3BAIGn80iOt2cBGQ
0LzemCwnSykRAicHJ7JnwFLMT09//3jJzkvoTVIANy0MDFxws2sp+LoVVTM677N5
Z7bD+8ubePsLGZP6oQbrO8rpYr72/91LLUFxQ6R73gqQpvbwKisFdK5QWN537WEd
WW6xw75wK8DR7onNcckfDm+reX2DAWrJjkvqCngcDrcb/xBmgHGGVvZXONahrtIA
YimVIpbJTDjN11pjESpILdGLucbKaY6jITsJVVHNOMUYfkQxQmUPh+fuGvI8iZ0G
7RfwUIaDMd+f3Y9FZ1emxpxrkoBWnMf1OgsnOHXIil12xWrfzmnzdzjNZZ+FhF4r
Y/iMBvz8VbOsnXO8eEj3S4ySEYsir8e7g5UgQtYkNrNG2l6gKF33NY9dMQ2ufaVQ
qRn6dyjIuqWVq/RAHBH0645Te3SYQxo8aka66PmK+hQxUUJPjn8lKcZ8pcUQ1b35
Qg4u7ieBQTdUO2aD0knUJTHyJfsr5t4ulK2fSMl6P3f6Rf6N1MLcxC7Xyo+3A9FL
k/B6b7l0PgEe4UdjD+tVE5R29J11Itxz9Uy0pnVoE3CrWRACzaLWEbA46lh7QQDi
FhVj4e6CEdhjm4z5iLTCe++WLFe4hmmrDu6vqjPZ45hAp1Y/Mfck7qGWL0QaHm57
dQxC8e2iSZkk1w+IckVtk/9zOWsPFGHJYq4yEDl5Kn65pozT0RHZoGaAQLXg4Ulp
doU3omQaxWJHJmDz4+o8CXKu1llDcrIDT7xabdv6hSo00hhNqPma2H5UWCImcboG
xInl50vuKNNp6XTMWe2xMFhoAuWyexpAbG7pc9xEQyJxBMFhUfjUOqGyAmzPlJpZ
t9kboMjx+XmoLuGr/zAQQ8eTNGpEP8NEBmq9ft6Y5fdOq55uJz75ssSv6AK1IjRo
XJNOCANGR49M95iiMVr+Q+Iq/xki5BH9YdCS1fJMvbZMVFCswyvedGhbZBAPJACq
LWnDZHVQk9wDFxsntqx+DUl3DOW0bjP16oAUDwMAxaChCwTiPfpgbtdza971KwK0
z5DPvMXdaG8TCAwcj3J61MzpxmtMz6KrXM8CfT2ZGORlgg2tPWjeXVe3E+2SD1fK
E//DCjT13su+I+richBlpZcfv89uZzFhng6/UEJI/jiLdcywJY/i9Vlgvo6L9K1J
KuBRWEriOf3pbNEXOwt9+xxazeOLU3ob3uxg9Hn4J6TYNzc8/HAm/H1eovZkfpvH
Bsz4IHj6FNgRIcXhyIpb92XIqD4C2OJJiqzhv5WNdB0W1TXGky/QyAHMsTDEOr/5
NKUg7pudoEvAQIOXIHhj2zeZMcjTD0PGXmagA6PbeTD1npxwFZGsdHdxFrjcQZNE
D1/tnt9L+tDtao6nVbNk1zNyP21apDNq48abZTu/w/BjqxdFJVKEALNGK9Kydhij
jGcGtTudoMuW2Zrp8sm+e0+P5mqfnA01QurdNHbF9ZYg5xjfn86SgTk5OEGEGoNI
TCrn6ReaziSAXs7tm6n/Udpn8iOVWcirwnqQoSMLrlYzNXSsRPXfrEncqB1FQu6F
UNpYi3xaCRz2ga+2MsKakS4yBxQdMCaIBpjwTbbSgjFNXqKCgnzX1BtjoYeUY7/v
tmY9XZCLKhRJ76ZdAlrHOEX2Ag0TgZwKGSZQmbQTtk6e2XAUfU5v8JANih4kfnPE
8JufuYef6HospfXmemt74EMyVEgDSN+3KTLqDhTKYK7wNzANUpvm715f6eVHyInJ
X3QfNLkcuQfNGiCbbfM0ZOquqROSRChSpFJqSPSRLY6pO7ECaUr5OdDeCc+qF9fm
QJRGoCPVwb/NCPN7YdnPPAGnulNcUN1KDpaneBAP56Yyt4x6p/jy/eFtAgNOI6TZ
+b3YEKGAKInjKwo1T3rPIOichd+Vxj6+/FfpmigqRh4DXWHF+M8CFFLhjZUaif9I
ST1CUWjvfvtalDIO7YKgGOqX1izy1Y1HktRwQK4J1jCnEVwOa7LykcFEg7lr0dEP
ro6CGqypDLti7bib4U3YiwwqxeqRa0B3mcK/ZnLnADvai5yIW1sW+ZM/eTB1B3jN
eTjs812mA4i73TiAmVb7htWw58h2q9Y5psU3fhlZp14C+twOpJ/Lsp7aWTwwcVkU
4QJnXgyxab5bd3t6+Y1t/a8DMofphMWTqpoNC8LwPqotlwPtWP8s1UX5RsyZUvBP
wp7z4q4PCEk2CaVuo/A2tVk4hOJJMygQSfvToFAY5syqLFmyhd6nIqFeJu6V8dzt
VIzCrXNVTl1O8CguMJ0579pbH5C46lVqqxdrh3hixJSB8AulgebLhYeGV5aO2Ps4
bJRSxMMZlFQZu9v1bcXA9SFeXe1MFEwU+8ZoH65KzA0DfJE4ZROODTYlkcH2JjEt
u5I+U+5HljIO/IWG84Xw32Oa1GDXRSxWXo9oMvCgAxObOr9LLF1EF1Gzd+M+rnTP
ZWSX1feO3/EFuUeWF7bj59h+R4kTqkE6wcOcYrNW6GdAL5unGu3HAwQcja7ZCT6C
KaDapYXYomGxv+KF3TIqFzGiBg5LnPETp5YhthY0s2fhh3m+0zCX8KYJWKJgFWqQ
ocdRclDWnxHEqhaZJLjZDxc6/wDEbz+2/OEluMGNEKWTCX4UUljDdAfOG9KXJznw
MLVGlnU19NpeGL5+N/F84WXhFnneL9dVn88ZCfGQktHp6j0pqoRd10pWQs8SVCjg
zrZKq2guuXmS43uJROi3Aa3NdHa59EnNOPMbkJETZkJec0wKLbret2qv2krmPnyR
kommicrjSNiyEUhWyEH3lGHmjbAG6cYAC8t6zBWHDUOxnVaUW2zm9jIP9Bdi+4lV
nodyKlDITjL/RpRqe03OeSfcTkCiqgqzqZDLsGjUPPzkuABbmfwsVZfplyio7DJV
a4p/u83yM3SdlBwjY7qtZuu5IA/WhVQ0GyVNjSjidFGq7YsKoyoEqpp+XF6NVYbf
iqAg84DsEn2oAq+puwbeU5y2TxE8wDEBsYc+4AMD5yNjb13m8332e9s8ISzwI/IS
V0NULaff+c+VHTK6BYIALvAYDMkYfZvHn9dyZJ1mHZdg1ntWtJGoY72nGF/VS550
wiykcCa9EazobVgZUEW/eiSX2eo3I3MJXs3+kdv040pYgq2lNz35ob/EGhHYJS6o
HqCXDmYvCcr5JFQGafLSgs1qsfaD+Y9lYap0h7O7NFTKj/x5bOvY05XLKsk97E3a
whhO9N4m8hqqLUCUjZCV3SZFY7f+znDmYJMDlxPM1ldmprXq4+29h8bzaDH2Jjd3
IT0rHo+3rDZwdOslDijJBGg5AfIV9+L6mliWkMSJu682w9SVr8lf8lG6MemHjc4+
AysVQC+8rT5rM01rntOLQa6TbUOnIeFTIuoBR2WbJgeTm9bpsqXAcmUQApwfqPu9
rVRdsKrqnpp8erhOx5TbstMFgKYSswGDjOMajeVenFX+SBttpCskzcBZUSnTbhDz
F1lwBR/1Htz/l6A93zJ8wzFDSIUmS8GF6tRNh6eJgV76zS6rR1sdyhebb6pbKAQt
fxomyHdd/KyVmOHkTpTSrgMr8ekMumFLW6lD57O9aWyozsJe8Al9Z/qMilfogg7T
3CNl/9fbckX2JdHhhBmN3BWgejnzjd7lloJHYTwFZVN0ay0dxvWj7L9+yO1hl6Wa
1OksCiByzpjnX88jBQ5+Eh8jILe1HYdk0bu6OYYqs7OM2WZ/YwyL08WCt9EVzPFo
yCcY/6qxeG3cmX9mWtvP+vBHyUX4nQbZX6sp0sP7Qx9HaSYdVwVNmiJTusm3E86S
qA5Ip518rGBkZ60Ur9mqJiffECCbKnC5XcPDnTturlAY72OpCM/2bpWGpkuPbdY+
rHMzYNRhJSREWpTmnQiBG9KxT35et8f9cJnqYxdgDSsS2ywayZhSDj3tO5lD6HcQ
nLf5FFvy0XY6pUCoEf7yxCmWzYKG13DXzhZdnWzDnVOoE2Lxvw3O6719rKsUCxNW
TnsmsWBLx4bYEpWkE23pz+lXY+2XdnSqy71pZZFa3K5PcRhLhHWFslVPbfaIl0lQ
neqFJ8mWIXJqAAs/Ci0NSwChE0fZtXpmCic9yhIVkjovzAeffnqpglKZ6WUpISTO
`protect END_PROTECTED
