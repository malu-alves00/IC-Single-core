`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vsITL2162FDfDkDiAS9n+f0JkmDxBMD6tkaQlzmAryaTEoNgE8ueohUwKP4PQ6Op
1yqQ6yoDGtA1Or3v7kf+suUZI9ycNRWTsjhba55DagSlP3wkw8vZUcIXJ922CYfe
IPKigpGHxjcJX0GLztoku9UEUWH7OBvN1qNaOuFIhTnAI2m/vBPYt7KHPpaTl28z
ldfrKUSwMNmEecNxoXDH8sL2U9umx02aqdHsu/HLbTTYQASchc2RJVF313FDnuwS
sNYqmkuvMzRtLdBP8A/MtfKkvGXiLjDxvDoDsw7XFywEJMb+kB2SE+XdnIfgspPF
2L7IfFwygtWU8FWGTdBv53kbNncfBAu7HMlbWU9YYGu3ymVYxd1LK4CYrwDqjKDO
AtocSEj5CpZUKaH+aPSnQT/SXiYG9Uj1R8Owph2phaqSt4gxIOsAQf8LkOwWEvr8
jMt+IhPKMp6hvtVGimTpc++82VOeLUR+ThrIESKq4FpbACEmVsjI7FOpZ2XB+nVu
koffH+33CH7YUY4WDEHrqEtM0Doa//OT4d0E5alei07Q36F6A7IORs/M+LZLil+C
DFl03pIa+ORCTmbwSVL0enBVJOcne1htZ/2yeWexOalPveYbIg2SxK0NSFOvviJ/
QSJ4rUeh2rIAuG3cTZGivpWCnrdD1RAhG4exGxGsA3SlN3xSWZ1Vm606/x4qC+Jt
M0Qj4C7ACKaKeNkn2bkoAcgtVouGlIMh5IoLW/Yir4bQU0DsV9AoiPWqfiXJUCxb
+nNahBq3DuKqy2ANWOW/lq3+P4TWz65o8FEGRTc1axuV8wKaRzWgpXzrNJ0QwQMY
qmop22ipbWHkCYdiagCex+PK+GDPeGmhGpKTLGPgux2vFcKF96joSMrhIUEHPf1D
xn2de7joHMUS6GqsD2bvBlrL4ia42NUE14hznF0Ngvmc+xI2f2kZ8lIO3GPHB0lk
vtLSWf2ki6F1fz7UDSt0YCzEktURGFhNYt5cL1QpciYiFOg2COaOi2ylAz2F63IG
+Iy4ANd1BnrecJUCWrdg/7MgX+IqKxEO7h5LU8L3CyS0g6PJqNFpiTn3ugioSNS8
avW2RuBc+ckoGayss59iSJqAhHgga3SVLxt4pqLbNk7zFQLF9H5CMZSiQa9P6FXD
G+yQkP9HbHVm80oFxMQG0raW1bGP9kGxbb+yjHl9gtHi7uDUgRWs0h3aqiWX2cbD
7D/AYd32d8ARVpifuWqAXVOC35GYSW+Mq+rOtSsI1691NDeyszpGWT95zSrA6HEO
K1pADSyGZImpV5V6nYxMZaSWTNvgVtPvXQ06Gt1n4W5etL1PBjseHHtoQ9VI+nsQ
Cg3okmxUBxgHoxxRF8q7RHSfPrphSmTMhvxUQLvpFz+F6yHx2lJfgSmhYcaEin0+
Y5CIOrZNrFLGy7TBqKGhRc25n6Vcjy8cRDiH8FaIy9+dIR+ynEdgQjKlmqioVM5p
6Z4qttjQRkSanfwsOYIDRyCckwftpZ+irARl5UdHEDLI6Lww7aRBhbzjs18tLqCw
eVVY6BNdHfHAl9U5klnbA67mTMkXZQzh+c88Mb2+jqzDuKG7DzYS2MxSsu2a6BHj
hVv785YmigtEvAiW0w5eegMOLSr4U90vBPYc09kSdxx7IkCUzIL4NRiVasd0Dw5P
Oe0whFeIGR2fiVpIKtzW30cPMVIs/zc2x3EHS5mkagIKKrG+qEEeyYEiHTXqZqXm
ZeI953bRBWLYy1016PVfq14ORsUT5DpS/QPaTdmfG4fKXElcZoP8gB7HphDZbOYn
FkDLAdt2cqR1nFMsXr7w3+bnCnST2m8xRKWFRXA0NkhzMEv0vr1NdP8KuonxsNNw
K9QDL9txxmujtfLgendCUQ==
`protect END_PROTECTED
