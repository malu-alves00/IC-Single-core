`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FzbYmtYhTBvmdlthF7lOITPiqjppFFZOBhvNytCn107X4XDz3XZtcKeWe63hImPa
I/MYu85tgXqVD3byihY+Vm8HUqHOy1yhNsLCQv5+wUm99T27bnzSAtizrizex2rO
uriIam5XCAntCaxNO6GtKuqc5XZmEOXntamztaTQybEcGHI0qTH6oW5opI3j+dBK
VKE6MQED5YFxzQiQPQRXLym2WqygSBLNXvjxq3K6X9DSicA79cW3ptAEjrWe/yTt
qHK3NIucNSFoxtxStHA26dcfPTA4pEZwe5/huOvWR76tFp6PyMDkQ00l8SLPeoyV
JwiEUtg4IfZSYNFGyNX6FMsR0OIxbYGSBnhmYCqvfMlaJonWk2cANie0ItssIBZ0
4UuTkKMT/4/D9jEjmvGzMQViWKhMxffjyxN8fiOGrqubY2minjk5C9SetdN6XArE
YI2hU0M/MEpIP/9cfGS1SFfkAjTVArTkRnth4eFL91AO3iAcVSprq7ieXnuPcXgC
QiGZ0YXxWOzQtgp8jgbC2FZoWk7DvVPioZ4obEz0amdXz0M0DTA/z3j9rtBAqLxQ
wFDib+ryhZpk4/B1T50XmHjN8WAQpfT4wi1ki+q3v0ox1JZ92/GGTDbuEQxLUmi+
3AlSpBe9T2pDSERXZPHB5aDgeVqNKaKC8godo0QJ77Gb5HlnkHrPfQtwo5Hav0I/
LW61nWryykJ5zPjcQ3UMc0/CbaqiT+YZFkVQbJU6zs8IZiTznQzWmbs+MfaZ9Eqr
QNCznGDnc29mVzIXbyltiKEyqpyeC8eKh8BS62dQdMyEgkvsb7tfcBq11Kfpam+m
OhRwtQtVvsOVW1/FVMYYN2DpE4qLPjhla7fue52C5Mj2Rf7Z9RUkJiOZhzIFqz6W
lNEmEfbo9Jl4sw0xkSfWH8UW8Vf2mBJZAC0TKqbKgMsN2LiadPczCNAbrtlfxjr8
KiLcVE2hf+2T32A1I6txJh67r9bQMVe2B11K/9VM8GoumijaOMygRW8uTLB8LC3t
8R1x0Q5fuLcwO/hp/xWygFM/Y/2K8N57qptdc7Pi+zo9P6vW69yEqoPfuRpvotbk
7TlcyIVMtZeyALvo8RpvuWIWEjuq2wwetCFSG7tLEtGp0yzWm0jYbuTpG4A2dW0/
iLulaFGgIkMiNQHpyc0RIGgL3meM4eB0L8RiqbhNh707E6W/ys6f3HzJZOxtINvK
rJ+64Vb8SpipbCwQI07dWd8Fpg/aa8xC+XpGSVBwj+OT18oejibxBq5O24NLSDP6
faaISiI7OxS1Zwk6oPnfE4opgwq3G5Q12D8AhcY/Th2UxosjnJUTH4guyLmICjHd
t1Is8WpQazXUkcOFHgWVICdqjoUWjK1Q5A+Nmrr1WYL1zLnximWx0+HtX88wo7F4
m3Pukqo+3lC3mow4p0Sqmhp47MP1RybQptvIGlWt/hCSP2XXygFmNjeQqnCkTzCW
qzg+ytzziI/5GU3cl6OW3yb8TLPT9R+KBfSP/G0v2eQH+lNMdyRT+6wgp6CS17d1
O/o3jwUGzfc1nGCgabRMaKxuaV+Nb92aKjBIhV71FX4sSxoVePtF/4IF86gVhjE+
NqDW1dAfXsfELVfcG4P0J07alV4R+XeQx4Lvv03BFxJDzxN8v32/r6tzJ2ClPB6p
tzWh+AyzE+uk3+Y7nEHgthYKjel8pewMtkF+hNAMQH7P3VUB70FRCUby5VXUARqo
211bzQRyDuEuGFcHf1F1iZI4ZnkxJ4qCVzGRYrNgYvf06ewvw1ZoMmY8AGGGdPPb
HOumgZeMQPvD/XYb2p804QZeu8dMMCiqj8lTXSXzrFuLl3DJk8QbmpI6y1rK86P9
R21fLhAFoHcPMevrE0IM8p5irkz01DpZnm0B9NQM1RKuczBHQ4tr2+EFpZ+1+8uy
h8t9XuK60M/7WtUcr8Pei62SjBpTk5OTS09I7Zj2ayZtI6ULm1k6h91nmKCMolVK
Ne5Wc/pM2V4L+mPk11/Bkc0hdHK+in0NUavU/Y9sUsMCEuK/66N0ocqGbtNc2rNn
QWpMP46C5ECedWx44dYiIAok6g8+BDB4FX1QgyBRt/LlyuFH0//rYW2xUopc+ZkL
7FM3LlCoHQn1Bo+4kvBcnYexWft87Z9fjoK2WxJvtdnwb6sKczg4/QwTYxcnRIpo
lfZhoWyNdSwK8Uoe62mIA7J+pve3PExfPzFusbEN3Wnj0fDUn+pJJuYYxuK/dvHq
R+lRS1aCQnVtrznpt6mDIjNw3m+4tMThyCfzbSvh2QlZgefbdzI+GSFoaBfT4ew5
dd8zMsWr5fBDLby2meH7r2ImIgVuuZiriN9NajDj0g6wX1T77+xpsz0Crd/hRkS9
zEPOJWi1K7K6T04+7VF5psoh+AzWDRe96M6Skj+fyT3tm3SSk9ouoWAfJvWh40Mt
+dWmAhooKkgEUGwlb14I6jAbojwvTmai7htZ2CpZOD7mZ2zVZ1O5N5VxQBa0HrFs
aYRMbWyRVYKrH7WLKZej2TofLdqrAHkrKZT9xrUlvDbuwsDG3HVUIaPwPG4kW/Wr
t7s13tRNjZ9ZfDg3SMwlBBZye0na9mMANB5dPP1mS0iDoUo5oLOnGf14OzFUJJVa
Dp2bTTLosYYy2clgl6RrBm/e8ci4RF4Xi2d4g9wjIsrfEZSgXBIz9i65A6vNrJti
u8/PzUkA/iiSh3VR7ERge46MrpRsBswb9RooBpvzJp6zZNCGfvIPYdITCVfFeAZL
L76Fk2EWZj54nhwv+pEXH5WkxH+kWQTD1X1heyFitTgtLusipJ97cIHpAcmz8BXu
CTSiQUFp4AfUBTKCMfYs2bKCf40Q5wg1jiOPUT2nhfKy+xnPcud4UwJlNUlGsLmA
nMsXbsHRw6BiQ0rAbpjsRdQBuMkAVg9VlNcmpdwlXIOwnP5PWNoEKJ3sxONZi6lh
6OdbqVQ1My3W3JJxwtNNIqfBkhwO3bM6sviY1sLqCfewv1pLpQsnMQVNwqM3mlRx
e1kqR07VPuoRr9y4G0gcgo1LTYAbyFn/z3Zz1Dh60BVL5nymYIXDLfBuZrdL7mUO
9TDcX5dy44Cdd0agPftInilG40e9+hNlxZoS7YEa3Vv/S2NjGNdWoldxbr2uIorl
bchENmS7xwoO7T4+IM9c+DJ7JmxDSaKfdX8v+bAGTjt/PIV7EM+jJ1Yq6Tdh9K++
MvJw9Sngt94u4ESBYxFwPFjU4EjASPr/pQhCKXrCi9mRAWbRyLGZ/9nq6wA8MNUD
c7i8n94mkwjzp6d2aWYp0Daz8TznJZbq6cBA308NrSnWhFwVjq45HWT/22Ns2Va1
kSmUdrwNfKIljlTIvRkkHvm9A3lcdkun+YHi6PwgtjdFQnTCxPTcNwAjaWHF/g+K
pRkpfbVRYNodJzAI4kcKUOtoNXG8kBo5GheAtAdHCPPLtInzNawavG87DGFOSwh6
DsyDUWPOxuAJ56/jdu4pjYiL3H4beijsYl0vUwpyiFz8cntwn2tmGW29IwCgCaia
jZZLJihays4nGBImR2WuvH00Cl23Ytu5mOM9wD+M5biX1/zS+Li36zIZ6OfBG+W9
ZRS7SVMxElsWzxF6g2+xbakbn1uhudlc0O653QNtH2wZNju3jf4iaA4npEXnnypi
k8pDYzoZeiG6h/sLVYb4vBmzUssVtTkLn3Ban0Tj2BQF8cNWmCXHpdMRkoWQ1KX6
4IckCzTzfGjOC8v1eEizc8/6OVwJV7qXOdbt13ecGrXiJRRE8uNi5mP335Xv0ynr
8DHWlBEkwz6xl1e9iW43kzePEWUfWeO2d6mw6XoRTxIE8OdWrTob5Lv853NmP+k3
bLBaSiyEbCledsbkzQkVmT5GNXZlxrg1AfE3nw0bP7DLdMCKFMhqtKVqxr2IsXsW
Mo3cL80RmJlX4j/gZcjwT1Ooli9k5o7OGlKN72YD1cn+nfZGgmJ9KKGK4y79Zl/W
we+jyMWNFThNYFfbSUYsHJ+su38ELZE779b+JrdAgUJM8nx/jeFtq0fUldOMp/+d
2vmc5TqjO3KWtQBtJF8Vp8y0ywrDnlWK64K5h/qWUtF3CMj803+HQK4TjhhBObgx
zn9AHFdyRjqnPt7IzII77GYNN11vYHrrVYJoo9zZOozDQpJLbQwSAk7x2toYljs3
YhJ0GcEEqwZsPsQct5RQQE39VGAUVN83xII4KvegAa8IvBFm1cW58N15OVWuiZnO
7biNxMBH/+uvOVuojC6zlmbLVK6Bjqbb/ydEahInmMnCp3BHfY4QDXKsvdZtFORa
NA7ftKZSswuZxlDo/ZnlEkEXHuiZDyXl2TYIv+L7Wt3QeKXBu41JagTgQLIUayE6
OHTRlxbi98ZH5Fh7jWwbXCVcu4JhjKVlALa4iMsTld4or3CG7j0VBz8pRUSV4VCv
gvLF24uKL5wrRcHE+1S9qAku4aCuRsGjonqiTKXkZxWrmh9CjQ86WW0VxylSK6Ae
DpHRv55lVsKcrA3UlfrOG4hRgW6UOjqV7kPhxA6d/WXy2xwsxlwL7Nby9V4vkvyb
7wSYqNhRC/kVLacq3Us6YESHgrE/L6C4SNy0JAxBexkKoqZ3YPAnYtViUZkRfWDg
ArELPO8pfTle+aYigUY7F3830fFA5oOJCEc3rvHhix55kURnBVtwNqAam1yVlYYk
1ZMriOjCjSugO/3ZS/w4MLqWzYDuMfHfs1bhAghNq6LJ0I4Sy/s4Fivh8IoAd6r8
sXLQxg2tP2XOYl9MoRUQWpU4TS16kJLjKRqOKBHdeDHSBtcUVdZ+T6UcYTCoczU4
8BlMQkFk90sgei/YGlUoGt/d7sOTp9Zi4pkOPpXr6ByesGPgDyseOWv+sqtM58sL
Sb65HkieGTDCzd6vHest43PETZR1oc6wPEqTLVSjZlQoYa1CBuOZHE2S/BlTbzOL
5efYDHO8N3tP96QejHZA435/llX/XwvDPeB6WK9GC74y3JKM4XWQnQX4KA0gYRWW
KPDkOd1aoVqD4timSiI5LwpfTwqvX+bD6cTfph4UxYsX7FidnBYi/o0B2gSCpMJE
xMuPlDHouD5p+Hvmx7KU291LQSb55mpzJqDyo0UKkzigs/JswuXAZYEMFY33hgdG
ORsO6MOaYGswiOQPJijW3cgBeOHuN/PgxorCtlxuW6kAhU/xYSLREGrabngbVMIv
es1bbM05X50HftGgAzKq5YQmOvrjzXgij/4H9oh1EGnF8DFWxSwtiMFYYfnsKwpQ
pPcbTfLLnCro3wPlFkUEl6Rm1te2Vvbvvhf5YOUFgW0yMRFNq6YMlmaWU4vjnfB8
y912BUb0NCoEz+cRJiNlUjOVZjFUq/cBJIDvvDfkZc9IoprwJ8RmiUNkDSAomSFb
HuVYORBV7Q9ymup6Csn9Xh2sgyXCQxmOOl4lS/kGbrmTHYaIKZL95wdd5U20qeJS
4UGrAJZl2s6rCMXjjrg6nNP42coowZG4Hh3OtskHyF+tJ1nGh7Tg5MR3ZOGJdYeS
UnUTjHmPMjYqu8CVakj0zMSuTc3HdeHswY1Z2CMAvddtQ/mNqLQGoLhcIdrneelc
m4ATQTW5x/JOFPad2Hi2z01+etAz0WmRQqDk1jMM7Pza21ZnMogVDQboH/k3YORl
ywwSeXVDfDjITFB3D4OYUhxUT+rSaRV+HZgYqT84hsv+2td1e55ccy1mSoBKovc7
rse8VKfEJiwTtHOnv4X3/euEOhOgV5JLcRwmWTEPxIKhGzscq5vdSLYvTQutPjLO
wzCJXUd9mlVc+B+y+U2TtOSuWzDhUo+7BkNXKN0nA3oOdZmxdspeAlLbm6td7nNR
eOBroJWsBQIXAg2imyzt7mjICnOSotY5nhf5bDYwQke506MsvCM94egqHEH7qwni
j/HpXMY6U1nfvyyeMthDt5ffwDwud6OM4d21viVhWl831QlDfXU+oU5GzzCwU+v5
mTKBD1Qph+d9tGuAhN9owXO0/GAdtSX+dUj2bnIYvQcr9JBUiIOJfWRhzhucAdKU
lEOWT8rbl3ms36MYs1rkWENYCe26wm81zp8fcW7IsU/9v/4SeMLvY6r665hlKhIl
TEf51xccAl1As3kFTPlUFwaCXC5PNQG899pcuh6a7rvH4o2+HwFjEnv0azrQvNa1
Q+Tity0YzV6KIp6KbiPlTSspNjVmx9a5ME+KXS6SiP+sUFMFM0fft5SyakuFo3lc
u/NNpTTJ49XgZbDkGToPVSsYHO98P2OyjscWzxhPydev9d1p7XixL48s5IB4Fmrs
WxTQMLt92mQkU8YMOtBSEBvJRyq+tkCy3FEo287ATf/Llm4TQ3YJSBzqzeaaV5oN
TEcosdRFJWs26XT49MNsu9ZP0oE/3Z29nddIvctD5PzXQCbsngnqIVWqL5WqrGCK
FnFQakXHwePVlQfDTumAOwTrAFlZFRvBZ44WiP0ElOuspr86FcMMZTgll1HVg5O3
dgCaNInF5DiNglpdFvIUHKYhVqABI1cYI2uCmRa608fIBQ0KA0KAudqAeuGA66bT
dsAdi6pGSsEMGpLElw969w/dR07FlXdu4W2/ICwhzvp35u1lozA9Z7aQsQ59HViw
ghlebGhVk61avnY5BaWGiNiUk5ScBQ+PEJDNW0TC3YV3+wRZR8vcwpvW1oldlSTz
oRCisw8Hox76Sc55c6K0y64U6idO7hLzLfglsfvAKr/S0qX0+KgCuSheTdYTbmkV
y+78EJk74lQGLg70rfPxCxZLlH7oeyU4c6fCEtooCympWH9lY71UGOCu8nR+SFXw
xif+XyGOw/Hff21PB7JTF4yZUS/jKEevBdbDOa5d2geSZ0cetdItAVEyxeKM6Inw
EOFVNaHr+OIzFaTtOMf2p2uTxGioahUQvuN6E6yx6dgVyAxG8Ljp5SK4xbDU/qj3
ZkYJkaRGWOYQE469D9jGNwxvrpUeKCbziPZepAv6d/I2lFIssxD/DmoZdESdWtVw
IpaSJaneYfGbC6cWQA00adIyhnjX56kFISpaaBm/hoRozPIp+hDrLFjl647hxbZ7
Bi/1WcZfEEhbYREl1VrXp8KaBS5UNQVtpee8OjOmoC7WEgacnptgLGu8ONBcJWp6
TYizby/HQ1479mUdqo3ljyLzaJwhhKMvbMM6uKX00EpPSGMdRtd0MzPS/244ApIs
mzMPSucleyT1L/2IznJdxd/UnBgfLTZZUOK/NIx6R8emh6TslCKmT16p+i7IP7dl
ZEn4cdlQptmCuQb21MGlBtAF9pxM5g66sxWrc2tV4yqlpskbx7hm3v4Mppl6Fqpm
9X6aUH0XPet9TanUw16CwwJrHdPxGVcV8ge0tR9tl9Jw0SAdakEoZX4wYwh3H3bB
M25vyQaGPueryNxTsbLk4iwnQEzsdmmDxcmWRSfiWUnRb7v9BoUpDVNBbafnoTMW
uLaD2a7BmUiiMXZMmd3f5ZpbqEgu1gYw/nJKvNRo/uTQD+q/Wd3/EkM/nk4Wksoz
03LFEkSP4dkFe9JNpkpcmTsjmngoK35ql43+Hrz3MpNI78lIbD9ejCgMe+M1QZT+
kwXgwGjtGNIVEWEc2g19uZkQr8aaWBuCZfpGwbXIih/3bOMUN48P05aefTDpkOtb
LGyjjsBkggTKmxOLR4IZJ2xWQ0ybRYtExx1jn+UaHLvBQe4Wie4mUQJm9biIno9b
dm8/4tuPZPRIiLqS45R+9vvULd2hoTfnXtmvTsMX2e2nNiizwyU5c9LBjMxghnso
jUa2w2R3fJW0DG9gKAPe6jqYCfnRBOW0KDIpfAdKAVXqeR1QBfSNvwgI/PqzU1tP
e5s3AMcaFHmCV9Y+fpgp+L0nb4TckRNDdXvze2C+qkjm7o2gt9X6qpZimKKHj+LK
8zLRBkcLbLYHTEe63nrIqZDAbvxodEtoJ8NHnNt8ifd4OhwsjUFx8H1SdbAScpJj
RpCXicmZXa2nU1vWSE9MQE7zhnKTc2VKu7UZ+Znt12mMrWoBJijhnnxe5cBAd1uj
cF/1z/w95rZoZb5lfQZtWr6HhFWdhEmxa4SI6faF0ACHVeTSac72+/6ULaaYxDSQ
t3z+uTbnf8epd0nizZsXB+LN7Zl4WDg8DF7L13EU3bO9MKzSF0nD+hspUxWbgUdt
dkpSWb+V90izQIwQ73P5Sd4iF5fwN94mb30kJKFwHpLHRqdkIcHkXCn0CYoIiZ8G
Iz71FqoI58KJgM0vmAR+yVlzCe23gb1XGkIde/hR7gRmcEPaQQCwZl2UhG1jPgG/
6Tf1q9P0VjVcD+p2LtlWjscIp4n97Jqbn84Rv2JtHXEcQZ9vGqrHmLy+rTbc5Fv+
uikSOAiokpjVAU5vWXTZQdT59tj8ABBtRPFCh/lWZkAdkFXW7877aCJGX9UO0ROn
G6ppN2WqBKZMD1FBHBWihZfm3dWdqCdt87ZJSbwsGRijBUz5Ld/Z0ZEjkGpUsJJU
bBEHTeezjwOuK7OuV4j1opD5NQNoXrJHEq0pNOu5c1C1RsUydsHeo2PzzKLoymFO
VPH85hVn1J2XFYEiuLoQdyigZsPXIHxHZ+GgYMOwfV6WfTSQVR9bN2cXXvflJdoW
u1nitUtC91nIytGegRdcb3ycSlnaN+rY75MsVhuKw6Lo5HXsRS3pbIW7RhVtXz6U
OLCTf6AIpIA/LHax+vdu3zT2IP03W88rMMCfRxX+ZqyH7BdtNPGlbjLcrDXmsq1s
jP3c3jC7m+KjRNU6/+12ft0zqAw8ugK1EoeIfFbwRmFmxZ48uGHhFgVmvpfgFAD7
thAgEK/v00v10vjOC2aWNHTLeN9iGjoAz5tAp5uBcKEEH9cOcrRi9b1JAT1EMtki
yki/aIRnR9C2BhQa78k0YVEfxD9s5Nom+EsJjT5TiwKmtk/0EAYN3XRPLdZBCrHz
hxVcGJUjoRlj3MPD3QEFTa0DGI+Uj8Yv1TXjz+OFPTiNrFOnt4c6sBgct46EdS0f
fRyMdJO0rQ0xLlx61oR9IG4h5iQIgfPIsRm5O9U1DbA+SvoAuDkbFgJsq+KOoXBa
Jqnr+khWbv2rM0RdXp1G11DxIZKHOhLHbEvAi5vSDgxoxbuPQz9/xJamCJtm8Dl7
9F3BKuBAP8eXwwV1+3OPEn6TN/VRt6ui67GHujteYKSazJmB6ewT9jlvKrHqgpQJ
LE6soe1WzCJ5rL9vn8TCY51eAr7pJRbAZm87R249+D0moK6mLTWF8H0wvXPPLaTg
Rt5oMX2uTjq1tCkgLSXMq/0vTsAntDJbE5iB8j4+SxekZzkBqIksp1VcO9CKdGbg
rFsngHwkazbFICBDEo+FhCTINjGfHpGVIDtVnMNOYD2rXmaPrIdB3y8VBNUOmV7W
/xl21jhqHyAJSnKgfyy3pFpC+tu+KNfvMrVjGXmXno6E4PZ11qisMU99tmfyS16a
KFwP3bS+ORCfzB33WxtRw/UQvXStwaB5GMh/GyCupuv5FN61xtM5dY7yFOKCsgr4
F/+hJALZfiUeDOFhZ4Fd4YZtaCBqLPRWs2IZ/IPxFC1ViqRCSbG1di6wQ1fxdi1/
iFal4VN0fjV+Pq5TYCykDQySvfSUTpyyE22ud9Jbzyd68iAYjjzgYBmK3aPWf6dY
XYrBb3xfsOXOJQV8eE3pEmwiAH8Hb4HpA4MLtWgGueXjxMK3rWe6HeRrEofhKAFj
u9IdSAm2JCbCpXVnFWzqoqyJguBBpEPgR0S3Z1UFcvMwfWK4IEHr+9RDE05uwCUq
QLKyrmPD5ruFb+ikdcT/48JfcZXRsjWfuWEClu5nmmj1VZbsnCNZzNy+jrm5ieDh
7uKv0r71i0XQzCRIDNWctv6xkf4yAdoz1lK9VU9QGSh5DzSmqbkOXj4vH8/6lhIO
H+yAlO6xGHcqQ7v8VAVSecoyGgkkQQyr7DJkdFSZis6bop82dUWoEEavSXaj/Eh+
VDrfHUhA9b2UuPOP4q2P8LjLqDbEB6uNthY3rbPiVLODUkHyqs18g9kwUIWF5vk0
WarSa00eO4lARBrC+NEagWbeTvVS3qy3YdWrGCLtHBNYV0/nnS+DUC7BCmB0aWdz
mFvJy+b5Z/ovDf+NvC6rZ0Ycvb5gJWV+XpYxM340l4WRxJY7wyrxsvszVrCt0mZb
LI+SkpLWixw7OIOC8WfQ+w2NEfA1wr/ucGnYIj313YDhbDtQrxfY5SwIKB3IAS/H
agfmbzReRdEgWKGd9HH2kBG/2dhhOkk4SCiOOlGAtEg5gsw4HrcxUVCjHeDabhsy
L70MwCWVkcsS0iaW3nV8+jxXSDZGsO9mYxgghMptugvcvEQmKBO+mMt1ejlTp2qM
DUfhxqSrb3pH3ZT+GulMg/1gRd67/zlGCYHUD4i5Zw1gL3r8htlo6oZf8vL+L2Vt
stw1HMA57CaNSiBXEhE9FsoVnnDlyqebv82ylALVIqvV06wVvAOcaxdtV7NYyF3d
KHl8AT5PcIDuFcuLpc/fCSIKqBJiMvv3KjVI780zfKhBtxkB0CylRPMthLwSvUOF
SlS5/JyhEAVDJJ32mFRS/YGAlT8VIljZdDGM/fSJyXTM76Y/MkmUBCUsEgg08lRZ
ZsQfCyGlqgYh/6eJhlzPktUMdpQvZlJcETuC0HBxfwMW4nHVc+amTbK2ELnNeMoP
eB7heuL8oalZ7imuLuhsFAf+6mNdfNwU8v0VvLeGxoGXsncFvkHTb1tXFbcTHD5z
cejLlnI+PzU7d81CUVpes8n5WZi1rFo53aglgQDhsHxMqsTNgpDihD02t9F5hFYZ
sFRu8DlzADsZRRhAS/wLtYreyZYY1WKeMZGdY5dUW/V3B0W/gmVV2R/1/O7SK1A1
w4x6+Bqo5e///6xcxyjPYyeA9/l1Pldkig6T0IzqE4o8ltxrUEAW80t9GANHwMXf
urCEfHIQDR91TEzV7dQwovWwsj29ADS86ceyp5osbjKDtZP2fNq1PFhHam30k0XE
loOK6LQbdkOrmhxH2rJksOs41/4X4YtfKx/dJw6E30fUWQMIwBN4BMVL5iwNjbXQ
TOhWK9IJb+ScdyhSUbSuKbqIAq8I5NzugB+APKOozoH/SSvEgZQFhDHzT+//CBup
7ISyy/9xvO7EzI3UiFqqSsl55NBFbeYdxeJTwGxv2BjMQAWTOfrH54JEFo/koV0O
S/wNmjeu8Ijt4WX/L0rEnTTCozG/GmLdq/0My4NwAseEF77DRDX4TyqJxBF9e3yc
Ufg2CVVUwx7suk3V8dfyE5CONU2UioQgg8FylDBhjKmgJF+V4cdafGCrmsv1CcCa
pg6unbhuIhTD9BMVEiAJWiA+o+agvg1GW8Kvqq1eJsFiWaZny6F+D0TnC5tuyEJR
VG103d++Nse3mDe7jGvhDLtnRCLJXv+RR/hYwk0gEo0ujjq9uY/B2oSLwZYaCSn5
MdnRD3ScGYZns9p97auJ6vlab9B8SfkpjnPZQB02zZn96Ys3l81x8ClV7vc3DCyE
JQiAWtGK6A2MofpCr+cfXv+HIDiw23/iVLPuct80zb5up4PHaCmEfIm3MyHOMBij
bJ2Tss9Cl3mFSd1CYQ8cQ2bL1bfjgrhGkgdDN9JYH4bBkkjoEKBAhXyA8oIFvvfC
49HfQgsyVe3Rpvj1ac2fQuHr23dV33Dyq0IwNqN1EkqWSn5THaF08ufEhEyKRayx
hvbwa5zLz194NEFoREvRHqcFDoRv5QKIot0lqvk0mC59hFfTngaMjMS3c11NmqT/
E0fyd/rimHfQaj6wEvRE572mASSjQAA4GVSCZR3smL/ONyP955KZKp2iQW1G2+6+
69Y2LGvnKUJiD/NOtkd6pbGzyHUoy8Ra79SZDAN/WGowDwIhTTHh0hhnGerUJAi1
IVR0Bg8as0cLKIRQYtpEtLlQMImRAMo+f7pxOWSdj5nQc+TE+JuMHbJjvOOqDcd9
PwYD3SkmNYUTbxMRWOIe6DBzXo9+ufHaPhqvre3M6z0/J/r1PRbpPjGMPjqLJxTn
XlQSjQEiyVxrfqd2LR/vtL8JY4W85GaNBkViKcjAtdPkqxrS8ZnB9ufG6eTQmKY+
52CElfLlFWuxgmltXU03MIbrOQu6TwR5b9q7OjFNPKDgQgDJBSSpdEv+1wn19xUO
HV8/E6PmmD07FRVje7y83/DvwR/iXd0SX6DjBoefXb3A4CFbqM1jB9/mtPTww7fR
vLJ2rb+3UA7AGJrui5aW0NjBV7Su163tLAwjxEtWEqL5vcEo6mu+pULRgTEoFjVl
MRJi1Ww3rqofYCd/9d02wvLzr3sj6wm1zkeJGtMLm4PSKPukJqR8Imdw5IymYhdu
8B/XNejJ+Ix3d+fVsxYVBKplP6wfppHl9+lDob8oeJk4HMQZhfb9vGRj4HYzJ2ys
dpasTI4Rmdm03U/k4DlhJXDgaTt7GHurxEdYxohdV/KxFDyZ9XCe3rIhtfh2fZ3v
RUUXNzXjK9lJQDmVa3hAcLYZaSVeFypjEBPzZ+b7uLbbgne4rO9J+CsTU0IwaeI5
+KdyRvZkOu2RufJ0gtNNl/1761IMHbqtA9xhNXSDdteYCrHSBhG2kRN+q0nxA0Pi
WyIIUyo+aCs8SzXCcXWflpeHTWmNK05csKHHd1b59yzyYlVTr45hsXqODFyE64yy
X2Tl/nt2qge3m84tHs8jZpAArSW+9ySlVhTLzFGQNhVf2XkrdW7BiPosDlbKkAp7
xsQo1PPumnJruJ54mDO2NyBRjXacG5nIDKRNy9djpIOv3deWBW2t+Ih1j48m7kx4
TazON1kKI3RP62WYBHnSZxWi3ZP+1BG31F3zyvVeYuJet+VmJC+NtODv9ipf+MR/
2+K4YjtgjXxPtCUYX4WcxxLogEMJeYBSpo6idcveJAaN8ksdhXcUu7NJbNGdB7qO
fzf92gXREivqXAikBwaNXU1vRiPS7d0Yw/6tdP26Wmc9LwyyZUBzX/3N3BD6jZHl
BP4hloqsJpqpw9a/Ff8zl5VCgHHItHHx864erA7Y1SrzCW4My+DQdLuH2QkNIjvq
fWmdoOxpIqAcEDT+5xl7yWS5UdPGdSKN1pW+fwtMwOxwgEC/8jL4+K6jqVJ1a4hs
zuowCNDzmzv/JCmHxBa1GvY+D1uLvBCKNXyvt1jQ5NScg14IKEK6x3LxpIbGu9mJ
C3Nlf7YiQDTB/MXZ0ycRjazpwEVdxb/Zar8rBDRZPmOtljCsz6TWW+lMqSQ5+FDU
GPN47tQaFlVzVaLye2ZpT3wZbx7RLpyzB9+rHHyNtZIQxmAYdw0+7M7UXq2iVgI4
6vRUhho7obo6FSH9JkWoILmLnJNkxcYvxkM66DUZ0TpTffyIdj5nzgVZS4Ilg5kA
5c/dFPhJGt26/fek0V5FWsGufFRfhrCPbSKNpzsJqvMfFHJj9096uuL5N4uNz0iR
PkBheffsXq5MuaVY15ZjkLbEin4n8XsdRSZFFdDBYb6dZow0yr1qYtpaxyDzXF50
FUBdMcCSs0bseIRRcGMxxzjClVTBcQpcV3wy3jXFZmIeEFDHzPcsQEQO1BKwt5lu
1eYq/5JpFcwlmm//Bnz4bLM8eSHM+EWm3pEaZD8Kyg3Zwwxdy/WGVQikp90858iK
aRu689xcaeE++yGhsJvCTaaHG8/f42GbYELivaSu2q2axyrmAfjRH9aq23m2rxqd
HMubev56RszXG+RoFy8bOWP8F4Kb6Z/lXNCJmDe/3rruJGBM/qxaRWv70TaHkpel
WA4y4Z3N8kojbI2bxMyq4urXUSj8fwEzm14Iw+viGFN7xpJZ3NVF908bn+E1Qnmh
Ph8x/R4K8yC4Ra0oSDwNEPhgqzeL8QYTSsT9c9gKhPS9bSSwHB1P0nLkoSGyMT3t
UaGJBJ+fp1Dd66cdEv2FirTQzqtjFAJGBMMYyhnyOW+e+MGfzbDolTR+YIr+kHbh
8wz3nKx7LSElQHgCrd/yaYWUav1XixpAW/aDQ+VOMgKIDLSRvXMx/ajAHlsjmRcf
4RFxjtdEvy1Zln9nXkIJT00Sg8oDRe4IxLWouPKapjrMTW8vpF+OMt0u86o82usU
kkiXgDeWIkDWP/h2DrYRn0sBYLZMPrpJUXUfpspPWP3WU7lM9FTGnNbFO6lL/t2d
9+TRpV8DnkqL4UaP+SW8hreO58Tkv4zohr8hNttKRxKy5ep9ME/cVqRgJroLk/KE
xb6idCvdEFwxgAaDWDx9ZjyuMD/1+cQIopI6jt4irV6CCAaenB0WfkLIBm5Aze4o
qSzEDl2TocFakNr900L8hiV0Kip0dHAx81QLnl6aJrX0PI/yu0Pe1ckjf5WEH4bO
xm/htWdQgELnWEZUFDuBJTLetqyBqSkOh4S9vR7ybcJymeDcDoVAxRHES/Z9IPUR
u+U3wrWZRWgA9UYOXWO/ocA6gcApNylgI8ov4V6Oe/obdBBDPr9XcV6MoHYkArWc
b39bWMvomtlJlc/VzRdT3dOw8ON+RfY9hcduEYV0dit4JSDeV1zV1V3evTjKer+a
lfN2tVtzHuixflgGVgq5VYk2URr0AXpK98/klk/LFDWDubC0LA+FqUQiwJCobrZ4
fulUtRq8Ehb0ocBVK6/x2xK3iZwYJ7SnIM92taR7DVdLCefpxBArwUtf7UJQzpZJ
S+n9CUCEh2hK/Rmf69+/0mRhate+b8/mcogi43VynV/rc8yqrVLJBaKK0NOFlByB
2mj5A+lcOHVtzJ0wXYuhUjmdF9XV6tdPfIDwA10KCIMszYmf/8okAsUv89WsO7iE
hJif+TBt0vMWyuhGAnbbBVf17upJageDbcuwl10dmdicjYtw8mglSVy0dOPlEfQ5
LcEf0gUI9ll4t8Ed+p4VZWfSnBKROtlzR6i0rAqyt1qgXG8wj/8yTDIEcPAl2RS6
pmgnUQtStg/5ul1gC2ow9p4gzCVr+o7o7w0ERYOW/TEYhrGVg7szID9WaFaLCt/9
r3a06IS145KqKLfYtbA9RbVpO3M6Ccg6M4w3hAyPpgTLvT95CgPBs+m1luxFWbsB
P66jka+jDkwyHyjoSMZ5/mLnvscTAfdNr5B5TkSCu7lnFhbsuN+vkcqu/j/eRnSw
wf+Sd32jqRNJ1TnyeIed23MhFaPC3S5v/PxqHoAXQgyL2agT3d0KfZbNvHokogRN
RI+AI5+CkhMm2oSSXgNMrZkKW6iLoHfgaGp9hFwJ+p5/0J68O3VYcPvlfEz4rHk6
M/sBRnPgjC4dTeVeR9aWn4PWoEGyjGk8sk3jfvYS9Q8hp1/I8n0u1KuLofEhDHyS
0F4tt9i0NmY58iwAbBDr7R74c2tzhAGR5TeB10sEXOQ0nvhrXvxKpcYc9AV84kwG
PmYLv/xFsVSg8L7IFf5KphDExlDqvEOSWaf/W+/9rwESq85PJd1jXtpzaPRrjVfw
/fRlYK7vailgtBHOhGsA8j057QGBZ8ThRmckYmZI9vz7zyVj48jLHRAuWhYiTf5K
5zYo0DsnVkBlJ0N7i/KNBxQdTOnwIhmM4vEsXvJnGG6CSeM4jD6d7A31FcKEsOKG
OazajD73gYHO+EKHel3dLMGHltUnNNMEg5soJxVpaHPFTKWUsD29bZyF9zdUPShC
zlv8SlJVWQXgYgRB2FXjFLss1m30TNPmyW9+nmivK3FO4kQloE+B4/pa097DsPS3
og/vlnboKdSmnYaoI4LYGAi1U1rPm6XKNR0cvWgrJQrgntbdrk343nHLkcEymVVa
xENwVXP0ts865a1mBRI7wjNAPuy5obhgORVUpbDr210Xo/0hbTl5Y4FHnVjnb/1L
cM4E06tsoDxWWSFbLWV8DLFdMIP+seDWlAsxlF/wsOGiCLD8LXHUNpxjIP02aTfB
Dt4xH1yhLqBYil2zKs6MHpVXuVDOcfH8exnhAjwFBGTHFwrWLWlFFnbMDZccYreo
7jiGvm52389pacM0onrjdxDyTzwa3fvgVTdKkKyA1kRX29VlxgDYD943QH1k/INc
jMdfcT7hM0RqCsI9Vm3PYzVby6SE0QqkM1VMt3Gk3QqkJp8sI4zPGaYvG0km2lhq
F7btVLUkF0nXsx8Yrt3d0yaTipUhDTs+Q1ZiXU60zGdBULQhO9xwfqOn3ui/5ycs
flACrUkKEoc28WkP1t025esPTwHTvwHySYZa4vBOVvx68ndD9BVqOtmxteGd5uoF
a9wu3U5PlOTRsT2432LBcakDOwXM674oq4RWimF/KcLeDzXrvDcWfQXc952uy1fp
bZg8f6PLThJBT7C6DzbZ4WwAKnMdXE7JiWyQrgtn6ighDfM/VW6ZPSThA8vU1lC7
LbYL9w3J0aB+mvK+adh0vdPJ/iDQ03PHyQZtPFDf6WkBkZHiAusRI4Gucejdytx5
1JZLDV7BnAQ8oKAPncJXudUW58hcEjaNJQhKl6nlWENc86agrEph6TgfHPQFObhq
Jamg758s1pz9bYOupOsaGI138SdPC504LqJbrVEZoxm/Bchfj4zExTh+TfwKU3eB
OS7xicRzq03fdkW9kHaP5+URp3TbHwCAgXsJ/htuJ8C2Y+SmJzuIgvf5Bmwtu6DQ
gdI+FR1nlLJdI1hqwAeDfoZ5MhRdTu9MHcAUYvQobvDxkRvxJYOvRC74U6yAhGZl
HoczVp/0oOztj2P/yrtzUT6BQs3xS01G3lPPzecO5pkpa/JpH9TH+QLPBfhPWf5Q
o0DpuwV+MJFlGGV7vHmLUvfgz21pPIVThFkFfw4PovdHPaMFpGfJWAwM6B1HQfLS
sr+aK0IshzLIUlQQdqkYNVm/HeJFWcq0OU1wTZ0BaT+gNvl1a/pdd+7pl5keUGYN
1oB00PCXyPOTJ0Yl+TLiupUYW7i1alwG0SlLTQBX1jM2XZvIE9Nzw10j/XReGKRs
B17QRBqEwEY/iMal2KoZQmJodXXj6b7NZSACW2rYxY8h2p41LSqbothBTUo243EE
Wpz82GC4dlg+84Watwd9Ds9xIHg2w5vadKcrpI+1+CqL2pAxgS1t0q4MwF+fWsHi
mWFBXCx1EotjqrDlW8lTx7QW5ucPs0dSsDVPMSbehAevHmz6xOULU/8SUMqec2m1
6TgjT5nB6HUtiV9KpTzEgSxQXE39fY1+Bm/LssApVvqYEe1dCUaNBPjjXm4dedQq
t8Kk0w/SLeO0dsRDMRwAW0+7W/UzQX1/RMLVzNCM2J0SwlxdKxD5S6QEn9v2kys1
cjby+k2FjdtrLXfJ+gjcpVoyl/tygfeXcE/JRROat/tQswdyyi9dX8286CiSwt7J
pT0ipGOTDxL4KJEHke9YIJsyzPzOnaotwJN77g+vEMlztrPtBJeumkUYirVATepI
/gf1yO9WZBbMgcXMUs0nIf6X7O9wpgnbFyLAbApFqs93yVDPvg+1iIIGGJZSpXgC
IAbjUR+5Z1AMc2UQT6ORZgW2ASzJJVQaapCHElY8Rl5Q2S+dfOhkJu3kRVrW+lR9
F35VbPLj47zP7ikzRJ+73vbjxx+8BHfBruHkaKisfM2PZxOxEsnRNOAIk5k8KwQr
c/yIYI928S9DaRb20qtmLM0kHGdDgfFPt9mNTAcLt6T7Yo++iRgRhQBj6ZmG6ilC
8ZZh4KhdHFT8eJE+jZ7imFRyVD2A8tkAFPRyhHE/o3NoQU79+eF6jO0kphGJj2E/
gwhzBo1CzKrVEmTSbiMQlSVyX85sFNziMVxQ3S4vpNVYhwAQQtI4ZXjJ78E3bYd2
NEchGBOK6S9PQyEa8IMtqnDK4kmJbfkJPySKHy3lAeElSYz7JGDIwiQPDms6Snml
1ZrpkM72kbanU2+XaET5yJz9yKIziNNWhPxVMgbIEO/CB2TrlLS2EWnM17eCnE1k
QTwaxUUjhDa06xwFmRgvl0C1cOXkhY8lEfeJ4RTeyvnpmTJmM0li2TW6njxaEndp
+zgTHym0QsnqxvOJlog+lDJyxLGNz3d+vO7sMatslo3+fFawdnYrzoGUinR7rYU3
A85ZYJlIQZ1WgcQ/1b6KFpcfERRGorReZVAsQSjSDVH4fkZkc+kBCy3kh3n/TbGW
z3yEwQRt2hvdTNTMbmpVMxjbekAh0gB/yThX4y6E3j4v//+z06B41bwoxV5qb0o4
SeB/LuOq8Nb1sRLy2mj7Uf0VJvFXn9Y3EopsnZnpyYbLOjlUISDTImswOkPln8IT
+ZMR49Kc+WERos+UnO4lQGr5KXpvT4nDECFRPbymL7gYehiCUrGaJ3W0j/o5FPdR
CwTDc7Dwdk9Xa1Luqs7l40EWSafdnuJOYJP6wqNL30Y9TYtXD4q/1N3cA2ulooD3
ad14ULNf+/tybiCx/s2rsqmtmD6ErMyMgnBScaYxy56ae6eRO6RXw6SSUbE0XNuu
U336EnvJLiOVcdykiTENpnvm6gJyp9m+qE4DOxkJaX2YwLbp3MX9WLuvS6N/V6os
SG1//6/1lpXyHivP/MrTClXPlwNrrZcLQZurSrOHYacVsibLsBIZ7E6xKC06vv3P
X8nDco6OtDKOVBrVfKDuJ4yQ+jl+fwu6K4+HHPeksZ5hNH0Ke0iMh8A+UYigyXk7
O2Zp2hB/WthUqdZshRAtmt0WiUz4ufg9AMEDNVaUEcF1eDhBU9oqOVy/rNAL3MbG
6xuZ28P3Dw9AfFoxdRoVDzPvUHLTsArD9a5JrHVnt97FgRlytS0i3s4I2nzzoNT8
Z86+2NbpJIkvY3RMDPHja5wXk7nwmrW6DdXNnFvMUJIL58g7XF0/IrOQsgiztkc3
9rJFNjNMTx0IWmpEhuG3zY9sgUbfG8eNRLSCoKsYgF56YHI0fbaT98QhiThWzFqd
OuEhF1EC9wLvEuM7hgV+VhnewD4uIXhWTToOtFrsUu6VMDZceHG99z5sIkM2RJmj
kvwRbk9hKdtafxCUcsUhOygDWWoMCW6XLW6DcQn0D93e0x2n7BFctb+iiywr+Gw3
tJg7CU/XP8NqcZUJV/Q8e5Gjjqhi5ygXtSuHp9PP3lH/PQbASqLRIVSXLw9LXJtS
XaBktlsmhjzKxyGYz2mY48o9Mp2yZO2E/v50PWPMoK6Uk/Z0fD8MU6susxbxn7oW
jXugRXdlp2LU5bmL7BjW1Is5dEDw7FnGGYk9YHcmB1GO/DH4o6k5L3GOvgaiIewk
9QQK1VbLjlKQ2s27eRfisbOf/l/M2vP6V/plSGVUdcpmzkd/y5bGRW2Iw17jf4fb
MMGQ2LmhKF7kWMRJc/LEl0guxznr2LEcyFHdhJget2ceHmia0gKNH4PAx/hkUS00
vR0GXOQSzkNAK7pC9IxBXFs7PpGbbr5XOrEYiQFzZ4ZMAp/L69VdxcroPetD7ME3
dIKOwKai/DY26d520Aqoh87+c1tv2ui1W17BJqll6rHRYlGhdd0XYZejUOSypXJ6
4i/LjztqitAvXyg+qTMuu3RwWsI+qIeye0b/xJYkQFUBBNK5l2qF1IjxFHoVSHXr
tx0F2vUn9H3skKFJO39y9b/XRApife3UKidD4eoj/pS79zFUrm1lyYI8xT730Q/6
AB6tlGZUmAuW0wC5NKNMtbu4q00dvKxCSx82HsS2MOOwNg3OVHo1vhB1f7l5ufQH
w9ieLCHjF8ZxbhzSNyeMGZiZ2x0RdZVwKm6O8e//K8qNx/BwJfFuWEGERgGHZ2ly
Ht00j+OPnHgEsuDu3oCqPPtYCZkWhWbKlv45CnjMDpjU6dv7Bt9H9YizQZyxMiEy
Lkq0w81E7pXn6OU/PazjF2Fz3k44UYTwVAbxYbPLSSQlPaeRAophUlnx3sGOkIBj
tcyUH7bvppDuI7DrKmIzbvnhZN4LrK+7M3nr2O/ojBY4EwtjEDnbMdZpN58oAImv
PWYWnc3APH7ctq6Euxrei44PH72PpR6mF8ZTlBB4ZMdEjQstZRV0UrKM7G5uqWRG
0I1JP7c8wX6SCnwD/6BmMs2ymbNcRIyiYQA6oMaftCJ4yB7257bmWtzOZ2PqIXv+
T2ee8vy3jtct2z+amzazSOFdfXDzNNMPeMgY7VNBi0CGbD42H95zZUcsvBKH4bk0
LrAYCFWnnH2+TBsG3owbBTU8p7IrkyMlpkyPRRtvIDkeG8AL9QKvh8cQqzS7hapd
yUK3p2am9v44rXwsQn79+UQJEVdnYGHxFCurcSVpNwiBCfyw4qpF+M9caF6KyHQA
DemjoPAS+b/EYSG5vKgsmwGjWPGAZLAbDEwXWaskz22XDyOydCagPpFntWCGA+fQ
QYM0j/gHUIefa2jd/eVqY2ykilMf3bpEb/xc5Z3O6GCG4ORmIL/2OKCLlRIBl1Tb
QNEZ6v7gZbz4YD7iSfnmURWTCBa6RALZHqMDlKfz5rSRXYvgQddYmgKDQUfbIBUY
gCIaKhRtb0UxpqjbBxj/TyaxMLpsNIVFCfS/9iYK2Ido4fmHAaylt9BENKDgEUny
MMpMJ5PDzThd3L6ys4rWmBDkYCnumOGzi7uLBH/EqYRUPEeam1vf48i1gVMTvsc+
qNpIIVXL7Ej192nr1+l7IpXZqn66I048pXsEC98tAw7i1UZPlKzXYsN269lwtTkU
+HElcUKSP17t0gb3SPOgzvng9qws5yvZklMLqu1YQCQwRh3mzwL0YXKodUI6ljd2
M6yvMldq3/b03+DPFj2q2DPhEJOy3UHw17DRQpo/q1QQSFh9HmnzD6XZoFzluqdn
dBzzbgX3cYsORQe/zGZqCo7lvsnV289wuIdyRzuxPNZ2Z/9yuJ3ZGPTarGMpwzKV
2Ao779CGePESYvcDDvBd/21FMn/HsUEsIUpGqigf1F+Quj2v9DCttP2wjTcWDiR+
p3LxTbeUT53kx/GwK3XrtRAia3kHpSSF5XOSCQRJbp684t2wg1At9OJxE8LKzWe2
BYNopaaCXh6aWOXkkJ/eGYLaarCCXhRBjZhVb2gtcV98/0dng7ac2BbNEUmm1c2J
nEDEg3CAUXWdFHOhZBYa472pYwop8lYLyYsbA/32ItOt2tGFQjSzs4dUkGZ5Kjnl
b7RQVAQHk/IYmk1ocOY4W0QRzQ3gDTRUbP45Y7kUME3wOinUPqHFXqgHnJ6xWWd6
hcUem8L7aUmV92JYg1RpeUz+6FDf6lpv9p6Z7BC9AcYQBndLku6ECtOKxytqmXVr
8dqksxWwyxvS8cIFHaIKpbglD8vB3y7HBddSxRHBp/h2C9YyiBtMMxVjO+7pIDDH
H/csqZeITpilr4EtUWnH0XeD5k2Kd0VViyqZgQpep7TV9fu5DiVCtU/dGl6alVcG
CrkN0gZxqmCBgAO0sIWFWjHlY5FeY28/buWpZoVmLOudigDhH8BgGbQlkBBYpgXu
l2awvuiYoDTC7J2JHqBmjH1gbSNUz3558REJQRSZAp0PZ/sZmDb0FihHMWQGEafa
5+tMs7oikd9Ec1V6xs+NNTruBtTlat8RsUkbzgZhNDWxJm+V4GNvMqzISbd/GZno
epLMOmO0oa59pFxHkcFbWY4mOrYwyqPWyNfXB/Z1FaV20HyCoe7sAQ6ZARfH97AW
4Qkhxg8j54p/kThYV96W9l1UoiWOW4aG9gmJNDbVVWGNeHGVgYg1bhXJ0fbzC3AI
0mSflvl6IUS6KOu01auH19ZzyKMZt9KhVrGX468Lv8EoscpQmoUjoWB6PTSo8Vuy
50lAzbMT/WBoBk6L9ofkIcTQr5TOAzKBrcNRiPjsmHGcZL4WrdRuFjwSQU58JXxb
i3yX7tN/5x2f6u1B8KlIhITRE/MR3Ri+toEOtHI8MpNVvGLMPN+aPloo2+gVt+Gu
7G8E4ayEoa8VmO2jmqpoaMty5XKIV2hmbXsfKhkOwMdxzPetTkK53tC6TS6T8Qbu
MCRoHZpDEOAWuvf6T2yUcks8zE80KkY7tIyUwrJCtGlZLplOVt51StJ4u7DcoMqw
VUVDlg898GXUIIuOQR+lrpeE5XkoUJPxAWq5vGnsP/ZTNsZUhADdZWJ+SlulQWAE
u3SO/ZiertedVtIfoCVuRZAhiihQIp9Osm+xtid3QgLUPPpWzvRsoNT9X3dpTC97
kpl8LQWxQsBsDvio1nSqYr2hUIEpsnnWrGm3IA127veeSSxrc9REjctrjPwUJtzn
XELSE8F99Rtsnw3KwOgPX56xPAZ55V2CjAk4ozLJvLdFd4BSIavPx5hdgnGQlMPN
8k9jKa+6TJBZcGaF3bIFn/1xxgjFuUQaCLOcLTbjAd8SY25Czz02er3ITAq0uDmv
0/0jbCFdQfLnmjDLgbnOLNmZ5kBg+qBmwBuK//JFSU/z1EkuhlGDbV/1BLfjIscZ
Tb5emS1dWLGNCVXa0w+HP8iWuKCl2LwpW7MWJf1RVv29j6U5ZKOiBOiXfJe7mItN
tZx4P72w2rnC/OKPNkS3/97vDK5G0+tmOPhDvkoM/HnPHDSK28p5YGfx/X/uxlkA
kq7jQOq6Q2Pb35LfEkrWTlq0QYizXckBPPXHkIEEnPnSzAON6JNxGHHrElvrRXpo
p0hEk7RLxsIKLs/rbUsZSz5FpXdxh3dCraYQUnRWWnhYxbDj3jXecuvgjt5KQWNd
c1J5Q9QRZYg/sYnhf6Gmij3XWEX+tWe2lKwofHWhzV7m1+DLz40gMJ/UtikqrzhN
qBBmQdemh8YZQblfGVLLc2bcf7WMpuZ3msXOpfNwIOGGM9jLfqRoadS049MqNSHS
KU7TcVotaYzaBUQqmEBiVZo7b3uNj7UgKOi1dkFYIHfT1APO3Y9xFVC9hmLgDrWb
3sww14/d1ilcGToODjUhkwThC0dKMW3R+ILb0vVZHxGKzt/mqr/BWC++TOVYoe2h
DdVQrN5ovcBPARZkqAmojqZiW7AIAIL2aZQ81QRfo9dM3T1hl9DK8T83/0rpNcUh
o+OVw9EAe2zu8jm3ve8+Q67cVV5kbIwF6qljEzU0mUwhBsRxQKEHat3e1gu0FL0O
k6uCwgbaQkRVkYk5m2hS89BUcyn4AQ+fiiYXESDkb5my33J7z/JCO0vbrbwzp3+5
HR3kr5t/uvf5Yr9B4unPRDCw1dcSjmnZJCj9Sl6ed0XLl+8eX1d6lcHMQN/P3SWU
X3pf9RXcYwv9w2vq4MvkBaY69mpLnne5+EdYBonqZalMIvoUaNIyEI9dg3zHk5UK
NwCZyVzPuyrbmFDCKG4YEmWYgCpvzBgZLsGFNShK9XsWmrsr/1wfR/iZzwY14qpX
g9sKHOeHk53JQ47Bh1g6qJSQa1fPWJiwVVw0BhvGDJL8AF6ABQvXrSR3J6DyoBgL
km3NOpYGaYqyETItfF+CTJb0dcA06fRCUu2a6Mz/+0eieabbdla6cKLtnlPE0KB0
WflPutoz3BDOhFPVkq/lesFXXXGKPGx1g8kwuOvFBEsGUUo9idRF03Oqg2ARbm1E
6RMEdLjKY8XNsB2hBGUZSzk9/jQKRjnVRNGtNPxY4YbnzcA0kCviZX018NVJhwt+
ZpGDiEPu2zy2fQZE91JtaPlwRk9T/A9B1wjGe36bQUTBzQNe+RQp8pnk7Pp9y8MX
+1504gvIJNTxv+qQSXvTsqSd9jf8OofQRaoXZuXCYM1qWtLqXAAXK1SCZNivW9Ml
Ii+rx6meDNgOxyYIh/kkephkhEJH926E0XXzH3gHwRLPvxeBrXetIf6xSyAFMe30
kQpIphM5Qa/DgVfaWQnfohrOIJQuBzUle0YKU5S7V1rwrvRBW5v+rZYvT1QX0T91
apt7CeG2wwKdqWXtXU6xTuLasL+IzSrt0t4/G7VqQbRPF5Jb9fT2kKINes1Nds7r
BRvKUKCujJAXMIH4cpAl7krKqF+2ydOxS5yRP3Nek5E9nnnrChPe4aAHoK5HG4Sz
iwDuwejIEq/Irh9K6dCdGMVjC/HdgclqFG5oT5rp1Xi0UomWV+Lv/ebmiJ8uL25w
T0Td602Sgrf/sfJSHtwhbTia+5Y42CBPRjJxZsNZqDzff23/Q9SGlG/LhgpBRPak
v/RC3crg5Fx21uL+flHatjz2WgqCeOol9IRn11WFSP9lsFB4Z9nylCii0M+Kxi9M
2M60nTDLJsB7y3WV6dEwOiU9p+x/iFhtHgMzJHNCFml02OaiEX4v2XPzsOv0oqQe
4GyY82+ajKIGM1KsLXf6remuQuB+xUXntETV29CkACdLVoB+LRuspg5cmotVYM/x
Y7lnAH5JHRoYlusw1f+4hyFZdWFKRlr2cy1rPn44jvKAeuLmgC5c7vLYojfKmJKR
lOJd6MV+nPpbD1DVYFcG7QBaA/+Ixzt8Vb0qwWeO/4qhNp2P2dlRGaupGGuVnJID
IHdOgMlzW5kUo1GClC4i8tVMgi4jq/NMEmr9wF3zQ5jaSpggeHXpqHjLsIDJOxcZ
J/NF9GzARhr96gqlRDP09zZqC92XW8PR8+H6zP0O3BWa1Sqy8iGtvex4pyrUPnEX
XKZbpLPQ3PlXqGPux4WaTWh67N4rs0h0bpdbsaoqCOB0AMujFW5EzJUmhMpHrFNz
1dC/7vJPyZ58PJ9/n3jeZXBP6AtJgxTbSruzWKF6TOkdk5MI7QbtfGT/lYw79bdy
1foxGR7kzOVYEK/FdH2tmzbUkvyoGdXpfZbK58OMLp1bnXLboF868DmJ1gQYE/M1
JYZv71rIPm8rUNf1lIoa1d63jpx256uavZp/3QwNgpuU+6NdvnS3FLP8LR9U+9mZ
oLPxiAgQ7U13JCWuWCiiYkVV1Gftp/XvQNTWi3otpNpfwatzLBhGyxjcksbjCPGc
u7Qrg/qCz10OKcPHP8tAWGO4RWvouvYEGXZUrQGB2xbvc9Qc8ssvGFFbYzSWtDXg
tvxcouQ0SFRMojFiPCjbs69SyGHY+qA8B3k0BI0T1p1qeMieSIzwcCtZGCQXRWUK
OKCxKrCpmflTLzi+5OkSN7Q7QSFPf3LO/+7sVOJKOahyis+ipRxOfUaCgQ0CSjup
6aJSZBAHGeD/Geod6vb2E68gUnEP0NAvLFfjZ4SXNKPrYJVqrnkfX9TKby9CukJa
zmGm+c2BcA25PI/L6EW27wgICVEXwZPVT6u3YTcC88nkiqhkdSpHQ8xkLI3LhWzh
hDT1mR8eP14NUMkfBAuuGMnhNYAYyX5szn/YpREYYHg3ovA2+1vr4skrFilGGWMQ
Pi6s6F/H6YS+xa/Q4fjbYg14xaBbTDm8hCBaMRjf1KKjDDLZq//IuBqVJwawFgON
3GYc3/jWWg6Grzd1MdSRwmGeCp8r3D2kznWDsWAUQd4unEyiUZmyZLRteueAHz89
As0W0UOI9L2oAto2X/CRT7cdUGNdztXjbJvd54eqoKEL54NFKmBlsrtWAippkYYv
3lz8hdd1lmGDX0mbpLkDvMFmWiks0f7sMELJFY7k4Z+i/Ivx6kJpSsrcNjcuDA8q
JUrEHkDAgCPcuXbIdRnJrpiJJRW5Y1xtzCLdtIZ0rFgsVrAIVAy2APymXO3DRaJA
qwcllIk23GY2Gn8M49aZjihnVUw+0roWfLk3edh5AFrn9GLt+6ASEQ2oV8GWSREp
xi34/bw9ZeMpCru54WOfDf3sOK4ZxuFDcqgkLK3ScbmDrq1adLc2hhdRi76qM1xy
aDYU8+NfGE6gsx2XWOXP1sfx1OzMmlkvCeJd/xLIc/muDMHq8bsmsbwt5dXpysRR
zKNoOC5yKL/JSILbCTiyk53RWRISEwC/xyQFfw4WLHKaTmXQVbSgWocKk9qcKqP+
fjMH2nEZRWRt+7DbYhmoQx6uXa0jvgtwjGN2p13Gxs2jatQjbuDdkJd/9Ryk3KV+
cqa95YEJdfzLHWGXJW3GhD7IkpvV99ssiPvL2rbun99lxWRfVRQ1zpq7yPxg6MIT
WbPKgWxRvJ8sDuVp88sz880XzuzLEaK9vyKObXX+HY0qSrVL7vgpZ56FtxFSuUdH
Hw0J0ysVvFA/TxV1yd0Quph9CkDnePB75HeMwPJvT2DuZH0D9Oyn0nxuA1hgwbIK
kVNxv/JL8D5UcsXDPoDud3dUmeaENHXbbUWdJU35h15Wl9cjawk+PXjemFo3xITp
RRqRgxQnzBeIwtNjnZQpvO8cVeePzwjnMR/MufQIrAG6p4UI+TOoHz35jggS41xk
WuJ5shz/Y9H7X6j+6cMESfMdoOBtOUZI30/vWK/lGohpKVfWD0fUnTVZQq+GAC48
l41YjxKd+06cHroObydtUkjHAYsiV9sR7gKSsvJQ6H3Ua38Q9GCuqBV+tHPE0b2K
p8izma6d6STuIbCAXkQSzwK79tuhyZStIJ0tJzA1lIVpz937ggo3LxZ2Kb0YAIV5
9d8fj7/6CCzbGggqsBpfiANOPkiPQUVN9Jp475xVe0f22gNQStJ0iQJd8ZM9lMxW
FPn8F2CPQZZMsXxEwylIdSUuyuXVygkSXvAQ6hpr7fOHSjue4Qi4om9FM25btA1o
9IhGldRyH1df3X3JGIvY2FOr3QI/QZvBDcKNpS+b84z9J1tB7ADew9LtJGd+G9aX
YqJmAoCC3MtGZtE2GkPpRH2/hBR8gjsUu2GhefTmMpp+tJZXrh6xcOMgzGyJZTS5
BrKO/W6kS7anUvM7qjC6S4ui0uj4P2FO8jig2sw1/jWkVr9R/p7ps+e2Ew8J30lA
JHVxt1DHzpI5OcR9xzYekA6VEYVvWbd+iCGWyObJWBv5LrD86c457xjz5cKASEO0
X48jlWqSbHlJEsd2hVLT3CeLHnHlfWxltv0x1jAKktftJoJSYkr4Hf0kJZzY1g81
rdVNf2oG8SDnTco6l+8tlddRPUFvJtfd5qCyHTAPzaYCP0khmUH27pBEVCtvGiNr
gunKBW9Ztjwkck27G+3b8VTvy+33dUT7hR68DRI4QrcgHOEg8LEkhxkBKBbwwjnc
bjXh7QnlJyjtTyxcU+uv4uG0UiyU6aqplphHZ2h+mWWLmrEZvcIbWxmzJ/Cqu58e
XFvb9Kc/qOFPry2m5R3U23QgNTX/DG/AewLv5XT6tc3h+PB3N0G0g+LZQu/riUUz
Qgtf9j0INx6muNq6oakyLNRxLRMkgIzb5kCR0cZbhtL8LbMbpu//MNxKA3ddjR4P
luhddISHC8KQunE1LIB0yqeILLqzpc7XbArvalZkIYgZnfhac4hGmGuTiTbcpbq7
tLtiYxTszssberT/5eMzlRSlsgnaLVsxZsKeV40NROM8TE7Lbh2ZozcG38ilBgnE
CJpmgX1HFh7K76l8AmPhV+D8LwTeur+f0BtgTo8cl9X8oDwrnO2QdHVHEMuoCU4C
htPClXtw7DQjKdM4jVYTBvdoHtcI060KN1ylhIavBuRJo+TtPv0GltGwIG5EjISJ
3yKK6gkPgZnnnlc38tzoB3cOKtbMd7itfstek+/yDKM3rZFHIdO+eSiF99kC1yCD
8g96+FTZfAsKQkBU6367fJ1HF0jHOgiPwAYZFUtO91zIQlZfY8S1flcJm7B0orv2
JnjXH7WDLyB2A+YhEqQ8xWDt/Qz5Zc5jKCocDAg8ipf6guwK2wirFOE3qG79MR0J
2TG+0wYrwqfA01TBMYC3wYwlPb2RbBbTrR0f0wTf2Y/DwmyH21vYnn7/cb7WVyfK
Grl89zsGpVtl2KorzTKYCqK5qfvxpv4tfDfoldsrDWJ54b0pRMB71svkwWOtGiaX
7dHiThHvhRQSf7jwM3zGKu0N+tV3zP7Hb+J25t0Z/x6QJqU0hziwhtrbsf8LJ8p4
PjEhoEXb8Mb0Hn4zFaoLbDuQgeA6vqO7zvUssBK2nheQIsGyVS8eeLToFjACLqTE
QnWKEyy0jbbjaNIS2EQyd0BzTWRJbW9TjCqhmjEOQd3aMZA3kEt125j9o6fOeBuz
b7wS/IFTdagSUkyPjjMwRxWo9xmdb6CT13rLSt2Oxm2tVozDFdLaK2ahpiv030EP
WFZsY4ADMbgtMSNa235ADWYvjEJOxBD1+RHNbqzQ6hgiOuPZdDV9BTbseth3bq1m
LzvcmXcGJrmD1gopioHiEmAaQTC/wUX4pXZAkJtdNqB09/EMghD7y99pqcOZC36w
LQi3i4X5UqH0T8qTlEL72AAQt+bw5DbJxhfizgM/n0RiompgWQxxiBrknk+IDPjw
2pS7EOyFMI10lltZ2ik9U4mBHDCEjiGpp3WwpO7oNeuv0BxDAco32RorYbLKsfqr
VM+aq4Djtl4IbBgSeZTXqWpHhdMFe4FqRHpYxes9qyInrgL7Cjo0NLCvZ5ElDpVU
9uc1N7xtLGyzbRDIHAvYnOCn1YgL+VtC1yGI6kCVnlGpmIfS83yrQe8skv/qA2fr
jf/6nepB7xT+FY1aw9Vo/PHnzBfKiXMauDCFTqrCLDKPAoFCzfPuAYcSqDkJnfLl
d98OY1Af1uJbB4QXt7EvLEiXxK9wDo0dVKHhFR0cPkjf8lU5GVlWf+7zJAdOHwYc
9S8KMSvEszfrKSFkWZOmwQt7drSmImF70XlSp6/oBzdLDNWcX2Bn/mUxLEA2bYcb
J0WY2T4aursJnxyI30PDRLMtfwdLCqjEaFmib68h9uqLHxLyiSZ5GxY/FDY9QFbG
Qk0ulAn8O3TOyBWe3mqbfi+Ih+nnyH1AKJWwLd3c6Uc3FNKQt40MtM75IUGrVUdx
os5RNhCw+nHpZI7e9Oyb1LE8nP9n7irwt5A0NFigXfxB7ZETbftu+ki4HrpSWLhI
h+mF3RCXjD04lSPFDRqs+0GU916fBtS8Mlh1rsMineGXQ5VoxT7cBgEa7MWBeiJS
k5ymoMQPCwISGPMua/MzJzS2JNelIXiOmcg6v27fnZUjczzEy9bytGMG2Kv5Exet
slUkIilAbc7TtExxYUl1O/F+v0UWdeV4sfhIRoXgPd0I/gR/BZAb+M/or5B5H0/l
w704ngTX/MfNird8BR+3voLHLFTiAyEv5tSIZq3sx/EmUjuXD11QIUT7EjsCj2DX
BUfPtyZIkAfZGWWhD2exmvFSaxOaeF7b7AXt/EToYiyrRzuV0SBPc6y1+bCrN96p
Tb5euBRApYlalX+u5fl/zjOevSVYU9M/xtY2UA097JBRnoxz3kP8WqepGNKM5Fw6
oBv8ImTRoMDfcDBVaQsU6Qmg4IhrYd3xV01aRO8jfwYw1h98VzF/oYyc5Tp8AZrm
D+UbuwtZFzqLJGnO5VCupXpEgS4Re56l8Od9fuhhQRlQkf09HmZRFhzO1TLUjcrs
uaLKQSnN1EIW60ChybQbFHm4RiIRJS861F5QV++tbhFHnWgf+0nGLcPlurnsJ4g9
aUnxSgvqTB3wK17NWgrO/BKBgp3BLqqQMqgJjKTMLFWmLWx+78SsnXwd/y4a5NBW
AguuzVBgcf4OhTDQL9vRq2MjVntcdgVnjqgr04cC2AQy3ZYDungOuZvnMf68nrpE
yxIGXL36Z3YCgWp3h2btYk5i0A74hzrH5Hgd11wULr9iRs3k506t9/xiyMu/KpzW
GVxAXxpMFtkbF87aTadw1ecNadKjigK25AROxJXEwoghturgb5GZDEISAflZPPvo
ZdxFNDfUVo/OLYENvZRkeF6ZXm0RFXwL+cqy/LGuBFeT5AkyE7d6zS+orGrIOug5
tQed0Z799ob8LfM/YrF+AUS5wBHodW7OgrJ5fvUTSnG6LmYAdA3ErienEr5W2/g5
Ufv0VKL/4kczwtWNEcpS/I8COl4sIoA7cbtlZhTbaVIb59BoTKwFtLzabPwZ/TpW
4TtGWa4xs/BZTiC4UNJ9ULVyqTyPm1HYlvhy3KzSOHtI9cMku0A3XeOvbACBCil8
6PHUUZ4qrinnx+r4qu2oZhX+ciWM5eRxdHL279KHLgSVfaun4Dw0S8UtFmeG0xQ6
vPk4vfKC5oE74R+Nym9lLJe17smpSsWOJ9A4s6bkpsJyeKb4um9bk0j81dvyY1d4
Szumhay99yatPs/xryaiPT2qJq/00yuYXo+vbk3tS+QCi93LVv+KgzMkgKOPC6FO
nhRRamZo28+3KOrWT5uhPClBPJXrAjN6iG88UhDIhvIbOQxn26xA2/gPn3QSX5Xc
5upa84iIrGXEcO2+fAl10ONONiXLhxB2AW5f7wyapZXggBe7K8g3Jas2EX2tkjTH
MsdvHJpx8Y7NY8Y0+xmSRj9mmWsw87zWm7wKW2d5KQDOi6oY9lvYAQoiWirs+46l
I92XF/hUXmwlZVCAxmWoCV4/E3/2xvA2aLX0nGxyOGXvPvvwiVa+1TEWy1QqTRq4
qswBpqZPc+UDLHd5PR1kkbzRZzBlnLqh/YBjsTK1oE2UohgbiDUwdkQ993X1kwSF
coFQS0IcnGq83p17YbkEeEyafSl98th2lDLMbSkcg+GOKEyZkcnPoSheEg8NPAWt
jTsdsI9Mhf4sMd/ANR0DLsU2WnfzMB3iS7W9b2GAuVmS9XYBsi1nrn0pJrS5uF/3
U6hLdQNyvVboBTKe44S5YpEl3Ag/vFKx68/frg2kcnu4OEPwpHixbSdqxtA4TySp
wOIPFDjI7uXT0Copw1RadOLiyjJmiUnsgamSMFNNGkThzPVxJxLFjRYwOTiEqZV3
9K8IE3/TTPng++YcFlpCF1eV3qFBpsORox4s/vPsz/TV+UNzH6c4OcD7W/jY8wW2
NGsGtxKmSD0lo+XRieYORPqEzlgqGe0e0Q2LtSAqnA9aAIQ++g9mS5u3F6Efdm4I
eDfXbsFn8mvIpvzqhq7xACRuglTicbJ35BvH7KaI8NU51bbycNW1wuBuAS6Kt5GQ
yQjea5vuZ0fgadsDXaPGiAuPm+i1KUwJFhYZjzdQtNj7deIOXHiBu5q5wT8XYr0O
r/5wCGpDdy7OZqa3ikNGizOhz1938Cxt9KFKKTIw67rQjYdzscZReBNiJkrqki6O
KB35olpaj5DMT8pjebrueb4/dJqaV/OyKyBVEHM6ndXqa4iNXSPXIGXVbz+UU9Wv
km6dVjuqZcW3Jj1anGkVyB80JcgdnS1BioOg69m5/m5lsUmZWRcuxYS8Z7IBNSFU
sDoyvySsGkw5Bhm/+nNeZdGzwcj6BrXAAAS/8E1T0r8Nv8lf6/CqZPd7AhbzjTbI
jH+ba1Y8iZDvOxo/LXUMI1Bcvwt3B7jU9iNNIXnKJMYQp/Wy3mTmO8KH6UjPlUe6
Mb57FtacjugwNJqwYmkKT67NnX55VVrszG5Gq9zLO+6+AkjDHt0RIY8s4DIFMw/w
JXGHbs6Z4m8XYfYjCXT02VyHPD3o/1tG1nEu6VgAnfuBZsuJg9+Cwk3t5EeGTisK
9QghkyEjP8mbBvg6x8bEt7yg5eW0G1e439StUQrp/qNrjuxDVPZr+8jp9YQCD1JP
8islBgp5unUsd6wwRQX+uZ805LXf8f3wzR5taorApwveOI3BawcW4Do/wFUyVrD0
mwt8Y8byFay6c0GyNQvdAL/UjeUHUXmgsklYwlVp82QB6PKNCjAV0jp7g7KmkjvO
qJbQjtafbifjyAlM53PFqyJyl57KecFuLqQZqETPTNjvBfsDLLYdda6VZH6k2/yh
bO77cpgguPTqyJwiwD/ohQ86vP1/EyOA2JdkO+3HYGv9eUGvHe/7L+S2OH80V6Tt
VovW76h82LYDKgYmMGIswXA4B/W+M+7zrrdz68PxTBTzd/TEb8V2yUIPqnQNTgcZ
ZOP1lO3fsRdkmGmWGpfLL1bbBteuAjZ53hF0hO4Bbhligm9yjL94wUY7ofKxvBsq
4LAxYUO8KPG0O/HyECAwleXGgD/D2iox4KGdjogvU/cxC+PivKNoM0iySeKUwawS
KcTG3RKtKmZfkliibZuTA8FY1F05/vKuQnW180XMcRKx2T0KQbqDSFGM062vT86A
QtEhTp9KotIyTL8aUnG+imruzbod30HkN715dG5CHcKxGtlOGVG2bn+2nrjhwcXG
w/n5WFTyLvjcSU4LSzW4tZus4LhrX1yBQbMOOoyl/9l4U+HvIhyKk3ME+sDvZWhF
fcNAilyAnX0IanezXqUDV+nKR4TYUFtsoJ2tD/RuE6vQOo/rh+vMPz6Qg3+WkYUM
Tb8IKRqFA5m2zB20NcOpHh1yJ7oIUzOsBKrPkBmirwZkg2LBbOF634thN6xC79E3
jlvcYtwh3LXvilJ7ob0mQcWoA92pvFALRSxvukYb+4FMdclj5VFUMmtJcM3ioAvr
sJKSqiQ+zFrMtgagQ+uYbEP4CqZF9kEVxgxWyO4mEV3qHFQBPObHUv8BW2ZylDLR
baWG8BHpfEQO05JSRAL+L4VdkN6qbxW6j1Zt3nSun7/ZzN5//n6P6zdENTMPWscU
T/jtASpzKL0wYNmEL55mDXlICWaP4/14BjA5UilsQ614VjzjPJB83iTdvcCqaDCB
3Sd+9ngpfbmgr7unZ3nzs5xILyoski0D7NqoiS7mowe+HUVQw1hClhdtdzoGGYyN
B6NmeQqDhUKUbxg9XV+N4f0mc6VmDzoEqf2ZckfPx7y7GjI6lSLCWMBtvKBDK2X2
Ob716uMHqTLvariK9E3V0xDzDHrbIlqfjTRh4JcTOVvS+t6Q4cY/LlwAebzsm+8G
0rLV8xD8sAFvSU8/3fgvv0c+2fr21reFlWreufzlgfYywpqrC31DWsV9KKmeMTWZ
yAlhvJ53Iu9oZlLkqtBVgLCcvDLmbNxKJ6g4TTYSh66E9V655tOjtF8QlBpo5AAB
IoaYO8nhSG8o7xPXUDJmBk1Dbgs39ozJT7BwEGU5vXE+aPyAliOnhmLAh0xoUjKh
rtNrTsooEesrLT4iBw85ws3elfCSxsp34j/cp7n7fHjp6Tzlay7APxzLKEZkwBea
HijpMKXVTq6866YB4YAi4GvNLxAIhgZm8ECLIArGw9wRoDdLmZd2eBBZ970m1maU
2MLMdVTMefB3jBV3UXmcQ6W2wG0vrTrS6snxmGuvYESD2ze+7famBoCAuhhbC1nr
XNy7ra4oxHaYYNOmMpuipWwASdVZRm5G+s4pPs1KUrx7JSYv3UuayumP1qCpWknV
A2bEnXGh9BK0vWMLCKJHoaK8j/U1RaYG4dMs14H2oD/Os5R31HdTVHqW1Llky/dK
sBwqXkCqVMCJAmfwh/D37WkRLj9QQIl1pIHi0udzSdbLkH6t81b7ex2xbKymXlzM
kAEP+tEloJkOb3qICtYbhvNhbQD3NnX4QVo3BvrPcs0iib5T1pchunWYE6y/Kezg
P7nxIUdK8tnd6akOeDSuAhlenXb5bZWmiG2mY8HAUdOUFwG3FnGnY1MkzYXuSNN0
+pGzNp7KZCxhRLgzK7ac/9yCwae2KjZDrGEj4Dt9FzZ2IIwCgapiOKFGXxuStO23
vioIINWVjiIpuHHCTCZ7/Qq5n6ShI9n5NamW0+wlKAtU9gbx0qCcMzMuTVyb8RCS
YeRLc4autqrqwQikioeN3yVIbfIeLiZ7RV1wTiTCpqG95iZhvQoz73+3kS9BaLjQ
kwfyYYeyam652mZrRYFTz7SYEHE3et5YEr6aPu+qMc+D6Wwl9zvFItkhg6qsnaxV
TVVl41PulmB3SMU+/8whJ+tC63UsWpzGPsIsvlpA9miLBBTokdtid5Az+PVOnWtz
6NpF2aonVxnEaVIpJYLb7Zr/hygZa5A9Oby0QenYsbHbRJKm4JrEVBS5xHWArVJz
95G4TaIzVrve52rZlVlkuBIZweAqXZmY8Uk1QT6fxvU8p/XVSHaoN3hqI0r9fQJp
khfWBC3zx3Rg1/sCle/XJzQy48muQ3MN60jEuRUutM4lVHnSqv7PVpnX6xCEsscf
jJor7ksc5ctS9+sesbPTifXiwvPX0+Qubx1gRR1+j36BNCKOG0Tmbt6gzfU3DTtz
yNdYmjtAeI7WqYoPs3eO8FtQZePWMfz9smH622JcRmROQJATwExSbUsv4QouXutT
qUjiNXQZp5rq7g55m7j3q2XWKbrThwbzJ4VVUwB70SHN0knkHCPCgdWWHrEhsACA
fNSielKcLJJvj9hAoc9MZihws9OS1xOQEY+ha2jD/N0hAkzW6XF5vvuYrhU3z3Gp
UxmkFQZeyVwNlDMlugnOhsdkIa+JI+bZNWVS770qrqsgJvcGzhd6636B9WTs/j4Z
x5TgzPjN+oFQgZAfWngfwFbNnnZgJBwDfBwy4U3PsQIuuEmQtAUVF9vZ65/kj5eZ
o5in1mv4tBDCJrHiz0duGvO8IX64zRL2jrsXCq3TkijpjvOrfS/RtAPAk5fd52TD
3gF2SKtfGBZDLb8ndCtqafOstQofE/4G536R0h78UwNRiUjsQs7oLo3p1CbIX1h+
qGJo0o702e9sDYXwCUId0p8ZobFycsCsF1oF+KUqNv+JDfuFBcjNkQvDnPg9cmiH
6xMk+vsyplXotMLWx8t7Uh7F7K62a7jjBtzPruT2sXWYx0cefN3yVVP5i5iJ10tt
zL1uRbJSYic8SzJ6LD+HYtBKcQEs3QGu3VpJfv943BD3Ej9p9UR9atkQBz1/TCnX
jZKhHQtcQGp+P3Ub/9r5MDD3l1TOgtFDxsmqxxG0dx5p2gDkOwyyODlNeS9CWu2g
WzzOIeVPR+xHszxHTKwcD4F0WTw9rgufqYIjEKYBPY2OGVlL+b2ksyDo1z8RjLd1
y1RlY7djlPIqziDCXTbT9VAizz0r2g3+pIAGLEevAsxbPf7iPDUZo55THgxrpYoZ
TapyaSi8+Locsr9aOQG1TtUYwl/sUKKSVwCeASbCj7dONgKSBoq2qWiTxeol6SzQ
EvV8sdFTdwgfxLHsCFAu4FdcPPdq/crSWiG995f/Q2b6baLg1yDXLBuY52YCfExm
bmIPsJsraS0TUx10NLsXj4nPs4DNsfl+AdI96/RCZEERrFvuRbQFYODGI2/TTnFb
An8MHQVHJgiXertmYYgCLdBOw6ZzRa1NUSz6B2VfHcSEQOgQKQ8aft6gXLivWpxU
wR6cMHVjUdXvw07SRbTx6eJwLUaY8OdIv++r803UFoxZzkDFMhZKBpx1iW0/AS1+
3lqCoGlRyH6u72HYZ3M0Cf/r2kivFVC/r0N4C8jlMBi+jomRAgJoe1+JCdXidV9/
KdobnbBO+drT5pmJnzLpFiQqjMeeMn8HWqZVkAK8UPiTHbf2EeaumWFOVltgDTuO
2TOOhCPM0PtT7wUJsgA05huvWmiu6QPBptUIR8E9BxtAqxAsTYHuvEbafSJxb8BQ
Q/BB1prSDUnJBGVmQNQFQTOD4kliW029rU9b6WdXK/3g+HI4rXY/N2+Se7hLCVrn
591GiR4ObMYcoagkRlGzB66cV0sY7ZXmIAGIGue69dVH0hBXIvQv8fI/aD9TcqjX
XS0/cauQPcUuNIoVxrYdZlyf38pjGZYJdTO5looHAMcZE+eClraapEcce9sPpcU4
w1t4epT6CYMIc5gN5imFLDtgbUKwNvl0ye7xc2cmbWvnmHoocXn6U7eDyI2xh4Oh
q2n+ASDuCa9G8BnjXzf5UKXYXQ1xeRvfJr5+M6oq66JOhwa8yqrsnW3PJWJwZ4no
uQE2Z3sYu1PHO/RPHuiemsGvts+z9AIb5NKVh7q9gtYXcEkjskO8IZTdHz5VVPDx
IzCa7KAzCuZcLzND596V9H13k3PlOemvUY4EVw1EeuIfbh6O4ym80LfREacXrDAO
5JtiDEMqzSCpfo1WCrNbPcsHADRyIcMIEuI3xor43zlLhoODXlPEaLXi11a56f0Q
o1vMkrUIb165kZ1lYn+Cp7OUS+aRj1B/bp2qppfejJwHvpnWac1HiNzl9RUYJLXk
w9Pc22OOA9hcpOMH/Gjt6RqhaOtmgwEYFBtQ/lTzUzeE/maCTG5/vazX3CKLsrDj
6z1lEVY3mU3P8YIGxvovaATBs7TKT/GIAZN8naLknVL6XHa/l7u9aN9MKVwncNv1
fN1s2L0frtxjLtZu3djxLeGCZ1bttUD2om6Rjh4GwDUcDSrjjh/4ZJ4nVWUS8Jma
92pID0IrCPkS5Nrdm0djE9/wd54Hx4qdagPBtsO8fuNQsdILgDqTroaNLgKydo7Z
gXc0oUT8uHSdZcFszgC8/B+KILYeHjfQv9P2Tmh8EYB5uRP769koeS0PUkhhAYOi
IEG60tUlW+CWE4IiwVLG22WJ/N3RJ59DDaYiLqbKSalvMQSyftiUJWbOaq4Yqpfn
n9K1EWxsBTHjbHn+QYlGqff1G8T8k4TAeo4ttSu6l9fo9gcDezVHolUhJkzbnrCU
IOPX++3zX10C+G5HhF/PEuvQCTfxWdJK8n+3Vz1dycXksJEk24zAubU9JoUDhzdS
K69gz5AefEs1pTqR8j+4mX6cS7IgUpjPjVaUviYvt+MR0q6pLUaAZqtYVFkzAMFy
d4JMdHVxPfgqAElY5ChrjGvCSZ5tyXDR57p0iHYd2PIKUZu6ooGJo++yyX4zuyZW
rsXO80GZWuEuFpacDtvi/rGdcz6ly8itHzdnLjtDHTfxlI6vDY1cVEghebOkCv4p
3lEpUuINfMjPFSoLSLWI+UN011n4g4cy+liwKCCiQwDdXrVYT97963YERA7MTV5D
W6uU3AP9mNuLNvEMe/pnYlARPcDuth3zzplxxjVn72bH95W0Iv3Ys+1zbfk/ulUO
cjnDeGnTT1jeNuG/Ml7Mfj6ZuYOdSdaoJDFvM64n4llH79j9rFXC7Sqjd+HNpczf
1qqBxzbf5dS32Ltnrsw+n3rbARs4pKRjeqQTFDevlD/B+kHXK9EOYdegBhaR5XDl
o8oVf7YwvQD4Kepsl9wJR20+SvBnOQqmWYmohXlqjPmOGRMexjqWadQIsLiu2tVF
FRtKWopO3VYcxpLZiOaZt5y6BLFLGO+OUBQEK6g9kEjA+0sFmgh40apKC4Ez4sMW
M95acWfrN/nyenLXmekkuL3zyBfTqs3Deh1KSEEhUllALydnXrB4UBgfv13xtcqc
vmLJVqhTX7Al4MggaH17om21CTJBgQiwJdXDCPEjpTApZ9qnOgIZuWLA/bteJDG8
f2M8hwjpSvvl16SPLs2Nrerl0cxIEVIRLHqbJmnNZ6okaStSaO3X6iVhUcaf931i
zZ3Rm3XnkbWqeavLwgWIQZxd1HaELP4Lony3QEC72jzHejbcv4ZvNZW1nWJPCOGu
g2fffRo9O99y+AoQrH+GAyCkT9TnYqn3ssfDtNCcQPBdrGH+bEND4BKBWqzTlQGQ
tHN0oRZsEdpGnvh65ebG/4aeo9C0bIKOmYe80sxw5tPZBa8v0Q5uJPhobHW3LK92
M+N4+T4qiagnPLrK2bHgx0pVKK+tRGHX+4vzJvMfsXH7BuTCvMT0wWleBJjpZVW9
IaCR/7p2P6/gru3K+w0ImvPGXq0xEDk7aOzZyyx6JgMJW1FNgcB1BPBtqJPNT9bk
4BZVY2ZB0ftaOZ2IFbfco9+6PNcM6cz7ru8+NR501VElc1d+d2OuUB68NE1lJoPC
lvlixYySA4R2sbKYnzHdgnW0iReCQA4gPylZhCtLbU+ULcEzKrzOmKI3/jn4vDiN
K6voUuIigaykhotQaa5346YufrVPdg47+oX/pwdrordqFK4FypVs9Lr01OiOVWQ3
DkZxFrp+dfQSsVQKL/5W/srZlq4xT0+432Fbw0lSvdrFqJe0NQZ0zYq5JxbOV5eo
HmvB0SlVTCBhN4MqFusWQVGDqALrDA7OSUeq38WISR9mxFFzSKGRVqBtBJrT8Xnu
UQ1H7DsrNY3Ph19eBgA+ZukrKb71zepaVYMeH7ST3MDaU5dyc58I5L5oMXHQOVNt
eri5pF/WocY4GoPPdmIKShQSZ50RHEaMrt4q5UZD/6XSCDBv3dqcegXv+EI+DbxE
njeFHH6YOCq1t5t581mPDqGXJXEo2E1/Wtipu/sOqR+viTOhXQOAvNzoiWZNe2K6
sDaniAoh9cmJreJtXoYnApKMEpuezPk23vrVir6sFQHIvowsn1AIcxYtxbcpAcxI
PqSZKvw2bKGgxwqx8LXDtIWlsxEW7PVLMTyJvvdcf4rInT4wtaFLqUunabU/cJEw
nnvhyFyENRElG+hhi38nqogM92yc/tmlbrRddhhHnjeSBNYBGqZ1Jg98n4AomGsx
A9n0CXc2isRTtK2SBJNyquoFn916rso3Xq7Gse19uyhG2Ap+I2gwL4gm8Few0iy4
XT5IcQfjv+f8QQe93uw4hKSp+TT7T1o6d6g1nldaFTk/BKG7dls3c2wcSYa37wyn
ENfPPxyyaha3bkfPJZzNUr0mEoMcCLExahyxSCQ4faOAhOnQ2ssLu9FseGYenrx+
hKNfBVOz2jLV8QmZx2Fywd53tYgniPQh0emvj3ZmaV8/2b6JgETzT3A1oLtlZyuJ
yw584nfbFK9PSjRI72ioWx+QkWedO15j/slL23JIyD5DUeO2dEi1vIHCEi9sstqs
PzwHgs0cSETC9dgSx9KrakzGxPSqLvmKARUWiv7tWYph5PA2/9kXxLjXs/IAHo6U
23glv0jGOnlQh0sMexpGBA250TR8y1c2nktKeQXlPw4pn5iCw8xodZCuJ5DeIY05
I9UktfFzNBE+VnQQXkCuPFGe1z4kzba4xou3/JeXqw/caY+AkYq7DFR1GlEwTBXS
pHNoxduhaaOZ2t6+mvog1IOyxViZBeWDXiZcINL8SgpAyZz13F/T53f5zvj3v0bw
cEoQo4ynYddOMfQr+e0LFN0ATwBBERnRgklBR4EKjV9k0hoTV0r3tliGr6S/SXvW
AYd9//8KLdpCvDeqrgMhRCDeIB+gGPLr5+UvtGk5bZ4pwx33zax37Rb/80ckI2fh
FsXf+Y89hE8PqlAKhJbmiFYF+qsTCsSYtMMM+TCq6BA0IvcRzd7DN/TMog6WHqd6
GCiqI+c9ZDeYfrxbGj6CeefaLujV9vzuGWz/J1DqrA/2hiIfntA/wNAG5DsW0u/J
lVDZ5wcpxpFnJ9WtXC8BJ562FOQmCqTNMIhSfz6fpfN6JQdJC3hcfrWuhokFWOz1
XTCJMwO7HcaJ/zHxhsoQ3IeufmLXd7ISlnvmKI8YrtvaOcYJQHaVPAFfLF9A5i9C
JTNB/m1SvD8TCX3nkeKHPbDcthxQmOIRyk+u2HoheRkTQEKqcswzCJdQ3s7hOXGo
axOSGYAG8pmHHtRywbwwfSfMQglYoGHSpoyexzNJxcUmorORHjw4AEd7oNM6dVFe
CHRjimyQpAVBWYduh9IzWHT63f+KWjfF+lOfKxIYeihQQ7aYLsFoF9fmhI5CIMXd
319wsxMvxMn/KqCU+oknaAhCQgHCfBCbQwKuz9LXyqVComAxDBuPf6l0URGutb1O
9bzNzQZVABraYJ3VJvUACwLqT912mWlUemoQ0YB7wBnYKPQ+adoAu50E1Dsc7NeQ
zCPrYNp+JbFrcHz6EsEMrvnTPV20yuNHoziXyZjuI7MMoSmm3fEg9XA1bxiTSFmM
2wx53zOGQM+M8hPAvYksRLrtgofq0MeGh7X29fVBE4UD6SGcFKGAGhSbYERK6Ipu
tlXEWPUel0dLP9xPRA7wy93KAMI5meQc+dR2khxa2q70UJfYAfbsQ4MSRJAFoW4P
YoSNp+0fQtyKByJkCgwwhTMQD+jQSOKBnR+RXX5zAM/YidgDPsWtY6GZ8Q3IitP4
q+0PKBL9CsYTcnvbpalMQOURdIu6Bf4B4TzVOcVUsMPfbVs+vaoEQl6PmDLcpMwt
p82wRGu3vWr8xFobk/6lExNQr0u+xX8IzhBUlwOjPQLNtfIWWu/KtgWIEQMjjRLD
ST0zaFv6bJ7kEMOz0NLRBm0VtyqpLCT6GOlW6jko0AglKdfNOYdF3iu0dfyGfM8B
jzlhg9xN4mgksTMJL+6QTI7fDmeUtXUTR8C2CsUArmgZCZCEy00urKZSR4o84RUQ
eDBz8sbgwNs5UQsE1UJw7HUlqPPMUAQ1feT6fg6maP8sh1kgc2tKd2SErOtuxSpk
y5IU03vLRQDQ3jZCYkfdMvnUYSoNQ5ZKGUfB80dwSLeoOQ/pBVNd7G0su0nBxNzS
Q+GJfoVhldPRhJ8xf1EbqxAIt1yd4Z7MTBquIoAknxftfjBsTWDofTczarLRlH+X
owDMIZr2HtR42NzuJRjUcbl0QWIWq/+rNTMVgYT/y8/aahOJwFIlVQ/Qc1N8gAeX
h+lZMuiQFdHFaND+FYuLBFzolEPLnZrzFd1h7278nFaFFPzLeeiAJevqmdhQXCum
xVgrVOlP5Mkpily0pqqIqQXtzIm8pweJTIxzT2Bf4o1fZJo083gb6Rf6CKuJG/3d
HwT5p6I2iCVPqbbdaFzTcZG58C/HXrecaIG4V4pr+xobGN72Gg499j0lqIZ10qB9
p/BcptItl+VgwlxrHcaWjtfvBA0yiRt+rUQYqxgrxsA++7FMKWZBHNelyHLuC/mg
iYJeq9Q86KcUFA0ENmvBuUII6wMNk5drhWGlg1XZako+wKcpxEtzvgb5X31SbIie
d032ed0GR/JsKsqzY2uTCkgjOHNImt2Hq3PC9/Kn0ChAINmD9gqFeCuwloDvUxoK
jNPTkMoTC28Le8FhgrE+nZsmjoKW8Da+T1YTasFhPi4zXGTiZvi7hL8jUVsPGwgz
WDPQztPfJwITt9SOHAWbLmUyMAGc0d1C/1S55IWP/8FfQG+297sDafitjt5RBYMD
73Us77hUo58fIsZMrkbOii/rFi68MpAAPEvfRfh9Wlir3NvIQAuxWuaMQholV8jx
QRPJTrwX6/w/eva7HH8OZA45HlA24D4v3J8vp3WC18YNQ3oCAT8Bx1Ko0l9q7jU1
LLSxSfX7ogVZUDO1Db3XPahx0MflKLt6EVP/hjjVLtKr+0m9ZJU6LNof+qddRuep
zTGxq2gB+bK/p2Y+u+nFsdubeWliOvU97kQfpqkDHsa+3SD6F+uBmuNpkK5IozQL
JGncpS/I8JvOt0FyGoy4Mvxwpz6G5kOBo45v+fpme2sbnb4Ad2EJoZHbxXBVbJTu
BETgawkgTWnJvq3LgWumTb3EnpxcHGrT7IDaJW/jTFk/xZrL8BlCgCsJnmS3ntU0
1Qwlb6LNUp6IINpMdHzlQMFJ8I9pRqTH+YeRyk6kvUID7lxSo76CjD5ieivvZNeK
cLJgFwrxoyOf5pv33WWAD0ZusfGwZviYTztkf009Xrme6zDqlOz9A02dTBqtQOkk
sFjReuis2I9CfES/4h1lpQLFcBjYox5bj5CKAqBtQ8Ot26cvHPWAsQQE4CxTkkwn
rEQ42fMYHWRmfL/rFHcmAigjo6Ml3sWz7o2lV5iDqF5zNArbjprJf2KshyZSQbGX
BMxf+7NxX2kbD+Zu/SkAuFaTXpjPWqJticrzow7y6LKA1amPNHkzJeO74bqa5UQb
IvFSOpm+3InK9tFgjbcJBOFO/U1Bb0r23CpAIWqfb8aLWvrAI6VC46INjw9AlZSI
S6ExJ4+Qr2TTSaSBSDO1GfvluTFUlBsblcyzPFpv/mus5Lh0lnLwHGIt2soq4KQM
Now3lHkUEDoFQ9Y0COnOyXRoVyqkp41QvnY4/0nc5XU/iJo3dFrm39rAfwZPQkJA
aHhjoJ1HSOYgcm5orF6D0dWxRGwHefarSc4hZhDAa2JyZvEZJ294gazJmtkULVVd
yTtE7iuccxWxFNWl2YmzwJVRAXWLvHtgI3MdtcwQVqwpM7/4FOB0qbiCpr5ef80F
ioqNKCRZGIKynDvNXS2ZOa1a/FAdUMD95uQCAQN5QEcgJCB03xqY2E1p2rsCck2K
+UfFAD4pFJe2cV/r6jlcThPIZaRsjs6Dhf0sgk1OlLOnjLh+GayGoZMlLjWbY/rw
MDfb7muoxQGxVbKY8SMyPsvdXLNf1FBqnE2q/zqLQDFeLhw5fhCmIwDGulhH1GAy
l9ydqED73oEOBhy2fo8ukqhbOtUsHjeftLOZu0GvAKGckWA1zXn8uYpkTyjiC/3e
VFBwMBJqsnBuHJY3QPy12L0mfGpWPIUhEi/CiTOpomjSJT6c8Bn0S1/xhL1XxTO9
Eq4JvsRckeq2HvEhJNO8u41iPgC03Q15ZXdK4wgC1RNk6DLSEILsX1MBkvBca9nm
4/zKrpNyqZsWdrIdlbo5cFuspEK0WVGr4Lb5/c7PPtpSmbtAf6Thr5+wYy2dsItp
ndffPWoX5ogYSiJttEPoErdpP8cqEAyhfGvkRzDANXJ1KfFrxEhuBKONJQOJOfl2
3EN0WxqYFqlCzsKnR3/3YdpqOm6otFttwGg3X1J1Swx4hGoQOoO8pUdFuqrBMT+u
lGyCLtUDHsQ+D2yHb+IzVv3lr7VvMHF6dk1nIaQTU4dYcKgSKYCgGQ/d/2DFb7/G
m9Pi44z74R22Wyml44aQ8OqLCdEBfel3ryb6jnYbs3mZXMPaDGvdua9DHwRIar3+
3fRcwlHpL97t3Pw8YHY8bAullcxERlOq0rdzR76n/oqcss3Y1ed9NOuvMlPgKrUg
x+QOn4sdBXG9xCiUVFfxdrX/LyeWtL629udifoy+CHWEUVuB9nIm/IP8i7fJXmkz
rkAiHfGNQvu0bSx4VQq1SXoa2H3vDfK49QrcJuRIQ22UmLrI9d4iq+f/F+LaHQM7
Pgqb4Ltaz3SbcibXNSsJ96/Q0YmwRvhHigRcVtCHi18R7CJ93JAPn4o2+armjSIk
R91Z2l6P5LEPu1WhXCvSFkByAGNlcxHZIz8YKLP46V4VBkbtysLr8iZ+K667wcyc
GVJZO8ie/f8cQCG6eh4gilm3r6a4Ha4wxpnx8q9aN+7BIvUpgPXS01X6zAx6bX6M
OV+HTVbAPjleaY5vHOuGcwktSvRf5Dwjs2gNmPfslWKDdPDcQba4kNuNF/3SusEZ
Uv8oQlBLZtvDcSGLQWAfGDZq+J44ghBSzbFvzycOnKenKXw9vXofY5kw/zsvFgST
SKyz/5NaDjkZAw2TEG0nqIowoFcCZciP9VxhRwbRj6CANLJywxThsHIbpOig2woE
cjIxb3uZ7R9jL73I+NxtTpnWAwCs/2XetbMZ2ouzFSeC1TMMoRp+ExTy+DRWEvFB
cuv53mAsNaLlnWvgbCFZpIzNU4dkSz2WUyu+fT1MgU6KuyoU4JUXKMFmocJhRnEI
smHRclqlv8L+ObjaBMrpmeIKwz4BupMZHki5N/UF8P2eDOB3eJCUs72lsaQ5tXM3
PvgM7iig08RAv8gCxAft8H8zuTUnRqMzYOtQJVEniaD6fEogfIIHr5n0WqT6o5qK
gXO7Sj1YqlE5x0rOEfGGTQ9hUupb2VG8F/MrPXB7B1x/I3f8hNzz0mfs0idV+9n2
jrswUSmKpvqwWt9hsvMTye8alae69isQyVER+JcdTWgdIcvtTHXGnBD4xEy3ozXx
LGFL/Ek3n1a2YZYFkxfQRbYVriwraggDjD3861iX3fVeWpxy1pMrCSklJjr+EAKY
791/vJQLXvnhLE/mLMMRSOXjdy20n2jZB/V8EniJyTxmx8JQ3AQ0G0JaglFLHZy8
g4W9Zb9TblP7YLT1z0Ut58m+tjtlLqXQmWCDlCiK8BHx699UESkUliZEOHpuuvSl
jMgXfQnae7T96CAZyoD7r5bNilz22Ey40G0ouOdJ9dhs72RiKGRO9Zz5ortesl/a
TTXbyHoU1SGvLwjMHKkOAuRndLCsgwfUnhIj2bTHI82ldxWDUyYJy1xWDvTdyver
lt+nqcs/wJ9JIUfCs0ulKLJG1qSYOLfHfSEM3kde+T13cZ6XA/pgbkPp557LfPq+
JMdINd/74+s+ehvju/yDgMQnRelDGaFiRUewghPumcCdKUNz3/qQr/HClQ6rKxw2
QUsR3Uk5Hd4qHDGqvQURlqYl89qVYXencahTsnzA/BxJmiz4KN2Y73W8EDqEdec9
qCE7AztJxg5GXCVMe30AfezhgrtLgon72Bo8PbfM4uNjqwMN9iIbil3TFyFmLE7K
x99mg/ACJw3sy7u+PRLA3BggSQFDhErqr6Hp/Xv4wBvU0LA7wibw0W7KBRvP6Bt8
ktrHFlqmhGj/3h9EFBbSlsN2iJQQPkcY8gr8J+TJpUqiNxmP1oDF+TfH0G1Z2Ckg
YL6m/tj/eBBhVBHJSxW6xyElMy53Fg79c7oyRK2Aad+OSe6Ztn2G71FZvDeqGOs1
eRMqrPXNaSqmhbDfnEgF2gX7hAPMRr/ArUl6x6nyQ0vVKfSPzQbtKIl1hS0IQ26I
yMnjneIZ7Y/G2bWUSwf6/RcnedgP+aUPDscus60FPS+Jtw6eYNd4vA4gAKQMHa0L
oC8QziDCQu3y+DqaLrKJoW/85LsZyuQHkNXUuFr/+UP08wFH5HzqucKUGiK6790o
eTCzqhCx7xiK2ubAJBGt+78Cgn4tHbjfRmx9UNM7gaP6MGv4xHhQKC6HZZOnO+kR
8WT38llMiH3CpCWzhsaWujEAxCmkG9Tfpjbf7t88bsSK+A6zTL8DppsTq5gyFY5x
0mly+G6ytkllXjCz0LurKA17aNbFwVPhUGUZYH0Cnqf31gEQWBqn05bCdWQxhwpb
0S46XoT1paDfIgo52dfbRK5nr+aVxOCU9Zfb0+TACvquxg+3rzmrv7fJ4atkBlN7
PwtrbU6UH2KKRx8VURfGcemM/IeAlWQ0VUJ+S1t0g4mzoGa+75rO8VmuoMJ9spI4
Sa8TQ86HUrNDh4ejYmtInwAyg2QZI/2BNx6+d5LId5TomR+bbhnLiGc2aimk9mFr
26efyqdpz8PftpUdX2v4nl8q9wwwuEE/+RMgpkHZhcVgCqX4Ok3xSkJeSVUvNDj2
WlaBYAP0JKjAZVzflWzUzX5k8GMeGxLjs0oWw7d1eVBhOJPtCjFMFXFg39SR5NL1
j8LVUgev3pTl2ewheNlc9tteBYJFNsFKaZKyESZ+dNdW9wFC1i84vBP1UuW6QJX2
tgscBcIvmy2EldFPfa8W/2gTPnHUYQ55Yt/mkRpOYqKMtwfJbc1ELEq36BnIQeEx
OGJbAA2eGL10iDCpBO8TKKH5oJ0Xtfxp+BWmml+D+lb+F1sl0Lz/kTszjAIRX+CB
KkpVMOydPLt7qpdINlAfntQK178GuGsrVpeB6+S61DFNyl0pjThRD8Uf1vLFP4EU
RpZYS/78cgn7BKz7ascJVnHrlNnVC7q2ldpl2DkuJansIHpOc7RnmI5c9SCwuxpx
Rz+6hEL6hqz466OGkCUdQg9HlEyyY3TJCUGp36gd3icmWW8iCVz0DzS7VeVpTbl7
hVYIWk9tqwHqP3fvB1S9b/KTLwlkhrbZw3LTj7muXzgote7kJfYdzfH0mIo5db2v
Oyic9UthkhWlvmXq0IPH4WWqPQ/9H2dejfF4/qWxLayspoCxAV3zP+pPdF01X37W
koe0WPb1jwLkV9ZTYRgV2sGzR1Tu2AZ+D2+t0A+pguCtxp3jhaLkpWJkEmLd2gUy
q5JaiFComaASkCF5AiviDQIKdn7iTLnyRvKV8ml42fk8JQekSTHnb+Q6JHHExwCd
5dYrS3GnQOR8b+mG9K/WaKV5CWKzqDYTpdwXoL5zx93KSMr1NgbmRMDK1fOxyuPr
B1sV96MpjmO6Vjy3n614qJKg4EZ/tHTtcfowvmLK8bOPqIXqAQage22GDyg8HGKV
TF+FY+DAVlcEvD9pT0BrSTTSOnWg6ahFn0OIMLSEruaE2dRyrUdiSlC5bY0uuvCq
+50Fdh9cVhYJGNFG6Ut6GQW/NPEUTEEITMuet16FgYfqhe3zQ7FKk2/4yJdVhKtE
57hcYX97eAv2tAJio9UBSXMYbYoWm7XLCFeuwwztPgx+Jq/99vcXRb6OsecESxAC
gTCb9k2//LwKV3iDCeJ0TRsV1pMV8hGMxc/ADLu94HoxkFt9tnsFqsPBFt6XPKsX
rRqqBywflWRMHMWzWVAq902MSy4iV9p9ojcnmWB21dPVdFhcIVR38g9XH/MVK26G
b2h0Ev2XTiNTUk9HHjLdgL5kQ+MoLAH3oWkejpgzd/DuEchLmvEjzhQai+QgTn9I
kfGQZx7JEhy4tGb+8dhsIEkAaGroEzjOsYeqw+mhpemdPpTjhMUaBPHlA13fjsPC
41QzqXWgNvRNYcECVnLTDr8xSbPG7yX95V3tjK5WvkeIpXj5n2baWbXj31ieHL1g
snQfvGpFyv3urf3/p9+FrxOw+FiwILvXdxjCYxsGg0Or6JlnyBpMr5qFJv7ySmhe
6e9mF3lqvIqDQTZEvrSblIPQ8wmnb8X4iL4rCi9WL9pDXATjFmDFFLnHcnhZCJ50
wqrq7qXRYFONrHeJas05Qtz2J6EQV1BOwEPoxmd+7cLxAxP8QErOjP9Y+WmnAIBW
biUJpeN7ipMSBJUaUZyGGtsG3p23R8mYEDlo01JBwi6GwJgwS0JoXuxspA8b3GHx
s5gGFiJnvfEc/RItDwCxwMdh81FzdksbeSoq0WdvS/JU3Tn1LIv47MMSb7+9R4f4
ueJ/EydXhU5jzjDXVX1RW4bGqvsIag7ICtwBbp/iayK5lqv/u961bAyh2YewR1WR
Kj1AgQAdeG/ub7WWfizkMzzim15Uf/f9FdWZfcqeb2P98ZPlMZ5Lkw5QioQEEDUE
2utRQlxMRtrIb6077l/Rd76SnZMfQcml9Kh75yTV3p8CmfnDnv4vWkvv4zY3Q7gr
Fyv7sc4wMUlR0lsEQYf4N6rFQp6R6RU+SU9On5lm1iaVeD45zKQzbrRELiEKw94i
t+DrqdexKk/+TVFLcVMoKddR79zckCJ17qtU6MlEbmClBf+PDhJcZf1oMWvVkA08
qaxIlNwxZkgfEVBCZQwxDs/g70OsAVe0npQdDGb1ds8G3neev/CBroPBniqKKUaQ
gx76tMLmjeWd66Old/PuTM2x5g/NYtx21LVB20ee9CKY0yW18/dDjzGDolv7QBhp
/psswEcOLBpPsWA/2URznM1PR85O79VfVVe9jmQuKg/htEi8VZf8Zew1AIaG2PO4
1DNXNaMzhydHmyHa/u9fPNiB/yqUs1YdMcNZFiq7BboWNDceHL7J7vDvrg29WAPY
wImtsAaHtZuWczPHIECU/eih6YZI3vmjdaJkotpJG837saSQWDtdRfmvNPhojhEq
xmNGfTj9Ssk7PgUeCjgz1qr5IUCVjki8g5Psaz3MgLxvYZQTAkCPtEvs1DbOPBOP
TyyJRcU8r4S4q3COK8apYQgIAE0xmP5svLQ8eouyddtEWew6XVqlqPTsm+YqMwfH
PcY47NqQW33oWmDxCZ002S8Ne8mxw5BIsCE3PAJA+Nlkkj5W2fChDO0N2+q3wFfd
Qa8C6D9eZBPT3/WevzOlhZ/KF6Th95es/yCAhmiwDYFgG88LWZkJnX5BheiBx8NS
1hLbPUCrHDvwVHQPgnMbICiodJ4YXj/c1cEhc9LxBh6gotVDfvdZHkH3TqevPeDE
1VBcyExvTC/68XAHerVSdoGwFaxONqhjxlXs+wa704YMLQLqTryr4srHjCC/exEz
8Jt8U+Wq2izWCzhuTCuCJhojk7OATvHAT9CY3d1yCixcdPi+9OXjt7D9H1SGYHbj
EbbfuqbPdZOFIlfp0Xp0x6suKmPYfT3EAZCOudpiv5AtQ5L3br8uIP5QWtcAw6v1
hyVEoEsfhVsrWF94TsDF72SIw+tHuxAXwOq5Ky+j7Na1nsj6HJ7V31GOeRAL1gNH
yJox3KImAnPCU33c9tfUDb943MVPqbhKss/m5oGCntUNZrISO+hs5C4lKGrXoRn+
FGVBhXQ+oPXeFMkuPb5UjwynVViwn8rwBifCPz3/Vi3lzGgXWa8VJrBaHiR6i9fk
sG6VbpXsjkQHSr5wLfG2yFaWwyjFNJQ/PVWs5SqVCdvmaH9vjWYYfyyR4zmRxRaR
uKBo1JJyIrvVhMXQA4ZGSGehN3zn8nDPcb9YbpJ0g8FeQ6OAgv5BexlUPxgqeFVF
EL874HX1dRWzQD4vWXfVR6WB8i7vJkiLolunoc9r6kG/2SRY+xGcR2xdLmDICVz6
kKMFdoXFCsWmMNx4I3Ma/k4x6/Q41wNJbDEzSHBtfphaVd9xy9YNGBX2SojOp+MO
dClBYhtjuENb5QEL+JUsvrdiqHHRGsEnfitYWPxSjU+/MEealOKcKAwFoXrhnsrH
puMWf98zFD5CQhyGbWJKNkxLewWsASlSw9LBC7riogL8uNsG/Gn3nPhd9N/1atNK
nop8rP+3ThXOVxS6Qg2/R/1eA/AZRfrslQc7HVa7Wj3HgmFyleO9nZnQwRUkNagU
EgtUHmI5dCzZJVXCahVXp4LJjPa3dPeWftysl9NrjhStupowZ+ku8cDC8K1UPmvI
ZdLCesypIqmDdXgJiMbeHl4KXSum1xZyv9dFN3tNCxNEeiUJBpiEi6w0UHofWdy2
NYUTkeHdqabeJnE4DYQ3+vHTZMo6dwzJd8M5KVQRjk/cxO5a4NaIA1ztIu5ZEt+Z
wzZNzFifyeD+og4uTV1ZliIMIMzu58d0dae4UXz5AnhZZkMFhFJfaHoeqjmRCSYr
dPY+G0IFDp9NNRJb0E8sIgE6CyDArO4rt6S/D1D9vayoFvELD66jjZlZxQN+Hx5r
y4V+Q/lGM/AVzgXmD0n5V9qf+lpNaqEO/SWEiRXingZe85KtpQYYcVUKJUPdANkq
DXoVem0S+8FXYoAxtUoMATjwXOoYhKOpq5tSumLZnqJ+5b2cTZ8tzi6q+Hvhio1A
Df7kTUNwneTxYqXwnNiglYewL6qTdUi1T+5xAZITrKL5ezW6jheQJ0DV9I1nvnlr
v/OkQL57urADj9k2mst0pHx8VAYBDLQbm0jzKUY7aZ+VyZplpcfBUeXklUriN2n8
GIWjMSQX+USQDqpQDYR0UqB8giI5pAUCryTVrIKHRqod7gcjJZG+EjwglEZbEn+7
WXLsps3SwgUbxIQLIjg9WGIws8jkvO35z1vgqRslUIYtFDfFeQLcgS/w/7y3IQUm
ckVHg6qey/uYDvr+ryDt31xhOFiv6DIIhwZbXleDaMCyOzyx/ExkxDX5WPQ8I44L
YFSOsMZ+s4EmqFqOMvGVPG4z0juzdKzptdrdoBLk7ZhbQqldIHnm3OxJyxeB6/qs
yaxGjiKVCYCj3QGEBeCMrsgU0LVpDZMF/nTC34nySMt5VAtaTEw27okJVnlumQo6
CRkuUQvVwE/eJjjoLOXyadKcX9eF1MDiuefpBkgkBUA2ZKdJmzYu1rJUs0RS5Lc1
OdPwoV7ziOzdGOQ4SuEwPQyrNBUDXEj7cBlPvazaKg+8iUk7pN70Pb1x3hRRcPzX
//RsH/ThVWbiGMWWmT37MEQKr9TFE7b1/Xo0wieTh3s8b4LlNTJgcBGqd0lTw180
aKcoxpaB+Vxx7OvxN2Xq6Y2Ui1FyzTz5wAtMue618G7vTe49rNJJmC9dZpu8ma72
4XDIZQYXlIUMs8mEtJOaR0XtQAWKupC5FOlCMDUjwcfBktpIXdY5oXCnfe3mTyU5
fDf3VOCJ+qOkBa/AJIeAXlNZ34jHaUAG7OPMBOloqdcS7AcCim8LTZUiihQrU9sc
L768nESHqDucuEqTT5Y4a/s29K0IEvWcNhGbofGGmL72aeCMSOhqxGZ2KtYSNG/R
G2viMFfdb/lWchmREvEPrMrKmyek5S1IGXclpQRFXq0G3ULlbMEL7bnQR7yLiu3r
GVnHOOQPt+0ly/AnU0sae9XOttuorE/nKuGHOxrZrJNA2Yt41iAQhP7bt8t33qJz
IKePjCDvGEEqGWx3PTFEJeqH2PvxBmWxtuMv6dTO6tW/QdCJ+HokcTsLY5M7WpY6
Fro7BixfdHOPa+LKv1gLRjhkc7E5ZDRWwFTTfsATuZgpdgA5USMIm3uk00Gk2EBK
yiiWercu16hjLd10lX9oJ0OyY/pLa8V5gQzPrUVkKqdAA6o75H2eO6jo4IpJr4q3
ToN1krC4sI6tT+DGeI578aLPkd6+wjQIZEcF7xKSWqBlmHZaqf1txHUWA96SEYaz
S+xhZO0pVeFhMhb8s5kulfmC6dzo7v2sGCozySB4rzb9ljWkn67Z/29U081mhCKo
oKFuW3lRjLHofYytOr5U8qsaQxf5d34Tn1FDYb+C2nbo/cllje6JoxsGmsc5+Fvk
S5rYp7p0dwGeR7BAvWYqC5siYK/cU7mMXO2VNo7GZBdJ3Xxu90JpKboLsVUmTutt
d9vwq+T6j8ykEs2/dANbYFcnmpt/o0yEB4dqCuRLgKOL8hIb2Cb3IxmQDtIcXGBq
AiNDNc6QolLk05ddT75xX+tCsgGqzTVB8UvwxB+EOI4vXUtjBFU5IoEyzPrhxmMK
C3XiQwHpmqVQaQ64aynWmj57QuVoj3MSgunohkty9SCLGYhBpl65wI/fkZumRrM1
kftdvZ7LE+0z143Tdbyx3i4rZpFUrar7jXu2/sEn1ma5gh4Xk8xQXJzxkbmGG50v
MHMQ61rbmQ2eC7T9L5epQlAkE72BG2J8itSJHS5fyEgrk4Omx0nHlBjbbtYmpy/Y
soDNkMs/83wmZRyClUNeEd7H0LgiGkj+X50JJ8TRolSyuJfukaCmZiXMr5a/UVkh
lanV3jHcQWZBCUFIfEqUE2Kfo3cDyRGiBtsYpzk/0f43rji9p1rUSJuq4oKrAdRo
DvN0vT3El9yORvRNDLHkRtGyYLfw45xTsc/J2uj/rje9Aat7DG0dKxhf9OqkbgFo
+LdGW2CbasNRkez9wkVimbCKWTaBd4OcZmYDkkujpMksrD4cQCwu2C/vekac4xLR
NVYW6wdxM+GVYLJBbVHbXtRYLVQ4Jbx3x6O7wVY71UfHs8RnzRrrhK/Q57JNVhzB
qL3AebOIJfp9r7XRHDmoDttdIMclAqICp7JDfqNdEY/Cfcvs7A5/K4YYY+Ej5x+J
XlQOnv1vX1K71ENgM4y2KohIt+fh/PctgsnRpoTQ1MEtsuApJc62TeYshwVXZvLa
TUTvcZ8kQMxzwhOJESMZsp55n52Da+UPcvuR/KVohQpNwUkPcc8u7RcgEIn+gvGd
sAR7dkRD0Anh+RrR/Esok8XibPwarT7RA9h302RzYj0lpmPTLx3XqSnUaEPiHF9H
xGUegzwTuNGSsrT2SFsESHsKcp/8Dc+YXIEdKZ4Qkp5Gzvkjxkj7fDAEwNoIT5jc
QpRbTVLqMj9POkbtFfNt91DktFP3IE4tVhAc7FfqrwR5p/Ym8wFvCP0lrGPQv//N
wd3HCPLYy3T6T1erG0YLrDt7nYEEdSIm4j+GjcqA2MTECM3/H8Enun13fTAYwQpv
K+IR7zf0qfJg3Z52im34Me/+updn7wH1LwHg7Q+xC4lvwVnz7D2ZHkmO+6pRrgkj
//K/OuKI/NQrcuFiZZQmsgoFHKerIlnEkoK6WyjQapfoa44Kse1eWuT/dUw2OGvm
2zw+6zMeemFN4bhA4NzDOSqFbmta5bMQft34/JOiduvAzJMIOyxuKFoinKPpaftu
rDQFKgNU3sM9Ume6Ox+I2HowElzhuwrgLQahaw02h+NbSw8jmoUypMoacIkL8cEU
mk0F58bj9fUL2sE3yaCQBuCOmZPQ1+Ce0p6j1mc0U4pv5Lc/uncyCQ+/vjm0G/u2
xeUfxlHlmpo8W6892bglba0wra8ju8wdlTzDxD9phXj/jbUh0V+8XEtwQ/GULxg3
9AsrbTljHN0JsvWi54rE9NmwyAUQjdCsMqsgTWRFfICo36qJUOdr2tSTXOtIKvQK
qLlS7lex+U38bpW0CmcutDoCUpYJTSxZaKN1pU4OecHZaFJP3TXyqgDJkwoYTn7J
Wm+yrkam6sn23i3Wos2a9B83XZ2rRmpHogUWWluHLM4TmXUJcfQjrcT/j/Lxumyd
6LVCmXVQ2I7gXbkXuUgPIF5SmRkySLYeRftPMHpCu7n524u7IoKsKOjy47vUn/lU
h7FfKhATW4AHQlRrhtLEfKh+gSykkNwdt6I8uzZ3wI5eNeuqbqvFI7MEBfzu2NI+
PYpT2wkvqLN6LqJ+shmRuyB/kCBRCw+hZyTGYFLHJN5O+AGKOoR7jIpcj7Mw8/hN
aGfQ6jNF+v8xgAH4NO48Rac7ijojyrNe6CF/l2MknoGJMBrP33uso+ON67R32Vsa
v+nax7bXT2wRHm/GxKWilNAwGw1bfY3SlwRVhlEQCoobwHIYtdpdNnaxow7vst3k
01G3cpl0EUp+phaqdYxXOM2ID+cP8NFcG/3zrV/nXqQck49Mw+C54dy+9exsMj4S
k9XOjKVm8ldUKK1oe2Oya9ddzMQvRyGSeCKD2oyxyBlkkG9SRapzhG+MgRrpu/QY
BWmQq5KJs2GAC/FoQ3Od0FNmv0iGLeZCzl4dU/08b7F1hR5d3DUlh9DPgch60jNP
9Ai8SPwGC8NQFGnJU1dFmtwpMkpDwRe82lI8VzytOaTsQqw31Rcb9iWLM/qc0GVi
hxwgB+fVj6aOat30zXSzXM+LSgy1ikG19wHCu6HO9NZVIgFXESfe8LBYdJXROXGT
eCZuAMA1CSxIWmLBE0Tq44Rhd7iL7KgBq2HcQTvli2BwR6Yds2GAq8CGI7P9XQ8u
apVkJ8ULRSXFskK4JTcVKc51Cqe9RS6F8E+NOqwvFYyK4xUguk0zxrBFJVsb0iko
iSQCOjdd4vbs/WiMnP3PX4Q6YsKOQyrsHhObSfa2zSpxY/0W/l9wa+e4dYrMH+xQ
JF5sRjjwrOPPBbve0FIgeTobYx5RG6iAI36BvEb3598FdscgQlGsA3InPIlNEXrP
zsyveyD8z7TfPkYd2A355P1a/jVCy9dO2Sef96QcXW0zsDkvmil4dUPMvc2ACQXf
4IxloqzbRw3yyPsbf9o5Vzxfj/H4mbaMNAiFbs7MwyGbdxrj4PDiQh5bSFEqxqUn
LFohLrmqmPjYvu8RnduDIQXvLZb+yRUru/ZXtP8V0pWrPek7lQE9mPFqZn9zWLJE
BTp9qCB7RDwIYu5bdBEZt2lxTer74k8DD6zD0jbHYAz/rQuks8o2i7Wwdahv4xB2
aYptK7WVq0Ow+Fpeeq9lzlSjdmOGJzSCpcOAn8k+ZRKQKjsHuSFyIbJFsnazAtcH
YqQNbCEeaF1N9IRzl4BCVg35skDGPeiN1jx8T5PPkamX9+gwkzXV4KQZlKKnAccf
hdwbpcwITqYHhYJQ85A50NF0hO0cX9auaHHIrhC3pOb3+atTyD7wujA2qhipwBeO
vlvQc5LnaE+976HsXGkyWeyBDgTRfMxlvuxe4tDrva6enVPU7luzK1+QWGVJ9/nc
AL2sngZgNpHcpKKls1+16LUkATqFe5kVxlW0j8zIO8CpbaPwFeL7fdHkgluipTdM
DHSa0qq40WFR2Ksf+w5ejmVTK0vjhhvtct0+AF3df8JXWcWNk+HVqBpYvWry+dtT
lGHxU8vwrpQCPZ4p5dyDDDvEebVIIAZ0Vvn/ZGaGi9PfkV/OqfkQEk/70Tpoc8G3
FaOOmZ4I1BBEfYzlqtaMy0xts2Wqab05rLUJIk/UMwytGnugq7ja9z2TY6bcVKsz
lX1AAjOSvbjzHDpMKLjndFt7gSxsnOWgUfH+TheVPTeK6GotngQGB058AW0dp9HR
q8H+CqnlWhMP58p1qFn8mXZVyYtjrN0LKkAPVFBJ3fJbHq/sRCLK5QGZ1RP+qQ2u
rSc0PfNAi5Gx0gVxLECs9R8kTKSEBm91YdxY+MBuOoTUbXP9xlBudCvIL/g6HBw+
wtFTwD8QLeLD18gIO0V+OY3O3CSrEehs/tSLYv1qgOGhw1BOM6btT1Su+fE0WLJ6
lRoBaOsu0QvMhhRfkzsnff87lW25tuNZVQaijqELJuEuvg1BHnbTDd8lIM01eMcv
g+DxtMkDun+rn4s+VE2Vmm0oamhHBQ03HSfwouZdpRb2ioXbN4WNKDU4BSzJ2nAr
EEOaHBcd25a3heV//dmHZbi5OELE4uf20TQ+vRAumsFna+KB9qE+pgxJ2vS+10Zz
jfAirXdKXU07esCgcOBp5g7YTioL12y89+79dn6PLCY/q+162IQ/b7H4Lwleva9G
SzLBastS+5LlSGqK/z0yh3eF4N6j99z0TLAHXVKjnwG8LtQt2zHh4q0k3udhmJWP
UeMTLFliXz7wX0ruMAIM0ZoPoopIIdMgY2bL8FSqzLrVsl7wzhFkaEJnfzmWQn9x
EBHzBlPu0bMjF0LVWHuPF/x3fgGInaGFtlsOc+oIaer38zvSj4gy921tMELG+iM3
pocU6++nTkM1Sjj2lsroSDxbb9U54mZ4mML7qLsKy8FtamfEE6q5oeMK/uzv3wXP
t1rcZVP7ZdAcEqtRwGVLJ+Gl8bwpMCqGaoWomEMd0z40B006Mp/QqEM2aNQKB/YU
h2X4U5bqpPl+tzYA0qDuuoSbe/1+UH9N857BSfa/Z7V02aMgh8mBJ0T0iWs7XVNg
eT2VkmUCAaVxcJB/otrxvMLEUz6J3Tr1e8M9hbXqjJJSoW9OSD5xgef15L3si+U4
spUq2isKKm9Y1FOMUB4dntZMMvoq1riAYSdWqfKAP7P5x7VBMyAOLInqU7JQkC1d
Ppi6gxsVeyMv7g03G2v56aJS6N/nslZiJjeVo87z4QAZOIgR+FJ7keKD/Z0lG/BY
R/zGYrd5I9swXt51uUbPsk6kNTOrshbegecwQ/VY472ImLrVtSTObXPw4E4oJDks
LbgXy2VEeBgxAKyTIyKzvIs3qXE2WDJlXmQah74ROHiRkQw5SctfO8PAecTMdKOx
FDdNJpYTjll08KYJeKvojtPZyuIah4XhE9sTZA4meuAcrG3acQwNDJa9fzCvEqmm
T037/G5I7ir2zfzQlJH0kLBXCYwZXcdiiOKXSMNBYehIo5gtVKQSiKaIKSJGCZ/5
dmkxXO97klnOKhP8+stO7+QzGyxLF9Vxun/MPIvLBoeF9/E6GO2E5VSlMgbSqnJk
V1puSCQ1Rj69enQ7h8oQ/9DTHUKuH53tD2VNG7KXCsHVo8cfzWgzCtD3L25SHGof
tJvsKtEOAmSOsR0NgTGFkz7BG5sfvH/pSRwk8pgEoFZzNHNNJlgkJNNgQC96K9oj
Vg+uZXOklSMEe4if/suav/ErHdkW80st0YF+mm6K+ymk9poBz98SOck7g4VR7kqC
+mpHrbLFNkEMWEN5YQqIL0W35Iqc1XBM+RKZ2CP88HR+qJtjGT6qnM8bDjBuu3Ae
PUtBhe/b95njH2QGlXOsanj9WvNFVAXexwrp0aVDOiG9G5Oou943dMLtPvMZHiZp
1bCNmm1cBRRv6fVrprGa2l3zu0k6SazI/6IMf5yT3Gy/bqfc1CRYOYJMEpXmxL2R
uLoShv2BsMrIQxLgDN2IWza9zXm28m3XibkISONnT3Xmhfw16ulUZBTBp6kUBWj6
4aJlRgLlsFTGClkf8zyoHaFDo2+i3yEp1Ngn+P8kdsWiuyRFEchAeR5HhAcqw3qm
8c65NTDA0hE5g+nO8c59NCQnDVCXVO+hIvi3Hc2kLw3unGLqIw1wUA/eI7+WEjBD
z5vSY02caj8vkFBqB2WJHtrhW0R2iKDissKpm9HKq1S71wbuUquTpPk+ie/k6s4b
rIpWWbCZEV+mr9zVo9nJsbf4WMeWPchauSJcgKEhmaZvV3Ro9Hfxuzd6pVZx5ArF
YKD0RwXt3a8C79oQ8OhiBbAXYKqvcbt5WpsGnERVGc5ci9R3YLjsob+ZOrhgixYT
b45BJ8G4D6H3rRiC5xhNRHVdxgCTPXcEl+L6xzU893XEpQFHgTskVScNfCzc1CbL
tWA2rJFMYXKJhso7FdlnkL2E4liSBsgKI8TezDkIw7RyZsR+B10r9xkEh9d7BW/p
NTE2kBHOAbHh98P1Q0BM/ooLFCULxJCqtbGXn1ShWG6+qeqC8dyTIUANz0pefbAa
9OJY60WluQtfX2SoBpVxg1oFhIBqA/4dRy6flwN2QaTjjb45NI12rWLjEz+j/Lw+
/Sr1ieia0sXN+N8q+qKyRXDgN8DTQChzZ/I3zpfO80q5+XGow4r0wlvQCIVXIHyc
Xfwdw6UMwrQX3zJObmy4fdxGIfBnodyFsmtjqxfXBG6fqga5UeeX6HH2rkmM2Oo7
GJoQbBaC2jgduZgekSzN1fQlbaitSfN5xAWcKvCSmajniSH+SrgUecMcbubSusE/
X+CejobVzKD09UaIiB1w4lW/tl2piapwW9NeiF9RbTcFVOXM/EEGM42lK+qmCFr6
qTD7h9aZmzFxkko/hbzQVQU/gEmRCqztpR56TX1CTYDSH4C/Kn2roZaeUhL6mjAv
4rA1Yz+sym3obZ3RGL6/33e5f4DB6By6UTpZF4V5rlJWSN/skWgXF5bUQ2kogxrX
TjBSOme1XnBWYNq4wGTws2Hg5cmTfej9u7+UWeEJjHM2cKkhwRph62gEWarjqfi3
3x5YX8l22Uim34UWUZCUL5yxy7gizVcc2385xsl/PxqFgJS2pdw8ALfX8668YdUY
FosgZ3Us+5AH02mRAVfj5AyPGhxDwA0RmT0Dwumx6phRWfyfjdJ3A3Zcn33idRw8
uW+OKv9vEaliOLepKMRwk8O67aW+8DUa30Uu33rFP0aDH3BHeAPUsjeGa9Ywaa7X
+CjYW1bf8+JVWms3ndyBBarHuWqP48rfWk3qifYuDIkZPzEOZFQCvvVjI9caHpam
dSjN2OMezpijeQc2NzvLVlZhrj3Xye18eQb7zVVEzCGuvHJgeIJoCnI3+RtN93IU
nIZ/0LkZNf+pZaeu6yNfbZvk6GAWnjaOo1g8GVNMV6B/2ctLf+tA3IGdfQGMgJDP
Gvy3P5ZKa3xJxtucvspIuwFJZNNfJdOlvir+AslY/EcwVJFF6oC4Pnvd3HCq5WUP
CWL5qLLusrhkB0hnRvKNi4yHJc+xdY8DAHePwl1LtjKK/kgsW+1AXzsWmZ6r1+LF
Y5tnf0habv8ZM43erXPSMMeCMJWk7Iplx5GsQV9K+QddnyJpNDf3RAstXnCOiGj8
aSDD5Q56ALsg9KeiMwKAHfuTSqtWcQBFlR4Uj/VaFROKCFbWslUSxgkd6qPFNZVp
aoUn7/Q6jVWSpJxHPoFIz8qGoXNXBOgaTtVj46S7u2Jzu6wUJKP3KplGKRSIl/Oy
FMsGQz36ufuJ7SqYR12V+T4w8w8bQw+kdMKGoUH8W78IvkfU8aJRiHQRxSLaia1j
DG2a7NkMrAIrYV0acNCV3wrkq8YL+sXyaGJHRe+EWObKIi5fVcXMsmLJuLrtsykW
/cDkSVJvEH543pI+Bbzg3+ZeLC3dU3KhKUPQ0GrVzxrr4lSEK/R4dz8FO1QhCRu5
OysSf+vliiiqNeu6W4H4isKouspPmEFV198BI7Mm9S/db436mSDOGX0BhAaUvT0U
Z8M4sysfOkFrRsPKXn3Nu45SepokThIUtdljBn6xij5pVBBLibCbfnpIp2syS04r
JykEnQWoG2sXkDU4wuwpV56GigBB9pm6LNdpYl0i4X36Rajj+YPsChsg22LdUFf3
gxfqzM0BYeSDyUIvZJWAvJGSvWAYq+rqIL593I5NeUwTevV8Cq5x3MVt0XGeTYfg
LC8zuVSSg7janFikdsWjmiSK/Me0U8JMmrHc2cm7qrMijKx9IKOSobwYTxN4d2U1
P6ro/A/4c3XV7sXpEZcqg4gF4eiYte+FuobADQgfrmChvxQbENQA9odsU0Wo+kfe
q+9jsi4pPB2Sz6SHTRfwndantBHd6wYuzmzx485OUthzf+jDaRU7Ub/lNEJ1mXZc
vHdP4VkbmVfmF6GAH4XAo/c1WZpkByj756BMUcExmSLWiYjwK+zS+I8r4+F08nW2
KqbIJGEiAFTTnSPBXObrcohUT+pxFGAbti8tEVQu9jpsoaVjPwqVXutRKDNFSrCz
bvfm7sBuP2iSetxiaiOEFqf+tGPEj99+ol0Sd4NzzHQmOUUGagyCvD9jQ0yEMm6J
uNwaRMMGxP6c4Dux7BejLeErETD/To29WKS/7zHBruBX24eGNQ6zND9E2xwRmChd
62KbanYdPMTMEGA7db064ZlI6RKgse+lf71Vro0kesQIytaOlNfBQGlKMhuCv45k
2YWJTotbIJZ3rtSgtr9swOp6vgyg85iCwudF9x+by8VKFHeNubolqzHkXC3v1D/7
8AGAS7VKv+ltTM8mOVARnUfZ54S83jogoa79g6cYrzOSwKfWQu1kEe6maRYRdEDn
T2LIDtIqAUnM1UytPw5DulsOSwhs4m3FIIH6boQpDYuLb0Km3E3MMUeRkYljqGXN
UbK5I1CvuGL2luxZ2jJrl92Kd1wklB7ngJ/lKc//JY5MDz/5Ttx9DvfDam73640r
Tce0jmvgalcc8sPcOyxq3hJxFH/mOF6eUSWXGa/DluCSEemMbF6Yz4s+Koi9tCBb
Z9qZa2mHk0sN9j8rc8NjcluRwggIaiiqml87QyDIs7w+eExMQFquIMZuwouV4hSP
YM5qoc+nVFO91Ek6abFojarPsEWvBC3YPp4wzm+MXpDqoN9nS+x5OUhTegXcxop4
rfQlHU6qNpmw51ys6ehhTcupRHTbPLJoG+J/XMs1M87y7sukgUMiL6npXOo4aQN3
p2iWhozwXIxwlkhqR1Vbv+vjATdLY7NHl3WcvmhQnqGi6MEPy79knHoBNDY5KAqt
FeSMvnWBqsKZLTsIWJZ+wIQnxUz966FXzOADFafPBwt/jorPiKRQQZ+3OThwOiiE
G2iXyqZWoKVub+U5hR89xKxG+a9tAoQVgmCLyOu417OFaoNOsuVbL+2Lnlhgbu6q
dM/BzfF1tUIhGSe4/Zxj085G8dtIxcR/ZuG7bLPRakLDsCbgX3QSviMJU/WZVgIU
00xXf1rkbKzaJMlvQx9N7bitL4a2bMEBmnesbZQggORdhSdBqJvdLYMLZCDGVfiw
f8Fmh2f+gUDFzBwu1lWH8NKC3S+X9KE3GRi92pc+tKgk3O3lUH4ccbOsxOk3UXqf
Fi6tCDxUMwZL8Z0sgtr/IOWH7Zr88xPIPAsoWLk6Ntm9Eh+yPZoWpY9zXCYD236u
bB9acJ9lM6lofnFf2CT28iGOKArjDJJ88SYXudBvvigW03gqX9b+N+DmJeoiF1U2
BLhlxdzhEpChCgrNpM8/MPrxHCOUoczqXxdc88v97+1Wuk3BmjblcOc61i8FEHOa
sOs399N9Gh4UGg7FFmmEhBXtbcxO1Pe5DhZij22COJ4FPLBUDuBoTtuh+isN070w
/jJu5dNgvyS2uEtnDSw2zYnKvnIw+wqRPQjWg2FALehr/q67qE1IqEd0Y86R2dtQ
CTskHNdX0tcUf+rpNgKwelALBYl4Nolka+fZ6OX+mjOpzuEzSK9+F2aGBY5Ll4RU
gyKWdThxVfPIyxvFRqHzxEAq4RB367LDwlMmmhxYXzMwuc/bCficlfGijVmXlddi
/Q6fctT69HNn3RFfaCiOv/eNonm/lOuD3mXDmuOIHKNTxTeBnSniIqoEWJOsDtF1
kRi5OdwLxXX+uZf5upKqFVEGx9RprLb/SBlIrzpZjXIsbf1e3yy34LZc50cnGThn
bmjtX3LOgAM7WiaaicQUC7XEXJ5vXBl/KGks4SfGWVo1w/WnoS1bYicpMjAvvz12
B5OoTwG4b0IqqUBukGBpvF7JKe9mDZa9VXY0IUFAmNvWA5JYpu9NxQdz5yEvAe+Z
EQSq2DPmp53Pyw7+SgJ0xPYdhsxdUICmIw4jf4bvIkqctDmXr/OO+t0ykvCG8KqX
KWi7m9v+KOBd8kxhbX6PYwweFLd1chfGJjiRb7576tApQtIAH+7AeGjUDgRGnbuK
QP1GhPxNHVD8X2ltnw0e+FziPltkr8k0bZ8ynVLgyrpsY3Wiwhe7BoGfBgM6pAtG
5lkJMILmOnH5EpjAHKydeVXVYdlA5R0pyKF+ZPBe5jv1u701iYSuzDW7WvdtWlo2
kyWxP1w1G3iuqxhMAdU23dREOiD8+EPX5UQtIxP1GbEzwbZptm8Vvp4PYCpaIVgP
WYHpjKYIZORC1HhvW/PIi+QUl+DAhrqNkWKC3Hn6H1P6sZpbD8tg2JoKZJHezyTp
f04YzFnLqU5k9y0vRZMBnWwKABtEUlEoBKJnKuh60j8T+kb0TYiQiSeFQIb9G5G7
+ox1izLJSS2/WN/2o2KcbQHCPVW0s127R6AaUO/cI9WyQvbeTp+yb0IJc3YDHtnr
sFvRdjMssGwODiKLrOjLsCZIeivlt0cotqvq18bw0ZctmWo3ACnt4QE7shQ2Rvk8
DUad7fQGeKcjZyJRQaHGTvZccOGYhlXTSCLq8L+00YKvzc4nFMzQ2PM4BBIKLrdj
e4yyHtm7VV4CjEwzVNt3ruO1HnNho/+oV9swoypZ/Se3EoFRkKPE4UHruYrTf8XE
clQYezbpeeiFbl7neh/DOGx5730objFJi29lHnQOD78BBoPWInE7PDjBbNpdOZ9A
ctxWB9MJBGS71679sPxzdJc8grm3pEp3covY4BW7BTSS6Y5E9Z04ktzTGSjf5bt9
df5neJJwmlSPkivgAqqM0d+tnZojwkA06xeuW28txAk9kXIle8beOdWCDIvtPewh
0xmGh762xfqLjnCJ2TW/stu7QB/go/hsAhCRfBczYEhxYtgmU9NJFfKLFo+S84A8
mNYzEwI8nkPhaX4TuAFdnhT+PWmokg0OBYHh4RnLuvICnsy2xQPRazX22ORs5MOE
c3GJCgsGWhVJ+4prhSDPdp4G/pvSFdDBmPZNfPtclJsHLrOE6kgMm8fw3KOKq3hU
CgdnRhqHuSusAB6uE3AHO+auSeHQR4251+p00GMqU4MDMQ2HtTegVbkBktO6i7GP
LtehAdgznu3FQpOAw9FG0lhhIiWW7LM7Fngc9Dz98X7bbLLJnEPeUeqxPb3kFohs
uwgxo3hBqpkZJfauwYQQ8t31XlNHell14ewISlepSjJhprQfWOjbSbDpr+IjV11r
ivqxGGIbQTNmTDleniO5fcaeoIeK4GCZdKoc7idN5MpSfIcSfi6q4fv9BAI/i/d1
KfdxEZCyW3he7L8+e7KlzMGSJfJ8yItnZKwQiqLGe42YK1U5DGaJYeO5fqVUR4Sc
SK8wXiFy02SAPz5nSdS8q3q3bb2DfeY9/pcLfQ84Y8afhh8mRtDcOy5ikfdpoFrs
XddMRB4pai4JRavTiYccUStUFXT/2MWIt4/ltY74ZaZO3xr6bts8h5lTwdPdBfCh
4yKKBL0XXxVtpHaAGz7iQX9dn2g6MmbkS4IqyysNYA8u1+iqZ1foLK9Xwsqi3To+
6Nbm3EbnL51sXO8/eoX2/QmRxbbW84TmUeyqAgj1txIngFQXWCaqtqqCSZRos7y9
GNSMLUpqFVnErA4wYQVmK0a0wk+yJPtzSB+eIKfz2FnkrrlnfYRKgeIeMG3ithxQ
/EtGZK9RPvagOboCvqHhybLRnckJ9i+PyU1AIZBvxDhoQR2nU3iE99HjsQcIUrnm
v+XoeokwvKAigiJyLk+ojVK0J7RUXQdAY/4GRv4bANr5ihBriXF3FFJdt0Jd+t7J
oYTaYHtOEUwODjHJX1ELtaopLKMCoUJZmu18dXkHUL4YObHxAZ0C7K5L6Hzuscor
YFJpNLJzJQPzDuaHaSQWj646Uwq9lhsN+M0gyinYK1kE2M6y1gu7ZDItVLdU2ZQk
teesYpJZ1FQ/GOlWLevyvBbb2xeUYU9l902cMzVbGA2baZqENoaesr9hr4KKf46c
BNauTcjvWyi2ULJWoWcDbsV1ygFWN01iMVRBxbmhmhXVK+JmRJj6aRGHJVpdf03L
JwC8ebB3hB53z937XrVt54LJCUK2cz6lKNqF8HlESgcHVJTRtYNE2z+GDWoK1f6s
pGfB5r7/U4wO/yd9dLYB3tKSJIpnO5Q4cXWZH2IbYqtNxVoxPNVdwuDf5eIKgoX5
J4UusPGIoimDQ+XH/RhjbgeJIXg91KIWuMJQZoNQFUoRq83BbFE52TcLXRQZPVzx
WJD9sipWYz6nc55EuuZER8M6ZA/RuIR4drL0uCKi9a5uxE06dSQufwMFJBhuGhn4
BRX0Mpm4llcdcFVsmKCr0cJp3aXJ+qUaUTGlnB7J7J/q8v3qHKODb9WYUsYIO890
u46tqmpXktUwx62MLL1Bk9fVku6WXH+5RcH8jRvfp051EmH4bPJiKU02E5O9sbqv
H7VdR733RRqFFwltUS8WifrEKuWxNeHo2dmsW2C/ZU9+TYGoojB6hZX7dkOy7UYJ
JUo/fTYWwxvuEpFb9vu01pFL3QhM26YME1EhGJQFPXnRUycggjSkLEAGdHuKy0cQ
OtdgP222NEFBTKqwFVXdNoNgZm+Z5rx/gWu/KhzckPLnDaaemr8PzF7LyN9I7wFu
hpN+gKPCQiZxjxZmlgwKxc7z7Ug4E86lPyXoIQm67AAbJ32RpCY1YuGllkMixewS
BN5ad1EPNSdbJvb7Oamz9OgFRkbr21fqBikck7hedOq3AClVc8bH3aoAxJ4NQ/9B
HNMLtoYtMJ9FGxM9XNqcqgAYP+FHvFdpK397hcX4zJtjCjiq+HRBMX8Lduew0Rmj
2qCwuAFtcCrrlhbqyOAHleWctv+92mxVA6+8V4dWByLA0MzxNC+AliP/3SYIYF3P
ndlYMTY2NMe20MDSCNWUXO6LBLJFHKkMW/tvPDHucrr9zXozbDNzJGk5FJlxZGfc
IWnkBP/We1PSmL//wPJRQrsnLebVgiCdiWkzfaIAEhtd4PgNcGYX8ntimVakildy
QqdMaCcaCFBhxqnpEWKjDEUQQibZ2nQc6rDwL69RGD6qChNO0SwUdo8mQCBnsMGC
Krc461xGixjqP0zDM9HBlWMEUdU52qKtjELtSw26kL0TMbwFB9QnaNgzXuUbllnV
Lz/YLkXAMPDm0gjVzZIB8njlXJv0ott/yDsZYqAWI9THbY7S8TkUXyQalsfoflku
WvdUzDLlYMhENlTnB5tpYpINh3xp69Nmsf8XJLsxsaP5s20VhVIw+KcAWxBQZilC
k08hdtlgfQPbFcObZCVvkIFp+OmPbm8H/BuVXQJgok55JbQ8ewWaN5U7BMkZrPYj
OsvOZARPcDcgn2r9qCAcM00llyauVmnPruY9T0S3ApLvXoOa4xsSkLzSEg1DJV8d
FEQI4Akx8E6jEFb+wdQ8zxTRQVtzIofBiRuWhXYnvFEVm5FNRQJg19ldqb9q7lzO
lL5nHzGBrsfr9+P8VirleS8fBdtSqcSA6q7G29bmiEwyRWNBtIglvurJUnk9LacF
EIm6rgWEaQPdFCNsoQlI++KFiP6xGytdz89NRFcXEcwZNA0urvqzAslXGGHvNuMn
d4z68qZKsDmvrny7ID/vB6vSFbHJSx0yTmjIyPfPRakbgj5KvdM37W/nMnziGK7G
OvoQlggkK1FytuOQwEz5jcERcuwqkac9Ggr43BFVXNnfwX8YjlNGypyCQnRig7WS
XRQSsMMVyWQGMaqRceUcZHga+ailE/j081oOxx+eYnP/xtVXe/k7Kiby2GZq3L4m
t64VOIK3jupDoCUde2nadh9fgy3DQbLh0R+/241P8U0RY4lWcMynMegBnSXnkijn
ccd7psUWgWdyNFyFeABsoHVHlX+Hgdve5JMHCnyjQzqCNunbJKeSr0M04VSFXsnh
1wT5I27jodvRd987ZACaHpIrPhev1mb/ZNQp/OP0ZbE5HLHWGeV+WiSCpOQkOCX/
qQENy1wUnzwc9NdjqpKZsyfyOFO66dtv5gvdO1dxDiKV2xgj4yuntMjz/0MSC+Fw
YMpOeZTsL39GCVuDEEYOLg9nqs6a2GV90SMDkCWPHW92DucTNTz7PqccPIpcGLA3
ATRiF0Gm8SqwyvjSsJDy4kaQKeqe76Rn3hbsYxUJFhHX+8F2JNXbBF0zhwMJB6BS
NPY+25Fa9KIwRDBhW9Uws9sdkMW94g8HrO1VrRt/E1wUfdEY3Id9YNPSwDzhh0LB
bQRhh+ea/ZEyNgxmoy+UVdOQ986EgRzKBwIsXRczwR244//2H+icOJq8X8BbzrOp
YlxmcVbaVOeQIzaAAOaH87PMJjtM8bJ9b3Antz576+3KGpNghNjwAcBntFX3Rsgf
3Sd5C8phW1fth0z+VtKadBns417gX8aT/uO4spW4d2roW3dpPlRO/nFipjJg5ib+
Yu0+Vf8rAX7FqpjAUcsJ5Ifwu4cA+pSBva50ubydwTh0S6kwWesfJuq3zKiALAEa
WplBX47lz04cNbvrxtEghVVsmMFZextyvB+p0AAorZXrFDMptVkHqhjVgxSxiTVc
18AfzgA1Vxm35KnWXEQcnACkZKI6LlKWXjjT2kF0qIpOwkLD6LkiVxVWWHGuOX74
DDNutHdHXupJXznCPDEVP60ap6ZTCuFGHdRKAxEeVhoOiAu7TnXj8l/KOqTpaK4t
huWptDHXblVsBUUUlyI/L2KMAoAWkcUiz+LxaBdHicUTUDb+W9Kdc2hO88PYtH/P
Z9jlO/Vxy7tWUQkFRq+0Bjndr9WGnZjeMi3esZSN9zVYb4ck14kgVZpWeCvIsK+U
dDHJX1alTmcHcSHhhSxvhkZcFUAcJy2c0OkLkwjQPbzGFuHfoWNnSTBaf7WLHcqi
THDSs1kGsZyHGmkpwV2rA8lGAWH+ZOeLw4BIECzqORAEkW83o5ASSJZZsXG3jDvZ
hldVijvnSM0uhPMVOBT3bAQClHCbg+wJLTTwyak2tqF2obMWmuvbDhGMy1jl5S1+
jBzgKAfjfqP78NI5djc52WPIgHr9xwTqXtsmS3aWX5HUhCn++qH0ltlhJ/OILoM0
ShABrkoZd0KnXF0eMQsSXIWzExPOn/Vg+azBWXlduBTUbQyMjiHcDSb2I5jFaXf2
SCbEZdfvd1Z8EKDmRDG5Tx3DgtzYUMHI4EChSoEZ+HDtJ6hLSkQN8fMtEnUrK9nT
ovCcMSiyPtonJYjVhELS+1uv+XNCw9X2z7D3qz9EXIjASZ6gIw8lJ3QIb1hczyqr
1GkJraX/vGTi4tI01iMZXRH7ZQBnq2ilEd9lCJoaTyrZaMYBn4/pAPaBTEC3n5dv
eJc07pPNcKo5Lg+lTJssqD7taI2ZzC0oSSjt8AU4BTRobTQs1eRs+oD8lVq3EtrF
RxwSDwXQwMEwsS4KCVybJocUPJjmbbEUseFHq5Bv1PcHit/QTH4JuRTU4/o+1OGy
S9eurrpKq0E0BW0Pzxf/rx8fGHO6fj5GsTxeyLGs4+Wo1Rq+wAmxittngA6xIPqP
jbeWea/21ABYe/2Xg5HntIgosLFcLTEcl97R0aicpNrz2TbrVHk2bygToQInBXk4
CvH+RKGeCCZj2wuKr7vH+n2hJ7ul49Lr6HGp+pE4GSQv+hcPhWGCBq6qx4ZQfQFa
ss6+Pm+cUUYruCpyS6etw0T0YcWl8k9vEH5+EgMSPdGVL0Oiwf99KGxI1hrVpGR4
CehGLpjjiwwfi9ZZzCcZGXVgz1s7yysqq3rMxJ5so7xtSHZK01yT+wN44a3bVbMo
h1SKQHApV8DaRDm1tDtABnx5Yk5rCdRNSWFnb6ZP6rxm5Pac0L1g3YoWgFFq+yu4
yYND7grfvE5JGqm9+ENv2nJJwOktWFVxOSbmRjuLcHtQXGQIeQuygS8XwrCZnd75
ulqV2ZwV4fHP9NxPJ4o4v8ONz0vHNLkXwpBX4nrZwpVfbNZ7AFl9tEKTB2qotBpB
+c7MIkx8MdE+jjZIkgzAXDhCBX5bYapSRsK4Qj5cfev8TUFR4x3R2atSliSiaBst
/OJnHXrgqiVoFw4B+fDFpNFjd+Q/ROkWmhvQXRCv2Ocirvv7edQ+ZQr6tvlxIjsI
J/5ZjnZZV6NUZVbUG03HtT6jhiMNfjOlSyD67umELtDKho7rIdbtQmLGCNMfmZl5
bbJPgCLp06ybd2hHy/qba8T3c1Q/QmXWyKhSvk6pHisidbXRCQmjYcrLG49ORpBC
Ao5nhHXprLuj7RlDMScUVOCn1E96DEj2ehi/KPxgrkRuJHLfvymmsVxaTy8rGkIP
g9X1/kJ7vdEIVsR7SzdSrKwj8vNut7UEGOJEGpVxL4cFjb6i+sXY7LOtP60nL1QD
S4lr8d4znELDTC1b+oWbfYTK9XOZD7Zosx4tLY6NyAIlTpR4pyz4Qj2AlwaIQ5la
+FXY3XJ4Ap6CmzMoUI2UcIUJR612Y6hzbPrrEAplm8tHIksIKPpuVW1cTi6h//ak
wq4W6pl1OtnZFdZQCXaV5zlLDmHbmIQuFE5xTTA1ygtZtVtJGO9wBExXUxqbtyMc
CpyY9ca+fDoif7qt0sypyFnWbT4y6UB8+rLJVcodQmJQzfClNTIUxPB/vmSA9OoC
8I/vvQOdvf3FBq0QU/grx/cXCmutzy8QCQebOfQvFj+djkg5YbVqAMUigMi8yfXo
ieeuoflxcD45yHRUsqTajqU71hS9KSxEX/4DM6f3pJr9A8ozemsK9INKCgD6ablb
SkWwqSDrZAIL5zTT3QSL0pH+QtCnMTinW1xHR7NFtg7o6FcS3wcWcD/lWSeSeTQI
KIA1HlEzRIPLAaDJgpcCiJvqnOKkqk/s64OZrdOFoK5p/lMdLMp1b1BVPvnzHz0f
fE6LUySUS9Zf3XCiku2FLxqTsOXn9wS7PKiBpF4WYABfQU+of3aoyk0YtiqpyViu
b3IOzgKbUA7nIH8F1xj7aJyHznKLK5+XluB695YdG55KwYUOJOmQzfNj8WjwT6I4
A2n1tZYWGGAZ8Qryqb5QqfXAfCFVoCWJjG8WU6wDYHfOrRfqxmRmtTS4Wxj4mMHg
etuOEq/pqHfkFkFlC7bHMasMP3kxYlRb7SBEtv+zO1gCC8hqmyoUzl0L8qUsQHwD
uTHqEaKBACAUy3wk+BY5aLu+1hi3fKc8rebbeAS7BpoGwf3ifL3hkJiQyaU2+qKi
ZAZjfncCAKdOYoGVFKDmUibTWaRWRsvuPLVHuDxB5L6DDrXKHnjU9lVXIEJWYSbn
QVx4ee0QCh7HMoN1D6s6mN1MW6vHN7Z2fJRcyg7HeEf/gB6OS4OohJ+Qca0QYmIG
lvDfjHhgZfSd8TCQLyH1ONahBvkTyOIbv6VQhCTg1pb80F2+mb/RY7CaM0OR1Bo3
h6+0XMY23FdgpGiSe5J5wBqImqWKKq/EuV3R55qUkAgxYezNt+IPyE9yaSgMBk4A
cp/AFXdiVlOwuK3bo46ZJAPAVURic2OGrzURfdPm7ODmffm37KmXuc5mELl9yhu4
LaKGTbnJf0RxaHxYwQkJ0X5qt32bMoyIPvb/nL+FgubU83u69quBG5uY5RqpglcE
CaqaL5CBTjuoTN1mC4p9uQc4hufijXLpW7/rB+ovcV+5PyMK0wOc29CxWQj90Wac
0lcTPkfz4KNBRSteiehOAEstSpBAU8elFpb9BjelaABtmLCOook2VosaO52CFaP4
3NnvVjkHhZr76xN0FIX6KF7FMd/m7ATSdtO94TIa20FAWdEbqglkHLcvidEwkzqc
YtVdd5DKH5jgyzJy2oZqSrZVTdZZ6JzNJhM0ioVw3EjkBBw6XL1eY0J4V49R4+F5
c68u/54GaPxW6JYX8J88HfAYL7Zp6oJqBlLZiLMv3kriOI99ComJAJigcZrWjSH6
ys0ozCAoJ2IBUcsU33QblCiWnVrhsFmpg2KbRgoRQS9sd8osaDOXRdrjZpXruhyP
XXPUOQAkyHsQjVoSRjkw6UM+juB8J3rpGO+N9phbNpAKdLwcg29m9fNLAw2egv/S
QM4aBBA6MDpyLCWwuUxebBSzDSTqMaJXTySeAufRq5PDh1D4ZwDcCU2jBlEMmi2Z
+uupautFE9580Rb6TVjjBJ+kez8L1/TBLX1AjaV6SyPGKE/G2QbES+1Veqe5m6LP
nl+N2CcOSbNPYvANQLewEwUo/+UlNa3rQvvyfLJPNUh5/MJEIatIV9d5p/bz7dka
UpapbMhm2YlAMYWPObO9RtH0BSejYsSDyYdJE8ZthOFSsVFUZZmaILCO+4uJp6wQ
hxhhlJpqlyaTOeW2a6TwQn6DiGokAToNpzxraaOICcLk+r7pTlpknY66ha0J2OPj
aCK+jmvD0oKMRKEqIr5fXTiS4hkXysETPU8v4xXG/LGi0Sm9f5k8Wqh5yLURJAWv
fHilUSd7ya1SA00Pa16Vj7eTKXFZT55Obt3K3MJsTly1TDpGoPk3V4ZALuKZVZuP
cI5DBFgsDDXLKOWjmtuqQp7nE6rkeUOSh//+mjmEw/No/RX5MXPzHGwz1ICfFhEN
bpT6nYqHYxQ1DxckyKD9xIYk/TsW9wAiEWu3FUtbyhg30VING+8svmPEGo8exTik
Q/K66Cym6WEXhXGGWlS/Jv0/phP9NxtuVSlBb97BDyOboDWvRl7i/veQSfYiUQRp
J0e6fUc0Wu5POhlcDtD4qlkjcvKUg9AAWT5TC5RM1LfThv+ynyuGAWDKopGonywc
W/vEeTRgsT9zOy5K8Dj+OihJMrPHgxZOquUtc4JRI9mjBIYiN0ye4TonHlTtjJrW
AMLoKSJInmlvv/2avltWeVwlUdLHmVOlb8G9NF0LmkxkHRDXAEoTLTiQ0pqdAmiU
4gmHaJ06HsWBAn9RYAuxejixvOda/fkYzTJBaGcNL47KdpczvFXktQmY4EevMhcX
G5WhqGRGmrP1vQj9eU4LpwjWsTAy6k+FSV6HF4JZ3GwgkcvpZJJbgQTG4q57f1c3
PlZzjJDmeDxOq5qe8rG67WxDkp7BaKSQGMsZ0PAXQWMb2D557E2Hk/FDei/MgzYD
DkyIAM1VMuzojEYjqpYH0d4wKvs7sG9EzagiyDxDENKlka20I3Ouk1bXJU9/ctjV
8k4iYlxJgL0GYT9We/tEmbGxEHYYj3InkeVk25n/zPI486BwzH6SO92OpvUgKxSx
O1T8ktf5MuYl+RLR0ilUvkOkCCMbl0OWRctRm4EISjwCwZFkhZmvcQ37OHWNOTm4
QRyuAYsyEkEqQAbZUsMfmLjNzP4ezbcKvYeJ59X5JVTnpRhH9njswDWjc6FivBOk
NexHs05vbNOpnGnUJfxig1Wc0FqhyAMTZog5YOrfEgjpSKpwh28FdFlQOz/ir5oE
H4zkRYkBVs2LxDGSie2OgSX3EOP5ZwweEl7fzlsTvMMdW9/Uczzlz4JM+CHBsmQz
CSewW9V02ED0rvtnT++gBXyluAn9vo/3kFNjdsfjw8DqTqYygEHi2GEH/b3EzRjB
YB0zcuAW7oJd4LueHANsQhWnsImUIFN6ogsy4b9PwShtLBfbp1qj+raerRl0pkSr
AhEDRyMs4q+4dj3wmqhTWrIaWAKh6Z65wnOEVjHMXeyQI1P4m7G7YXnIMtHmT/eX
SDd5sp5ELp4xvjdgLHUn8dZJjHolQF0gfoKxN3BMJg6VRqEkSGHW19SdUY2y4eB9
iyCVXy8QNsI8TG0UkESLikW5isPlp4VE6hCCHnM6WqsakEEJsZrd+oOOlNzswbkh
FXwEfwEwVic6hf/PTpJhUPvufVmITTSYvMBfcdmfZsBFVzHzWjuLijfEqG2gldoh
tafY3L4+6YtLOMwoONeDHpIDPNS2sQOCveo7huq0G/PriZS2aUNtkSXeW4hDIoXO
/DC/MeQMhFULEYCw101sF0899E8WQyIY22MOGa6+VQ5GKKdRAHFak2GCYQ3tmPUr
pirUY3apYjbGja3XQJtcSTL7Hh66PpS6d4gqVWDeZMtMey4/JlgxrQ0xTTCjEwEc
GoqOrMxsirMvEjY1RC0wcBuyBY8YLlII/DtWPfByamd2Uv6AGBfdaGMy572fslh9
wSm1tnTdZIoUJWusQHpgvuvykFITjKk2Kiau1SIE6i9ZXegpnCnlkAMiYa60hwcD
faN6x5SVwf8K6Vu4lEi1opDwUjOzdWT+kNql44xVomdHICoOzT+gbSAOACOmP5Db
L65DwYCp3uUrtTda1DEFjwelqrhELr7LZbBLE18ZG+4oFZxrf+pmiigmlLvwBbKf
KBmE1dlAG9My8NZZo4BvelVggsVPFaBYluPxG4xMNWiEVxyPrPouILbqqq694gH+
4At9Tl+yUYxjFTqb65D+hjjXyHnYGvk/DwAICE1oeCJRhWtPY+P+X6gv6DfCC9zO
cgnGCXobKOujenRDUrskxPDgnbm2l62ca4MNc+miX7/OkHvM/EpRR+xHfxEqxz+Z
sPzN27UMx9M2U/HZUjx79R00EhfPpY8E6ysut8d1Oytmdz8yJEvWhq8whikntd2Z
YVW/La4bBD08LJWMAbLxWa+BlPSsvDl2vXTlTgTKXRLVB3ZerFckudkgeG7NDdaB
D9bJQDdrf2PqXLbvcqZNNwM3M/6PHtKB9mFfLqkTadzEOLJ/tRiiMMhxBpnhtXS7
yDdNcneWYR8TLn83G9LvQigqtd2DTND24KmqofN4W+NI2Ct8wHtyi/o4C60LsUaj
60clLyOvh+IshEBqUVH0eyXF1z+Fx9Y+IFsg7DLiPIHKXKpsqUEXUSpuMrwNCKLT
SHNMgIM0Ehn6gTweHl8Vxv0i5x8eh0PlYFs1NCxGgu1sA+/GSittso4NfEeIv0VF
qdmbkupbYC0ur5C0uUALoCe/wLZ6t19h4XiOECN1sVLYH8xntgdG2L0QAM1R6RfF
VPJ7Q0SRzjzI2SBbmfmF1UlWmucWxjZiUfz1UFPcnTppX+5U99+3kaMBoFUgm0lq
ooAjO1E9KMZX0LABC/Su184NorcKZT89MXJhw/w0VHgEwXRJakhmz54UF1B9/UmE
ZzkFFc1r0Z0FEoZTbcP+Y9IyvsDrHjiqjn6VgcKoyydLIIoslWJ/Coq7TTmKt6iP
WRAEhXje2ql6QcWx1HbTWz/C5CZ17xkmZNt+Ujk+SCaRgvAe4Xfj6uB7SLSWmJ/h
aTaNcmvVhJGpsB/84V8QU2Z5m4B+JzJ+/MSR+fOMrE+DDnDVI4RnWiZf/W5FZGqA
ob9oETFqtPObbHO1ygFNj59fx68ImzLYz8ZPBkokWS2NXJNN4l9xjv2AixrY5ngb
1MoXUiqhHHUDyevC7wwE2EtWHqVeQozs1NgxeFsIk+9umIAVCgrmlx9j+5SSrXnD
UNui85gc7axh4HYeHFg4T+lSTX5go2lSavIYx4T2cMGQ9Bpmj32SOuWMJ14vMSLU
lNMUdWmY9VdLpPpNp46qGpl7SeKTLWRxYsRRjxBrUV4LCuie6GInEP2anW4l0qHJ
Zn6EAuUgcnrRT/76loNsRZxRgJPvo9FKdiFvhkERu3tj9DkSBICoHFMjcPsydH+C
UzWxrmwgG89fpqctebUwGViFmGKJT/4opOSWwjbau2dOVTz0w3e/hzsjg2q11pjA
YSc/hoxAJH/8afCsqWGVIbU1ZQWy72CsiHJzZwFk8F3i9X1e7jcHKmCYNEWoPHwE
SPSRQM6a99TowJm2TGPLll771Bwl6fPc0b6p4D0UE6qF1CJDEs+WqAWwidWMxKpC
p9yq8qD4GOSoR4cj/hVU0UulGh/ivPOWziXR+M0LLr5zoKugefqhK5dypH9qJqPT
aeRSWX40fLhBshHPu+VRadAt0jgzUp+9HAMLyeSXZDbuZUVKFU/7WzXS5O6unH0Y
1/9tJI5Mz2KoZL/3kzCjUK49s2koi0tkFt+G+db+OGS7Dhu2qGj4JJ6vVY5GXXEv
OGvxZv/7VT9CozVdlIag9hkVe5UoostbQH2u8fAP3B6nK5KMHTTRwyrzHa0FNVs+
MO6U3kHUnnUo4Dm6I9VWj1QfIxroGz3VB2bHJIxI/MpjLqLl6bsMoVWIhJAu1OON
bMXLvnLnNqoZzlB3icEeWM3cj4mnPxpCup1zBcILUntQnZdmGbUwRRzcVoDE6GGb
2Sj2KlQfZXBdkXVt//sdBRMR5KmDA90q56SxJxoFc6yBOTmYt/P9d+h70x2PRMXZ
5xd2IblcjZnlpyEdeUuMgspzlUHivLQF2zCIari68zk9hPKk9BHcG9kLzVCIIWzm
vG0NNyRbuCEi3iNAiizzkRETi2iFFO1cphMWyqDxyLdcvVvxJBEqmKObdCDkI7kr
csitrkBOSW+WpfmjtiezpZG0bzIpFCYw4NsVbrYUNwRQ0HZnKWJXY6fHRTyUs5q9
/JWFVm7gEWYdOHTbk1T4IwZuUG9cxm9UlaUTjtfdbHpqHw6fpga/m9+SWe3O3AW0
ElAlLWl5u7ye5ouvbrcyqVn6UABjUmknnproCxFYW0xir6tSKHVlz+eT9Xbzx3ck
YtoYAGPvYv+mLaQXwLuca4bIw4rpjWGMzABB6qLvZXSGJHQSq/64hy3oJErAuwxb
GF1vqtske1kptdYJU40qxh4LYh4PJSqk8b06WuEtmKX4S7Qib8R3RBTFjgedLSno
aJtwDHo0adWMdJ6D2P1tMUXYHyJebctzqXFHpIt4edAEh2A/JZsu33pYlAbJuMnx
qS4yIJLkwUFtgBxCJZtannHEcKVjZ0HWw84Mqh1YGFj1xLYyysI8VqVZB1y2Glay
0UoxSVdWEB9H3Pai0pzmnZvfHk/LJv9ZrCM48chOUveiZgx6MYsCrKsD0yTQqgDQ
DZRpSy5rrywCeT0ty9J6wZx+BD6CimKWs2OWIBL0xCX6oCORlYr4zsrvPWehIpek
xIOg2G8ywlRTxyUekno+v9c9IB17WDVsTLX/Bf+2gD/XIrT5wjIXiFLCX4n4QIWN
HNCJwIwSHKZfaO0kU06b2WVSxoByaT4qxIZuw7OqREm+4ShlpXfFKw6W0Yf6Wd3T
7hD+0jp/guNf164z/aGh+qMmeHrw+QPNF2pAksx93vmB96TsjkU3moZ5E0rlsjEs
AUwejfvlM3NYChYvLFcd7PnDrT9fBitAb2ghrDdqknRLUmpLZCtuziK36+hOXPZ7
hPlWN8p7BJEw8XIv3T/B5gQOGY9T+HcnNov/61OrtnjMVZ2w+RYH5FsrYilgzKsJ
wCyMH/q3wI7yK17tKsNnSzbELFcxiAd9RdMeesz+RPnCesojw4awB9BGcyQfHNfI
2Jw/1wpyVA54161OFjFe9uRCRObm7TEJvsyzcY6QS9bwsHsUyMlfD/jejI4YiN+g
ELQuXm7VwM9a+vC/5wwgLR9bRIZ7rjhFg8dx87LRvFtELpdn6JpgMqZyl3Un41ik
ZE0Qr2UtcdNAo9x7mPxjABODA3yUZydZLsXYp2MbNSG1RE9REToPaKd6pU9MLeKc
TNM1AysUOoztFF+VfrS9w/BAA2OjUgUJzrhSGJ2efGc/IMpADCjAmprpm3+ze+81
VhI84UO9oQ7HWAMTYKTkc9Fh8WYxThIUoOeJn/zlZkWC7eLsSUn1Fe7zrajkfYPX
LKKczbj/9C73YKYhEduSFg/qi5rzJNdTJWCrKgxl3yV457jd2UvcHgFRCmxw1sBv
HUU84wwxONWdhd0rJFQcUpzvLKJxcOJU536d3/6gxWWGnyxuqcEl4Y1/pasCwn7X
yY2NTpl202ZkdonKIiKL89eQI9XDYSra/VwczkMTbtStqGATEkXJV653ltyBMxUN
vI8ctky1X0e3w0BqrpQTvPpF/e7OLN8B8GdVoJhKsiBsNQ3QmkbnQpUkC46l3EQT
2XdzDB+5d47bdEih4GK091u98/NCNUXMjhkBcNy0g1nHvP1zXxFkjjWbZUiVSlV5
2F/k9s4NP37GjScDSZGPbqqg5iuE6hZtHh/1sYrF+K95Fr3bLcpIjNH+std2rfu6
OTx0CVweO0G8/4Mv0722gmEQoPi+im3BP1PP5tJZjtVzpydihMDTEH72TnC+TBf5
RSvcSsh6fcdJMZx9l36u0dZ/RGCgNQMiyJtXXLE3YsunfyNWokcTo4LSKh8jCOiA
iKfAYJ8dT6XUWAOUFEN/kcd8zfcRiZCcGx15vqiw5qrWmdF9oz3WgS0sKbyfmKBN
KoF5PHEBT82dlIL/X8glDvJGdkskxSgww8yR4w0dG83Hn4VB9PvMWDe0meUp78Qc
XnKnDvrt4BfgIuGE/a/Sg3QWoj5N8wN9RG3lmv2NDEwPqg7QuvPWqmlOZMJ6/YSY
BLoeL5N5TWgj/8dwxHq7sQgrRuPav+q/nMciVp1h2tMALTkAhkLn5PIohwpVBMDe
6iXNzLD4knLONzUOQ8AMsRQlnF5If48Q4Q4tT16GoBtP7nxSvlpumxOX421/zvjC
GaOJXRRL12IQAI/vvcGQ3VEVC9B/agKsrlV8YogThvxLHTwBp/wYJuIYztaz3YJb
kbDa69lnO/6ocexGa/y8e8ZcRCu4E9XO+QPpn4iNXpvQ/l/Hmhl+Nd2yfOK9mflh
3+l9ExKi1kwUfnnSyIECA23NiHzPEtcZcZJp0kc35Ibf3yOuTwjSUXjGZegJAgYG
cbFjru9742h70LdgOLxKaMgxaW7VWkTY6u9yh9Gyo97A1KHbEojbfEK+Bx7lZBqd
6Z3PZN+XwGQDF/qlfhCk1/DT/CYOI+qKKGTuJZ3iTr3ifVaeM1VlPFLvocv1Ccno
ijdNRh02tmhf8LetANajGqjp4XHC6qQXCDLl+DHGAYNZ66AQy9LVvvao3jRbyRV+
4GQ0AiJhfGzqgNjp4zCC+A65ftVZ5b17kyTD0sPaszWi/8ny/OxWH2iM+UJJMR+v
mgXOjgkrC41hXN+LXJr37hPnAzCnDcuMLLbxGQD5RUSwjzyPlpyWa6CcKHtRSKph
xtIZwUFa2njmNuswe91czHR8unTP3/anxkHNLKB1NMa3ZSvnsb12vGOVcaRYZA9i
Ri6rw7he17csrcnsm6GHujaANQWDd39eP9egX/ElacyYLnpkTIaMfeyfwN53OQkH
3U1sNi2ZaiKS4nbG2DizdoGlLjSphTczzLYBnmovEg/V6dJ1jSI+qdDKOEOfeaq2
GJVinvMK4VAY2GY6BRsWreU0JISTnMVg/mm90dwkvgnQtIhbRZF5MWcSroyIxtMI
oxz3C/z6FHnrGBKzO3FZlzwGIWbrVXWxnQur6j1O48Fxnemy1BGM7NWFASqA+dIQ
aT+ytUTn0oVruJD1nucEJsc1Kpk6cgo3VQuHvZOmzj5wyis5xBC+9ZLlRyIpf8Nq
FuulPHi0D3zJWUaOsJjGK0FzLRi+28oC15y5yS/g+ePv9aE7j2gXCVKdWEUq4GCS
GzEBp/brwVPvpDpm3lHZK8m9plOzVNMJOfgxUyE1mnICMsaUGGf1+6F0eJ62ZkPM
g7y82K5ksKll9AY7k1PCiK5/mfsII4ldx5Fba7hQXX7Y4V7F20ZRyI5SDb8G8oJH
BR5vHYk52muPwb7X4nppIqC+LfYhZPb3XWy/WVqcTLsh1RSuAgRLghOUu3EU3tVR
o9BamJwJZ+EbhGmCpMfw8YuI+2N3kPblgE44RETL3u/VSz1gLLIZbNTwkBjigyZy
n58IMpLOBlXpyjLCDb7UTw775kLTE+rzDwFHf6yyPzBZo7WPTVbBghRy+rIzYwX4
eN+XRgeSa/CIHEcWGeFMxugjbQWI0wTQi4D516wMjxtyxje5pNZU5vFMoTJ1cTUT
GUcmelb7XSEsl87dtCT1QyciJuHttUYRvtTRwMxVO8gtbB+7egb4+Du/5FbIgPv0
TIJfNp+AnWB2IZfazWUjNGmcEa8xNWLUMHtOn/hTUbVnf4O20r4B4QJx5u9vMN1M
0M0SBb6i0HsMKtWUyswZMbxiTPrQYCQtwzc3xJ8ucQMa7WZkz+qopN/h+ECS05+U
KxXDQEa2zGXyDe5cLTLlYFgPd0xwv9EboFQn4dnJYK3gzKZY+l+aytLdUqdwwq/x
WRU0aRxto1F8FMsRoBbt3SdhANcD8PLNdzo/Tn0nzpgH5qTO6rRhnrXYUZiKVTrO
1HCBa00ghjdamEm4DBYPNt8Iv+g5V4wvT/hlJNjs1aLwaBxbakD4wHGnA8umpRwl
r7ehye6PmTLH5Q6RiyH4sJSVtH9ZQWzDONjuq8l1OQ28LiXK1Fr1H1kB/sJzGQV3
R+8W68Rcpps+tvs/ewsaubjUGJX1W+aJb/LrFQ+MeokefNZ01ljPdjjUn+rPGLXz
ZKxeurfItMTWmmXp0HvXt1V/5oFcc+IO/RZr/WjSxe4fBZM1STtTm9JczO+Ae0LU
t7Fnnh3Q24W3axXDvpRQQFApA4gr5mfcslGecc9EpmqeDqBKR99qPoVI/eDfiRCZ
u3LBa5jCOoe1vOjriKB/x5tx84q3ujOf5u6v1DklUyFzTPKQ4fCoGTneRksZFzoj
GhHT9IC8qtqQVQKRvPKpgaiTHY/F38cUllq3ZODvdCNX1pxxyrUnefcsAGXuv/WZ
F6xwFzGx78wfWmV7BPj6DCLqUgfqYTtSJ0xSb+eD+bDRCvHnR03YJxFTpEdNHBVq
e/90gQds+w/UV0wm+76setjzkMq8uHKJz2p8CO2TPmrmbGa3ICEvW2u2yUjJqhip
1emCAcOmRHR0RGM6zQ+BI1kDJY/9l40OnqLyNAhm9sSe17qgzlMpH5HKF/7kPpHM
6Ftfnu7xqT6294evnCil6pE8ARLAoBqMoItCwJcg1XdqP91/2sdnDvnmYVMceZ7e
iTYiUfu3sbmWzqtf+J/pFMgW0CTCS87EYNeORz3Zx8ARckWqBYqJPFZfB/uwvFlP
N7Zme6Okix5ioIOkQXj2DPXAo/pcBC8WVRCLRp/0DUmETWZJjdx43A0VwgDzjG3E
gG3SBYhvH2sk0fHzIwL3syZ7TP03PPku0EPjru19i20duZhn6WqbA/xXEL08afjz
ZqCWobMFk9jDUGICzUQds35R1UmUaks4cGsfFl7pTWAkh2F4js56eRFUUY4zqJcU
lze6y8eU6dY/sQnUdAEXi7bxacZUDjgMsSAqbgJrbAZgfhXEXnlnqGL/dfVnpgHt
fLJcdCVWZxHQqPKt1lyCcTgLkbGaOk7m5avAv5Uo3Ecasu5qrmi2DB6Hdgc/85BV
VQevLGDqMcZu0YAWwKwpvVdH/65uXbitHVIODU+yJLUtW1hxbRjOpvsVDyhwTJVe
3OmoNzo8U0IhN1HGMRvq89bRGkmpHI2jg6EFMufWtiv5evD0bjZv51ePtoyXHdEy
2HOx50KRaIF9DqClFxegaYMDoPVf16N/veDPK2fUDdFLVk5LDn44ejZEzUONqiFW
DSO2zq8RnwjN7FU9Q89R6CDB5ZaLfDCDOwdvKZyaeI9PRsedo/RNkUBztZsSg9t4
xd0F6ji0mWm/nPtv59HyVHlLSLgr6Pj4MmNk1+3GfZ0U34ADCvL3BMzXLDWfQ0Cb
3AavxU20UChxxqdDZnA/x5JWw0pA82t9sAODtrWWk9sFmJ6ydRkBhlZ0RC0/IxB4
wx4gghigoy4zfpn3xu6Lq6Ggvt3ZwvZGFSY2i25B9sQb2QZO3GaV018kitx6TMqF
cnwFSwj8j+ONBuQ5PvSdPhrdF3Kf1OoTKj19ioboUjhNA7GukOJd5XAOXiBkydrr
zl3JRNAAi6aJnQnpA6tSxQzGx3vJ6BsynJVi8+IXiNiUuUA2mJU0WyffF7kaEu0Q
yUwuDIqX1N1vHENRzC4bqIkuBAMBiceIabJNPsMdA5OUkaTRolpKr0y+adbtr8yB
PF7NqCSYHd9zNEGwnKh75ml+H7Pj8DPqKgnV5xzVlRqD5nElTPt/mJm0DVUh6E0x
AEU28D8WtM5VPYy7gnGIrmlf6rhDFrdyWrVUV3itS1IUAYeZmylLVzi8TXi/xuzH
ONJEZXwFzU31qZcsoSZstUOuwlMChf+ivMtOf0sFV7BOh1yZEvk2nW7ey3DN/eyt
Bv0eADrTXMyPegXMOCkiOXzcssJnxPPkv7Sp2FMI13ZIhMB+Rx7vtR1MWJo7VC+o
RIWEfcWNwgvjsRkDRgAwQN7ixFsWVSSPRFVnxE1nx9GUXjQFUDDrzEvd3vFFt/li
zazliPWNGUTOZ4aU5L3nAWs9anUwT0MGNqkuPFT0cXDFPMa9kk/VcXKqgVXu5bWi
d/VjYxW4K6T8gsN5SAmgCf0mRSzke4WXhxh5avz8gj4iLnchfPMZrvsuw8+WWgrK
BVz2c6TKdqEQ0NACiXj5W8cxn4MisV7XjR6Io4pRHOc1uXBMX3pn01oARCJMhfRB
3hjbQaJROOkxj31MrGD6ktPu5AN7Vk3PbK3wzRGg7wc6EONPFG1KL5+Er/DzYfY7
jQ+aVvLOo8Txl+gwxY8kUYSeDn8hf/cJxtRudTMvWDau5iG5gs365ADgjfSKVWgh
jDHpYHXCZD+3FG+hKx5vJJGFiC7/dhxK3BPfqZ2vYcnNuiqHj0kyz6qtrrG1wqJ/
wIacim9xr8gAuPT4OZPHP3qWJllLwQPXvT0nkenuOZln5H609S/dmJx9QtpIqs5m
sHPI0c6akNKZ+09w6KQFodvaMtoaOy+rJgSgr920AsuFWaYIlfLjWxsWV8pG+8LH
XKHupkazQqN/63y9rMBKZ1dsmJ7xFDYtFbb0oft5A9ET9xgvlt7wcZQQMcqraIb2
ErgTI6lrJMQsmvPlB1SexUzA9076YsuThDgQwCBTDUAB1L1bDkvyVjfQv5SNs3Zp
3J2b1xNb7qiXZw7qwIV/yzHKIkH/naSg5tFbHGKO5z5eIZ15O7jJpT15js/h9DwH
oJLMj8MazR3AY7tK2e1uIPgJ0QWdmp3+W3BCNT44F2j7UqTR7XeiapIyMBl//3Vc
xocCBqHw2FMRpZIzEE0Vd5PRufRmRdEFFHPYEA3ThjIU0hpw/8k/5AKTnSL6O/LD
R0T1rruu6FHx41FiLGXODrSrVNEHJvRt+lJ/mz/mp6B6cv/RYSvJxmOZOm0CRlcI
aOH796gZQnryeEX/boXh2rFmd8afsfhMonOcoKSmsSxn2c4cN5jPDDlo+8Mk8le0
yBm/BnWK05tF7Pz24qs3ls3Cm5tnuSTLs3sDBV9lyYZrRFPPdXXb9LTCnWAUYPno
9lKL3h3gF9vyJjOaotw2avBWt05ETDyoyDmegEdt8Od9lF6VjqXczeByGRDrpbAJ
jQPNS+TntHLXBzPkyNxVZ/5ljVakvyZ/1CThrFDdkHq1x7lScRBNj+astTPXtz81
ha18p1UMOqShi5od5QexpBZOfkjv15OrQEjPxe+QFpJAydYl5Xoqqjmz3V1DHjze
4O2QqlJN23B2sLDvCr2dDXxUaQhFaTO/ftS+Nv9aS7Zk+HXfpEkUQj0B1Aq2wxgk
UPaD3h1aLYhurLfgxciPySXhleZuaea6SypCNKiAKuMh0IlMQE4jPBd3QRKXL6jY
2gz3zZ9e2uvnQipJdMo+lPrWW2ygJPHBxCmIQnkSiNt4bYUhd0vi7AM1k0QqR0qU
cTpPXrNvcxnabxg/OyFaBNx0RBrr7YLVhbQVU5jPN9bgWFTsUCb6iDrwJTm0k9Uo
uiUN47mR6yosgZWaGxMfdO9W55+qe6U4KeXv6LUnYzWPOV6HOKauSQ3DNTTwKiwV
khH99cGelTWcVH3jT0Vu5Uks8jETs4cyt6ANgBmxyYQXPi1QiQVcDBRTf2F1BCCF
sO+HgvQgenj7XCuvYb9EvKu0VJC5InyAwZvk2pMo+Ak+waRzouhD9XEKwCWAUqUV
rlFKvadrercZciOc3dj4jL1BXEuwWKuPZ1PboXq6BW0x1FPfDe44TRQDb60QWYsa
rv3wy3ERKXxl+httEM3c8YWsW1jCZS49lGtz7vktNBtTrHUZRHKXWiV2qow09938
QsKzNXz0XlUYx1dyqgDc3GzlxnG8UShoxBfRni54ixnbZ2HhhQBqrJTpiizskcx0
Rf7+ZFJNmjmPsDgAsQed5S/pQLpwT+X5SRcWY1Qcj8PrtrporMnRLPy22+AGo25G
17dE+txz/wPAG3vCEa3gSfOt3Ke6vG6T4/DqFciXovnGiVPZc97LXepq1jLtOQ0b
pAaIZaqMjjniQTzEIHK50iz29Xdyj5VTTK8OAYRvJpiHx/PDKK9Yd6AU9HxC6Kst
H68e7XaEYNAla/yEOnn3/dBvBFgGe7sAPRcawk/eMnALsEQLJUuhdGGeUt2aUijP
yQnOQ2bICKTvOi9U/WO/q/AoRQiEI2wqtBvRWdLBZzQv82tURS8w1g0n5Y6RIzIb
ME0jxVpX4Tu5DGovmfhfQN2tSec0rGpuyZbzmZZrX4nnc3eRujcpvpvWcCbbm0co
nkRWMGxKeDG1bGpz3WHYxBDGz4iBRo8oV3MnbIGlLavWE0nM9m5LTf9W+pxrCHwS
FArmHnkbjbyECUyEzsGwgVc6wIopZST5R1RtD5nbKt1t/9lT4IVacYWGL24LTCoe
MIg4yZ29vv4iDxHy15q5eCa3+3zMDKSCOTxVn7gpdIbc1q1cnLt9/OrCFtJtniQ6
WPZUF46SL2gt4SIkW7ybbHLBAHW4bVOOuO7ItBGhhnhkexxB4T1SXPDd4sLgYi6U
a5BzyqIEG9FfxiGxhRjY9p7U9xHkexxtZGvgULTY4FKxMf4nmZ7nwrXkO+STJ+xI
3GZ58D/6xNbJiybgsqVIBtwst83CCXeJrvpSGncbQPxzM/hASDe2AZAKHJMjIKh9
Uq9xvyFc6nx6KSbcJDMN3hBcH9y+qKzIyK1aKb9eDcGHqjvzdO0vljzakTaHEShb
lvtO2/ro0JFHU8wYEiOD4DAVFlVJnkP5HFQA+CQ0o49rVFV06oSuxg5mIND6luKJ
wymWU1RSf1KbSv4bi54AQae+/WEr8s6c3ftDBdJrOpFx1VsjABRKk6CheizjM6jj
YcHst/UNOORs77PTJrNyaAc3ggpIiD9pIetK9sxw/1nScpeYUl9KlrdJhyzaadKw
QjD2FfMz4CpYi8N/Ur8oRc5grq2H0GXvHQjIF1ksXszZCidB1VCJnn/U9C2cX6LD
W/PjmAZku/gAtAfZ757CvH6ZUqSkekkPOQpCAO0Z9X8LKiBwPhoK+m+Vhbu57V02
oQhB3ouc02RZdEQ/GVPVtf48XtzzOBG2rmF9265ZdJYCAqzqc1Yw7LNsQb+hILZe
ZDvJCkCJdHR4V5B8yxMp682wvsOOtV9ZdIh9in8FdfgGeMV6lmtACL40Yy58GQ+Z
zV/CRaO/fXaOiGPSB9fAm6M35XTsEZGe0rTnwSsOiOMx7h3HfxfEJNKmiis7fN/p
JaMatAm4UEA/SrBZALYLI1Al+v4pjnF3uLePsKBQEsh54GP9aMgSyUvlcP3xsP4h
B6sRf8AD4U2CZ1QNGpdzMm+uThsZTnM164Bg9O8BxkC7UD3zJ2RtqRAlltfALVt6
9HmO+cW/AzWU892MFLtCxiOxponh83XzyZIA204h9mf7rCH/Rorwdk3CynXjufQv
UpL1iFdK3FmDU3d/fixNlwqyvk5P80dfdmMNyAirMyqXisppoLiASjSmOo2N6OlE
RUUoU3wiBuKj2R+yuliUwb2ZCnXfxZnW54tIwkW7ieEHgFR0WrsezwakYdyrR0Xo
HG01cnhOjxX5/Jt5S8WABJVx6Xs8TTbPSsF+3KHM58XksDReXIXHgwQgUsJJuitT
3TwQIpyT5PV8rY1fqcEQEgBKF1dYjQp5Ag7gZmlLiF7wB3cb3Krd2HjkFutf4ftb
99mzFlfHB8Pr6u3GCT56suCMGDFsJzijgXQZdOfiC4y107W3j66E9eCabjGVas7c
lhqVpuPUfsUho+19N9Xd8s1PVgEQjLcjXEmj3S+AW4Ht9fG2XMQWKVwTjSsSCfd7
vPBT+Txe0wykijk8ZgR0/F1ns3zXI7+sp0nsjLxMigHt/edmYvbl8r7LXn6rgonN
jfxvkMsqjeRlCakJW/vqLwqn3iHh/kBEFp91Yi9kgNR4oA89Q/XqBSnJybcyyBfW
YOLSptGVOxiobX2aXokmgjHmKiz2/mB7tKPBXEdAviNO7OlNF3826b/SR6h1junf
zS7XLYxNMAESjxyPlqYrlPdpCTgNx2ty+u8Y14oCY/VOZo+cptIpXIXzvYuqYzQ+
LAMdmj7mT2aQl3cGtUOVB4cH53/p2eqq535Lufcks9r804eb3kz13Iy+Yl08RA2G
NSSqzA5P2Lv4M8puvshePfKZJQs3Kl/0CKIYTfIGsSh7wTz6uBdCre2jAUrc6ocD
6vYOPxLwHZOXvYu0agUj7LPIg8KBtLzSKyNyr6RjztuZ0tMd8e1+ZoHUafaG/JQC
zOxyKObZIiIFeJ4x+o2jx6wrWa97p/NqdfLc5V7DCfXnO2kxddPwG59zgbDBXZ9v
wBfjN7IzYtq6p3UcKJArBxwwTd5HD39w3nHzFqh7VCOiTtgjnT4ZUAzSeM+DGNbD
urNI3A8qNERjwWaKo6nq8dITWAj2dEfyb4kE1ivFsgUgpecMBNbkUMZ38XN1nNKF
fH00r14vkY4ONXUcHWDgoSzpXnab7U4kMeta8450QwqoBGCZ+Z6VT+AAA0uyryGq
Go3j2Dfo0PtmAzw50LoOMpweByJrJLO05yGcMzissw7rHvSNchixgXMknlldO4Sb
BlcSiRwJvuwI3ve1/5upDb9M1hnmzUVUYtKbM+9C+TvSo4GQnOi87zVt8ToRRe2L
iR2WYnbhnqm0p6KBb4l+WVzsPgE1fF4RxpzZJ/kMUWzR0pz2Tyef0GBl8LRPnkaP
ZyZPjOh3/qe0AaVBZYUjrqT/1jJodDGQXak1NAxcUwafy5ZMojjfKFNBdrznxuEe
cHxcCFuoeVINnBIN/ESdcVY5N5UkEzBAjdb+0fRlT8DnvTvJYVMCwAEDNFQj6HAC
10HlZYUIoF6fzqmJt07eRLOobyoY2/DhC0eI33bwjEFSkQ4SitxBzw37Xx3RqTQq
Vr1CtYPsJKlxA3FVcdh3lrSYLbnXKmsLtQjtiDeYL8J7dCQWY3mjcrZytmeNRIkA
jJK2zElwz9I5Upy69WNkYR2sRVAon8AlX4wN3/+7kAjG+p6+LJ//8D4xZkukbF2s
6qesxPY3GYEtdXQWNeTgYTRRmYnuYvIR1aahSpITQniNaouaGkJ87vwEFjcc8tbz
ZLI5uK6bpZm1WXvt3RUFJNgbY+cowSFgzF6q8xUS14xWxK3w7GslpufYoRK4YN7F
mVHynbcWLtMCiTUOGzYlHTTliOmu5tNpRooQdrpzC+u0GC74t2Xpa1af6QIsIqgs
KQPnhxA7bLstJIV+H+h2gdEYrwx9hddBsHm1GcBbrqGWEUzyI2pcy4y9W4NSycz7
qr9o0qIAQoO/iJN+yxEWRuOYaDfGIArSot7VpAO2m7QQyMFkwLxpLGtZ99l8G6L/
egV+pbC2pTXbmaFVIeeXQhgvj+7qQlO+nrsxU1iVaFifWvTHbZZum3MJwvZ7mj6W
gS4Ol7iZCwjrhpYWdFYnGvoxiNQl44T3JHkXPj8vjiK2BaLKUTmu0PAt8/Kqemd4
Lps8nDakHTsxICG5RBRJMtCi1zJ7Bhou1IdfD/iKlb/WcG+jel1CQ3T6m8my5GYn
msvkj0CIAd3lD7ocAnSrdF9YnHIgPRaX21cYTTuzmsL8xpcCXESQJrntuc/uYfKg
a9yB3Y/Tqn+ZwZch08SXmhZZCCWhiapc3lYcrcg0Iv0PbkIAPvgSTzRWGIxZLN6V
UtRaCFgpUtkHiApfgF4hkwnkH+wDB7d4splcYAk1MAm2qJhX19Vuck3J9XflvSOL
UUib0prxX8KaduWjLVXVYZvI16zzwlt7gYJ3Ye1PJ1CPUScyzHriqyLvb/jqwUd+
SIEXY6x2hZ5Ki7Q48lUd7B0qNk4660+bt5RlnFVRJX0Hy9lX5nXGVLVGBhjK+IpO
7jpCKhzGcJ1z1Dszs9lrM3LMi6tYG4Na4DJy7bbjMPj7rX9S+OIfIqbuKcqVk+ZE
e/Dvi1meSUBS3CvcHp+cd5JwfNHQsfKsjvf2l9D/H1HLTrtPp9DxGbfmDVToHneP
hrDsKS5tjZWqftv8KEr1yaW2VM1Wg15DV5+dF4fdF823N+4d9Y6JSbWQZXzflgon
rCI2bvBfk3N1HWgVDbopX7NvgPkN0w5fas6NMc7Og36sl3s9Es/hbvJqIs5QP7Mw
PmI9zSjammQf84b2qEUx8Rhw3iiwTnldm0tK6x4ikZlLaX45dUO1TOlGqVD6nvYG
QlnelFOYRpWHMAWRkZKb3i3y6dyhaCbLoynkXvPFlmKHeSoeCYjOj97hW0vT1tpr
CUfcyZRx+E7UmA7UFGJPD7UKzvC1pWWNwEJ6RIdXHfat/YXLz0zQKgcEv1RKEM5U
lfcsBnwiaOhTm+XrzN0eb0kakNUpXC3IKkRONobo29z+cX29h25E1R2r5Hycgplv
rNsWBszaarp4+bl+9/nHyCe0Ra5Uw4hvSqI+qsCBFmVXXMc3/JzY9qM6cABTeCeF
apJk94VtbOjMoQXcjpOv9hVAOpuPLSNVTJugGHUZjq2CsEI1zHbRZzgU97VIuwhf
yUiYxx/O4ZAFaVGctykpvoXUQf7KSFgSTtY1LLeK2IJmkBX/QUyKQzaX8dgdFuGU
VAjdJQnWCwTkEG4FcR9zsEGGFFxXCQ2sGU+BtnMAdH/XdhzXL9SZcWq0JCqjE4pN
UatXzPeIAKZ9ThHJOdx9vVIgz/toroeXOvEvwq2Wc/7FcqiRKN6bTVVxqzVbLZoi
abjhruy3+cKOnI2hU1vZPlPW0+dRU9uMG7DvZvYoKfosINX3GhIkgW8fqAe9Hsqx
wfOgiAqjZQIfm0SF1Ick7iXrP9jKY97CduMAbqiq+H78qKRYyzSLYhMS/2geC8KJ
nSzYrO2zYINdN/kI4n/CvodZjuXfXY5CBu+jJERyNvqcoEeu5OZKtpbxlodHkfgH
MNBc8KGB7HECx7eGuIHZRqI1XUsiTObVYf+FMkMgK0aHzqES82n972JCPiacy+eL
OwhXorCxmnwnlCd3HlwQjvI+kt8WJ4lk6v/UZe2juE4cjuTIHqZLP95aS1GUSFvY
1nwt0Eu1U+kBKeLksAzFiyf3G4gAdbQ3LQxSftmHjK3cnUJIfcEXJa35HWnNgBWC
9RhrA2HSaOQw1jiFIfWPjTUiUO6crXsZXvC6ymCHK34HGrxwEyj2Lk4VNHNvrqfL
IEwU5RIC/2JB1gPp4zpRuNU6oOplL3xJqaBuy6zE17rikgsOeZDBvJIGc8yrWbWU
DcuRMl2RhsbfvMwxWBMEYL7pB4rZ/4Kqf/QPxYCWQGBqh9O8d7DCJo1uZ5CqR7l7
B9KAblt0BNsuLFL37o+EUvyhrIQuXuTcMIrLGqcCz8M8quvRUoTdY4J/Nli0hHwt
pwX/EJjUi0eQX7wDz46tZ7uFitjCoXDZOpMVNTvw3msdqAGHGOiG+VP0HWZ5NIIA
5mN6qvHUkk6gGz2wQsenBBzh/6AZ3PS9UIDegCzHtTSn294BsXOn59Wv0tnc+IYT
vMoN4NCgbVeaaD6Mmw1vMPl9WCNukZV3z3ym91+TNKHpSxy4H8eRs6Iw+gYtjYch
3hbuXfxhrJv+klFgIsqgiZAnE6CqKyLtfJBTmknMfag7sX/nTcrmARnrJc19EOMm
Eo5IiGHBoMl7mJnJGeJOaXtUOb7DCsJ0ohQEymjQReiPELOtjJFtAlyf2ve3MTi+
M6hx9ycB9pJJQSZR0f2z17M+HG6FwyVR7SdpArzGR7yuTndoxuHn24jsMJaznGkL
lIUAkTc65f5lWc9xeonnUnU9zsizXM8EctRDHStsOaMLcf6soSA+fGOAh6mVs/8x
NKKjZboE6Aa16X0sEswxovnyCpg5tOjpER0o5d0su/u52UgNN56JOuRHMYB54T+T
06WfQc3RPG8ta+uKkaGWPKJkO1rX7pOBG+BfAkHf89DaHUCsx3dZrBZILKq2b/r2
u58SfLsJUgEkHqvyUw24YiVEi45xNUdAEIWdzyLM4kYiY/uWFT6Gh9riMPXQOW1V
vbn78xSnYwYleGznLvFYtm11PR82VVIgMSfvntWvDLQf4124OW4QhiaBT7Ht5+Gp
0Newu4SibjVoqPw+HkZqO9kj/cgZ7wrf6cZ4M2qO/u4Lyi1ykQTzU5NqwV0H6JYD
PL7fO5KNAY+HlFBJVsEI0ueS+dLl09vCbpec6UHOgvOXdxGi+5clMB/9zsutLYx1
TshwDwlx4DLVC0FhQAGd6MoUpb7tvBBNwUuwXB/5QW9XM9eo6apMcb6mHsuD8uqX
xiZxWEKKn+a1d7mIpCe/qDO2ruC6fmMZdYgXNhab3WDAPzDJ/u7hO1T2zOyLpQGq
NeYZ3x7iWROFDFQ1IA/A2lsaBQHH+Bz/M4MDb9POnkWcplDWCzSId110i21Ruwai
0qeLud9QEQPrudRGyBkIMl3bODeZcCXg58DqdOwkFHQ308eYtOtxqh55tyZLUqT1
IAiGH4sKd8Z4Btncte5wUgzJqo4jPRTNwRVbnYBkhucw3hkJGdu78YTL2mn/GyRn
AjYfp833Hxw9Vaynnn5vGwSAgD+Xxko7LK8ZGDKfE0/C12euaNLVd1XLJAa/n0fV
jYzeTxwZmCxTRARZ63AJkf9nylnn49SWuXte2Z0ZirG/mKfg5JI7nyI6+tyhm6B+
BajsyJUKOD2KP11MCKSwP7DA3FYFUo5IQ9pbpqqD+FCMMrkxPC0Aa98rPuWmyr51
quRDNS2YKCJH8RM9U/OizSgVe6C2qCZl1XKiQxRYrFEpOFZBGo2pcTCfsW+G7xpr
2iRrpNiqqPoJj3m/x1+ACM5cM1Qh9xqbQCDXA/EXnLUVEM/wT9qZ2syyJglR7lAV
yZto4a23g45SSkacu9jE6yEVtE1vZ8P1pCP/afiwPLwa9i04s57s9yNSRGLfRWfT
66obSgO4g/5oAZ5CujSgoA53SFjJwTI1mTV3lKLCtbFJf+hAZAL8QDpts0cNEQGe
nHTVZRv9UfInZIWf/EtMkayMMqlsoWlKawA8HQ420gzqiugy0/iBpoOLCeq2n2EJ
+wohZzcblAjGdzK8K2cjeNUE+rJ8rwEtyWg0bLyiEX8JeXRG4RoKCxGr2cmArMkw
/5RDmRHkW678rMj127kPy6hDZzdqV670UmRV7Pykso4Z/AMybsgL2bKRUBw9lRuu
8IOWuwMOR5pdC7tTL3NxxsA1PruitXDL55V18gUwWvynWPLp6wK58bVE5gg9qVqm
0cjCX1JwwBM85q3cchj2Dd6ZR3K9AA2i5y52Z7AxFvGu/LmKqTmLt21kAS0Ki/6L
nX5V/0whwP1EwP9JAqHNJ5U8wwLc/i3V++v61t9iqiseS2o0/KIDc7/gXPh21sAV
dIgqnY+fvuK78L1VMcBMbU0hxxdxRA9Sa3L3OTAZ75sLkPMZuN20RE+OjwtlGx9L
ys2Po0ChIaWsZ0pYPjpxK60XMrEwgy5u5kCZtJTTr7rlOtMQ95c5sFgN22wieNdJ
D1tRhKsIWLm58wbtYlXcNFPK/ECxVSDQHvqSIN50lmB5SVabknIAu1tSCMNu0Ozp
umJlVQHCrUPrwjdO8CYpuEBaSSIV3eOSaHdOBKY6Nwu2/5UlZ4drN8O9By8NFs4V
x5dVFoGO9zkwQuSiRdR6ip1BygCbZzQN7I0E8W3b8iLficQ1Qj7LODubr2cNdx6m
jCLvKRmfG0DGmYFItLsfBv3EgahX8hEqUV2D4JI6VpTXjuZBlXv3eXNaB7VURVin
IG5F3aNQR4AVgfUijG5vS3BF99nR4+XRvADc1z/NPEb6sS1bGyJ2DjxYJ1PkaSHG
IjWqBFZ7zXuIQv1fs7pWQr7pGxcL/nUST/tA+GHZurtcK3U2baGQe74DCOD9boVA
62MftfUdGkLkGtvLbrBtCJxrORI2VrjLTVeuNQ619o7SMKMW9pFQ8R6owuaLzgHC
FklB9uOgOHfrrxE7nDZS8wupdWX1/AZ9viw1rXlTKIHWDJNatBnYESimm16J+e+M
KBhM/DaUvH2zCvxDP/9gzmuB9Rjy8CcPGJlEEL/XpB0m3U4lJUsGKAGKmwLhdc0A
r67EU2V67s80kFD5eyfIskQMYt1wObyrQoodsuoVEP8QdN8eOfbm9xdo9ARX/Umu
X63ADIeMV2aRPr9WTlg5O0C7TLEgkMX18rxerX+Py6Jq5Le91tyC6hcA96IYWTFd
Wo3WR3XHEFs+rYWS5cFCpc3MfajTcK/YbthQQbjjyN1zW0Ul9i9dyL1467l2//Ce
C8fxNHV0hDoKaz83Mbz0NsxvigrD1hEFphiKam1HQKwwBwxY0WSM5SvFg+5NDLe9
ygYQT7ARO2jIX0r0n5nabMVU8jleW80FN9HlysZiDt7rTugs9nt4mYPVXa22AzZf
zZQb58VhosnG+PJB+lKY4ko8/er2eUsnfQCfrv9Pzn8iqpNiDHxLDp/vkhM3tQlU
dLVTEs2MjAW2xoKapTqbvyHnC9s4Nf83Y2Ib7SfyzaYgmUJIeDJmXMpUsC+JTFfS
uZfIzVHyg40gcVhw5wn/c0KlhoD8AmYBYEFQZ3wfElsu2tfpoUnLERXC13JDIQaj
pxRVLlEyRAgPkg94uJw+AyzWhHM9wNrFbvst2Rqr9+YKLBzdF3O5TGVRNzOT+CSs
OVCj+dlSoZRCvCgwaVHAeKMEFGlg9VeBH1SP8W6H4hWoXenMATNbO2R2HJiUCqor
mbnF78GL83ybo3egLU9gujRnuFtp2ZBhizqRWkXjGy80dBG2+xMSFuiTAwgE+GnV
p63K6TLTsqKfYkBK1Y93pVeS31+tMAzVCieuA+kVDE4YiGbwckxTKtNIV00lwXey
lHpD+NAASZpn9lTjn6/RBob5kCyMiYeYXx5FqEQoxFmr9P0mkouJFIJxZpAdl4Eh
Ft/jSfqZ6wy/PDUysJUZpDH5iQ58SI81hoca9s9x3O0sU8F9bdkpL6jX2tIhcsSg
oSjLLT+zIEvRybhPejdg1UkKLCdR5vTP0KWiyyln0HRZ0cfu8JrEQMQnxL6FiV2f
FhMb0XBYON9EYLnamW7c8ZBoMl1+vSh3Mr2Boh3uDIGZMhzTkkVXvFY6DRe8wEMa
zghqMXRtIPqdxhFPEmBWAHC0iv/NeCrMcyhv43zZSY+/ennaxC1bFRfY5vVR1LlV
inOiorUYYtnBpm6x87DlrmRP6dfhQpwB7h56V/c2MfvXaxnp2gJ74IS4ywAWwrtz
oSxGn0PFj+xo/qo9FTusDFrsG6AnwjI5pCWn/wRLreyjEmJ5jFlwwQzxkuCluWuk
2um8F2WbnGpcnXnYGxr0C35hRlE+qHWQqugF0W2ubyEDFyG2jK2eEDJ6BgXLa2Fl
9eMs7eVfUicbeTDqP7z4uolS4Y38owsODualir56KTaPN54SpQcDTCDaehO3fFQk
oMBVRw3dn3WrTdUkH9Uk1ytbOLgnE9JZjLCkVIkguxIoDyz9yytnHwaaNcSO5rBU
0wsy0xNj1ESOghADpyeBFAK+Kpia7nXShvzxkFhImSpvcRclpg8XVeXy07qo6bvM
mUnAhR3jMQlBCfBMFdZD7zDQluEtCU+vUZ/WAFxwSmgoY3ew7eEkucJtOaftvfuZ
Zfz4vjZPNJfuvYsszcSh7YaCgU/wekRSOxcy9u/L69+c3lqSrnRCsAn4lAMBEw5T
si5kDDNQ2s6YIUgqYFzdY+6vuUDRzq6E5zGXLZKlRYlvVtC8KfugQR0B4XYBnWsl
7jTCdfFB/3xZm3LlfWG/8HH8AXg5Y1p/ZNTTfdky8yn5MKIRlexUMPaNPKxpnICI
OUCJNd4XiuBLaTfONi1dywjyu5BxsRzfmfnOOjUWznEvcnuV76EbwyMaTF7ynVw3
h/Te+mvcvH3SJ2i+oVLTSyrBEj0cKydndVS5gfflcLox3EeJBt3oS4xYki6zxSjF
OZa517wj7jlrRc63kGqh6jfRDGsR8Him0PnjFDo5C0yW8WDA0fHJv1vgTnA0AWRT
IkdeiZUM83sgKzXmU2PvB3KrnE5LMLjUlvkGWvknfNqs8aVt/UFgiznGw8FrGsRs
39dXkZhAF7NZYBUngtbZiyvM0rftpwRkkTs0FYZHQszKSBa/JguHMfI8Pzfx2g9a
zWDa/fWzi+NZlw5Og8vF7qqo3ofeGNSnTJ9ngAyLhvfIIB4iKqRdXyW3FXeaQuif
dJda2EWdRAu4OGUyMfaYvijKCdtvuzRmumwJC9OATgK4YFqZpy1DO3Q6h2/i41Cp
imSKZUrE7trnM0IHgGG/8IcR2kMbmBLp4GZzL7ZGHkKd3UupWmuCQaOFRn40CZ9l
HvcGoZjOjqJa2wrdpnFSEnUrYErDAMZFBaE9hd3o5r4vVBIiWtQDEEmYwYkzAMhG
DwdsBgmiURhAOn/xarvMW2fwCjlDtBtJ0WRQtAMHFkDpoJQqbD0otLPJ/nvuhFr4
Bcf8tX2bUF9ojYKfFBBjWcu8AxweMjUPcMVT3IkJNLPk65Vv+DkSxKpj/3vx7sEa
aKBAV0tKahW9WWw39yPRJykefoB2sgwMMxLs+Zd+PNBUV/UTbiX9By/aN24e7JRI
z+CFj/OH/JEkM/v47WveSkdQXl5HKtayeT8oy1g1eILxljOdFpzyiELkEONzIzpk
Cw9DtqdlPej5IZU6RQNGx77G5bR8BrRrPqJk5lYEDfiRAMMXd0JfNjOPeH5Rc1PE
HKDE3uiMqQCZ9x8+yc7hTLcLyPFIe7yKsA0Bk6+kbQz2PLrSDTkX6mHcIk1n6PB6
CYo1asTdo1ixiIM3t3breIHPd1InD2FW0DvkDTZibnepE1Ft1/K8STSokAW9VZwF
fqP77Jmi2DKoleGr9XjIu3l7nYwiNnJVlh/o02lPq/TnblbO8YTjSyPmdlcdRv9H
CAYVx+BEtlpez7SxsmDnkmq+6e6u47f5K15BA1+nkHXRPNTWvyX00xPFYupEo+4u
jm/kdueNoB5SDoad3CTFKOfxKnwniyastibae7OnsuUVUWVUUxyCNkymNOLROuWG
AaiJZcUCExBjag/cI5wSJF/U5MDn3skXxqiHUTIo3gBMZmBnZt1d7d7r5TCtJ0aX
hbXY+uaryyzZfee4JVVDA58t8iEgl/vjmF/DiXi64+TfBIGxcv67RQODUbYPw/qh
kC4R0oQ/G7lFt8SZlpdANH8d14u6WJ9rg6Iup6OYEXJ11ev3WdR2r4GXJ0i2rseA
f7+DtIt0tWmIvNAlYLwtvMpxTxJFfJKyaKbKfTck59UIUwkxgLZ6HT2uNIECljXt
uPns9P965kF/L8BCKDsR+Xdqgeq1tBMHuWfGPRukGFcGjzbhXaD1j91HAnNOuDW/
wsWT8XqrKNODggtlOxDlxw97fYu9/tG5buY7EBmG9Ia8fFDc0NzQNNK/HopgnBfm
IB9ASE3OhbTbfty5iur741pDWPTrOgfB41iCPItqYS8VrOXzq3QJZrksh0mD6lYX
pKAJf3FnQO0PA1ff8Vp7pKWmm/rMzfBF0tOEhSDO66lYXMQZLvOi8X6yxT5xXVah
58HAeGHJ+KPrBJPkeVeMKlxfenv7aWBtnab1cV+/BZwn8U0sd7kMJZXoVH3TcbsV
HMEbeDyv0Vtc8rqwErwrUntmRwFNBVeAK6OfXngo/omGa3Q6MTD4U7NnEj2kScMN
HOBCKNY5JJywiuIcocGSt+Oq/O22Fa950YeAyYXvdRElLOd6h8YpgXO//MUnzEJR
YPJPE4StOVmytd85MKpLCNau/Va5ZajrSxQuYrasCyCHQgF3NuovvR9+orFeyKrj
4MTET1lMUHVPhulqsyQov1O7apaAHk7IfIL7XF57sNmDjKLTogGnjlpMXmenAOHV
+n30cTymOEmrAHd/DncNPGq+/em5XtHPzlz+PAqXsI/pdoIVKfuPEcSM4MpkRJri
c6DTIr+8IpGH/1xdoCFNTF1LFMoOOWk3h92h9fYXcwyciVI38ZNSF0Mzk5XqVWQO
B+DR/W//DaXohdkOhwJ8hCJmtjD9oYuBYVzkcMQuFIzwl+jhUPRUFqb+FZSKxFVB
KtxWidUVjP+392XX59U1YDJSoTKJFviMZuDgfOPWX3NBefgi+V2TDEijepSW81Ud
dh+RjaAkHnQQTtYi7QPCtK5RmPPxrrXi6PKJNEHzhNWMB1l++tMjdF5gZ10YM2gl
1Qr5rq3rl67VY1IySXS3IBaBNv0A7hNg8Ik8n/s8k3fWxcWdagcMnJZ9IuKkraYn
RfevHinNjnKl3DB93GDMjzRuPJw9d1TUKA63sKNiPZDVoxKZrs+TTJXv7LebMyE7
B4eBuZITY2efM+FbMqSyvW92AutiE1mi6O4L0c3dXsVLZ8CBxlmQm6E7lYg3idau
lMdkbyuMUZHqWgPqTp+/L6/EUHj7gltrykkYsc4MAeUmfXyXRd2Sq8evLSITFCL/
PYX/O9sVWXk+mCZPoLNbMxcjf4T3wJ3c8AzOlvO/fEAnaRncjIhOED3g6350oOXS
niE8AGYnmU226FcIPloHqMAdkvX+Yxd4dcauw+bvhUagBzN6PyhBgPcPB0kQ8KXn
vfzWDKd7Hhzhw9pZ/2LoWi2hcN2har6xhpM9s0QMcuHfamo1SanNhuwd3wdjEWXV
+csLrSzsRMmQaAe/7S3avNsEVDNAd1KPFV+X8dfZKcCZp/jeP8oI91ZUtwgD2egp
Qo5EXA7QjGjTPNZfaABuPi+zf9ZPA5Zfb4ZPq/Yz6GIh1OFDD2h3C0PIqLTb6TfN
VFilzsA9IExqFL2KjyHXjc0+QCFztWpaWTGHsBnUC0bdQMdBvqrDAAKk8Uz9tdRD
q3OXI/d6N/JRBS5crPucy1sK7bq6sKmuU+49P33GWrEMKx4oEPop16KQXB8D8+zT
/uQsgX9/dFQmdy0j22SD3O9d+Q08UEGV4kuge8qgmHnHporl1NiosdS38KrLk6+K
f3SO+WvOpcV2/9dER+HAwiMU6LOAVyuyC0IRdOrKta8kWfvrf+K8Mi3d+mUrtLPx
NhhkmpaeCZhkkOBAOcQnrC6wKbLtylae/SpjmG+gJW3ZkFrs42rW6GQMXyHNRYFa
K0hhzQrlc7N5nuiAjdRxDU9HzvoeAMzKX92WyyD8EeI6BuPRgAPiCPjLAB/7hHlu
+oW6K67Vjhgoqv7RJNrKeKDxI1AZI7OPQthCQYeGiIadi78Pw74ZEroazYBgLYSJ
vhftQuPpc6G8POecKWm8wynyzqlge28PZuY2tX9a4SSNh8rucR8cNYU6YtgR3lyT
j3vMjGL/i81wynoXQQ29fPGbpWYIIwn7cJ7JMvn1Bp9/nKDUeEehcNuk9za5BTac
NT/ML1W9TBOPhaZVjhIV9NJB4kQPQpPKsEyFS0f1pqhJ3Xg9gOJ0l3fCEErj4VHx
80oRx0pZIJ7rdmKA+9lTbp7BMP84w5c/pl44EN9cIJLlyK8530lVQ3qm29C25HYX
gUFplF1HjtlsPZikVaI9Pw+p6EpAbmsiXT5uT+uOkMi+NrYf/NdGtNso1W/BZdEh
MvqweiDIbtLEt3DRUjB/dAZYZs8KMTSZ3Ay0MDmzctOZOfa/KuNJO/SSIhjnCPhF
4rVelOWCInCt1s661U70Lwiugf8mkQC3CU8W0wWP7Zkr1U+nepxffp+AdSSXH0Qn
GFwDyqErNeNDnW8iKTygBNA2tUxJ/YhimnU2Ax88rJa4y1NVgou68E5ET6ZWPHKE
bXjvB2WXByMi6AbnAFAc9tZvJ9awjIAzqbOS1rcdtcKRYkm3sDGZmdirrJcbCpzc
HSaVjktDdjuLd0g7FdmLek9Dp/RxXUntTs3rZN0EXjuF6soyIl2Rrof9Imi2t8eX
rkIQ6Tnw7EdGIZlVk8B9F5irlHS6GVfm3fBINw5zVdcJFK9kGShxh20zbkFP1F7N
slUJYP7nlJnB4dv6wJqQYHN/KWYxQyhwOhqq4NS46ggzfTh8s0eu7Xc1XZxGB9tp
7ZDciCD9nZhEOCmv75hGg7Omx7DFUBLH9NjHEII1Jrm34NSysHKwKhzESDRf1DiB
23ce2G7IYp/kNQhYZnWVTzcOyeA+MAXy06eH5gZQHaox/xh+0V7vLSnDMVyCa7/g
2EQ3QuNOZYUU9pfdU2XZ7fcoEB65Co99coRueNtGYj3RXvzqZCeYnaf1wWL1VUOi
Twl2QzvBTq7k74z5H2GhFIfRr0uUihKkWXujao37+GNXlngw1DbS5ayD0JdApbLB
1N1k5Z2x/AXjCtJs6fahzVLM9rlBQc0+2HaEbShqaOiUVFNlwtPeWiAXCKSZyGrd
KO5lm5y3K2dYbNCX+KT207oho0GljnVdaz5uqPYzpiMxylWxfB4wMEKIh6chMiHi
OjSOzMLHquvMpn9CZAthl8ra8xoRw9zHovKpWiUCelc6vdNheMx18Jg4NpjmnukA
MLOpdMCxI4h05TfKMHCdFqzEGfpiOmc1h+0Ea1k95w3uQ31DCrDBYL3S4UdlE/lt
7mxxrDVMWZZbLthrjpQ0QU+Z5vKwgyghEJv+UjJQjKogp2J80sTncw9wkh03O+//
mrhqhIQAmNM3kEHPqy2HmxIrmF9RDS2NIs6IrCPeuVMJStYpnr5+rcZ4Wx/xZVHK
7HoRxpAprnog29esdbaTSRrLNm66Jl+RdnZpzsI4XIwePu/U7gD+BYKsXwP1gh7F
SOQdB+D5DyjN9rbn8pbMyZYwr5M5d+OHBZ9NMGFA/gaoaroTf1hgURf8WCdpNYq+
4RwYJvzVVGnpdsjxnjuNB3fwZEsbcawySE53LdQgDaltrOqylsom3aIOZS3McSRX
UQ93Ws+8URdeRzKMjxsMrVRS+fbR/ilZJI88hCSYuXuylJHofSQ9vYTteQkqQJp8
+wYSHQxq2YOIX5jWfS2q0q0uokfjMlM0J8vsTXVustzdqLKcb8aJUHK+/6rA6Iqk
hW1R3GLlFo9A1kBDt1gq6URb4nwnlNaBTA//BFxRTz0qa8XKaihti1pWUTRKLVa8
UXWjdec+5IPiucnrE7hbfUJJyWyS6h/MDRUMd3e/xuwrf2LU2ymWUJIbRRTLQxa5
aKVGo1a3DIrKh5bDSkfXhYVtXBoa3gsrtHzviNsd99lUL9U2J4FH4y/ASKMKoskA
3a1xMpPP2Rk4UyOy9j7NDCF7kVQeBSTK7tYzqyKPePBOZ1A/C1kAwl8QZ7apZORJ
DYBhhy0MhjcNli1OaAcq8nNDdGJTf1EiOqa/S3Oho6EonWs4vbjZ6WvKKrLVRifR
GbjKgPFOLR2f8qbxfw9UH0kqPrjBOYXK3eDvh+acryHMt1VB1+wLiHls8D4lNU/G
pI4xjLP4vljvczKYTG8xqY2nrALVetbXsuVj239vcqa3vuqgnYOy5/zqaWcrV61R
RmKIj2Lx8kdER+cRWfqY1WcydXwzZaZK5Vx/tiRngKVIr3mK309jwe8oZMiTcLhi
xi39hpXNSOT7TqFH6QF5fa9n/srW1qrVTqKEDO4MArAnH3tCD4eZyiV+VCWlyb5B
T7Z5S1I2lXsCpYueffsBG1KqBSyzk404IzA10E3b1DvIZ5SuklA8BOf/f3O2h7qI
oGHQfuQrERGmQBSJSO45DAQZ9x/m6xbTq6aPdyz5VRgFT4ofqo1aenTlIyJZZ82a
EzTSZ1qh7b6e50xfUnb12i+RM/hhCyRZIeBwlIgIUsnlY13WkSOeNsE6AlqCxtOh
xP5F3t85Yv3jBrgMy8Tr1qYIne1udrZLk0fSK431FPLDWYEVf0iIt+cwh2EnWd8G
mz790mA/l2W1Mwcbhh3mFquNNNcsK6cdTu8IeQmo7HB3cEMS4gzXsVwA/2RpV093
vGaNccwNQKGP5sKdDuk44+lK27dqDuFBZL5lMfjDdL0+3vWYpu+PxvoAneSvVdDt
Oo4sBUEhbIQFUeQyR+AJqIhoKxfJviXvbmTuCaLSX17ZabylyFbraP2yyuPIajyg
LvkOfnf8zm3w9HazJserety/RKgSlTEUOA1SQ/gBBUgPNl1XfQLwg95rdwcqdZtw
H+KILp22NuqNlLob5zznQ6WbEXl1m9aZRaLdnRtC31WvIRv2GbG6Jcpx2X2adc0l
WX9V9HTVhnbkiNLHrVVVrgFwyslp8hUBRvlXDyaJilKuwmel98K/BgP4C3I5tC5S
XN27b1dwiVXicMonLeNl52AZAF23ZtX46zAjkBeUt6UkAvws+hKEvssRx58nbz5h
Rr5JosZBYPosMrxqQXoKTR8rf45K1oXRZQ3sPlRFsjhsgrfcKBvuDkDwfTS8Hmkv
L+K9o7qX1X4fBULtZJ2i972gr16BO0woL8CPzfoV9WzSblpkhJj2+e7q0ocxyGT8
iJ4v+uKKJ3qxBI6GBNhNZ5diCxdXVIucFeSnxNwoL72UJCDDtMme4ywNRTA54e57
0/VeZAz7HBr50PEkF9Hq0QMuX621owns/FQtKtzj8NTSPpqouYm/T8dGxcLc5ADU
43qqrce28+H5UbSsGmb14vx7FfneFr5hUzh0AQE9r/tXKZvtJfpb9i1y2Tm+kALE
UshB8ILtYyfn56MTkVD/Ptu7IU1ZbXCCPSXNLet/vaTeqAg8xatZP4epU43S33m6
cRUjl4W2EZkwCN2Bs3bBGkdJG4AxbIEqOfyCRmoQgpeWi9vFQAh44HWXFyTEfXTk
U15KDbfs70NzmZ5kctot88ibGCClJ51CCdopZi6nKDLdbebcTyx/hcQpIUBQvsZK
U/M/PrIV4LCFzrKbqwzUbHVxCUtYCpamJVvFMN0gnctl7qH9jxM7TuWviupM43xD
uCLdRg3Kk2qcpI0CLmhb/BHkOL21DDro3z8Zzn76OfpZWvqujZ5eRQ0Ac8Yt7CNz
CoBJ3AWy+gNn4OfL7yNnR7ydSG7JOqhe81zuS2bR3SXnNxojnutDKxo1rByhiTAb
HBi/3Kzgfwq6I5BxLpfpRSlJ4YWniMto65ztLBCL7SOWtxt8C5l05Y7JMLWf+H+Q
Y1kjMb1hjseBVy2CFXgmVhcX2SDlz8BAOmZ7/i20Bs/qIDE9w/KTQaa8yE//mylK
MutjMa9pNL8E7aWajnwEgY5yoWu0zUBNleBRrrn70G9rB0eo5JFTGVIhDDzg7ewH
p25U0xvcTZc2WW4JN3QmTJ4rNVz82poZPTERHUOjtTD9E8yytdhngVk/22C5vwc7
qXv1hqjG19+2PcTAz9halV0vi8G1myoOW5J58H19FsBSKcHemcm0bLyOlNGKJI6A
h7cK9z4CYxFkBcB+B7UrYprvXVSSA+JM1BV681KzB9P51ZXUNcI9iEnexKx/s+rT
iNRZunt0NM7DzSHAiJIPUdJ3YPhky1nzoklf1Iy10jeT/HJT3LwXo9ATIFeu4HOw
II7VqNeDGCz3ozmi0igm8hm128y/PX5Kmly+1N6rqN2BE5M8nqnNfcEUl1LmaVTW
lfWWb/VlG2+cCfqQ/DgDs6V+fpDeUUiX1ebleNe9ZRSsnT3caJidEoR8hfK9ixT0
j+bxGKSpuxDdMBMmnoby1JCDQHkvCwl6sj7WE5OHVzvX7p6OtYbT7wHWw+laD7aK
bWXXKeIdFVJO8aw1wHx56RjDlRgwDvTH91AELPtEoiRzkhNvgLqj1ksafG82b8Qm
Kj4x8Y+KabcHUJ8dfASsXxkUKArjjYGq9qmvsZisasg8MwtSclaLnYrTro72GgpK
br2GcvJhZqCZ98qtOCqg+al2dckLwLEY7mrC00POqD+UlZoZ4bO/6KcOslEaj1TS
kBqlmABy9yvkBU3HdNmheF/Dc+8Vtby1dEJ/mxtQmHq4+sQoeWc8P30+XhtqGHEo
PCDTrvPcPKn6G+wyaJVhRzumt0XGKgiqnUT1KJ2ML14Gth+pwk28itamzDaVwjtD
fB/dfQ/U0wTcRUw4xsylQaSL8wttm5IJDiIGQSc+8eS7szttPrPJKUAIqrf+86lT
S+jftwCcCEuTl1Tk15f3yeF35F5JYt68IKifJmwRvn7XO5Mad9iF7wviwigcxEeo
IFoGsAPufCEecVXCDOwUMJd0MDpI1MBjiPw7efSnK16CvcoqLXAOv1/4ViY/KD2O
2FE3YbTzbTSa7N/s1aKQwsmBjG9CyLPipRnNZpKh6MFAV7Gesjwbc0m5dATxWQYd
JLITmC63buWlHCOoaL7xINKgfCT8mEq73gvybACGJ7Vkuzw7uDMJrTvVyXCZ9/ku
j9kufb5Z5x62UmrO/gMDBh7BtzV9GWSS+NGG68OK3hqLJ5g4sAQmZWYQfuNnGAsx
Zar10elGVtm7vZFl0li0VNoq3We7rdFHh8J4uxMB8HOxOntZ0PRycLZZwh/9CYlw
LPm0o7nxD6D4PkWqjL3Y3CXq4TDWZl/SdcLlBBIBagWesqFAZsCrSgpEXH+ihINT
dqg9woNXM2nIBMs6N8f7ed/P3omu48ktQYCcGskhaNBYQ1TbKYW0IsttKsYyHUDR
ESBNyXnPFur/SB5mjBfiM0xqgHEV6Gt2XRFfIJSgF7pP4g1o54yT1tfWUV8itmNY
iTTvx2Lk0ry1aMqz2BlI3LImgwwSre0eMoTGTvQthpTaeYtT35Js4Ccbz4oKJZF2
P+UHZ4lmCVqRbCcPFQ82K6lUcX1J/+PHORQq1UnKnyFxhGEf3R28HR31xLrnK1rP
7omijrqhldyMwF+Xy1MnFc4C0aJTqm5TOaiedXizIzJWosi/uG1X7+NdY71Hl90w
nt8wIXgchNKtZ+Vjd1F3pRs5MWWZcsFqc6oio7kCCeMYQPqPfPoOHN57izviqxMR
IngZKzAKLPpzTbkU3YtsgKZFbzaDP2J1fJzsLxTYrzx4eWdwnVryfZozor3sAIsC
HLqpfwikcQYLh8k9Tkl8hMmNNVQhzTRx+xr1klZ/TucpI2fqPmmPzecZittWyruk
C6SKCxUJx9YQt/Gr9of8RMLyF9zTD1ni8o5Sgl7qvFawE6a+01waHaiT11ekr1zW
jB52BeRCiBWwsL0SawfhUeUSIwuDufelcUuuV0kTSAgK1LWIk49pp7nMVMTIQiVM
MiQc3lHDiF/bQ+P3/IvHubqGqLaIYcqB0pUb3roByFXe/RIUURY/zLBEZnlJihIj
kW0iIAP3l7O674RwbCJc/bj/O6z0QeEOflkD0agEozGcUmgKykpEm3IpzMmW+kGv
E7EspsjTYZ2MDKjfgH8XWBvxr1BtVIURShD5bAtmt+OjPk9wzSP7YqId3wdjeOoW
OZpIPL9V8iUMEDYGXT61CLzzVl38ZJL5TJrcxSjB75K8/lTIVm9wnVy3IVFTFQQi
bzuSgL9HgD/yunUVdodJ1J9zqRcHHTrWrboF4u2r61+kw452huAGSnoLU3zqgabH
tVAMWM+sG53oFCVKPYjsg1AFXpTl6ZHfZOt47LNvKwKpa4HfYzgBhWklj7D1tIBZ
qNJgd6uAOcYt0W/d5emVBSSw8zVhrx/1T64p1tX9U4kMoTmwHm1aUV5DVsFWFyNy
4VHLMfYQA5BlWQEHOwIqxPldmmxbNXlU5HyQUkkWg3tR84kqebl9x95q//LuRSNY
z32PcUSDl2O2RVcbPPnTA5FSzfnMjNhofFhBmwJMros0ZeWSjl6zwodgC37p3UAE
YlTgiSy8DfO2aVRihEnXMjh21zx/g4bf3vTIk/5mDlLU88rwEuV1UHrRVWHgmSHC
ukvt26XNjBXLlL/Pa7sOLdc76pEhXxQGInc85n5tGmNYx0elcM0+NYOBoLx/vJAB
M6uC1KA5aomjTZOjbbDmwyGqMWIieLAODkz8dd18nWqVAVgtcqLz7+8p5CajVGEG
dVyxbzy+XQZeB35220qmP6mi5Vi2VT142N9y4qTsaRdVESnY7xXwy+Elp/6W96/3
ZU9IBdONigAW/RjoDFbWUD5Gcj+WYo/ePCfpKDHinU9rcWfa/dvgQ7j77syIMniF
09hQMmd8x5pTIv5ZG7soAT0u0zG2ZvugnFFdaQ+jPBaxRc2M0hPRua+N5b3Q/jRM
SPxkPxwtULR2Etr6ebXp6YwLoGYbMzMtc7gH4j31DDww0eBzY5Awy7PxQE5NSWf3
NO6otiIRnOvdOvbNkDyg5X+LRmcnnr7ysHUUxHFBjCj9Sv6Zxc8P3DRI4XH2EZDi
fTbll68WwbL8VfWkXZbfc+n7IBRzFDZjMDK9Rj0p9h/KUhuFQFJbj+dLQOX98OEc
Pp5XsDpWHzrhfmUBmrSqU+Jr8ROnAebvYhdlSI1hCuzQZsQ9fzUwGJEU0vP5Kq4u
tRWgY1Wtg+Jf8B6IK1SskQGT+KGR9L0rkDosTKqfG/cf1xhrV1gTi7geeSOMG6L/
Tj6BFr23j2ku6mxvzVl08xsdWUs8Aht7G37Xa74AHEIHHgf1zCfFatLaTlJf9NxH
kkVpPM3xdrHrbjA/NkqcLhP0GXLaSh3+ItRxoGt5lDtn0cvrcam5TylXqKcPgS9S
U8QQPl69yN24drFdpt256IYEtl6si1EsSgwGG/OuI8Omj7PUWQ+XGe8gSzr3r2F0
Ouaae7mURL9IWUXcIPtqn/327JvBMLpegIFANYmExRjNtzOhT5bB4RNquYMdWpu4
QvF/QXXlgpN9bsF/LTJCSVD5AB/fSCkaXW9zUHz56acf1JSUqw4TCDcAezn59uyk
3iYLAgn17cldJ5CHK7czsHBHmxKRUOBSKYDeZ1oNciao9DBF7G+09m7z2wh1ARNT
ETC38FS+JlfjEtSqx+TC6HuTbqloKy5cXp2nnrhkYVVzXNADAZb/48+OKoBIi8j6
5qLncX70FLcQMSgc3N6vhQta+xJU/vBQOM/DkKIsIAp3ZwBc8sP7doeBqPH0mmvc
ZRQjz+ChNt0IN0o3qMjdgilwpWXMWzzoF6PleDs/6FBnGKG7uccUB40qJ4hgu4an
jhaFDksA+w8TQ/J1La3THoATaXbH0qK1AU1/BD/38AYaRiyAJKOeklpygryMsEDX
FcoCvq55bRhQEyGG4mO9hR46HNQSeDQYwHz+FcDGINdVR3xO69C1fDM/9z2KUy8H
d25f6bMO1zeTyycOnbmGFvs9NwU2oYQwpHwBuFE2w34Q3Zeoc0HADAj3z0bN0TJM
fHPs0xpZVGQ2ULpZc+wpKcq92vgdifr2gQuIVewlUmGNYog02y/CwoO67Naozy+V
SL4dIfz0EDY4GOdDh7GUEUik6D1oiTLFdcpJg19M3bV+Ps456cibCrINzKgt3Pu5
Qq/JMry7YzU3T+sMOrRwNNRXBNRlaz5SK3dQQaN2h8G1ziAUGgJfR/BL8AbJnYNC
8EhxA1e6tAb6vOgKbNlxL0zKQCVcA7iTpfsAjSWTqdf9Z4prc4bIEb6pdhA92tc/
uneql28Tn8lf6rfA6GOrG0rGcvX9cJilQLbVfIk+/N55P9JlHPVuC9nXpPV+TqTF
gVlSTvlLjHilXOn2GmBoryOaa0jTX+hECDBSy/pAMksAtDG1OCwqDt5sV8c8STZo
qZbIrBWDhMHEYb5fkqIWqbMfbFDTluwmEksQhsmLG/0zG/cdZb6zSAGnspLMR1Lm
WQXFYoEVl1LblIZtEE5FdSswTwW3o0wGtjX+/Vh+CmynuSJ9/s80Zm5ta4KK1lAD
t0IFCVk07ustdssItiYfiaFmndd1OD3ecJPDaQVMKk3U1izlVjBi7f+y/sME9UTU
0dT0DLU+JRFKjiLCVoBk+wO/pD3r4AeV1W4WnZVZTVhXF/EjeX94mHQXpTVhDKeV
SSO9IWWgfkHcQGwZbaRS3irelvrDaXjuYFnkxK9NaR8TexWh76502iG16G0NkEwK
aZ74KxxGzkvdnOnlGJQ7F4jizQw85NhevsPEC3ySqpcSHnKvbjNWiHEQs2oOKN5l
/vR99RYpJ9VWOerAP98weUfzuHHDfQ3jJmNbE4/11NxlECHFY0IYUF9iP2t4FDiB
i2TT5lsMEEEqGLoO/ZVbFb7VJ9u3oJnVGJ5J3tG2ToinXILP4hP5KK0YI5uJ0tJb
aCJqmgkbumEEDBA1siBAaxr2UlmoBR4R7/IiwiTGZm6KHZd5N12AIF8azyVCZagS
57+v96TlMjeOyhc0lptAYla44/sPwI8FY5f150FJuTSGBNDN+PTe/y1/5mgK/rF2
g+Pxvvw/wQvvqLu4Q/YSBdSEx0kCSSL8ouqVRMOgUeSec6iIyp4X0X9PIAZ+AYyK
kovbij9SRv76emT7IeK6c5S81vVPGOeA2MaIZlMObQHsDM4bnugvuwdyr3lL6Yus
WsoCp4st9KFqQx81AI8ZQEqUmlA6mCXmnu0Ikgg1+3bJRj3UCKk8xSl9QhP0wbzC
b/OijIo/z7jB8PoCVmqggwOwmuur8oKwB2mM9+g2wRoblf1h7jx7WWqE2JedXVGL
fcInSBBJNcmw1yknGpotlM0K+7uzXIYmBCEg57/UUQWdv321dMHo0NL9aLaBOrRs
1YL4j/32d0zJYDkrb9P8kEXmnBNTJ14I9JGVBKFf6JMhcFv06k56F0xPbtn5LNlI
ekLm/FNG6WAqiDEuFVwF0R/VE3NNWjRpQn74jdwSy4n54w315Ra9SjUEut4urm9j
XsRZmiAHLJSm//B6e07Drx+oOh9Sznn1Vhw19LZUuVSNdH2zEbF5120Xpc/kHjAq
4eANi7U2r97/iC9gcN7sZWZ1W1/0eBBMR+Q6VJs/u6fgHuqAx1WtQhh+7aL0OipE
cNZO4ETtYOpvbQMB1l2LkVcbRa7K4NiJh06AJSuUZta7CGSmt9ByntNK4bVQcTIs
yA9WAnch0P6n2JJn/zNTXM+p47IPeMKTXs0o3hkI+O3rDVv5kjW8ov0dWDXa4+RJ
TNFDtzx0QbdIcfg9U6a3wZ0+kTUmrMuetOoZJl+iMSZ6kREK3mUSDQlM1EOIpXmB
r8m0uxR2DuX1H+9kSAXJ9K5MTfKcWVng5oGcUprJndX8OIcS65cZPiJvuBY6bePq
lpUg55XGdfpPaxPvPKcB2ir/VPfprOVifD2rFZynsrV5ToZLhonwbpkamRIpyz3N
tEib/NdZBnrclj3TEkdVxhuirSbzjoH6osL2L+MdOL1GW/kjeyfHBVuj1WwnyUSy
TMDqCdyeH0Q3m9IzJ2wz9O02tizWiXsvCSeQiCktz66zVFchbFxTaDiLEAwwfdzW
u+8YVMfv0/+d+5ZoSNJ77s8Ll5DihtlketfMfrclYf6EHUCLZzEuAvZxkHGn3RqM
5Cf59Qd9tJ/CNRiYrh1sr9aRFTzoAxV6txPKF1iuY2SBhRWY58Y83gzIUXRKT4lt
jLpecTK3WEmT89I5My4DYkSHQTsxt0BeG/Vo8sDGzvC5TcFPbObVd78dNfJojq5W
qkgOMLg6MQQSg0g+JUMxTPpwU44Q1c/1Ei0orgLxbNjdsXD7y7BhuZ49/aeSdTuK
VsgGKT+Mn6kJDkHOy4v24ICwGTExHgNJb7dm4l5zo7RD+24CMUZsEBA6ZZXGY36k
XiCP2/QyZoSG2WjyJ5QyBp2NauI0ufX5gNsYKZEqBfo5yUzJhxXh/B4YU4CwS0mq
pOYSTfXCR2QmqoD8zPq4itfdjgYhorb3vEzmHCW+JZ8VXRzgGm87sxjlzl4CjgaS
hQVepBKvF6b7qiMkSSLJig8Jl0Jmk9SvahHGM5V251/0dZvo9aGBPL+roW96TzlG
mIjHlhJU49OiHE5fmiNs7riHeJG8fML8R7FtmTvqPeupn6vOJ2NR8TXEfE6NX9tt
LGOd6rYl3ON+tnViE7vM6CUwzrAxm4bqiLsWtraKFuVb8PFHFWm1HOp1CBKZoYl2
rjeRWjxCBex5fwoew5HhCZrZT+xp2zeBft/q95IfVEmssgjnv8fPOa5a3iP3ngB3
GfGIhxXHZWdT5ioOm1YKGlfh1b53oOzC+fAth8U4uP9UkxVDZm/cUJ5cZfB0OpTY
Ab797j8K9QjYL9rXLSuHlSgVeNWuRkgTpwEHDUKkvoh+wL2+LB2n22fG4XUxK7L2
0ee7RNjpEYMUqrt/X2tolh0tiC+Ip0qotYBng8ufZX4aW5kXKXnDge1YxKd3FqHC
5iUkAawCo6XEBlBIJb7zixCgiT3OYr/J4vsJhHChvwTofZ3Jq+bpdW6AT4+xXAV9
I5JFI7YW7EdvzdUAqQXbfA/pZVez/EFrE8A4OL96GqnPcVeL0n+oe2YmQ4etapfb
cU8GQtCM5fz0bajhSO0A+cOmJaZnBGu+98kmmGQR3TThj8Arzx66JjgR837ge7TH
zP7/3/ATSjA6MIXTop66WINrbMt5iPEBqNywXoqGc/TXvFGFJCLA2eJWAUUMS/IH
vfLhuTbOWOfXpfjJIQ/VQw/VjLNJgKN29gT5CCjGKE0Qz/lQ2kKsS3zGh7vUWgfo
td4jxhbasznZFMQpyxzIrplXOa+g4s60KwAopgPbDu77UIVo110sLZRyr2Zc2yS+
EIm6+QZHyou0OqfjY998bbYpkeZT/R4lZzUFMj7DaRM7TaG/USAM4V1lGjTaupzA
9h99vL6jdcmsuL27spK9cw068uOoD2TThP65v9sZEv5+k/wAI6Qwo5AvgVJgUef1
VIY5MIZn/IiEOvZu3jMBE399OsQBY+q7xuid79jqVtuDsyYcteyB8d+kWSFM9pae
270GIN2CiGUSii+06uLPrOUxTC3FTbSPNOy+Y6pmQsQBbw/6bXDLSL/7n9MWxdoi
3+QG9D3CklFRdWaw4shykj8z6Fy0eKWSM66HUKpL4QP52C2zowGDvG50bwdvJWPi
Cy/Q779X215P2dP951NIBW/2rNulEJ0ma/FhgGK+cubPkYx3O+iaGawi56XhGlJx
Flc1LUR1v/sl0RvFWs8Wonhgm8O7So/sj/XMuKbkvKHwEPSZAFC4QeKYxTF+863T
JVSlk3j++r9Zq+Xfv+v1C2DIcCQgWfAk/tu/vVvK/LSFq3f1hGXT336iz9/+jtW3
CegWLOe0Nnhk0pGyfO99MjRrPi/4YZ9tit+2TL+GoxBGuBaEM0ipwNybSB0wY82h
MocPpZ0CN7BsaOYw2EaQ1JTlD7F5HPZwO63vvQ6l3BXNs+H/KXpyL2J+bLjeIahA
+sgzHFe708CEfXVA5bPcEcy2STAGBKc+X6JgeB9zUIJAnxQ3+gm0aBIsna+rXFZf
SNRqFd55XZDCuTgcrsOUMoohBO36PvvDHv3FVnav8M4fCdDbMxAqRTVP3OCOywZD
DRfqke8eOj9lP3uoaMfO2pb+NpMM3yms6xfYm/xex+FNkUuo0JwivoUUc9a4jncC
Azmn9oye8YR4PHIhiG3OjrKjbGbHqCrAozBV8RprqbY97oEfxVwG/fMA+SYx2atr
k2Gddml67SjWUj/MwVDfbsRa8rTWC8seC3bWxsJvwReOjHp48BYBr0Ku67oXbsax
bElTjdUOSWje1Fm5A8uWbp8SDfG9Vrwt5PGhYLD+vHTZITxPfo1wS66Tj09V7bBj
bx1fYXNe2AX4O5mCVDu6BypZcXha06IONM0vncClh/frysiPcK95ApFWlrxCKypn
z5+/0nKHJd1YSE/x+59OIUI6oALnzsDuH/oKYjZGIB9I4cGmYYmN2xN+7M1NqH4w
xLEsm8PDFlfjIpThKc/xknRNEi6sH15y1YWL+FAYc+dhI3O6FIUz6DwjXnfMz214
P/g+xv03buTlOX9T4XQ5dPz33R7J/dXHmieXOe+91VViGXAl56VneH2KIWGj5BcS
5Z5YwMQ1nV4uCOoYQH3XPwZCWP5gyRh1sr9saWtK6DAEpCpKEXNNmTpIiLk9TYUk
v0zCQzSqgbrT5nZlDnL2k7rxb86zGX1jWn+EhEekJeXNwihtKCohdk1WGBmmU1y/
llvg+ujO7E59umvHR92tIOEmTpP6g1XTCr4u6Dznzx6dMfvY4FIEyKK5ZZjG9055
q02LLcrgOoguS+PwTP1lEoNQbw32aFb+xg/lpvSuGv4NPkA2JfWKOW6wpRz29bNY
Mzx9e3qK3OYlSmLCfPQWPhbXzYInXuaoKbAnVF1duahTLK4AwLu9IlKXDquYnAG0
LlCU58QB2ojvyt0yHsstMzXo+jdoHzrgoPxve+lmKZ1TQlsOTfWJE0fX5gIsi7bB
8jSNvZHtpha0NNMJ0T3t7pVutBRwzPXi3Pd5xf8B/a73eJwVP7JUDp7XjSuFzGYw
Hg9JPOkm22t0kfS3cb5AS4Hz36Lh5+6U6fFHrH/w26fouNqYdaEIA8bIbjNcZBKF
lhrTsL6EkQFwkLx27fO2Jl7YUKM8w9j7kmun2env+1OFlDAsI2lZYOivCxD/YJEz
8WNEinPfmJUJ6AAHvN7giq3ogZYIZrW7rOo6Ke6XGiRZL00LeWY4eUdpS7Dbif2O
R8ypHbs4KSq7EC2QFsDOThrMVzNNCCTx+8OPBEcl/fRjWpIfznYKv68wXckAimAa
efVuwF/uLKNNH47MTqGi8poenqbzSp7/FtiPMji9MOvENbtNvwKzE0dkhtN+7b5R
aQTvgwQDxBOqac63Oc3CcaYTcF3bLeVU2GmQx8pTPnn4aj2TTOkfuTlXBzW0lhsX
fAoEixDr28b5FstCf6rBlNND7cKiC9XpUHkICs2gPPxLiHBFuIVc3Ma7OZJod3+5
zonbqDQdVR0RkLcWTewwcHrnI8SagnyeVNBWG+HAyBQtvRjLwnKADml6hyOqXNf4
E4Cy8xzMXgTzNA+moUAp3AexoJHNBMUW7a0KOtYBpQf2ZdFR3nyXGXstakZeLlbX
IJrWzmSr8ugyZdRU9ca4oEtnpcJli6QtcKvS8+iZ6tSBO/MEDPU2jGvNiTq2u3Uo
R/P4pcOAJ2tW3FRU5TLG6QyZsQ21sS1xQcEf1UZWavK85IcJWvwI7JzYdRc0lXaG
clUUbIBCk1fS2ZOM3nlV/lhjEAwLCVKRsQ1JAMj99WjJ4CNnLe75YFcNxMLBRBE9
j6oBidLX3BrWPyAe8wIJzm/h+iidr6GBIkbXiaaluOBztIbwMC11AUF2yDdJvtBT
V2zC4T1nsTz6eYP3SoRJ4+BxBTuWHyV11OJP//bwPsAxSLKcclpyCUTdiMDVkVcn
lJJsGpFfCu/jlKdJE8khrNZXnePjI7WW4LjnwVVUE+HbwfIrsJoTt5rM6xOqQbBk
2sOBsMWNDvrKemqJL1e/yIn6gneNgFZYd+Ie1uob0MeLa/khFYg6mdai/EZzO//Q
FWMRhM/HqhiZnzHZQApMS/TbynnWvtVPBkUjDT0obmOUuxQwJZ7pdYHMuOquBc7i
b2u0XpyLilcr1tac0ooW08nkPwTeoqxTTA/CWqq7AruVNvhYhvWX9wG2LywPisln
fHvv8hpc1NvG8rpfadd59dOpl0fqh38OxnkSp4wsNB1byiAPUjwY4zgTG9yNyxvA
GIB59iuy8WJcWkgXgeraj5K5IfwWftm13VxEo5jcPBQoC6vYn/Kt72zdPvt9dfKb
LFsoyS5kGFXB93bmZwC7ZzQW9+Ahnjwq8QqdJ3gib8vD45fIwbwOZ7AeZkgzxbpa
HOR6uBOctzgnetmvUx4TOwUNLvpnIBmTxx3wbWKNIno/uDzpG9HxbQV5oFyrKm/9
JwHjM28JTv6REcXb3ituntRP0QH9tkhFerjFO3eFI+vou6AuY++b5uVxAkgJ4us9
W2jMYio+SL3v3QueA5WuMTOGTQ6wA87GyxAwaLhhU5BBSZjyPPSPKb3PbP3bL73z
drITFgEFmmlnW1Wc+mxU+RJZoTU4xdXfiTyzUWA6Ll96wQHNlwX8sJLXneTmp7+9
jwosbk0f4SdRSRMdT0g+uJP0tccGxF+eXjpEETvk0p6CrREyYiy4WMAmRpY3XX7u
1PMWnDJZxej8DKPwdCgGLJjXvqN5hRlQT2YF0j5oGqSmyIDV6vXp2hfjN/Z7Xht/
3puHXkn5F0hHB+EtUGK9/VSs0c9fdZEArbE80ETiqlShzbtZ0q9kva1FW9jUfPrA
lTodBloxblLWTdNLEKfJq+fkc/iVBVtBEhQyzbUrVUn59b4NsAy3WqbUudIDRn/s
f9TAr4BQ7Qbgc9+5TOwg1LW8ALK1I+C9kVNzAp2a62XfMZ0Uu0cBB3DzEfCW7WA4
DUkKJVLDkOmg0tZtVHgdDRo5oQTZsjdzM/03D0lJIpU4x7yCIBxAtYFLUgZctgej
gJkI0lOGPcWHcPOF1hB7NlU7WMGfCZAEeUexNqlzGUsnVGv15lOS67eU+VTfbW02
N+xkkcqcw4dNzeuUTEo//xbVC40k3TeHeA8fzPzA3Dm1Tvw38WBthNNrpdXipGGx
gIlQAeBEppOHbPo8Fo95QvigFoNi/7KbspvA1BHp58uiAHiJgcgJBzqzGAQWpIaW
HpNmBezKPRfyy+dgNkLW5jgw9f6YFhcBaO2g1S2wmVmVL45Cvwt4ajeOIpjvLGKX
lhwHvaP8QY9L8igGFu8P0gzUak2KPcfFtMrtQekLRpf7LsTD+TvCk7GUbz/gYluP
JLdIHm+1Pkx2UJna48a9tuN1wzBgZ5NZ55fDKzP23T55/yz5/En7TAWVmgETiQ/h
V0Qz9bJwTtBdqSNW+9g8SBrE7yLKGbb2MUL/j5l9NDEjm6LNBu/Rt8UO84LUQtpE
4S5kzIA1j91dc8Te/waaHwsDAcbAv9Qhh6T/aK6Q564Pb81HL/PQbTS0JUF2JUyY
xwIeL71oMYarJhWRzZ5Nj3IQBBOO6yEuT02kdA5Oq+TVcXyHdXcg0Z9Xe/h87D9M
Kz8cRwwD4MgYHo9sD6kx53u6+4ObsIImjuN6y4UeOzU+fQTd1Z6pgo0WNin/b8Xx
P/Kp9DfcipfBJ8/RgA6io7ep0t64tqbaVxFs9twJ0aL2FysiTxpWR7Epo400J5BW
4If5jOY3H8fJ1P/aWsCUEbQ4BmwePQ/eG6WBnmojXSlno/d+eSyNr5MgKoPcqc2u
Z/jpEwUX+fsEqHhilHvIewdoC42ck1+ykSqX/m3VY2R1XUIZJb4YxfnSS0kXnEA+
b+4a5J/D+Q392tEkGWT11hgYFOGkU5DbK4TvAqBvxRHF/56egcba0BIl5gjTMw8T
yWx9S4bAku36W0631Wl5OIHgIhOBX5MFZ6wM71Q1JaarbOMEH/PK6qt9Xar8DQQz
63R6HqryBOM8OSX/mkTNrCoBGMaPHN7yTIUESVhA6+Yl1UoJdirAar/qkHCc86kp
svyiUsX/5Uj4cqOilv7kMDLhQra+ttxLAQnnvpR1EUgaUqX4xNVfNYr2/w4KxDtF
a1tl2XdrccJZ0SHkUjWJ/LqkjO8exHEa3QO8Pz2DX1WXi7QeeChX00xAtk642FvK
7FbCBIeHWkDA4NnzvR45FRYCyLB8SDOtc6vqMBm0gyuDirAbg1D1Ge0qpgBRMc5N
MPhHU6uSL+T5cZKkyX5pPvrkamjoR8QFYThvVVUm6ZZ1ACz8Y2dmAPqu4RE0OzbD
JOlSrbSkjqKwVRtQNq0ppC3+2zoFki3Fnn4Y+q2ahRMvZY6qrwsCgdaKWzVwdlGQ
3hdjCXDcqXSOd+zgccHqlvvLQ3uAqgM/7wuyw0izYyg7YfrDqNdwg5chSa0SrKTy
UXbbTiL1HIakXAt2uyJ4Fz29bPzTGOqF217XN5kI3PmcRRMSVrZcsoIcQD0A53+w
ebcy/xEzETH3nS0KjJq7A0E6Gaz5U7BqBaDaoQIB9U9UPI0HZvzkAaDGcxZeqySd
rJVYn8HnCFTRoDTeqk5WpnJOSFcIqf+LiLxMNuyxYZ1HzGnlPuzn106jTwKE5pRQ
XYLZYxSVHRo1MmEmKtfUYO47IEULATrE9w8Mjq1RaggXchr46wn8nRzaEIC5iDa7
1yiRly/cKqelGB0GWqRoEFLnZkXzg687ioz0YJH6pZtaRTdP98iuk9Zozlf4QD/I
9E3dvzvHw+z+8YEDTVm7WjjeTTfAWaFffPte8qj9HpkDz6b0IR1dy75tp68+cc/3
slbFxlXr/NWbvcXBxc4brngQEXqfenAj3TaJVIK6Zk+l0khnledT5LXHOJexyEK6
JG9kDKwvNcSDkK8bcv3xNrqVC/Ucz7I5QCUsfDlvoh4y7P2/oHkNEJuxtvRhsUPv
O2OKbmUXcBA5+cwRp91W6g1YnBrKZ6IJzzAtvvmUcok1rnMLb2rhtl7ZPwxzRbeF
WiIc9BcQeoQBeFpgQRwu8BWYuvKL2HWLY4f8u7kImHcJkHGgwW/chxd70KH611ut
2OMmCQtVKERux4/m9iAWjRJCPx4W+sjJBwoQYEXu9BybVLIb4URRs5s2Cr4dIJU9
ftoTwNl64JMbTLAgwVE8NlFC9pEV9/hh9WEjzumES1sP4EMkB2S6YkifgpP52AEu
5p/8zBjCngw/FEcO4wWtaTHhzU8zIzad3eRux1UETCIwZhKBeZAPWgg5M4GcPxPS
NOnG2zZzwUapSmQmntV2+A77A14SghoEW4bF1LXSAbgU5FWKkQ1Rm5Iv2z0QqNkb
TBmw5s1LmUaH6xLmHBImjnHchrVGCvgRKtcVp0Kx2vvGg2miGvAo66tYWefe+HuF
YkszX02G+TcoeSzX5xGIyG9+SAZ+3Zb7Pbzs4MUFJjU27vxZInmfnpt2z2m/38nv
4d/eTYXwMBRVkio1CZXFGkkpCTvIotYADQWaTMqfFo4cCbCe6HxQvm9Nfa0n74YR
pNncvKS3/DA6igj1pZr1VVdOdeELwB7aroDQiVvx1EGyDPrWmMWJnDyg5uSZCkTV
u+dNya3lIZxmyWi3mTzNVl2QQI2lXQDuMxeXkIDCSl1jlU9p/eq/VbrjgR3VI79I
lGj+Ep/WYAaUJxrcHd2kC0VSMfsug5kGn7gpXWehSCE5tPgeurtDmqkwd7+sN4Yj
onqzZMnTLaOBIM3pfDyeGEzCxG1MPfAhW+9BydxxefbvcramBuG9bOZoovaOgRaR
MboPcN5U2TjoO3/9/qAgbgjqmFPcZBxGwtzEonqrmMWptZV3AcYCv3ZKC6c2Uf4z
sNeInvo9wA6Q3mm2ZMtiJhOJvyNVHhO/iOJabmOh0RPEQErQUMbzvlMbysJvDDuQ
+uB7vVjyA3S8ewUH1YPJXzhLeOPteKg7I6sEDH/XJjtwIRazztOXqNHhyJeJrmqh
S42aGCFDaWaZh2ZSMh8farmdMXnyJhXSvfJgUz+TAkeEogHI+FnEWPBlO9vQLOQv
WTR3oYdmAL2+hg+gn6zHQkFR0RS5ZRNslMp2I+2EwHj92dgyIwyqWZX2UADrIt/x
/96Hu+9iLowL+kZK9wbx0oObBHYPHphOURQRbAtInpIIWbLqTSlA6PMgm13BADKE
NpEYGBcfOUFdIC0uPUbK2/YSqg9fJMFCgPaiJwbUt/PwZeopi7wlzNerWiXoAVAa
WmQHAJdlyo0mv0lnyOuiXrjgUTusA3hOYNxrMTfyZs21ic0W3l/FM0uneWzRnhYO
si8YOPNoQg2SCyg/a2ayWXTuvXKarM0pSoFAF09LkeOoUr2jqTZ0aDapavYmrN7H
astpxYbLUd3CSBselLEv75DqbYalxGUdf72sVXylO9QnpThTskMi5YogR7+/gL0+
euZQ5LitzbWTPmJpxxzV9s0VqPhWkActcSMYeVybODxDYKnhX9DA7FnMHVJRbJdM
Ty+nw9gu16+h7FrpjUaXCN7QhSjNKrl+/9n2m9ylVyTcd+3InJ/+ypkh4DpPpM4W
/PuiWB/fcnS08QQsBdRQDKKUnPmnXgCg5/KigW8N9w+72xEe9UhtU+p7qIrYA42K
NW78SkgmzORa2IUnsQzjk8C2z0yl7Q76L57y7hlDBr+0ozOPfCxImgxoR2x1Ec9l
desq5CNT+ty1CYNl2c03qBNu2RSf+MZ+3KvGTlT8lsQO8UrpYgRCvztEAEfE1jC9
lj8fk8bvxfcTrxAuFp8Yy9Eep53qbIdEZpPnazn+LF1Dgh3Eazv62BXHci5FWAM+
LgUcZlib662Wc05To4dqL3LXdNkvT/CD+6ZHiKwoXdTNBycrNjWT5dCy6+z4ZS5t
YdktGVqTVmLlNXI2O+1diKBQP9TZjLWztj9MuZSiFXiSZKnoeGs9m3wIp+GregXq
hINKiZenxyDf9f7+mZoaxDch5tDLPCeI1tsWb+5amvtreg8IsXsKyNsww9i26zwj
I3Pa7v8g/C09FOmQxyqCaM3bN42j9ut1hjhZW2EXqd7U/0ZUFwHbZODBDP7XuA9T
JGr3Z3il1QyPf5GpPXWnf4WIdn7XUgIq8qSrvNutEcf6lNtJ88pQzF8vBiklO3dS
pJxCW3Y07PnaVPIoH9kqEwcqkUZWcunVK/tOIVbmOrsoH8H0tG+6zmIb+fbP6+5M
NjFcEu0JO7YwofvwqRHdFsrxN+PA99kb/ihKG0LUKAVJEjummUT7QSE/TkLc6Mql
LX341BXDyEz3rkvEjPR/N8wBK8aYjJcrHRd5VWilK+dKG5hemvk5Go5OElNG2P1O
bG9/pxstNUjAYGR3rehpCdd7i8PBOBk9uRydVS6zzVdiI9CPPu7SrJ+eWkil3gbM
ETscgX3FaibNtRPtk/Ue/R2qQrr45MiZ3qwRELoyeHs5HFlMuW8oyEFm4d76fDGO
xvb8Oe5nc94zRjs1l+ItxEhpEjT8k1db1VdWXTu7bBsvyqkW4lUKBTN3y41n874o
M39e+y2gVfmhhaszhpMJtOsqVc/NFIZFShgvr+oxW3P9/n6eXgYt8O1K9cureYX/
oXV/i074GJv3oxd1FSOLA+7jH+KYn0Y5sc95Rqal3Us/KXTMcmZaUjq/CJR8AwYA
LdDIXoMKcD/kjn945wNkHb2ajAk9TbF3kmEREsZnK7QBic6jQz3Iwxt3meDB5Gie
JKy00Eo8rBfsVadiTFYmGHs1zoY1TXtIEgXE9LzuUN4xwqQCNfoFZ3ioOf/wqMPb
TOMTBjohxKervwpV5R3jJv1jk1vOJr88GukGM3vsEdesMiWkdW/Yf1Hk+pIzbTQd
M+UflblmxDRV90CPR7LCZUHgfla4tJmRwn8eScB3/URumWfqu2es2Rz+dvNm91em
7QhF1lLa4Xc1c9Qasau64pEZORNRkv5+B1wxqTsnlA3c/8puXRVdth5x0QIOVIMt
fBNfPG3RC1CGphHYdPngyOszs8NC6iwFK4bG6ItMBbEQDcVmZEAC+Td1OsQ2DzZO
tp3pwNSH6Oasy03xHnglTmuHjiirqdc6lfBjhhYrNQhQNfzdTkAs4QwsSz30of62
FcKr/vbx7g9seMGlpcu+bGcopdFZV0I40kQKvaPErGoL1Ejd8WMCOkK3EQdhMtVw
4FowMxmJNnS4W1W07SvmlBLX6hQhiuahg81Mv+bM/tZFq9oRuD1vIs4gOFsEgMn1
oLzRi2V/jhfYhAC8BvVy6E0Gl6YhQHDNr62T2NhE9eqcejsk9mebCb9aEf4+7yy1
lR0xuu8o9gGgD0v8Udv/P8IgFY0ak/RpYBYZ20DT/eiV2e/SYicF8wKg37995T+G
hmqZ/ScoYbtUC5nGN2xM1Oqdc0ooOLFdPANzQAq6L7xmDjJIDjVvYvjWatd6/T4/
XKTkxdgdI2A006qGaXZLzs0WbwiiqW9l6/CzKmeltnNU9xODCWKc/dAcLkFg+e4W
0BijP9108Ld+vmQvnW6C5flXIu/SzDSYkY4doVvdS5veUAyOiAcgUzzyUXilGe1u
KckhboLl1nFg94QDEcFbx2QHhKqUah//jSWvmE8AmGq3LYgP+sWbFlju8+HSRczK
ZibmDdBV/eanO3X4c0C38w5+Yk9KPtrDnZhrz78u7zl8Sg17FD7CO6uw+GkLMd/E
zsK0x3SYaBF6vKshQp2puHr4SbkMbcGeme6/7GpSvI4+kHy5jy+x6hoUZTZgYR0z
J6c3ZWRFk3Gzn6LTdg6wg40phu5vy+zSfSCnk+sXm2BJTPJ0k5jycx6Tls0MWBFS
klh8LMjy0+PsEdkj+4e28ifqXlY2dLVrIqK//TjvV/fBT1W3e1yfpx8OK+Z29IyB
17ahsKAi7owqwdNIpB+nf/6Nl5d8bZsoTxVuPL15SLSKduj/1oqNa6WyWFUa2G8o
Ol0nnmWzd52NeO5Y1yUkD/raQ3inrSb+ZubP3vrg/v0GNNQPg6mnUWyEA2oOsfD6
d9va7OKgJ3B29PHvWSDjpuIvacpo01TmTAjz0rBnVpXNlykCEZUPL+le+vUWyIqV
YPYJVamQJy1U1ua22qeieQiOe5oAIe5JM0w69Dkssuq1oSvj6bEqOhyG77OjKgtw
HrayHpPliTQkuwvj5mUAAzwwowFux72zbqVVpQA8p9ZCHIGglHvW9Cq/P8pzWmre
YxGQp9D/O80Vq+q5hxqqWWbbUXhCoyvywkSfrAwM38bOvDCZh90fiwip76dgsjWN
fxtEOug5+Hh/L1s0tj0DiBP1xdtCcsJagqJGIJA1yFX43w8nI5jU7sWh54pn/M6z
W09XKwrOKeogoAXG6IVdfLDirU4yg6faxy9/QowcPrTIMhd1c/mWdfeUXzmHwi1r
+ZE+BXTLrPWDHzXvOMOwnpn/Cch7gMwsFWS3Hjr7BlzFNWK0W3yGbX3xlczyKWFa
fya3vyv/Pgt5YdwA0siXj1pXDyfgsVcOUqo1O6hvJ0ivvWXUCa05LI3IHV68g9yP
jwmK17BDOlAATqIBVL/So+hVVc4gEOfh9sMZnd7xf5JDPWDzkiSfXzof/ATJAKo4
rnbOElSUnHzLzJf9rHau3heb763j1ylO6+jbIz70oewcYGoLizf6EFT47wZHuGBt
hEMPBAB41lSGk2Os8nVKB6NpWAjCT5mSBFHxsD+OXBBawPgaTfTwAfzmii9V1zWc
Izl7uZkSTnifIYxbiGkTbEiJmIO9mYqIKlIIyTv5M6euRo86q8LJaS1unU9J5rdR
isLtG5wWALFBU5p9F/90qYpJKb9Ja10ypH0bFguwDBa6PZlOdEAhlNugGHk4s+3Q
ip7CIQg2nuZDlb9lxQvbu3POFX3Ey/xC6rD3Km8BQnRgYq3clitW/K1fDBr0v/2x
bD6UPS/b1eLz0kyVSef6CEWiMJGRovMsvqcpmRFSfeNvkWF2rHqnpXkhoyZMyykr
nxWcwlS/gwGvWaDYo6NIBenRerSbdjzfHlIU0E13xIy5R/X/x5jXS6I8NtFZg3Ki
jXUOuVW9SHlCFp/JYJVuJ9d4Gw4WLWz1Kojhlhiok3tv859nYd+kgP8PzxR+P84Q
9S7GetlafUguE5Hk7ex1TjLDVzkgcDnd/Q5ptzh9kpQCVa7E04b4Kl34DFJr0dYV
lVHG8S/cj3lVYKiIqWtz9p91lkDwLCgpI6N7ae3Tb3efGxUuQn70WEaScBD2Dj2+
XGvyGW0aZLwltol46ut0wIChyBq9bifQZ+G7acwitE5OVpNdoK55kTkfbxb5Jb2B
pcyvLhUwyXTSjgNbxLJV1frgdLt7D601itXDJXNxz0n9XLY62zH8wbNazZioqjGB
g0cvBrbhopud4TNvslCYOwk6fRqQcZCuoPXnqDBI9eglCAbc6An8+/0EpFETMBv3
0aQ+W7JXf2tTLjkDr8ZBVsiYNCaxkeDTbObse3d2JsD+ASqaYHnt91hxiKZKIuSj
ewP9fdhojlw8gPCk6ygSNg6IKDtcl6WgwSpSlDpQTaNygQACz7zVFSRrbr0+zbXx
M0xFAFwiac+g0CZ5zYWJLAO5OemrQu3qvoghRF/97IBp8QuEMVqXeUOKHa8RIkV4
MIP+uPJTV6Y82zn+96C7Pu6JWh4RqU3/mrRfZNK7pcvBgdb5i/+/sz+UihQEEEw8
T28N6BhuI+vcASdy47jwWJTKjGTD9+Eurl//iZkmfwloyv3M7ZXB1WCFYMdYJUIj
WuDubd89sAOQlHv2HKFhdv7FI5fPZRQ7pmuSyFw7a2MLwmvFQfHP+uqKkaB0Zbym
MSfHbWssFE87lwyi7pjwwKDPZBxCCiTj1qmIl8oZP28pRHIjuEP6NSa2f7LDfB6l
KiVXpXJeTUxDUm9P85w7dc5VhlaqvNefrJqHWLnQf4JWpjG1bXNTo0DpZQmzHjMZ
5fTd+7Sl1VWRfijLa31ZODlmI+7/AdfWxjQuyv7kEZ2YS7KwiEEGkvXvFFWFAmVB
UvctI6qMQJVZPXuHvphUdRDuLc7aw1LujzN00NmS/y6B2PsTrbbvHx6kDX3QdAJo
O24lAsh2WkabDWNErUk6Ukpv4J4Jn/RXAJooTMq5rpa3fuLbh9ETURkTW6g7flJr
/8ooI9SYSJrloD0sTiSBLrn122jueJ3GsJ5ubCRa3mK+e6N9i1vKhO8wuDVErxiN
mxbv2uvaigsfTxxZKTAJ6xNaq6booJAd+dmur8iASQARaYTduvgA3hjPKppwAHwa
GSSNStYT+MfIazZoYgqNwEpOArRsaQbEWZJqzA32YZfcy0uOjkF6IO9k7/Qs7BFB
EvJX7HngvUCWIppCJSJgKrF1hk+9BL+G7n2h2+u47xe+C3W8DZ9cJNyUQsGwGEmQ
lAFctzmMDJinFW3bs3p29Gm/WKAd+IsERht2YuErf5LFZNkeAu2nRM6/Gg24p0eM
EFEknIZ9zXFuet7ynkCAa1qQHVi2nRCwZgbdwLfDcx6cAVuq3z+2YDGJ/njopMh3
8ddeDIFZYvHLR+vybRMOVZdFU5Pna/bywFWSb40qbzGxFj+JCOvvWZsmQ4xYDetM
gmzFZkq9jsJZD8CLd+HenfmcRWPgKETu2/+drF96F8Hp5muEm38nqYIbgyHbqudF
01OKu4Fkjz6FoaBulZOK6UNtNFFZiBTGxz0jS8hTCLa7ywBQ0o5+Gaq0YlMWvgmd
4dtyLFwTUj3ZwqxwDxBphAfpb22njMsdsDXt2hmPNDy7t7qaVA+mmbGpY3D4Zb2i
X8/T6GkS6yV9qUqddaubqITLH+HL8RfVYTAgcGcgNxiAVwOGu5xJ8crATl3JCis/
nv6giWos5ObpMWYAaFwmYNXrFlQZMlJ1kI9Y9kx5IBXHwO6Pb/g4VyMVZpULbvdo
Ja8mHQW3/KzCRtBZeTdrlXOjeDfDdBMAdf32qcWEE+6li7tUTqTXwHaoflDaoTRu
Xl5ZP7m/1vDLyYlZSx9n2Xy5E4sAS/Q8f7B4ze423uJ1uP9VcXlbacMa9h1ENbiL
buzXAbAQduU3Q9KvBqBs2KxP+mXnlx9OBcYPLqpvQ8bs4rlUOULoAuqOrGOUpA8J
sR5pbAzaNEoE28Is4gYKYIe0HkmS6t5l6LgxKRT+uIpQW0sZZyVIQNIYyygRgVsp
cZa39bhq2k69gjKw27oswMTCfX/qwFVJXeUL1utvRnnBEjlPa1IFnRZPd+BzFeK4
jv1tiPOoA3wVzcreJM7aYmBTuJKr2CAbpVE8kQe5iXZ68+YGbre1i5b8JDq1xr+1
iYMFAbv0G7+GAK3sPgE0+wQyB1motmt5GhuhJL59ev5xdbBsI1daVwyLgV64Jm6g
Yu6OykcDZuibTsaXlnWJ439nd336c0ncFO4/NUt/pBylyTuEvATTJpmpCLPOsaks
JVKa+uwHj7X1asPxbvymJcAFXUrbEtUxsyoh+kKrSX9DuF+Ru0EhMOoZOnJrj7Z0
4rIvdw1hUXNSlwvHEnVCQRdftK8P5KUFGvX/zOGQQ4usWhoDnw+B6wBWfRhgtBnY
8vwZjuTj0N1peEWHXLDVy7oLOVHEPsHzjKgJt2DXFfx0dqJfrU97J4HP06yXHe+Q
QKH0T+EdO7cUOqy595ukaSVrd3gJXw1F95ptOPeLwppFdmXFXYU40afTDjCcMkSW
4iVUhWLeRRIaLbhLspgX9ByULEModSsRUt3TnmaBQ7z/ga6cgbvTm9dwmoenZrHh
k5NDTqKbn/NEermWQ8QtPFTgOnJOtLocPj48ExnbyRM0ObASJjeRiE0kaqhdvMn/
JPKASqIUbEROs+kJSFsKwMzEF1W8NxMrIijEIrujK9LRjiae6wiV3Hv0Fztu4QQ+
FP1qxjukdvJtu4pKnjn7bxJ8pdc3cKBqICtVI/37HwNMtimOX4e0oqBufpxXJy5L
9MsiHRC7KdfAb7dam7v+upLW4VXu5NL/GA13atHIQhpiOeIuyRUJTRh2tdjSJcxC
aT3pqeGRiRqlrtwqEE2OD5O4/rv2a3j5t1dLNNT8kPzKQ2djGnjYhq0TpOZZdvid
eUdOcorphOQ04jh/3J5XaiZHDpLjuvPOFf7uCNYdG6HRIohb4/J4DJpv0nMLfbfJ
H5bSIU7cRixUY4Wu+W9hZZlM0XNFlVVAVX1qLBYl/dWQ2WntlMOqHmk7jN0+BhPV
0sPwE+l7XnYbx2cLZvHfYAXxs/MqkIKxZh1ZzJijtN0kkzidPtsDK6jZ4jRO4uuv
zJgA0koNp21liN05EBdZItcWXl+Hd4qCKuLsx0A1kSYWJWDddywyzLeRZW96SYBi
mLi8JZovdZffN+yWIPn9Wj17DgsGF1HjKhf5OKuUQ1x3iRL+J2LIeDkqxZfo+Ht9
lFLGqZKIEmDg1ffkmrnlu0qyKNNYMW9CdtNHPLF0XNtRG0SeNVN/klAj3M5lV655
w/Q+NxcN+C+QKDjzr3zVBSlWEFV2BktlItul271IlR3eGN9+98OR9Fb/oS6BLuph
9PvYKWurSzudBGO94MpWFStjs5wYKR8eCEKNBbSTQGecEeURm5ztCOxlzOP7zYDi
VhRIOtIwgW+jqtl0EBPTG7Te90dGGEMjRxIMnWUjT/bogxS+mqWkgzrby1ScoqDf
qujv92C4svnXhxDd2KHnXsRO95lxFGsB2dhRm85wU5bPCiZXm8je8Wxw08l8hSiY
1R16GnPKyGypHHTmqD1uLJRifKsSdOEnb+uNJCRIqEH5y0gt8reXveZAQdjHE2fK
EgNzZZ+Jcl2DsUOYtacRyg12OiCwj3A+jePnTzs2HQeqV9gSgFMDd+6iei/XYEgy
fomaqZHc1TQljRkj/8SoVIbVNb7bfsdyHPu9ftdfrDEfUseEkHd5qpdwFxdCfaJj
hb3HFInIaZsqsA7IhU/FQn/GmlMndWItAB50BloSs4c5scX4AOJRjUV17YeKpUx2
fx9T7vT/i9FqYEhNqOm0awfBeb8XAX9XSglRiW2/hzEjcVXYIaG7nminPm8Pnyjo
o4f+NOwKCxT1rvz6d1XnkkrhYthH9QsUqh661Tqac4MdPeEo9B4VcRMFa1yNAzPY
/Vunk8pHXQsWS+QXEbDZWmVHk4QK25TpFTNMbNgGYHb/LcRGH2+ABvHxsayEbWdM
xciFoJuqJbFhtobJKNaErUbhsQg8Qnq39ADCGLUHsAvvcLyOVD1b2rKRW10r5GpV
eR/PKzet3gMGJsUCpjkE95xjEk+xI4hDeEc35AE44f84tdxMphp1fQ2alqc/f4Md
xSyhQwmKo/7zsUoZEDUFuC1RUiXQ/nvT6fZ1ne38aRHt9Jmr29/E1WFoedmOMfJE
sKAnkCuNnBefSaTknbshBZIdGqj/ZKTrlhfmTBMusu2Tby+Mrud72o51dwG+uzed
aa1Au9NyvxDEdotgfk/5//+cfgyEnJ9sQgMJLhdLBJUXEFpmiNfQ8bz+plgALxIC
1S7Rqk7G+FN7wEjklkvXa2iIB/yJfYjPKoD5kmuVot59DcJ5ky/guDVKDD6cSryW
/74l8A88ouvcFYkveXKkUSmYl1WtJ/+rs7lhuRH1LEjFWVGkCqKHe+PSWxG1znmm
sWWhSWdkhDjnZS9chCL91eue9/p+lGn2fhYam4PRCO0S2OWWmrYarVr6DGsZ+ODb
3GSN5kCJQmQeXkEN+fXKyn52CsNhQeulTfNP0iwiyy4ampUK8zgwfDHoDZaocaVP
3FT3Uk6WcEPebv3oG06IxG4cmB2qcUzHH0/hnqAwV5RYg1/QKMsIXaF4ztpGk4PT
HKAEZE6C0gDEz3S6Ou0PTsGGrnMvBC89cFcx2+bZbTkW1Gpqq3PlBkj62vITfsTe
+XoSoawzcjUlBFAxyw4IkhfGgmWMRjx27Rm2Db7dtFSLmNu5kmNCck/iuzARKwT9
g5lt1OPV2YkLkTOO5CEyrxy+f2R5cR36caPzYdouqNnXa44fCuuwLcP7RGGPQUtl
1N89kCbL9foXlEq3kckw32AUx1tyPFfAN0K7GCfkrAjrT9+ciuLGJSZGtpsF7xDq
6yL0F/cjzhHXOsQOhQNK+n3VCEWFEBH3Bgyesfxa+gW3619GZRf2BD9NxBaf03/c
ikleOIGH10rV7RGBGFGzToqhfKPH9mygktjVNOWO6Pdvi/xd5EccEHM7rWud6BW3
ixiFuxp8lDF5FpH8QgRF1wkg2hoxerryI92FDXVO5pKkvIyalR0WW+BxAYTA2g+o
WsUWCas4V6149dIzL5fU1avJIX/o/QFVMw7sV0ExzEWPfmxJa0V2ecFQuA7+ATE4
nno8Z75ztnEsYKJjY+X1spXdtt/WLUJuoqPgmtPbxpNzqydZcgygQzH7/2ihp3Iz
2nN3qzdrvyoQNbFGA0yEgeIdu2mD64FXSLbXr68MtNjE4s96SC6HWg3qlxpeoFns
oSZnXvctl7RWXJYcBbx7O4QN1FZuo0wPejKFPnS54pKC9EDlgNq0nYEHCAQ2xhsQ
WWkHIajvrHcvVQUvFzx1egYn4nX3FSJP42mR4DRycZmigyMUuXTqx0F+i/S1Mm74
Y0cEucLmRs0/EVOpflxgYRXLa3XJ+kYNbaphOssKLyPCyb/Ej9HJsjEBbJAiokLR
boc7FNDF4k9cBCy2LC7KK1vymrs1pAsGMdS+vQdvHgGh9J8p9bq8OJT11lvsYFbu
oorNA2AIyIPueI+UqaGA32GxTSw2I4i4dpx/F9+fiwbZX1K/1Em72/bVDfoPTcOQ
kZq02nsxDLT93P3ZAtpBE2nKgjqZwL9ht70XcprTHZ2NF1x0aMwzx7z7Da533CKX
upkGjOOJVCapEuxnaE6axpe66nZKULntzFe+BM4rALXTbANdCwCHTG49iU5pBMaw
qYJEArwbajU23Mby4OiZUEQ+b/WhOHhU4hnKhlTgafROosNJ5opg2bQDoDSyxJiF
Ql+RuUOS+54lFt7SSOp6WIOtbQft2ILpeK3pbBYDoXoI7kYHqb7+gUzYa8hNz3ZL
raSIIibkkKbuhwLCwM2WBETDS5C2cCkW2450IX92Cgc5yFRc5TeFgQbJNLjUwBuf
BP581CNpShTILYxdmy+2ut5IyRJ4qcbW+VWrnEo0ZSRgn/A+vhM7thUi3fO9Up2y
oPjEz5yMiUxgBQPZ8zN06TesuKCxZLLfkZWawXPQfrTiikhIif09oaxrjbdldjFz
m/TbZ0RQHsM5LJd7JhokhXHXaBdhQTh/r94z+ew32rZ0Ul53jga1uGRJ/W4teDLX
8gTaM8ubXzNOBjiKEQLAGyuaKXfcFTjy7YnotdZmDajVFnJWA0NtRPJLrNe6KQ54
86ZUWBxEqO+8WxWUX1Q/OUv5GmSGPQhYKCd64JBMboAGB53zOhxo2jrTsYFyCZwO
NHS+DSmvSkBTgE8MBVsQu8thX5ZWgPx3wxzTVYxApYaGOvG9z0n/NAjme3YXyMpG
dQbsDsZvSEn/uch7PKSTYqZBMs5958waell3p8Lsfal/qZdmfdsWIYg71oBpk24R
IQtoVZDqzsua3TaRvTFenY8PqojKrsqwhgyreLEAn80HegOcV2uJpPmVN1S/6uHP
x0zQvOFDOhfPqrq7S34+nlfASSzCaoXqam7AZBan6a8NKrZS0UyCm/Svf2LwRn7J
ayIpnZkFh2hsR8IpLlykmMSv+491UjrUoEaUqeVgL84bSw3jlwSdZrj6GJyJG4UJ
R303JCCxAizevUPejZHrIEGcn9Age+V06dT9h9LHERfLHKKr+vh8DiI978PgRBCK
Tsq/XpTQEEiki/CRWpUuNeaJV1ykfyNelfFSWpEQ2mplEKaEQlvqWePbJITzn1j5
wvgQHzAl5j0fBSEADDLFesxStajG7yskYsmDhEKJgnlsTctbsuvaiBGF/3vwPmBO
8AsdFK2ejW5w/BpSlNeOWapb8aPqbg2xnsMvs0w3f+dEF63/GGOy5Tz4Prvs3y85
GISPulLOuLNURrD/dtRLjSH4f9nFvliyc7drYfgafEAbGpVE+KjD/ZY6Sjdw6xsL
50+G9PV1+PVPsnoX7WfmtzrhgqN6QfOO2WrWw98JkIkW1qkKIE0ueOxTG8x4V+dT
RF7V3MPZCGvbCN7nsGth3CHtAlzhPu7j24tyMcaJfyFy6NiE8YAjFDJu57pU8H5r
hRxsqW4MzR0nqNdptilJcj5b6MjxzJ28ok+e5+iUW7/HHiKZsdPlC2V76uXql1mk
HryUk0QR+MiLgVUXL4qwbrn87MG8xfbga/xSMaqsrkQpeMcf/9wabyO6QKyqn0OB
NLoldS1hOE9QYwCvLTk+j3++6VO9QxHipbGaVxl2f1PMs/ksI58Kp6pgmno5IgYS
fwlwfDqECITCo3L80SmhCyo0IsPG61UQ0n15Ct9Lq+WNIfgLnSmXDqCeZMCZKFY1
sXZmZ19JEd8VwCSQmKvbNwCAonz8lLoI5eRL0vbsig91ojXn1W48Ju19WoH6DSvX
1xoWtiBZsUvT5efloORA/YUCejMfIho2dlUHTwbLyVMDyOKpU4oMEivsTiNQu+TC
LckeGW2cp4BdY61VotIwR+wfleqVxLVZFmJqV8gzudCcUx0JBF4S5fhWBBtBhfQs
XxuiknFjLCgkP5SyE4Du0AokY+Hwf/N4uxJhyexbM8Uab3erZml5GstrVd8/qA9U
5dUDg+f0XB4AiufnTFrcLs6+WyJ4OSdARgbX5RtaGXycRf0sGiWqay35c6qXrkhz
cc8T4Oc4WYVsh1xrva9I2ArN4A639slFMkIVhFVMHWSKW8cXbwUN2Im3sBR8bGUH
J+SbfR9Xz6f0X0XRiKX1gZ60T4gt7HK+9sTWM+6atjJIHDvuqJk3Zt8LoeY3iTzZ
mBHO9g0ZRC/i0qe7cAImucWTQyhjRgg2cU6eXyysdF7wJYegPTXsAVes9h5Ntclo
seEKTlyXtsyHilq28+csAixlG4Z9jCiREm4FVs3kAppabIkKhI4ixxhVhRadNIuk
YkbLEe4IiNneVO41RH3hIDRvKTYzW6bkPQRDZpz2CNp7WhqzAIeH7Ya0oPjmqkdO
QZZR6QiX7vBh9wEXiZ4SQ/VDd9gswlQLI4vXoUlX8ORlotuOf+9sufLRvrrcSnis
UILGWgjeV2SYE69Ea2dxEjY4yPETgPt0ET2DSD5HPEn1kZYx0vQvoVdCtJF22LsL
7KNc44vtIvsZqq7B/RUcQeU9XY3k9hbE7KZVYERCfoZwcDiMt+0kxwb9yMYBV3Ih
wm8/uMpm8R8cRMlAINs1nQfoeqods0b/lNd9ha0s6UHCiGtqgaQ7pOTuZdbQk2AJ
upo+NboOcfl7VCSjM7Yo7qBZKt/oK76LYqV9O9jyuhTqZ2UOwuXHOKORu2RZucCd
xYNRwosJ/bDxfPKvHT+8E0U6T2vKIg+TLtjmtLFdB1P75zYTp/MbkSH4yYM/XOBF
pzMEw/B0i7oeaEoScc20f62b9rPl7torr+6hvD3oPaGjn4lX5nU0zeY4ZoUpC0+O
b9t8pDyz9cA47bRzS+Cp2O3ivLrk9b/S2SMJ3cMPDcOJ2aYE6j4kNNnhJuqQbWIY
zSy8vOvCw7JpUZiyShdFmotZYasyajA88t3aiIDX+NAriwAVKiS9tazjVQ2fmh4y
V6R7af/RuK5nl/3aRAiB7O96pPWcY6RfwFv8QVTlciubiLkPrJ0NnVqluespyt2Z
fI69QSwkRlzSzDYjkr0sBdI6YepBm9FTDWSz1VZ/Sxifi+gSrUzUYKnjrerM74lc
HhQUSql08gKAst1gQRaf0QwoMIjNj+WwQSP+H8pZHQTFV0j1Zjv8i2ej+jEEa3iq
Rx1Aq16JBZ2yb+gRQN0ROGo0vgKW2MJd8A/A4cnk3XIVPmRCt4XDGftSlSznj4zL
qQtBltcKKZEpvyVHcAHSo5HT8l22YKBYxVuu1AOObil6J/KJaazSMtXCl8Wt0OEm
iON2PrnlpKA5RYx/4ej/rEUFREAhY+JCeDf8dxroUwPomze5MVcfK64dGGxNpbjQ
0ExZCu2iHSCK3mWB6yMBJvECf4W011YnyKDNTUA+uwLXR/lJHwWIaPkpP6OkvvSd
GMb2rF96Is72kw8x2kSpjShzZDEL9CZ9cxeT37fCZyonMC31C6w+wMBeIhcVLGjm
WjZkg/ZRXHPgDq2FT58jxkWY6LRWOtJboyactsE/pcKKtwbpJEKtMxb3W4gbGWJ7
MGEj/5qKxh/MA+AeYaP7JuOsI9uQaL4BgVcnWbU+kF7ipq2btazoH4TEE2auYYDv
jrC8X19rF/X0+WpsaV92k7NkV3yxTDEnYVTn44cf3wC2FyzN2dHOgvAbj0+tWYrl
aTsL8nHW7o0KEVeCG9tj96/SvoezXynPXmxh6eu0lC0Ex8P/9jGaAkdHe0xUfOeF
4G9EkuhCjSgtnzvHpQ3VqRFoz/lMCfq/tJ+3DLpA3w8lzepNvjdhwVfkEcZDCr9F
2bsOgoaOe71ZIZaoU9wPTf93pMh1O3CXJmQedu6A8Uc6DJqJ4DHsD1O56P19F4xT
dAgB3GLUW6+CUWr5dmcN1CWNkJxqMxGCfA6IeHYVM2iRc0snIZuCk05hfiLZ1tDY
xlSnrmtIgN6nm01vKI3clzsmUKBA03cNkhGwwHz9QdUQZABodkYdPb/OLhMMiBWl
y4ak+xJGJ7v6OB1AmYaF/Hi9fe829oXDxfVBpXq3fdBLMF9lRO6wzo+oHkXAWsNg
sRp9CDdLfRg0QbHTDx8abV2HueicNz9BT59l+T3haHAWQcefV1eQkqqfFjWtPh4W
bmaVSqKhfMhQRkwUeq9Bt6umyFSVpaoODbv+3bpziS0i0PJmQ6voGQYnZt3E+1b8
3Y7yH0C8N1Q5xP6ojKDMKlLTPUkJxCLEcZQ+g9SPbmkQrmSwZ4O0RmS7ImZLoKdV
ry9ZYUM0XD8GgWmVu6YbVewnj+YPVChqygU0zziF3otSaqHxRz+hKogvWvw6r5vN
/3+B7aG3Xo1tcgC8fVdJJk5T7Br4y9VB9AyYIqVX8vk+HIA00KHnznVu+t0xh+J1
ClBtaDZSTxooyIgGUx+M0crE3KdAN91dSyNw/n1dJ8/rZiZh/3U/kf6yK6Ly+a6D
xckKo/uKVNvnIiJH68YLTaYY66BXyXoJ5xikBv1UnK2lLF0Bs0hKj/oBDF4txGzB
Tvow58+GU523NO5bSyo341PprmNw0VasJBn9afN1RNF8JaJLwyjcWmt9ObBivCAR
xmOmYOMdgU0Mu/apNZJBSVS0rv2s1dkpRZI3p7kbqp2G2IxDWWL94mkIKZv/5WCj
Ekbj72Vd2k+2SvG05AxvgJpGjMcwB1NaQYC7Ek8MXhexXmzdY06onmXpabujDDSI
HqQfTe2M1+Kg6v5wQ/BYMSBOjHlE9fTwwCSy+J9yDaP/KQobt+7IMPC/yCKXcsSL
Ujx+F912KFSBgEm5mNL8HmbMQQzGnI5G3t+LotGWVZHnwhQQvvuGp1dRULaS2orS
wo5jXtD+di4z+79bKkIqsxBt5QcCjF8R+kfIJzj3rgd6QkgTwRyoLjmyIq7zQ0YJ
q9kaHMsRexZcRMnep/cfiltEuJn9HhIY7lAP1xvVrWdvV1CnazZmiPTozbySGIJt
aYm/91C/1ufgPs9KmwGn0lH2oxiNgkrQ74MdD+q1l/CR0mrApyVhWCIIFOubXepP
vtS1Ez8mtF0MGrgYdMNzPhbsCi+LnxH+BzfQB8FX0nHtRz443WCjWJwCKanIF0lV
KgVj3qLicPcaUcNIPODhohOods/XuBbzclO3jDD3o2/aUCafzuywYTU6c2Kr6E0t
LrKLgXfyAVVvbwOA5pUdQq157l6zEGESp0NHQ28cNvuj/45zyWBL6qMWN+NWucsR
4MZ1uJamTz2gOrqc7merbXzLZ9XLCu3rZJcab1prFZzRTly1Y/Nj5oSKukmo1KHS
1cmLr/1Q2zuivuyqjLoi0J2QdRKV+7YYE2kc8zZmbT3ae8QWWdPN5KO5jS4cEPEM
5pvQ/k8LlbsyLR0lEndaSI3AfQ+MSSWIk+008cPY+cHNIL+X35s1U5CMYihAYv0H
nQHnIUnfl+MhpZHdD/IXo4Qbd4BhpcJ/2mgJQBxzczFi8RhoRN7T+yaOakccEzPo
aY0EYOVrJU/RyHuaUy1NxnMMcVlH60q1dThZwONzbxEwht28nxPU0HACLMRofZ8I
o3Uo+VWjMBO0uLVALvQdkt4VC4THxVItQ54Tx1PuQibXopWf5QAZIlJSHl0A+PfY
z5a0ly5WQUMi4eTui0jNc/HH4TwTIXxt+kJy6Tu4xkxl7cJ/FbcMKiP6DS9iGYkx
2a/6B5R2Wi0RbGB5UXZH7Ke2+b7mzeJEX+xJUrJz3q1lUpe6Bn86RQZDanSYpdJC
FA/1b/PFlQEVQlQDpfcXrzx5H9VXGgqJGJvCqraQVTnDHgqi6/i8ROlTarhwB/Im
SbTA8Qrm40tDagWQcqF9wAb1gyCIQASdt6CNuS2x+4ZlaXLQjl4MK0B2jSoO4RYY
ikNQ23cmOFb8wtImAoQ93QJl1s/UbrHR4CSVl7GxGJzoJCgFK0o695AoUEJczoG8
kYMbikZwr0ZL/z6WLDuIzAcEwIVQVq4RL8nt8h61WH5SbcO4ucR+jAn32mtckwlz
Rw+JWSSxM3fk90HtKQrlARog7kLQpnkSMPtbRoKlbePwdw5i52C4Id6S3ZURlilV
Z0QEG5lPBhP0xVTfgELzxPiFUhYmv13a/67ak+H3GeyJqN+YUbMYCy3qfK/C7xIF
UBKUfZiXpkewp0JOE24UtDsA5UdembV7/8vjHXHEuQNSjn68V5sJkFjPxaKe5pIL
0erCSiaBWMV844pPcy5OV5JDPdl8BFnwMhrPB1x1Ddj8gW1Q7fyl/xlRgpNf62bt
SyJgnHW+NfpQP6HJnTVPQ2MN8dU0Dvn0nobsiKxCkEILqoj/bPL2OxmhmKGSKoro
lYcRtAcnixZcT3rhmMEe7lU5F9j2mGwBZFMCcH4vJ9KeOIk3tF9XDQx0dRaxpqge
d7pyqS8Ie80XKa3rXjoiHRKBHsg4/tw3swnYAZNLJI7VD267mZZ0mL9Pel4GPSm8
IuAOicl32IuUAinuOa5LSBUam0hXh1OXmwKZLwC3NhkbBWwflVPhB3OEobvWTMMA
LVjKlVsIK4HgcfEaDp/FmCE3rWJYDftHmiM/2bin+HaC4yLPj0A+5fguOw4fWf+0
PXUiLWdAgLc56eOJrmiAxxzag0HWlf4eo4NDgUdmA8ZnyedRdtb/UOxWs2qiI+4U
C9QF8JYOrm/SecHgEB2NSbJ5S2Pel+0vga59HWEk8U7dnPxN+YIoatFEJXn5AVZl
fk5qmpXjGEKmwgl/szwyo+CZnlVl7hY7IzWmE+g4fQR276uU/EZ4z4c6tUoKSu8u
mQN3llubz2wR7K9gI1sYyrMHO3YnEAqRC4CdMzCPjoLfNmALGKdzrbkVzdPGb7LF
7up+pdS5PYQykhxYU/JmCWhOF1wIlFyUcR2AmpxnilOVnH4wPMOxzX2Ae07YxmNz
47l+aYKu8oQKGhbnOj9LoFYbz4555jBnsx6DEavlmedooCf/fEko05AHKNfF+OQw
zp7rB/ukr4TR+aHs/Qf8OWazaqJ4VwvglsVySBQEZY2YdI6TiMS+ELoYtPYR+h3K
4IfStCQr5JmqmTXpToLQBLyXboPXjcQqC0Yh+6U0MTJjBkjsY9NtdfgpA0lW8bz+
IDrHERXijo1wlBg8GXmjRH3dXyHfYh7bms+ZSCtgHh1qMt9y2vQ7gjC8KmGTJEOL
HyswMFN7/Ql07cSN+r9NneA3rQi/c+4hA6orszvDZ2rDBfWiPgHfxcSP1bfIlLE1
f6zTuuonht/sVxYqOEjOh/rIIOEFa5CjYpRfJUHxxp1/GI6SusdTTDs0sYUoUfDJ
QvDJISa6qfk668hzycH+dV0B2FeIC6a4RyLls3or7OXtCA5j4EXsNtJoIr4JA4mK
27uwbzT9tk8VOCfZPxtshV7mJ7Cf+gQhp+LTrnVGPuSgNVwjp/uelL6bVpG+AU0d
6ytDjSQAvcfTK0GkAcu6vV81GoGllUdJuojHJB09bnCl12nkV9QguZATpWYZsJy/
SrjoCbcDlfEuBf0qYFR7+g54t28EO1AGdPuUAG1HN3u0cCEzdQqFC3VCgk0yma2P
+JEExVyuSQPbByL1vKElBMzXPXG4TIfujvLVM4Wfx2HoYU5diWNxW+Opurx1hy07
ibef+wpid5FwqVW25Qyp0Dsakam05RqKMo9uJJCeM6vM1ks0AgAqiiYXFOXVifNY
1oMxFLBt1Vis5QHbAlYSqnf2947e0ODCFYJ8a53U5o/uhO4eJJ7JnPi9HY2q0vPa
gRr/3OLFL7Efi5MqMlw6Fad84U1xlzjSSq8OuD+xSWBNNwVSBPctzzhH4XceoOpB
ZSF19u3k2daAA8HdAYHnGU6Qk2hSNDWnHddv4DbDo7XCnus85b0+vmI4ODUY/Sza
hMnmNqFVidwnksTl4UVWI3kQxBEnAoVriTlHE90WfyHsxzqKZgur4AHRgFA/KcUj
X9hAonR4ZUuxdhVBiwf51lM4io6xBWDeaA8LFAcuek9LZ4VGIB/UeHhuB9x2QL3M
uAy7YPPTLzXXAdIb1Ul7LGAcCYuVGg/Dbjhic4r5ApHqbPShCwclUpTigaE9GNJX
scblpYwYA0JZ5oNlJkM/GSEJSzvPQK4VEoUemIQ9uGklKesccHQXGS/uSgVfb9B3
m0AlDBQPuqmO1DNg4hIn8uM8VpTytei5IUfLyiEJUx9IJ8iklJC63QPVeUZVhB1k
xZBxlG/I+ROvgumFKrZtojsKpXvUhp52NgCcrFVMYfTc+IjAPaA7zXchinKG6NGh
TcBcva4uvDAoJ8dFVqZD+8zRb/cPNQQVJU0EPcNG13VGmuoUVTcK1fJG+kVoVhA2
uLZ74GBc53kt3eRtOLQQczjhB0297VHTFqrdh6xwKKPoc0vW7Gm3AdCeqdaqajBb
SI4gHxhvjd/Fe1FTCvqKF0WIfxvQkZG2h5WliK6pOxm6FyuQMkFjLF9czQGWkX87
JPTGKjwwDNBPxhYmo9xY0pqCtRCJExlAi371/xARvw9xu7XDWFPKyEOwweTrFA2r
7LAETvd3C+cGAx2NDi7RRIIbLXNmBQGVDtlQGIQwAWoEcXVGQmzVAhsqfPHAGzVa
Y4SlYKfk2e2R0rZdXobgptHW0LSSv41rTQSN0WNA7mKZqRRu9LsF4A+1wDHno6sP
tQfhl7wXbEGFP1jFUkhBA/Gy6Crnf0eagmr9Wb/cwBTFVYbNLShv4gtKUS9z2ROX
DbTm7CAcUiCKWSi9xnDI7RhyeiKBd5lO5s11e6Mb1MrjKJKZ95tZ/eCQR9ivO2cV
a42R+BANHOHMGo/whxLL9vrLFcaukwblHzehZAn7VrefJw9JMftsBeOrIPGiK981
86eFFnt14ZpOnYtkOZvXjdmj4e/uDC8pbQtMryvNLiWcQfauWD6O1yb7plPFO6Zp
6BFcqG3YMtSWagVxfpIIqHvG4N00yk60Cs/zP0rIqt/DAfOAjs8oBn3GFooyw3lH
inxECzptn3UjzUsbu04oz39zDEIxBXYAM4zSxN+vDwRtskNU5jWT4KbJuP+CvpDO
vu2jjbK3bQ9hZkUX0EBXv7HqjiUR88WRZPISCEXdorzNB51oJfqvl6iSHN+TFPrx
V2pDc3ROQ2iUj2c0f/mDsr9j2Imrs7n9p+34jX0qou4nAbZ1lIPMWtIjJYAgcWnj
pkvDn3cxKuc9eu91hU3ReHnvDQcCEOnmS2cdVRoyTPficZNL9YqA0vtrxZhGwBVR
lJG9EvFOpyIQ65pn7hTfxDejnN4EG+9PQs2TtCUp0UmPHAwKiNriCCXJvbKvhHVi
4Qsb0uN++kVeaNe5/t73KTOQMZHVEcholWJvMGLIJGEtpDgjChKFuZ4u7iApS/DJ
6d9qx8kSkhMY0BHnPV0KBj+GgiVfETkQUARz1HqiJB1oGzf589Os+63nMPACPH3E
oxQQLz27IbGttGcN5rK0bkbh7QsW5wiAaAuuqkMzNQ4biM0y1Gp4rYCBAQ89mJSW
oI5gK+mQNlNmUvlSG+Nf+GPlEF5XLjKzJmd94gLM4gZd1ePcZmMHmF2hlD6LSp+7
Dj8n5jWPo/CrwawET9YHC3cRs8dSEWURngpmM3xY9DVssBEgHfoTRdD0lFmK1Xh0
oKCRDkaEKRO7ia5629eGZdSLiibUh3OrnOhOOAEhq9Dk+cjuj2I95rg/6W/x4fSk
QHbni51yrIBfafALkfbTTcWMgX83DTLCh4pylMAVVLk5P8p6a9pGK3ZlG/aIVv3l
wm73PPD8rrgiIxYFxgzJ1Lm4DizGQSyD8hXZNzKveP7sYJgRetgGiGNeGfaD0cHr
k4znLM+Lc4ShNBnhz+U03khvcF1gZh0hX1IWdVyUgd1oK3cbRZh5dEvRdN7mjX4t
uWSV0HH42rGK2YWSA49Hw+jkLngVnrBXDeceI8/797RnWpG5+HQn9W16OjLcWuad
oEavv8YIlF94MyEbQA6zVZ/fYpVN85yNowTWnbxd0TOSKpDuIAawY4rspxZ+HYem
jaMyEJtjwtybu5PzfkcW6OpI8aXFYMNTy2a/VG5GlJ0iF7hIlL50apA0RraWA4b0
Fd0YOgKkyjz5MT/N/b+yH7LEq/lf6mDl6O2MYM+kySgoY44OZHVGcEh385lDhD/f
yWBmF2A2FiSJnmArfS9eNWQbdYdToZ+ERzxSa8fOeLtPcOIVPMmTtt3H72wdR7sn
B+fUueaf17t+IjI79pUysA876bz+Qbz6Ims6XdpHU35k3lUOqxgpwr064YYkxgbK
2COdFl+ZwQzkKiNdVMtx7VUcqRPh4qDGN8apPSzCVKNQSxRR5Rpu+X2+FM823O63
LsddmQEBUHr20gT0sSm+Mp+Z1bX1ypXaKAoKkwLrIxOC6I4IAvXZlhya4VV2wnA2
OEDThvi6QfIjObXGAUa+yaTuopngMIVV2qXmnE5lv1kw07eLHgnWqW282Usv9Iq4
vIlBqX91dfoZBFZbux/WkkjGBZt6chniMtrAitsrv+p6YmAvnZbreRSDth9TTgT2
px6nMuyPKKUTEZ7OslxMPsrP7LvTGf2vGjOcFH/bmzOTGtYAkvJUV2T23ojE5DwP
u2FFVxcJnX5qSFNo8uu4zWxI175M8d2q9onmtEtjsznu5T97Plp6WNDRbVzFMrkA
FCtwgdxDJEWiNRJ4oSUg1kMm4PqrIGC7V95VIbayUP0zb8hDdzN3baD++jSNaE99
Q91RQCQYWQD4/BmaKy4TdEnJ7JK/VIJgO2Qe3RYucoL/jboeZIlzmFDoVQRcTlFu
e8HVMw5RGRP5HeLOF1sKPcPITccavTxVdgnWzbshfhqlfFvfRrM4ppNO7mlNjkg/
iKanMtGSIpRY/bOMC8z7zkK7k9CZGvaD692/zq5pPwayAEoxUK4MdcDij6ZZYLFL
ArZjCOZRHSmTrpp2O4vODqNRs8EW3M0+kNM9hJU6TukwpHuO70Y/XyonH0fRoHD1
uQDywt6Pkhx5VivJg12KDA4latGlZeT9h33i3ara09Fb7175mKaOU3EiIcuIo40t
ZBaHAfAkAIFkpxFTBcchk9zyzUzMmpjLwCJ6rQw3K9CuOWkvWuL6sb9EZZp9WgD8
uIUEVd5BpbjyXgItEZR4pgJA6rRH4rxbmve36A5TS4rT2i0O0VwkRTp3O1pfqCA1
AvkpwlidsKbAOCTguwa5kUrSYVn0IBnAzYcR95UlZBd6P9WjGvsARkVggsRTKQf0
jQ3SDSZ0WOifJHKWzTGllVgma3fflaOPOxWxQizEIx+jmuVUBDoQnP7RodCk80Op
SOMZ4Il44EMWCTzAJfwZ0unFstJmYzw7VHDAQIBCytdzyyXPiLsGkKpfcX3lFvI1
YXk6GfuF7pNM6yrKFXCx7t4ar+DxBhwgpsumTJp+dEh/8nl1H9O/4dtKiMgEoz2s
RJVD+qf521r5P9Yap+Nrwt3SERNHn0If1+r9c+ddDZuRScun673IgcOvQQ3C2HoQ
GwAiyDRKFrDGCGFvMJTf0nmq3jzPxz4z+WVvdRHqpcURqql0kBRDlkI0IKu83jSJ
kwa8b8/8EZettyEe4lvpRhNd6WL2f/torQX4+A0tTIrRDHLJ2WtyVXHrsF6lyGD5
btJjtgCnEB+z9kaM4l2xfVvfbFcg1bhuGWOQP38/IM/V8icBp0tE4NePhFa1s5yH
aGMLA8acUE4L86iah3bEIkWv6uEmCRht36BYmwm3hJ/VD38J25BIk9VanJsEWreq
YL4w1sSsgfHCDnQLKFvR9HUASF5l09hRvRs5s96PxxUmmfZqhjyIk3oLgdz0PVB+
dCQiSQgnp/zyiZj7cxusWN4QtfHgNkoI91MUixdopZSeEJh2SxL157YmI1uU4C9A
53T89WKaiTjTnDHxoLrhX3VtQOoHFXxA+UzkNNC5EnGM88K0si6p3rL+Fdt5aUqG
cLRbvLxCaDNnZOo7KGLwX2xRf7IaHFTG1U8lxiwex2yD7ysZfvC+utNqnHrymL48
AqiwOwtHEuidHIywgmpRFAj7t54iRAJPd9G2O8mBBrZ2wFidzE2Utr0XiF8Mj4x/
vwS66tZwpOI9JXbfMoImgya92ry1vO4qhjMpShkjh8unKux4N23hTPemSMhE782T
Xcs4XG3iqeV2Jo/SYHTcfbYr1U5iu13441zE2h9j3ABRAeyN1/aVjREeGWwC3yIF
d/j44OKkfgnefKwRQFkhRDlk2QqAELRJqYyMUJoWwB3gUKDK/U6Ury2SIaADLDdD
gKFce8yWhVa3WnYCfhi2mG30hjAvaPjF+2X/Ohod+WOIYqT4LWuYhWTqzcnELcZc
VqOU7BFy37fx4HNv4/FLgKL1FdaHRbjhZy5ZD4kDHcEDU8BQD55mtzPgFS4t2Krd
S2rJbaQH8SABqsLqLZ9GvohvV0J4TtaY3tB+eyQYwpT/4LTVVuO6Zg97HBNSublQ
+PAEP/c0GhpbdeOjHn/u7hGfOvWJFEg+Y3R/2haELvowz4zNvywQnSWFNxCw7qeC
MWaA+bziWj4GJrDVKVOD5G08VgHx0i+omdrMi9Cb/ePXWIlIsn4Yp148d23y4wAO
pUa32HK1XOThoyqZ7OOL0oby22DdRvuD/UsJErsxh7Yes7ZmkVW+8D95rgR0Hbxj
AAhGm9aistMO8JqrMKIl7ieXCFnygZl1vOoDNprmeJ6r512JmYqzJTAvzQbZcCG4
VGCVf4YMunMwtQXBPT00RrM8dB+ccR2YnQDciJ4yhgRc6EMr5z16iz3SZI6Api+X
IgIDdnQGscTDqNQcp3x92GJyBtMU5jb9Rd1afxVQAp5sZNT9w2jZZkOc1ORk+siv
/CizKpVt9NswQ6c0/fskvrjVmSvOseW5gGHgr0aSZM+Wmdo3bvZZiCSuU35X7wq6
quPj8xXepEajDb/VnbjjxEVO/+6mk5/GeW5b+/RP0PRnnyxBQsMWbkOVGPlNUN3w
x6hdjUH+ZJp9yF9CvtWwxBErNXLQFHBUwjhb8mGshbjl4o1KfsLV2BdD+Zny+BVi
eOabPg2S6UF5zMUhRwxtrd0VdCzVc992xHYS1aws+5rdfiWq9m0oRHHblneCh4Vy
G++1APjAkbDHH6AnEu//mpZkITs64oUsXd/bbeSeHFhZd09FtPlUtUhkrgpi4LYV
P2p2EtHKDf0Y5aJs5SqE3d0Oavm/iRuEj6ugymqS7lvXiZJrJOHq5DoSzWO2acMD
wXVdTv2q8fGmE9M0HhV5XyWQ6ws6aYKyrHgxuXxpI0nA8FCZE05dpK1nmxoyA+3u
ZUhyikHHnppzz8VulUjwu8ABl2USAOhwsH/+2JtWiE3fA5ZPoJKTM2EcS6Wn67/4
bJOY2dyBQZOPXyVJEppRt1LI9SSll8pmsPLSd2XkYNI9NsDAo1XzBEReUCUetUHY
XrBlppPX54HKTCu/upwmzt0rw065sFFcF7c1BxG6eNJbIcUityduyhDYBT15uHob
ELHZmB6LpP/P0CKBbblbp14ttM8SEU6o0xWSKHWWzS2Gz/CW9BJktkHv1hgKeDv4
qIglABanDkiteJv1p2rbTvB8Po9I5VzpPfWQKrxFISCKmtUHvT33RmWhKl6BD8hW
F5vWTIIp4Ff+dkmiPAkCOaGZvm71WPWU2//7xkQcsIvvg2FQvjppkEA6DmeHmzMg
cN79SKscCs0cYZJ44HWJn8FD+ZSvxoTrYV7yyQLfOpU7JmwSSqkN1+4fxIiGm9bp
xE9WjH5JpfATwj7S4OelzoKxjZ29fmxM8dM4oR7GLB21NcvVGTijZO1wdnhQajjY
WYq6vzQrIxDAsB1wVhmIMbcB7l4AMS0K05v9qr0x/iGaXjkkbqSedorDR9pop01W
zTnRq21jrYU1TbBTIpOMV+/KpjwuYXSuTi31Gwv62jB8JbLhQo4ZJ0Hh4hgynni5
aiNGuVTMmxo6wd891mfu7HKVMb3JbyK2sNqBz4UCFqtXMFEaD/Z1yGZmuDkUgnXn
Ob0bnND0wC1sBZ3gg8qgTKWBTpM7xXUC6ZJ1svwCCU4pDCcPcFA4ewzyjv1NOOpi
OfHYqXoiL5znLQVHxxVfyLqbKt+rxE0cSfkxw8GVhgOUhvXKF6U5Xk2HnQPE32TG
33v/DAJU4Hvr1zHo5P/hi6gPnp0iFjpC7PQwJm8ehHDsqRA6iYSeuSjx+eA1CEi1
Mr+0Bw6Wicc4qx9GOCzh1LOQyOQrBaqLPJ87YBwL3sUdxxUPl9UCiNdEHjfJ5Y9+
WPgv9l8x4W5Y8Kq5XywTbJe7j7vM438tYUrA+HY4odu4Tnoxn39zjhYbnL73djA/
6idmjnQFlwAoTMlQUuUEnST0SkV8w+CAcI8NeCnQyUGQpRSGK6JBstf2zBlG3tCZ
H3vU4b6XVf0vYh1j7srguXYLo9niYOmxpxchtf3JccWBHINgjm7P758jyeaGzwco
UyKgxzRf/JME8STco7b+sse01M7Im1FCBTnTNlpE9UOvBDpOYXNQ/DsigqBu2pam
Ruhc6u5rhqqyHKgIJD8UwJwOX+1bpNzVO/wf1HnzBYYVBa0Lk9UbwM9nYhfiXVdk
jSwwVaIvMkijQKb/+Tfd9e1TbAj5bb0v85PIGqKpyUvrqvs8UMq8SxRMeAivGBmI
0RnXSHyTwrnPX2wEOTQQVpAjOCDtlCAwIajVL3EJes2ZHOs11jy192dSyiFHIo9h
cDwWBaM9ER06UMBhI2NCODC5jFDdFiCxo7mlucMoNNSgh8oq9N2bJ0cG3RwX6Gee
nfh3rVINO3qfymiYYaJKC8/yV1NfatgdDE27rad1xm/weHQgG4BwNEGEMkxVedHd
CvYpSPsaNDR+Qx9Adf4DlN4GPf20YKUTL7H3043kkL2dzO/XpNnDGxjLFeNxNH+G
knTUXPq4tSCLhICdjNEfElQ4vg+qSEKQdcz1XJrTFVtKOj6ABVopfPvloGYAoK0i
sC2KUKBLtxn0Wm0BnugY8InFrwqu5N+P7nR4OqTuppa5tyjHYxMP3qF4qd2/oLra
hjhpmtNC9staP/+R2BR4/0sfNMPNctb38t5yRfnYGY3p3PlPBTjbvwB4v8/XmLHt
U9SwXtlUbsWCQp7IRvOoOhuh2XtewCuVU+ND+LP3T8wYnm2CESeD5NHzX0MPXHhI
dAg2dKSA3qmnf69WcgbjwFQ3FZPzZgBbD9sky/6ZlRhUJqhtvu66n+QGuTfriXSq
R7THE4u3nyH1t4ZXqAXZ3Jxgc/0CuP4x1lPm5594d7X6BoYeMwiaGJ9Vf4h0WHUi
1lxS3sBDkxIWyjVd/9irikJ86nJvALEJIyE9xCvfaIL8eI4TxjSuCO8D5r5dSr4i
8tRVk2Hz3qnYtqgSjwCrGfFkyUcHIUJWRUxs7WmDy9s/FNZeglKuPOJwynaQXFih
qzMb/KrMj35wHd1aKHpi4SWyMK7C/pUEst8zDpzd2+anIqo73mxjweGWwnmEEH+u
/zNWFJQNaOatARGay5NVhA4bx6YqYOYys2QHD15OGkMDrxAKNL4LExMtlJRLCTE4
qMru2vgy38cB+kbr4/L0T40jS+fnxfRlHM1Mj/5liNMvyOZScNLFyg0jy0pF01NW
mzRtjdJdG3ItUxN5/I5YbW3FSX2HhgMmmEdS9XK0LLwGkUpyYoPOlniAcIjbxgu5
r24VA9lPZ/pbVgU2cJl5rw7XjHvUaCJwVkg8ivcJ1IU+sunVxy0q8rMpOJ5uxmiG
n8uDJblsgjrA+b5djCvwKwnjQ2tsHV40MTCw5QEK8RySJ2yQkZbpVANenniHW6lH
VmZe3BUHLELKD3BJwYGZlNOO8+OSJz2r925uPCuN509UB0ovNyEXmnH8DZ8wkccz
h304d++vBznCFFdWb3o3JQYmx0vdyZDOVm98GA2g8/69ZZPPKACK/9sjS0C2ASUU
hYM8JAZPcViv4c15tBdoAmoWgmc10YrnLleDZ+gfJdgR6kkiD5d+TL0MmC9at4y1
R3VmASGZy9JYS4wMoThIphyWDwLhRIwolCDItxQ2iPCUNGCFuTOxML361RDAlM8R
46744pWBrRtoDfWPAySg3NHUcsjxnJpC0dRQciot6RrAo8XScbY0oIEzMHzQHTWD
uwgbB7NG8jTL6pHY+ZtaLmDALP9wMvpqzn3iRWQqKAw9BqSvislkLMe2KjI5J4+I
Yxx2semUXpKKPbXa7pPKW861UQDr1j8k6WvzF4oFm24/faA9IPn3hxBLnPSGDT/Z
hSHIG40vFgKexlcXRmwUzWyZkuilquoPc5sUC+1QpPYvJfi5nLvLWjLSBDrEnusm
RdVL/809rVA5Z72SWtC7lt9WV0OLmhucyf8spfPG6W6pQDVdXZo1JtuXDftdigUy
ttnxAZqHv5NwQmGf6gUlSR3R8sDC2Cq6gDobxN7mmYambcUSete4rCvHnR70aNNW
d3GLnGn7a/ZDCCgCAn6uUGYCZB/V5jlD32PYK92yMp9uI2vNNVUJX0+BvxplOp4S
4HrenqBM7hEXI/9+2e5WH1riE9MZYE9VtZRaIqvhBUM5h49q8Lygym4TICSW7VpX
rMeT7KSD5vJr6wxxUzKWB4xgQsYjR+oskyp5aAfluhYCs0ol56mdMnv6E+0x4udX
JZA/I/bcTIwuO3xbkAb1Tvv6pTDOCMGgrvLtQarmQ19dxnMhNj015ATbnsHs4zOj
H5G10jmKX6okyROzoCBaw1GPJM1ecLbkBe+Wc8PxHD2+C0wproHkFAggod1urz1b
/gI/c2VNbUE61SDv1AWjPWuIV94Gz6hSg1lIrN1GrLsSXz2y9aGyFlQwBe/zESYv
ZmkpFDLgwq0aHWjZlFjZOEztpP7NwXIQguZEpCQZ90a3U5fln9StTUHK5en6kT9K
Id/GiMrDer4SvpqZBh6zL9l/ZGCcEkb3YjyG12CPqJXwRVDC1UipQ6kH05a7XvhC
5VnyeRLMqPLrr3bO4jkKGK+WkPIshS6XGkShIKtgw6ZWSbI7WaPruHJc7kIIkMWL
a3Pm36NfewVhovH0OkyLtzo3TiEWq7LPHnWVdcQvE/yGtxVn97e7WmWP0deZEgMq
Li71oFew0dEdq1WrX+xWFFhIIEKaZsEHGn2oprR0EEVftZ0pOPp0aRLcJv5QCOGc
R4V2d0NvS+yZMOwASn11KbmsnLZNIQwN9Jexdq96RyiBaGlMTBMetd04MvlAs2TA
7/86MJlZ9j1TLqswIE2LsOLBHfAokEQmIQKb/4blpHN9NOCN9fYP2ZLbztK2g2TZ
d0NtlPvu1R72BY6e2gl+eUnzsSirbuCoQq4FOahaTr7kgDPQRNTQd3tn++Jsc3bc
lW0r5SlYD6ghZVFXA3pskM06gYDw3eoI1fc/bM5OBQVtO4K+gHQJZh2usoY17wnv
RuNVrpM7PJRMF7DeaAubbBVz+FUE1UbJfOLCBSQaA7r2yLB3/K7AM0VosTs7gjoZ
lqXy5q/h8gNXO9BHoKKVTbJe/GA3axfAD8W+R5vv9Nx9+MwBNgs2pYUyRLeRlADG
FR+syL5cLHOUUDYXOeK5v+JvXLBn7UD2IsNyPrGFpXXKoT+dz57xKAWzzX+1H8J/
AbyDc65Fm41GT+vluH8N+Ajz+qc9jsbEcFVIgnGCFhmr42dfzlDJ9DJy7bg1guT6
Gf9mC7IAJ3mdBIQ6gzNszdtkQVt2maf7YIXqOYNDuNStaOMrcaPXVMa5AT/pajcb
IVyqAyIap5d7KP2dnOLu22+rUl+NxKTMh6aSbx887z8dkcAhqIVSWv4U8gdOAo+c
AD7fZ1jNsxewHSFsZJdVQgug5+Bac86mpmkWjtxharv7hoJrP63Jk0a1vuOm0g6i
zPM3jyawceoZQZOob1Qx0v/IJCpl+wPuqGRXSjYfEYxPwIUpyDsGnZ8bEZkX1Jz1
0rgjyygf2DZIlj9+M5gTkHrcytViApAmoSfybjJIE6552ff19AgKnNsQnNyaK1Xr
kOQl/f9WdYi2qLIb1ZPOup8jjDE23B+ecxFTW2+nFFT9vv6jOtB4IroCK+IlYmqL
1r6RBHmiRg1SBUdnUFYz/4P9R4ErBdamBHyFG4QWU1BzTJln0rLJd1no4+GeWDVR
T+eXlO9ZjoPS5IqZa/F1ynXrdqNYVzSxEKHkbtjvpNS3W8RBKgR0lv20Qd/8jcMa
3FVtKhRvnt6v5n4U2hAB9CgcnHRXiXelytgaQwgiDz4KvykLbVKiprktQPiofNVQ
rxNvsXIzq/ExbL3YjxFjiG1sM60jyd63MqA0tYQ1iB/vDfCHPxfTY4uKd60k7Znf
XeY78nQlb56ICnt3U5GBnP79sEZSLO2yNotueFjJMygikTYOH/3vIYZRYJbUEcUg
cfJKQ+tzuDKvp8vLFD/02zU2B9YOkJhO/J+6Z6yFscHNmKwrv0Ex7o/2P0uS9auA
+fyzTi/t5u8SfBOcIoUwiUkxWIQJYIb6s01UAQQ8x7VbQ2FOQB3HaugkDaQRW1P9
nH5dlrzAGom1RxsUpDExtp6iOPrEq9Zb+WCfirNSbLC28Hh7Ramh8sxzNbqtqvjt
/ocblxZNhdqh3nLrcl+ui40cN75p+Uzk9h+eliI12BE8huXGHA/Hm/qOIk/yCeYe
rKsH3CZKGW4yFbWqVp8aSKuGADnVH9BFWT7R/iRl6QPJEUdj7ZSXQ1fMlBSGz+Sk
BGt+s2hUrgpF4skIAfzcO1ilmklKv6fY3xqA+p7496189rHU/Eer0aqXOqghQIvM
H8xmmli/c4N4C6wS+oO9o0ZWepTRC/JmOJYEH0saZbD8WWTsN4zdzotwyx3nvVot
SHIZegKLSi6Hmog2Q68pX93frkwFzbqqxC44q0k7pdfYQ9NY+XXSvOoA5Gksjwfl
sBZm1oouP92LSFqKABNBUWWiTiDpGyydi25WqlJuQEMhDoiBFBQyQuwmOmQjvDsj
H3IwQcKh21tLQ62m5+Lo8+3bf6tANXcjAwBB0uwaY4Pl01G76m7cUzw07aQwPpuw
vatZGAOH3RGPznjjPNQJKFsSsCeIJi4tXEBw5/klZrtD3frFF1vOUrrJA4b1fTgu
nRltJlWgqCD0F9o3CRVhM/9Za/qzljf7Dh0ijLvKGGDyEy+pk8klhF/AplZw244p
lDq4I7tmeJal2r8Zu7/2wcPh94tEQOfVNfi3bw3OIijSiUA+Oxd8I5kT4LuZ6REZ
/bo98+pA24CfSZBlQltGHUx7E3PNkgFqOlecgQnvtV1dgWSitVWsFG+8zEZOJSM1
kRqNkMsmwN6kE4MIYfif9S1HB5u6XvcSgu9uyExvx+KyCqM3xujhoHz7gVS4rTlL
79ltqMkVoMBR/62BM9c0+/kj9lZAa7zGcE2TYp868u93vg6pKc8ZUs8IqMyZ0E4s
DD5Pa4tic/Fm2VrjQBIMcsscUVJy2gF7K9JQpoR7TWB8GhomrKIKVt04ZiYmmZyZ
Ea2ZyEBLEj92la+vvQ5FAZ5QmGn+PLG/J+IBz3GSccdWZxcEivyYn5LbKaIR/+Aj
7TbqIGLQ6GVOTWEDu7OvefkQchdj9MrHCUWObnLrzFPnzBvIjtmOstEDDWlbJT6q
Zpc9eL5eoFo2VI4esZ11SBAGJNvn5y2EsoHzm3+1dxYBU62ny4zG3ej1EBDXtzNy
IDo/6wktxQeie5V8h6Z0x1pukvPwjVC0A8HZmHZSBlf2voShljv5EYon7cU6sy6d
8AIHXlGtWpACs6QRHxZ72PAE9niCZgZMAzuhWpB5s69aK8fx+HD6v+ySV3nKnZtu
ncy7dZcT1dhflGCIkoodLCUg4FYBUTLV2f8Sj0QdV8pLgqSaEvhc5vWh+ViEYXQj
VKtSxdK5S7riVwh40GGGPJFGw/I2Bh7h6/uCrdLSR8yy2Ooj2vky5VO86cBXOMsJ
VXm8q84qGSs2SY8mIb5XLfP5XO7OvtGGwN7gGZlXne2VOi+dkLGbwNbaQPSUomp2
TM788Qob40Qllnro3/A0nTH/z+mwit16wG5WMhCAe1JM6cn6b731rFxvWylVXipg
V0cNMvzL5fidJlnti5S9EmJJG0W0Rl+iT/yd2GFapmKLLjmp0req9mFVLSI0lpPy
K1/dxmpVu430O3cRez04xVrbJlTV0/7MuyR05yN+DJHxlCxgK1XxtTmVB8js1G1T
o3w7zm0GwntTadLM2BXqbd3IN9URvI+mxiejYKbDB1/BZdKg5vdelVJ8eNqN+NW5
VfRGGO3wE7gqW9oQKkJoa1o/748UrHdUFkh5tuZ1gzZ7UnOoi9X20cmetIQ7dN1A
PCDemXPCa5ws7/AAdW3EZhJlBE4J8u29ywXNPYOcI74T15MLmOF38WDY5amHoo+w
FB+ad38dzi/ssK9Dts4hot5ZcqmUynjCM+/8Os40fcrlvpbHCQ52r1hb/h4y6UZu
u2lHuCjuAaajo3EQv9WUhQQlFr/JxWpkKAyHQLtQC9vysJec9GHtpeDY+fyJ4d+o
Adv/GHvvix1KKH+y0790Uwg8NKp0tQiGDJ0JS8mlrCBrbbP+ueTaPJnoHH/jGDUf
ibCP4vHOMIG0CQgUYfNmN6QYeFmQTqcRx2y0CPwF0ezxEPsSRx6D7lLD3TiXJvtB
yVg0rFr9WpG8FmVbUXv90XBDeEVuLH8lWrZt0qVSXsBU7kgHYfDAgPPFtYxO8hs/
YzVUDgzoxWoxc2uwqtC5Scl3ydm9CkYim2VlpzTwyLx7wZAlqCKcAsWmJzCAl9ep
+p0+hNOIlHLA/yOGjd+QMbrSwP8hlBMyGQ71nO6Zy8ibejLUXHgZ6ijKxX9K0Ckw
CHcVcXDsCz2eDL413qGE/EYNsQtAU/A0zvzXf3BpOYh+Q2vwQn+Vkg5DQncx/KDS
jE0v/x+YJCjmcK9JoU/GM0qsuQ8tUQZLUuO7zB+I3YzAEx5K6WiD4BGVdQhPvOpE
eF/ShincdvntpeXrNPzibX16XJcZURIm7B4mH227Sf2NfRwWD5nAWIuY+48+P/lw
XX///Y/pjNFAm80R1MPCQ2AeLC9isL8Pmb7/2VX87z7UniQTjaV6leHmTL/+WjL9
ojVk/IiQ9DEjwSgRL4ncvaIqxacOJqy4a3Wl/7RuMn0Rc8E4aQg4moWItDgR7q9f
4qS0Xzq3+Yr+/prta6MAnPw6ol6HvCQdg7D+lJjrwDtXnKDAd3Q4qhslYd004VH7
klZR2mScW0/g/iWq+Hzv6twsTMmAuDdUcgT6VVHd+/s2UNPCiGyGNY95ojl5j2VH
j2QKrCK2TKJdM6aDjT0EHFwUh9eBOHtwuUCW1hrLf+P7nixu4MoyjA5ys89fGjc/
rp3F117Qb8i1Od5ewCGt13jnpVDPTa1ULI7d/0FbMoSw8cFiysvAOCINjEaKBuK2
QoSJOJIOZZmg/ge0buvF9NqQ+zDna7sgFB4IVDckQQl2KsgaJXY53skpP8deiH2C
XXb7SscFG3xgQmz5xsWDVtW/wOzsQei8ntgwMtMA86VPI0KG9rTwMjwhubUYNvL+
rbFJtZzNwA3JDzS7F+14Ym/H02sptRp5McdAqneRd5w8lHqJ8IvMeOrffvIWhxhk
lPUzFyqmYVKk0cSA4kw7PPsRK61ecqgaooGa9NT2OagNEtqDnAeeI4K0rP9VQpdc
cJqgyiX1w6mGabSZN216BMZHAH1Kh8gcM23h/jD1DhVubs3EI6qMTn5oIriRJBx+
QJCXrYjg39HtQHwqFpLYs0DVG5xy8HHy78U0pLJKAEcoulPbFJ6kW8dV2UwzOEqJ
fLuJwnRHKO9aGAeilKjxhG/DLfLnMadc5xw0/O6UGHBrR0P59kxbG763h272QUwT
NJEI6VBMTQVuBGu6YCgBEZ74TxopSxjAC08b/1BhAltxfRTbxvfhty2mfe0UHTyJ
wj1ranuJfVFUVE/9ZIschSiwAzsPjzkVrwZ8GgJ5zBVM5aSOxf+2x65AFY55KJ+j
l0OgU7NkfFjcocy5S/G81piPEh211oklTENAUXn0NSTSPisCKcUH//LEMrDzGxOG
NdYes8i54MomgbgqWSE6b5DoXGVoTC23vmkKoUvXsN3QWmgivkuTzOzcbfXp0pFr
01r6PD/NyvsFMkwoDSz6XX0LXufrwayxo57jzNX4rJJxWx6HcNbsucubW4yizV4Z
RD8NqcpJCRjJ6IMTJLXsraoagAVT5/WKzZqTDs3v5br8VPtrBTAEASkkTBAA6vFk
ENzBYRWiM+eDn/fVqiTxe5CsHjyP8na89bKj19mA45+zsz3TaBKKyoumo4GQ+ybu
07NOtF+HrKwjIk3RX4mLihGYlsyPTXygq+KTQcD98VWE4jyJHkKFaTOTa/fqRjIK
EEU40BH0jjdtbAhQYGmY2oy7aN6aQ7X6GmvsCv3WwoqD8YTTcsi7XcOznh4KmaeC
Lk3wkEkMVGLZlMaivM7fRro1gnpsAtDShSvalqyQQE7aOL1nvAooKO8O5bfSI9kX
jc/NFH5jImJ4qzxWrfCbbNATBBpqiLnwuTWD7DmEux4+HLlR35L3/yJ6GkY149ss
M2idpc4HzO4y7uyw/hErw0XaalXDP4Pd080b4FuaXRZ7Rlw2JkyFBu59Sv7jF2dh
Teq+sk7z6tehuk+eCGKxp5dV9QpJEtIGkeeBSuHfCTitDKdPyEGdgpUPcRnjSw2X
NxJ4EoULLsJH82VBJfJSGttezWEnISC7hdoUojbgThsqL43S9pSz8Fj8YwuBEuM1
5IHPtTG4XpP/amEGPzjmucKAk5evU1pn4kDAsSs7yZHZRvLMDweffQpDfIFHK+W9
gAmR0hpjXMLhjo442DJMf5Ye+7QwwdE/7vhCmBj6Q6vaT6iqT4nJt0+LWmuquGJX
BOrj6izhrJAS4N37cWsivCLm+9bCLGMzZShB6R0h67lPdL4pV+RP7gRNfnYY7Mol
xxS7Jccm5WnrWY2VnYNZbA8k86fJXiHDBhrDIQHFbYW29GkBML/gXOSt6yA2SGMH
UiIgiY2HKGlyqSEzxgSdsHe5q2BIiAvcsDm/GAM5F4adpb2yjarGXhn2RySIEeDc
Astmp9O/6AZcxua2SWZCsykZj5OCi68+aIqPHYEbXj4HrCy90GdR+Chsd35ZiyLP
RH9NM9evQtxsXwxht73VmLu7NmBzi7xZUrYJ3SA7sisvOqR2omzpPPQOM10gH+qO
Q/1n3lBX88RlKcYQE9XksSlVqSyA7H6qpXO8SLizh1jwmv4SHfZzDCl913dFbiGz
QhmR3AwludMPggqfDSj6qu/2yAODxhlSJ95ydLMTVYVHGVBr2bxCueu+rgjPB9j1
5Q2L+dw1fvz0cQJbNpXgwVLWa1pTf5MENh9FUWzdoxpJW076BvQ1lDGagKMfMB5+
wybX3zJyt3Lq19NgMon7Vss6F98MzO2aSj6pN1RrNQw12gJ+Xo9GnJsY7NaQu4+O
9c6ZJTnqgABgba4Jc87aht9Lox+kAkEfdhjOWZlqR7ev0eyzmn6bLtmB7I84MnCF
SU7uIJNpvzhd7hsvkBBllay88yi4GcAOPEVOPQnSMHz547tyZ7gDkAEezK+rysWA
YI1WfHm9d2TskkqWPgtxbQzqtBAntsac8TpF1mBNqPighC4eZjRhS+U8vSSVFJDg
NBiJkC9Gk11KiTwyOGGFNIgASNwRaxRnz8kIwMF7rgqOTPgWd48xlH0TyBnaXilo
pYpgsjFwLE0PHlg990ITTS5BK2Gr66MrG51qjMM2AZcCp6NbnMJlgPkctqaKVTs5
pORT7spKVYcaVU11ii0FbvJuR8c1hKlmPC05C0zls1esz8bxP0yXqnQXfXNFR5yU
BRdD3YEBxuS0WW7OsUem97F+41Z8K5iAf5IwKMQFUub/RcO/Z11PSHsls3RLrmdk
tCyrQhQqW9Z9sOBnLVqdOBt8fkNTJoat4jJI+nRc05bk0kRtLLOq9YnaFcvrVZo7
Ve0dmI8qfe3UQjW9rRkBQnGqbnh+lFXGLRV8AtArtTh7PLQclAi/7TW0DSDoWq6Y
2Hezg55PNmKAECa0dFDeixjuNKMkUWc97OrPQIqACFK0vh6Fr7HiNtdlytZ1lU4l
Oln2bD3lpFyC2xiedUX9hi1ax6CIIthdMQJ/sq9SBTxTKoxaoHyoFVthpmoYwQSx
N5LHkQugFOlmy3Vb1YUY7M8k7Q+iSkiywfKF9RYjcccrIvFLIuGF7ndILpTEw+j0
7GjPN6ojl3UK+2dvYWumEpaxtWDgz0bcitjYokTqGKuJYqzUeNOc2/EsNrBSCFev
OCEKQAOITj36mSSDqAOvKWehm6OJW+maoZOn27fppO6E3rIPh9vTxauFYclIG3AQ
FH3nq7OkNWDjpnu6wczSiFda5qQZjSyF8+MrDPCa6ENzKApvXgS77Eq6rrcK1iJY
wGVdNz7V912yFPr4bPR0elVipfwNrICIbHUHQRk2gAHVXAomGQs06Ja8NAaCGQBF
QY5myDuYTmmMuoLa8AO0Ea4nhQjS+5bj3r4TLfB30lVu4hCwha3nXYjU4Ak/Ojlm
G3yH5p/mIWOUDK5yjoP6G0EM1uqHMl/1MHvhX1h+0Ry01MauTcRqHYqRrKEq+1Em
wJBtYjtYESycMTnWu+F8qJadDf0BfK34rMjXJpu0y7g8gm3SdiCe2MEc9RVsoABD
x6GIpDFf4cHnD08fhePOWr6gNeVArQJwfQVoXzukoSOBuaDlOB82Pnje92CA/2tT
eaVccnnE4NWWgyDbAt+vwAKbgfKjAsMC9o9fel1lsil+xjGFapLyV9dnASEO8Vm4
UoY5lgOMbkQD178V9kVDqnEZSyP7WUREilCCQZPBE9qHnr/CBzA9wyBpCoMbVkxh
QGNRd1z09FSjz4ZcxUal0Z0Y7AffE7uiepCHPf9NRzNzitrQM6jvwQlfjOrpv69t
5Qz0ndepAimuQbPUTHgVnrEzaWjlJTQ4vNhnbFjlvhoGLdyhUbQB2tUjAtoOqTMO
yUVccGTDXVY86/AcR9iDiotDlFcN8jgsoQ4h0tEmN5oR52TcnyDso+px9PH+m+Xp
NxdRJqOBO7VcGbLN47pK4eW3hGap3V5Zu887UdneH/H8bFT72x55fTavy16R0R8K
Yt9AgoM0iOCkQUr07WbWOS3bUGKSI1tCA9hU8yA6nKgFKN2Jgh8od+hj0aZfhGlU
3Yi7/dFHFUHkf0NKCRj24fmt2edgu60EyXiICL+CklgoCRQKdMsOs3PFbsRiOPh+
VaNpzdyG5ukCs3UUFp6RyHNT+RfX4tTZa268HjYkSYlHbsBUYJaJ6ZbT3ETQLblk
qmTD1Z1n8A6cSMtcfF4N8BZReEraIqrvQymmucU8qFwpbdPqF/nWU8KYenNTJT7X
vSg2clFNJIC3fM+6O1Q0kiyOsBP3L2/7tpcp0iiLDjYk1/QmzHiQiv+FROLcOr5c
1ocAmJDxp8f+nsbz39T19F+MFpI3+Yt5xTDjmmGmO49eUy0uuDKLN1ofFgIlffII
0WBfP3V5teF4HSff140LUvoUhJGc3lD4bpeeGyUxcTmSemQn1JMUVm/ri6SR473Q
KB+U2wUOR0yEw4KCXEGiMjR+5WYUOTeniyt1AYMMpu+7FLlin+o+Y4UtyP+fVXWZ
KicNdvLMirVd5XyAR2kZEf/VyVHLgxnjdZsv+ruxOVQ3xUrwSaCByir7EcSWO04q
niYZoE//IPwvtl6ZnE6BjnMlk323OPntY0y5TXfjaA7scsH/WHzJ2KBW34DKzD30
OuaLw8OAlCG9mMQV7zkouotzdQv4xYzvI5rGzwVYXwsbIsgy7ZBht4DM64QFtgEs
gG8iC6aaWuQnqqfbiZTS0SeT8xkR6RvIaX4Qbc90ZF0yee0gTHbEG5KXF5xnW+cL
DEDT08vCt10qIlTVxJ3z+nwgL5lt8JdkLe3ZREL8On9+AfoOF14PtOr537cUAQeB
pqnV+zV1PE6mNZwzVQFwFK9BHQboohQM6pWt2a1zRBktWdmH8WfYOe2sJMqF7c4B
3cO1NcEr6BvEKV+R+/4EACAjgRS9r8zXNf20Ptwbeus7OOb2o6klM7m9Ya4PACw9
X/8MdUmOJ+o8a4ZA0GSjPGtjjYp9DUs710M2dq3Jo7GgKgJg3WbIqqLcKWIyMb4H
NLV5Sj1FVx+mzV+232W+sf4jECUpTg6pFZZwbTaP5/S03KnrQyEgRofi9ejXoEFZ
cFncEH2pD8U2SkeOGTs06n5apNVfrm//UobdssuWJ0DazjaFyRFS19E5j9Ql+Enp
AHJTWTpZVpRAof1cedNNJPyUIdmCf6BK+dbTTGJ5dL+V0iRwSJ7IqScqzAKwUUio
wmNj5GR+Pvgplhob2p5ERB26KxxgyKVNC3DaHjbA10eGAZ/vqR+8GnAA4KX10cIL
uHyNoRsYdViMcB9jM+C4IvpFcq+fJ0srlPRh2gtHp6K0TGOvyPLJ/jEnH18C4WiN
fQ0nziXj4EMqiq1aohlro/JbRXQMa2+jNvKhKZQ1A419AlIOa/L18jsNMIqEQmaj
OsPqb+ckRpdegJA1cp4DQe3N9x04GJtEvwJ6lEgTshFPMKTKX83iXgmA7au/VKGI
VRRxnchMD9svhq3c+BQWV9HeERFM6akL+WHo8NpKEsGAXk2SpGX1ifNA+FcDfO0D
SOUdffADp6hY9nbxhadXKwkWTk6kKBN1OdicC+OzLK8DUtSPT00EhNelIxDxHoyr
jHCSPdK9H0Pk5EAWn62+pu6FJgmnp6Szv5yuEH2bjMLmrvr6PcEOc3E+xPXamlTJ
Lv7eBI1zKYEW7m+tCuNhSIiHrpliLsRqB46Th3qY7NIUNF5oWXeD5lIdL/79nhjU
AxRw6VMZ38NV0zKofwWgTQkMibWnBbRknJWgUVt1pPTntb/hgFc7dlewQ+VYAbez
Wm+IFSGp00F9TFKX6Qg1l8sXKcjJNGjiIA3BayZpWCWZD0Df7U2lZqMCfmTYk26I
fgZ4YfGqQyJHIag825Emwgy0iXhUWPb3jtGN4xi4A1xs3Yz5yCkPuHZWtyvSXL09
6tJx1u9EhlW/pMSFXpXCkq3KZ8L3WMEf6x/FGIXlZ7LOM/Qs+3N5IN5xiQcnXhfm
CzYPkQK/loMOZOY5Hv/V+eMSyLr+zxU8zLvKFtde9OYpdKzbvbGuc78rz8jcmy8j
kPNCcHaK6iI+OdJIWT+hGz19efqfx/x9HF6HALYg6aca1PDhw5BNfSp97PS0N7Pm
0N42O0hyJhIRLcc9uM7vnvg3RduzqJsom4QGZY1QYi46vWC4aIlVjJn8kvwPdcHK
qN6wAyrv7mUTPKX8iXerbiF9qD5cXu1ZelAVVbZ5iotiAtGjcXPTvEHKSSS3pYsu
x2WfyNKQdPIC5UpLbJl0Ul71Euo/tesQDKqciZ5DR/DRsYO7grULsnbWFj0yrjFO
x41Aux7oh37YaHL94q8qNmi5KvmAUjaj2+Jk3kIB8/+k2UEjiM15Cjl8463iSPvo
QjQl0KCAxY5GcBBr5ONKnRnvq74/OEN1vTq6mJ7nRSqS/nAJxYwHk+acgSypmsDY
GpwMVT1Um7Wvm9mKCTVMXUUMh5+kdNvkiLP4ya1knwNkz/xBvXKNfTpG0MLvVaWN
ygXgHmKMNGKU0OyKkzBjKIh/Ag+pj3euHliaGAfmJ/T7nvKH4FNC411dbuJ1JkIT
ZW26QcuuxYqrJNkn2Mr0yxiBbxRGjNmedgaDPJFOz4Wkr3oUq7UuoYYVRGZXK0Tj
3BLGk6/86hvrZ+RrKY5oiZ+1L2cP7xxV6on4bB5mcEP/qs9bsc2TsOyoCU67v0AD
weVOXCCDBW7qy2J4oq7xuaw9npKbaTtriSnCr/w5IEFzYpz94vHkfdlDa6qzeAm9
N5/6lPDsWOZCJz3wuav/ETfM/9aib6TLkmJjh6/9oJn4gLipVsw9HBMHvnaJOgtw
IrXAAZIaBrgrWsQOmD7/6Lq10KwlhyFuTOR9kCP3hkMtQJkTQ1Ngh8e0xqrsC3fv
5biTi9eT8QPbvDqB0CKcQl3yeu2dIzVFKJcWA6nJhDgW3sIy7zPScHy9+uCKf4yG
WYL1ALIoWydScK+utKVxenH3oDf+N6wOikvHA9O3oavbl0k2kDmDTvVQaT9mQFYG
lCo1Rto4rIecm2ubBixprg+Aq3LEI84Km5hYUoPTx6dwIN4baBVrnoDcQK2kYDkS
QRP+NGJIqP6J8JlDkXKYUQTRMZzDwFpXJPILgUPb6ShVIIxch/yxOQ9luB1aCjG7
GSuqC0yVGPsciIbaODjTdBp/liinR3g7epf4bTAezTx804dKG017V+aRsENXYWkz
489qBMSfUiQ4PMR03VwrwFAW7QL6p9X7HAQR1MkwOftDq5rlKxZUMqb3h4YP7RCP
g6P2CO+hE8uyP1id/39/FctCcVj7ONHKjD2ixRdY/MWCZyDpmaEPyFsNYSx/5bt8
1gyBwEU2KpXiREezeZsd3g8gY6WbEPpPOz8ML7DOtXS8J3a0cXufcBiftN20Hcdi
a0vo3eXXRT5VTlJvN/6QoS6L9JSMVe/NTAArGhoNO0P936DzNhngi6NzlaZFHGJQ
7yGtRuCxAo2wUPqZy+h6UrL/GKiwjPdLa0oq1SwvQX3bmsBrQObsISGHoRUEKdr1
YspfiCruFmaP0SrVMJ8mtnDMHX0/XXcmYhhSsS2quRb3RjbwntatdsA/sSvw7UQX
pMWqNAmZgxaT1jyPk35UxkMx5J4rPh8zXBkx2BE15lCb/SqEgRwAbQTs+7vgbBEI
sVrxEB2sskIkNU/93OUENCgjH+JvHwLwIBSIO22zF6/mQy0rhHiFxdAJzzU1LwjO
vXdqEKoCWMzzbTFKcIDYmyR2k2BpfSKH8g7u6LtVtBoLsfFGmVnUMQNmkEApEbi4
7i1U48gitxHy9D9EnAgn+buVBQU9OBwExZHRKcgKG2ngpom/uh2lE7Piad6vIulK
CJEcChK6rVuBxsQksMCPrQ8DSLq+3HpyPRepmXTWO405Stp1XHP2jAWGSIoFyiO7
L15S4VhaLlPpjTATG1k9BMMg+DMK3f7o4gfmAhcjheD/gf2PQwSfVrLJgoSvZjN/
c2T9NV3d4Vzo5ihLMdV7+I8Kbo0AerdL+khhilmc4JhVwKwhKDWjxXLQvnDMlc6m
IT+l4cFOdEkaherKBC1U1JWk66hluitGM2aHg0gVOUJO0gfEp4N/QfVC709gfkcI
WHYb9BBuaMXRkV/2zKB6TMmcoWgTwlyRnKUljkC8F8lE19Bh0Er4kBFdevKtB8sJ
yp+Vb8+Xc6JgywMzCrao1BgmJ1LFcrdzOdWaT/Kltb83LoyMWuTw079r0YXZk4WC
Q8kUxjdpeuU6ITwPfkmAn+yA9OQNEjQoPUU/U9Ge41r6CmoYlhuBUIJb4R4HSDoH
Q0Q7gDCHCSK6NImRAusk6A6q2w5k2R78uBVGoqUHIwVCCvLOa61nJJ5LCdoqre3j
56NwLSbtmlpw/O0U8x6+GcaPE9kXMEHZgkjX3ljxmYwEOpecP8FRM+ksLzFqB/+q
//SkuIc/LH6mO8SyCehhxZvrvGPuk9t8oYqqNOsIN9DQS/qsXPLfJwWlcs5ztJPO
H/98YwkjZgVohKtV26nOqZljIGj2RR4/MNUytUJDKNJleoMSxnqv8NOuiA9jnpK9
xQ20jeR2C2GS09x4MFEvzHXuIdsDjZoKCYlI7I3R4T83drOJHru0a43sKSqzRs2r
ELl0rMqioj54uSE8cxArg33+gshMLb0CJcZiEBm6PnkkgBj1VKiv06mAKNBuXwzd
kf1Crm/AC1JvNe4si1UV8qNqnEMa9TMWnifHBi3dnJU2A9J7dizCp8GDliad80De
XKeUBA5OkTTHR74FPloX33n8Z5ZqOo7fHFhe3fumPqPPik8qI5jZ60tDuy4acQj4
F9Gw6KMoW+WXqzO7bqf+yXp8TUb00cqYW4Jqnw+nGckUccPSzPKvp10Q24zftmCj
wRXUJLhPThLmF9IPoM0N9i+KGm57ajNHU2pmkPnqwz0SvPEPggEgm/IBckrPdmU0
ruW0HYfEac/0Xp3TV6MgQ3EcA0ih1sD21x/e3jiiVKj7Tnhd2yXny3gmvJE6GYZ7
xP9HXpTwyYf9m7Tfzd8T7XQS1Vlj8Ia6QFDzHSdlIxWYu/YYTYaIeAJXo0nDDogo
L69fkes6z0xstZQ6BescJNVfRPgBw2ZOb2JpUaOg+JnfNWwXmu3LF7R8BULuu52Y
Idm7UakOO9CisymeGDlXbhbdNBPtxS42HDWJJ7QIViFToFnztcLfok+G0obi4UXB
Z5MewwraPmlWq8HW1RLpBhtcyb4rZ3Xlu5NmGaRmwIT3UjIOiXYzMkgXxjzT+LrA
V63SrE9PA6iPVzNur1z64SbjDLucG1S7ZMc1/7cuDgCuOFO3Npe5xOhzBUqy+X2r
Ff6s6VBVW6aXgW7LkTtXfq90CTTb8Q3ziicugNYUJ33OFUezsxmb/c5M4ltMp0bZ
o1RR376zuQHQl1soCVVSC//EuSos3lnhtzvA97q705WXgF4ee7B8VgeB6ZS00ALw
fnN20nHi4ltcVMdVwgAmwWPLoDwPhBWBdUEPoMH+zdNreOIrivQuR4r5UCHyukr/
fIkuKa6i60w0QtlvoOVe39R2P1WijYdS2K6dy7i6AnbNkATzcNodcqj1BkmID8yo
I9fRxU+xBxo7m1Hm7C1GwSQp8Zmr59WmidAsoO0SLF2Qs8CsI84WnUGx2OtI3rc4
93VDQShv+VZ9vy7hLO3hOq4hdfkbSljZUDFvJCR0RvoxgNlA7OJtdLT6riDBJpzL
4wat8+b0BxPm5azP1mgOf7BxfEi6Ge+8j3gXwJ3gBi3tQKvEaiztKaEbTC69sLOv
6LahBa23/LyPTWjSDOEFAzC2fshST8d+f8QMbH3pgX7EbEZHS3pV9iMjbDrHS+ZR
bXbdgCw+VA+nQa4F4kZqnAkGTwy6vpswsoAguUCO6OQhbkW7ELgYl88jk0chTqUW
ggch2R4UaRowCmb0vUVynAaypNC3QrMr7k+z1sR9S71cOggEC8y0EbzRJWsQeh4b
koMQbBkUmNvcz7/JfnCL6gTD5Drbepr/3MckDm2zas89Z1k2yh+JbjvDxn740vlI
o84KMskFV+ySbco1cqsh7SJFXevx04ofqOWer9Ckkm/lFoPO6yf5iVKxPqBseIM3
+bWe+CA5K39MDW88SJAN9dPIortdbY8DEU9snygFzbOhsakcPciUxXn5Ps3EKKGf
7KH1P76WNTg7KiaU+6Kc122kiWi2lS4IEFaqtPQBAg/+NHu/aMfXOFbJnq+nJxlA
RB9XXa0clJn39NRSGR18tR1+sttJKzh4W8CVN0iGQqRLuHt9NiNSY95yzJSqdaaE
2SFKtpCOfzA+ZrMkfuU0Pq6hU2elHepDWyKZhoMwOES39dmY+Aq5vRx7OwVEzvO2
wykK6eocpCgrMsKSjXE8ZZSPxy9tcXR7B52tF3dg2IauTk9v1xVEDpazIP+Ky1HO
MM1PWAzdtUICVl7D85ZDjlLflnGwBMSuAjOAkmLQ/BuBSl0e7dpBcBrSA86QLo4d
freC5S174eNhWcEnR7vEXdT/K/+bxZevMTxxx1McGNBRSSwXku+0k1TXBdKeAlTr
tj5nuDkeAzEZXvOw94cvgW/GyEwHoLaTQ8tqBWC0u/5cMTppudhBFv3H5eFkUBHj
54umJd8FHC0WBjIwk/sPoaps7qLjJiKebLoB3EDoEPToz1aF9vCae8tmzEd2jZth
90EjFptMBmxybAwaqoW24yP78+atSQmDVxvLf1qAkVuIllCO411bJRWijNoKNvGM
M+MkE4nxeRfrESjD7SHDvjPACOriRiS7WCBFgZtvxpfUql1RgIfhh+zr8qIM8MDH
aX/FbH5XhlFJ1Vh5Rxj9+PbDLuf2o8YEthHUmR1YWiokScweSP8TWmQIRSQ2nQP3
arGjCA7wE4MdKD1uAqWtipJWuJdn0Xl2v/F45lvkLmVBXg5k5yZN8L1tgXcgxKsK
aMnvWAyxH9sAR7xWH36Adx3LNjvaTZKWSNRWshEUueAKsszKfLDGNeza/T3VoNqk
zYeRxsyAMUpa7YoW694uPZDwnDgtNwvTnE1RsxJeUydOwutK1UtAugHVy5ZpxPd6
mqCz+o0jlI18VGKvnKkOJBfrpq6Jr039r06CC72reSgtb+b9NJUq7P5FKFs4FSFQ
GanDW0cKZalaUgJsgnwuOFnydwisa6RqGqNhtl0spOZgVQMaYrIu0aAwrnPxOHah
Roal+W3SaH7O41pvPY5YPddQdroP0VCxFm2qOTJ5HewdkV9+XNfOPCOTLzsTKpzi
sGetmXhVBoYKRiWg0PP/DGvPTC91fNBSZkZ5JPtEXq/Rqt8pfC5tZ5e/175dQKIt
IONdYMl3oCgBe6V/SN1GOukLmL6lKkDWxNvzQQ4BU6V9pgtYfBQ4xU9DA4oCRIyF
bw9uDx5kctNGAew1CfIvVMghM1ZnF1Ru+9t7R2VLDLRSVfY/FiNdyov/0Bf9Btfg
WAmpYaLIb1eUm3HPPSi5SXr4h/m+odm3TbkxXPEOKE4RKxBO6O/zjqYgLhGFbt4G
W/4v4R/4+4IvUUy8yhQ34Vx88ZUlhT7LvRksf1RCii/tBtPJ7Nxqxls4BE+5mJOh
QzDKqeEX1qDkB1a1EflGyggNo+B4rd8uch6EJo+nDWUDmX4ie1cYUv0loE3z6Gji
RR4S8/+6j2x6WA7I7ugtPcLcyixPSJtpA3hUtJxPEkfgCmi8w2vKD9PD7JskMpHu
ixf5t3o6T0VmhDMW4Xf03DumDzrpS053AmiuYfWJ2QLHPSxYaVbC652xcZy+BeSH
Wkibdl7fGhx0ywzpY8p8Yy9lOr2Pu/iVE4hjyobtq2SYoaGcTzF0rT8DwFzSRYN3
QaRSHw6ca3vCzcM+qCvxf3jhIY3VQ9AvaR8tpQboWpMeIGHnLqlp1Pganpk7jLc9
WxUhIylQhZrjw88IpgR0ZIhllKE/wjvEDdtIzo+RQgQe7D8HKwFnO1Vb+ZgRXJ1r
Y40eBuFudLYomJCb+HpQvkYZWXg/gXDr8vaT3R1y0ZShiq5jZP5wEmEaYWlVkI7N
Khwa80sOigoY1Tg89Hywq62Xc86J8ThgLQfke2r9tlECjpUidaL69Tdtr7ZEaJLj
lImikSSHIW7aawkC2ore7TDFj5SdRXfqPJwMey2BH3K6E6e2gHIUbrj0wDJEmniL
52lbghPcrUtkHnCNzUTM1BJilalN6XfvhXiBGEmgyMe1VpfuGkRCmKCqRX8Eew0P
UyfSP9KyN4ds56pThc+8VeCpWXS/oeocXwrHw8Z9p/dLHJr6LqW0A7KekizToaCR
7n+c5eD1yVcBUgNar/07CRXllHNYDGAJU+KmiBgewYSRzbZPOs8U9PhaxPM0bWac
fBuQEB3mkp0Q217rV7SW+pIE10BJeI7eA6v0yVT/TTk+B9hlAl842EeavVtT4YCW
KM7+cuxYteJ42Bk7OMoyS1Qqj5Vmh5mMv0gjYnVO+5yMveCLBbFukxQsAVHeuxXh
IqcKs7+4wDi0PItUyTndr9k1WUMGO//N/EBb7d4IdG/pL7EEBXmcYnhlm3vByXYD
xopq2+geA0EieUnqI/1iMeEUnpuI7seyTY7hyU8nilDLnoffA/J4U7BjVkc5rvQ6
7S9VKlJM/qERN4LXo2U9vx0bvIRbSRYAO3ZcGCeCKG0PlZm8/O7NDlzDrqr2E/YL
xsOIUQu1X0KAl/W0+t7Myw8EFginEqG1L5tAlyKBMvvufYEhGfL6hTp9ZPqRwsPS
QaZm0tTHMYXWWgjFd5Vf1PlmSOQ9uJlUmtIsEtK7zWZ1qnmyuC2RCzYpiPUFSjoC
XUH1AIYBwCcLVnefjusTnVcRzCj43wFITGx/Cquzbk0ngem2lNaeDVH7Nz6w10Ne
m6J5WnDxTpUDO2SQHgCLntjtSbFL6JwSfS7XLHvwIo3KGUnmuTbnF4ACIL7CjT1I
KU1ExgTCLWTV3Xa6QC565trV/cIRTxLrrzSWmI5V4dtHzqoltd+9gxoGkBSvaK6A
Dn0TlA3jJCJvToJNseotYxqbiqjiYZkrfifFzA3rdV6683VKM5SnfJ9RS3lBgXg6
eJbMLr9ZfHV4d7SA0GhSUzb+qxLXUXl7b0I0XyO+sfzfYfuMcgFmnLmA1ic3KmtY
HHWnsEEAtO2tjRZo+NSl6mcuAW+TV/+k3jYddsQA/+phCHeXePBodk9+Mx3AhxIi
owqeSys3tzYyxhLvplE9MqE/Fz4qwKIMJ3YBla/pv63rZpwiVZpMF61FVF1fAY5P
MQeUJRwW0+nsuDrk4Rs3Jog+qgPSqTCLIPlpPTnnNNrJ0cKg3nSyBaab58lzBLPI
g2cDxHmWb/6tvRoooAXH1pNttv5JbWefYP67ZO5k7UJNdLPqoCn9gT9iSTDiom96
SMEcRKW7Rzxrn50IqU89VmPqB/cUuMYihPvYCqA2AjV/RVP0BptfD/a8whCaGFhH
ylzW0OVD+yugytHi0g6XraA91SRbY+fE+sOSnxYc2w4oHjI+b1P4H9xt7/LnWbsF
R4OCDWW1R/XSWYZQMVhDjNTR9roWKyddtRB3EsPNHkkJTt6wzTTxQ82a5zewYICu
epIj3yCb/rNcrQS7hkWf7WvkgZqjCleSOOvlhtbyYUltt/3RYmHUjuT8QyELNCgz
9fuVA+aM1o5R+jJ5e4kCqS4PLoy9jM32GmA6vtKxp7idC496EJa5WMFnhmPUZVRm
NvWgShGbwi8dkrDPWAn5PSak5IB/n3KII0UTUWvkygWER7rjE3QfQrZfnH9uJeez
mVAOF5ol83vGqUKLowu9QEkl37dFO9yffdLIHUslrD/iZI/lOidD1+eAc275Hn95
R90uysaPgZ2ClSwIiv5TSV/zkKRd9BKeGZ1s9eLc86+Z2Jpvn4nitaEUbjn3Ih/6
ns28iB/BzbI62k1ik07nkSnQ45it/4eQwAxtP+HUARPcUNY7bc1z1rzp7qZ3Vwzs
Kvh7I6mY3fwgemEglga4X/abksuaF93OkXO5bUU9XK/JYHhEVoZk5/GvmP7kxiWM
3lAYFYz6BEKsH343KKIeie4hqAxvjvAJ4RaAOTwi0wIZVsaV1eVoY9eMfD0WiMy4
kbA7BbEhlkEhHFWGXO/l1LmOxz1cTi5rh+x6x6flAG5MCNN1ObMMcEdsbzoHDYdV
nXIRXtukUiLPGsu4MjIxwWNt/V5uhCMqGN/K0t2ATL2pygb9zAvcL1WiMIOvH8/s
2+YI+YC+uUF8svdpRoOCREWrTKQm3TfNPBB79LmzdsmPVdJO/mrudfMJJ5koU8lw
mbOub+Ax3GjLvRAtaM0UpWZ6rodiipzGm2P4MCZfenzFQQQUYaTUYbktf3b4aqKt
TKnDeJE/bw1o87MkdhFKNU6lZbSK6wqGj+UPHNhQZPcdnzt9bnXIG9nS8mN6OuaY
37TVjxnPk3iWoEggXbijKSxWaGfp+PUV4Uca5djYN5kkEPBG0JU7yFQ+99lSegUu
dpblczyueqwhzuTtjcuqsEC4iMP4dTlH/XJ/Q0xE3CatkrwE+OC+AzXs9x4qwv+q
/P6AZ3KHGjdUG6gi/WaEWDC9pQZrSlUXz61o4XMsHpdI9Kg1T/0LN8AST6xuO9Ys
iqawfDPfkfWavRU21UoidVzxIviStybYizTK9G4JTbX0AiB/fqgcSezoQ22XjXcI
pQbwQtzSzKoGvgk/XhX7rTRVIIQJFQi+GBcxrWYN8gNjafTrL7R1qoyFhIX+4IHS
Xs09ZsON2XyPc1sBb8QpIdoCLaCC974BS5XeWUSHU47HSQST6nbfS2SQetcckk6i
7v7cWMbxgS3VoMik382e5vjYYNfttRadnfMZ7uFcg+x6dn3KdITAs0xlbnkvfkDx
eZv9Ey6JzkK1KD1R2P3PO3qVo4l3lQ6JHfh2Kpp9KY45BOnueVAdBE0Fdb2kaYgF
YfdxZ0TaiRN/G7NSQzJJKdPNofd79vB4D/sLkZ4Cb4mqDoSnVLPQYFKYZpi3SuEX
hOQy+GA9IycPojcBgmd9vzN/Fws8/ec9uTRDy5IWDNRBdLy+nXbKWODjRGmtw7rW
ecH5Wni46xJlM0pbXryZDhyeGuZYre7yA6p55KipcmtTXGTXwfTma+EVwXx5LAm8
+JpV8MvKijiFLXI4tgBQWDougJlH1OSUnYZMUiS3xdh51oDy61ZUeKiKi9gMrtxZ
eNmoLYc5E/3LxHNtP1GF2skL1DlhW/DQawnOetSDKOqmBxWwBHDHjnFi8Wl6hj+r
VHzFOnTLlYTEzDz+bP78zdX1WLp/xOW0KHDY/vF/e0H/i6hPii4YfPW9922vYUE6
Zk4nsnmYnYkJQLaSVynWu2FdY6njvPd27UfYrBxkMYNp1eqAHkMJEpw81/fTCwk+
epDeoOjU6Ku3Q+QXTq2O5UxYklp/QSNSBy9wzvJXpmnYRkBkoJ6NJ5YEy5lfThy8
1MLwCaj5LU9neuFknPc2HYWRjtpWizflY1mj+Vs5+g3r2YrGw86BC56Wxo9keWVg
TrExlg90Y0Oi0HjG6xVq7u0TCRCk3Qy372UzB4RBOj+IvNhsCwqslUcxEYijSI5K
jscIvsVQW4eYDVfkkCf5luxh7OZwCkfbXsfgRsBV1vuoRnvjtQRRdY5NZGf+Xdg5
T0FQTI0zGzHogbEjwox8Ob30oI6804ywS2i2iyUh2Cvu5cMjNeMVbZ/Tm9w1jvhJ
zUtyOjZX+FWTFQInOD0o4EfkRClsRDe4drSw2IotSvof7Mwt4BJmLd8nj1oAOkq8
bACMjYbj3hXpwqSXbSSqxUULH/tU5y6Wse0BY/sSdyPDu8AOKcT5h+9kQvu/z3M9
RGJqwj2oyJ2hDgpoitbxchVI8+Zfq5Wlc35nKUMlaFxVgrBVcyUnM5VRzVi8Oo9p
p9NW93d7bhffHZHY1dZ0TowdztUKsOteqvV445ecbBJGOT8cIFarx2p5YIGiUEXw
anh/b4qDv22Og2SH+lxU5kLC1X2lK64qX6UmupqBIj7jpIkMZ0igBob+xeuwHbtY
hcGoFOF3ohuVSC4VI94G81R5FDTkeKqALJQ8nrseAN9VHW3RLn4wiW8HC3CZVWcK
cRPgLdI3AVMCIlpp+jQ/BmdDt5+9Dxp4474K+bXajfOdzjhdWihrj2bjtQDkYvFO
5ilHVoH3iOvuFOlAfmoOw+PzVhnTKx0O/IZDS58623yAh1ZBEyKew2ufiHSHV6qJ
MnPLy5bD+vGjrgBfgiYbp92RIafRKe3Wlb4RqMs8lW1yQzoIjAUHbq+Gx6MwRlm4
vkMsQLJCG6ubf43e9SGvii3deFZs50JEn9Pp4l5v2Sx36eu5oY9hBJ7OnBh7FyCr
Y5F2HS/DE1YJL9IfdwPo8RRjSHNp499CbC8By5adD8f4H9DUnP9Fo/Jgy/Tpghi+
vwkGQR2EnGevqFLn2wOvyKOV9MS6Hgwq3N7fJhiQN2op4x+DOK2kstUDdYFG300d
spMIGj/veTXn9RfAZJKxxMtcwVwK1VOmWLtv9xUpTbnIPXwM+mWwlwpJjL1hU+Oz
uGAHeOlLjtsiav3MBaUFsolMWNWORt9QLlr9UPFbthNhTiUx+CnrJGPP73aL6MvN
1zLOAndfZOM9b7s6YWBsbB3nXTWIYDhFxHVwBb8rbfxUqvUIWAOgPOfhopIwvwCs
2EIQ3IgSbR6aT4DXnbauj8PSmd6HTFrbgvYMAHMLJzCizDKMW28qADGEQjHqkwLq
W6Y9qlbQWDyBhSc/LI9t0nOdXAF4RormuhmrRkeJJifOiLXR1J0rUMn1jdYOwCJx
F0d9yno1JPm1E9RSDhQXYv1vk4cyHsGoTFHi1N0QkoldS0YfUtK8YHmmLMfpwrf9
/2bEXhp5JVR1QD0QnInNaA1LDdnvRur8Gbrn3M2h68WtvXl2Q8OUW2CT5fCv1DQb
n3rkgKoNMFeFz3GsSdxRFTTJuTErxQ/lK6m37NzosZ9T6erH9VE0YmFz0P4bJYcv
wMwbePUxuTYoG4tV3OjWHUNKR2wD9CsV4/hW6tQqrjLszt6xyTAWYErTr7iUFs+F
cztP0IpsH5jBEz8BLKF1LxgI6kcDMUMO8g1yqM2Qt9wQf1K6Fu24UBFKIqW1U11K
Z2XiuRD2kPMX0Wr0xPqCnqXx5py792m6r2lURk1N7wRkPkgKtOl77Iti+FbxfyWP
OowXPxONjAn9tIbRmaJLkioK2dO32A1+OssW5IW+02rVEMjFC1pqQIcr4jS7q92b
ucrjjKPELhkS5MVK/kHm5i9M89v2Zd+pswvqU2br1VDUWE/zoNJw1jTmzJ8BrQRZ
5A1rkDNNq4OHsImlsnyUBQcuk/DUaxGUdePkg9VPv2UIfiLEvkb9zZmGvXerrNfr
3SPnA8in/2B1LG2lLUElytHWT1A7wglH4IemJGPWakHXvHGPdoC5zbbp7eDsJRJL
XvYpW1nupP359C1xevKGvyooxnAB0bSPIrDwX3iGyUck8Lb+HrLxDjdg7Qw8OaOJ
CtuNhgjhZ3rOKsrvNO/4064rrBeQ+5wWwilutFcGSQr63Cst8j77hXe30+PiGTDi
8/NHMyNbwX+Q9KGfTrQXmxBcI6Fw/yK+rVz9lzuBKqndYVE0+YULrZJRu7jXecb/
SYsKCYTCNxra3XXNPzmU+BFtKANYPoETqWn9qXClwHy0jy6pVVq+agQzPqbSMtmg
7bLVl8Dty5RIPwmCppshz8KKhdipps51oElULxOit79BNGOuDJh2tbSfVzUUeg0S
MFZjfu0WDGSfSGoMGvYDAI7ePPEOyTxRzzTZ7xvhmVvQqdzeeHZhjpCPT9xQsDcY
omoW2GqC9AD83etaAEpy35+wp06UcuLS+lLy81KsTt7GyfDymCv+N1OdeQTuIMlm
klVeYtx/UCvxehdmguJa8c5iMYvpL6xwDmFd1PKbrSYr4uel0mroT9mQb9gtG2CF
+HjTeTW+TWp/JsznyYjB8Gbhzg4MoTv6vt0rD5Xa+xJi4EmmVF5QEtZSJlEnyXg6
2c38rxh7PCxwyWZ18hh7fgrduiPPBnlpAhrH0ZUNR7YR5t7VgtUR/nXgK808+Lw8
0GzSCPhBuAgU8e7XYPHLh28w0dFgVDlcUl9K0KHJTeQZ/Z2g/jodkq84cjjqw+GL
FMxvkxDWrhxCMmZJLrZ4vcmbvbhOKEkr7C8p/DEOKXCWM0OeWVekWcRADHMTsQ7K
hVjjM99f9CzvP7DiZy7rZAl0hzfeGjzRfxfsYA4TGCtCWCR6mX/Dws32lM/NaKqj
ZX0IV+C0oV6ltZhNs32+8yDg+030zYQiQaMyCYe0+hlhp0DJBy3y1EQ6JaWx3QSC
z5CrhFJTXaRm9dt0e5WOkY6uoMS9m/ypquQTkv078ATLGjpXZzGWKLCxndDvb/Cb
n1+F8IzIKjGjnvb02HBYj8QIFFh+2ziDic5EaV+m0CvIXFud+Zxi1SCAeFJOX2Rn
6SpWcaeF84hY/izqOjqDfowlzTgDR6COAgJUR2MjQYfwvWDA6fdWblQOkakyfms0
gPFNSW+u+KUdyCXgllAC6pUWRv5OGvEsHt9fHWYHBM/+1pWT99OQDNdB2Ugc7zaJ
amaL5b9wlRcxe+TnViHFwpNY1vOQxhtWumZ/5pe8BIlFQfkdof4qNKm86ur2k3u8
qhjQhFWAPB9IUF9qcOqLEfpVh2tb9nHLt1edic44zYQZvoGlXUUcfiTQBqvxa1y+
FhUDFg2I9i9w7C4JCKPMjtx9i5+LezvEpKI9OAhZI/fgwwLsV0ntu61wR+upYpFl
uc06WkVAHg8WEPNFPMbW0fYmWaNAnlJslT3S0GWUeNH/HA9weJ62IdpJRvFHNqeJ
COfTDnXRcMK4YJMUEzROEhtX8yk6OmaoKYCmo16JPunHka+tqioWv5KsYTqTeSHD
te1ywhuTB+mwtR4X6UzZhrizDFgbc/vNEaduKAs4QsdTtzUdhpBZ7MNgf+ty82QX
zjkjsorKjHli/guabNR96Z78DBcaWHSGWj0h1SKEXYQw9f8Jz843A9dVls5Dnwhf
A/99PFQEVCagUcZUam5quxEGrZTeSRzcaALeYiWyV1vuGMFmb20qv+F3fFfyMqMg
KBox2Zu14Fqzt3RKgj0C/MY8J132tW5N999QQlrSMM7+DK6CwZXPdYqqcTrP+w1+
PLGM2h/Ro5ezRgaFJYUX9FqC5vuAiTnq92gBB8yE3X79wKFfCls8V7XMkALcCadv
8xXM2gXpaRB6/RUJsXylr0l/j3YzxFZ9K4UPeGm4D+k/4psWWQ0aTJ5fRO6oTxkz
oGV/PlWsQ+LzeJrnPBVoA1gdxwblM3OQzYgfL+pVlUYJxJz2oH+db92BEZaL0n16
0RMg0VseP5EsDDZppQMZkUPCZ2SWwKIwegzzcapqb8+66bg1c6gPV7HqqozZfqNU
fh5b+A6BHYcDfpGVUiE9PKSPDesJnOQ0UwZPbbD0AWy4Y2E5uLwBPhflIVy4BzdS
WGoh4/MnYHx3HZhKZduJRKeSRkAJGcq9MbNRe8kwafSQ3kSTlVxlQFcVPVnyxoRr
3LMB5QOhD0bwsOe2fcIERnFZIGKhiV4SP6YxsuW0TMz0zoTnZeYlr5cQQI47Xsnl
yUtbi4mvyh/JgZiq5uM/LRPoFiVU3peJ95ElA2Elu6w7kca+bBiihq9F5fLKBjVn
aIk0K3jriTP45/SX+3D/+htoqZEsBLDZ9sie3srZsyf674QAaeAPovAl65xKaHCJ
UIY75yacAvFm1k9COmf8OcUtC4tPiuZXURd4dSpGQfIMuprC+uGqkxgIyo8V1r9N
YTOXiUaBqkPKM0+zirRjJcGmV89ycl5u+sGx5ak1PS34Ez2LN7w4VNkua5y2KDL/
wkDPby+tbF9uxwocnIafOj6SVWpx/V7JhSLvPXfNUrJ4x2m7TsbGLpHwGI3CY8V/
0qf4tARdNeb86NVskY0DZxeZY8+lyEUMtbz/vYZVkWTI1RHszjWxqIY6sGWVVLfy
vQMmmsxrz8Oh9xfL8OqbtNUGMfpvbCaku9FA3gWMKZEEuxP9qbTl99izEQpq+C8T
yjSwIOV4CCnmsA+ce5tleenfY23jeTljbh/CzmJ08i4N75l53v3rex0MV0iG2Lu4
MUi6R4BF+HrCOqVGcl5QwV0DnlNFws/00o+I4lXu9hV3B/5XuiYLXrnsiAr0whn2
tN3l7742FeV/4sKGaOKyJvAylvc//b8DBF81YBIJOtvVq+TfA7hVU/erYn4X79nJ
SjpNxvTN0vu4vhqzwQp+ZgFWtfiQ37frcRX0kHdToVATzVILuPtoXlqE3nIOI2pN
lm2cbjh6FJyZqSWMQHHhh+mzOzzdG4ovcNYlJ2hG87REqIHELwV6Q9O3rHFtKmgH
iqx0efTfAoIlbboIfzZzYW/OxNhH7udkQgo5Q0oW+dL95kBI4pMr7RctNTa3BxLo
jwinLrLQEbsKUv8PIYCcb5GgbKPeHaOVeGwDbVHoMhSAoSCDexU1QauDHAftAz0m
oHSyslRvl5TiXfxyEsKDs9xYbvFkPhDioeSbO7igw3IHwIk0lP+YdgP2jixihsB/
LikohcZKqt8FAMLJPqAI+bqPCxXJy7J4seFOwZwwZmUMh5ruZdIynuV69kJt4/UU
bt2Yri2vtwkbcGnAxS87+zk1k/2be8UZcr9hA8bp4FCeL3hj/0EBrdMX8Xwc8Z2n
hxLiNJEYmvl5tkNPe9G/nAzmT6GFwKkUrHnnZPLOSK0BUDUvyatmHB5ho8s/cI/4
MWllfoBfX09JffpcipQ2YwDW7zoqaDscrE0za2ZYf6GXNPDX8Xf7PigZOBEYl/iD
nh3JfXXzBwS5hpQ4X62kCvWPC1wK83zs69C3mqq0TnjscQ1TzkQSN97l8K/3f4vx
rutVUI/p2WbD28/bVulmJRW97yOz7oQBJBi2PXIDbpVUZEaSdRCrFSVfY1CPMZQl
lppKpJJl0yULCxPgWGFHPnfQuNFgD15lYzyI3+amE+BtyULQ1OjwrXFIhMVSZ8hP
a9CbYvaDqiVUFYxfj+2wIrIuvv8xgt+P895873SXT7NvniptaWJL/3Yc85WpqRIO
kZ/HkkWJ8HyJy6S7q+1JOZIJYjiEa9Gufye2Di+6ag8s+RN+Y9F8BotnOQvjpe8o
PFQStHR8a/YLOidMT7WzvStzWivxhpuKY+yVtNr0dmhsaSFfGY5QdoFbB+t2r/7W
uDYq83fSCh7VI+9hI1qSb7MKxBVqSJWVL55ICrxlyvLwyXNoo+qt6gm2wiObWZsX
owgezLi0L+3qtmNFKCdxm624HAI2sR+qNDNFR4bHk646gk8uPJS/IH0djMZR9w3f
xqZeV3iltYlQlnlUqA0xGeciHM1uiYVYEKiuEtGG6F/nWIF3UZlnJ3DxuuXFea1i
LudSI/OaLDm6CGiAL7c4PC9WOWvmgwd4bFl06GzzhkBQHxxNtaTFVn4GeUWUKPTB
ZEkWyYFKDSZvZAoAQt50YOpsLbFuaFQcPW6bADABrMBBWF0pWhPihmomBQb04CpR
z4ti6yxayQJOU0hcbFLX9jGGnKd0nAsaJSmmJPsd8iOeu+Pf/71/GmCtOvIc0VnX
ANUT2/tWIZtuzXtWjuBTkxeZMzjAMP9SzaD+ons2HooqROTJMX882L1rMfUlcmp+
xrhK1uG3VRI3egbliYXn18pUxJykuTnYVk8mw25HIOQrROqzZGiXyTOP84xXVbHq
bk2hJi0AetnopMcakkRd1N+NRVm3r8pnRZuGX7VreL6ixo8WzEtPaoAzHtLtmPe+
AjnQlkhtb+Q/pqrgJFQCBmDaIH0mJoORRNz6y3AIAa1NnNVrEyi1b6Uffw19GsGu
s+7wqyNcan1tdwVtbRKZlehqfOZQ7xK+ZvdTokrJeocY6xbBbOrM9ufv7yJmkaZI
WZe1ltIAoMbhYiC5P9rnQnJureswcmibS4Uss/Lwy5c0QqSbVvKogCRSnaZ4IKF5
bF6NL7ZBkbm7ryKh+LPu9glecSpyUzj9md79wjwVHvg2957/GPr/9WT6/WJR6CBh
60XUlQIfvK9gu7Vi3YXTCrn0CqPuhiCOnmblUUzowOyzkY4V+TSAiI3CXRW+d+yv
RIhR6toM9U6EC2usfF4T9S6hC7pDiWa15bf9E1d1/SZuBITCTJ9PssTPIdAtZj1C
m3wEucfjX5tYyTniMks3Bne5McjuJvoyRqLs/M7C1dfa2DVUId20lL2NLSBMbACa
rFG7NBNIQJ76shP6Yx4e2j3NBFvqBRol5cU5WDiX/u21jRVTWUo1Y+sBIqYBwxLh
+MNOSqZuw5YUhepi8mCQODrUegAu9SjuJuuy4mfvZBpLuusP9hwHj7mm+yWGkyR1
Y5jA8IpoPw8kdgU9SP4t5gMuxL3xNbABXeER4yJ2aNLPz9lpVw6wGVdiWvVJJ6St
jWtMZAs/5alHeOuUhtClILLJFj36aIimmkYn0X4GBnuLxXLiY+cVZ0LOGu4xVLMj
cq5FMmGKTk6GM4z8QBVHohDof2Y+iPgBDsOHakCRhef34/CDOEPQUp5eJ/lC0VQd
zEnwZ2cLQhXkmxKEbWoSfPlSIPBI/vEl1qM2a+8zApGRpQkrkaqyfRE1/GsnxXMr
TLj6pIcorNYE+K41Ndyiljat/4v/vo4X+JZzF/mBKLpsp9tjRIiAmlFs5wuo1vgJ
n3czfvGzMzStzH3b6Abm/NZl/s5EtF/2w7+LT2ImKEBjHj6R/O31cifj4unRHsTB
6XKMX+irm3ecK/CNNtjPZzsJVxCWPtVx4UPv+NU6yNunmC5/m9J8ReXPxJc5yaD9
F+5DdLAp+NYKuJ7APWX2Y4rvjV0eE2ZB1uZyfNIffZ0Pgs7UsA6qJxsbNjAH3hjX
1tD7d0SjHt/APbU2pqJ6lldYPj81dALgtsX/gjQ/Whot6M49zWpYrXKZQbrwKRXR
xBJjsGK0ho99k3Diu55PMPFs/UW1enqUS5qipsUqprtS+rliveQ1UHJJYCW48Tyv
m1w0Yg9kYK+KQehRu4+tR248ZjNxiPWZEWtb8zSY466yRPJ6FrE8DGvmJl6r/RIj
zH7Qrsg8cPiXhNoJ708lgHDBskBdJDkBvJ1VD4cPDtgYQPjVBy+Y9qJgtgKIfaYH
Dv7MGxXBo6WPPcFqbkcv2g94cljKEe18L+eWK2gLg26nHgW/mpiBNdmcWEuj3IPD
T/hQF361wCSav+Zd54pg+1SAUTgex0iLg7rHzkukNh3zA+VctlUJQJuT/q4I1SgK
jzljGrJVEB85l5K6UsVYJ0fqfPl78j79HG9HBKRDTpLSPBHu5VcJHO46zyS7uHDq
9N1IzznQoddXBYvitI9jXDMhULFSfjhGw4m3VOEx8/a6PJmrqzYrgxzjuWcte11A
67UpWjhtQ34fCikcukxagm4l7tBEPSn87g9IvI5nZhTdZ7fHu4xucgcjaojeWtFq
HcMiGpgxjcoYQUmxJBRC+xqW3YQL7z0U+5x+25t7jSdGjvyTzsEKoC7M3nPZDuOT
T9vETbedYkHY2pUncgS8wU1AEW+deexY4MsbZkSQasmtPqvhqwj+tTlIn1ayBG7L
oT49E7fKEakFCPQWej2oczhGv5jmtycOpA6PtkZKwWZq5tTjL9BvogTDdbjnFcUD
0kJ/BxPCWwroh78pZstFVo1EysuQ9IlfJXBeNw7GizIdRyP+edYXmY55KLaHq4+o
Wfy0h7nagHPM1Dvb82oQkFqKCnXANLzkeCA7gBX6P0BOi3361FEpy60Od+Th5xLR
ORl3x7YtojlDNEAC9z3pst9h2aCFKzeZwhVqmH7zMOyjbiANw324RA/IJBDi8OZv
u+zyrUWjWdoAmQWNrSSbiCl7R3+K6awHOxpLSXPAwJQU6qjMy27tq8Kq6+JpiBZ5
CbR/byr+0ZPM797mgnct7ivh5hMYwlS4KOqXDOZcL1b1QaPOBNZ+glpgZKrIP4lx
JmnNxjmQ92l1riylA46rz3AioxG8yB6JRubyH5Jx+CVh4Vdj5hFdkWLgg6uHziNM
FybViYycHM8d6tvX96KhKTFDrssmSgAY0dt0SKfZQwK88B3jpnxBvP2ZcleVbL3U
5lU6rv7jfejsYo5anj2/jyKxtlqBnrWDmVIUFMXnXXe7TGnniIW4NrKGIQ7EXH99
CRaFanVC3Ld9SI+HUihXK5+eprSJRiee90YDm0T0P0sI/qvQAHP049wsKbr5JMco
zOqkNiMoTJ7kV/uwOJlZujvElC+1T2FfVPLHrBdswAJ8L7EZ3CWglrQfy+ofsn5x
0522GeKZDORAWvN5K/QRF9Mc67qdPOVrkVwDs5WN8A61EjQv/aI04+q055EESiYf
MHAqjujOWmswZNhUhRfdBvzwhkRxrE23ea3/syo+cAQSeOfyDRk0eTr+IUs7EI4N
KiRyEsXNMRT9J9Wf+yK1rxEbGZNCvGM3KStrbqQIjqaCXwvv9X4SASbF580fl08w
P1U6+PMp3AQr5sbWiB3939A+QaFrTmX2KePhTqcIV1dlXp+N0CVnH0MlqW3x+hcL
vNN7W2f9IlCiPLUpCivtfNGygWVJ53p99IW5DiGpOk6exncS+IdlakGiHoBpQaz1
ZP2ul/lpHq4Ime9RBiqRl93XmYo917xly+LWXS4xwqljR89qFQ20eL9spzkrOEu0
QXc41yBf4AHecxUJyfUd3DNeZwjtfqzxMIvAZcITm0TEGMis2ollgi6P/34AJSU7
BzlKMCnYFchGU48+reQRphya0hiqU8O7qChPJp+lE8q8aihsw7rRVUBOioifE4+F
9rQMVU2OyNfZLWvO9EWsf7gCvBTIUI5NbaNRHcBFRreWkL9+9G+TzKM0JlUy9TZM
AICnvdpV+bEQqDVv775be0rOWJlHpISl3tSZ/seOPqZxzkB5Q1+WJbuTepKTlhTH
j7c+TckA87EXccqB9S43qrOWT8OYRVgPx+NL2QbiNfGAObttsnZp9KreSuVDhpDU
UXJI+O7PN8uaUiJ451nEjWJH4ZmYjnZkNN1uRaKMFYBN2KSigTPEkk8cIZU5hI7z
jC8Bb9mtjubZrjpOJJA276yQxB6P/KSDg6bwHGbWMcWIPetlqAW8hUZOcgnJe/0d
ZSiYREWa5BCCGq/I0a0U/ODhE23z/mnb0RdfGa8cW/bhPKG6zjRgrnyDrHP2lQ9v
s+zZpAfqWMmlr2VCXqQBIXsL78NH0vJBhBM7EWAS7tlOmLxJH8Ji4PtKP5+MX+Ov
+u4oNaqiS1hs5asrzlWKObUEwQGoLvTEb1+3RY2ZvVVXDiO0L9dK5GbfXcb1QDkQ
lw8wCoZM0urQVZzfF8iJXSI1y6XN9+OhhuP454p60B5KPt2yQB3gLVZrQcPui4dR
0nVqLjISirSsjZFnrY78a0qKuXuPlLVuwljKCcdTe4Gv2FJjsS4/dj7m4KiGX7yg
DRbrEmHY6UY2icym7FzUTWzxH2pnlLyxV+vvhfuaiEEF4M89Nc6qpnuSiFDFtU48
tpYRGsPqN95ARWuvJhkFQY7ifuzfsTXw8406zQU1JSGKXHgI4NJ6CnqoFw783WC3
v23DD2yO9igJFaqHWAMWNHrJMgm6R+zcH8/jPmtpYxtmd/IUBSpdgQ47pQhXqm3P
UUNqABxDcxwIC8aeqOKEWrWsKW5SjEshaS+RoEp73OqD9Our76TqQ+zRRJeXBkOX
ML0xTRgOffqClasEdsxzuQscNggCCyIfnB7wnjG5ZIguQS0N0SEpHKC3xIzBkpem
N0kabU0dAKgfLkFT2MB89lD6zZwggIx4Vi8OR2uCgtGi92gUcmtGDALNbuhaHvFn
bl9pOiUH9T8/EukRqogvgVrWTZrIo9319EDuDj5A2DFRYcLe74HwhdCBwFxmOC1v
ZSZA82DDSz/QNXrSdrz2E6+NWbK0IMWE7+OstFDTnm/ZJOVsI1kwJXCFZyj7ATBC
VLO3RgCbl/kmQfMfDjROXR0Rw01dMTE3yQ9AbesNc98M1UXGUm0ywUE7EM8q3Mxx
xIKBpS02kWzO4bil/u1uEL+F5zOPovROADlhP4b1lv5WKUZnw/Zvavpbcwx2A8o/
4qE4Nbh1CfZg7BG04AzqHzd8fOX83xufMgmWYda+a/KMGT9kyEm0hQaOC+EUN79u
Lg43KV3zrhtGrg6p6PSFARvXKyF/LenT/eFI7Y3g5UniqpZbK5sF2JaKgdZTQa0D
toMNLS0coW3R/YMUpIfrHevENzAMTeDVvAGyVQziR+sCLhESqzU0d2uu5R8vwzkO
hdfYT4/StGGjBE2UzICNrMaIoi97RjHdoZJgngWJhiktocl7lnGjCk69xdkg1+Ha
1Xgff9upOAGqiY88D11uO6Kj9KXnpQYCODU8mxFR0czPG6aLjpwfmxndOWKmwDxx
nXtpLLaFGiK9bVMkTFL/IQDNxcGlKmfLFgK16zjoZ+RtIrjzxm5O5RG4d7+eOxTv
jvG1VCWRlJ7Y3p3KpQG6DSZMM+YZtM5sR75E+c3E6pUHBKn2tlVhdjO1euRZTR/H
rC8wTWvGZO74sv9h67vgtgDZtxB2wZM6MS4+0fpvBUyWoBxUGUT7NvFiPUvxmMIb
JqRoEo15sgx9zhGBGJ/4GeAQzSkztBqjCQrqxp2MDq3Ixi3fuDpD43cbi7O30wfg
C+xyUb0QqTxINaPq32ZUtb0u/xDI0xyAlp81/XMimwMRb2a6CL4HpoWW1BPN4806
kCE+/kn1L+HsvFp87TOrNux88UkEohRNN9nfThUWwHjLr4WlspxbXkc1VYcTJRCP
6Q2pEP+HDd3+wtZkVYzLnXL2W0EouMfvWBD+XpaKn1NcbZWh28MhA6FRexMDbIqw
uQYMN2AM2SMigJ7ENtRrm63bMVGc5RcLEBM1YQtimXO614bPYsOm/JBBekzw4ukB
X5a7TiK8knQu01bFrI99MRPMXKjsZ0m4prQyNVtxv3mxzJbgVLgaV+0SNYa5yXoi
aAh2dNnygYS8Hu/hxeZuzRpyZeh9/UY6Rc+bUM5vOhvUkKJRaZf4UKKF0zq3EMSR
saURGhkzV3GZTI/S9YWYmZ2TONhvOXGS0MPuuiLpHqRBkG81AAwLD5GAz0bnBs+U
JHXKlvTIDjSX11CobAPGBRFedGE20E88oG+gpzHCfclekLyhCFKxJ0ngRqzHGrek
SXOXrkqxQfD7W9BtBQrq3nIEvm1WS301kdqyRzwQ1TRYTf9/qlUTdrjd+KpJU4Lz
R9/RQwj6SSG+HrlNTTiqZIzST8M1jxT/t37QVMGkTZK2aukGhDTjGfw9ifoWvWat
xAfF+uIJLz4MSCdS83kuFkUbfi10KWXMAq+YWrFrKCzawBDUxBdC9E+E4HYtN2Jw
z/kp9fFB1RvhkcsEBKg6ZNsMsZGcwZfszXFSeMP6vTjzpb32OlG/8Qztus7vCtKF
srNYTADXuYJp9JWLLRo3B0e48vCg+aOaNehgEQh+QxkH4KHCx6VzzOHxR59DA5Wi
ZMSdC90hPKDQsas9RADnfNDTZElavy/uAH6q/GRdCo14CpFK8/YF3isxOEnJeMh9
nYh1pxS0a4kRtSbUfqu22m5JlVcVJzEqMJyhdsJkYbfhKwydlUkrZWMlJmG+hLgP
tlBZ3nwNL4yqFglJzNU3QypMxdFQwjndOJFdmCIVpvuq54AqUx2qfU4+0H2RCFgk
G2GUczVZlzaJZkKo0ni36pk9+jE5ZtxlB1S1L5RB5dyU+sEO6VtA9W8CCRDLLMzj
hGaiSrJND2Iy6goNovruV7AzG4sassRgs/h7xPwEPYOQC1bcbc1yd2dciu1NaIgY
FIuwpGSqy4HemKF4skzXUXvtAsCUxxVBtA0AFqAu9D6iOxDsEq3q2gpUnbN2Bf09
MFbqfqfy99NZplNH6OTMrBOiOzBzkNzFL2CcwgfIS3tKcNFchRV637diRGIMPfVx
sWroswC1Na7ZzDq7DU3t02zJQcmfZ4vNZgeZ8rUjeVLDFB/B2DRGSXkYZIiFgphL
mOw3Rs24oeXRpQuhU6tN+qClGF/PHz3vHHXDhfrjKETJAz/6ve+MXHi2U+fopmN6
5+IkjcqKvJ0+syzVonWRz+thyyroxQBqlXKzWgPjN6c2vCHEej9iZKvjJhkxbi5O
Fw/xv1FuMGffxRa31iiLBarhtOhljHqBzBnfK2dPbVMfeStiB4yjUpAqX+uRqJq2
M12TkTc8B5jvkuys7V79okgnviedlZIvDGC5PcRYq7pmuk1FytccCsq9r8fajtda
8iscA0rMzPySBdBy7TxqGSOo7ZKnnkCthiFcLdBOk9+2XykSCcxdCo3DZWVcq9zH
OzUgkCqUjQRvivMd8ZiOMh9T1kMxFhqwjK4L5kc5SB+EdFEUoUUb/g33rRmWkCsn
JiKi36wda0kReFxcHTKNizgdFoD2NL45vN2qL3VOKLZGwxkWb1Z07q2M+xYat/cQ
1sbubga+cKxhAxV0pB/WC9pXYBx/MVSEtmvq50MGPfP1I73oahap8sXS5zraOoHc
5FjN3e4HYxfyR/gv8PB0mpcG2ZDpb8qORRMWeaZDXKHssQfcgLiEeYuKbEgoO9ni
TcZTtihIUbW5my7Rev87N/4KOshAdFD/+8ELxXLhPS9QbkkInwak+Gd7b2LPmShq
i7KZlnjUz8XcuG5Imz5qMVZ8yA2JG1Oa8S60dh6KMzuXyRQUPm+oT1Py/j9r3opf
nz8wvtdtzTt1bWRM6z7qANTw452gDNL5XTXasKUpOWVf4Y/8R/vw9nzuxp1cHEPs
m0qzMRGvxQkTTRmrDLeddxgBqtneuON6E/rMSM1ofDw3/jqTILYmbFMHHPI5my6d
ZWeageamEtoGGBq/CdZnyzF49AT1tK/RN0RhrFjnymW1jQs+v4eXykH5sypc5oyw
2dumw4Bu5fRKWyqSnXGS5VkXZlVzVFAGC81g1tijkSJilPDfga6ho/shYXG7+bG9
lZFlSz0uprgoUZOeaftS1YyuA6GuPDhCDewojY+9fcNREIsgZ68eDHelujpHARsd
yThM+HjZdKcrfB/PS7ROzIJOMPzkKoZZFzfZW0H9An2cHNZ6U+Z7JiBGQDIm+M50
R9JhSNyYP7+RXJMaQYco3chuYhyQ5CrtqXMZ9l484KOEpFge+2XB08lZrIDUfYFm
YodCwsuAl9xw5bhx7KkEDz5WWlYBIue8VEDY+JTVGCmo1bRaucJHIDhwxtM/l7h7
w3YG5JJzsNItCS0pPQnx17hZrDRY+joAvP9LN2YJ5uVxwLTE1+nwqVRf7J9lQEN5
ncFDE7n2wCZk+oKOYiAaN6De07N9pYuH5Ic4ivVnpso/QlJZSFyX8Oid8g1EHtU6
n7z8GxBpoFpS3fcUsEv3gv+6j46VweHmm+9ZBPQaJ9m3Id8lQ7XgJhRe0I01Mwvr
NTVdV8wEA6i/k/3Ck8Fg1jPU+ZdxbWifT5X7fgTfhGW6eGy8XIpvVWWQe094zCDJ
FJ/Aml+sZe+7V5ibQbnQsdZEoXYCq0TTMD1at9CUgoxMj2uzUTnVuFKwuumEymIO
Yep1jWXNQDGk9VlTfJP3FYNgIvv1C2wkDphCp5jmwD48BB+jLyKbzx8YEUjVqd0E
wpSDcoSO61+WxsnLFfP19x7G1NAV80NwvM8lFhU0yDxUGOWk4aKj5Ok1L/1nawoc
cjdYalyVdmczdhUb9oR5/pytUuTE1HWP3CBJHxD+rK9OE0rxySAscdC1XFj2gFQK
xKy5A8euIsfo+pffvZ9fVyWoUCpXAGkjGm59r4FHulWpWcWeEe+QXu3JtFFzQaOI
dlmeN0JtbPsYS6N6jbYTCTifpDIr7uZ1pH7LmCbS+6AG7WUPW8hLdfjpy3SzwY+I
D5MuFENeQydWqRUkH5fxGZ8Vw4LZjCglTatH1gicH8UL7SJQkw2+ZzrXfouUoKKc
8WJLzwAtzCznav1D7ufkosf45ulC3G/P5Qfu4a4X1j2ZdYzVSQA7+mnStEwp5+uP
Eu9wo40h5rI+19Wg/+1e5VrZR18bRiGuZc5Cukw5pjp0fK346MRAgJsQmS9uS13G
Xj0XcetT/v9hHykCDdiVUvD+TLOuMvLnn9h47DnETjPTBQi3iV4KUndopKn99mkZ
bOcAgGsqTzgWxjUs7dtuGxr2MGvYNr5E2S1JGY0D7SK0yAdMAd6BMtnXGcOEIjO8
z1Y1Fqq3IYd3+fonv6vJDqOKbcxhBxf7EB3E7ei4ispi/VSGEllw26a+RmtIi+iL
B/JaKspwCy2IkAv7yuGjBZp9HHsjCoEH/NC32qlS4XSbCXkusS68aKu8MxAr3+kL
aJ2WHT4XHWCLexuZsghNRVrx8QSReaLfx/yVBKkFwmO9I417He/gNQ16Wg3msPYK
C1VY4mRhmgzyY0CfR7fcNcL91BWj+8ZMl66ue6s4pum5sandHg6NWrTjzNLpkytz
aC5Tp7LQlpuW4vGBUTF7xSc9jBBy7aBkowFRPQLSduoq8ouSWyjA4RR5gpVGynx7
JIrkbprlVMkrYXJgU9juT/CsiLB69fR5805OYBokvaASZIJjNJt0bChVtEDe6sey
HkmGwsoXX8KGZokF8MWHn0jrtC0MDEvF0uEMD6MD0l2tOZ6hWnZzCjtzBQhaKj3z
H8TLexNofWQDJfovv++VvrbpnCoWpYTATKwjcHuaKpLSBVYZNsjvU0QrBycq6tuD
82A35bD0ks/3+fWL1KdEtYauZWZIR25wKZvWZjliAvIwD2iottwBzjW/qDstOFMT
q0hYkhtV8yo9sO3Nh8x0RmdkiAybzQwBoiztRySPeESTF3F/tPzF2K5YxMgbRmtt
2yrk47sM/aFn7VfP53x45osQRWrLwB6/7ku4PO6r47GSE8xvZwl9WpGNTDcoAAob
jJqLVw7We9AXLySFxOW28jRePM+4SXPYlXj8oUcBGO4Eo0UT50mgod1ecFvVMjZX
gzBd+iDAXWgXZagCm1I5ezwD2lRPPdPVHAfxdfnZ3zIL55kK0ygJqeQgiMcodnl5
KP7xPQiXDyPXGIEO3A5zZq4BzCWpc8hAbUnoXG4fdEAqUXe5IHjNbWKaU4jEg2MM
eTr62fIIbPn9/dQ91Q400ZUbTjT+eroWuAj1hVwWh1REJCljm8dFdhHF8OmUoaRG
F16vy46tRJETkGs5mrTN+NLL0P5VlnhtbIswkyFMwJDfDI0SQazRmkxsjbH4v0dy
lkI9CWpsMfUQ+iPF32I4sfJk6KZXZRHOrmqMhauPZsnksc75jX+68AAtMRDnuHY7
GFMwrg/eirDp8uhNgNlT2intkwdRJLzAnyMimzDRzi1GRg5P/dKrAIpl6vf8nyRz
1QhNmsKSZbYeoN89G0LY0ZpR+I68tKbx8rdQ1ZELpj2rozbPV9XcZ7sM1R6Ij+sP
cPTr2hDMcJmxH8Oc0V1992BVIOn0y3obmIGkLrGi7vKNTHTGYbsl7zLR3cxuCbaW
HZcFiFa/WE6TNe/wLHXhxwjCm1I5vsJA6EVMg/VA+LWSiDODFjzMGAP991Xa+7BP
Rv3TyZaBZulOaWXq7T3dnSTlBnAOcbaEJgc1pLAVl1wSbuwgN/ZFnVAEfNbrxVhw
ol7ZF4uOK0C0S72xbhxXAjWQDQojE/DCLwACpvU3ShW2wd7oIjf/H0zf1xieT4VR
ZIcjRpxpLxB9uk1nBp8i/daDIqlQHBb3rMfpaSMl2fiJxxc8o9Z1PVeGncnkpe2T
8hMETMfXZ3V3FgPdYxKmVJQsja0P+MVbVfBy/VDRDROBb4cltE3GJ4SNMWCRFU4S
ZFYhr0BLNrVMIPLCDGdNLy0yb/FIGRTlbX6wfxSx4NI8+qonwglxrMHrndzGU0Dx
xY/8o9Z63qr2tRrXIyfv+Pky8ZRTCRFR+Omh+OSoe4rgmdZvz2WKM5LNiFa9RPI7
X4TGo7I5uXhzA9bN4ZRrdnKsevcU9+2GCCHb55jw40jA+ASblHxp/ABGp30q2Wfm
/AxAvVHx7aWXHi5zdVtkg8qWnTDbBPvlD/b0JDN+NQxSQFJqvPZuHGk9mY9LQknv
ru114Hardplr82k16EEbHwcMZaKiN8/gI2TFtTgYFM3weJ32tjGe8aqw43RRQAt7
1638drTDO+LnF7cHaZ6g/btJbCHtpOc2I9zRheCH/T0AwfMJiXBNrZfxBfKxPeBZ
L8J7u4mY5t+wcLA4yHO1SwT3XHmSR/QoY+WfLLfe+Naak3bypSxzLFSPH6O/LVwY
Khr167yHLinZYpal4357A1e9FSYZN1fm6BFVgLV4jvy8qY32v74A6bV1n7GUCbzG
q5UxkCLeaXb4GobxDhz2HsrSaDcfxClyIHFq83eiaP11ddJvj0Zo4poPRIsZJoWu
2oKUe5yFHC41UP3A5ufyoZ1NFHsFyLCWT6DVnd/S0aqWErQY4jp6p2pqteA0UHRx
JjiFaoLtKm3x/7hAo2MAhNcwe/djzPNp7VJI8s4il6mby7AmEAslv0PnNIbEgPBi
VykYwnpv+b7OMAHs15/tPP+eLVrxxjpC4+VsXrZ3N9B+GGffrsvAGPZRyQbfOIvg
2zF1MKSOUe6sUs/z9c4elebbneCIEDSQNigt8fm+rNAxkpMW5d7kmXQsKQthNHDs
h2QTbt9z5gVLeJKdy3pa7zs2pswiAj+YV566qUzBnMIdCeAiEgoa2TTf4BzF53Ue
foyWEQYByGQk7v4ALDC3Ifj8gI0JLc7df+LsBtQN/yjZ5DsU0ep1I7dCb3S80k9P
SNsZmc9StsacXxqVEL+GmqLbSiEqERgTMn+Jwn+S1lx5qd2dEdtuRG9CxQLYvts4
jdYpOGNbD47inY1iyHuTsZXy4SYgOR1UX/0LYq049qICyuJpRWW5aE61QkCzW8ZM
wbKy5F2+rGHHW9HCPgPmeIdlXUGpQrbDFubJDR/Xlb0IpMXoE6rAUOAovBc2KJBF
tAZd5pgENr+llEpvDWIbkOGNGsAMlZYJFBA9MJmuBoJPoODEh4DzVDPKwS+Gxw94
RFNL1iTWeOk7OcJm4vJfw/owSYULg1mUNDQ2W/H6F0te2y8+f+904e7rpRPZZz6F
OYN0TvUxrvcJd2TN1VUIqOdwjr+9XYm0w45GFNJNdmuY9NsOz8M6Z75TRa0BfoI2
wMQyNrfxC0awU2ob8Lp0DLw6BWVbUpIzgO7dodteFljO7NfuhKYDiI+S+D63N+3E
s5mFsoIUxRoBV0DqZKSMdbQ6lcJg3BbKq63v0sbu3e4u0Fc7rcQkEe1K8p1pGCx/
ZrdYwcutvlkCHjR28Xkm+vgiffIuhGQ+c79oyPQpW4QG9jn4XlWve6ejaZRDO6B7
s/zYXWmolMIKrD3AMftdQ0BXAabNRySeZJAPHjrXZW6P5XL6LBo0p5WOfnQRvAQO
4ATEIA4EyXBdBMEVsVlcnGLbgdJMQP4qARy5KNMcd3iKlE+2LxgswUyU1qGMngOH
wgapm1XYFsg8DureGDp5CYq00kIop0dq1z2wmqNNItLWi92SzRpE6TqYSKGPkfvp
I+IadvSbtMNLg748cbmHx/5UzXvzTjDj5FQyUXgW2h1MQBlMs0YExYbRpugv3rHm
DKfL8UCcodQLD4nsJUhBYym7q5//r68Lv+fsjaGGPgegsr6S1DoDiVtg36ik34Ep
o+SiD7lm9mlgaEAA0tFsJp35oXwS7wT/K5i6a8/D+U33JEfChQar0TiGKXEI5rTm
QMSEH7QjODzmxFF8aap2cMyJWzxNTkebyIpAWYyK+Nzmst8kEw0Om5NiLUW5V3Tu
neg+/XR3JK3CwQeDOhozfkgtwQTUYMJ8vVbHOilFEfM6v+k0fnhJj0/pRMNXixdK
flAKWZWktd2oGtUDtkNBjgZy7kN7Uq2cWNPSqXWD5ZeXDev7J32DELgp4d83j1AN
gg2znKGqNgIPqw9kSBYbfIn1BheOWW3sO67jsyGobbqhB/jsuUVRq4tYRa1TazVx
MSz/azr6upGsOjPIcl8ia+pa2jx8kavkQtzp0tkeaQqj7OqJEerU7dQx8C5oERZH
Oj6VFZ5P/8wr5Q3AXScasOe8YKpJM6p/lBeQMRSv93d+dFxW0JTPR0BGLwK9Zbx7
aADkWUZtELjyqrUARMGYrxKKKFy61bD44DftE1XF73Qig1WQQUQYLtdOYYC8Ver+
5cUfK9v0ITzrnthOCjSAJNPK3+ZTzLPS3nSEwhYPFkZ4hTwtFIzP1MeLnDmaDkZQ
cQcFY3eTBVIE4t4zfNznqqZUiWZyqwO2aY8lFncgxUpEgZHLI3Y5QxPD2WNC67YD
nOejCZGPS8omH6PZLgYDK1DhGUSs87OGcii6i/BvF5nltMvk+Kmd8klkEl12Yi+Q
8M83Yp4aG70JOuiIeq9uhmWA1LH5WBj1P7aI0KLnoyGPc9Mukg/BhLrVOBimGbeg
BLhg0aIsJ5qJJiz4u3n6zl9IrJOK4/R6AiyU4QJb0ino1fR7idJfN+TsjtslUN2z
1nhaGljDS+H7lvdfNVKHg46molKJSDJJx6UVymVpTpmiW2IfXrOLPzD1SIXLIkxq
bf10cj7etAYgDr76WqIf9dC7AXmu6zGs0ImiAPNizjtz5iVWnqQPdqaxAIxhFWkE
lxqIO+rcRtOWKHKPX0VrY0gOREHgGHXBrPx0wog3HT4ktjHCMzENQCvpaExKsPjz
dbR7favpD41Nl/m766uFj2pIlY1Ux9MVvUXHYikUKK070sC5dvsrltlfXsVsI0nD
tvaFx/+AIrB7zh4M1pKr31cMrcVnuECXtRLtnKKS00jXMtnQ6pu58BXP/4mkTxqM
SGumnCBAe0n7Z85ygMCAKZQ78d9nHGi94/zULM9c4wX+1BpCXiLQRVyEHxWM0KYV
BBoDaXEmyn2pqbVTaZCD5zhnbUaIzjI6B1OGe0gqW1ZRMUUpnFWRdmAQDYn1mXJ8
cxHUjbOqs9HaZmTIjvR6bQshnEHhg/Wi/4SIs9n6ykcaLFmli0ybHf404Gps/tlv
6f1PaVlguc8Yt7bLnzkt6ZYUy4AfY2P/O6vRK7E6BQZpM+L0dcACO1ww4Klstrys
9+cXo1PwGfecShweYasJXqdDTZl2L4IGzs/fzyX0KrqL/95+RZJnU8M/xzNblBHX
yzmaqSq+wPbVP8RrD+TRZ9bxgduB7aYx0SxqxQXCmj6rDR4tpfOAd4LAqXiabdlv
PC2tVE84wwC/BkBEIu88dOySQX8yrf6gIklyiSPt48PZBJuTTDJmSNwThI1C1Ejo
pjWK4QU4o2OKR1VCKxE7h/Q+ty23/GG0NkCqZvcZEkTLm8L57P6PBC4ILTBoopnT
kjf9rMtD5vGoIUoJ1b2IHUAlh5pgisz1AX20MttDD84905NhIRVpDrEbtLhr6VQp
sU+Mpv6uDFGHJp8u3dQY0zk05DdfeLDhQoTtW0OPY5xEN05MX363MNSSorKXEAVp
8Spfizs4YFQRPgX7sCF0BRKZpZlZ3wUEDPqQL8DFJ49MiKOxduKDcZ+ixbm8Iofe
y29Le0/SpqslEwjDD6etTcvNax0V9QP19mOQMBCHInpvl9DY4zwNguANlGcdJwGE
7Ye8CP0dWP405y7PjwzNaDLZYgpfj+LTaCvxcfS5OmjrUSbxV4BVocurt5xfYQ7g
FwME/Zg1G+c1widWVXpUm1YUm5UTN/BQ6rnOSGRp71k961pQDxzR5i51syegQmuK
hz8YBQFcxue5fnSTvIoYlMSJN1xwZ89se3Ad2mfc6M/18YVbeg2RFKkIPISSqqPY
7R8PMe5IhE7IjxN94hLFRtkfmf0HH91/2Baas9SoU3babvOlxcVvNT+MIqBeQI70
VAMDvSerVeQY4nzBOUbGbryeV/kGxuGFYDjpJJcfdUgahZqhpeyYFOvfctxW6Qmj
Ct4NLOoZM2+107EL79l0ZmzEnde3dLqrdmXIMzUqUVGTJ0ddK0gs0zgo94SXl8YA
Rtq0Oinw8B0dudnaDPVCBmzb2RMiK1N+nY2JpETzO8St+hBIiguu7uIYpXyNqUbt
WI8FAp49YfLNSkk8oV7vh7z/Eso0GCxR6Hn5hUXNz3oWP5aHzNAinINrWXV7a3pb
fObSZ/b78hSwR2urR/mihqMtOvf9DgeCrphfgD2G/IzGYyVWh+Mfucx1PJdqIwvn
EwkaygM9Vc3gLw2M3Yo11id1HpODYopMZnN1xEYNKokxAkTruNmRCnNm4aNytgJD
9nBh7FGR0lZ5K3gurM6u7CIr426+/a0Cia8ENGj7I8LQeV1YUW/c619fahPqulTZ
E2qC8U1QBS1kK2U9ve0TWkvyIashcu6a1c0VAhDPsLhkkNV5VaaslYV1oSLE/7A6
9xMH4qwSqqJekGVnOXw4gyGEFwlHyjszloQIxRmLwGZnxxolz7qFdJ09V4tIbaH+
N9vvhBZhLHDht1LkOG01mFzuTWhWXrN2PyMkMf8K/h/De+WptFqHmm4z8X3vMHGG
L6X975MvWXmn8Utg0icPCVcE6l8asdreYDsl1Yv0dtFLwDic1t1PAdJVY4uhORtv
2QtP3ZjDgGxvARcI6KK1IJMk1ysDFfPib4aNdO13OaTVxuVu6WFL7eH22jKnCXMO
qcq2R15/M69TogkVHxLi5wJ04yHxjve48w9nNJw2XqI8M3itecPPxHWbmpI8PTLH
qQvGOwubpr4k5onczYbwpxZWmueuCnM2rzaHHIhShZB97xO1IWJTc+kc39xGKDgQ
bgBy0Kr4H1blE2WXtOtlEqnSFIVKZNnAXK1QZTu+rR4gILNVcwJU5a1YJ+TiNnJS
2paDBK1SkayuX8mm4Ftr7ItE+ckd1FzduAnAk9tXp+S+OXlhNsmHkH7mzNDOV8n7
0/vuOPedrURvVRnbx/Y+bInbtDGRW7ApINaB8dARHEw8XF9EBnCQik6d63lb0hz7
IZkcGQNT9djH9CDvEceFSAdbWyWrvFAY1akMQDMt8PG+2Xy79ngVSLhMsMyue54t
7fPU9aEczt277TJlllBSHjfG+eBIQzThRQdPA9VZc6/BI1Gkdk6aE7PTr+dnOBHv
UCc4KdOYBrS/R3fK0P1HYD7IRu+k61s3V6x+s1Wm0faDNVWoHH3tGAndOoZ5RuD4
RaLgZJbdxyK7lmT5T65y5000S2Wl0UftBqSWU2/y+PQcHbD2X78EaLhV7U54JMY7
OoD7pUWLBKGs/u8LF27dCVt4IYUV6bMYe1dG5m+5SqU2RAI8tuVXyu0bkR7x2aSB
VUMAd4E5nKoK52tAml2ayA4mOjWdxKop+Z/8xlt8FbO0ZP2rN0NjSUaLEi6+8yfz
AkO6Ia94dYalcACD8Js8KTNg9kPmTCmOyT9TC8UnVGkB/YN7cjK+jLzTqKobZRCL
qBVSIC8/UH8XCa5zTY5/7WvnOo/a/CLlhgrxdW7z86jbO/xIgBuI7s/Hx2dx/13d
u4NUsE01/1sQnSw5R/1dmr/+WcDHCa32f5BvXCOD/XYgUJoOY1E2rLAbWCgiJ776
uFh6nVgROVVNqwz2YcqwlrZeYZyiRZk6M6hmQyTno6zyDB/XPgxqj3P00tyn/aEh
/l/Bt4d+Y8rGV64aL1ky1mCXf+f0+UZ9ScsFZqD31vWhMssifG8phbVlFH76kEIQ
GY9INL1P4V4WVOi5oJOrLJah9ACDtEC1ZFKOrwIK6TrI1aUwS9FqivZWT3uopIlM
s3eSglpBcYzYQHUjMxxPKl5oFfYi685KistDVTTZvmaznILrcqmA5GDh8CIirZ91
61BdGsnb3fL8zZuEexGRVyYo32TGeGR4HLSdjelcREGyV3wHSkMSMj/Fsx9X2kNo
W6N8pX9C0Erqri3H2YrWd0r/meTR4s1XPNhK6ep6Pu/qumUgJgr3E5JtjumWVZ2e
1VCvInNvzk6UaesyznuZIPyQV/UxzXKt3UIOTp0XX9xeSlmwhQy4vUkGl1xY7dd6
p9P996LyyDAWlKirIFQP4l26DRrAuhWV9On8L3mOluJnzvGusDHT+BSkqARPK5ou
ThUDQ39DyFsUJ7MAPtWgAFB/eJdqw2sGbPhpawAjnCNj55A7XEhq55KksbJOtg8f
U9+mqopMSgBwsjsWZ2Hcj1o+NG08REbnkjGdDH1N0mbuuG/aOEcCJEsZjnBb7KUp
zMDlpSevvSYf7F1gXl16a68ZHCem26x8zm913lzUeFR0vVnNBreLGNs4WXWlWUWf
YUleiH7Wwyn6AMH9kDnwUrkSkvoUzUhIMUHZ/0ZZRJWq6hdBsqwfqIbrRilgVxoV
tPcmw869ZQGVEtNRDCFqVbOQj9CVxnMc6+C9GO12PGRVrUvPE1aIdc6vzcxZ3fIJ
9YeNk/TkS3r8dxBMCv4IlWurCEgeHyp3xDii6QWyY5CKxnJJzv1BJLxNvZhd6dSB
h+3lZAtL+IJJ4fFHnp8cin84cx3i7CGDhSH0dI6Rq/CdMT8XOMPzISupoux8baLf
DyP3gTQUOo5o0m4MyGfHJ562/sHTB7aob0IXwcB0MwELguVZ5RuFD2WdYZItCB4y
m9cv6FgF4tUFtaponAO7ZPBoXXjqon+Eq07uGaYin3EQMVxTHxfwalOsCADwJxUF
BV57yfljuEHXkjtI2o1iKM5FYCv0jGLBUHhZqq5mgf5WG7l6MxnsbJkuj+QmLiKs
moqjsloF6R2Y0A2M6aByazWCNs6Pvb7NlNrIfpkhPlXORKXK+ZK9hrDT76x4yGnm
CL2SD/O2kU8cM3BE3zVFzIEDAavtCFQwRFozCzFtcL3cPdQAn+by7m7j6Txl626e
qF+JUmlKgq750ev4s15AHMOfOQRAlBgsF1HkuVKCHBLQ+H9loGgncGzM01ur9egb
FEeSXpQAztg0R2oxUL6adUNMrMW0cfxMQFnDpiN6kJ2dqTNrDSGja/j7816iZsA6
JzuoNrY71E0MryjwQ5iuUoOlSDPPLcgvdn0Kkmz4Gi6zlZdZ3t9Bl+ykcOcBDRmK
9r7sC62v3mMd/d2xVoXPLeI5ouRVuP1wHvoVqhFMtqwZYPERQi7IwJ75hW/Z+exz
QNEWzhmt4bBYrGcGrjcrHn2BEPkt20E46I7xMoEmlLnAffH8m3yijhdu36TrL00m
OLpHHQLogjBt2uFjdlc4P7wlyAMQ2/8bZDNlV2KlK2R1XR8vhR69/oa4i9TaCPHM
mx5r63sGEbHe/jMKpHTEHVUWKPq0Gqcu4Y7Oy90SME1fNaJHNHBJGhQsIztw5zJq
OKgFSgAqVYciw31RY5xRmp9wST2LLRx7UTZI/sXezTKXlk6TrG6Wlv+kK1KMPMvT
MG9mwoUwFss9q9hhQuC3jhnuA4YGsUyN5Y2Fo+x5hjdBl87ba41szhUg87QQ6I3J
qUEEkyhlymzlqJZrer2V5k/SSj/wVLJv9m93O0y9XWYtKOyG/uEbi6BZTj8nbMMM
FINiny5b1qGWBq2a89Spb6WZUZf3o7lUSsrjfEG04Pa4Jxs02++UyacTIL5voVNg
UAmqeDdMoZmPmclV+fJbZrNxeuYTgT4RZ++kiiP6La2TWYUnpvmZ8rtsAdtWvVsB
kJjW+xNf3AV5zNjx7T4Dab+8YheGyuCuPK/0jqa0zK/6FNtpLO83uDpDZnlLynvX
HSmg7nF5VKddnKnrABciykxpsoaiYtL9KEhV+OEjrvYmIh8PLFGJg1YPWZ37E8lV
BBs/L4zFVwwdbhNyoUQQmQ3dV0UhFKZCooY76cHbZWX/Mv/TINHeUeUZbbtSwaxZ
IZ1q9JK+3zEodwA0UvpXo6gHaTOFmaHtqCrc5W/j9pS4au4STSBOqF8T5Ym7ub0d
XDj1r7ePOwwmHl+Unteo6+yHa2wPigRZKFNaxQEsV5A8QIM+N2ViNlsXoNve4ZY/
tz7VWXMXrq9ZvQANND9JXNfLluu77BclcCdUaSUKDff5+gfezzGxLgK2JkHYE1XJ
VSPMJc6iWw3orLnUoNBYiO/DAlMFEOUtV+PuJWTgvSCODZOT37OOm1fyCVayJ4JB
pJbcunHGTnqLs8Y7d++pvc+soHY+5o80cW2GcJt4Ar1z+iZX94XXff3FQFImu89/
ThLJpMJyNNu6E4KKZ8tV8ohJY4Pq4E4/8ZUALYvPGY77/eFO+duqdZmPSjqPvMjG
SjJqKKh4p8505JJl5jOgSDhCVEuHzkpxQn28pfSpRThUf35y0Ib6/I3NOOOlB7z9
LlxH4iKxpWpVHeB9WPTdaPtgS4MPt0snEUBEiAp4HWNMCHid+mZAANgw6cItJFUb
3sMgHBytgr951I5k2cVkcea0V7Pe3RC3n5gr72VHe/Rb/3lgcvFeBIHWbaEY5Q/6
C9WO25TPiaflydmXOG4R06w7+Kxeog24Y4UqGsJ9JyyHzCB3zvjzO/b95Dn2F/st
BFREVPANwtrJEKcUTIXR7E+bnAF+rIc4afhDhP1LKB73QRFl6sfJbdCs0ORFPNTr
A6Iu5pK+LA0NxMDItVYVag50ldmrTBLCf4VSBjrSt+46SC+kneDg1JfwT5HcOhAP
3Ooqn2mYW8xhg9yZKfoZR+zjkO25qqNg55J+Cp/lTJk5NFdiczhQu723lAymuzvo
3Tr3wpzqTnaiSl/H15Y38pT5CV9J1MawNb85WZ/e8L8BwQxyX0328+gHberhyowc
gnZqZfuYROyiR9RWbCQo//ZPJtkcL/2QH8kYBacfdRBzeW8fNp05KOz2fMAv35Wb
njK2CEiNqEb4NVNyFcEa6YTdUnfc8iH6ZbjeIDIb0nI3+dvIonod6yk1u4sz26Hj
rTbSPWjOuxqvrdobabQnuULswW/7PiBt+HaL697ybGuv6pXRqUdMjqDndLLl/03B
nUwsB+6Z9aKVzgk85/sva5Lg8ybfr26RXWdbZJbsT0lJK/zpgqpnVtpSUSysVlHw
S4DNt25kkkZFBhu5ZXqn0thv06tgoPXzT+GIipOdbmO6TOK7d+CoOutPlio0gJN/
dFpxCriMTWk5yFEigxLkAOMgBYRrVaXMBSMIMLssJZIUrU1VVs5K/XSjkTrsyXND
9Cvi+ZnRKttPhpX10GF/sn3GQxHEvSDwb/h9Li6q7aJG13dm0RfyKlDfDQs/vqTn
4ZB02WMeBIuHdyOm/k2HFoXZaa59O1r/0r9V83gGtcziLZOnC6o6h5UgrNHnkCtA
gA9zKIDVCLcmpgYdTzHW9UGY5bhB5WseK9cdxkUQpE9Rxk9snItWIA1oBhqVp2HV
TLqDwVpeDkCoxeHX2FumskBiA2/3hSd65t4BY9hnK+G9Hu5/j4Ms8xL0d5qP/LoK
KPbnUGHDeI8P9YWtFeau/FMwB/17IflPMoWycV8ymEldlILQk1HWC6KMHc7IHuLL
0V1VDt7ZfLIZaYfgRsRh4mDtaQUdQTadJMQswd5FxIN9KGzoZjsQ4caWBWXS84+V
TrkBHlng13wSHFhKYI3kXOyfQiKW2r3Wgmty/al+nETxT9h9N0bZ9SAS2nZ3bC4G
4px9X6vER4PwzQ3t9upF52FO5YJVkFYlb7uWhb3Kss6dSC3AYKGjfOTdRSR18TJP
Bl+HI+OJORSdzHz8wnajQ713Yshl9eH75BtQqPZobh5/L9XP8/W0O/98ElSxVHdc
+m+a1MIwTV1T8c7hL/rO39jSBEkAooLpqTtJ4+Q2hCt2+e3rbwm0A4MbDotn6D+v
AvfpyaUpF6xKZp5KxiVVZTsNeNDkC45TPvuP+NfMk7l/8fCsYSf+bsIf1JXBNN0X
Rl9YFgT1qC1osVJUiHaNL47UOpByXP8zEdaAwelvSAbURvs9CaTs1mqE4fZJUvsd
b706zbOpzSOz+iedvFhAWZPtlNfMtF2gc+fUl68zYNYkyMLXd85dsJ88wkOwfe3Z
u38KEuWxkVNq92FtsCt4JUpKEcbTdb3bVeY+sxGWzfstMZocFat9uM+t3Q6agFE9
Ssb8bPKFii1d6TRjM8bOKVqyaE1yBdc1cquHt4/VXql6mYbM8Wf5e2EJ0GEu7yvO
D8bbvEKVS+3Tw5rOGRz8dvOc5KmwRQCfAHx1O6jOU0acDiQcjPJUX+HYjJCMtqoE
LVQSgjJNaSaeiVUJMThc48JgtKsqm70RwI9haLqbIISEg1Ox+rqU+jUXrwGLDoRN
QU+FRM7zxg7Hvb4Jd/5a7IPpC56ySpTZ9oNafyHs4rxKPaL5/l7uFdOuOwQKAna0
mXMhJFobn6+WhRAYeRybdryMfhe5UM+ENW/dFn/Nf4NIc9z7ggzx+0f0pEe9I+AY
dVgrg6cPR5ZBZMMzc8YLtwZDKSY73RMoakXl36NXJEvhA90I4XwLWXaFr6b8AXr1
EneFXSSSEeKgHVmVaargqerqmXv6Z7DoUyzxWCb6+IQxh5REYmLfU80GP8XTDjY+
dbKn/BUDfc/UZEgcLBE7W3ERW7zGuErDROi+VKN52ylHlRxXH/0whsjuNQOU0sD7
EZ9zA3U85s5du5Q3FZ1ipzNfXPlC+wP5q6sC3vuiP1i3WJAF30D70UExr9FnvJJ2
JdT8tv4nS/sgMYT4ANFI8JzH0+Hg+pPwpAghxJ5Ons6mzwNuSQrDT215ioO/LPLl
ZcKfVO64XxiQEnM27aaQo4+6IRXUqjwIErjO5R6+OGxCS6OmASEtcq++6fqavFLl
8pZfjcrynLfXr8jI4gvDeVNAmJledAe+AKb5Sa9AFxcLevAx6ALwG5CQERYTdEmz
l2EygoTPmmFiEhRXBrUUaxfL6+I6ib1Cmrx00Xt/IDqJUtTwLdq7agrU84F7IOWU
+kvKGvV0kU/sDtwlgmVb73P3v5viCo92G8P97C5ldOuP3/eaCvVjMv//cIsoF1VC
FAhzfs8hsyS4isQXBcz4agGc1n+vo9UpGE3GsgKlKvrJ6Tl2mFq2lmJQ8PAVXC1K
qjWU7Qi/WZnkzqbXbd0BwvLgML4cAISoAnnNbyOUs59c9qnkG40cC3MNS5FgXBOH
OyAd87xmdZMXD8+OYjAUS0BD5GFdmliwr9gx8n79IgdoYBMSmqON8HE7oDDjSLOZ
FqGygPSwsHhCdFGGe6xBFCO7jg913Oa/h1wsTbJZbiV65gBxv6ozyl2se9izZ5E/
4m4vO0O3vAhhv+yNDBBry3NqCmq7AcR246SvxiV0RkMnMdksLhE4DZEDzSptkWtf
TlHvnxDN7AKMh+3pZYcmJtp9Bzh6zfgO4/Uo7cnWzaAQIbmd3Du1UqYd3Dig/KX+
5yTylTlvG00lynpV+nsNw8bF9AMVm63NyVkfwA3LbAogx2LcyymJJozwnEX7wuhm
tgvsloeZmrNurSfSl7mTfnrFLc61BlK+a0zrl8dJ0oTow7xUlCQa1Qmux6aeyA0Y
r4d6jInr+NJUHWPoHzMTY6j2QPz8Q2J8JRirwkd6+GFh4Rt/2TLOwEvgedPnQoxB
nXDz3hP/3iqyb0OozIDNK2BBmXzBr2ATPgAfOIVczdavAmvMySA2nUGk12lXnEd7
1fi2D/jYvCrNfQy3DE4s/ePhQPkzCcxsZ8AkhbEsfTYuScxnDdVVV37uXtaib4to
GW7ttMUP10ysQ5LL7jUGLMS+yB89oxpiDOkXyhzjI686AVC7cYwkUmSNFadsO35+
V79KxvqiuH3s4EIEPt0y+Eem911wiRN7/35wkggoKINV5Au5AsTYjjNcDNmhdH0F
kn8Tubw1hRJw0F9rEyzCiWwWCsB3mJWV1V5V9VaVK1CD36NE+7DbMmC5kK9H1LSd
qx5MfHf1aPWn/duvnOkAEHBTX4hDy916hwhzhYacT2hPlg2h+vc1jyl1ovYRCwBi
NaUsfcrgWEna97qe7DncTqYoNfm/408JnN9UswqbTqs0aX0+EfOv2mEh448FgJtW
RZ47Ij3fItttBmtRToN4Dzeid2VIybRDFOKZZU5da42ABGW1pCcSQdcZkpJsQGRr
pRhKtNy/Rl8EKWTBQQFl0MXpvTTsAWiQsvoBVdJx5ZISmts4qX0c6Fq6KjtFRP8U
77+tBLdw8EATGPiTykStH8a3geLPfW4KJvNdaMS/v3AW9BTkti0KZ4r1J04U+SAk
2xbUghgzAa81hsPtlhsd/hyYXcdJ938xsawxZnHlgCAJfMgxaND5Hf7u2Hm+yjqJ
/7+tBT6ymLyVJOY/Czan/O/9w4DwNhVMr7RucBFnJTdMrYrEFT6uzQzshHR36bS1
Z3+AMJL6lg/qTSGC5GfpSweEW5Wg89Qo6yVA0oFcMGqk3bVKYwCC6rPOvOswaXK5
R6WPGhVmcN3unOYudK0mxAYznpOTksdwZSBX9ioraQnjz/X737LIDZvwZy+STGNE
xsBdZuIRgAG/Kpzhnf47s7Btgp8XLP4gm0FaG7VuiMtPUAOHe3r95On7o8hLby8t
/ZJe0yejwveWgcKRzDoWK35eX9hq+HRRwzpsJcupU4L7f5tuufnt5P6lFVBAQMK7
5xGhl7c3APZ91YgNqRevdTm5x3MjWXMb+/IeZDiKE1EAwTtBdfwacZPybuMH0b16
YsRn+ivop/tIRyHMmNNMZdm5oDKyNTklBCW5FjIMu8I+R1cUbh+xvLQGYA8uHCs6
5oWQ2mSzeA1M7SyuZWaR6xUO4+/+SyTPKRkbGdWIMvaEe9taYCJLgNkrl9b5nBr5
7hIJUu9l+P3BDzgXwwYlQYaLeQMnW61iH4wHm/rwcDGokLcTn8i9K2VBRZ/K5ws4
W4H195sLx3xlQe7UeLtGk0SgadQycfFmvHeilh0YilgyFnQoKJAU6R+Bt7Z8X96Y
8JugYls+YXNC4Qr6yV2mFFHwhD6AXix+aIbciydbCxq46vd0CNyVNM/eF1snmviT
Y13qVmmw7La5Ff0YvdE/H9XcpSl5cdN/qS8mys8hj7NqauqhHZ/2HtZ9P9vLjSAF
I+9hb8swAzcKve1UpANXhSrAn1W+wug+CKHYukh3y6yQA+hvxENOQxSbNa6m7Gum
z9L93LQeKkxdAfJAQKS4A5IbdHMgE01CQ4zyEGBc0UfFPtjVIx2o4kppmkAyHbHa
etkNBkFDmTcKBi01ccnC2TLTFABnuQiq5PK1iCLfmmZ3rsAYtQ5pkzvzwkc+g4eA
vr+bv4bfdAO8VGNDIUSeojQ1vid5ugmsQ7rpP95frC0mz8ogiY0mde3Jb3SdCK87
8WKyuRkp2wuHFhwvO20ujkfgQSWVOW0Jeoym1rDsb6Pla0108WJR24HmtQ9GYciJ
l2mG0IALLCqYVzgrylTPakbvNGtoQwjN1pdvgpKI0GkX8g44ZdBpf0hQECz8uCl8
LmSkDPt0DlIjIXsAmMlyhgMhCmY6vyLbAfqd7fE1CC8=
`protect END_PROTECTED
