`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KYliZpVkNGYoOrRWU3oLh89yAqjI4P8kHP9ON8iEh1oD7UO+kCMwQP6Xd50uVYvT
AcskYNH6x2Dp2+GoMSfiLstsjqeVdpQgZUtxf1X31EqvA9YZpUE20nIl+wxeyar4
4aYoxSO7AKxYrnDTygp5mIW4fYQr4ODH3K2Nj4Zzmu3drpcsCCd/Un1nop0RqYqi
IgIg7WH1IjPU9i0C6XIZmQaiF9DIoxrAvX3pXtO5sewjfYp6QL/EO55G2/mglGia
mb4TiRc4+2Yi8BHmEnhoIn5RA4hKMsBgXetc3th2LhTNKxkwgdlH4SWaGFtsC9CT
Sg4rtyyNIAsYJFR6o9aY+1oFUT1uA0InlYMcoFyS2kMSWIAcVOpFSBY57sjS25j7
PFkkV+sgUeJTiPVGGyPXZUgd7umuNsUz2j5LDRp/wlfdDDQZ83hc8u5D1tg5Tthd
p7eMlOsEuZN1gdXe9sw1j+mn7ncHg91zcPAG5crh1hl6/e+m1MDMccotssnUvGC8
NHFlsnj6ARN+CROsB7gN4/DB9jy+dqG9u7sB94rsjMYeD/Sx742OOvq0owWSHSOz
QHcFlHWRLPKDdwdmjZJX/oU0HhHj7wBm4fvEhSz5d+piP8yZSdDUE3Cqvp5nKj7z
oG+MYMgPx4YzQsrSj8WAVUtQQJGUCgzXSUvtU5aYvZU3+YPdC2iNyBJFaLybzWiL
QJV1JbdFlQNFMg89R4NfB1oVAQNaQQ/lUHNR6P4IiS3zhVGhDDvNMcwG2dlyOFfK
TTggoZiTdEIAJvPHmTxuiw6NsOZkcKNR0bDvu0yMkD+FCb6oLgL9xeOBUVmpQegB
0baRNhuXgPpTy2TXGH0ujuywzYYlHTBqjZ1DSxOKLXhtFqqsaWHkniYoCbsEk/vo
sysJ4o3S2CqM8UZt+zafWSySyn4DWe9kpcyxNenWJypzyhYZI/Jn+ol1mW02MeOk
n9sAldi8kdbHVMYvMMokuH4Qln89ITcbfOO138ZJ0enGZl5l0vHtyKkuiVqh9/NW
8j+mS5vtHHfEFkBSxFwVHnPiyN/+oa4N38z4MKsC3GhIi4at+oC1kOjTBia0VKlY
+y4lRkPtuFMz52J0pLg/yDdBjD8cr9fuh48rMVlyIiYsz8mSf882qmraLni3MMyJ
xYsGemqBg77pJKL4hP/nNPNuSFX6/RJLtR+IGuJqbZt93owkHPqE6PBL4FLaADQh
kDKsoPjMA5/mRWJsLlN1z3Sxsj/09AsRwjboQ8VJxewIIn4ElHmoL7l7lWtOcmy0
qgwR2FIEd6ZeCdCCckxQtOaIZ7jeQ7D5/+uoFsKk7sqKqXxu8LC97b8vXT41XiJi
BtiVMq/WTGZqdioj/MM/QMs+PYgJjWkSWz1jH9HKqi+JJ66ZjcM/Qs8ybXCbK8WY
QoagkRLfvqVDxWacnXMX8Y0zeSHedRIqxD6U1ByYmpQ=
`protect END_PROTECTED
