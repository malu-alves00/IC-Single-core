`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7t+OJCrHX97TTZauSF9B1lJayf3pkcv1HTmnYnSEiIqQEu00G3QGUpPhv/MnBYAf
VSOBA1LrHjwti9DHEBSksEk1fMj9/7xjaoE7TwCu5XTKp6r7z+QHpMNcM3vvhcxh
gk23RyVbrH4Hos8Xb/EwV7u1UT24uLArHVuCeClS7hcdetO/tSjeIF3LnTpinWgu
hwKxvTr7lWcx5qBcwLZprqCzT6Kq0jnRqNK29AKfyUetOP7DepVG7vpKnqfQBC0X
QwhUCBk9FOGTE86YPrTbDtEe20NI0JKmEP7AdW2ae9TjkKhKyG3mtd33kYyJBG1y
Vzltw3v1iqMYZ1GSAAIkcRIebmRxDaS+nKX2EBvhl/cTuN7zEqRBOL4+TtPWEGT8
k73cqGxqFmBMIr7HOZ+zpr/04TaDkO/Ki9/eHaSztFFPw0hHCgzb85bcudFeJZo7
xWzstgQZcq7iGxYg333BJFf1wFWv/RcV13s0sWYTeepuJIADDe2U0soTsm2GAW/2
VQMvmkrcL81PSlZ76beRlf7/qwsuDbE5l5d7sUxOcw1sLB4AgO8hEemQ4RsG18bq
YuIhLfdyEYEBfWCW5nBM8yuBBEn0jbuWSdMLCZSUkX/PVveuSc7M6mPo8yXL5bE9
clk2J1G8KvZr/OdFY3fLnUDOE1eX+Vx+cLoDcWEE5RVd2cPqmiq1YE2/kTFCi0YV
npeR+JZNIWpQK5FEKCI9MltiSMuqWOdjSN4vjwZqJ7kwGGeVNN3jtQ6Lbhf6rfN+
mwpqBN6JLa03GB1uIMkLH/n+5hPLq1GEPddUwc0TTf18Ywkx8J+taNv0sMDczCCB
dRxC/jTcHFkGNcaE8WJQI8I1DvAFrD56vU5TCXQ797EdZwPtlIym+IHUiAtTOeqf
lnd/p0FFJvmGf6EIkkaiM2O4y1qrAQvhSjZz80wAcgXINS0l7cmb5lPM5p42mKzY
Xv/65wl3G3mEnIDQ7F2stEKV7LQKqO43Ke4KmM4SoQY5aK1hsX4FWMAaHxGTB6E8
bBe0CuE0PDAjXb9Z00B/R2iBtA1jjnxuhf3y0Ok9kpfoBau32tJMY1KNe/6O0Xkg
3BES913eEX8UECs4AK+c7NPMslc2uc8Z5B03zeemZwpKu6oB/3hbWudTAEj2Kzca
+hw0Y0Mr9WQAo5Z+ss7SUJrc4SiMcHYfKnPizeOQu3RlhiqpVmy+/k7Y4yB+/9Ue
XNBUMkyrRK8191+pC+XWMPO+ATfd7zLNgRWjrNlgtKF4aHQ+/sBpo8okGud5e7OM
CH3vC6oOcp7dTab3sQeX2ft0LmW2a64m0zVCc78fYvp2KEqo8UIrpkdgdZ75T224
TEG6fN5js11TSY//ZfzXcFBgBKsViCabjyCuUQagLS5C/koNLipjFp+L0Iijghhm
eb895rBe9pqlanzc1vyTvuT7hVBjJHoPtJXV/mBaLEOjqJe1HXheXLJo6uicwHd5
nGWfs9Hy4fM3cjhxcFBKJQM6nRi26t+5BWlXQM25/nRJ5nPU1t4nU2nZsdEZa3g3
1KZ9UpvbQuEtLWZS98MF0gmqUmDfkGW+55vLWjT0jfCBbpxEwFhnMeXb7myDAfB4
TeBf3mVjg6KZS1DUJjdylJOM2s9H+iAIfwpqGRzPDK4bB7dz5mjdZm6PoUgvNgZB
DLQN5C2yoO9YazFw9JLCqzpNJjmOkQ1+8kLaIrmBmVgoaMP4/bWueh06XxbqrdgP
YuXbQ22amzuyXHCjqNin1pHX0nlMN/pEUKb3VaYKwZwAdKC50eVFMs6gUaOmpZeJ
vZ0DQc236TmKM68/ftlZ5RPrZ5uavEOFG/+hAsAg5KrnbgUZlXKtrdAlp+ZhddFK
hMRY5YjAET4Kj+PJitGLUC7t3fMxtFHS13+jWrmb5PXkRosw4M3e3M3oIoOlbyAz
JchzVyIWihWxQQSefEX8Npr3qKvDVQ9UNvWgJzejYBPox4xVVZwsfovQDqegL6lt
VNUqdQ+/oCxOwtBPNp39+C8bZI3pKXorzBNruuhyCeoIAwwtM279BVa48DKqa0nZ
Ut249FnjfVRnoKxUx1tFeSbNgifwhAkT0GG1+FOXKzAwqrhzyOnc3IycyjkFsJoJ
04IcZAwwk/UI3cEpbKi0o7LwsArvCshO45Jxe7kjatX3D53gDEodOlVv9dDMRlj/
9AbvLbiP9l1GHNoRWk2Qtsx+/A2612JJ/Zr113iWh0QvDfVgvkX6p1xS6Qm1gTaI
Oa1Q6sTzMcotW3k0QsnEenuT9j4Fas8y8V4KoN+3mJLqkMFJJ6ujtpaHFYW8ieAG
EHzfcrhGbfyNDGmmRjBz8AZAgu4vwJy5UvZpDH0zNtyQtquraEtee+N42E97MwuS
`protect END_PROTECTED
