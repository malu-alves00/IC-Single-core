`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GYySeilyEO3lo0IXuidJKWLAr5ks7w3m7KtnUchGRVt6ahVeWtgahYi4DTDrvhX6
rJ3eExA7UYMeCcwYnF+2MTBlN8FltSpAqVF5GhYgiEK05B8gxW+FvSPAjKhX3GuF
RxU0TJT9+GtZO2dcSDe/yLjkZopBHU/2VsRcKVqrWABNm8SYDyLsKxoRdsr2csun
kh/zpF8p2PCyXSXZMPNI0r+PpO02qfNz3zkwdnCyOIpM8tWVPE2UMtZBb4Gh3Xxg
m5PrCLu8LqFSN8aON45fcLyYdhuL+GV3PUENKET0goM2jMuZwBhIDqUa7OM5FRYa
vBJ4i93upoi61N3GlKHd0Q+WXzYNHfTFIaoF9kvY5OZQ9DSqPAfejGwr9m/gBQD2
bqS5/Z5lm+SdlLSA/dJPteIfrgels3DvONsFmb8KuxP12K1GnXAl1wdB0spjdGwU
WQnUKA+jnB8Z7aOHtS45sNV2dKcWsr7AgXpCeDtHVzHisMViPvfENy76VmgP+MpK
v1zyPw8YDe1PQna++kjIoXBq7R7SqBk0I5yo4hP8t749VU3vQkWmtw2Wt0olEi2X
ZvwKKS5IfZPwJ99CXTeV401qRk4UbZ1d2GQkselRGt9RrJig/iPoiHVFiQVxHQFi
NKVpWTmOtH0ykht4yo0Qsdp/trbgskl8EKRgh4Hcz0GWk0NJnfNESz+Xq72e4QUV
xj6pMWcSFV0YYsenPygW43mLcbQJf3+nzybn8CxKGJqrtsjSNujPoxmRjGU6jLDz
FfY1MOPmxbk653r9xEyS+XHADh7bOohvqqb0jgv2Z8NwsC3w3cOidoLHFOUtWBmp
Svl5ipCf5N+Lx6Ei06swrtSXb6ywnXG4MpDwebGz1w7Vx+EH1r59kioqtu/IcPVk
qSUzQr7kjy4CGCStICXUmAeNzkljaUj5GrGmZdk166HSteCLHfgwR1vRiFPMwicp
dYzhf3GNpGAr6d+JUSXrJ3tOGLv3INV8RCS3whEoTcwSz4ldsa+camGEIpKHNaGv
/5Vo0TOZH2Tn0pJMdbUbkGmjqKTmskSzShqlbwmNoGquZB5ZmuteNtlEvV3D6Jgu
UBnEr4wBvoTs3sJJNEx8JddgYf0CnO/ZcbkwqlaXtBJf2uJp0uKs2AUF/2waESD/
51LNIJU9X1uG6rzDJ+ptmQUxs22oNhqlEuPp1nE4OcJRt3WAIm6LlqoQ3q5o0is0
RRL+TYyLev93LO8jO1aWSaK5k9j0STDwioxnp02FaSKa1u4Ffh8gck4oXyKdQblJ
Q/TbedoWmdoLZaO83OUH8Oh0Hdsx8SHv8K8RNCpITv9tzntBWnAgeSzyXANaorPj
63XP/kYjY0/HCVaT75/MHbUhBHDtnoEfd6tNwnRXW7c1I7hArZriGizg4xHEFDPb
F+5sbGu/556GpeBmMslI4z2VQdGlUtyUTLkmcV7a4MoZfgcekW+bI476maepgql8
aLdAAm1yihqVxTp+zQunyPyyyAViAqj/gxl/ALQYvhXknUC8v09Idam2G5eqIpLl
9vbE/7jPvKWd+K4YPoY77RR9Ah4xL50JBle8qHlyJbQT9aEOQXAFN5aCIdhB5VDW
1tf9xDTbVl0qI/RxqWMRtbMCmg/0dlvQqZIH2B89HxVIFPhVjcmSmYXBysrlVose
yECUUWapLWGq9fPpLTYJn7fOMPiTnhE9ReYfvPrqoZ4Zw5dZRk4xLObiHwUTxaEJ
icRAXUI3meb99h0iDok3uXEa85+rDnRVsBpQzwmQdKa4ebaTZ/tx15IZjyCCR7HT
cQC98pHTheHRMJHiT2bCYENgf6cGIIU7Kjr142aAh636rP0INkMYkoEzRMtT0H7Q
EaErVvhVoqxu5IBeVWyyDGaR5SXHFrj6nkIIA6pWgdcccOPiShfQxirkPOiYHLIL
ftk1JZpcAtrRW+391mYZY2+rczADcD6wGur/L+eR0lD1GAK4weFFFaqPUJDG/go+
Ij3pxWlVb9ZRhsTZ7gYIAFhHPclxs/XdeoqZ6l6xHgZGbVGFL6JGoxcFQYorZygf
JUG1ABf6qxZx/SywWBi0KemOJhSOzSalyLKGLkrD7CTSPgkvoZ4GcNLmZW17yGma
x0Z1wwdOL1eKwzRrkgAx6VjoAIOvCGKspsDEohn8huBWqw9Dd8ucs5fFbjeMQFCX
rkbaPjmll3sVO2a7nCDUuB/MGGhuYOFo0+6TrMre7KfEXqPYuafpKkeVWXnW+gbp
rPyB3Nf/Q558NXFb9mkLZ11dNFCrInXajJBKnEeE183R0eJNyI9PCAYx9U8Ch+wj
3PyjAZMeZ3M3Q93GiJuBKHD8rc+yrr0spQei64Xs9OOIbOvtKhBjNv49m5s8QXeM
7+28qXQi+Flm2uwGptHlBZXl8iMJ/6IBCTjtm1EEvUb6dkCJuenNWShdyIIBd7aT
q/Pvsr+H0XMNxRGktIQcQeHJpE4oY5l4MMBMKEfmDXiLbT0wVwBTHnQKYr5I0DRj
YBSClgC3rCMxP92WI81RYck41WcaGVHPLxQaeSPFyXQcRUENfmJtcmEWvuutdAI8
yKx2uKJut/xGc3pXtoamqPpZg4olxdlrn9MIth3+Wx6CmQB0E4JdjTCmGoSfLWKv
6w4etQw+FXUXESoiBtEz4Y8f+7gC3atm/eZlIIGNv4DeLN+tR6lDEpqaTI5Duxln
tdu7/x+L1WMCwzYuVb4UOrOiRU62hAB1pAevtCGFtLcSJkp+eMaU0mXHo2pWUrIx
2AZwDXoSYT1qQv9Etoqi3rs6FJ+ObBiLPNxtHrDHehlzjXzfRQQ3AAvLzp3y+Mp5
87jXvJ+TCvFVY7HmMTqbRozE9vUJnO9AVFxxhwthj3eezMCEFhMl43CmPUBll4nZ
zqn24+68lhScGOYIQPbfDux64+9V9UmhvI130RniWq9lImjyrMfbOiTS4Kn+IgHc
97D9nWwt7CGafwH2fuep5OHh6uY7c0fmR2meeCPMLJhb4gBdVsmKb8mir9MTVu4i
cib69l7aD/iGFoi0t0RUtwgYIeIs77MgFiAfqT0rBFPPvFz3ptSo4O5ktiNT8BDI
ZSvuK/ZPbv3MtffkhUu+Xa6/nal2RZwzjjcrEZ7gTU0EIBtMqfk64YEc+Jp1GdEs
C+BTmOCApZ9034ZexTdIcBjBgLNZ0gky+WjhfbFeOZi+sW47MKM/ffUx9/VS/HUf
nMtDMCmxk+mvnSyqZ3PYJjURwQhudfVBJKhF5voA2epfTZvFOuvQqgU3+ceMNlVM
LBJHG+WW2q0z7Fs6iEC+sDEW3vzRkJNs3l/5huKGiyE/uKLSFYcJCEsO6kjIUZz1
4sDjgmvbK4G7wHF5eDAGj7C9n4Y3wtb9kMNEdRaIQJoZPR7B2MAzxl+RYSnhksSs
jyCh3/ruKvQKn8ppiNA+f7MfwS40PBOGxidW9+y9D/Y5rJGm/Ukhproka9m9tpns
0aJy9zollF9GMFP0cnWYy1ikznKW/dLE/Bmg1jDDOtNNMRYl+4PNTk2IYi9MNxaL
t6DpdZX4inUkVdiL8+CfhRvDjGjaDJOlFetDOjBsi6SdKGWHl0HX21EzFWY577Zv
VMPUsCOyMFxcx35g2TQBfn2wMuwDhiKAdnmmkf3OkZeL2S5jPtBZvK8FL3m8+Dxj
sqWJmYdkxgztjI3pOQWs5QH9RNG+BsXWm61npY6JnhULFRArJDYoDcvgE6n/hHvw
ZtYf//NPK2kzyUF84IToRyvA3b1JVUK1pxfTeXsGP4gkHilnxoJPdw+InIUvlfi6
iW4NyQz7egFASE1V9ECmUI2sKLhl7K6IjUnZbfVPuDuhjhMLi+6CUFhFcnppqG9U
p9KkvMmHhU3golbZmFSKO95HWNBVbYeDEZEutDvXp8MsCw206UCfypfG/415M6b1
dSVIw8cwAixwomM2VxEiEuh4j/lR77Wdkv+92WP4SYrQX1iayQlo1d2V+i7w4SQn
FyDafhbx1vSjsdTaLVroljX/kYLbKl6MzCI8NzMuA2Aw4aO4RNq836anGiJyZKJs
YtdfqLAJI2wKH9H9EwJXA95F4hIH4UEtbXXswb4mkwY6lw/qckJTvv3NVQNicyIe
s4X8wMvZmcNCGGfR/FG31rYpjEOWFoa6zuCg7W6EoDyADksffqslNucDRPX804Nh
t2zSnBi4FtkbOYUm6YHhzp9if/j+HKyxonee5/kJFShPdZqtD1F37XIJC+Aknqn/
QSlQPyA0mJtAnC+iDuv+IjD6LB7zfLlZWnjy51J/yc+0kdH0G1JYqvp/fdVW0QyN
vVtLTyStcf0WAHuJCyLOvFoLEuIDwYSbzx//pj+fzd+3sDzA5lzU8g5uYJlpmdZJ
a6lb85WBiYmq72F66J/dniF0doOxNWBYTOdBoqXEhDSnJOMJCW8WeYTPn180yMW3
TUv5ES997cW7bl08EsTYXRhDueDbFesisybpktE63GEGcZcA7VjgR4BVAptunqPU
/IeID8to0JhMx2eVJbO3ePZiHm81Aakemk3s69uwUfkZpRG8aNJ5vdO5sUES/xE/
wvT/Pg+js+slhBYEAW05JFbXlHlZL75xInxequ87fS0cryTnVL6uY97SZvCs+Yj7
xMx/BAiN9tP/H6vcYVCTZ/fkadbWCkYGiuEbobATEuWFP3fgS0yX9UaXqw/i6GRw
qsjNWRQfJJjtD+ukJxISm8A1aAc2qHdz66MHto0FGOCcGmKtLOT44WFOyeppybA+
p3q4jiARwpHRr96VXVN6lw0LKxmco1rky6Fl1+Kdhxfrkh1itSf5/PdaiHO61SaQ
7W/YQ/8Sbkqq5vZrRNZ+HjFLULo6dzpVN/X/iQqEoPPJFLtePebxu7UkNAKN1D6L
Wvkp4R5jvvOUsdxYJ34tTCSa+ahLB1jmzRKDDoAeBBeD+jQrM1JvlOQLLwnZEFxu
g4NBU5nQMi6p2gusHTkXdlEiTLkR670bF2x51WAFoSGM/pgZOFjw/1Sh4yG8iNu9
J6irr+i6V39pY1sVk+ij0nizYaOtFo3MTWvORBmXxD25THOcBZxH20O1Y7yJeExm
vMQ/snFpn+YTTmNMlv8hbriVW1yEoM2SE8GMu8Y2hFVIsUezrI33+SyjOpVrB04I
rxIyRw9enVu2IIF6E+Rps+lPKMJpG15N1CLIgsffIO516m9RYsSA00IocJDeTSi0
b+CiOpJ1zMwniZE0vdu8qzmPJVgB1sz8/D8Q+6C0XD8ahQLzB6igBQdiP2lNE3k/
C8AuvtMOS3n+txD8dok9evD3VPzd4XmvrX70bgqCzzU9r8ci+ueuGXC5rXMRw8ey
oHZJdFg7lE2fzfvRjGluXXRWzw9jNde3utG3krX+BOhKnvy+K65TRv1P4j5Frbtk
M+k61s4HSpDSzoerExTvqudlfIKZOVTEJfj216nIemsUsKHUSUuw9ZcRk3/RVw1q
KxpkuxzGPitgsqntL+CXkpEt9+SOpSMIS5fz4u3ODGRX7GoC405mlX8XogkxWdRV
aSrwtgP/AtAPFWF7owVQHZJd+morV8JWTvs0co2i9KuhG99fkraQrO7rdS+d4EBv
NxcpKLoZbG4zSzA4LlIPA75e1RpJhzBeU6Nq3uFQy2pp5n5YQOp+0JtTf8nfPZvL
dmTyZwj1jGB3/6MtiQUyyT1NkhnxP/slrWrIx2wWN9Fz9B534jiSVsYdp4FGdp5p
c6nYDxy4cDR0x3S/yWTosoW2o0ru54g9YBVCXHXO8M8056Y+NjTJO0uO+1DklYXT
SZvndq3uF6I/jkOFbwkR8cm6D4EgI1DaJqpXoEwYmn7m3Bo7gzTSc6t+Tlr7Y7HT
6bNPgbx9hwDP3kwN4YqPTgrUkj8z84X2oFhuolW4DMVgQrwKGOGtpoXQusBvaKHI
vIgE7Q3lAaZZj+4fJW6lBx0/dVJSdCS5zTK17YUTNMSqYk2XoyZw8dBUm1xOpYbl
dI+WXGQ+jHTbvgnUUZ2ikCx5D66ZeK2/iqcdXHx2B7XE3Ymgw6WDDERUwZY7lpz6
YFj55N7tv5oGkr/k2iM8Id+dbB73IisNtLLIefd/+homT9e9CCk1LAianaNtBYAM
n7VALGo6RAzol97Geo7Nt39I10KCkPfG9DhTT2WPUaowbGwusL3SiAfx23yW+Gv+
HlovNvDGLyOVGPfrTcx972Wq3qxQrt6XIFKdFmIr0RkU8qKL/7Uu2KxUBxVVtXZc
nC2x17rWKAvJzCKJ3v3bODK238ErL7XzaH8kyLdSsx5omvQCKFwami379UliIRmW
2AAz0RfRsysGFfW/CYlv/3HIocuJuHbWpWP68ZorB6Gylo7KcleeD1wG2JgfeHUQ
dqcPI02bjefn6nXPfc5pQQ==
`protect END_PROTECTED
