`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YfTXUZZKr/aQO+fry3Dzt1avEa5GAz/E8BO1wGlqNOH6N7SvjebwZjzdb7PAPRvu
Bc928Ka82H6kEgsyl8OioaGiNbM76zTwpY37S8Bx+QVdM0x3c9uuoTSNUxRQcQyi
PouUjz535R7xiMycZ1RDpV7yj6Eu/cV93+plb58S/G4bFg5HsnKX2uKitcxq3X+/
EdeOz69XEr6jDybmVyxIADu429n2Pf+lNooQ39splNa+apgRm+RnDbP3zbypWOeD
NH0vME0tY7xtbWfjS5fE+CxXHRc8HMLQy01rKcd31bZiw4R5AcTJcwiDpUzYSjSC
kYF3xzlT9qIQbWE3LGEFpTaS9tndhIT+95oHqX5XZLvY0XMS2X+PGpijMtqOHViH
EYw13oLKx/kkCUtlBMCgomzjVKraHS78hV3BhZiP/eordkZ/sci0oVqLpq39BTbl
LYc0+QFCyZfiy0UOaz3SELoRapfe0C8yRoLOlxklvkKdX6QCmTeHeyJSni+i3Quk
UaAIEdL+wrbIAyIib/F7i5D9Dh5ok10RLOwBOa3/HZuSWlwGwO9jUXoigDMKCIkX
4XES57gR02/uUUUpaoIir5HI4VVRLdSe4KW0/pj20Ea4/7X6XVJAfu0xnTDLbIoH
YWA/J2SnF/49ohghE3i7S/j5l1CjZCHMB+3fsGbwPc6kYbdo66l3bsXAxDumtkK1
R5JkUUI6aIUTQagAOzRv65wNuAdupsYWUT5eYdADNYpxONA6ZXsqz60Y7xQBWemi
8cUq4OLYDBHBecOtniVLgZHP/Ujv75GwmIz0BqpoBGN8Mkicf8qgN88QfuoZ9NCH
`protect END_PROTECTED
