`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2wrBh1OIHo3YpFX5c+YrVnW0Y0RSYYwG+yk3DUz1uwuJcMm6zcEf5/MLDI3m775w
0EKWnzwMsmlPVa/QT1f3j/bvywCJ2NjNCnNCnNrXSxCakJmTU+kWJLcAyDhoFdzB
4hHNSYn6p/M+brrrRrWq3LnBVNi9gQwpOAUm0BSnjnONLLCedWmSwQ7Kcc3U7ewZ
YnJ1wckobH8WafSMmRLsRiuL/UTSgyULTrIAfIJ+tksKMJJxCZcFgMueai0UoltS
x7Lqyqc9zesHijFJnw3hCQskiij0WuEQgvNl11bg4osccEkZEQXav+uCtqVScmcz
ulvOBdOs9q6mVSTRFlWzU1IyPOHj2HwY32bfCcsvaLaLv/szDrg3F1SdH8MSLwcc
duWGk1K9lL1hFwmqkPMBy7sIWdBNg/7sNWIaUM3JoZsQ79wv+dxO6PiilpUXPuUs
fpqgDPuREkk4ogmcct/jhmZXUs3FXDt4bIyc1QxnmDXSymkgpPHqG+s187dRHuS9
PHO71s57TkdrE5IicYWvCJ5uXs44owLcVQXZxaqyZHeDVRZW1xwLIP7rrXXOFdsC
7Dsk8NTzY9oVJwyT+HuEojw2zLABFG/1uQ6lW8+2ZE+B9VEq2vY8RuKnLA0590ut
sr6baqSU+KPxjj3uls2XydqgaDzoqwmp3rEUVyYlTAQaDyluaEjNenzLzsfYV61O
zdoSy0TpsG3qCywQz9Er7m9t16+KXLZ+/d6Z9/LVctkBn18gwQv9DunY2HbClQrB
fiMW1NzS+6U1anvb8ih9VwOVc7yZ5a7SA1+fGONut60ETqZgUycSNw6fgMN8J86r
kDhl/bVgTKDoPZQbn+4KIQAGK0IJxEW0xMtgl2mUcBovsBPZSzYCu0YkmlQLFrxY
9NGEhXwtHismbMC17abewKenLxmIIy95zXUaof6+dOk=
`protect END_PROTECTED
