`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mHpNfCPktC3jn6mTrrFqthZvrwCO2/QjOH2ZMFjt7woUYnaRj7OfLDUGlHotNu/Y
09HdjOh+fAvJBCCIRorqzXOMdxJPWzB8QksU9xQhHcvKyVTuxGTNQlp90xXag32L
KD/vfL5BXK7p4IZLaLL2llDIxto1lz9qbd7DWRDX0euf591Ye4z29QFTVKmKR949
d74vBUCYhuRGjkUMGLt0CMwEQ5wfF5f1s8wxRjjKvzYrQqxpVrGiXMJXG/e2Tmgu
XUps7DJWszNkltFvv/ppnFWaZtciprylPmQ0qFZVHwXZvuDMEhkXetUxTAuNCCPq
NkvJpWSVM753zHmxlNSfgalvMI7k7m36+WN7aqxx6ZXzn3r1T7FOSdYo8ADHOOGc
2mbqrt3zN7CPueIV9d1ooS++iEIpwKbC23iXGHYwpA+zubHdDQgY5Xuy2WXKVfSw
`protect END_PROTECTED
