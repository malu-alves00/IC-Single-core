`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
19bDu88eWaa/QXN7vFxVOfABqL7nQzhG+cgjt5wJKdaJXMZ/oWJbcIY+IICnruBR
3w1ijaz9EDGc0OQHbOpWshjygjyVmTylIxqpW0S5bWQOgOqvwZDDuNa6zxOJLgM9
WwCzDk3QbeIu7f6QV5MknI4YKKLfWboHL6ajCaApUCNX1GJGqg1YhUPjZ/sJw4FU
+bOt1ugE7q+LqRNVhh7mGQnj0WE/Lsu6IIQRb99Topm3lHZFL29VNNPu9Waao1KY
D4/NopLmRcmQ3aG3nSUgjUUVr/6GNCLWr4cn6q335fZ4KbhDzfRonwHGhccHTCfM
YaN56YT7VfUOKoWBgJ/QAj/EixxlU/jzOdNYtf9gvw31aVXY6WjRJ53woOIshgs3
EqcCEKIwIc6bZKbrvzf1oUD9/xI52Je/T65N+yuOxby99PLItETTeSEWbJNu+Knz
7FNyKQNDB/zY+A1C/koxPHKkB1yuwNH3VkLqdzku0Nyt078vuYalFTwaDTFHEuYr
U1/cxrss83KHYYaeZTF+aGvTbxQ7fuWSXe0yxLYc3vpnIshn5aOC3K44ST9VSTnC
rthCeYwYXwPK2uVNaJDYyw==
`protect END_PROTECTED
