`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BXgSpKsh5n2D7RPSWZ+gbU6mQY3TwfBdX5TdehJZxVqHO91fAWLZc0C5DjlxApTC
7rvLH7JrRGijQOjeqYVAAPy2iifkdbqjBDWLb2RBMmF1wxQMCeJWjJLaLT47mjf5
CsxLKjuB6AwY47q8Ki0kijjkFlHZlhQcUDuzjTmofBIikTuSh2jQvp2ufWhSawiZ
TzTUBwv2cE9RngQHrdqWhIM+PLJJ5JOL6u9wa8568gXO3lEDdAJzULRJOEubZljf
AO3nxCYKO4zbOIGw353s2SvIlWvDkc0QsNLJdts/KkiUNNBMpg5r8R/O5TcSWFeK
khnRey5W7v7uVI9SO4Egw6PveP6Tn1QDNSz60Q/0tfKRMBn91W7RTJ0IDO9LUbFj
RNAttJMQtQy4hje5tK3q0vL8Ln0i/5Bq1R2CDB37VyGPqmEoP9m24vd9ClkrPR82
EANKk0zpoEp3Dnz7FDUVQwqPiO7NFQdXdaGdosU560Ok0Y4euPOaMaI3eUA7+pZG
C5LCBPH3UnGt8Gdia7rUg56u1kI7iAAwwt7E96nZFFIiHRAqfBrLfpN6v72LxnMc
Lo7Jk1lMms87n3VlolB3q/fdR/R4AJGygBBBkO8VyhXaBVRn0aIvqC4DIWEuwbEo
96NDWzr5ERdThfvhx3FhXLqUNL5GhcCAgtKyyeFVlBnVKcIeFGwpPizLRiRVR/5w
41JZ0DHQ7pQAkUYV9INoIL55SxqDZZJdVj2gn+/iyTf1rcPOSpQGCtKalPFsd8er
Fdw1cLB3FZS5KKuP8fQFCbTGCoQkVMcuCLb1vNKYEBmyOxOypsTMjI034I4/SwgN
Nn9YIFoBxWtfMrKRSvSvKYjTa5+0H1P9xliddvy1kSUG7axes6ugoWOhi7QGwrfn
cJ2JUBTDqJ67YC/8EF9H56WpPywEzLSxOcduHjTJcaXfUwJ5NdW/N4RvmAkMBfpB
lsCD/O9eraWo24dPtRCLMUUFJS/C43OtkOZD0PA7p20/duQWyJUssHqEY2SDP6lS
O/kTipj7mIjiR/wFh1J2gK5BG9BknV9EmiyZ91Va/0LwN/AcppBMTTe7dIPIYbNW
YXmdNLu4vU3Ows7IxU6OTntwj7jQrWWAaZQSkztIYAnIP6RWvQfp3ekqQ1FYObcp
xPpQmLy+mYhkJ8ZAOz/n5RCy7X0RGKWK4hSVu2mPYZOsM/jD90Vru4wMqId2/VKL
ik+8klQOYPO6glCyASV5fA==
`protect END_PROTECTED
