`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PTO4dgWwoEzwd/tPUvYhIjcpkNmlcP1eLE+j8qjnFRt21e/X5PLfZSrXT+wCLTXP
kB40IDvisvJNFOntcrviHhCfjdiaQG5CMt+m/3gXzmU5xsEPs3aKmfB2q14/OlTE
SSqbYLekkLQub3bRuZ9Pzrsb1z/seFEVNxkSAw7UV4XAkFUBp/b8lodi5/jmAf1w
qi2Ig8lNtFWHHF4PWWx5JvYWS2u3YXetQP8F2O39j9VyL4AeftTdsQgF5BbZNtO4
D/pkbVD2qPhCg3D+IIz4ZOnCx++rBGbRiNygwcGBM/vPPP0fb9WQW1qd9e2EXtdI
eMa+zbeFKJQsb4hHCQGHlC1cHx8l4NOS/m8gXTgmpH9yWQ8RzeHuO6uc7ipMoU2m
EWG30x91jIL1AfOD8ogSLnJZtibQdw3IcVN9LKfBosm8ehNlbqZXbECEohErCgwd
2gUcsANKEvVL8GmJNKeBwmbAJ6DSMrJdEALVnJEf5FQq817WxSWS8B2EKXTs9hMR
IDDqSxUrq7gNVsqb7ZB0/sY2unzj501D2PRDF9h5amgFqx11M03TqasE/PqRVqbt
mEVN4Ry6Jy+EaC+E0APCUJ9E5FRGwBjH8C/gykcLdwciEl2p1MKqUv+7GTI1N9qw
CB8ME1DN5eihZfqfMiV49BQ/SCrQXW5sfOW86gABZcLV/AOsrycZiDx55swMUfGy
csrdX3VeJtq4uzs2V0PI+Hn7o+ElHUoyQPI6enw3nX+BhtKymK8WIhecV9FUi8tb
K0cWW1xjBycJ08UypCUAMOnosYRacdd8NoIVdu7JIt8Xf4WeUIosYvBZrmP1StkM
d8P8WtLJppR1P2j8cvKrXQJrWHaEICjLw/qRxFpTkNTiXi4YJz7+9cYFQvaVlzq2
W0N8JqBU/0zohKs4KFhjBdE6GlPJYqaZjNKPIn/wLJCWkplFVpFB81bLeQdf/1Zh
lGj+s/jPa3E7Zl7nMgfxSjoSdHX2V7tNFEkZgHDVXUQ=
`protect END_PROTECTED
