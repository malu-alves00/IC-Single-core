`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9daLVavlH9+2ZGGVHxBdzfkaL3BOxoevGB0Pcis7dkgQJF8YpjY8Hefh/xDqUekz
6nZDHZYOlQHA3pD/742RaL7OhdKEBRh3iIKlI3pbxA4nqJyglPQdiDxuNUgrQetT
YUZ1ItwmUqGK9vppE6Zhu6FUR8BLW7YkFWbE8zN47mfK1W94dMgkolnk8SfWlJsM
HRl34W3mEOvbpdipKbhFa07yVGJqkJaT9JmNZ6biH3ramspdn/37mQoKrD6tPZ17
CBG7qCCOWUrl8RAwjIt8R96gC/PY65cWtOQ43Jh9g2p5nq5/1T1s1NsjIf7r3fbK
gHQA2yKqRdbuzDqm2QPEFaGtkfrq95kV/fqHjVwPXhTBDK5N7C87plu3i19IFAjo
vH2ogYqMxcOIOqfBKkavou2O0a9aU8p+a22Y07/vnDZOA85/8JSU58Lygv3mfCAk
H0xHtVEnRRxtTWp6Y8dv3t6k3fdxY7lxPPjw5kv0q8JnT/au2toEbzfSC/s/ZiVb
MuG6tQN5Ma1Z0ZxtG+pYELucMdotS75/sw1YGS/L04DOJVP+YcVs+v3kAKwtlDnL
7kkM3gl741N0TwkmXmGjwY9/DR33UvKyetX/8qjgP7Cnu/lNRCE3VIGyPnJ3weu/
wGQnc+4NGQ242QbCQDHuU5Hvv6vZ5Eh/PLfhJAlz3JbKKMSqL8J8cZr9lQdkAUTS
NRD0mClLVUdxO/lEnip1u6vB59kUfBFqEIcG6GpbZHO42HCFCqO6yb4IbBDPtTOp
CwFeq1t8fYECxZfKk8aik6km88aXbS05+G+ftuNLAMI9l2gNU8BS6ZEVFeXs0oYJ
`protect END_PROTECTED
