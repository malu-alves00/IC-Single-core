`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AWC+cUxTiy2L0gSI3mvEzcT1/AaClgdKZdTGBBOLOB3hHKTzXZi2iGA40LGJ3bHa
158pk2OY2QVCzp51xiRQdVB2C2FLvtwMPqzhNlXu4QZRau1uL3e+v6yEtRkaclAY
el3M+Dl3Lz/ErCAtnqidJrMl82WMwXaMRsZsUQz4G0n/fHHoaKXq2d36i8wqZZV6
Rtu4HfwpF50gQIbbEkTLZ+Lui9d6XLyk91Xgwif9kYJjSwLIpyAsUX+eXB30YZlW
/XpuOVAwEduMS5g6TyCmwa5EzWEkLGBM2up4bGPoGGmGtQ5Anm8xaaeznmM3XfQr
fuWNLUKdT5ob7DdCTYDrYf9oZq6+Shrju4NxaN9YhK0gG8IGV8Ja/bqTVa2O32Ov
7rYh6gFR/VkS/fR05VLJTh3gF+NBZuvVgYrSBL06z5jMonkh4lxVuBibAXRRSEHt
ea8KopQivcqmjBgVzvzuIlB2O8CCqQdDzMpppvbyX1pWbeOtqFzNMs9wfzGC7Zsq
jGodZwueeZUPgzHJ2dz+hka0R0ejVI6YW6D0VqAO2m7DVTdlCy0mQROyEyGt6vNx
tFxDhK6B7N1pg9swdJr1tW8P5QRxjwp4eLJJonJE/U6/Jue9a2GV96GGP5IVjK0g
yaU8qu6epIRiNlBsloY6RIzjR9P4xXINn7EB3EcMNMQAbD7TOR51wvfvNfyffuZD
2HQg+4DNEEaI43rK94DVa+EHwQ71eFGNufk9zK/miwSCyaC+77yYVEFvWUnVpfok
PQjp1QNL6QKa7gCV2vVptA==
`protect END_PROTECTED
