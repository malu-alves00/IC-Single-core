`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YOAy8Qs4iWIwzLRjjOUbRLYRR4VBIkeEurLC4Sbmj4KA9m16b/T2xLRapEsJLQK3
iISwRcdeiK0Rp6HFkJxi+CBWkY7tJsONfJkqx1SwEBGEnW0UZuwGVDhOHQ+x3QP8
PZTNnccz21wgFhxZhQ6mer4ozrGz8q5V/7IJwRLijdg7zB5AlYevh2YywNP2i6xt
an8RD0DQmoK/BWS4y+qJpWEGG47zatPe3xYOB/9ImOyWuUOueiLgl74eJlKNcibl
vcrs6tV0MkeGAHhqTmwykN0NmWTFs00eSU+Pa1B9hIiZ/arjUPiAREfCyqGYRe1p
IQsR2EVQd9w1BuFbu2TAOtNx5zB9aKvFc/AW1UoRF9kivQ06CkOmtC329ZWa7YEu
AnGqxXMQkdYGUiJm10eCZ7eFKU/Kl0q0vQ8H3qb1bh152cWV/no+R6eAZ6WOImgS
eJR/KKVNaG3QvmfXao+zF9s4XxLQJm2Jq4XT/roLQbmAJTTOGaC7GHRWsWrOljJc
i0ApPhFTm4pRMEC1cVBiImfKM0ZvbFkKq1D3ZkCnrH8Q8MiRWKXGrQNkBuQ2kTJ4
2IQHCxDtZnPlqrNg5zhFpvK4Q1Cvo2ipB7sqF4TIVxsfO8Sef+T+v5Tm/A4bTqik
0pJIkdfTdYRcRjVFl2EvKb5BkeJJSowxr7cVwa9kKkJ19VbX5uKAF/I3mz+1qoAh
SJuCQMwnqd/IK/mDjN9jmPrBpaBomFSJ6VryYkpRlFNKL27ZtXrEDaeEuROXD4+l
BaFTyLRHbEjYJHxR5d4tOiInM5kNkitKeTMnLrqiQv7zBgkmKAR564UIkKuASrZw
3/hBQXf/VPRI3KPH9l/IfaZherZ2I1HQX6gH9enx7YZ1tctDm0iuiPyo90IjqJdw
THsfCfd+vNUrQ2pvIkn8Yi89c6owe8r2FTYi0FSghZ22cWO95pDoVRbjs8EJFNQu
L+eFvbdgsvVFiRaPwkSxS8P9c0siUqsqmSsbfu8eSY3XGXZsMdqxN0E1qaq2fWyU
XgbXEbhpexaO1kWV9wXifeSPdN8Kn5KN7lsZm/J+Aqm+uIe9WJ38OhThiccJkueE
z2ITOq3xxhHZuWkp92YF4Hue2qYBEkXnr77poYkKFvW3Oxj/G+4yyPPtBEtbDxzf
0tEJ4cZEMA2OoR1qajq/OG4g5xub5hFfk11rSGguHe/ZTBF09ZM155xoe5/Hge9H
m2BLL7SjWQ1MR66pvwh+5BsLozha8Paynm9EO5yZpoimkvQ4xE3UI/4lzGIIRVmx
Js0eXTDZLCQwrRdL/iNK7+yle3MpZp2pWsFhoIeRLnfd4Dlj5RtqPnp/YjfGuE1w
xvtrWnFRDGVOn9wwHA6hI5+9Yts8cG4Qe1PUp6jzmfXy8FV6ACIaEatadI0f9Ius
BbXkwnaTj6gLBoJk1f6Z3B977Fx3pz20i2uCUBUzjs3PrCMOVFYdgNg/3Ysx1y0p
SkCeeA2zyS9u3lAnfCafVYkl851HeO3oDR+EWMgp5qiGuEL4bDvpz3ohw3MvRin4
j3HuDL1mOR669Q3+trYUeBA9bFRjj9IaCR2Hsd5HD9bbeRA+Ps8+ahGUWNO/ju/i
8Mmi/AVXERON1Xn1sUf6hPY3mTCU2nVQcekY7oxOcyY=
`protect END_PROTECTED
