`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NW8zVMVNWAErgtLim9m4tObhO46ZaZroene2IEOysYMjog1+S7o3Bvpg+c7ou8D7
vvdN4rURFtn7I8cLzFcIXMGnGXI/QdKBnSNqsl45FUHhnpM3GqnKsMfLFdyOjKfK
8KiG+lTw1+GUpv2SFVBuDEMkRPuCRTMdeWfXzFLTgxqe5NaGm9BaUP6yex0S/qOX
LRGiK855se3z4bz8c3cpobNG5k7pLzEPQtpzg39OPHn+vPRpbngqwpOfsRXfq9CK
lmGuPXFra62+Vy7vzCH8VQw14BRviCR/naDoAoXXk0JHqYZ3LhtYcJbxmn9bUEfb
WvYbiCJyfy3iaz0WfArh5BPIejcBtH3XRLOtLLxUvgOx2QL4zXQ3GEE6g7NszRlb
9yJSTd7OGryJoCGnvm07IQworwDabLu3vTrNhTOwfNj0xb5S+nubBesgQAuB/3WD
5GWMZ+Pebq4I61CKkKkkYObsYxgX5rz8hVySCyamewLggeswJcJn54cF0HV6cius
hcqL/4SBTRXUs1Q6IBQiKiYJR2gT0tv4Dvh99cwSbrD8+/+epI2si3bJD3i+IbNn
ZzSCsG0mI9zE1IbFMxucT0oiVlb1KOnJBrShN54fHWnZX1qSYZKJVtqkqlQoklnq
HSyTOiKXK+jetlwIdh3kmC4WBxt0i/uoG2jlHEKM4JsjLfT8darup65nK1fEaMxc
HzW6vEWGXCpI8YS1me0dafL88yMF4OhyJxmMcH+XxmwRJSZIJf1BWOShZGNfwP2k
glv5h95acepg4ulsZ8Nz/Xd6GiEv+kRt2pY0ZX6NqBwKrEGLcYNVxpYvuenZfOHZ
Cf+ii6MtXsE3lYgVj/GLLj52p20OVwfdTerVC03F+Hg=
`protect END_PROTECTED
