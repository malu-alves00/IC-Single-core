`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jGYIPtHD2kMkxnHdX7CP/PG64MQh0Z0W7KUTWu5nyYXdkBae0YEkOZYC6VvyNZN2
CcQhLaUy5CeWxU2CyBC9ZMIYBKEs+MNRMHZKTmtZwIO1s/god9PUUqxISKiFnh1d
IRIGIzFPlZ8eNyzOjOA0/ovOPuMUTwku58/H7EPQCeHfV06rdpI1ObMU9iCUvb7y
624P6dmElxLCMFIVAw1+pE6VVcldxOwLK7VncPxotbR5KyrJkGnwCHek9LRJ/GFt
JADJzOUcNZ7GgTpdgCmh4nkF+1WOpngJi2p7RH+mXOO6IAUUy1Nv7Sv0RqKojyh1
u6bDbRMUQOQjgTYU5jzqy4sxOXvT6eKtRBxTut5ufakGTziE+oiCxvaQdSrg9InY
LuKqNmQVlOeG0h2c1Rjy7R47dblx1zKgy5mwqRO1XLg6vLCeCX6QaUJXrX+Rdgze
ko7J/UOwa+EfHMvHaCzrTrjVXmOCZi4twPyhPtT354ymEYnzpEtziHp0wLq8SGox
OQwe/XGnC25FQ2jJyseVmQkOuQ/FoqkE9KTDWoIG9yWpU+UwBuG8o4VmJb1l31zb
UeZa0Tz/YYin6zqdOpBEzfa9vTAAh4bVrudYgbQqWZiS9MRWtSdKL9BIHmaMsdLc
GC2FFwYV9ThKb0gjy7Hqv0sgFnUtLmdUxRBLshXCOrNM93EqCUb/9ESOshtG2CdT
`protect END_PROTECTED
