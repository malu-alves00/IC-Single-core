`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2mf4D6y1T6iFv53yHXMpO6czHp/t5Qy6ml1Zb+N71sT5IsWpty+mlqHWcf9MImFc
GIJNIhtbPLea2oIaXtuT1O9jP0iIIsFPYzkqTB15bJkblg2Rbi4uPIpSOCl9k6J1
hmbQPnZxie2hYOuLLtq3+u1W3Z3FySZ8vsiZ2JksX3vpSXmfJqwQXRkAlB5eOfEQ
wZO7VFppmyvqg/HaO9XMQUafgA48jpQ4xzdh1mt4VU7/5MHJHVO8bNGvXRF0O9va
ePHq6WVycCByhVq64TLRuIW956McN9AC3023cLV7V+7ycRGMktrnpVv5OOYLMOl5
Xzcf4+TeDMTELlJ/RgRew0M67MOaYrSc+ueU39EcnkUKbtmGxlsnlewC/eREzRuE
OJNc+LBCcs+3+P5f6Zhc7KS2SBDJ/MNzjEIjFihPcrU/nGEhbsKXnQe/Eh+86rIx
VB8fuXoPebiuBw62bEUJqVWDhPQ0MajhKWPj6Hm4dmlLsgLBskz39yvB5BEzfh1e
`protect END_PROTECTED
