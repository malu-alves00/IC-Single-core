`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lQtXnt/eoAtTXwpYoxyGXSzjODby3iZQTa+D7IS5ur2xuGwahHBqZ51dPbxlQZpy
CPvgUmD8+TwfHcdrcbxJL3mhWn+wIAOAmvJ5E4OONoIYnT115yMAWbYkiVUE+hLw
I6/xETzl7Ylty0jWTWGrgiaIxDGcW2hA4D+KTGKqICfGUumDwEPH2KJz354gRiz7
Eu4J0fs8jXRv6YkQ8DAnDMduAqbR1NGn7FICy1YOkZTbHNAgT3GrEyU8rhTGai+7
T4gg7aU6h5xrU5dMixL3jYhdUaY55HOuoko4vmYcKG+y8W0vZWVZxSER7Sizwt58
uPY4+vNMRCGdE+hVLl6E9nQj5MiW/N6wVDqVf+0DP1JjjlL8Fq+MYdaIdzjcNVxV
1qGml9a5HbsgvcaYyuM/jSSnPsiOLAmF2grd3F+WUjcbdhg3eNjPjYtSxCPDp670
6nyzCIJcunVwQlADb2DyBA35KZJZhUkbsR4EwkWrKxEwb+Dd9DXOWaC82TTeVr2x
WNmDZse0pvp07fbuOSGoVbAjt9IkFdtYGKf5gTvfbsksvKZRDzswU/b8mrDT+zUR
YfiDnrUpvnCpI+AuaoskG7/zt25h/S5oEZFEWEO3JO7ny0yVrKXNjRXsJMDT8MZR
gapXdWuuK+0ISlvFclnYv1WUCMH4wEDrya9xOrEcFeckKEA3jXXrw0bve/XrjWXt
CJLRlPToek/kBR1TG/Pwov2CboEe5MU8m3SbjGnSNtarAUKmjDc3YV7/dB9HP8dP
h5KgfkaxQa/luG0kTEwUS7qXPgnbIBVII8EGYiC6vXVBNtPADA8pj1zmT/nVSlHK
YWI6dHACMch182NNVxz7Ogtfl3qUply3ZNEN5gYnW5//oNnxDwyB7NMZdF1xpUWL
8VgoQEFOHxwGodqQuiEaeZfPe5TgKIgfn5wzwilLtdIkC1q8hMtUNdBSVx+fD5AZ
nbljWG0ua3PE3UO5VEfcDogMqyjcEohrcCca28VJmmOaDnKE7R7FRrgZUnBL5+gI
cEZh4QaW2XSl3YhvLJWIKqfHgqx7B1IaS8HlVTGCnmx9sO4vh4w6tTRHFLcE5lLt
5DbI61k1nJuo+rAB0jzYY53kmTvwJQmuv5m/JQ+5WPyG+BGqIy+CRjlprhvNdoOO
eFXB09DSGTvoJJCWI7G/dus/0poEUPI5UVYOQ0vwDq+e5zCfbZ1V7NXp0nsiAi6r
iNaLZh6WPXPn9IXfzby3moAld0/B7l0kfGfVVekTdlAnFTfIkOBInKNVW1mRA85/
dYW64anC/27L5OyxbcCzKxa0ShJiS+pKULlYRPHV7949QcasfU+51V6Ij1olXckq
e08kEjzkafWU1yhbJA49hKdArw6DzgQArk+4H4Ln/LtZwO1j58VVYKzxXDjyW06l
fKdTLHQQIOREuJRbm1f255ILDMPfdAsDXHca3ec+bs69jf4CobTpG48Kdka0o/KZ
/WXy7ghDm1GT+VNUDe+6ow83qsRhlWnWgua+2vZOjpJCJ3QVVuS6HoslyPWmJ1/h
hFBXk4x2xBay9G0bpx7Th/e/Zs7eUzxfH8ExLyF3pROuYMRrvptFH5G3KnRZRC20
ZSW7yHJFD0CbFdvNwh58jehyHsfLqWWkg+wFXHsPnqsv9ONtrTUIbC1FL/yz4+te
taVdgF9L5dz/DtQLUKJ+0aXFN/GwncQAKG1FsRgkPWjscVoKG4n/JZCroVhaomEX
+FQ4qZUVNWZUCS9JfWUeKfmHfjBrnn98AtYrVzkgBuZDeyrTuEORIpBr3wOf4Db+
ZksWBSFheX7Qk8jKB2P6m1zj+MPrIvX7LTanf1Ta8AXrCy8Lh3HGss6Xh5KGfeMN
U9G4E06+S+ktd/nq15FXWuILmjfW9wcJdbzfSHAgYn/F0DhtnkhfY8joZkGotDSG
ZwTtOZGO5b7k/VxNBTkFn0N5scwvIJ18iT6xG3Og7K9X5zp4VD/rWea4WD4ru0Ch
qceoq/xlv3slzyDJhikA1ALPSJjUZO4MbZ3y00tYWvDsamlj2tNdyMlNW0QL0NtZ
l5FB9vy3f5J/6pxGSqS+3ovP+t0zruXAozzTToLlJPsvnVw58IPlRqKt7mJxVLqc
tpym9GVVhqYYPSAQdPCIW+YruP73Kb1qxcN9wuGn3XnkaRnXt0W0jILuo88Bp/Yt
i6YfI+92sfCNQMxJ/l+sy3dAvitRxBDe3An6Xhs8jVJOV9zBN4cmAulyH5AWBNyS
RCpd00uUeI0zmHRxxukikMg2sLF/JdZW7R2mSmOldYCM6MLimmuaFZcPjmqv5FWK
hbucDddkjol6nnQv5RGpFLl2KlJcRzNlT7hTWGvllRBOH7E7FwfYTYXAIZVEZNhN
g8DTfOZhEM2U9teY5csbr+LXvk3a2uqGxZA7lJMOW+8=
`protect END_PROTECTED
