`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GBS7XfT1dGz0KBkZbR9MAnuNcl2hDAhTS1kZdlHKeBmmAc4f5NuiNEbVHAnkQb+a
XGa8UxodI6Azi4YpcQVd6iOqy8+MKWcAUPJ31fedNwp2BkCUo2HE8jBKTwUNF7Zl
nv3EoOuSt217hbGgyaFkbq7AO7cUdc7KudOzAxtdKbfJLkKx8Uwy1YgOz0K7HAwi
QIfVhZZI7Y+8aLxYEOO0lURqYgJbv/5PO0+gWJigQplarhtGIzOe4Y7r6evUGAgt
J6Jpq3QdgkrvDt0oxs3BT/H0CSuy6RyqZkAhiz3grR3pQN0pHiMOstAj0MpkFxsT
YhNfJyfRQmHJ4iWch0c+roE+sgVQ7HwgDXFv27pXyRMYFiLm3PSWSkB6UIwEg0BI
i8YKKXGzFyqw+eg8hJmGOWMqcByP/cAZEknOIDzXjDHe3lmtsEmhJOjiILzjMN8D
5to6QEmrOsYyiAHQ3CZO7joTiGkCPA9M3F5lSyOvmB8cHMqnAh8et17/M1h/D6R6
YKyTd/rx42as5U4vqbjqJp+vL31/Icu+d+RMFY5X/x/Olzeb7dIKusUEmNWb2hq4
ahgnicwX0FoV7wN47sAcU4CDQgKnQl/lhL3roWe1MJ7cYaEan1GAL5SExCvU7kkE
o55caP+5gAS7g6zDuP0Z+2SZ7q6qNJ2B9jrd5Ytolqz6TXC3lqyHPizYNKotTfCr
VW/8J98VLVXcfdPzHp1O0JRaZbrpd40ldAjkGEdKoZNdbmHrRiqgebpmUtb3RyhQ
HTNwuW8DdhlWnJ8/xVh/Pc8auqM+V4xZ7QPnsGjQcn4HOGkjDtRiCjcSZEONGQdx
i3+Qf/jKDUFiwCSo7dw+qytZDRS6AC/aM+qptXvvfqUuQaQEMv34c7NBP79Nek5x
hegKEVDAbTicYLc5JF/R5dmOyDtQGO+ZgKyXAzGRtF25f3X4BKNGk6zEI2Zko4Ql
imFJlACrOEvTF2DjHBRPtRblloQCAbRtRu0jU0cG8HA+PoKRizMrcP02BIC/Sqaw
PsAuFkiXpSvd5FHjf5d+rarCU/d2LeExU1w4vfEkL/ZmxHE7w4avjBq+bKH90YDD
hgUoeY70Jr1gkJsK0MbmX/blBPDF/toCpvJ0uBRkUjj0n790zHsYZraOXHMaCuP0
Z+81Pq+XZ1D+CDFbkugGUQ==
`protect END_PROTECTED
