`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
j0VqA+aF7PYsMFUIaAgXL4uUfLoYnlmAV6hUAjY6D7VlCPpvbruzY8ySivWklfGG
aKaH3n4bmhhVf/de33+GYI7r2lbZua9/t+01FiJeR1fo1Iwt2z/i/1I0hiKIw0jT
sN2Rq3t8ZW9LGDfrEA6Y1g9WHSSiL53LmXJYiY8aFab+A1YFbVjaORJdK+tUXoxC
TKvImqEkPiMrB0P2PzEqtsu84sg1NTvOIGR8MWYHwtWFFGqEiZCXXo5+sCzsbewM
q8dgN8UhuxrH+goSdsvI11fmzuESdVj5t+N7BLJcLI5A8FppvUswtTtF9yJ8bA5F
nPPhoSQV0kdwkwxAttNZY1pBOkqKCsCv5mTqDOEQ+I4ssdtT+kMJddHt9/zncVtK
wOtnpnU4FSym5TnykCC1eanUEhNUPiYrRXwQupg5x9gagegY8Z7o6+E+7rXUiTsm
GgdudifAXcxOiNc4XlAEA3ZSniVh/VEwaileFCoP1h8V2068wrzoOy6vTD7J3rPa
7K6FeREKGXttDwbtBkylwOIKeF4sf5baIWGlWlrQi7CA7LgzfU/gqFof2P72sloE
nvol6putLe2M1WnqowB2Mm5/3MatryTJX25pFiErqWd8Kv5X7rTzwrSkbezE7LuV
c72mUleZ4M9QT6J751eAy2GQG5dyYKN/nSGsBuhX2nomcBFwXl835PoWQmE8HTS0
vo8JfNMrT5SrJMGCUE1OWelrizNoFY7LEP+yJiF2+5IXID92Rnb2PDQ4raK0Z7Nc
ZDQSUfB9UAzsw6VVn6wDKAidLD0uP66hmSGu3FFESiHUDbCc4Wv2aU7+GKuixAHH
rG4bmklpDr67qOQnzuyqpmUoz3tNYTDBPzFnCX6he9wBYOhRizzUhEBSHJtpdfyq
k1AhEHBn7f5syiA3dXvp5znm0DDSeR2Kaan+q58zxr6yKJ/m8Ylk6XfDfj9+hiUl
2vgOOUujybRZkTVNq9LLF32PtY9bWsIwBOy9r4QPCULrxfP77joqKKXjSr7yMe74
DKA5I1FMmealzIdScMWM2QwIK47WgYuH/JdA0W7/Bj0ZRK9qBqqPwslnoOPz+Eau
8OoBR2t6o0PH3sZIR2ubQOr9SMw4/iybZCqUOTwEU1oPfhNpHQSNqOOUKRDASH0t
QTQSMLMJ4uEJD63WsXg80+KqS8uB2nF+9SJZxD4GVbOPyRhB8axXwB741/tfoKMx
qXFZlk7KvvK0gtXOUr0BBOlBLLBgTLTEx0Bj/8PLli8uXUESbo0yXfH8aM8OOYX8
5uBQnR8XAQ5lVhP2oTJIO3KpO2T/uSshgIrvz+img4+yTR5rOmM7jNdraWljqcdM
y8hz6NIj0AV/RR5IR9V//53OfzXEfvn4/F3U/ngy4TmGVfxXF5KG3hfinOtfx6mH
h8xhb/D07I3pftkqSFONuVcn61I8bP//LO/ig6iJrdaRTO2zT10KkfR552fjg7/3
rY5ywRNqWWpry/5TE5Oa7/EO+U2EVrnGioH8eSNPqeHkO7mUBfv91GcTD5nYaSfV
MwZGNd0GjLmsPZLoJoWaU2PNDhPPBhQmP8ASHr7Os9A1MKeVbOp8ZA3tcgr4/nJi
ZeVrYqS7acoBfUxMQ5WPIMyplvfH+CQWc73rtH4xLJOY1AytvnOO0wep0R7r6Caq
UrVnXfloyHdB7xzz339MEFD5eQ/T/pH0zZ/ChOP2Ju7Z4Ns9GRFM45SLZtv3z2YP
3JR7Zq6rDZ7fgOaAXJqtcR7j7keKhNUJlLuYswME2grInvzZKNkGXtodbLASl+B2
mPprODtUGdxMHbp+K75jcPBlAjxkQLQc5WdQ3jv/BuB7xaGk3DUkOa3p0RZ6sdwT
hc2OLL3Ms3nn7DR/Wbso+PGF/B339+1oqUe08WCc1fU4yYDFF/IJhx1vfgVc15TU
P3NyUKXtAn4pxxypnWb2EPQ5sURbXBwM4XICdT0vWcd0+Ibjja31nqsLg/EIGHp7
7XTBzQWT8JUA7RkeP+YeoY+JcQECBzO/uRfSSdBo8E7pg3mBt7JYAMfhVehdNAYv
7km7QT2CESoSDxF+AqU0Hz2dtCL6DvxgdV4Fs9fs6Vr+ZSA+/svTi0bBSKuYZJlI
Y7r0UJwSyLpfqg748zHuDJeyvfqizqU6qR7F5XQJ5mu0tnhzQMrYfRt2Osxp1uqC
z3bxUkHM4Z3anpLaBl/7E4dFGLH2VSCfhgKwTVvlmpSdhooWYYNd2hJHudJIPapS
BYuXzsSwpQEtvwZGsIIxUBXolZ8hnwHs6HFwnS3Cdh95EMsuaKRAfmKl/7xV+cao
4CN1Bp4qqUtO1qoJWI1L4uxIU0W516o3gI2bk+GFZZgPoKNc5MmhM+On1Ft0VY5E
0YkfqFwOAO74wZnaAvjwaCobUv2W5CV2dAnCvLupkLCLBQ78PY0UEQxGy1B0AB/C
jCqqcwv8a6s5sB3gbBenvtbdVRsrEfDeZTL2dAPwKYnnqaNv9JaSYbGvnpIwyOl1
jCKoHvuqt5tO2SdP/i2Bmp85p4Z2XUyyfNK4+gH4JS91Xsrjx3aL2rbpzF/Rqb1J
Bqv5cE0QA8g6oaCcBqkAlr4KQ/87W0LbPpnfJCh9Yx+Sw7t5qe1iId0aHGNy5QB6
cYJfeTidQRLBJ0ETCoL9bjzySLrCzYOi8ZDCgSSysCU=
`protect END_PROTECTED
