`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ve/PtpVds6Y1iBsfT9bOgmEwRv/K/umdofwKiQYPeKVjmdVyP1dHDJmdu+MslEwS
U6QJlJ/lSp75KDipLQh4W4r1MmI91EyCiQsKPio5h/7n0J0TuF6anJUItDwXFMhA
2LS1jmjPznvFRbrzHCiLhLezFs6jiVHFw+fl3FadF/OhLtwNAr8Le3usvxW1pgJU
Rfnp9cjEv4slNh6E4spEkL8so3Pq83PjyvoqKrLYOZCepcSuH8bRjMRJBbSlGEfv
kCQ0EqhOEomO1IOhm89zmYGITrBwUq7jY1AUj2dHHgCc72El5Kbf0JZ+MPblj8Oa
fSR5v1i1IsaR+c/dg8gDH7KKRB6qzYJm0BQD3NdSlP8LT5Cj4ZXevv4ve8H9HIU3
Z9HyuAKhiE24PfVz8vpz2jO+jIJwxaMokNF+dqEA/OrDRaqLWUQgpPdSzwJ+EBiL
UdW7erIbQIBInUrBtNntRR8YikblWrU1O3AOsd2KDIaEyah9lHdQWf8yBBxF+xGW
Nlz+KWkkbbehkv4TI8E9umdCN9NqCq8w1L09Ih9vxWZLjGlB5FZdI92XJTMBNt6V
BpDYLSLWLIRPeNtVi7s8Umbu1h3kq9YxWjBjVG7yQNrG9vaznpTsYIpme1val2BO
QBdTO87c6KBtbf+pTH2FDcPWXcIZvFCe9mb6OBUNF5u9Ke/O4dqe6qCxRiSR5Lbp
TcnhF+g5vCFnJS01kqd4J9FODKXhcb6Z8wH4+yWKJnA=
`protect END_PROTECTED
