`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7gK7FFLKoQDSi83/xtasxykTqWwSsA8owzKKsomUUtiBq16H3CwvK2/Kz1WBdLSE
Sm9Z2NT83G6BFFVOEa+YFPmZQgLx3fDqY/kf7N4KCsdZOFdBFUxoLFptC5X41wsf
7rdV8vwKTjbvGddvqvx/RtN1q/epOSFj2zVPpPJufp2Lb1swovs7xjB2V6TcUzru
h/5htovJuRY8rkjR9uhoY1e15j3W7nl4Lg2V2BC4Ubhd/fcv5T5k0rrCzsi9yAq7
x5P9df/9L5vsBJLBwm5LCwxHb+xvPubPQGo/+Z76Bg6/iI1z84i2ftJ57Q0+lC5/
nEfcatSu4EruVPghbYZ6ytwFLUqB0oTdbQUMUKg2+FOArdVSZSWbVwPBg6gYrxH7
9FND1hEnA7sTjXzvSb0SIR5tI9xQlOQtg+uZrWCaueP4aixUh39oAplMpX8SBn4q
zYaR77Sm34b66QLijG7MiHsqkSVoIEOnXRY53uhop3r1RtrQ9e85/q6oAo2eMCRZ
+UGr9tUyZoI34CHTTc/FlHLACxF3L6dR+3I6zgzrXCatISOq8kKHO7Ss+VkEY//n
Ls7Fq/4iyQstmn/Wmug4S5UXeuxiE0JwfXfeQw6zJjBV/1bUv7tNQGVgk6iPDtSX
5wVcA2jQh1ZEarbjADikxjMIc/qMuscM6JNm5LUfNTwG971IPoWMN+6vTQwYWpnj
cByRlXnJ5b/hSmsfc5Tqin4UHxGgiXs7wW0yrj7rR8QgMWKmW2vCBb7O3hV83yXk
8I6vZCssMDtqVl0rIQKQ9ZBTs2EtXzA3gWfCN/7+wQY6MRgiYRn6s29YSpj7Xov2
k7lCk5wLTREz2R7JlywlQ2HdSroEvxGyEtDi7vn0gVLRPFeUWvTPyipvKluWKDYv
kec+4NKP8VeYaNK+MjBxg/Obb+o3CkXlIPfMidwrDcHxZj/Rqz33SOUyPKUSsbi+
4HcsoUFZftlpd4EKX8V17H33YDuA842hsXsLfr9ozngHchn2WcPLvc7eElytEEYW
QWe1FhunfzoMJ4ZamrEWbA6uSSn7Rc1GF9In3z9BG37U9ViAf9dUB5ubQI3MxWMJ
d5TZonHuO0gC8LZ29VN4/WBwCdOTU1zcJaQUSU013+uIYZd67MQDe6Wye/tKOSVs
I8DgpJWQ8Pc8aZ0E9VKdpxALgUjSsNFcWdKQbKV+YkKxNq8sZMpNu3/FZ301VNGz
nK7eeY2b1h2lejxBgp4JcbeJpcpzp2wy5TkK92sJ0cw6AjAtqUaFTXyHRoIxts1b
2WoB57NzGSmCKSPxZa5rTJmTQThoWRNZdpmXnoZhF5EGbMj/P4SONqE0kkAOUb+n
IXNj8HblM/RKQx5S1ctsUFGvHYfNNEu98ZOm2H2NK+YhH3jA2+3PT4UIdsz5Szw+
IGiyLMIi+XpC9nGyjq5ebuKuyspnUGNCxB2rRj+PzDHu/+eQab6tfQo1Ncq0UvyG
f+shY93WB8xgG4mOuz0XdMOY6bb9PqFAgZ8zF5ZdhAw6jEl6dbr3D3Wu94aReLtn
pNlDC6wpMc4Hk3rHJRGF0foVDVx+LnqcBJ0Gpf7obYVdAJMoX6y8RDer6Bx315Rs
TfJ2/rre1QPd5/KR0Ul5+7HHjrnJNINB2pj/plGBwviH3eBTymw3SlkNtSOIdYjc
bXoXlPTr1x1d6uKmhDOhIyzSV4IXKpO8wODWF8OaEhhPAsjT+6C0WR6gcQKnyOk+
bpydCXXldhtJX8JopUNTXgvJFtYmvV0D133UmLrmEP8hvIJmEaFHxlPp9G9BQGRI
9Q4P1QkNNJVFl68e7HuMQUvtx+3zvxPCPn+cNH1lESu9RTRNClE1gQxBgJ2e4Sh4
tcIPqEj2hDgQRLUJICThxJLk7Z4ifcmPl3w7aAGPUdobT6EJxoHaoVnHOvCzi+Ty
s0OHTiy9pB2vKh3k82EeDaPmf27SVy078NnJNbJqllBsLgsapeBPKHS3ox1Z6pGV
w0VaUFzfUp/XKPZs7v5u8xTodexz5v9qiE3yqw7qqOhlLW/gaK+5EWf87RaSwYd5
a/zeR6NddYxmta+aQITI0/LniA26NYUJYZSdZOyU1RtzwVV53P0ish2Gejt7myxQ
HMJ3GJXqKLJ+IQeImyVZD0lykuFPtV7QDYf02jZQnBcUES4iVvR8KIuc+gSmKgT4
deyhbx7hZfdYYqFtWoQVGPOEcSCu8tZmSQxWX8+QG4w=
`protect END_PROTECTED
