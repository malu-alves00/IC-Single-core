`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ml7BmaMeJauOKFE/khkAmMAw/8UjCMMslGbPyaxLWR3kwkVKtEKf1H/L+SrLj3Fw
g588vF/DotDF5ewvcAgMVTxRCOib/3YcH6jBhyh2VFql+N7CiaJI2DlRX+2I7XuJ
v/3GBiJI5KZrnFHOvbOOPT9mj7XpeL243Z/zFzR8/yCzuhiu/T9KbuFqeaDy8Wdg
00Gjo3sGI0+U9vdGnBzDTE2vnDqNoMATuVPDrmJgrDYf0GYul0AhhjlUvsN6Fxe6
mES77CHLhm3hCTc3YcOSy265gN7bwAKOO7F23NNIoVjIRN2lX60Vr0tlActoDxQw
jKrpHArEQ27djQ5GP8b5UR/5Rchq7cs0LDghEBKKt7n/UT3ksZzkKuODYn3F8edH
G85637/7xVjwV3KN19xzw9XKe1PanYJHzZYuk0yBByL/ik66mtO0TBuK0Scg75MA
CNh3u/qZY54VE6cFDy5Q+T7yN4r6kVJKWjtggKUMlCcQoHwSRqRvux9H+vExibg3
ydwT/PGbHQdAWpm41YHDyaLHbjZuUkgftTOv4Y/XZ0LHXq/tWlJT3aVDgBEax+jP
8ZQPFlpxE4AbYrVUIEVk/MuF9UBh74nGchvaJ0bIRUB8c8PFJJ92WEsmh/rOrJeW
CIbO4LmOSpQIlhGgw8djfdOH2BD3mnYswIArn7xd0Gs8nDhTSKbNVDIAGN/ziDvv
m9IzarlhFLpv6a8lTBeJ+tz4Clhu0Oyd5rBGoVRxuRY/hcR+jyt6Uqlff2dHN65T
dw2N36+Bsm128Dr3gKlBi1+Sk69BN9ssG8SEISfowCZIWVIOChkWwOvI099/pGwt
3LIQ1GtaRWtLHu+k0jpPrIqD6xhiDZ3TDO1EmoDhmZtUagFFmUDsxRGLO1JjALgp
oyBz7nK77q2iXcWlUMIatKtGWG4VyPHqOCE7Q5VW5uLVL3+jJ2+eUZJFwrzEudK3
zPAQKqc4eFvrmVJu0ncUe5XqCks5KXRYXDsTVCf/y6FHOagVxd64v7fD0ZQM4Jr7
K8F5efnRSTl1xVBJtxOmjTLiLz9pdcvtw99A3dfPRRuEPICjyBJn788bRSvyV4jQ
6zKdFQsUHnSbc7qTOLU5y3XZ5H0LnrM3+GaGmWLl/vd2aiClzTz4axXHL1hDJSR4
rhQi+3UAmAds7ypu4Wn/y2KQlGtxxKb97tHMACyYjpIjBGRbtOd90BDcmf3SFh0I
r3UaLEWLmNWJm5stxtAB+8JVUNoV4hxwxmP0ziPbwweo2V/QPDPwG98P2SEoCkpL
9m3zN+KYmwloQhP5CnRY7pNE6MZmCoNEqaRNrPUCKBNLWFa9yW+nBHL+AiPm509q
Dmn8qXvx2E0ms8tzVZjtDY5Ay/ZveHdrf1jtlnpJJ5xKmt8vxRLRno4gbWeBkpP9
qq7rpsjkpXVYq6kr5BT8RJTT6AxKaXHZxesqvzF4vfew9jFpAhLLoVujryle+EsW
`protect END_PROTECTED
