`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NRq3aHQTJ+Y6c/57Rv1jn71dzf+bqHCKIJKqTGaw9rrddBrsnpf/pgOg8GFOQ+LM
FGInWDsWrWMoNAN5xaGhgKglx6GKNxdznArN3YZJCcc9m5V2gfJAQ5KH008Nvd0j
RKBFOyYYG92H9GhXKk9F1JysY1uqQJ8mE+T4zn4U1YGv9mC9HHPDc7Kk1595eh92
q3m30gB3HXJM51aF6ue+tlE5tL0Z2QAwF5uWbUK+7DblClGaNGbga9ATYhd/X15z
zpchx8eBJfn0qlg+wJmgyJp43EOun4smU3dJx3X2npo0LJ5ZL847huEdPLHZnMP/
0B+JuabI5Gl9RGDHM8ejk+cxFU5ga0PfTp8r3oWoLMDHxSTyqdjqC8tdYMoDz8wT
yZUZtMfC6vMyCWuBfYfkdOXkELBcToROtKf7ew7ljNkq/6XAv2LnVDq1KXYNes6b
BEjCjv5l8LFgFLIJeboVbxmYolJ+L4aBNR5MeKiRkXorYcZ8hDlxJ8MT+h+wfw4m
X2I0vFWCW8w0UJ4hI88iAArQwUYBnqi58wynGSPSAtpO3qZR6Jao2aYqyWo+XVrf
E5T2zEUsUsrnq6guQOY+QYv3h8xy6SgrRoiLDLjqCU/nm9Bd3B4ZRdQiG4rL7olt
m7yRuf5x3jNPqJeFPmsG5VRaJU+SYyVhOTLIGRl57UPg120LbPs7umbAofoseFy4
xWIDfvwk5AuhKZWHsmOyG+yzSZTiIkXWZ975iUzq6VSU3cVxhBPRBICDBSVBBgyg
NAzZfyCOfW+deWCw+X9lSDx5HzyCG5YV3EfotRnFFCMZGTO8XqJedz45Zwqd7CDr
z1LumbjzzkA6PDLR9DQ8lXfvV+/bFGEY/0O0hgeQWRgjv2ltdHf1U5vQ/OvETl4y
Bz6/rLD5QzU/eBCRBNLaZyGXmeyHCNHlh1AyNg2ezO99AelHUUreF7TKDDBxJ/0K
praELRnIr0U3nv9mnBJq/x4N9F/PsQlv4Nj7RRo4hwA558y26mdulghfoelU0ErF
Q+D89PLiij/AfCudP1fiAg==
`protect END_PROTECTED
