`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qCeJPqcYsyfwAFxyU1vg9hVIky0DGJBRpB5LlfdkW91+U9R0MN8rXyEm22e1/Q1h
RJZlqT/BM/P/yZqqXoJd3xdRMfaD8l4i7qOFMOvjlhgsla4qFZkzcg9U7DWcWCSy
jUWsGeHz3eX7SpMowtP7Gtykjp87GVfo6NBAq0KuMIgnqtdODbfhEhk1sM+UQOCo
yqrUHMWazt5YBcKZL/qsAnt5izk4IOLRRucFflfdYpqQY3gHFrGhf9+vUksQepst
SHKAxcJT8HblLOdNqVOH5WhapNJj0RgfMvR+aXTBxpGpNhKqsXZBIDjsVZ9MOf40
r1xv0RL/8vh6StzJ2XMRbj/ZD9l6JAxBdPngp00kjdNPMe4a3dS2sYt+0NghGeBE
LAy0sKV7Qkn+4KJSWvC1MNNI6z/ZkpT8IdaG3D2h5EBZmKL/YgnfAp2o1q/JFoZr
QXYIN4uP36XTNKopI8vnRIaR9sd79VixBXt/SzAsflnh7RQ/NLx/VZma0NQ7mCOk
ZQUQDCpAMTU/G1+AVhStu1PZS/GZzFy7EE6WMC/LQyRvzUHJEpEufF8Ad2LtH4JU
Y4f535YlR5vNDGDGPEcMjUYGzT7tUJtmFuobZL7xl9ZZrkHatOhYsB1cRQ8he+FB
TDcEurRdel9T842qPUxSlxSYkgotQUL9Xirp887Tx+WB5A/6JlOQ6NmJ1ZsuvZyi
xHzcGTbT5gPAfn9k3VpcdEXOwmyMthodE9/GYtOR7lO+K31cqa7iMa1X2FcqZRuB
R3Eweg50p/3MmeZD28Ks0e88B4FOWXyqQkeqDqVFpGnS+/n7+HsoKILdqJdzlgLG
lie34gS0Id4GxcuGZ3F73Ab4SiWxcRbWrwKyTnToTZzyMdccrAGmGX9ijBsrE4As
dZ40YHq67KgAO03e6wsydHm+pbnKO3m+tuUBmdVKKcEIt3ClvgIGJ7qNhzYPrLLl
icS6N97lS6G87ccd0qFXpGhQbA49TOVD4yjhP41LdSseZ7z435fF31EsUqaivpVe
YsGqJvmhGlpKxv81+Knnpqf1/6hnjeQcyZjMEiphhWTlmvszAkmwAnUlrvemixM0
XDV9o1/QV9Rn9IAvCeNsqs3ALUEKiEWi23BPrCdZd325epcQJksHi5gVefTJGUFs
sTkwS4qeyU2j/Q7Kn7Yk50mYllvkdPUQUUN2e6JJQb5PtY68jLuzlgj7Pn70gjUc
REruMjzRi6UmaiZBnvoYM14fyu9X8ap1BAFQcrg/OgrjsFNmxEbiyNxH8bklfhO1
qitskt5ry9uNRgi/rae4EFEXcJEoCxSdpVb1vHzKFIRhewWDaaXDUUIUSzGLmBKg
FFiub6QnJQLEJfs/fWd3tp7vhrQyr7UpOqtF0rMBI1ZEv5rBZfu7kliP1pVNuBMb
LG4hgwtngDq9FuSQ6yZrqZKC3U7ZIAbIlhcxClX8bfdy7nw/wo4nFHy+9amdNdni
`protect END_PROTECTED
