`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NV1weJr91caxF/hhJ6R2aoxxm1rsxQyY2v5KF5Lk6n6gQGMb/BqD25YaVpKyGb1m
rr+s8tYFD2YKSKNWERsRljvipOQwMOK3BSsAKuVzcB47zhWXU8xk9zPSSWN2dGo3
yuzZ1+Hu/Hr3qvcXkNzRasfJHCdZw58ZVrsTVuniydpH/MqNINEjgtj5bzDI7R4+
nVt13BOKbQsJuy1on6vZFGrejGlBofHl2ZSVSqJO0V+a3atFGA6vSVbK52VoM0OP
xolgRQYCxJAmt0ADPqCc0AGtEq7lQw2/ubkGKSOO/PYlrNiLALFaqKLVfQNASOum
9f033B3IJ05KnaAftLN5L84hy9wxZywbSikiZQPKaVjM/luv9iulW6NqVlXjp3ks
/sZeXMksYGm+z+vcCqj0+42YEcqnOBIkaUMf2v58o85RjJIlzFocfewWB2wVf68C
YA4PQmo5CVx4Fwh9g1XiOj8FRQdq9Jd7oCjPx41oZxFHy84pkQFxoTevTWo/fGZO
hPf3pyQhT6X+pRtQlWMqNkjBWQGLwVpCQUKc1DygPR7xhxIoOXAHNHQys5J5W2DL
0PJSjGD1yRghehc03M/Zr/qInsBHipEb4tNK3l8OIby40fkVvy5xbkaORejiPw4E
cM+40QrBZ5vhvQsTR25KivPaIv0/OeRTOZSD/3sgn4kQ62RJI0IZbuaFSJC2H7lt
n9eGkZrhappzTwBZphHO7FJcbx6HRspb4WO2u/JYuK14Wm05KPeHcVKqTDvEdKnl
ELGgUJy85KHKZVkIb9o1vH2T/aF/+F0avUHjZyd+M0l58QbCETCyW0sIoqh7OKAC
MdTxP13rkvl7c8hDj78Q7nXXif1G5eOWP7MmZylz641PZhUNAv6mCxFSU89Cqc/E
pvsqgHMsoBh8fhN6QWNaXuRbWiET7A+VSMAH3u5aaofJbwhHkZUv3aqDrFq+ZVsf
5zmdfvn060io8Fqd5UyxdDbVnFquCkw1D8rQ7ATFPWocc3ZNkriT/N7scTsT6gH4
z8i/S/J6lHGHjhxW5w0lZm447I04gbXc31W9b0niu80xPoXBnzwxRcV11aj8BOKk
sZsiu55dBaYZ2M/kudYjJcFDehb9Bt6UoOLTQt7LrfkIhOc/LtlxXcO7qx7Ek+Zn
L5mXNc1+zHxElKy9I0gQ+yF8jOc3cu79Eb7D4AjD0Ahm1FNSA/8cM+OeBqQyHYUR
SJlkPqZ848iSAxLTqygpckW83hms9jJa2LKKlZB3s8iRFxQ4HWJwafDGhxNeyZSF
lwlBqZg1LTHU+Z6q6yE3wKy+tSSv8Wr4IL3oKzhE7FEpOoZYCOxqyYyHMxvQITB0
o5XTwPPx+ESs65wzD2gUWXAQQDiI2ggJEJC8zG63+j219vxJtnjSkrD0/J90P372
lpuqcOo8UEhJAZp5dU0T3UMdlQRlMhC1iFf5C5mi/5wUcEye8a0t6xXVI8iQXLvI
lIs2aw3WGvASFq/ziVBPcQq7GXXGoxNLKHLlUcYQKrfX9NKePutgTyijSIC4KaaY
udZ5KG2jNt+hmOqBl4clMKOxpmbswE7/ixRj+4AFUjA7hEQfoq+rEqM1E3BRuDnu
UNsshMXcw3B+LjmhF9xCIfk0zReNjKgWDSBUZGkf1oddqXcE3T+7yvJxoDeBUxBz
pn0o53jndRDdonE68K969tamjvVPpL/E4xt+TkzVdFeLVt6ycc6zAS4T0/jgAMxA
0dRcWvHjhDG/U2L4Y55ZmSnAb4XVSczfVl24eHdAVBL4/HiASFADqLeagLxb2F0z
/u+vVieu9UVl/j+6VwZ+WB19A04FXwU1N4XVUjh2qP/hck/3QnREjoG1G3mC57hR
kPBDWUCoKD4+NkjlTqfQGrh0s3L8+Y31ptSXbttlSSykhfQrve7z0/XMhYRMVGWi
AfArbLk8ORSmPC7SPdgITr4uAAYuhH9Ef+cddVrqa47N96LGW+rudqslLgbQepIo
WzNU+gqLUxHIZRBOwVPBkqVDxDyChxLmu9sACAEyFZ0yg16WInqcUok9Yeoh27wH
eyI8mTcWBxcJkIrXHXc09Zbex2D4Xwf/WXetO9ljywYBGyxIAdImuwdFVCZdUSA/
qGa07171Ar5VIUol0pRpI0jIRfeNpPsJHSabf1IXc/1QXWVZrEFIaAmC3GzONfnv
SHdOZW5KM+SJ6XcPg/pLntve7fq7MFsL9Ta4UUGlZBktcpbrTB5lYjvKYglBV5XS
IkJhcoNhM+IzYieT+0HtGXr/Aq9sypynsSvQ6GYuv+Bp+tHsruIU/MNsNX3/v7b9
E65yO849k695CsKrYEIQZKel/6zd17GQ6Jo9lsT3V9HYmTerpAPMFINHhb+y8/pH
ItMUZJb8iA02t4XVao9QGS0A2ogyiRKm1Cnjr9PCrmI0zHXL2ZEna5DoBw4kdJhQ
SL9CVzGp8is5XeBWcgiOyAR5fVCOc+oG8r3h+u8/7cVRAQqshiwJ9qhes59VjHT3
bVrMq3ZCNimsc/GausMb3V46nZsFxUiktp1hgtIB30I+2g4ZZxbUOS+y8gsA0QWy
YJ5THhc9UKRhjbjzwLr8dfDmZYUdiQ7OY58G4U4Re4yCGbeqbS0jLDLt+5vi8oX6
az/8b6rkUtOROH1jPqKIxYyksjGx3b9A/J6zMtd4fbxqZF54pO+B/gfzoRw42I/j
JP12vY1299r7euzksSR/Ubq+IetTVxmhiwzr3SvF7q+qUCKnbNQtkwjlf7OdjwhT
fNy49WMMsTzljUYfV7vEliakxaA4tO+jT6VmoFCOOrai0T3XSU4+Eo97pR1fSKae
gHxU4B9p8Iq+tn6r1Ssmz3QI2ScUEiIhgD4HZg+QpEj+QccAGb6G3wPt5x6dqnfL
QPTCQonZHl3D+/U1BWzCm/c+u4GcfhWQjAEH1gfe30WV48kcA1iS5UGjPxb5pDgz
IxhxegBigZupbDCp87iAHNjfpzHDhrRK5Jkqnci6i2y03lic4PyC2Jvd01uvgVSh
LdRL6ZySA0JpB/3gjGkBQndJ8Fx7h3O5evYhhM20z0X5pl/gQzvbFJme1m9zLfmB
UoaStFPdtAHu6MjWnuNNgdWyzd+bXh5frFkC4nT72YOVFNCMv6A7ug23wB3HGyF6
cBPfAd087ceU769l8w0L6gRGqK7gqoJJT5OWDdr9xe7yNgdyzKBkFGi91e0tLWQ/
2j+BDYotcWX5SIDfbE8iBHAJqUtQA8XOWJV7prhNA9B7x7goiUzkS0rLYl6XzPid
aCScF9ZFwJIb2zRJtZrZvwtXeW1YZIgZWXx2rrs2hhgJ7PKr9mkfvmT3At3uB8+E
oSIj9RGtasDBhJ/q10GjjuIm99o0FK86trRbc7U1dw9M1fRUQLBgol5gHeSiIG8m
mUBWFANOpmyrr5J2ks0nLH8VwQeqm6PVNiqUipvS4sLMB/x8kSAk4dWV5H5c9oF7
CJB80zAVM1sYeKeGa1bB9qdaBNrds2XQTX/IUN2W/h3aoSR+QfjDntzbu8aT3zGp
1HVtAYBQ0IpAvgcMt831gnqNhC/BQKRMPe27jBL5kqlwIkhSZjP+eYG9z0CH7/Qd
pDgB50UAZXISmaNZuNW40AWr1NwBARBPjtGkfcnHtULoIyyHYJeYvKVvOlOQnyng
/0nEkuX7SCuOnGCi9/nfo1LGqFAvQGfpasW8yd6zAICO9Xk6KRsNJeVp/lsXysf2
N7LaS0vgVjnUQZf42nz8OF8HnS5DMPp3ID4tLfNWxscam4XyWYK0Ive8stTLsWRd
Ui2RIlzLMnSeOUfmdoZ5zh4cAvn1qZ2r8nnIpF/uarqrt+OciYKNqp7VZKOMVfCB
o80cFFek1Hws0tijTR2fUFYZRIjz2CjNyCOQBt8SkRCJS6Y274aFWIb4S+mRTWlL
8My5u+YLa7Ta91ZtjtsMEX4hP2XiikOJbZxOQQSFgG5BcI9V4FD+BXc/vtd0hQ8C
DF8XCn2aBazwDSfGwWACIbFXpTkQ7ao5ItVTKln+a/oURGqDVvdgK5evJo0qJb5C
TPfv+4eGiZB2KOUY1/qZsZlVJwx1I+C7YydELrnFFpvwDuh/czTrXdUmJZxy/rkO
kj1m2LZc3FlDx8pekWqIRivOG3DNW/vhA93juyoZmd+kYyawwdT56W+uvCr+YyS7
a1iUDSPcbMn/sXTjii8zUsoD2Hmn4aGVSt6/jroyG8zY3xQsjkInLJXhdLy+mLvd
ORh6gvUBrqd987Bll/whqCQjU4eGvCRCU/Gvnu2OX75IhqDZBSjrCiITvXqFJfMk
GKw/rq9Ez1HcMNnxlxgJ50HZGmq52Id2np/jraZwRVcYOdrQd3W1LTWoV3CXWEP/
bqEsPWstd15N6qUPUHZpmnnEu9yfS+qU5UNzLeyXL2FTBNixh+RHC4E7/gwwfLgb
roef6ziAHRV39/nH9yPvwqqH80RFz4bupMwo9dRRToGlhi6R+BfPLPWqpwoj7Dqy
7VwrHdtowBBieBgYlPqTvQMLPe9RfDoI8TpXml3oLwmiZmHmZtHn4CJTM8AtZ34b
HJF8qa+Y293jfoBijJihNuHee/QQ5/yGYhkzk+eCItPQmohjS/hxlBnqHdyAQRVj
cWYcUU8ivdtYa6U1To4kTI36JIifejtQK8rVDI9MVzAJ9IMSraWcknBCnx+6xcf8
jxZ52X7wkfUPwuZb/Nx4yA0WXNL0G7ld2LGPdjFbV3XntSGp3YfP2beJ9Suzvx9w
ZVZwQquQYfL5cGC+llCqxaYBBeFnwqnshCLqdMXcRxjksamoNKcMrTQKWiOvG/sN
3o0opF5JBfLpdk70pS5rSN7JVJ98YHva92476Fi1WQu68jv3tdjoxNh29lTZRhQg
J/Jqaoq1i+K3o0yVkICkTEaBHrFwN2FoPVYqJIgCgjXpqyGnzUP16ldxsINi6fvZ
`protect END_PROTECTED
