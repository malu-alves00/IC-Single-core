`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bPyReAKti2FuEMIt1hkVkNaJN/OSZ+LfihYIjQdTQBoCT7vx2mH2LzT5bD6+ifpI
yJxDXyf/AvS3qXyQmFbLBtPqgY7HQDlr9i/0kqEOBKPUgVDM7rdfgOeNSYSkYMbE
3WXyfulrKy5tsYs29PLwsmhF0TY7+goTPtDnUdAtgjmTcMrJjfc4bJsn9MQxmM/O
FTXg3ZlzzHNzq+/IZWk8miHWmWPPGG1NlD9MhdHnJ97lt3139HleT+cgfsK99TbI
kJb/D7vZ2G/n9h0uXJrU3D7zZMGy45WTLlASW5D5WswRgu3yweTfF2QVtD6zY1pk
yqPmyKS/dkB6Z/B5VacpM0N+drh9WDw9H4i5uGID31urAsGttc+NXJgnF0qj9cYs
Kf8S1eHheJp8aZFZRAaZWFx2xQR6TcyqiTrynDhro2qErseHdul+DwNS70m2McE8
xqdh986mWwJs3+NeCKkaxIecMd8L7RyvRGE+jetmJhc=
`protect END_PROTECTED
