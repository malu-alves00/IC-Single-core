`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8OrOejKElbmjwIHFGmnGbhSolGtr5v3xAVy0wKtVri1uykb46t+cSFNMcutp3aWi
TksVoDgPL/DsSDyJPm+9mLIkbDDdEYtty6UZBrfWHavkv1O71G4+XklHxAPJrfa4
Eiy1p6BEAXFjzA1YK01A+tclgEWnLf4B03HCZE6w291wl/3BAvDQXQkX0ffzfBGX
f7CItopImqBeb9BKy2uYr0UP1EzlVQCcquczdYeYJSHLmHYDxxpIBdkkMQnGWkjL
jLfoI9cvTseO4O5K2qjBZTkmHVdnPazUQ2+3k4mVmtef+9LBbf/zIuK7kk5dayN/
P8GfIq7hN/0tzYAIABZmnePRAONzCxCNaW8m1TVAj9Pjs1/KdfTV6pwtwHvbJ2gE
hH2lsDTO8NHwsQtnwTcWIPi1Rt9fB+3BR0TcfhdY+kzdoc5UPliP4VLFGvaHzGd1
MBASyRhRLhGPdkgfhhuwN17hYnQJSFn0cqHe39RmbXNUBfT7iqFX13tB9luTs1sv
bEPCjEOFuW+1Tfn1JwSd3XSX+Fn2lcl6PP0BQXFR6jy5XFogkg8d51vkv6b5j60H
Tf/lImC0aYvSVSUFQ2j/JzWCmamwz8mV1sBKcMsJEXk6hHR/Omh+yUo8ViEEVlPH
IGNe5kcVKeZss5QTWkGpEA==
`protect END_PROTECTED
