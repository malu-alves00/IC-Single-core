`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NaCnUZuu8G+XiuNIfKFhMVOPdaBbNAzVvUmuOgQDjgueqFRw8voZ6PCCMHZgsIBq
7GOvGmkwb4f7SHVG7L8YAA3CadXMx0unzNUWSksAPZEaxJ7FpsgSWvkx3Bwj5HPY
wquADzZ90f2k0F4P9B4xHUqh6abVnaemepWkdxKL0IO47hEzQo6geDUpw44GJLp6
5yAdoCWfpWG/QEEPWPybrZWfxqTbsvzmkhpASfYLoMHKEXi0XABQ7NlEWJozFe2v
L0ingTO+EHeWi1vCLCvPL48JQe+7b4xMPU2g7Wpw0nf7r4Yc27h4it5/LwZUKuxk
iPQm13mjBd/p2lZSm8QM4N/ZAzeCGV0U37kKBDx4bn0gQxni8J/a6T6hNGaU1UHi
sB2XUNOv+EoNZxL5w9fYQ203Rali/WuIbhU28SMHbH57dcgqDR42DH1dkdTHBa46
kV4vbk5ZCYwrWnOsE7c7ZPyeck44NXyy3dA21qppLGghUlrVGIzvfM6OVfHEtOIs
zCVM1u6AVNzrHtgRv9+hGfVbbJQjWwVoANFA32iT40idogJThFRcCXTGvN29re3U
QmWM1ZyEXhmF3s2Nha48UNyiaupcyqzRmlDWhmhAiuhAPSSJUsAZIyT8HhDYii7H
X/tqF/swh3CVK1WLx/94cTX/POuuKHiE5Xoqrkb6q8uVg1nuWaEdbmv0QTHX+mtm
H5YNj7kH3TCaT1ZTj9UJwGbRCgS1n7sjPdGLvrRhprq2nqnAL/SC0cRxM2tMTCxv
70HBe0NacR8aaUfWhlVfWYYr/8G5WFGXgEIv8CVRxJz2mwUI1otPxy2Y3fHlNTH0
AlPmpDX2k8oUlcz4PJO2WDg2KA70Hxs+vJusAWGSY6VhYan1WzhlCjotF6GDWFKy
mBtRX0eYQtP0T99O59+bkT77/+Tnd/+pwDtc2bYS407sgjgEj1vezyeXgSSfTz5t
lEcIAc5t7bR/rfY3CRzlBkFdIsdKAydLj3zHkcA3mGE2ajA7+Uo5ExJBv9kYkfJH
z6f+07j1JRSxzty3hQGqLlh1NoBN0nqC2/+BdafdCctyp3xREPoVmMfa1vNLR/Oi
0RO8/OBwqmn/xJ/jMkUcVdRMAdspCReY8Dt40Sx33yshcZJIc9Qnhb2H2Ntq/P9b
xJ9gR7Qczy8zdbRp877cyH5VeU12tL+YSuR92oXvwDFyyHhPvuJKICZOhntV/lKx
KLyY1WmD/MdzlfXA36Iy7IEFs5aB7h47qJXwpDjsfDgPe5wqveA48mp/0neBywXa
JQJWav2qy0KWUxsofHdejtPeB4yhMKWDSW5jvw2CuKtL3nunmDa4h2ZVCPSXvp3c
HU9w+PmboGQPYtRDw/aN3XnJWRLnEyGBP6fIOpN7WzzmXDHlcN34eimHnvf3CWDC
UmO9I9aUeZaA0juRhQktaOD7kPKFT+Ir1C/FWXIoIGrcHOpYEkiLqLS45RdUIFHV
H8n0tsEYTXcaydZgDPp9FMbCq/ds/bi1yFV6Lniesb3kP+UkwQw/jUa9lxwIhmlR
r4KBAkDhP1ccbrawrIlWfaseK+gJX4TJHZbeqInsJHd2HK9sb6IqN1kVPnU2sNGI
1qyv7LyX+p6XvP0XfpMW0VCOHfNJ0CmkmnM6t8d9lXf8ZNtj5Kyr3DrPxUEWTPka
aDvKSXNeHpVXARJq5jph2nfa7L7YUI0Xpauraqj6evlMQ0S9iNyNxbjUbXRC0dhk
gpzEZt0zuxNivMRBmCV8cDzRYhutP5AvdUdhBt81rQ6NlE/L6YQeUo6T23hvnRsY
BKRKrCn8cuCh8rxZGSZDfsnChfd1vB/vb7ZykLmmIxC5Y7g19Alm+MIGSiDcsqG+
`protect END_PROTECTED
