`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rGSXLsu2xal2SGE0/pMm2EY9TMc9hX0QHriAknmAxCsi8uPQK1EEVdAoCzu11qZZ
74EyaV52UAgwsd/y0mL6O4hYPFj4WXnTTnhIEvfrl+cITZZ6T0cliEjvMAw/NYqc
O+hEGteOabyYbdNAImvu1x/pKKbRtoCzXLpLdCifma+sd6YlahGc+oWUkgkt/2lQ
snWqG30KjsgBeyvZUO+KcDPNTvFY1USFbliwxI19fOKGTiIz1gjJfJZAYyACwHkn
TaG9kUq3KkfrV/FVJ6I0xBSrBefG2/3umj8893re9Eais6WGcdxu+x4OhTW6ULMl
pGmyL7WbgQfFHTaJQnSv7qAzpEg+p2ZhIRM1bO9AJekFiOB8hE2JfbEev65lzQCR
ozM9VbY9ESH9kZE8tTNiWn5yVlfN8NAcn88gbns+T4S+VOV/QoBUlR3sVnq4M+Ul
XvCKMH9gu39ofqgBDKmIqtpWFimbU95PRm6NegpCX2oJOXf58oXDkTI9ycHxjQ3b
t/KuTJrhKSo+CVZg8/svUSXs6qreyrXHFcQCXN3FTp50Z0Qou3JIEm6zgNB71NFf
HQXmSiAPNNA+WRfOOvpX4OmkIE3XxbexAJTbx8LIGVVaNX7VpqMyl5Q2yOqdDeo7
1o9ayVNCKTNtUAIkf+R7bwdzU2oCgW75oFkETfwCroO+ItP5f0mCycpFO5U9IW+t
8Id5OH4a8TI0DDE1Zu9yhcY9xy064YwJkeS2WSoJqrzUml9ImiSuBQM+CHSMmn9y
mujaLTisJGGdiLtBEJmWm7q8grV9+EcJtoB2IkPkQu/4drb3T71+vdvOwd8fnN4w
CSkp6bBET/9+tDyTbbrLX7bFr+ngaV8OS8EtXLiPvLB0olzJioS0rZf0NBoHd7CU
3zjq2+CbdrI7o3Kk4HKnpOAO9lrzghewmkdQSGJ/ExA=
`protect END_PROTECTED
