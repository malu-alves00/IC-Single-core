`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
78njwnO8kHUizOpJ8vXMhDYbpgoMm9fcK/t+lCQJN6jVmkErdVof1RvMs9IUQoFz
MKKwDm37AqjBDOfIfrtErMnfGEEzJwatfmSVZttunHnJRE4Vk6eEf/RcZQjM2IEG
9+m2DsMaJAJGhCAeavEYyjPD/zAHLWUjMii0URremt611FUvlrzmn4Y+r7uWuVHq
645R3FZHIBBsLNMblzhhGLXEYy9mqrl46W8r7V6jTFnwBn3TWbhnSUTehOD/dyyM
dAkPHWdpt3BVb/44pAPuUA3QCsfnmYxvOVq0W0Onkqa8S4t3AyPWv5Hl58C0JYtl
ZkOs+dAyW+L2id/urwmSdNM5P+Fym51TJD03FOYOGaMzXPQvrKqkijfNv/DMT/S8
8HQdWLF2xFHhlIKvZ6xf2I/lnWpAZx+PHxLDTZkIZbXx0b2Mqfc8uwFAeN5D9Nlp
6DsvbqS6SGrY7+g47UwcCAMzPDvCeGIGSE1v5bsL6RhVQCd3PiqhX9GVHUix4qhD
iaBegOOXB2OVpNbPQcIduCiP3ZG97F/rQOoqdmm0ZdLeco5lwM/fhCkRUKXgU3IV
4VULpCPtZfy7iqgZ7f5o8WemVC+3cjDKxHINBgk15JJ5bWAeFlhDYMH83xP3rKqZ
XumKssYA2NYlrgz0mpuiUuvBGPVnC1XhwRgkotxdIsNqgvna2lUQHuHAcj7jh8H3
rzszDriZwPVWp4vVqW4xQP7xxV0A5T+Bshs38pwPBqYSzB66vu1MSLeMobZpxyZD
p3kz1ZgyVzKwtZLxW9+IbYktAbqqWp4kVDTny1nu2g1jjs0RwOABSeZknIMIdNv7
/uk/Y/rU8GlQfmBjkN68jqbYhjc7g+DZv33q6hdknL0Rx4GXtaDuZg9FcYKcD6+1
TkMCeN8aBivgpeKesk+xlXqVbZtJi684bjab6Sy6BUJnCnn8Q4a43r/CxgsPtCTV
P+sP7uW5BFDuHio4n1nQVIgwJbp5HzN8LMiEepGSif1LxHGLUV1ofZyCCF2r5fDi
re4d2+Id7RWjgCeEyRxbCkXkJU8J/ZQliezMHtPZ0KAMcEquQGLINBCBV4HvViZp
0dAeYQrc3E4uyE8qp7QZvTCVSh7pRLmJ0N5kzNDUN6RGk2HIBFdfeHcnrYyCD6Ui
vz1RK4joSG/GId3GDAON5UEraxhOijwewxLoqkXYTmbhBnAkL8S2Pd5ThqiRzMTL
Lx69gU1IZojf+ZZ2VDQx0dgRihG9f5i1DiO9Rk71vfSo47Ih3rHTlJ7LtJC0JEFf
hH1yXp1gKTBEHJoajc2YmUZDW4+euP1ZbH6Ihye3nSFKpIM/Y5mRrITRy6A0E/w7
HiRbf6FjhsYq5v0qKDcD7fYpTi9Crrldsu8e0l7SZrqQRq4f7IbmhVkZlJ+6QQ7T
V6DeUP4eH7rXpU/PbeZLHNVQG9cpSPITbwsGNHDS7cJ3zf05r9Bi5MZr5j/DHNuN
iqItsJvTgHMS1xuW+2ODY4tHqht4XEagQzWQ/SSz9qx/5xorLxav+gVD496C7oNl
J+UlI3A+sp6xi81X3CKcY5ZAlkqrmbEqx6k2uAF8uzIpqqJ1qnSqbP57HxtglWHa
nRlh4NDTF91C4w9TbrmdJA8XDA61zuU2R4tEQ13SJli5oiuWBrr2soT+BpnExmPd
RXpTqIAkpQZefl+5y6Agr9J1SJaAFXYkFU8vNLY9uPDWF47EFMwXat+fwP5afOVQ
mNBkup9uDIAlb5o+glVQbxX4pQMkAKNlApOxpfwa36rr92W5P5JrYUAB2lQT1FvM
mtH6mIxkBaTyle6/DtDctNjHFiN31JyAcNEturOQ3yX95OF7kT3IqUztRl7QODPU
JfeCxGB0y5e5eR3eW/nKYsYm03HtSBnRDeEr+6BhB6Y+h4h3k1u5DylfVOlIX23Z
D6iiaTJqCqEfRKpvOld1j7tGdiM0hQdhdXFSzyH3VpOv0tV+3sy5nieWLXYz9Gp0
qmXzw4zLkA0VH5Zzz7pvPLrKnzLNxjmUZkhPEvspW2oP47GIWp8XnLzsXWXaZq+w
0d9vRujmeaWLuuBQptsEgWSCL6vX2EZXXxFhXMq9JuDNdwOCSWd95dw9OcQs7zYk
KFVImhkNhW1ZX7KaUx/1A16qcJu2J0ai0n9ZBowSf713lFvTEJYhQ3IUpB6vbf5z
aw8AaTtvr8m7CN3+zwZfwTpBKCPJc9U5kOcESfnq6ng1gHomqVMVdr+Ri2K3MM8v
YhVWE/pvjWVbB9dr5+WKxEu+ypXJGhzbmyuZcKtpNOmraciqQnoDohjKK27VYaBZ
T+CE/4W8OD/T/qzJgvE16WnUo6hX3SAF5SVftM5ne69x1fvCn/riefaR56NLux+v
ANnQf4KilOBNhivlyxSqhAgfnkhQOAriec025Hm/qCrAjv+9js35wV/rxMDz082A
oWdnN/6fJYq7WaptILm7tHuiR80Ko1OZfjY2VKsAgUogRmIKNB1T9jE5q497P0UT
MgRdBt3pOlTVc3eJTTzCnexZaii0xAo+8Hj749VK3y+2Le63hqwIBX7scHZ3iPlZ
uJ+5L2UUuqikpQ+y9sMExJ6Yzt3fjomkrjPmWOB3W+knS0XA+HWnMRICuYqdx3UU
4JzV5OMct4ITKT9+Uo7D4dNCoVnyLlqsSM8pVdT3aryzgRmJ8aLQ9JRKoKvgvTfm
XttuIWwXHQjwXg8VbBvAR8GKGPiB2bc1FNmszBJIp2oETQXO9/WSb0aDnzou5Tfy
4wjKhixNyD61ss4LHJmOTKqs9ooqFTDFZSsfazaWNmsGZ/dd87aLAXaGCu7DM+L6
/s5fh/6oJK9UtdX13uXHk8yn2w9cfoNXGFzMISHfGeED9x+QipZVYbG5/SLIa8HD
m1EJ4HUhMcThYFtNhL5+5WccHQJ2rp1pnkvOsRsuf9qN433Se7xNlecu90qNGyoB
+lwKr/FP+UNPAMDSFuFEpRZhSqprlbV8eat5G0poMTirIQH8gPtih06120tlmjRY
GJb/We/LNTzUeHTvjWmv5EQJBPaqjv0tDGar2jAOY5TAyylRy7L+GEvh+l/eMEio
AcafO4yi2M3XS7CT3F6reGRPFlG8t83TsLoXx8wgzXMYk5qeT/6H4jsiVopjS2NB
I1Ox5pGDDUjs2argJzKs0AFLbGKOqq72Or7yETAbyrcqwaOT/1za1PXrCKv6gkBE
1wxIsCRXQF59ALhfxRh8HuPLnBGeDSTYJ8dR36ZDp+CePVov6KhGcvmwoKEWjEb1
psy1VnBU1N3ZBuFmandqWLaM+EMB0V13xjAziyVw60W+PZL4iYgSHg0z8vpQPxe8
VR/zY5Px8bp9xumDtj/5RIMfWSbOltNvKNNcDXsW33XMiFO2cmnvf7Zi3VUTNP2q
uYyTk2pmEVVq5AEDcSUGe1k63U+kLAGA/oAMqBPcI+bfqwxJcqg71L8uvEby2/WM
n6wXBDkmSFNBfwYAq7jdbAiFO0qo0QiSXXXRSiWBx0qx48jk0vxMSd36PdT1sejX
TklBPJLTehebI/C9wFNh3r3NAByLRAyCJPnNqlgNLxuokW6DoNUtHl5ja5x5AUUs
4uNO22oa5HGgx0QnzX4IUo50iJP8bUXo1eVkPOQDdMLaG1nbl/xGTAkvoidFiWBY
AHpHGOU4f9UPBLD+9I1Nwi3D/xiwK22qamT9Fbd55qO+6NY4gq4yACX2AsvFZp5p
joPe2VOL/gSipi0ajwd0q6XDihqnNJ6kJYssNUJA7VqhAWrG1ZDfAR7vNkOy5OG0
jGoseG3i2c220wy0ZyPiOmajXEkIARv939SNgA0CYFDfYr7Mpq3RpgFJwvynd/pj
FbvppBqzs50YenjX6hV08femHtWgC7EiE+83mXlE6E5beh/pOCTmi75yOFzlDfI/
pX6ED31m1jtCiwwMQQCSC8+ROPWFmN+56Yqoeg8bKWHmliQcd6k0QXgJZz4eoW2a
+X8fADzcg1KdCaPIJ2kPw0Nj54XbV+JCLXO7jnaZ18w8quHfhUPPzApAsw18nAki
yjxNcZufJNd3hH6HsaBs8ILjnbNYxcYxyhuOuiXMbA3or2fqU8eMrP/LMZ6phifk
m91OgJWD8t52KxSm5sdgVnUnZ4oLp1jXMoKOlsfKse125IHccTnc3UpALPAdoC6r
hMXX1vZJIYr+eMnV1joFbwodx9N9O37UOkYbWCiMdQqWvgjQnPXEsYRGLTZHGI8T
kO2gepIsVKDsdMPYo+ZA+peGrTu/cWwbW0eBjzu5xZ8QvUNldJvgx3VnMeFUBB5p
gM842CrWic8vjas658J85Ky0znFbCjHkztjTFkrkOVmM4M/Yufb5qCWRabpH3srO
/9eaiwIZtXmzeeUc6TsGkWcXN+vy3O3pYyBsHg+wUssBiK4q1MWtzC7eMRI7ZL/K
dOl5sh6XxaCChNRcnrJjNF7lvTAR4pFm+EmrAAWWtxRvLTUFVUnrLxzjWFCOFZke
0X/q4Jk4DXOO7Zwydq20JH3uKkzvv0Gq4geZyR9rjnw408opayDcLm+p1mUPsc/z
IB5fY/oejpdwJi0dcWiLFQmlkdbO7ZwGApBR0RkctDZnAmKfgxdfNtBpMf+Ve2w6
mcoeRgIXfJj1Dj2EcmyjFPG8/X03qS/waW7iFUxuaYf9ZZt10T+sdx/vrP3JsW2n
bEsdd2LTGxoOD3AaQ9LBkhG48rgyNiI81fTMwZu532nl6SVf+HL408SJykEHGf09
9hKWHt1wQ8qj1Q2xJwhzsSsVbo+yzCIyXO4wNaMmuH6DgDodxcmcVnHG4guVQGR8
f8M98qjNL88EysoP4qws7QGxYHdrecZBbXPTU6ExvGG/nnQjCvWAuRWbsnFHcKxa
AMW53f5vMKiaqZhDs+XQwvDFwLg7IiIVxl0awYWvOAddZAXIjNdifDrAtchf+iIV
OceJk8UfpzRZYIbJcUDxPSRc7w4GRr2arDlDSdgoGbPiqGNZoMQ/372Ssm794OVv
xZxsHulxNtdZlrWc4q8xT/kTRyVn5sE2w44XkpyWllCngBEvFXDtmSEWUIExxSWi
rWnvYCL6wm6byNYGKmS63a3Ev6oAui/eTQu5E6SpP2Zo5McBAFX4YK8INPxd+d/u
gNhifRp4naFAal5NPPeyeKchK/bUCGvBC5+FfJaJJBZAABD5ldZRvnFYh5Jk2rKo
n6kdWRikumYG6bLGz/TJXEoJGqZ1llaxerNseEVO/D+j7NzOT7u47z9l9c6B0lYZ
uD+GJp68n8pMk5SyafzsNAyStJ8WQXeOUx6cs/dKLCOtyjird1u+Si1JO+8+YNYt
/3D+h8ogmTlqrn4ixyQGIhjfbb4uEuLlTxHcrx84+yF7ODX/9rEc3SuSQNajaqJ2
92wDjIcoWsNltwWlgQExsDAX+NaLkGZjQgmaSocuO0ujzQYeB4l23GrK1+5fldZ5
u2G+6qdA4BiSC+pMIQ8m2jVXCWre2fyNxwQ/2uLVGfk48yIyjaLf3NZ7SzpWt43e
iwVSWVULV+QtM+tK65YN37aNLV1956I4fKUq2B3wYuDRfPm7/O5IMFx1urUydN5w
OiCWmPdG/MO+IWubwBLeS9C4g4+cMEuOypcW7wYjuZvq+7QtAYEe374iAYdz5CZP
o6B6pU9CjqcKDF1Y3tq6hBrcT9P5aAF+SKl4/vqJK9oeu+QvBSbaPuMsoUfBo9Jl
ZI4u8CVowPesV3zE5dJXUq9xxatRS1+cPCzswE3/Iu0rFPwoRH1whcsBiIWFJElJ
LwMxDApxHdAOy8/YGS1AIEh6q2kENe37lWnDX5qG/vsR+8cXoLQbA/DPu7oMYZ3i
0ENxW9kMjRF0e/WRflQtxt+MAAkRHHSvCeff16WTZoPfNF5x1jTCKFPypiUPtFrM
V9wQQSRlagU28Hh/ayP5138008x+UMoDTvT0jyWgE1xzQVY5g4o7+A24OuFbemfw
ZSVjAN7tijF3JKtoYPh8w9q6DupqWGp+pnikXe8CeTBQ9TLcZg0bys0tbb7Z6h8h
+f8GbzvDpBZrpoapmIF3KDNLLp0dpbf6/DBuOeI+ctcLLu38qbyygW8f7VoGowtu
L60u4K9wHm6bsGkxVY+5rfbv4+wTX0VR+K5yZnMPUqMo9CNA0//9pE4TeljZdM5W
K80AxunMcJEXFONMZ0iHxrEuDiNefoEPvSVeqnFuq5qvH4LjIMHO6btJzCIVEpaw
Et9V33DkEHu2vfcokmCK851qaMzbYNyjgKQ9wz6Ec86P1O3sVt1AdYRftaoaELKZ
E3Om7vjpaKzsN9+95NMFfNfc7btp7PY9kBG+83OSNH1rNCHAmrKw7QFF4dKK0JEn
/36PQhhxYAAZH0J54+dIlhTMlX/fWiQ3edXerDx3Gk8ozHHU2juoVhGb209iYcqs
JgbMSlYTjj4k6jARt6VMHVwtRcs1qHzIpDx6YGTDPlBN7RD7witOhk6wUnexfErv
wZkl/hdTODAhWn/nAVV3SrGt29YkIm6mMGKYIu6QXcR8XzT5lJ0p39QGHaDIco1o
EfEllDoihEd1cv4c8/i54NIV+zpxLMaDrXXzMfs2aipK5dk+gHVu55RFkA84O7Qh
Agwkdtz12qdvjQSPAmqpdGAQBrUW5ViXNyJwFCJH8kUGepfI0mTptJjYAG3xYzH4
CCXEQfJ0RsTolSPdnCCEwSI5OqIIQ0r8Pfp0VZPaC8n7RaMb/QINLsCOj6+TCGKQ
Xl/t7EbP/8qtuA0ahEHPdfSUwMhrrubaXW7LDjbdNIMoX8vRbaIDxbVZaj+3m0qp
EVKPaeE7lVPj5vOTaVPQmOj7MWHXJUVstxLFJrZfFYJSZk0fE4h0GoKgMBa/82j6
ZdifF6SLc/++VWflVUnuvPpdcznbq9FZSvlv1KpxbvsTs9ruOlMmNK6oBwKKmipv
fo/u57H1bG+Wgeo+NO9DXaIaMz5/l0o1dPDtqn63IZ84orV3NnLMpvxJODUcIoJn
q5lo/YlL6GDlhvvN+/kVOcrZYnsjW0GoMpaHP3RPPac1yVgqTe1/b62vnjRSxFjN
Qf7uuV23IVz4sO8Pb6+vSsT6BS1zDzPIt/3WUYRwDaps1gBApVyMKCLUgCW7+qxc
FnX+hX/BBbVq0B1KpUakuWdCDNuCymB+0AOp0uYEX775qUk2iquhji3mFadl2sVf
k5bQunuMOWbQ1D0+tslD1/352tXNDNh1uwqt72OtieeR6HY9DUOHeQQUeAX4iXTv
rDjQwSTIboHbvTLiF203cUxEuD7+j6NxG0kxGftj+SY4A7NILui1PtBZPi3+FFuK
vKXcdKPN1VKg8PlAZK7Jws/scJVi6QMlWuAuYi84536Er3BGp53zNXtIEVzcGwjV
2/h9KMpB+i1yxQS5m4QGDbN7JLaS+w/Anfcag7DaCx91jV3gInzEVITf0AtEGiNO
E6qAZ/vRs+A1209DGuRj5AUWQxLaMXqlG+hnhyHWlehnSJJ7sDpcWcxpCnlaxcdM
a/5Bk6CuuFg38ZRV91JeGmht4S+FEoOIFo2GUeXR+hC6iYmFLE4LvcsYtJma+vE/
ZldL42AKPlmp3rrZpNAEDZZgREzN9vCy7CSi1nVyJXJrUD/d26Y6LW61+BgWSrKQ
5YffWtLNCA2knT/pbE4c/MDHsywY+h+VbHz2w+wBGTLbRSPN2KivBMrJs7STwOBl
edb4y4C0avtbSnfFq+Tg9jjQ4GNlqLypi/rVu37ON29kFJ5AwrhGvT4tRwe39J73
9WnArYqpglBKje9qSppVl2unxsfuA18rqrpKNHxVJqRJc8naiNoYzM3SJUGzl4o7
yuA/L2QeHw5kQSWdmbEywsZ+CDkj/z6tRVJuEcuGbJtu3BxF6IYwXtZxSbMVxj13
jsj9BH2eU8X5ai+ZZaYUZS1j/vyfHHdiVLPe3mRporKAR4rhbDApRuY0NP8Ul2He
jYHNMTTt7aJF0EqIcznM7GGRn6fGwQNXu7vAxiw2jfVj+TMYnxoiUpoHSRywJh0J
8ZBs1fVfHAid6DcbW6FPCRkEWjUWFZ4v/lBhOcAWd2LxF3F0OPs93HxCORY2gvRh
G8ACFVOUJZ3v34sFroAjY/CPqRu8F0WoeVmdY9KXum8YNOsFB99Ie3hhn1eTEPsi
DNH6ZckJtvzkCGF2eUzFnoI5NP/DkD6PjvQ6jg8v7pk5fFhCJoIJ9mpsZqPUy2ts
oGB/LnKf5L0162AcErDBM+1OO8R2x+frAPMXsncjhMMwZGUqaLGkBOqEyJxIakXS
qxsz95cZiCOBUqM9Q0UF/VTATF5f11jLnNC0heSAxQ+fzKrz4DATIavfBbNTCn2X
VsYlzjEz+KxHCoDRJncLwgRjWzZN+ZiGKbhDuwUd4hjUE9YdwTYkhCYc7rF4MiMs
D1e9oeDxhyGak3G6JqWlb2IWf1mkKvjIxJdd+zfjrfPhcFlzSeQGIhV+ewhCkCV+
CX00F+dYQbtgxbYwKuhsVJoe8gB9lQxsCW5fQ7+CemHlWN0Gy34irW1h3FZqZVc8
B//ZVknuT2S4Cslcm793ZlusTnUlaeebndVHGMr9brazkeRmaJdACwRtVIKiR7pG
yz72YG8NMo9npKVAxIzWCmKwHR9vqE3WNJV0kymSfi3COS/dBwuBYxNqI+7v9E0+
B1fSOXNdWSQa9xCm34f+HiO1MKpsAJlp82qjoTR2oZBjv5nhcrNOItJttMKPSQJs
7HJDk/0ylPpZ5VqkX/bPG/EmIGOvmgyDerWJ7yrziptiOkPSEO2GNIe3za0OUeG2
OPYYRIBpjwACjQOg/5EGr7Nds/toDe1eRKKpZJ/0DdFgDOqc0byj3XPpWx2s/gut
2ZWUV5tssrHl2es/sChJXS8IICiVVy3CmOEUl/7dscQQYnCURfAkuUasGZpDAzAH
O8q0w+ZOt5KTaBqHsk8AEzyRmbS9zS/ZGj3gv9aIT27DRsWyKJo0dvHin3qDRvAf
KYHdtD+CBjs0yEuvR7XJmh3u2iiR2yiedBunSY1GhmWexSZlFJ+lvTzufYpDDfG7
qMHMy5pGZe/JEKniJzq0Jwqo/KSJ7jrz4vSe2c8HFscqicVDABnaJda5T6SiNRuR
URvxJoats+eXiagb03saUjVmo2FFVhClFOaD0TE9bp5gbShJtQMY6SoznK5QKKbq
wMza3/jP68MltYQvbbHAWbEIxGfM60FZLhJ2d5FiDkgtQqwP/yzmvR+G7Zav06jH
W7JDyxlnuooRcEgDojw4SoZZpZ/xNQdx5I7qggfeUWdYepeJgB4gBklZe29oRHIm
yt/N4tj4BRgC7DyPhn7opwaZ/TC1uOfxp4K6d+q0nHPk8guPFN0MgVJ1PiHah3tN
iEywCY34HwiD5lvqH501MIGjFb2Wmm0DuIBpwFIrmnHS4TJmEJrser+Y1RlYCyjv
0d/+9rTLXUGpACP4IpihoKWELWW/9XIarD+udsNGDixvlPzPPaHzab+wqn3dUTte
cWc09NYFgUYfw4D+znaLbioNJyj8sbjKJKNilpkyObZAB5oM6X+sL/xMcv3DdigU
VVTiqIwtgACADavc2aGygb5q1QsOq2jJTUOArjiaLqll8uyQHzftPuN7xc8LeUnK
1Rb18XmL1WoMjw/r0OEdVu3DMX/n6hthlkPXh2GGIndNQ0gIWnIqih9b2E+GovFI
Y9i6pcQ/rQmfJ217+qYtcpLbORIR5Py3x1un54pNfRBfwAcfcX6K4QvzKa9755RJ
YLT+vxF1Jr030gjyBHT/j+Zk0Uv2lqDbHvKonb7j3miKzz6NrFp6g+X605bjYxSi
6Vj17J1/L6xacV2DPxz621tFyvr0oAZXcCQRw0KMvaf/cYlojL3eA5FOUf4+yXgW
xsKTbYARGohon9Ev28DOquJ/Nz//XJl7Q/zDp1K90+UKJheNPWNR6fzp41b/Pz3o
edHW6feGmE8I8NssujPKVPvNWcnMk9GS6ARsdk3xN2EMuvEtTxpdiBVljMRAoqZR
XXbDtrMYBVrIcbaCewdUEM3IjavAZ4tz4dLEQIM6iyKY54+QCs6N5DB/0PA+3Mvv
ClebEyWJp8tw+N1wqJi0unEX/zLr0iBXkF/cOqUm0VsyErssRDvUXhMh7swfETPo
x2Kx6eomW5axlWXElCA+6YZlUNi+r70fX8Wi8OOk6D1vZ2BDgzfVdtWXXG4b0Xx1
YBKCq8lOV8SSjcyO+3+9Lwgd2/lUhwTnTAFvIpHto5Y0+xy/4bDTTw/w08siirx+
tJkPyK8PzlHnbq9ZLxz2s2T+FGLFTE2hOxk4Gtcc9r3bMS3pfYWtLAdKOE9dLzyv
8sNZfI8G3eEQqjleDRRaR2i6OCi2zjpOosaMANMyICR5LBYW2rkwl7Ude+8KtvFC
t8/Aa3FrWW5oM8P2fE2BH0PqPvT6KskD6UrVgKCDgSonrjExrap4lplGCec1gFRu
xV3hxJje9VeINZkeaN5xVJZeArmZtk56oTTKhZE0A3F/6RQIA9WY52i/vq2Fl/QF
JwDuWygbL6SIFZ74WujGa4uZElTqFY4s+ZlopA9vQ/e0HTlh5iKpFLunKhV7IMdv
lXkKV/lermQJbdm950qjZudSIjTRawQimImB5i2QaT0C7+RLKYLIXcqZSJXXZ08n
5Cg6OV56SMqtjqCC73ARz9tRpmgqQzM7JqCqGaEaTSicqwXzht1Q4BhI2FSIukjq
MJunslKyFX3gmWxIDW8scaqeMxHovn2OIGHo/tSBdNnhp3t5VRQw54ncPCyZ6uEu
pDpO+o8lUfLfmaDAJnA4Vkv0ntWYXm/xjX8Z4VuzfiEf7RcaH1ThXjRrWKwwU0FV
/pqG/ttLa+F2dqphFPvCCGS1TDz9epwJSaWuw1eK3iBzlYbyEndCPC/9Hwy3La6Y
xq6iCGq8WcBMCnUgdHjbYgiPHbyjP6xOa1NJ5L8W7VDNFXesF3KGp8jw8Rsdd/0r
Uh92oNOKzs0tyob14xCK2CuVkvfTOiVBMaWrHjA5brF1MpwFSlphVmS90eFVEZYK
6+XL1Z3p6W5S4ODmjF4M7PjgQk2gfY6hPSuqfV7gc0fcEcd62xlgxK3Beoq+iovs
0LxnRYIzdKqUTw5Bb39G9WlbB1qRrdgAMaT5NCqG2MnSoRV/69c7QJrcrC3gf5fY
dVu1Tgv9iScxkA8ZnoRpwvtbLoU4zPylOfo78sKeZT44Zo0r8f2NEql4SgtOH090
/rBJE4q6VKD0XGOz+F9EuI+XeMiBMwEXV6wLEFCkaDY8G7N2zICrPcqexCbtLbpV
qkCHXtHDVarzICNYWwYsZcdAcfS1pJxdceOagD2nlb2mcO4r+xnUpw8WTasdzKWn
v+s6pEE8qwCrR1O5nof4X2FZnyGTE31HKd+QxOaeJC1D2KyNo7675hh+4LWbjjKF
QbDRWeJUTnT2vOI++KVtuUq1wh11+UCXH0bKzIThNYbc+1jNsH1iU8S/C/bKKOYB
lbXkSXrCRoG2kKYJwicB5eDQxcgS5X4awB4giwD+ysN76ikyz1XfWqQr5i6pE6lJ
sqFmwDzHTpQEbbUInOY/lh08QGJpF4Gq+5sADmeVFLenpoHza05y53KvYZPPXLf/
AonlraNMf8jWlEVqQxs17jO0yWfXjMu8nlXnkrxn1gKlGYvAtIjXw1VLlo6O0ibW
HXpEwu7qrJ10SyYRTxPnVY48R5UaiTHx904cm0My+xkeuDvm1t65FvU/mDL4kR0R
tTIrmq/xNAulX5jkGkGbSejwgUsfoeDbhF4nN1dy3rGP+bBPUlq2wy/0YpoZl8/H
GLpv9vjmvl+ajLXm/CNUA9AkqKpcSR6afrDAWLrxfHozsmoKJRIgwupBU4Xo34Z1
qi7dSN/b20TyqnTga511s17xCYIq2IKuJ8T7LOoQT71H9AOlYGnt1uQu304C0cNt
wUeRtD2fdjkuiJ8Yc0IAautSQwgzOTUgT3jgBN/pqWQbr0ywKfsjT6U8WbN1Q3B0
gYtn2XW9GgmfZmdb0SkvmhRgZyq5ofGRGwQ/lgK58cuICJ0ERdNwNw2xM5a4O7JA
JYO/8R+A4f/x2Yuss+JT7Ou9DpTAY1IbjK6DG9EI1pfKfLRfB93MTvmaGDG6h44Q
yFNNfZ4p52lVsHHFKi1201TotTLpPyyE3m2S6T0tU0wpKSrbIsMwca8vQOhLmbhe
ditzEIXjRGSIoINGBeAHtfnpW9iObaMZPwtmIkB7hRI8sNv95ps1Ewjved26GMoi
gtZCWv5OyK+3L7n3A6gNBN7+6yiUjKPO5aVlu6RMjljWyjzMp85/qpX3zBCb6UuY
DOoQ8o427yoGmRSgv3g+J+JpD9/pneEyDk9nLa6tDk4oQmVFipWJlFGuvv9WJRIA
V9xP9rSgYw1H9Lnd3cytx1qUjojn38zFAMngYuawKzaAWkdt2hTMwJAZKq3Rx5bx
EmSGrFqqUWdAt8iawkdQPCsY6Tk0JddHrwxm+omOUbsAQj5f9Jmprz5wEvx40Cuw
/4gZPORQBXc4Dcc3qIHGL7+wdTvMMeUfbCLTOKsJ6J1+3uLVOR7RAN0LWbJ2GQAI
5l8lkwuGB0VWOa6rII7T9wp1vOSm1RvZcCb+nnMkIJPjC4R1T5tiiZoF7KCdEB7h
dfbgchoOKpceGiUHRLMmfpp+NZ4nv3VmbrXnQEpLtrn8XLUvKar9KRJKfyeGo4Qc
ZUPpn8fLVVSf1mgKEuxG7/BEGFGGpGzsBjRvXdpliGGF30/b+EUQA8qRUVu4JaJD
8vf8g1BuUsiWFLfYfubrLI2O0qAGdc0b1oxFY6x37km20PK/0bL9XfuNvt6ZbNTV
qjfLIAmm+HwokPIvWYhC2I8jZBF4DREEe6afvY1OvtERF7pe9KVEy954NgfC5IWw
WE6EJWL6i4jEtA6YWfwkDYHhWCHiHA+vYTny9OfCuNJ43pDPGB7gRgNjjht4nsmZ
5bEILVEXJoAJOLGaw+Wn05JLLnfWbb7tRsKEV51hq8AB1iZdFPouHRsJCfYTM9ce
GsFzYvkSZ0wOi9oi9Sw7PDVr+vp4sX2pUy1L0WImlFc5jihSOCQlh8qlu+kyUUqI
XN3PiWqqXJx0TerYVeq3EWjt3DBO4LB6gJc36hWpudwvWJU/7H6wd3YhSWEurSeS
5KrEHomPIY3dwlxQcJ4JDtU/MoTrvtWa3Zc7CvrfS1Cg35zY/Xf+Af5qYPADkA+L
4ipgIfU33NMoNP1gRiBomukfj+Gr6DGnpAhGOJ6SW2zHSaPLICjAM9Vf0EiP0lty
zA3p2ra940hoaO3GNuCD+HDwIBE3SzceEaIwkIjxtwJfgs6uboeCRFQY4rw6fLjQ
GQ8RtaVV/y/d7L7BEpcaXoti/Y7q2FQ1esKUZn/dQNuwap8HaSfY9JWsBvmkFOXt
gRhmDsacGDHmAuFOW5uniSoNT2hIs81PwMd27RSpPwfhZldmHyVs916Ti6qHJaN2
3xDnJ5Fa0q/hIJe+Cf+1SV8PSwTeFlEotcRJ/TrupqCJyptCE6kWgduN5oTKKVeT
Hi4+k6dEs5PyI+KIAFlYJJv9PBn+8vhy+u+0hht5savAUG/F0rlzWE57CtrCeBSG
Nr/ehxkfMwKe9BiUJajGWeBr075KyckfHvCrVRA6Mb1SYev92PgRwPDexGFeuP4p
Lu+bfFWM6bVUko1C6nSbUXmELgEKVYnHrUo50M7w2O+Us0L2gPf2oZJDyqizbSzj
+uKfunBYxjGTxuuSLY7cmFUxzeyRRdVA9ZU9uDB6tIDHg6Slzs7cshPu6MBphoV/
xM+lg4Z45PGPoGSRbsgDDdKsnTopPNyZp2DtFjQ+xrEgQ8/X0qm0YIjnxJBFYAPF
nhdajMBUI37oIq2bha4vaG5SxzeTMmOiHnvC5YjsMwkLuCV8jwZ1SoE+lF5j2sN9
Eq6qNE0+bjswYFC9IUzdAmRJSsbXS22XbSTVkZuiVJVpIOYtDoUeMaUL/SDPxUGI
v16JG5RMHPXTav2qA9EZjXTmow8myZmqftISr4J2MYCVG3Wgy3b1oAfVZdrc/G81
PXyihWlBGfnAPyqGFA4KF34w69X2EvlS5QApuEIGU8zl7jP4HKifFSyOcJEsKc6/
u7JDQ1z/QFaiv5sozcG1na2flvleGvr5q6yAdmEelaLuVYfj6rySXnnDKA7Y+491
0xeIrlp0MqFfRSZ92A/+hAfafbiKulATxMaWZuHWZng2eoJquCH+1TjqT/dsi71w
QtvlGy+EFba/dA9NfREwiY2Np9nZbK6k/r8DDb3rynBa1JVBQczZWTb28Ad1IewP
HsKrIXNB6ih0l5ZwJBNDjS29xeg5waBPJVmKgYzOjuNN756RQKpVwbVaTk5Tp5Tr
PdUY9OXRC5Ax5ZPWMXoofjzaxWCUSfUBJIPF4JPWGJRZbWX9irOwRaWf9Nsaa/u9
vnW1YXsT2HXaH8isPM/0zsVDQehHx2jBSpgiftfgRCSX2U/7/JFCye1cHbM33VF4
iFzdeq1IW6+8vwAqtaADTMs3Wk17QI5iKL7Hh93KNkbe/e3+Hoj2TAGSgHPWCHBD
0GbeU4IRELpV1YFsZArzFOb4lvIr+ObKS7t7xeQtTuJKreUR1ZerQDcW545D9qK1
8c6j5FyZJjxm7z3cUCUxUXJloZFAQ33BpXCE8sLVGUfdwCN9WIqhXawYIZkCyf2x
1/nsrapinloOjlBJv6aGczi1HjifUKMXcS0Ccau/ONkY7O7N5Rppq0itDlMLUb8R
30EMEz4Qw0jaWdgs8Frjr+gBcF3zUmm3T6+WnzBa5GIlAKnQ1zwRg4MxsNzsrHcu
+qimobeepAylnpVMUrZacCsHRHJqxlQjtgcd50JdPVtZWz3m4sBdDgI+JZ9CSo9x
IVKybwkQuboIuwn9FXDy7bhbS7XkAEgyucGdL0RsljymY7O+UivfNthdmmPmLyoW
Pwdf8KMEDwM2kKjqToYX8i4C1ZbjzSGGEAFlfexqw2nWBA523bVihQPAKbq1GcTR
6a/VWgm80W721ievtXYzuulqDKYgraQ5weQpLik2T2tlpETUU8CPhs3VtvJepU9b
fHFg3xx2rN/2oEAa7Dk7orPcZzehTYFbejdMsrNBoJ6RK7q5zk+EXO1Mlsl+HByx
bRpKtOJT5SudBOQOCgBtAld80Rtst02HIQllPXJBrdOt9a5Cl8A8pWsUIup4dCBD
sRvbmZF4PJGcPGvnts0ohndbyaeF5zAe9jonofdM5WfvFbD2DbWOWVAmFfgMXp6L
CBssbxOJkRPPXdq77Ez5GF3HNM2/SY1AGL37iW2eFfpwZu3v9v8XoqOtYWwQ4xAS
jep8AdRUn+RdL8ymcYgIdbwZMWWozd3d71D2s0VyxoYQrygbbhDq4D6OpULx+nYq
J+EWiPhvvXEpJmgeOO+boYJjLqsB2Gzafb7LJJmZ1EZQPiMDKFeqMlbEuaLmmH1O
lNirie/JYCfG1GCUVBAZftH1MIxk9MTw5HGP5QvGP9hEF1B1cbX4+UkJm4/3T6qG
Sowp1lhjDfNd4PP6eeTi/GeFVkFSPYGaxbQbfbcm+AuuFqSUSlE8nlgmR3e0A7f3
i5FRME9U7IGp74oAWYnbFP3CgiA8pmXqkfhCf+354td/Z+enjpYJqL803N+oCrmy
Mw+MI8xz4luACxQDGzCa8zANNix4GZ7v1IONRfxOLBtjUwTmXZi0Pa+tgqax1LZo
3ZmbMqn7tcSNdKg4gLG43gNXYcs4kQzvpp2zjgiFwJmTw9NgapGt01tltt9gsPH6
HP+/LryENWVPDuz4o8lMLdHxdhfd3ydt/WPxzqZ2z5J07GWfL1PGknNNS7/z5nnt
6D9c5lzENAKTR/XIy0bi24ZsK+ug7ZK90hq8ilQrKQBN5git7PNGAm7oeBuS8uDi
2peNLhUA52xIaUMJUIJ+HM4fmoczN1qM2L+FVVbRe9qz488gc5DGQoRZdtaeCUj/
l+KZOK9OGbOBE23MvxBnr48B7FYLuA602H3DLtpBT4AAXAvAra96D+3/wpIGcMxo
sOt/Ecr/N9mBOupj0OPpw7EzSshyuZulV3OQXHteUMyQb1ViFKtwL6FYw24y8662
/tebS0ymkk5voQoDer/tsw37TatlP8Dog8DLg4Ba4bkned0CumWOO+KFhpCTLd0d
yexmieKt5aBXsXBEccRb44VURVpcp/U6X/s1YorXego0+huibXJpByB8dRSVl8Zs
2zGDibQXJed55iqJ6DqfEh+2r3gpOHQOJ6ny8/qmYR/oqgIZTA3mMKykHm7Ru9Rp
bAlgbTJGGgaBbP83bFsDi6Me+VGoil8/f3WHuDoDXjAQCatpLVFgUJaQ6ZD1GNw7
LOv8nQRfIAKudsirIoFz8REI+PDzngx7DS00pET9ImEDVG6v0qthgParnXHFEeNo
lvssnoF62j8TxY6bH2URMejeANRcKwJ93cz3KqNvEnWx+y/hQ6up6WKuxqT8SXEC
HK21Pc5A7/iQlRzgBdAcF3FEGDTrDyyx523CcZbyi9ALcpP5iTg6HkTUvTABiYsb
eW2uiJKcS/R2r4yaqLI2BhVqUWUSQtsws/GhfEjrvY7iLVlj2QNdFHuagMWwP1EV
TjfQQ8TstooJo4cyHS3AlTud7meijLyF5nHFVfd5ejS1s2yLNRJC1ASG/nariVjb
gHiV11O45+3lfvSN2M/bfyOxJ+fUDqx/osv4RVt2vJnMjlaUj7o4n7sGP/SIBf90
oKQToVVrS5n/JiK+38v8fYJByfC5B+Ws3SzEKgeXbg83l11RrxG8hcQlK6pNTPfV
ABd81FNCGYr5sY1QrSkL0VOVEG3WcuaxS7ah9IG70tCHWokZz/8+2Iqv72ah0f3w
C6GlMaz91zexEt5SclLpdxgLSIz7rWMeVRyMX9tukqgKccExRVtfs4uY6kRNFOmQ
iaR5iOpq27pXfwJE/lZ4zMBHRNcTz1gkbh0+3WppSwCkBAzNe7fy3L7OK40UT/15
BVnHZuDU9udx6u1OxqhltMf4qZtD5AkoVWf9OTGNAL1YBUWd/nonr6RkSzUnidyy
g8rD8yzbsifvv61f0qQqTyYYDa9QpstgNaN1AlZEf0haB3yY9/+U14OxmsVb3BIu
PqvBodEmhAw9Odiv1q6wBETEl3DXTKVKs7bnnQhjVwtNcdATtclhjBEilffXBnSD
WRqslAg0IbIgqWL7AFilhUkyfCW3WuNs4hA2+7+YYEVfDSpFeFceL5O4YDyKmpD7
qOVNubqfrzmXLPGIGC14JU5I876UPBVIoWLBR/Lfq9IBbNoHbP2osFUroSBurEfe
825y4XvaKkfe10sv24rStLinFRlZDVfhwcsifwtNef10p8O+LF3ubsKpZROJoEsd
YVUNnPR+u4OCGB9Rapn5BKtQ4Lm2zjFr3BYx2OHWVqUDczAv/Yy8icawIhRxiW/M
9hcnZUcSXIXlCNiVfeP0aljIWoBuy3mvXsBdJWiihaWkx088J4JxnyEBPBS4tJsd
fAWmazOmvPMjkCQ/mFs1dJibGnCaZ4vomOtv8Kv1K/n0HlXXF+IBdNEWHyjzBpn/
W7HXPPjZn1bnFQQHV0J5PgaoqUcEW4W4qpclmgddwqe0WkQ4x6b/ilmvpezKr1i1
Si5VOsI375O3QiM1cH6k1g4PSIIy6zoDdMK2m0AZBo6o0mE7CTUPW4m3Da01nMu+
kZ22pYJ3XGelWc9rJfodb2TQDWRhOjVtPjpIwpFqBnyGaGtCZNfp0QQvuWNg71WP
A1wMEc7PO0LydkYBrZnCMPr8jgw4j7uHA1dJE/l+kshtdOgZ6o69IDfsxd4pRnNz
ZKGbDqwLgw+ASYuGhkkqz0Ku/saXGeHahts70uk7p03lRdPxyHbOj6UdM7w39IjN
jqbDtQL6/cKWkCVRlaPHSF7bswe4VIcn/AYuss2zgOTQb51+6ccMRgeY+73YWfwd
8mD1JRPswXmPuAAQxma+PCMkoy+k9oiY0ZNI78UzKILeeQgvzQT9sWKPEgjX9OpO
24dAFT/8+mo5Pi2LCApaE4FR2w6qVQEDqcIlMsBZziSEOKqmfGDORmWYHme84H4R
1PtaDvqUDg9ZRGNksKHK/ze/jhO971Zu4sie/0Jcoay8922FwB+wPA9JAPKvygb2
FzArrn4WBotdJCn6XOK91wh1Rj8hUVCf7oxFTklRWGdS6kW534E2OHWb/7j5h3Qu
bYx9CrrqmPY/jOq2kGsYvrDIoo9GbrDcjSQ4GBWfyLcZnuyjYJiAq62uCIJp3Ggj
dDg5FSxHrCpt+XrY832MQ6r772CMpG/F9Po4uD/8fxP2r1uX2wPFbNCTy0OoIB/i
4lxEdIbOUSFgcrx9FWgeVjTE5+YEyqMobWoNwfXv4kG678/eivaKERBtn1ck3kDz
/awchQ0DhhuEGQVlMZxNfWHIf4wa5qrd4DQAGB4JXAIulvwlqtc6hHxuRhJ+4+aB
v4I/IvglFGttYT2J5l9ho4aXukzebII4jvYVSFc2eTjQFH6M2OUlT345S3WWSvui
W4o8x+mJpgpdZgyDmfrQSKe+PWFW/hwwKlBymRbB2OsF/dfy9Z8KAk5SjhvJZR5f
VmtLEhoh2j3+e8Wwa1oQO0jb8Jb7BMEKqIc+G5aVOxUVby4mT3Jrq7HWw1GFfUNw
dA0VmpK1YWK8LRMrCHpOsI6ZgKxZ8O/WsmGSwxRTUh57Kh3GxHL3I6ldaMwI6FLN
ykq7nyK6H7gnROy/8cH0BQdxo6Hgie8WbqMvwzdcC5bK+tMsljgWa7C/pGnKTB/M
pQEgGekO+eygDWAol1Qse/QN39m5z/BibvYXt6tFse5ZKmlZBqEFmgFHSVH4KY+F
J056PHv/2MItEVX9Z99droAcz+MbWmOIF8Qm/nSRpUe/rxK6KUk0UiYB5kCnKVDH
h1TFGMalYYQ+7Ercj+tUDASpEe2upeDy3FacvHnr6/ESvZfoBpUEXbE2PsOTuuWm
jn3b8nbwMRlIb+DKwePXm+K40M9FvzoHjw0h3CSagkS38kvYrS+63DLoWwK3bdPL
0PkPdVuMXasvkcqWhIstwujgKqpbrz9OWSuFns4f4wWih1mtW8wdVll6bEn7wsWy
Q7TefA9Bs0zsSW6HlPiR8Pd91+UayjmNFIaotEp/Jazq42zJdyVWpYc8xWAW44BL
grZF4TaXIcJ/dIX/+xxkcVt+p9XYbeIFcJ9Vau5+krzyBJsJBty8zrKusX9NcTvN
bc+6IuwaPDNIuenxaJFW7Ca2yvOKJS81bFIQ9ZBm5GofLYHMtqWbN7Oy2c9rT89s
h9TdNbhuMWw42cu7Tw+9LQiD0Y3YXEx0vBEdZ0VRFfTMzVwJRCZaksFL4Q+Xp0za
sUtmmD0JxBw5t8Z2gM1EN4cHdEzUXRcyXvwhxE/7vDk0Rd0vDYDUQhECCnUDHKcP
XmthOfFNg+cXbMYhIM3xbLCudYG7nxM9FOzqtyV2MdKTYotemcn+ls1MVlssIQed
oGi0Guy506Y1dKvAeuPD2YvFqz+zGc57ctflEoy1oMsJxxU3Tq9Rbc/gbk69Hp5z
D1nMdRfyDTsZQy4QmLLmEg7wXRm0Qq6OG4BFrU1OA/XEkaB9hSNf0YpXOcqivKuL
V5ewOHVYpPj1Ol+J5338BRBWRnejxTqYOYkUeLraVxca9AZiri+iGv899QE5xy62
n7L0/Jz8bEfK/SB607lGM1FZAdorbrrRaJps03GhKuMsyBG4K/lCr7O0DowdahR4
FPuSJjpLWkqA9oqhAtSQlrmUSVcYyvqNCXZrwAB2k/sRwKLS84lmhirFVohEhI72
4+96mssKED3GfEXWAaGSADgKWFCm6u9JgGa3T6WnW1/LtGQrpwfPgN5KnXJJw8MB
syW4ydHr8xw/M8WNQ/QL/9yThv6vKFDVAmwUN3lrzUibwzX5urFjsKoGrZaGHJWI
MuIIw5si6KPaIcRKLliXGmoP/6+rYHfdtE/gNQy3BDoXr1bmlbnGnxq3A218ZuxC
OJU2rHBPmWthTh9pktFZOhMuBI0ad4i0EyH8l2VO6MsmkSpVC9JWl9VUe67GAmOg
xE4ylGxEaf71FdXUXcufur/KXixGRKtPq/+6BtGJv2j+IWySQIc6h+BEw7HMiBZg
g/9UG0lXMe6Uqeigz4BcmCXUDZhrxy8U9TWbBZHETpeDqdao09gPPY9+zJf0NoKt
ClXSBPwhMWPU4xVrZNZl2dkO8B5KpnhG1ow5UNPdLitlLV7jsJssWm2rdTlArvXZ
5MCfej4TFVFjbkjEphSg/Q/Xf7vu3pHKWPq2PBYoIugyez2PQkQOsc9QQwzoxmRy
bBgQ6K00yrfni7tQHdKfdm2L4eS8KRPYx2HMXApuKLgFem3x5k+lwOgbXQcJzTev
JI4o+OwudBJQQa+SOuxqUYiT5tMC4ncQji4W0xIKlm0XZeC1W8L2tmwBnU/awp5y
0g4XySOGmIcDddXMeDML67ZRRVDfTjTOljgnYDoC1excpR6bubGCLDxQSQwEP9Uw
swsN8rIiPjx5Umdy9qY/czdwR1qgAX5LfDDaO/uPYMXJrMWxH7KEgxH2u/iWQmh0
GU8Hh5K9i3Oyh4ehIR2zYjN6jug3sWvjl0RurQ5gWtGkU/HqhtQ+DVP6v4XikkYZ
9aZfB1tG/Rod8GdCFGNVwSTOjzKwZbWSJuKlhnvWGYisrzMsvvDLRZhaiZivjfHI
CDw20xKBIzLSTf0D2sPmhctWi13ebcCsFgvIOqESFZq5eAaR/PZrf9jM50Xf9zPp
jlXvVyfOCD+73vQLxRkt6Ei4ITopkZA1FBoxUKco7lL7M1ms4tjY2/pFzMpdHP9q
GolIDFJkurRtqMSv9lBC3vNM7ic2lGB8eI0o5BNycEOOpyGO10wZ9JQjPZT+aJfS
EGZ0ScmUfmtqJE/kL8VOL8TR/OieAwCdDIbZNQCmRhlcoK7SvpKxc3gval08VWw+
gQytAUMQHbmnxFg321EcHUpENOnFQ0/+eAQlOu+1OsA2CMlkvgrvK7wxiUGpl6Wd
rf5pRSUv5z/vG2yDMjTZGKPrt5sx/vaAdDsANBfO5u48A25/jOx778bW+rb+RHdU
GK/wREwnmFnOG+Jz6z+GSkGa6aPFrQwMhTeKc7/9hip0S5x/JxZYiwG1Kop38mI2
2V7K9Xa82IOIsAgUxJDPU8gnx8cKSamluuJZdmo95g9xGFXtWICBRAuNra6LtDp3
N0mD7A0prgt+qjcsnKRArXtaVFyIZEFjC0UhKhnOgxM+6OCerV6euW5uyuH7CLi2
WLx6AiGcOy5jdnEAJhBFQhPkNpGY4gniG0I2oIOZhwo=
`protect END_PROTECTED
