`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sF0usUs8uywUtxNJ6kZTg6nDnWEIOFik6seaVY1+sC+mFAkuAOhJFGhjULkplKpr
ZZq3U/djvI8tyoJDtaAnz+AASPaR+QRIsNT9rlsLjq7ID/wyf33cYIQgUOI7+Acr
g1IBrj4dX4/c2s+r7LG2pdBMMRUgTi7mbjyBd242xw73FkYknmaRglNu9857yQwK
TVLe99lzeDsXUu2GWvJ+IIFaEd3YwrXTv005tBAVaXVIXuPQzpfhax2LKTt614/8
1IboJjQwIApLYZZBZ5rizhj8z20nnSdaGeWBybj5cbC5cxlMOcNrzgbL4x/8RcV2
W5qd3YbliuICxwoMhfrvJrv9rzkJPt9cONwnBLCETgoJaWotlNT0I6rXpU6+AbJg
dRA7+7te61sTO2Uo6sTfieDfABwE1q5CgvilVXSksLdLloqY+6JA7oI1E37fFTeO
lHNFHdO3W4H788dCkrDB8pSfk1vUF5/W+iPDPAXjKMST9Tb0I5So2lIbQkypMaTP
TLF/qNumQcTlMqGCI+UjKb1PyF/f7ifu7nJnkSCUx/3DUZ9oD0E0+/FaUByn4d/7
FLwxBhWriW3otq44w0GnZZ63SK8yC2MbU8eLFZdt94MT/PX+JPvGlv4yq9lQRSLj
4HcVvcsrJNCw4UJy5ZyLgV5LrjnC9yO4dtyoJs97GJDQ943YZn1aV0fjrWyZBwsQ
xBeaFl4jBvB6biDbL83jwAcj2qiVYKaLs2TJ2aMgbgjgEE2BavdEAOzSm/jKOXQB
ggioKqtHe8PU7T2okG3Pd8KM4HPfvK/pR3YHi7GPyawhhcGM/Qz/7aqyti4kfL62
xq+t5uKdxFA5WEFkC+yRA0QwExohGMbdi+aXbKdvAPSaoYpxFeygqmni7tzTX9AJ
zgnTZalaFq5vA9yAZMod6/3MSgzAPjHQkiD2FVsJnMBTWHHpjAceW0SK13A65bYl
NQO6vAyifWpUvw3tv2PoaQDuiGP//5o+VEvNckfdpvd39CuId+wZD+tX1jhJeZa9
6lSMwkDKOcfi6NgkyOcjGH7Q5eNZnJdOXXPQqRv0M5MlNee3xti6juEn6flaM4uL
7sYsr1cooE/IQfH/SMZEXxYT8OWdsX0vquYFRbUpupF/bbwn9h9Sn8w5anSRAGLG
5S6jjyN42jUbVOotgjZexl2XuRhxlYUeLLYjHZXNeWEFaD0ziHe9jkTATT9YxgMP
yvQqM/82ghZlD9lFeqAjf7hD+5CesLnY8TH9qQ3NT5t9cp9AxqzgJY/fnzo+xbWu
uaWbNy8CeEVglMhN2gLqwfcXJCL4wwwOj1M2UCVZnirPmB9MVQrRMy0ctNLb7vzg
cWeL/6kFsEJz/c5MJysWLh+xjvMTmowi/0bMb9QILWM7fR61GpA+5wVhU3p+mqID
PGcfFQ3OE/HgbeRLcPNtKmKo+A/Ph4rNFCDfDkyzmVitF5NtVEo+7B4f67Y/Qpt3
NYVv+u+wErHkOPY96pmfDg==
`protect END_PROTECTED
