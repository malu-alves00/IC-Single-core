`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
brQ3eHdSphx9vlRUkdZW6/Wke/x3Pz1YuCLB39Ir+wwEQQIvZjCoKcAD9zCqtSls
BKvitlaBfji24pPd/QWGYVbaux3S3F+KHTcwr3VvUG2dV50Y/udLxaNPEb+H1dDi
3UuwRVIpVQE5Ea6+WigPM8iKDQh6cM5lH0u6hc1ESzLejjtBEhwqiY/zlMJlGiia
YXvCzURL060gKWY82irdlUh+fUuVeYoLbPPVPDErnuoZRius0fNC7yjymlxqkj5X
tlbNgsyqM/J7x3Gz0HQG6SdIj32Ps+YKxB0ru0I8oDsPYsy93JdfH+2FsxP3Lb8b
wuzzIeGGufJu3nveNu5+n0hJhT5SX4NelRoSp/f2kcAdzcA2rRz6fjEiAb+tPnAX
utVK/95iGNykFJhQxIkCyJ1IAhhR5/gZSlpYmFjxf/3cC3HorbpnxDM+vioKQe2G
EBz13eCtl7xPNaO5KcZtq+VoGZddTbfKebH5hHa0ipPhq2y7YQitrBS2S1BtL0lp
Nul3N3EBSc2tdH1SavoO6Fx+7AjOd9W3UYVBOsguNbAJPzxtOZZFOfENKM63yryl
kx+F3ZMkAy1vJKylrYK5C09kOium3B1OogQEBUV8UieW4QFV/q4IwpgGjiTQWGY7
FlGJ4UhA6wFhFcz5ZzHYBomW1+ADwDNYnRKnC0M1UdFSUKHY7/egawNbuovTT4M0
4/Df4tkSNdBXSCzFV/A1/MXw8klJA8TmlHcESdo/yWEYb+nAC4JXj3XO5YFCUXB+
j37gWfwm9JWOIp+TyNkXUvOjNchmBK4PJsF/A66My94l42wRttKPXssjfBTdvNxb
xxIx2vF7wyaaERfE/0T1t8GmgvYs3GRogex+pjXffC233UpTQy/e5YjOIlbvfG1/
ZvNPgTtqBHcNOdi620MktzEmDqR2O19mebHjt9k38SNpGCmYr362qVWUMND4kmBr
k0Yd8KXY9AM5vp9OSSHMVLdRRAXB0hbcwqSdgvs+roaYfgEcJ9SDNgILNOuusfXu
+G8VVIVKMCPJVQWLtu0WTBr1ATi+Vl/hHRhIAByOf1iZ8/fdN53XSJ5LW1HEz+2X
O5WWdeuDW2DtZJPN/PmvrUmQ15HJZuqKe2yk6Pb49EiRJszNJA1fY8y/uTlpxA0j
UgQx8/RvSIXu8eVPVmIm/AWpYyMvJ6FeEztntSm47BntirGddny3Eiv9N0ufcj+L
LClkameFilUeZn2UWV7jan7sJ8scXOei+aP5jPE4SiQ=
`protect END_PROTECTED
