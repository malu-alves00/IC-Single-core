`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DNmGIfV2813cEqX/PPtq5Oodzeks3/eYDpPdsj7hAM3mQ7f8FqRIb3oNLOTqO5rq
5RWS3O2+bKjrQS/x+5JXaLj5rLHpg5Dxxxyjgb6zyKlgKZ1KJacDc6SJiH51ymA3
r3IY2QSCrdgz0oAFqchbkTM5vFoG1/PLAPvvNy3VzMJpFto80ZlU3P3jBhOS5YyU
PC6Et3zTYPCWdj8mRYfU8IoSuKNxvXjwomdfY0JIGKlTSM6Byoo/eBZK00RKbk9G
JpHwvtF9WQ0pNsnBoazMcfQSJdcLB+yHuK/gczohhcErErUnzDmIp4lzIwNuZC5w
hTs8kI3a04y9uYbsZibcMpGYbAPSYd/OrFl0Wja73r8iIcpEhDkqTxx4u9JY+FGo
vpP9iFEAueiimEVj4iS4SbTnyXWO6WRZmO0IaDerYpFGxndPSk67JGiB5Q0bu7qq
jwdeQPQ0AGAOT/tbkR6Mf272ZqyFSh9zeESaG9NAGVqIMCz03/u2a+3i1gkJQKHn
Tc6NuT+Lr9IfGYooVM3QKg==
`protect END_PROTECTED
