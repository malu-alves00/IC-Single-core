`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kXMHUsoVrHJJVQhtpPT1BspMV/B/5YV2TjaEvdkKVFierEZqANCHLx0k0AuMM7Bx
TNOqXUe04dkczMleLUoe1Sxcde5aYz9mD5cwbQEJJZg1g63uUBDx5OHqNwXhSn2F
3btFX4SY3fWo5lUjHYaedpRXjiXfgf8zfxwn8LksJC9++2r1a2fFfyTX5clTlPJn
5sf7mcnIDSQCUsVxku0HjpGWXAAM/xlkKpsUYdfdtHTmCKTzxkMPrk6QwmZ+sKwS
qJW7kFY12cHy6IU9cqVj/758nSzfva4Gy8X3r60PEitm2ZmCNh3rSoEQMRTYNtLT
qZMmQcCnGBBeHNvcPwaqH2EcAWP3gZqC5DQWSIsUlgxe8OXGzreZOIoThXnGUDZC
HGEAMteKSkts1gfM+al+zT29Sac27vkgYwKyMSq768I4cjt8VD8f61ES7ORpcqr4
sGg1FXOFlNAnAEnPMJD2wS+I0N+mUSkxk+mRAJec69HwD+WpV61BiXoOSoJW/ejy
5hFIzQme3g0Ri1PbAwRjlEIuQh0z/ZHzrSWIAB5giUKqpprkwf2nZJZbrofSRpEP
kikQMcd5gSRiPG7se+XVQBdC0h87uhds2bYkEsbQ5VvN7qsLelEbRr86mlgNTJOC
NMjBVq7WuSLcz+vYvyoK/tj3YjoX7Dk1JVKGkW00tWbYBm1dc7KrQhNd1d2fEgQY
2r+mEBtWGbsnCTvsfFG1JqOfblAlChdbd6e1PeRsWa+mYOx+B91s3wFSPwY9fB7O
5baLph/AoAJCXuYTiOcFU9HYzKhqf3rFnhWR9YtKzlb9D2x5WFoNB1bD/X3QNafa
WhtxCqUDQP8AR4x26Oa6b+AOzZ1dsTcIwAWcZaBFxY1PYL4EDw8nSj02KB+MJWgf
8sv5oGeIE3iwr1wijEmeBfnKbpgo4bekOpy3C4xcmF9AhqEmoAnFj5yA74khIotQ
MveCloDdMOxXeert2IPmG+G2YNgS7UB2SyhkBZMdnBlmxkE0ogzibEJw+NZET2fd
hFq0NCuEDFIRAU4FSl/FDXRe/wYnXby2mZhtcatSeUDEm/rkI5e8emlWFgHrYkjV
TwqqbYik8Bm8FasfA+sJcvyfYbU/XiJbf0nlHzOmBmsM7mTFXo0RWca4yzr01ShX
A6MAxHMkYSMtM36q2yUFk/7GrjbEN8UQL1yhs0qgmwlD/4djFQ1nIwmMvoRhSoJi
Yt4nQVrRSndfL4EvpT6gJeO0A7WFmobcqsXplf3LcIxoXoJN1raO3X8x5qdwl944
iXHht02J4d4Eco5QQ03jBqiUOlYj/1wj6h80fx0kKeAfbFD+sv6jk6/wl0BsXakA
T/4zi65//n7FIuRXhhJ1Qd4DLHd/CySste//s86QCyGTKIf4Lp0DlTM8KCfTbrqX
kXUecEUPUxEHWKX9Fr903RL3CsIr4UyYwhJHY6hNnRJGhUCA2MIv/P29iS7nyR+h
9qHYRhHBGEiQgEFX5QoisMyjeTrThokExIOGJI/qGs7y5XE4TqXqHOVgvdJDpKSx
q275JSH9AGnXuSOqgN25udVp15DFruGKZdzEK7uc0UVFuhBNDGPauntwk45qqs4L
C1jd/5Mlo4PPYnth8kUFIhtBnnXYsfot2wtWliBrIBGFCMydosGj7mJJganOuAZL
hzzw2uTRpM4Vf5EB4qd1RB4yT0T0yUMrW9WlsEF0FNNOY7pUKmzOGcpWUfLVdpRj
+CNHv+e04AeRxBFvzh6tdx5QFlyXr36hGgxuzlMIteRHypx4yhiIWYUtUfeL1ifQ
Mr2ug4gA9yyszkeM5+hOtY2GNk6rPEcTGaRHgeGPZGku+t3PtV0RV7vhbMqshDrh
Y+jcG2YkSGhlsvNu3WWqWwJyIofU+JoDJBaE9q9T2ozL8OT1ja941QUN8E2h+u1/
ySYS+Qrbmh7qxEn/s0RvL1EQp90K0YsjRl1UpsuheGJJH/Bbxd+IYGHDgaClnEWi
H1x29dvriGnJgZTBMQEOB7JiBeuSpFz9z+Ttf5+lanBuZGz1bHFFucvGuY+OINUL
+YqIJVhlQral7989l6APoYxMlNgKWVeU7WfnNABANrOYd7EwUhX+CT/SrkPN8OLF
FqVWtuZL1dq73xhUzEzacEebkK5ZSzpr/7fPHfmpKhdWfuOHQENfjZuZwUlVzf2A
4LqRX83aL91NUiyHWy1yE/XQXmcj+AMUVQqKVR3lT1MDzhEtD/maA/3EqDh+QSx6
jcJ0DjNvjrX1Z8Fs7HU91Zp/0UweRXRGshIHRSZIDMRUZPYirYz83vq2wzdl1U9i
vLcfbN1YcxpAE0VKJVJUvi3KQ2/b6ZVB0sE8nH+nT5wC0Wxm7AJ47Wtc9GhR6b6C
CLVL7IfmrD6JKzEaU5RTDCIMeOScPpF2QmCS0r5pXEZINN5T0JWzqCvezHaviJmh
9Av4SazJ8/fUmTLvSVRVVQCgkXLTzskqK/bAY6TXGwpdTPrJ7wj2ETigVeeRHNNn
rbtxlxCCmYItvwgXWoX+GqvQd3p5N6Vn7bQU6UTDV55tvFFVzV0chgEGO4pr3Rx8
byWPpOY1XMgg8rdTSpJQnQ2BYHzcQU1gX7N/goxY2zBXwRe/FFH1Pi2mKhxWl7D2
n32Coc57IxbDblZP6ARMSpKuwJMPtqM4rPXBScyR3Fc1beOMg54hQ6xieL94fLxP
Z+dmxyXaFZahG12YWETVKe6iJJCFdqeKbFD7cBxl970GRUVXwAiw8P7GeGxFek5k
FcZB+wcya8lz9A6AKsVI37QHaHjdejqOBHmCYDnUPh5SzhIUKQtYCtGIr/TA3Xwr
CTmctWLHvzrpgigzflE6WWunBVK4nXrDuWiKT/nvkIXxnrlnWwsucHWPqdjzJH5e
qovLwY6gxHnEDurdumuEZ2CeRrl2WDcUu6jjTXfX+Uo4VlOhFK9U6vhtmsql9w5A
78j2KbY0Ye23QPtvgdH3AT6SYkZwoGMhvdmBfNDE1pRrQVcX4OjakxHGP6jpoOCb
aw80eQYY4mHr/czyp/J1p8FfsnvEhJGGgFKceDDvCO7yQGwnnd+9qTkHdnp8P28j
PAdtEEU7Q7Qf3QhwXwcCSGO4X327HuX6zHRq4UA/CG0lxzLWE7hkxS6ItVrEIwHl
eeX1odKZLyG5Ktx/MwNFigqUH9D1DZt48Nmx1L040AhZS71Mb4w63whUZYXrvqhq
/XcY78zi8dT5zW/RfOMninCIerGENUIsbmSANFSWewWLCSEwUuF08jp1BkupdpKH
/84cXh8q0wApoT5UO7KBZGYVZ9e1cF1JPMq2cEklLvgzfYRYMEaxMNuyzzdfDEgg
T8ydvl7ynRBxXs7gbS8XIYWQNSPibxsTkJDnBz4jjj82D+DchAcmGlepJWwCaBvJ
t5x3HKtYDzGxFBwZfnuuBES5QSDzDmatlcRIwJRuSEbwuWErSuZmFpMlhFS3ntGP
geR9Fe/Ggq0bGnGkHc05kFjeaYF67yDD4P08+rYQvOQ4iM0IzLDOFONg8442GTEt
TKVzKR6K+8YKvw5OQ8hNlMUv/RSbpEkYTIwBMuOU22dZ9xQ+9/pnFTPHla+8ZyPL
x3vpIp0y3g0RPRdxkuB231pFKNbogKXMMJ3iVvBN+XS4hGTLW6zTIERq7NULE25v
E9K6ylt7Zb25f0g7IZfYpfeB3N1A/sz3UII1MCKBvTOsieDwaUi/ugNcXSFxCCHT
Ge1+/n1ro90keyi8DW4BbCVt3mJuZOQF+VINjrQcmZX9f33z/3FCbv6E888BGqsN
IxkZKgiD1aphodXrd3XfeY/Utp0oLdEZN8X2VATLvDMqLEmx3XdSl3Ti+TUQoMrF
AtXIRzAPuoogJ2O1KsXWEOC0ScIGMw8gFOJJ6Hc+IOpGT2jCx6HqHw5tL0GguRP5
+iKeAo6kFS5gjW0gRlgF9R7klnAMnMT+AJs5VJQLZgW8HNKHk1CltgTR+n8F02KG
aNruWh/G8qyZgiXLNBI4AwB6c0sJN39eCT2nwn+brw3DZQsO3ld6BoOAq0eSPOZh
TePLfUvFgfNS/CT20tG1vJnjb61yvqQmCihYDQfkHG9IArl+g1MrxdMxa3x4ipYD
o11i59cfKikLs3gimIniyaQMpWi5isDMgaeTnfqiFBauVeqBuqewEG3ZSJXYQ3uR
AGqcJv+tIx0KPQj851DKinUIuibPB+5MBRB2K6epe7Wtj9ew1/uoPMdCwL8dHHUl
hDjMARiZi5vHwnnRM5g4/4XXGNzWcNjQXblbXOehiBFFrOd3x3tdLT/2U48F9DNb
QgwUciAH6BTVDK65pzwsJrdGms4jaOZXvHtbTkbLhnswiCnOJADfVV1Ns/f99Hso
V2SuGYNUYEZcYqWURWhK6yk7T9hHLnirXLzshALEsJ88GpOZVUNbYDnNnLeoPUFl
gsQx7ImiygYeM69XmwDVeid3XF8gF6IHnyENizG9yOx+LUfHxZBcHjz//p+ans81
5h5Yaqx8bcoJgMkyPqoZMhzU8HT3XuiORRZSStJ+eTFnHwQzcBQWIJdxGad15gag
dLnZ03jQfmXW6H9OkH8uk9cvP+SUQwo9nzEUAaurqtNZzgso4Aho0LSBKaQBR94B
89sWcywGv49Z/kHFvZpTitGDBcKhU1WUM2mIZrMr8uLj7Dd7BT0vMyNN4FVsQa4M
gP5F7Uh3kBY5K3mT0jzL54R6fNkmnliCRLrI3WJCIY2NTiqP18ZPCIG/MWdslyOb
/aVBpHN2IYQNVxc8tAyZsZrrE7BvJgnhMZR89a+bra3TgQvNHpAUWyNCX/AqIHke
`protect END_PROTECTED
