`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yecW225sHEKTSxKa6vTZkvyzTd2Cc9N5fUMI9xLYFIUBAMzn3gTQlgmiL1vZqLwp
UcE5CGOeDiQueOKhFdA1nQtH/2mj8m6FLAtD4HZbiVCOHgIi/vBR7Ek1KbqSjBvz
x9k/86PD4AGmsayyQWhdLJvpvvOmMl2pgoeKouxJ/ZXkRR4UV2qoNO4XNyJmn2/W
JIpDPLs46eEkj6+mm2ikwMBjONZ+05c3cKeAUpPb1hgp2mtjxpUu2GnHTmhHNLgZ
Kpook+O4EfABnJiXntSAMUuMPB41l0V/6W2mVYd+dDWFeSZLR9OColcjMm3WHHZD
uUk6AtghbbeG7fhdSoG9Va+TA9nhPsZzHOlbHJfsyWtQggwE3o/5P26Bq5T4rBYR
2NzM4Onk7Gcm+8Vc1Rk6aMSb7fx0QDKxEOQfi9mVDHi73zh7cHkSZaue623zTsPb
FSoSvlsWiFHEq154uoWjS9mrM2vYg4up8bH+eYtnlvGVqDz8VcQloZ2yRu7jGQCZ
x/nWhEy+pHYioB5gXWpFp80kJU0c/pAc7AW1F+ybnFPsF4GxUAtv/mNRkh1RiYF9
dlH/tT+EAk6k93ZT2JDRRQSdXF1/ygfmigT3pTJb0wvFFW4UEsrfD95lzW4iaCMe
x7oWI4R3OgxlLmBLfINSPib5l+2hTQZ2hIKhEd5+uKHeq+7sPW52TwDeSZLg5CJ3
4CfhCx4T8HnGgBSQFCDuR8uXXQwnYDZsIO+wAHLJy43m9z34ZUEhw9RDs4jFyfAt
7nZHDWoYF/4oFHNkL8v3rp+FVIF6g+R7QRVrV1bhmpq3MeQn/aNBWBCys/XtJbWy
V5/Gl4V5hsG7oOE6OPYTqnJ24/m7xag5fC4uhP1u4N5uHZZwyNWm1nr+gNCupw8B
lzrZXqUxQHIjd1pyoA6oEtZVCEc4nmxAkrVn2iCTrcKnWesEnTZhXCZ5kJ/UA3Q1
`protect END_PROTECTED
