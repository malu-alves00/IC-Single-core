`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
i5EnqelpOPODOnxlmrNNEaeTEgPuWm023oeyhedzlmVPfY5zSF9XiVn7T4tqpXo6
016Zhzd/1SSqr40vxRCjT3dTLEhVEqjf4OFbGnk7L+Ou7QUbBw2W4M3YzEiEXeT+
2YpZFppxfnJ4TX6t0uIFxux2Z7nFs3wK+1qRJCL8GAyTQDpzGIxo1w16+/Gj9aMz
MWYSITHlBjS4QhpjmyUYKB2ZCYWkt+0tEKPomqouy6HJb/IE/uUJw2MEhXnAyPTL
GQFgwNSKKBOmj8VNZAhQpeKpHkzyU30q7SqhGqGc7E5tU465genMdp1odF3xo1PO
pXlx1KfIggHtC1UzwAqA5jlz0wDnSqC1kpKomnqFUnv8O7I5w9umjLTBMlFZaIF4
yx1PK2cFEBK2ks1FwPrP8GCf+vWj4tRva/ocXpyt5cbCQxXxkrwKfNFHPdSoA79u
qU5Caqq7EnF2/4xH22qDt5zu1zXy+7oLhpg8tfsApjtybcZst3q2HqIWUw9/A2jI
H6JduNjAxEV1gQMvxUgU30+tNYt9Keh4cH3fyCFq333WPYJx7fUbkFBFhKqrPuiH
mdibqLDpQTCYWu6S+9LZnMWLDpd8IXVlQzB+jfSCcqNaWfNlhlDWfJw/vnJ/dUlS
BF9SjkTl7nbI5/4b087rm4q+xEuCdqsO98WN60NL6SMA5i6n98YlMhKpXyZuPt/1
2p0sx3BsX5w1LZdLeHjkSLgk00bMnq7Xj2ZOzGmWL7Jg3JkrHRDKON6ULe4z1LS3
pNWOtIod1HFLVWIVDyXgJ+sOL3IpI8aIv4cp138HKUka8ouMhtgjaTz9PkUCbSIK
IUGac68bC5JnEc77fWwSg0EsFrtHommRIazg0XTg0Jn6xuBme1yg7Zwx+M3JdowY
Pzcn8tCC86HrIyzBqTUFt34qQuoOIrXc6Q7Awlx5VdwrTExIAj1U0BqLb650aexu
igJAqAH/hy5HCtFAThI6f4FK45yXjJtuAmLGlbLP7jRbk7oX0j5u8+O3bJnlo4ky
XAgM7ohzyPbZ4ibxHQRhCgXWcupPra4uZyyjYLLbFfE9edXIozHpYjdc+PUWDe1O
A93deUsjWqjUcAxknlQwgb6oFU/MMHCL7UTiIXs1zNF2sqUEym9e4vXW+H3KHtQ9
P5RAvVImhl+nYKDIoq2DXgbSDweybtAzZPAgjyhOb6/oQJWL/FxWBZpd58LHzVUi
vT4UBG0qhwlFRm6A50cPbA==
`protect END_PROTECTED
