`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CLLTS4yBya0Ax+XoXV4doCsjey/wTKypuIK0MeFLBpQJAntqdyKtiAMD5+VJ/CMh
lsgmPtQbHOv9cwW4VBjBQXLL3Eq/CdtbJ7zUXG704LpHuH7pojdcD7VvNDVgUF3K
pbwUuackqBldqpnC5cOkCzZbdZZarBXD0zHMiwAbnHPQLonMBTcBzcFKWg/nRuzo
Snnawyep5BX3x23uxNnN1uo5dHh3+FCG872Ins9+9R9w3NdtJQ8LyvY0aI8C9LoZ
v1qKFSH0huTsE+HMCJsbgG7ifzCrS2NDHXRB99sIKigN3DIXZNYj9+Ef7sl3GLRH
iahX6ugu2untrSAzPITYJAOi13G1t6WJw91k6d1uWZF/KKkRkYUidECmtbJBEAqL
`protect END_PROTECTED
