`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
huf+KrSKYKnfvqZNYJrl5KKxQyn8IaTGcYo3mW2dnplby3fAYpCfx6ESkb1r5a2L
EhEgUZgVc9Vv2P7Trt8qPdWnC+rVYgG1/38iXZzTGO4JXBZjK80ey4SQc+Vx1A2z
QAb2DiQ2EjxlmMKw4iKDN6m4ykFLbxeSStNvkxXCAXaSbzuVaDBKLJiNVEoSE7yL
I8Jxa4ynQArOVHYlIenb3tD5i303EzmCdW5f+2NLIY8rv6I9yn3lA5aHRNYO70q3
qBo2TFkK3zvCEWTFZLHNOJz5hYWi3OcRVeQ/AwqJO5xSr7EmrqJko/nPd29Qye+K
ty7IsURWiWaXLkHJqyBm9hI/kclDembTYQYy1LFE0LXBk71WpTIGeqve7gmSPyH4
v6HGrAu2nfT9sCMNd3DrrQG3MwxUhFDl3sWtMcEUvI4ctFbxaTJ2LjhW5ex8Hp34
PXW/ZXRYC3A9pds5KA9+geYN+zVWtTTcoNi1obkdODS4TNe/3yG4dgGApcJNoTBs
ysXA6yFNAvt+3NoGBmAiVSHuqY1azlKKcuUG53vK6JU1BxbAR5uRRTD5C1kpJzIT
kjSVLGvzrEi2VjrRsjRTs/XIEqwdM1iIMsm3Lspi0NzOTMGawLZOelRYtddri7DX
HV8aNi8yuRCpjowEUIShbzAdyr+kVTVlsXT+GnJkRKc9Ke0RLBAKP2qZ4ziXh76D
8GB9dRykUr46fA2afikQzlAMjiki8cLtI8B8zsd+xVVanPt4CMTe8z/EH00ug3U3
qeWmRV0CMeeBmd7dfju6C/HiJCqrVrJd7ju2qS9EFnN7r5R9D4PfiVGTt5KvInzx
7JI3+7RhopDL5TQWnq64uI4JP++T4T4puP2tZuLCHTi2GzO6Z/2IA/pmRyaWANXq
6F6VtsioOJm/7UfDI8rmM3VViwLf0S04fIjGr/mVrq14SHov3e9cZxLXh36tqiMA
sCfFyry3IMjI6BZO+hEeGy0oZKnSvVtQixG/k394DU85A62UNOmxMrSkRCl7iTZP
aafdWbCAmhV7Ok4TJJ4rmUv1huQFIbOPfBuVDdk7P8Oe/WaR3nsF082ad6IfOTVJ
fNtWtPQgvoBltE6M9CT5sdL76VoFUSDdE/aVBek49LO2IV9aL8zTPv/R3tbW7LGh
R1pHGMDoSQgDxl9HLe81zdlM9PBdc/AM587XmKLt7m8ckTiLuibQt27B3/GFnStg
thlXfKHBiF7BiHMmqKar5SaKPWMOvr5MqcNgBlT0BI1KJRoJphbku4H8Msa8tnew
Am8ZaRvT3gXTf0ZEqlam1ku89cffQATHxDQMD1LjUTxc+Cp6KmH/DcfJ0qL6ILOw
6MBcnPcN6utFvUxI3u50M+tssxqRRvs/j4rdHybwMDqoMvJ11Zx6wM+ajhpErxB3
MT9JqHAfy69pMISYBFEYAZ8CV0rjIXf9ibOpFzb5/qbZIqjUT/IsFpdcv9bEn2cW
1mLRS8uBJtNCDauWWKYtkftTpM3XUdUSkP4MVliyXxo1LocBy/jE73J5icTT4bO5
ERh46NRvhL0w0QAQTqph0rfFAKXVuaeWlv06TKb2Q3VE3041bCgeAtEqYtZSnKis
E45JtWcVRKEaFpsvw86AI6YookI9lTQ7NGS+WqEuNHd13Z8ajcYnN6CIRrys8YR5
5aoLN9P9DqEfV2i3fmzuvfyKKCVXFj99GY4qzqDI89rBy9eoHqlgHfsLtrlQ1uuv
4f1BlH+d8Ynur6dRz14LCUyNngm4XROwjpxOdRwuRmK15ArJfnKPH246gXHa5eye
VfM0vd82McJ+JX5Mvsx5o/sZy21ByCpiDIQdqHN8AmhMVjUUD0Yw2It9qGimdn9z
7Mxgl7eI+EM2rRDGpOFYoWm/0tz9vuk32SuzBYddZnyaIW/nyXJgg1eUmvq9mNuh
3CAWXfSnXFP/cCeRN9V7o2cOegYN0LEIlLMEcMLUJSvFEGykBDhgLLyW1BkllUDa
/lYP3fJWIb6RTTf0VN6jwEXfiEx3kFlWpPTyNB78Bg2FXzGwZtKfiZ3DoMNyQRrn
0AlUPTnTyBYFKbpuZ/oq8Cu30OZZfT8wqy4cJNSmPLf3rJwsy6n3MfH39wJVcGQT
ImR9ta+ZgOxDmD7Kyzo2/0dR0zK7FAMSWFsA9iMExbCOVefHFuuLTb3h/NuFvca1
ts0uvyR5x5jEPhgIHYZLAHT3SPId2C26uNQKvnOsXpRSFNdD1g1EBfd5nphCJJ6l
lhrClPJVMBjo2n6dirQgTVMpY9uRYYRHndsTA33Z1yfCeo5YOC+L1nt7x8EZMfW4
tKBbUnujqQqRbl7gJ3NWKKEIyQIbyUXqMkqK/z7R3iVvYWwxBqhMOwSl9lodFfFI
7+VIbznV6Zm+Pth9Vj3FyB+ChwiZnWjMvF4jBaoxW9M7YevUa8WdDQlyrXH4rNRT
bCeTMQNQ/Tu4KvBZofIsBCu9KbcUvUoBZsGGUDYoxqzgitlCG/sS8lrNL8oOHrCt
U+0uUSodp/l9RxSG21dmNFxwfLGfvMDZuzTFnPQMi7TTmjvcRltBDuV+crVtGLyb
vPlAByZf/s1uk8Z4SSnqY22/+YwgOE3uuhuZVnOOxG0KAOhP1uEUEkje7a/ewr8t
Nw4U3ErG3APuxO6aKJkqGGu5VPykLQLYh7OGGDJVR6cHzXj+6NPApmnb72XWhntZ
oZk6KBdq2BS8uwB67YR2HueYXFHMFwl5Wd9h1rLByOy6qWM1VhAjOjZXgxDzMKL0
it06BGwqUxltSQ3H6BK0F55KdmDsCgojwIiD3/noprx/Am4BNkVuUKekMhdoZCK6
CoUpvCeH1+5fjayRsQB8EoXOPMH5T2NmY7jeGhr7h6BmQuHTOWonTrubidkoA2Ew
zrNh5WLPoNo2M1iw9G/kNhCke13PnJOO5bIesPqrWyQi8TlHBxUsLw9aHw9jTKXt
2JdT73G468N9gg6cxCByS4L0zSLNoJICFjcssrDUtqHZLEfm/5/OE/fbW2D6yhnS
Za7vSV4+p7iOTYHsXahWbXRI6UBBxRfF+cDZIHzdGkEW6b6nSFXa+2rWHsuW26yw
UUYTfvJeDTgcUf9S4YeNT49lTSyyIunfrVblZg4cJap4YNmKycgXl3Y+9QbVB5Wv
l753qKrip6Cdw0a2kwhMLl0oftQTN73MU+laOO6qeALtgp830UAGUQo1LgyrmPQC
50nHWeHyETbUyeDr08mU/Ixnn7vhxMTCsxQPxheE05bC0iVddRu1aALsDymWetmv
0TTxyTIQNjX2DacHXTAFvwtRt/iu8ApgydNSwPPyFJUWNQqiz9bOn3jo/N+ecwjT
4a9lzUtKeGQZPiVmENmHJDiDcuWwRKX5NjE6jgvBt3/krsBlGufuNWpbGihbmMWB
GNingry4CBlq0dcR9U3Ye6gKKs54iMFjJfuLPm8coBhGmSVNAN+lg0kbphRPktSu
wrt8kIyjzHee51Ol0HDs6i74ouvKy0iQ2F+GtMYiT4f66y2bPSD/QLSi0MwPF0kw
RNoXQEtV8Iy6ICUTvDPFJ6onXtZBJAODRjxoXjnIcp8oKh+RrJ+8oFcEr3O78spY
SPzTKjSVpNi8b2Ka+249qvk2Zvn3rHoBVsniAlR2Pho4KOafFRtFkZwi8XDNTLgh
6ThKX6RGj59Zyy3W8LGMjlPWUBV4E4E47VwYUmXeNtwc4mFyT1oZ+uumUttwrV4x
GgvsuNisE/VLV41U/07OvHKFjzo62GpnSJM7DdxAh1Cc7hc9VcihXM7iaw2+eY3g
G3jKXVGIs72tXy7OgLJZ+EufMT/C51u2d44oU2/pGY+DGrCEq4NUx8YFnBs1iYXq
bcF2zguLtTefvhJmxct+ycFzCeUZ6u9Z7hW6N3q9/e8jvkk383so0T8KMBhbvKKA
rzl5e3Rqp6GAMvZOKofduGCgbUxvHRdBeE1xPVtj8MjJhJJpguOIKv1p96zaFOnP
MDIjrSFLYcSWyUZQApoodeSRslbEZvF+PFyphskMj1Cko43KTKT7UAhQW53+FCSQ
MoRGe3CLlX/Dc2tA7nxHr8tk7UHJh+606AD9bN36hfkfBvxWZUAJ9GqiXBmQVfp2
FLBnOrinyLkc82hQGT0AroOzXnhaVFK9jTC9kAOqvFLbPFDXUpT94ZfoM5EaDK11
8V8BM7Q7k4hxXjUIF2NaXWN2tgeYVFoCOsXcZCcvE54ZGgxjkFB+zjtSu/kAtRU+
Yo6F0wexRbOtSkH0YNltZlYd1i0h2hrM7Hsp2a3w/ikYuC8NCsMVxv1ZWiXdrTBy
ZKP7q8G5MlcCUZjazwQ1Qlx2Ahsc1QiymJA4zhZjMpq76xbUuBCE9BJkVaMD33LD
6is9baUmxFjegJRo0xumyfvrrGq2r/341DHsj7/c0aWuusjPuajwhE6gnLdy9voI
1m7aIHJLYiBlxS/BLauafNB/OUitbSg2HIzZ9cXAzqgFSNc+m5bXKryV/3cFC9Xr
4P+/D/P1XfwmoyEFUsZp7SX3/AK3smFejGH5fhO7h65QXcT3xzUi3p1lQFRb4hAD
T8rD/F4iTFM3T855Brc0XXkjYjheLNqqc41ONkW1qhQhX48Q0dlFfZp/YKB+4O7D
XyPjkfQ+Wo1lZmcEGlOPzPJrWywil85ASyK6v8v2D30z6iTwBGkB9pHqjcqRhRvT
jSW0oZyb4I9AdYH/u5THiFLTbvw/6oxCY7iYwlqhSbeKJxdC6peYB6nFKLngDvpa
UhRyPtNb4cWPsBF3n9PvOe9YX5CmE+N/m8GBipa1Zs4y/fN7gXlTJdL8XaJnsGEp
sXTK3lkRfpSmMZWc0ZUcYCFdFw9840u2EwZt+9Xt/Zbgbuk95iL5r5qhrqopvRWr
1QiFdgndMCk3uX4lb8WYGWEWrFPraN67wO4d/dbo8K5jMt3cubxFROo4Xxor8kIn
qU/I3xGiZVNtqK0en9JAf1pWNwnw5UYIi1w/qdGXCsRlzTjOpIwjv3KtXkndCCI0
WfKD/QiQACMlFEg+6W0679P/M0E1cFQFRSy9U3treL0ACavJG/yKt36g5lHjg1cM
WqE4AImqBhUAxoabo+nVYoEQtNG0IhsePjhW8Pj3CnUxJMbzuN7K3stSUBRLr634
xzq7hsW4sp4/5oWFD1zhOx0DsvNyYteSLqTJKP02DJZHDhM7dTAqts4n136XUt6A
mY3f9zki1KozQKwD1UkFH4R/suQFuwZpa4Ghp51/CiPKDZRXFGV2rjcJHFEdkrHC
YOG0WGKHmXXjxAmlxZ7QFhJTRFZbBuNi6yyIli54GUx9Ek51z4CIAng6es/QMJ28
YUtZo9oFug+usZtF/HL6dThK0t3BPUTmLZDsM3jbD1QRRBAf7WLrPs38VMgofj/n
t33wxNRkF7rantyKnbyLfGfsy2cWgS6ex3ZLnXti7a7BqANjIrcyDlrEi6/+NAeb
onsc/VSmr77b5vh9wIpj1JFM2GBXFkl7PEnw4A+2etMJFGJ7JvS3xD+mekJ461ik
V6q6jBhmGdxk9OD3jpHXRYt77XOF3UPPybGE3/5dOc6yPaVdBfP89TfykSVuwdVz
9rKVJzauRJqZJIgYloI7/64YrjKzQA1NcNrlFLVaWZZnSdCnVRUIMHFuZzhWKrW3
VLxpMxDWtwE3UChjdwTeA4aPRbS/SkGHB09DKqq0pFrugN+MBfRJTiehvgcMxv2S
MTk4h3ALk2VLZscm9UL/g45a4pHud6uBXL46UeDlrwizzYtmzddFv/qdcOd5iMbM
1IZNzCERwiIAqSIdqE62eKtLlM9WLnrZvWzf8xVNtM6EMud7TOwu6HWkwuTqVppf
Q0zm3Z/5gVrU4P83rn/7/iHp9xREUoK5PBfPKEigXnIxu5dUEHQ5ZSAn3jaCXier
hONfeu61/R5hgyIL+O/GwONlmWnA/Z52iu5j0WL30fqe4u+GHV29P2BIgGwa/QsW
YnKPTuVFnGz1qWwOaKUv5VxSQFQep2fv+IorSB9jY/jjBPTTRIDBZ9pTK9bii2o/
HvIA2AmIysrocEjXMVth2n/ktAplVJp2Cf+f4C+EU/7ZkKOw1YHiMWDWDkGEFpOA
JRvzjWWRTKDdTapAlFJ60oY38JdWDSY3Fygm1iO+cUAF5B1if10x9MppBdGXUGn7
4ArtOeGmaS5vdS5NizM1xdtfnMWfiSiJtXxqz/8FEKZaVS+yXLzIojVvJF5136XJ
W0vUz1gCjIN+TcZUW98aMgEn/8gE5vYSsY6EzxSx2/CcWNPf58Z82G3R5RANEhRp
yAcrt6F4OIL97O/LhjbsTD8V9JpyTwft4+5M27gF6DKihoxindlJMyeWBu5XLBC4
fa9SUnE65VoMvZlKJ0Ms6Z9Wkyli37HFIZSqwNBArVBZdr7QhmrN8pmkLiEVqood
U/pikzX19D5wyNlqZBBZZcUuuyia6+K4D/+xyz7FCRY05sVynL9wNWwx0tWyzkha
R/VH5UPhy9il/x0/6MpZ/Hr64zTVtvaaJvoW2+lxWgdTkOBtQgES+JhdAEZxsmIe
to32iyfs/4DfTZUtiK7qOfuFOW4iPEcr/Ngj1p5Z6x2n9Wx8Hggs+eBmv7yCqE/Y
auuzBYs/CgRCrD5ulSEp3LfvPGsxdGlcAzno7kzBJ+qZBFy+MJrqULrWCm1SEXas
AObvtAgtLp7hPRVmOlQD7YtBW2EK5wQ891Bpiw9Sf6/C9cLT/Ks6kva6VMtolMBH
bjDY5cCNDFzEh32DkS6gCSak740HHmoDgkMAVTX0Zr0apILtM0jBPWit/9z//0Vu
2KgPxi/thhP5lsl5BbMWO0B5C5t25OlEFAlYVmrhm88/MeoUH6m5ta1FtGRjoKPL
7/OFWyBzh3QDhoMG9NqmqmsLQxtdhX1VuYjMvDb1l+Zc/g0AAIbG0ItW3cRLbzwT
38SKyqJU5tTDpFGnJFIH6TiE/XrEs7HdUp8E6eHj6SaVNA2rhrpCQFUiBTgzGeo8
TlzFfsrhP/Ze+eVDsDhB0vbtOMtkDSB/4i0qDI/fLBkBY21LrIufRQ8YGa3BzLTb
W1329lBJBcWXucQKkrL4s9ArlGPwhdiSIGCtNelvC/Hg8pkmC/0wY0nY6bQvmVTh
CZxRbZrSab16RxBXa2btgRTfLSHngKfkNrJtlx0C5HtrFuINMU3XZMSMWNGXhusz
lOxcwIEeWQ36AoXnBXpq8I/oB+PK+5wMMIlL1bZTI89VRN+lcGLf+PAFmjGsqHWE
gC2YlY+YR4K6gt3+uK43Wu/7fVi4n/Z+gPNaCA1GEqSmrgXhRzC3Uqnzxi2BMHzw
rsYDqZBCNEciXIe/dyRLAgVUkWwpx3jn8VzPUQivcno1OA8ndP4ko1g1x1o3aDM1
tnXAbk9eKEySRuJCB2S+CDV3nlpsluwGVKMYcz7QQmarSVs/MuHFDGF1VyJMQK50
gOJX/gv3bbt1TmpH4znbBjEB58ZBGZIcaCKkx+aUqjFQeYk6VqdXB3u8tNtDFz59
/bYoq07xPFCyNY0t9DpoEfeUPA7Hg1rf+qI+9wVgZ3cABLV74y7yFG/Gk2Jdjmkj
CuUK/Fu3PPElrBeWi4JK1foPoghHo1JHiOEXKpwGt+ockZygXYEC/hR1qhVSzzc0
Tv7xH6EQ321v1ThpvpaUBjBUjitJBmM5/I2LoqX4nkP7PCikY7zdePim35xeXFdq
sA0/oM/N0CFru3+yEV3dpEhEvURj+Axpz5Rdy60mEYnoGUCKmJFCFktGbHw6tzNR
KOjre47LplIBse38ts5+DK3h9TP0Ftcs0kKJJqytKG/JgRGs3FAKcLfR2KgWpr7F
G9tj/DKS1TdfIAkBC4t4QjCxvu9/nWJ3lu+tHgIIHWWDMB7Ls6jzUZv45VcMfzCP
sIw2rYSMPkX1YIynrP7WMkNrB0OIyP3fPfdQEKFuYflYrYOg7wRaUjixf3bEUZGY
RdzdAtmATpSB9s66w1e3o6xsCKmY/tKBJVaJznE/3u4RImJCoWGrdz+/QebGyYIx
vIKkXdFna7NOMGEaTslcueYcIt1dyJsGWJgD+GeOblrvmuZaAFF1bwvLGkAZBKjl
bQt+iezYFbEdvETgFo/9F3IqgBP9zO817l1/Xvcdd6JoXtghP2KgDU6nvxrUUwPN
qVyBXBSLAFfhAFYRFlU6Th3NTAt1Q7TfNW/7PBOdyHh7PSs/gDs0HGM0qIhYyHPs
7ys0WWDmb5MLADBJGOw6sZpt5c0jOqyW4lc7toHDRyX4kV+JR63NFpEWj8piFIaZ
8pe7g1eoJ5UmgSp2Uz/zeRphVBhwsOdSMhvLaEB2ickO4omwYEjJCGBUTUNKoB2/
rHIjYHJdSw+CQnP0fTksBqhbVZrT/SgBVfiEQNnD1i/sg9B2SM7bLPkftJ4A4tbO
6QVlHiLtLsDTapLUt6OZ737Y/twz4vhfpFmHdYgFFbbjmhUXK9grSpE84kDT+lNA
rcKoDF7GiEWXronHTEGLOwaCfAKvNTiReylbXqY4IHGhCnkCJSHaSrIKXfCl1Eql
aNLq8wOoxV04EmE5TacVD1fFAzgHFue5VW3s4Aj+pQ557Rc4TJzA1+2KOMei1LdI
CExVJ+1Y83BV0QLWJ07JHFL6oSL7YeFfg/hzKSmJfRqPA+WIayLP4mdb+KptInE4
mpv2AlzZvVthdFSH9fpMTL+H8RPBAqmg2RcM2E3GSV7VBez6t9yad7Zgy8kda+EA
exC1ZBZiJO3iNmQvNJBH6+7UPKw6EeFjaHood73iCTOL8W1kRYzTZPdq6+yerTHq
0n7FlozSPhZocE+1aie7z56P5bIb02lEHbYNxELH00TMQrkZog6OuOIUs5XR8/0Y
dPW91RTHlMBHoeu44pcVR3/5L/OBls9x/wi75aHgNLppSHmJYvApVPGqYZzw/nWW
Xd91Pbec3LBCQY7uzAEr/SVLzmNoMoSSUHRjvIaGPQnDw5cJia2ItlVttypRzty5
coX5WF/vPxXJYlrWevGd4OwKIjFpDPkGNhzKKC9nedygbXg0gSD+8R8y0HTTkdNO
HxakoR9mmOuIWrNP0dJz0KFhmh1wVSkXAVTYIkmsq5Av6vTytN8eT9JEebQ9Pla/
rR6S7xb89ubpNJ8FonG8u9wiSHFmwgtiH6p94vOQVkXVkDIk7ydy4XsnYu/rl1He
TbXOswowHkSunJdvgHyf82R/wX2RdVEZac6MdkeYIIgQttaES0hMzoL1kBxNR0TL
Vq0/RhZfx6l87oKCrX/lkiJt8uxvdfpSmwvywu9NtkP/J7Eve9g+F/KbkR/pmXR8
/EAZ1EZY4ypBpFPYlRftZ6KpCVp3ZudJRSa1d/C9UMWJRREdmnEO6EiY3U5/rJnA
/SQWqot2EXTLwdS/C9Dc3hhUQU5VfBsE9jpK3V5Cz7z8YovK2GA4Lusuogz5yQkU
hQg5sLIiPvOFQ2pI0JvAepzb9JvNLtUIfbmrfblb1wHvGPrXzLQG8UWh94Qr7HXm
pwKwWrDUP2Dlfgaq7CCqRej5d3KDzrLhTB6DkKtAjjhFPudl5VxhIFa2dqyd4Uzf
o38YnlM1UXH9yoUIPa7WG3wfNTo1mvo/uQdUfatRnl2BtG+11qQBM0orsTAs5XIG
H7QExHqKIuSSpENY6fXjjzjknsxK2xULcS8nPjYFsVR9y14drFsc6b4Ey872cZ66
v87H8REr6/zMqPde+yC7ZXaVXK0e/DrmEDKYRHC3yy19hBxyqlVpbR6H5Ex/FBNN
OfWTdPl/wA7lA0usJnMLHw7WsVYflydueN7/1yDam3ZV7qfRE3OmmIRxDGu3j227
kolyQGGBLrD1uqKWmeteCohzztk2XTZrhfdR4GvToc2jMYBLcCRT4tesPUOcHqmn
CqaLzZufINOjXRLFyHbQWNvg9iXoOvNO7chTFiEfiVk54B10VlekvsqaW+tnDdb5
oB6Dfu4zhuZJ+sQz1RyAuTPbtSMQQoeztPd/rPCiCv46ovh+lmqCPIIkHz54DR4q
ho/sO3tkyjCJrjMpE9zcvAMjpcFOd9Wofgm89jRt/WzlBYZoqvdW5sH2yL1wHL6w
jh4PrnbUBAQsWxq9PWNZmcFb3clJy2ecs53HQMrgN/NV0t4xsnMqad0+OqH9+cYq
CkTit30lPQm1/NCr8SONaNx8JE4KggyAmkkzOQz19f0V2CHo8/7zgVIWCs0Vx8Bz
9hc4a+J51vELPWy4i+jYmlEQVZS6Hbmd3ueg1SjjwJUpui4JDShXHz/y3/NwEhUf
aM/smf/Nn7yUFoWITMIEbgEYKub8NOnMcYEB+n5IFi4C86xS1j6iaMJipjHR15OL
kjhGFf1Y71yyzl8nMLhA+umQp7kv4KsSVjSuTK5WV1iShGJ/brDrpBgCMdW3pCh4
SoOiiXoX+GEAxFf421Id71TTjGwN2KXie8G/3SeDBYXCi/jB7ibgJ72qJd1HuQVh
zJw9+JgtKfGHiInJtk4/KthJ0cyNCKTNpsU8NqYFSI0PXKYUhLkwMm6hS6O5Fq7x
/2vD6cwI7k+7Kjn91dsEvdYkmlNt+evQB/3p9w8cbGJrbK0W98ap3duuk/m5j6nI
NqCzLmbYH71V0yTfpPgbx+RPXzlJsf6mc2yBB862t1/5Sk+2CAe4X4ppeg0fbWZh
Md7tv3+A3yyKPYbLLWZ4da9aH5aJjTZ4RElYHwr9uXeH4MeUy0ev/AioiVHwwawE
rm5jvrAgQN89x6wwojIi3cSGQ3B+l1uPGTNnFwW4XS0d1eCMh2RlMCd9gaYYtllp
aEpxb1GKI04ohnV/l8IQZW/Qmuc4LS1N6EqwDx5SmvEaHwZpioWE+ogQ6lHYloAK
vi5pKUPjD2vIF3BcQieQEVvzj4SLYlyDpUDu8WgzQr0xdYNGPH1JsJcA6LowzkJ7
Lkss7Wm8CXxCenSMMJvKu++vQslM5hi2FH3t2onRgFH8uQrSsK6F4MbyNvk/plUe
T6RYUZVyQNMcagt4lPKr39TdZ02MTdfIhQp6/KGxheusHv3j1uEiaeCQ/VD9lSlK
Rv0i0poeyQBBJpuQ3PwyyLLfA3HFyAEfA0QqBbme/S4VriXkczXC9tU7iV/mN4vz
hdgNb20MP5ux6wMvzWe4JbmdlhU3LcnAoOtod+73TbKE0OI7BgLj+Zskk/8KrPX2
4W8lxOsudfRgvEiJmqulV7nh5KTx4kO5RVzY5kZ2yTPSnHXquiaZCXb1Yx6sYBZg
QzG4/5Lx7yXJjPSl/X+7Dmk3MVoHWZxXmyX8/8FacV9I+uHXu8BX8uUnVX0bwSfE
I3pWUY1O/5RxGwykwhYbEb2JpNnz2iG/zWSIScS2f3+POeYS83Oy7aZc5tyWzHrU
fLkoJgCm3KStAfEal/Yi57bgx0Ueh2xT0GQMTsgb27pOw83JZTU6IqEVAHikDKMz
hwzuBpkDiEHKp/oWtCszrBmswIEVAKxUUsiiECuzmdjLvWHcBvmhGaZlgb1emUyM
yMUIPNWMab4euIfz9oAAvtrSWUaDlk9hQA2qJ8fCm0Apo1oAw/C9EylbDaTbkI98
iPHvWIYGY5Ii5ZUx0N/ejf3mP8ZTQ0j52qa9mVCtE1JKleG8u8Gkm3IojRGyFlCW
Zyr8ibfZ9U/D6OWOp0jnXxhyVRxi/t7qjm54VbgbW1ir/a5KphQXur1wfMoPOd+M
zUxicCqFzA0UGP3APQHmfkfNGm0/+E1+kGoXs5u7QI1twIdaRbqRoPx8MIzG4VvG
m78pUkFE9KjKn53H70KveET7s95yis7W65kC0sBJ9d3PSj7Lnd5ljlaWnMRMfdn1
RYTcZiBTF7zSHqOfC8q+aDJLO5byp3poVWchSjo8xKQDt8VHYSULhca1kbabPnmN
bhWRpa6cntvkHyL5XHfzBVIkZY+XJXcORBnqgsEXT2btJ1L8imCgl4WkS5aAuJIC
oFPJ7xJfOaXJ6NTo2bHwOzRaLvYL+P8DFWu1DburAFJlRjsotoQmxscL+8F3qpsL
weIq+CGFSyDQE+0LgOBzgFjd0RYuDyfCwVRc7XZ3B4KT7P1mUe8LBcEemIjPaXDC
ZECF5JC2Qo02ajqzZh6o0pxKUlWWmDbrsLxBLUYRME6fgI7x3sq38spKU8V7Bj3p
PgZkQdeNMQomJp7Pf62S3H2jpea3vcHwrpGi3ng1e9qIQKCoQS1IgWT8t06IvzkX
EtnVVHYgYkMz/tFPrfR6oZENLnya+pc3aDPEgEDDUhjxAlqdx2KMtLDWpC++HGsf
1Um9vGGru7cz6r/KRgTOGhFqXVbiFc3iYj0jbMegLYWc4NEP0sMAILzyr7nLu81R
9NFjDtsV0YOX1uQrq2MWMZXP7ekwfibksFwcrFOtNofp2c6WRke+vYI1xMG9Fws9
Zi7MMSm+OAWzvD8uaUhjgWlkwWuhI2ji0MkT0NUVichKH5E5vThbvBEKSHU4VVEu
9XbkuaRheavYO9oxqBG26c28hn/BtmeOrV2kYcKT6fkSeRLkx2mjfhbffKi6wzWZ
AmDLhk7D0gFaccWBlZSmWivPDu7oJdPrdLGHQjABejy1Vyd3pmAoLb1688RiP4JG
drsGAa5T/bnQIosAQPNzg4G6tDbxwk6+jtlRP0H/brcIoZINQ4qrfIj/3w+xtwo0
b9cvYS9CuX8NrDALTiA2uYY+5ZyY0SqQ55FL8kFrGijIyQKb4vutY9uIVxR76riU
dQ3DkuHwx10ZpZwA0vdQ1jJ/egaObpQoVLH6KNBLa0VQZ/4iS0i5b3ybuo8LjV1Y
Tx1QxH3D23JOLM3konE8F/EqmY6Wiy4PGXaYh/RnscgOyTJovptN+PIOzTZXe4CP
SGGUv2kLt6AuJgEHHd/rpLHSsXHBdQCl9L5uUQmOQ1+b1j54qB6aPq9qJN+lQir+
niJnivjQVS+jDbx89bjNusFy2lJDNl9OTXBznRKa2BUKv+Oq2Xya+ldc2RJm+585
ZoIBm9rIm/TRchIAF+KXD+wFMp7kGds8bQsPN1XR1djCXsn92Y+a4aAsRa2a/9DU
Gz5b47uoHTzKLDMmlk8cpOFuFW44l3RZAnP9M4wBdYu+7Ql1i5bO8MlCFDShQKLb
yrMDD8v7NsjUrCoAnGM7DHtt3sRQyWjT/VyIGezHemvOL6456gkMGUkkQ+tD78CH
KzpaVwc4jdhQv34NquftnNkMebYql0xWIXsAOuYqN2tYLrU9Oxt1aaPQvAFMcHXJ
c8+Pk1GHstV+e7XpTdv14Z+ETPwo1cM9szq/vU5ZNI+0a2tabxcCtKUHx3yzzYnv
YJhsw1PgEPcCW9G1b85PiNmo2cRgvL+ZsR+aBCj6N2tIogaL9YZfi2n821azysvF
EzbZrJP7DHkcdnHf+US1bUnRkgVu7LhTLv0vmpoJsDTLhRUrJ/iHUSxuYP6Y+fOM
u4LXXddnDiP+ICk2a2jNcGs7Qm8li9I4N0tn0z3ito5iKRlIHp5/oFUkH32OQ9Ol
b3Ql9Xd6qhU0vE6dKzZ7IC8cFy6NCHiLewRN2KVp2R/LxFYLvlHDwMhWMhmr4hPF
ullvxZZdsyKwAX7F3eCi0tKz3Tcj/iFwUojzAXsjsamCOA47jQEQcNOYfTzDtQMT
LtsMMPWDcwNDJZgD5BFl67UA2vpr2f8Wcdwm63cGacndKn+5mv0k4j9zODct8H99
4Km1USqM9nYPieS3aerwXtmn0FF/tREbcFqiKIvUDDCX14BwTaJgDRmxnIsEduUh
A8LSrzbRLcxRzZFq7gDlboCt8PXflpalukZM3Zdr4mlJ4e1Zer4JjPRJ6tos5Cr0
6+Dqc4Wr38kSQmV0MUuxn++TmXgASW0u/rXMVyzmV3rZCLj4lnr+vr/pPUzPV2lC
i7eBMbgSi9ffqLtmvFnXRXH4V+zEL5LN6f46SPsNp2QxJzaPIiUPQ/vtbvZA1ban
kWx9qBsvDsly+VxqDI74x7v/u3uWf3p8DLNVMCd6NcVZ43+SZIItgMZ/K0ZVuLbW
urp9rx1jG1PuLYoOOVY2Ozx+tHU9bQY8wIEnTmyoFZyqiH0TOftNmhw/k+zf0n5k
W/7DLyvlN/haXrNMryZjeEIBjrk6ZyzY/EFE/eEIL613Lh+Cb63OehMpvp1hcxR/
BzxmaS/K0/MZLJafIgunM9C9r/bWUe72b4RBltWF2jVeJ0l4Lf5F1L9vMW6g4IDY
cZHtia5pTFVggkAiprob0vjHx+uDoq0SWzEN3XkSitUVwARKR7pSk9bKJnubtCMc
sdriMPN0sDUFfW6Tkq3pfz/fXkEWxcrWiCZuOQd2YNfoiWRjVJNKi6FRVAWjEj4k
xvXiQ3DmxeDKbusAVeQJ665Xd37V0yCnG5aap7z/Z7UvS4GFTgJ9IitPLQ4FV/gM
RUC5raEGF89d5Y+AY7N+JoXdb/S0Wn4rSy7QrvDF0zICbe+6QrZrtMKTMfRl6YEg
+89aiQlPYm+TD4vw2ybbdQgmfsb5MAkxIcsey332SjtI5ReX3jI+FAY5KO48FFtU
ohMLbhI365mn/P29lJLhOAQkXlrEdCV0rbC1kn8DsODUARM7tXUkTfcx2grdD1P3
VB8S4+izQYskx6KGSfpRWF7jmfkhjJZJdeEvGfbcdAUyGcUwRdH6yf90BhERTSSz
evvf/6eYn0g9+kbeGig19WtRXmNfQrPFiAqoDAOqRL8aOKRU6E/hKuSQUdGU4G6o
tnYh08oo4Re/10f+UDJzK2STxKMihe3YZ/+baFFiDKGNE3cl7O8l69tOGjrSLAyl
xTwgU2V2+vUFcD6vYU7H5QQzqGZDLu060gnRVwrD3vZ9aowT+wviL2FxpFc5U4Pi
au0d9XDuSnitxgET83wLkpdJHN9SQBi54JJKTOvN83u+7z/0KwoixCDSRpR0PZC1
9uuLexuXM4K7UhuFG5CSETE8MUteFpEcZhkp3P9rpmxw7R4hPuuraJNP0+KNR18x
LmoQ697OVCF2nYChu1Jzm/p9u0ooH2qSgwpDkcRyZc28xSxWmIemaBxbWToPpuq+
lDKf55pHZgXeE7QIkdJnLbnPTsx4uY8Mr49XGsAcCEaJ5pJAzdJGymo7gBw1pIFh
614KPwDIObwF4QYMvf5eZuiRftjAKc5z467k3MKyHP5DoyVWC6tnyMg9NcLgOmb5
o5GAqPCKhYP4/m7nzWeBJZhHcbqFdy/yLCUdY9QlAEAD/C2T3ZwyvA7qeGRcv8+J
ZL78BO6NbgSK/ecZcChkEOVpC+MwwzYTE7pNDqQTyGLSTLr4qF8bmuI7JgX7q7aY
l+0eSkFW4axzXcNkksVJkJ9XfiYwoVzFZInbKQwoA27ZHNxklEICRNLr8RCwafQ2
OB8U0yRWT8Uaj0Iw444NHz2vDFUoDlNxhYNfZwqaCAI6kYrftiaEG7iPp3dJou2E
VVm2RrtBylM0wMerKRmvkNREmSwlB1cZjdWafc8z/053eFlRJTiOZYECyOQd5h25
9dbRFKz0QCDi3r9fWTN4cykfjFl1IPUJRQuGa5v2C5iskGxBFM1lUMVtos8U8JjY
x9hoygVQA5UrYSQk9HktgpjRXS0/lJQXH1QjbhdjDlfeXNpU/PzdqNfl4e30b/7Q
fM+fAu9o5E4AbVVxXVL1263fzigRbXfD7bHNY0eVBqjr5AExgQhT+InND4GUVrwZ
Zql/tw2/b1OQnziiEb6bl8beeQMqL/I6E+7OmJipqvuf0E8NSNjCFJ3ahDiglFbB
kmkNNrM1NoULsXzleuVGm8EFSdajgSvNCvVyfw8qhOdQTZZ1B6jXFYQ+DGjXniwV
NzlY+n1gM9NdLGV16ZjUpZIRYOxznd2RBJjj287hsw6OOUu2Um05Ahh1B2n2yWil
xyQApgxYunIp5q10N+6JcRPx9DDmEfC3dmn8vCJwRQBviFehdlhZetDb6pcuYLxN
sNVrN1mcjp69Ax4N2aoRm7hPQRqMI+sbGdKowhd2rn2i7QfY2KpuyRRXG1U01aAO
wbbZDDos4IlZ8QWqwfBoJyIyprxde3BIwmNZT495bI62epL/DNN6lseXgaHUHZQb
uT5Qizjk1fxvxPuR4zs5HQwZKSJC3lW5JhODY0eD6ltoIgv+TilGU2HyS+/wOLkn
f8fkrodFX26MC4K+JiwUq9lYGtonYIshe3RnzR8HYRCqQqrVomSgXIY1arc4n6Jb
WcllHeScsTyPybzeDgDasZMganjlkO4WJbRVPBa+IFhldITP05jil0nNqme/J08D
V6uF5r2LsZcT2SvW6RMbu25/WCualJhjaLgE3a7XNdxWEdTAyOr2O7fSVrC2NXww
DWixxUiEUk4z/mCsekQJZU7QGdhkBXvU6hoDCESOdGBoRlvSVvueikUpKtWF2y5L
/NiP9DBO1qkp2otyWbfWYG1bUzl6f99vPjrcKmRJ35lZ4Cdghe2E+4xcb+3h6wkM
McPXBuNxJihF1GMjI+dFlVDfjnzrSe6Ktib0QjTfJ7xqSAAtqI9HE7kWKvooiA74
Cc0QvPubAF9rz3v5INwwIkvaKCFz0n51gptwPEB0a0NBSXHZ0z5pyfPrPoGBq0Sw
7ZuwXp4+daqA53XnZRbQMKBao/4C1u7L9rIzPxu1DBXGGP2yg52//x2ARs8Vjpge
z02aL8eWUQ7v3v3wKwjrvgHG+P7aHwx21V3lonWC46G50Dd1BYjOSvKJX81qoXI3
wBr0uj2pT7rXIFpxCVME7iGCeXM/jiWygJHxIDddtqcxc/MU/Rfyif0+liojHnwy
quypWxdhQIjI54pSyg8Gycc7z7V6C4kH3dHYaAkopj5viIiE3htVpYEo2qZlxTgw
4Jbb1gCRYm82zCMYJF6/O9OQJSjg3OMwNysIfl15F9r5zaeV0cLlFhNFK/4d8rXw
ecdSGqKUxypqH0bm5RQu5OWoqtF39ezErSeO+BnfSWbEDDIwt01bETbRavLo1kJZ
Lg0Fue8k6tVllLbEemI8DnhNswi8U7ojelygLs3W1KOwKe0SjWAM8mARGQsbP2Nm
8uT1ZX85EnzNGGe8L/SDHk63NTNO2mxiKwBEJY8lmxKGLq/jAJlbYISsRg7ALP4V
c+Zpw7JNWTHVze+U8Q7Ilaw4PyVUb5zk5m3HhkV8DWTf3iPCOTFuZ8a8o+1PsGx9
rnXXqfvqF4fteWxkCeCIoJFFXzHt5f8zbkG4E+2honzxAkqKLg7mzV+jTW1a+Blo
AUcQ84iE0WG/lSFk+uff2LclInUh3gHMorRSpyd4ZbhQW/l6hua3Vc7NSEQoyQDQ
PBgd8TFSOkkyDhhgxgKqDwYom9CVhij2id/3Af9ku0eEL//e+k/aLmmzLvqdwjso
goT2xiVQH7a2ob4jLG3ar+TnoB07fBDwXNgULuv4D3f8uvjzgicxzjb82eSb7VP0
REiIoln7Ucd5cUTflHczi83SMGgzGIq26OinV5MLCIubs6RqK4pm5yPkhGoZoiSY
Dwvi+GBpwmniI+GGBn4fuuxD/e7xjsW0IW4vmPIy11Q1i+aUAieyM6tC5APrQsRT
tvNPwZOjrDNnZKBkHCaBZ0jx9o7LcCcMa5owHE8DDWqSuqj3aJcBQ2o+imuoQgdG
u9Vwgvsemv6zHwELeRCBWTLCeeI7E64Do4jS6mr5sbAfLNCe4xD63ntf8c21vqNL
9q/OPoruIxyG8qpv3pvHFEp2IS98Prq8qG/Z2K611juw6S75iAODvR9kFYcQdHWa
Zk2bh+BUB5kjoxDsFLpjh0iNJ1x6YAM2xqqLmljqp2k7TCHdH3jEMG3szvZ+l5zl
4R40n0+SlzBALYgBlKXL6Jaht9f0kzHLJGEm04nY0lpBTlpCt1jsZj+qCglz5kEG
ewo3obGiSGI0lkRBiDYfFdCRdXBxQgLJPbARez7PaiwwMQ0qtvwXV5S8KN9bwanO
PTpHV7i49LMZa9a+eeadKaWCve9EY7Pyx2LKBfoRm6USXj7UQ4B6zmr2Gen+VRu5
gPnl87Foj0Y6az2OrKWG5r4i9NB9+u2htR108ceiI8hlSUGTFihoS1rClLPqzr4d
5u3tpa/BPDvIhMGGqVUCiP7asHa/pTGWA6N705nMDT7R9vN6gXYVXB9c/Ti5GPnW
0HnfIoqXscJDltj+8nNEF3MwwqyW2RpF5aw/XKPD7+mvantpvSl31nmX6Y3RGAKL
dYTSX9FOt/kMnpdOzB3LKta7fgkvCRwHtmd/I7M8BYq7gaCyBWtHH69CMOm7oJkQ
z/8EFG2CSPclWTvi8hzzDmpe7Z12+/isjAa9lzJ40kSMbutk5g3HzIezZn4Pgwh7
ea3uG6vFQp+RsMq/iM+U3kHWlEGBya7Q+CDfro/F02cVcB3+bZ1m3KXAQNR+C+eW
RIfb2P8SQWdEOS8bQXNHKF/9gM7zuX0Rel6R3JiJ52WHEnZcg2/MrXzHqc470cNd
YGBZKWnz23iNYHe9mr0G6+XcIX5tAO6cvAqoullhEv4IMtSMrTYKhXIfEzWrfJOy
8YCPMWYM98tLqL4S8UqSSxI8KIRk1ond36HRJdAipvfrjkPhFFh9YFspd1tOWQAG
wXpQyjeVUTqKGcyKSIO9Qi8J0AmdW5rG02pazS0ttuwFHj2bOThAooys2vcJbnUA
qGFL0OKdn4ZGb7ul8+BkoySirmu3l35EZR6N2LuTsE2Op5++UvvxdUv0W3Mis6gj
ZW0I5dKQhwcchR3AeUkwmKM8iGMM/zoKNuA4Q9nNjA1ic1CQIy+jK/nj86J97s7J
jbedAVa4FGYu/A+zkjx7SH1Gfk+b56npKHpU6/e0y2VHOS+w4vBqDQLKRwRnilh1
yGD8fD8WM2u750Tcr9A4O3kiNT4tikn5qkGb1w0IP3pp66ODkWQRtDnRqOVlKkqE
GhtZ3e6Su7lTg7xkKr+fNgQ2PCsoW9DgUHCxWluV8FZma+tCGIcGhsw0fU0QcPZs
xWXt70uCVGe580B+RfMfyRQ+t+fWEcF5ZdSvg9sryuwGLXmaK8gYgbt9dTF/ahIi
3y8b3KCWZG6G8ObZ4AKDxP3jd4xdiyPv2sii86dHHtMLMIe/rfAwxvn9zI/1c6+n
J9jscFa3/V8pzbUoBEaMMNrlmtTSf3ayoKj90qJjcgQCx+/22htftePUp5FProxI
jAqlflUBf6roHE+uc8HwJucwoEBZUeMS/a2gtrmygV3p9bxSru5AsL8QeqhT/4AW
cd+qTzX58d0Xtdmy+fXPHL/lpB0Fk9MpWucTt7/Iu2uzoBABHOmAXgxU9Ov1tWGs
Jx3GiZcjK2d7pOrph7OKmCp1+Dt8+JkiTIUPnAf8ci2b0qWUMD3PmG+Md9fc7WuB
TbZnPor+Z+jLEDL4ANT3RsgZC749Jm73YWfQ3faVUjEmsJh4bfmAVZ0AYA8szL9s
UwV/4salgILSVTpxBYGMAfFgaAI02AEXiGB8K2wG+do4DhBFaSkWUhp1sbUcD16Y
+5ZNpjNUUqk6X0OqVEJesLXR9ZDkD1Q0ew0V+BJaMq+kDa8XGvLEkUFXsXwfWKug
C+J0F8LSQafzJGvY7Xzsg3Uf51bM758quVM1T/ox0/ix9vjB1+v+ICk7fwXTcmoA
rlsgTBy4E5I+RRlKJrZ/oiEnzkP0V7NKUYFlIEuZyDDIdQY5EC+afIKnTewQyn2A
sql8OkU3PRXXS1oj+wXvAkGVbKus9c+gtPQrlPpjKANCVvyNQiYzTqiBUj/YSRxl
LoPXXJ7tHQWrP5HE1Lvd0uK6R1IGRn4oiw3e60keajXJwicmVkjoyT2uMWK3vlEl
g9EghfYXB+eWEjxU6U5QMehHMGKWeH1TtBtMZvvx/9v1i5OL9bDYxiKL5c4T2nKX
nQBGnHJLmstmyf5crRaecOYIm9aIFJ1DrB3sQ+cUyQRNxSf2pCnYIFcSf//p8IBR
OTpU+LjJPem0Lv1ac0I1aMXHT7kgFVp4LVQM6Gq7CYMXI7T8s3myEOIlXcpwOHDe
je8y9XiGDWAAw36bTtU2mpDxOX5/3uD+37q60j1hfA6lDKEKqUe9/HUJBQ+BuIRC
16P7234y+M2xh3lVu8G+VdmjFN4zihxuvF74reh93KDP5VrEnH5wjVlg2Mg19Sss
x6lt11eikJR+IKjiBEAchwop8PoDKFWDalE9uB5en7jR1grrIFfrzVMavDXniHnS
Kcs3xnglO16agK2Se3Van4ORw3x1J8alwmm9D0iPxGpmc/f1m8NdxB/sFrsO9mKK
H/7foPUHQYBTRKI8umlxBtfg2lC4DAhDdJ/j4qwT/hn5tq/ONRfUJU7w7sSJZKPf
dsp7YBv5CRtY0PSo4unL7SD6/HqC3j7IPg8KN6Ngxd7K78Yl2u4KoExTMCKlX/V0
70TylBruVoo+vf8zAjF6EyNGSvahm48/Uh1U0tyAPvWoi5IJKrD9EssSV61PjEUm
zqOQ9F5KENQCZ9t8nktIjpCy/MkJn1/A/TQbcg1A/fIIaNOvHZYg7vZ6cof957Nc
2i1lM4zdMic7pNXPdPV6ZpQXseI6cHY82WjLNK10ph8tbMlKmvVcS+pFvvJ66MJA
OH9DmZOJ15kNZULvQGHH6TrvzZnSjNNrj7hl9W184y6Q2E3fl+8wJcL6B2+zdGVw
VqARZip0o9krLfOZdodd9p9zvAeLA+Bj0d5kSXtGqxmMCJ1khMY9eBmdbeuO5TV5
+4OB1JGtegbuyGG8DIDKc/cVuSTwpz4SrS10U87bNxkaAB4J98BJBxNWwO17z43/
GY8N3nrxDjcmQKTs2wP49lKVr8aHUvjzfDYE0aWSAjZmEin20h23lAnQtjdZfT4c
03U/jo0syty+A5U+mlbflCCFGdW+nzfxQJbfDyAarEKdI0hSVivNpaCPOADBnLVE
s6XgcLQFrSrhYCAYz/4n2KZdMBX36yOmOyuvferxkFfup0BGIA/Zqd6XRtTrsPms
MoXpLs1aLgFNY48dAraEyRIihyx6X219ylobgQjGTx2unHfou231y3o9Gqoazvkf
Ozl3X+rYmJi26un2c4aqlRp9tCwGdM/2h4Q39I9S1aW2dVwkfhZ6AuYlvWUNbB3B
0flIOKDRhrORWS1QP2TNHhsLap8F/hUbhfAEEpeOPEZuUT9wmuzAX0nNx42tdpvV
wgOIUvENBczmYTDSTNhq6SHqUkHNLVvfDQUkurILojx1TCdygd2GdAmErPiGmB38
KQvpwDVpDRQJB58u5CTX/X+LMwhkTAqIdhB6VFdGiI4cnsreXPcmp99T+QRG0Y4b
cQlDCsg2i5/OULar7DMsVC8hCzkul2Ym2L0SPV3WElilcgX+t8QRoA60wJCrdQBu
3hDhEuZM3u9Tx/14uxCf2CUr7T1xJfHRASco2mlMZnR5Xwl/hCtbSM1ACMrqANEU
odQJXf2C4rio6Col9r/rrQ4eP8aRMDu0YJzxW+6CvntpWynM2kDcWnHcc9Oi6tEY
b9Kyf8igSPZ0K34ZcB2HY+cn06OPwl1d6+kgt1PDnmSfsrhRY/eEP84aFP7ttAUu
QMXGvq8DYJYWJCycyjwMBa4LH1MhF6KtS2uUVpbtoFEUs2iDAT1qCHE8czpMENlS
/TEBQc97Z2grjkG1jOONhYPyo6u/rA5sURNCOUqW2qGLlKag94PMT8E1l2H1rZ5A
WmkcnEbrhEX8ZmPC639Px8TiBzQXf+v4G2MRPJ/m5NSAIC5FAFFmyUAbKgSnmEIh
jWlw3lk3ucd0DPpJX8AnlBKQL1a0bsPadYmd3/O2/80r0gLqRWSRqlOjDSxM/0xu
mXR/VcCBxIHXIiq8tkBFXZDiVwQ39Hkw6Je7xsVGMAaP0gi1euZek6LzxS3+amVE
uAUVbj5V47P36pptaz/l+/l0Hpc4q78ruiMGgPpsdmoZczX/fjnterTkP09aDwog
3s4jHUo7G9cYcTFCGjROPHrsvDZfO8U5GdLpUgHtOf/coMjdiOGyOQb/KznNJfXp
ILfYOwUqPvkPARdWKIp9SemCiUjPq3nDfECcbKK0J8n5XueA382nnJTCgOKwlx7u
mJ597qIpUgipeaboeIANtWbDeVFmynvOlRxY4VDZrXfB5/4FN1mSA9LTtsmyFN7k
5MkPlL75SWdZ1Ps7d5KWfcQ2BW3Sf68LuIz7X0b9D5EoLAF7hnBCsMOrX6bd8Rjl
CqjvWKJy1v59+DzGaAognwOmRPA/IgE4naCo4pi1+ObIQrdu3VQS/ZsXySZYJPiQ
yWD7qTiLH3qBTcRXQA2HMgePJQbWaL4VexrDMEZHkJ3jqub27lYWHztgzKsVmlSo
3ppd4zKTxmVkBlNK0HaL9kEJ1suMnVJTKBMxa8INmmPal5S8/+aQv5D4Pec5UK/v
ZuKNXrn6mdqVwrb0vRS7R7ptWbz3zp7rn9QePSkU8FypOmgTOpwQyWqil1N1Zof+
GMhJXRbfDhD7n4HM5KyPe1KHiDUs0l3VKyuALqK2nQrzCs9YlRnxwdwXKqMIYjcB
ygp4y1SMmHFUspnzHyHJCfvKWn06zqO8bVtr2PeTiJiF/ruqTSHlqVNcDAsc95Dp
VDMVmYmeOL0wUy+EoMNSNwtgmqOLm39p+vjtuu5VjC6mtFOBNbS53OJzleSAD6vO
NoyC+cIsBhYWLduyqng4ERJxN4tjCHB1eJ02/zaHy5BiTnV/+U2SlEA6OjRK/Y7V
/NKWGgYTJX/j3yVms82RyajFt2a2ISfssvVuetUIbR9pIsc20eQ1yQ9yWY6vDbr4
bG+U/gVwE8Sb1IExfSBHkIMAtIYGZSK0qo4aDTO3q7N3GRkr2/SL/u0fMwY/cm7S
tczDGzjtWdq+o9UTGOSqzXutcYcLA8Y8tuP/CmH/Erqe05dQpddfdmtU3PSOBvvH
nddhWiK/Puu2lOqd4oU9OoYBE9zIvzFT3v27GBJQmaSTgno+I63NMtDnXTfkEBFa
n1LTbcHFeuVHmD1HbEjy4HUFOGVCfhlld7L41uL3Frm8XJH6Q2gknIrmXzpQF1/W
Uj9CsX0hO0Md2msMTYO22wprgAI8YUaYeQ5wUyHkDf6sOMYYOJDrwY8Jhe0rNbJz
Ma39WyQqxi9Nr0N2N0+c9Hv4ZVlomdrvQKrYFe+mukkItuwwH0lmemSBGF+uXfLo
mnJLLsqf2uKSjaiKMbfHZLCFsb/BRqD0OjYGORmxu+pZZ2Fp+HXjkovjzsSSd/vM
BURtZda0Un3F+6YZrvRfLTfUM55egPBDAF7y8sCs2Gc0OvIF4movTvbrjFmzQNTG
nE7VUzE103mhdIsttnT8PB2vDZ9quwzFWyYOZFbk4vsvxau8XYqU8gXYoWli2hck
D114qlfdc51nv6Sr8+o6CUAICcbw2yfysS1joXsjt5Ot1rSvFLiRMJuQukvm/ZEu
MNX3DtfPMqe1XrEiamkvBV0MrjEYRyfmYIdj7JuxS0jBVHTb0uOdYsDbG9K6jE1P
e9KR0+eZmYniYzNRbCrM0LwY9wy6Cr488u4MpaXdQK14tu5BJmwHuIdsBfbd+xoK
mgN45qwCVB49L09JSSAMfSzDEpQQDsSjywdtpwPD5bxT4RKVt4FFsX9TJblkGpPu
NhkI10xD+TukfCaRfv6DfwrrXLDXKMA/8kxhLyMInSMcJWee9LXC+BCpJ4Xpk1+V
zHsQf+bMoztpTa/csRk1mNvPXc6cqQEt3NiT1wFudJUc3A7E92AiFMB2+OP3fBap
/p3d3FzJpFlOymfOcsDatwlLrQhWdHrXVcxGfovvl9LJ7Re5+gzNx/UjaK9HQSA+
SBb4PVScbXKAoyEJh+72rfZVCTTIecxNdtC1I1ucWECCBG2bLsi+oZoYWzImt0rC
JDP4loyp3NMvAP7bW7PojHnl6mZmUqTHoSSPGeXYo72dfZzXKRBx09BrMC6xwkIS
LzFaQ/8LW1QA9S/jyQYE6tAonJ9G/j56iEZCAWxqpzHmNUBPa4o6I7lXF74v5JED
Atu7GA3wpbDycioi2pYjzyV9cb+8p8e5KYOnR0R4zDla2lpSpihQAar4bcfGuYs/
6gjsfxLfg+jcghYujh6++YIFvMrc1OL85rzMZ/bgD9r653dmtx+ol5se3sh//P+R
r49PDHhDPnA7pbMT7GaZvNCBnRjtp2yVGRzwE11A3Tfq8UV4lRxgC8hh13oIoKDT
GKropbOEBQnrqOHYkNn52BFTflIgk873fy4WCdrH3OIluEghsoX6DPs0MpsLQbBT
Fc3FUlq4fnivuvrDHKyYeZcRFVwSTtzq8IGJUfWZaXgEXpPsiZt0pmo62Y9t+d5+
JD22/cwp6kZgjgiwaDuVah6SL/V38Ho7Qqo9tf5shcqfzRNJUb0KkVtjH8HeBxGQ
sCeBYGheLOx1OMCogtdVSiI8/TeP8JdNsDXPKalqSrzQBVROdLXXw270Nr8pTyfk
NeWWTB4BCoPovWTPAMpY2sR8UCclXhfNalY465WzQ1QN5KtItztNuaUQpR426jX5
28HwwmlYz6ijLJ097FozRiy9orpqditAHtNICtILL6Ar+L57nXBheneFrvhc0gyS
xcBxW9vgXji13ge7cKA5YOYtE1npTD4OdoZm8tVsK8H4cPmsRz1noFDx1ZIwaOPK
pYhHH6ONwDeYJbjSd7OUpcJhV/fWngI0ztlf2ArDOFX4PCJ22vs5nYE751w/Ecpl
/I9y/zsSNBRtRtWPV/RpcqkxNfFL40yvmT+kkc9MrOxCT1YboWeqbRtzJjDWPrSi
ZzToSKEAcyKJuR2VNxZtu3GD/NUwyuOofKXn7Vty/MhcKQqAJ9aJ+6OPpU555eyf
S9akymsHoMJ1sxmOQTuIDycOoSVkYDoFBZnMDItPRymgs4YHzJDdHqF5C7M1hx39
E4D21l4tyHx6JhvGxl14q7ihUY69feAi7xffZAfdEcI0cyY8+ugHdexRuC4r5oz2
wHdpiTx6b3mpAWfWx0rq9UZfVGcJxaozhf9cbD2hMuUn1GOi446NWYu7ZHs8aBJ0
zl+lQhHfsyZb9+zyEwTT2/TZ6uEd2IRSuTxyv+F99KXcFU0h7Ju0SfAjNj0c29pZ
ELBRO+c4hNznv0u1q0q8Aop8obElByq391lbhV9zlbu86+CMmpkt51cb6xorAjck
FjYFwxydwTgVW5H29E12MkWm1N4xv5RulmCGPWeUuig/SqhSBwnkIerJ2mgP3/HH
yWm8u25yv1v3GKqb7vx0X+wcLeynJ60erlIrq/yx+RYMQ8/byw4uTsEDaOyXxACP
gT1w7gIwb+EHeYyS2gI+G8AxU84CImCSVHOe+H+3gsDhQ8YU9vQVdabCeHors9Q/
H0SwIWa9hwc5L4OPDcC8wAKkd0tAOeIbB3XlDyleKCHPqjPD1WOtBPGJ8TdZQGXx
h04Oa5DazBHXtLnWLnKrxhzLGur7rd85md4kplEY23MgYg4KjHSqebfewkCcWDPN
U9LKicanPS6cqBZQJ26IwOgMRh35Kwv+zeEfndvIFwLz6Lp7ZJmR9GQupEC7fvJs
sKzy/t3Dmpmmqkb7Prs9Wp6FFTGnRWzvI9RzwUQ3POkWICUcUj5sJX70YQkFf52b
5SSKd1www26zVHYtlKB3qHAlUxi4DY1gYs3USuGHYSgwamPGBBurV9drmo2SxyTp
tdTJJNUXkNPOgqqS6YhDaHOOOMy10yctnGJMcwM81pjOsK3/6Kjpba7S+eRLnvUn
LSgBKu0i1NilkYBS0ht0P2B9P35TfBNWYIXqqlwdCU+UdDCNzNXwz0B0qQ0KD9VB
fn+tHDLEEkrmSiaF27RKEkZkbWRfm9ys4AGFOf8E9CMgR8wpqquEIV3XDLQUkY8V
vJA5wDfLemvJa9tNZcnPtaOFyzzpeeM4VqqsQUMLlrJPdLgU8bxDQ0EwTg1Fbmbn
Q4KoToGC0oZ13lyS540V1Bpa63fz/j5VgbzMe5cTU++DLaIh/8Mgz/gdEq0suMYQ
nAbZ5I/UM/93OC+cKD85KwrNYvJovePprvQIkakuwUFhw5kgMURwGefzB5Ij5XE7
bTXj1GZZD/3tImXm//PtDvMTwNSYe906HmdHU4gnx3ezJSZKU2I2FA5edMFGNlT/
0N9Cpt4kSI3jIHyb93GeywewZdaDmuUQtn2kbPlDJ+hVFW/vGeTkhqibZPDxIL37
yTlB1lJtrZpOIgK5/KQnYisii4knsYsRayfuuFibnRc8K2HZUclj7QAQJSGnvpSU
QDKyco5WHSPjVa3aqfnxnCYqAtWKH7K29ju8fxWL6DgUrQi52v5AZ9a9j/o3yHCg
d3rQFwkvUfvsL++igPhYGBxjCY64r2lF6ZatnYAzelXKSjI9SdnnLB7wVZXPB5gJ
38ng4EjiAtJp8pAef0Qksx5bFKYD6XmEgiEjI2Rxfsu0MwtKPZ5eYzWnMl0tyhS6
UShIEtnGa8b81u46K/tpB5Bnd2QzM5NvJl9reQAZR6Kyk2cBEWrawjEfe9kduyQO
3thAGlzXoV/O1nnOUd5ZeTvCB8PjvyOlgDXLW0ukmZaD8UD5wCLVHpxlxZUHC9D3
M3c1MU5zg3FIbjmRgdc6ESOgOW3DFgDylKYUKqGzSIRfwu9orW9XJWZwJysnlMEV
7T1XIs8BIpjTjkcto1pBWBjp0t8SRwhKPw0mOzJWAq+Bz0DNxjAIdvN2WOFspftM
AZnJLUmfa1aUvmIM2yzLDm5XiqeistUr1kfYPcXCx0bC1KB2zAp+PBmh6HsZg+GX
OnSKN8Z0h59lReeOIcsjdBb6e+jQnaAywKS+1YMxcQDeHZeqlvk5zRgQURveDGUT
dUq4L/28nFHQ0+mwQDgVKyy4PmGuGFrJusaMiidyo3M/OOidvlTxGLerS97h7quZ
ZT5iw8tzidHNvGGKnxXXgxBrOOx7D9oHbOYdkDU+t1rdMO6iv5uqgN0n5HMLOL04
x0JYz4jXAZVxZaaQE6Z2xAboCnx2HyvXvmTNDVVQt+Xgwq7zZdo0S+7zGn9R5SN7
+ZRKQCnvFp7k8TimG8sPiCA6uHOFZRukpVN6WnKyCGs8+vrcnJHGl6mPpvWW0bXC
5NnRBUMliROxP9VfupCg1mqMXDKIHkwb4IGdOfZD3Y9NGKd15+gpKZDJ4elTZ5V5
e9mEmJAbV1+AEBYYN4600Pe6xWfLL97QURWOCGFXmj/ZBM9QPeAHlzrAajQKC5Qg
bP88xg13ssTGVqEHd9uwnSkOoJKUQ23PWBU082tdvHuIMHsxK7/ZXiRu+CR/RGYH
H4usRC88sBQxmbkrWZbCSxXFfZ/P58tzhWStYAPTely4c4nGU/N8MxRhxbvviECN
Dp2P2N6xLwiLdm5L8qNZd8xR6aEkivQV2vybsotqrhPfemGs/IZqaA3xsPTz3Ug8
wVLjhOUH9oK4HstckGsIRsTxWp4kHrsNnf/f78mS83+OIgWuZ4L3f1rUgO5IwCq9
H70cxj0xrXFoPR0y5IQUTuEsnJrRSLJVmDo4dRjSL/70oDj35U26nc2oRXVzH7e4
Z+r0AV0zAOKQ/pY57Fcz7zBVAXlFsZARLV4+AGQjNvHWmDiMov/9Dvm6O0mA+7eG
Ie1K0Ml1wa9bAos/HTXxf3QcRGqt7axw+I14kWFW4kn2eeWcSV/MELPYdnvM/ej2
YLfw3cuCI4i3HK2CONX3dJ4Q4KfGVW4oJdRJDo5clUM9WR0qe1SjWElkBiERDB6Y
oJLmEPrml1KRvXsQ0fbXSJlIrtf9K/10MGTN7O/UukpAXRletIs6rhnXYRHG/tSs
KQ3kScZhcvT5VgU/Tbqc+oSzpFiHNFWNHu7gUDYkaGs4+0Ok7MzssCIO2nw+xdgt
+slHbNNc7yTeEwS7s1MFslfI/K6+zLIRtV4vHt2H8r7Grdu7ezr8POue7qIjljsR
sI9ykRt+9RbBqrh4eyHE4BV4JGKNubKL6JyXGnSnrBtJIQph7H7RtYPx1Y1xHvKX
x+Q4G3oEEFPPAlzyl51xgmvEJLrh/CRoveqsjN2v+UlrmEdoVWHGt/hoT46XTasJ
63CBETqyHDrzb+SokMToEeql1tDTOQERNOhH7mQ/ZIDW/USX1Dxdzo6Lpdaf2r3i
mxl+Le2gr6I8HLN+Tzj4gJgYHb4D65KNsZYQEzLihmL0PGvB6FxUbNFlMbk9Swgz
HSEPtsNvsEvl26A98Qbh6Y9mOkDa7/X+yLeYvkB+O17ajHK4fVfPd0i2xb7UowAl
GP5TW1fBEGL5Dr007hsmRhxg36RVwWrJXqr2WHaXgAg9mTn1artgknLxgvXHrFbh
bfoe9BGcS0kX3boXy8gVkXNwh8j0OdlXmUTVVEVtblxBVvNrTc3aL2LM1N62QO9Y
bmRSJDSV1jOkWjvP6OOmMYz5IGnogMboGq1vafJMavUbg+D9uILOvk9Yh3vl7q+k
S+MgGKPU5lXELBGgJYT+vnr1I4RZrF9rqw27NdE7Vvr5nxlAbFqJz2oh3cqQvF1j
C2Z5F2/DGfsd5D9hhnHtWNtlEXeGY5j3O1Fxf+t1qKkW7y4l1J9HyIArLoEcrPJt
Go9uWfccbMTew2Cf85Mc6aZi18UQ0bFB20KFk8T3vbjhUoEADB8LKvuUGxM7eUhC
vJnUqx4GqbJRejscBd2R+0El8igRfVdrMllV2oMKm2g5Tg/Ecmur4Jmt7NWNKOsJ
1CHl+WzAFfHP7iTc3F6zFDXFI1Zg/ChEIAR56eVSe3xZ1ydlCz9bPr4dzmWiWiQN
lNZyW8RutxNVTnPaCX1TrVlM73JmXF49LZKujlpFAX77aH+/sgBnNS65mJzoBMsb
U3AloR9mviqBLJ6xWJ1qZIVSyIM01PLKk7LhXPRqBdpGzY0O24l2aRuCBSIVAZF9
j7PtKjt33tTqO5+49KGcBRDCN467z/bo8JMNWWvoQ1krmMpcQYELqXn6OxSrX3I8
cL4DysuoGDbshKJeRz3rxA2zcaPtjjUD+b+G5PHkWvTN0rVHPP6T+0T0wOi75ef/
BvjwYBuLYhB1tsL4/JFdjgHEi+lPUpdSMSji4s6M0IQlc5SapHklQ0YB3XeiMQ3Z
AWhH6ZUM8mGpfyOtUcxDHQLnYsgtZ/3qYOfxHU7VqM2NTvIWU6TvUZeX7MxI7PVu
RByMyNc2boUzrq7EYLsrLN2Cr7tNckQad2pyATF5dnd4yz7Njfd24FVOHXm0Gcgx
eyjDoXoGxHhUhQfKsgqDCfxd8psOdt7H6dL42OhqP69U4WF7a23XaPOacyHgBPLT
NOyuaWNUd0ZHqbuYsdzDUZEpB6Jr/QFmboWEpDVaRojacVjlOfhJNAHTRSQr/iWL
DrtG2+zCUfSPInUP6z98+XMltUUo7ZMlNVfVFuPwOa2siuZRa6f8ctoJiQl6SbPr
KdkH1CG2VEJWCkxkeMv0QBdsYnLRlEylMcLMCs5G+jQmehycxzpYP2PZq4XXuSYN
6dcw8mK/cuYFDZy1Wvl+W9DT1QxvG5PB1MVpyQfHIDkecE9tKlSmj+AW1mw3e4TG
CjBKjSVQsuJCKwX/Pj00qLCkhCsyYxbrvl4tPn0V0yph9bVC8eA1dMXbNdBIB4R/
O9EfJITi7+uVaJsoN01JZ0lo5mdnhTq+LyUa7NLGBP3ZWJpBNRBTE6m0LkZ1RZFk
DWF4rX2SK02sZjqgNPTDMIkmVP60vhZbBRmRtgpRi+myLu+YncNrcjolXQiy5Uy1
7wzHQcqRW0fFDBYCgh+9ByABNAgZ1as0OdfUIA/WDz+mEDrT2etB73+F0X/26k6d
zMx2K5bJ6xn2f6MOhp74A0BmweO3jt4pt2rRSKb/OUSKWLOGAJ1TKDFBGJJcE11q
Y8lDf4D+xzEnMEc8MiBEDwT9yezYsT4NkbFyO5wyylznz+YJSZkcZ9vIKG7zXshp
EYW4/Bm//oj8bOpCkumsVo/FIGATuavf0d2TtxmdKEwZsqI6Zfnr3yDryRqUtbE6
QSpTJHbcgxb1N20vRntLXqDvRCkcz40g8++fDnjsUSwfWR73ti50iC/q64tTdR7O
5kheYE3iPffF1TkOQb1TGVv4E1EaCmqLc7IP+rwCksVIcfozZz7nX6Zw/YbHAqPk
6Jupg7orqh2oziw4XB3s5sAQXqArkFWtMtUHzstOofPpSb04r8vd9bTXrFRJowDt
DYAmZLIiWyHg+c9AvPv19a+Rymc5gggxyY0ODBV77tx+I8gZ7q6sSWaHfyi/+oQo
AZGs+63AbeKQNxhDqjDwhJJNQMEUWwTtTNHdez3bNAoK5l4YG+c8ePyVDE6Q6lvo
b5nPezHmEb0aMXlWR39Yw5hZjsd+7JOd9HoTbr/CJ7msoBX/bYV6Ys3Eu/EWmTwQ
mk44/XuQTraBJVx63x81K81a6Jwaiy7LOmLDIm6VNuesvdhUmo4OAKGL7E9f/T2+
IuzihOtOWhnrpKebtRXV9pwiiYD1U07pQVkBzTUiwcYDsTP73GONeKO7LAZO3YCR
OJ4eld8X68caCmaU3xi+ar5TFGbOUo7Mwtvdi36JQI3knX1rWqxTyozi+by4Qsmz
vfo7g5AVcuNaxAIL2VCdaij7uB0Pmejgw76j8pYXFxcZ0EXl9aGCzig1VV1UCaiD
z3UunX6xufwcBx6OyAplu/peLHMvaMNw3Wm63aOOP50TNco39zwgm+hvNbK3i8ea
H2icDaSvoA3PkX2PXDa3g2iq7fBwA9tE86hJR3+nI6PZ13F+SVXvSAbrsU/w7Jxr
qJrW8xAwpjKYT2D3CKUjph4l78P7gy5UHwlA9XTkHPa1jOcBJIpoUbazIbFHukMp
eSaoSKuNsSEWZMYAJOrYd7mobNjRuGqAiaPd+iPlGkOmzxLpq59eHvG1zBVLK89q
SsE1psKtMBpI3zu/EX5Hbq3NqQcqT2kdM8Mnrkgqbh5qbfbxpO5++XChfOISjhEm
OMrk0RKEPSkdazGdx/zFC4mmSh4J8pjRvogexHGhT1wHG2HsIRio+j6dAHCjwhCu
sVMz8PLs36SDbCt+4+wnrvE2Avaw/7MTDCU0ke1Hfn0zkNAd3koqDfK6kERlAdkg
dkhHcNv3Oon1+KN1bExsff+1YysNpVI5zLUk2MpdfVSMquCIF07sKKCMSbjOZJ8o
lUgEB/QcsWpqrccOlDHY3bB8948H67fdDTFujAqJB13LhK3clJ1GXmYOnGzERGcn
qBUHAs5e4HV/jCT6gIsLEv68YYF3my1BI8+UFC+ggEQlBi7OA42RRhUC9W+U8qzg
L/YeKlZHnXhpBfdTYDJbpdZlsctnQBsai4to7bE7nNouhG8xH1JPH2WgRe7ZA7Du
ODFiGh0ZCMFoquXMtxK4qL3rzCPDdhE6FGQ+nKOZVwUgv7BhPjDv0DonA2bYbBnP
i0659qaii6ix3Kgq9jV3Ml5znynxHAAo8y/ifcXypbfTIVIgDgWRnjeh655RzxdN
yfzRkk7d8cIDipkQiLvRbs8OygOak63atJ+bWbxtCRuSe4sIaY1O7y1rUfKE/c79
w52/44mli9oC7phh8kyrWL7SVBqKlwMYq61RCoB9WGRQLWf6uSYMaaLelxFgT8OF
O0LuLCZ4wGzPzixA3ya10fd6z30NPsFJcINlyQxZfNQc1VTn6isISzkMncik9dSv
AbQ87qoF4CZqRCpYGR51+FtacIqagmNshsndT9HaTxFck5RC8Dc4gIVzMwSrf7Hx
wEX6IVqvu91Lzi9C0oNrPWorvt8ujKKnUgJbvJshg4I6NHNx0wPGOBsmIb6j1vuV
vVrUMTTSeRnIw30ThYCG+s4GWJBUhiB6mOisbPCCB+YY2XZDXExE87nDhUTaGdQu
90hVjam4HVOkXqPdFXd96/BT2Vxo/92kkuQcu8EHHVlGLnh1pCf3AfUNYr9pgbX+
rXdruldTyuZq/Mr1c2caxNn1tFFfDJCEXDI1gGiiZ4Yyj/rxIwmd7hsZ8SVtebTg
WfO+QX5g+wNofvcBk/9BQ/NK2aIKGC9kWT8oTH9DwSA7/BKSdlDAsb5XhxlO4oXf
L8u78x4nTll2fAjCGQR6YyORtnIqixzOSlREJYtsiH22q1RfQmF9lKdc903lHv++
xYdWZz8zzjZCXLh/Nff966UUfNPZ2b3KqhK/oE+EqUrB5k8aEkhrycThB1apVyM5
r529SycE2T6AfnnWvoJU2WYjIto7FlpVTqlwPdcjsE73LA+81FzUrVV5NSxNs0uz
S1yvpyvqEpYEcvxWFB972SdIWP8MDbyqoRIIJii18x9tkL7S1QMraZwT7PeA1Wc7
V/2k8QuxuWrp/RQwLTW5Ixz11AYCI+oZJn63EOaXl0l7uF4+SdoYlhCWZ+PdBGzu
bjrPtH/uyxUbY+aIlX6gae9xcZoEj+BAJ66s6SGy01GPbRqSsDlcYh20gOKSHX1P
LZZ3snN5HSTScGRwaUgR2zOh2DYwiAQUfVXRcCJeU8o5D1gEA3d0twtwwmT6M6is
rA4tKFYIAoQ1Elf+SSGNkFWA3ahIjrFQakU7qfHPptoTVugNtPGlUBEQRxCJbR8u
h6UIAIVXsKx83Wxg92SlVxqXKNbKg7DUJK0ACY2qjT/X9XJNQyFV1Ab2l4kn7bF6
PaQpfX7rtf5gBWysF7WmwRfK0MieVJrh4cZT3Ba+yLbrp56N7KGYzDj0VnDljnvL
vzaCthrmdNSQwtgZ6xXyfSN/+eevrqhpHuvEJpKTcUTZtcun6WMAivIqpw3KHDX4
r8fR/SRPGp+p+WP9JLvJ4QSBoA+/3nHzEulAHugs4WP+pUwGMUMvfYnVT7ctRUmj
rT3yukJTfyaB/YNjt7XddQjwaxxhf1aJVupRDPgpQQf7OU+wu2ufm3fpryMhrce+
3EbzYJdNwwf/vnL3IE7HF9WqD5wKmCkIHfFT0/MdzIzSMBTe2+hATKuNmYkAiuGF
chMPOS1bv2oRu5waJCuLoN3AnCqJ3mOUDYW/2y4Pfyxr/8rjZoLFCuxnLkfzw0SH
Yn4BEQQlbYixh0+KGm9P8ARKvONVqg+GpoChA/gPX537Dw0KEfFmdA3YBWIK8urB
eixQU2IKqCAVu7Gd6hNCCcKhEzlSUTHwNxUkZ2YUFyYqZ8oY4ye7vEO1lpz6Kudq
FvZObHGiOi59Iu9RxsEhVE8A08zz/AjcScq7DN/jvxWtXyTEqxWSHQWqUsle6ljv
p2WB6MmlJHHTiS/rB6OCOa9CBlAfxshUFJcEl0ArfwjBGJ+1pbdxzwu18ZsZD6VZ
EkSr9Z8Ij9JovaAaTTDudf8xrS+TQrKzqLri5P6q6pM=
`protect END_PROTECTED
