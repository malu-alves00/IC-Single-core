`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dYWhnOZ2GhrlVTE6BIAIU5IHGit4AYDBXKo4oBbLQspz06npi4liPN1PhNLEQXDX
31gE/wpLdm5YPn75cRNV8aRrhk4QmMthhS2RKx7zdBAVEaGPG0M/twUxT6FTb8d3
3hlms5zbt+7d81nmwf9eofeJ9qPVtn9rq/u6uoUP/dU6Ty2xOuzCG7X1E8piwnHE
StI/J+Q+s5hWBle+QxJdSuadZVjXou3MTfkI5uaL4X0isz36x4+lfSgn4mjmPqW2
5N4x/U/oPkcadKqmy4Mx6VjZQwlXxO7jG9sD7xgwVBfygUXuYWAp3tjrRfXLTdEg
TEabjK4jiT97TFlDLvDRU06D83upHpC7BnEGtcudxj/J+TV3UVdxaerc75UufZ8d
FWxA0gxhz0Ywq+vAKF3mxpaSVog4hnqugt45y4k/gmiAfbTbuUL/iGyYvUtJ3Hjs
2AESLVi0n9+6xJ56UBfdrumeYFKNt+pvKfR/omHW1SWWQORIPfUbr9hciHft5P7+
8leFvTwfNyqxLosjAZphAXxk2mzhAQHYs6VvoxOISaYe0C3OqKsZIueH7lzNegDh
MIzrD9GIYzllkJwO7JKN1hxFzglJazSM9hSOuscLYDBz5EnnpabTcPT315EQ0QCO
a0QHBx3SfHXyGij+w1sZybzSlZoxroHy3EG+/pMds8b6kth/WABGiy0LN/bqDnHX
yqiGeI4fF1Ob23noPw9wTmNT+vF/bcGXVQ3SNuTvW1mpwRGv/QppABdFAPLkl5c9
Op5JFdounJQ6QzPU84SOLg==
`protect END_PROTECTED
