`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/GaBjNRpKPiubgJ4DIk9lih7q8kQ+RLYDO1+oJ04oe8KNUZ0oYACbab4P3voRAwq
5x6j7xjyaMD9Its2A4YPOnp9unWLlWB9FG0kiWGtpJGVLn6ypglqqbi10qHEudKP
XGHdoBaeMAJce0or9Cu8BujxpzxjynKfR/mekxLN/5lKV+fYcQEISjo0/ysyazu4
LafXPu6MX08NSbF6U+Au7E+69VJfk9VHBphHABhJZKkUxHZ+DMvSz8GQbRwb1Hne
WcvTPJOZ0x2tFYqAPSTC1SVvUh8uZgA43nPomr4KMzqIx+nnavqQc8AGCsskDAv7
KqkHZwxfhj/fCTCNyu8J7gq9TRmi/kRwOrmNnkX6fLf1zPAgUz1O7QnUdXDgjzyb
zt1AmlfRd+SalVyt4KZhCK4D2KsUQJZ87mVTs3ruRT6ipp8xuI4VEST56ZvXxWuc
7o8dhKeJE7Ixnt+7v10Of8JXZ6KctyOnj8uESteP3wq0pyWPzC6LBEiVbiD/RShD
r168XICCQ1tNFLgB3l8tIBLfe1IG3TYGs+HS9iPafv029PCfnbihqH4n8tc1uYBw
7NJs6602sHem8wUljQQGOvAGoRbQjH3Jv2BaIXRyx6sC70lrRd4MnDM39VDO77ji
egplR3FCjIgj5V7O8DUFr+eI6btwn38k6kE35YNcBz3Wi3i0GMnU5R1O8hvPhmy5
ixqBlysZIm74b+0Z8QwhGskqDiPmZo28OTb0aaMDtr1CIP2OkYRxlGVSUxvHaZ8I
grEdS0J11aEhq8L2+GygGV4lro+m4lJAPYg0cjB+ZE3FbfYhIlJXlXDXvL4mWf5X
IqkBTThYxz9ELNhoQUMdXIVa+EByTYVWTn0neZJTf5ppl2EEBpSSWDhBs+zwacmu
sOO2eWU0eY5iU1/R6Lv9dLfnA3uw0UHJb+A6p8+m4OYqNREhJoju6qHBww1zUAGj
d78epByVg+FzapJAV2Gu9aBr9eHxgAZrLP2RxeM6AmR+psQaJC383DNTgSSjjhB8
6O4H+ZA+9tOWyisUYz8yngjks14ATqLZ+3rXCnHFpBo=
`protect END_PROTECTED
