`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ppnqLNQffahA0fTMTpwG1WJfCRawImjrMCJsZSWxQgHllA1wBhlLruGHW9Q7QQZy
8STGG6IRmuraqvDAEujsT26pmPaGAm/xyc7VJtD/CkIhU41qLdjZgP/kn6XFB9vA
ZVa+/OkWN+RK6mRg5ITpLBOsZGF794z14UUBQS+glh7OJq3BJP0vbCNIwR+Jt06G
uKhKzLT6JmjTg68KbiQmudZbsFq49gpwj2KpuTMb98nNkjPH2u0dtAcl+0ymszp9
IJHkcSLFVki54YP8qxlxSwH6C9xaJmgiXfW6hO66kja202hEnWlZtez9QZdltmiQ
QcEDBP6MvTrpnjnyFAzloRL5bQs0FeuJiJiZhJbExRnipi99P+mgllvNvAz7wcH/
xE90n01aln5Ndd5rOWnGrHKH0WqgvkxdaPF4LcJ5GI23AZMinj3IEFkV5YLl+v0h
S6u/MpZD5snYVliepKOnfDkkjseMFd26aEFBOhFhS4PW4KOigrTjABkqQ2M3gGeU
84/VJ0Fa0DLDTGm6X70KuE9TkqPj2zwkv3cCWLaBK4WZH+tf9eRhQ8yOucoBPUTy
RZI/YChiGefsKpR37JrUHu4CiBFO9FMO3xv/NBdOB9zbL9bUeVN6ahocsrKeJlcC
U/0pXCTiWIg1SfsXqR8k9b9OVJYXD9UVLmPxVGPxTPhSqNtXCpUlzG/vxlt4K70Y
XJWE+Ggi/fFyVEv1UX1E+ZGO6zUsXVL5NF4fS3RM/v5bO73miT0frUEn3Fo7Aoxh
NN+tpPt3yWm3/seHWM4mb5YSY8AT7pXyPsigCfK4i4drw8LOrSWf5pDHiDwj6IIK
Q08hq+aOcIhxIqiS7pfNuuo5wcpPcn/MJ1ZUIGYZw2niRsXpxS/41D23r+qJsv0P
aMuVUhMid9Fg1KXlOj8YK23K8pKaXtBrthxQxOV2zFmHwOGMGFmD2ziwES01QHwx
i2irOBSEgoPtnDssh7fAjDgcF8F6U27v78KIPRNDDfJdceELbhqnzcMC+SBhMGlU
GuNXKN5unFGXibSxrN9hG2r/hWkV4g5Ujjx1/hZiCaMxZ0aG+M18ab3IcRqVr7Ji
m76eedGuA7Tfekws7NugrXW4gMsr5kNInbDTyQXRnnJ+QTOBaO7e+4N+jnUfFEoO
xwFJnsN9xRKdaBuT6iVV5EOCo7gGsIR/eO2R10ChSJKMZ4CYSnf0sHAX+DZtlMfz
R/pUYempyGymz1wFtLvZitTQXHFbd4xPiR0Eu/JgjXie4w2tBPoLHpDEnrkz1RD4
/UAiPqNy8JZRC4tBjSTlVUf0NFl2SzUrBTYcrrBEgWdidmN7jAs77cF5s3uDxeMR
2QltTeBIdaCtG7n9MUGG69RiZ6FG+v0QuGd+BNQMm2TKJ6KpS71nrd4rYCwdFXTi
S4e4vGpcg9TbQaO4EBAAD6Qv8AQwc8h69MHrwzI24/y/mcRdwtVG0f+r8C7CXwKb
CI/7ad1P4jIwKmaT/qcn9OcHMYVLAiLysIXf9gfK9823VE2+SsIPmJrmNBOGrB47
Eu0xNax9yb3HryzgQiWpJBa8ubQ58o/C8OUioR/KNyaE88Dz9gMRiZctbbSmPkzH
pv7ijtM8V7d2X25aTNK9Vrla/h6ZS6cRKb5liVi6+vjc5AYcRKu+wkbYZeT1m2Yz
ba4rZzBdq9gHD/BSKRzW3SP7YGyxV52Wm6/+vYpJslpc9KmW+ErtP46EO5bZFUPZ
NlkeZdNqcyoAPRww1iN5bevvbL6E/WT0cniIkPAquhtP7wfABlHxbNprovyQqj9t
TgzR94HjgA4gDFe/A85gHWIPxpaRR3vZAxOFQdlLEz3Jo9JbimWr1cM8I8lpPW8j
1qoxTKoVJ3VWEodSlGZIAWG34ixDniNzSvFMt+pJ+cjb2TypGZvjXbzh0oZbzgaw
Pu1pxZVwxf2bZhXY+kN+Q+xwKTXM6ORVtD0YNSXuOHj7HjWUnRisNxFmp1bnSUMG
wvYdekR6gcVkJSZHu28n1XXiv2zav2Z2tN+nvIy+ULbqy5OwzS8ZL+X0vxKxi9hq
9SDUSout72DZw/qZCYzIUqWtUJvzU/NZU/qz/pT1Tv0WvHblSVdUdJzjyalFf1IN
W9IU5y2ZniiVn/rA992XXTH4twA/DMJ0+JbUtCFSNHVQgEBcuAsN1Pn1m8Ke1R7O
0uUyw+LYZYaaLen0LzZ6uz88oaGFLZOeQT2aI7c9AhYxylpVhrtCj0ZbuQaqQ6ij
KneEXEm7jIMTpEAz8mlUCbM0R6pyZvazb6p93WHqUnhMicnIm211Gk6M5f6qmxHc
e2vdEmKQInai+202LTWtXr4OiyebylHBVoQG8WnML9UvOSn1J6iObhdkf3GIBrGB
sdnrRsFbyY/k1GkafPCr7s9gWCbh2IISwyCJHrRi+3k1IoS5cGZDHC+cJiTJ0g55
iD8zPXXDbj3GuIo5qXu91nJr3cx0/Jh0ZZW1C/J9IJiw/VBY0EFJ6rHO6Sc2pvUO
YLNszpyNsIbVsLPfcdzE1OI0tJCdB8glgmLu8Gzxj3Z1C1i1pyye8sfWv8Ts0GFU
eZD04AlRrtWrAOu0xOD4fB1hq7D43ioWom6uWMr3n4ZOkS28wojsOv88uqryUmDv
8osyPEdMXJbSt8gw0emPp3QkAnpeDWCBmsUt58YDXrN0Y5pwBNVGcPF4lBSAu/8n
eWFLY9ez/leNwXkEDITf0N9doOIAmizUqIlQP9vtQCgERKIYTBjFrVGB7uotkhzC
`protect END_PROTECTED
