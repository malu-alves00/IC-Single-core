`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AocBsy2+fF9caJCjwXiZP/ve8LMh8rHqt3/dXE0jzV/bj6x+l02fgWjenhyj+lqA
3ZirKZ+PVRzRs73igDsejbnGxFOz6J+uK4oFi6A+Z3lxB6AEl4kLe/BMtkIpWFNY
PCV2GkWrGzvQWlVfrgApLyQAF5wQJtetutQhNeZ/Vf0tOztk0GArOhfeuq66SRJ2
Zq56jAmtyaUtdaNcwFJCU1Vhe4PiR3S/NR6Y8ZCGqrk6CfnWeOGxCcV2qvyOuEdz
mY/w6xJIGsRtdsq3pK4bXMb45KzoeIujIUR40kt4WNPVzCOzkyB8EEZdNVZ+Ild4
/MuIjvfM0qEcoI8eU6BWJ+BWB9YJIx8qLLfAwy3dAE6D7Jzlftr9DxXqRhZH+HNj
jiuLJbLE1Fg8zoXTxHlMaKsjHv/o4xcn/bJTgUKKNdLuQzNxhkmiVQ4rXwSMpcO7
300D167UqhTW1nGbW/akNIwC+KNWPRMAU+ai9371kA7LUSuNiB1KQf54QfX7yVQ3
pHISjAvG6V8HV7Eg7Xawg8xyTxMuGgz5H6fPZoJLu0e2CueGGuW6h3wl9JFTJVKj
i0uC+s4FyiF6ZCZONo7orFZDIzbJgPEpNYGCmQ4eCOKSFSgHk0KD8wajMdNCljtB
3JP3j/nEYJdUlwFUkOIgXIKLcYCEVzlnAkyZE59803SzxuRYx2MC1YagZWsS28bv
3dFHXyhkN5RvK2/Hzg20BwIFDyIH0daK3UHOWARArKIpjSfr8Pzv3sJRLjL0A+8L
2eWIpqsLbuwEstD7WkbeQ0tzxXy4zuPebsMyR39eRwljzx58tkHaBhY3lOc+Phvd
aU+S33T0AMp01Ts6XbmTucL6dMMJPGE2oOuPaZU3crPUUhV8CglVjMGIFFssC0gf
Kf+DxcJ7mK3YbLvJ3AVKChDltp5WCEfXqembpGpytTmFn8VhoIHPN96agDUUU2VS
IP3nKIyMpmEWMiHLtc0juA4Op7flLO6YbGg+Aw+FhizD1U29zCBnwerffrDWvyeB
uQXjPpQML6xGMQXLW3FmvbczNV1gDQP0AusaM0n5D9a5dMEm9gdMAf6teAzASzIt
F9O12dBhtIdNxff4rCef6ss/09yfASkbn+hfJE2zB/b0NvL0WKYjDmEyzQwibJ6A
ut21lKyivzBpC5/adLTGZOTn/wpeTqSCF+pOZxMDSQS95Er/HrURRH4bfLvJFsCQ
IPcOk4UeK7/MOfY+mwMGgtCEGA5NEwp+oLLMXVrHxvasBt8mRzSabJ99LdV2GVHS
mUVxN+74fc+GgGz0MoZ+ehfKKK4tcyWhskoRm9tjo/V3edgl8hqbZxvo3AOFa/y6
S7fCdXEKUQGHXNhw+H0yXBz/YdyANVBBjBHvjPxhA6SyML0q0sm78a/ydVbld92L
lvgIIY9erxzfbyVItRtWqGdGacPnjSx+1VXyQMyfntRIdIVW6IOC/4CJt4WNAWT+
m8PWV7eDtMFwqTmi2ED/sMVsjSHeaicosY1WnELtBp8tVakgUbUCqVYu553lI1tv
xDhxzOdup0WsxI3dM1s+EZdtEAWBoX04if0D//SkDFI2l2OpyqWRtd6sjfQLePQT
kGd+HSMxDIFofSCaX9/uOGJr3mfm04lqTmGW8cMotYrFIC/XVXkHzxnIsFsH4yDM
8cNShnVeDTV0KiLYdcdzbcRpgIQLwifYqtOm7T5RSqyBc6jsa4URUv7e8kVjyigk
JhJu4eHIXn4wXTwAeSBZJbESrbgpM5+jdvKLmv0layWHV6NRz2fe+F7nqe8jI+Qg
pQoHi2Z3mcb5qFZqx4aUCy/1hBveLu0EvcabFngPLKwCPVGYxqhTNyFTs46Snfrh
5EkoxnN2/D9wJ99yyEd2hqCbwOLuhwzsguiTbxekTP93J0juyv/Ak08OjKhHsYOs
V7v3vz76Ql/87LFbSSRkWA==
`protect END_PROTECTED
