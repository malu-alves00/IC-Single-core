`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Du82tzWMZiVa0TznizGrSUhZsSqhoC7ETxvx5QAYdebhk3CeLzoNXyod7oSl6IGS
2VJuEfgkSdG6GiVePB6kOmoOiRD3Mp+RU38t7t8UJckHIV0nWgihsws9coKaEYpA
NuwHig1eOYAvw6hyFVq20BQyuebzWYvlgSUhsdgDmqsdhTXAT0RF7FPl26G06WUb
gCNW/omr7SGWiq9WI+kCICkauQ5jm0Bneqzk9Nfap7N6kxwzJrrfZMjb3/S/glQS
jd4f0KgI7x36XHimF3GHEOXZHMjBhx9ArnLPjxT8+jppFssIol8RrCa8PdpdhXlH
XIpujcyJjJuVqea6cTSzRUuEAezrHmuhzNHJxflOBazUfr4hw9+CIsvLRnpOsOHz
l6p7P2X/N5A2XiT5dKuIiElz5cb+V0LRNFu2SSEhAh5o33rK2+LCN6nQvOHumEqm
MR2uUoq3mwctP3fcx+tePjIqueh8qLxzQ8sf+7hcmQ6uBB8TbVyO0eTDOqxGviwZ
f8iB981WYAIf88mgrMl7+62xiOZ0JnG1M3OyhebY4E/YUtDCkjprQ5S6W55MlnD5
fWB1ijwyBYOxO6XLOBww0U2fAs+OfX8eLf0sQuXQyrN9d4jAEE9qo4u1gQsEb0Gc
ngVXtah+nq8eejqvmRJyIxkppzEhQQjM86NPl0MNbCbxwWxVoKs+Q9DGJjwg4J0f
arrHAQSYTulRbCI56VL6N5k9xDkaPuqSyix+C4Hwwn0I6BHbkxTlNDMrspyEEcIm
cJKrL0Yu+3tBcGgypLxPwA==
`protect END_PROTECTED
