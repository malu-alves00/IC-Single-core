`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4sb1okKx34JWlwAanaSj6GKpmOhzEMtrTeFzrmrSN1cmRcHlKXVTc6TWLF6D30hq
8e8T/Em5Ryic/Jy9FzqPKVP2o7YYCKrTiyWhmX8ebFEaPfxTXHpYhcgfEtDt0Mal
HrDBbmOy44Fh1KQT7j7qFPDDKHMZFwaJIl0UCawVKK+DfpZqfkPEvzDj7DWbiqs/
08rl+8IkZ+7u9U5qQNJus5/CYWmxeJuLPy7L0eMXCbxJuwc+dHgzb97Y5bdoDGlc
5z1Aidt6RhhsPFmbc4nnXBMdyQdOKLgqp8kUbpPfwh+N/jMGwmkKpctdXS9Hh8DY
i69hB2lunMj/265GsdpPMel0nEViaD93C2Ay7QL49ZEDXsnW2IvsM3kXxx2KV0BX
VyWvdxLz161fMhFlhwopH0H2owAH8PHD2OFjzrqRsq6J87oW0dqby4toJ0BlUIzr
5KdhCb1heSGMPFEtZMODxqLwOxLTSdN963cy17lm42BuHJR9P1831PdjpaGbua6/
90m7Z3n8cXCvUSb0vn1juymUMzCgWzUxmLy6blM4A407mGuNwaezRSQlJSREGAjo
LoKU9cb++8HGTQRNxB9SZXiPv0+WoARgotsqsq7t5PsRDfwDw3661YNbvkjBweH+
tZ1Gb61OCnziqenWEVe0RboJpHCQl/24Ck76zT3tbxzSRgGUfax9fWJ6MEMNdPET
pmtJwed+aJxlhmTifTnW4rZUVpvA0Bnr9QlhbtVezYYPqWHu/F5yyCwbRrCFgSss
kzJdL9W9VhzRsxyGz0NzBtrhTus+tFKamolM4DSkVyHWiG6osO9LLOZciKRvLn9K
B93ArxkakKtt6j3ASKdjyo0O7XgNLS0BInzCg9aNigsFePmrCVvqf3b6v5ZZZkM6
ELAMbIafX6Tf71GkgqmUsfUyDUOpKYfahd+vZiSTMRFua7QtSXcoqk1RzSbZYz3d
cERRfKwKyhu0j8tSEazxoKndjlyECZnkxRkDGI4wAdqe9UKB8QaSthDhGiUpLXy/
6ayiARK/QywsmHK+Rk/ZssiP0K4QAuYluFFm2o6baQonKOcIbbSBBXD7XQV/KqSh
isosczew50pwbdXnCMKHLXQiGjQqU1+UvZ2qXQ9mvSJE6ylxQdqyPwBQrBpXx/5i
rsc4ndVnxhWte1PW9DydOvrmHO4b40l9y7alAQwxSAdB9oZ8Mo9N5rQ/7FCg3L/U
E4wQfgJ4JDOpGkyrOBrFB3aiVBX2ZYCNKvaRWdKPn4MQ9GiTg8FFVMHCX0eycumL
cuN5bqRywkQ/DCCzRS2i7Kb1ViVXRpxzzyo/cgI+JTj60c93XbLvzSeaXN8xXFc6
dLjvk/6LZG49mUlIHS6rX0Ll36JNrIkTOqEfBsJxLbMUr5MZUwhmltAwVGlcuGmL
Wbsql0I2/aTZqOwtpNxxt6c4cD7Qb5ATRviVltF/4IN9qvAOvTZ6jh+aY8fkBX1T
aK155zJa3FjSeEM5SLUE3YcJ9oW8Ynn5fKU7ZXYEcnvbIIKuC5fvKU4RmBKLSUYt
pJoFV3gukWFUiLgA0B4k/LSKJ+P8r8K7eF0ygYiRFjJHQzpqkuC/yTS746VmSQgU
A7XQ6OHKUBFOcUB1wiC7ZGYVFRUmzYC0zFpGa3Ufxgn6H1rsphuilS6QZ9dw8gZV
ZNzZWiSu9UW2+WXx3y6qrsH6IVraV4EKm5J1qduJEaJcKTn76/C0APi4NguWyTGP
n7KIJtS+15uPWRe3KmAxOqUtaihg1A1nI5eGccYnDzS5CwIXfyWytl0+kp///OhU
q1r7Q/CpBPYmqRqPuzlt//blrCrmKubTMkw5V+U0zOvrjlhX3Hibnofh2Cq56Kp/
c5R7gZmXuLzDD2/swoZR9bq4tYv7TCgTuib24sKeeqak6BccdkP11qF5K/wm3dZm
n3ABk0kKN1P8XJQsav5LKtv6SvVv0qhlZ4hhilb9W4MjHNDkUG/yX1VA/ZunjyKy
8i37hC09GUE0SabZJjdQfQES2gE8JHdle5TlYCrroYltlGrqh8BvdPYk0og82rSA
ypjSCQKOl4LN9We8NEuJDqeUTb+N+7SHqiCm8xev0GLdVL0zuhN5YHWXxh7Pf5IR
8Boro4r3lu2ZMyCDPuRKmPC1eSqiULh/jojWiPmObGt8MF/YNa2QVMx7EAA5gXdS
dq8QavhSH75xCRWGIeyF7qic2Hd7raa3AVmVZSuSRlt6KIbhJBA2x3qenNVEed9g
yRLpZL52G3Gtw9fh3OgNltS6NJasD84/UebCW3/T1No=
`protect END_PROTECTED
