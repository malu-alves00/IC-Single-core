`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5Q0GeBPBw56uey+sTIYjJhh1AS9uyC4ZBRv2nDHc3yW8Y+lu7nXMyb1RXK5v24cO
WYpR+ymQzcNoQaY3kghI8+DAXGWahkjucmQhGro3r2A7fs1hf3rX87JiuDcSUhtR
66N7D6cCzneE6FbLKu8rlaYQHwPNafLeyE2led6ytNXnuFkC9XrgP3cCUvrDu2BW
M0whjXJv3u/AJkzrxw6wsGLe7JjZtnSL7KbKGO+lQwjxYEphR03tehDzipv0DouP
5+ChaPda07/6nt8ncpmEViawpuuX0VUm3QGFljFYcF8zOO1rB0nHMB4k551W32Vx
ww56KgC1N7HE+Vmyi/2hz3r5uFGFkCmD54mOl6vjzoNRShHFiy3EIkszUTgIcyMI
fca0ax/q39YkAqSG+n0ZBvKijSG0t76IDQujpkxHC/CuVEMK8yD4zGH0e3WXCDBg
/nihYp9fi8bf0fcs7bizoPR/a6tw2u74CwBOsAVH+8u3Qr7H2fltsFp/R4SPYPSl
rE2DISQSVbEnmRzApohz5tYdzPxQwnXlejRIeoO1X2a2I4i1panV0k/7kVvL9++U
2hDsyZSsD7BblZjPjfmWVdxTl46D9xPqfwFz3bTglXHIZsyq165KlsnB00L4zqGQ
Y0zTL6Zbb5/nEBJK9B2w5+Gm4XMpbFMoJHR506Rmw6bJ2AcmNeR4QqkBVacafWyi
G0tWv0VgPIoYGhmnykCnSfiDonyTyb7A8OhQeFUjfjT16lunrsh0nXma/2t3Q90K
b7UurW45vsMuzZ2U98uTw7QRJCFfW5Inw/6KNyeSeI7aseRlLvlmgGuY7NnLd04G
kxDJ5kevItLNjkZmA8E6jTEgXRcR0wBuebadR0hAjUSFHg/RuugxU7zZaGlBbCDT
lEtbnErD9NCOKxChz0uWthrUTUjWhTV/Xyw3jE2oW822PjsA3axl8+EAD/9R2dr5
Cd3kjpWpJ1zLR3V/CvE4suYQ1CbTKGZdl1K09/XwXRUEnVTRCx8QrfDA3QZ049In
I1n1AKmW68iy2XAvqwVZdKui+4YGwfb/OPPiC9FRrymL0maQ6FbgwZ1k2QDxsEtX
L8E0y9pEp18wLmci4/8xAl6RnGWPUUtXGfX47gtpCBRp3qSS4gYzlCshkAKJvdIl
CH4Fxv8I4x57QdIbuEG9R7etw9UjWAB5Cs9HJvsvvtDmD1N2HPDHSOKo16fkESo0
gpS3Xns2OIKmRqawGeP8SPVStt1JL7s6nIBYMOAopBIPhmg9VA16Oj63UGSOV/y3
SG0rYVwTPL9QNe4MgT6M/2Bi1PBVYUK/MjC5sPubSGYC/r+zP4p7+EgImb9IDJl0
G7f7KmhQFvi6aIu19leICFFTlSSv2bdhMU8yGR5JrPyp18Cf7K4Eoff9JRgJ0eE3
/+PWlteJuYkeISvKzJKb+4fqHiY6XJglhYOH+C6QB2zraP+Xa3BcCYWUFfgjm/R3
swbNh31hNRGr50uEfsh6UUNeQ9MooQzP+pmEB+SshXQIYvAVSNSOx04/L2C3sLq1
a1F+wqY2VRT0z/fRn3Th24b+JJ5IcUbt9nuP0EcM8ENc0S9XSUHbysVgkzCjMYcT
iPpa71HB7j5XDOoGa5z2f1R+X7vqx+Setszl76Um/+jPjj4IIio00v8YXKS6e0KG
QLcW/+ub0/0BgUYj9iydWCDhrsikjNQ26ZsuWmm7WYDL109mFWYjHpnB64y1jgOv
DWCy0n3y4RipFsXh/NOupq0YFnokeyV8ZjjhQTklVPBHuuXSOI6egubDktMoJNDq
AwKcUUrqAcmIITj7/AtFQtJYx2pP5/xJCsQYebkJIcxehl1lavaez3WIqHW2m3xG
AaLSahsQF6ACD2qKUVI0cU0XLF202RIT0Z64jkrrItzr4aiRK39uWXoP8IgAUUX2
FJVjmbniyUVfXIAAJKK88Xo4COqy6CdvwV0xyVCgQPFBJ+bwM9yGdQrGIyr5nW27
VTV6kt/ihbTXSv806FSivn4PAwOconPxUsSmyZ62Se8pAD8QbZNSF/CBoYOsuYIK
4IfdQwoSMTQqs6h+UCKjgyyAVodSYUTcMO02mermDMdOzS2eD2DwoghpxtN4JM8/
5Sbn0F8nSGRWUxZQhyl/n/YouQcNB3SENbH6NM6UXUx9JFqYy42KFAZFFve8ubCC
0RkOFkGDwGm9bHWn2cBnOBYD0s63KOlMbEKHywvNlB2w58sljwCUqGVpk7i7xspe
5dfzFjVG6A/a2maTzbTkDGJu3cXRLkKQnOt7jWYWS2fQu69liT+tyOGsWbfiLIk9
6EZpB7zmcABSIycPRbYWVotkccF2h4Wfx28A9SpifMmh5FgYsYPc7JGqndxvNDuB
OQXlovdCFrwBeuivXyaY0XRBjCgBqq5CogXltMkATwHRR1NHr0p86yerlmMPPlom
vnbXoueSgZ6AxC2aiZj9+9VFIgY+0HqIDjNfmgiVcD6B4HXhXptJm/Kr4ubB0mWm
8WD5sx7/kuTOgC8vDW3fVe9fyLkPmdH8rqjw+IJHW79aB5kXmSWAmSSIp1TnZSLK
N+dmyw+xFpxMeeQJinXoLeRxbkW65AFm6ZZlOpJD9IOYCfg1LUnzOoQ5fkIf4vtF
XmB06z5dQNN2OQ00gv98fv5AAJ8rZRWeWl/mq+WNzyQMEXKwUZXv3srFPLW/4zIo
O74gu0JqlmRR8jGg5MeY4bsms9GM7ptu4HemutkHJBK3g+aBcgfAyA6Mh6KnByxP
PtezA0aRyS5/Cpb9FEIGTLpFDf/4FtbBd2lwgVXYPtwUu4u5jYKF4PQpBVXwMTs8
IAHEEXJm8tyAg9IB9sQ7optl7NnIvp+S2Ahuq20VsiBBdrYxmJ5kViZ3QLrTLQ4P
wzK6jl8XgLq9qfEiBCvhOO/Itx7wRkhnZShKQjfTI3iBpEbBOaJ35QME46CZxpZN
/MLtYU6Cjyx6BtFLjNwXF1r4bD/otOMHV7sK09BjiOR/RNtq/ZMbuUNbrcn0M9ZQ
dCJLNjw5oCHvqT3TaTIpQ6tMxEHCfuqmzDKotMEcxWMACPDPBpDPIsLpZBiknGVJ
pteyCBR7VbBclQr5H2LgGBbGlCd5JF0E6w4I/qNOYYDuJdmmsILV28LE+iAdVDSM
uNo2xQbOBth1I7+wzFk2d7KTnLXwxeKMrpsUEBzzqFJzsUlA0fx/F7VPlMr6hn8x
lT7BBRsLTzF+gi9oLcld98EqsUEEcA1u1nAB8UhuUOo1TG8cYRmp1CfkgZuS5rH1
qFt8hnL16mMofuFUgm+x4QrXR0Sd+xR2InBWtsIVE/k+9hzW+dcSdC217Sy+qH7V
Wb+S23TZDRxIeuwuOgKvThJh1aZoZUbONizbGMBHnXByEZHaGcYXugK6TYCbm4ym
ogbRAn7DS7cztkKcRXpaIg5qDVrgado64DtjTw0ld5HTng07GkEWMrhOmTgueKVm
FHekfLfXBckuvr9GAnqnvWkc0nrromoo6trWtRgAH9qziInJv74yYrRLqD6VxObT
vcR0dChljc89CChRa1+4Y35nBPdeF88KWo4IN3/AoXArLkwxMss/fQgRyebMWdak
7QWcJ1uGM9LrcSkbhSnloT3uXhwptMZtWui5BITO/L2e38p/nWiXPql+XyGFwsnf
ZPCLv9ZDq4pL0M3T5Z1me6/iCSwuBLcqOwCKOXLkCrxH73eyUExjRUoj8lxunE7s
hiVGOqH3bFlzMjupXwE7cCuzV+TOOF9bnMGSSl0E/rKkXMDbbXA4YG5sqXIuvIW+
cuSCk2zMKNVZ95WBaoNec0Y+DgZvOUr8OcUAAJ/OwvYYJxPXxRC0R7jCil9kGdmz
6cr5CzfJAbCzM/wiRCtoL18iwX5YnEm2Wi9fUh3iF5FU+Ze+5Hno8tS3Sd0LPBOY
4Xh6VUhyANJ4PFgq8B307fRKfYclpSvfP7mA7UGtRojTcqDuddn/TDJXsTDCne0r
bMJAI7xSLDN+PK3K1m7/zXhv1AsuZ3o/zWGRlmf5e583R+dXCLxNLuBoDc1KWoCS
nHTZguHxvHQBWmZTSi6NNkNp0DO2q33kVIZtWu42P9wqCUUT3zNTzVVcqhrWul1Q
ejSLySjdiRkpFFROyG+Yws5QQCxaoJQ92A+/gMNr8QnxnzAr2erN/Y7sR1oeBLxw
cX/ITeIP6csdbPhd6RVLxcTwBeVQQnRZx9fUXRjUAma8LKQE3RLMWUv5uaZMKMMG
o2XstDoFJV8XEpTNsMnjERtmIJL5v1/69ngB7LuvBUdfYJ5blYbfwCAHpTNg+tO1
2vNHevUz6f4eAtuIkmpfvxwniZGtPwXG0UsYzjuZaSWj4NF6j3ipcKo3kgO5omhn
WkWPBxbU+rbwrqdBpqaP/8T6Yws/qJn4ladcSRXBC8xt0pjovo6ATd/T9eVYVwiq
h3NJ8XJ8KfUSirhtjCAaOb8iLQ1Ckj6lR37Y694fm+VjWvIEHdUqojZ1+p/fN6q9
VNb2uzsIWEqjzvGmxzdGs/nXkNQ+8TSpHl6gXYBgMBks9Uu/UiyAJHflNsIaGu+N
MVwwi0aGua8MCI8cKiaxuz9vyGJ4lkdIWDiitbJ9GxWNElZ463KTqvkbjeO4tL3S
907TznOfif8ZEo7GMbGl4IKNYWLU27C+vX58kC8xYaGxMwnLSp5MwphLYLmCeB9t
VzNyf8OoQuBCcGuiq9RX+0k5XIBt+il9efJRO9xLonYyAbftEItlXB34YinhV8Jw
RUNIH1mOBwIdIE7aA1oHa/zL6U0g/CO6xA+Z1ROFWN1DvTCn81FPwttgDHFpVkTT
JmfFCASBmemj8JyOfDqsXANBCMXsyTmHItGeRAePHZUSXOL7+3BpgknS3fhlvryY
ZrjoRu69TX3fRrkSfYyM1cVcdU4obl1SDQ+o2noLbeQkMJjZWACOoAc2Uu3r5nVM
v6JhqOBkhkAOtGV89+TN6xCh0XT43c7bR2yqxm/hoH3IjVUAy6348RgMbUwSIv6R
7apkwllB6fP9lpkwZlAiZu8Y8FnP3F3nC1D6m9i2/gqeHE7h9LIxXQMwZO5w0aPI
rIvunCzbiqJNHMW65fHU+T0BjBXYq6IlPw49KZH70swrrcILyHPfeQzXPBuzJ33y
jVsD9Ess4gBIiYw5nSD/pI8IkvCKP3yLm7mEYyQeF26v4RjFUT25mXxQLkSDbjE3
cSn+5MI5CbGaOKGtB1iSRSiu8YrAb3UDjE8i2QmjOJbnYlgh1iUjWP0kEUku4oTS
383Q7eFe2XXpi+EgD5ymLdDsyPDE5JZT81tor9GuzOuStmXnsDtYw7Py88tMYRkQ
gmo7GITmwLu39IuU+tGwnMVoVmWB1gx7s5fqHrN5SL8wakVvp6RDIl8Cu4HBAsi0
pIKhFSC7B+RDAAwKBbXOLj+aH1iJE+dxlqkAvhbHS1VZpTH9gLgelndr228z+A3p
s1jHJUJyYS9bRhmiK+HIeTfwyZc/8otVkeQSGNwaynt3xL12JOTMlonewlwaVAKD
SzdhZk1uIzUlKFmiFqJ4y0+be41FmTZvwClqD+pDCPQJvvSo1OGkLX9SjZo4iMBY
2PiamatXrFI5iz3DMifkUuLeMmvmdqqxBCZEcxYpSghU5CxZoJRT/I8G1kn8YAxg
gi3pbeMmJc6i7nI5n7u6S0LCG6faHcNnamLeyfBWvXlg18XLZIO6CqB6KKciJjkO
piED1wfOK2OVX9o/PgHr5lGqLsl938wu0JTXe/houo+WAaEnOM6Tayj4nw+II0so
271Mzo5mhrzhXZfMZZpkSnCSC0Xph7oGI9YvGH4rgg2mU5JYKDGE+IGx00/MePzc
w/x7CmQf4A2wgL3XOfFLm9NTJMTHAqP9HWyBNde4hccj1KmCkqrpLYrPKe20Q+GG
2tEEkqsrE6ugYfGk9pkg6AlckFFQne9AoZfYUU0xqu+aTWSHZYed/pHoUBANfm2+
0e+jddX87nL7ULLlU0zYF97OWQXk7d09ZPSs9DhKJm3rubLrHdIMtIvCQgwESwaO
xJT/6dV/rGCoYWHzlrUwWq3OGnyo01tiCni03adhZAHd8Kcz6E1o2oBz+C/oFp60
lLLHRFllvB5fOlZXgDGcBGgt7Rw0jLKsYeIx2sU1T1styQ28KcqkP2J/IXLcsUhj
1B6e/kFR3A/aihvcpXYSiYUZbCttA3ooo09kMfje5Gg9mlbAMMPlyR42K5iKuvJG
IFAHZUZRvpkYbu6QndBtketyNJ0HScr2zin+7JvxeaBa/EgG9aJzByDVSRw+TcZn
LSQQfFYrMJjKLbd8AjU/nMW4LT+nh+QvtBQelODolTqsOfMcC4CWCX0zFUIwEeZ4
0ETjiRO21CxSLazPBfJ/BP9GyG5GoPpzrj8/hZMCx75H3owgGwnYwmdQ57/+wb5W
4tsjlJnrNRk++IBWoTGuHN9FjFLrY881KhhbPmFYBbaMzRaYPnnXIsMsoHYBfK79
H9MlSHBbM9hAi34EmINolMTpqZ13ZALnzdi5PzlERTO1ksDQ1y86abAThkF5Sk4X
CJtxAKX9qQEtjunwlBa6wSvCq0pxwNYCYdsizocmqbwkStOxY00LwnxmtYZ4V4QZ
I9Kl3wQNfyZTyEBlBtH2IR+55kl96F9XX7EB6tdDTbJRwOiNjTSo44yUtqwfbEor
4c5ywrtjh8dPktmg3pqiNkmecPvO/tysvqJ6X4Me/qmng2K06ONv3frZhwtJRTWV
z5cGe9C/basL7VD9CbQEbJK9zLQTI7Jq6OTBm9y4piyHlClMRStZ+bepfzElaIYU
Io+XVtRmTM/3+FOiTKBj4l+x7uILdMKpUImaUSzm4+tug6shobX4NUtVLOhDobpl
Fb/RS+WFixzGDwn5aJz49cLpgrMhDDmvNLBoZPOp7/lJham2u4lISM3CqAYSSptn
/ZCn7A46FvMBK3YHUGhlYy41mgTzezfXDSE41XsH9/s1psO6HqrGpxoxQh5sk6tc
1wq1cqRcj20w1frKRLDtiWkxt6TDdUaKtmAnrZWpaqkmsflOU2Vko/GVzoWNCo4F
I86z+WCVYDnRxwxtsqLRVi4xklqPmTOPZE7XvrpWNYZhz+0nH8Qd+BiZkQt13eq7
OOXn5CChr1StrV12pjN3fqZILxaK/iWLGrO50SP8a283qBBencisH7I0mFiJzoqi
4BSXjcMbpuoPM3KpN/Gyh5f9+ZN3L4aY43uwvFKL+3ri7rRr2+21cEFmhQEoNcF1
B6LyT7rtD0hXCpX4u13rVsaWCE3MKibGceBRMHggku8r489m7bdNHY97dmkvRB5g
11mCN5qBa9Qx8Q7rRnZhL/59WJPrdIj9JYjah7Eavbl+PRaZMsPmmPSZrdGSZ3Bp
Djd5Wb1tqGYU8gB37d+4OlpNHC7T4rCyh9OKAhYD78PyUtERq0Wo0mLpJ6y/mAS3
ODmA/Roe8mHtg8LBQLNTaziyaBN2F1RA+AE+Xc2811sfte/Wxh7mSVx1w2mGfB/D
3q6j9lYaygjnqrmAd3NHcmpiufKikcuiR9VAthIsyOmBpTSApAD7cduXyoorT1qZ
R++mhyCBVENL8EVqWv5tlVVPOPyYD/BTlAmTNiNunOxtiDF5VJJR4hCVaLcDASPg
1WZHNLjkrSPQODwBmd4//4Hqj5YhGeE5GzGAmJx2IuzUoFMPQ0ApvB9yZs+9LXmZ
mzoHNe/3Q7D6JZjRv7ca8fk2yxUYvCo1nR8/VxM/EaUbyim9pQLaeIXyXNAtJ0rq
6LuLLHy9ByRafEegoiT/yIxjAqymMx2XeHhTCkByCS3rHdm0AfiWPe5f+WYshrKc
xPg5Xg3RfDy4BCE+umxgqpfmkadrl0jd84DNfoyp14M=
`protect END_PROTECTED
