`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tNb3LQhanTbF5TvsUDaHyfs0HtXw8ZRXUOFOtcFj7r+miR9nxJaYtyCkncn+9qXD
zE2WISD8/BJLFhM1+ktV7oM2+qRnb/xStFwFX7GPwIn+VHYD5BD1oMFMiEAhVerv
uPwlE4K9k23pKssTSNen58XY5tKj8BliWJ7vL2kfo3JBbtiT+GUVj6Fp1a8oGyRS
R6AzKS67Ipfih9ig/Y12DO5EJGtABZNdcSzySJlhqRLqkWwEdO7CTPL0ZCBYGzqR
qHEpTCvI50hP/SyZw7PzeMaVYFujKPLUFVvIlM/5oXvPrlO6XbVbD08+uRH5L0Am
T5iHkzLuPgdDyuE62Y4fiOXpaGDqItd4E7e5cDVCeIKTU3zxTyf1Vfof/ERbBAV+
WIlUnQUqGKLOT8cSQwKDzwauzhnScBazpcAkRnwBldTfzlj3ZIZEF9II58DsW1+/
6S5OFv6SKXHMneET7Hlv4kK8I9Hm+9LJg8QHzhhpsrNx+/cLEAwqk5+m2GAg30Ru
4AYoHCb9BZm3LyAKSx9lPcMUaisbN+kr+h7BA6+hmOjlrfarEsOS47COGZN/lH/z
BemjX2mGRPUqqVkmlNZ4ykQVZ/Dnh4xrDZmwsaNoApvNswWEUuAiJkEQbDdhy0lM
WZ6wk9y4Vjfi7mUNwnObYrFxrdMD7KS/sGSW4McV3bDycxci69bxfUpfuqFzk+QU
FGczs9ARbuVLVkhWwCY1v4rXT+1TNyHwjECBN+N/ABAEo5EQi4yfFjYh/39qHZD9
Du1hevhips7f9TIJ3s1yQiHJsGjVcawqyiq3MCAZDTBZ2VhvUWmndorC7NiybCx2
i/dEGzxStKEkFbDA+okmTOcZKFz1CGaEK8ijntGQYkg+u+GNSnkalk4D3B7E6tbC
whQeGxDwcfr2PAfJZex//RkSVRLNA2hIszxCKwb7bzKJPtC/FF+PDLC7WPl8ld8/
gFz1rxaXhYAh3rlf3SW+hWFTbjW6al15OyZ3vS1fHUYBag9Y/LPHNlBc9YMPz5uu
YwM3CXFqtsG1FkfWNFTiyuy0SmF4gU4VlKZ2FiCoshSTN50qYQ6p+Cr8rJp4VUII
+9raKIMPwwB5v+R0gpD5uluaXXMJNrRXqfUNtkY/2gFEGb9c8sVrQ+uSLfwgWLJy
Ktcdk+y+ppCCNqBHc5PF3B9UWMpHcN1sa2Ug2r6ofo/6o9FnbCprA1WbtR0Avi+A
mbykCso6o6Ca2F4pMwpyDjXJlZVp0lbEgxo7BV8VjiGVGOZXzFvR/VRerMlmZu0h
sF8LRe5eJvnM8z3ZbCkN/b0LgrH6t6wcMSSCOitoQC7mFyr+jRpgYYXmtbkdF08v
5w9TSEetsUy5Ukz/7jH0RrHS9QltjOVvWVI/6+m/OAxp3GKznk9TtzKOYTi8WlS6
juYVlL6wTicbN2e1l3/zhcZCA8FOXmoI9j2lfNYpLApSq+MAIpwzQwzicNUZ4gYQ
`protect END_PROTECTED
