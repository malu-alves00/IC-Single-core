`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CmAKhQyawL6J0WRFC7pjXtN22/0r2s//HJw+pSIfMX06JP9EItKfEm/K89h2g522
2vp1EVNYapLhp2kABCOyxM1URdTngQkpDlFGoLZeJiyYQRzYrjfy6QBA7ofC8ZHZ
lM0hhMPsa26HFwFx6K332lBduVxR6LIbEfR6tE19VCsZn96PDl4Ptxct9YnnDj4n
uO3ghkPL1QS32ut7WyJGL0P8ZXmp9nEUJvhrNy0UubOezymKUnc9eICUrLwWXsCB
YnJ6jtSZpRgwZc5q4YuTpIjjHCYYW3Y5AbkYkdl7+WvaMtZCtrLL89H0BHl3UxpP
UW8dEW93zUa1CAw0gceSx2Iqgm3EStStCU6ehu313ps82Gjp5lzyNf1lEhAfZpHe
V07kb+sEBO0/+zEdV7Q76XEdPhj2ptoVYX043AgDF0IUUJDdcOWcPNsSp7/XLUyX
DLSsymZCun4E+a7s9DCys3ZzVaZKaJZTHRAc+GFEAhLPGzboMzcJ+vfN82Gn4VCy
fRiT4yxory925YPnZJqXcp0gHnLm7vspRZ3DATE7XB65hz6CaDt0ej4vMlZTC/vN
mOYEN0M4bXrhP/yNddbyqg+4Ze/hHBMBj2niwHXq48u5DPwZsQjZVQMabpE0zKoI
aTnJSXfPV7zUa34cs7wIXH1/l/ENkx+BVTmhuWnO2V4LIkhmN7IehnQSLXz/oRxt
W9mnfX8BdCJ+4SrXVe4rk0l/19xnYUNaRZcrkbUjac1GePlKKX52I5qw2xjWd5ZU
8iMPgOjzFSfSYMvOCb7rnMiu9x8apGzd4o3e8pXRQ6ZUJ/iZ8zzqNqsy0XZcQ1GO
`protect END_PROTECTED
