`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4qcpP3QyxrF/Ps9KDc+aZayD/lDmhcsrO242C0DAHLXMMvh+bUcX7HDUHQjO0kXe
YySGui0mtMqymg4wq/8XZXhnawoEwx+6GPiq6inezWdFGhpzF84DkpGsGpJhql/p
7RjSBfpt6lhofcMer9cYLuiQvd5rQtli5h7co9VpMLA1kSBCNqBuMuYWxysh+HOz
N4+92mQhpOweBvqLOrHr/DZzoBd7J1LNFm08QeOinCZZDea8XP4cQDs6gnRvr/85
wFjY9zCZIRpwX3HhUKtQcvG6aIqw6RbYC+pEZa0KH7FxSX681CvDqu/IQwSwM+X5
ao+fIzsVk8JR78O7FtRsd7cLm0/NDEB0O7nQzthbOKGopDXFyCj5WniRYAd+GapI
jM0+AipVB07ulknWfCA0xu/HEDAMqK6xkiIL1qEQot8+LQX0PTaaepX7wyJayAq3
73JnauV0Z7eWpWslkPHU4bul0FqxhXZGal5x7lwI6BFr97ut0f0dqg3y0yp4YYf6
kj0gYvqXPJzhfrhwJON1JekFeg2S4wCH6/S02dCtCTChsfvvQ7XwfwjFPmEQ4oTA
l78fx8Vt2XLnUH3uWsD2truC2jrIOVw9xqEb2ZCXHwy5Z7caR4xb03VGTj4QYIHF
BhFPRXxUMEQim+NtbMU53rd73Xul+CZW4cBXr02HxsMN41qCor0+c4XxtUCTFsec
OVBlhzzyXexow4TvmUDOPhI6eUuamuDYLNEFT3vhtL3VegI3Hwm6fPNnd5aKslif
Tos8cGKFDcqN4/kHL5ZS7y6/5SRP93V3zO+hGBzj1VBXVKMN9rB2MKAzWAOzGiIV
Jt4ZsfsLj1fl9uNQCYvumAXPO5eU+JphP6d/c5qQRi720At3Fep0Vc2zO1h6SduM
Uy0qkYpdvGWjrHLEWE/8kQDAPn859m/VK77Cwh3Tqt5V/E4IcYp0EHPn3bBXc1M2
QQ6JCpWzInrEYRE2r0Hr6tAK5mLpyKODTyGQENlzrbf8CpxT8krqTHfduF9QanDb
5Vn9+p6D/RyxcwvoIiW2IVI7eG9oO6g76Ah5vDYHXOby6FUHPjEIkyT2jy82d3nO
ARHTg2NcChU1XBMBSTIY6pyJnHSAb0riF6CLjPIuqNBGLIojEWtJLVHGnnsKxqb8
ekiFrgcamwA2H9LVANkppp4egcvaFDP9Ho9klLoSqJq6iifJFo9T6G6bbwX9coSE
Tap/WcyL7zITpcuNJ74SZldFfJJ5Vs5a3FE+I1yTS7TpEJs3XvhvpgOVn9sZJrTm
U46HWg3/M+J0W7mZKFtqriLPS/4Z2r8aWJqZaWuwNQRH/qciOyPMsKyIKeyUpkSn
KaBw3o+Oz8Oo95Yax7BG9BXiFn0CpwP2ih6Svt4Khy+DNRFJy5/Q7+ZWLC4oV60U
F+TGJb3Ak7wKlrocqB74GGXfw22Jz0EnsaOFd9lJJudKcKmi2ph8BptWrtkiD+TQ
i+GfddG+Vs71vde1RRC7cGlLFfp1t8XV28601zmjASULp7XgDt2Ewevt/oOluNVm
0bspLRZ5qmeWT5UTSmP6yTNltnwYeL4J4h7z327Xm0//xadoheJ2+ajfgmvPGL93
17taR+C+aOLAg0bv2831tf9BMSpmhEI70+2as78EV481dK/CvqNQwgTveC5dWgic
5A7AXW44PYlhQf65z7lmD8f6kxrKkrSRVjkBcsPiseeEmTvWOHVAiY/cPJIQtpZR
ajZcVAol5aN4Rhf0nEd4tMQShlyf5WMfAQAW7Mf7xNRtvd/fBzKyBFyWhajXBhtP
9J4Yifh0wKwuOh8XDT3TlxTCQ0hqpCC7Vv9ZLlqX/psEwlUDbA5/Eyq8SbsxD1Y1
pRmAhdDuaUOytWJfYGl44SlqCV+ElIBiLcMCs7mz+gkXeW5e0M+vkkubX+U3i5s0
/B3/MEpzHPYiaLSOyIff4Byod+1hi25c6RhQZ/S64LpRl2vqzM4sgup8mpJr+1FO
8KYe93FF0NNecQIiJdnYmEFVRDSDPCVkRpYn8G38CN1v7cF8m2LnAwDbUpFxXfZk
Dh38EPZ7N4BK3tkkgzIkFr7nSZBum4sP9zdPPXAxgVTfzcXT8jz6+D/2JRrTojmz
ENTvcXEcoam4TFWJR4QzGiY4cYe1NDFe1HI3pciakI7Lc2DPSIgovFgUAsrNblas
GmFzJChwrRsU+cxuVnORnYv7XE4bHfDfAq+Mkjs+LbD7SfsGh5jS7aDwEC9lGtrp
AMlcJD5V0xhNeqZWdkpDlBzm1crKH/30Si/Ic41H0hiR37arEJIquf8SZT6G6DTd
HRak/Qzm3s4ly/fP77lXkcawY6gG8DHAk8XBhxz5UrREzUvcdlf6WYHWnNq8g3K4
+LL8+VvCLxJWNXsTWTNOub6+EYWF+q3VbLdau/C1TgM66rFxt+PXrI1xTAewfwWV
9vGxMj9ZMVx83o+Qe88c2uE5LlyXB5Ei7x2wheSful1UrofGomKO/qdu3Lcaiwlv
fbJN0J4LC738wXG6wd7wVpTdpQGbMVAzsBfsP3CQHS4DutaeZUJOkDACjyPF7H3C
ftNw34YKfW9gM8Mj9R3V028G3J4xuCU1GkbusjRgA9Y9EZaLJp8j9f3mDMT9gJkw
Qegy70NjpW1kBcnXen0zfgClq0PXtUcfVhu5i6sBL52Grc/LG3Z8V0gtV65mslKy
WUyT4h03Td5A7TgpmVvJmX9Xq8UufmhimRN5cIBPSatBdXtcZTC/oCZJgla++620
0iYNirCWjtAdhV/2Ng9Cpz8p/SLMgq8a8R3EpBGO2kdX5ofvGIhYgJWZ4L7NMLSl
oNvm2bd/aBB7RprZk1q493KPyMZ7buz/WXAwQ72bVYn4fNsOcEkX/223u8Qq7euE
4VCsq3VX5naM2qpuWNvn4KJe7uL0Pe+vJA5lbmKmu+607Bh2QgWhk5Mrp/wybn8w
N+6mnyG3bY8kNqZc7gs7zCbPppBypLexoyQqYgAdJzJJ0hzrEr3mXD8Nq1vddRg6
e9wHnkqc29IT51+nvewf07ElcrKNjwA9mC4GHo0C5xgdWNP3BA99Lb5SBE0lSdYh
gmsZnsC0lCTRUZS9T9YGbS5b7LCjVAQy2xPDI+GkV2L0zNWXYyjxMn2rwvb2i0Fk
9xs0eGdXsA7Nnvfq9MaveLSc4QaELe0vfD1T8+gv7mylm7OHh+2P8FreR9NAXK4B
WK3XsqV1QWp6D1fZ9ZtyZ0gGrawxoabQLybPs/GBstZ33IO2iapHSrrmCeu26GMi
YKeJWghHuje6iHqIRKJAWBFsWc/LptIelrNkTXTWay4YzhenBuwrN1SYk3vEd9AJ
Y1Sjtwbxxs9F40+ZhhPqltT8G6jmlh8quxlLSnkdRQ58mzg/RXNwIyK8EEpjtjRd
/GxxTzxBLcH140Xk3h9EquXDI+C2+DUGhIUrkDCn9+5QiSEMbqr0AOR/okxC1/nw
fBUwVIQwpfHwJ8gLsVG7XHT36/1f3Up7r5N1brDACi85iwM5xqsVFSxZ7avbbSg3
U+JUYMleByHJWCX+zxW9bCub2LpGNnEbyv4ldqg7KFAk3mjy7YMjVssQDAionbEN
OjmqVJ4kfGkweq77i+SWdiHjKWEGUx8EnqhDED02ql35OgD+4B62CtDFWKNImn7O
kHWACsbNlagzkRj9tZ9gYJyx38NAELx8i+/PujOMbL4bUvw4Vc+X+x2ZFXIfhNIx
LaUahUrnb5DZtxrg9lDWKHq8ia2F7r0ktMrHmN9lSmH9ftaQ9d0bBtSG23bjtoqT
pMmbJcF0HsHmMlEyrNAXXCPxrOVkwOUghQMAGr1lFKqF3OBqZySAD7c3qbTKmrdK
qpBEhimjB+tlY+A9xtgt2cS/mFrVPpXMFDlNxkTO6SXqYVe0w+CrcALkYWsgGh+3
xhpwWx2zwxVFVF1t0UbmKce5vS0m7+F/cReCIZhqyrRtiQn7a+fqsp4WvQhkPUKq
aUmAg9gkcPuBU0mEBVKPKfevK72qiF9Ob0vp5xfqa5Q8NCcLqLwWo5AXDQ2KKVqe
zDQSUu7THwMf/eiIlK9y07qti5Mly5ZZ71OFppeiRukOqRd/V8eLIuObEDOJY2I0
VxlHfZ0p+nbIbW/nIUPJTlfpkzd5HgrtDafPLnEGwwWx7NpbuQAXWHqqsWN7mDyv
gM+d2GxZW8JbbOYbN+A/Z8/itB9D2eeaqLnIsrPrbAUzxR1YXdo/PgF+pmiSmTvd
QaxhbUQ6nEUPiuQ0wTDotlouf2QG6ws9Au7LpFUmRHi8Hgj/uqkl1GwuHVR74esB
vxsCu2PBo6MIECFwS+MEevnvXYCjxMW5HaQofBB/3VNc5C7QO28j88/9awzh9AeT
Akfdn8nR7RQFYugrMwFlAXwODb16HFjVFPgrIVPIre65rnlwxzCwzZGVBQs4k+9H
wToAdJWZ37vvuvquQC6pqJF1FwLr7hrSevtfCGkl9WFIDYCsixoxfz6TdRHDw2hA
aC252Lz7az+i4uQwOsuIKbGHa75dkuP5NHnDA6RWRph6gBGX6bl2id5tX60OPtBj
ykqWo2h/7zlq2hr3/I3U1g==
`protect END_PROTECTED
