`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kU0IIqjHoIttOw3t9/UNT+A19KZtqWBQltOvjsRlgayfmJpqnR8lg3kLEeg0C4hk
gzCasqrHnComW8Htx6lEH/DkyUXbenqRlRYb1GUGE7ZbrBSx3nyVQ1+Yvf7sYZ0Z
iAmHHoQnn/Fd0GTfK7QUCnK689v2Q101euOYUR7izXD5B7XBKhxZ9+V+mE/285h3
cq6bhwm3sTBcIq+jWttEEdXEwhVZSMjav2cInI9sPUILiNe8rKykz4wXzQ5Z8/9J
wVWBydX4O7hzIUd3RqrqfUgYELoIDNSiPlRR8rFebdKhzpNUb3HjGYLGMxSHM3hD
spFS4EpDkokibAbl7SmwIZgZllDaYBABEmjHmtx51/W4AQ3PZ42Y3QRCDlUMQyaD
wFQdoI2k6PRJ33luf694wQPvi8fIxvUDKAqfiGYw1Zt+puitRXPtrkq8d6BO061Q
uZD/eg+Rezufq1h+jQ6eZIvg/w+/g9df946sGAPgnSw5q4281pUJxIX6/gigSfl7
berKr+4ZuzlErSRuIc8CDpyR9Tn776ZXOtBWoLlnDz4qTkAQ0wfi3Js6IJVeqns2
HMOlgAzNzLfWREhc9ys3hmNcu5tCmkOasag6JQYbuBeY7aOqjogURt/irWLDf/pm
F3Js/qFOT7IhpFZg3UhyPlXLgtVop7Kp2aKC8hpNWY8kEozJVRJPbIAWaOPcKirp
Y70PZyG4xuKtkDan70J/BT4wTS7C5gDVF2Cwjnf3aB2Rw+v5ESYa1sVvMt9xIF6h
Y/OWzy/GbNlb1K2ibedHRBXzjBch1lbufNUjgFWH1/GClxbwtTeGL78HlSgf0AjU
UCrtHaeWrBys7OKRKwhpqLysZuAXGTpHZ2EFTkQucZM4Z0jdhu8RropkfNbEnLzi
8NgNB+Ah4spK4CKnhF8xktN8+WCnKWDwGT6MwlSdOyML7ys2D7/9/osn5Top5H8Z
2gUKf0Iug1kE9hgpZS7FVXB/vd8JtmXKrC/7enJ2tlS9Bzw9U29+mn5de9mfuvY1
VKKI08M/fdft7LfpQaxLXaZNG2F+88tXR/BsPfJUk4Dd2tIJtUJntm8Zn/lyjgqL
IMk2iMmxS2Qee0wMFL+ERgUdtNSlw6aK7eiuJCfXYwB4NGU9JFLHesd+nfrNbXZB
gZcFtpMLmKpLId5Kd2O30GrjEGtZKEShh8BMPeSsqDO2ChqjQRAjm5fhPPUBuX+k
cOcsK0mICbXEQzT0Sb3X3c9bGJBUg9f0PSbVXgD4l6R2q9VlogULIRnpoHVBTjCh
4Dg9T3wdv51AY5zu6h0ejQpaSYfAw9RVwFQklfdHcg6iYYmoiB5J2mV1nJBR34hv
ew2DTzdbflaKX/Feo8dX+Qr/8AMaOwsliO08Wl9GKXdqzFXsS6s5EtMyps2/kK1a
7nsT63krYAe+ayipGLmS8V+zbRiod3CqoUq+kz42zDeM4g4KemkbQGLeRRSRLbYi
qDsc0Wt/DihTbtVNn8mQWjB+R4kegV9fieWTaiXyBGtcfRQlcmDbhUxzztU9tPVH
3kyg3pZgbkcvAfYmCMKhixcfkJcQDmtvzst7kO7dcn/YABprziYQbMyKiKaQ1nkj
dETFEBKpAIfGH5SwOASEkAkGk87hG2Cj+PxlUtUupYd60F6YpB/+S5Q2lASEeO03
B++9Fr3m1q2LS1Qh0io/YRZmYLrHDS3hb0g0QLyo/zvAUafEQzQAU2n9G3BtptLZ
kRElKhhkEc05Tb/b10RED0KVmiWYBGyN2Y8kd9hvEuvhskvNW5dRp5wLCnHok8vX
l40tiLYkT1L0D1+hoKG5Qi8lwjsATQhIMAfmprqwRK7uUwEW0qsiFN8gbhKOmJxW
qSD+r0Kph3U1Ye3E8lGJKvA75liIL3MclBXSN3pR4QQyzRl6f50NtOCeAAQ1e6Aj
fBSehj73iS9BfNvlS+Jyogbg5O8x5zrTj1EFS6mYXto6rQLwdR5al2k9EX1I1fvP
iFHZP2OVwzcV3PFAMzTdbaBNqoe5icZRvGSo2RW4AG0wHwgMEbaDVcDO9tGZd+O6
8vGccgRZnQv7Q5stEGPDkSGgwa3zCgwkebA+qifzLwTRTj/XJynaOJgQJWb9Eobu
32f3lGIkeJ2LsZ0KJHffm+9fqxE2DiTA+wbs2znW3gZh17/ZZOYY05f3wSoD5WEj
aD/AB2YNiEYNJDkd/BwpgOJrkHyOmGi1OvXm2uHBUrkw0RDenQTg6Vpl4DFhcHCP
jqKbGWSNLtoTA0tg6Ze1mMupq0NgOZFEp3eda/9FoYnLRo/78wnoPDldDQTTJ6m1
d4ViFgkJvCwAkTyMuaG0/YbxiOnAm50nHMfNzULIWwoW6kaPpIyGTnAGCIyBmwK5
fpPdcJBIrEtKR6okTxGB7GUzgepE8eMgELjzU4qWIs0mGD8S9NPP0P3ZTOJUl7sF
qgy9GTEHJo1+5PKy9ln1E8E3p3W6DlEN7R539e4ArfoURAsVlU53U3HJujNgECvv
+JqVd4D2+TLXontvWyeHUv3QT/4eY1d6Q57MlSJnIPshiIUC0yyLLRNJJH4vexh3
5YEXSs1mEagohiY5ReFTBvg4MaKHBq+cj7V8WZHz8Q/bUgKeks0S/qCS1TsOkwyw
fozbylQq5LHx/qNf2gFd/XaUPveAIUWF8g+JXfO4w33gXEbpu6IGny/yv5v9dCCz
IDiPCRFJgbJH5LM4JjAvfO0ZZBs8jDlclIkYvisdpriCElxklGXn5qEngKvTfejK
7mds7uT68Zwoa2rAqN+k4rwi7douXsW2UHELX7l9cRCd8pMeIHnrcWk3Uz1GTcPY
kD2yZEc2jqymuShCKSBmFyWEJt47FyFi8vXL9g4EbUQ/Q+wLNEASx/VkOcEaK5M/
2GUKbyVibuUbpHzNHCj4zs8RHfKggmw2L2ccnO8T7xlMZgthrW1r9Ev4Itr1kePc
Mq938Rw3PYNgHL6mkczGwQzL75afJIQe433HaB2HikrbxcV47ztcqXErqBts5SCn
lV4haO+le9v9RGD2/oRzydDQ43VG6/aXOjEF4J/5SEwX4u9E59i25ehkTskoV7Lr
b+682dy795NuqckpfKVRsLg8vUkRDTrb2HPfASvwwU7Qdp5WWDjXU4vrb+iKRK60
wuzEZZ/W6b8JRb5N2DvMb2KXKpkKv1/68v3Utuo5cFYLgURhfjDxkUV3VNyPBRXt
sWOg1c6g+N7gRBYNFmxhF3RoAq6XSV76WO2O3W2XCGDHet7vKQi7xsk4ZvsDEbhx
nZ/mnvbDCW1ey7BDtPXRe+mpsR8aPT7GBjTeaEv+IhajA1Tcdxgejp2TZMamQcVX
Ujiwe/TdW7inEahPmvjAWQaIeoxmMNqD1R5cBpyMUFTlePGVpq+HiyPTfOlSHxVd
L/Abl4GqVtOsgrcgRcob1xTF4pk/Ww2vAVM+D6OONpNtdbriN4+wFRF59K4hFA5o
a/zyYWBZgpQw3pzhiR/kX+eSGzPtRe4QAgVfGhfIuQj3FD4tvzrgQEkSgRcS1zJX
S6XVMJz+xdGrJDtT71zEfAmYO2wKFxmtFh9/Twra5k6+0gdOEiZqVeEs4NUavNHo
GSXUbxIzVZPbtlzpbqKwTvBSr4XOF0CP9FpxDhcPrEd2OwyuzrJZuQok4rIi1EJK
Tf3kxkkXTjOp4CgYHrRT3LiNXDELr2v6I16H5IDf10crvdT5lqugJdqqcoi+MGOG
gqyetshEy6TQ3qzY4rRLOdB3HBmc+lhpcJiCsIUR86A4G7AhqCEt6Y+cND1KAFf5
g7fddYcMoccRW/7pSrrGcmqkkzjwQyjsqp98RKhzPlKwhXqtX7Mj2puBfSp2ejui
v032Da0Z3OK/+7x3ITlPjnIHmNU8QSrzeeqx01vrrob9xzJCeazZdY8VsCD5v2Cw
cx8UF9ne9C783RNL9wXMcJH+icAmEvACGNlzeozjLUDoWkb6QZXc6n1+OAXH/f85
hMThn+OFN3dsPodComAQOuZyb0ExxU698Qz7fDwmMuLXo27wtrZHATs9SONfDkR5
jJz2R/S778eUTWCOdvC8m5OHLbY47OK1Lf+dn0fQX/wCHrGD9J6ek7xb0uc1PXPy
YFGsoXJNgGfM+wSOtYLZuVRhPDRIF+W87gzRTfExVQqm6rciWcEuwMqlARTRv5Dz
DutKQgmrryyjuQpS7GAwWB/XnhtUCOo+in+o+krnvjyRek98lwW8pA/43HWujkPX
XT5s30F8RL+YFdVPgm8p/V79cJNuM986blv4Cfyzws+57jID58r5hPRRvqwIXau8
5YNl/rJyApKH23LxFdsSLEsgtR4Vqj20DcgfLOyZx+kv81YdD3gQWi4L6w64BmYf
OSqeqphrStQ4r82+rwR951f9V+xm+CnBBqCACY3Sel+vI/T1bWBxHGvQTppZw/gT
RXXSQnoJXL50g3XjKMvsOL5LEjfXV5Y8p1viWtrMFIT1p4LEUiP6h5cS1gyIpWvw
SzNtgjf13LMelEjVYKh/ou+MCROO9bVng1++FCC5HzXVePqw6javflI48hqDKD5r
BAt92BAOoGb+XhJfu5csPzpx+AeWcVesAczbLjUY6Av9jHi6Ggqa6fAyySKMiSH7
hu8iIrR/DQ0xVg781yKyvl9fNKkFsz4kcEJPOD0VPQrGzT5HdH4tAgLim50ufthz
txp8H29VOk8LKkxh0xlaw8LDQkUYPS4w1MzSgRXH8VMbj6c6q3LthaZJqdm2KIlf
Ak+2jlWfoAszI7LjB/HjIt4fz9fKb/c7zr7726gNQtk6ynRr+MPzpOQqPQcTH1F8
Dfc31jWPUZRf31huC11zAiOAvDXcDC3xE3JUuhj8dclfp0at1U0TQRktP+1R09Sg
wptxI1/1haS/D2FadZWtMcmsaVvIQCApCxAJQFthJHL7vsmpi58/7umelRVFHCXE
BINhMUZsUPVAKNF6WJi7kMpZlcPauceEE57H7dLYVhyOZQq73XUaf2bt2EJL6LQl
Crp8Eoq1ex9FiXIWWR1q7/3b+FYr1WFXGyE1UvNuOUee/lkWRKBqMXEkaJebtBTe
99Ue92w9PcLF1XT336LfCgtvpNf8n3zWtdtZbg91y6PO7Rktdih7ZbT9K8aMBUtu
/JqVwLm1qXQ9f6rTBc6XbqAjdb6s14x8Dz4omOgoHRyNE5B0Q4V9H337fTuENS7N
t6UUYlMgjuJqoj4W/0BDpv7BaklB+ytN0grbRoXe85BRETXTAvTjmAXfe4hDu1HV
7dqT+lHHjZ4zJXq2Op90VfOeEnU76DYXOzyY3m5u6rQPKU60ByLKKEZVwNCa89Jo
PjhpVu+P5iURVHenpRGrWN/Ej98aCtgwXuf6DXkmifrtDPIcI53VH5gbISHIsVCy
NpsgcPZqXAjSPqYfcmeaBmoOqEo/oW6RnAjsxNwDHF+i6DrCUcpL3aD2Ql3i7sKg
wGKbHI2PmkBn5tj83z/X0TAqtXfUmhX8s7Z28zB2y6nwqMlvOFztEabt3bAEc9yT
2oaKZX/CNt8j38sP4L3mA/14XuYeHmTFuxMYMRRpo3UvqT032Yb5uw/UYQvYTy0q
rYd8fA3swqJmZXMJm/j6mjQWz86m/41FC+M/NNZQgF1yRoKTJ4KpG4BUsEl2xcV1
j+JlZu/0oLnrZYNeYPWp0jTGoc1ME8pd2UR1mihCTOPrveYalq4KQnA8uDHd+cFv
Q8byBTYwBE1/fcnkDiqYB0JgdGr0tdBBye9eMXaNPUPX2OfceNC8KUZGsvNCDE8w
Ro7C1FHNS9htcPv7fKbblgfHFkaKVQ0z3YooSYXTJJElxLzsxd0LINO5cgZ6ggIZ
fuOU3TBxFdUuDOVrywhrxjQETkIHz6K26LJGLErzotoaATPoh+pFefrLBlauclOd
VoAx9rbqd4JnXjaYdbZPf1JP7O3PJIywH/+SMuzcRbYudxkCD1pRj/dzR9ELCiCa
4PsxpIncBtXF6D9mkmJcItYujTDl8uxOCfCQorjUnxKdEXdRVb6Hy/+9TsTKEEvt
KZwr8oAFc1nWAfvpOqE6F2PCv3IFko6WeCoTkfkKVi8=
`protect END_PROTECTED
