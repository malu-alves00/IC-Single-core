`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Eky6r6/Mgo7ZY9xnlSHIoRcPvufwzpuWeOVYUmbjTrVUSzBfGwP0AL7gTNHOcyuu
g9WQFvPpaSsLxDNEK57T7tP2gJf6xKtJ9uouckFOaSQWGKXLAXP4xhdJRqUvQHtP
BP3FsYYlOVzLamWhmPt+Nekf1RUZl4oLJY7DZJsSRCcoFvnPw6CtaRfd4Uhd/uGf
Rv9qiyddhmZDrjKqGJ62re4YL8D+Z+e1/D/LmkER/O/3/TXPXk6ixUZDMFJO7m1Q
yK/r59+vy+jYuduYnTPRpuj0FC7XeEG5YOaq4cSdCq7VQrxAtG2CFwzI8WPATZhp
w7LqNLRtc/QZiYFkQcENQgA5+BgzrDFVZVkoRUVjvy7s7pRYnYfXN3wLa83RiVAS
VsuAa3YRRnxNvIsqh4y8O7MUY1njoLHHWE8tTWY7wT4V/2vtIxT6h0qbhKS1JMBi
rveo7n85b0zY3WuqH/4eCatGSx1SoxH/5rg37wVt49S1CEUMSZ+4/iytMxP2EULQ
`protect END_PROTECTED
