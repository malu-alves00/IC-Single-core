`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
J8jEdEanonY8ye02Pd1d+trsVYZm1qo2rUpWLwyoG2opyR4gEnoNUwTnY3UKR3WA
inLWazbpefRs85/lg6c0ozk/jtj5OpgsYfUfMJcIxhPlYun1QENs86JMEx7g7irx
8Eu6NmNa0/5oE7O+dmh3LHGCviUS1VgHjQQhrrKTCYakN23l+e32EbDKk/Lwuq/n
vjpDvoFyJvwVcSfV1GO0VF2d/Rzc641hYrNIDP7nn93sFoNyPWrK46jziW7XOEIJ
/+pezDJEYbSe4HCXdUsHNIF7qU0Df2tY/oLT9Nl56+eRH2dMj1CBtZQECRO8HT7N
I3P+oi0U6b9bx1I+GYnJioRPDvl2yHMnj+9t9uDS4zmdEs24BSgqhEsXwdFg0VRo
oso9NgJknKWKSx6E4XtllaDGYb09mTj6lle8cSGupmJ8H0bArar+liZ3fvtftG74
TnzaS6cDxcnmCF0GFZHnBsUVCMfkIxnqrf9dIFtoOWzDc3NjjyjFy506bwN6sFCl
D8ukxr7vDDi0dKTCcpv/XXXgmP8SXULEALOMe0z5pXBdrATnBBm9bE+4/kC20XqF
TYlzRP1mjOl/ONZsnUhEhk/j/ii7qAgfmJPRvJ9314swz0FmdAAid+8GDchTvCDX
M3uADB0i+lgASTtyR1QJCOKBCFtNOjIbOY1sD5x9TFn50fELyNGXhkwrOvVIWH7t
5N9ky4f94OqyFdMg2Gv3ZJb1ClCGfHfsx6cQbKfxIrQASTiaHoMi76sp+0v5RAge
VLWDJfXBniGqt2vMDxosOXm63jsR/Y1K55ufZ+uRFgQcGWMLomDABZhXbN9kNtLV
k9yutLejQfa7dl+RXCgASWGRaCKvwYl5H5Ea5RvQF8qnw8XiplSb8EA3yfjKBbCV
BixQ+Yz0x/8FSoqWnalpcjm9XyABdZOCOXPD+ULXxSKKs8zsct2erCRfslx0QM7N
ipAYV4dqZOh3kOCSq0MCDjhzPlyJQ/5+SMHRYVBGzVIYO0NxH5liG5UiBjkD0XyC
smNXVVgfHVWnB1VXvpE77OWLb1iA6tzWMYvgtMuFhu7C+2CL783wqWz6Q0S/fR1l
4Vw07tymzXhoz8cJPX8+RCdqBMITV80Wi7RAgo4UvFXbES4P2Lav/egQCQ7jQo2G
E6q2YMJUv/J0349PulSO5Fkh8BdfWFtz3IpHxsWjrh/X7lPd87zMfOrNDIN7fcG/
rLGAt2vYm5O7IKwKOVOX/ITzkEB3egzb2kF1p/Z8Wk1ZQ9YFCoBvJitdd1F32jbs
MAw7yFrQjcdvibaGr5PZDSzWUj0LvV6WUPLrUQFaCYK+KF03/zfZ7Yd24yaE3Hw1
UUrwjbOl9S/buqadRQq9jJ3vTjoli4yPk9XsaPIpgKjwZuInSsGRWBkD7uDvc6Ow
9VfbQOstvugpOhyo7NjBRNUETOLoQiTj8zqQHvMeTJwCUeIuOzIrhKFkGxW6+6+9
OW8Hqg+EdZSEuPupFoyDnR7ifB1uD9Gut6Foq0V8Za9gW1vB8OXNYLoFtXB0ND8Q
kgAkAWLp850Nm2J4cRWkNFmsTdgJxXt6ixU+UtMdAxyMN0DLlzHHawogxr3XqH81
xMrNBWZsMIdcROp8qnAz4sB6X+3eRfFFa1GAPzfvp7bHTlQOXWyV32zpvB+u3GwV
RCYzXV32ZzMqsNdpj7iYOYwTiotgbag3ThIoI0J9j5KH6g7tdn056osd7tF4BRk7
Kr6FI/pIfpFDPmdrTA4NA2EM34iuXGZi3rUZRrcMUucDrcqAJ3HlKOv28/X03CxY
8cJDUzZeo0TN51euQR5Evelp49UF73MsdLUWlL/e4hv0yezouhtJ0ApoDsfdAzW9
EshtwAATGKRHCdUQsjWAWKQzS1k5nbfKWw9cp6TivOLgo9SldOvBhv7ABmEmekQt
gFDyoQiBX9aORWsmRBnwWaGK4pSL4yHkpfOsWlVc7jS0K72BlT81DPsZ5uzNgIFh
OzksZxR0/CQf6f6JUzpaSeGT+OIT+q8GN5Y4eZVWIleDYU2LGhYD3m+PasGAdpFY
EQys+E+QXVYR5d5yW2cS+VtyjagD1wadbPlvIU6+DFXoVep9ks2t4Erf7/lGXlV0
ST3MrbCyKAzMRhX+NkSteE5MtddaQlpC8vKTwZLus2bYg9LRXfN99fFivtCsi0Vl
QqjS5rDLGB+aaP3S70rPnuytxOuwZHtNyzhhOa9t5FSIQ9yMq7d+PMMtbM+WI/e8
VIek03O2LTurgc4GbLDlRzFZjPu1HUgFe9h6Hl2Hl06/awziLmU0C5vmV3K71f8a
BkuJ5igFhF160xJN/zjuaNv5JWiCnTsMnNIAd5L74vpNxAl3NE0uDC3Cxz0Jgbjv
Eeq5MXnWOFNQO+D58L1/qwIEF0YUoPYnl5+yJzD0Z5GpFZuKwlXDJN/Ni+36wnNn
SmkTBETdG9iwzSZ9Xdb3HqHtZl+Yxu2D/Wdi7XfTCwTBDKnXr1iAkxP/UHGLwHs8
jtnhqf0Wt41hZEXcFLrCoGp2vZfjVu1PDjujjB3CDRa6lHLN3C3OU6M5Wx2HdT/k
op3pSMphr6lEC52g2Jh10SatPME0fjxPr3He6gu4/RNe8eKZjp9laOV425eTNzfB
gqWbFtlwQ2FT+GRvb0/xYOJzwGGf3ldkkQYgzPoubnlGntJFZG3eihEDIGuMern4
JW9QByzdMIINW7dSeLdII/wirS+8JY28p+aYDETqH54VqRnytpf/+07hM9f5fDzj
JoY4nmqHd/uLGKwpUiT5SqaKv++sEEvHZadSwGqbl/XYn7pBqwpL4P/PHvLZ//2R
7mA4XEoKag4FQ/xha8SK7kgQG1ZDy81bdDMLN+RC3HcAlYcJDZr9jd0ZjdpaVif+
nGlmipY9v8PbbRuiSmP/WhN0q7rHHuqjuWYQlPJXSjwiove5VwKRh3PPch1ICjyY
Sh0Y8n/aWIlCP9gust6z1Vr5Wx+w3ezOsD1lRaJSzPmp6U8gGSNw/Gsx/g/XuchE
uKUuAFns/V2QOhnDmakV87CowO0jo+M3D4SzacQ+mbtqcax5RUm28Ohe5tS2yr3m
RjjlpEskJJ4Bmr/4BQ5vtplgFXJAxc+NFHT26BLuObOQ1CqCQzt3TiYP+RJqCVnX
daCtdw+VCxVxMqboTIfDUZNMcMZdWB+PK9dUSiRIyjSUSD0dPnsrBVkKT6Ucix4i
j7PD5JrCUnXncq9Hu1ArCjDstPqoOCp0q6mlxMBjpQE1nXoJYs93dj9+YuO208hF
yEft7wlAKlbfSZXiBoI9jx4TQ3rdK2qbOMvfJXjEuA+6a4c/meOyOjZyiDA9aNmi
aZqAeN3L7a67wGqHCWREfN+5LOVvE4iS9O6aRn8fHcXDtcnSbbIY8MJe7MuDZ+00
n5ieSPShbdMsfrZq4qHps4Av3FBt/ckGYPywA5Ig5ZclkVaDO3jnLElOva0h2FDq
qpwa5bl7cUrFgruB1HBNxXbRoSxQ0FHLV5Bg+PuuknYTUwL4L+ois/HTIBN1AKqf
hVzhMviCm2e0Ckc8KR7ZcxL3QkTY97pn7/3TzCUi1TvqlY2ROMziDMmW3KHdjvpJ
8dyeeBFqcyfoCQ/nsWMugTSAmbFzHthLFIjKWpbY1YG4JPGz1XuOLtYB+VXuSjRQ
JMU1TyrttqhlHtnlHVVWAvdxpYlhrNgy7xy1F0Wz11YDGB7FKcBK+wGEeYe/d9db
k/5XTVNqheRQhigan4TdxryfBNTJnuHXfddn9qFFCxvkLC4QSWZhevSAXT1VvNhp
1C7Xs1lFWdFTShWv7tj5JFystKdkbqM1+u/X0o9cYvutlIczDyBeUIdrQx4LM/zN
JuVi/Pt9AKQ9zvR1M+U9BmwHuJ8XDUtva3IUxAeIwSUwoq7MciMXufP89R9ncyCe
zO8HpVcwl3DtTCFM3DK4NTwjSdKsvL/NftnYX8yXo+35+Pp/1qdj7Q6ykcOVzp8a
StAGAHPtPE/o4Iz4nwgVjF3bFu1QxyXZ/DCz3/gi3EL4+A2d8JfxJ3EOWM58CAMg
hn9snCYI1/lG9x0CHiOg3gBF9Tbt6AcuLezVIPltOUXNDGb2SjNN9fI/0rCm9qMy
WwdOETDjPSkbto9aPHaBD1GirruFXkZmexZwdQXucPC92Vr3PosR+B44vG2w99qJ
X1Q3Lk6xnPZCfXaZVA1IGbt+GMyMmNzYEKAOIjqRjUCb8dDIA3s1QgcryiAe81p5
RojBgjOv7uBXwYtSryV0JZSITufZo+bMdPx2+4Md8q9rRMW5XvM115qZZZSYoh4u
UVY/QvP0s/7X8vqnoViaBQTC5JtzekJ1UGwPTltQZSdBWlgHSVSLk/vIaC1anNOv
Zp0ci6Aek0KXUu1wgsE3fvImzmVjwJnREih3OJNv0ZE4UICoUkgq1/QSp4Ez8pWh
Isz7i/RliPsUDyJMZ8UiwKImfpJUEpJ8j2NANKWIVOwqThcRWRGYLYtxZ5O34Zw3
WQ9Y4ie61zm/Ow/0LShrG+ZDOfYHnKpIaXvYaByj5N3YgI2GOTiHyr1ivS2GKLsV
fcYU/wUkYCv2cKUVri/b0s0erxSfC5dALSXcEIQLJJNo44lonTKbXDkPCi2LTo3o
6jPm8hsTKrxH0/Sl92p8tqm28nQ3gBpGmfJEJpTHrM+P16uY8ukAlqM3TsgqEbGs
hjMLOTS/mG8bFgPLtTE6b0f2DThZvleBK6wNxjC8PLf8IYZeZG7egpfTWewLkowx
F17wBoZ9PwJNxfhWtSkNOj/YgPuUw1PL9V8M4Ax8JpZ8oAyf8itXe4ZukHZh9iTh
H2w1/VVIIulbLkLaavcybX+OsTfruH49jm483HFIF2TvH5PDR90JW5vd0QkUgrfP
IcHbZETFKxCT5AugaYMy7Ckm7gD2YM4PJ/3pFEVLk7j05ZCB51zXUUXwfG7/GOo/
PJHsRbj/M9pjEYRAyLx2W4hUv7REq18IwMGc2vHcYiDfgrqisqggvbfsuktyBbUr
XvRVw+oAZBQih68eUqElggDK92jfzH7hHnEGwQ1eYLKij+Aca/qp9v9QBEHDY7cZ
ow+0xx8FosdmmXWH2NyESlo+WAqzjlZkqAflX3cP0QD31zvvru40zgBJigg64jzp
3oI5eol2RyjMrbDLc1bYQfjcdPolFDEknjxp/nOfMS5BukJlKQEBzCU5i5ucpsNF
15RTZ1446Xv9JGu4Gb9XJ3zmYZVXorM0cvK91ZyfRvOskhTltzO0/3Os3+6GZMB2
5Ay1oEBQ3AvItdm+0rTmOOg9m7Afq1TZwPJLClTpSu3V+tbrj7eNg9jJZN3PQyuz
IIJF7RvjeBl+hiJiGOQxrk8eY9TRAPf+JUiVqs8Ut3/cTj+ldqN5DZMajYVk/Chd
FilzOKM3QamthPuSnErPyLe3N+57qh7Vw84bqRtzHhT0vq8kEztaCbOdQ1ZbAKLo
qyyBN/hJx4zKaDnVA0cBiHtVbNSNRWzXpY2bGv7XrLlQDNq2nfvI5QEZWgQC9QbR
h9hlkcuxLh5tTaDM87SgMGDc/XIsAV1TX+I/JcqBv8bnmqVNcTMPPBACd+qMllsg
2kKdiDEp6W3ktcbZAR/kTpQc12c9lHCGElFRLBMG770uiTM4IAk5QloVhOMVAKPT
gOh6UxIwwGZwJe/7aF9FzyYzpXCoJoDZEN4QKvpdDYaQfElRtDgRGjR6wVLTOzNk
ALrwuC/WvTEEavtGlTZCl9up3dZH8RdPGIth9JYZGdp+FerPxcLgsQ2ebGLN378n
kBLi0TlMrRzW4W5xNu9Fy1Fw+jgspg0bYYJ0aHpE5HF0JTyhhJQoMRrttO8MJXZP
GV9vmBqH0QIIc6icSanlDVR4Y0eDLVIVhz/XpMAXFZFdoiu6ffnbvBrt/sVbYhxX
1pWZm1bDzhqLNdsEc4l8GjAPjJn80A6jTlnt2wvAEAdh230j5+qoJpimcmzvRyiJ
Mw65h9U8Hru1RmxdjepSL9NlbkT24IXTQZv4WYUMhm6iMZmhoflDKaeF4U0eXxS9
uzxba6jahvODpbuuqoszwE3/Xs9PE6CYepEznY+S+Q9LnytPH76xid36J9dt68rC
dvrgwOStVT8znGcXL4uCgG0UcgpqpW30h4vZGnHR0inDenNDsWJWFr/AEpy1AV5z
GuRhSfuELE7D31zoZPJcoyk5tR4n7cR9b0cXBlip2dWClxeD8WT1Eda0zzgszgpK
DoQTtOerOl89incQvvt3T4aaBrrYqsfQP1AxmhVFG5Ij5oBRZyIdN5lEdCya5AqF
7VPPPuyVqLGJt5UjXGNuxV2Twf4Ei5sHeWBDSyLQsW86fK8sNWeuUnOGv1F3Vsq4
Df8dlSTbPoLE/t57jr0Mj+i9TCW+FTFryhU3/WznAMwQr2OepuuNArpapIlMFSP6
MoxB3/dKk9njk1cbpR2oj/fw8jaRhHkOnJC75e5A6EKYLCirlOqzAX5KsEZKo2Jn
uMynSBqryuUPlHSo4CZbsY4Wqxq0WuQPD1qykXSFHVm5+7lL1Os+qfTGBX23aYjq
gwljkbuv8JVvc4CAAw1/xIkXYfQ3XgPU6r6iFXXCZLSZSKW+U+2stYmZPoHLYcgf
O1/3y5rTWOH8xeKWHvCCR5W+VtwFRk3sSjrWLUk3daq/XHJ5UeVvqb7Cs/oJBiQ7
5N0die6EkQ1rzjZsf38RpmWXjWTC2mALWHNemGuGKuwwdMDfN0cHmJKlQCTAkg8x
XaozfMMiGCL7VsS07WdIbZ8Rq2hFSDkaNTd/iQH3PPIhY6MOUjWwWB6SB9AIh1QC
fldncjdbtukUZ/I/2QH5Eo7k6yL4nB8YuQdcDbBR0+9jLTUuq8B3v/HTJiFTg2PP
OaLejeECpDkTZPGzUXDq7Nc/AeFyO6bHv2CNilQ0z8wmbGdQIhoEvr0UBO5dK6xd
IZtfg1wiW+Ax0A+0ZmdgfP6Pn2j7Z8TcThWXEGG6d7zAxK9THFCk4iwxbABMJ+33
SV/nL1NkKGfQPFNDWwHuWfrre3WBdG+2d58IWv5EsZZqWGm9FERa4GsqxnbNfqWI
1mC60i/+DcPBzk1pL5LCeN3sqZg+rBKHkT0szS+02kEnBmyv7xCpoGBZ9Ql/+wf3
4cR7y234152VFHFGl06hwDiNXsuvLAyAbUv1bBvLmnjY+aPTeTuHJDPemTlZjsSU
MykhoMt4z8/FloOs77u8PHSiovs/tst1zez6CsDd0JlxpZS1RY9rwmsaIf3dfySf
4TadhfEaulQFMiTtqhEe4hRZpVwZ+TtZZ8proMCM81mdPTanle7gMQ8UxXRs9rh3
qFHAlVWEDhmUiy7r27DKE6sPBFXi/7sN83P9lDLsNMs/vDgdnbrwwxKUMbV0qjER
fNq4yWHOnh2q8Obu0CtHWEOt+ONhwWwTVcVkJZkRm++GBQvXQ8+wpcj+PmtamftV
C56M3hOfySCN4N6rNUwGvZ0HOG5DSClxJl79jgvvWiSAQE8+KRDz8re6sjmLJdA0
q78rA/jTjq2AcmqWR6CT7rIKSadqEvluFw3nKtwojuUXfIV6DKmSVYqMAYSslUrJ
P9WLS2oIt1mG/6euCr4SEGmgIY+EwSdiJZLrFkDIrkwlQaSUFWnlAXVeBqdLUyhZ
0SfryUw/UfZ/OuAXMYAB0QE5p/vVmndhc1CHhHFVBhW4uyPhO8VM+GpWXxQeifjk
dLWXK1u5+sb//odQ4xnrwiU/PoVQ+ApDUy6kyBQinbAGeAL6OYx88Nh1NFBvc2lL
PmSZTa3y3SxYOMsd2Q9WqpcC1mRKD1OtKw2mlO8Z3freDNAyw3aaDZ3C1MvNZhyY
GyQhLOlacy8LgRJx6bs2m1A6b/w68jxgSlzKuqi4W9esB25ZtJUxz1hgAkhGKJeM
DDkh37tr+eiNfTAgbhXCsmnjMEKL1wmgNIptdQwwxoHpp0UA88s9HPXzKZJ0VNLx
hVaN1BpCCjp6cWHEnaS6Bs52mGP8VKxZJG8XEpZJNPQ8J1Km4zbNzpLqEGl4SSav
Ft6l6dlB0gF7Yb03UcoNiUp4xnU14RS20s7UOa49l1cBR3ygO5usj9XZaFMRdIUy
okhdhrE31/x+xOK6x2puS5DSA+RP72BIOm0KjMKDdfzHBRddpZMfwDMwO+/Fj1Iw
mfUwlHvCCOlHzfFrKo4F+Ueivm2WvXQP5HDArQIc4Bl/FtTEUweZF/Ew48opmzGI
bSSeo1je3zRqYB2tFZk8WiXQKMuuhiZBCuiLzTXAfgPmnRlJwo9l2Ub+bEcS1fRF
V7M84CR4kZRvMHTFHrkBfizEnY2feaSL6XI3lQeZ4+2tnR02hRRt2OW0qQov1DKt
qbbOWjwqrgv3b1yovUoNpGjfYTnnfITamxNUWW9qbEFA1ko14yGn4fPrm+0AK9zq
XHsk+Zqy/cmwlI+st7BpU+LVj3r2SaS080D745as/y3o7dNOtpjLlDgMm0lRt/Fo
ZIDqedUm0dP5psFqPQKh9hvRL9wvWgtACNhhOmkqqyva857TlY+B3c9lbdwFX9cM
zc7f7flK0xJ6Ip7HSYIw1YFKhUQw6BioZMB8pBsMhsskX57D6S4Z1+kCpp7Ns1ms
CJtkrTwOvIxEjwzJZWE1NBfS7I98W6yOoEFC1w4efjWGOqMjVQoMADLRWyeAydCl
iUPO7IqEOF5sJIlZ8gYdTfI8YQl50RDSWtSpx4/9+TzAt5Qke4dIZ9CnbMWDTBEo
afUxie4o/ljhJD2CsEvh0qA3/YU9IUYUtIFkthH281xmzE96vktpXpHD4K0ndD/1
QfO7iQXPkHpUMBBWePE6+77Ok71mNDMyeVBGH+mC6w33IgDWCaa80Zxkrvh9mGfM
NfGq1te6TG+Y8kT5j3g0D03QvfmS3uxks9lDX08aM+yk/3FPa3c0A6pdsZd8Chqf
YIgV/mGkRHMBLe65fJQnR83v39OwFTVpQ2Ox39++WS1d3U0/8MaYSDRbW704Rcy5
4tF62vTcg3cNK7PposKZZm+fNTu93SYlhmGM5NWrh0bHcYiKjqSfPjx9kD5O1RgA
dayi1EmbA8h/vTMZh7pNi0ztKhUt45rw2K+nNv3dUOF50pmFHfWVSNRA8X3Mjtmq
4yoJMLFuYncEE3/u96DnmZjpENodhfvFncqoi4/ae76A2XGbKuk7pnEHtoVaWD5W
upB3OUz0wUoffUylvJsZwNvlE2TMDTHK8HZyoFF+uk0VrqPl4fks3Pt9p2G5gd/u
DGJsuH4IVM8fsrL9zJzkJ2V4DfDTRw/vxLG+sPrUqydL1XLotQN3qwtCOZqWQYlZ
XddcnKJTq2Epaah5uzuzwgm3ohNm3DX/1rA946sNKoYtLnz1firz2dSz7/18EKCK
dZfOkDCP8MOoCvVzl2tjbgo84TekP30b7vounJynCVpWOkYZNN27mmL4/2Hpqmxz
LWYFIjbSZWeCLOfp677XiVxj8KajBv3QdtdX6jtrVDOVyWdi0T22PICOVKVk2PWt
KB77N10H2pKHCnClposmYU+7XnPq70880R3gXUlNfrANUWZJajUfWy4eraGSxu1t
73ip1tYziBE4aDSjessgxAYyTfLtxU7URYDDSDQurUTagvijUuGSgc4B/rvuhcLY
b4Lv3m/vay6lCR/clUj3ZRH5thVoO2gaCtrGUbNFPMzvWDmMOGUlN4PDoWB/xMmF
3yMhwgkilKhmhLCihYc6RT5swd481b3J2kwwrJUwwqPRZzYffReS9uvmpcmVA/a5
YQgLg/jZE5g6xq2g4DkXHpK2tBUMFAuiR93h3hjTbxJqvkVP8nIqIfj58PFNRpbu
GGiBdVyPNzFeZ3qWVO5cxQQYbtb0Dx1LAZIpA0Vo76UaiYwzamvlXQ3wLmJirwbq
XBqfaYOgskIBYnjBviE5xEl8kdtiBWWRH7dQujOvhMluxcOOuDGaoLivpfeorQKq
c+XikNg0SpYR7D00vTKwa0VEHHmrl+4bWgBusNiXNkwrDUp8I78mOPl56/g1CZfk
5+tH70Wtbg/pWvIN0rw6kEXeHk62qv9iBHOufPrS9ZATOeYZ25sEshtMt/4JE8oV
rj7VTSlLpZc1Bnomvh/R/EKG4iOW3f6iLqSKHteY/aOzwSo5P7aCNEudA6YhWFc5
vSeQfYYEWgOT1JYcyx1uQPTj5a/+/O+Nu2mIMzjqV9LtthRcui/BSOsLOFXUonFy
3TtsLJOBX1o35W4PAHqhW96CIEbq5zxnRGNxWMGKKVHxjpIVciDzXrRm1ACGwa3A
FSxS7EC63RDKDTsXwDVIKUuuMutHSP31fobEg91e/Yehld3fd2m/ROoXUMkBAOHl
nwAUq2kuAVq2MURIPFDbNlxXXgOXDqUlHS9V1o+9p4zUZXaa5Aj9CjPIOmypqe4d
QyaGqxif7YwQhhVpIaLkDJs95xEdh95oP14rzC0XuboV9uZHXwHcrX2UopVUXDkP
3S2fT9INPN4w8apVF67Ygs2FjTnH/tPAVlVAb1rs74O2Q4GabyPf7iDzbC88shRX
dqC2GrGpM5P4DIRg9FMdueok9WHctuzv2hWHD79SNx/4GrGMf6yfvfZLNmQKwyqG
K3GyH6S7s+B3uNnGJ3AvCV7TtLJcPK16WwroXwRngXMlfQq5IoyxW7r7ME2C8vu9
OvokWeuQdyeyNe22rUUVB35DzVh13K04cbUnetXx4HD0vMSnHyfQFISGpEnfGDjT
KJCRt+7wOvLKTxBaIvsCHQHy7x1ItKlOypyFEjvupg9eMwjlnXJJq48nxna/nec7
boRSttEbuTnjiDJnuCv71w730317ev4JPqivHM+GggxmE4tDt2SHeuzOM+bIKwAy
YHcMaLlGkKdZ/O5PL8vkCTlkrmsUKpoQeyBXyCP0xF2BmUkMXFbXOzCeHTH7sJfg
HTQhhhZzl8igCkktB1kfI8E/jUP8paWZHwj7DoDjIeO0+Ahi548CVIB3EIB6Zk5c
RL9ZwZfWJwjXQYksK2f+qDHA4qMIT55GzbjDls2mSUuPSjG1G0wpBUY/uUvp8V5i
MzkHjLcJzACAsP/OC4FpV0qJCwGqTrjPXKSA1EXtxA6/Y1CvX6FlWH/dOmvpozWH
IwqOdKbf+5EcdltFGV/krzZm4WSORqLJ9qnfJpneM9cicUuITD0SZUi3jtFee7la
JCOtPYepexG4fqqS1nrivE6hErpzluiKoNvgiTpaLn6HT55zvQkHZUZpk/axAtgd
PPSHuzwwI9FPkmp0mPory4WLtZomDI7tQNYbE05Tk9/NJaeUIx/SQ6p2K6r9D6GH
AA6+zmYLv7+2xtoJsLycW504MBVrNi2iDAVxJt3TwLeryGw8GwicBTzQL10Oam2C
bslHYp82oL6gEfchPli3kjxhg4ShGjfvDHUUbvxJ8PA4Td9bF6LgcbUOZrTlj7xq
KkqltjO5qLHGEtW7A17vov+J8arNIVcHgO3rc4lkSxSjFPT1B5O2T/oN6yOCDdB+
SbmsWLuD41K/fc5c5eWKNUC4RdKd3kzvJpIxVPxFAsHVgVcGDKRskRAOHgXAILW3
ss1aLtAiTmkhZyUZnt4zqtNUMUoqBJM/nCvynylibFHkYgOsr5NUDIHUxhgA5LIG
49XUy4Nh0H2lbJEXGXmp4LNyYzC60mnNVDeOY3/2KpB5j0G0AVilb3sYQY6lsz1z
T9ekwhULqeIk11M5H95gseDjYwFwkMTTpO5THS0nrm/ydPLs962/ioE9sLqAzNQ7
lrfL0zdMUj1FqDmxjHAeKbW2+CPlSJUBJNfX2IVpw1rxUeDScNgvcesY92+8I2g+
GIZD2UM9QaMyMaoL0sK4BcjvMYtT2ArIRPP/mrM9njKOJU3ANwr0ilLHQysPcAbl
Sf904+4J9PExPkeYFQiTNx/BmfG/K86ImqafsTw9sPbwndfcDm3bChQyHqKPpyqp
MXoLLTmR0ubFIsyYEA0oeWBYw0tfBsPehqooSvW4fNHJoQQ7BiEIy6FHndnbf/5j
TSq7nidRQ7uzi2c1YXZ+dVUpvvvVdSKQcyUwE3QWnTYmqXhupNtYs8Kp+keP1q4t
lWXf9FE5QBMVtFGzn+TRxjN1pKTkNco0G7eyG9WtzXYfOFnXt5pVPpttOMOM6orn
sKy28ROj2PDgSdTwcqWBNaDXq5WvZ7KBozrn/5ZRDonOwTuQrr3Hl6TxMLluyVAp
UmmmkgDON2bKaapRULZW0b02oJKzx9KRjH7h2ZGZMmpFW1se2NNwMdsCXIpbRTHJ
JR+R5R9V7S5LPjeC8qQs6ABVuUuDqM3E0wrm0O6eQLo28vpklaGWciVvIqMXGo65
IFoHQDdRPZtoLAoXFzvPCZpDHysnqXQEGsOxF4hPtvlW1PMRim/x90unL3RRfB9m
DM2Or0QAZezh272hZ6OE9yXOA8XAgnhvF6tdccH31LP9JsY9MbRNo5561Nd8mSCa
UVVhiNXYEXF6b5oMf6WAmndguWMAWzoVIksgT5mK8ARl4pxL7xudm6B7Im4PNReS
ZfZqXWb3sEHHLzh8AQEA1A83xiRCskRi2Bv86C9hmC+WhbTwC6cR8ooNwH+E+MzE
dYwV3UjhoLU8G8dcjlAPvbgsYl/zEBbWjnIXCxVvihkK9WG6GR0XOLlMFPO4+9qb
3Pjrb31MleP7Dwo1IjnDoymf+zr70uJFVJYbqWQ1H1k8mEzgxuBjCGd8YRui6omD
BwgmrG1drMutnitKh9aS6600zuhEwNDS7e5y8LIdZy08roRqQh/nseW+j5saST/V
ddETXWYSDuhizcnONjRWiXNff09GUPBzNYFSkPdn1cXj9zM2jSPdHVxdi/0n3Pd3
1YwF8nAZ1tCDkloWLGKeYAcDKKDl0axhfHNMGAjbA4bqaUjgzbnoO6O+XKRPtW+H
aUAeya8iX2hNVWAlKMU1rdAeMId3Odi7JTcAcchIfICjTFT0Dju40mmd+NyzH4FO
dewIl6Y9gaPU/wLOY7DX6pVG+G4Cc/GX9nnePp6dOpqrer1VF1dhf0SM+VRfDnXY
KnDCzsmHTEnZ5ByNTiZ7f9tENfGwUcyXX/Zd1f4lJRCD8NLEB8lp3Pguhulmp4I9
2/cEtWccOlEfk4LBzAB0dAhIXueMCNmtv5PjDu8TQ8OlJAapx7xWLD+22FIFopob
1XhI7lpUy4rV5v//Raqo8gjReuIcUvsBWo2PPxqnyaAI+I9NdZqFtvgMBx38+sWH
pY3zDOOoPL76WJAGXcnvLJuPA8zdeocF5sQfQUPN+sEOw5jR9mqT/TEmoG/vPzJo
ZJUWJPVgDNtw75hshsN+AGNV7H389ifak6SJdc2KniVkHMQRChvbgfJnM7Zuu2lY
ES8zAU5JT5XMWEgoUg/DSelFB96oYM0g4arYxEzfkZ3//5Hdi0BzBEoLhNATuJH6
dZi8/SBNO0Ht0n/SU+zf1Wr7ECBrv4eAxFK697E+lXxQd3vkG5Dn/yb7qkSWoRqn
c05c0qKGSLfncXujmMfhGVbhJ78nLR7L39qpqu0vAu7EY3ybqc3PuF/E8KuKZ93R
xHb18wdlN7zfAVYtyf4IDd/OjwTa3yRq062M+xk52JDZm2wE/xctIhBMySOoJt0Q
uZexTYsuM5lQLqGFi5oa4faeH09nAtYIsLpTEmFD6pyA7M6Nb2iXaWxO1UxBxAtp
BBT2gMq0bnQePg+VMvkAJCeYg0IMo8Hdnl3wvEcpGrZnbnB3+obt8q+6kslP3d2S
vcqfEJ+I8NqlkB9eSzT2mWRr9pvzrGdndq+Zk+WwoBKVKvtmeeahv+rXUZOXOYAs
2//xjYwtobevvxAC8UjYBzK+Qf9bQIj7BukgcxsjKaRNlrQw70p4rH3z7WnH0Tk1
jNmBxBqRXUi63rHlgfjVV45fn5AM3YnqDpq6EUjD672y5jCUq2tVXPavHDRh+PSb
xrEqCDr+d2YPSLuuspRrw/y4OM8DNKNbHsXCJqFyUHnoy7WAVeAgBfWeoXxUGm1x
hBSI+eEEhtryFU2tbI90VYaiTjjwGhM+jQfneb7QfnHW3ahzKJkPMy7Igh2Ny/vJ
9sZEAQJCcL4nOdX6fj6g+efIcFyA7ALPd3S/zPQb+VbQO1ibKl3/7is5vvnH52tK
/4y3e2JJDfM5gJPqzkazHYa95MJ3vYORRUHa3SGaNJ3/OLbDMuSuU/pKTOoXIENk
8Dfa3G89+CdiLZHrOL4dTkvZtFMD1seAFC//fTfWP6XXQUOcKF0Wn2uXVrTppctI
5DXHD/HVQ8JZpgDXGse0GPB0k1n/VtGKi/9kvn4BxBCkpBWTGQKIOCH8KqkH/KFD
cwg5zKO9RzhUEMygsyiXKEavDWR/oqCmNpBo0vj7eEI9ETUXObUtRqRamO8XSHVJ
5SYxproEplSG/0m0DqPNxCUuzjw6SjIAFkrT1oRkMFb0wfqnRq2m5++cSAzTuyF2
Hsd3Yqv+qHGAEMyyYsTUpOjLBdzRe3Kmlgvld3s9aEzlO6hnwvfa/LV5N9YECem+
ulFxzZ0Vf7HEsOs+ed7/v6/ZYlOL+13Nk47i0l7TpEzpDaRt6d6g+kulYk9ZugX0
TxSMznxzCenZuTm2YhHV8I+GGLzMHP5qEsk5YpiwgiA5YG7Na+gmJqS6sDwcvhgX
2l/mVYG7SCAE5aksFdQ/jWKHdkU+BHJjuwlQqr6YzHfjQWQFQ+R5xfUVhkqPLOF3
6kcf4wrDDGPVKD37uh99zJp1mfHV4L5EAlvoMUcGo/AbCSrfIphsSPxCBhCah3Bd
XPJ+tjjbOLd7HITnST9N/AwlBAFEHyswdGUuiGFTCeSWCKasNyjy2e6Q+AbyLWba
Lj01MbiJ90AerJiDaJrWvE5tI29OCAsH1V3CH43xzQ742TpgpzTyd2F2agfTlh8R
IIksWSDL+J2EJfsClXpNmnR0RQgyy1dDhnlXoJpaZ1tqt2yx7aZIUjfy4Q3W0JVI
CG2qzGXZKYrYwjEuRnk+Twb2VuEGVrgLSa4o2omLw7gwabkp2oHWDylLdVo0ytU+
qaUwG7N/hxo0OlvGT+NUMK2AGXKlJHbtoYhjyqRrCcCWsstKtX1mSM4aNym1ocqj
v7+mgZsNnYhlneqET5cmf5JGLhStS2nQnlhBFkSH3tfWEwDv4qwIADdDe0NW7QaY
r6ZtepI5Vv+5HPz6tIKcyDd34ijbzuKSfnwtWjeB0GzFaGBlHdZXPbHX4fWjGL1X
D0FsrQa72JpfUV3qkPRPbFanKF5x8kn3L2x9O8+Vsg7s7Lht7Zku9b/bEZWs/M5h
+Q0mPj3R/SptNSSg04Y7IGwS636qKfYa00ZPMufc6qtQiVMWW+Ro+UJrqEfZXMfL
idxuxMRP74llb97Dg0+8kf3tuVmb8Un0BkzIr6CzvDBmu5W0Y6j/jUWkfQhrKvul
Jz+6ECtMfwveKoiyOYN0R2yc9qNulbjc/PdRka8IBRXMl1simoc4Akf7RlunWi+J
+M/nawsVp8R3AIZ7KkpkMhy+T8FK8IftR18aWTiYrvjxAFB2oPIh0aIVTlW+rg9Z
a/z86XNHv/MicAzM3YjP5TXevwVGxrFT/rrHOEyserHc16pI3vUirkJP5IizKoJl
3E/2Hr07UA1DzbhtysGNsGCD4LjGtLg2PKlY/aRZgQlQpsu9Mck0+9drUfSrq5yu
XlURsKSyZSoCChgnG+l5hOMz0e80SG7rjl/ibGbDBojJBRBOhGxc0EFIwo8b7RGx
PVaOwiwL7HsmxSHXeAFhypa/xJv1L/Bi8gHcJPX/T3Hk7mmpeC8joF1v6Jxy3N3n
xZvyPb9TTgJ+wJoy4PhGGmnOJM61hr6uRSMRsCXfha6BqqHd3vt4g4Kq0zLmQBke
zjRibVis1KU76eLf80qHP1njJiUvf0aLEqlY5AHD5bPs6Hga+ST/YiIxXZRiHa+1
3OwMT6ujZK5nXSD7A5Pb/3236zSLdTVDMtxHnb2vd2wQU00w3vRKV1KagayTkUPV
PwcB0YQe8IkdgMeVR9PHpi+6NmcVahR4v4k5/5wsFhaEasdpJ7yah7tPOiQHeIcv
Kl5Q8UD2X/3gcHxMBPyUMAtDjOzbXMnm30BgGC1FIYMTM8SrMBFhsuqlHFsJ+iMq
VcH1S07S1DJGlJARgPClaIkphTlemEQqV8kEsbhZ3WbjBoRXDlKje/sUZIzDU6qJ
FRaY9xkjsncrDUs4kGkdc10W3DsFGVA2J77/zyL8X1To/eJvy02UQ1dq04VcfrM1
BRzacgnvDEPKcBqVBYQfXdrDoVtbXHvLfkR8uT1sR695LgE6FifIWDH8OvcjSr6W
j53yQA+zKbOpKHonRbhx93D3OO0XwUrzflqBcXEcjOCpa4oi8YFc+sI+hv+WSXzq
07y4o/M3EFH1aVb0CowHTg4aWoJW7bri9RkETdoH7Ysq8tsqQ6Z6+vPMFoNpgHGY
iKw+ZgTRuO3qNrHvvZkibwSQeCC/DF9/r/A6lX+IjkUSaY09C84yWiKXBLLNxsIC
bNNCJzPO0gY02NVKL6lcAcRG+obQok58eM8vVWfupdpcLJzrmnCMqjhiMYdLcsEJ
lEz/LyMQL4/8hTBlwgN6xpXskx1bucXt3++yYVcTAJREP/gdVQsOHlwFBlNcWQmU
NyMXSkoU5ufjMtgoLiXVQKk519raqyn86t0bCj+kUF6jr4DWZk3OKWv3EluCtqDO
64B0K4aKEJxxWsFbUGOfyvi7Q/mXDVWK8um0kURDQJ38/VnBsxr8GyOOqV1oYo/8
+V6cXs6SG/A/3PdwjwD8Wd14VbSZqjQEQOzSzfmUCDVzRPnE5a0bwJbhfC7nDgxt
7ZEwp7wGrKW/JFDwjqFq1mJ0Srb6d1iMCES58zsdurmIw7MLHYQrvwIoB1AggWw5
lK7YwOwio1H5adktCFAL4S6Hi+yAHUbt9CPrTFX7Go4ygEdCGDdQVNNl+E9sAP3R
hizKeX+Xo+xOvho5reYT+BDXYKEjRvYZrxuRUOVRvF2rb6im40eOJX/sweaJZUUA
T3cxo/PyweHoed8NtN5iR2+HhjMNJnSbUoULKLs5JiH2huD9GsHeB6+CUtDWBnXR
Eny8NgfkdNW9IAH4Eej7QKVvSyDYvyMw8zdDCvjRsSaha+zaQ+cekpYMkfw0gpuA
5r7H05Mb/f3hl7lvYC33tMLpB3x5LBkmQAYpZaWyChoCRXaqkdwBIM+tTcgb9ZR7
NEq2YpxdcerZ2BT7t4Q2eNMlWKKeFaL5TyJ6nwFbZGZBLVYL/nsITHPQVRovmm5Z
3S5TVdbQjzpTXkQCwMQGht3Qt4G7zDqtThB4DcuJNiLRPMk6vzWJssrgFevGCaOm
q4rRQG6XvcO4pzAUEE7LYNztgfXY7KrjLwGa3CzBsELzo4e67ZiBtFuon4dXCxKe
M3/YiHDj4eQTFQ2wfUkkrY4SfZAb2gC6tjzNXMK7PpsTRv7sdXC+zJKJ6BSm2z1X
QQZ0tYmODHKOpG2or1ohx/IWQKw70S2ovz51+h8Og3AHeSONgtD9CyKQ96ebADJT
bKG5HnD9Pqk+LCRru2ML2noDWYqFR7sxvFN+kh1RVQYzCNrR/hfwG/u1gnoB2fc3
KvNqH2skLCTPsVJttyHue3rK/k8lTBpKMJzF+JmTHWZCyIMM0+9zKLyOc1REBIfd
smrLZAyljbWL1S3pz8URPYR7JddaEhzHwOidZ0b7uerTKXkyOlfcWdz6UPDsCBjZ
LwNRAvE+v/xs8dnSQCiWC7O3Khl7bS0q3ONROxuw2vEZXmiX2qrmkkHpIY09jHOI
p8F2z9agxszylEovFr9cfOz6w1fZPEf+DrJskHr6T9kXO3IhPLiGNwpQptzBpQSs
50KGfCJS3PJBvTuffTZ14JwXpFZAlLU7e/KNlfnOLmi/ZNYbIaBnQWSCKppW7x9n
QrwuOktXqJY2Lxx79pRvmCTQnFgB4MipNVFus8hZ3Zk9TVie+1jrqEkt70/mXhG1
y1AGTFoIIvtfhNYYhE/yKxrdNcEVYnSSSWoWpzqaa5xRjkLJGVxH/NU6ghv0wVjm
i9YWBg+28Hwhdg+2VqLn/F8q+Mw67SziQhxjHdKE9HKvP4Hcc3agju9KkreeRyZI
gdAAePqcoDxOYfNdFi1L2rvu7aJ/vfUSM64FCF6zKrNwqhJRJnOT5x1NN/l6hFyR
3JcNyQq6x8xiboJr+fvKvbdEn5Cv0FAehE9lq5TFgTO/ggOLzy8Q/g7VtQCEqpmp
45HYrvZVsor5C6xsnRLILgKFcOHOiY5E35ECqfbSga05pwwrAcsGmCOMJXAtBxMI
0cipD+UIfylggJkZJ3I+GbcdYlR8l/CRLDdlhSWURppA+RQ2JxnnZgQ9HvAbo3wx
OV6CmkY/oryAqLjkz9axaUcFX3dtSBwTzKBiTOvlQDP/rq3x+0BTcMj7n3CUn4EK
7BOVteihxrxpSynJj+xbdP+Bk9yyJnYKwifk8AI41GZA1wrWK2mckfHZp9kfp406
DrUo9D32r/i/c5WUfzYt1M95qkyGpmyZxBoicuRDs8NSSHt40mzbgWDuwLIwlgyM
xdnO0Z9vHJEhiFwPn3rbz2S8/DHIOyGkgwLtmWXK1ZygvlWSbjH5My6eGOI9lbbw
QcToIi+i1LPTrbvZ9Ya7JJdJWcThz50apysh4ZcHyGEGcMBi6+ds+AWi2m8/5TKm
gwJD6y5d1tVZcTriJMAVb1K7VdE/J3J1y39SoXOrv0SDU+olPHT5gCw50Y+oQJGh
Di6jZ8drErQzukXTJzNYLfLHsU9K2pVgga5Qo680pzE0mZnAQAj09jiY6CxysZoo
085XYh5N5Gn19ZDf0u1ab5L9tieOoDMho2R/EDKfEN60MUGe0Rwj1MaZlfKsK/Yy
5Ag/8vL5PnQJ7nUsoMl8uwksWNV9umyYjlzFKaJmuARD5jI7tO/aX/vKF38BZYn4
jAS/RA6r5BUDgA1FMcv50Dyuhm5YNwu+p13+ih4EvRGmWEKowj38qVgY6fno2TNY
G+mcM9mqh0dSaiLNGVKrjMHMikF/rvb9d698TKb5xHCpQaNHK6tIWtwdz1XhGWFu
xjnzJLqAvdLiCmVQXBLoO9vgGmVmh1XNISK1SzwdG5PXUvs3001k4O8e2RVbWTPv
PsA431QX9wupwvKqxuRvbWnNe502e/LdGtigAbEbxpbVhPKAYAdnyBnJMg4lg5Za
FTUfdVEheNL+2cVBLO3VW+Nd5CSUYNHFLDOLgGNFwq65Uo0QgaPsLwxFLSKhDAx2
Ert2YZgSIGnuyusb4OpB+URorF8+bQOZ/SvcpFZzli81DkMZ9q4vPCReMWSoKUqC
/SqR1Y0iUOBrjTus2C6O3IEBaa3UirzTmedlYJs7QIC5D3aChzWgxIq5563bAw3d
/4o5TTfYp4WVn7vo2zd1KPvO+1l0SuY/vhD2wphaI0ah6uDvZsGEVdpneDl049j4
aRzx8pnftgxYvoWksq80SoKTzSXJnaZi4pqlVc0UHGK+peWSsi68FrAZCFYqjJ35
OhOyrDfOx+dTR9co+4fsggKXws1zRJevqJ4BaCiZ0zQeW5WPVUitz6rqK42uQWMe
tMQP4xPZfPVK/z4xb+FwZS8ds9dYTmedJNM597z6qFEaAupjDKIORm25JFbEIx1N
3rLPIpa3HdyU1o1H6q0B32frlRR4sXXHG8fKwqrNM9z7tuOYdzqpy9CiJ5WH1iu+
CPxEjXtK/epYCX3kg+pD8TIcMWJVpXBfbyuAev0fxLc6jGQMCgc/9U1NheEFoid/
IaNei+LDQUrVoDSEwcX+MthdaorgOt9gJo+PjugxvDNUMohP+Mzk2HatXDbXVi9b
tJftgq3x7EI20JgXHHnvp5ryevfjM3tYSFD8AZJ4Blbzv+ti7x+PAAB+nKAio66S
/hETs1+eUQWSnqo9irWFWNj1b46jx/hStDxCm3EXObVlVDsl9u6T/4PbHNlAfMIU
nDd7LnWz0p9EGDYSxVX1atvb+pGWviB+m6YHflpQgm3M6wZsN6oIZ0eGrDx5/L3g
8ndIAFZKK2+jCrPO7nMT9VeEn8GyTe1aq9y9r8Q7sH1/t7Oj4zYnXJdaWTwmHGKN
hL7G2oRy8OyrcgHaoYBfh0Tl7b6Ns9pUlPAFkz8fFaU51+jm8sEgJN0J7mZtNfzx
fVo9eVgc7ltG2dzBGqFQwoN9HvrtbwMiwdCWwFeLx9nHpOm1DiGcBh21V/1kYtmW
Rdsh4JJFX+AuIrWQw3GU7zIRUPK4682GrFQ0zCiw8D1Hkh7sKyCpMCQeGSmr2X5s
7uqaa4gkpFTFCkdz0yxe7PI4NYUlPDkSOqLJfP1Q9xvlCgxMfBOGepWSS9NZVLYY
5SAPrtqwjUSTwlAJ3b6mdJqoYdDxQJCJ5KgyrdpSXtd9Zks3HsL4Vt1UGgw4Zio6
D8gXx6+2P97tlOuF4zZJmcXYYMe/SruXhXsVxi5SYTsKDOu6m3BtwvMtTNaYlrX7
zNX2Wx3u6cf/fwjAYg/DsdbTPnXxVmLA4c+gP0b3uSli981JWUVkj0chws/RpGcj
PH7CQEO6ElbM7fXT7gRYnR4cF/24gNafDM+IKzcoLSALDVHrLo7mt8ODCCoBW78c
S00FgajJsGAyNJCbtahuhFOrbLrcZ23gDqCOqG3vEKYVQl5qE6DiAxcj9KAocSUl
goUCw2GX8sVU8GoCMWKKw0aVjuyYamitAVAr8wUIOAo57ci2UBqR0Z0ZW90WMGwF
ZCd7pDdg97hoG3A/0eZ6qBTe+j+Hv9De4Gtk9NS+cf3uGhrkVCugNkO1GTUDYOIZ
I0LnYuJpdcPZ7QbUlDPu+gconULWzQxw56CbNDZM/3M4PNBb0JoLKQs5t8yWi8QE
HThdoiRUGl8s/MAyufrepXXEuyP/ho0yyN67Jp40ZJkWcfwK+J3n5Td/+UQdSfeS
dDE6U2UBMkMMdvpotPdFWCti+xbqfQYBVs8ZK5rbKremGK8FT9Plr48E6QJzCpQX
7VrAdgiX+5Q0oEW9R0U/+bsilu6DJ9HgBMEHegSp8cNdAVBID4gnISmiG09n4DPL
qSUaN23qSr+8e5KWv6Q+UOv8MeqDg4QReDuMLDU9YE1CKrs8iF8Gc9bQF7ZZpHaq
qM9drgkMg7vNGXDHWMVrfGKwuhacy0TclXGtgsiic7O2F67Ng+460ENoo0ek7UBA
vpeskq/OFYLHlS37vDDnzVlocCg6hECFKETcIlbTqev1yiLFn8XW8H7bVTto6e5P
WGnBr7JtvmqtpIzPw/NUImGEBVEj8LoGTGMZTJCXesYh3eDWqAlAh+CzWajaThts
Lnc45ynyAKcKTYi1e7x47iJFW+zETZNdDdegJEH8w+DWrmaf1bXpOTeY9KuunxGl
gZKCcj3qJOByyALqjrRqeF6vBWFrTg85WWilG/K++VMpDCI+YA31lARIln3b5B3T
n2v9g+GK4Z+HWgaRVGVeD2T6hZZGhBwDaia/+7LhJ+hweHsV4zjGdqguqWO5fuDk
5FisCSatWuIL46CeZmlZBOJzOWfR9GbIJNaKfp7ojhLNq6euD6IiX1AZzDoOUFaB
1lPcnVKLBFgW/aOyIoSj8sVNQe9oNfn54OZQW/HYpLkUF7ZIAjXCXorAHuSsMt+z
lIfW1laHn6mlM8PY3hYOGs6048AZzvyL8GzuBijHKaLXWtl7f2+tORIk/Y/KxcRF
7ou0SFsUJQ4bYcITKywhM4ZiOaLdEcL32w/f3JZzsURtevHjUfFRHQl8KB5aDVMo
9xGbnUKMdRkbOCHVXHptQpTVVE9EbLWUMZ7VnPP0xTF9VawSXEVorWUwBxI4/Mdu
Elg7UJb5stsY2gIZZDpZRmXd5KLdAT5JsBhf0FOXxHCyI+HiP2sND0YUBApGmay7
v3phiG4thdKEwduXmZiEi+F/U97TtfeJk2gJT8EVwV772KXpyMNMHgN1Z40wJ/nt
J9vSn6VPe+ylJHLCQxinLrG/I/pJGr5op188KH709AzXBmLHJV9IwhB/gL0Q6PO+
XgC59S17dbdcTOqMyBaxE+d1StRh5u421tgveDlbXGijxiK9yX0c180pCYhUoJ6d
2wxptgCo725BlyzrwFdGLhOvBPzxvft+9Mr9pr1OoB4Gkb7V8iTAq0anENZHwH6S
xCwvQ/5hs3RzthH0BVq7lVQGOV+1+vDPvJ/xmgmhiLv8+Tnq3k2JnLWXIye5rasE
ndeCxc1ZA03kpWRG9gKllRT2hplv/uvPvDSNgng52HKcYmVyDBQYuhXUnWm9/+Pr
8fFiA5xrWp2oBDgi+iA7uclqIB5D+2PzTVTdPqPmm9e2uO+VZ1p4e/uuHMSTDkyL
NOjoOr6K9qmFKGpg5Px7rSdvufxZt2/0ZfhOrVLCA9a9nZOiQ2AbHvl8bFV/7+L7
V+3wvhoDPEjG7FQ+oIn9YN90kPFLI30ZbPlNHEd9Cq5QRc0O/61raLbNnUi7DQW3
STphuHTQbJoRe6IC3nuymq6tx72bkHZoBhMkIw6yo1XhkO1agJWjZNIOEJ1twXZ3
IIGXs+MFJw4WLU+tFWv+TGwyOIzjO14Md4zt+ZZG7yMhp56TOndZgj5V7ru5li1s
FOZnR+8/mSVpVzO1o03zchnom7vs9HpIvE2HO8ty4aSWmYsh3M1OUgOqJK6/xsIK
PMl/dM8/jc3hMG8IT93We2u+ybL+ZFuYtS9i2CPvi5fVM4FaHQnBHAXWG/LgRhDF
UqD9LKQeDCnTtAp7sttvhkaa87Vahjk59MQpPUgUzMDF8Ud/Csc31gvKdcGs8wB2
PhSscZW8MHrg/t4AleQGhWXMD15HycPNrgT8Q0qnjqG87BswhAHvRAStcYZe/nrq
WE5k3DfsdPQMB+7DWP03rzhLqZ9cLDr61bZAyq97OqGoBhc7rT+rx4Hq4YKbUBSu
cz9Cmht7rCNp0LPyvK03iPNJYK0kPV8yYXS5GZYwYNj8I9scsxoAnW6XDePix3sW
Ks/laFxanQT4ILlHyjoMuvNfxuyYO5WEBE4KIWgkh8sra5+qD8vnB4adYSBXRD2a
We+8nQRjfhfUXQUYCl0fVTcCODzuy3lzjbYVlTSC074pEKplIv757noYU5n43kOK
HTOQKXTbI7y/H9RcWv5e4+zpX4vl4pBGK6mmAGRPlvt/4nszQDojP4+X2buXER9Q
IjU26t7a4PFbYujAAXei/38b9IorYRWhkMU9NXwEqh1vT+XgVqXmxBdj6R8ugek9
BXXoO3p/WPGrASe4SKPPqIqh6oCVrwOXXmsDf3ZV4JMMr02gcYg8QMp76aexaj8O
W0MyIN/sh00JS8HlKKdqL5wHv9NzVDPYJFjeMXUPSkw7Qv7UwFqxhT25O2utfUjG
zNd62eoGEHHWpBD2wOOtOxfyvJzo/RYOom0l4kvXwGFPHnWNiVrO3HJ+McYG4Exe
CFfo+rDbPy5j/EJYizhmZ21VM8A6tWANHIUd+7JFaTNN8aONGWo1tTUmf8hN7yEK
FIl4AfGRMs/jDrc3LllCsE1Jv/objpZsO+9wWZ2a4X7aUgkDcI+WnQ5BwAigtKaS
BFC9EJcoBm9kjhZricYq1zIaILzZDE+Qf5Mylwj7846Z2e4JKvTxmMnEo7UPkO6V
stxwByaEqN+B9AZf+Jmf6k+KkMcJtQgwLslxW1PMqEv7lxEOJfCSDEwdPDYQY98z
Ydr2BR5AXtM4d8A+HnfgoaCc/8Qj5EostfvpAJ3vIw8QnhvV77fTSblY8itRKrbo
WkEfFodatfiUVxXeAdZeWLrNZKcNJEzfE9M0+lnDeHpLhtr3FzqCKDbEMiQwKzt7
5Ct3NRgo3fKehWK3n1TwWVygOWtg4QImsyLNjBiJCvmKTtzrTQwjaPnK/ttVPa7y
duIwlV53nAq8WByDyyG40hN9zVCtb3XivlUWbxsAiAPrLeji9EehuPPdw63/uT+r
P7zceuKmAVbL+LHccfvD8G+UkxDX9iA6smph2xahkBhKICcGEnqI7e1681Db9DY2
CHy9dTqVbi+dQA2jTHO6Fpj7fDQeaTFospWLIcRJbuOzK46+xuQ8siZb6JOxbwwN
ur+JuEo1tKTzu9de9NNSfLHhsJusPEWFkguZKfkG7H7/EYJw5DOBjTWKnq+KG0RS
uMcOOkX52xI4t65R0bwMEHWHsoo5R3Wip2TTHSY242VzgZwJj9IWZ379VImzq6gf
rAc5/ceTXemMLhs8q8j34nq/ejxfvPYxFMFsdZ9UodKIjowZU12JjhqsHXx4OQdY
ipBeHxwVPGIu4HeZB7eFLHkSQplLMsGWQb8/FfNh1JG4QnR3K1VLHGd0XSA19OsG
AWm6sXD+4pDN7FlIa14boS6YcivN75ID5P7ZBHSyvKAnmqMsh5dhpD2EEFKjY9f+
yKVKGEjj8mHr/BozdYK4RDWpgdo4H6tbZxIpFjlLKBjIm9qDC8a+QCWxqqBsYeZX
qb4aV/QOhBF5R8cnuq4d4Dtr43QU7ee+wRM4t0IH+TV4nIG3vi338QQP8TBmIkge
y61jLKfrdIqBse2wovb2qRZXj/vRq5FgrQ672QhLvYu6HPtHcYuUMstPDYUOb8se
wCq3r2oMlNUy82aauxwKZAFnZ4RiTsOZgHg/qgfIRmBo6BMA9Ehk93CZfc0V4E4g
LX1+hUwQ900F0CTO3le4ayEsDzOaZqiEW1NRrugVhuL/kqkkFbrq6XSp33tfAtOw
EYo0DoGLSX09xiNdlD0cCHpPHIlnOYD1eFaYtWU9J6+mzMzr6bbo9I4Ux8TFCk9g
p6BdDFFYsVraUvnJNujFjVwbR1De0uBVrM/4yIzERc+kePkQ0KGiE58S8qyL89g/
wLaK1drSsV3NG2qg9knaSB5f+imOUWW8zSLp/ZWDdRBpBs7hDCWAN6XPP4CBZdKT
fzZMSU9f8BOebI4fqCRJa6G9bA4wkAUKgz3GqgNsObEpGRxNzS2KTZ6pzNlg0B60
oyAVFG2HsQiNeRnnHG5AGgur3kFobCk2gNZVdogVSEAFEJkPzxMulLm5dOaBNP0p
NpW4+vTmCvhCfXeVBQtu/B8FgWzAx/ruMobalt67WYrKW1ZU2rRneTt0FGJ0Egeh
uv2/bpWP/H34i2TKVQeo/ucqqnZXCOL/BIlXnn3hFpzi8+hlI3ADZqMHNEPnWyDa
+XIa8PrbFCsDY4UFoW+gPiBhPYkVNy7lpEcIps0qTSDYuiKq7Z6xgfwul4978GlR
Q4U7/TtFgH3nsLHXQU1O3rMGBh+A8UHrXXM2ZpSmHbanQ/AfCjTOr6guj4aRm7qK
O5IIg1lDJDldahxXHyVeOH2LNrw+bg5+WTjYe90k9nJoQpOJoDdTP9R71N+YOOjF
l6z6ORf1rzA0Z8WpF+l684K+OSY+Ug8wUJN7pEoAUx0KRmJKS4ILtaoQUjJiTJv3
V+NR+x3iuft+/D7B3Xb+QAiFt3f5/iL5ggf829iiCnA5BDQof6m6pWZ55+1NbGdr
NoJ04KgH24KrFxUfMyLH0FFrrbVxwgqikl676zD6QPvSuvvI/fYBtS/D1Z7TIoAo
yIprtXbrdE6035Tjk5ECmtg7gFeNJ+mwoWFHaw3fgUji8lPR7Yrs/rfXOd2Vadlx
rBn/9c8Qco/8lp7gHhaEgok+qiH8bQSEq44M0Wru89IfjF2MLIJXXbGjOzX3elWA
ja6EaLYuBNSQ/3qnl6aW9KbldNa3/lYIsa5Cp2JfrO5xTUZZDA395iIgf8fsXj5N
47/csbnam/K6iYEntYDR8m+owpxUPwGwMHNSV0gNceA1IHzKah6ze2whqvxcRjd2
pLGB8cv78f1tWi1Br3M4ZOr+8LQ4MZ1Qz5VNE20jb4Sky3SIdD6pMpK+EYN1+HAk
I3dkr/Dhi8y3KoSzXTYmBXzL2Agxx1zJnabP2eQgAobuDMU8tAHputfPtw1fkhW3
3m9SnwQJeibPfcwTMIoTKbLbwmqjoYX4E7+AfUYpXZuk7WmEEoT+yZu280OvxGQM
9BJjZSLlKMynSnMRv9KgF7bHaVS2rrMq4EfXG4FCuZFWh19IztyhCfzILG3n4i//
N2Nyp/UMTOc8+7nxAb7jTrYDv0Y5uSnQu+6M22QD3V0jRaVB78ofBqKRvFdXlHFf
rZbvd3F1U8uW7RhxqYimYXnPUXF7VZ1x606L5mY9/P47zE9FfVU+NzGVLs6BBJWp
3xJmFIoUfWyqPMNwHhN7efTe0MPsMr6yoODokcj1pj9pQqFgIQ9E8iWY1ZxvuyCG
g8BQltiBncZRLDzpFrqU5t/bSvsFGgT6esfvt4OnByvheUCiF91JA88Pt9HuGxml
f9rd/rzeLnGzsL4FQesICbITTbNAyPN/Vd/dfIYL5Nz4u4UWeNkACH+d8UY3gbEf
a8HWGvQsztC/nzRrGlU9XoC+zq/11ODfGLEgKsOwGhGzVpZDG6MIFpvO41C6hpeX
vgG995kliSi/ywJfAylV/UB6NgF48IWPXfGd39+DEL8h1kGsHB7KsQJsROHkGEi0
l/fMSjd/LvvnqqVHzJ+jLwCqgAkcKiv94Uz9+tiYU5NJ72rmyPoEWU7eFbW0TL19
bZatKjEOHsEC4HQ3UiJseB1wv1GQytZ6cSiuxbxR+PRDXejNJn8cdxS0OM6wJq9+
jk2ybdAyswGYbpwLoAgswPQI5YSvfU3Vfwc/b1RF95zQtrhd9bWeZGmcmcw5MMT8
ef6m37QbM5X5UhS41Bhf2/AqzzgixYgE8wdYleiGJAKRBFybzLJcl6fA1B299/K1
Rsk1AvjTb1p1klm+VOFHDXFdsoJKncwHr+9PENJ6jFsMgLpX+FEhuzrv1JAMkIBK
8iODABKMyuq8dnfiypl3b7bUUOXGrgeEOIzBW8E3UT/0ami6zhUFvqTz5kOyCzy1
v6WDCBh75fs35SW7+pRWGRZI8U6IHCBiQPj66jgnrkID06c5ShlNTlF9SHsc3T+b
URm0e0/KOznk56RdmISXRxYja4DHdlo76G9T2ETYemweAxjZqWAnpXuSCRwYtEOq
w6OCKjU9bcs0QJPGjbPTOk4JKg8h1EHDhJ0SXD+alxWJcTz5Y3XKqjLBmqCFIIe8
QzqMGGVe0Jp7s99EGkVm+EMTY3BfowM+1tQMlv7ViCBMwinzvCc8pTz1BkK39cDw
nBMwVEITYfi9w4inj9yaUTTJMMyBvXbqEIlLnWyUA3cLY90r5XHuj0ZDGgerZ4UA
fL/9DQs2j/UOXL4Df5b5WomthpVFeGU3dphMxK3BcDOBAU0td3Na6hb9x4jWqLul
a5POxiMrImMMaTTCHTmxHHSanX9siVT79+oy6T7qpZdG/Q9AGFDaKetXf1mw6/Dr
ZHhd2HadJymI7ptSqIj0LK3pTdgafB2UYQl/ajlc2hTK0GnChvosqjIORoSQzRyA
viLJNvd/Gqpp9a8g4u8CgtKbM61TgchlnTyLvYk1PkxHcSIbmcarB1krFzqDOnpE
I1cA2J7mrSp+MofSGx3j3cy7aMD6BJqvlsG2lx8QiyH+riwrx4hLhbGnQzLbj+hR
Bp9qrJ+Brr6u5AdCgHyUq0IwIiklNoGbJMZFoAyXi2YOwXSIEME762yHXGPNIoMd
pjOQWR9yaw5zsQIQFiDF8mUrd6wUWzuS/2emTFwq0e2KTiR3jST/rcCG31w3vZfG
wWJPLMa7kygOOAm0Rth9v3TkWkcBbMF+LTjMFeQlGJeLtUOGnkdykkBmuFA1xm7x
DvY3ekDFJkyG/Z6dirlOBwHeo5P0/rh9VG0tYv4BR+5wHydyKlCsxQPid+c0FzX3
fWVkvcjVSkVOSIsbHQ6imnUSf/VTuq5ZljgwydoQ9xdYf1xJMpewOruFe/bptltn
l88N4tSHv/ypHhwcesqOhrp/dCyz4U2nVfy9QpAdk83vvtf9HRPtYxDTxcUBvOqL
QyUuOVsKODNJ4C1t57lo6pp5LGoCRiL1I5JeexVud8mv6cF9E8PvSgDsBzso6tOm
GqcuBd3KUYvAcoW4Lzv8cNFjHZSou2VMs0stNTxl8JLHYaF+7k9tyq95RMu2CZDO
uOoNXpr52WYEt4X988PwkzaPrc/mioBgiwwZCyss4838uKuBHAfsg2a8lmuz1Cea
1efHCr9Ni6d6bppQ6G/6FalM2gyYbjQXWNZLusEOVcKlDMPZEiRYqWaWuxhURXiF
dx0Rz/PSyTQAmS/D9NCt60dN8bdhkAmebVVRS7TSbQF3oTTYE0T9XTCUu+ku+mph
90jw5LhpOaIYhdPuS/R3VPvqHbRoeANB7pagCZeWzqlxMzRzjL8uww5pVexXOfUs
Fdbf8k6kvSMrgyJCQMHCK6e+nziuAt+Fr2Ei1HWjfhllPlLxOayB8gx/QDac70MK
RhSzPy2mGE/NNhPy/Fi6vwo90dj3JevEcz65S6yinJTIDrZLrKj4FO2MjqZTQieM
sAHqHWFt+LcnOhlaPTJdW/JL1WqR+Y14T97nATnOZRIEeirEPkfDs/5Lsypl1Z7t
uRxzGj2usvSCVx5Ig/DkQ2IdIW0k48SdZGVh9Rx4tU5NrFhIbpxQZ2XhGWR1/njE
xjPkoJG3TWaQXnv+DDcxqxSQCH4StngX3p9+f8c5x+NAq/XbyC7dBjvzRumSFsxu
up9HUsMDe8q/5RLsI+X1gaONZsyPGWccRcvOXivRpdZ0fZlDaBdEYP2pZnXP86S2
I4lETX/AxMikGkrPHlDNHotmOVEqnyl8NWEa9aVtUbTTfCPoz9+MiSK59NBPV3y/
tMOSwwrWhX3G5Z8R6E52IYvnCBlEjiWcxAYiJ33IQsGNZg/jnqOTS7BVr32i0pJe
zzGIzUBYSc4gtlgh6RHYD2ChFfF/CtCqDgL1hvfpoDOr7DbG9o28ZE3fgdGrPvH4
48b0clX6lwCtvxTEZRXKPVP2rtxZ0+Ko6i35tQvFlNABHwleadNQkW6esUPeF0oW
uapCxdLPVU3EQOUoEiYNFM6/6AMB2u1JNxcM+WqDnd4xhStyCj0fJVCm92fghb+J
KLhkCa0HsGisonSUzVQYsKK5biFRWRznCyvO/geq2nq35yw8iv+abcmVQGKsuazG
NGgbz3Zh+GyEoGl/fAxS0fLN/o9XSQl+zzFptrKgG8Ahr6LCfdFzzCeMsChB8g4T
aeuBnEvZTxb53/aYstxjZPqTd7T255GmH2BdGvotHgGG86JwREwcFbqOVZq3qSJh
oHuyd5M1hKAHlexBIadgr2v3dQPHSJypeVA5iL56dvmEbfFPLK+U5+YKrbYYmIDI
Id8agb0ZqyFifd/ZwJqKhJxQpWoxU7Q85+MkUvjj7hc6OqUDHEYQtXdG7XFh7tfn
sz6XWPtqsGwNxdEQnkRQtdmKLXKQphaiEozIPladkcSm6Y13AnSFQRKxgxRh28yN
54ah7j8J+3/B0bZwt6XTIpV6NevycWdwjtA2N67Pg5Hedk1EIwIKggWX4QIzQZ90
FJdCNM6z5qdCYn8pwmv5PuPnKOfdJh5XKvhTlTQ003+rzRTARegXrRzWl9AOqRHp
6X8b8f94XfDhsMi3a5v1YTb2oR62oHb/5J0K8Q+05iKfdJPPKjeA1UHiAKoZJTib
tzUvP1ruTtndgqpl8dlaUqOKUzMJ8kZEfNIQaQ2nAFoCTi2yLECtXkSn1Q1htZLl
tTVfU+H+6LiktKAyybe0VTHv9c4fHbOoDG6UxnsIdvZZDNgz8aEj//R7jaLofAoS
UOvydkC0YaMpnSIr4IpEMTzR6p/NWe3ez3y8TblpbV1OO2cyf3gpEfL8geASQqSa
7PlpX2VPjPMxKyBa+htb7jzodyeA9SEucl8xYnuiRh7txf6XCmPzIrtdSnxmQCnX
e8o+V6yY9sJkFlF/ri72SWTFi1MhAC4RrTHrWSAob20whtdmHzfMytt2abNHMCxs
hzzin6lFclUyQYOE+nfZmSXsJrM83ZIvZJ77pH/f3zed3/TIWfAS5V5lXccGEJRY
9TlvClH9R6f1TXoLm4CEMhnbzR1mMqizKL1oLiyicRVuATQe2h2h9dXQEx+W0FL9
n5LA/GR7Rp19Cu/F5XhHfLg2Ykf4/wpFa6HrqiRZbVD0rAEgkmFAH0mC1FUjxRi9
zXkudJVQWZQ39/BZT8D/mlpvU6jnQTdkrtmb/S2wpwLphMgE4IRsvjGwxmEQNIw8
wtcbtTymXjD6HVLK5Q1IByi92Qp7avaNxXvtU3KjfPs5w3uNFZ1I1/KymUzaTkmx
wSpuW3kFc9oxqxAp0EQmd2KVKamMpNH51ea6aDFEOnXQBjuFDrJc0hT9s+oLcsmK
1QPu3+Wkus+NBt3l559Fc4HcwsSLrCamQupuJVqJ2EQC71Kx+yrAdBC+UKrXt9r7
q+wJczJ0k7kqpjbSQsqZ/trVZGV3emOSGapcfo1l2GB1y9WqyX4s0W2QhNdQJLIx
ee5q4kFV6U9jOAp+RjOZ8irswMVKlTdpO10vIRRq+3XJNPD5EhfzmIM7u08Peg4/
EeX619NcWFcR2er1OQ2kXqZncSS9GQeRZBBH+Y8L4Ro8HZfffC9ad4NiUoxRmUry
cYM+GmueKgA8+RCHodXyLSfEPjVdGg6JYvkafR5zks2iGhaUevMQUaZCTqhQAS8N
NU0Uk9s5oicbvYFR+rUtgWYVXqzFMWy7/kosqK/HtKEuEcKNDh/N33oybVqtlcCL
/k7Bs4oPCNHfyOjvdzrUCXtaWzlNqdy/MjxHBDCabMsMQh5gChK2ildoEOF7GC9P
H35T/FtSXYkzhaeFYtt/gQNMJ23N++SI8qSu2HpiBashIwp0Rx0sBlMUrnoaLeW7
1u+Ls9NemhJbr6aUc9SCYN/OKZIqR5g3b7vmINbova8cw7L8xBd0EY2o96BGmeFz
Tzeyvzt2egva3I1RwIFbQ7KUBjkgCk1Lmd7mqugvZK4=
`protect END_PROTECTED
