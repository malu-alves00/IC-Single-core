`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
X/7JmpFpr/u9I4ZNvsbCLAjgo4FjdJEInA61LYMm6uDUXF1ynAYQmJ5BWsHQQimu
5PLqIs7qjelZ74TUNSdzLB1wvF0MWKAREq0rDvGiqDlZws6v9OVWHCuPWL8V+J/t
23T2fZZdyZPeKVvnBg7arIGHPA4wrbQZ0vdxHKV9sRCADKCYuymheICUsOFA/3kl
Uhfz6RPFmpJbmcBCWFR6H7sgFCFH6Q5zn2ENKyIsvWXwC3WkJZoTHtGnUDqcDy3m
ztB1kCmg7toJWKXeJt+uLiFNC0bYJ6p0+dT11P1RaRWQTR5xLNPucZ42TN1CoeOe
GuW4s5qjYukfFzukIFgtkCHCg1MRVpV2cgKZ7iLHQkfn8VA84rre8moktrXsjgb0
7G0S5p0yQodJcvxlmnh5wmrdYnChEyK8U11f6FfB+edjTzVjIl1VA8hLDIWmmz3w
Ca6wF+cHQCy8rcmjGHNQAdxmFW9PZJZgifILyOMRlyoNVKZ4i+dmM88v9NfnJuCF
`protect END_PROTECTED
