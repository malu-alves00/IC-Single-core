`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
b0zvMYpTW7d2sVN+gqJagj2V3Go8e9jW2Z/Mh7WdDzgLpo6O7DSIiTmouEjRYcvg
CFB1g3waCcpkh2qTi56dQimC6oHjjFx/RVX6Bv0peYqMj2/8DSp0yjec4e3iEnDt
kVVXxGUSDlseUztBy04xsavL5tjl4Wn0n+reGq1w9ggV+P0rMquvPxcJIPcsh1Lm
Ba4xuOdmIbxQWyBoUae/dqE0I/FTkKrJ4Wg66ODRzHH1yWPf1i4mUfGe7jWv6iAa
gFt93PF7hver+V1UqC5M5w8/jhe0u9dl33QiHMwU7FLzvKp090PRYi/sdfE3RZ99
738nBRizlwU4qZAW+x9Kdz6f33BzVxyHxch0xeLfWoIwXETuoXnk5PgGloya2iU2
m3+wzVkPxeAlC2o8tA8OGqDxgyHMNlqXXTabS/wAAiWfdB85dinRv/iP4opDikC2
Rcj+SNS824/0GMt6j7KEzFKqWkZd4E1N/JLUT+Zf215TStVbd0DRFDYkLZFVeVu5
wHha29O/8WLsY7KZTA09DA==
`protect END_PROTECTED
