`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hSDwUBN0DxGW8rXgi3QSj7ZKuhnNQt6q8Rft28PbLA+MZ4ibAZfOKcIY5+1maCkR
1LEgwaNjYlgoHCy6+IQohnmEXWLuEYPehYgM08zPdEXrTc4WnQ2ExjM8HX5SPHAt
F6SgLfenMIFuB1O+9heupTKr9RtTUGeLzJFOmfpNmEI0yonNqbMbjzziQRM1MX/y
6jbU4UmoH9TX2D/qqT7THb3ZFQj5/RBywMLcgkHJwUCpmnNj/V+HipfEyhe1lYOG
nrbqHxGhzIXzrgyuLbwmvSTPTGzsgn/JFMmr7LKxc+xa6UIj3ufafVm7wxqmNfiH
oU1KcYrWqppb6c+O+ArwSC/+YqNjse+KJL+zsxZywKVbRguIhAR0DaNZZOvK4YbO
q5g9DhvCFXJ844yc1u7iMEU9bKbkO6m6X5Ldw12B+yN7B3Bh03Dqcy6F7I6xU2xg
aoF+wXnMue8tDPOz4zhjY4guE69btZ7ko5MOL91CTR4aw1sASsWypQIkbaX0NT/p
HXvR54Ac9xLp6pTGk9H0taSAU9B5N/QgCt9RhjOsfy0aFkoM1SME5vn02zTN2SMu
CFHbmV6rhyM7e1AE2r7qU50E4eDbWnhHQbiSY4HNTyCiMtc0rLfzJu08nP6fUU9I
5ZOHDwqk7Q7x0TEXZJv9tVO1jlMsc+8/L8NPKGqycl+cdQDEdyUzhCU+ILrA8eQF
tLHFX34I6be3/YiDtx1j/8W4UeBRFdI+UXKBVV2DNBrhzK1EY7AoWUsQBoAf18+7
5jfX7AIeR9UbTNU0x1ThW6I+JJgihvna68gxpiIQceOY6E/+eWKSn1dUG9lVcj3J
5FLcOjSfA75yC3SIpzwxlN0jfUi+2kkDTBjsUDzrd6T+lByRl3pZk5FTrDQ2FSL6
cv1wm0IDd1OCPxQuX7QUMKyW4QBznho0wmUxYPi+1c8lBnOpv1b1hF4TMVfWlp4h
LYshMsUYDQw3UNhblVuytvXO7MYI1fu8v/n8bF8ipfqh9tkgo5b1DzfmpEvoKJLw
StjPVqa4btHAWLihtsmE5LNVi4gAwsnD9FUkwxwtf7+MnY8vGyfr2flO1Dteokbr
QO6nKbOQDlt77v286wfnAVkfDsfG4rC1G7M/eOIKyUSI0ZO4b5geSy6z9+zlCE2+
FD5OM5ikH7FNQawlyhVDqJdNG8CkLs+U0JEjWHzN2i2ZVFsJFyEEZY65aT+lneOs
zT5J8n6ZcmfNZFxBWwWMvtrXsYnza6d8Ub+t194+KBi3zikel0yLL+F8xKoWCznS
FknUM7l/sCc9EHfEQFrr6MtTj2GJi0Mx3Qu/iEUJDX/mRqdevruG1A/ODpvjBuDT
Lt0yjLavUqn+TqIEEUvCKM7Ab1HWAlrOcuAqXKNxrkFYsPgayT6ZbYKogO7dzrGt
HQKhGNHHgj37MZGd+wuTMQRZ8541S0BKlz1Jo+lB2r+FOYjY1kF2XpMVc5NZ8owW
B9H3Zh+WeEWY/hHPHdZwGQEUQugJd3bLB9NgxfLHGbWAF1PW8vTR6wA21rFfZQgH
4F2cwbIyj9ze/Mgkhj/QdYOOfqAdDJeQMx19+xQULpEXk9zbF6hMwM8v+2GThCc/
9/DRWqUYLlEXksbDsVka0TAeEB8rfeX46kwuSSQYtGrfUdjYmXXEup8f9f/PHjLw
0pjlsffyMIA77koYYoEIfkBOvS/DNiD92J+u/vfQXkJ2xfYq9MIAk9nozMMuJhfD
SeO+fDnpbDTlV1g0CgCRUQuS6AOwhrkGEzAlX/Sq7O6Yr3c1zsfRpBSIXu5g/rU0
Qssv/i7cvnfhr7yJvQ+HupyMiIG2JcGj27yeDtFWI5Xy1gp0TS0zap0YDveJBuOI
LpxrGA8n4MF8ie3N08T3ro0EAzC515xLnh09bY4Nde8Cy7c9/NBdluCBvJCcDL+d
j+C4ujbriHUPh/PZmuL8Q3Sa/okhbFKbeWabLMmLmsPBahZU/7YBm9vuV/5STMnE
t3DPa+3VSof4GsRX9t8Yh9x/mBoZHZFSunsrCcXwXj7SYbmzxzxc7DaRrVXiFwZ8
kJXSfdwltPzNTWqXDENqB1/FPbt8AkSohigSM4T3v9joiwXg2apbN2YfYcyG7ej/
k8OE4IXv2uHbTeNEbt01qFufIeli8BAqLB/cmEmvYKm+q3DwH/1YA+ko1gMIF55E
t6np7Ndr9AeVMn/oyA+Lm7IbE4MYhKrKzTWZuvNyfFhuoDZGZajcS7pyjSALZ6xe
4ZaV2w4kEALcP3vh1uY+pzADq4R4ObnFTqT1G9EJDEKiG5VcMGwmOHjmZ+UN4SFL
r83FqjtRrC7HhY4QwE05dZmRSdwYegTaZd0IRmxO1rp95dzRpDgYgiSuDBNrjhg/
4GoE+jDNfmJ4D4jemqJ58MBpygQtnRy9aDCEMcb9g+klViHZ/DWEgwvlpxp1fc55
mgsUPv1edn7Z5Ye3MFqMpGcnCzeAGnS99qOvIXz2OKioRlSKcNvIlr1l/ZA5rLBX
aLsamtq5Pwu0tTtgh38xELAKFwBKonVwTTZ42KcCSUuRAuBe4n3WJRv83lzG9gvZ
fuqd9+sxwJ04zijLqjDm8TOEoafNdraTXVMQwb77Q3QN4zBpGUsvDkanFEVdb9CK
u6F0Kk3TsSnt7riiBZcBQDr2i93tH7hJBpEtxyQgAC2KjX5HdNiiFyUZI1MaShNF
z4Z2hZYaYJguBwU+FyMTWTwbD9m7MxNHg6+NE9zYGHSxO/cZR/v+FYTVUxtfaAz8
tRHoEYE2UMHV4/3seYK5AAWUkiBt+1elQCDwfYwuM7p+a3lwaOve6p7B/pCbUcEj
SUSmfP8+CtVM9G+5J40E9tMozSAtmo5hCL07ojGXD6Kff/QQnylT3vjRYB6YiSnD
xgkMvbMfmNro51N6lIfzK4rpKmeRyBANk5GAznOZSlq0C9h3be+K2LVhya2YtXF3
K/WqgiPqC4kLsALrfIbUjWsqiOZ5fXETJhhBuHppxsXeplXaNaW2VWXHRzcSoThr
IyiSB9sVNWK2sL3xjvPF6Ag4r5Lwf7Brr8YQJjZzfWxNMJtJ+bDRnH6Z+gBizjct
6zrhAEnehc8k+NCRK22poXuQiVuhMS8Vzt21+FV1HnRg2dH2xL1cXsmMlWyuPGZY
I7eK4y4knHWEa0kBeYHwQaZu8h7Orc5ICOPNv7kRbHTWMyAGgVRHEQSI1pTDT6ri
05tNG9TFtU3M14gAockqUWQNRu6zLWSZvLc7+CfxMuT4AvD0xElKjpSC+LiapKT1
VfyPC0o+MLvu7YE2f1GJ6uPXl3upRy/1vxGeZBYerV3cYt/1FflCO1wD/UmmyWDt
l70c+8rruTRLCPb0cGbzapdapWw3Kt3VBCRQ0M3jsTlX5vVhPV9EW8Ce+TQYLmwy
2vqR1Aq+TNHnmCbhqRQsPR5dE5b440EBArwfL484ih7J5J1cISFNwl8AfOLqDKCa
qV/CZ3m5tLm6qesCMc3Oju3anpAXESuENTvJnWnWaglmlpxxxkXr5PR0opisGEDp
4fvoCxBrSZM/amfFiL696PwICPtVQRXvuXxrJ3V0BpK6cy44eUisd4a2KEUS70Wr
Fat8VePVFNReLVhLyGsoVpe2DuWHrNnrXqnvaNcgAGfcYZjijM2OkNd/4n7Mcgk7
nO/DmRs0ji3I/DwdW41xLdFcCiDLaR+FwES4WbxgyhH4Ils4lkbFOkyEI55EhpYi
ebr/M0fjhsGvm8YqQkPE31pbz3OwC+kzzx8t4XKjZG3TJRxDPews5N37s5JwVlIt
hcHtT8QGtEjNHZiPswqZEPfpzHu3ZzfWJj+NoGjsokVmsD4qsLetcICTl4jcEq0Z
CoajoXgzIpZaoGStPTErOWvr5sDAhosxEIJe5uoJd0NmX89E7CrgKCSIc+3uYjy+
LZORikN6/dl4bn1x9sFIvsoj5cy+8y1x/CPm+3vJS+uNrwfa246YaJBHxuOOFOCP
lbcQ6zKtjlAT50qqEQAXAPABT1gtRqqtfE1XCdinR634h4b7czFduCA8RpmZlnJz
qqRLil6Dxxli0gkBUGQunQKmprriVdNqYzrBSiu7L/Z/vtDzOHwsV2YHycJkuw++
2rk1/B8/fqmnC4x2iBW5ubBpZPXo4K7LbW5OmYLJLErX6+Pc9Jpy3v+ejeypqsk6
dZfTnn/LRhcT6eTnaBeIgefO/x2AmmD3ciIoTP8OKN8pLQUFZfXSDEa/auWkC9Qi
PhLAcpUVJMgdUzYQR9rAC9VwVhsNtRM1XcDv9/i76q3dLtVr26V9giXul2MWUyKu
mpYgOWkx8JwMPwO8fzYbR1TwiBRv8YXzkM/EnWj2a19F1rfcnoGZTUEesCFh8TOt
NafpetmFp+ARWST+nPPFAeH3ww9MTEOYXPlns3Szdn9qFghq5oFWHVLtFYTUYZj2
OJSToAxIVVbREsgsMmCnkSyOmhV+QYInpqF2yeKleck7s/4Tnc42M2nDIkDXHnhC
/HFDEzjlPchUEICLob35cdg6+eVE2xawfos2AyyKEscXes4CC708xOcjzBEdLx/v
hVXPpxwIWqsB40QEhzEo3WCNgmrDTJCzu2hJG95Itwbho/bfVKBMTRItMVMkQipv
l5QSVJA5oXsj0YjvfBzy/gnWrfw/xepywJFA4ECU+VvVJYHHsSL0NokwFwZrr0cU
hrkkmLG8Nhv0fCkkoBrQ17GyrHOQ0muzjsS58R2Z2wrQQwToSe1cYC5yfOmhBX09
qJWWVkSRd3YK99WkwLcSLmmIzKwQCJnBSwJj5h8EJFNBshkBHzJn6ggNvVHiM4X1
odDS7aqaJncGEWE8xV3fhj1b0Ss6ms6qnRYsCFXBBWmCGmB4x4Ab6ZCuXIQ9T0Yc
ZDTHj4AAgyU10Oguw95eutg1Elw2RiaQRZOPZ/uuQUh5RhbFV4Tiq9/hqwY1OeQ+
pKUOPEfbWfjR7B0OmmAG8PpPirKR8PmgdSkKiY//E41G5ng8ZTRvg1AfF1C90dZu
YKzvZtPd37LimIcHWMCz2EZAj+XvoTSF04jvJAxkKWWbu39rdRZALQaCdJzAaadv
rMZkbY1paPDrYVhJJM1M/BYDghSI2t7iIsLQqlBhC6z3w/yNbL6kQ592iFe/YhAT
X1AV2OpHmNxmbFasyB/+cItiS3o3S1U1Pq4cr3AIU1O+WWFfMr2r+XvW+iguMF3I
WbfCvHeF3LtUiqLY04MXu+EJ+AQDEIIB0TKVH+zA7tv98sQxge65CkUtHoZIGn8i
NETawxOZT3oZ/VGP/iXn82CkNpJd+wwH79sjs4NIxzX6gJU9c7wWv+6yF3RM969S
Xe017J/+7pAOsRsCwDpuzDFurYGLt0nR+yp+rFmkMgyUxqfElr7E3Wpaf/w9zsiO
Oe3eaovHk2hFb8/gt6M0Z4IwepjaCaSafg4Vpw5ineREQI6XZ6flJ4TjpXkfduSl
tyXx+PnWZU6UuW5FAeHxjqs2aV1UuMpSbnLJHrI0RlJooydMCBuwuf+06CIpT1c9
QBlWLrWbBSBKlK29WdUXgSJ8IJ/fYBurU+tbyMjbLpb5QXZXzVswfvL0YODMRECX
sMqpv5LRGsaYxmdjp82XzS5ZY7Rm70JueZnJEkirME6tF3KmfkozUQ4D+vgJq5eI
vR1hr4Vb4GJH8Wh+2IE65Rd0UTWIHK+gXq1b5lI0JCvwu2SJ9ViCIZJLAA2HBAOD
P71iRU38aL6o64C/WWafz+35v5xe8gkmXjRMnY08CDQxDj4IEHtrm6mfXN3NTQod
ZzwZg659j9UrIr/fgTKEV4MIkyy3+rgqHuQ2B1gJbyEqXz0eZqvQiNreISnTdeKb
OSHnIAyU4c9qEaptp2g4UuO+1bIzyzkiDAp24Cr0afrtDM/7wIN+YCBJLT/9cKtv
WCwh8GZvWrDBPPbq00fPCuGC6Lu6pHxds0zlMM2StcBA1pNm3msnetlErXiZcdqM
LTXaeh9vTm5X1SMoLBhyNnE4+EqCFyaLjFyP18mG7UGHB6wXf9p2xy9xXeIDvvrX
P6NuRciAmKDmdGkh4mlcQ47oN+YHgb0JRp36eIzzg0WGC+uktpt3APqdOOaN+OQ6
0YQ8pwzZCq3qSdp2LzEFpTsmXd0njFi0xAuX+pA2WsmyQ7lILYzbp5mjZ8FUllM3
2dCDXzr1YCs56IgSfcHPSzyA5T9NM2x7bvQhYP8jH9Z5HUl5NTFlFI0KA2/6r9SK
+n/ycSV4FShdiEBVLSR8yjQYV/fO8wR0yzfGO2mGAu4m6zqJKoHp8Rfwl1BCP08R
V9Ldn8xCZ7ME7DBY3EH2ff685MYGFVz76xwtYQzlAQQXCxmBvy4q6m7nC0X8qiyL
0EptHsMR8VGHfUPOc1AV4cG1J3YxYzMO9HtH7WqA/SacWj4XCB2C79PJW5V0DLVW
dXUBzE2UM/mMW2XxDoJN238s2vIPcgPQlkMETiN/4+Wv06mC1Wvau5g1Xo0YxacZ
Vqb3J6Asvor6e/0elUpZQwm9buJnnNu4AkRqVz0jxtspF8nHjpSNvP8cjynBEX7o
oQgB7kpDOExD6LwnKhmDST1GVmStDy1DNGKoSfzoQXhNGL2MGL797ZgxGa4J9J+p
jd94aqYe8Tt75fg8kvnW1m7mJ1yDz2qlrmwibr/C1xhMpI3f4a5mCtGvhJfYJjs3
/5yq1M9mIAWU0DFyoIWEkqxYdvlCHRzyykubC09CPvt1zf4lWDMujUvsI6jEnf2d
d9dBHx0vnqr5AF9491rs7SfhDO/8znKs/CZMjILjVgEMxqZMnbaceAJv+3SDEHCq
34VTE+kKsJP5kGgaHPK+lzEKXyFhyDKO3izMM5rkM5VZttS+Xf8OoxcRCc/GkJVe
Y3NIhZznV/zxDRMJLK6WKL40skbrk10gZXIMJeez81E1b5DSG4eAEJJ7E/zFTkU0
UHuTuWj0tx6g84/6cj8jcf/V2qbiYthxm6YJsNE49Z8itZZhRbYiZXPERs1R09hi
h+XhX3WwExx9RnDqtPdTb8DXhTrdQW/MIXcYgtO2c84+BFcnpZyn9DVdHJuapVgd
jpZyxqp4gjY8KdTRwf27FHUaQUac3mHUuhF+ddpKdsFr68iq46y85O9TGQ0LKWI6
nFK8/9N7LeQk6rAtPExW/Of0shJ7+3dkXKeLbjaQdfPm6DDol1j3XdjE3fzlI/is
IZW+y/s39joSn4JkudpRRYAn0uXsQIKM9ghRNTZXRR3UYaO32lvc491U3JB2nxYb
qQmK3jsdRHpkDwz8AhZ9Hr8A2/kl4Z+onYxcF9XuSH80MR4y5jmPw/v9hKPgGUyl
7tqOre1bh9aV9a40cKF5WsuseVYQXXeDVAqVWL2oes7NG8i1G+jvSNfefzicgsvZ
bj9AzARJpBkO1oFFdFzXkipvK2smADeOy3pPivIAylv/M8IU1LvbMnXbKy1wD0FM
6wJ32GDqIzH6Q9d7YjhLxZVyfI4ST9IdmULtRyWYmrukufwzlaZORnH1NFG8L+nI
rPN7jxmYj0MR2C+IsnbVd58s+idHxX/AVAWoCUrQxVOEw/Sn4aU+PjfTAMumgF/t
HQpDbCVyHDh1ewSI0uQTg51ca5AEI2jOPRxQBces9HJzbNja2UNKbYRd3fbbviP6
J0mmZYEjJizaGZrT697ew1ydJXJZJqMMdW2yjQUx89TaMqUMBy5J3VfjyXqC+e3/
d5Sw1f/jAXrarC1I/jrZr3ryyJzYhzYwmdSrVOjBlwLqaQTCScblZidLHTMNZvC4
9wgYQx8UKLic6N6K1GtDNl8RRglLTPebibEFtUVrWmj0heA2w2aUC6po02uNaRir
rSNmOMdl4R4QnIlmq5bNvkUzpvgJj64JD31Zeq+ghJv9kAIk2TqB3NRAhOfX5Xal
SQsKZYkKgPtmYe9NjiJvXfKzAgqbqPp5uMJF9D6SptFAgHNK+T6rmEKKsNuNZkUb
nLfZM1+LGURzKjO4+CPrAmajBN6gX+Sddg+ecEZpqsOhRujTkYlqyz0+synLfF1Y
la6R+J5kx1xq90tlTGMaMig7zAwS9B6NMN8updEzPEAoxGuOCkzksEy4+Vj4N3UP
58IUzPK4GcoL3k1Q4r4Ht/M1iNXGUgr00ziMLawToMk6qq21Yno1eM2SMAJYr0Lv
R12TFqkrny/S/vWOiVtm/AsBMh4YiyPJdMWa8mAYHO0/5wSCyOzErE31ANW9iRLy
BRmEO2HLLGS7Y1/fId5Wl1OvN9ft1wHU5FkOlUgBpte58YEz1LMnkhs69yfMe4Eo
zegIPK99ShGqDR1vDCgaZYo+7ucGHumJP71dNZeWAaHdpETIb+S4Y0lpDl7/xvV7
2qqfNMVVV+bpDLBHpVCjA/CDrUcjEz/4jn/ARvC7M7U/klI79HIcskGNam7u2I3U
DLodps3VZeCzJoBGD1QZ1S8DSPuYHnKxl+XNN+igH43RFFRE7fh4mf99ORFRRewT
KSfyYsVoA5af2v9lHIPYPa5tuaYPTjoJ/lxVPX3wsxN0ar4HPGxcvAo6ijZeSLov
xd8hKVr2uWyeaggK4rtCcAkRonYarDrWWtA3cgZP0pSQnd04OB8B7yzgBTVhcZpJ
fVnt0DHdyV8NUpXj261xy+14slgc9SPzoRNrvgpM5qfOCWFI4Su5pw81/E2oY+NR
YfxRHX3jIZV/G9zhY6n9AC3OqvJk270EKbBFoqg7PwOUBmj/3oQ0uVoAQJBfT749
OWC0/unsPc3uutzWeK9xeT03JfFbHB+FqEk5McfzYY0RKi53EHrfSNbhUvMNKfKW
EL0P7JryOgZ7FlBsXoP1N23rfLk5tHCkTVmK3AA7u8FSiGLl417/6X9LeabtKMuZ
mPfySPQqNg68RU3LK11+/BSyGsS6fvS8O7un4AIzhGvhQGNswv84ZkR3HpYjvg9o
Z87MwlKd69TuT6HlAzvtlFtPoRReQi1tXnryFlJo7+SLcfm5WTqNCEatDsEt5brM
8ZIGxd77peykS0ouJOsr8DDR3OxileDSqi0YgWCnx/6xZ2DbX8HTB8uvAvzG+uUC
MTQVh001kIrNBwI89q6bs9hzl6YbYGMb3acPs4gaSwbwHOcmIEZoblqMgCsb4ewV
xR/RAqHs3H2WT9kXLuJDpiYhzdLJ2WPrveuKhbFbjWTY4NL6TKpNRNpHZ6HStHN5
C038YS7gsUBISx7sMofgFnbI2CPmOGriViNG4hF6Ao0YMlGH+1qe0ZYW0d/Xh1wO
mRT8c50EP1bsNQF68QAQ+LVWfOQAW+23EuAAOV4khWJReY4BSRyE4rWektZf8lWw
JahoCjVWqPQR+OBOZITbKNEikYhegXX6+Ua8Z3mNxMawThK9274PUWIWmxfrFRUe
cGV6Y8BHOhxaaZ3g4oP8T2a4WU4jrlfmaODCkzZUrGyrBNA6D0vm886chbxTUpMA
6BYoMSY4Q2IEj0wLFj2kV9lb0yBGewDio5C3Hv/sHoXtSKmbSxsfo/9+gefQD4h/
AM9aFQ6Qs7/uKMEMnHh8ZQPmSZZA1dTbcoXBeSN31J47dN7siIKI3b5ALshrd564
wAel6nFVaATvhTjx5EuxiyA82Y0xveIhlYCyqGc5GFnZoOvHriQ3uOKjV+M2zxj+
2NBqLQJer3mtEy6fwHPKfGFqnX18WMFq4lcwpFuKlCf0+KRrEVE+VUyQSsGz++KR
mEFWf2Rd1IEFqKtP6mNP07O14Pcu9br9KeRysjXFGEvk9QCBnWnhwFEUx8zRoWTT
txL/D6dD7Y5wXZSKkUMFYWGmbUKsHcJnpEmGLmIeC7UqUtClHAB5OgAlCx9bZXSg
/fRhTYE5iT1bXi4vS5UMuuQUWtTujK/2yxaOO4cWh5NSU3HdaglKnxv31qqydtKn
bGlrW0jfn4CfA+2azfGCCjiqS8P3GYZQGVH4GclartJk4LjcnONEY2XuSK7+SMpy
5X3Ruis5yncr1s8tvqoUUdKkEAhqq74EBbTiGM0QJSmV6Tc0tdJUjyPqldvVJWUJ
+LJug4pCbjGgxoKmuHq/uey1lKB4XDk3GPTOcw24Xa0ssGdwReAB/VwovZpuZFGe
lUPiG5bAZlBPYiAovL4zxsuXaZQ7XBFlZi6MzLUUcQesO+rZyFhO6DB2IWJL3sLC
MBe8EglBR6Vfy8uGMSkTOlNPbKi2LJvhranzdWYZypZXJcFdcqnFZUralhzwOj9t
dkw/R4eC4aB96sZW4+pLl2/ge5Q8lvMGuuAFYcmWGziGcI0kaxNj+t2kHi8C8MgU
kn7OTLywaBOunbQVizHUhoXRNWoNMRwUQacz48eKlYwUcsnVJsHN3pzsHQKAWJTX
MRC2Xm8cJglOHE8GpuCOJtT2j+h0cg1oLFcMFrRvWrfUi08Y3lUq8xSTg1Pt/0qa
oIkJXrQQtFL7GQBxIPYRu+uQz5YhcmQlS2H78pQWZeMdP+kdA8+2vit6NwX3nXR0
QBJ3CzMOD3h1Ll2Efef6PYPUrdw2K18k6FQxtqVzDi+a35SBsq+sQ7LgnJT0MM5Y
cykHEG46OCPT92paigfI9rG03J0TpVGfi4OMkBOjIJlNDzEC3SqtS+6Aho1o3DVI
mX57XQavbf2OiRw8lg7vYEB8vz393NRjGb/hDkRURbJiF5kUU5B8zBgcuIepDWXx
HNW2sMo8WwEuGB6qIzv3nDuO8oNSsmmbiyqd4EJzZ0JhyStCVuzH3oXVi/m0/5Wx
xL7HbcSQVcyeEiraBFOIxzu727z3QAKH6B7X/usqMW/7wP9TC4LQ0rhmnWIBrG8t
LTj+Tc1+aB1L/2uD/5tk1pKDjyad9W5jnpy9cgdkuwyuSg/m7Hj+3jj4SghAcWZu
eg5Oy4yU8NkGWNH8fN/7rkSU6TMTeAzQ2hXjmioaa3mk9Cv6arPd0fYI/LRAIF8Q
UYsBx0zZPd/fXvuFPwuEWsM/To8Cjzn6433U2J7Ed3bCxmPO+G3W4DqhqcpEv4Ey
yIgCytwizIVgPMlLH4jnpLwOueGg+bTRun6yfMOQRwGQ/ygIqtzUOau5TUlWRWDS
b6082SRJ1y8OYYLncwpvW7ZgF+YQkVbCInGPRolXEDae9n6oAQsb6zEnZvVMzhXn
ySNmnGH9DW7lYjKKuErSGx2nszRfdLjPIjBYKFDZguEZIGjW9t0PgYUW2hWdBEpv
H6uRyW3eevYLE8mJ1UVwvFTGFZ0S+vpraAEwvlJfVPwrydanxh6WgTtKJ2SbPlG3
MbrgcsmAYtgdJmcIkMUKAf/wNz9DdkgcpdjsdQeP8K2dM91rIRaxDzwa/dYQf07E
kfsxJPYBiREWnz4mQU+Wr4+oAvo3dYOxcKvOdeQFvu/5/87Qq6CFxC8KH32aLdY2
h51s2tnhrm2wr417G1VaIza+auQJytkHpf1tXm6WtTD++3mkW/Izk5i6Pxwk96l/
5s9isL/c0ENIZjhd0yz0j+7No4D/n2YDcB7CyzFpx5RZonS6EGHeoOOofJH0+x5B
Wk859ohwptdDpsgBjGQPfGD++NtYD50/PnLRAi72cEn+TT2qjwD4jg3sk/xQl+/b
RLo9//xTUCG4AsuN8nCwAbteMUObzEM43IIfX0HxEeuRz7X50s5KNmmJksBJap7y
8vazcJGjiuIAtc1piwudIGRrvwvbY2KRCiOntsRsuYmy45130CSthK5Eo0uNgrxb
DbajMp2U1M8rhMLRoKN1B5wDNBmkr6P+w/ORXeqEhopuRSZSf9A5zeNlMTS7y7Ry
OLkQQpFKnEz8kU9HjBJjokBDnTXPCClCfMPe8WCpFNO7UZ6LWyWtQHWqFRgOiZuw
PFpVUpX9G929CE3VtH9RE86DFpa8+KgnMN7mZuM71vY4/mA6OwIf70+EXspr0Rdl
mZpSkMJVCMnMBpFMMzQJO0qd71pEihnk2uvVZe9YgT9Nc5EKjnkI3txC5mUL4XF5
+p85VMAM8t4X4Ve0nPSbEysnKZkw5sljWZ6LbQs1q+P8/5OUJbZe72YADEVG9GA8
C1iFjWdbcqQqc5xREVcYIgihcvtW8lCLtKOix73yaXIJDDr3FOcBoIuICOUo6Nlb
3XMdLtqLxjbQwbfYqKfFpYa5859AblmtHff7Xj9ZYRXhBHTAWDTC9uvfOurRMFi9
Lyzp7wISd1hiuDLG1oxDHK7xWPpq5WFCJzZdCXFw7RNR9BYl9dugT9sZiZFj0wdB
M5pU31TvQWXmYxqvYOjacsumMpvFtRervU/5gQBj3Y0F0pu0avH9MK4gqfPJdwd3
mLPe2k1gSiF+JH5mhpIK3daDp9r6LTBHYpdu7gj5ZI1M+NFhyn6s/Yja3ggBy4rt
lzdSxjX38vAF/Hzj15Dl8jZESDOKlc9BK6Q/R6q1F2CvzADhS2n2y4R+E8fQNATs
jJuJwKerG2IP9wZOAkmOjMOqyU1WR3e/hQtI+tg2/rzwmcu5ybABE1nCo+xeIw8+
c9yoUs/XDZQkEbO9NyPqesswc11dhsJTnJWGpHMOWEMlplV6itX72CeKNltJUFku
OV+oVxuzbHoODti28k3gjBr+XaeqKvJoMXeFeLI/d9i1wGpKVl29a9n7WIazkI6w
e3scGte9I9EeMFfzh7GXdElCWZUlqTLb96bqS0cNH/w7r/6GUX1UrxUMP8ihxfXK
3LlOHQU2Tt2vPROeuehmZigJLf4+c7blETZtrFEc2uGTRcQXlFlI24dLr7wV6jnH
hq8R/snj4joY+g5WF1rnuMqSme+cnGVPQEQRS4fcSNsqKeMYqIWeJ1lc2yTgSJpJ
GdwJyu+4RUUaHHseXvDV7DE1VG22tW0fEkztqK30g6tSBLAGp6v+vNemgQYtAlbs
Bu/iA8RBVzPyQAurD9gd6yeexEDzph2JPsTjNbBNTsYsEamkkzolDOnOT1ahZukr
b58D3hl2TpjHmOyJ9ZQGYuyivt8W4PAg+rpff8/eb6Bq5xJQ9uiTMBJ73ITg2pn+
3leH7j9DWjZfuXFHqIKYWEVK7ffhAFuhhUQBzaLgOH70jsBJV119DQCStGxKktud
dOpo2RTTuvBz85jOMH7uUcAnTlB7XXhrc2rKlX/DumOeVAuirdIOo4OlQlvESgmi
TL9MaLq8av0IpFuaS7qZBpAKn3u6oBJQK6PYYw1SxeCtcC/H1kIN9f6Zk6WYx7cZ
6heIeuSOjr7V6us7aupD1N1IZhMvFZRWh43BgOy1r7jaK4ZKGA5jyMg+w/wgYskQ
5kd/0GZHoEtlKNaD2MWtypTx7nhh6RvaHCIHQwvp1cfZsT03r8pZutB3wJWE7R3I
L6lvzJ3HZDGMlHMYAvu+Gq1StSlw8j9FHf/sBWGAsEXK+llHxIjNhaTk+3IlbzVX
fpej1Qexx3VW6Yi3u+riW/ixn0O/38U1152fF+2aP8wgILUiyy+LgZUTbKOv/lHx
ZsJfP2Afz3N3MixJ4iSR9LkaeszvhmrcYIR3xCVvlUPazvlgqjH3lgyJCvWntr2A
kS5bJvM/EDw4/c26JVb4LQBJHFbtufkniYMp0a9pHw3Q/ypteVEEZDIg1JDRHNk2
3/Tkiw3n2/eoBniSrFbLffoj9JweWEK5EY8xf/20LZ9UTO1AUctm9XmPjxv9aRJT
ZvBK8lwcXPTdPk5qLgJf9GvwC54okARp1+3RE7dYONDW7FDucZerHpyUdjYZQCHu
T2MycDDXvSj5gjwuEGhWccWsP3gMTyKOjHKhyEhj+qXbhvvUaW0KGPY6RhVmp+0z
gQZRPwhXn+NbJooPOC1gsAHo3VCMOEi+x0DbCMbDAoDmrJLalTzMjYe2/oXHPYK1
+nYjuOCHH41FzEJgzLHUDLXKRiArBe4bDbVZffqK2X1LS34t0WFdba6P2cb/L7L9
p5vtAa90qinGYFbLRo4hR0hhOCCc8Nc7CWacAlgkoXolOyh5zAKBNWX4thxfpF5b
PIq4qJlzrFsefVxcyGfICzepCQvILSWeN2A51Yt8OR+0PCoEXZRHAWR6/qX7fPeU
23ih6KXo+osTO2nW+aAOVjaIzWWn8JVmSTHLFWvdUT6NQYW4V6NUkZOyVNNFfnbM
RSIr1nmdDf+RTtwn1xsKzyg7HGt5Vs3sYB1X3HnBF+RKrWIBvo3CfC6btUBwbpsR
4kLLlak8h9hmdn23DALD/BjuBxXFjr24UhHCqXedNbOXPT5EPml3HGMEsmzpx2H2
Bjgce2aSOksKRsTSdqil5jGT+4rooKKKSNwC4fqMIKFKymeWDi2eDvrLFQ6ZlCbJ
gWDnvu4u3O6n/U2SAKOTpDo8syTFV6rPGNe5FQghd29Ma5ejrEtxO2odZssv8rD2
G9PBUqmzpZjR+MjfGn5jJliq5Tv80XNAU4cbZcEZzQ/Dt1ThOz29u92zd+h3V9Ma
xLQthQxMQpQHYxQhRQfUFGHa+wwRrt40PvALvIuT8Ug00K2wV3TFYEiiQQcv1LeO
0jnQs3M1P0/lV7Nq6HJvb4Mfk8WnBgWb0RGh/T8gkJkzELxUWj+CplEEJ7eW+zpU
WbAI/oEn0IrNK1eeDeKKbuM1zUOnkN7nffPjboZ5MCMDn+9M7EBIkNoOi/X9Fveq
gKZBR6hspVcGjx6b3NsA49Ql1N1RDIaE1uy6DXoKyfr0di5ecpPPIceSWobFARPl
h9bfIVH62UZzTZf9LNe6abWTsZfr5+IQm79Wg0jW0vV9fqicfMYQTVWxSOK35vqm
eM9NowDMpZEu6V6ICO0n6Lv4X6h8NS7IkCMY9dYfmV7gqoJrxDyZ2KTkTiUyUFRv
OkLrWhFragESHZPsheZrK1R9ndnRwpYKCFSePMAl5mpmdtLSOiejJJfXsUeaiWpk
4WdyYY/pRYZDgg6Zxjx5v4uU229ih5D6N10sUcHq27VayXtM0N5EElCgebjVo0J2
8g2k1Udyj4ypxpEmM5tsh0EEq4jOx2YZeciqTrdSXx9OHZNtH8LU7F2jJgCBQ+3g
9fp1tuwbYqcMrtWpCT23pOIm/yMC/4p9VG3ngskFc2SCyhDlPWd3wdC4C6d7iire
GnrIsAM/JXFBbFeg8Ty6L8DKfEo3K7pGHG+pWyReonx2zY8AW0xEBQ6qfYP/afsn
UOidP7B3nNVoo2f0o1mQR5SIoUv9JBYFSej9QmmTvVWkZzBMqzwpZRjS4zGtXTn/
bnI4gv7tsWNidZa54PBdMZXjckZZXFckwOU6FhyL3RpopdhVEgFojbGP74JiVGTT
p6jFT1ADH5KDweMVW6Z1jUTsWLjq0ZwKBkSW9qBw9ayHXGEzM4xbkhYGYFPVRjxM
Gacfyc6VYv4hfYfljINvLOf74OzerZM+mokn1wznxPgiQQFuo90P52N540Pd177m
qecyIC2jsPbe0uhfL3DO0DVt1jvTBOcZvfc8gNp1TOUuK+4RdCek1Tg3QSeMQCtD
8s9JkZvmqd5Mou5VEj2y0NzVHTjz5Ilmqi7Z5Fl7lIu9crgcDXlPniOPTiNARc3U
ZuaVK0pzmNDlKqRRqtIEOkN2RXQvCL39xf/bOXNTfPr2TmRFIMWQMezGoSHguC3S
hFdWfL6wqyBZz0kvGtBy6YYA8hlZoPrVB3MRktiyrAP8LWdGZwTGJT4yyA+lyVkS
kQn2y41IxeyurmLIl47T5lQ8Tz7Dj1zprYZvv4SjBVsrLbINn13aXFVJyQEwTc/5
jr0GID3OfAJHAoe4IpW9NdzJNlkzZ4iKULQ7/3rWhgRldybioLHMtzo51ugA+Dgh
6k5D0M9OA9NVIOIwUpRsDCJfwnjO/cBn/dPmYeBsKT1TPfgdhL1yWyHkN6nq7g1o
I+r7aGDtZds+FJRAJErU02W29XnKqG5VKehsdfQOlFE3spMtvOXasmp0tdF3DICq
c5XaiqdzJf1Kd3ZYOCHmW+qwq6oQixKGRMbPhs8qKmc2fFBy2kNRTXT9+SpIt/s7
8Mj8/9JuSYiEG/iDkps2xkUKdtfHkfpUk5ANoQyxy4qFq9bDcFVl+oWGwFUT95Y6
QDtk1/W+Y17YEKVc+zQRwMKcCiz56tPXVS9jgNGd8leESSnA7QNcxdiIwWERt8LL
8b9EkfosMqqw+tjReXFNjUyrZA6c2CvIMya0GPrMRSd5TTOwx+jiMS9DBMEB24/l
hJ7y+ghU+Lfzsb+IEjILq1LWNojbJtglPi7xEEnrcJrjJHf4e1FkHN9IhVxb/vZO
q3SDwUbhwIQ6O9Vk3+bbWw9eUqJFaxSDuyX3fgv6zGCPXvGWp3b6xm06WC1UjKzs
bGBYJQGmNsmwldFltSzruPUliDR9TqtZS/cVpyS9xcMXqnFvAt7ycpY1xD11QpbN
FS5MjRKAmwzzLrH/2jtgm0YU1Ggm3HYi7XnptKysnGdsXv9IuD1T+K1K3s2TOt9n
M7dc91f4D4c9PzipWAW23Lv+xUVSjR5YhXVcW5/ey+dHX3B9wrFnjE3Hv3aBtFQ1
cJBcuClXuU+rkSRdF3MjRIuR5f/eK1w1ETKLFNkeRoU3fEB5BjY6UPXh062oSyUu
SClmWT0TeAnRdklqJIPVfAC8ljnmXYxccZhOI3iwL5lBqaFSDkqBhVrAGW1sNp3x
sSnE9upiXFmWin7txIf+3OqUfBT8KnM4MzDcm/26yES+b1rMWN1s/A4a6vgwfXSt
iT8Kg1VyVC37t0WtBKjXRzt90IxtGrwJWHLRo8gzwxq11F4CPFu5+Xw7SnC1gIgA
D5uN8+eRz+TckUI+9HJEO5uwOSMsA8tFxumwj+LWwg0cP8NtGt1CLKYHbRJtY2kz
O14vJOBIx2SUbdXATnWOhgSmdSUvDUdJKfcx0p+FPkiUGhXXQjDiLcww42H3kcIJ
yFcmTcoCu3V139/iJD0p/c9jbIaS97WXCZLmHCou2PBdldaN6kaGWjCBs5f7Cc7K
mlrYQp9/Rih+yVFDIy+IfgyMGDYg4t87f3cIFXQpJqwkOTJsCLXiuazpgOyj48C4
eNKuFhgFu+6a8djRFYkCojWDxVbY4mBxEuGH3hBIUjc7/Ib3tKZYDnoOYjlGfsW5
7zxbFCry8fFWaSNzLrMk47wCtcGSmfv7iS24JRvTBZ51sE2f97sSfPK8D9KepI3J
zcPs7SeFJfEv8IZaBeBZDV7kOgtj4UF0lVJ5fbkW/IoJP+pNyHgB05Hoo+O0rZbD
FE2/0T3eTr9p5ZBFG2xqNxbDRJcoSWBeNwikZOlcZaLOtZrrz1ar51CHaMlRkBNc
foDRT6bPvUzGyZeu6Wq4lyV0RBaybc4Qgt3cPcXf8Ti3wn8zwfeGTd1BH9dGMiBw
UqdYnYp5PF49gPVA3Hk4B6MwwUXOoJo2TR3ozn43FT1H1nx4LqNmHf4++GWetBzJ
Dh8PvcdlxHusdCXIychWU7CpbPKT2b3+2KPGnI1K0N+LASOW8lSnSRFX/Bg/4+u4
UT4XPYuQxEZQ+cIf0t6lc/CiNmyvhLWrIDOiVSW1HNfYZ5Rar5zRT3GevM+OSOEK
NDQP/xbQegKQDzZpU0Bq2apVfb+IT+5ZZL6zQaQS7OE0WUnrEvS9InjoccH4Asym
tC9Fym+oDNYQ/hclxuP42br3YvgcwGVOM+/IwSPFrgVvUV0fN+tzo2/4lfwgAM7m
Za9CY2LO53Y8vYpv2jorAGanLEWCabv49x2VdNuR+/wDoHgq+3pS//r347afGkYm
9EQfUmxYrLh+GzCMvXVOzE24I1gnguXqqAgRriRCLn6DsOtOKqq2T0pVsVV6qqD/
drvJqbtwYdkmacpTaIpFie7e2UZYuyj6kPjOKOPk06yGlY3yyaopkiUVA7jU7+Sj
63K0iHF0VYSKfwrHUiUF/XoPF1c9O1hSJMAmL3+n7W9fdxDV4BpQehKvbqBRXrgC
xcAVICyCZErGG8buCDasRBA8W4oYwVfD1XjIw6SuzOHkQ1niOGOGUrwLnvuuY8r8
eZ1mIFYmR22YZ8Z0xTLWtO5ShDuOt8pCrPm31TTJ1Cdl6VctE4psn4zMdy8wFmnA
Yq09wv9XxdHSMkyhnVdNQdmEfuWURdJpYOUU+UPCXAgLWvC3z0eqTXFEP+KA79cp
vt5mqPSvyA93vLSKL8T6VPu/o+eEVf5WvG6jOjH7SCcZPpRzidWrRuvF0/3jf1gy
UVIpvTs+B0mFPif5prP+4LUI0NwAujkNWipVifZU+C4zwj+dmX1e7q/182lhp8bX
5cXB8EKuCwvchVoK/cTR2ldwYIuZQKaaVHMmqQ7V1sUcBTlK8fIjMy7r4nk17pc/
NGMNVlCIahJwlYyCSmsiT1hzTi+9WSOXNh5+wbhuyXlLFJS+7KUpWcfH0ddcPWLK
L8vgIeDL66A4b6v24hjRsNcKQI5EIxVXkrX3VgcpWRjsUOf3FD7T1qdPEdt55hRP
/w16giQEm8C2dYFjxOlvZmJz5yId9yS53oajtHIcJBwCmGzCmwA4jB2GG1vxkSVZ
h6tFAVe8Rp7ZTI2f0WSZqJ8eiOtkdEgiAFcKCuWAcNMc8zHZDJXOa5+HP6qSBbW0
b3mHKcdbJLnxeb8mjB6ftSyLsGW24OTRpb0ka1Sk9bJcC/RtfAlqTMbSiAgsTZX5
Udl6Y+PrTfygQM/5h8ECcZXdVLwx+dLd22tXwGYGF1ZU9n9Yd6zL/38RY7lBd8YM
4UmmyNUqn1nYVChu/m1p5dZ76mt+VnWf5InfEmZny8J0J/VdoevsfTQ/70rlhl79
lfBF2N6C2DIJLUCCb06F7EO23rAMAJb+EKmHCivR0hD+Z3pb5KkG+FoenGFPXuve
N7zkt4pstkJQzrM3eC5w8UG0gQSK+M+iW/8hK624SOpx22gEK5UJY3LGM5JGyGUz
Pqe7CZYKByv4rrA3ZCahFwxICj48AVNAY89T9u7o1kntYpSecPidpLaxIeNPM77+
xJN+jSOwelwQlg+RdXjTCmjI6ZyYncQTD4hn63q1mcHckZ3svdBhBvVZzi5l4KKh
a8TynzOPrJoWopwBL5mut6NRJGOn+T8EE7nHvrRH6MqPmXjYO0JsQMp/0oj6hHNK
R8SMbaT3dZ4AWh1V/KW18ifCPKWceAUJcNUDCSwUk4+Pv5dVsF3EauiNos/2lZz8
u9n7I8jjOld3+XrGKW2nSSHLePNWYDunvWwS5yNCde4kLFfKpX5chyQRg3g02jHD
xR2qOvRBGv6eNPVZRKGpqY6Oww9QFcUAz2IGhrf+7gEXeOjTvJz/H1k2JC1LgXIy
3/e6jSFABv5zEB7Q2TAnSliVHnIRVX8fv+65r7ricO9K5e43c5u/COTPMHTlDnGP
6YuOWegb4RB51R+2xW4zLtXMh8aUwK2CS8L7d4lj+ExWupSC5vRjWSYCC79El1NE
RaT7zKv4JwYMVHPYg2rQbJk6Mwp/T8IBNeWAEY+LTaru9PmxmGTVahB/d2e8PtVn
GsIUoPKevMRy5PQSpX2KRbq6m8uHYJxyu7CKCNbtfwm5JqEJQRICT9UoQxCEyM3j
8GV1ZMGKeL4kljYL0xoJC+He01ci0tSDImN0o2MotyNqp3sVHHvF98eiMDg+GZ4I
v7xhoGxCzVeWa0iyGG7oZ0v3jNrUsLdten1f0lm12KKfY4mlhOKVi4p9GPpvbjws
L2ACX9GmwXeZgZKttYsp8S7mtItaWTwbJhB5Ird3EjzzNJMygRdcpjbti5EfaFUQ
75GiXPVND8hVsqZ92r/BnJYrnMz0UKpT4mL6cKmkoB+OKdYTLfwxxelQqVd9u33/
UMJfMLvKkIeXzgqqdWN0PwW3vj95GtBugk10o3GZeichx6BsTbOednjMydTT6Edn
LcyKmgQO+nExVxVTci4oFuvFZzZLWXKFZuU4ENPGqa99wwbndqsUXx6603kSfNMP
FAsHVUuq7ZJqzQvBjpbUsewpTJTMFPOoB8hkicmkm146uJLprTBzka5J6xbQ2Pt0
07B2zvgng1hvbKxhb/cBqDrfaxfDxKy12MNagZhfoFidQbpLDRfRLiHXnRGEhPSC
QVs4ai7s/Arme2jyKw77O41bx2quUdam83J1yMSB5npF87SFuepmzEXuWPU0tta5
6T4Texspb87avF48lmyHbWwMCr+unTdSC9G/fFJ7xVLBHpAWBbhSxsxEMnUGezSw
lZGT05HGgazJ211SJyYWQkXAbwmukf0CrgQbqx0oR/vmlEWjA1qojrS2Swjj+qHq
gr5ZzDaQUZuINyYUrCbbAwrHOYQSaDj1EknkgvyWpAGnGXVLZlEmxBCEdEcJqQ5m
tQcnfdOmfJrE9G4SkkSCSPtyeEO6sTTGLN3MtwW8WanYL4aB3SnJpnIgSCyV3ReF
sxgIBRX5DIswksRHwzW50CH8x93W3vwFxo1XLhhpWNW+F3o2185hrARDbxl4JlmU
mmMmH3Gn0jGl1M/iXf/jyqr2oqff63L2DZBHkMgt4dmEIsQiuSt9BSbDdHHJ6xfl
1qQK+6IMhONePgslyUDRniNPyjuNKYoGBLBKjkFIP/eKTAzl2JMkpqnM+GO1YajX
LwPLSFeszVsHyEIySREx0MZm0rCLuStoPq4+mA45uevk/fGv2Y+PLRA21sbawDBD
euOeSnlATSAoekf3NiZ2uhmLS4P3/ZmNKLZaguV8XUNl6jX4akSI8n8hci/WYBmV
m1VHT5i+1c1pgBLl9YmP+LUpqAI+WIX4nJxjgg9tkGCEe6dBL7fh8w3tqm8Va1n1
tHw8/1l5dltb9xYlL+lNsvqFPjiX2gR/LCwLzHSWHIj9NRDm2/Q9QIJXnkcmpvQD
Smc0hoCg1qzhY6+r5TpgNOAdVHoukd23riLbfJ+li00u3qacGXburXIrZQ+ueipX
nQiWo71m+hF9QvQUejEXB9Ybihb3duUuhOmWKMws6Yl28M1fOU4BgM8jSRWoxb2c
4vaLOE4vByRf3yaNnDYuFZlWIet6uGDr1qNa+tpWMjEdnrMIUS+8hN2aYcPrvKg0
fcYDigNoKIu0Z4UEc9VyLBRVblDD62eDz3hJ7Pt2Ps9XAsynXNo9SAuFIdo5JU7O
vL7Mob28et+CNAfO0X7A5TtUYKbwyf68dJGJtOwRVorYh5f93geYoi7kyR2x43vA
9z2hnUQnY6xWBs3Y8d8hMhq1gJC9YXk6kUbhs58pVD4JpJcc/YKpfIAtHrsK+I10
x3AFr2IL/VCMcz0T2Fev/5oQiLuUoOkCccZ9ewJ2PK9CcbPjexWjLK3hpJdSZ7YL
Bl6BUnoIrwxOprlYoEh3FVvMgYeE4GXoDSwzDh7SsVBLVMjXqViKySQX5MSbMsVc
uXxOr41kf7/ukUCyx7BfMinq4C8pMTM/gdtUVqX9q9Xz1Zfxf/Og6dv3IcfVIWMk
BRezKQ7+YleGqqSoWODIyg4u8eqfVPFVIy6dxrpvqQ/Xcn9An6D6uh7BPLOCgBag
T3Jg9Kb/Voa6nuvKisVpHKso+Fceqavno5dhoiVdNt25JMBfVZTIdWl6WVQRoGiH
dy3eiRYK2KP9jBDdtax40ffO/Rzc96nOeCmnVIR+5XlTK+m6R/KpHZozq46koh5p
qSSIpX3VQYbsFoUGdNZVAIXzzvoC/URE9CY0lDG0jHy0Ddq6xmNavXGhGqjXnjK2
5+ExJqJDWxR1/yN0Clx7wOElBSswxROPhOQAyO1A5T5/DYJ+kRphoC4b48aFBHum
Ez/J253Wblb47Ahv0B08UIFSh69MUk7/L7+Dzv5ZIJcesnrayblNqW7jw8v6M1YE
tdtosPmEFDdPZ9eN5vCHcV3mitOWQKch2zl7cwCd8Mrn/Odgw2pS7/TZYh2Cjsum
pq7BfOmi3ssaQLiW/yZ24nfyNlyum4mYRcX+R3r88na0X3cza4IL2o+L0qfOPZGJ
Y20V4SRBJVqKCnTR3RXMcApm8sg93/rUQZx/oGWDuMSMx0c2TCrAiDeyqk75NGPP
zfI5T/YnK/QrMQmy1EgudahWwzHBMhimpqgDurVvvqR8Bm9SQjjlnZehnfFNDk50
sxvB+5eAhAGCcv7h4xWL07QKWnGCA0yGzPi6vZhBexTc4qfQRiGky33bha6s5byS
1eo41BAPqd7ze8aVmBxjFsFqswqJAHtrLNBM5LHLw1XzQmsulAZdIpHISnK2GaaY
NafMBiOXxVWyM2bYeHfbaM1+ktDQbmennPxryQmAYtMPiLX7ray9aLFYg7quT3Mt
pAY2aCKg2Nor1qREhcVYiKIFjdSedJr/Q3meviWVejmPg1rvywsHnlGz5LoHFwZU
ZUDebeXEiFWTl5G57eYT4JYIXiG8qIAVwXM/wOWFl7CFk7yQliF2DirDelUMvp/E
+/wSOAP+QYBB2AUooaCuVRnwEBFsxtfvlen8/Q1g41MtGRCQNlxKT38Rcgw95JA9
eFPqYvu+wkbW0TPwJfP9bEmlpA0emCHgx+jXL82IG0hI+TI2p1cWtxTzOTa5Z6HU
FfhxfKkDIDONF/mb9GsKhImrUtbgqRIQGZTlOHG+lbXvbioY+QHu3zJ+hLhOCAS1
qDOrnsAPAtLQhPSb+iMteElz5drTBg1fYytZBch2St7dygFGBAvDaTYE4nn9dln7
63+mwfnZoAoKMieKrEijVKD+biCWCm0ksrRgZnLW0OSzrRDK11jf3P8hvOGcJXXh
1f0BeuVLyA4heIisLrP/Rc/t1RLI2y2brmwcYez30v/idJQTcwVU9GmYCGHKwgqL
BV0cWYBN4+FsPdOOUjXEijmgZy/U0RYMRm2k68O97xaEgYAjGgDmMA01ya4Vu4Df
tCsuL0Mjo/CuCS12+ez1nsP5LlhRGQK1dXXUm+2sYvo1Hj1Gl6hBe5t0XZbxTixL
GIkAYSu/81HEtExliVJVt7In904fBN+ZEeI530+HMGBiv2ubsxL0z4B0eSdJgwxr
+u2awPacwwqbk99ggkAQF1HvRjRCyVZXsYxAsQ0XPyv1DNVQ/e7FG42GIE+R6p1F
FhG8X/uTOESUG9B3b9cPYxAEgwkglj88OHl5mDEb9+Hs6AjV1NLcdNC9qZ/wvJB9
9sQBPWnSWn8r2hrJcKQvJvt4boYpyOcqn6W8Rx8IISAXC6c2MKotTDN4DHOpv3ZI
W512AC4wKIwHj2P/+HLa2fqdifJISlIZ1eh/ICmjEnzajMksyZMnILJtZfJDFcfm
YVdrhtMc480frcqOUdc8c3Sfo26JwQd+/H636QC5VyZthU/282bqgpnwY+suOyiH
Z1tfk3/PNkwtoW2BSe6OKEe8fSzzwUMhjM47ZucyUpMKc04LMVdQFv8WCNNBW3Gk
DhxdouQPUrV+YK43X7uX8nOFyfVU+1shf2XwZOkTk95vfX4qoysORs4oz5RC5ICO
MKv8Wvh2YCfFnm5QtVl01a3QUO8XQ0IrlBt4jh/lSBAFpub0sT8WPUvFrVuJSFWI
PkeoZfdEOSUDdDLjomejRQcIKkASrTxqjvLYYFfr96rUe4CiMLMK6rxd822KX0vN
KV5yWuqLJcENM9rMqBT+I+JD0OFiaOj6lbrY8v1xRQWzPpKLS2mQplAMrHseIkyy
wfB3GJ2wCunbhbHEMkEVQFJpxpvvccnCGnpmW6ZB4OdkJ/nyMj5PDdWH15qYwW68
QJVNNd+Gc8q8KzcLtFf53m3CPYXI9nEvT9cA45/zCxOLUNfIKsvcP21KErUYdMEL
ZS4JjwkshmIAhq1YAXqjWEFfzhAzOV/y81e2sJd6/HYKt4sSWWmklzu2N3j+/JQt
w5WG8yT89FCKSknEytxY9Hkrqzi3qA/5uxLb0yFleXde5u5O5BiwvvIkq6oM2Sfd
sJ1gWb+UKMyzm5pUk/vCS0buB/BTcDJ6raupZ3ozNF+lycI6IuIyiDI3o8npJHkV
ssGichen8hy6zQMKSHlAlsqVDIJJcaah2idZqcYtUzbY+ywNKTfPxF8wMw+pTs4d
JCQMN7Ni6VCSBBuFw6GsPTat2DszCCl/zNtXYDUQJxnHsN5T4ufoYGs9YCyDD+gV
+OEB3+TtKYIz99gMGfl+HK6OSU2jAuGMqiphQVkm4VlrCHfG+FPaFoZ6ZqAp/EhP
U+tYMsqiSefFHkk7DXoj20DOlB5MAJFDzbFO6eBvZghS8y5SMwhE6jyCyKktudDt
r8+9iZebgEsjxezEv9XnpNEWzbMRuNaC0y7lOM/PM/vRT0PtGjDqq3ZFFOlMp0U2
IhJEi+0zY/9CPKWoOqIy/qa1+J0TEqF8mql/i5WDL1rHFO3L3QlzVyCgcXWb2XxI
JgB8HA1DgHrisn6vCScf4SEkSEZ7cTIGtss/uhUml6JwXnrFuV1fw0tYp6Bh8wLB
mXS08liCbcy7GTp+aQ02kXso/xOxjvCFo7X+nVxvW/CNSqrJjwW5ET5tlkYIWqSg
YWlW0mPxLSjsfX0a9vsNugo+JoW0VrsbdIC3QzDNJLuLcdojIfEQ1pjR6ywC03Rp
4rHX6GyGglIzaP65gkIBfdODutan64XGiNTfTwvWfMRpAfofdxdK+or8fy6RX5Q5
bUaTNpIDUT3QGhjRb6n6NqnbXsxLbtYxYwHhqVf1Z+Gggx2FlfFUkUmGewqPg5mF
s2TVshCQhOaXVTyfJizTs06aRMy/NGxLEkQIPUBwOLBDVrKX/ZxbrzFifyVJsODN
DBT0hho1mok0U/JrhyWwGeDJAwatZcdtx5AoyjGB2j00Vm+PHtWZK9uWL+VjxBWz
dJLLX9h9a7i2acNJuca/hhkoSIK6FUolFpVJ/d9F6VJLJ02s8JBRC9ZwHqW8exA1
l4Jjgjd7LO+VXYazpce/0mm1TZhCg++6MdoQJlhFF2IbQHR1j+mfCl5nNVd4asJG
fSg9gVBKths+C4gNa4ynHUeEdP81rTEMpiug/uSJ0wiUEFDf8qrX5WHASMHyomb/
+iaP2R9qryyToGrtpQ016k+p+h496UEgtr371ZfstJavh81DdDFY8Vi8wzL7FaXZ
MLNd44//QNxnzL8p67Jc8UghYIA9GBdywxaFvG1OSJohpiRQXo8KUBQQob9zfJel
Bz/JjF0KYoILr0nsaol4BHHmuX8BD3V5T9ddTIMsKo0RaGQD6YYzsgMXNGPCPYbx
6AwtzuqZ6cqt8SHpdJqk3DlCqNozTRBHxvI/BVxfP7bDey/krOGedbn3/mP3qO9U
+VbQ5wQhMHPlmosVg/fltgze/c0Im9Ow21LO+OKvlq151BdGmD10Fsaue7Cfv3h4
w5hRjkkrQJTaOU1160iTL/t0S53kenoD4Rg7HBkFNF3HOtJaL+M7ean6sby0wuBH
8V2lZfg0/OZtlVJGj6IywTPvnb4LTNiqYnzm56aa9s8MaaqW/tFvW4dctthv0REF
2MUdMaOfUIrFGTimH5P0rkD/2Yil1mUHUaH5YMS7f1hUEUnPvqS3AYbVbmirBWd8
RU6ttJyS4hsrhqI5Hl6r4+phUNc7kEYIDX5q+VB+G/ffopHPForJrDPLf/b5M25x
S4OM3VYdMcifbfKoxVcSOwdcyY0V/Q2OyewB/AQEpPZ5U9gojruj22TZX7sO11Rh
6StB8r6HkSMNv9IneBf2667saCBmxik1u1mxN9OzKhArfBmuvV73LalXugWmiFaN
7f/PC8npouCj+/26z1/61eZA2z2lISSlbyE7xXH2JqhJpPTAeWMjgxPPMjeqzM3Y
l+ixP0lsGF0uFgqdGO3o7wwCgFbGsThxEEafJ3xs2GgVH/bIT9krdT8UI/aSfWVd
54PsV5eNLVdZdjLbkUGcyH2wTO4dPgFjJ3fSFSwryugA5y/K7nqs2Ojq31MBo+nl
LT4ZyDwkSWc8ldGJ/PkW/y7xAcII/mrPL9jON3x6DS/HxL9xaSBUSPiKsRHQkYYn
PrG3t51BaynzoBQ+vWz234ex/2gFmG4Lu2w7Y3utd2B02BNgJckn9McN8hnWQuhO
pyKu3Do0PfDDCU5guhGJfJQ0A4R00ZmpRcC4r90sB6h82g7KFsp3padf0DIf3lIb
ZlFtW86+XvrpZQCa1QaSM53It9iASvb3muvg1Qe3JtTjFXPnPiXGIpxX69E6r6r/
EP+LSQEXUu6f0ndJKVkrvMsMsoe9pcrwqN17mNRNVcMTGBO0SCeenr0Cu1l/4P9U
zm3gNDsF1U3OZ0C1ioVGFRP7/EB708/vqr83cOWaQrS/qfpHkxvUEkdnROnr1wOH
mLtlJ3bsiKhpF4kcl0NXCx1IrqsyWd/sjtCOteCsRFkJkpq3gsqzwz9RQUskW2of
BABMiBK1nthcikVGed1mqiX0vI0B5yBQdPWGyGTZb9/Ahog9EJIypmfBoTAVIjIz
6w7A+L7D021ejPWD4crf3QeqLgrVMtTANskXdIKvWQ1GMwCo220O1MfyXZAfqbGr
Cr+C4jhG5HzKYnJeJN+fxUJS7pi84N8mfKmuBAPo6Kwe4mCgIiWUzeEtKIEXwugt
aLPL0kcHoqEMwRSuOjexQuR6Bcto6A8VI5KZkB4f08OROPaJyPmNPVVBNy2L/vTe
OrFL+IfDkce8pvGwkESNKATiyGL+IYSBDhGikcAb6bO4PqlCVudM1YFd4NG40fF3
uY048Eu4OSJZRlhUYkQMTphUid3N2cSOU6TjKuxBMQTTqKY8pGIQtbKe1iXtVz8P
kfZ7MBSjg5gmYFehGHKguLASThdnJc5qq/j6qxjropGCMuBlAMRRlLgdAPyw0e4y
HVgawxa8JtJ+hd869WzeEDA5MbWgs1lrFPkcwIUJBCVBtgn8DpTfxQD6t1/f1leL
F8qsSUyw3hob3foRLY58NUZjdbSxmqGXuwfP4733pZJBZFfDDJh4UzE60FodV7bt
VWtky+ak/vi0ExVjL5ihz9SyscSJK/1t+J6Dqk/YFF1XKumwEyEHYMSbNXSMmiC9
+3zB7J0/Xl07aIUGk7vWRL9WNm8K2ubZYiDkYgkxpXwmlygJkI3ls1XQ72FYc7Vq
/pImzD+0xz2SR+ba49kVxiXdkO3JrOwlN3zm6NoA786Reve0GvYKHFRDpFmwvAPH
HqyvL9eK8t+ltlt4cUTKrFYHuVsmKAACdGtehJyjDL74+WfqrwxbwDwSmknFJH1b
nZDpECLFexqdEc7K4aS59UJaztomWeEeN/VyvoUlwftdg00S8RG/R2x/zH2kihck
wJC/vHb3JMsaSB2rpkk4V0zHiHZgZVvjx0HHYIVqEQc9KyYXhP1Kno7SKqo5EDwk
MCLmcTvhcONnmq3mYUTNPe6KbyQrcmPyoSb1uorCnt+auD2L+/aYZGm6fjbKVjNc
Y/TaTJh1KPzuqyr+gwgQd/vopA9eIzIWnSLTTB0foGAjafMZ068wj9jpgN9HTvFf
glYcumKbl0a18yECUZzX5r1SlGlGE1I/JyOTpmxCfXEKYPtEcOZQY4rUUj5tNIVH
gY+boxj2aBfXXvHl1zMmMXosjD4RNg9DhGX6MHm8NWcoiLCoMQRAO9GJtn15dPJ/
5PZjrraGCK+r8JLv+d7Jr6uMyawt7o/cQUhmhnpdMzK4wYRqIgzvfRhPxuFycqm8
vpS3PnGevpAvgQKbWJbXPIs1GOWHMU6FFTzPIANOl8LiEOddBJChOi+cgJ5pZKyj
anfcPQjqRxQJOTRTI0NBF/K1GzgkisVY5S3a4mAtvAJeZ84Hq/Hf3n6LTpJGR5LU
MeTKQc2IJy7wUdmYy5J25x+9GQbh7KBwmHV+yfFk1YM6nagqUmowCooQGF86Vfjx
xIIbQ1VRZ8TIuYAhgZu/jAbhelP4xknOECnNe3BzvuepqRlzGxvy//oTKJcy1pdU
GJEGK3eJDUBzxI+NKf49+stCwczGTz4N1Th/Jd3vzxpRCAiNLJdpH119ir6+QwQV
JWU/Y+kfpu0D79HKZjYFbLGhxxnEfvLWyFf5pTV13aSrEWazcGYKyVWwPNrA4cjs
SlbEcLabm9YZWbGbXI11ColjngBykZmtkVrvwUpuFW2yKlBu/jpUUoYvzqqJHdnQ
UeXhgD0OYb8OLnXwfo+SwU9fH7S+bBbnKcz/rmRK0A7y3Bx9yvuPCn2rL/hCnV9J
U8/XU6ZkaRMEmLcqHgOwiucmPYnt/BcE21LeFhObj8PVdl0npOHNIjRqjtEt167B
v2VDj8wgQCa9GBgTHyNHv06ks+U16Xwk60Sqzm80fVW7RPwpoqfbjMkPtYYnnaDo
/6L5WDFrYTEZba5nbTO4/BV/JBvtsSIy+olK7tXPKRaP61JvKs21emPGVHBp+gyx
1WQ4lAutlA0dmzGu2BSr+gt/Sfx8ly7QkFlH0LnxdDGZwsOiBZ1B5Q/AApHVbDXi
cYzc7iVphtxki2rFq3pZHy3cqSJJ8zy742bOe8FyV4cyKHTdDNN3kYZB4lLM4PMJ
Fe2YZOyzwcRViqnxJ0IEz7kfWC19HFdizDBCR0jKBDLMreZGyWgchheu7pdM624P
1665+qx6Q1z2h5xGT3sJA57wV6dV06kb95CiJNCrsmajSa6Yy+nwHff5DJnX8o1/
WDdcQ4LuknECvvArK0iw1fJrvLIbB2G0g+EC5N8IpjACC4a65G7SBAxfOhgJSo34
GJRvTXIwdNNACruH280QTjdLLGTdoCC/JGpUY0u6zfeR/t07mZ6eYmTyFRVzxpjK
68lOj1S6vJQwhiKVsTV2Wzabz/AuMwHJvQeryi0imMUcyRgdG9X0mOyKV4KzUPli
al76/brgNdBoNc6diBuySZy5x4WiHzNKKBQhs6aF+2oTq6/A5YM6IX5vNRwAKYMK
2Sdrz+KHgcngNdrym+GyM/Kxeoz+Jviw5k2WAWDI2xgbFRbBI1zLiwIJrjcuIFQk
Vc9U7jqjuKYhdJjMiGhk+fNnVbirweZpXQKafqMWRSRkBy3KHPMzFCek0P9GLUyD
PDYrekXNzHK9U15+LKgvpXlElZEXUy+bcxSzalSk/ejkvGXLkJWbU+6oFdcsT46n
`protect END_PROTECTED
