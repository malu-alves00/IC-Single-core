`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iFbMFN8Jc2jwjxa4m8Hkfpcg+dGJQgRwrKpb/R2RzhqQcQUIkC9tQk/AbAUBSInQ
sUgPWzeMJXNgKXe1Qm303CtGgJ2FXwwbqhVqBwXQC8ezO4GMKZgnslHpH4092080
XoeJBQXk+ZWtTaW3I1/XMt8QirkwCN2RkqSLMdMrfExG/cz8h2PQGem7YxjEOwQZ
vQ4lfrAVCQp0eBKBjlPbgHBkVzKyaD6/ZGpY3SpaHDmY/q8Nj2pLWCsCD9lNf0pX
ml6n+ex+x8Zb81/4wJ+H9ncDP4gFMoCJu2Enb49jVsQhd60WCaPZgHEO/yXv0DVP
OopUfyBXRNRFqCYOKKD4biH+bonBD/PNPhGetpJ9ZAdCygVINeNJHboMBF87sSuU
pg/wkHXdpIpw2lqNtw5El6j5AjDSL9nFMcZ77hzX25avl4z9ykFpw3gFBWyfvXvy
2c8O8KlScNoqxu9fWtclVE91/IF7sSE9HOoFGVGY3DNLoqx6dQg45Y77NK7yjqml
78TpbfSRSAhQ4zG6L4j9Uja8XhtzVDGfKwr81CxtA+Vpk04iAK6K6x44t4fTF2sD
`protect END_PROTECTED
