`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pDI97276KY2bXC7y3v8GWgVcERniyDrBlj5YYvSnZcsnLgb5GZAsOU8YlExj29IQ
/Tr41LoH7+Rl10bcNed9Oegz/xLQEjUPYnm/Gjw5u+fymWJzAhDyR/4Iuz2jG125
0gSfJRP4iprOHbIL5q7lAiIaeL0TCtN7qXjofvxVEs/7UGzwj4OfOj20dh3T5LC3
txQ3lQLtK6dqZVHdZBWJy6XGvqnG6ysdu8pLKZ1LLeY1lcVuXDerR9uV/Bpp21bM
BUdE72pCYRkqMHLZlpKo2jOxJUTf/O9cl9n21VvWDJJk47eKneAeJG/JGaUCEzJ0
qOK3bqRYY+Vd/ByotTH6aPTStgry+FlJFi6l+EEbBeyG1wXMQ9UQM3Z0Rfionc3Y
1MKwtoyuaJqm26YtsAP9GEFnVj6VIc7LiI4aDe5X7BMy3pFU++CCpEo5KCePezT+
YNGYni93Cik/HiOd1YrajjOv1KhasSDWNaCvwAmX3gm9/rkWyC76DZY48ClCLkzK
B9398mvN4tpBNaJZbolOZXr3gYGpNw37e+LBk3+wptgN8/bAgBbYOfiTwPpsed9U
0cHD3T6vFmN1d81/kgj7JkMDzvxqw1m5KLRat9Wb12kZjk7UwoLPX86U+cZPRciN
PIlx7tSayQb6SWNzYHEnE8+bM2n/Z485jnc/izBC1jAf7i92qWryWq+TOkMAD3oT
gCRCX1nCfGrmNl3DQIDQl2v/JcamPcjV/Y+VBY7fy3jbeJUjhXsfIuY8e+vEvNDI
+v7hBau84H3NItDYpd13zwlB47iawFyDojE2TJlbXN4b62vFxooYyQscqr7Puayk
OUmw2DWiLy+Lbc/nRQUKNe1AIJlCnYrPLWHmbtocHmGlhe9NzhhJnufYdO8ygrVe
04JpSTjXm3KZL1Gso2rKneequCjFd6VyAeRdkiYospR3KOGL4G9EVxjUgPtGvluX
WJhiY92bc8WgFnuB7WVnztP+YC+sb3ybE2hacnQikgsgnVkNgtAoZwjvl8ZwaJg7
uKxaFfpRdGK8gW43xdGoU5oRAxzTKP4JUDdx0tp/AVPNekOUyTtsjCa21QqAFNIU
N8GcnGDVgrxsI2FxviO/ufzsTUWCAwr2idt4GVzrqeoJrM6XNJ98fXrrs8ckGL9J
7U+6GFH2s8hFqSk9Yqo6uSFRXdIbcLXoedAV2OrJ9wipH55PHIC10pOH/RDyOWaV
VhYIyi5/FWjI0ZFco8ZoJUVwPBFeXDS4OcNfB0Effigb2WST5HsbaDbymkc390sU
GSkGMSsjUhScgVtjeOFtxX66Z+lqOIzYIE24+UyErliMWRB4/87LAnlFffg4mn6E
uJNzeEk/6PuiUYbk+AhO0DAvsmh1Adicdj2D3f6bWV8KdQPGCcMUoamGCdvwBcfX
faj3IMI1nojpD5x2tM52BqfiA/U2ouHuW/50ICsnI+6VzDpM7QN6GDcNdCtdMGab
ceHrbdIsSHIVnQ4oRBscgoeM/ThZJYHFb2PZAyuwnk0zRzB6a+MrNEWEChFBkPj9
441YL0q9l/Xr9t0de/c1oavhdzcOZfc0NrjP+1tpaSiQyHGu8Re5nPaH8AMy4MrS
pPajXT806uHM32IiVdHCuzaLrkND3AF8KobnygL4vxZBPUb90z3stxaQqPGvK7QS
QL2ogAOfzqUIiD0lTxauh0BvmD/ouNPThfcsJM/hTlVFp/MDbknBFF/ohLy0cbiG
sQPVaUV0XW8CJT6LxIQ2F33qhNn6tO7YcoDaTi8B5Rc4o0hIpgpsUIQN2nxDtEfz
f0/J365Ix6yCQL7vYlVK4jQZ2S5poU6v3HWu3NL0ldyeAY0DOlQWHHykKYdHsmhb
/Dzq1aJYk7aq23TQUuuhuLrcbJ7h3GmoU1qnrDKBenuuEzTSMQ+mYziyRkK0LaVm
rKwy/GMKLkJIg0W0W4Nh9Z+wjX9yCpx7KEXh8BvFjhD2pPbEKs0ArDm0bk4foqgr
DJ6hIDOGKa1pCBVLXTXB9ut9OwnmbHemBBj09JOZBNauD9p8sdII1GvI9HRdzFcf
p+MWa2gyMNEWNuwNwsx3LNXjSklsaM+pMxCgzxhR0nuqo+O46DY8iK8uj0VmuSWQ
Fx4Op23SFsysnGglX/vC/BDYyME75dHduL1c+wicRYTX04jMsp3HqJfSSOXT8uHa
x1ryjLfA515JtHmf7+aSeok78hhCAgy57Kuh7HJhNzyrEy01HO02M/4lJXwkOHvH
XtXhSa+I+xBimxsaLT5wDOzbTBwDaYOmb0ElWxKyiXDzWQBXkepA7JvyYDV/09e8
5LxocOgjksJXQlNrmHFserUpj5pLQJBeLnRkjvybcmdnl1DHwp7DPAIelZ+5DV3x
uS/w7LgloPr4xCJLhP5+CgQCD9MiL0Jh80fEeeJPgioiMTlrePVBBMzg7FVy2bZu
VxnWBis9g7XiWI6E+PVGlCxfHYAir3f0+zPzreML8YP+/cOUR515Or+cIg58aRo7
GgqVnCEz2tm1fMeferIO+Fwi91iDnkUPMrIVeksx/6N1ShM8/hj/zXdfQEuO5AaZ
ipN3pl6Ag46D86w938Ujl7UpV9WPKWhwUVo/3e2AM4nXvRt8iltoRJamMCLr3O3S
RE1Y4ijPdu2lYjFg0WQnXoCrK1H1zQchve5qVhOEF/TZpvZurBJX/N3Kza47idHS
HyqTd5Aqj1CpdJjOGb/QymaDZOLShrS+LNOn1okHKadwDWfrYP6Gonsdqf4KcBSw
XueuwuFF82d0y0qOpe+e90YNKFv94zYBGdNGWGl0znxONdmFlvBBVZqmlVLLWUyX
3isbh8NRoz7Vm9gHmLTigwSGhVRTlmxMxEIPsQftErLOzbe8QsHaeYEfD/tuwgjB
ibcYR8wCQwtbyFSwx71Da+Z/LI27v0HL7k385jhc+wyFwLlwkILjB6QVyvYs2kIO
QjS4gqqpN8gR0OYxNqvwH5dHokyHUuhjh1IdCdRzs2d2wfuegu3tv0UsLN38KZEz
FVnMoh8JfmfT+WdIImO8K8mgo1MXZNDXBBXGoCL4OldmMtQZ16WXF3DhV/aHjB0S
GXGVnCsZpujXie21zcOt1rMgsiQ5z+1c4XCzKZ3pM0cMkUhXqFh7aJ5YIQFSySbX
aOig0yAQbW+/6zCHwV7I44c1n/DMMcWo9oHCO73hNQ4Iwr6Jbs8sCLpUj1p+b3Tb
J5y/RXCwnOYQLQW8WTnryGW49CV9Ij6ve0D/jlNMghgotArUETQ55jx8T/mmo4Eu
eZj5EYIAdsiU0zasO37WEVaV3vmN5NZyygDn722Fm8+JMQ4Wfr+fUITO6b84UfQg
eVIzyAAcqzS2IfhmryvyeVQwwU44Vnkr8PH2rbqHn7A+BAoOxRNkD43ttsyotOBo
1op7p/KKkUet+Xz1M8qlu4A34DijKugYihWzczWCD9ryeOhuwHvVccxVFY9kmdIn
cj3xZvh+bkX4Wnq7EjpLrVjJnr3Dt3qLV/D7nysZULQjIoCouj/ezXKt8AK6Ipr9
8efOwvhWFkrpG7puiaHtwDzI9Vm0+6VPzL6jKrbUGjU6aKvHxa+R2uB/RC8A+i77
0jx2tkKOYQqzKaVvykcpYY9TlWbFrF1EVGAEmCOXxPN9uQzTCAKl94I8o3+XxoJO
orQsoW91vyxMZkiG3XoHpuHK2tRBM6GCmeCXZIaG61cxwiL2GtXyt8ztUneoIjUN
55JSzSEpnyBnE6SFc/61xw88noMZhV67VdrUKLuHAsAGFPVWlF91sgQkpK0MNreL
5yk64nza3MDgRWWYg4y/FIGmkwcdChLZ1yGdadwa6+wvLxnH2hQrYjkJeuJxEHuA
KE+hTV58uJxES913nlwwOXmkAeK9fY2tL0lBh6LWDp6ENzBwNTnP/icYexOTn+UR
LJcJMRqCad513QRfn3x1VHxrD+rvycY3oKo1yU/ixIxT1FfANvqmuEL2PEGHsM0H
6bYe40wCqy4cHqaPFAk2R2N0JNmT8jUUjpdn9Cq0Bh75LbUYUSIuCDZwu4MsNZM+
0POguU+FWgvcj2vE+tVj9hA5yxCMANBVFLIBgB3EvezoGz4LrysAmKU0WYiCm5B0
WpJQM4Ir6Dwid3H3GtlUQB2Cq3Xieymmnh+q9gyNWvPl/YJBogiirUqD3w55gVwt
9MOD5uFrLsb6dU9KcZDB5O2EhbnIQPgwGHq0htHxym1XEUN0u8s6r8rFeZuuUFLm
tbcHnFnzYfF7QUSXQiyc5sgTsynKDQcfTV7zLEgqiwqKQIRQrm6WSw6U2MvOpoCn
Xo9m80/uHzi1PsTDy5iSdsolbOxU9oNROwkteUKUmH7qZDiISJxrny182FdmfwBw
RGxxrCzKceOxhqz6xZ+qKWUua6GwQWNi4oSoj/Sm0zLnP+rKJSlVHlyo+v7pauFq
9iZMMVIDWNgFc7BQyry68yPWDRA83iMrAQQX8y9Hfscx+twa8+jVS7Lu6hSGZJJH
zROqWPzL5R2zz+IBOk99+whd+NfmUI3/qy0DcVKMIdk0H7H1vBVyIWljC4kCWY2M
rseKBFCZWs33OZN2hIrP8JFIZFvsMowirlcP9rhwBvbGzzO3ZN1ZOzq5SzMlp1Wi
u1tgQ5ITvAH7+15tLCrj7flJzYKMXyr/o0MTQfGWHYD5ZFMgRByz0wrfNkrhl3tS
iFTtLzjXycqUrhELfgW4vYwQKu5dvd/naMsoy6f+4cHJ8CeqMm2mVvAYwAFMG6iO
29njTN5EtggZrRhS1G5uTIiyAmKd9eZc1ZCiqQoTd/8dXItpK22fOFRO1VYBMfma
N8e3vzzVTeWvQH8mK2HMu8H0fN2WhrEccv4PQH17eAFMYNetnm5SUeR76kZXPZHQ
YT3o++O9oL09JubPcCHP7yppFOWtf+NJtcyXHa6YkU+NRtibRU6QT9voLay+qUSA
5BVTONZeCPzFb6Ndd2Cz77Ub+smlWj8VG8Jg5vjHiCpb5f+pcOnhLHqTI3EdYxxr
vutrTi6D6K46dd0beXsvu9Eltbfl74PNWDlAR83xHbL50EBvrUefSWTGbZzuXsmG
DSxYQVfvJHBimsUv+YFJVVUsA1ZuUncN+48dY36zxtMngVaHRjs0dEQZi+nAbM9c
77VW6hE7mi+Sw3rJTFSxlHIhwvrSMZ0Fk18+MqSOY6JFVPYu8IGXbZMKLmfK0Hag
mcfROx44+KmlZAb6tuD53JPBtq0jetAUitK179nge+dh5gd7L5xDszpDDLs36lQA
umvNsVQ56sOIJtpxRH31MIjrpbW8wnjSec2WySD2ciVmGiOWo48z9fguWR4/OcTI
4Jfj8Fb5/itni+tru1gLJy6QlsWPxd6VbHrHJQ5aykXmu7LVtWwk0nTAAvUR8LtE
UCrnSHgtYNvbrBnwLflxzwSrs9Q5e0Q6yJ5JzD4SNVq1n+qYvXo+Pw3E0QTyMxWR
cpTiaqhywNIyiutK1TC815B5UQ4F0qp1LuXsEbq/lRscdL2OAIYI2yXVcmrAZAZC
odt/mdQtpXrYutMYM4b8HLoTX51hMWvKfOomFSOBzUfwCIdia/YZ/2FquRa6k76R
KmazEQFPPQ2/Qhx9lyyEIRpWPBr3KXEiu3/zRwWtIs2dLWAOQemrFYwGOAv7fDJn
ERGMaUMrgmfg2NxFyNe0Fxs41T8QnPdEOSXLPamcdlhSSZlY+lrjWwFHWIu4WL5l
sXXA97YweDMfNo9CKAh1FnSIakjdUQ3/Y1hruufXbFvSM12i1HrhgombAESp756w
Gi3+wqB63GVaVnYCuvm1slSjNoxVKnb3Ae3RtCOEa+v7F/xrCiuPCCsW6/LdEaYt
Fvt5uidEmfUuNg22faO3tpO7XqRdnB0ngvd5LJQ2VicKQ6X9LIXEBZo8Xf2DcaYg
VWCiYnqlPa9hRVOXJDrRGBWIETCa3j63cDn01sPJUzwGymij1183c7eaibfN3H8m
lD2NO5yLMY9+TBt5pyxPkIqYHkEBXIQbcckW9BE3CqDBpYXfQRhR8HTYUM+QGIrm
oFiFcscskAoC+aoUAjtJ+8WADvAo2sACbUg12M+TC/hpho7c1+lrznY/KOtsw8my
YfLVGqVeFxJi9izwWGUubX0q/kH6DF5v86gkuvp5dTtWOm4PZHsl46W+EZuFR3k8
1RJZ0GnHFynj3h7SLEN8j/gRQnDpBKWEaTaU928mH5TCSsXpH0HvP6Va0A2HVCsx
yRrpthHPooje9RiB4LbVw+LkJoYH1vmy5ybdPAgrbV5Z4MSk0ZtnJ/XwRkzOeLZi
UvLe042v9vUkLwYQbCw1RXxytFC/RnjVPjiJm/ld5/2Jcqe1aw6+qfdt9yMZ8EtS
usAaIQMJeQc4oGaGJEwl4jZDv1FLeXTJN/NKKgO4WHUnFuut+daT9DGJC0HZ1i+o
CibMIMgVMtnBqeIpywvBvr1YzUXLO9ir7nHsntM2um93G5JAdv935cBtWXKrb/I6
wsU9AoYR9SREpb3c1NfXxqBM8XnT14bh7+GbDZkAMTL34abArdFwg67GQ6oRyiLC
OFtzbwIpTrNmcUcPZvkfKBmVa/XZXrU750nvmEwr38jYgRSbhlbHG8L/1phRslUf
80C1eFsBCgZjhU9Rogwiurv4vXnjeyNJT5JgohVu62u4mgkWhGxeB18oqA9c3ExC
8cpKxSIebqSg0TUyeWI0URVYWxYQ7msYuithvKQd2JROl5RkPJTpQFuTLFV0St7a
bUSAorRpx8q9zYTVA8BoCCOGBV1u88bTPeKnENGI3ZcTW4SfCaqTLRUrEM61My5C
VC18Oa13IA+I+ogtaLI75LB02CKUH3BQmc9Z4HeWM7uHLf4TPCyYI6hEtuQ5aKg3
UZNsUymWIkRIUdZTo/g2lVBIhflFNm97mi0Bacbe297kf8I1FHxY1WRxPM0ZCZl/
gqWxHWgCU148OZ8LvJmnUZbS5qlVkYjblVBBGq+2JoTCgISGIw81l9CCUALNEkvT
hXdUtBxvIjXX7h5qouZyAEJTv82rArq0OD8ftEncwLXTyHyS7y6VE5jlDZ87GTGp
5Mo+TWq7qGw9DHVnHPwlwp06y8YzyYYRJaz7cLlwqrY9KP0uaY3KCngdCnPdxXpz
CDt+5dXsUaZb4snYayX+ySyX8hXEB8ItkAJvMbijVXYKkShON42l6FZPXj9hqTmd
lcnd/fXiN1Te1NkgHwfqSXMESmJbuijYD5XWss65IzNwzzmWaI1ER4ItPCbbfXqB
+HlegFBQynFH2I4s1dkggCVINLfwP/s5kvpQgN9jCBc9vaMen3PNYnaCsoQfSKIb
F2Uge9xSNj/T1b+6DqtrTjA29SCnEr9rEF3mwz0el2K8hGJrPeqQlmI60/Wf9yTw
YnxpkbcYrL3N/8WlDx6ne0MB7UHGxgvKNa3Xv0xR2AfSFpg20zAfI8C8jHbPEpbu
XkLq1FwzOeWOiqomBmuXbuwEjzzIEz+PrHMu8Cy6BPxeZq0s6+bOzNu51WNDlAyE
migklx2fJMKyEEENSrP4Mh8U14oEZNqddEO5OctnvhuWikS59Ddb7vUTuw4rfVuH
Sr3V8ym97dGtgHbDKLGC8UzWOnlYylAhufYP1cgRrzo8/Un00yntaD/89fBgeVXP
wOwUtnxb5UwJh/z+rkH5bGl0pKoZdOpxjrAJWqBC/cgq+n1Ot9AIWTdzP6uCMD2d
JO6mz7L1s2UEnhetnq8b/j1DgRrIio7TI3iL2O5k3OTJKl+38Vkz2dlgA3qiNx+w
pv3QYNE43q8VhxTWDnNToPcZtA6agSXwq3rN3yfdARDhk2ZHI4TfvW+aiHRen9Z7
Mo0DtI8zmkJA33zO/uT3uekZi+l70dl+geWFmBgPxfNmM5pkXhnRIoM24/rHg8iS
fA4xbUnKqfA+v4qDRNfinjVmKvphCACHwAfRHkaGj6hzKLvel67EViH2zbOy/B8l
5YzM6CDkcOaaqQkB/GsaB3Y7iQJTn4wGx+3hNsQhiozMUsLnaPjechiA7h+aYU/p
oHo858zd3OTcq1sDqQacPwP66iI9cSaZQmdKbUe9Qw4TaILh8CSqu3g0mweweie3
tD2+J9e6E1DND0+WVCtFYkakQGBiZheHD9D0ym6atuGDrsJu6Lufpy4HtFzUzvFW
3NcivlX1XJyTkxbptSYZm+jPMzqQT/umLjdxS+/DdWBwOa3PU3Qzv/501y794thm
zT7BfzFN79RpjOd/UNfOgDrv+eyklaiB3cIvv4JVoRpMkeS8U36Ei7Sd5oMiLx+Q
In6ozGpMySA+PUJ5kUHFSz9jGIehYLvHMYAGGwbYGfdNzSGTjyDUx3VPUDrjkl48
HCTVbHTNMQgNkBmrVXUvis8xRPne0ksDVSuCTjCYS3q/0PfrnGEb4++FKCiVBNfJ
LYwwGRKPjcO0rSbf8zQ2fQtOAm2eLMyyxJR2cH4gVzYSXOkmn9Xp6Mvi3wOyrxdw
FdeBqA7TWHF+2PCdJssHpqkfdvlG1L33MovOtyMnybylJfZxZ3xNvynT37UUGCod
TbM2Q9PmzLZgYgLI2LNbHfVAn6r+S3M5PCMS6NM93rHoQyJyiNJXtANjnaTI3dc+
5hALQqBwEpxZ2Id1r68Szpzf6sm/4Hue95ACMNnqy9duu5RBs3q05maftliRmES+
9p3vOVGwk9r0j3NN8k/snJgJP3HDNGaSbcXfDXm6oDDm5dLS7q3qCZXMZb6CVUuY
65VpBeBhOUWfJ7wMLxQ3YmzUByFxa56XEXXjjSKwiwYvbDmibsjLGuB+dc84H/QJ
yX5UhfuZ8Bj9u4vnYWCBGajOIdOrZ6xTBpkKhMeohURt/MyAavfX57MQYXpg/QcY
/hRPkqRl3h0rXApkCz/DSkvw++yewWazpV5yPLED6Nmm8vFT+w36K8WwOu9UQh8I
tSKPCvXfQhJjtckG+DJfVVXVK9vYXdNOgPHmpTyUzlUtiZgXvkHp1Mvn8DqR6SjT
x1Ak7P+eWfZMthU5OgnFDWoLyNW1oiqeNtoKofEZ8n4S77Kjn2C7m/jAi/NTSc57
RhU8RY/mVLgRxywhmBJZK3UHdz5IBgPbJ2BSDAV1c7WbcANBedcyo3atbKaV65eL
EPJIw1JvRR+NoXYNOhWXgv972ZI8NlQ8NNC76n3ObzP8oqtqyALpizOWVGMxS/CU
V/2PtGH2cCVqyHaOUg59b5VTJYWuPxF7Z6k6I5zVE+FkrzLN9/F7kLvE8GGqEo2o
XTyiWF0LuPtcR5kRWg1GvufhNS/Mk6JE8BcM5UwRVdtfRi+lqScZf1+k1A1YSFja
YwVMzt/wamAVGFe0AlZyzgHdG8fwnrMDGai77Wu2DFBaDiXNA1oClmRVdERYsvoj
MRTiORYLsQFoj99HLZV59f4rdWXN95Yo4kgbr6NY0JKjJyDg8BMbwi+tqbExc9Lu
QP53k0TQtioxAtbfW2xBAd60r3x/9zaeogzWKXmIVrpTY/YYwx8kLae6fbv0sjxa
Ax37MszjCLG+Oo4hmI4IwiszUDCHEFQXm+Ic+8iGM5gxEVDjbkRPK+XQ73pXPjyA
n47f8oxEAjwktpw+HtPiKGD9rtQ1Pe9Q96jHG0U7Y3YLuIEyibpjxJMvXvCU8Kzo
FZkX2dAXZLKIvPPWcrIQMm84I5vBS1FWpeRWRH1rGDy3l8W/gD2ow4AXy6wdqX0f
FRrCfgVloqWp5a8drBZJXyqEBLhbsHEkjxzgCiTF2x1DqZuOoqHoRepHanHIuVz/
smD21MXkxE8JNwD1Pm66fZIsF//zdB/gVW75uSoxnJf19z1eFZV/3z5ZPfw9lo/7
XBWPZ19Dec0ViwFN6JFZjcTT3GV31zPQjzN1FhngU5x6IexO0ByvfudN6yv+N3cs
+uv0BXeFDDimsWo4+cBkHPqS9blzYeMp/R2uzUSxX1E4tXOdzJfU5WPb983f90hl
ohW3ob8ysg499QCZvLGmczRfSHh+1H0xB93YFWtg2e7JCcQdhBk5uiEVWI7KLe96
0OwWlH8oWUG4uuikRRUNiJnS8SbA78D8iFtJtVoHwxlxUH1sKNjaI1qHwkdNbKJp
ZkMLHbY2XWgst5V6Csnz1BNIb9ky88opxVNPYMuvutuPJH0g0msz/Rt0VWuyiutE
UeAnOqdD5S/CeBETBekm+nvmEe9zP63BDUnKib7cANIeOBvawtv9kVl0MPW+98a0
zzOAaR/jzf8LvbgmkTwSb84zIBQmHreOR7weKlSqNSb5ADXmSRiinBxPaIrUglP/
dV74kKzsbT5qa400MDShvv3CmWQfL1MlezZC65IyLARFgHogsTlKac7TzXJKzKvq
A9a7e7LP8sFzJ6buYFRKfEfloDuhAABjkQhijQAtLH6YxfTAkIFvtxz43fMUtQyD
xjiW3NHphMBIpc6gz4da40Llv95ZT+2toX4nHG6030R+Ybz1z1rZLimfORezGPoS
0a47Ho/W39GaOI4lZqoxtEIL0Vbuzr+YO8zc/QLiexoAVaHIjGpL35pac0nfknbK
pOk+Yaz2uvENVjj9CnRBid2uhLrhi+WkSPhT/H0grRaZh03u/5HM4J+v4rsJnATj
CPIkuzFvSltDNZPIWISQB4GZp+ku7DY9L2zj6qX1C8wf4n/IE2Nxn3yEDpO4O8MY
zMJcMwoTjnEdyrnMdUbniP6lcZJwOMRAry0Q45tGCRGgQbOwfar9JGSinPjAnMfC
0pNj3cxc4aCO+o84ch4OmKPC1iq8lMkrC0lqJUGQ+U2NcgLaD7mAdcjSX8Sbg2Jj
ZWp37ORhAlYmcbr8z4XDIEzn6dTUbtJFBt0/nKeb2+1ONbaxDTAdqqE5zF/sYfHF
edhV9SCf5sfszjl/ZaUQkA6NzbXFBPqqzyyU5hbP9a0TBUt1M3nov3lFwFP6efw3
VKzwxMfBcoXCp0elhV49EQWXpaZ75YUfq8BoleUuOujUVYB7zSMxGPbqAtralRjH
GjUlrzbDvb2DKeiCZhpK+yrAV/fAGjE8exa1O3nIIejq1Gd4/coUL6XJOtdJmkdt
t7h/FA4SAvkQuMb318UYBBnuRRfU2SS3WHnnNlPcDm1HV4uVI5TlEOU2NoDEOlbE
dTTl5qEEzDditcPA4J3g+mreuAqrtCEa/wPOgpal+mRLJQjqU7e+b1BIytE0Up0o
K42p9tOzPjVT3tBDIGy+Gqm5hz7rVZRKrTAaqIh9n8+h/zv4kPB4sQuPly20SowC
V6/EXlV3Jpmn/JYMhRcIvUj8o++FA4OoDu0VWHvuqbXDwF5ZZpGH1Mfr27qyEQEO
HgiXFdaohF8Gpn7LRY9yNjhou9bZ2ZcMO8jTxl8CIGB9r75hvFAyUAMTR8c0g0Iv
XOYx679nl4r6HjYydUliXiYZXpDP7UIVYVkJbBIgxr96bo9UWu/4Bq3f7WjKYL6m
mEZ5/d/P1mmxLnRI+TA54a8nC6JlP+dVheQb9/sYkSZM2L+ByjhHCFaZD8TCWXc5
Tu3hr/G4PECeavBVd0fZ8SfvU9ZGM9P1gAMPVchp9kJFlDRNkUycX9oQ2K/XXAwK
KfW7rl+KQZp1c19oU9zUQzeIlxoi3ZO9tyHOrgimMBN1hCWlY53W82buZTPobSry
zm/A6s2HkZ2a6d79W3w6sGdhxCG24BMWW+7twb+peSZgYmOKlvoTe3f5SwEAdg0f
x+3DCbAlInkNoXgvkVMRHIfjJZRl76pBqr3rrNNIA0U2kE25UeoXKQ5KSXrGBER3
oTaV2M1NwAaiNyAfLUaaDFdKBRYdSi1PJV/9yAzaFSbfG/u+I5KmDgdPOPTCxQeZ
/EalmvMdIVSKGl1OFd82EAR6a8C+a6fa3aKeYLnExyYG0EQ6ly9X93sZ8GM/OIcg
qhtJgoudJoVI+rVwRpH1KUoGPTI+HCTQIoO4MiK1grw7QA9mR25Md4fq0J1YOJWt
AA6FdTVxhA+nmAJjPOSkihoF/Y5iGawxqdVIDKRdU3bSidEWWazkKrT2wJgF+UJl
bFmwnam7FVa9hRyg7Z+lSZrWcGsWJXWlantJgV35Z6k+wbC6RODLlnfuRo6cJc2Q
nv6RId+MVYFioFnkPeIDJTnG59qANezFQ3jWGiRuoPLRiOCOcErQjcYHr6tdpbXo
bRiMiP+D3ShiT+z5k9VfLv58FZ1xcn27YunmiEp6iF+dsXuRfKb2lLDjxD6V8ThH
1Dc4ikCs8feWBmV6BAQnZTqy81yDeqsx/vzbzXFGYwiLzOj+9H6dEAJp0LZ22zR1
UX/lvzJWhZwgRtXZAk4HMWtmsYSr4+GVWFqkNp61MGmK9MeRIYEy07ECfvaEq79z
wDb64ZVWLpAqlDDXcTOBWVNuye3E/DWITV18RPrQQvnbXxzTClvV9WuMGToBZ6es
9FSV/wK/RZFaWUn5gDdzYr+rhMrHTcei18xoNlISQIKO2fCXlECQ/RZhnzKeCuNn
L+prE/r026sEcef4U7b/9MWjkYv3iXYN8WMPkLHnMtII1Jq1saOe6GGOlBhYGPJ0
nL5fYJhIIA3ESbYMiFhuUQG7M1HNsWMuLLvoZYgKi9KY8XL43qRp+UIXki5MNg+2
ZRvYhAAhqDppOuKLLC1/rHUIFnRn6j4TJfbnFr6u0m4iJMFP4sBCBDP+PMbxPV52
52c2X2P4ZSkoHl86+0iRq4XAFyu+RCDq7GnvGwCX1oqeLKvzYMtoPzcGzwXI6KUD
a7un26KdE7wcsGRaYNQHGBMf+wYy0Hj7aJqTZoUCRvIByG2S9sbRHuTiYGzOfjLF
Wy+1yGFEDXgPsIOYwEzWzlTMFBuVzgtSKMyL7zTfEslAsEYHJMdvS1+8lACsE6//
ZiXZZjSOT9uTH9UXBzyUxADVZzIIiivgJHKdhAU7Zdw77zBAA1ni4bqg9yiHZKiw
Xfuo23UO1tAruHJo7TQW9fnyzPfTvwzlrUpSxHfCGiOIObH4N7lqUEbGRMv95Dtg
eaKe+li8VJEOPBb+8dIJQ7JD/5seoUTCaUJM83lmx7zt25HFLCmAef3yEX0GTL5O
maMXMCi0PH12grXbrXgt/7U0JdSnkMEjbjNVeOeanbkefpQw1V7LL10rH1oma+Dp
3na3YGxCfqGP/1kSxxpc20rqhvOg78kOuXsf8hi3SILfO/nyxboEScvq8yoD20A1
BBvKgnvmS11qwXSze8idnIVvlCKDKuwuz1YsE2y6Ajk2kH+3ZNYrjEZxOz9evKMo
10phVA00u/p0OXJRSr8fduNQOya2hnAXn2TDdLsc+KmgsWETQ+IMyOOV0+ilrGxo
VVnHKNblcUbYhIx0H8Y7Sp7wFy/lVwYT5c4G2EBd9lXCagDHPY59HZtASGdpA2LI
3+uWMXKOq6SfAsKCMNJvPpfoOHXIGcUE51rd1rn/DhSSOTPV2VSF+hazd5TjRpDZ
bmEhvmLiYDLnFaXukiZfN6JrMqf32m1BABCH0Q7ZfwxzTSq/evkp6x13b70IX9nH
OWRVFHgZXSEmYdbfI11934/2igSZazOVOqadBZH8bO8zFHIVSb8XEj6N3NdiTauG
697q8OoKArqwf3YJdEc31MLyr0FLx5iaw03hG7+ALPDNje/ArLRvyHEfEg3JVm0Y
/71Fv31/OziF+d+QWut4D/podvpHvWRIZcZlr8J4TJGUaZHgGymdMy0ObYjDuzii
Bg3HmRRYoFPczAeGROFlO2oJHFUVj0NOviPLkvxW1bSYcG4UaLL4ObnZjzTC9alz
u64EDfOYELX2uizwM6lijekd6KWkly3OS1ZmJyk0om4tzKFYbpQ5ZtvKNLJxU1zf
qLWpqIJHxc2WqKGAEZN+UlfaP/xuaX+vnwxlx3iIpYmOKB1Norn5Q5AqgofbgBct
x522/CQLFhwv4ciVJr+Frqbq+oBUeSXK9SGybW6Z9bmW1b6fyT+xQc88w3smvC9W
Pg/DSczBuOBNk8BY4arH7A8k+bKwtQ2sZ1k9rS9gxbwr1rU123eEKl+SOHny1TF1
mmh2ZqVLteKCjWwVlDoAAgRu2X2WXFjdbvxhG1jv4G1dSL9QSf9cduClFYin/ANH
B2Iomkxs1q6OWt2ndxpvuIvViCNvfy3yw17TUyObcEB/G2/PtPAYau8zUtsYWh7E
2leBglRBajrXAROVsJ6zyhUAFsFSDwwtAah42EmfoZ9FnDAkCGcQaecxjbiKS//a
QXoQFi25dFuK3YAx61wMkg5CG9eaQmvnjOK7NXJJshIzLKd2fIFWLZpcbrG7tKq0
+HXTRmbpiGiYImXSOrPW8hOjWUkwinJYIKhKquKJVO4XN8SCJp53U1RLy1Z/iEwa
PsoLZG1IDJEgGrG/cKm9j8g+Uf8Q9L8opm3JmFAsV188Q7iFChCLUUjgkIbC1Q3V
NadmzAI6blaeS6wP5wg+qOZrLEDIxvrq3TSHQ38STNa19r03aLmSDlLoGwuTVgA6
XzoQGro6P50Yuksz2SsKc0xa7hN2mX/ewaK4XHvwW1+kOLjK9m8NLXzZgs9Q3dha
ww/XXfK5Brotuz5Cz8CLqU4VojFLv+uyQV3CahTPQfI43vhTrrGbM5PzGoLw71wT
D/J1SnXcw9yl+NE1dxBGdo90t1qActRRRNx2r2KUZuvSiZPjWzsoHHglsyFJ+BaA
iiHb50tNk0aKaQvqLlm/wpIoAhUICkR2OSazjP62wKQuXxHVItEh7u1DsnttDqBf
SgR98Bwi0RnEbZRBuRcBwaXAP+n86tZBeLw1E7w5xEMRX7tuGVfrt+t5H5Ful5rZ
7IY0F3myywWkkbJwPg8sE20x0K7Kax28C2oXcvewyO0O4Ka8cFVuin+TbFBh+Epq
pKYawhnmV9KVUOu+Ul3t6r5opXt7XMELj8Lms3m9T7b2S0hJl4QRz2XkbhYqNKnW
gOxgCs1PX8m+m7nUg9uBn2d6dENqqkpPjRxe3U/kiaDCE2t5P+1V2spLNtSNu8lS
RJfvF9sxAt2MBD1jcx8r5zrr2ztYD5UZKHNF43D17hNYreI60O3HB4CfFbAAP1rz
olgXhq+aSNCUc06NWJ7LNKorvEBdetwfjL1YXab/6a4HiyhMViAm6Ndo5UZwfj1R
1XEa29CzHYZ6Qk1PdJRf50dBzwaomZ1xMkJD9az+05dJHEkftf9ni6VYRNNhpNF8
q4TfSfjEAMH8cdW/Fqa4rqMToVbYA8k1DUAcuJyjU89Jk6KrQ8PvfPIOrKSsBUbm
zRciPPMU9LqWQV+uqV5w1Rx4b773DqBQxnrfZpGX0QbVjnAdfFiKbFFvqoLilI8Y
tTijVQH6Vb+uWdpWffTryxdWWvoMOortHYN8YvYi1+fLZkrOhJwexaFS/rcBAKfY
3mVz5sAHiOV7tPP7TKe9WWN3mrc0otiWXBj7Tpx2F57HfeHDEiY+B0fDMESLMzq+
4tWcX6ZQDLlZpyr80mVQgIbkzH86imbH+gUVgOVMf3uxziVhQ3mntsisHoGl44gp
f3oH9lZQm5dfftyMHUUY6U4dDqzpwHFEOp0kKZxiCU9c4KgCajO+f1d+6pp7IR0o
QBSuFxBiiI+cmFbffj5Ceaad9TLbb16koZ1kkYD3cVDrIjkZfLpzpDKL+eEMUR5S
QxeVP8guMTZQBhuoOHKltgLJWx86Z+YpSoBUdy7p1FWw8v99QeN+io7Gz8mHbKvb
REy3NxE1oWdt5eWxb5JO9J7WWHYhtg9mJwlJtB5tVCkaBf3hm4BNTgNqHuyZ3r2b
saC9TjqnJRu1hEqV8ejNdOi4bEcNbazCUIV7C34KtDsNo1yC/QTpGOwz0m1Y+Gmc
iXtvYgc9arXaEmEEps0mgAcmma/A6FPAV8rWUK0xb78GbRIq6im8WHoaj8JV8fIU
tt2LQbfYPM2tOfx4TsfUcYG7ayZbGNUu/7qqYOB5oBTvtFekeNuqNLOr1tXYy2N4
GZpkjWF7lC4QiqUAUmqlb7UzodmC7hp/+y6ej0zx5SB7mWFRkCuJUTb3Hf3gUJKe
o64U0oriIo1m6NCgjNDW9eziNEocB+RyWNHS53oVqPvTWhlSUfKOaI6DEJspoSoh
0IYlP+58nP7Zorcr+XmLn3IWSkWjtYxOhGKCe4KO0sl3njS/u3xUruUMfQylRlTB
l5wbU1OWM+us8LluQtROzXoNLEofKRxnJU8BVxk86OLGGc0KjaNMZjqVxbV0IMPU
i55S9rQULXb6QJsjQ8iUM/gEDUf8ToScDaV/Ykir3e9PlTO/dsaF0oWeDzdshR8w
oX4aNpo/60cB2xQTVelhUBvVC8GxQY1kmR9Nh6aq1uX+kLl0eVBRiJQ7IedoTSJa
ctSFWWZE/jOETrPs8g+DD7ffNE9w7HR5/5TUIc1sL9wj7QKMwtT36l9r3TYGUg6H
3WjZ4WH4X31WmPlbPyM0a9+e6L2EWBFPI5YT3rTwXrdN0GbKKjmjlVU3AEcJJkZs
9M1P27mNEts9uEhX2007iX+8SQjc2xNntWUE+jwSib76ToD2HUKmFBNHF7Zr620x
sVf3DNmDEOnRpJAvRDfdpL01HZ8gNtN2m7h9YtdrI32pEboSUM+i10uFBGFNxZB7
Z1MDjC32dJLX8isl6NgsyDS5r4xcnVPMfGh5xMjhtXg0+vRGA8QC2CVhXUwEjKbv
cf+SwrFZ2X5YXJ2Rii7PeCMTSwW6uhlqumAnkt9ZQ7l/HumRkkkeHQjGyI4qQg5f
Io1ujHkUk5j09j6Y46VlI7pbgbKujV68XwLqnsmUna0=
`protect END_PROTECTED
