`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qJL6gTBv2Eo1IJnD9F1auCgWInHlcjSQk5MAQEFXAXrV5vTqh0IXbyPzZbCbju5V
r4G5tAdfnxiqagOATGZgt5lLjrpiMXyN3a3SYhPTtkAiuER1RsSmR3JuY0+EHmeC
FHYIThsZzkdnn7wAV6EXzlg+MXtf2BlQeIjtovlAv5e88Or2+orqU2fglCw3DQJY
ztKxt5opkPVZ66E/F8dTpDAeOT05Y3MbjBsXQeAgzZnPz7HDH7IVPqD2Hl2Io1Pv
+pQtp7r4lD3Tb7MkQ99w5lUo4ZKUbtC8sbrxbxbUzKt0Z+6vWxx/aOPMjTy8ujEN
i4VqPKrZd8D9wMLh8TltYyhFDEiYSfhZfCX1d3KPhu3j1opyXsgVw8BZJ0jOYpv1
vsgrbMK1/jlmPI0ei3/0xbFmSsmKsKgFiGiGp3d0+cz72zcO8EguaOOT5jhMBsZ4
CfCXRyy6m/x6fWBQbwvLeBjREVJArr5C6a9K0NKLeG5Ioi4kmj65ODreIycb0Go7
ONghEqlnr5Ds7yTF0A5UTAGt+gLWrP2HgOlWOvEWUY2+lpwbDnhBBgQ5TqZmx1f3
hmvFYuQH82fzklMOHwKdIDOrouEODVb8clONL5vlcSmqA1cpaKWqEZwwOHhEUMp1
2DG44/6Pr69tuOEp2JNbDpvO5jaa2oTubMU0Y/qSGxfQUWIJVIOJMLYFmtkX4bC0
d35Rs1BIDzjM57JYe/Hea0oZxavDb4jl4X9kSzOvWVxwJUoHrFHqAh1BxpNCLsik
d3qGM3oQrFXbffEDMo/zJNT/oCOGUVR8FwPvkKK07hL0ENLtRmEd6LuIKa+eY5lG
Rq2keCp1TddXcWuN3SFHzakQ/H/Zrg6l8/AylsRh1qFnqhElfggDdSlVRbvB6ybd
FQ0htWipcoTHuuBhR+bHeBVuHKjkvExpLcPh7yD9+gb2+8xmjXohlPm+p5KUk3rg
P9hMOATuN0QoAKpTfXpxsdDl3nvieUaS5+a7C3ceiu8bvhkPvlzLelGxybM6a+7M
/MPenkR7ZVkN3fEo6CGGViIEGINXkZD1FlQLK8KDiRVoVOIX+ugUedBAMmJesU1C
OOCLIz8FdOKOCX0Qbv2FWY7oqfYd7YHOingSQimztLrcEWAhWfSXG0WMY+yRhZB8
QS4ukaqYNdmWgXFsPylGjRhYZDYntfrHeutIMdRK7oAG4jpK4IFXNZAb1Z1BN2jI
jtiAZqtwDZUkgEW6T11/N7RYJyr1buUn7s3BXZ6qxXW+QKVndbIKmnb/OC1lRueN
rc2RvnYdnf3xeZamIBzPtiYUVRzrMKYdfAVL8aH8RDTaVjlbBmTFkaTiKdbEmOH4
2JdrFBJlZB2CuyP7C3WPOqGlA0mXqiGRPdBPdSKGlVVhYcBB8Lt+psSZImDpWtVP
EGcZgO8Igmsu/qfffIw9qw==
`protect END_PROTECTED
