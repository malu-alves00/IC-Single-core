`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ydaqvXHZBgNp9bEwWyVMKN6nsy/etxLlZzVGYpSFonnk6fRa009mLPNdl8sMClpo
ODTz4PQsQW9i3yvhYM74b6MCkQIexjH6tRK20QuEbBxnQiEShYDM28jMuAt6V+Wz
BVOSZWGMpihN73mrZWWLkpKdGjJ+cOKKWxJDAcZyRvyy+X0XVLbiLAA+UBGDY6Xu
F4UJS75oyAHtaU2M+z7mU/akggwfUROtS3K4na5RXiu4cXyqbRja6JME5edrSBBL
MKsYPczmPl7KFuss3tnofgF7vfZs+LE/R7vyhavg28DM6tCLhjsr3H98QR9iN7UA
sEY/eQuVzvZdiu2InZThrGvXxxAd2b/BhpKiVS5+5BR6NJ+FTVD2zVN23MO/96eo
9arNhqKSHPK9sH3HL5FXjP24V8kabMaMdbT9O9XlD/7XQYwb1nxLkBIlIedptRMe
K188NpSX9WoD5KDH4FkTs64HwSQIUCDNvkXl3PhdyEvSDnbI81SZdbP1fuLM8RJs
8Twhhi57BT/xEiaMUSs+vfIFVhOTJv8kHX1wXECuzMc2FV5vYjkjjc3vQI7N9syh
rTrhCf37zqXmN25YjglTxnCYgWKSbCAAt6LeM5Pqv1hbbY+nAh3yq5A/SCWd5FQz
i5gQJHe06Ozn1d1dxoLMNDXeyHCvwdOm8yKoIFpOUJyXVAYje8/AR7FtnSQB6kGL
aV4QQCtLuNEuKCfJRk+20TgIIrKoTIDxkuLgjxr/UKTd3NOcxCaiv/0rjkD5tL7t
IK0m2241xd8lsCLGfx+7e+tv3REUJQg2jdTioVfLNIPZuiUxKv6HzvYnQ9PkROml
pflTw49PvHJXP5HV9r+NUtHvCq6XzHMiJjZDY/Qb5+wghZnfT3qDGGYYsmXIogMZ
WEyj4s2BtwU1mQIjog8QCaSSOBjlIt0OdPlofJ9eQw/dx0zpCaSBUFIQivkjggh3
XJOo/fqEBNLomEsBisx4mDWRdjKK+LX2w1Nz+M/9sUMjPd1Z+kl4EIP1puurStNg
OQlxaIxVXiZcQhwuh9XCwMppcj7gEvX7V8alD0u2CjNHQnMVT9Mpv/QERL+JKrii
`protect END_PROTECTED
