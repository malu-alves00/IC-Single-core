`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kjDcHwC1k/LvPl9MSpBi26PpdpuLbPk6Il9djBN+O0RCFmUWVYdqyB1bHwELzU1a
444DE6fViPvNxDIgCKlL7KQE3fnXhY+hN427cI6DOBzZi4VoQujUE4/AwHq2+jhr
M3Cgxu5gkp3thEQaVAv7aM5bKLUivdTcZENG43GpvNuN+UifAVrtJKu2aLKKeuBO
IbpE0xhVI14/9o9CswO5nM8LabOLXZfP7BoVVhIeAsmOBNphY/4CzhhAAkxLbH7o
8h+rrI6D9Vc9W57UQFzw4F+JZhUG5iPZdHw+Eg0b1S/ChchybHST24eVlnLCfC3O
gqR050Df+WbVscn3b9ITxa0SZrQ/e0XNOxPUK38vPkcfe6488PseiXhjLOSZLG8b
cdB6UdHsds1XoJGJu19X/+9AebY7i/zgKDxAHSGyhzvrDUIMg2n48KDigILVx1nh
3rBUGsQSJWE8czaPs8LCTqKGiCN34ilFhzO6mTDnIHrbR231FNvBd7m2LGYXJVV1
vE3E6IGhZOvt9Z52A76j5ez14kR0QHaVXn2tCfnaKyMLsMBtjD5+v2h4QpcNMGiH
t1SCQ5nt2Ixoyj8J+EQrYQv08SvniOKfDU/VhR95dApY60Q7ap17DecVB1GQ6dYt
piWW7oS3jQQ1lIopw+q3kQJLTApKMM4nVXcHk6+8CthPIgSQLSOUyQJbLSEyu6SI
ECisJgn1xkLCx221bYpV+Zard16bSDncF9ivSz1LDReVM6zzYSHuiUlMn73fR/NM
60MlFyLG/0M2twbjdKAOg1EL32CGdzc4PdNQjaCTR6rFgEao5U/f37E7Ik1YKOWW
+vjAf1xtxlK5SxvsKjOKk8V512QcltRgaOqST1lG9eUb9ZIP3qB3xdOCFQtQC4Dg
NbRRQe33nr7IiOONd21XAE25ibkPQTlTA5uWIaz7EUsq5Ir/duHHP4+DZNAerU0L
+F39oqGFoerd14lS0y0bSyfmdfZ49KFRMPrfXpYEVshlES5I5T4tat8lErlrDFti
3ZHeMLyonWOlfHrOBHIR4k0gagRM9snpvW5O9Lqhg356qnFE/2fRp0WR6yLbEq71
V+KFHnk8SJsovSyMzg2aGZqDMybAn423qJ/OS49uUp/zMd5aeP1RsA+695oawmqs
Ebld/E0ZomK+1Ij0YSdsJoD8xSuRZlKnmk4SjtDs1JLKYumoUatnnjWpK+SAgP+E
htRHlsn/lOloMqGarn0ol1M0XgcTqOrEGqhRdx9skCaEygt/qvyzAEQo2XJ8xJ9F
JXVvsnN12IEBV02mW4BVzzuopgD2vKOnCxO6iG2om6DoYlf5zN2WV7tx7sw7lCrM
yrYsQBWOmqtgaAdfHGW1Eo4tpzoh1sHn0aG6YiYovAFaVNFJT40jEAFgEZRRYxO8
5AjjCo4M7OUlfVsXEo/YUMUn361y2Ysw3nAoyLS9g/wYRPKmNK4mtT647u61R3iY
/LqY2AaNAXCTP7lu6glDaeRwGkkHjcYAeAl5thX5RiJSEDr4J53RJ84T8ujfUf1s
SFwscEOwggeq6m7wEkyd9ME3SQgAcL5uB+GZfRumJyKxwQslqwSrUirpl93AycnI
NwuV1R5Okt2LsqQPrSd306B+1UT6UUR1Xj4WH1pTJEyJFrX+Me+j3VhtTHLuOnl6
EcUNmur12FrZMsiJyhESvFmyZLq0Od5F/Jr2LAQ8jj5u6/JcmMTXtGxPlykMwFwp
8VAHstujUUQYSbZ2KBozz+2MWqZ/D98qCYvHKaWSlt0k506E+6JvBrGIqU3n1O+u
Um4o3i8RjTQ8fhpuC0bDmCDAuf894VyK1kNrd9Q/vdoRs8wHMMW2fvVj5N/RNcDl
LuJKe2az1WwmOWKNHwQNbkTn7Jz0oJ35/i6yjgK0R0CASerxdruMybs+yU+91Wmq
zARdhZJ5pEqTZO1PEBPKCUxdsfxpL7RH4gS4oL20tuPu8wUtq9yLiQbLdbty4wlJ
rkvtQWPEdULeUjwNT0cXwfMGWh1G5PgXO2tPO1Iu6HdAGZxATc9xOoBuJtObiJ8S
Do5LRotoKe23nJbl/e7wh3Gk6pHBoZkhPKH4yN6Cg6pp8puhSUT8YUMdrgVsp84x
jxljuTA7FCTEmiqVUM8ZgnwjbeT1WYxH9WcKrjfo6+7OR8W8PinufP5DI1hZRNUu
YcsVO9a7luAVXfCXHBEJ/h7f25S7BktNQtM/ajG5zYcCbF2Y5qBAmy7LbjvvZ1ue
OKmUi2HoXA0eCiC20DilNrRKxhUkfBIS+UZm9iRwhp6+Egv9n9N7/64l6SILsCDn
t1JPT7NhMTMg0EFE3apC+yZR3R53uO1/rfZ8JgQsi19+agZ8/83DGo6/O3nw7rBO
iMVXAQ4Rq3VpuYIkpApnRmQyVjd5wGczzvmjsjPd0oaEAm76AX0WxzenOiq68Fax
Xc1ASNKYbPJBeK89PMYykkdTaNvGdSTfqpycsAi3Q4pvViJLbHgGWG6z+U0/F4g7
boeiaAVbIzVlySXkfV5YsniIBTFRYiLZJsbvK8MUtfzW/E7byX18imlfH4L4JAwz
GRmWYwMDgPDi/GQb8LjbOaEzk8RiLlujynAlHF78td0v9Zm6cwy7vzMVPCNBFJhv
t5cKeiSqFlln5hSl3EkrJ6ltuctex0p7G5GJsI2Zvhwmz8cw3WWQBgEnWRBlaJ7w
WXr5FP2j6tsBL6iclHg3YGIW6sc/EjeFWa61IGe6YyuDIR/9020I9kQQyMMuN2Kj
Jbkv9DrXTbLlQch7lJkCeETDYXPgLw4Dge9sLjZv9cjrRbqklKUS7zjbaXORrqQ9
s7e2XbX8dOjLcTEJerlzpueKvatGqWFO9ssy68eMLGLDkzMegM35rcMSxiU4laK+
x4BYy3mM+4FrBAjMrcD6yiLvKV4STVqD2gRiSPAdq6qVhSSmPtr0KPCsdlY2is/q
IPHNLVGFDQxpFhQDSxkuolRxUvC1zxRKrDflrKMTab+fdjrzjleQmAoiIF4jrTQ9
phut7/Oa5BRM1z7hl+OJJnKjFlhEIqsUtYh/ERkr90QIzBLfPXVqyufY19E4xgbs
7bbXf5yFl7qG/Vq3reVLShmZpzvU1qkpBPEoNswg9vnVcoRSFDxtLvjBbExBx6Wq
fnNGr6iLgx+Sf7V5s3q8aBLQlIg1GVa5n62rrBA4tlq6twr37iD3sWN1gDW2SmXx
R4MajIS614I3ouHDKMyHq7DwOkpyGqvo8UstBMlQUmS/2KYvXIn53Q7AhTqMYFFa
FY22vHPzSu01m8gggbj92BT55YcacyrdxPwgRukDfeql7wgJWX1Da+0a5lrYiTpH
3OaraAnFzzmfDkeT7fIaff0gj8YZd78Aj7ECYU82MaX4u6WIG61coMjy/cvyh+Ic
+F3svIikHxLwyIROM6+X7099SaZ8S+b0HXAB0G8/g6I+jnirpfbuYlV96DXzxeOb
BW3riNmwEk507QBPTgoHQAWQp68bcVSWqQJpvOpvVrk1LCSeAAtLJvHFIP7tXXrE
/WC3yUwxNoPLYcmZct15f9+U4BLm3yzXbIXczMj7Q4hh4i31ZrQMBOkJbPYUBsRf
dI6bv6+HCUr9vJr0ChAG8pZO4ok5Ff5XqO5Ie4NV+bKh09ZUTLd5etWd0w4SqTst
BhuQJme1sPcmrAl9dmrRmHv8CNqXAMPi5uoXceqnBUpvKd4HTVjO89tl3S+vcPqd
4LXLdG3cLAGe85f/HGrVHGSO2pLyxsaMhK3jmGzhak0Pi5txcB1rFpUxL9Dowing
IKJGqvs2WYswYjOK0nrvzaCJ+VhWgbdZU56SdADF2piONihc7Ei3+t9AUt6FAEQY
ZaMTPY8wKgrMnHimSqJD9Frn3pQ7zOKLH6L/YXzN2F4AKn17Q5EHA4c/Q2CCl61U
btnDuVi5InUIXEz1+lmqAEIXz6q/XeajhtkfS7bIgWZOnSQ4Cr/pSK+re33xpgQQ
Un3nyKaCZQhvEJmCRG499NR2bcgE9UuGdWuDe6jqon5K8SDaFIWTdwC2nBXG+gTW
Hr0HSvl/8I0RPtrWbAINcRU8rTIeTc4CVJAzevs8XENZ3sxcE4e76bHBNiIuny70
b9DrzPrmfH62aYhf3cpJQUJ1pRLMc+8xJHnKbUqDWIBVsCAyjJ3iJu9X579i6M5J
7Ijajve6VChdVUOr6TY7rC932vskmY6G+awSsQQlrByhbPxsVeM/rzD3MHuI96i1
R50/AAi9Dw5suhvkh77wiORxI8Hy9ykTrRcn+DKchM5bLuiVIjCD+CUHA1YPmJe2
+11KxeUjDfuCKvYTm4kR8eARVkYA3IYfH/d2XvDNKqYo+Ym9ApeEmsRV/e8/vSNL
0mmCGBmNKITVsk3cxYR90KYuLOyLfgPHz5MwIhmPjMeHl+5mS4T6Oo03pYvW/jH2
5Hndc+pv2QYGnns55ltEPj3PCunsVmpPqf7BDwJ/7NYtrFUTOIg5xNrwqj/Hiudy
D0xABDMDWo0pQGnevmmHGbJow1qhbI4SCGhCsZR7XeL0SdqZZPdk7MwjLT9kqzVL
+7pe6XGqniQrSAiO85eZ/BeGbrNTS2rKEl2LqLngOIcCfvYQEHQAPirR8yJtV1WP
tBCKIBdvJjhmw7hiXl8d78d9lWx+ay3USSGfk/lJvDxWtIZtyOvhcLqPeT2eZPO/
ZWllr5KXbuE5alGenUPkhqYTCJn3oRubDlgpB4XHfdvRCD9xmvkzlTIbn6glxDaK
NejkTmctVPDkSarHhVkXmX3sWEOlZsOFi7kfARt3zlcOPauW14u9DCqK8ba0ZHFC
L6yRiUKi6pkJM8QFl1gVZ68YEZ70EUxFfCyISPuWDdOz0V5e9w2RK7z3ylrcPnh+
ayuRJQ8/mCmGFBEwTIV2nsKVYyDtHlWJEuxsOitd7QRI0JlndjbS7so4pgmPkp+A
qXGnxboinnz+QtbVCIT8rFYhS+z8a9OTV0SpmKfc+q7LVCFfbjHEf3FEb/nOp8fv
Pdzec0CcTsnPhmLmeDcAF9n0sFAssO1D2H4699R0HRpKghwWDkQVa1n+le6n/JJY
eptAbD9Ii68JA+6RtXOEaq5h6kI3x1qKNyci5BTIg2OXaDS5xNMcRdnvEWJU+LDm
mOLsElf2xMR4gbGiqNiz1LDNwnA0xq2kN1BuIs7niOomeHkoPDEtsSV+4jjMdS2k
/sJ7g7iWG/b/ZspmoM/yQ9eHpMysR8koXGyDqi3K1wG/PW3GTmSuDtwlnm5KiIll
yxjXfJrimSQTGx5CVBxEWmbGw1e+7Zcr1Abvbjt/BazuNxoibQ5+TlX0+GJT3sHb
YnfJB2ZtUJnAP2hhhvepf3xCFzoVDP4vBxANEGsVNEqwzseTiepE60XBV+6p0nu2
5CRVJ0kW72PZWZYSfXoOg5AiAMCDFmHV65GvcHfBY5TaVPBo/+K1F1/4Kt9c6q2o
VubNsFYqHALrAeouFnMa8QZzi9WcA6fUWRdgUbNTY8wN4WAyzdIizauyFaIxCd7n
uHEQw8Ls6nHt8HtObkQuX1LcaXWinSZXRdNCJptNLc3qitZoI+EkuIbMjF8u7fKr
MPb2fKTuqPFPzdwr7oA3r0+EkLwl02kD/eW4Y6VSUMvwMV3j7tfLV23toMmVZqNE
P/PAuLQ3Pz0p/wb0seVWjDKjYDCRFathx9oP3N5nxEu2ory079aFgE39V/0++rJi
IB2T9hlDr5Y+/Il7akxDfSbavMZxFU8rgoed21+s4Wgtjh98OCT4y7hxpnbJk0+o
S3kkJHxQefPJH2GcRTE5Z0ALYmab+KveJDSm3XQKI0snoz1lmpoTUXYj5tDuXuDD
I8BOfBtSCP7KzQROrv3CwxRKPrTWOnY0JdYFiPK2EIESN5I8qZWeVvwr22QOl9rU
GZKRLbq0hUINXxC4+R6QorW0j02H5u5DEPLIXVcROaJVHcdbKHKY2qHAD67qwbE6
F11PfTjnOpoGWsyQpDtTiOYROrwVjHVtoKwoZ9KLlQ70SPnk0PI3ZfVw4yqkXcgC
9rVVRGs9de4rannUrz8JM0wnlEJTCOe3B3IniPXk9UKtNtj4qBVWChANtPv10BCu
YmaP3/SArZDAt/Z58NqGXKr6ghjNs3U7yhY5HEQjssv2ue3DGQBdqokh1Gu7+upQ
uoRxYNFSOMz7BQir4E/tMXnrCg+pYTp1jk/9rDOsfQhBmeS6VG32UITmpnOR3qOc
ym/F7vrMXUUcIcxhSsHBNTaaLibGy+uxniefLeQgU2Z2f0HqrpOAIGIxUIJkYCO/
T0+N01w6dVvXWZs/5ruNXGdTXFPD+1uk27r/Ou6Ukz2OkimPd6rhpt06ogdp7QqG
DezkpX7s/ZLd+b7YFuU5kbyzjK1gOYVBKXgRye5e/qw0/j+ll5TzBEjeeVS/gk2t
iLsiIqYiiNwvczdXclKCC2QUEOnmPoVnrfmmexgtFTFraZwb40gUx2uIkvb1cuS/
ND1pw4DgR7Pvmor+JrH8QPiwOivDRnt2O/K4AgvkCk+GL+WEO7k/DF3k1KPxbAEt
KBBhB8nabdAvpoNj8XY/jy2EdwePVfERAPByVtJWFgnsZf20sXToeG8wKvAYiiiB
uDiVjH+Aqz1ALwl0zalbdJpKmA7S5Vm021PHFR1L5qwltIDmzoxgCFvqJsVVbss9
3OxURPLBnXMGswuh7SavvpuhgnNue0M5L9U36lP7rSz4jey7VePoHFjZ7xgst4Tl
KOaxVsEX3gD2ijnWMaJd8/Wuey5uHLiNprKqgflXZuRJ2LBm4YZeQ7mxgwE+h3Lh
fRQKmGUqV12aOv18DWbg4YWuU0XIihsNmojP3tpIZlUwfrmGKHuyObdZk9zTjtBj
j440kxIxXNQF/A+TZoJPsWxBbcZ2OZWjU8InJeRbIINSDTM61NEp6oqOquI49V8J
zig37CZSgBXhKUwg9GcKpflEBaP52aIhqQI86wZKF0zQMLrI1QpfruleIZ+Glwah
wGzh1qFquk8aeOywpV+7xLqBdUweUZ3FIbqiFy4i3A4JDgtDajRUYkGzuMMBsUs4
51NYcNEW0YdHsMdB2UPPWCIUIwWE+1+7LHGOam8n9bxgxatEIgWdYrIdKePmZJJx
SGQsdpf/lrgnIhUEAJSPyi5uC695L4GRAkap5XgOO6FaEHrPKjwhNkrjkdJjXDnx
Pt9a0+jYSoT+Yz9XMS9ylPVCHfXyJKj5GvKd/V1asNOK/TVHYS6AuA1KcIk8icj2
DLv7mPhPGv97soE2hH60p77qjjWOJOmSnuV1GFg1OhCmqUgQY5Stpf4Pi/rE7FAb
U2zC7hRRQZBcQ315dIAu5cg5GeX/pWHRp8WHB9FzYVPxkodxf+drFWpXQiHLNl8W
sLgFGQ9o36FA5xfOZfRiCIpByvcsoY094yswz2IidrHDeGT/MTu0IzS7aszlgEqh
v1Iow6rw6RzHI+aiCJ/l3qq936ZrKbKt2/H3qSTzOsPCsKQcyG/SvujH0t/3iUXN
hbrM4aplPjKN+70D7c5V/Yg71pbFsnT5VK36G665U8+VqC8CgaTBjeE6laq+r3aU
oTllrGisV1UmSJl416lqSYaYRagEN0kiAd5dXIVo7W7htiFazLhvWAAgd4BQcNrN
0dn9vEjD53GpQKQUmo+C+dVADw2BrXhwbYqggkYOcaxtaAHOjk1rTYLXaCmwTTzA
toCXXR9PZNXaJtz+RY/uLiIUW1Kva6WGMf3j/hBm3cXKDGjcLWScFmUq34lJMXpy
2t5SUgeYhE4xwFZpwpCDBsmgTyKlQnJmNqfbUaZd2WyRoNA9zkUIQO4SXWvqF1N6
9mZ6/JiTo5KWINjW31dqKBjl6iNdR8JjbqQX4+oxvN8JQHAGvC645SUB/sMyiXnW
15y2ymaxdGmiMKsTR6iInOnDFhbTLhmTlqcXLrHTgdOxqtrW5Oy2vFdkNM8SjZ65
spXvL9hzEVJfdfZGrDhvxZm63Im9ZIBxtPR2t0xA6Vw34wyQoLaJemdoQSSq/Xm1
dy0j2mmeXW/0hDldnZvh47gJbUnuNvyL+qTc3HdxT3SytSsecG+GUpKwb8Rp+2Qx
2R/fVPVkpFEg2zZJH/aRSsgM1srORbGMJehQCZZHexVXlTJsm8U+fRnBg4JddnSl
rt5LdavxU5e7GJDM8STey/UoCsvct6iiaH3W1l/N1sruouSqAGsATaGDnnEuoPXd
WQt03N/bRpsj4Gg0XocP4x1HjWmadRYFwQul6H5cRJTeE+w5KD7X2H9kvMjW3sYp
nH0uNBsBtVx/s8IPK8h6kSnDNG3xNeQRXjou0Jnl34SO2I5r2vx29fXLPh7c8R2n
FDXDyW/MVwfg55XZo7hikp+vPT+Z+qAtF8o86R4LwFHmFXVQpmOdTCGyTObCr07P
0kbs9a8yDr3oDHLJBeAB7lj/Zk9SHsDIEdUvMooVavyzFMF9NtcceGdanCABYsRm
VLwPXxujXvfye5mOVWlvko+Vycge7Gnzx3p72BH3MQMbffNjeETf/KaB+RdNoRRj
DgpTvdPspHIPC6ct/J5jtslxC27lUerjJ+dQ5ajia42nqQh5fJNRaOw+n3LJqZID
AV+NRhv4wdcvWwq6nIcVAKJJUlrXSk3RHA+axumIH3vgswCoXOu1AUgglydmJ6SE
wJW3wppTud8ZTkLYAoqRwrB3E+t5y+KZLqBb545z7aR6CVsqRtPuusyNHL47NB9v
MhK15Kdo2uiP10FkySp6FFVZLqSlm2TDQ0EyvrOeKvQaxtgPoeG0Fb0mUuR37s1w
3V+x3AKb0seMytZuQg0BS3NOFuZRl1BGe6xCQb+2gnClBE9qHXBUCUjGyGmF1Xss
Ll2niZ89LEtnM0/8+mEwv0b3jX7s440jcxqL1d6TVXaPxMG4C8b4ohkppZHKGKxD
mKo3rxWBnnhhX1uKW5Wh+rSskq11Z5NHvSpQneceoSzuQroToig87DEFmyAfekkZ
l9CZM6NvTw9Bss6Mly0pRR9FJYJ1FWQIMzP2D6t3AYxjgTd7zs6G5ZZpkNVZbKrm
VHbe5qy1iw+nHJT5pfTZSYrENquVf7yB63RTTqBy8kfhNmvYyxx87qUQ54JIysey
bwyrH2EXtimiNyPXkNXZsBFlb9ZSe4sQ2XUxkfQv8D88wnT0fdCdgrtvZUhOhRm1
kgSX79qhxPHAgy1eBVJJriVlX5WEYkw/vO8DVJV+rKzZETa4feG4cfkqp/TuapOu
LZauo/Z0JCVK2WBLaBTnHuEbIiyFGHYdnGwJoSWU5WOOoj/VZVXfRIdpRnWnySJz
toR5EAm5+xYGZNMPsZbtGENPiS3ZoYaUA9/RL4g5irGbEPqMdZa5WvLxkK9CrRHP
Ub4NRpxeTgYDC5ettvNp4MXEvYJrzSkQzmqTLa3CdQjwvrE9j50oZwO4tQlwK3XA
UVqHXHVeqk+zPaCp+OJM9tg3wq4frWJhikl05ErALBoS+T5exwHXkhTuErxwfHGF
2VOUORUrf/ncLDGGlff4U5EMPq6TpCj7OktARv5rk2agixR6w0P+Ep2eNY77tCXT
is91B21AXDM7kP564AUrI1lCPAuFrNGMWSQVbXvS0ssB+9l/bOfFffqLa8AuSrCu
m0FLXv6XKdYtVfCO4+HfHf8EFono75YJSqOQ29+9IrOJNvD7L7VHkMUEI6uV6bU1
5DqAy1vP4BkxGSbWMrLgVak7cua2t+CfS7lp370Lo5dV24p94Rp0Gneypxlc/QWP
sNCqa3FKMuNj3sDLVFQerB/J0ttNS3QzSoTfGyYMyQR5D3L3IzwgsYGGxyVkoWE0
ykeXvtJ13RdQjEz/s7uv1mgaMHxwu9F5DCF9G4bLDqYn/8n8cB5gVJaLjwKZLRsG
zYnP7yHorH3P+uIiNQyy3iSdoMPZdK2ODB+JX+DgrLyoxqbA11OxpD4i3omM9+CP
cz5+q+09Ku6dmUnmKgQzz57STnhsLFZYtpQRps+YuKxSnWh4FdnnNGLTSymaKiu4
s55KHKsQQ1J+7t/VtrWpxBdvS537yxP9dRZZOBfzbBjuHjsoy7cvmNT5cyaniLth
4xbY5YmQcz+6Ux81ygb9Bf1q20JMGwlXt3n67OSPKGdzWs4zpn554ZgqOJ4UOiX7
CzEEc5ouAsC3uB2bCWtfMc1Wlcc8yM+UexTdLPFTuupKOEqcsCoXHDOxccYHwy2X
xmngbmFWKEM8mpVI8CYLKxrTavj7shJqG/M0yiEkmcnK2JcqV7Ch9/ogdU/Pwe2T
G6IEzjrP+IBf/WPP/5pHgjH5wK21JIY6ad6DtJ4qxiTZLx5S85VBPBxAEXcapnc0
Um03Wmi7//YfkBd+5Gob0S/Xg42P71cRM74AR4Mrt9wZD1GaSWE9xLZqh+k+xa+9
zJqg1cIi3RE007hOnMnUGq3KsaozD2YY1R3OFZq8g0DZiIsbSQAuoVbo5TygIt8t
q39GBwknEfQ1eUZU4IzfxZfMLS+k/Z+uzVp7NqmlCg3mnWePsNaQKQDq/RtXqT2/
CnKoojVe2a6fHt78xBwUHKWMdoTPg0wjp3vgHIYKSxsHqSkuC6WqqoK5WWU/9UcM
AFWReQg4BezbrsGX6ywKGwTEKFGmggt2gb67hDFK+9fwPh3Pj/BXH8LmP8wjzIXn
EDwAPstBIKX/xVX/Gnzv4Rb+ibJ2Hf5CK1IhiDXR5mESwV2n2Htc4FAPRt+fro12
Zl3m2uRWpq3pxWSbWPHMS1C8WLxVMkwr9oCA000bb+FB4tPGY9Z9wWbUBQcFUZRd
AaNSaezNyF3Qlv1/19oXAwDx/Pfc3FH1VmjNiTfS+gHhgFGnJqjDQ7EzLvySdJK8
BQp608sYyPWaWRHlMlViHi8iAZd6w3CH161k65mB1gSjqDbavrD99XYPF5QFJvOE
d4mAZea3AB92DaDFotfKAxGliiWU4LYXjrTgpFsMDpyGB0mV0AQx4bn5kVzPZUfA
RDBOgsSz4+bK8p1IUVF4GT2i3KTyRUueHKezXCCSDm9FXib3oHG1enPaGcXPGWeR
HemxB6/DAw7gqSYgPXNBF+kEiJcLFrtPOZH0yrhcQGwTE2L8hkW1zU1765ZUSUHq
QJOx2dZGi1QqzElWUB35bP38MkGkFY1UOFa8qhfLQb+F2OIekYU8llsrX12Q9qhl
y2D3EcUEpUxLgkj1gkqvnAEwR8SeVyOpCBNVgxy0kACnODbyOQB/yKigPN2D5Bbj
eHno5nyCbJZ1t51lQKCHY7g++Zsdr8Omnd9Q/vpoKSPpYOcvj9BmCMxolLiOp6rK
e5GUEphYcWi/OW45GU6feEgRpB0J29fLdWmDMwmFMRlbPrcTeceGq/eapjB6N8Jj
WBWjIn5n0oA3NWQ6ay24w8SxTPuNvfWHqKGl/rBYGwF6CRm2AhkLDro8EK/C0grc
QCCIAcFlMVkxaFBP0NBSSR/pnW+Tn4f4VxFVlbjVum2d2QO3KL4eBYtuRbE/AQ1W
XTRU/93vUhTCK2kGSmRRN7EgHZulJuzQUnj0YX+rXRLuagpBBnP9AmcNkiDAD1nj
qyDtW5fHGrLsCHmLWqRbo6Y4DUFFv2uXKj5q8uaKAfewjeiIGw2xqT03wTFtOjYN
K8Hc7BKCARkrpMrv/dX4i7EfXidh4OcJhp6Bao6h3K4ZSLXswVWlg5jVdmFvhN8w
zQGb2VSTtik4V7PpOJ6psOG01q4R12mQf6eYIHhyu5zw4I6cERi5GSNhpwUzciEh
TFWrN8HlAIOcxdOd4kP+oIAci2JThm5jpdQdFgB6Cu8xxW31DmXNEWdl8RxDTG+C
hgDOBly0kwAO6f8uLAENbqpa+NsHWW8Jet7vXf6k65W66um/I3u6+qvSn4M2CXEh
ten7XZ3LgLexqne2aIsUw+wJmnU4ZwIY4cXqzQ7/1N1D72WWGxnijWkyqDKqcuXb
l7zF//VYOf0QMVJb0e5/xA2CO7WVzZmif77CEV8YqKhL9Bj3sXwokcgrYwLDOpE+
3AW/6jSZpf3iEaKWEBdf+Ev4zVYIDkH22XhU/QKUTe3np8uEe2ihykA9wIH6nUKv
9AIG2KdPQWuAVf9kqMDhjlzz7bTNORyk7VxbBVycrs7x8NaFwDLDWXTMW1o2HVjb
PW6G5/QdbFNsjg2z7kSY1IYbOCgUmlLX6EB9BN+URV0Hn57e5a80ZgUza6i5vP8c
mXZgiPslTGqdyXB9kP5iajBK71ujLon4IUv+p1hNQMOurrvxLRflOCQzNM0QxFHA
Csxv8t515FPdPQhbcYFA/ZHCvXsKlbPuWaQApMqE4COzeBhZZSGu9eRM6j+ys6do
6+xpqTnrH2qFHci/FABrGFUyqNK11iTNO8Q19nTYaZcCmogdlVvNPm3iBvNULPf/
6I9+u2EaAH3W1xW57M4UPWZBsK1L2dz7+KtMeouB9sD82y70XjmV6iuDHUr3aXaP
EtAhpp3hAAYW4n5sDlUv3H1+DDKbOaPWiN8gLEkCtlJEdyX1H9d9Pq2yFw240Iqc
wlZu/bsiQ9F8oFYnjepua1TfdNAEoV0mQwGeM8LY4y3YIzGCvAhDSIlT1+QVdjmR
jrYyGAYBWpKQacicP9HOY83yBDb0yIRJWx8w+cHsQ+aZQH5HiIOWIaAggnG00oWz
SUSKeSsUD3eMqrSxB52nS4rLLtNgRvVwU6FeeOWWipdop7vjjCrKGahYKFQntuZB
w+5pTmByusvH8C+kDGWD0HsQBH+QskIsQ86ssVwl/9XC153LtN0/yu+Dh59Rpx2s
uy6P8l/m4PlC3esv74w/fNu5c9k/oXFyEGTLMdL8DihynYqK7WjuUrO8q7xGKUxS
v4pInXuYrdO2JjhRQlTtxHbLt5npEz5l3l1pLvkZAeSurHM6ZwoA1LylaQ29lYll
4qP76wdwbvmCT1n7ecwX0DBW132+PJPJsGx58gzGA09pbpIazxbo6suP8t0OL1Hg
VklO1EjW4F9a4u23YEK/nZOqpzsCf6zWwJLD5srvffSFaN0O/awpcVmsLerc5jt2
LKNiGCvvs7pvqhH+WRiMffDSj0XkCj8D3d0ob7Te7qdNewkHrPUzcN9+QPwRaN2m
ZcOWM5T5HaRAwewjZqoZLF9gbSMQvrlNRxTBonOBtCA0DdtRYYnp5rnXJd8uH90W
SN68aUiQKtdlzdjFFwuMjEQzhHIjdXg3D1oi5nptSsoQ8BmoMC04PV9jCdOudSqG
WgUbt1OfiVlpD+WSEhAZNdO2xsJXrmNSo7bE6hcvyBlfNVT2YBDklaY4VzHisu8a
TvODDOIGhR7ORTGcZF/Gz6DResUmF3xrINWTP1Jg3bw11Aeoe7dZOV1RpAelAV1m
jyJ714k6yRjhNCmJDlcJq+bmu2jBcd/3Pw7D11Vpa+C5Ou4moqPEzXvc1YHVYT9n
A02y6wULM60j+Dy+WJBFS+Rc2tRg7GiBzfE6d3KXuS+B54cQrciNEfdNRO69n61z
PFO701EjJibQXDBDgdwBOVM+mEwcX8zs3uxCB2SXILLMK0A4Xtqio4AMiwQybyQd
71psUpgP5vcoKMkzUTrEWzj4DUyIQMwzh7NjilFGl7gZQEpdIc2yWxhrJFkSfcN/
ZRIcvnH+vworml4IG2Bz0XUJX3Igz21wVH1RqeFUGbF9xQ824rALq8sGu7Uo+o9b
ld+WBcJKaqM5x+8RDoaGqyf5BtXDJ7J0lasoQq17cywfHZnGTmp8pnkvt/vThz93
3HnJ7k2jMMC7xdFOQYU38oNe3jEqzr0lmM0JNCw2MUchJpZG9auoVfdxnnWi4lM1
gakmkeJwEnueNXaXFLvtjQ1pTX9JLdFuW0OhkXcjXxxS0Wh7Tfo4M8jkJCf3ivza
hQTn92r/mcXYXnCeN3VMOG/TJoDWs2wLV+MLiDZpaWkohxLUu33bO/0oTomBWdZd
2ANgqpUgLe6KgBiGBqJqKy1zsgZdFQwmO//so3fNv3jRrS3h5xgI8tgP5Hv1rdND
3KsP47ZeUp54Qvm1uwCKj8bno8XbIh0EYZb9irWxZdgS9y3ov4OycYUGCBETyyW4
rsUhaOxXEMgZaoithLFn0cgpDDFvc+xmverwWxmvyorrPIWkE+7pV7pD+ZVEhAk9
wc+OlZOjLpxsOhznYBbTeekeVWtOt2NiQnyUp6SPLD8+NPxHB/O402CQqbzck/JT
Z2tMe2dew041KtLx/1jl0hEemcb30XrlfQSJa25XGdhD5G70/6IlF5xCRj7mG+sx
312zSenyMfHc8lNpa8Of8VcoCRnz7lMO5pTX+RSilXYrUYdyPn0AmnY0CMMCu8kk
tfJwjGHxbGVuM3yUdlpb070KepCU9yrT85HmtVNNHur90xmpGkh5a/YNPE+UuXHU
PuFfgPlRo2MuVDZ3ODg1p5qVJjri5l5EQhcFh0w85zKXGv3QbgDuEdcfGbhgoVDA
SNbi19Gpt/9UPrN/1EO1sErGj94gy4g7kQ/Ag67H05DqnlFoW0iFxxHAPFDPfqpt
A1iz4PolQLOXSANuq3plqYn08NRFRq9JYpWyHkjxOopqvsiQvbGrDQM9xY4dPZ7p
1g1HQ2011flBuutvqOwapn7W/FM+Vs6zBZPSjHDTu8nljdey9wNujL2QgsMXoFmt
0/6Q1xGv+tmiAvf+iV89K+Xe5VUzta2WdSZoUvpPvuBYhzMdHqOiTUz5jsNf/wy3
KvNLUQg95H8TSEND3f/pzlxL8ZGeBVA2N9XPUgER5/qrkWo8cKNzujLxtvPLnF3d
neaHUkwDGARmHeRuggE2Lt9jOX+6LeIHW8PdBHgamtAS6K1izkvi9ef17PJ2/fQN
ICLJIeK3e+s7LthXU6hg4QMzOnuOFUiSK0gcSXBG+LL0D44TRozv97SN3+qwUd7S
fWrfPR0kXoYwBTAwVrlodF7ww0SFEDjA8O8TRmvcfgxxBUaZBEWiesO0o5IQXu36
WNM7Mlbgtw15IEDk7D7XK2GBhnvg5E79JHsIeKB6hOreqLfxv6x0UIGjXET/ZveF
CucrG1xXDT1YPZxnyBgc+tflebyT6cTdJ2dDmrwLbLVQDnA8Tr299ncE33j2oI/B
vk/m2xpyvXR7+jC36/oFqkNQEaDxq9Wzr+SIYmEuhAL2j0T8/nyqybA87wn2LVvF
ZBkyytsPd4JDPTEB2P4E50SuXb+cIJNKUetXLUZlLRvTW1CSz1cugqbHtH5t2D5K
RM2HOXSpC55VT/Oa+AjV9Vq67Vn4yykzBn9FR67sDYkbrL7zC/2Dhq7TiZ6Pf8XP
e0sxcPZdB7IAoN1GIz/fGtwmNV27NC1tYRUq1es38O54Y5aTg0e5o0LoekfGqZMR
aIuuBTUA6Nt1QK64gA4Fj5hEpGE/2BESn8WMwqqq6u3DoQvIvEXJR0lXNC/Cv+S/
2eAsLDiCskSmNmpzYbJ4ACTLz8cWqJK891G76h5+dZ4vClWzUDtIKmvo5PVcVGEr
AuUUbpo7/VKouq75OPkVymlfpPxlMst3w2ZwLVs+S7U+Wuct/yNQU8ehOtrauL27
SnmW3YsGM0v6k+hRgbFxnvxPwGHc1h6p7OK4vbdWVORq0dMDit8pnDHivL87K8a+
ohY6A6eC0jVOoCz5oTKoHQ7Gg6iN0Ng/GgOK0r3EEKFqo1rI0mkdtV7c/eJI+kZC
9gZzHCmQ2yYsUKVPIBbqEw08TMZAtqQej2jZzwW0xefrl5fPz05BuLcT52eI17kn
KPMP+SyC5JsriZptYIGpR6xVjYt5OwnmakJteREvmIufKNy+82ZmwZqVWQsjkEix
ZAfahNvF/2uvcJmk4Y8dGnTjkCSR2RNR5cPDb+vCaCXELBuTfdivehSFPQRsSZOn
KodJgAlTyNlRxDy/CwHMQzg+zMcDvUrtc7eYEbeBRJBtcF73gRU6kYXJxfIE9vcq
jhGq0B9XITcIEv5csoedqB9NMOiLJW4AhPRKKB1Z5QNTzWPH5rRbtJkA4Y7gJVF2
BAd/RQDhUFeifHos+rxEo9luVQeVzNYEtwdB84U1wgkzSLBmxmgWj0qRkTtRZnZc
pAUzQrXNIblimZqIis5xAL7twTq3B66/nPNRWUQ3pNR+6EH8GFwlhyNgm8xSEqLY
u7SFALzEWlTmwcGX3OpOSE2jlJ383OiZ+KgMQNpWPgy7k2Zm9PholK0k5KP4lKr2
I1gnRHuZVgf+P4Awvi9HCzIheSBLGR1tvN06er3L/C+I9/GaAMpMVday3uV7hE32
6QO/XYl2OOOMPzYozVIJytti6uqhCn7tpjK5ZfIeLcq11WYRvIh7/azGcnv7sFpU
ptrlKf4/69tYyFFX1omAquxD2+vUk0TMEcFn5WpnYbMK1RWOj0aaM27lmZoxa91E
K0+Yus5Rk4BfvkHpTgOPghp2/IcfnJ19o1aWJkg5ks44EPgYK0hxsA5QsQXaIswf
jyjtQbn8m9LbuQ+XrL23h1KCDXLMbbUDmHm8uSONXV1tyLFEhBxRDsEsmEb7n5b4
WSiRoVAkSnAaSUAFORfA8HPpjF7QQvH5OxubSOJ7VXK4m9aJE/Y40sySKDO3qrwE
E1BlZ7vTMJ5DWx3joucJH32hUEsP8ymxps9xFwl7KCWEoAbEyMkct0I+71Sc4vPQ
aA46kSYH2Mep8+Nlif8VffJm/izU0tTBxvgVgYLBgyMJgz+Xql5myohNLlgyr+te
eUd+Lqf+3MgDsuxhb3U+hRTc22nX6lUXPaPEdDYdpuIxTCeE0WzQVsXjHuDxCikB
sA42bmTnwJ/kOs2sXVgeEsk4N+uj00v52iJiTpTdanE1ZftmkBppdI2T6p/+N/RX
76c4OnnP2QLYYpXQ+qNG6RnbHIT42fZ1b6Z00Ol+JpnKKuDvjcBZWHdki8o0aKpN
IZ4as7GOssIBEOXykZ+qjd51VzYSpzr+HilY4sjHEeDks7lk7IiU2Jb/Bu0aWu5q
P0yUdS0E0RekVyhINnzxVWQHxAsEezD2mxkMMuNOwLsGYKEgghhFfuXGzZhtiuMq
Sa5oxcHSumTu2VwGkhfROF+5m7d29fGpqKD7B5d/lRtaG9E6C8m/lRQg9W23t/tK
g+Y837/YqaPyacyowXx9IqozZzCbbVSv6Q9Z2I/Q7mIQgqPHXnBU63iVAwUp6av4
O6yAav3BwslFKVR+dVCtxrm2gJgFKAPan5NwK2sFpiwwVex/GMoplt1Sa9Xrq+f9
DgDJxS/ls4bM2g6caIgQW/OePHl3bLQvIHsTJAwcXqssjEJYHEHMDTKFR4U91dxv
ICIVgsjufahNRbt6lmTK7DqgPvRjdE8NPMQhdD0bjGcaeWuhO9kRvG1/ZvjLpa8/
6pvm0Og0QiD3El5BmwfORVLRNo5SZQAEA1WHlqOgqONXAwV5N0oA1UJeCJuz5lPv
2RWiZleSxvwt9wMh6m0x4G+1uedgDszSZKvLzE45cTFOfnGJjZLALiXfBEL6lhGS
EhK5BIoap4e1/4jB6Jv3QdPTNUXjIrQnUCE7+syLy7ff0ZZCylPRxKIQzR7+iOie
HrKGPw4xcg7jQyd33Rs1uv/8JyPEXwJJmgVQNYnufrXP0X9HDXQEbtd87YjB+UCt
7DtqGt6m7lMMUcI+eotg/r/Mj3FtI6YoXduxA9oZAfHenry6FGxRPAufQAKdXNye
EFzrIGkQN1SmYxS1Q7YRK1YHtMSnvrx3H/5gbfkre1HFBmMlImQe+LW8ZUUfSyhq
ZAOindayZyx5VWB7lKxZ679oJ4A0NF0uRinS2q+DxdVOE/hU6YC84TtWqnQS6uuw
W3/UA9oSa6VKIehq7me5uYnDcH4+wC2SRTTANOE4F3rvLWyOWCC4zK3NpUW2zksU
ilF4vB6F7fujHlhLTWFNn6aaVF6HHjQ9iDZoR4vnXMSUXRyYZysSUMlwwn405lTv
QHOLkqCZqvDGve5H0TbRJCc6Yl9LUy7VjavYzry7+kPgiqu18rO2SsrU2KJU/FWN
kj+ddxmSMUv1l9ZB9oMBjWQx71m3CLw63s8bgss0Q/+SM9h3JONmbfqR3cO4ATNq
k3zeM7CsT8uWn81Nxq9HP9s89IDMA9s9FnXzOdLs7dX6vvk5zW3ht8PZQ5x4vOWj
EDpco0RMDVpLlibq1cE++aZPo+vej0fdgWtmGENKneA8CXIJpxrqPIVwxZpPS/u6
poBpJ0TBqoHceQuoS7eClFegfeowvZQ48CjJk46Ay+b4WlmJL5n78FQiAhV6FaJ/
JrQJHKRApYRybUdIHL0Mm4gmWw32sjVxfeK8wljnuOd1V6/mYZZwmUe8F/ggq6P6
pG3MuPPgovufLAj27G6zmz8VROJd9k3WGUC2zOdPQJ5rit0jQVBR2fwJk0zNUFED
cezfKHnV//SW2WHsoddQHzqj1UqPXkh0DnzcWckfT0fBQtMX1qOm6CiYlIo9Gj4c
4emIjHwUpaXGjmf7S2NBwOzCFx9muOYJ8679B+tXvSX3Bxs/lcWowVuGDY/uYDMK
ls7YISWKGNmmOxTJUQNuFcV7YzPY+ebotwWRDudhvvzYSHE+3WaOxGGfmo+nnini
jw0Wi3KqDpnls5ZQG5JFfHbSEjBuKMBpHdJEGGhONiQp7qY3NK68JYwbKNH+pxYm
2ReTetCmDqeZSX1rfxuExy/A2s1W5c6JLvkAEaFByWS4lRHjwape3Gg8dPnE9Ww4
tLX6gxrOogGN4Jo1V2g/9xbEkABLL6LWmM0cPi+J4g1OZuTK+wdfLCuXmwLUP/37
e6Gl5fB7svZ8VacjeXHufqrDtjT8PWTA3qUCiPCKLSb+c1Lhofou9zaOLcs1mGNo
Eg9VwqcQzcBQFD8typfOoqQ5KE9TRw8qiK8eSSfPq0+kj6tByRXf6kI2irndmlSb
A7z95zEDi4X9FTWEN1aQMoirG6aDCeiog8dS+/Rhn2XK+7hGkTglt5nNRk+9CFm3
Z2nELKrwYMaHA1lwbUZm/OQFMEEqcCXB9vn9xPAK+DJalHuhq9KEoh4rM94wL8XZ
NP0EU/v3hx/AU1Jz0xCxv5SDU9MBO+UBjJRPABzq/pAgaLZEhYZF6YftpDXz4Gmv
+9yjF8wFZTNaIH1qTzwwDh3dKTa4Hytqr/nDYhkBKQ92RKSJhXJLpOwDc/ctvYxM
I4Fz/pZ+GPGaFBmMw60nd424Q5RgtRbWGp4S1xD62BqBGfU2rxtnqFn2DRnVF9Rn
uCqxJteb6j+za8XcHR3gLUG8T8nX6PcT117V2TisKoMLmtqci+q6soa4CFBtB9wV
cfAapv7R6wAbjeXrlauvZpL8Ubi2J2rBwRcyqozcue6qVoSbtOvhTmX7WyFjfubt
bMFbNQBgDVG3tPM0O70IM63SOdyEyxnIxJjVD/nDw8MiMhI5mRPAm5ndLFj+YUts
KfWaURIvrmFOQQvTgJDF4xtgpGbFDcHaYWVwQ62XqMcAu63QZ9F2IIKwb6EPwmOo
EQfr/sT5OADF25j9J+5vf3otgIiwOXKiV/6KN/B0mkSb1EHk6fhJxJlIEJKGGRcJ
JmA00fCQOcBzbjvPxHkIf/3kHXDPCPuKW6BDO+GcVvJiwJCxJul8BoeMFXksJb+C
jMfaHCHaHx7k01ys12DpFwWz5uKLs8bBghPU5ACEzT7075g1j3XX55q7lNZ1KZG+
GA+xMqV/t2ux31arNx3eDUTX719eitwEzDOvMmQPEL529KUIs4ukkJM2RBBZIflC
W3JhHJp7nmpeJIzf/CzNrTfoyG5PCsJFprKXNzfizDn/FfbrneORuM1OLY79cFpY
cebZ2tKFb/GeefFzEdiB2kH3H8S/dLDjMbVtEUBTNoh5/29ivXOlqIiPkMfnxzss
YIddRltrlnqfKvaLF0jL52zmY/2eL8C0tqRFmI94Xt3wRCV9xGtTsqjerm7Dw260
4rQm31rn7pjeIyi34gsSvviBFCGxK6pmEjVPBtVmmqwJPHKsMrfRXT2QiVjk/iKC
m3mXOcnzk+xtfNyDBYI/q4BpiN8j2pSbTLQfIXaeSg6rnoUP9Me01vH330fsYd9H
JV0k5FAvTWucqssUjrtbpppdyfxmMNcvh1kurAgYChtWnscSldY1VbQjw5hQyUZL
/UL75N2bTazhiRyeC4DB9WE81A9fC7IkNoMFhSZMX169JfiktfoEuGfdWYxJ8eHy
6Ti4xTyX1iePmVPjftgy1UClkmpYvh026IYv3pz3INuIhZn6+MOlC9dOZ0yFs/oD
AyGGfFbZugjfEZ7zyQPvV9OB7GrDLO4XKB+AtMdaEOSxNdF9LISbhncfmrUnnXmE
w5wLWcNbIdO/hNbqZRIHdxLkqMpyJw1fWdJqIYudIqQBz3h+0vrgnsX8Xo7a1p1B
1XlY+exoUbCpkFbCadXr2UaX43niAGnpsZqH/4lBhqPS4clfGoKcHO8gJELsI0Ps
ZX8dbmg7UnAdWYdDbYS52ZzeXG+3O/AztZIK+ZKmDwNF5qfnTHtOql+y4s2Qsd6y
1r9ABSdAJCaP2owd/ATPkI2nvZjIkAI4G933nWO/e5kX3sX+tjH3g/02x44JZA0J
zyYKrxayh4jvjI1NwS9f9XLxU8gtDviKOjC6ttWwNQ7bB551zQNWQq2Sn6DVES2i
qtcTwU2kinOThqcEbXzUkwImmUivGJvxHIfRIJhN6GnJOzTeKHGQKXB5slzdO489
+lW8WOnzOWDNW6j+LUPMoCdOJ89YT4asUf/dUnXYkhIUbXrbmZtgMp62fT82h6B+
BeXJSk1dFlgVkQ75datXnbvJnjTzTEMrJpKpmO9zUbeHzTRYYNoqmgmXN3usFDxe
oTYVXlu2gtSOF0L6uTMzNCUC4sYnt9Vsktm+uonrhQeUI49etGpmeeT4q2z6oiCH
e9QEFCh7PcMT3cltJDWLe8TXuCwxSizhrkjvHVcD7yap1o/kt8YPhhplaJCYObv8
wmYpbKYIFgNKenVRVle/l0qNn6BuO6AHoKeAi8greYgSRzXeKwuOMFM1Qb9uZtis
8tl7h3LDyfaBbyFkvPXewJ6YKBnmV6Ve/lRjrwsP87wuRKpj6aSjyJjMSyShZgme
XINFeO9817/UJqW12BvdxA5MEmxZHQ7JBMUfXmhhnKuUJtkVmKiRafSv+jsFhWTz
P6bm/IXp2tSuesSqxcNsQ9URHIue96VGAY+XRrgvxAu19Vobtvc54IYPwUJ+i9VW
5NGLLusdJPA8Vi3s3noK9iKQUrYuIG4LBgUDQBPfHKy0NT6XmXZh6nkBmMCCD22K
VBN9uWFqaWeEMxTUKtzZQDGqAN2loJELnYmVKMAac5aY+quxe1V3ZbDSsXrzQtYm
Fm8VGMXD+gddqnwmcAUqwO/XU4oFO8UInBShhJ8ggEQNX6zXWyJ9O7h2eS/Jkrp1
eacgmtSnr70wzkuvJ2OQaJoTU8PF2jrTK+gPlVLRbVDYKA5KEpsoJw5QrrbJ6HwD
Qqo47c78yqO5X1CxntcPf8D+a0EkEAStWg31z/uiYyB/bZPxXGiGlNq+FcuW+GZ9
c1jGbjFDg6Ucncacsg4yvAFGjCfq4q/SotTO6ApTEUqD6etBEmWAJ0uhOqQYb0ae
Qyt/1eY0kQOrXltQFTf/WVwZFWUzwAAMWawPdPAgAyjWfGBrM0u/B1RMnwQ7Yrsn
COD5c3tjicy1n2nZaFtK4AOsex5EFYCe5wVMHOd82yyCZQDhyInAjoe6LdYRMwss
r5nHrSzbMl1awQbR4uE3POFkayFts9cUTRuXbAw21LfG9wrWWCnkx6o23EuMkg6U
VuvjEOD30Tbwbqt1M3RJapdBDweawj7gnILXahcOlyM0YuxibLbyLWz0DxLlHj47
71PPN2zWK5TkaUlUZBKHioaQbYEzMQklTRQDMyXH36JHFoe7xIKfzodY2g1LtTtE
qNisahi3nVSMGHz3xrYlewto8CeboEXTr6kGGVw6KQNM8G70W59z85Rvq/XmbbAb
ZIV/+KAUw/mGG3+x5eRKXyIdZ1YxoAROsxeZIAacGJ0okoR2cRw/4ftTqVNXlmd2
e1wJ3lc8AGNFHBBWrzHW0A2yA+sG4zG3RKrhqrAbJPVo8wOoEuexrlIBAkAWC7iE
liNWaWbRZ2bMLK8ts8V0xHSF/oclXkRLsUZ6s4Uv0Zfp64+x8JZKcMsnTNSkXTKD
GfgaQLpjilN78Q13rkzsb7e390DpOOQYXIBIqL941Y0yYXp6lHeyb2nBfIlLwuFp
UtJwSQxESSM/j9UcNef30w4O/lABPvJhl9D/PH3TlKHDe2Vf1aE+1XjFsrVPbsC1
kBeJqoaq6J9V/P5C27O64xa1vVpzuOj/1C5QDflVDjaPz2mpY2Sexml9kL2GN7TU
h6Fr8OLuGdHL5Mi2FSucSBhebnvKr9ROid77Vwg1g+G+6whXBHz3H9BUqNEbG+Hx
k/Pbb0HC+aW9wNHYiW4H5EsXHrrtrU9Yun8ROLZrlSVhhKDNWGbSnuHg11k6jj/6
xKYnDyVYsMaBIbPUTHccSLWIov9R7jgIgQvk/3j1pWP8cyZ1AXvepL40q/z7UXBG
oxuVi8V0bciw3nrehVYtyIhZ7vNSpFR4m1zKM3aIdzKIwak8KEb64b13CNU+p8Jq
alu/Ow9eCVpUEBxPmNB1UQiAt6matwtkxq4WJH9g4pvVNaou9+EukOhZGy8hErzP
+656Chq1cRMqmCMY0sXNgtML3n6DpukJ5vJTJM+9py5+YkwiBmkPqrScgDdYTnP4
2lgP/OTzY46tKrYo+MewVUQU3F7XtAKRpHn3sKeR9K47oLvNefBmWh7fsP1Qk8NJ
lRGQIqCbh7nDw06FQln6bwz0+1JTnbUtWcty59JKqRZFjE4KSQ6EVC1ZWW8q8u+g
lrnaNOgS8Ds3iGV+ooQF7AYzXHjg2ypL026X3qzW0wjAE9d0C2tk6d52WiHmvFWe
pw/EqVoxJvQ+eRKrPh9cIIKk8OCjQkHsWJa6TNVHx9upbHwiFiaCG1LKK8V9NT3x
9TUx5DqzNZSLK/MjEVbIkWeWp4s52VN76KYgAOkTkhiTTS3Rq/huZrbSekoOsHbQ
ZQk6N7ujcM4RGPbzTny4sQVfkLjYVs60I0aiqAfIM2ZYqjbdEloPvkPyP4qDVoVZ
uL4d5kNAhjgEuK2eFufPuQHXu0it1XL7luhz+ef6NWa839ya9ubZ8AFRRCn7lSQO
H9/NGKS3QkPijaCnmUQaQhRoyzc8YwTiJCFP0EJX0cpM1er6nmj1Da5iC7n/7C/p
Rwmaabb+wpqyftNUGF37RzQ5sBj8tL7OZ6nXVFxpyQb0foKeQjxsMXILJj84Qf5q
bH2Fm65B6M8H3prqZXO38vPAOiaozRihbxuQTg0iLq3L9ynUIZEssPWCiKUC7bKz
354gtWQstTrKOcwASLcl5JXFMS4vWP2TOsK/RJYnvoMU5ZY5irVQTuNNnJIxwYS4
4Lkf41pf1APy18UYCBFVOFN55nwvKBX4VHOhVVakw44Wz91qHGLwYmf1oKb5k/eR
4pVznxtKEGmn2wciYIDan5TKUVSx98JjTefyXtl+7F8j7mn1NvzEVHZ92OhAzeZE
7T5yPTA9bGedwv4VuHs6SK00jVbj1iLsz7rhQFswy3Ahh02uTn2rcD7nmOFgi7iS
EfzfLpEgJC0oCc/qtQTRvImQpZ/yArPXyxc6hS5ivxm68HZ39IwFLctu37ceZQR/
iMSehuoXZ6O3oHCQlIZe+oiIC2+ml1Hcm3mRKQ6HuZ6TbyuVE3O+JtITeLpc3Ofx
BZZnDtcoBg/Kx+yqrnZgCYfji9evgDytmP3Wloi/OF6+3X6V8mVUkbtQlfzRmab0
JxiKAnv/nuxFAOMtG83/LwtLIK4GFHQ2giGyNIkgobA/z0C/Ep4Csjf+I/G/dsHS
NPUq7kpp3NHJD2wQn1wIoK0eFUtg5235PBrjjlFaspUg77C9hVH1HUhXJbFNUG33
Tq/AIf78RzOMyHrjrpR2S2J19DBDq8jK+ZRGok/qR0q1NqhGiiwM+4i1JeT0ZE5T
mmr6I4EjmFooyj9K31Ghm3KiprcNoQRpaPJnHFGvRw4rqY82t5nYM7+zO4C3sCqY
UPZgdqE7qfMT5TfbtpiO1f/bG8Uzb8+ygGsSi4jlWYQTmV154YhKJ3FodYFfqbAr
p8cGw/YE0BXcSDHL2Y0dPs+k2XgsXmg81I5nSakODItFKILIgTaMNX62M2dvGnzr
73XOBCK+W/EB5z1EbrMIs09fegHpkccO958i1bh1EfDeGwsoOxJEXsDW/DyP2jx4
3WQbzpp63KoL/K+hQ06nD/3Jfbo9G6YKImskDEx50HidBNKcQsP8wgMO/zedwjwu
5ay6gYHCQGmKatTY9GVVwZGmmRmxzFO+gr1duQxwcJMGyxXEn90Q9e/6kAhyCzRB
7FLLO6vv9WZK2ALbG7sghmmAnjB9GH5ks9J2Hl7PCRmqM13CEZrsStQ8uHW0Tgm5
kqf3jSsSjKdJRiPl0iulw4aPu9/RgJvey3kayZhsihvaE+m43Q8ZggCHXSp/Y/6B
0cuq1olczCI6yY8xQqhtjWW/iH3/6koVALZjjV/eovVlCCqzwIjkTf6/x3a9Ixyn
mhAVWXC19GLLycxS8V/gryeXsZqyWsbFQr3Vy1MhO8WKDZRiGBjR8jK0IsSVclWP
xfMLUQ9tSDrnfy4L8KoalBRhu2OEyALBihVEE4EvBp1dQB8grV6g/NO22jvK2u0p
c1VGux0FiJVmRhHTEJXIyqYeuU3tS8WA5VQFObD0VV4I/oMTmwLJ6T7xWSW7IoLC
bKs1CQnNWGbfksed7PEjhxoKsDRw1EY1eQrO2RejqRFonWjfBEcHa37sXGdu2pSR
krbEjRphdp9rkzjg8MMjmnpnK2UunWFE90Dp/oSGbYhGDWS6kORtFYHfYOXSVS1l
w/7xhHp48XVV5W9Ba4stkNJBrSd2/VguSTEVnkBvNELvMMVSjOQ3+w4PJKbWxVmB
aCcIAQxJwZqBJYbgS9+wGbJgyPbUwly174EGJHs9gR+ok2XjcDLEl8KVNXXKisVl
spt8bqVRLyDSZBtNd2evBtTGy1A/Zago8uCeDVWzMPN0P9jy6fXJ01hk5FFXowFP
vgbZaGaqvecPBK5TbdQTX6udtTNQY1NeXsDf3thYRYw89IL451HAdK8Ce2uwkyo/
pipawAzLg1oEY20UGYwuuhMOLhw4mqfd+FJO6r/iasBD6Od7zUnjLvCPpXI+4onk
jZvK6vEIwemT2vxhQeKnTRAwALWMjreC5NCFEdI6xA9bkuEKTI4h9c5CXqiaxzfp
yOOVDfm8RmK33V+IF2ihrqVCySh43EB7tJ+zS7m5citcnYnPXqYB64276cJpJoMl
6Who0j5u6l5j7wo12Q7rky5yjayD4Bal23FZDpkyevvq+JAKm9qtelA8ZxDronrN
dGtgwBjQIKIoAW2qVzami2Q7J3mX6qC+kXSYWQxda312LPOUytdJZrki4XM1mSw4
HjsS6FYgmaZJg3dizpJe8vNSWB2W8ULDSb5taPIp13DR9XCI2CQWD3JQpanPL1Zv
MDwveRS2o8d/ZTQnKOYkVP8U9Op91UqqAJurI1c6ADflT2hJAvQZKEzEZjZ5FIJQ
J/dgtC1XnDychGjSGcK3if0DKCOgntetVPcO6m9pIvUpYq5IdeEWIRQtiuQY2HTo
OT2vNCKdKUdRILPD4TOAyJHxLjR3AflqLWOyuFDPhqWSpitf7Cx86c1JibcObKeQ
iJ7t6GL17EEmEyi0/RbWzJekUm1xc41FSdJKiMbroYhHmQAHbZuobPwa6s33tfUN
Jdrz/cnE9l15IUAWACdfA8Y2Gyk5SptW85+hcbwFp3fXFjx/zrS5v6whSjJp3dcO
3T5QosidRw+decU4igdlCF6277SI47CDP49dTjCCJkKBd7PrvMVX6rAbJQTxiEtJ
LjrOiAs3As0N71e1rNmXxlw1RNgzVCwNVyFca5hQEFUP8MIjHoKsiR8hkaAsJ2Va
Xk4i53wVSHqbLyStUbbGIQU2PY3LdoRYWGkvjyzljFAaoe5gdWLRA+QPpJtdEAKf
UGtAEk6FWwUOHcCokRRsByKJr7B/AFi/y4YcUHr6yFbhqE415vRu3mtdkDsa0oSA
IppQfrndiMWifngKEvapIZfFrLjgRqzpX0f/H1lNKeX/bLZWqnBuThH40ZPh76gl
AhjxNtxUTI480agUrOjH1ngipp/ZEJ6od/1YkqCgVZhihGXi2ReZGt6l8tsz/Dm0
R60oYrERjxantaqnkxvG46wMcvr3Zi6supUyq/Nq7PHEgQaBUoSDjB6S7a7aNalW
zbqAuGna/AfJda8JnebU2n51cBWq0zczQ5Iz7T5BodOa/gVUL1v051SId0ZXM2ms
ywOOyl5KpAIp97G5fXL8LSqmQvkmHiLn+eK0x2hfh834ZBhjekS2fb53hWh565wZ
wFYKy9RC83jWW5GQGWNwrl9CiwWafnoSzxna5gRfYFep/5GyVsqVr8rplXEeJIAL
qd6GeLxfVySGwUDZFWeus1UnpGsQ/z0uf0SnDK0Z0mFMoeFeVORvdXQrPNyogFyx
BBc1M1d8PLOhlx3JoBrymyFZe3E3dYmNkkxCnQAj0B7oSB59ZhZRnILOfDSXv4xd
1I2mcRQ3COwHa7LYvajsytZ68Y6+xs9rO07rqfJtTLa/SHIuB5C5gSd4DNo60qiA
N1KdkfwNu8RpCJMm3mafSthujKuEDwWLZFX9ZB1IiN5kkcff0XnUive1qx/fG/UP
1IbrH9z8g4FNjnoEebV52LxJBQwoGgIOeXyGwzbN+Yy+b2jFk+izJZ8ppr4Hj0gg
HNVD445lb9YF6KDggVYQFexre94qUfdUvHyoHWCK/wE/1fzqxvjV1HkWCWtDZyX/
QyCirsoCTEbGi/zaBg/P4P7utC2jzEYU/mMwcdtZ55KVvn1U8ZkxxifKtjNm07jX
sajF2oMrklCul7MMYR3RdxeQj4jk2E1AM3SaR0tkW8Qga5uDJ9/+DtZCplXseUVB
FxUkgngLbwjWTDJjViUBDrP5agSD6+SGK9EL/YUnURc1+AyXyQCdp/kFeSDHp+OL
CTOZSNy29xVWYhuHjb7TP3baHxVEYXY+fLgw5qQMVvpB3kbWmnWIvVwDVr/5sHoW
N8P+7RCpnX5VmabarMbUx62WJIMekj4R8KpxqXKcAPrSsnOKrhogAkrgUSJhNQFj
ynfbr254SfEuac9mUIYRWcn8uzvBmtySqv7bC1alyUSFxYTKKApSu/n4Nl9Bcico
uSuzztXMIOISyVcMMFaUQKUzngQtIPAu/4jd2jbNt7VIchw6nd+kYAmYeIrUYAj2
LfMUOwzRXPFbaMEpgckZbGq2tWbRX2pa4Z5E6gLLhbHtfHs1bc7buhnklTzd0ink
9uJEDUDVC3FNec5PKcPwjUncAzF9pmbmQBTG0ITWDU/d1xNElv8M/TtVx91BH6EA
IVrBsPZr87q0bDLc7bEnh+mEMtFO+ki4HVj0GRdEXe/vvsOElxa0DyEqu6FuVkqx
5ykWvvDX99JnMMDR40UeFYafdznVzywjtZN4uxsgWgBVarwMx2zFsCNnm6IRVcug
9IkpoASRgRV5A+aMSXN8p4LIa9kzd+hky+Xcxc9gxIEWB7GHYkY/kYz2Jh6N1i3R
FdGMmNP1dcp8b9gmnXfRB+mL5MV2PqJFcVzjNRyqMoyNuifwtjRl3X4pFsOOSSso
C0glPdp/KRl+ZjhwaxxEdFFmQA+or4RHVCwpTBDwS5YdsBp0eggKI2zqrAr77vpY
toVrthAJ4ylYKgkas6zyqYycAxotcRvoskfrL83FQsPbNHd28JEVwoK8nS1ffCYT
BfHl3LA9+HWyBRZxaarzeEia0smhVrSRgEheOh6Ebnb8vSA/PKgtZK+SZ6UZLPJg
W3yf3uuQENu8DqJnFudAQygpgnbl/xk2EWObhjr8HIMFQDHAvrvttUhkvJ65q3ss
qKDeG/OhVfhVcxR2A73ghvLYM0P/BbjUv5n/hTIltMM0Z/gtJ6PlRp2lszwVv5QZ
LILwCxkDUOx1cx6LYek67llMkAy3M8ocdl9NzmUxLQUCvJFyrrjm3JXOvijHgyGF
fCqUyu0ROl54YvFtggk3bS17L1K69W6GC5y0+eenm+bivubnRVU6WQDTLxcp7XnA
7vEnOFScqL/pa+14LGRf9iXxnDftxMbJb7noKUDgWNXY2V0gZr/t5qv9H9kcfeR7
lqUrxI2nSyTjeslA1I4imyCRzfuckmGGvnp1GQxNXuJLiVYZBeBzpvSMKMyqLJ+x
0QTlHQxn6fVmFpITD6+YeOwmNMFEuSzXjut4527DYkTFliHC7Whcy3PWHwPuqdD/
YwC7fEWQd2EA1KelFGijLxPTd+EKUqzAyHPtlmnHZT/jddrnFfu5oayj/OT8sh3y
bvl/uRjM/47TNMEK1p28muErQ00ZIRdnf33yarTSRkHh0Av3XQcXL+9cVWkDirBg
KvR25HKv3Z9aYK8PvwrcyoLAqks5iDK+Q09NUyP/yS1dVEv9GSdD7NQpj76CbPG1
WiyeeTEk2B/rieP/G3/6ZsM8M6ispDd7cs9r7NC7f4E5eSBcBGnBxAsn3KDXZstR
OUMEEAQ5hxZMXIsmlzYeQjIcjKgmMyrPoq3rL95T8Sxk3GYs2jCHnaE6AlwkmUfc
TvVnrZ7l5llwiVRT1+CXrvIfmvhudldFZejyC9H83tqflSNGudkE0kzewsghE6Vf
CvJaiEMAQzrwSf2JhReLy2JsMzREjRrVPZYSJzQ2wmyAA3Pm3wkD0b57+o7XIdNO
sFVXpR9PoQAfk7L0vDa7fh9CC+kWXREUlO60Rrl0eIlY2k76VetVs2PB/RHAu5Lb
v80jGnlfKzXOYeSDXQA7Ctp5jRPJk0T8vuLvB1w+uzYKTm4Wbz83HMDVcxPaqbUu
MHjBEV9h0Nf0EJODHICVR1YJsz4feOkbF7n5nGtE1WTZt0nO2KyEDFK43ir6a8Oh
ApR+Er+vdSAS8PlvKzWV3ELtlA74DCnbs9n6JrII8CyBw3FXakjpTn6D+nXIYCrO
FerNEPwXhO9xSaIa1xzfPCLMN9r1lwGnKQluK0S1yWtDHV1H28onxE8eE/NWxMKH
tRag225wKkA7SpJe8H+2fD5AT8l6GZEgmywpRMCfhhwOg7Lt7IkPN3FpDnqrNr9w
mjAW6Q4YBARN7HQKlW9ZqcJSBGSDhI4LJH5bHhy/UbJv7bcs14VhoR+xpqLrhtBx
za/fVubOmaTxlwc7ILwOuPYxt/l2NAhKwq5yhj2C2mtLAbcRLh+16GWy7/dwPNTO
ElV2sEvP++ljIedFJxnW1h19CwzW+PUmnqSniyI8z1MoLnNXlNnTVAvTOyYvm2se
gxP4VgamLGkHIrRqTPee/MewkpLXdM7sGvUEXHQa28SOjW/arDhNf8MerOk8eII+
3NxWE5LHIZd3MYlrpAnUMFs0LpTUshNrUk9/tl721QDf2y22tpN2+fgkzYAHdte5
VGn64QUeXz17zt5xdqLEv3mc5tljZMl6TfaHNWhQAkVL09diq8aa/krFpO2wizJi
BnH0VZplWERfi0p3X9UxLJNYDsAx5PoIN4B2t4+Uvpb1vKcjkIPd69jUweKLVmSj
GUa/rY5tQs/SYPqK2xyGFt3+HoUffMHOhcOF/WPuzf2qAG+KAO7vq1rrqAViWNeX
EBITWJ5RDpvFoSCphR//OYNmqURajAMKRi49Xqz7542d6tu0HMgLQ7SqjslsxbP+
EYCrGxW4ST9fvGgWPz9yW/3kNPxH8WJGsN7YkLNH4wjQtd3NyzQ+RMLexgmE0teb
HOn0iUKY/Qj52AuzNrnHBVoSmxtYFrorANX+l9sr2GCrrCZiECRWxMpj4U6krs0e
TZmdXyFDPD6bIGc1U1cvssAbINesbrvlHDNHXjVPrUjOmg++vwW5321bXEZMRqPS
70n4lVWb2jwousaJlGgm0gtvE4Z/sRiAhDPUduijyLygVFs3uIArvjDP8x9rRQAa
IBUF3PoIdLdqMmDASsDoguLsL+nVnqgLg3tiwJrxO3mdROuCP9AhX3u6fQKARenH
ruFgurSqejV/ik5qy0u0HA4ra+SCp0mDVcFornGKN7+F3bMkNsM/HMXqulrFyRhm
r389y/69nd0+vYoDqt05AYkK5Tif82D7BK+1egk43z9b3qCB/1TAa9MT7jZnbZJv
A2D5EUOD7TKoXx1Ojz2JYsi6rIkfZa++y585CL0tsUYc+saf61Xd8xnPq4DLwykr
92AvfeSuD8wyLpbRRh7gr2CNcMW9veX1DtNeHrTFGkRBK1YoP4N385WS0D5OBfPW
c79TNiybua+EFiZtYxrpf+bkFvCLB4LcSLWEnY+u+M1F3y+swyHtlYSuFCXz+96l
rMa/ffA1AHoT5horY3kPLzRcTM7eHet4S2ZDI7BKZUb+q7n7dsiZ2lxh64jRGhQn
IilHoEm2WzPFD5kzHYbGGktIG90NzdHyq8yC+MS4dmBi64LUkRbXbLaEE/nouNAq
WQ/hVm+A2vhvW9EyxyrUSVMmHzf47yaoI1qC34dyrqO/m7nyAl4zWBndxhXQbizv
lgH3vKnYlwtlS/pBSVADMejh7mWmMhcyOihIQEgXmi55qXKQJ3ktiM9xRq9qOcf8
slI3l3MY9NqWXc7nSMfCNkrKXk0ZiInKlLgBlJuWgmSdEUTbp2+DFv6ngLgHW+5V
Sq0HuZv/BrA0yRkqJqzuEK7FPBLenVEr/nV14lCv+1AGPgSnSV6UkKh3dBrTKgqQ
3C79tEAfY2y5bIdb3rJ+qZ1fHQNjNWzPk+3Uf9eneRopa7i1GbSJTWzv8L/el9Zn
0l/nuSr7s3vXxbB98W26ICtpjMEDjuvLBCXcMzpAsgSxMd/4kOZOCZjKpgeVTHCz
WZKSOGIvZr1oIbCX0JcOP6HhuC7hzIIiSNkub43fz8CEiYFA6nCcBPAbE8RBKrqM
o19ji53aIidf9h5vFTtxXTaIlFJRQBxQEcO66bx2criO3N9B1D4kkQVClFDsOetp
z8DYsrZboh3cptMUjzMiwKjs4MZiqq+j3KkgzQ11v7M4XCWMgaeFxC+bc9zZZfFQ
DjvCOigMzMHc/hWH4QDKmYz/brmV+Yzz5ZNrfeqnNkhX2UH2QFs8ebsWz07oHqgm
M8ti/F1K9O667pyi8z48s9n5oyTSeIgDw1Wxz5gO9gHc5mSGVJHNlbMw2Dm7B6ws
WUWV+MvLyxkf5aJQKovUHfeblkfwy/FJyaYjEuVZaCFVEu6MUYDkaj1SBtyb316L
djm3fZ5+5N0p5MxonXv10Ih6M4BqUb0KDeC2j1hwMtZnC33/Lkf3x+Ob3UR96Uw7
skCtwTQaZ7JVLmpCkhs5a5d/Zw62cTpWpiALz4BXyToR4dhB/TzgZFtXZwakbbV/
QLjM/+GETantQ+Heho+PW1y885jQEz1TsmrzDEE6yf2PpBC38JoSKOCeysXY8Vjk
autmBM1/9BwcIYN/Rs2CsRrhkOvCCJCgmU61x8Rephosn1G/UcHmDpt++qkUdHoP
5vYQHlt9Z5FvKvKo3G0xDolwn6sYr13ZqHtaa7gAuDFQ3hmis66rAhZNIBvwLIGB
PfibCX2Swt0gtpE77UcZAO/Tivh6Qkp8zz1SWOTma7hQPTn1hApe3HP6W392HMrd
8DzNwrRCwD+IBIiRlR4r9QFlbkBA0/E3ABkdgOlvoIecZgy4ZvI9xNL8n+bL5xcg
p5x6MAZe6IKalf/ZDK8Cl/lKOORTkIcfBPL5zsaPJ4PChM+Gn6H1cbN/LTVFg/+T
ojYI47I49yt5WbSsM5MBWyAhhZZAl1O3izC9/2clae6bi95wfJKLAdty+ZDsqKx1
NYskEcKp/bFCEUrsPR+D0sbZveQxukRAS24iP/pFJ3e9D0DGbRuZNBLfYJTqby3S
gG+FN1UqskkKv9+c8eXvVSYN5mEAHV0MCFY57GQKHDOzy0p7eRUEshdnhzw4MOGt
wZ9OuQ5oCX0FGuOvtuUFcjP59qn/dbH4JHa+9RXDd/EB86J5rj1PiC7KCl6xdC6H
dlACNlY7hPWXhvUlEU6LWIOl94FCfqJU9PAuf5FlWXGLzUQed/oJS440cj+fChnW
hMmq/2n2bhU7vQ1U5CUDIMDtE8+Y2ewdwpr20EPf/PM0gv6JNXsJKs44zBq79g0y
d2CyvnIuCpMlndCeyMJFp2oMSBpAQDYSeCh2+GHhOwFhe/M4S+O4fzmF16lGrR4F
RRpLI4xp5lgZASkUPohOocNQ2ghVALbLiSdrWXkrHoLs9uDyP/KifzQZihs3uP1s
OTOUsjZ+T+T+28O+NDb9++yS820RLTHz4Zvb0AhBpI/X0kHACcC8pgq5vpIwns2d
FOnBJFMprOVyRMVWgsvCJthlqRukloKNdQaNnDDbEa7sNGkSGDq+fwxsH189nF5p
qyCxqPK93RdgDEFFxlpEYK7KCnY7fd33P9OdXVL5JBHFkTOyAp170Blf3Rk7HTc+
RJDtj99/Eb2yEqgkHWoHFaZyxL7ZHlgQA1RhSSQ6yfem3KjdfgY9dtORiNzrgtG+
/5jIHubBD1bu6XJxV9WVyaunsnzwuyUq4j8/kjGmfdHWZ1M6WB0gW87vCysES6sl
jR0zKWvrbVSa96Rf/cn4hYrI7hcKG1v5bl2TtWBIuwzWTo5Kp2GFwqvJl4+o3f3r
gVLZ3+fur6hAXCawKIPfGI6m3/2vIhOKtpYWb0axumPceN1hq21VFPRtdzhEmG/o
ioqYqYHmS33hQAO6E09OxXyL/PoF7YTQxnL4dznkN/wS4+azEMZqERgIa6kmtlTF
L9LnyR3tjiQSz+fb7F3aZBl7ftyLvFsA6HUbUZDiQHupviIlrvtWdNGLBj6LqCEA
TvP0gIAJhxeT/ceKawimpIjkUWK+P4DS4b460V7u2h+6r0bG9lgeq9PbM4r5tWSo
CF0Swueq34Fc7Vj/UnYUM8r9y9ypIY4G2iEtHhFlozz6BQI8c42FbEcGikchdtKD
HZvMeQGWESNI7X41vh6PMPXOXmvMXlE9QkcsYAXHAEawn9o06+7TTBw4tP/+leMf
UaoKuYAq4WaIsJDPZNtQxddiA0nvrWOAGq0QzY5JQ1itkg1/SXVnrZA6viG/IumP
HNncyIKVk5vUbNhCnM73+2xNTtLEO9QKlS+zlZ3pCt7RyPz2h/KFuoAMeDPY5SOJ
XCon8C50n4/uHvJrwzdIgau+iz0+EkiJkHlz0gKXjIPqTKMhFtIxzkHhfFSWoC5n
T0abjWJ3e9deL0N3/Mk/L7sS3hQr11PQm6qCK+bs1WtG+1QhBhea0atsLlVm7zXx
D7wpiQkd08o1zNhyocuiSBf1yoUi21CkSwe4xpDp533eo/4y4aPKub/YIX6dT5kf
p+K1Mp//m6kJgijU0s1UoUQ9hzEruSkmg/Kwt0rhCU1wT/oSIqHjAywYVCniPtwZ
HNxrB/mCpYNtuMu/g2Jc7q8lBnOOyeUp3UKwr1uUCjxgqkywN+QnjZczN5nVBvDt
8qIUePmKCVzvMVC9O69fy0EyFtFesgPzIGGRgUDbj93vj5IX6i1+aOWKK8TyDge5
Q2j2oOSq4XJ0gW/yqE5JleBsqlYBzGczICXiOIyCVPQgQO5Lqg3fPunq2qk66zNm
SqW5fzJNUaoKieiXMILVtnDAY9J8JrnrhfjFXiGqqdM5uXA7yl3zjkvmmbLaPoil
DNEx1UGzN4ZRNsTlgO43Dl2VqJgWtDriNkGlFub6rJJrGfpzCH/Batq67mfRYvbh
52cxmodbg/Kl7e9wTleJktfgx133QwzR5vMre3QaRDUbzobZSpcnX9slLGZQLvxu
M1Xe7OUcZXpkSbwoDRSkyh1TxGscrJ83owA0idcCze/vmRvLUsT0a3bF2T1E9ujf
7bCoLHmU7DLn7aJZdBcuv6H/SwEySo+XfA1qoCWzicbzzXOHe0YNre9TFmuPq/yW
LQ+G8B7hEEWFflPeZkAzZFQfbmvI9k1V1SN1/uwnv6waRbIpx1oNhUhqiqm/ClEU
tKSsPh/c4zMUD7OQDm1kX4TArKfjVJDWdFobk3peNPxrxix2ZxKQ4yrrs0TzN+PO
rzmqzHbO+a4wa2BM1uM/uBYLkVOgP8hy54kk8JjjRvRpzar2uZUXkAEVpEsXWRG7
iS0FYVjYa5unLFAGJurKx/wrzNNZxs4X4bcfguxXbbMw7YroBHYcPyNKvfS1DwWk
ZFE7TqIz3W0O2tBVO340JE1x2upodcoBLLsNLxnUxpo3iNlcclHvGOoDE6/qrGpS
0li8rwuhF7rp4bL757kUFyMBrmHRLPftqsR/Zxvba4fMxi3iWrdgmPXGE407aHiO
tl7azAcEiFCkJIEHYJYVt3sUPDdyHZPU3qYnCPr1GsZc4AVbaTX7PmrltPmIfF1b
nPJs0iBjf/9TC8Aw511CDyEQQewuMdYZ4v+0vzJ9HvDMdcOSz75Hzg9W6nbYJbjd
AbD/h8GULVah19CyNDa/ZaJnp3VqdkpZGFe4aRVoVOHmqE6ewxei4gp1EK7YNbKu
mJmkUYS8fBTWYKxHCUKwJNlpYisBVYCUKvNlwtkcmfx0F/+vUXD7IdEut+wc85C7
TQnVnIpDadL5LH2UE4nSLEfnPlMPb5unDoK3HECDWDk0mRylPrSW+DbE5BpUhtss
hU8PbfotABQmNhwwIJV7TB9J/g8VAlGtb3l+rpiLEaF7rycvnO1SzCaWiPICHR5D
dyLOFcM4NrTwnyLx/v/cvrjN8flH4vzMnq17XDA73KQ9YEyscxecSRAEuSE6i1Ol
crpRZ0XidVDk/uh0MRJo9QIUZmkx/eB2RPmFx9Qyg5FkJwWBGEQOArjgkl9doQ57
FKdN8izsJ67tZ2tkBzK4nUm40xI/V6391CFlyXQvZYRqWqA64MN0GHQwPMctU5ZB
+VLf8lqxV0Ft0ZzwZ7egWs69h5QbTHjKkpNKrLiRVAHP6uO7y6W3oF5/RPxuQ234
UUGhn5fQpZszUlCN5lZ6gPF72LG7mwRifGyIPXvJFEqrPlz/hn7fEhZCVCk/6WAd
1EFhQ4gHtn0drpeGnnLFHFPyTNNhQQsIq28K5BIfjMIEsbksBVw94oh+YvYBFQku
5AXOZG6mxSvaU2aT0mBirK+AGg1xrBMfW1cs1daq+pQ2G9FTuGyQzlDazaSkLzeN
HjdTAs9aKDD78KCppw+gWY268uqVdZMA0WUBPqjQ1sLuwziuQZBDON0/H4e/9yXR
6bth991xluyorggN0GFWMJpbV9nOcP/IEhdt9s2yKq7xYy6KwG2R5PMM7Y42XFrj
IGu08BO42jyRxbxlryrlqlC9juD+cdfjrZPxdhXqMLkyIKVRD++/12O7k15jZowX
k7Bo4Bwywn3xOm1A8lKvCNvG/egybWl9G0DKGYPi7f0nSq7w8hhw6zKUh40y9w9U
WNlTbRfhE/ZBi9Lt1tV+e+FFR/uI+w7/GCUYjdoL/qvVT14gkaEK/Wjr6y6HNL1e
3v8wzrUQRkESWsrrbzelkQgCNfnNYqTCOZXqntYb4UmrVDxTrMUQJ4DI7AjJxTmF
NUpydkrSiNzBEktZF0CckCGM16djMvoZnLgd85t7QdYOeunEObjuFYmSAKvXj1St
fRlrNla4f4tiaFlOojsqhqdkpUfKDcj/9jyAZN7tUcsKOIWwrCXcIYSH2cXZgmFQ
xhhEYvwxbYB1WFokiyCGUipZ9DPsfzAK79/l2Jk92KQwLvR3UNh0TBbR1flClfok
B8pMGYvIbjluNAiI2m9psUdZzfNt2zGuUE9XEC8SkMyQGWQ1XiPolDf7dD5yN6IK
w5SV1w0Pm1jCfEAJ1UQuimxEyx5XOs1kixqVrMUxrBG10xtGtBBEe3i1CSwT/uNG
WyevMv4iScSMnlYRpwcYxLVDN6AEPp4TXBa04lXIMjPE/1kvGXjEntcthaIUB32P
wrh7BduCeUj3ER23F+meMdZ6uTG5CvnMOM6UQ/RK4oZtv4sYSVnELxgTRcjIu8PA
zWlGBmfIaAcqgh+ts6BRS4HKSzd+R2CNsIH5SqFFlfbsr0pnNwKxKonCCdTEclW5
JCrxjjSQj4Wtn43kJjRV08+c/ANPl1/BB7q3YD00mSRiFOPIyTN145tYN+/gDDkr
bJawaA1hw+vN6Dht7ieI51tQcXKtHYpqwc+5QBn4s44CkC77IclrAzO2jRMuQR/m
L9mv+Ds6hQaGWq5DSJQIt+Qc4whItU2Sp55GTR5Znc6dNju1Uok2B3bXSfMzcCVD
tGvPilGV9JbzQrRMw9rjCovcc7yN5xv19rkwH9cgCywtplY3CJoz91zES5wZgk2S
PgN9vKDshZmsS/TooL5O7hGjOhj13/kO8VYbflc5xrV7dtUL3VjjOXbmnroBGkmY
eTn7bQB/3ThugOvljpQD55l7jy4a3eZ47YwCr1ju/JqaoUM7z9MMmIvXqgGb+VXO
EHlY7plsIppMrW/KKsEPYl1QWAv7i8G7yj1DRol37AQe/wxnM/MvHlr1tP7dmOtp
PNP4qlGBdowhkK4TeoxjJvhAHuy/sMIhyksQUdXhM+CrIwJujz5p6B9WJG4oaWKg
UFcVNgmCheLz3uDO8l20DAF/+BVxCZNCWRGu9t/lP0mWndQ/ikI4p8szzvH6BceO
uJGXkMg/TGyQHDBKx02bm0T07qZt+s2DX7VG1Y5YIDCiOsawZZFuXWNZjrmCm22d
0/wju1bcO/jm6OYo/v0l0RvCQUJck0dwJDF+EnMG421rSGjK4dsy9rRpSiaCvYni
uacj3+9fNnPBr88CN3G8gv6Zc4MQ45eKl42r/Bfl5PLdm11tSRoWKwY5dPlpO2LQ
MIn4SL+KgdfyinYUwjovEPbUHmFNSZ3SJGd5H6eOm8w3Jo4ZvB1zGiO7Xt7lRKaZ
kxeGFIyPZfH7GlA/OqFhjnjx8+4HHMK5CmaPDVm8NVxp/Gx7rSPocr4nHPeRWiju
0YyChKmAwjHV7RvFT+5vGi7fgvROwGQflmO8OOK+aLZa51HDgTLH4NvkRFHYXxJv
PA2Br3J6NuhnHXcHvLZ5K1DwM9Z7tdWCPedr6fA1AAVsVPbpu/HWU2gLJr8+ExzF
sbc2LLY7FFaJoJXi9P/OUplF5eyr3we7FOmUlBuNgQ4OjLnuZXNYRx+fya4jPxc7
1Xh241mjb7FsMSboOjCfjmWrbTsguneHV0H5l4T4KAiGWNADwjiLtYb/9k842eDO
st+ZDfA8QP1e9yKPt4TP8WFD1balLeRKR2mq+JZMtIQn4piph8CQK+IvweBZ1B65
ouRQ5KF4dFmmmlW2LKMBs71Kp671Mjfmufm15uw3udoIEAbJOIwzkghwUKAY0CF8
2tAKIthLiqxYP9EpK1N6/GGXVm+gQkdMQ2l70UugPhFhfEoVIJGR8UxIaWpTvWY8
jX79bwOpxNzfwtvCT2zt0OTJGuYDAee230YoiLWL5qoVPAR/18FV2Iv8F5SD+vVU
P4nWgFAsH4eMge+F4AfD+VBw1HQAdlgBIpNjgASy9iBrIxnns65sJ74ESAvWVv5q
PRyl9gbhzt1V7GgABOZ2cPgEmfIR6Ex/zqkDynXXolw3l3m+Cm6V1NPwKsdSYYr5
Dn6A8JneU8vBtIyQ1nRBnpauF1a07A5Nuj/l4+mgpBuwgE36UrYPmoSqP+/9ho7h
jas+13iKEk2EhW4QPtWsP83A1M6aUNeuXKi0CJOeVGXahTRhaWdScTaHU8rwt37S
/OEp0nSJEc9/t+lkt9sCDmsoKqtSmCpF/FAoTmWDwVOW2WpZaTO0dYV3+zcpHFRw
kT3isy76lW7J2kgHrT5kTHE5XihtqY0KTcJ0nU92PLgM5HHIsSTFw8E92UgIaIrI
eXMqIL+3BRGZOynrhZqcHfuu6RMO0A+6TxgWhzXt8YPMfCi5OKzcngUiTl1hJ9vg
+YDa7fwMjphE/lCszvVYvA2keDFj+/U7Yo1NgDdnoUc6dScNIKiV6FA8nLKjghHx
hZTRH+PiEZasjPaymaNmt16BoNzKcFtjA7j8ViIauV09Ss4nQfQEctWNI4RCusjI
DPUlqpAN/uCLhmo4cA0ITjN4sNjm2N4P3kUDLF79hTklG7HovYxt8iKsJ7IabSqa
lBkuJi2Ytmb337cZ1bXLW41CO4U9C9DDbkzheMbGE5MUIO/qvj3k6y0zI0m/lhKW
CHSRe9QGl7U8JeQxFYrV3e52CxFWji4jFAdxUz4Y85Ik73oNOKits6bBSAkw5ZQJ
khb/dHiLMtbE+V3TKUmuj+QskDevuoa+EpzAeycqMfzyuBjAezP0cDsVc3kDbd8Y
kM1bVy42LWj2g2/dnrk2x4xsQd7yEjaOgaqcPlt6EfLrBHvpdGwfo9rasDGxSjet
0PkkQJwr0cgCZetLscDCarn+e4W3jI6dJwbUkskgv2uw98NfcXgA2DVWHDxmBh7i
32yGmWlS9AgTQeaL84LfVsKPCKMtCu+oZrX4Gw/NAJz2hVx/+fr/v1HfbAhn97vE
UMmZTcDoSxxudb06k+UYnrkzqa2/U211nGUeGT2rOYwEbJjdT75BZmI+xg5tfMzM
o1EP8N+Z2JtPbniQ+U5fn8uEjsLAFipir+Odh42tJqEeCgwyfRZ2Pz4+U3S5yMlS
UBU/YJzqFLLttR4zskDYHq5CJbjL+5TTA19pzNWlJ0ASB/UBH93I/py2d8HmABBN
lwm+JEA7IrOtovyljIX8LBuEZvKe0c45BW/iwA6DnOl7ZNZ3Yb3Amr0IJ8LZk/Uk
xYTzwCjCQWjKAkQ2FCuRJAeAY4u/wnXUC93paSvwTVV8lOriVFOxvlm63dHowWtx
JK45u3hjD7i0gp1++ilUifod91BGcfHsizEixjt2AY6kQH3+RnprqkQ/5xOTa71z
lw413NeADZ8cyCYxv2cpMKXlzbQv3FOjuSMBJq/RB9miNlkeXkc4R4PJdV3OjCxq
RIef+YORmbQ4gfBd/Hq7gsYZxQDjK/+fQrK2mtNlSXn9GC14TVIQ2L68cNuI6v16
VPcFcjve4Qsh29hRVliJBbeGHhIJIQAQE4GEekAyiyeqlo5YrUV2ycfvbgtlhNBw
K9t45bg/r58Cc2grzeXqfbJFxqPGC6MGD1YMwEeI9K6391iWkAG+wfpr6EuiXyw0
E0bGaoRzbnZOo2z5jIF2zmfccsts7S36FzUZBKtFUSZ78RyiMcH1l2heE5GAsEuh
Yyl+PsHoNhMxLEWU4FiaZRcCFs0rOA1LP5Vl09vy3MYswYnKzttWtqrRJzQdTQbL
bVyDhLFsUDlJFoETiEL8C6eOSJloIsIWSf2NQ0oSGZTGKB2UtXudisPxVhVGp9jf
qwB+ygN8iOyTsY1mIPnEDgE3FE+vH+8R8UlKGSC1zZHIsYHCeimsRuSLeBhmnec3
zBcV213KbMXLwQl9FNtxdRXQQ7dGPcp4LDr3hh9yMvSW/11gCPhkFra5+N6A4MQX
/MeMW7on8yh6wAKRBRmLCjsipRm3ZGRniDN5nwEq0fJEqczWWL0Qipi1WRotm7so
+dn0hzYWQ4qHMFHhyJS+0TwfTJzjnM46a1qgEKqQ1AfME8LYJGN98c7kZ095cgq7
GYPyqFESSk0bH9q4vzDW/1teFH9pC1u7r/+bbzHKoe61QYkjPaZKrgX39a20gnQ+
UzmkBysDMtJGpw/31jh0wPWLDL4x2GgF8qTJglpTnml9Ajp1h3krOCZOA6gcNEzp
QiRqxrO5YzGEAAWb0LL5eTCYzYRpXb+oKD7s8HBkWrkxDKQhjKMHK94+1L1e9eza
9lmJhwzg9r9+irB7it4CgBAkB5ViNzt1CBbseOokHHtuniI+3+5aH0m2jfEBgKKA
N4aCDCjzXkI4liNQDWX58M3Ut336Bq0dhGlOrf4EVjKgmdxuqqUbNO5jE1oTDNpb
nKi1iSv/vV35mFT4bhJqoxhFzuDv0ihvHe2ZUAQv5a2EPzIaqyduJPuXxQjbBSRD
Vkm7oFetLFHw3zPbP4giogNRVo76CWaPD/AsfW5f4VffePGZiufTtkOu0f1Y3r56
ZSE3mU7kf5MDv8Gd91Wl069QBlsWbjL2Deqek4jBNBPhzS5s/WswTaNLB/5C0w6i
x1ZSuFMJNUXhC80+Gsnd1g7KhMDSJGiqrOQJCRAxW/aacmLBH6RrOTwVi0XYdCmw
0rzgb/0gPYTd0RAcFIn16af6uNgMMw2q4hsvSs3Iz/Ba3QRdqmeGufkx3IJ1JSCW
ZudQ8d0Vd2xX46q/WvWcthFwT786PUAIvdFuUjMUf6ykvRCJ9Sx4fypRiJvVMYD/
sH4HND7YE1ipljN5XCrava5QBpS0Z70fofBNgId0grSXGW/Z3URD427LSZ+7HMdb
yUy9eekGC2VvfovH/yD6JWtsxTFuuNM6jq2vHQVQkGwMtnbMmQUen4c1aHJSNo3X
a3gZJcWLn1HTsChq6gni5N5goHKy9PUAeSIo4N50NzWpzWsA1FyQTdq4bjIuCEJ6
L+x+BrtyLR9zTeks48H/pQ0xXFGy62YnX3XFMDDitTBgcZtrBgdqF0F4vLVZPiQU
iXLpB9H5dtxEv0ojfDyD4SOoMZvUyaFlWrnPu0G6Ac7FfXI3TpAazEG5l0gdv44h
FC11Gf0b6VQIsTPuDzD710D7I3ykcYfcTd0E1HkyGmXjPWH4bEY2BnfgHRyAYNsY
pwYMi/ZpeMsyuumHweQ3o9uwsKC0NIC6PDzX2w83fQsREKfLQXNU5wVOeimycLde
ePyIQfhSkfFN3cmPGy3N/xFFgtKrr+sVqjGfjZXRCeclBzM1QIZQl7SOB76TtO/v
vs6rhcujleXImcZzxloviXwGM9Oac43kV5US1B5TC03q+D4aUq1Fi0YHaFE0CFsa
DA9mAwqLUgMy59+wrfl669EeFjJp2HyfH7PTtvmvWxe9hQBfsPhY6VRNu7q0IZZW
IRdXxjaw1HSsO/pKGfIjhzIpgxl8O+GBluBUNQKh8DQooLVoLxwhl4gOttE+V8Fk
8Pg7mpJEqGnJQOe/SSxSLbS/Xjj5yE11l7guCA4G9VNO+Eay+WB7jDpjCNaMv5aB
6RtKtqfvS5hqi6X25VfhGludnw+W72FuKmikG21QFfHIUM0QvzHU0MSs4SNah67h
8MyAqUd41s4nQD4r1d7UdV0ptO4+H0ztmlG522JuhvP2V38DUUlpwksT1LvTH/ad
MUXuv/quDE9fm6xw+evpSYORmbTyaNortujipTQWc3D3pxJmvDYm/P9e5Fei/PDl
BkHegv4OZNSeFf/wCEugZaHqrYxfwx1YeCW67G3KqhoPDGrIOLBAuiW1V5Ej5Suw
Ife+SwTnCSVgOy7UuKVcZ2HI1gc47lsxBbVW+pnPU8iunCpxSmHOUt5th0d7i+9a
MHyfS6hp0QMaauyqtsp5jeGqVuryv0u92s8oV2J4Rc/WY60AD/WKCZmovisJzlCw
AqSdJwhn9e3+Ti/W3B0cb5IyCdUZexsxKwzZkv71lbJqTE702xU5Is6esiL9koGC
rVKb75ikE2c5zQgh6vZjxqOqCdqecoQU1FydBt6NriFN71I9HjW5kcRr7q1nDIWT
r/tQCyENTpbQKpCqkAdgVsdoFySZTzFsQtiDUEEbUD9uHZSuCEd+t4lG7lHskMme
164SoV0rymLBKDePXLymuK4SgpmmkRAL/xDCAV+ldVZMtCRzCrjlh2uQhCWrg3Sv
ZM7nFRYnhzF4v/Pib2+FZZBbcTaazryF6UR0ENriGxojfFyL1hVXglh/0DEeXaX8
a6G7UEHgk9YBghYzSE2W44g/mzePgzh8BZuPWqw9/awFeeW3iay/WrwBsflJrTB6
Nh4qAZWL097Px2qZWs+je5bTQ5+W6ZV/Mq1Ds6CZV+Kfa+R+PUiNOj9TeV+ULRIF
zJ7ic7CN5+LgN8MkCNXSjpReysnipZCl95wK/MVsYbUkJlEQ9CJwmIe/rI7nvIYt
L6ZuRBTtKc9gEQL6gvPhwwc/Jr5PzvxFm0RJbKop11hI6oybsgyOt6JFfX26KwVr
s8MyDd0/U8mkxhtwqsUXQJJMlL0ubMzKq4EhhIokkjxe8y8vPQWEr3eUjT1Je4Ci
2BNqOSqmueAP5jGh9xKFnEY5Mo56b5pSqiJ720eh7x5996BWSHbV1CcBJMgj1C+X
f05Pwg2UWW/lD8ppnVCKVLIcAQonlDfbWp7aCgHdLI6d74dSy3g01YeziyDbDK1O
EHS5WZ+SC+ApweZANerH7GkLn6aFfXWAM5ny25SaKxSQ2RHCZBuhxXMjTK4vj3ek
3PUuqslnk6SjN2CLWasY7HNdCU0Bp3My+QHfMJccyj5WsARDzHCoRNc1KGSc1//A
h9pyqMCY1aSUkDMbRYVhXV6SnOc4SZPVFWag+pyowUm3uDjWcWwngqTpnBeW6RQv
tGq5UElNRisaPA25/Wm40b0I21H5nl1HpMMqqtedIqxDgQAeTDKgmjTW61kYF8LR
J9QfK5kycXrv6m067E+fVQ08ncI6y2n4kNhlJEFnc+goREwotKkPpywtsIdDLGAb
24XIN/h3B/yiQZr76GA/bXhCozzfuWQ4fOgb+3mjB2kCcONxVtbttM5TYCVhlNxe
XnWtTzM8IEun7XHEBoQq7Iw/jV1Xbq1znaljj8+aTGMxLQPPXYOAfZQW/4/OLaTO
yqsBLD8rB08DdKx0K932HKeA50uLgF8h1sqgwHj7zpb8ab6CpWtR7RJ8uFJbcYyZ
O6Frh+f5thzHTil4WfTAF6R6EX1N4W55owd2JiBTJkKachXiwxD0O0r0anvDWoVY
FFeh5WJtZo5DBdkuoeID7liuJsrn2GgZ5picDm4xkpAndE5mlftVhZe6dB0wMrfJ
oS9fpKqlFMdZbcM4Jq7VwGRhfX6xoO+eJsHG9sy1nirUjQGVPkeb6S5dSbG/G4zh
Et1p3f0bYMc9liPsBSH3DIjOBejiFXhn8QZCjMqrcQYqOZdAR47cUw3B8j//sqgN
5+Kzags1oEuvwwsJVQ2gbVSK7WoTdvOiMqtsR9jVff0smNbAeUtQgPJ6KmtwXcUq
A84haK+iKD0Roa6klRhcG3FcUrc0sGgqC3EkPxgByA88onpeqlw9AqlvW1i/jqLs
4f/usRZzrUKupuPOJFK6JWKhvxjrw355+oaC2hGInQDzZlKgzU4nLyT01scmUiPj
OvJJLFbsG0oREBf9I82r5f095DR0RlgJi3AHgeER1B+syC0PQvyv10Q/opWSUo4X
bILqBwzE4WA0waH71/wt/M5ZDwHByRrAhkbaks7NZ0lMjfRXqnWXezefTbn8DlH7
CfVuwatxPAmbvyJ3s71mP14cbxxeLFt806Qf47lHmyO/JiWs5GOt0FIAPe+zDX7Q
2QjCBGew04UVRgXLZhQkcFp95tuadsfmiQo0iUQQH3YLIyqwYw7hxj5waTmr0Ap/
6Qtznpoy3TDqc4ihl2EGDfDbfC8jMcVE4n9WktCTTvcsJ8/zv5IvBghzKIxFMxBR
v/pyAG/1/2LgSI+/GiTX/RH+O1Th2bbHer+9gEq//he+c839zNvMSvMxnATkoM7y
+25gDLhtC95Tymm7A6lmgntq4w/UxWMg+Jy2WyYca+dBD9Nqc5oeEQKGwIRLH5J/
78eZwKWCUKLhkIS7yb6tcTWxdTr15OThw/cClJc2o82aUA1aVTWRBlN7uxK3kzNO
K9OXnDajxkzxJyH7Q/T3jhZzZSVZXtGZ28ejVFzZkRMy8+zHkJg5sT0QR8rwYZpK
32/mKWcNoPMbf/HivaIWReF0edfypFqN2Uq5kvGi/RQE+siZGl31gXmaE7NFqvxu
H/xgIj6dHeQYaJ2C3ezM4gNAgnDnxYycQt3N1HpwgsQGkNyxStlSPrgXUYZ7vyK7
/XYKSutdZmwKxhbDD22gpFnK/Fk294/fyTCWlIE2ukoH8C5EkRpBirgxa//KvltB
9K3QJR2FJFEHcLI4iIVznmca5TJb8PF3mAbXr/Pbd9KrwwVL2oUiQeBVwrU9XeI8
vD+QlYgwl2VCx5dU7HSgmUSALW3ki0j59BGqjcIoQ6geROqNt+ngTG4XlMkRSEab
f0GCnXdppJfljbBu36kXupBQvI/twl6sRyN4wIoD/XDheSKTbnMEU8e0iuzdrLVY
08Fg5PS0iCbKI7mPayrL3UegtunWeztlxgH8zhgEoBwZCFa0TsQEtFyKBrF08U6/
wIPpES8Av/PJE65IbINy1gMJRbk0uZb6vIpwg5DYgcYZTkZHgl8w3NF50TIm/ink
Hc8+qHoCG/TQK4hNZonwtztaE165joR1So5gfL8LhFtDL6167j6WCaTARcMLztt5
H6BXKY9qZ4rky+UxcEeZhUhpAusdCQ/DK3Ehu+Q72AQBEn3bEeLZhmwKjJ5RBeVl
JRO0QBmpeC8ccn7gAzrzJ4WzT+n/KRs0gqXl9k2NTAbqme84LFS31TWKzit9PzUE
2CQUak+MfguLpm/WYAsq63xV/LH2Ow60S0PnmPuMcEo+bUVd6pgiT3P9Y4v4TAST
5Lrut4585r8xx/ChIBSX4Zga0+4Okdi7qLsBF2urpRaiHiVDY83kcGWUSSaBI9qq
QJl+BT0yTwsf+Ib55xQFW4xa7nCaMBy7T6buPFvCIPnzv1H0VpGtGa6tFvHmFA6U
/MSAFyJzjuNwwUTv1Dun8wnjx0SQZU4w9aDssqkb8kTI7Si5vLdTBILkg5CNlN6V
N3DZ0uXuQiSaubMCXArWGVGn5KCZEjlg6ba8TJh1nRbvYwxXqkIMP4lppgkPbXVv
RQf3a91qyR+jtFzkfRql+ThiexQcQcd3ljmzp/Rw/YJ6GgLBhKC25pfcHfJkLP61
n0glcnOLskb9QdgD+X2Oy3Vovw75bZbX0Uo+mQxHzkrn3phJP3b983Q4K5NUmwLv
OjdRISP65BGzR0Xn1a4Gt1Ju8LjLLqGzRgcVC+fquB2bjh3q7tq/vB92v20hvPKE
eouvrVf1undcSwrYo/0CyQkTo2xweT58UX9n7x32i4mlTFynW3Sv8jwFe7vXD7TZ
+v4wpx07iMa8VXIxIekOhnciOC5fZ32GuDp9JWxZFcmZjzZSIbwAr8hpU1quLST2
i6r9ePvrd6ecM9UjRO8jkfASlfzZHYQIlPHkOWHsTf5Bs8iglectWUUSpjM2ajop
mPjYDOTCYkt6fXYqXjXvbOZf8c7d0/IQ8LqTaG+Wc10Vzxz6e8HNf+SARjkrqSOP
ZbOmL+50AidhCCKHPxcLnOchxBuX6+USF1YgPxavoEZnpKxkSLAN3pHGtkA0QqOx
nEVUe/uFZa0J/aAXJBu4Xfai6hkK4+oU8lpCbZBW4WdyAyWg3IuZmi46ohjvECon
trGTRQXjXpyatx4mgcRz5c2GsjQ+uHugT/kJMClXdvAI4ZrF1V40+vgiQEH4E0Wx
eav+MR6IWIe870MNi7Kk1RZLGRM+Bl08CTeJw0gGMp1C3FRryRWWoIAC1djhHQMt
mr/jBGX26+z+TxpkZeLlsb9SUeFu5651Pejf+AUXCGzMqr6/LLJ9/0YX1TA6+tJh
5LLf+9COqlCgdCPm+MtlSaBqAOrZW8v72InKwMHvy5I159mjVOJ9ooc69IU5GaU7
G2OzDDUMuIQIOmClmtnQv9huHu6odUDXzGvfjXHQfjsmBEGeQgskUOeW+P0YbIRt
5BfMMEmK7EPKmBoLF2BpQH1WHqj5cter7EFJbccgJIRRP3XXZ4P09huFNBUULeEc
YtxxqMCebuDrOHzSNl5x4J3icgTZxY6ikzwLqUNNlQ049SEgtRC3QALKcsvu4PjH
7uyf3qp1gxOtLPDs2iV3IIFdhWvxp+ZjfF3NIH/gMjcYEEXHpymzcUQiIZF8zM4J
I5JpJeMrlFrFTOuHUCxW1ayIUin7fPDEgMpk6WS1z/1riljhi/kjqPFNgpwxA9bQ
BUMULF08IaXG464m5thdIHKjVQPOQL6rHEAFC3Fiw+FKc7DJE6qdeUWC8mcc5VI7
lft0IMHEQbnBO5tkyAAWqdfkB04kdoo2vswwS9mG1YyE3GXeqmliQK5AcHpFGt0o
rVEswND5mS4ifbAjehDPc2DIzJRtcVOFGqex6MzOu/Gr4Gt+KthiJZ1C453JtN40
/eE03ID1nTvzWS2z4nj5QwYW0msp7tWnASZSz/5pCT5qCTCjDwdTWUr2f1GN8FK1
c+VNnN+BxlWDpw+YN3CERPV9utBxTcCY/qfV79xBsXx2pT1XEaEgfB0Jf6yvE4xc
l8GPtxW4kG54RgK7KDWJ0ObYE46mASKQaw4raHOVnjXWxwjOHVRMvV0Ik70lGOjj
5ojCjbg3NB1HVRMd162R9HIQxs6R5NmwIY869ExLLzT0WYOHm9raCap4os2bpp56
u4tCyADqzOkJTiVfzPn9kvj/6TDxrFWJJiTJNfQa/4rXBMCIOudZ2JIMsCuGchuA
0W7AEEZS2n/1QOy/1pfJykUOoGLlNdtfoC+t7rkJnvrx5y5ZIZURI8TBOetnQ2dv
TAbvDa+v77iZ8wbZiYaQZPAdi2pLUPuUd3iIfCuXOXL01ufkSnmXAEg/USUuB2/J
C3/qXXLpprnoZHbkEraM0H+r+hZQRS0I2DYfX9xLsK4+F06Ll90ItCQpYVS3qj1M
8gbRXXreBkXTYMgw+8wbiUT0e7Y307ju9yS8atzpVYWpPzCxt2updTx2GiGtfz5q
rYUhGBblfOZui3f7bowRfvsIBHrjhxIMJ+pA8PT4uv7N7QExaYchC6sFz2YcJb7U
mzEssStmHMm8QKtp6cj8f5J7Qbg0qwreALNH20agFQiWeZ9QtBGfX43mavu6vE5G
y955VzfvtYmmQMVB/UdtiIU+Nwrftels0hp07ODkDNpeNDmvNp6mGg66mY7fZ6M9
YgdVA12jp/mZE3Bl85zGbbRb/KEV953LekIlu5x+2PII+5bIEmtDO78wU8BC3T0M
3lMo64pwd2Djs1DjqQA6QjZJLqmC+xj5y/MmTMS+QHgot1nshA0vQbfnhRqlW+XU
bO9EymkrRyrZ+9U+H5UYpH1yLsPs+6+26/ugjf3pbPwOxCxAQchdMLgJJV0cxHtU
tw1akdZXSQlm3GfjqsAEyGN8/A/P3nP3WGT9OioWSL9irnXoZKUFbjkENV2r8yfW
r4ItgjYQDXgTAn25MA51S2MADj2I0yQa1A2RkTb5J+sDFgp5yWVpVJFscLiLsLlz
v3saHdrpJiMwJsBHm+wjGOFoszy53l37Cn75N9/+imgOO3+xE1LxgP5p8MslpvS8
P/RZfLf7DJmbAnKbp3uZhZ6KaiVWr6I3Q2DXl1SO3/EcHeMjuA/lLWgSt2hrA+u7
klCPlkSxsD72Kgx2xaMh+1eJX8zA941Yr6pOHCaUbc0HE7NjUJyX6rca9zXW8IG2
XXbuhIl5idWgutu2fBZ71DOlxIhsF2zg6/nbz/L+0zPTy7Nj80TwTNvuKgMBTpGB
ckHlvyiHwxTZeu3uBXd5akkVJjKdNWOZGN6+xjtoRPAFwADlZU4W0a2tGBfjDI8+
l2P/7JGbgGNpZSyYMjPt97RiWwmekxsHvVHm7xIbH98MErJytB5LaFYmfascqhBE
5pMYGCCx3n8Y5RGZrYLyEO5G35nW07XWSkQDz/XXbgwQgWeFw30wSnfV2H0LJzmY
VwCZVfyn/Ftmoairj5nN1gslvMygKPTmghXzJI7bX+E5IrYoJtQ5ohPhFUIagNFq
fbQQg5RPSjmXGFhrCbBLg8QhmsDfIi3cyd6gaDn4r6QS8/0iVR/DFilxsGVXJGcp
CT/EUWnjANnms3xGZQFvjuVTq70icA2V1nM8SQ2JkNKDHaOVDdRtZO9iXpQVr3JL
ymjgUo7xO7EN+Irh4QSU/qy0NV9h8zqnpJGSgxyzvN5BUUGZ+kMdFZKc2puSjznt
6a3eMWPhxVNLgyv3FSgF9t+S1f4EExg+P6xcIAVpnkT6RBkQUHEZHNJ+y9FBnZZv
pzCAgkIEQMpVzjjPIUFOdt3N2D7y3/nqEL/rA1FLQYcZcF9i1KQ3sc7x75ipoCqj
8c1sJ5FMHT/7Usie267Hoa8oChsQ+NOgV4J1rb5pP8adPcPmMoDgFU43NbN5mNkM
zLSlIU+Dhw0y0AAUrffBvvZex6mxwmEQOEsePe9hMMpxy32WUP1c7RD0iVjK3hAW
FV7a/7m98FgT6BiQI/F3oixaLQD6lHMHsZrKwrYLcE7AQSSilrXdCgkGUsXl4I33
cQ3qqYdXDZlMn3F/ImIH+uOcsQNwIzukI5c6bILUxee2xPoFfigA4AgDKoQt3WvK
P2dAFVd7adKJnmAu6a7nKiRAc1HqynF4exWP7qo15ISMSmbFa6lnZTS14+nq2EjF
BUrWPoeeYaKCYqAYfn2UBBehSd+NpYJIf81QtxpBedG4nvGief8f5IT15dzHxgxH
ZkDz1kBVm6/0AzRK1O1fssDlfBo6ZlLivr5Sow9soadniMrcaF4dP6Ch8I6mmY/L
OKSxm+Eo7REcJKw2V9akDZoaZ5izTHKYuk8msUgt2rdxh4f56yn8xmI7XNl104ux
a7z/123sA6hd2Hy6E0IRmgsMEXujfp6Vm2PHGQlRwKRxsOkzGmrq8swYFay4wC5R
g7979NZwZb8CRbpAmUrRSDlbjx0YgV5vFaFdLJ56IUx6sBhn3eAzKj8l++qXDBoL
/dqponTwj9007hOtMpEfXIML4LUqkRXFML1ImCwSoFaZi/MoD3e7Uh3pToqiaBcV
2LGOvAWxLKPBz90REOMUs+jvG7RHNhNruJr292hVCcLIB+8/BMlu4bTy5FGVKhtb
n+o8snjJNGnyYo6mjbzl7O2hK36Z/i+TQzUEqrF4BAeoApXeVKpePeOKyocHKz+q
npUa78vknmg9xRZx49FfKm/HwQ2GZ1UJKF6iCKvllFN47qo6YqO6BASjTY/tBK9M
BpAEtxKjlVldnKirZa0ZBwYZaIsIl1V9ph7t5y0Ado13U/GHSnzvTOEslVJ8KrNO
QYL8KkNSPIf9bSopoRBZNWFZ3/NRjAwr5Y8HNzUSnZyDdQ6l5iDaRSnbMWUYMJIi
kDQbZvtQglFKSwoCQ8PMMjBO3kP0/YmO4gAzdeKecPtNw2YNyKA9P6iUEgs9JL0B
PnwGOwbDiQkD7o0+zFZpuLpQ9fpTgTmbDllRRko3FcH4qJavExWgbCaGhpDBazUx
GPHJhZCO0r9Pb7J0Cfe6Xnqy+I3P+p63AzXnxIqs6JBtKlFPZELTs+euzfNUv0Js
U8F8z0fo3aBjas+miSWXsVqnnlueXkrLMM929/vUPuNX1Uebpi5OusNnBzUZKgr5
J3eA1rV/RM4KdRBPznvGt3OylD5M/ms7MptBKlPjtAlBCotvs3BbEpYZmrPMfpqP
CBPWCwOIkoLE8GyZtSSbV4GLqP5VnS3FTw7ITRvYHuNlux+o2eUlz0k9QledN0hY
MurfeHCTCjTaJMk2PckzVPwcdr1nv5Ye1A56GELoppJfJnv1TneUXzuWQw0AUjsO
T1W27RzFOJ06lRoM7SYAEL1krCtChSrjXHWIOVX8Z6aYP175wkGtq0N/3/sNcwg+
6rzU690Lw9Vw7OouMFFzvA3u21SlakhSD1hmizsiq+SeN7uGFHpJCtFB6p4956qb
qs2UPZgUSbf5CcEhAIfJ1KgvdXI+GSv/eVqwoc0mEXz689G1vr9ek2MNw/z4246v
n4A6aoIZUUC6m6bjj/LjCZtI9ZMZqXhaMj03yv8kd1weAhnN9ar+uV/rTTqqkFKH
T+0NtasWpPo0KRMSukg2wTX6W4MwBqkzO0YAbNlRpAv5Vy+PAxq3Y1Mc/fH0pa1t
RSqZ0cNN5HdfusEe6H8HYSdhCoKgR8DN1Xuod0gg7CNrYEJfs22V26LZ3YZoZbg7
80MCt0LrVduD1xpEZnj1vDJGZKJQk92AM3wFhbuPEnlp3Q2Ee+/Od08Vb8GWi7gz
gwPc/0AeqDXItBDFvm5pxkFfd/FnUTjybRmY/EQje0vESgGQS5T+bGOgotG4oVua
nf6TkkCDhmLkpWsUxNEfdInutWH9eARgkXQTQpn2igl/TVCq9FqCRi5TCRh0ZfvW
cabBPvLF91Smpw0kn4KYVkZhWXqX2ILzPt5JPec+8LqUUSdzVpVTUURLs6wfLj/P
2Nk4TGY0Lw2VjfSGaQpYrSSnuBR0CCvG394StQIbvRHNz8uGzKho1YuzcSnPw4BQ
8qV9+QuyhtNmbm5ErSVDD6cl8IP8Y4da5Ey6zIJCOy3ceihU7atFykreZFHcQvGV
AYJ0nCLLvvet8bbSYZuuXisht1Tp4fv6HeDwFFoY9e9WtEAPR4qIPh2h4hF1c7nb
dXyEuT77JUVqA4GYGVch7SOXo3Sy3WqsZizqgSLcNsXZJk5ufRw4bqFy7cNF0lIe
EFHKFiiDD7CZW558DUi/4u7cjSfqEAJC0H4W+eCPtvziijm2G0+uDwPF0sFwszxg
aYhvWhX0wWvxqnm8MZMeCZxhh1saf6+c0+HkWNPNUoT9oR/bO8kqVcfupULLClpp
CHDXH+9yWMFUCS9rjUQNnOzHAO0rIuq2/TBjiHzfUIFoLuQLhLHBR+JXDuBpZ/Mm
0WVxwPIh2vJ9cCad0BweiuHA5KVrbJrtrhIgfoAQVlDx22tfjGGlB6cJFH03XEoi
471kPeFMmq5uXjuvsPxHjgwT9E5B6p7G+hY2hj3bXt5c1LfgwuQX5f/Rb7wQ3bQI
GXBffq1pOatUzRDyfExbNQGJqML5NJqgJ+wSfiO3Ew+T2sMyjriUCs2Z5XI59cXO
AnlUrdT4JLVWMADJAcerfOLa+NcEMSihRmB7D2GthgoB2mXPbcmyMA43G00w/QUz
dpslY8TTSPX3z8xVKxPN8lpLpkqAj0KpksWtBeee7a7H6XdUIHedfuY6WqCYvZ9h
L8TSZlfofELP0Shl1rJ7C++tzJydbhF3Mh4pQn5/+oTcq8z0Gc9w2/jSLQQySb7J
kU4sTy4WgNg5TAOTZqOtLyGVLYuOlPqEZknGBSZqItcXf1HAVq9tIXyhj5s6sB+4
4K4gbMRC2U3SUTTV6AlI9szDhAsTQGnk3bkqsOPeEnOyL5IK5SNmE7n4qGpyBjCs
zh+jRn+boujVmY9eEzeygB0HWjf2S09kfoRHLM62OkXDVWkwImSpoPgniK9G5nc4
ZyRhrx7LXfQ4anhnhjzktvp40b8G6b8oaVDJYr12lCoJPYhavv5XpKEDlC3eJ5ER
3wFiwvYadfpvAmvSOAy6nQiJWu/Kg8Bg2qZoA0xbHoLcRI0CS85cPYP2sOws92cW
2pYgYZBbOS9ywyj4+JxfsX1tUMH85ztt7Vh45OP0Fi5tDh1rLKHITuwe6o5jjLhi
YlOkMdfIHsZgasaKW2jw490sNufKO8rtF58dhybTQtWTrFaMaCGquya0AIHJXPdI
yOSJoiUeGwNV1ybinJKCXW1XRzDNx7IXeWqB/xY6c+5XOnWwdV7veZOSBEwUF7oe
viIO4O9c9Wr1jJ9+6y5kCkSj5ALT3otn+0s/cD+CV6IFNqW8f6ODq23fQSdSKJ3t
ZcaZcuhLMcL8z8Hk7RQuQ4Gve9ailU6d62Pdpuai5pTZ7MdcJSBs6Jnbl4e6/DZr
rrDRekP7RxyVyK+Jo+YL+Ft6cFlUKI+JbzkQ+vFLO3S3mzWtNcObbK1zx1AlIOMb
pUIyeLQD4MXrHHIKst5dQwIWjq58Lz2pOK1EQjLdU7FGmDx080iZgWJTadEAl4AD
tTjpblf3bNbp6VWoGLASxNOrMZEXSgPgbXDJ31Kyl0PpXfdkCugEBlUxYr6ODXXo
DoFPNZF133i9Lq8Yo3zOjgD9a/UGzvWHdI8RjeMf7JaTY31Iteqn/GtXB75DutNR
W2slWrF1YDvPFW5puUzmQeeDG3FOfo4nzH5HkJG8cuq/+R2B0COyzAMagAX6Arvh
qofRloQvCxcIBP3pTZYFpHRY04urAlTJlkUToflSLdCXPTewf7qMfTP048uRG2DO
ajaaRXxwU8W56DV5QgMI3jzDWGgN5foyoRicfyBc7NSzSKZiTHDB/crKpQySMGj3
AgPrvdo/saoMtCcb7JeknFQjLysaRhTJSlZfs7FGeVXb1HhQzidljGGWSnTSwKdM
qP6C5BRqX0LB33NwhOTpaTShkByKUcGiRZX/Bmk5s3BYndbQ/I+GmWIA6gUeP15c
ZMvsQkhKzZ3YL9gSroXc3IyfOaSIA626GbF+gwm7ztmdfQYymZ9ccuRDAuvjL799
N3I6SIbRQ9O6f579UQKd7sOm3/G067T9AUo27Jk9/72dv31WDTsHZzMj1i8tu1ZI
DpyRD8UnbjTBF72JaCOmPFwbjVohpid71jGXQrNAK+njfVhyG07o/ASfyX69VwOf
G0avFE1rQckhGoAOFE0+0NSksi1+Lv/VGhSesAvURgSz7rtspEWpA+3IoV4+HT7M
782NA2znpwz+lZVu69bU4PXcMU8MCUP6GL+0nuRP/+g8x1ythvU2M2U3vELsFd1P
IYfdGkHO2y+hMTxHHZ1gis1tyN3cpzAja+InweylmEpBAXrQxw5khxmM+8CY/LWV
VRxEjH82kjwqLqQzEr3vdAs5Gi1/v+htd4a+4to2i137NfUb+WS8NHA9ZuC/bzXX
mzBVYr7BNuHvqJ15+Hazmzy2txrfC3r4MoHk2wA78MJOFbk8Nw2pn1pUWv3LZh/K
9weB7nWLe44HLrAY/IHDSJOGeictOXymkBJyYrSPnQvAjcWVhj8QeFhIF0CyDIlv
1mAOh5wofQtEq6MohQiYn8/psIzcGM+6EBHlnFdB727uosXnSocu6PdtNamfqAuF
MgZIolmv7plxHtQl69G+ApvOroMplE5JpMxRf65oUzOAWVqNW7c17X0GwvV2bzn5
vDkVXlf+cputI3sAmQ9GxpH+RK21ALSGMbu1wgW2ISK6+ceaXbBW1H6lspp4BbN0
2FFxp4T1GCh/UklgkPkD1oD2Gpc0GhFuMvKd9EpH3I9gBtBD4JX0BkDTBO4Ys4xY
zUnPaFGAVmDoq5S0tn1X/jgCCkiWYnYAXGLcoEBMtACo6Az1wJTfwYkKWguvlgq8
XSnx78FIhDlpd/b9M1igo5OvApp163nuAe8UvDVA4LSQFTsWRNig7F5tqnOjgXV2
V2y9J+w8pB2DudUf9luOkF488URj8wH6ZYf8dUdk1ZHYOnUxYQWj3LqZaUi6WpFO
TX8mSjcpIBlyPtyrjnaY5kU8G0QHnj5REfKh3TGN1UzjT76gitbLE61J+O93h0v0
2xBKNhYUs+55UDTc4YyWEjatL/zxxAuTrwo9bFvJjicKWxWma+h17L1MNurAYkOF
d3HhD7EoRpNd4GdWdgrTUzFzEL8zejYMRZMbBYHJorpkg8FQ3pq0unBf4ROxFUFB
v4i0AaoqOM/F2B+qUKD4hj/XR8P/xul0J705yaG05moM/n5uMGTelq/m2kxPU1BT
GpRTWgukcP5ovhTtiv8fP4nfvwDpANTlHvxEY+5fW0xCVOpptHq5qaneMUKcaU4H
AcF32Te8+ViF8Kk78fzqZPEBJ1EBKM+tRP34l8sg0tQ3dxt3Iy850tIu8Jw+lHcR
j6fH/IS5tqdtNo70yPsnmiVdcpzA+lEYCKP1MmOjsW76A0bAKvuZxLoNCLa4R6LC
cWDuPTqk7JKGszWYXNe452oJ6yBNrBV1CYNFqjIR1UY2G1b54LSWm7PLHhyA5Y/b
YFx3ZzNq6gN5ThXhosoGrJKLOxFllAo/tUIZQFL2IFUnBE148cANxcEg+p0LyzDt
jqufaDdirBuAFWWkXAmt9fvww9WL+QH5YNuU7ssGb+j2TY0gZziUuNyTQKiznRXx
otM5F3kI2FqY0AdboXI2gTyKkgL/CsXrt0tcF5LTKX8qeyPTHybuiw+d5rc3vP7j
mu66kVr5Esp786lZjfGrtlQ0RvKb3zr/e5nGuGA3mgJ+V5XR+eGXNUPbfgI9XNsB
KRPWPIA0DtqWJ2vhvZtYFWRp+GxsMdkSDQzJ9r46o3k2jjiX14lpG1q+GHO9pzfY
1BkHMF5eGr0e/PEjnuj7L/Go0MXDE1/Kc296XXxqgieqjfsbT0Uy5IrjKOj/PTuP
YquoLl5/79DsDnoEXgn2Hre5ati0c0ZPDYc/njS/B2s2ZUxclwWjuPw2V3OpIqT5
h1PnNSZe3dlDeXU+k3GQnD8D4vY3djB5Vbjk+hYhZW1PwdI6Ko4b+xUZ+JlBpzVX
48dtNahqnhgYpQ0164p/m0QUK6OiCNJA7t3g8UCopmdb1UrxpzjTd0mcIn75VkeI
54lNnfQbnbL39O10/fk6OYdb8KDhVrhwm2hw+05kXz2UabN4o9pS+td/1kcFEnY4
2qtMnVaxmPazX/7n5aDLLVWja/HEbV68jmnLldauicuZPivwRs9/mRNPCuU9Xl1I
BlRHpLDd7XmqlbSBoywLfh1wxn7f8dvnwtk9kclq8eo4n9/zcKJExB48LIypNjlE
2UdKo9gALu5NIMnS+SmWQ4pEJDVYOvMmoj3KInjG/TLftM2FZ5XYiIhBGkrIQPP7
iEpC0durBAL0uIGo1t4xz8j1kufC1LeMtpOMDnLeJ3CCju7HCNkDSlK1Tm5BGaYv
/K7UFDwYA8rNXRaZ66nfb7UKYSTwzX5voWw2Bt96TeH86UYwvZnRqRxAagKyWptB
Uw9rrx7mq5zkiFKWgnv7zROk39eOMPC9zGr9MINntyChhzGLhXJxkkc4awuCZAyb
FJD+jHoPxdwMqKbvas12VLfGCSMi5GtxtX/cMj9lF0y/IIdTedcPliGJbYxv0NLB
xETcFo1CXXIzgPW9oBCEKdkOj/BeqN7u9wxrgIsY3vZHW5kz1Tv1JVOUVxMD2BSx
7T6cXQ1WXANGaSLKnAkjnb4bF/EAdBpFfMsXreTUAGSPYfzY9Bz+1rqOMSq3cAQr
UkSCf3SMuGRJhgDLWG6Co62gaUeyHFv4AULPmExFOV1Gyozz24zlOseEztwqA99U
UKyWaPs68urQyufALXheNsrC+toEOf3o7ngVmE27jwEkOYrLHGPXoyBo1Fn+sBsP
g0ALodo5u//euwC67G3axl0MvXVlKaSQkSHPsLfzMn52tV/cGbZA3rSMHBamj2Tf
305uazoGBW2ao55US4CkSKtnahpq+d/SSZ0eP5+Hxlc2lAH3UHOMTeLeCa7aj02e
T3vJ0x6qxmEawn3s9o6JvYhzaoAgDTiZ0C0UMUeqY8Le2xbPBFIthlzxgH9Bp8DX
r5+T6EcnDbr98CURHGg9xIdrphQJxfJY8TYtyqJ2IhptjpqtdfLkh3ncf1AXEZAr
BZuk2MpUTI6LmOVzT63v/6wnE8YuQXCic/n2AbgzLkbZhaxRi4UFnj/uD25JSgm+
fx4QtsUPbKC1ZLLM64Ziv82ydMoOFxd1Q7BQIdsiTj1F4u8Fj/AgJxYMbcWSW/Li
omLpFPetH+xI6uhareWLzw42WLvg3Zm5IpSqAvo8zVWGrxRUqH/OJ9+jDuzfDlXQ
THM8RAaKco68QPTfXrIa8hx92TW8OOd+ZF++1+iVkN3T7iaVIzuFXNYvcXltF0rV
u85oNYGd/7pD80ScQrmClX13so4Xm+KaJRtpS/74rZiFgXohzGgvfpgn9zWg56jb
1cbZRYHgT6kjUONWx+Ksfgb908kJuk/iUaFmsVxNmnU5cY/5Dw1OSxpjmifYWHEt
L6qIQGo6oUsqzUw9rKKjB3siNtm/HpjrTpIwYqSsH3GzaWwPgGQx3sQUHap539Tl
sHZ6IBrTcNF/Jh3Q8c/FwgWFLh5L8jZ03xrVj8jyynna6qmJ15aFw8K/QNTEk6J2
Z9pZUmPPm2iCkCJTOVI16Iqv51U+S3k+ExTIAmeGUc9WrJyXSVQAHgJb/hxOJ49S
lPAMJ/zYDcWj/KMTFB/i2sQvQ3HE90dhYIhJm9rmbvAozHGnD2DLBql2ZjcggOVZ
Cl50z5icIKKT8oYIJ6kCc9wnf0dK1mFPJ8nvqqPcfwMI9+48/lGWt6ookSCF831x
OzgDlo8tOqeiwxwgWRY318DEakVn9gK8wHLyfbAb1y/hSS1yB4WiibWoW0ld9JB8
K69IhwVJx/Cg8KixBE9KvO5evNBPpL1x6mnu0mbcwAPpVhkeLe25U0FwNlnVZHLe
PgAtInbSZFPIDybfhGHiGtT/I/D9w7386vN+boEXD7lpQfPqPvN5iu5faqSx/rV7
p6aDAaEjY32AABMCuJZSpvA6bVyOt2an/nKIc4KTD+lIzwo818gSYR6fKgZ6NEQZ
Dw8MuBh84Sf5A8pnH7gOC6AXI1sH5OLfhcys8rjcQbc/cAID3Q3Z4ms4yKf9pB77
ogLf9RvB7tnE4DMOVhPmduADwCUbXZs0OfFCQwiJKcwIsHoBibWwjuT9K4Rn3wRt
R+W7h7RcW/QfLul4E8zOKAzTf3ljQOFjaEtmp5fKCXiKpsjN+D2+dta/oJhsaawe
niriLQAzd57OQSS4HKNZ9zW8DvCShe9zEbzDXGz2sFnQegAKOUGxkWjurkYrZPDc
K+OeRXM1qFPB/R8/dOJTxTCEkDdJP++6dvesZYuejbwKf9YP8/uq1Lw/FWbFruR2
qTUqy2J6BOXdMbl+o4x15n+ChEuYYMZicgQCLo/7lfHZ30EmG774HWzbo3hhhxpJ
RrY1mNh8qUu1Fz2MdDa3KKLRBQfbDGv0XS6rkZc8wXtQP8WLz5DVBAI4PJeyTFd/
NUpeBVu2nfPPLn+MJkg1gqwdfMuycZQhZVlh/N3xWa7OfTLGfgv2zxodzZF5Huak
pMtmdwGqR3q1zLR/kXQT8ayfZDQrG1d2KurfPg6jzBBTGdDgQ1eVogASApYdpouq
LjcUpuQXvZHNeKQEFHNeJh50LvuxvE60wl0GAj0oHPlNXib2GRI28jfSiU0SGX+4
U/gnSP+rHFaZjAWrn5O/GYo4XrmoKIeapkiZlL+OIZlsa3xsHtY1UvSiJeVVue/L
rlPBzeYMpi1OTjDJMlXR7PfHLeS4/K1QaunGWmRrj5E40zP5jmsTdA8RkedHjOq+
c6AaDdRjYCGmy0ASObG/UF6lriWjMIunp+sbWoTGwJKWSEEkNiuksJkNfoeTWSqq
A4OVhwMz/wYXkgPyaitcatw86NyT6P4riwVTMzNcABK0aDlUmMTYLzcC0b3zBzNM
j6jWkSnJC40MwAHoSOWCNPWiUExnOBk1Xdfvk0hDHbOu6nkFCUGA3DBGcZV9mgtC
4e8iRe2mb7rPPkZ+OZSl1rVgx7UZZEK4rOUi1KKksk0THEYeZvCdP5j3JCDlggR8
VpD4cXrU2+PXDBage63pUILEM7RVLjqKLAFgBW3bvEOzByy0CaZ0LNXUhWiu1UdY
jec8vcwysYiE9NbeBaeSS/8EVOLnM+P0IBqRPsTsAXrsdMoetzwX0Cwndjm7g14n
TOlzj/lXU5/tUCA4F750DvG5gJU4Exols6MRVo75Xr9fjOJ6r83ebrqqOh7qTZKO
pF51zyQb5z1Cl6uekhbLxGoNzei5TdYN9semKsbwMxVfjjqmm4xpBDz3cgRJM0Yt
CmSv0lG2RrYC27lv8BCo08bBxwJPv7LjBq2T9P5FqNP0Zb6zGuTyl5U4we2n0Wfj
24zsnnqYzeJgH7nufCoOvgRWX5ZdOKNuzBNRKORBAf/br0xtetKBTSIo9yDGr5EB
pdIXnjN1yJJj83X0Ilwl936JnLG2azG+dTMsP+VXTCHvVxikNzD41xmR8VaoZEmM
6Lp7cz9OlEpKsTQh3u0uN8Fl6k+OdkcBAjj9FJMWwcpAxwwm/JhkHsG5o/r6uIS/
Fcgzuomq4pMRM6l8Mvsq8x7YAmaHcULyaajo4Wsp9G/GYVAF3YxV/eLwDXQo3ZGa
rjWH5UhHbEnBUhlAjyD5GSqPBBIYGLtAswtiP/Z294035Yq690RRBIFeskZgSCUZ
xNHAQseIwKwFNDq9PCPsIlKTwg1yvpHj1Fp1mpygFU2byKfnMivyLBu2eGA+xSgW
Vks5va+CfqQQLp4nrK8EwUhWOP/Fq4GUuZOyRDAwBqftYu6/7tHvskCSKZTcyD8T
AbQ+p3w5YDAfL+zRypkaa3jF1NY87JEK6o6mFgSv1fF8nTezvxJXBLlWbAurHDI6
YSJWE68h6nyz7bkVz0sUw26gpBFbcKfhe865tuCeeSovHnEk/UR8Dk4pWHg1gtOT
RWfYmkEnCubp8gbpj9XM7NNswD39LdDpidWDNHjLoDY/dBFJkQAOgsJjNHUtE9r1
xGyPeA5oBuqXnEVhaXc5O/UT0U3Yxzy36EWVjmgOX6z7was9BxGCifpmD3rqKKir
SI56ss0KyJDglynzCcueU320981MjzMaMRjZGtIml3yP4XV37GxCVYHFx+tWEQDs
Aj941Y2O7bCWYlVm97zyf0sSQ86HPfl/UCLg/0TMP2SLs32aT9/sFG5LhtgNd3Wo
CoCUmOxelNEu5ZYCqG3zC1yMTyGbBUhbza5VzfvxlGvVpMyJl2la9X+B+az06BmK
iF0eghKvWCxX/L45+XgXj1LhtgYU24rP1QLxT0yPwIRqI9Nm8OPD5qr9kZwTUZJ9
chHo+ByUPJ5Zx6vkD+hJkv2PZ/EyBmbv8MvjDTYN16UQJ0FCKJEMppcp22WsCLO0
4GloqfR+pzd+VO5R9jrz2OT/EjGy1h+ez5Z3+j8WkXEbdqC5Rth4KboBxH+bMG9i
n+Y4GUhTajh5U/Eum9y9zJ2kcvSVhvMYN3yYM3q1kVx/M+WooMJSqmfGifpOhCJB
a9TsUda8r7d+02sK4262Iry65E7sePqG+LMpDCqxpACRp74Std/k2Va9JUS+St5A
FeocO2Pwa9F31bj/tmVkCT76PATjQRfAi90O3f6ggMslaUTpQ+hnDSI45X1Y4BqS
FbAThci0H58l0e3deBITw8g2oROUIa7BRu+E+mHBdTlfnOf0ju+uWa61F/D6cDl+
IST8bVz1E7KE6N/BYDDT/eDJuNuTO8ClFq7vYdoYJapRm1VfRE6f2/VJzbhDZaTO
0eY0mzMxUdaSn45q3Nfpf/+7QPgMkgEo90TQi5HeG/aui3TUEHcS2biRFrPfTqrL
LxuVBgLDx/Yt+rDJqUPckuvW/wRqyi3OWGmrsZcrmfEgrx8rrnu7r/0SMV3RZvuX
5BPoBKEWWil8LEDRwcMb9288BiP5yaJyWk9FeCdA3ez+VZCeU/7z07qGCrx2kjsW
7b33HpSLvaRBYqZB+EFHe81i7ff/SApmjnkl8EzbMrtK3es8289uid4/VHBFVomh
/MHglWdGKfPufNs4vdvnjNja8pJsr4YkLDKqwrTbCJFgGjNsAYUvpHySJDc9e68p
tSBOUixdc9S82Ym97pSQACjQLB8nPtCU8k/1w19hraQttOoE4KBB0f2swI+IvLzi
iFEcTiL132reXF17dkjXreTJPmNQ2h9SsrDLeqMkSeT90q60K8tXT7jaNzd4r+5Q
OFzSd/lSh/6rtKHuG21PkMFj2pQ3rdrQ2KEdkGP4yy/Xa6WQVyqjkj86zRPHSFk1
FQb8URX+Ke8kWcr5BdNvN6j69NkCOp5D/0Wm6LdhNyzn+eiRGAd0r67KZr9BsGx1
jfn896q3B38wwvhp3MWMgHKhKbB6wgLmiNVSmHAMYOmm3+znDvBzfNCkucj30PpO
VA1W3ycZLk4bgsdNFNegwJ8ye7xAkAnGC0X21C8DZyINRtZ6BBxTzjKDZsOj/Z2q
fzrTuyyBCIIhhngT1kH53tTg34bFOHjnkuIbg/KnhkiNzMNtsHFcYx6OTQoSUw07
W09v0D0Y/m7pie3YPKRSMZsMSekbKKnlcb2WZZ0NX2wCC24HWKarJHAHKQtJyLx2
sIgqFWLGXgVghrW5pUyKV6qtq8i5p9siVmhnGMdf0FTfzmwCIgxETt3sYnyqIH5v
Y9cSsCapkIPSEwQptDU4PT5QbbZ27RA2lPZhTgrFO7kL3K8jJhwIpzyhYM/0z0ey
jzf8L746+0MKNWkhUpSvu1jbvpeYbHw3TDE9nKKqHkxoe/23KzAyEayBqsY5LEAt
QxBVmFhgnJWYrEBHAts9el1M4qTOCREwo3Un2A26RczDZ3Pn2CcyCN2bucD7n3m5
haA8NNQhKmpCvJ2xETgylDhVcbDpO6NPM8KqRUTUOmHIoWMjPh03TeZKl5UO0qvX
95PYE8oOenjYJTM+XOzOPYopc5nnBKUx0NXhwBaCfDsolC3adokNWJt7X08bFQcv
HS4ZZh2xFp7im7ipH6VUnppDJlMMFPWrjuKA4hPartxqZD6FUbpR4j6htAxa+mTg
Bsqrde0muhmviiIpvClLEu8pbZ++VqdIoQjT3Z9qToU0R8ZLyOKhubKK2C/pPflC
XesBgCfz8zT+hu7bu1rXNQo3DEEsnuaO8MjgJ+zKp6zZLEoFltfA21aQgEVu7nKW
zf7E8lL939CU41xWmPMJGholuhDKXwXya5t+4L30a8SS+l4lsrWUDbovOJz1kkwX
qZ3tWcpaIXHRrZL0fSwVsbUO501uAwOdnXfzSc3MakrdfGFpXu+JxFOgr4S65sRv
3GZ+vY17CbFlZPRz9VA9fy466rqdYw4GFbH6cgZdnXmTIMSoz+sUN3FqKIcWikxq
p2SxFNI+JiOScBKJlVvT/9sQ2H8slhnRVV/0AT20y8QbCs5I5fHb6IcFjDRjftdO
vkt2o5FL1NklCtlOjAvWtYp7A36PhUVHN9IDVkTfZZj2Byiv6KSnsOVaEm7fx4Je
CnVByKTQTTDq2B5lKkPY8UtqiLh7Lfa6hCza8D4PWUKACXrJiRTpfJvbnIi2N2/5
w3NWwpQEXFmZFzDXEBPwfGHJoOwyjDKcdRjeefAcptRwQahPtvMVGlUGiY2ikQ/v
k8RPhxwtHeNpTcNn7zIM5VIKuRIrUAAd5xrFnNFVzf+NaZQ4J8WaTwUm8kt9SskH
M7qKIMprSBoqBXWhY44kcbwK0HpNAZTNkbJWbLGT3fvX2lIs6m4Dsh+IzMJlp23f
dSQAfO8EkDOzpFW3/v7Tsr0Jjg/PMvK383ijcpbZwhvguqIeUXtVCSUb4gsTp7ly
wK2wsc7RdpicKRCPSKkcWM3GHu2RheRbRgLRjsYsN+khS3jpu/W/DsfIgXSS1Zqh
gWE7d4QVYZIJlJwBzrr+7G7ieJC50RJCbsA18VyUWEU0bNNLdVkJn/yZ/nOB5oXM
70mPIj9H5OQp0i+Z2ayVbgJVznRNvirwARqAu27hkYAvnhvMeq23CYOo7R+RQQ9Q
s225PbmdJXlk1UVA4TV1Yv4p2NRx9UN4MQBbE+gIEcndWnZO2h3F/YD/dLMFS6yq
`protect END_PROTECTED
