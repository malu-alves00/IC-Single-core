`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cfeCKzYkLySy6nI238iNEH5+5UOM9uicY7GCqIwShdy87UnEjpN2eiEqqwju8DDv
tzWxWYkkNlGrJKdGVwWENMRNBWBLzktePMwqJUAoIEdzIQdy+YhmWTarD+Jm/nNc
uvKrIdkmIcvTdJLHeQipHKKdcvY0hK/WBNavtOusjy6CGY/vSHgox5fi0ftk2buI
ggVKBlkGeEhPkQGO7SOths4hDnWAkRSmCmlSE6CTMETZ+JzcogWNobHGMxcH7Kvl
ooPmqRoGhvuY/7bexkHrPx8v5fEaxgXOe4X/jY+soTO/NxUBtODLsvyfwkLjUu03
cZylcUndMnmHhg1Z5h5jsqfnzwWq6rX3B8hi4oPbl6Y6bsxOAPPGEBmFBZ7gYXLL
OQvbC5LN5VUrsrhKC3leazQDGt4ObPIPxgVeUefTSaxSIMFkihZnCcjbrXwWHrnZ
4rpEieZrzduOuOxmFnQ/fn0r2V1LhpbH08tTzlsxG1o2BM3cctFoJ+wytmf7wiMN
8BpyLobOQGixQBQfUSH//K8h7csvle0lJG0nuD2+GVY+rGU/PCk82Rf4aRoDvtlA
Nup/zGR4scccZNrKQr3GURC84WTyGXZsJ+OA2fDQA9fEKd6kf9/6+9Q3weppcuFF
wKNM1y8HovdX7D1Fj1D1FnnLnww+o04JybWWBsG5MFnHoqkhTUhWycuwtY/DfWIw
IlmN6A2wsNwn0CGI14/D6OMTb/U3TNezQOPQmKPegzHpJiuROL+y1pee/kl4ojkx
BKGzog/r2lvXKNi4dvGo7DHkxNG3GL8KO2zLrorVjGOs+jC5rJ6cHOD35wjGPsTK
GXDsQZD0PuRGQqFGB9zY1t7VIC+nSahptMaSIw2Q9Ny1HQ0HZ6Ey64wCdrxzyTTj
+cVCQotQ2VkKkOudW5ZmgyJ4a1rB2tThoIDqRrndF5weJe/ynOy2+3fkve24h88C
STfFZUbTRlDYTDjmNvUBdMP42RNo3pUzbUoFrpiMnDBrA1e8SqZ6EVH5GOKFph8A
mSCq0PdGwTJTVPF2+miTjijvuCSAs6b/ZzkG9nZ/0tk7EbzneRrOrQUdmCU85HqJ
UiNtKWSiHEV8vFjhvLLZRzFPK+wUaDTOclRmKlOM5WQiEdc9C3hsp2lL1xeSRyCa
jvYq28NHJZYfq1YCPjb3zGSWMlYRek44QCdb/kDDAEwjCnopG3cteQx5njgLGnJU
7+fUPEJYalBAzZvJ41Jtf0E3jVsiuKhHKTw0oIs3mXC5VH07eTB1wR9wIWGYQXE+
NEt+1xIYdH19NWyrn5XudxnC/0yQoRSQB7i29d6pjjbTXhZYrbZHqMtnHkUwUGMq
WnwbeCGmA9OoFnhrDgjgj0hMT1CcrtiqR5oDsX6fdNi4F6KqmIn87cUnoxq/JDw+
5FmKfbryy9vwbVFLEayybb85BXclKXB0aipSAUqzyoXO162SUliiNxAwMuPD0N56
FqGuU87MLUwjvmm9abLKzxF81FakrNAuKu1MhdicdGNqm9Dc/hQ0KGRhEk/poGH/
nXus8NGGsnWwJBJ04Q6cmC7Fc7yk69VZTLgC1qYZGIqp+TID5a+GwIEVltdN3JUt
rIbICJvZtvLp9TgJiu1BDdADMiWywireIbBG6GeJcrMoF7hqSy2KJP36yI9gTZOf
rqRZKhbaTFHdXNcC7BeDWYvf5/Unw6eMcf1DUwsRm3bfOT1msdgxg9zpQy648Sad
K4rW2JsHRj6NXQZfMCKyyoXFItLdybIisuy1UlehZBfTUugJLi8Qi879LiqRpKcZ
RXZOywoTAJlngpRTAjBtAOUrWGvK1BvS/t+VqtQdzwJrysxq2xo1drYYUM/r1207
oiln+SXzIndX8LnlH6h7DjmzmHX24TgBAiH4Ls8/StVL+3qnrIIsuZWgANVMT921
/+fUw4gIrcN4XAIhROStxkSDZWoo5PTcmNUdeUwzzJCZ98GJLnF8TLZbMv4OzKsW
O5AanmXYIBqeOq+Ko7v54/UykNn1dpqOVGwD1/WD/2cFBKLUnwD8C5U+zUS0VesS
U15ZWpbvdgOuyIGP2TVBSlum3oMH3xPkGe8gb7p+ZNFenjCLkHR+8dkLdhnACHDl
CxS9uWX9gJaazaPV1/Ni94LOBWZs8P78Jg9YeFkyczr5N0F7dZEVkqjrGw+/AULR
GYljESqaFEjwpijqVl+YlIAUbJtEGt1zYeWjxaVag/QRe61fB+cCPlCM6TlnPtzv
zJZhCxwMnL/eUNSkr2ZnO2LN868uNirH/mQaHSA9zJGzVvxvbfF6GwmtvqvOm7/Q
3IJfTH22RKxXawXacsdxbTTVRwkOxyfjhE7f/+0xt3fhx6zns/7hZC8dq0QC7L7c
6VEYZiYE36n6lkkZ3jcz5AvISd70ESxLpO8kLjIBRrJIxZJDBFS2GQztgd3aGg5s
bvVVkb1QnkGROHT/R7xmQQAEgklwowCnUkL0QFRY6rPTC44WgKEQuCw6RA/kVl4+
VmXXHvx4GLuvkHM8u+v/P4SgkU0oMAA/oee9s2DvEzANXqh4/ctdVdTUsciWsFVl
og7LdvE3d7aqozCOP9cX6i10+gAfSkjhZkelXlDFdleIM3o/tcE2mXy7nPcxk7tu
zSj4+Kq7srI9LO4lNpphVBBo3ACMn2czg9/zBr1l9bRqbYJJ5xU/FMDPJxRhp/D9
94/2MEuo8kG3vZ9AX+7bzfY6g1a87fCmgBsKoKNWayIU1VNZq2xoi48jaM71TRGy
VHGKpee6btgf6OQGvTa921kPp+AXUBG1f0LUtQGYMH0OLTp9skT4Kz7W89yQQ7aP
wfDQ+5HdE5wIgui4F7ck3gOGOTMYPsxPqGCVRRfQei8TspCFrGW3SezDU/5zSB81
VodjE/AQK4Y/YyDI0+xfES31wa3Yj8jJS1YR/vrY/WZJOmJz5qu//qypU9YZ0sbd
gw3QED2hEFoOvROUC5tFiqRk1rxtjc0wtUad/o0PbqJ3nW2IJA9RrTFZuPVYX9WR
nAmIJGq34Xwe+eiVK3fyh/lLeKGrnHW4U46rw0o1wJCLNxMtcwZ3LDrnxTznUu06
BZDyxer01YkvLwf0vR78zszDpDVcjF4vdwlkEO4URxyds6+lhQVUniSKqmCvF8ZT
fXJmIoDsnHft9CMvDlmMRRJ3U8qzyPw6rVspFzdb+zjDWzo2ODR3X79nKjbUL/Et
1ratSdrd8SP7Jhben7AwWrG2TcMHhuGfiuQd9AxiK79mFjkMUGVylu5win65hpiS
HQbhwk1kpc5T4DdyChqkdcDLSbkZM8LviiMQc3oMnN5v+48yhrs8ry5xB5GT+Bum
JwdFXeHiTj83lzOFL4E3sf2poxVxENkR+DJ5xOWC+X8ay8pbKPYVxOMvMZnuOzAb
HK1YikfAuS+Qn6kXnYltoTaMckyBspl96Zr5d8yzFuzdcIZUjmBn4wBmvBnn2ys+
expM84Sbcu+Q7uzZSCIsmeZsVAZhrZO6iJHR6lLrhdCaLEOzMb1d1inCXdjL9uW4
4/493tipVXuX6+gK6aEct2375XE84f5HsQbPx0b2Zt+apOJqGDBGXf6qegFYuZti
QuxpmfJb3kjWRSxM89CoMuc2IeRq/j140uFjmBs099818FFyoysfjHsS+a6TBnz0
89HtHpskIfwzkNTtTuHLAG8nq3Mk1V/SCTMnD0tFxqJarfxKH17Iv/cdTxjFvz7d
3LmgPu1rwhgPsH+jXMniwfypVwKMnFg2WcewvEelP17S4+E/QRsRUdDgbsbnFxfP
98ccdYHkHndHuPEdiMBUd2xXMLIMEAAtyjAWn22OqjoOF5aF/68M2nPRgNeWUKk1
SH1lPj9YF5UsGSPKjN2P8vJbx3dK+xUOCRbHDjb8DlxF/GfNuaKnsvGFvCnCLkgY
iZXuTjZ+EP/ZYCCQlzBWEC4rUDFbusL/RAEGtarwXAqViBiFsNu0Z4EBrkIZIzNL
0k6G7jTuR3PAkn+V9U5rzEmdoL+rcoAGJuXsFGeuu+AeRLEbNLHYoLf/XaMrs2hY
uLytiGw3afhccpKSGrbvssvamY/X3T3mANpM86gwU2kkjR8YwiV6rgqsAHRaxpiu
6jS7soL8Phf+tNsri9sZK1mZFd5zBQgHLWfQYiPW0Fey1DiPhfZvinO3k+Adavf1
ktmEVAc/zBTokaS9HWJqfYDH/i3UT6SdMtuxh/UbXElkT9vW7ggUTW1/rjzE4nvB
NjxTryLyrbX2gj6IZosPCQmho/OnB1lqRRGIRqAelx/6HDRGsmie1mA85FMVyV+k
Ybx6DKNsDImvHaUQLkpOL943BkreqzVwea1W5P5iYGci4TAnbwBSnYTP8aYUZsdj
eQ/anlV1gcRG/TOkauOdXbMWLDwFd20miX+/bSjN+xJeef2FGX7BoAXzYtJQzVQe
znI2ipnLxFfoGXDKDB0mGqwuhpqdRnRsH625WCnLpGv2u1ejA4HKCiALxiq27nay
vLbLRONe9rdM8mDYmLkEF7utDgb4eao+EVvRXBQG6KPQgqrLMMjan8t3ozHAQKEN
gn3GcVJ5Q0c/YUIysOQsxVQXt/3h1phFZwdR6CZKufi8a6tJaZ0Mpo4RHXcQCG3k
+qqTNvwQVwEIhHn67mgij8lGa0tjVKOgnNdiGKmF8a0HoXODZRzr9owYEXNcMlSN
qvXpu37Ztb5jicDa/L5iBKRFdoH3ZXixuM8ts8Cjd2NWjmrmYXgO6rnZsEBf7LaX
41iJlZOt3jzFntP+oPWDRKxDQnrAzlPaZj7eUoQ9jQGIPXpfsefqkgYjn++tqToZ
l3EUh0E7VaXu8TchDKCbj42SCyzS2vWnyR/oqCjmxIUYdbOhU/oPMNwoBSR+Y1Vo
ZAKjazeWhRztukBxceH89QfyUrHmxexCu4Dj10o6KAXCBtY/a+YEu0adO520X5SL
rRJzZLmuT38emB9wda6eYn3vt8zj5w2iDetwLFLCMEaKLBoNp/5WBWY5LfD64x8J
Y4agqHAmTC+z5oPq2G0qkvM80QfFQEH7fgdWSqQWD4aGvAfJ+8xIu8Ox2UnvhMlM
JqAfeSiYV7M6e/Y7pn5HkpWM2y/hP9sBlN85NYPtCTf0SehhUVxBH96nbjie0DRs
rVlGxhcPg7XLLIbp8JgrrXmjxFOjyeN9AtM8OHfut7rXkCyLekIx6E21sytVaSo8
gxbo5BTuyt9mjtLp1KjeHKOmgNhW+qzeBy3cPHuBMl/fMs8HLgsMy4jQIrQO9QZE
eIIAKhFZul1inq0YSjjqlDqaKtlJZwIXuuCAeFaw7sNo239ODIlpmN+aDotHGE6f
uWcyu6+QuSRMl9sefKi1cfpEV1rqFgvs04cvBiWAsD8ilUUfu2a9pC93rcm15q67
1pr383zm81V8SF/UguRNc2AmbjVRPANXmsmwemmwIqXNhI8sqe1CRdGteRc2TGN/
ucZCfVVPpGNbJVk3a8ZHQX/95OqHqIoZ3vkYdxyd5A3bviDSUGrizsNkJ4ypQ7kT
RclUP/mqHUZY0wh/yi83BtuWrgQwxr4hAxOk8Q8NvF0NjMiBwMsXsEDHZa8pn6P+
jgoHaFVhUBkbD9yNbp6c1KIPmhmLqK07DM9tQklJF4airr7FE1LTieftgiqOgJgL
gn4M58AWoepYEtUW/gltWd0HKshYJRCIjl6ISJyAv0fP6zLotfuK/idYc5BG4bIL
c29URNjtjv3sPW3fpKiw446W0GzbHrRjaZeKh0hlacZVBK7ADnwR0+k0rr0c9fW3
WJPsxjqR5CH0vEM4U/E36zuTmHyEzmM5HWHcPS2H0uEoRYIlqstEf95wz2QAl6VN
RkI1wXEK8UYsNv5uZwL0haz7YTRggx2ZE0vfQ0/JCY8dPbmho3WXrFCwEhisi9Vj
PVldT+FTfjiXqK9BH42wE/tXk3qusLrva7UXymv6gQCFXbE3kn76UyhbcGXen60s
FoT6on01LpZm2JPNsR3PofpwfKLARJDz41kEM6xtBdphUxBo7P4QZ4wckkYjA6dM
YxYh3hnFs6capY9kkb1WM/78G6dhaFwLjFsHkVWRY3GxoSmRVQsCT96lRoIXm6ZK
gERN6wn7hYhXWNTqpixbHORyJCizwjFrqudmzQyRg3v+vmzvD+SWPKEckvssbv6X
k7Ytu8d7SPAP6Qa5PkgFVo75w5wDUB6sG2ibIlJtnRka0+WksRyxzf7vx3r9L8Fz
F7d3W/b+Wp6ac8/wkYAlPW8SO/pN25GG+gXx9aOmy7HDLVDt5Wyu551DyZKa8Rqq
7JEoamUWZ/gJhJoC542BVbXnSW8Z/PTEYPEaKIYt10IzKWkDW69Dr6Qx8bdgeelo
`protect END_PROTECTED
