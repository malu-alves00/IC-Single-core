`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
B0OHvnmDgUgMegHaf8jCslBJ6Fsw6tV7pbv+LJIVb5ZhNolm/pmdmQRQjkmmIrUW
4qTB9LnH7+qSMW2mBvhk3dd/ht9gdsiHTeWTH81UqHC4qFcFdo42qqrW1f7HtdL6
WOssBGQuayEbils2rLUknnTr4F/KGGxbKCCwErHF+zHiQJMYMKlbeXzJExik6aJo
/zSrYMyH6W7f9Ozyd43syLQXVVSiZSkG71ULbxSr7O+96UyhcyJ1rFqJUiyNSn8Q
yLFZsQSRqyzwrAswi8CWSArUyXd01BOVeP4dBOTgmQT/TwNwEgvWOm95gUQC28ns
OhKknnmrTGJc6DtgTRjQP9jVExia27vhOppSRLHhJnEEsNlX3kmLEFjgeLOKMUji
k4GgdE77aRYa2uConc5aYCGP8WhPKY06+jtUAR2raWbFNZ1F+DVZ1FIeYgdPlqhj
CsgPIQ9Ai+JDEvz+jLfdMplgweXU3lExc1+VYBA1Fwsafj6Nrn4KvDWHvy03iXpZ
ZIJPBP2ODHw1hiFuXDAkjntVo6DQLz29FE4H9vhPNbrDcyb9L8qlNkkU72U3WgsP
z3kUm/KG8oeaY3xXa8AUQdAtqzmHa+pgNgX33fVAOr7s7WYk/nlb9j1SzSWsKkB/
4R8sQMJzwdEOfnsKZMQW/z74Z23zmGz+iNiryzcHcU3E78uZYPno05mzdKN1dHw+
0IQZmBrmrlzXyJJEpLE/UGxAJjxA+q3tJ3sVJdwWgPtTIrhBARx56s62eAAPVzf2
ALPA16bE71O0kQzsynGWUDHwuCecVFu0zWiozsqeGAk4lB+/kxwjNoiG8NDOTOSd
75SpC45wsKGprXfQsE3AZwH+pDlEWfk4syVtVbVb6yxolYLifQZeMQRnBXlxsZ3Z
8n9dxwwns6Caf3vQgGBaX2JjOm1fiwDpoR+4bbtchj8aHH3bg74x7SDTNemApf5H
HI3oNWnn0Ep6fb2mn2j1Yz+rCw14/wbvX0yfgOllhX+xkXBdIeiOxaZoY0Jc3/8w
DwlZz010cyZWQxDZPzKvrpTiEL+KoyDYv+pUnnx71zmp46okcrWIO7cwfKhx8g8/
d4SuOggNfTsiNBlbGIaabyaHaIUtCLt/7bcqAwsjGDRpsyXsTS2vawzFK2UvqujH
VcoQc6a0NfLBSk8uAh5ow5bmineAnob8QS7RYQ+OiM1m5/jh/Ls1BswEq0mPg1RU
w30Fa7EA9AFPC4DiWJo9KOUNFSitRkA9PWqMPSr3xm22cSx0ADAYGaMNL6E3EZzs
5VpHB7lowrpfArr3gBHbMimtEu4q8psIX+Q9rA+s54HvjINjSev6GTk6hVZYJAm9
FiFV6fVUbpye/EhzKiSiFKUPt6mdujy6SuTGzcmODdCe9+46fEbn1l/W4BL44kyi
vRhBTboTVtfnQeEOLOaRSq39nNeWe17/xo2ka/TKf0DommpdjpSMpr0LmY/sQAeO
EWxBlBHZBg7FJdvltiA6d6w2GhCAFomki1sc3Pk+GzMYVmZula+pG1p6sCsscN4S
CnBKdWhBeu/S2KtukUHPR+KrcdT3FKG543Vwgu67ANzIHs3ljkMWtoAruzFbmS5V
vojbEinWiN5uzkpfzLVlv5GHVASyvCXhrUiL2FOL8XR/h++sFmWq4fTVOItDAFot
YBR34ZOrMOo/Aied73ftSjBqsZ+2Y7sZO6Ko1ANGUdSBCVJJMJ2fKtqDjm2zRS1u
pJx9quzSFOBX5iUteAk33MTp31qp3i5wVkbUeBHvpy74Cxr3CGkALc/FYnAwWhtc
/mhSc1Pc8k+ev8yKs52kI7LZv8aZLyGwZdXRvS9fAGWp5cb4aYTfg2F8p3gDtSU5
KAFmvtp1S73hku9IXhteejIq0r1C14go3IeP1TqLRlD74AamI6f0IzAZzjhDE8Za
bBk6JfKN763R7M4K6yfFR5R/4WfbbGdWJ9+GIjkGXDwjP/aUxXXJEQjKUVt1ZKEV
4AgnLSOT5Okt/umeiVrhv0rSIBPkXsHJobxYNzm1IfqZsN2mkJF570izQFG6I7VA
3FWhXKoNQTciJXnYnoPQBpffyubFZdOLsFWNSWOjBdVY1cLbTPuIvyX3ivbFn6Nk
1iSHjne7BMcmP+0xkWpkuuDvw1dLAhpa4WyOzG+M8rjtik2ZyFbf17OuKOM2tJt6
dMIVazAxkNQPgjpdzjg0PRYndksNTqfHX3GZaCwmYqs4yDaHW+JeCxl+aUR+CSRy
DOAMRZCrYV258r+yqQAAZ/aEaYrJ2SQevovs0WrHgl+J7hLnOr8lFj8o1QE0TAg9
mnHirzvgS7QD1o4uC026mWlXwLMPp+yBUeqj2ir6Va6lc5W2uNbuEG5l82Co+FXg
cSRVdyFP8Jd33UgW9JMxsb9CPogP7li3/WMCVLzEwuMG8IKZbcS6S/v3BBjss1vW
mHNnmUms6+vKmuRzf5X1Ypo+DvDEhIdZNU57tt1gdlhbzymV2ZLLJ2bcxYuJjQfG
loBBl9P8q2wSDAR1Av+7tix2OX5GKR/VZwSsRiIJc1oe9UDuirXI+fb3ZUJXH+LN
ZMWNtCsAZ9+yGtNDfZQTwBs1UvXxL7pK5n5LQziDQkw1O0jls7I99Xh3c86dZnko
t04KUBJWdmaZe4B01RhAClnURj0ysb9XMjibH7E3QD/Qnn8otGjmA1vIAVC0Cjwl
upilW6zvzxXaXtIVPC9u7/3SRe+IFfponNYYxUM4XiXvBJXWuwIk6xH5Oys3Rw9v
YSFwBQ70Hv1h4LHgnAnc0CeFOrNn7vUF4bmZJOdns/VdT22/gf0X4j5gBkuvzlRA
7E5/PhQQM+mWqOEbLXUpGIU5wkvFXQccSWKIOrUg0bh83fINTspCTB8h5DNICZY5
Ffbko/4Sz0VZuIf0F8s8LPtmpq/LYxlFFAK6a5ai4mFreELhS9dzuFzUmf3MBtyi
LEG5kC1ilFkEIhm7JGHSIH9YOX18dWVKte6USN+ZBv+RK3FHE4SNhWV3dShY+6TV
4oFroN4W/XaIQnJa+VslX+QSXknffPLMNy59ah00LcCa5id5ZGFAUj6E7u+Y5AVT
p8w4tu6ZcuD9f7S2MgIDSM0wTGv3UARkSdzFoAXoPoJ5JsjkWI11lCpweO6qvsjQ
rGTd54usjVjf7JXqbtcS7Sf7w38FQa/ML48b6scP/uOQbqi7sDkuhr5gU/s/El8E
IqB0+UdW0T6i5ON0Z+0Qx/bhHKzEW/WzyJMOE/ChNUD1x4akTi464ZR60S2abG6z
Jc+T+dHQa4PeGQ5kOAw22gWBjAUNuAAsqCJ9opdmUm/iYuA8zV76i1xAsoZVwt2E
01IoXh26MwmmIVut1secZ2bgs6dbdHOQcL5k0yuEtlBjuvskQsiV8vxQKJ/IRHap
dauqaWsNlrH6s+EyTawMScb5BCfqqayUlX5/8EHjLQtpwUlsFrxX8kiateXEbJHy
rP6WGFtjKVtPfvxYoXYO9Q==
`protect END_PROTECTED
