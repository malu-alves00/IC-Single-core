`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rATw7JxTtd8QeU5XqqR96xJ8IS1OuaLYpZbkrhaCWJbHgVRUq9bFwXatwONBDf9M
aITeQIncoh2misWxV394uCUa/VROe3hoQrIuueju+HOM50nmKFYX6vCj3CongSFb
ONgWz4gnyud1gl7TePyp3FRPxovKRKYVen7NWp3eIdpfVSmaT6qXmWUDGAXVjh4w
2P/rLdk2b5KmrwNVzC9yXwozaV1YeaUmsZy9KViwZdcOXqFcMSd2LxvhcT18OQPr
+3XmMfLRv8qJwjvsnyCyeBu8WpL3zd/0cnWDDIFTxhW0TePUv8taboyzRrzueRe8
nVQYIBTpT0wIPL6jXY5GmAICyi2SZLVqSwCkrTlvSmIrqLqDulaJU8PrUj9WWpom
rSYUmh3j92k65BbXtaiZsKVtTsj9fpyyh209AvOM/JuuDzzvhbBaPwpuvnZD6qY/
SAG7RueEHINOc2HMaUff9g8gH827ZWg2jh9Ur9h/gqtSeaFVd2oMBwLQMnjpn+YT
upzyq+8nF35JxCs83PQT9U00P7Mml+ep4MZ7ReJEQTBBfR/sEGPdWW/PPwqA1kLs
UDz+fp8qxTL997/f23I/jONrvviqci0wu3JYdMngnCA5cCGx8sRktuY3uLgvPe3M
dN2scDsqZcrpFGb8ONQU4jk1VkSb8DZ++oveKIEkBVYZ9lsbVHnhPchQ9YG6q6ko
m9lVfG3aUZQwmVaYch8ngXSJxI8QmJKOpC5i8UtBis7ildM1yDCaE50KZrDMiF9l
oxSyzV9IJfDZSjDLoOHrQLC42hSCubYvH6JSGJlCs6yJtgfzZmD23np87VP8g9a2
r2Q78E2HdU8tw7ZCivzcuOh/wLPr+wICbO9rhmkOFRh/SB1krW0EsmTYIUFzbRYx
k+aEWpIazk2uhWGu9ABTbq+Z8Z4CX+WdDqPUqXa1HajPL46aU6bB53oCbu4ZmBJ9
WWEJk3071ue2ABwHbP5YomxI0lzFX3EJ/wpaX6eBZs+tFBAP7x7wQybAPDFJgL0Q
LvUeD4jX/E32C32wfKIqY46JLkW+aw120Lih5QCrbSao412Dyxf/+ywbce0bH6v2
tIzV53DNiuUvHEro85+dv5r0KTzIuUYKcPcGEusade1sYMlbXoriZeo3Kq5Zvbxd
ZM3qP7CW/SY4GdYYql389XfMPovO+352xrl1tu1ItqrYon+GZ6OsjR0cewjaFjkl
qlx/OwaUlvqHgRXHQTRwXHPaKQHwZ8uxtl0aWcN0eZgS7R+Z6VW1BG9N4sJY0FQ1
aLE7SEe3NNJfU7/uQOMjxVKDJrfJqIk20kXL6JZqIAqilhGejiuW1+JZ+u2CsHb4
eXkOJXN+Zc35QWmJ39bKYVCpjGtTjNe0seCbmUVaU+dL/+zv3bmBQyT/f7HeMBMv
2LjBXLfjPbnjrhaxG9z/4w3kL2gZYewRGtD1tLfPYNYC6wVeAVcOBbXOCAjkEWqJ
KRy5ubb5+AyeKzCjeAfP3QSoUlCTNqjk7u53uqYT7rjrO+nLbdlx2+luGw/Mf4+H
HDq8s7f/SsdbZPhSemNmI4Va5Ftx9oP7LTI28jwwYRcizD/lHbRkeWndyys/GpiK
JfQJpHl/T09mVD0cVBTr6VF7PuPKWYvi6V9DjRQmZ5BlM89FInAiouQB3Zgib24t
bM6wQJat312Go8WnXd7bQOWws1hOiHxGnD9Ts5i1KWLdTC+nGgP/bGPrB1fTcX4n
I/8p/SoZlzGXEEnwB+ZeCh8cdUrT5/VsNTjgGV4PtPohyCVNtEvA83j4/K244ymG
ioWJa7N2WX8IbzBsvReufwDkHbM+obVdsoD/31S9hNvMCtF8J2rK3+Hr1EdpYhJg
5yAusoHjOdqbfnqFeG7TueJLxwVXTY+pzgRRe9GBQFZRz68WbLsAixMzLjqP8570
JKAmzcXJpbnHPLabLj6n5LPQ7uO67cQUpDE9JkBB3vg/cWtt68OOV/fR62pPmjoD
hA67ScCCgpeeYFrz0itq1GIc9tZWMqwdfikZ+/ehYda8IH5FnCEu7IKJ/nKVH45s
zK9zRWvoS7hwo2S1dASZQHyX8rZOc9rWA1TZesRXoszJI2aXbnhpCE06drFPiuc7
n6uPvhseOXkDwROsa81AMzBl+FIa5+uBepmn/0SxH6yMuZ01GauR7Lio+lOHGfvl
nzhfhuJ91FDEj7csMBEnhzlrMvNMqoKrWJyymbO6ghbRhRB84m/M4rkJKOQcaPmq
rbPSHfRHLOPOtLur2nl/1zGH5SjBiin5ja4b8kgRa38rDuVUqVWp4Hb40NILkPER
yMtJv+fmZzmMz+j5WSJVWfl7TYtOq2W+0+9sJXZ3U1EuaResyXX4+dZJKMrBh+3H
s4Nkv/lsVnbX6V8Hc3SoIWmOlvkCcvQwnRI8HYZtYmlkHgynGztBtbVOxntgWWTc
PaR9SfK1p5Zez18SnwQ4ustIWxEx7nmHiQKoMRekw3gCkP5BQZjFRiwrp1t0bBmP
3pfmy5pjVKhN+0zOtmBQ/8MQjSbZclj5VmVJlM4uxQdVgHzoDVEVZxRFOpzYAnQ7
PyHFF6RwAwI1gytPjAz9sm38LUPNU8RlUeMePDI3OXEKtvNeQLNxfyh4TkNEe8J8
pFg2GauvDNevf5zu5wt9LPh1NA3knt83A6s+AM154byMIeXgs3xpkRpK0uEjS2t2
R+YBWnQYejXcpEEW9F+SY+pzU0DvHyhce/aljR5Om15Uop9wpu3QA227nQ/h7et2
iDQ3yr+ydMTnKNsB2/aTWMBXE5GJzKXe8YjicX+Ag7h0PkBH786bGofArr7ZuJCp
zURrffwTnYXyfCaDNQWszmzjGpjncgZrc0ndcbXZ+ZDkeT435U5KtcK3uWF9ehyF
0dcuIKbF/lEeOhtgE/cfTpYdOrhwBTEO3HCIuW7FrXKUpb0QLD0TSOoLvgMIT5a7
fGNaupFPgizDmRZVEBzzfqPzXemb5w41nBXObZOE1RJxFzKQDM8JNcna42Q/VTf5
2xmP3qLYTrx7+dNdMUmVDirtsJF2VhENcRm7GNeZea+CwstO76hHPY+/ZbquqgxI
5H9RE2FgPPnJZ4j07Eirm1S0fmhYGBB3IsD22MW5uLe9ZIG0G2N6pKYSDBZLkNE6
G4UqeD1pKaioxy7EZeoB+0BSwdZzwh2zshRTZWfq3ILBbicqsG8frc7SIGRuN5mb
LuMf7o6hsi3k5gkHiem4aLd3pfWjlD8PCZRQ5suL6XOb2sPaD9MRiXdx/ZBhxKeb
4igS3V2rgvPcRbRGeF/XRwfO4rW23dy9tmqvNw2TSwDJ1wkFFb4XXPSvZZNzex2X
MIUx7qRS8R0dxrSLCCl+S5Dli1V4sSQlCeXx6wz0X3msuugY44+C0I/3yfmsigXM
6K6Url4bM1CkJuTcWgjhnhrYtEamd+tzFgX1M+Yjp127LhHWUkRGK5OFDiSX7cgw
7k6NrUOdMHAH8lTsOsRln63hRUZdN1GoaN1ZDVGKdarAl23cGJhQFr4p7zz0WEAC
kaNUAeLs9Rl2UXdr9d8XqlMMlmhxepDTZH0yDDbTIZ27eLnxfkqZJQGT7/7xL9n9
ZcKFg/80Vmq+6Tz77Owgsxs/JMDBEAFebDBAqDz0yYoTISSzQ1P2M/o+LNEHA/i2
ZwDLQhabwR+phkX/w3tBCuDCIqrzVlOMq/0lRkaB58lvkmlHS53RUv7JPX8XyXsN
slSDyMU4Lek2faXF7i4UkDGWcWJ54b8ytXdr+zQQDVpuiNtWDr+yZkrV/APbhK1L
r0Rf7O//bNb9TMnRJaz3tfWHL7EhmcSeJtfeghnJriVzOj0aUPIBBe6zW1hrsxVK
xlZMREN6um2idsp18kOJeEXxpisiWHqz862zsUBxvlc5toOsG11MymBp8F2k/YqK
MhN/B7DcGng/8Zp1k1JGV4WjBbvdh9+/P6GeYTJZTGsNZDjVvkO4+LBQg+C2MwWQ
GSmHRCYNgIdM0lhxvThw8ZUSOYpJqufNKiVmpEEuba3rfBOoZJ1ysoR5exg6OxzK
doYv7e9c31hf5g2BOc7KqwEpm4/2IWdKmg/jgRLX6RxSQWGWEaOvDAjrbjCrKGdZ
HEopeKwDlNjTbzHKvQyttt4yUYUfiLYOSkhGyfaEhLt7j6vf6Z7lYPy2zJRALT8L
qVOcQ80FkzGHF5ZOK+ct512F1B5j2QPWDAOlwRK4E4l185Estt72ptTmmVUgkqvw
pdlV0CXkAA0G+u2Ght3EbZeWvkAnNhSssFI7gU3yQMcbhkvhOkRLtHur5Otpvf13
vXkLmNkssNx0WJFkQK8PyPEU13hHE8PPySryqbR1KkYIJjlaLqhbI0rnpfw18Q2c
zsmkUcjIriihI6KiM9WZ/5Cc/lyO1NlzqTe/xEjwfk1QE2odM2n46qgzbjssmCvW
X0wFWRU9r+Lw0+nMN/0fFAm334xy3ZiA14NBNtn5TRYguWyWqn7mCe8A9lGo908D
5pqRFozzidWZwW4/ee7n25zTMxk7pK2YioSfdlswIPoajjMDAgXmlcOoGCu9eQB/
SDc8StgkfbO9b3DT3ycpY47HOcyCojaZ0HeFrc80ToF84TJ1EGGMwBnCeWzbGtCD
vw0hMRVMSCtEjkseiokLMAYZLthr/vmpt22CSRA7l2q19dWo0w+NzkP4d0/BBG2h
okORcupQEBSmAnDub3Kj1NjJinzP21D03B7bZ9q6GqpnxbwA2dnoKVJ4SI9SBayK
gTyrzD1xxVwVp7potUzYjW2+w9VKutQBN6FL1iT6+bX2n/wqe0iH7WzK4wYObzJ3
L+XyAcj11k1+F8l+8rUb7NxkZ6HKryBLN4v9xzH+UITEgAk9LnMslTpleK9dMlqH
3mW1h+XEFzv6k3GWOiPtfk0SkWjbPRtivICHXViUYAvGAL5uyqRtwQ4SHub+SjMP
cR47rHmV8U8sNKqGrB5t3zpdak2jamK7vw6Q02ozWlvSqmfGFf6PhzVKuCEujzJT
8fMtWBRTr34QBuuHkiI8pjBg+8vjJRXBc+FjNL13wXGIRiP03Q8WLn3pVsV4aaDn
s0cd3P0fHW8a0Q0LVOJgr7pcdrCfRT6Q959VrPh+D8jiwrQsRewunRuWRHAR091C
ZzT1uf0qRep91wu/QhXUGczHnyzKWTtky1aQ0beQUtzdRP4Wl9jkBy5Tb8Vj5tzf
GwXZS3ybT79YD72btzVcevRjEu2ORWSerMeXBW5UB/5fd7fjNHAsZ1d1AKQCKxqW
VK3vfTO2WNTX5OAGxkM9XLaRYfstUJUm4oSe6mXHp9c6klyK43sqS2FwC55Jjo/0
2VrQqnZBeGLHMiBL9cLIGYHdc5RRamf4oeshlI74Y8e91V0ObzM4ka39YIx9odnd
WiFC1O54EeG1OXxYDJagAtOpbg5ke2/sykLWR45nH3taSZrgO9vL7s4X6PMAjdGJ
eAvEA+9moR3iVKN95G53DHbhHpezpvCKZCVgtmShAXZplZ2f9ooYMdeH0eN1Nuie
uJteBtZX474z1NtdZhnL43g8BsvHQHOiqvfL/QWwIXSl+Op44nxToUc8GUBy6zwp
yWJViomkJMteGmWNwqahEZCpmkJ/e84h0EjF4AHYzPdksqzjBZEP01VT2NG5zsZn
OLOqr3BE9cb8dx0yVJd0zoPzdtnD44bkvA6k+puZOYCd1HxnscJdYXzA+CoBwrUl
HOsdk0In4ep41HIq0MSF0r+WIAdoaIixs81hLgGBfz3kCs7LFJ1+we8tyyIc9/qu
sh6Z5gFO+/F4xlZh9+Zr9QHH+k/YIP2FZFjA1DCVNwcEvjIJ8ngZBz1fEjQo/y9/
pwPOK3ZN06W/4OnB6PTrTS2n6vJCtG8xvUxN9L2/sZ34d9hXIv5Pt7tpJ9zRGNP7
GLwEdKJxzemfnVCRd6Q6awSJCgu7aJOMaHix9ar7L4butkHZ8/loAZr+cinoeevI
y+Az+/wDz+bLQ+OTCvyEwUfBxyfBc4HCcII/MCNuP8jzAntF3qzQLvp/w1LgyT/c
sDRKUqOy4E1KZlWNbcXhWfCegJro7PvX6Vshw4JU9RVcTmIs8daOt5sP+qaT1W/s
Mh3bGHLdxnT9zYsznwa8pWlAjO3Dl40OBUNVLyk85PuhuJTOwqCJnVerPc80Hgjn
8d1vtlYbIHX4uqk5rGkEezdMe1Su36XVUV5D/vJpbZPXdsugJIRyfd1GEMh8XHYc
uE4Jgo4WOswfOgUeUOlhElVtUmV/v8+nT5+J0EM7X9OTIG4fCdF3Nd9qq1wy1VlE
BJqQf1+8CylcxhxA0yj8U9MQcNqWOP8NC5axvQLLd3kNjCCdlls4z+PTKvdQKL5r
gGmgYyvZFL2KOuS396i1xA3LUNwvjD+iXjqoZl/9G7KQ6/Baoo8/wj9cp3U/HjIR
IbK4FtZulwhNbe1seskMD62JS9UdbLcv5+o5PYj4Y+4jERGn+1qg60KCugMQJFrz
RLKEBZEhJQ4t3lVVSiCkolZkyODH4CCzGyMSw1tAlEg0ghI1Me5WhrBvn617LIWl
C0i94ZfIWx7NiOOtp96qAvbFG/9MeAUck8IXAo/PYmad8Gk/mJfGHHLdcMrrsAI1
C4SPEy2RyT8zlR0FxJ69DK9/YqUr4++2JMXuUVc6iq4diQH8UMFa6L0zwmRdnfP1
WoGFNUZ/2mFEicfFKe11GMHtIa0i9rBTnodLIGdzx2Jkj4nDOh5ztUIYM8MX/Zq3
ApWlvqbeLs8HCGZ6ak3PH9d6TB9aOxSN8qubtOYN0rTPPrJBR1Bzu+nUJhbsZ9mG
LwLzTtf1HLOuhWrfGkoMWV9ZEQ1d/ksHhAZGuteAzqPeetelP4AJ3qt44Ql19hI8
dPuiYdwm3iLCQRprwNUwqb1CV+lBkCzCmf+dyLQTELiEAEeIf6/BguEL4OBqB7tO
ceS9nVZdhcaznsmNTh+Usp79jbOJGyQoXWOgmBXDdvdz4H8NEKTRJ8mGsqubNWH8
CNYgyy4MpRsjzznmPrFyalcx2+b/Xg89+lpE8bkt9ihIBBY4ZIwpLfXGGZSQWwvt
O2vL8NFlNDtICHuUWP76i/akP8IDvIuq1nxktyUDimXHAHXugvEOCDJ8UXdVB68C
HrFY87423nrdz0wyfzvhNxImjWgvKLRs0QXw96fXCixdMpbMBCjgeDHQXo9Rw6Wj
9fHmNZHCU/yhb2aDGm0HmkW0GBL0d//qRHmLd2juqN0mXhHu9XoQIYjyOUhGOqxO
dR74NrQb2No0xL4auzDNu3p7jKKEn9PvMWl6fVN3CjSC7i+x6cgUnti7+BsR0QRm
bIE+JIoiHNEwH+uJtXIjAWOLdCZXR5bhiBQ18gilC6633VbpQiQIE6KF35b8vXBI
W5wHI3OQjaKciEBornIakeGC1nwArslPQAsDIZYwiHGuYTv9mY50vKnRoO9hb4Ok
HiISpEO1xyfWhystRQ9xhK5EH0IDpaeP9JbM/gO35hcHBIRxj+c8+3Vu+ntO2/1v
KdvSxliyAJDwKsGButud7IzJUOTMe6fMO5ZSU0d0Jo461xexSNafBMu6vjepGqPu
707dv9IwGhu97M8fLW5icTIaVHgnN4HRg2WJmfo6BwnECgW7dndl6Voubvw5iLyI
dh/DoYjFcL4TknbklZqDLMfZQ8iOr+cxnhkudws0Ig8+F/zViYaMq4vfuClSX2ht
uvhsH5lt/M7fFf9ztQ9JXXyY4K304lQRzuS0loDrfky50wpBHg0sKmSfI9132grt
qgAlqk42R/Q7td2g7cBTWAgJvsWlUS6HNyp+YCM4NTYHI2+3e/b3fFTj4dlleYQB
MKKB9TGOdEMqwRLaJ8NS+BYFB62DO+gRie+n6GDbXIAyFfSeIE6ZVgxOPWeGse7s
cblsM9lbLKYeVlYwmWFOGIveQzhUqHISBs4aCjgLSAoiSq4PaHQOF2WHpruskR14
F7Ksaco4hE0v/1cfCJTO5BY3DEYKZTTDUNC7w0UCSmElkdWeAWSARQr+jaHg5BsQ
zDYLfDgRokepLYZzQdAEQzXs9WBTLw8EDoUkuadUxnM4+ZjB2hN0pwiPEI+dm2P5
4Qo7T3FOjj0KIgPBKU7O7uj2vtwhQy6fVSiKZypa11wp8cmHVmEA0MbE9Rox21WI
RQG8cv2/5tXIPqUnQgixyT0/2bgtdN7YUi3bvKFTFcGlcY8cjarHHtUSjlb6GRs/
AvG3JP/Y6HGI1Jl+xO96eht3VkOyQaPsnpZR2ACcYeJgHQPpzROWmz4ZTbziHh1p
SadL2MNv6Gf2yxHxlH+5dCNP+uT0Grt1Nbd49G//nbHB9zRl0sTLr2S/UPPEnqbB
p4b63nGF/r9OB05fkc83HAcjOkYx9QxlXeZ34fLOZLZ/DjpNt7g1x/KErg0MhhpQ
VagBrKRKKuU3H0zENBYU2ekCwPQWNbSFxBJ7LRoexE2pvWinXIJ1ERQzdkCZTsgV
pVchTWrEm92Vpb66/30v8KLvKgGLQXgT9t+iPclprlijdLjzJs5DBLh/Mv4ek+tu
ER25TpEJNSJpjHSo5w3rrVpr9kx5Tg5pyD7rdaGfJxjmAGevNT31Bej2qU6fx/rX
55jSsH6gK/z9wsEFpssPuTfxTj+S1NB2O42Y2+h16nlNbbcc5F0dAOYdrkwpyg+b
TXe/qibM2MmINJOkE+RUro8kk3vKlYQAnOd/p1c8mLLvzW9YEhs1rXZQh4S5gwRx
99SR/1CML5QP4E+UWnudGpPRdYAavY0g+g0UWHRwmHqfToH3OtIiVyTWKTEY6V3R
7txsqqWp+28CO0Rrbwa1whW8MGMlCumB5BBz9e2H6XdhOEtOkWmO71LDcy+Gnwlc
LZbDPlpQE5JPp56qInQqZEhjyr95qlMuithyL8ViWZ86MPr+Ywl0NMgpqlj05wb4
8GYhi6QvBv0c/nhhxAkiU7tgcql++zU+NTiES5qEWl5eM7Ph1xHrjh0MA1U3YNwt
xaHE1kOfjoZnjoaa3uLMBZN4E3MWrGT+r5J9d8P50+x0qrgmN+0c9Sk0ucLqL5e3
zIb/qEBUSZ1f0JrBD/8y9XVddOGvZpmXOhOMwd1vz4XJoiuB30/gCl+I/gm43klI
9T1wV18KL9iF6/t9UxctTXIpTgxciMrY3m6U4SX90mVX86U0nP+nwNzBDFfU+MHO
I1W0fl9/y+uvKjtncEycC2h/TzaA21a+YlzQZiEn2Ph9xwVLsfOqJ+GU2hZTpJhF
Y4bfFQZ2/4kV/zZqqdoQTZLf47YkMFEeRLNfeQzPdHofv0AzT+wbAVZp6EeGsakX
CaS5r07N/I7UZ4bymPXLMhRSc/BLPFg4N8miyaJI8bnuVe/UeQO88whRQcNrW6r0
g23zYl9P4NUZUiSvhSUZfj6AuH3KkIk6ohAMU6vEU7vXCHgRRLw+k10SJXLfpWjX
ClSh2Q01ARRy5gCHSTN85zEy8RE7wXqL4SWlDKLpvV5lZ2F0RxnP8lEK6ChjdApL
opG3KvYJzaBTTwaNdaYSH9H2e50dkCzYav1PWdNZ5OVTdHPOWRmOMt8DMqTRYLVm
ZA8+PQu4yxnsjLU/hGkEUPv7jOrP2HEoS2nCm/r0R9RLF8C9pW9sWKpekiYmydiI
ZsYmkbvg/lpiWqrrKgr5hkKjOvPp6P0AnY9K9Rvkktmr+kg6tvJ2m1RfY+LRp4p7
ZjtSswr3dQmJWVtUUa9L6ubOy6vLMlzAmeZ/oeZ1I8ucU72PgSdL84m63CgeUrB7
xT8e2zszaKWcHUvCf2jkVX71s6cdnzlV3J7GgtOOxu8zn6mubQkUoeuEV5ZILFpR
nWc3DM/Y2wHiuiWbzPDS5WvN0cfbtM9s/0fXwjrJ+GuXXPz8HsxQ+SSJub/Q7kB1
/887Ar660hBmsE22Pa9OaMENdLeu7s/z8t4KO/ME2BMXPSrXk0Ku2bEs42W7Pvee
h9Q6zl9w+fjMs0bZ+2amrERUpLgm7T9tgiRR46qypLX4kU98uIb/xkmQ1jHpG4tx
DkbA0ejR0GJCev9OvVZTD4NxMmE2X2XyA0iln+usqvFXu0tep2TKBBPmei+wQl1b
R6LKK3qRDB4AzQK8xLyofqQEvMkhO+TeQo5e2ZNnYR1zgHe55ogrxFKwUjP3BFaw
zmE9UeNdqAIkQN+c5tJxwJNhamfYAhBUa/k8HrtWQf0P/94OtvGmiCKxASX2wCl/
b5lLxqGMnO6bA2CJaRgSojkgcvj+GxzuuvrXy8aqlD+AdEhdI/7GG03MSZJ71VIZ
8CHbNxTBffv/gbeMkg0/vvJ0a6tw5JHdD1xxceHk27w9OxYWk4Yvf+r7N33CfNgC
cCHo6uPOPZzOdVZVgFE2srb77PA1/JhkB+YnUrze8KVT6/ccOAkMMDtoZ1PKTB5v
mhwPxpOq6TW2txaTUJ3TbwQZH7b9Cy4ShPiIAzR+DBUMCnGEBRC5qqTJk/ZyeWCC
vkHZ/VFoF8Z9FvHMTAihq1+rpNDCyM3U0wjQ9OcHmi9ED3DmUsDlr3OgJ6soPmWI
GxbWiZQg/hXpFqe2JWvq7PoJIL2fvnIIbEYZDJdjwA6t9baR740qyPm8tEs43KJH
JQiXzZd73XDKX1014LSmwuLVeAu+g6CB3SwviMcHIlTwq01tf3EkhJg6tZNhp4pY
b+b1uLrFR3/Lr78fq0A7NH0qF6Z3+jfMewkMGNvtvwezmjdp9m1yoY0bjeqBlSW1
M5etPaEjNmIecspxwVL05Y47JudEi9qRjw524YnkTKVReT8JSoPPYovcCEd9jq22
Cx6ovkWjn1GYGUZOu7sDIQ==
`protect END_PROTECTED
