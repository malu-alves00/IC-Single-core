`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bZlTQnitCqt9QJTOOpOGEeLBrs5H4eFd+oBEI17VVb/AR/fcUPzQRgT9/q/9XHw8
6DI8r2faHpgNjjg/f3E/AlnotLgbC/AfFBA3ZimOP400zeqhFd6HJ8whL1vUSAcA
G0Kj5z5wYA2/k18DDfovNY7KD1Ac8+DuC/uXA/x/TUoNnZsWdX7V74EDxBAM5df8
hvFYTtb77C1z84q3nIAwt+4V9XsBa9X1feYRtg/PuBOrxuyco9M5eD0gMEyuoY0v
0XXZ2Lsa2Tv/ORzm4vVt6mmlsMTfuJPwrJl8/m/hahND1y9jpX8HoY2CwQV4RuNR
9x5RpYQrT5cQwg0tNTM1tdWJGfLLIujnv0ZEgzKK73KGM+IcFD7/oMtLV126xxMU
W2wxYhP54FekIcl8yCclFzckRBqcYbQVFxIQ+qXTBgvgycsrjIdb2cUSRF7Rm7OL
LMfUEuKJuFEj4OXaajJFWx3yrOd1g3q426Gg54KMRRqJHCgyHh18ljhjV7tDHqTv
UvvIrVF0WA5OiIhe2VNyoQC/+gpB+K31O+6KtzJ/ScTrXMmoxiNn8xD27psHV5Ur
Tc3i2nufGzPgyWFz0TGIEEXMTvSupCZL1Yr/AHKAYbl7cWd6ycH5bjK0Js2XgnpE
8qCc9jVHqOIfD0FEbrNQyjeuVvyzVEsZz6jYMpKVLTV6inVE6P2tLNYy0pK8iBx2
zwhz9Ug5LcbJ+MM8SxIq4sota3fZFrKrb+boKv6tryAe+hQ58gTobqqDeQdVJEMZ
Uq6AHN+/s+gDDvZ3NcYgk/JbLtbOEwhUP08ole0jOz5KE2HOxB50y39EQgcA4wvY
gFLsnQKrRsnZvFI7PeEXBQt5Fyw532putjX0jCk9/+R9tNptZlS08ElPcQCOxW8K
GgtYk37Vs+S1DMj1Ki4gCEdCL0klhINoyiBbOj9Y+nydCfAkC7U95DlDH2AQRShX
Gkr9xf4yOrh4yevuItVGRnl4vCHQPlK0fwbHvJuk9+gMILsf+TdzD67uXex0DOJu
WeABKRVmMaHgKNp/waT4QZ8AQTihk3/vNK8u1J+4vJIyhxAOj69OHOB29xFPI6W8
+ObQLfSvvFKc3aI5/RmVZCpNG1HGKFwHn1I5nH+jt74JjE9fSw/41w2y42dhmKoF
CCfPJBQaFZoyn6jyTnkV/Kt5EAMzm0uvIyq5bfgdB0yQUuJacbcXLb8u2ax28Hgm
S46QP92pJ9e1Ubl36ZWTyjjRjBRhpXTk2L6KeuEWkc8xZF9ByL9PwyuOAFyotAlw
JQbEtWZOVfHgXPNvBQl6j8Uv3sMPo0MCTAt+FgTsqpjttJBSCMsG6UzW+g0obeVL
x0N3F9xLOBo1J5eUvS7w1wzmfn+uAWOb+FYv8/t5BvVE6qP7KPVAXXU93RtRxBUN
h1A0nYAa2ljFZ8NqCe8wrCzhKIyJJRs1kltsfbzsKX8YI86OUldbdpZvL5/w8s+L
GNzRA1jtA6HJt5mABNJtDjdbDAOWRmR0pfCFjdusI6fS9/62LySE/CfIG7UxOHhM
0DfrPf5gIP+h3nUjOOMSiXglR2Z5lDH0f5plW2TBdPrt55oREyG2mR7aBA7581gh
iFSPbVHJ4n4XM9v9I3d1J0ZLD/3FIsQFQkShvzTa1nU=
`protect END_PROTECTED
