`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eJcwMKWEgRuXsxiZ4G8RcnZ4dC6xsbpFgzKo+WQIR9Ohe5hP7kJ/qRW/6r3NVYSN
6R7ZpLU0TVB1I8sSc6dfeUUzc5aUorY5ANhmsRsJGCXDyC0C8RZLV2Kg404oYk3X
UQUPR7Z6SFHduG2KwY1wMuq5x21aURWh7uzOKM+NuQn73WaKARxqJAspS2LHK8eg
7BJYQfbYqFvpNLOSk2BMSPsfnEeajukw8Zvg/scF4yMTUeKOML2+o48aIZlA3Ah3
6+99kxI3URGdFlWEAMm0fMqBh6iW0R0DbSkLegaCAxq5lVkYvlilF9WCpbDP9nqa
SOlTZaNgM2MOgCBCnxq9ZPnM7x787MoHuddRPriSc2ZhA3uSJCylubtttYFFiEEJ
7mpPCkWrImk4C5ntlUIWij16JY1ODCii6bSZxKRaSblk5r5p6uceX+03jLgf5kmQ
iH4oruV3h64xr8bvKUh2Cpu3qzUaY6ENxA1TF6V9b/FtJGk09A31JPmkT0K0RRRy
Xpf0efq3mNy8mXIfI4JzWkpvqqi585FBd+dJVIpJKEneMcS5LtIdVilS4dBQr4GW
Shz2Rgqwxh7H4gxdBJomlC4Qfv1bSWjjOoqRTaV6TDiYyDr3f1YJ8NzFQIwcPaPj
3+LhQ3TT8QGgLHqhZVMzwAGbumhcmB/pXGxToKtwgAAJNgMj92381aAIW6B6a+Yw
paMoWHICDzidIi144bMgqglV+iSwj467S3NPWZSn+nngC/GmPXfwrBuJVM2C6B62
7UnevH0oZxDVgKXD9sUXro3Z4w405qXlWXaPn2ObcSyVIMFMnUJr5AknipEnntO1
jxNPC6GgEA8txjXHIt6dvqvQ/iaIrYGlLwZ4tlktVMc5a4Qcps+Js9dIQSKKGOpy
q5cjh+PwpfC1Y7kvxXDK/y+ofcsfBzZTUVlSzysWfok3/6+P0X1lXE1vUz5lezJR
vtoc2udn+nhIf3NBLbPlwtoqgw0HkHe+31+qd4ID32QSRGUpZ/PvVLsEMFAWDrEX
AVz0Oc8A/tyNOxyJdn2eZxveey8+FFQUzPcsqvqJz3/xYoaTGp4RrQF4qbTib2MR
9uDdg4T6cF5zRFTF6ktqaoO1xDFngzRB9v4ccbGZ8r3eOWClUhByt6Vc40lS5MIS
`protect END_PROTECTED
