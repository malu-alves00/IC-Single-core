`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ppg07ZvZToEDC7PQ6/6q7wUP3uiOAax1ugCN6aOvcJjHDiv/yvlWx+3th+WslkdO
QwJDHmBqfUW4b463vqQDi2MBa/Hwh4nFrFt/N1lgB7fuCHpRjNflNL1MEJZ2UhEA
ztDeejHrxEBkCq6LxI69YFdFwdn5AOZxh3DHN2gsaquIhEpf+mJzd5ddzLRsiTtC
2eDKLhrOC7oDw1GzkcugfAJNkUkzMN5opR4yuMUnweU+CfLrrR5CCJ8cX2h/aRnl
asCXFGPphk7wV9HhrpXHsPC3beHWjHlwTQ7dJFRMLgTtsfNcojORd84/918ObXM+
n/pjeXdUeaDJ56DJ2jVPL7nvsKhNt4zV4zkkGmD1wRqH4RR5r/QQ5xsAMrzH5Cms
CeIuRGmezrEfr31Fi3YrpZHZ6JDCpKkBZQJv0c48HnQi5mWYL7+0GNgsowUp8D78
A4hAJJ9B9LsBI2hoiDN3juy0QY/Ul37V/IzWxToM/4mp7isTPzk25eqQW5z8oKWM
rMcvEoYnrZhQdKaE6xeaUc7DBtYT1J7dVyjNrM+VLvP/xrKN2P2W1uI/UKaPXZc+
xjxnzaY55cRu6DmulVSwSoXZkdfvt9YQkhWQiDPvm/K4FvKQAK3rHaaSL1B7DczP
xS+TiO3CO6lezq0trM6irrU0M4cC4Ys/zhOclX9A87OTnIvSdUgpXK7a63DG3vsj
JYn4D8zwHNdpigOejsUei0KYdtl8cre4coAwSart8jDhejrH/mvHinIPD/hpeK13
Ok6yxLdU7PJB78DnkEjLUHRSgracmBduQSdPexvNO5ZhOei71dZjoZ5eTUMCaDS7
b/37RqnY1rjEsKCaPon8bz+nh5NSNE3UZCVIl/jk+4lGvgL82LCmRqVgaAeYFDbd
OValgZb66lXYtfDFOpkRJ8Cwq/wTaD9xiff3q7eAljM5cU1v/9zeF+cuaNjUGbu1
Cngc+naqirTAZnb1XiL+96dUvdzPI6/8xZLiI7DiQlKjOmbP072WDC3aCnl5AfMI
q799k+KtUc4KK9SnNgmEnmsOwirfyLpDRgV3CMThQV0ghHDsqnkfzUi3eunk/KTC
a+ollq35a90NMGPC777P+c1RNnVymmadiQU1F7XESyAa/YSOA1K2N48pGrqKHfIR
JHW8UiydDCZfXES2lQi18emjAVLbrGiXZ5XwH6pwcKzU2ly4Em2X+Tba3CrGFgFo
VsKhliouWlXVxAdevfNCChRT/R8lNGn0hqd45ZwEejT54OctTkeXjWZfwdsDlfgQ
2MFybxWOyzkgHNOxdF9EqcrQc2rzu7t8NS3Md8z1EJ8D6NeBXD63Oh4oXGTwaPO4
OgTeqeLzsuVR9DAJKOwsYIhxnF+mRdYw1TpZPBK1RPFvUu2pDUdB1pwnnHeOW9cB
IjonyIPT62JjGeD7rYzKHx+7T/5k8RP7Zj+r6XF0e5LuTh0HE5Y/JfPg8Zk5cqVm
QBAtm8WnPrMJ5KhcAo6E8VBsfXOeUohOo9ZhxP20h6p+NKzO8ljyzCR4wDXKW8k1
cZpuhledJ05uG9tl/67nFLxgl1kauJZHsPjC5WVya6JH/YymGJmM9++yg3ujQJM7
oGUY3FIrF7j8VNvd9DMq/u2WFllf8+8YrDpqPUHNC+I3WCPYe7Y7EZ7oxF0pQMkB
9JExgDq2/rXiX2pZ1pdLqKJrDc88pRPqP9zljmWhQn7O2yOzOmq7BjWAEsx+Gcnx
evwQmbl/bKylAvl9UW8oX4FGyF5+SweWlDi+YUjxanaK0IFAsbm22ZRDG+bupPQT
CuJTdS+S/i3LaSAYsZ7aM40zcXX0/HxgJqWbYqkAgVA24Ap14qXOuzpNi/wgqWHx
YZmXOnpb0S77LOC82F9/eZR6ds712N8Llx+qhgsSs4CdoN1SM0hVVM4rNAW9OgJr
h6QkOfc4F36nlQcT9PaX86qDOaOBJC4fMeQeYWp63BJKKHNnu9pgSH/SFL5Z2Jr3
WqyBSd2FW5BV6nEZ/KXGzHMJw+1uCo+70BDHsJ6jHeOXCbJpoiSnuFKPS9W8+TK0
uRTYDfyIvK0Dqtyqiz7KSTEV6iN/s34qqCjfbG4VAyC12sHGx3BSSpjxHUoBcCYZ
ZQJ4dqF8COfxr5UNJrMKIhCarEqzWM5aZ9c1YIGxdfKbF8WiDYm205kPloY0EnDt
rRDNCxYV3jdiJsmD1dJzHJr49NXj6sFb2rOx6IXPVgQLUN6fEPkxGsfLrEMTuheH
vBM4vFPxmolNo5MWhR/7C3Bx4AJ5FpZVpH7rwWsv6clrbO08Fnnc/ag3Tq4N2hdI
kiF9tJ70REgIAxvjejRSavPfd/nE6YHNVyX5fo/209eSKCWlNy2kvHw76LraaTie
8uGavgaAqgqHFm+AchPILNtBPHTlRiS03RQRn0uQOXp9l/9hwiyzLCP6HkAP8JQE
83fXR+kmSBwh6gT+Jf0AlLCKR1OOLtSiPop5NbYvyFv8ollZomjJ5CD621iL6Hma
goQr3jQBQtOKtIXF8PYAFxSyyxqzTFeOQj1J5FZp2xtC3I089bpd5bxNbpiLrZBQ
0Qm9gTPbxhkhE25/svLRVylIvfFGQXPbqAKGyt4rAGupDuCGH/rtsxKbnM8djI3e
I0ctkryVZIHCcz/aXjRjepB5a6A58O4FG4qv8x7gMnq+1TCuljTHcgmIlJP5EUnN
PyxAOYlyYL1A5d0FoGhBcsvedWGQg5RwIljaemampuCbke7Eg6nBhaDmTuNKL9TO
4Xf37jPs1Ko8UmuBDMnyuxaGvTDmUM9d3LHq4HNl3OK8fx1UaktiUhQoc2m2vjZy
5de/2UwjnSQavPISIKeqmyGf0rzCctbw0Q4NFHwLfQ7cVQMO2kvDP1ORK8KsZzNr
5G9jQoOtgNuws+SXlBnNtbD+4I/l8yZKkVmRDY91/o8sdXnHl6B2zQ+UpJWh+Yeo
W+nw6qSQGebHWDJBLDX4r1pslUgBcDzRKdajLftJ9oqLXthhph6UQ5PsgQC9c+WN
QcHvvb5JHfyCUQtN/tKAl6B/YhdUUvbiZ1Z4kocVjPz+lvaM8LS0JN4CQFzkemSk
lvyXe641gM7SFFoWCFWOtbfKBljzEpf4ubWqYdzp16Igp+iBTeNLkv7xJOXhKX+s
c5CHKTzROkUUfT8WsyrdkV0nZpilL/cjEdFwfXHjH5QKS7oJs+cOcs+ke7tGuMlC
7/44b3zMGWDj9gev978dDCtaw6BxbmlzUqkXMZCXBrg8nAOnqb6gIhwSgkJVg82W
c0jaSpdAFVA72+V92/vDWf8lRxUj+47Vc10FglkmbVdUWd7psORoSklATb+tnVmG
86Mipz6bnl7kUIzIfVnL2DWKPlvk9R/9mElLPTqdw1s=
`protect END_PROTECTED
