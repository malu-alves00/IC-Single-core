`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ASaHeR2fYDNlV9kB8kypz38lBCI9cMxZq49RmzfalnLHe0XmUQmkOhSrX6ZVT7wV
1btQ/39HdcV0Fh1G6fhkCMtQVwNoFGtIKadJPA8Qj6QSiR3PJYAwe24uJ/LlEatd
F6WP72rR5fKCyzkBh1/+dYbsph9CZz5wtCG6hUXoubZm/WB5KcJXlUv8yvvsVuHD
3ZfvauK7uUW6/dDZGWFehUyEIWMKuNaNhqz9bLB2txP0H6alj1yoog/OARVfKHQ6
k7FsnZJOIksw+mCt5TQod0SfjKdhPhhMPrbtjUFpHTZcRX3Gr+1xj2wZ40r4bKNU
bA0ea2F6yYO2SmZkLVyUdSX9Bot7iLvKgftZ0W4ypgvoyMdhYq5sMXf7wLOTBc52
ylB1HzDt/a9gYD9ppfwUcImZLlzTzSG2F08tx5IWKvIqQi8O2YjtuJSbJ6o0d2fU
pKugEyxBCrHf0tlMh/6jeoQbA/XUlf+2se/jMm/cQfbJn3BI7rUByX5PUR6WSSX6
8jSnhzqvdWas2bIL3hrP0mo+x/5caO8D2qVWSRgYOqTkV7mj3MZs0q24lutQzkDM
uTdKPc8qr/YFaLtTm+3FF6B6M6kMgEnTfkYXk0ZvpSdU7w4J9wLSfzSOSaQaKRUs
9BdgmE/8nJ7rJ87y635vn9t+D9jbWjFi9uVCTiyFWWbLJk4y13VAfMUDHjy/63jO
lanxCDa2HCXBDcG/tjZuj7sgAMiCfgOhERSRvv00KsfA4Ou5Ef07LNatnZkdOyGi
G1GIHvHpazg//Z5cq0plO449JqTgNv4PrwDnQhqM9mLdyTYT/eMNm++a7XfzZsIz
ebcUoMwBe+7OBZGZdc5zkldbvWFrxNTEWf5M6e4PkSPWtzLt5DO/mZu+sXPQjuax
GH38tJY6TsfMAEvd6UX7HMLh37vQFCl7IcwLDdBFOPCgKRHIPgzhDKvtXlyP0I9k
O1zLcGy/WDoSBwhly84wZDCG1ym2o3Zuyp+Yg78u0Pp+PcQxvrQrHi2eoBYkI0rP
Ukkjv57oI89aFrJwBbA6p9kWVDQvVDglfpUQV7orFwASsdtpQeX1sOQVRNvxQvpH
pEUmRhWNUQPN4kYEKVA+IR01ZFhRkRF1v+aGHh7ztMbQr48iULQwQzReJwn2FZRZ
upBcXwAfRj8M7uMKGhb8p9LP/Sh9L1rnbLER9P6IdpDAmmiEoNrzxnWmmtuOcot3
plkVX73Kzi47K62bcDxvSz0pGWi8xhgq5HrZhpJNQVQAcG9SVMOVJs6/ksfoqvW1
guufqzTDFCG21DEw11/hjI2a3161jODwoZ/Bzw+UvFRW97xmhweI4ZtVzARlhvsR
52pcJckzfnq0t16ZAk1s4bdIQzj9IzbfaJLSfg3hP+Mvf2j4UiqgChCpXwmzAn9f
mWI3G+20bcFDkM6o4Nb1Y2cOerloMOtTrtf5Sg5YWHHVGAMMBpB6DTuHTd0ndFxN
vsJZVsnMH+nQ3kKWStdhWr1wSZZgtX0qGufJF9C4a7CupE4qMr0yeNxMP6oNfkwJ
VDkjLqb2J4PfGgthbQYrSHfy4N+6MP3Qo2alduQVte6p45qc6ngoaYv7/zpd4I59
HnWGkjbhifXrRtk35JsfSiqJRKOA9TRcVL4mKS9W+DPldZii0ItVVAyK+uUWEeOt
bdNIzPjd05N93v/7Va0Al2Vf6vglJHi7mLarjQvPWpA3TtXVY02p16+yaHQ4nZhj
KEjCfzcWlbrlMvHdTWqjckA7nRM0om0E8qAUVvnKvOyG3YE3IBGyT9apI7Vyy291
oswznrAVhPxSKbMmrnKcm8ukFQWwdL6eX55o5meOvFeRN1wbewQDEmFs2dUFEy9Y
rGJN8/EpnwUdZUQ8OYOEhA==
`protect END_PROTECTED
