`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IMEen3A4G6nbuXUs3fMEI0Z2STuogqwP6k/6bD79495AnIvFk78W9inSwUx6wfUl
RqGw/f42SJpJpytjNNfgjPOGA88b5XeGwPnxqUWjcK2XgZq7aQ20nVH69001+nOr
4WfwEqYYyJomx/fli8KjO/q4Ggl8nyF0xKQGX9thtuvndVCaeaJ12nVdH8CiKuLd
PGovdubXf4v4krhzuTNOPFBNthC6knxhYt0BpgcLTsQdl/zMz8PhjjjlGXv6zUVk
D89Nwi742+zph6KN1onccKR8gLMU9AbhdMsrrl4j9si32cnpdpHVIXAxpna7aUcF
hM5KZTPeNwve/8TlRXydABNpxDWQKM0h/Fh5seXar9AjMNOUeN8eZRFLhikVDZOR
nyqons9MnoquYUHeB3xnWszQZTxgShsN2dweQpc0Io+s2/i5ezJxvbBPezPpNFcZ
XiH7ZdJz7jy8N1H3xfPzcpC+DBOFabquOxijO2sBsueWBtxmKhdFt2ZMitoBZbfY
NuXa02EtsWJwNST1Dxi23JolXiMAHr9duNuG4KSjlwcE/K9r4E+F8Xmov9ATK/zQ
YwjlBwhfnIUvJJQjyywBCNylnygjviiMRkO5KSOBB162ptNn6BkLy9RqRECdIyLc
/vx53N9MGElrEoHRKUrW+QqgukFAjOz/ZQO1hcI7nK1tluU/yaXKCuwuTqz9Nhm0
BMmTLZICxMEvWs4e75SGFY5Nkvfnr9QkwEanXN6+a9/OeltoBrL3qv4BRzk3jHaQ
GiAPc/1UxHVvu0jDC67e5lJz4gv9xOd73M3ciSBYP2qmoVo/GhpDNhiUceAhytqS
`protect END_PROTECTED
