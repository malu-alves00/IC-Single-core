`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
E0nk+MnRhroewQ5YbkTZElZOqwtopiNyq7vaHD10DzpRmNkELNFhcPucBn3a+2Zc
QBHb6KVevJBhvoNko5+cAvDmLcNvrvd1CRMprjjMTG2ybbz2VhFH+cPNI1BELCpZ
2/E9hjWz5gvav7O93O3jop0Zr3WDXWQ+K1ib7uXqoNRePxQsPJKZ9q/7+cK+bAFM
CaVy+hRvXH5TGZ55Hv0qnzTfHgwHHjxs/HncFu8aRakC2SjuJie+FVjMSbY63+Ky
e+gkAYRDn5Xsl6UNjlkA18MQf5Tu1vGH8JvgPXtPzEGSOhu2YHB3cYcCnnTqNhDj
mftzPim3NUXEswhg8XBjHBxEXUkUVwyP+PXfkG0s1s8mVGl0Sw2MnTiqFfLw96xW
auuOKp+J+1B7gJH0FATx4VEgLEvUDzyS4XX/PTYaiFaJRM4i0C1/LghTFCJ2wua4
WUX/tks4E1zefGqLQl2VKvPNc5JYLT8KphIud4FobY5biB209wuDC5jmLout034e
bU98RUNzMBfG6h/5GtaMPmreqxDOk9fESsBkuYudzML8WZiXnXsNh7OnCxofjN+B
6zuHG3xH4MU47vwBw8DHIkL91/YPHOtwozVV3OyZvnnD6BN1PHd8r/gi4v1isCq5
tCDymGcK2ojFw/3wMYj3YebqTndamwzYAsaj1SM/U1L0BMv90aWMiNXv3ACnhTM+
+Naxv50lx0eBomqwgyHfujtSUuYGfBAWGs/e/kz1UGOj/iwZO6mOumwgxXKcG6IG
jkicf0UOSWmOiq73sCwLrFnnNomWWuDq53GribGnlXEwx4aJrqGbLc5JwepnGgKQ
cgAnmDj2ElearLN4vnlQx1W+Bpcu2bXrdRHC1bT3UTp2cmWbtNwyffCVlAaaLZRz
qQkuxZPwB4SxV8DRB1HAT43rRRWaUeVwCG5FpkNKxhRbZbc6X7GJPqm3rLxHP5pp
2pSFM8l3RJlgvRFCZSHJRpm4f120Vv/SnMq4XIMff5MeSdkwTDsFd0q4sQohy3VD
icuexLAInvHDy64Kb9CEOX2ccfLhAy9bosQ1DGD2++vhwGsO0TQ2zXxDpaqJ9Em6
t9BbcmbHmA+79ehncW1uUfpRidiQ3HuQiGrvkb8cUSG0s8oL7mLPQ6vWr7ezn0ls
bk6KyJeAsUClLKGGbFBiDBm/uXa/Ab+16rmwzofNZELKXj7qhOzvxFyIoVltMoWo
Ad+zhyHVgcYjCbwzdFEtracGnvAm6Q9loEP+fSatsp2XznV/Cf2887SvVHJ1XJN4
U4IMt5OM+ayTKdjNbXyUKmDyogtKf6W0b+sT2JaSPwybAiGH3MK/7+kZ2+WAA7EX
VUy8urN0J2Ha4yLxDsM5HVSsezC1bEV9nUGqLGyCzyUOxnH6Xuw4oNZlX8DpB9K4
OdVVOduwudg7rpGwnqmp7Jbi1jcVh9RwUSOQ/CL/xs6828FWO1HAai8oS9gRGpJt
8xjXyuhWWDILYZ3xgGNdK1oz9n3wLML6rJVWB2wPnZAHpdBLqQvhngnQ4LkRlN+k
FXngVPZtcEyD6ajX9be1u4IfYTGnnFsibPmcxhyfbZH0IqOwu64+bxF1sGFJLpVK
5EBJYK+xtw9aMkvX6omXkSacJ4b3EiNRP9btvNozlmTXPI3apVbk3ipbgtyQ6ACK
cB7bKfTxjjrXNF2pa2U7i2C0InNkomknpGSA8bxtL/+EdPxZ8umSswD03wpIfROx
U1247y7+PNnyBfx1lL9Hc/YPV3HXPxVmTtsZxGYYtNhl5/auyZUfz/t7v8rpOqOq
zjoAhFrk/ctcT+CqlumqEng6pT40i86hNxD2/ir0WiIb3br21sYw9DOFir1r/m9C
Ccnye17he1RxpFGpIifKzvy6fClbzuUr1aLSOfOQHeNqAssIpjaZK/UxqibQ6Jom
yJGUEncHPQJvE5pfvFMkVzgsVoAHIkq2KljnPaFkl+agQmfptpGAhNTnsRuVQLi6
8btxNdJoThc1eQqI0aepOKM4GK6e0Lsn7CUgcctaJTu/XFk4LJdh+YHoqoLHFp2l
4HjAHglBzVCUr8n1zLI41MDybuHKXbWlK3mjbqvruOv2GfV38yBpsdF9XAHZb/VK
2YS5GKpadHJtWfWMf6Z4rFrj9FfLPcgZRkVVm/YnGabVcVUaknLL/grdd7lDsQ7z
avurXiHjh73SibNymxTCdUOTVd2j5XTShtFHw/Joo+pYzoaJpQgySHve3DaprLQE
H7cut+xzNWNHaA23LLTBOv2BBmMjNG/a57+Eb9FuqEIgefkOVNcEqWvTGqyOpNvD
QAA+0g5U2jVtsbfX6YUEPedgSD8vHuazHBH7EqdiXq81V7V5Ux7LP7SB1/qaDpxK
qUlj3euimZEy0f9A4BLaHkER63zh1XjiMT/9oWdFsM4JKagj0UTN55cghM86bBdl
Snc2g1fvyAcG884P5AE0REuE3Nz4DyvuHTPJsaxkWFRGie/H6TUN0YWHA8Q0Dt1V
xWoqqFjlH4bXP191Ppx0bW8ZbGFK5uEs/aF8gV0BNbG0kNx0rlBoc3B7tbKDQnlv
nmuU0SqSGKdfs2MfE9El/Z8Ey3hfSfytvqjv3W+IHz1XMLh23HTrULa9EfYZcEFS
TZIc2/e/kDhdSG0fHk/NCwDCyoZwMIyovaOspDfufc2ObSus7mt4q/hqfNzWGnHt
FGTU9OpAC8m4xvisfbjx89JIspqiabZITNlgJFzCBBAVXtOinRsoctbu9drsAHH2
Fs45I/V9URKtW5FSnLY4O9Mo3LBA1GwLHrzeOAuAbWlxhSVLmVOoNFcvLKF4JZji
GmKKjb3pYzgUrHO2yX5hAIpYLXWA51lpirYggoMtZc90aclqhqMqqawkPxbK1/RE
3zINmD8/B+hFTaupl+D0Yu20VAYFKdGtJ3nL5N+G8R8rhzPloxrlEFHfvzfpeVj7
Uu8rZvr/ht+VjU8P7YVjUdSchi8eqtyAnx9eNEI3dSc2flgRfkwisv4KN+ftKT0i
QOEZE2AjdnsGP9bUFiTd+ib5nTaas3eBtwiqENsGbos2EM82hUwFu2kZLAtdT/jK
FkfKEtXYECoO+JrYdwmXRWqXCrinH2BoyANXWp5p6air8YVQtz1Wubi5lBYfxQNC
kVVNGFHU8MJeEDc6+EL1L8y0/x6Na5EeBof5dlMCQB7OL5AYCV/5BU26hpNwFc9T
ljFOzjiS+f7rcayslN3k910tL0tA9/G8PsTqhuCD76TTlJMYkgZyWjNQZAb2PTL8
6xLMrRLuGw5i05LP4v9neOYIxelpTAol513zZa9GI48rFlOSqhq9UxMZcQKAvUaJ
ZMYUcp1yeg14owfALo7E1paEfp4Ho+xFIw0ss4gqZ3jpRVU5NqbOXWgih96/IVoQ
UtINqKDFjXglaMCNvqddQOjWQJdNgZuVx0kcj89gAgjyeGlvaT1/QbRkr9dyuvo+
ZW1RG44Y0tlhqFPZEFvfX+ifidBFam0d4TKjYd/GvBntyEeXF/ioYsxEPq2dIikU
zLuFVUzK/WRlJDy4iLPKNV3a4aMkmViTD+C8bcmC5Y2iR6cw64eDhmGag/00t9Pq
IJaAbtV3s7s7aTlHp8H9sR8HHsAvQ+PbNPUHJ0Q4/nZ5dG0foAuXFbLKoFzV59A8
rbFXTV1mWnh3cR7jAgkA1teZQO0mQndIftuQ02CN/u1TmyEVh0ySwh6Z/gVNLFu7
Tf9BOqNUg7McwckAiyxIgFGml+bjy7Z2Nnnp5Kq0IthQaZs55fRlqFDkQ+pLqv9E
Mpam1NNJB5mYMDUD4Qameh2qiq2QDioFeBRVuSGfZjF3XFOq4YyMiuA1UawPOexi
+446J7/UW+BNrzZGXh4UunR2k7beAX4sjFJEsf3ngY7Ybe/XkUgYMIaO2rf/rXri
Y0HAbRDSLJD4uP3e8V+i3ynLsi/d6sA+Vo8PZ7Wb4l61Z6enV1OaYmvJspAQGElO
pBSAlwzXSdCsfD4+qQkutlWb8Zun8NdYiS74oGJ0wvP/uNlfDtsKXY32kPiCESpT
8A1tcKLYAqMnBVYZm8wZdJxI8rCAXj8fc1S2Gd0+47pg66G6p7YV64lRaunM2zfA
UBxQusKUWr+JqDR9PToGjDHT8lNod1mFYHoWTM52WjARl2u3OnV3OPUhds5INVpI
4EAed89trXXhjdQzwHwc1xnxuXi8ze9vgjn8Qobm9FRpt4MOFcTXpE8ld7X60SM7
m0j6QnVKLnTpNI+kENFgH8FcfiLuA4ATKi7MIIAltThGdi+bmfIBzPuGzVVgJvJw
`protect END_PROTECTED
