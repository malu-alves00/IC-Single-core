`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4/7vqkPei0zEvEISstEg7HaPvpn/pnRYDTQM3QaWqMeFYyk/LjZ05bk2Ifx//2rO
Y0pvTU5+J5fnPUcd390BTpW+0qS9Gydtr0sgsf23Lf2hHm/PPjaTO6b1E05HsXZK
3UNAIIOEyWKzknX8HtVOgcfBazMnrGGSlOTs6YA8H2si5cfW+vZ57J/Eu5tXZdex
gth7GE8Q953Rk6bwR1BENbXuTa63SrUQPDnuZ3xegrLbjGcYbgK8taaNCjngxvwA
5A+JYCBemEfXEXrIsxxNsl/y/+5qRxuneNoyHNr3KtOwtyIWT0z70OakgvpyKCbi
/Piy/lnvzSMEMW5SqfnflmOa2VZALyJfS0aLk7VNWWbDOBdtjYf5EG3BzgfIcHq+
On4rVt5lRRaSSgk0Y55g3e0gIh3fDGreGyJOcSvIZblorv7ZKx5sR8WmfUbcVIDz
KG4u+5P3UmTAK3W6PzNZCpfBL9PMdVL9YqngeMKxG0c6wQjov5kNwNb7taFrqwgI
gdWZEbPZMWqolTor9pHgjuQJpLET72VyFQPmQUwAdIS9WbgpauwssLGgl4dqGAkv
wnSWCMsNTJXnv+QkxbpUyhP8xQfitSnz+18XvcWE1FsbRmLDDxmtxIvUIsBfYUIP
+Y3sqbRo5j8LSW2l2jlDPe50jfj/YWMIvN07VR6bspxzPkUCTsDOdZtzGDF3BhcQ
`protect END_PROTECTED
