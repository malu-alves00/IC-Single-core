`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hLkW3zbAbTgStvC9VgvVYppNHmxBR27rT7mVwdsXXK5nRh4WXGZlXT99g2xZLfP8
E08Z8sNSlPLBr9xUUnUGdvTT8zCk3KYuSj8zRA4CAqwUC17QGgNwPrCk2la3g99T
eBFHaaBQW9D0gMjs5tCYPT4kf8+raDhnq8cZItf3UGsye2tJcfiCUJAMBUjeqBK0
0SMFSTyAHCxXhGtgituGH1e0SvGfsgw7S/hFbFGRx6SnKkuMnlD/ek2900EJWTtY
+YOVDN0oOoiUMw7lWmoPOmtHSxA6OsvG5fdL0kDA8HHaYcwYSzns+ZObfuu7vPwl
I8ecgTt1INkc6xOAFIlXBUhfRKwIQrRUF7I17AuXE9OmqqCUoN133aysQ3M3pBlE
eb4/IbybBZOTb4Nzh47sD3660HKS6t35tgJp/4JwZ3+Rwb0iSk5GxzcK9rn34sRm
+TfNbd6+ImGxhcWnrWh7W/l4fIWyKrTpUZCUELAf+Ui6whoCxRgAqDrf/nfMrCZ3
pm3T7ixLJWpcRFzqUfTehAg2uvvA64qiJOF7rSldIgdHVPI4nIyuMxJc8iQEv6ak
0Z6NGXvgLVE4l7iOoQTw2mqrQHpBeFxQVKfM+XoJgtDcA7XPczS4T1syA+59tIyu
OAtKOuVZu+dVHw7+3UWweCHyNo4pgUtnhYC0CpmkIDV5XOJFh4jQDDQWTReFlbtp
VlRt8wOzxMTQG9oYTvXXmFYMrk9ph69U3QmySRTXf8c14d3do0+AH+bxL7DChPaT
K+eKOGRyKKOtUSUd5Xizzw4zabLxVo2Zhkkbrj07L5YX/A3X2uMIomcDBlYlbf0g
BXycH51q6gCxpFPaVGBMC2EzdBcOjfwKerYpV7daIQKgyKARfy2hgIPpqZNQaUFH
osjXBHuV8Ce+1LIy9UYzvPbVcJDRWXCVq0jYCwDqty7pzKOHwsBWS2Wp/TG7gv74
`protect END_PROTECTED
