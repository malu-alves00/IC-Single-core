`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lwvIbJyeznFJ2Ntfxv0MbvKPRiXTryD/Nlu/4jMdBZJ41WJbLGIhWidQZ068EU28
UNagJgVc8CdH4lBeN1rhKnnaMVf3gpAB1B6A+JfTELvTASfmbGcy8e3u0sr+qWb0
xRftwtY9tJCunC/9CoJeYQISnh43hf170OFvrQqzJTGTHZRmCuBfC97XQV3OAGRs
ama2VMnTxMSsz0KTjfLKBVtIXRsqtu5h/lbtsyJ6RVyLc2DUJUUYCsWSdcqGWVxa
4QzatfB+ja63DatN2LDsS3la9w+52qcJKacpH+bMDuLFL76VYEU55IxkQF8nj0gk
husn8lLhte3L/65pIjgV+SvxOqRkz0ESECgeBLtCBsE/nyiY8AwY1bPNbTZWomzO
j9gB/ejiRTMQPEsHj6Au5KoX4hc/28HFKePXRqHKPbF1w1rFjT4mMkF2bk3H+Tj3
m9I13z4U40EtVyi7TW6xLU+Dtcwmt4Dr7QjwkytBaug5zaq6tRwgjY6a5mJcVORt
3ZEiD4Khc2uN+RU1z9fh5m0QMhr0dTB8P0JqFcnamh7baOTJ/U+crKYaJN1GFeMK
SK0UCNknTHu4pqiyp3PRu7H+pCSNQl+BxzN1r/ZcvYYYLmOTxbiOdbRT7kiuYG5v
O/4IVUUHSaVJw+vUjZ7De4xxzyE7GiXwuAu41QqHK4EakGenju2MoxuPwSq3KLQM
JdSnQJ+tAZmSMDXmz8z8/GYed1B0ImPYiHCFRDS+jefdxZrIWO4IwOUtLWT/Q6Lz
zfF4pj8d0HkBafrtJvGCeYenGqXssAF6TGBUeszMLRbkQh8eBSqfpFLVnPLpZxP6
9zsCuGCTyxZ1YAOoInLVNCagsD1tZm1ptHv9TudwbTof3KWwkf4GgUYJ5zgWK4p/
ooJKHFiXHtJY6rioplan5kYtAydG+t3JlRELkb9y5MUx8ntL2X4h+wFxZlIcxjjo
pbwCOqkCGPPpOI2Zu0cVRbvoggTCub9LCWgZ0BMw5guPCl31WhPsPMRb7B0EbuEZ
F5pUqyusErazWSnDtSXkeV8MOXoixTFldCnf6sKNZ9dRWRdlPhxZfxwglTHUrOy9
FyEywRwqgVaZ7uEktctCz84505BYKZVce73fgjV2yvdOAvq04rh5RiOuoRd306kC
wxuEhqjYBaldjq9YFsQ13zMkyNRNIXT7TMzgfg0LieQLZRe6bXzs/3nJ0ZOx/FgQ
bGB5MwMAaYNElj89Q3aEfFvVePEBWR85Af5vqv0M3YrysI77aIafq3zMFE7sCPsO
4Gin0OllNJyc4n9QeRgNVWl5MMh/uEnOT815nCFBfur67JdWr3pieDtkm4gdLR6c
nnm7JLzgThu1qEX9LJd17tdTHynSVPRHLFxaXewCVPEaoOZu9iHpa1+PzGAK2WhT
Ql+1WcUizvzYLiPVCHE1z7gITzeXoXh6b3/RdwEFvNOoZwUZ4Yfk+XQjQWXSsE5j
a/ijx4PpbpvzEqCuJSkbhJYsd1DJerv+PoOmsBvDSAUkA5aPxMcszkU1J1ucKDUf
1I7DMfKOlrtyCVJPNDvQrKNB3t3H6zU7kLd2kL0+EX8aRIoUzfLfyowB9CME6FvE
5Nw4XHjPzHTWX2ClJY22eZHphaYGWX3CpBrtXltu5r7hVIz4sM3/74kXeLDCixUM
lNsIXLBCYLOuIfLy0OxshUVsHpgzRX9GZ3SIwSAfa10x7UtgbxAfRRXW9YJJQXUn
xOpOYGTSjmKF/lHlKLok3um8Ko454PRi4rKivCSVxEWpWclvTbly3P9X2elFO/lC
Psb6Ms1EVJczBmwf1kD3aRtc64jXxTkaGmG1A6GzjWBhv/os0F9m8bapItAYDf2k
3rohsVXfB3Z64CwV2GZL+PBT+fncPgFZipVUFq0spTmtDf5IB7Fa1AaG34Ou9w4M
Tye0LxJ4eGO4K6ftZx23YYtdfYOiQJtlSsnxd49hY78StdoyhxwnWEmuxqfs67sk
DkYt18NU7EEEnZriujkUlIK6nif5bo+PcidZDhWTEm6HuImQrGtb/79m31w15c8i
VrPcPf39//gWHFxu8EOlT3iAUexcKU/Qbo1Ri7HiCV8JH8J6PSV3zQaw3vRycldc
gHdkvz8Q9GIX63/6lENU3hgCukjf3PMsFVuN2bcU+JUswdqNF4Lr1+pR0u2n7rxg
lRcHAv0S85056RQS1OFQke9ZEVeJo08w4gksLWpDGMKnibpQQ1uK8XfdXzLWdS3h
y2e23NPFPGITT02TA7gv3cXUs6VQez11cHep9evGDE16q4KRD/jmt2aqAKiTYZt/
X6/ljL84GvcyoedI/Fn7AG2EwUZp0hRXbk7qDHvyvgN2FGChlTqHXlmxs17cjPG/
h511TgzgERKHRkv56a4M4/Zd1omNYpkY/Em8Uh5RaqkjDNssW0GLQ46atYC6eRVl
io/HF/WJCxi6D1yIt/1+DX2SRidSkDJhG+TurdlqnysEt9SkITbDSaWXKj1M9DC+
p0or3Uqc3jyO9CY084EDSDntYhcRdxOA0P0HAetfkiAcSUj0KlHrF3D372MiO17S
CZ9jFkCSF6Zmbee1DD3Ml/UjLWlEdW/9D87C09zeHS+5BHrzPlWBrYR48Kk9ZGQZ
/BnuMVrwXh4jsCT1KZK/vDohCyF1yW6sPYD1DrErJ6j3dNxWI0ubFDU1dbB6c4en
H+Te3ri8QvjLM5Go5AzGlCcMwX4bEkAXKHffGe8Y1IvLyUnFRgLkmCfLcUz1ybNi
3cPK2+ekGy6e9txCR01LzcivBHqZ/RGgIgqld8l9c8xt37mCkeItuy+Q/0ewA6aL
T2aYLs9zl1QDtDTYui+7k+3f/AzfFtQ/Suwmv94LObjeNRZ8dkHo5pSZyPMYNEIj
1ngrE/Fpl241YsjAIyO45NNyiuev7Gd28vrK09C+GoFKPqojF1aN/nhSujDmYzAn
ZtHd5StJ0KBSQjgczao50EEeB1OssZqGq/8o1w+3UUUT9RdidOo40aQkrUG5+qRT
7Vstmw3qLknHz+9lhFhhlr9cy+YiYjKGxgF14k0mqw56HaHC4rXZZbkcOSJW8fpv
e9PoBThXlRMsSuMT16sk/lwg0/4uRzT2tQZUvu9JHjY1DjWs6psPH8XT8L7S/Fnt
fkaHjcy+nTu2m2hcNRssWa+8JbNBFK2lHzBNKl+dTfQkWjvDatWYj4iA37ERDCz5
Ax4BI+AtE88SWwfWuImWOIUHCCyZonYoEBUcsBjE52k0YP3fDUQa7TwxdEg239Rn
I0gyUIh6m5g6AM8QJLxz1X6N2PMt1OrpNkNNfiN3hgaiWIwCSGHICq8uToAs4zHw
O8z/aAfWS2UgITIYh5aCRyS3epv9Jt0OOfgrnHWMKsfLv+dQDFwowgPMK4g5h+Rp
OHyWGs55URIvJNG5Au32vkUCxXSOaq9N5VJip/gIFrCXRLQG5nky0Mmq0naE0Fh9
Bzg2vl1wUaRcQ6QfaOMn6iul7p4wZnxTmFRr8vNhHiKvsuL0EnwCaF9FB4QTpZ5C
P7tYxUIzpcnqrE8ALQxEioqMNTX7PrDRgkh/fNVmqxN2vJAioLg5mMTXxlk3w1ka
o5CM/aN5NPHwl1ll6pthDQ2gzG8A64Vk3jiVvTJCvZWzOo+TlvQxJCTx9Gewjirf
K9zf6lxOg+hsi/zmLHT3vgpSmC36ecJb5dtB71+hGv4R/2gjjZXFPmvcFO35x8q9
XmhdQArk0V6h5W94a82qEN07uVNX7kUqwgaJvQX3PCVintWNuFNkf8L8RGMRV+Oz
tcOCNWyEukNyb2+sI+BbjKMvIOs2GAIrGZ7LR8jRdG8wqkwhGfrwgQNm9A8rInmA
gLZBA2SJx0cDUhcKsAObwCPz05Xj1pBxAarGYREDieNvFFgBZolqv0H8bau1HGDZ
dnMRlPoBImhMq1A9D3N7hxKE+EQSOw225NlMn0xdE+NoW0qqlqO4oqNND5YATULk
jZIS0nmtxlh2lmLGOSkW9RIR7CDGM94dd1+q4GEU43bDrVHpJ20vZkfDB6d3SG6P
eQXOo5g8OPTZcMHunw1kdvB+eOk1bH/EiYoLzHDwuNUymnFsgZEs+Vavzn+yrnk1
ZaG5gvIyhgEViLuD4h2dgMt3y5SxyLMc1/D9uiF3BmpowtM5iREfusFtkgrN2qk3
egMSAT3LDuK7xsv1RUi9mIc+aBmf2NEBE32MkHf/yZmis21k8eD3mQjGr3xrA6aw
R7I2nWUd1M6Msrb9ApKe1ux6i/2gce80B6Jl80nT87SDU08GDMPhMB6O3eQYyPX+
W9J5AZS7CNRvsMyHlIUlKlcIab3wvtCmuJITCPwpWu/AgBB13wlippBPNv354acH
WNfTI8Qktl7/vvvTQqE4qHBd89wHaWdG+vztiQcJvY9Oj0A6ZALJ5mVdsGBWhVjV
hVRQhDqsAYIcjZNjTvh2WZKZo926AqKZMRitdGYcQJetC/sgPqEougaNp6MkiWSh
IjIAjAW5v2HG5CELh3IUbnCaV9XavVJhdWvm8TBI756yVM1XMxyO0eu2ZCKft1uT
GR8xI6ZxQ/aAEHzeuWB2FryWsSKd/vgcHfCYw50WcjI48zTvgO9e3EKc9/ZJqxHQ
FkAkL/gX7OXz+Bkdr+sQGq3DsxWyY4RfKyu2tIgjHLYpxDAtN9KhmFFk+5v05b6G
GTHar3ch8diLf9EpCtYuy9J85uxFd5W9Io2kvYXGcAV/EuUUJeAhnSAvbD83qHpV
UKgxMtCBFkiHPJjMWu2jJ7Wia2oq7GzB5glMHyk8rOhjEBhpqloJddkodIyCCCxz
8Jgd4lsZRdRZWhwXq2LYsD9CVLc8yrHoJFc/pUeTS0O1UGb83r3mZCPmNAtPkOGh
+8HCchKaXS4BiZ1GntxImkwDjrYrDs2b46Rto/W46UzRGBsx4xydsu42oi+z5054
fKXt5iAI6wvx1yabtKogsuAqE6vvwqtcrrI9zKUVQzw=
`protect END_PROTECTED
