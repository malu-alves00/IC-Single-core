`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sqUu9U9L3EwVLNd3JzliYZAw7+n2MOeAWmAr/UWREgFjRoEi0F9nfng04jh0OXnj
4DSJxfHZA2Ro6/hCRfowPYTPR676YOfR2Rfi6I+KdY+gM8qgl4rZ3c/4oWlAuCvx
eQ7cBU1kOnp+ZvM2F/PBQOXaJqujzFKzXcieceen5cHJSGX8CL+UqI9QUdW0gdfU
SD5HceunCwhBPeV5QU4qkec8KGpl7RweqCy/nU80Jtlf+L96oGji9aAeRrhyBwbT
vZwvnyILaPJIDoMC23E7+icXXgfOCcJwQQYGiRBRMsQeug7qC+3yF/1CdV45PpIB
91vDmSsCUGL5QIuQa5YC7SCFpfmy/fHVJtop686mQyfxXRtpOUcseEBGk2OQb3V8
bOG6prOXmNV/3GW6zlPydxiho2Z5NOfqNnHSSg6vV1WVhG36KbRSOrCLmOmBHfGf
ntuhE4Oq8ZekbyWainIFeQNTuFVnaaqijRuHkAZEBlNzYWN+C+h3iMN7UJWreufR
uymG1GnhBDJaSZFxzccQlM8LacPZT7X9Izskc1yncxL9Jp6ujhg+yWpiO1y/TwRN
mybJhXDea5DeeecsH3iB84easTVXojcBXFdDgGikOtTtFrR57+ivY5FULM/11mg/
QhkEac4mr/eFYqPwvEyIoKgZHvRY9GMSZWwvDaGr0fzEUcV3MXzVyjj+j5LdJHwi
lJI8jbXzlgZIWKyn9UJ40Axs8Y9CQr9MU7vLe2rrh6s=
`protect END_PROTECTED
