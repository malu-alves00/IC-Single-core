`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9J9rDD8xQrG9a+5F5QeITnxyKb3t7TnArHW6h7eD4MEQdnmaB40Sj0whcaWNCzgf
DPnJIs1/GWMZdFM2ZN/BCQnEfzD9i4MoEeOjPk3OTYtLMHvUIfCOz47ChyuGA0YA
iN+jhVBTgNwZZ8igFX4H0toqS4u2GjCcGKepMQmCTSEPimj3vVSYwVwweZIOnPJd
qf1CaiDT4c2/5WJvs1EY0rYUxsRdh1i6XMbASCN2utns2PT/ludzKbUUuK0d8UkP
SzoaEBSx2QEiA1GV6xgvn12DuLF/0VtIdZC+h2aggfTYjSgb8xKg6r16a51axYHt
OKeqeEa4SGQ19hjz/hSkKO6l3DHpuv1aQXuPHTRXe0GHACVd3CdRgRXBtEtrRmXP
iBincCmT0IbvcPSYYhGWFZ5azMCua1ZQNoYONB0CFTSopqLfXr3FGymfDGqjwbo6
EG3jqGGjK4ALceaxqAY/Qx1aiEr8pkdf+QZioB+br/ekfjNNrlkogR9tKvYH2kmq
jGXIPr5qDNiu5Z1co2yThYLH6n5RFsw5zciL5LmJrtoCr2CL0vHUWmqIMiLYMz9b
VUlEjE6GaeOHZ+wmXh0RjHE3kZpYlfQJhtdTKqt19UcRb0hZFNoTRUveqesEcOnM
N2bePQ0Ckg284D3VttpD2PA14onV2oSKV0InYvnsa6WL9TEbVcZO2p5KFYwaLOFC
lqp8Nwh5dKVszVMxNsNK8PIR1Z1+shK+yMHcPY4TugVHeTvNMfyB9yn0mYR3+F4f
cs3MMEPJcKtgC016uFEfpp7nVegMmmtv2h34rdTEZYs6HXyE7kTWjFXAKqpuOD3J
GPl3REUlHPswmpYrVzy1dKrH263doyIWnTXMU5Nzwpsoxxavl3SIaVOEP/mCgbLW
vUk4CY+0ZEDSvp+sW8A8hp3gYMfXydtRLF20UzwEMn2zbTqzQt/pAcvdrZGC9Do5
3i9FCaWiZyeDHyYn1usM3UdqRvPCnsIPT6FRwtC6pxLMNdhuuP74JvqUPsj7PmaT
/Fycuj38qaqwtQT/SuhOnu3t8toGlp+A1SAhuA0lZbhSuBpBrhQ0OEco+Jbqa9lP
jcWWcsnynawmMauTHX4txHoeZ3+WpnKvy9FfHeLPQaaUuO8d6GGTfgSJriftkXSi
gSJfplpGcvKQCmqbJZcZfrJYH8cnTf9Xlwu2en7yC82ZIM4DwEPxk7Il0FfQZt0z
V2puZKKjd9Pkg63EMu9OYapzAW7NRppdysGKWHyXc9Oh+RSROAp0Y8w7in4nZFvL
ZW9AdFuLnbbrCdAdhZbXwn0YD1gRDUcWIpLPC7CSmyCmIVjPkS/SotPUJEz1Qimx
iKOLQvOI5LLL5nN5Kj0oScooxgkb21rd/A7QYao9rU7JzlwQDXVANHPhbbBu4DLo
ZoMpQCHGdIhlmxQMHwcb3WqQQ4R2UfEiWKkU5FpCZkBD719E4japtVx8yfdERtqB
ycUimlo/JGdYwF8q8ItLutYKFU2R3sT/qEQi/CutUYjdJfpasPO9DATFCVA0syZc
CgCW1GDr5lkeOKm7xm4ZZoIJfRzpVGGZBb3mpIrUmPwpwCg2ZmdjMT/Xce4fy884
twSyRUaawTOmkB/5T2QZ9USbCnczlziwPf3EMOGiMzBu9ji8SzZib9YBK2r/ez5F
bv5TRuAxZksqtD5wppSE6FnHvVocPrac87avUjw7LyudrY/NNqKIZVkKmoSFUvDu
a26pKIZGHwZV/VKggYYli4TxedEwgpED4I2ceoAIRY72nKjbWA52NLVRzSaiWPlo
RfQK9boIm9FdqN6iR17n4FC3zgKaJEHbo5curLsVrEarl+oZCg/ERktef4YT1NF4
RX88c/p3WF7YrloWogoAHYH3gptjbW1WuUIBfasURT10BiuLEMFNkopY589DebDF
TVHIpThgr6YmPZg2YpW8aMG6e5uZaBQyU9wKPXWyH9BulVJdJXZ7FrFWpQqEBYo7
NQdwH3h7oACYd+FVs8bxJhn+dQq6nEX+N0agluipbBPDE7xK+5JGKgkWS6A2fnNo
d1A5umNt/NIljoAJeFCjgcrmHYiUUvwsVPewb2j/N9NRgnN07MuJSoXGqZWtdE5+
qwB2N7g+zw53UB5562yH1xSYEy3nijveg7BINUQbfEo9V69KZ0gfZJietYmgLbRh
/Kp5sYmYwdwsSWbfLeqDJ5kAnM21o5PruR6nQwM4J5PCOCRWIhZ6nc9gYncDPGza
6aA0fWsmgNmIR8dFbC9S1m0yZH7UPi6NgUjM7BtN8yJUw0IUHAQ797+RBRdZZFqw
yQxeVk+Ykci+VtjNoUhaTx92f4zxuLm8b1rnyfl3JBuShgCnDQtxW9iAKM5Mz32v
kK0dxEb7cTGrwCxuXfKx0G1lGrjAJmHN8KxHGsbJQxzcpkCgINjOwBIr7xvWXO/R
cyMfZrDJTtQIcDyufJZNxatmxWUgQcgtQ/BSeLULb9bNVqhlFJi8OF/YAgFGfXKN
bkMvuGkHOExJ5v2czVCQeJwtge7GtSbLyfnoj0I0PPw3RPhIk164ym5ActSy0gnj
rXbVx++/sn4MIXh7g00Qj40Z4HmqzyvUIvMkXTwgYoDZwdU9z2S8RI7zP48yY0ZL
ce/t6Cbk2kk0uQG7nwMPLxYr+sHXE92gik/f2ekM54XLMoONiB7n0FigqDvV7i8U
4Jbl+uzMsfokfxBKL24GiW41usl1sDhiQRb0iSe2fhybIc7soH2nBiu5StTFBX34
oRtMXUfMMYJcw3ugGR/3Wk+t3JcxL6pc8TAdbTZX9lJAu8RZ9uJr8LApWDl5ZXg3
lWZEgLM0K/GiXoekVRx6MhRkNvqyouhC5539Y5ndyZgEsmqDsS09t77hM6IxOK1x
yJAbGer0H3yL6zo72pRZv3aCAgNfLzjKuxxNT0463E2M4bqPlGSUyooTKHfsXDQr
Op7C22axvJIA1Veqj53Hmv0VpvOBUaH+Ib36CutmCFZNB7zSD5T2xldENOeNuL+c
jMn8fkAWWD/T+cvXOu/Zg0l+NoFovztSR2LC97xklCBG56sFLPEqeX9DIGof+OgC
vYHjQSpffHjPAzmOBpjHggGOVlKfnq/YPCGnHGkhBD6/D/USoLBeUvI6dfTRMZpP
7Ro1Dta7WtOY316M3uGf8CYkt2fv9IgdFWdsCCSLviUspsRN+8NF4bIzBehx287G
yws1ttPuSq/iw2k57LDSeoDyxVzFJd90Bhk8CfrZjYmi5CmCiR14xcjM+Rqh8P77
r/bTlWhtkXz0biOfuUQF8tZPgp3Co9qhuWP5yEF4MhfqUEPRXDg4/EfE+GWC8f0m
sgR9OFBGC55N7cjmz+A4k8rY7txgHtxFz8/iDYcCROFPqcHV18he7LXgCIzDtfoi
3QGow8fTUHMmcFYexBBoDvPfEYpkbyqwpfxyfy4Rf8M5pVTVmqgPQ0XQASeIhHYh
2Fq+qf8IYp6ShSgc7PnQb7HY13pNa/6AHyAL+ghrJ77CbqAqcmjSEihGlWRC56wy
DudaQChB1UByvncdFuBk9zxTgCAmDcSOxhtFBR2Rnd6cW4VQnlDMv7MOa97l5f29
amccn2NCc86EHcVcjgKsvgH6AtTxaD1NV8pvf09evaGAcf7/cfGGnTcF8wl9zwvI
ThaXeE+filQvW+3VahN5fY2KW0Md6kM3nt2xYwq95clfBY6Sp72nNUnqAtqOZlYz
Qw3+aSpNirAeupExZYEpdE2WwRuHQYDtuLdHCXapQrswTkiFDORCZJ7kkBBihao+
tVAqLnompaQIjQcqV+Xg7FscABdHO2GJ6/wbkf1iZrsOEdGE8g/Znreabm4ZgLk0
A9ZCTv+tuggWq+zmxvgFahe+C//1IhNQoDmrH9I0rxOtAtkoYSlzRfwsQWoFR63a
l1Eozcl0LsHJielGghDNPiAk+KPNEvKlp8j804c0ynnes3dGVmq1sM9JwnhIcjPO
qFav3hoUi9QX//GsffGgW0KFf0KPWgafNzc1cnR/2j7THVhJtsFIkKb8dRBPjjdd
eOBagBSW013eI0cVBN6cIeWSxtegfQ5fDrWaWFd80WfFxOGDbLKymez711TUw7Pi
DUyhIJmehtAXFhx1UTFRTS/A2CpmfWYpMu2Q7aKu+Y89x9y8JarYI6I8zCOTKXnT
3Af1yt1goImkTcr9D8LHuUF9zLl80ZN4Lwj8JU7CCfDcL41DEhop42QpCNN4sY0b
7Mn3yeFftssiZcrD2bYsn8QDctI7oDZvbI3xZxvg5pZkOFsFZdaDO+NZkZXGm/v/
g3/e1KLEapIFn/aHiQ3FuZGTOOt3okpNTHaHNLo0CTIHOh67kdB3tZB8PfH0MdtU
1qgrnTP7Bp9QhTdQDHIJMEdzvtiaVZGMt6WlZnwTb6v+rfjj2lASchp7ixi+a3ie
ApN0DJFKRGZZ/X9G/tBPVhH4nKfdjzwqpFUkDnKYnMEVuouEfe++pEWz/ucjXQBJ
gBlcXtgVHbZ98tzwdGrza7aA7wEQ6aiwvAe4AjozJabZu73XOMDwv32KqyP2VoEM
GfnUIGm3YZ6XTpdahCJTIeNcO7lRhmlmxA6y8ELMGPREftPOUl2E1x6uJ1k03gS7
esH5xoOmtb+aLzePu+7VV1njqEnXaJL36MBnEZsAQrmZxeR6LOi7gvKX09LVobv4
sIvm1NJyKv3h1r3lyRaz0/3H8GJvBp/+Ljsw/1zxng5yfTmKA7Jw5rcRB7yU72eH
rP0OhSaEXJD5ToTOr3jkCHLzm28ZP8dPKx2hllQ9S3EAbclPTkGdH2fzVlyj8gmS
LHx1QC2a9GbJsTwOr55kP/3wcM7qY3CIshmXkT9+EBivdv3NBo1Lx7OoXpVVadIl
CZaWIOqvw2Mf18u9fRdVxlaAAqGjWUhjTE4+4gbjV9dfafvS77Jrb6ClYEqvOVXU
mqO4EZo79HgNnahTZQ4qwuV6GomrXhDq4orHzhEmoV60s1s604tYyhQbOGIzdCAe
AUvYyJmu3LTXT7dGSNWoUJUaPHYd/jy4ZKe70jJCoTS+vBj9wcM8ZKw3qfsgdJwU
aj2bLLA5yJ6irnSgRuJ3VMmutTvTYIE4A0Rb0hWUgwcEs+aulF2PV5szWXvjVmuQ
kTXqjFB3AiTeK5s6uiBlscgyAgOBwvKli9AeElOaOfTAmNljaSIa2Gr4iOVR2L1c
ZsyT5/cFiE0qgqAjmTWmpV00AVYqqIenWRIQd2zKAN7Lvepe81b33sxWWpdxMmC4
rCccPTQfZZa3kTJ/3s7H/ZryyqGg4qPladuF8r0ZR6j7G7nD3eHJJ4UcNoe/aLrN
GzmrKh3ifHCHw4WAx+VThKcUtOmjJtV4Gk0c1PEMjfZ4MNlA3tpUDZbouKV8fTIs
hjvcVqzv3i3O52VX/z4MOl4Om3obCaKnQN+7x5gn6Zjql8+ojfsDAZVCndPeZu1z
HdDPLuQdcwInQtmunVqR00g6u3SlJ9t9DDmYXvARDKRUjLuyIWlBQnMEEnc1pjuC
czXtqbVCsgCPoQq5QPqztK6VP79feNV2KmTez5RWNt4P8wzczLQ9TwiT8CoHSqmn
o/AgOhydKLJnmhIIMnb21gyM3uXfwbZdKvbKadWm1lZ5PEuCdr9edeyxwixvSCc8
HpeB7qx0Thz1GHN/Q6pE6q/1rRn6RF0B6Jspt9J0Ql9QQMW7ibLSvD6HwLetxj4o
NZlskjunmEhkyoKQK4HJfa34lBoNUS3FftjHbYkjh6//EGfZv8b+fMwCLOShHd04
V0/KwwWPOgE4NcN51+WI8laPhZC37KknezlZ6yF7uEkrn6E04SFtHF1DxXSO938f
oOkA81+0V9UtLe1QzVC663+6gOAkLfxkRBqMuAFH2BJtgALnhs4keD1CRE4p3ZH6
s0IBVO4Cpn82Z7Eu+0C0skzArzawbMrCQZhAZb7zND9oJ8MWe2VBkdGF0D/PlSP+
msFr0vH8j1Kb+Al8UTYPAIxcjv6h6ZRTDPL7zrAcQsO5hz2iZLD8A2RTfs0t/jeC
S7g93lfPuBvFMU9z8Y32qsb8Y7EBEp0GAktwmFYEpzaiHM7K8shsAPNLI3N2gHXF
kz0lUvjaWFSbWFCV2IYa7Z/dZJrAgD1IY2bPb0GgFm3R/ssro+h0UWCoCZcmg5WB
IMiR+2SWuxzKUcdUlOCH2KpxUN2Zd88YqsUW74IrDpOyGOCeU3QsMbrElBVHMz95
0gOsK5JiFJDHE6SiNw413y90Cl4v94PEsW26wNEspIDc75AmfTrjD3sGIgrGPC0n
q87DGZp34IdYmm8P47rbm03kWgl39ZjUKswZp7Zw9/dgg701wBxYiyh/vgAylcPQ
zqz8vaJXmnceaCFzZ9o2DhqNWHhYnH0SRie1dCQ958xFhd+DZcoGbciZs9kc5Qix
WId9Fg39P53+btKlkCJQx2JUpzEt9lxGB+ISThiL2fGdCorssOe4HZRqBoOUC9gD
kWbkFDTDCVV4QX2uLVZcjvea/2Rss+Jff4n5n0FaaFin8/oQs2XTFXNtu8m2a9O6
NNUJc41xbsL6NWlK+txnu164T52tTBfyQ/rRzAFNBtX/VSnwxthtDSN6hNrUfwTi
rGWobdyLxPnbiS0+qEk0oA/Eu1givvehsDJdUKbNHPgGulAjSGmJq2z7TzaFyNNm
zdmTuB1h1STcBKNFYAf3Ma1gQl4Q215vpllvfMx1+236zTCwSvKAk3pp24bqKk1g
mAWJDR5a3WKkrLFxrPidwLnzmdBT7jZuIXnIiyyg7/l/IqyxiLbhQ21IZarzLT18
GTFD3e/tJ+uRBbEqG59AujmsvX8Vjfmj0OVlmMw7EeciC5o17MKcsPzGwcS7tMu/
AFk0f1eeUcRDMfjs4iKMphtG8QuLA+V1W/jxSBMK+Qw7Lo5nFRBcsP79nUiGQKcM
Aw+RSVqtVxz+qlus33ReTX3Nwecthv1K+DNrw5rx4biP5BdrtsbVbpGRWFu/GOCW
gev1l8yrqlynvKFeSCX48JUtl2wVU3DRy+PZ8oe7trBj2bVvIJzZubYtdmB/Pn9G
J6A2/i+ytdPGetvPbh0WW92uV/Zty2DN6NRMLcyO2Ha+gSX6qojKo5OTQD7cXZZ7
EYpcB1ClhFLZ4OwiJrjkLECjueEJwcfABk2chlMdkNQtDK6+L/4CVPeE1cPNjh12
D4WP4QetLcCCNSRCy3zflck2aqo2gGOSk/4mjYlKiHVnGt5+RyTgjWS9JpPSz7OL
0nQ5GjxdQRF71RTYNZxHJDkTnNET4dq/HaVMqIDN22Qnawt5DR/gwq+Wz2MZyAfx
jVsg1PeToHjmr0YJPBJ9kMHwNOE9O3tTzH3iogjb8uW0GNDMoR2uVUaUxLBqCqFg
Sz42fhqj+9E1pcbQyKB7CnA1E3ZQFnoDrmH4L1JKS/aNGO5hEsXzprOloZMmyTb8
1QcWA8w4hYPsOrpgA23B/L0rXQ6qEaDnUC3vDiaSPJ/ZTa4v8lvse+8e9XtpaDtI
WMTVfQX/ST3rLxDUI2hsvX0qSIvty3OBLrO0ogmfnjRhvbwDLSn2r7/bzY3qB1lA
gBypwWkS12IrRthfHRUznLDHLXFhv4ypATb8FzWRUiLdCPwMmXRAT3wXFKskuCt4
0kJc2vjj8CapGs/sTpEF12d+d3x5WuFb9uJYcKkYR2asD58kvarFTqg66MS4ZS+2
P+DQBKhzF0xCkZSr6ZYGMUf3fN9+JmRHXUsVO4c1vPKH6XO4uk2Tsq9L2Nukc3qg
DBgafvvtR1b0aJnK4zxr+UPDtA7Gcmg1PsVJXTPFlRDs6aC7lxwPW7myt/LNgD7U
oKGTqXmdCxdbVUy3OQKU+Jyb+fCLa7h0UllaA0X1xgf4VNemIlvp6xPhzu2FSvnA
FuMDeiPmPBm1b/2ev6KiVjamXedrsY9UP3eSlhRIzM67Z+l0Zemv5Sy7RuBqXdkJ
fUngVFwjFMkhzzcyI8avfJfnKQH0BbN4Ih6BaeCA9Y3Fuplw4qOaF6FnEhDb3rGN
A4BdPOId9DcVnENY2xvkYAYKbc2CdX/hcsddlWKVe6ZyWsABROhFGHvSS8yuiAKh
1f+x4bU1OOTVRnjC3vhB3/XvqnQakZqosf/isZlmUMcdjcw1UKbGL3dK4LAY6ckH
`protect END_PROTECTED
