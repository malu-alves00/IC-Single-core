`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2gVYO2lz1AKc7lTjph9+Q+hYFpM1VExnwICFY9bH7aS0v2KB7ROxM0x6lXIBzVmD
EeQ908XJAGsib0hBC5VDcX12TgNV8+1bbysP3Bn6eqg6pn1T2JtQGsrpvxefefRp
+h/AnXA/uCqKM+Hrn7JxgCnqBH/dWI/ExBvgwA9YXlE9HOnQ40IQTXEygR9s+Ckt
m+ghyvuxjrwYGhi4C+03FRNy5fu9dlRRfmbFtb9++MMv9nEg9uIJ7rXyqiosyHWG
raSLchaFofh8ciCyMLgqe8rC2e3qEjcmRhv7g1nD7rtEZHXMt5CTNmEgsN0eFGNL
Jc76XFMDGJ/6rA50VXGaK2MjmVKv2eIcMy1ugnguvLEYfalF+ZBz/qozYxPvS6jm
TRom/AnK+UsyZNTLPINEk91oMM8qg7SLR6Ip3qoK92ktBOKgEPoNS02LgTpjcRRR
MVndMYoKJ/xHoux3qXGdJvI0+FGCnEEeX0Bs+NBKQyli8b2swg+elceB4QLkP1xu
oghYVvu9HD1KwwdaE2ztZBG7/iZ2sv/Q1kWKd9IKtgxwPEZ8gKVTVqb04GoaGjCT
8WNAEKqXfr4rIlfvOWAcJx1QKzwWe1eIEHqRiU57lS69MqLygslF0/hp1bkDMktx
QtXMeArktRVVfcYFSlVGvsKqfPraUrATZoLk1oW21tJ9HbdLmIDSuR/eXYeM22uK
XTDPqid6msoxhPhWohU7wBkXX8u2T3aVhcgx9Y7Upp/ei2nz0oqhGe8eAkJEaq2b
4H+V0+Z3iSVilTGgLT3DAS6+2TJttm35/mJ3elUa0SV7Jw1Zf1jvHoQOxZTkTSFv
HO1xc6LvyMy5OnX8ZjFvwFU0GzFusyuKOSfygzBZKbfpk3h4C/lzSxwkqjYrUhh4
I6B8SfKV/No+Dg4RgwbU1Flw32cY8iy7bavfJ4nb83+2B1fhdEoYMnKkfIK8mCcg
FDullQVCE7o1ImZHKxop3MtLE+sOZdaeUiZf4u+lhxb0ud/TNMayiDFxexMEX4wT
jgc3uVvvnvWXIurPEdUQuT7cH3KKwNM3fgdKd91FVWCX7b7ICWt+E5P4ZggNzQVD
P3EYI1aRZNJzKJ5jLw6WGYiuDdhiEX7bvB6yGoTKanzGlhtJKUjim/KV9xDMyBtp
ZvNYD69F9p4h5z/w/lmj+TcqdoVrHHOb8+j/rC0UgxlrDukzyOc3gvEO7N5ypbUH
DG+LAiTfXBDUYDULj10m9diMJcn97M8V3gbq7VDacv5sUdj2kdueR4XeVSUxsmz9
NtIlG3fo0Few7gBseC6hvAiP1Nseci/qvSGOJ8VFHmZFSDQ8CmlYNbC/aArA5d9f
BaltJOGkSJRz8CZ89b962b7yHxUSiidVYni8rjYgGH8qN4BrPKSYZffSl/BVU5R2
gJKUqoG/06lLhV58ETftd37rHcqAwcwLAASQPu1RovU1FhssuToGDk1TthEahcZf
aS1O8ZsKc5idPnUAlwYSm80Ny493AfNF+D6F1Agd3vkcLQIyJA19DdlLQcC0GANl
Y2qQReASIB3K6YO5MzyvbjJT+GTfnDVaBG9tPPRBWYyirC1C/CBwXbB9NioUrun5
aYaTqAlLrbidO/AbXkZ+JjlgbuSD32xik8ttxSmcN9TO8bAQasAXFxuiVLJpQts4
4xD32X3PVBcR2kpwjDG0qfUPG7P+Y3cr7TlCMSs7rUk0LGrzkqpIPqPXI7n0dLTZ
nyWzrEVuZXzUL1B2p7tm4FNRYnmScEW6+oLb0a7b2pt5ouzT3Z5B4uvg2IBT8YAY
nnlVkMVT7d/4+xxgprqHtaRpFiK+IKkROkcDua6XjLMTidoCG/VSPtX1tKvhOA9F
ZMPYNNULc6CzNU55/QQhLwb3fzJofG7ipGpMYoDSQESKTYtf0hOTjmSqEGRJZKPF
rnKU7Wlntu6jcUGkLufOp5K7RxZdtffwjR+pZps6L+vOIF28X+6oF00mag2g/OHQ
+T8TetdzRgoAcWxcYj4iU27Y9RFwx0SAuMD57tbHuKi4Z+Vyct1955hW5sueAXZ6
JMn5QrbI3ru3bqlQULRGORijRHkEF1HiRICJLgNOTk5o+Dd0Gp3ebuVvNIL1fGd0
650r3yrTqsoso//h8nsYWpnFudL4BaS2JA9/i0bpN1/ul9yjdn/4URFT2CVZQuIK
bPDq5ElLXkQIIv792lrKVdIvSwAhuNKOYrZQlOHPWJKHNxgJPeA+stV1TjeSRVq4
R8zyqsaaAivoXtL28uZKIWR7CrjVl90i3X9NB9GOynYDqwERZPVgC7GUQytxYEzX
wX5P8XlQ6FLw5yBTxdph6Lyb7RbvxjDgzVDDHpCcnpBHU41NEpZFuo0rgK2zVE4p
1IXSpme9cDdNw55+KAyMlVTKatVB8dyCe9Cvhv3KrFcQcFnQ58K6wrmwSmJCKY+x
3SyNwGLD92Qiz7YBaorWdySSikxRvMUdZPKsL9GTEJB2YHYcCN1pKpHDf0DUijby
rvKroyrj7b6Fcn4t5fQIL146f6MdeXlrPpPUNJau99YUPBkePUV2BXUpCmDFvzj/
Ykf3NwdnzcCWUFV1g1WyfehfMGoV5e/EFz4YNPDK+w+Kvlzo3lTh/+c7levAnepP
O3QgQhlkXHZ8t79xu9QNrnepcthJaBz8bIvZgBdpjrJIirVtnBZE8Imhr5I9s+Dx
aqY7BbZeGNQTOPcDoG+iDTc+jQpzk1OspgZBWL6PnnSuvCNCMrLQsjTHvh6Ne6rU
q8C7KxAC9ih+ZIby2u4kJxDhpqepFYZUFMiW4t/vSXilD8Atq4O4/zRTf4D+Gld9
gbRBqnJ5gTSnjkE5tvPEHVRYy5+x3Zd5p+zf7MoE9/s4aN6pLcHMXcarZd6BR1Ip
oL4BJdid9BMwqtr/cyICM93/Y0JPxtvtTuWeoZttHGdHQh5ZNqqq8e3ciXPvtGIY
vKRixt51PC5Q1wN7QEZs/Kmr/B4+fmU715QE4EEOfJolzjVyXyxXMGRJFEUorvlr
zhDqfyCoVijSWebwaFpOzNp3IdEfeCG5gjb/nqCrlFtPmviP0lDQIsu+tJO7w9rQ
tVuOnwDciycJ6EqB00kM2A==
`protect END_PROTECTED
