`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sfwnkcmZLs+hKSNYHiiGzJPNSg69XYYPp+SsTh2OdJXeildEiVgrXSpXwXZV0WEc
KEO0oR7H3DXA11uq20ENESKxyMfPO7pJvHoG08KGd4dxeDmGO78tiWGcRqzEba7Q
dN+SjZHiX3NTNwrngPdw2aWxT3T0S6zjUjAXIRv1l4RSkOUKfH3c7/fHOoL7FWsw
bRFKiKOeP5vvD2OASewzulqXShTMPjlGRh8v3jefcjDbn391/56Wm087TPisnVs+
i5rhtddZmo9zcLrMR4Y/ehWdWyRAgUTN4E7TpMstUN9uukRaV2O+PGiIM+O9UPqB
5ymYKpLnrEpcwCX3I/5b8Nom1Sb2JZxEKWgUtEnPDc4s7ASMf6XLmHPKOJoN0NYj
`protect END_PROTECTED
