`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kC0f0zat5f8L5xCLtu0UXnGhyoJsd4VSk0tnNauUMBBhLuTLVfUHA9zbaprum80z
vPGNQGLhoagz97ShrVImv89Hb15nS3Ut5Nqnpxp4fW10wgjOdqLIerinczBnZ9pm
NV0wxhuCM4wlQDnPq/UR6tSOHLvrRR/XaULl3Cc5f5+768Wzh5evV/qrVZy2IX47
KRN3eMPbuAp/FQKYkik3SvzEzFpqeakCEJQP/LxtmiQnOXMB5eV5IFMB+tet0Hxe
FVcZYpgG92eoBksCTge+lAKXfXAtEQWCIC9h2oARG5bZH5kRw7Dpjfd2uur7MuO0
d7oF9TF8oiN/YQ/s2/U2Y4sk2JabefVj/WkFBSGj0823lpVw02R0I6i/yOPqzzjf
EWjcQpRK6925ssKJThrDcJLs+1MosDAuPDFXsdU8JQbqiwBkJ8iNuyhKRgRTwBgI
kn5E5iRJf9sm63NccBcCRW2rKqCUn8T2gtQ4gOYitefzjCWRKLICaa1YbpY9VyFy
kWqW6p1uugobqu4yud1lGYRC7uO7F/fb7gCFWbrFBSchSo1xikyiVafx1eds+CcU
dPuSYBnXEFNpwKfc2hp1FKNiqikQT4GtkeREWfKFd7ICmBsDXyN+dpkyMzJjxra1
Op9wB2LkT8IdHY4K5xpkNqre/DBrGZUiE8v0U/IqResBcz5O/+YgmOK02s0ACFf1
ZWQ77qgf8WkVBt/RGR2tvSCOozvqPCUDEsfMHTVjhbOVi8sL/oX8FRinKz6v0j1J
f2lKHpoA5dPY8n5W+Dehf/TYyItcqmkRG0v8/sWNmDAvgi36XDki6dgSxM3urMkk
qzpoFUrWmoFlBQfQ/HC61czDz/l4oyADxHyHm0V0kBgkyLPLsyxk+X5x0i2BaWGm
IeX4/VpZLrx0/8luJeK+jzdM5FSe60lEW9V00uA5N+XPElTzt5ZZZKHBdQku7Jpv
1imDh6gNFjdQ0LlnOaSzd6wR8nS0sx0zQfQQoeiiEKllZcmG3Tz491jE4pIWLiP1
GoHbHqP4IK69sfQ6IzimAbuiZRrub9nbiOzwhavvoUXjzbp8XFP2AZ1v8k9lJK6I
0nFdQ+Rlghrw/sH7bpUJroTlF+dJtmj984ChnOQ6BVf+xsYwMPRVZez06gsqm2SU
p+yTpOb6SqEB1dNqYUTx5oVRKmJN+nsnb7DLKC59H3RIXArvPluDeVztszY4vwif
JAfP1HD8+CnaMykUw78RTiyCW1aaSVjsCMnKa3ire1TPB7hGinDTESIVjWK+DTps
5jdSez2dBHJwm+e8HyKkI/1ZsXDwncXJD62nYkseJkQ/p9y4iZ2Nnyb92XuEkfUT
ZOXUHaK2niPbGBPGlXJszxp5NlcwhgxRIhGdcOuK1foQ9u34zSHuIS/K4jhpdFKv
schVYpNqyYJZvtax93J9dxnHsA9zh2B7z5NwwqfE0NZQioHTtvolZFykfguZEGmD
2NubIXJc4dDwl+pN9jEhbhMHqamQILyvzWpeGXCKg3Tw89Ius4ZA+7f55FhSgAe8
PKWSFNJL838tBbSvvn/GrTW2vd2WVTs9/JhI0IcH8fvy2BB+rSqSbkdvvY34H8sh
4n4xjhqVTgssD5HpSCkVvm6ytwc4CP+/8R4MzErcA+DXj19DEfnneKMQa7heSLwo
IsJJ8tf8DkBL4DsuIfxUkPj7agxJEwIutiFSVdp9cbp1Q21e41/ECNcHQ9xVuiPd
ByVUdW0MLbzPBVRbrlIs1RolPv84HrWLVw7lPa2fB3+809eMyyLClTeybQPiJRgw
Xp2h1SgEHpp3RA+9fLTZd6whca4Nu0NqWa44Edt0V4Y7LVzlwtHeXScVSqgs5Nv0
pKXo6qUE96Mnji8M+SkzDqZlu7UFCiXZbneOD8G/NaaDMXeJl5s09QasptuvezLS
v5VV3oTgh82yDQ6wIy6AAaSJMCWQTsfKFSOtC9wrizkm1JKloCcYaIJpmJNVi/Jg
vpQ9sH9RMPU0+nd1M6PD1cCGRcrSKABhJ7UsxJRo7cwL1hDTSOk9YIiocR+bNHNf
vKOY4L5/PD60zlc7ZQ9WafUcgpK5x0pyDmhRpUbssDndjmwpKic5YTd2zZ9XWyvy
ksxLYfMvzopOfQK+XC+yZypPRk9U1GivnHdgpYDQslv+9sfg1VUMQd4+0CjVwk99
JQh7L7+e7nQDg8HzObLhdsGo2uQHc49Eqo/zCUFbcllVA89mzbTzs+uNPOHIK1En
w0CxGCzkmBeEkdlHQn82TxEEIRlELKt+tKFTX8FL1rZ8M3VPOwAPWQLq73el5eSY
NGYYD4+A8lLjVUITPOe3kkVy7IgICMoQyeowNIXD+F9yBnZ2/yExeZJ1eBPPmYJ0
/9kfy4GfxMTZXsQf3oKy+VZeiTxnq+kEj+v1fZy9X9rUvJnF4I+f5uTMJZJ9B6tB
KeeOxSt+hIKbaNAXe5Y+XkDBJEXLzTUSRuZeNh7C8AQyzXJHwwQhF2QSwHQAaWp5
igYmTznuEzueCSPQNs7nu0ugd7ZTIMLKc0prlK40DGxxlntI/wR34xQCq73lIvJq
n8HI8S2euQmbIoD8CTEIC9BwhpTdCurNTzpcBBT2rgCrxbhUbanHV1Uv0P4ny1ut
8HgiGL6C4ThzLijh73Y6OjUQdx8vOKgKeLU6/lJs0fsLuB4P9ozl7EGhaxs/k57g
LTrqLMWLneWr0fkQ+AbwQJLDNk3FYteAWLnL19u3JBhrAsQl0I77vuOdRh6+vbrB
aapsDUw0/FoqDuhLrNdz8W/rEZm3Y7F238itLrE920plffTAqIqx5l9BDTj3+kc1
WC5dFuA9NOOCNJPELcIlz6wSaZOswkYB7EkOLoO4JD5XhxHis69zHfdCP7E4/yvw
CnQhTBHd7P1rxJLS+X4lumDCDY4pk9LoBE7dh9aHUjrov4UCqeBrSsss9lsST9GY
CQmjVyw/3+wsaWUaSszKPZupnPthYmfzLO2DcoDa0F02Dk9DuiU8Wf7EDV02oRvb
`protect END_PROTECTED
