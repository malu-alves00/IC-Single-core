`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SUQPAbQwuH+/Xm7W+Ndh4D+r2ybIv8jEFskqfCSik1nL3x5w8PUohMIR0sWm7JCw
4dnHrxxsWSX2Amr+wOP3sMqXNOeQk8qj/BZ0i+n5tJ4HE4gOwU7EhNUpmpvogc2F
mcYTQqJrInwgRg1Y4z9zIaSq8y41PN92zcD0CajIKjXNdUzsVd8OT2k+r/sBRAtt
5w2RDAfnOMCyDwfHjJFblne/CDsHesUKTSI4nN449ISsWlVw5oSeEYVFM2XfUCjx
hUPL5zPA7OHI8/KyhQI5I8XbhEO1hmYQcCBXYkQJvn883afoK6Btku/cqzMfVOxR
ojyFCl3ZWKWjCiz3/9hLrQuWQ8WJZEncYYhEWK+vlUl/vrkE+wZLKddycHWQZk7z
s3A9CU7hHYYQsZ7VcxFVW1q1EV3/RLe5NftoUqCkkXc4TGS0yrpQ78I36/2vWEta
J8V9VDucYG6xI/8Cz8Oz4gO1PNhrgLTrmnVEXZgA6FUP8bo5B6VglwjnzouluBIK
sLUktNJCOLwe9OixAvDEpFVwGOkXhcm162Bitzbvb2zlfNfv7JS4tV8YA83cJgdC
S9pOR89LyLk+d18m5hUuZrncTDqLbBbpIhrzX4X6p5hu+CND1zp6rLC20CI6Xepr
9PmBziF7vEg3cZnlgaTK77/h5gdMZnZN11nLnN6j2LA92qXp8wA49KNVDmkJeG2F
iKNXpl/5eIcnVUC3/aVrAdBHv/LorTZP8xnk8QT9j/9kZoE3Ruan4KP6aFMg9egB
7Iv2T5mM4W6pYULeXssUvBB6rqjJ6qE7tZ54AKQSl6espWZtjv85cvWMJdZvJKXo
voa7HiLgWaFwlgn6gyVjzBJbSxSlsupgCvNftbsarqbWC7knd+uvUwAY8ZMJ4Rng
oD+Cg378K8Pa3llIWS2Ag4wT4ps/GZDJYPSugTy8qOmIJ8HVE1BnT2o7OBb6q81E
KWhji+cXLg2c9JAhMHkfe2SebRCTZ/pTVvQ9jKbVpjRv4DHEyZW2UnWypYDbSFFZ
nxD5M9aHeIeLfySr7em22cCrUs8aLlDoACKmW7+DuyX2uzrQmh4/+jnlBwTKVX7A
wzA29QPkGnX63U4MhdiCmtzMN22xltLVZPFpgtOtCNh5kbrwiuanW2ecGbM1jWql
L/uFZxJ3AO3yIL1mqwB4+G8Kcu+fMZG0kVl3Ois9QurmG2yyljLJeTnJ6yjAzmpE
5Fj+GTWzpMoEWFjd3QNujBCB1QkjjC0OpNzT+AS9/QEqKkti7tUd41rRdlSyt4wR
4M/l5OfwYjz+agd7IYSkDK8uCCyDMSZ31FbZQ225zJraPdYosSy+m9EHyI/Xe+n9
hDr+nzUkmcA0PJq2740VoIlJ0VZgAc7SaWEr/+oFZZdXOX2dLQ4EQywHhisA/r0a
aV5wXNLZbda+gHgB4HgubZpyDfiefep+T3FgAIS5OReU0Pp2CT6Y90ZUygxW/7JK
xYPrr+4OnMGQAk2wEcjYadLhv39QQUtaDnELfO8558a7GTPixZ0gOhBsXNNeiN0h
zF9jHruNMTMaGm3AmCHKuYxknK76tentAEDQX/EybIqhPdCnxMIzJ/3U4Yv/Svfe
gS60ddmeAYV+EIcJlws67aeaDTdU96dKwFTpu+lBufCKz8j08IFXaTBv0r8opAl6
B1m9Vu5usEsRjMB1HejmHziZmyvrKkQTcAxhIAKO/DKlfLCeCwjRBPUYRNmefqrX
T2Xy6GSON8xoPioZGSg4jfSSLbZCCocjVBXi9peczNcp2xkFJB1+SIzhUCAEDP6w
qvXiuqKaa7OaJhpQ/TrvhSb1PrO0m0i2gldgA8MyxAptBipNcauVk4n2OsXiCg8b
CJkCCz703u2qfnNjb9VAdVUwLnM4IP/hXm85VHYN/5ACcvxDVbungp3+D4q4755h
selCRqwu2hkXPR954zEutg1XZ8c3Sr2vmm20Ptolm/lx7M5PMKPdIKz03sYoP5a7
RmUYbkeUQb95Vs9c6dv8ETqephstCH/LsIL9BLZzsab2+/VMzlv5aPTSzvh+ZnZt
AnhC0Lo4GagXn2dHMjvioFdgC1jV0Kf8w8a0Tv3ulij1gIszT1lhfWnxw2WukOe8
2MLiByz31jtqbA4/cBIIMDkBYcixeV4GavIdAaioie+sEH8d1lQ8HF58QARjz5Kc
Fa5HMlHueDFWzqnMpq+O3MT7ZVslSsIuglYtAOHLSr2/30ZCTJ5IzcKmG5a6mlvH
6ewMLYp+09JCUfjHiR0uktrEAYX95WZBR7lQXK6kyimN41efg38dpZLjEyQb/ewp
UscKm6KopBSK1EX0OZP9hUsXKsgXMc+Zm8fP2qQuGAYcZpPWoMCUutUWzgjFp1zV
+0up0MD4jUSXtbxdlNqYRYf1xLzYeiqM4FQCQ/MqKW4NyLxptUxT6czD3ucSVPSx
ZxC0GoG6ZiKhdLawfjktvHvj5HajTr6WM6ep9axaEDKCL4w4mVbuOxgiuTwx8f13
R2gQX7WjN6lTPMkj5bddbbBLelNYVbmkOf56rKfDkaHcrwBoiYWJWf2bXNAoukLc
SVkNn4BTJmb5vUUIho4zlr47Hekn6ekMCmoaT6PcJpE85lFypPx+LeuCraFiAYj/
MBKCQinwj5ftw91HSvnPVt+EwqO23S/c6dTxFUF3bjAq3VTjOhL6k+3qw2hzEvff
QYLFQty9UQamRrCTrftL2Q5KTlb8bco356RQ1cLf5icRXH97QkYmLHadOBPtczW/
fZ2fmCqX9kQQCZmAB0gLbJP6jxY03YIDE3M3Qx+0SVgCMtmI3yE3JrFGrpUX26jV
fhsXUKp+AZzm1QPWc+yo2Rp/dxLEX0mFBz7HxHhKwLFBeJMFXMvTDZmrBfhuRkFI
J25I60tCmefMP5nmAYM0wr6d1K1W5YaxCLCgdlBanCZE2cjPbXCHmoGIIonIVIe6
OxSrsP7pupgStYhAwQlMKh391CLASeo/ljo2OyvFNXxbn/Gi8Zf8c0bf/Y59rOYU
DARlEk+rQiDvQEgM/JzOAXGLcuIANVZ7qRsVOGX0Oef03sjaP8lAEWWEj0x4rKzj
4maXn8r+SvQYS/IFMwd342+WGERVlHt8thOW6RW2E0zIuyrrsEsShmssaBwVRjOS
kkoa1LYn2oIWUqdalALAK5oxzW13pyi/zUauUmrjpLgW561iIw45jQuUzHDh4y/Y
p1VAqCFB+2EU0HrSFq9AEE+rq4Nhus8JfrlZMVT3SSBC7jjB/cz73y+nwUFYti/E
l/1lb2G3/drP9pm/5eRH4ZtKvYgbhpzpon2dG4XHARPQBCfHEXAfeHSFR2bfzmP6
lFrbvW3Jl722wfWPUCiE9NzWAX+H9aaNJNZt0eXcL9GAWWfsJ0aPnoL8AaGIIt5P
snCo15pUfKDL2tN13RKzJ/bQHLAzInRy8LzkIEfgb6UinF1j3/RFFRRtMFbsClQE
4FqRLKnDIFxAx/0iOH/0YMBf2X6ZJzYn8v2D6Jy95U07+6PCxvWsNuRp24tR8DGZ
Kkh4IzraThj5zG6/7MfQ0WU+kxcGX8p9Zc2/JteFWYBhSPxSz34YT71mEGQ4CLMT
16dqtV0pHNvqjL6A7+qjD10vuFMmLDqtnt3aUxlJDxtCoggnE0iOEzGhyIupK7Bo
BOE21+ZgcIHR9ohL1NM8v3MlZ8fPUJgREfSbkNDGoiJzKeXJ+YKCV/vuHz+7zA+J
O7SlvtEoll4HjOd7iAW0xM7s6HkHdrs9FYhlD7ZMfZI9sYinx1SQkmIZcRpKz58J
Pbwb6i4Ixvjb5N9sAS7m7g==
`protect END_PROTECTED
