`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lw7V5GMEJP69jYImNXpJc/jxJAMZiigPmIpLMt9cZavSiSdq4RswpjGtl/zriSA1
OQtc9U5FIbU3oobBdcIPo+J0dN19c7tZFD+uI/YggoSXDaMIxis/Pot2e/TDpLOz
GQFBQSAKuxt6IlxAR+N3VI+MPhoJrnM7ZTja8xaew1l18sfnyh8pz0mBfX92YhjQ
mfAmm6vukI7rnE8xewoI1725gRdG84h+ApONdwMrCQYObxUno9QBJXXk/GnS6E7G
ZXuDOROAhBcNIz1bpsvVpCP4xneev8LY/wcXew558kntiW4s5u35riYnAwxdvGvK
5iD/BT/1JXckuzDP8elFFbr10H1tK7jLT8QwCrWgXFiZRy2zUB33jencBrl3Rpma
fMkfzoAoJFkvPv2DoasGoE5D2ImV1RYCGUZzEqP0loJLUd7kW7y/3LSCfXTtUzfr
ynBChrMjLyhiFNEvgqECvowqiLIqzH+1dnhh5HJYB7DQ1tEFaDg1t46O+lBiO08g
VjeBypK0c3isYyWQNPfa1yTI7QL07Y8oB/0XknG38zXJboPn8rypcJuiiNF3xBHW
Q3KS02CANJtOiAXdQxgWUoF/DZFiUTRjRKw1lGL1alVv6fJGtdsBOT+lyOUP2qHd
1dbm9LgJmMwpecAZxqLnA6ry6fUP3qdeZxyE47DEmvbdctgex5WGIakSob4wnQSG
1H4HSIbyNpX6vdFyx4ZKh+ly8jr8U1FdSCfEORDbAfFNmGw5xFbBicN/aX+ysIkB
eMFxGiah/kvv1yWMZGWgp3Mc5vdvOTS7Cd18uHR7qq+hdsV9ssoSVQT5kW4uSQcK
/nlO4c/Bu7lTw1MDYcsWi6haFKkbLeyoQ2tOzk9jemOFfuxCivxuUQvF/PzVRHUr
gVg+VmNGdulnOrc0AI9O3qqXMWRsUwyJzMjqKlaYWqVqN7azDKob+U2juGvCKegl
UsRBERUPaIFZDbXooyQEWkQaHYHr8CMVduXpiHltv5x789mrqiz4mLhAWpMKRVRi
Ofny1R7dnoA7F5OKl6BcH4QneOK9MNZpZ5QyHoxwKXBcHaMNnlMWFZNRiKFnKZC2
z/nDeVw9yKQcKiRxsoYNTTdxOA0AGt3MIAXwB4F2K9ktz9PgjXIq4ahr/AQirlEt
`protect END_PROTECTED
