`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YCxIKV3T1G8UrsbDsDBTA5TGIOW5Tdm3apxHcx3OEcO8AqXBzOx43DvWeYPcYeo2
4egEnt1fsdHew8s0rSn3TaoE8PpCErzYFeMvXlyI2yQID67ZD0cGQhvxIWypvGMf
GxSRmVbGHuH/bEJji/EBZHPS089VWClp81cfxyF3g7luDVU+Lo2WDD98pXHlMDi+
mfxFfVrPV9hf9ves+IGAYoicCOC6VFkCu4VBgJe93kLquKoyxmrv952znPQ3wTLl
5Hj/Aw1RXHmxB7LMj6wyPx1y46K27iaiTUdgDDia6M64hDn8MLjTWL5lctp8cnv2
e14b1doYTHejwbl0dZ7FnYzFghfC9LkeI85hg/rCcc8bDv71iwjTXZQJ44wVC34A
saVrXV1vJ+2KfgsmexJDuGdGqj7Kl6bKxmCriHWJolIBpTUtEbKZl44KXYIwC7/6
flO5X2rN/klBZ63SUpjypsqiqA5e9+9F9lv7Ga/8DKfnCrrDho0ZqeKvKHUj8KJT
7dDgSP0yTOcF6vCiYU3cJle9LM11cQnYKYVLmnvG1XGpCKEN9cfOXssWLZFMzvlX
F/sGrrJWmf1/cYqIPQ450w8cmOVMZmzujO87oOHVS6s9qTupP2Y2A7AIEMU+ulic
N524ZPUjyJ7OokkUAGWAiEwo38VsK4y0KzPX4Q0xcMTR0UEfpcgTIDD5fGthYSJ1
/j49cin7WbLkyklHD0PkeOGvfcW+pboYzkUXBW0HyC4aw6XCoeBpm5Mmtqh6tLqo
tT06NJxEWZwoTYjfrxHcayDXyUPiWI6r8kAXhmBQ0V/yfFu/RahDSw2Y0AC1Bo+J
GPPKeAdPYfDEajU/npbDF4Sjoi8KkPq1FqTuAx4fbJDwetjA+v2npBePT37BwHhq
FQ2sPDb67pktC9+nfLL6fUd6pZRwFk8W1+MqhpBHHRQ=
`protect END_PROTECTED
