`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
StFpPnT6vp/zYHVFon15kQlUUk4RHkHq2pao0NkYJu0SZ6eH/9lXaIY5iYE273ZK
sZX4V7pInPJGAKGJ5KA3Cqu98xFDtx2PgEGxY4SUddtR+XsEmcuTnFper8cAiNJO
6+f69OVCOsvIH2/ucvGi+l/W7KgOD0ppdsmlL8M7Qa0wMy29tfRdXrbyOhz79dEE
qhuTVHUFEKQaPlCRSOBXDNJ0uV0+alMtVaeJE5i3TQaOOmEZ4iIp4yNKNojC/9NI
hEaNv5OJI7+8GTkVkObzzuTpO0GIwVJJHWVJ4SWgrpYCqdYReI0vC4sEjTlVrhGV
niELXq+4Z+9EI9AspuWBDES2OjtS88zVICBzoBStBmL6pXL+7vwgEJ6epoHzyJwD
ZBIkb8zz68YZExRf65qXCSLdZqv7EgaMqOYbYyoUnAxPkezr3+m14r8TJ+o4aaMd
cso74rS6fXSfb8ILBHal5hT9VvpqoxP0sAKgiGG7s7i7Fbq1WraVhPuq/J8VTTVd
Hu2irpW2KgfTaKfcE9n6YcIDt7Zz11DxsQbsakaPFYcN43M4HHCGNacEO2LVt2Ex
zeK/UmoCg37GIrXnZi+yaefHadNoONWqaJV7GQ3+m9CI6H6xpvDFUNJrdZvJIs0C
nXg/KGgZ8bsyYMPe7QT/i/FMHcY91QAiCaUgewBdIGHtSiObLhBgAW44ZN5HS+yG
D4uiaiY6WsVJx2LmdTU/bXIQzY25ES8VNOyPp38bYgyovXzYaxp5FD1St07653bS
N4OtZHbor8/rVl3vZlvmr0tYoWCXg7OC1lEt8u4Afyyav8rlXG3vQIsNYPYvZf6O
HP7z5MecttwmBAK2P3uAmKmv/vocNq6UiNLgK/XicpKAJ/igNBxPjVrZs1fJW/zw
xxvEsmr/78czaawUkRk7k59VGpemjPwlBeh649qzHyRPfNxf8++SObXdNx06kTN6
/L8toSKnIuGhWjix7y49gdV2SiX2NL+/ckGy+O3EJW52kjgdF+nvoTWNT4SnBxdQ
nNl9AScPfXEr4TBkLQiKuQr4ic83ZY70AWNp7kUJTImYHW7c7YBApkoZLoIpiNvi
gAy+Gp/BZnwTGNzwsvQSlxdOJJo0nnB0uYa6MZy06ssWKzQ4O9jb1YqJGztlHFZq
kG/rQPThNUaU8dwJI04EoNEHSuhRd+VFMD+cx4y2C6a/rGIFbK5JrCMie+lwpK51
FDfz8/vIrONqzDi80L1yNXqwBKdgMAFAHh0RRzuuB9URJBuEVbhYIg+r6MM+nnix
fBSvBU6T0tcSmfNF5OxEbnmZ0Ly76KP+gBGjnJEHv/dp9kHvYuwaG73u7Y2gmNfl
`protect END_PROTECTED
