`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UVhdWtDWdLgzmEyVHmItBxRdbN2Qgh7S92fK4IgiUWUrxNcuPA71M8fXVpg5Ud6A
3HFffRLQgCyoVy1g3AenBdVSGG+EqsjegGRUey2Rx/W7n90rox0LPMjHBJSnnHES
BjL3etTgwIG24JTMwRiNpQZVw9KJusaLen1P5fiH8GCu4dpEHhEyRuqZTWFcCOUJ
6P2V8WwICZluNSzPn2gU756qwykbw9ssorVixro5kw+ZcCBm+K2qVwva7o8P/FC1
LBPrERzGg4y6CRswyQNEV3ibYlJRxsigVf41e1eUigoOIcYEWjUc/QO8skL1ZFNv
9twI5PfU6/8oBkwNrqtbSmhwJOw/qO8PEBI9pimPrrJkgPaNbetI5Bg2A2BqBbLX
68zOTJGzc/lBcPFLbkiz2w==
`protect END_PROTECTED
