`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+uZzxb1huregME0xB/yOeZ/86Q3mApfqZS7F+UYIT8UFkYeepM9eEO2VZv5iWVOl
4AvbJd7OAumvfFfaASnfPUBY2JsjtXIjOSRlulJdrwMh4emZONQH+izfV7iLeNFv
zwTqEiqnv8RnSbG8/d24vD9mCVnyrVhgcA4XuS/Qu5vSf1O2xLku+RupPM8Fxq5y
e3IHq756isO3CujXtxWEU8urcoIfsAimNdcMNdUFi+n5Ir2UE9HBRuiPUWyjZPmi
97jkaSSaVtQEhzx/mrboQap4Cucs5skozh0pWGSFQiC6dAKJQw04SuNDdCq7bQU/
QSGH5W72tZ9bZv+z5gbtmhQajvpzg0ibK2gZ5MyA7Iq+eeY9/TsdetsA1bnPC++9
Ru21BduoojDzZRV3w2Xa0Q==
`protect END_PROTECTED
