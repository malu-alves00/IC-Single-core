`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DWfSqmZxgM4RHYF20F0Ri1SGcEoBMF/S36LdzTZ4ZKS1ZJYaJ07d5x7theqkzLB5
hIuzFT0vSB8E+hMHH/oDsW2iAYbhHsznTPt3uS9Xc2By6bAvVLUg3hbEKbK/wbFF
FEQIhNh2fQphANXvGkXtv0zqGQSuAU16rzquGyy5T5OxURByv80NCDucKWEdw+XC
AP5c5Yza6FAPaEico+MaxmkiMlkxRHqV0mpgXDNAIbTqSN0oVPbQGkOnZwJ8XOBm
o1H0rrrYGc5sxPT+GbcFSf98JSmYvPGNCYnj2hee62MsFpCRHpu4B+MWGhIFX5ij
k7wDyZppTxHbH84znNdOCW055Qwh+rAITYx7f1GPeExKhXjrbWzIHf5M+qMSLHF/
8DwvxX5jw9mfsIunUxLcLaYwKk0SUP0HKkzpfFM+CVEiJTVmpgd1226a8TJRW1+R
j0kIQXBxSzLxYuRT3xHMIaTt06AwWPii1xYxOO3oQwQw5SGSxUC5hnMKpZsVSiAB
buDbU8dNFeJopQVrGoNlX5L8zUDILVG8jZB1vmsDVpcqnp2w1ZYe57HENTYci5ka
3dR/G/7F7SMUICOWYNRkQSJhTtMaxBHbPzJ2AFNbLVE0UgiXvTZZ2ZkxsnuCEX9F
GnkaOgiCECM04H1M4iSqvl6bdWNcUFeE9R3VofvpjuUmlvMDSLWx5tHpobeOXXsv
grEmfJiybD0Y2/WO7x9iJxh47DOIoPI62dvpcw/BPvMEOCoxD6+teU57C7qe/rvW
/RFw9p30GsjDTtE17KVWPk4R9MKwTD0df0La1JCT8i/jEcwBzR5PRdje9YELY8xk
bkTS0eyvrCabe8amXtSq9X0Dpke22hFd8TA4KZF9qgLjPWvPTaaQrwXcl/xSfNRW
yqR0Y5haTwAFUXEzYr4erivubdWKI8Tk9uypCoM6Yms=
`protect END_PROTECTED
