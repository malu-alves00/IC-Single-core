`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9wv6Kbn9G1Ozbvysu6jgwi4G/FYry3o1Esloi5AL4F3B7OBhOHBNqGZzfC6FM6fu
fo7Cr69Uji0l0z5vjTY+OMuEKAA9m/ZK27J5D/MvNkLSvkNYpdMlQQIX5X+tHuFT
6956yXw5WPR9YMJxxstF59y2zXQHfybrc+FLOLFMpfH2Xnyy+beOtVPTY+E/phrY
Fd3qOhbes8MCR/Q6/A4X9zrsWzJQR+s3JHW3ap84Z3ttZobpkqG3Oe5VHYA7Iyy3
nRldyISTMqabkVCkS/I5yUZObsdEo32WDuLFtPlvltwdfStuZRgRC9GOa6mB1CkA
msvWhssgeLS0ra+Ps1oGqRhJbgBUKNujrgzGwnuvZA154pn5VWFm42qLfr1Z6gwa
A98SHDVyLHg1WaOLnwRihqayDt13ipVl7bHmemo/CaMZgZUZjP+uv7kQP1uP9ikS
r+Lo9uBfR4opHq2rs4gXEjKdcjGdjUzt15m4i40jMiHbl8TtHo2qRQhvLk/PYTzf
vwaX+e1Pd1PwihNcbpUIJ7mLotABAH3rcWD2f40sXowspTAeTfxAZJPA0fcrg0P6
SrYQEqTuMeL8J0R2PXjIN5ifOWDt/7rf3OT5pECKcSwECvqaWPPCVg1KAk7iQw6Y
/hNJzNDwlPaiWUoLj99BMZjnJGAPtALDCJ/PWqYySHFN4xSvZuqTcjlQzHeNd0tS
fB8Cq6dIHJQqjbV3CBtHdYuZu54NyawOV56OvLtDPkTT1yi7SQW7Iyol9bBOwKvG
OQj7pq79pGmQZz6dG/ya34m8viGZ4D5MMLdxh8FUOb1M1x1y9J9ni3JSF5ccb43q
eikQXfKzkmL7Rl4KvChl+0Of0/IYEfTeN9jDRWanbTRE5kBC24KJBuQPZFbqsSpS
tsGlbtCQfD6/Pb7S3LwQUGn/4N1WoZnliWurPT4VTgfjQ/13S6+ozqhZGrzOBars
z/FImG2rEF/myeym0oUwmTOvleUjRmcH4yW1ltobx+L7TBcVV7bwrTCskKJV9Yzx
imr6HigaBCNSpZcqiQIgajx8uoqU11Omkj9codsr6g3Tya4J0GBSLbbmN4wrRELO
D91hC0WZwq0fQt7cokb+Q/mWDFta5oJ1hPkkpMgs9fSmtoYpOys8I/yne37wf1ew
dbJ142aNh/y4IfLuLSjQDbwqZ4UKVfeT2uNmst4fqzglOU+PIgEThfGt1a+fsozv
cs2Rhc1tx7Flnoe/2G7Td1pRGh7JRt/dBWBeUVrKpxI=
`protect END_PROTECTED
