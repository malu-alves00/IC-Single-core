`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
luPfnprNBdWWKXj7Y98eOfCmqTH0nb5+aM74uJNtWsW+zKPQ/85R3nY3H0e79jHV
HW17MCGrHppdsztoDXtsy/YucKl1dltfnXG715W9WS4F7ddbjcLnJ6V8WGDyGU0f
m6MyW0xvZUnSbY01h9Fnf5TvcDJKA0hMsDxkA4Q0MPLjQL4qzhWVWFmjnOGWOTrv
4sZw00yFheam6h+NbP15DQ11yhPsDGi0rdEmiWnF54LnTJlzY/RljljfBXb+oh8c
wy4oLPFTjxgG7vntlg0yQu0nbTm62MWMDY8ydeZkvn7Een+689OR6fLhEh4pynb5
EjGJ1e3szNh0HoO9o/0A9b2LrItPEgxudMa/dKsnbJN5Pz+KqYHQevKERd2AZXE4
1Z5Q3e8rM+2pO6zDKBovHpUcMw8E9Mi/IhQ5Z73OnkUcwe/N331+4RXO/mMH4CE5
zg7ijI/UMXkYGzwu+1XbNQ3361u78PkoeV6YJ9J4Z+gduZcBiIpuS7DrNX44nVKs
Y87AHmvnQCYo3xTuwExG0ciub7GORwdmO/ey8mNUCGyq9SPakdA7w895/I9KsTts
fRHgEUB4NFI3yD12lCPTdH2krHa359FMD25VJy0aXBnJLvO2qJR9YoUeTB6qcKjt
PuKz5h/sxXBsJb2yYOgGr7Jj1hXEhQ74XbH6eRNh6YPstA7dULJe8pvKL8IkBKtl
321vRzXSROWrH4Ny/8xND6PudZwB6LRtHa6guqKINZdgifGfopOOT5gvHMggKtUp
o8wv0bmHUZbABr85VNa5Ho79NZqBsOh2jy6ZHZg3ggc3zbwPnn/hLfii+LhE/6eS
fw5iPCiTwMmx3u3X3vEcOMUTzOg6LujS/QPHb1K0Z2KBHpxtTss5XD64wKVBwruM
BrN+sl4exbiM2q8EDXiDl2acX49qESR+HVwl3b5y9thRm7op1SndVl0lrzHXzcWW
CB67OFEYlwsKLGg3GBg0JnB6zfm0JTScK3Cr0QeRDJQTUuFGfXepuXXip0dYQGci
qiTAnQ7wwKqrxFEu+vL/Gj+FliOuahuvcKyLFe3p07s2iK+PhLl5C3YBoCkHMmIW
8PwGgHheGjmKvQBz1cJwo91ZSp3JZzY80TjBlEZalC4ZJvh7wy7Vgu2SXz/RLz/i
HMLZwhi4ESXuR0NeMaIN+lHHA6+cWty6mkn+k0l8pqt0rIbEMX/KhPLk/dm0/BgY
eV26bTnH6ATsonW8bt6UvUbBfBQec8LBQNxLt3DEJxZjoQNUhcVeJAh5DhmaZrz+
CJtT2MV2Xu6HPW/bYNtuLMQ4Frv4wxYnFdpJ55L30vH0js84F2H1CTjPFnhPiYFE
n0t9nxGFWufRQ/3ZN7BaK0VWRft9FDkTLGUJ7oQ8IpinQrl5RFr9mE1raDXIsfP6
74iOvlmvEFKThU6x5u71K5HXuhj1KyoqvntU67h89Im3jVXWVnpvtjNKPga5ndyk
prHHZCNzYgXkO/jA4G07CXuHsHCq8dLMXmxT5+WE/SlJFoJ7gkCs6eWkcnSLcTi3
ocnw9WIfviLuz9KSYAv2OUfG9JbAAWUEWFl38MAXeQqG18vUdX2ClpxG2kSYKxsB
FYIiC4v/VoNXV81QS77EItxu3nS38AjSKupLDbJ1OgnsXzz+imyapqOguiL6AuYa
u4+f16wlAc0KryOCnqx6p77hYvgqSf3N070EzXqX7kbavwRT8qfT3dxLx/hWmGYi
BdSo+UvOWftGksnR3roBuQMjYjHFqJo0vLmlEVPaOiPT9QbzypLmssHUfgnVjE3/
fnclss6N6b3QnHkXtVJ9ia5H0mLx9hS0j5q0FUyxGwRtuvxhRTiy2wprvKlELvE+
lpsIR5191KHbtJEHF7hT1kUXYTnZiuzTrhBD8XZ1XGNIYWp6SdT5Pnb9A3HKTB2f
YWnBmjg/Mn1kvuk2PDrMKQ==
`protect END_PROTECTED
