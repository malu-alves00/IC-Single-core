`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lsAnBxBZtm7jqKczrM9Qe3+Sb1+MqqEPRL2Mr4B5uOTHj0nrW3o23i3DAWW1IY9f
8n8eQZhW6iC8DvwR2ZYPApiy924mBNTBnefDrquiihPvKujLVUAoRL+8qvH6E16H
X7UDi0peGhQx1ixjcPhcCMk0+5vSUhxM6jk1XO0lKZ5f/v3+jj4Clt/+cp+hsGQw
aZstOvmfLhQ/WzRdtdCy3sI5kCR0SJepEe0gPEiZoEd2KfJkk4dtdZNBYGb5TEct
9cnMJA6QnwtENu3fq45Z3VUvufgx+n743Fi2X0shmloa20vWp6/I7eh1vXv/qcTR
hRkT9pYMyXa6Fom5mQPzIoXQo2dzjnPlSV9t6Edw2KWhIdmVOeO1eEN0Wy+znntl
3i2jG/mAviDBANT2JvZ38Me6+2qMrn2oFxGAIljsWcwcJ830OrqmbYvVqmXyREtM
WpQ/WqbauhezcHbtOClpazfcRKnh7J0o6wsoBH0W/nvRcdy0mbTVDsX2BVwtjPYa
t+O338UHidRMkN31fDoblm7P2jeKDAl3ahNOfmKAXXmez0+Vp15XddVAvpI0jUzE
sr/begJMGqLxXyBe1qV949ylrwcxQ08oq6rYXp98SiU+Xh1ZOWEF439rK7PbdJc3
E8W7VtCbd3P/3o/zA+rdq1q7JWri6bbCZN8yWw/UEAkdBvqHrdEcUGhZt5gYuwVV
hMiC13wVnz2znE1Sx7stZE0kelRaD7ltYd7tndCA2FmtUeNufdTPJ7hmy3uBe2qL
foJTIMDCk5ijSkqdqtBNO5+2IQpJF24XrPXElq9YIk9p1/aeJa75Sruj/6WoMTVd
/yXDUHD8hnavYouAQlV43UPGImjtrmtjg2c1kjiPCZrrUwMsady5MhcoZ3o2yhQt
/cKa8VFcEO2OH863vysg2/m1E+yqlZHj4gRtlnSkeYlWdyhrNH1rO8I0VzOl1Bft
7FVs1dsE8SNl5ILcVzHiBYJpt5cIcvLMS1wU71/n3TRsW4bCy0NWzKZLESBG5ABn
CcWPYVC1rL5Jzkh1vrTLgN0ImdYVrFrBG7dD4590uyoyrcfINGkNRsP18MYskC4J
Xks26fCQ3SZGQRizdOo1+53NjVlcSrTKqdI7+dx+Cq2y2yFF7Qz2JxHPZTZFM6v9
6z1K7fN4/xeaks8TfFWCaoyADR56OTgIABtFE4pFy8o79/UAjNiKjgJqdoFY1mlt
LMYU+JhJPeb9Drg/r2cKjqZwJ++OkshKpQcyxFLC7Orf0lbA5Ddqcd6s/EFLoH8R
/g0lWN/SMLk2E7vYPMQQ+oB+1strQDNKcHi+5vd26wIX9ZWQS/SVza7cmUfSElRD
acuw22YsoBvUEPvFnuKqjYgLlQWAN4m18OX1/k+2OOV8K4Gm9vsifRzKGwMKs7Rj
WNHphVFPmtyUsyDEXwYQeZCjfr33qlTdLJE6taxgLdfHfENT8EIrSq5ilTxfIFcW
A2dJNpGJNURjUcl1U9YI6njyp3dc78j/EgRP9SaJSvM9jhmfRItWZDmyoKHw+T1q
PmOASnN4FFQvG3OKvV3/rSI3bHCC1z0fX9Zf53xMLjy7NUi+3+V9P+M34BHrA+wi
mF9636bqBpe9JH2WY4igbi4o2rzBShka4+9T1r08LSX6w9Jp8AUzaANrmV0eolE5
5s3z9gK+/a1RD17/fohhPpT3Eg8WkD+IdjtgoEicoC37FPXNHTYo1dS+HEbwPDBM
tJt6Oc9bWXiehSD9Gw4r15i4qkP3KvsWK0GkzEPvlJedM/RwcZhJ1yqmEr1h+E66
/CcQV/osBv8f1ymrkua056zP77ORLYKDkmkomyV3V7RmOdGMDOmpJi3HeLkdoAB8
oHAQD2Z3MxxrpfsnZrokw/GtL6wR6ud1JHntZgn+OXcgkeDSUfbBtHND5kHNopEz
zyON9YzzgOZodiRo64NZm4sCs0oqoVSUOZNZIydErd4H9tM30alZo69DKbSWc6/M
3E0VZ5HG5yoFLNBg6fQGOUUwH46qvZRK60rTBoVxGCv3zAPdAgEz0HcARIWrl9dq
CpJCl9d1zfyiBo+6xRCeNzSx22qgV9OCDfnCYmbSpvgM3rdab17XWSEGfygsHbVp
J/IliBbr49NKiSCt8dER78LzkGtaTPJ7MnsmXuUkj2nWF2Q0I/RugtMLaJ38l+oP
kKRNNzfZDPxX3GGXU+z7V0fDlgbdZKzvUcjms/QuTcbZvjBb6pb9dl3jYq55bEXL
Wznvi76lFl2CXwdPts2+pCowIuduhzSYFm+RyhXYLdavoq5/rNI5F1ymr0PxblRj
o9nw+6e3JAL+nr/8Bdj654xkr4dlu3nsTOJ8tIv2+2tAXS5qUBrWrPuPn0Mj+30F
0gQ4yjfQjzagIu8HyMokkHq4y9NYqQK9ORFSESmbiHBpktiyIauI9qHliZvJoX0Z
VV8VhAL90S0pV8VQElVNWogdMvOFwRf3rNLZM0D1zochRphdun+UUqMXh5EFozCV
EIwnMSHa78WpWzhndpZ7fY36D5iHEAjng9fJKThFvbn2g1ZF0UYPhYs9l48z2GBD
BCb71PcgE9Hrmm1X9iS0V7nnghiB1ljuTNIfgOnQpAlK9hysfhFjVsZVjzBY1MGo
D++HN237wD5uBohMfx2opfcoCEd81EC9A9uxepeO/SBhH0LaDJcUFeUZHfLfNZaR
ZHl3WTCrflsyCiHpMemMO4LNbxFMehyd+/FHqtDHfvwSSj3W+0P7ASCL7wW2c/ZK
7l7cDMxXzJvFXEHFgIT9HiQdWsRNNyRUnTgKTm2Ft3WCqxLzlcv0aagyyulac3Um
qZQP144QlLpB8FPE1TOeLeGCP5Z/y2VhD6DCFEZir1n82GgHOT6sT4vdwrGKqfM2
VNkLVmi5Wt/UzkB9eXIJx9DNoO29wrCqpOhyhzxuiPo4rOlTnPDwkhSdkTwoE6e0
bbkAXzG0slQmSCgZugsomVFq1YTOp0EQ4oPsognH+LyYoYOtutMu/Xw25ZI4Sgga
cHW9GdZiUaUQChdYtmg6tvGgzW7gmSBFCFRSl0mxAYDr6RPnqBllPnV2/FjvxbHU
IAnugEn8raH5DRxdTBtI9iI+RgObdDg2DtvaXjczJGRBUGSgf8cUsNaO3Obids/A
ppPo6th2fpkPNzR1kulLNJ/E0RF+tAFZCG/V2lsT41bfSzZNCgfp+dgIS4p+ihQm
V8qWjmVm3wLmp65tJCieTXMpUqrzMoDCsl0mjn/CF5lrI2+C8uHhE4+l0YiWTHB1
+ImNItyRzE0bZox+mq6Nc5P7lVyTU2YhZe8UJnZgHsDQy7vwtgHJp7fy2Ji1n+LF
NTIhfWSLH5tCLSohsmDnio8UNfReMAibPaSU4yUx25Rf/KQihfuR+/XSZ+yCD7tj
yE8iXc/k/SsuirwmGjYbw++8TO2bYs5b5+KvdVISRN7wwMN26zmVxQFhErufVI8+
8bbs3Obplidi3qt/fq3eTfe2RuqLontU9dIVF2jr3YJcXMRbkxpxJWugRxyAK9lQ
U6+7yW7aZXI3XxuXRI1J08huISmkfilTPMaHaM4c00/P4wDVhXcVKW6qRcUyvke0
1Lf3zQqiQob3qojVW0edraac1AthPQV6sCP69a3KEudPHptwulaFIT9arwwDdaEX
eXKuUJxgEIWi5ld51tKeEi1W2aRgT7v0e45mly0Wowfb4TzU1Cu8G7ijUvinRVQf
/yXYidBr6vWwxMOMyP/zA7z1TXl4LjVyWZGeJmQo4PQw0hBvmu2IcNzZa3Wbtnvk
U2igP7zcDRVS0URGlQisEK42UqvrOm8zWYdkHLUc5dVEZDBGTI4/x81upQgO/zoU
rBLgzWcjW7v/piTjgycuiTvo7yAPfI24i2K3SERm/QRSUDp02a2f/cEIj2FR/+hb
PC6EBkITSxatvaS/b9b04c7+0pSpxzVyaeYHIysr2Hl18JvR+S2kf2MWUagunR9r
drzfzkQ+EN3TZ25oyxUyD4IaGYWzn5JCx72OtCJHrgxQ0E9npLtrmb9F4/BCOe9k
ny4ZVU8aN5R93sfodIKEYVkrXHsF3VNoOAvq0Zi2/yHAKCrRew29KvPMkJHAUgay
8Qkg5UGXD7m0neN04mnUSgDHEzdbmcALdoOCjnUTeBuCM/xkM8SQce6NP2Mfv4k6
G4nX194PCXK95+XacH6+8oIIq5C8XfePTyusQ4Fza0CjnE6mNJTx5YiPzLPM7hv9
Yiav1dLPxgAO9QbxPO1dWE2ueZNcSDZbvaKoe6U8nO7BqzsOp87JEuCsqUznPoQl
0HIpTtPqWh5qgj74tAym4GrMx7VqzJmJNhruMfbNeut0//BiwOv1cwpIPxYst+S0
c/U/jXPfPfu/fW8pGrefdm6bgtP+Q1xurmH6sffM2i7m9YeXfssFZJhDeO88BKwi
4rMzERhlaqFSLZF6Pbg8JSCLv1iWtGODPupqPhsy+HvKfO6A7mcsML/Nd1eAiQNl
ks2tqMpgA8rqDfWfhVTPyoX/Di8eOCC8Rv2z3493D2yozP9EAdlD/LdXZqMg7gJK
miB0RxZR/r+nrlKwqyxWC0Gg+viw5vDoG95vXfQaU1V2hHpuWag4LCuPbtGhFPQh
uhBe15xszR7G8KtocxT/I0P2LDlpiJYdt83gdqGI+Sov5Nm3iCmjFWX/aQGUqk8b
vkYovdCzGGTFAzgBdF3Bc2lCHTE8ABEbopQl7LhiSEndBQke7j4Ev3QZNn1y8ngg
Ias2oV8tdb1R222LKIIPNdWvpP/6Y7JrP8hm7rZU0yvwHuLa/X+BulrjDPmtPnYb
jZqFaqMvmlESxvc+RLi/Xg2YudAI2eTvTXtKmQ5tc+KVv29KqNMfqVoev2gc+aha
SLb0SpFR770F8SL02bzAhXkkWIg48k2g5sub1G8tm+7Uo2XtCvb1eMjcv6buG1yq
mgeETeJCvgkEnZFErQmXZ7tBNbAgrhCvC9V8O/vr3a1rIDSOU9WxYkgzSOjUj9uR
/i/c/wB0P3LOnVp4mv/kalMPiMPmdvMipedgTFo1AF04eVSM+IMcxTG+aBSznuo6
3NDg1suM4R+GIJ6g9vUqHa2q9pJIvty80hnrBiakroBPI4jLlqTMg7rpVSucDjNN
qURV8dPE1V4oE6WAGac4+TArlSfDPslH9fJZgMNj2sgdBLFa5nbDT6w93NMmElfK
u7gvhm4mcbTqr5hMLiH3qzdHD2Ynx0bYyUmZRiuaF156YdDrzmyJ2JtX47tkYz1P
kzyNWFBJuTeGhVSSrS0ifEsfo81q5gYGskvK/Yu7mjcw40k2qkAx0ZNV+3XjP4+8
nImLGJloRR4j09kdDiCp6Y85c4XpXCLDihMsFALgM3dWhtUWVdIeCY0lZd+s68/f
1CvgUHiIkhXHAKQbPN7ao3pfgxE5QOKA792xW9zF7C4fnBxxy6k8PnHSa9hWrGtv
miquYvH5Nnf1ehAKBAKPg+SvX9MEgcM/2vOUevcg2xuoapJ4wJIIVQyTbWdhCBia
F8OywwRHUxSoDAd99pmhWyYrCxeO9Gsma83xv222SnXPN4xun6GDhNnTDfUumMm0
DVygEd6835cYGOeCCHZXzv++RA7N2Mhjyinz5Mr9HtSBmZ9ZS4/FhGgYxvvR44J7
teeuUj7b+dxBT7dgYDMlF4RJt6iT45NA3K1Eu6xYC+E9z+6knXDF9xfvn4SuWiDV
ETr0e6rD9p5n2zLkic5MpoSb8vP23Q2VGX4XF2z9kHMisMAYHFQbhfzYV+gGiIgt
5c11AWVEwZJjI9nOk+sGMAAyPn2QddGV5puA4/aEKUd1oF2OP1GlQFf3DXmLPuDA
pFnOhOkm8zS51Zl8Yzqv5QuXDpwAEthli2HrQt3353WhkM+NhaIiRK5jai5Y80SG
vm2f9mDk9eZql/4zx0lSkDvWiB3XjrDLkM4l1VPqLdE10gtfdGpjkKxRRLkbnZbt
nHGRsLOClebQfClqnNK9UyML5D/ZkDGR6r3+RR/pjrg45v6KlOrkUXxfw0DqG+YM
Ad2LS7l4WFEHhK4S0XOi8IbkWDOC2B7rAXkLXaecHXMUjzy6DB13u38Y0aDlpZlx
D7FpZ3h3N3SZchEJFfflbAdFmgtGEI/lZekzHUlc+kfmot9Bp/8AhIKyRhrrRf0N
lX3Y9D0Ec2j9JITqp65Me7VtUJojJhOnZeo2ZqMrXPavMIBHoPrHIPhAGXpbFTfk
TmjpGwEec3gWGm2bpN5/sx85o/FoojETrDGDx2yfBF3di3tLxSaH3gxy595HhlA+
MWkd94X6EhaSlNiVkyt22LFizUZddRBOfgXEGTanc0kRad0xn5RdoLuQ+mWnrKkK
nljPjBPt3Q+2RQkUy7+YWJ/zQmetESRUvEnVLG0PLOcBT9iPObibdnMGvJ5gdk23
RDov1Z+lnmr+L2EURmZPoPENKGVQc3pwOADfmfuAlkwVbfqH5yI5p8hbu+Jqqt+q
rtgw0CHB8TI5a1HQACWsPdFdfP9IqhKMUB7Vtsr2kcrXtSa/Ye9pyhkh1avqJj3W
zfgCE+MmBf7Z2kOD8C/9A74H1v+2TtCP4oFTquY0vei92gusa4NUF0Q+kwGGJ1vx
KamR369NciYbvxku6x/qM3iZEBYXiZav3WiS4PacmwwLwVOGAaB+pqH4HGanppO8
csJilGTq4erRNiLX5dBZf29T0A8WBwyrmJevKGSTT0X+YDraEE1kpnvE20AfAxoY
ZIXtGrUa59bzAvLZzpx68ZKg2BVclnWsn+o4ZBjsAb1+nPQmntMJEfd6CmOxWsVo
8nAzajYQ1RmAIwHLTYJtkeuIeDKfB1DLK+fYtL5loFUw1bO4IcQ0033MQ1JNfuLL
/Wovlfmc5ATjCyW0wkGCjdlHEb3p/pbdIq/ubo3upEtcdev11mKNFqJyIseSBAOT
3gvJYF4MoA6c6QhLBuq+uhFzb7y8H0FnY4JrrZsdVQJv2A+a0rDN8LAUQMybUwpG
cOSDyJpNB3HnltHEQp4IAI9vZ+Wv5RIp7zvPfN+dlrjVsONuwcuL00Yvbsb2D7vh
2GjuaphSoKzk6pKU5Dm2GAmfIHgEmF62VUeHal5Nj2rRZXI3HgklSPnQKCay1TN1
1Q0jr6rFnXawdJInRw1AXtGJa9Dc4IxCjzk0z1/7MAlu4bQhdb5FJQPnm5gy/Fgq
DKazZZ82+W0vYRvSzrcjKlqGNanVyYh3OgQYSg/McAH70LZonqo90YMqmvXVVNYO
HzmKgwJ1MIPS519Ra6VGWeLLcZuPeF3bB+Kb/YnQmH0Jg5wLyr6ttcnD+wSrHomE
7FMWCBtpdpSWfyJs/TFD9jb1Wd9oZYRJfHkNgT61HSnawP/6rGqoGfsYZarTm+b4
E+NMKR9pPz+psf3XAdrEUu4fcHF4i+4tnwqx95boQveItwGqqhMzmZHn2zgxVuz0
6A3oOJT1ailPjP3QmX0JNIJPFeNJMwKmTCkHvzebdda+TLUTdwQwFnyEcKzYq9GQ
iSr0CbAr7Fv0kwrx1zGiXIK1VbSrIhQ2y+I7+ULTHutjK6/+VH1VwaSKIuuyr9T/
Ab2mCL8wVPilj0sLIww9ymcvvV8NN7aB4tI9Ouh1kwloj7A+q5JwQQAgrcCUyfbw
lUGc5Oam96lXuY5GFfqWHy9W6PtY84vRv1htEWHlGNjZYiJrRQOLwai9SgTvw9Ac
7Psi1ml2Q2V71lcBQEvzrbd85/BtIc4lVMSamELuX9EZQGBpzVGNCTJq6kqI+m0N
9SdyoSlpESAKvmw9/d0AnnILgxCF7qrJk+qPcCYnPifLaGv4i7WqpodpxkXIfb07
zK7nZe84K94qteqivPcHOBFJ7+N4ycnKzdmXR2mM6yVaZjR2V+PtN5RYInXjiC+N
qZuijsLwLsK2FLnO/A9iXvxe/+76jDY4AEYI458K1N97hfsTuYkmjA82p4DsETok
9pUsjH+P9AcXZJjdTuunk1fRzva6i9RP5Ofp7fhvLsyysaIYBme/ToCgVocE1sdT
TQAHTJFTCOUKREXaE4dMDbryHtTwZtsyehmrvweY1ElDHZAsx+9QPq/URP7MW+SB
aTPNhuzdFYfeHthCVdnngNm1rRavYni90sN9oZpvg2Bxvt5wh/dhTVjCa5/SprHC
AjkpnpyI1gmnoGN1BsjXfSKXrSuumXPdm1XFCOfCArqtFWX62pc7beqxwDOVdVvo
buVA9Ir13CTDGCkNov1/aLjoL6FJhRzI05J+etJWoz5J2RghCVhfw4TSKbNa7bXx
6lbXCZenO8cbIfsau5x35Le/vq3joPgwsmsvTyGGB6ISh4msFvsS6MBg0Tw0OSgH
eDsJ/KcnjgB07cMnum28QqS23eiVsN01GEV81j7JOtQIJ/54UrcGUv/qOpLy+Nuj
hh9JCHJD0Rsy6hI/3t/O4JrU9G5hRTljR7RwfrPYotLjjwbmcI1rkZ6qmT6igPCU
PrRDojCfDo/CmnqScBW2WTY5GxNe9SogT1zIk6UowTGDQ3c6pXHfk5CJha4XsBUu
4r0fdj/ZgA6WYqvsikmo/Tk2o56czGlMYxyL50HLgtyZ6fiDopuvnpNUJgR8VA+3
fjUGaQR2bQLVzpAWOdoBA3ROzDQNVZ0nT5Y4rsZQaKBXXdxVdjtkBUH/8L+a1Mrc
FXLYk0KbyaT1OHHpHQy7qdXNk+4rLINV2DI6we6M8k3Ir3z0rOQpqZHIZv8c0W7u
5pRm+eUdf1DpZezgS2wHynjYLNOB9JIVM7fjHeG4DdrwEfLBZv0+y/gYK9Z50Uiy
nTXEtn6CRR2CK9bo9onzGfgZmcUyZm3f7i3Mdm9625cAjaPhxnS6VT8BsL1B7gfX
BrCI66bSPBGs3TU5YvkRQVkHbhKUyRlcomY/99j0dCMMEa21elBlMBeB1Qou9bRc
y5RBRAizsKlqBg5pea38fw/baYk2L1cY/sg0Eqn5U1dAEUuUVQwrfvFKXYGiyEZx
oj9D3BSxS6iogWg11HCDvQaqxr4wEf5K5sheCNvWLh5CRYMpdQqiXrPgwCUvQpM1
xjq92RRJUztE+4jjKlCjGL9FrNs3jH/uFJjZvcQYww4oSXltG+nfvPMRCpnt+/EK
IcgtA+byixfzQ6RZKz07W9o2iJ3HNuyea3y7RWyCdLRjCxjvVi0y1ZW90prQcYms
vOMcjbCHLlt7uf5UuUW342KVJrdDDXubZeEzRvekiCyQCdSTI+pHzE2qCvyBuzhj
3+HpWpORqXhD5srWIGHzZhzSPFGowg8iBdp8KgV41hebtr4YWomkQjfd3wVSGMjw
4LWj081NQpWLFVepQQ5k9e8aaavn4nciVJ1WEpAAuI/Q8l5vjo61PHM9HyQX5SOm
YOREsgCi5uvMHzqmLE9nus3NMfdXhlxM3siQ9SXOpt+G/HIWiiFHyDhshSKbE7WN
pG8KDcvWr5ip61PJpeu3fg/vg5DcNQa11uNOsxLF4iOaXRO8wp/Fm0GXfBi/8Q74
Yhl9xTfjDJLfIKIUv/1dZlMMqxwW5nvI2rGsZlZNsh2CQXgsaZrpnGN87tj0Gvfe
xEPwd8AMMVNXl04LpGDj01b2XXKSWYA/mc2SN2s+TkCaXti/NzzysaAwKxQgj5lv
ZNrh3YCNHBfhfn4bkAOrLYRVf4qWhJw2mBRd5iiNCn5bo/GFdNTMlQ++WhMpGGNP
j4Dw+fm7koZVZs5XMS18AYHu6VzsEvbLP1AjykgfrJ0cGgA4/ldApKFT4mhv4/V2
YGmS40oHLJJhmMTYGcVZAG9GkX7iQ+nV+AmEEtZwJ8S2O8HgpfH+zBLu83BgJVJp
g5J1RItcs4GY8uErNBHSoCcm2Ga4wFMSEVzpew1uhbvhknaxo8EARdkYQ5Lu2sqQ
I2G0JK8Vo5/zurZjylZxEC5yx6YnTzUYNPYIlgQOBz1T3SeWBSj9ZDSKmvcNfr/I
EV07WWGQQrYiXAVuni7zGZCLY1fKJac1FecTfd/Xl5N/7U5dC5NnEl2q/qso3EX2
VDxEfbPhE1CVDWJAYEalS4Mgid9CwpSvQp7sEJ4W55je7m2IKAzY79rCkuKemyYp
GFKhQacNm+SG5rW6lWRtOEvgGRZgNjnKGFaYGR7+SkinyyKvXczsmbbCF2CCZ/md
+uuaGLer7M+hBbNNhwmApa4LJB2NnMR8jk3HFjZSByVZqta1i8WWrb+HFjBKFhjl
beMc1d6k+sYPFkKkXFeni70rVeqGy8OGkVHnX55Ybk/T5hVkukan8WTrZ0znLwP9
qkczOsIIWpLV+yZ3ZhQ/+uB2qnxod5D5lbUhYsnD3dJwDI/cUMMxV/WZSpBNkkEp
pW1ZNtnT+S2EANdDIRpWSBdYoRk6xTjYR49H5fEbfA7pSAcGFvCyMo9ZXi3k9SYn
TaXL4Ai4K1FhGlvllt+df2WOt+RD576vjqMQu4FI+uTKmmnAZMZczV34bX/TxeJG
HPkPOTMbBBfq9TRmy5VAGFGi7tOEVqB6i8RUU8MmLytZynPnHQ/10tTwmzyuY+Ru
nVQf6gBxOjCnOa6aZ1IFEqIz+RIU6y8HPh8Dq6ZtrqaEPG+HM83q3GBqIB6l2kXm
9In+FpFEu/1p9iDG3FXV34fERVhLtzLGkaUzByaULvauHyCLi8VLyBMCfTd8BZ3e
wcAC6E4+ABDukNGtBqa4xb9GeiHJ5/oQI6EWAjcV33KUrv5wQDJZl0poW+c7kdMy
JChDA3/JtY05FgOqOb6FHq7CRuyxBceK/9n6RmXDbK0E4q9UfEbe0MKR2NCFfF5I
1hTWz2rVFHy3hOXSug2fZUJLUhE1j/2gUCFamX34MIkkeBPyLkys3sOfxkWKuu6t
arZkB9eXt9YSwQ1Yxjq20uD9itYevPcHZkPQFRr8xfzXVRw8lAfbQaVYdNcdh4KP
FoYUeF9FfcQcv63stOygWe22WHwtNqOpKs5Ct/tMXqsmfbyhuoSyFrrMxj4T8SSG
t5/ncu4ocucn80TrVWdOQNlDhp5r9P5wjtY6qqc71t6VkHNCWmBUB4mUzkblCWHg
vZyirEcDsxY+D+XVJqIIdvH92A1KhN75KPm++UebB5Pp7j6ntbqsVMQs7Uis3+Kd
z4JMeTloPdX2A2mCtUfrzzPBlEV5nmLwVmyqGtXwLFKLpjKH8R70JQCMJZWEBYpf
dwzDMvk1IED+DxokAUFuNYTSLsCNJtEsjPK9ZxU2jm/URZV31p4G0/JNRlGJ09FV
Z18GYb0CE5rPa3rOYVb1izpVz58Rm8GXT/dVYzIrpSqFxkd7eyWhNPd5oEb5NE59
l+DwawBiK20CNsTaP0PloHosTehYONgIX6+CdXmP09abqjhGrnXb6kUu/4zkUWlx
5qcMJ7XGLjxSQxWtHMLGYCibCCxwJVwg0ktqCR2LmeflwRj4jPPiYE7m1okO2eaU
SEf7kzGEUR+2JreZMcOcB9tS3dE7KJOxduWOZkt6KShPRkw9ToxJM8bU5oihpFmJ
UnSiLH2Wr0M/VagNSq550Z/Y4uLqEVgBNrKDR8PWmgURxXhiyrrgq8SyyCw0DQa3
ipz6SViM87z+G5ckreitpsuUu7w/hGXOoC8mDtmaG40i6/HnG7USu+4n+C48USgL
Id+/Hs4+B+ODZE9OikABGyiNCvryQbtQwZ2fUwNXX98JKpk49yQh1FS+lQ6+iQeJ
jOsVs3sUcyhn4dY75JyHkEr4VUsvlCikeFWriC1gmru+dHJunMVhGd0hCEFFKLUG
1KiC8zh/rlD+k1tonptSfGt+NYrKjauf127SWK+ILFdTF/35tfXqbMxQntDcrZC6
m+Hhg4eQeMntU+OA9g8cxZ3DtXi8SpHbZ9vcYG0HmiZ9OWJ5FkhYVnPQFhwHtztG
7qWKc9dpK/lsjGtKsTXrYxIOrKohkv1wXMaXxoc+kPzJ/vo+zauYY3pVSMthRoUM
67CowLv60KSFc4UsFPEBruFjCMCnyjfLMS7AJlyg/Vmx8p6vBWKELJ+7k16p3YqS
bWYWFEwMUQclnoFpqjivj1dnuopUlyV3P7eRnp85zM71U5aOZyGnHu7HDdU+wgQD
A7BI2NnJn6HEi1/zln+cQtl6smHUhtHmZNUZwCPlsnU0HwUGxnOERdzW5qo4DqQv
xrXuzMA+EKSjpYe9XBPQXEDxrRGaxQ85Ek3REMbPFNItglbJRGIzilEByHpwrhMO
NjYlVXz0cz2U/+1Ew16HuQ6HIEC04rb/IqLWjLVVTFx7qRiJvejnFTKzIMyaiy8s
07IekdaGpzDGCfiHmxptXCoOwTNtxBsnJh1FthfD/G/YYZEXQ1owWEXnJeuntXlI
tdAW2v/V1FEy0IsrhzMFDTEeTxrrVvnWMC+E/jz1DOHI9eFBLrh35lOsf3BSrsB2
uk754I8aY1jc34uZwZDc45OI7j8mOdUiSKkFQhc12o9MEPH6HkNkUT8GcRTT8Jh9
jWzoqJo1r1wNbfyzwIAlZl9vefWl8Cb8cRDOtUnwgRaW739cvjfv/1yOidO3hTd6
DIiXzdcTFe+9AcJvkx7PdhJ9J0XPlSQPfLjUPdUYmSwa/Qq9qa8k1mf5r+t54x2+
xgolad+pqzLBMPdj2Xe0gnYmuZ3JG3qnnUMBbv6+UNEb43gSCM2d+QQHJBUZHzK2
Y14wpoyie5c0Sf1DuadjmSDe+QXBVrmlPpP31HVIC4APGYQ2YoVqCx6miXOzcQIO
WmQN8Xn5dQlkeQkaXQrPHqt6DnxTwUpz3V53AP1vPcgf5BSYK2rfNOUmx63QFQDj
Rm4Zy/XJ+JpL6FmSZd8l8noDobjiBH50HR395xbWP31qy/SA+zHQoySwjRp7cI8i
gdZRW9+AQInoVFSvcnobmdlquPGCcKJoZ9SIeoEY6/zzV3P5bxlWZpG31YpNPdQF
oVBf2dtSgQ9LO9EEu2KBSI0wnRmdlf+CbtCRcAxcYZ4b2xdAC7SGY7tL2aJlYRi/
0NYhjrUfxPMgDcNEp3TZOzbTIc3eUga/zsrud+1UnpDvG2u/4VR11lIcCpWlaxsY
Xb6/admmNSl8AEyu9JH4FhNqSEsYujZ85lWlwMkyYkg8vXHI3QbGe9vn8+CtvaW8
OkZ8VYP4cySecuA70L6s3oZ5LmAB9XY9cO/O+iLSQ4cOjEEqTA8XcBYNs8EQiw0A
TkoYXX+LHVpAHbpGQrOyaAW66VWdPn9H3HW97kQ8PEr95yGKH/azPza9Xmstbwzi
ZsSFruSEyjUgLEFXIE0TpVtKJ1amt2VOSh8Z8eLAUt/lExvoMzx/0rwX/I57VDR8
v2IWQa1jTHnwuMfsvaNbdbXkWJ4PUo9vhB/bH9a5gFWRbI+2D6dy769dmIXZtAE9
mMRUaL+xJolMddNZP9Zi4zxcghj2KqMhuJ5j4JN3EANFhWQ0fV0XfYYMe4SW4EaL
VT86OZjdLwiap/n4aK9CgtIRsZKqFVYYuqlMlewUrnBA6UWAlalTjyC4V5CFt9kX
1X5VJD5VNHjNDsjygeJ9hKvebeGurT19OEjUVuf9Fr6Q+SRasodIqrt18fqB4xKy
3FKKE0WuP3TaDMpy0H4RdzSQd3pLY6xH18IyZG/65NswzttOSsgBMpGvblqZ4Uc9
7bPJcxcEv5Vda7VVhzZiI7YQ2p7ikFg3YhsuYkCnYHk9QjeO/kL/cfuXm9DcJpT3
8RWdv5+hIy5v8LQf3J2u5sTN1inyt+vmSbEedBQxPPAF3S7rRLmmzOGpwxP5EUTS
nIZO3hJ9QyA3mq5Pre2YS4IR0CZThXNkm4tcOdKDhDBpnCrejaPbPCtPITFos3HM
tiUWbvOdSjHvlFuPcVqVWpUflER5xuI2YeqIOHvB0/aR30yQEJdFB/rdZo8NMuIU
SEkhkju6qV6dKYN6HdDYlFds6cy3eS46RmgfAdhtmIONG9EJOMqPo0IdYd4h6Hvy
jLDFDZCQSP/LXBaO9UJ0NPs+IvLpt5wxwUbb12oJ4DOkGSl1z47+5bc/HRWzPMf4
2/Fh5IKNa/kaKG9aOoHd0r54fdOyeXk8C3Tfswd3qaP3OZB/QuDzheTAPcvce9IN
oBpLJo1fDDzT4Rq3U0RMmF5Z53O6eIG4N8/hc/h36ruRe3evODRH5nYJBaM4YT0S
2HFJKFj2E9c+2J4zxcI+9D/7V04j3r0CGFqNarp0Vak0xQlYgoMgoUaapiM6lbH9
VCsCiA1FgnzlGWekwXZVly4GCstLSHbXY+ORBXUhFIy7GcGEsaZPAh8xoJ99W7mx
njnLSjBox/1OPBx5LhXI94H/xD7nSzqJxl8/dfsL5RDn/PLTOn5vLC7+gmdWf49s
laISM70vLF6o8RhvkW/xK55tlSrXjAPJKZbcA28PN2saQpg5le3i88RTkZQEKcDW
5YYg91wDnhnftbO4L3+5gOagHDomWDVysedtLonTLtwIntK/2xoQZOA213WvX60a
g/X9PD2dkcUrU0K9NMz7YA4bj86sJ5nr0iNr9LvxAyMclpN3JoB1ZXhIqOLdxQis
ZIA+GOO6b0HB3Qs/WaRDsTS+6syNIFaNcA5U6vQS72Tim5XB4zh+dwdRsO4IpfBJ
my0seDHDmpBy8VPeOF1Tlda/NDFDL2R1t/jHUzNMXPK1i5XrH24o7pX4QQYll7Ec
FHYI23afSsKIlzA48VNMwvb23B+oOULE4qmlRgpDmFOU04Fb2LTfZCdoZPrbvrfo
AhWfbeMcphHf8uTryzwgkD4OjPgG3faG4fc5XvITOJsmuCEmkHW7WvGNQ41tjrx3
a1Yjqrhl51NSY00BSayWlUinuFjid7ch2Iue2ptLOY1KYWGyOhPcb223OzlKm0Vd
RDTFHGeBINDkwqp2QoJBdDT97S4M+o3iINK/2P2QLvBuGQmiI0LaHeVDkM+iGfyX
My/YktIOeiG/dR+debHJ0MuBU9uLyd+2sgFVpWugpccZJhzAWaJAArkPJrzxxxfW
P8Zi82dCukyiETYw1m+Dq1xCh5V5yDI2nZuy+XdsQX9BoQteQbQuUlTof0UM4ELU
`protect END_PROTECTED
