`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oAXtemYr/0VurvvyiOFPQMsF1DFlo6+3gjP7wBv33BmkUpr6y6PVW2iR5H708lq2
BntyERrPvvbEB6DW1asm5XtThlQOI1l+abPHYCeLi8dPsjbT44dJNQk3r/jPWUcD
rliHP6kyHsVvjM7Jy+2QNXL6m9TAbS3DvGxQCTD8PRy1DxBPxtJDX/6I430J/Muk
M5Mfqrs+1RunoJizmoUwGZEevkzmx9bqrAvY8JJyDVqJrNL/qO0vlDLC+d9bzyqH
UKXWPGYpI2LT5YKPlJjVrfa4m8gjJx7MZbCuu9eX+XUV/2UFvkV+L79ksr+YCI3B
cwOLhd5lUdUW90MB0k6NlVN/SuIvemmHrekr7/3OclGYeeP++vIECBYEPaLvIv0H
351oUnzt8+0pyUsu6iEVM3gy8XFSih/6UHRGfCt0+qtb5M6Hpacmw9vQSpwSZ7dQ
7hswqdCCDx7Q6ALCI0IS5ZSsAZCrQOdwBNhCF4nVZ/VnEuiKo3WuNiswTsdxlUNj
hJOYyPEq8umEVtvc4uPKr6LeZWpOk8sWMa0y86bd7CHFsmxlNAmzXaIeDaq6YiAT
ELAm9hfSiwrTQOw6qHau65seK3QFGL6zR2+CmedHOtRDN85ob010R7ADSArFuKPw
Kf9ETNDhuxh/VzcXaPXgM8Lqjt01zWid2+hHZ6zLyC/TkzS93eTcjGM1RxQbB8Do
5FaSVcvDTHL1/W6dbPC0TCzAPONJFtCOYMYBAeB7tjzT/iVYid2YWHm2W9MgdFXS
wWZFDSrULbVXHJFUPmk08kxaaP8kOjf1EWcUg4/3cOroPEwv3zZep61XKvvSFzbD
Rx81JHL1jhxhdzP1u/m1XprftLVRdGP7wYh9S72O4rXVFDYzOt03Uv6au7HyloBV
jq6wggbqm6ii3PDRu/1nZfpcIuhGWPwVu14eXHpvECQf1zWDFsvqtkxHAhwuognH
O3ol7Ef0F/GmKgBqxGddHzmF1BPfLI28cvLC282rXTdBbLQxK8GEuBwO/A55lfBo
VAbqiF4ywDyg4I2c3oZ2AO1i6uxs8jhTf+HneYgpAJRe3JRd3PjkmUNhHCnp+UmK
eA1LJTPoV+9mDHUcEwgw+cdEOq7TfAWQk5t8awH9lV+A4DnOdeILPXe+aVMAzYB5
9Tak0RFTgwsX/ebBvviPfJlronqA5RANIH6Ui2rassi+BxK25GfLTNo3CzIx13v+
fO4vpmtCiAB1VrQzx2MeOxEl/bZeuM5O40azS+6YHXRBgOqseluU5moUpaWPMEE/
2S2aJ6fRpltWEDLQ19Fo3WvBQr2yKee6uhnOrKSxuqznDyby+n4CZL4qjxklBSTb
rVh2FDyYpbctxzsxt/dvqmLLwx/Sf4+X2O5gysnGh+BIVhl1MoAMfxwowut1baPI
oqDoTOLM+D8vwTqFO/jP/35UHHMJf8Km/FKszxJ4lChUj1/2pNA1lK9W+NtabXwd
nFA3N39DVpgpaMw5NsDvtqEWP9xbr+x0fxDrz8XVyeWrp2/vddeWfbjF3xYrWnFQ
y+l9v+poKuHsw4iX4pFI6Und9o4rMSRFTOtNM8cTIEJmpOpU/AhllCKMlJhwOy6j
5Jr6eTDJZaTrNTDzwJTYdW4ekMiQMvcGA31Iw/2boZkjRisapOPjXyT5xFjQF5lr
1u15w9SmTPEX26JrFEvAD4/1CH0Td0FfpiINBNo/PFSt+1AQ9BajejMYHZUt/cTV
ykn8k1jFSF6NeplnlwYAreqQ5tDk3tMouvjCXuXv4kfTt8dGA4NifVXl4D+Rm5gI
uBS/Xr4708iAN6pYE4fzyCQo8SGB4m8nxOOTiPO4l9H54Gb/yO2I7HMhar3NDki6
yJfL8wLsp8Bzo2imPJRQuySHGfVqFDrcK6XyfVxBE3N0lSh1gCgbFZrCNrranT4k
Gfw9FdjSeR78Kv2DwycYPSVfk/sFCxg7AQpknNLGPUyq62X9pNGpqNY9OBSYEZaR
HmBNcHhTt82GmcXQvGZU8Pc2VvDCWeEJZAg2dM3Axv5WoyXGDMwuAmt2QvWgY+xw
7H6Qbc68RmsfZgWIAS6a5XAej3ET4KU4SlQW+5oLU1xLHrofGr/2TuSmep9qY9Rh
a2mtT2oi5xOnIvzG1T4ze39t0E8XDn6ar/OAKDZ8nowFnMAEEOZ4oX8ImZk6T+w5
cjbkmt8mALRZVw4282q+CCuiopxMzbwOLHz1ea/AauCJGMcf4lJlfXj5pymjRh79
RkdSJUSv9OXRLo/EqmkLixPeGQyNwiyNhQnz0mV+nMsmM2waFsC/fmlpxQ8ifRl/
R827fj+1SMkMIvoEl0f98iSTLpjivBr+DTW9pTEOVmQvVefkZnh8q6n2IRXigGgO
VkLvBrKsHElgS4gzn5V4jQWU7IQMMLpqSjNl2VLYPXeE/plNZP6WDirLCLv7zHXA
p7d5XfVsFfo93c1d4RFiwkIz0Ynrz63MKu7KTMQcM5vHCTMluM4tdjl8AniFi8eP
TPRhxpkt7RjYwrIv09oqMPgkRRZ3woai2tIGyL+R+o2VpDt2cWpzxPsF0D3B4smH
nQPqg9e2k/AguCcSqqIlGm39KQqEEdIA6tgt5I8bhg6TuUQeub5VeMIDB444o4IC
UrnmAlwTRBBAaOpmUwc0P14QFuLBeF1N9g2IFrPGANhAfpXy8vCPD00Nfo3A27If
uX69u4LpPmWaM9hr17LYV5L8b5wwBRH/jz4LaGDiUg+Mk1UsoBcvXq1j9IwmD438
7ORZHJZnJ/kdKvF1e0xSDizvj/ZgW7+Dgnhpu9sJSacLnZ+ErV5LUyF9EDnze8xs
wuBjECKcRMfXUuRLy8AVIUKhsbi62DDl4q+uF9NX47xoIAkfrEfEPA6MNg0tw6AN
T/B5iq0b5hApNxMCZpUD+zvtEhNVoWX4o3eV+MoVLHQ=
`protect END_PROTECTED
