`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
31hasM+GWDNwLrGtkvUNIG1+KyNyVdxOEnWNrSScD1pD8GzvY1Rl2tFGuCbN13kR
G90wW2SZQymlq8z3tmfaeQ7TD2h69KO5JTx5IA+Qoeqt/vN+lKgZ2hU5XmZaZztG
FwZOQspze0dLWsD81o9++LF6X1WkqMYfemmA6WNzHS1BQQXlE0/tRRbcXuURUU+a
jee04olf1vELT2F30caGzFCOeLMOKXS6ZhrPkk/Lfb5Y8tuhSDliDL9+i0iC6DRJ
2oWrcjXY80Zfms1ShCV6hC4vDmsnK+tsFRFjxOfvqUhYK/k72Y3TL4KX2WmNJxFw
d2UvRHkLfqxzoDBPlCSXrYze32H2eUllhDNkck3iQPJj5Qa0FFSbjh5YJKD3uG/S
U4G09mQIotEnBq4QXiAH0Yt5e4/h8AHhPEwtSmhU5/ifOtDQixn2YS4J0Qt+Q0zL
+PEpH+XGPxTP3CJs7r5fzQ==
`protect END_PROTECTED
