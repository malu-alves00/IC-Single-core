`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aZUPdFIPxyCAFNounyYDKS2lIpkLVn2GUuJ1RSGhVR5XDQhU+oUIUdGQInOsQozA
MIg6+0qi8pnE5fU2ZhmRVarSkVYmOFSmEVywwh7vSOR3LaGrif0MB5TUOBOQkg/e
anZ0eph3acgqHTMZdzNsEz5FIql/TtmSnrfccch0VdMJetctmqjdjpNcKr9GuaSR
JosVZP/injD7y9HUlPkKjERMN2b2vYeXcaKV6wxJmH+OVAObb/nb8UEwLXJB4bZX
jQc/Az8wU3HRlHeRSDE+TV/kFX/DMiPZGbqs7WYbkOmq/j5FTstvOI/i0bXPPEn6
PZrGR4tE539zvLBgJjhhbVZ0hypX6g1Tx/blWoGqIm3NAWTxY/bmeJ2Wtjc+oXiO
i4zEDtyNw6HwMC8eaLzJuO+joxR8S0cUf7cs6zpXwP7bUZq7+pXQoSslEBc8T1lm
hi0EukaCN0OPFym9yAhR46QUOwKFikXhdjnfFSCa11B49rZr7i7CmUC/MGopvXem
w6Bd+XckVyMmDRIF2Sr9oVhNkRXQpSz7s6jP4/ekiAss2Av4KxIC/sVW5CAzHnvu
oIIAiGvnlUsfxSoNDU9v3tOT45pxmzIGF6IFgluARR6ls0Rd0iIl4NlmiZepRCjx
ar88sD5W34ISUryr4zWZITWzwKQTSVQHROdaO64cuKHxtkynYZ4jbx1srW0H8IgI
oBBnE9hUguN4M9Fl1ieCwtmJo34gS8J7UPDBCxEJmH+VYdMe64fdnZRNyQziOePf
a73VSVhZXnCAVyseMDVUuM/iZOcggHfUiVADywtillc8TTS/wYzt8t6fgFM18EAH
4pDk1zVFXWMOk//W6PeC+wr/PB9DVtXO43sGE2E9BNfmDJDSG6XKYjm6lMjWc+jF
gieETvjRppeq99yHA/Dhzmp8o1sfHM9gHur78zZ3WpXM21IQ+a2i4cRho373E0hh
edEA0u+7bxXnz2Dtn1WKig4yZiZ/29iWLBa5WnFlEelC86N6rxRXhf0hOOnOCuel
fGBDxQ3MHgxawU1AGDB/HCANZQjXbDD/6VGPz8qW7ijmgOiZflyw6T7xsUkMK+4P
PZX1KcZ2FB5o90BmVrBJaEQbMurlF8q4efRWyzN/cDfvtRDKn9f1UyCLJMDzU5KV
4sFt72v8BUjtdd8d/hWVp2qq9Mc6D54IIAQoBG3Bw9bm1naQTK1t6UKxOURBROVw
EaDj2rf9M9HuVccsQStTgwabeZd0pa4r02QpiGoYU7DpJ62FAOPwVDPVX+3aE63g
B2bbDZy0T7NFp7cRmJgC60JD9XE+STO/jp3xA95qXvC5Dj4pIq77WTll20rrGUxy
7lqJLuAWqKxDbVYVafzubg4xge8mWEMh+mHUEXlT5ASlRWE0FqkWjZdl2UbBq3SU
sfqLZT1VeRWhFINEXowd8xsVqkH5kKMWVaPXRyXu9VZ5YBp4LZRZLNIMndUtq+rC
tKjPxMN3bP/rcFkyVv9kUEKFA7ZiaEKZbskUFIVoJS+oMf/IONk+fJ6DKJO73ZVV
CMXRTMjsFHpnEQTzByz934ddKaQZYFn9Z114Y55FVk6bvH+QtDj4Q5Jjtb4/9bFi
OzF2NUkyvWtKIBBvDwyiBQT6enKRJX8tmz26iaLKYK7ltpm2K5/8S0rjsvg1qvi/
Tpipgomyu05IA37qbr/H+Pv9LJJt57Xa3rMxqIMITRaluEDjtoDNw9qtfbMhU2Dy
WQFZ0hKsc8kk6fcmQni6jqAtXA5j14UurRaHKa6+xHkxzJ61y38Zhoc31AoAavbs
2KMejy9S/EujuF2zsaA+QgR+ZDl1ocWbRFrKWQ9aX2GRPQ95c6uFxe/1MM4udS9q
repJkdFsCdjihB4RBcKUrUFuj+QPPFwk4S5xYOAF4lbxtAVPNIfEuvBuBucSSluv
aXFkFmRUgGMGa+LWaAQPT7Y3o7lzM9Y2LoGZyKGhDJKGgCTDyJuNNSdSOL4TYB3s
pJuIkjBDBwbuWbREbiu+3NUzn+zupEgZQ5qlZoVBU2cZzGXWso7mgcPtfDwHMjEk
HoGGFE4A6DrEQsoZljp5OKGUlWx31PxC2StPeJl74s/tIgeD3ygU8cYUQU0FEoW5
/elsVS7O8xkVLURROomjRWOu3rlAlF6sCfHVSkQipSpIfp4+4vGYOcfQNRik1nz7
9/piqMwlxZX/0BZie+oExYE8nD5HyDu8IqCYBrQVEDvahI3ArfEQJqb5ccOVhEfz
LUFN7KkTfVCg5cKlKhbZpG//RwvqMJTNzlXNOA86106P3PnIUHeN7P5v+HzpzQFA
U0D2uryO/vAE2Lefjurk6DGYQpjP3juTj4LeXR2ValcAze4cBXkss7A4S/vot48J
OuMta4/6LvaCLV2JgNgZc/V2afP0N0eQyQssqSKX1j/1KB44NEHuc3V28e5STJCc
hOjEbd0eYGILXqjgfNyTpgo0UhDCoI8wP72/2a6+Qul9P7575kbRzNHFvpLEQg/Z
i+Oh2LxbAaF4IXpBiUoelPMmwiLDaChsjk4RHDeK6wY9fOJ9J5C/0duMS++1aQtl
fEkBRHHnn8YRd0dsuik7cMWtdNnXv6dFvJltlujuXM71n/Yfn+QM6mntjucVPC/X
MUrIIeM38rNUX4alg2J6818jVgsgM3SXkbbZhJxt2F4=
`protect END_PROTECTED
