`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tLkH7bI1oYzELtJB/Z7/LPCnMLLYeN5lZQTkL2U8F9D3Mvc0WMiKdE3meVbFC+BK
PVHZiNBHZzj89W3Wd/ABXY/q5twLmTwlE7DISsJkmY7VHXNX0PIvN4tPDwDN7HSA
07DarvSWtPOkdI28kOIrGkfBIOQeDg0WAPYTNlVrVwsP2VcbIt1F80GSN9iskisq
TZ+S9wGHFSUEomNhBzwwG6jC5tFJCmBIIydbw6TmJD1BTJ4VNxdOIKXXhZnS6k7A
HXi/kt6XdaAJbwIH0nQ0o4bndXZsAeOBc1gP4U9vQc+CmJ+ZwQd9/azR3N/6olrL
2hvrFl4UZLdGMo40KdWy4jYcQRWZjCXEKX593BgUQMd2wyuxptSJt3F91R0TySgq
xeYT2zZbhYCvUeuM8Flz/5Xy2Z5pBti3Ke9r3QR8fza8yDLkEXhjMsc2xFXAR28X
gvGm20Bwojl9GBXX3GLYzqCuL49rioGfOoTlkwh8yjSw4LGrwtxv/p7aC5zi802g
ME+qLxTsZAzXU+Q72Cehx1UAeCuQf4+PGzYYrdBM1UGus7IzWDmKSsJ8ZKd/sKKT
3AkE+CITi63cC+Cu3eF4nq3DAsBiOtrWQnAO0DuVlEU72WgWaLXira05FkXYeCMU
Kja2nnH66IUf3he7sRCZdGGFaRnE8z1tWJoV0kOG2LKd5ayLAln1wZTLL1PXIIhg
JZhpNDC0Xc7JvDGQodSFGqDK9IPtRtJ7i4qZFBZRTYojkXVaF7e/3lhdFYi/fDaZ
mBqYbWiuzEMTYsolQS80xXaHmbOrwVWIz+QpH7LWyV6UvPgwcjuazVVVC9nueFWt
MK7iHLkDphhghIJ8MVZo4hF0kF1MIRiqBqiAgm5938nNiFpWgNY/UfJPv2g0rdN0
kxBBKcCDFYChOkNl0NmX11vhyc3LuEHdZgMQdd4I6RR707Af3oC9yEm6lBHoSoE+
ieYl2lC0B+vPb2C4kbC54qEm4H6w48REbcoOvyLL2TZRyJd/j8Lo5ke+FFl619vo
PbN0EXqL4bYpnLWuQJJYmuBJiyNRqo3yUiJ0BiUG1bLsT9yxs96sjWnVWWENfHlE
pD7u+nLa/QiyMqSmtH5a30TWCGQP/hB1u+NevCfivaw=
`protect END_PROTECTED
