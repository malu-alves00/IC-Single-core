`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UleEwA7O6z8eoZLvd8/vwUhOk4HYOprISiHu1gbxF+EEerGr+cBv05GjXSmQHmpW
eisUXfc8IzVAHXyx0tLDmZz5mGlbtb1CV97l6OmU/Vkm1gAnFpPej+vFct11GBSF
qD66JsC8HbB16x812QP0DsmDIQRsx3KaJddiJy7c8qWAgrk8Q/11XE5pXRPqqZEQ
Hgl58dyytBupp6NSFveHsw97d/1x52KO7u0iKMLCHp8j+fhfhwqGEG2fjc7qMXVW
XGCJnWyVp6gqfb8VAhaZWSW+5hfS8fZXWNB2DQC6x9Ae4rwXYwJoTdL4lssiK7Ei
gQSyrWWjUuFJxzFet6TMjCJbJ07ASbg/0sKKQfTQc4Ziw6LLaBkWbzD15ST+Cu08
IQCqYgwRMdul3NL6lbQwKgbj0Pa4uazgWqQn9CP63O2SLTfMMGExlA6fvXJHL6+4
3CifRqWSge9LnKkzF+QHEPafXcjVDt9dJjeGSZ/cQSPSp74P+HOPzoJ1wp4O0E5k
oZUddeW75lEL6lxUk+HTVQ2T6OrlOKv8Ah9L1Z2e9udIpfy4wbw6ak+DOn9r0zFA
TYMfCCPKpnR8P/J9FoRGxDkW2S9jVtsQhjkdsSgIsI1lqwgnCWjQiQUfVtDlqrto
LocF0Rzlrgi+rcw90wwMp/bYzg0/A0SY4Qmb7nniTDbTOM/8YHY4rSkt/x6HJSuM
AWFQlsYfzEjUXfm8vyvAerBHaNc9qVFPd01iWQHojqfQ2rWe4QeRK0mympLkDhpV
LFvvaFsw0Ty25sjKCyzCzzTi2toU99TmAj0YNU/FRE1a+Pc62WrlkYD1ItSYT3Mk
vpvDvEbt9u2AvNY4IprvSEBCmv5Ho5luPYuP09ERzNxh6jkOLy3scPCfkgPwjeQl
Odd4ZPyJe5zYL4iCS0kPHtBSaIZj3T5f3URhW8MXQUjd4b35jcnyLa8nLj5zG2B3
HTnJ1SjMRquiYqrrrb44vIvCc9nLqw8NjyJr8IJP9Hl9mVzaasM6YiarcC/v9nRJ
EcRkkRERhJeaqrRoMOittFEpVEi6gq5UJC5AufD33ns4p3e78eLPRuKIHVUb/KfZ
HrGXDknuYmgDwyK2LNILXrp1u12aU1TFqkvlgyEkXs9+D2K12QXhoxdqpjqrcjwc
fMUGHp780hisNdPlI4rR5zT4cA75HsAX6bzNGiLthYu+Cv1btD5lvms0xL8LzY0Z
Ndb0gOOvDExBVkgnhVBt/CDAhwHdgEiBS+UNFrccwUnuaK/RpETUCpEI8bc52Dte
Q0LEBSmX+k9SN3ogVx2Ulzj/ZmIiTIcJWAsCkPgG7/z0P+LYuIS1Bp8W/I/HlMGm
nGLwY4lKEeIlLs/7Z1Dr9mmIk3xbGsTToGKN1t/e9abyzU6R1RH7R70dZg1345uk
1MvUk5UZSm62r76Ix3MFLUxiS1ggFH3MDCBw44rP0JE0AL5Aj1NEFQoqPdfoJHQN
eSGhs8H+Q88p0iAVUIqSzNOH/PEby2m86Gixtav0vZVIr6mdJBUxb1nmswkE0IR9
OTMlYmCl8u2BIdqpVlzgg4MgTWVb1AHsipTozjxRYTKlQrzkWH4PTWtEdMOgodXO
VF012xsK4cK/vwJKq7HW+vQnehs8MNF0uWpPdnU3MF9lZ7J0wkEmzxtvdNTRI9JH
2Elk5zLHvqBcCH303dw0cR8gRd4yLN9jsodSGMolcdT02ibyBlnLvV3bxDfJw9kb
fG4CsPYDltNmerjBVkxbZ0TvxxVpGtKd2dMYkhAwOiZqcLZN539g3RKDXXh7pLDN
C32e2ttdFHewwuuNXJLU4OkffxMo3vVamlOZpRbKnCN7iZwYqrFn+ADRpxXMSVlI
UeuALXdufTskmWN5PC4nKK9scIEN+TsR7xdCAa6c1TVS8rINLqGlx9AW9skOkhai
D1PUQLnjuG6B9xKtN+Yw4cS7ZAjorjsypPKH0fkTHOI1zdi/yPEmRi6O0o0cu7ud
wa/r2fFLjK+inoCfLfnlnS29jcg9O1UCSlw0xDjmHodQjby+QoG1+V5hiTxk4oL+
fnMibo/B0kG1hFvqYadUjuEHzbc+PSgy2a5c9dpAuAMopT5daPWG0nECNrYkowq+
XvjoSMwWqbSCJeBI3Az+80wWWncfCQFkBrz6bg2y3a+0/Z8ufU0fK+SeaO5mGtBY
FykwGrmyht8FmJVYhDpoNT9yyrq1AFd4qPyKR8NtmilkgtFNTcetG14IPQ6d42ll
PprZ7yReJhUBOew9BjNydfr4M9B/EdB5TE6WdNzehcn+a9YJMIlaGtppJ0VsmuBj
QTel6qH7VcE0A1nj4YTYT6Brah9Zg3hncK2IJqjO6VWv5FmqZ6sUIaJVIG5YM2w4
FNuqve2buR2Kjn55uc5wgGs8PE2UReuK/bAR8xhDuAI6jFqM/+0/C4zKURNFkfXG
EbnJRXA+bnDrQioWzVbRSmg7Rl0pbKK2ZbDSooE+mFGsVIy+SPM4To9TCV3Mk28R
0XEiL5xZBjBn3TikxLrxPQ/VkQkbYxjTK5fUGXiK8D6Gcy6ZhpXmlAcMN485gKMr
fkkR94WsGvkOMoDz2RXOT7g4EawcCjZZe1lcLtiFPZuSYc2Z9pwsMz/3vVVYSQOu
ATAmLt8wb/wEEjRp2r7Ae1aDuTbYw/mBIOgGnCznBcLvnmxSPcX46XeEE0jFxEi7
MWbFVIZTSO93RXeF1YFTmt4WXDP1TvLU+LFWQkqFpoYz8sCghNgsagEZNmbWBgXy
7j56fralPxMB0Y7B/j4eEGDi1+AtwnyoL2uBh0/+wFTYq8vfj6yzxDKKtFqKCnIw
NW0VJJy6oR0HFbMMND8VZEJJpWS/c57rue+65fOcyRG1sjmBXhvTxl0dHZxg706F
0tA5tgO5TrF4fvNpMRBVpb5INs35TkePHcoCTF6JWuDeUxmwegyHCT9DUcZsyjVU
8Gv+lltq/wKRfgBqLEXA4ebySM5jzbvj1jxiHN1n5GKffeQORKBMBu4nH1meBfc0
K+Fb9Sh8hT4k1+JUtmaY8GHGYee+EPAERCT6ibQXxO9S6PTIhkPjhkNdMco3KZ+i
qq78TeVBw1IB3f59bHWDP94i/Hbw8bmKD3RyoSg/gnqUhsZSWioPj+JXZSncteud
9BXbu2xXcjiF7g4y+wFObYfBzdj6GYKTeKP5F3V9bqJasCLL3eNUbD0YCJ5MFndp
E0HYX8r4wMLZ+UFRKsEr0ErntRAB29VlZxD6spJbulbyMFwBAsib4tqkMg2clO32
Yg3LnIXOdRj7a6n2rT85Bys6VmiV0R2wMg8WDhkU4hDg5Qop4GjVGo28aaAObMwI
fABf+c1l6v1yFEWY30NMrNlg62SZLM+807xdHTAA7L1IZXxNuLBnCvePhLJOhFyq
EUGu/ZORdhQW1XyS1fRNt5zfNdeHmYhjhUuUgVRXzlgxV+6UrUMeq86L3d+y+kyC
Xp9LQgmX/JsPuQ8vx5aLJrHNYDLIpNmOcUtwo95PpibW6FE3zG944kYiqt6ReEO6
KA31NDBnsDe9AgL5mjjMNNR8hjtAOrAGpZcqqPvPhD7MqpunCpQOSVeerbpv+xZo
5TuQ0KAw3F1u+XVpYMy0SyrD8hMrbO9IWH/JkmtuFyYFQnGAri9MKPc1WKX+SNZg
lXYf0nxoji5wIv3MG6FCfS+alcj9IfBx7eYRMd1D0EAJCDNSQkmnF8yLtMtrtMrH
E4ui3NS0ZpAbHFqx7a1LziYvoUPtri/6saaDW6syljdOch1zbjOUvhYqjwdV6pdJ
msyBaLu/YdAWyFrdp/UxaXfE/0enCiBXljq3roRV30CZiQe2MMWDnTzOqMayLOyf
1GIPeiLkXM6NgNElC8ilLkVy8fe+rSsBKGuBfpHjMyQqSfvZZtA0+vcjiR+Zq7jP
5hRH/pHSpd1XkNqUNXPf3SdrzGvr9WSS0h+SAYNM9Myv8s76UcFWYkk1kvouMruD
Fh+KrEU6CfZK9f7veJls6hf7Dc2XtIJAW1dojUfiNa4uQG/b3wNGgy5gHeRtleth
kAKZN8Ks47jC6/KoHcPEf4OXhiQWQDdC1wdrGO1uWSjqjV0DLZXmGQxTQdo3vPS8
FWZss5tv46ilpYUYA2YYalWLCn9rlisoUBBpmHczkO9rMtUvuxrWn2k2aMRu9jho
4uvr1tW1Ilv61sph5F/0kp/Q6wF6LVWsffhKQcCl/EZwdDTSk/VMif/QqlKzqILB
RqH/+WDocc2iNBLo2Z0KtGAZZpNn9VPWmurxPIJwa2QHYvzU1qHeejWAgeYpCTFM
vk7s7HV113cv8larmI6Ra9cZd7BE3WkWgBvNGAGsvrDMLPW6KNc5nQjx10Kiabxa
8ML4YHAjniTZpTV0dAHvQcIZY7ylRR+Kg2YBUlkXRxBb9vAsAC6OwqNJtmw2WD/I
2Qc0bfFFG2GBMvQBQkuQjhP3vO13aHGbhYOiTXUxKaSjXBwl9Cq1JvdBpera/3Uu
faN3H6Tz1a//N8BmuJszarT9K85j/K9cHMNDphRgwtS1qIwZbZkJ74ZPZrWvJ63I
XfBzT6DD4ijn4/J/AVTlPrfI3ZDv2TXjsLYUBsdHMQ6f+tGlk8Eby+3REt0QUqvW
jmdvA3z/SyAWwqYDlj4kwfCHY9A/bZbalQ+oersa+G79HExDUBqXq5JYMkV0MZs/
zMocBDT2Gz4x5dGVBPN9aIT4++GgVt223WyaKnuz7t6n7m8A44RDisKnLwlRC8+m
ZZooSXYEUJ5dgUa61GXL2ErdtgWIEK271ACjb5CR66en6ugfB2gLBlWEepA7i7/9
uRMhZJYCXxCp2iahkUYCLb8MC3AGKpbJnFM1Pa93kITspWzrqHOUSUVZMVtoynJ5
zZcKAKn/VYc1XPzGFZe7n3YgrgJIDn7qNur/1K8Hhy8+9EACy0728SNKagkNtcIP
xH40guUytY8m9OXmUwqR6EzqOlnTKL+OvpRwyrVZqC7fghdZIUx7B71p++qiDa7X
BsB6wBiITqQVFb9JLEHhZF5ksunsjXpESZK+ZYpCQEO9UUAd4udcgw3dAPM6NciX
pw9zKGRzvafzx/UaeerFzYOdWBGJjCveGqbOn5XVU8hjPb8b+gKocrKXFlTaDJ96
WipIcHzaPexRnrDvyKCF18Ret2ZvfXIpYRFJn+6f7uZTPIaNGafEhBJu2lOxqROT
JC7LcLY54L7USlaGvO3LB1X1uGsd5WpcZL9KiTlVwkEYI1HcufF4wpaoLL1xgsoE
AI1Hn0qYNLgTF1ypYv6SwxtCIOWyMTyWqqJRtghabxW0JBalJg94UuUvDhm1Ly0G
ni3GjbCC+fXIk8Cm2ITIZoFJSJ9oxG3+TSAmoYmmVPWmb6HF/7nmX6Ej0OS6EgYs
E1Tilnj/ljjrxbOxT6CaOVeoBQEVIQq/cED8wBi/Wj+8coYzCrbLjs//dSyvrDwc
HPLzzIeKWAWygs87daChXwm6BIUwVeddfrmn01FSN21hPuuwBam7R9+OxBgImr07
4sjI8FRCDhdm2O+3rbB1bEWvc0Eax7OaSfS+6DfasQTzZu31eoqrjqm6qM29qAFj
Bu7dBREa+UIOtesAslUrBGzBRC4jdrTA8QtBNRVm3EoG37KU7XOfK7/jWOR4glye
7OUCJh9TcpNNX9M+9oDGGjOfdJIx3TYP4PkHewP9zc1N1HV1lnut9GLWJVLyjtwn
6gfBryVitjHvbkc4zMuAUClfysUSHQmrKRkSsjFcdwUXnhSlj196gtPvaSAhtrhf
ABvLIh+Po80rK0rYj0QN5m3A287/bb8H2AUL8+vS7jEbij2Gf4wAnI/X5WLbgJlA
dcjYsa7+NKPgHwsmAIXNiiyLXlbg+uEYmpsesmtYpN6pFn7vuwTosaaYCt5XnaQt
fRkPfvYCaa0nrFYC/DQCR2eictaofGTpzJi/yQjhU0NW63e1KcLopX68F0QhbfHW
akk7eGcTyTdHDekdi0J2KgZJ4JO7qD/qJZ0BHkA2gc9g1f7COwJaTKQq91b+2/fJ
adb6H4h10kEPEMoWTcTBOc/u9lBc7633VPFSpetf4KLJpOo3Rw1w0zwsvCHivNVu
g/IaGsvx/+l7/+Avn8tukg0waSTvCUL/2cVbaatZIIXIRnGtnyF3C3TFMhurkhwI
oYrxovfXpRVJbSxnXzr/Q2Oe6HfECtXdR/H30ysGDlNGL0yJvjP4j4BsyeEzCgPj
Lh1fDzwOwJn7S51KqV2cHVUWB6Xlu3SHsOg7hcvf5mKBGj1dYZnBmLUTtsHAnHwh
Y8OT1PrA0wwhZOW3c5d75pF3bszdADn0BgqWI6g67hX+TkQbeSuyCkxI8rvplJ1J
5hDp/ZvSgjRVAKFq0qrjLO+dGmQaCUOHw1CiTiYeyiU5oyYkKlDUVo5LPtCCwkqN
yCSeEe3kP5lQHq35Kczx4bISPRged/zouLNzOR2tSlhHVpsMDXNv5Yw09ZohlQQ0
d5CKFkk8uLtnjTdGXARcotwUNLmL753Z8RiH5bJvPs8S5o0+LKU+HbUemJG2BDE8
fLXl3J5x4OW31wINTsKaLE66qkkHnEmC+uuN0QEbZfBqKQbTHTYWOLtA5/egbadT
j/B1m+KReeI3uhHbHGXf1cQDCH8E1Ie5ob+z1J49hoLM68dlmkKaE7vNH4kcNv5x
bKsBqJDOpRcnxRTyU1ohXA4suCxpfmCp3rDTW428gWogtblZZNCKEOXp/SfCPPXh
j/N36DXMrTg1q7riAX8tcU1jhXlhnfcy3QiTM1CvK1bp7pv4MJ3NF87jbC+4F9X4
vO1JDjF5rNynFLG5ovdUZe9gFijp/oEkPsk27QmAXRWmdRepRM8j1lzAj0aXN+7s
DCSt3SxiCMmgCeMsX/UMS11jDXOFOyvKAmW6+s3ucboD3If7c+F4Ms3Qw6iLcQnq
yGEUMuGwOBfDKw7Qld+dQgi1WLc+04CaHnQelAuBSQsNDKkPrUeXTnv9grJEHQmM
u09VTz7Yigteo2WS1jlw7hVewE3JR3Q3s1AGjeMEF680z144IIYpJ6t5Vs5tvQAp
ocizc6WpOv9UqbKgat99y1W2ApThp5OhEYBp5aTbDmYX4aIvGNil8vtCvsDzVSwC
QD2pyzE8WYujWefE578ufzqwNVhMa6/+q98e95L7bIC5PVNWAEcIXq7vbKQKNBUm
X00GvX+86tjAyWBvU803z8qboEaxFNA96jYDqI6jGaqbIO0gBFc/nW/+7Kx9MXWC
jnE80MBuhb51Dm2dJOITngFf4dL4HwaDsgiJmRgJfkhggXa/jluuxpUsw1+EwRip
T01Fdl/UainTJLko7iNkD2OXuad2GcLu3USuxxGNLvb8/6kReVDdZREWyJllAWsS
3Yxt2ieQA9OQYyf3DNabsTKGx0PujvGLdMD5ve8rb1dNkIoXZUtOTDA1yD73rc7G
BoQt7KOjPjYZSlMc2OpinORy97/vZB3f/wdCdIdgitsLFiaaEj9qhf108DS2Qb4E
zZ3/6CwRhRutsw8FxPpOyfJowvKb4564j0U/aRSdXZwUxH7w3j1GxgW8rYMcqOif
M+b2oxvVumJVxA/90WnF13rri7ZmsOQiviTB8EEcdSaGcXWnzTKQZyCffDPQBDF8
Mu2s6nlyf76iC5CEbv4BBx2rk0qUnvLFYKfM6p7l5Qf2OS4f7M0Z9KCAuNS2GgIi
+Rv37PyKOS3FXxFjPS7MfS+xahNfZnMGyFagPSSs4tJen6vhQGFq9LxV3pDCQl6F
cx18+ahuW7N+81Z7NWHlCWvDNeevUyeXWa7H0i5A3x1tevh6GLumZbOhbpOTTNet
lZy5q5I4o/ynfyo5nZA+ipExnt1J4a5/tVCCks96nV/H8WXHqXvh1dW0Vaqp2cRl
T0235uLX2CIY9Ue49cmVsWbSyVg7jHg/eBtcRDdcp9IFuQEj0Z30PT0qIk/nZxB2
5q4B/MJ1BkGmAfWDQU6z5znJzH09yUJm97TFnxVi+2K8GYiTVREao+8T2g4VNnK+
JdQvF6h0kxvTO2ejLU4tjy4iE5vA/ojaLmaKz8YY2RiOHrDEazB3fgYN2CYNZGSu
4bXwcd/DaiKADXp/ySR2n+F/1WK2bJ3HfNDtKLj4Ye5uy689LVMygjpXjx1uARyy
1T17a3+G2egK6ZAeyosMIeChqNfjWv3ju1YQTEY6ngybrq51yjXU9hAAjgabq/68
YQiXPwLGGEKThICJXQrwp6d7o7NxQhE2W2lTJ200LX0QhZ3QzFnIyV1fzNPMccO1
JIff9W+2sP+AziKaXsgJ/g8+SnkbZihBfOg5nyXkXpAnmQPeyuOFgpvyeuamA4UA
GhnKmwcWjDL+30L1wgd+747VjiaIHZMagsuG06XyteAGfYMaX5mQO4cklajuyMr1
6cfJp1w2j2GjVAP8v0dAVRhls+B5fkKe+KMeWv3vUX14tIDJffTcn6WK8Ps2C/7H
SxNydklDeiiV3ez5LViDHUV+oEYwSiAtgQJVsH47vSkFzOOhNwvwoiw0EBz8hoDV
Ollb4fDcSDHZjJx8UvlMAjjLJeG64An1mgvrzrLrx3eiLf2CJ8KvyjaOLHZ8AtgT
llGshxwACbIhbn6XhtFRaHBXMfBgeQU8VRpwvM7UByvMLfU2XuyoN+CVjU64QUr0
WDv1pHxYPRCKdK2b2sVw3E4vfHh9zyGhJ7Wy/4z0DTtfLJi4IQMV74VYCEQZMgoK
JsDdQl7u7oav+R4OmT9JOPnPoTZeALffDJdhqQkl8auORLlfkDlaL5kMaB1wz05H
UBli/O/JPvF0lTv3xeUYszg3nGPHc97AWfEZH+WHBlC8N1XfiRe1SafI77YjoJXT
B7WX/4OKZGhAyL0lBTYMmLMTZiz8KmDMa7CYGWoW8WcteCniSh4Uv+lcxhkjTs8L
6gk91pBsNnfuWvLvY7Mas3E4hV5JbJp0yxD32m1BptK9uSd9myqMncV6MpWjv/EB
L0Xrx5ICHDN4EB6+LKkAW6GBb5rAltwujxl0cZUxqkg9hGeGQj4DnXCR4ey2A8AU
8P9a/lb2Nd2rjArIr3XGPRYsioqyYjCnUSSz0uSlTH59SJ+sOK1Bop5RfpJN5oj8
oSJhOmRgVnKYsq7X2GcM0wxWEibc51Ic0w+TK9kGz9HJ/TYzaXU+7t3rCPrvuEtZ
XacycBmFyKhoIepKBaTU0Tn0J7udhEfO0lgWl/6D4JxBKquFG8nWNJ8J7TmbZLn7
gklqIykukvZeg7yJzqeieRbvtvZ87FXwvffm3WQmJA21CjvubeAvXreDuQDbGpLN
FpnqSlp/IfPJeQQ5UTh0zssxtQ9nV1THxqgppMXsbU70khfA1y0gCqnScDZCcmyD
pPhvDEMaNonbboIOdmvknxQ4iF0ZCHrdLtupJ5wF+u4A1UfHpUp3crXWbtzTs+Nk
nqZc0jgzY+QwpABhELgVPCwV1E1xrKoEUon85kMfnlJpD4WG2XPqafu63eaA5N0F
s1cahdoqZsDhwUxyTnU/lsP3mqv/V+7HkbeS+mnyrgC4h1vxtGVfrRlYhNZWCFvQ
uKjYcKAOojgv9RTM8vTC7e1dItoHL4lBf7i7C6p3nWwxu+kEI6fkhY2ybxvXmp3b
mvFmWIvNdVrfeRCr2jIoxaG2HRdhN4zco+9cnHS1mU7Xg+Dovif7TDQFwNqI2ETt
LOH00pSnCl+y2+C9c+phoyIIfFNbbkSOqafg7mRAe8KJY8JbNGoTe8NKiUbXP7l4
XbOXCf0er7A9gGG7itvbb/SLuXsBZhqCTXq946H2HRA5lLnSUceyyth1ZYUIdOBh
pKeZ+AbS6IwupX+iNvDPTabQbizuHN1GJsk/vbdMeNaVy1i/NpbqJqmd4OrmanT8
GAFvxaeOaE9o4Z0jfXojtiF8+h4/L/Mo1e4LUZjqQi8//hhADwQLEI4MUYQ+hjLk
FRUi1w//u1TaStwqAyRRbj/kdRoBf4uWeWMN2K8FynnYcxG25RXsBiJeiyxRLDHm
tam+1foxvBB951CkEjBu8w0aganB6PKqJX5L7b3/RHhbWPbEAeVaepcbUA7TEnWg
UAOoQ+nmyyyrfxExxS2Vc0BiQPkvv2Fyclsj6iT+q83xI+zU5Aq1ld9d3QcAKwlo
hxVLYvJ2R+3H+Dy70bfVJIT6WzVnzfN965AuUzEcjK+dnk/CimC4wUXneQ7szZKm
ACG+upgGbGRgzNSD86SirfGLSkC2WsiibASQ/Q1XNDH8wesUeLDoof1Wj5sg76UR
4EbtkBZeOveyrC/HTyRtJnFL4ntqaQkkU7oK00MZjiYbQ6yi9P8yj35yITYGca2F
sTW8CKDA2pzESkycOc6T7+c4S10rKhbYivhKmPrfLPxmi2fX5WViSVHfgVGTvi7V
0K41qnmnwMOYys1v+0gZMJpR5w4VWLbeI0gVPDpNW2LVbZH94UIA1ITQeNGHqr7S
m8AvhxVjr7/9/OG9TKhlustjtZxJlugZB7WFbEvA8Qu+OFWhVALGO75q4M7Uc+50
W9ghs77lQAmvtQb9feBE2B7RDixI8puu7SHvp6Za979O1P/oJEg6FzFZyRvtSS8M
doigfVmKq71LHc2OsGVY6cqBiuXiklrZkZWa9WeEO/yCsSrN2f2WTQJrd2Yn5+hg
4G+iw0sMuWCDcorA1s+8J0in/qDBoqzJWu7oxQeER5RHwAM7mnMGJlr3VSrAA7hJ
WChQV0ofcSFaIwLIkDcTz9+w0BfRb4eeJpfyJw3b01yf+FbqmSRi6Mb9l25VC4M5
MXr5gFhE5PcOfAidLlvVc3iA2F/ZicvYvvEIpF5DFPqk1VVUo+7Kyoaz0YayQC6E
gHCG4h4PpYcM0hYomlFz+e9r8unLXlROfrPJTK6+dJHmFP0Cr50lkoNykag6vZjy
qtyMxhrDYcJYIm3mAAQSGa1I3runtFR1mZILHNG+nsCpcfjdAPxUa9cfJ2k7jiH+
ud2N3EdUy5UTScbWN/mtOOYMSEyKL+DkW5sUHMEAOWti9nOIopgPzG3oohxQub48
Geq1QtkIzHxhlqdsLIcd+Rjp+GhuBTjvmh7sSYScUeanzM+hY8cHvJyY+QgJqoDA
eGBj5AjNxNSi0S8hNKK3FSEKqH8Das4uL7v3FMVsJDeo3p8V0LOoUddnPbjfE35h
XDlb0PDRlSTPSwjMf7GmbKDKK6/k+Qy8bNiEaviVqVo4EocbdPVllI/O9HDwCobC
2gUTlKaY8VYkcBXwndPtqnJpAluw4FYtyH7SHJJU/x4/F0h7dL51TqwbTJE6dUmm
DrtbtcjHAc5sXaG9msWM+4rgeq7pR3cb4UgZQt779NbxZugLOee0W0OpD0F9BIg9
b9omZsrRjulbrSEQAJSpImndWRgGC1KerYn35sXd/jZkdL1FYz5WpMzZL7d+iNdW
4d7HU1UvmWKf5ChWeurehQp+sU59rzggKPZDqUVhn3XPLW1DZmwlOo9VPxfRqT0h
ySzUnqDXckaGxP72JQJnIKqnydkFZ6IM+dqNpSANHcC5ypfHwsiQJ1T8nzQpAara
lfnShSviH5GHf40mqQ5DzYMK0X1pL9Kq9xvr/EJbaMrAcMTZvOnDeDWJNL9XaT57
flxQh1fNYGQ8t4TjIp1eI4fkjlPbaU4hWc4aqv7+Ktepr1Y2oke6SLju2CAbmbQo
cdoaZXsPkbkf+9VVqu30U2FW8/uhStiPym2NalqBI1AzAHnH5jKdQPbZeFn2nTwG
BBi870NeZVq0nXkgGxahWqpllzuvousS42XEvOn8ajUJECvPnhw12vSOH4X2FLrj
OuZ33IWO1HrRrH7+O1Oq9sQiT7Ila8fs2OdqjKXIMbXksmoMI0PRVO4/D7Cm95ra
5VXLeTPOOgrDl8pZLKipuAhcF8GI1Xkj4hBNEUP0eIg1t2w6YInbBXEh3aln4pS9
OMJuP98jeLhPZOTLzvai+zoXl57wjP6S8Ok3AvDpfw5Fok/1FLXFdIXukk7IJbXg
skZdkPVje37hwTm5bnDtlfeXKH+JMaQNYPdBCAin3szPhK9dk5mWk5NA+LcePjRd
JIoWv08+xj6xbpSNyjp/Zw0ORD+YVXjihKzccOoPQrmpPstxJyBE0vwwUmB83t2t
iNji1ePuwaob48XEe+2VDPpaPawnAcqLh+lBV2hY3i1Y/UuJVgaeMhN6bdyWWrnd
GPaBGO4GUPd5g9qpk27lTr88UopMj1lNU2EC3KkPekJtOnEVgHgNUhdjmH8ykwKv
6L3UxwZSsF6pRreb1AM+4vxZo+zhmtJNCiG0Ovpn8x7zw25e/j94OxQuJjmTK07M
T6lHMIiNIdssLdUualDiBbxfC3PfTJ6iFiWJEY49eVF5/DAEk+urKS+dVshcW9yn
ckxTEpZH7JvA3T/BVfSF7NDyZ3TZMwhzV1+7Q8fvqIsS2buKOyZKBi+6+LsFwa0I
ELrAUKeMUENqVCUb/kEVwOMTaQJLwCXG4fzkL6CSI808NH/PGmW4kVZvSP8X7/bO
o5BLODAuLkda97boYrNwZaeWw3KXiZRgIJl09wztoEIv5740/t35CfyJ2bI2mkQz
gmJSqKWYSuN9UvxtfCN635qNoBDPgMZ+kyPOmXeSjBMd2sayzDEUMbn9By22t+U7
Kxoe26ApLUZS77D8RDp6ppeyNrnKvBg2yt16z/10f+axPzdV9LjWJ2RglZO79qIM
4y1aj5Nt9qypFDjvdWX6Ws41V4haWMqM4XgYYchWGcFFchh48j+0nT3vZk9DxVij
YLArJfY+ClTd8rQpCWHlMhQRJZRWyeFfvq07/HNunDnRFvnWseoayRXy7GQxeLn0
aFaggvUI3Qh9OMb8Y8zAiTxTY/ja4BhKUnTEhWCkVe9vJ39tBaDzraOCnf4s/Qj2
N3UxupUtGs8bEX6EPLNDPfUUnIB7y7shFifZykk5W63ovyDtAulrLk1gLDSETH1X
NoBh4JJlkvFo6ctzeQQ9VQ6NLFGkabyoZ+lcj/ggk9YeRj4/LPTn41hcDIv2+5e3
P14KIbd4b97az0FUyvk9bPpPzu5Dc/EckoecfLUeLqJSQUcqVRH2yUUP3fyMCGA5
O6jZJVBcy905B1zIlqogNh7mn0NYGd7mTPz/8zbonVPWiubWPIVOuFlEMM4YsthJ
nz+MiJqptA/tRjORepGW3ks+kT5ODVYgt1CB8aKtJ4gGC/7ppXyruQyA/4ijV2y0
h+wS0uYc/3uYNihlBgbLfjYaqjyzvNxf6NrVDGttNb7dbfwImhNkoflCV+PrbUdo
BdDcp93gUT+j1qfmOaFg3T0HTBj9LsT9nADJ+7OLpHfsxj0i64Oghad5OTiRLy0Y
L4GM6Zzk7qE9ynXwnaqddmUKHNZ4+z/DlL6l93OCQgI0r2pDOhWKfn1wDeQc/Rae
ypgvd5obXnKm8hNOhHfRs6rjyMK/ZDYzKbFBM3DM3Yc7R715ma0BVrPkIRdE7Kwu
ReyJ9dt7/SAel8kWClyd3L90FMV+ceDJo8mTEUJh3sDuptLnG2SBQWUC12x6xdvp
C2CZI1/WJuQJ8Am1ch/q5TvovsTKSxz1MCGOT+VBiFJ2e9jElILWWNaR17fa9Goq
9Lmp1z4aZ4yrTu1w+ltv00H++NoH+hBDf6PVPrGqwfNqVZPTk3jqMmb8WzS68zuu
VckZUEgIfERp3dbJsdJh61p1/TUmnp9YNqEWWjyfGqW3OevKuKtEvfEdDBKdGtLB
L2MiSOQ+PJbjzd+YQKixZLFPnoJPQOHSjVXHmuovNLzjOeUs4YAEZY0UkF1LMYXJ
SumMoaVzbVQsb/WqhOHMXrAYVVBGwfoWYkKd31yMP8+pSaq+FnBr9lCa5/G9dmV+
UMs3L4F3HDgVRDaFMEgag+6adJIsbNfXtkYd5mHF/+czq7kKn953FPxaoBsTjlJc
s/UwXj26lgpWTp1LInmECTeM0tD/Y9cmNGxxa/mIWD/aBL8VOWWNRMWYX69Pvhm3
EKdKzcdivhcvsDXP9kMwwwpglNb2c0Oz+Ek7fe/btFMuQ5hLnVK0mJ1p6RssntpF
7Vrw/kCHuCyAJRXXw8yv3p4P8HcoVEGlEvB/zcnx+8yQKB55IsQoHaO5ZY8T4nd7
nDNR6I+30Wa6XEtjpHEOxo2qJ33GR3/6zrPxRNWuU8VyQ0y/P0KNDprIh358ihaa
new3eFnJqXqJgEUppSWJFJ2FIyV6muwQMcnQ4LBdUJChN3eoi4ChSXIbCTwJJmiU
L/q6aoC8HG4g9NSbeeu7oJO2e17xfjUKGr+fs4eLNhQShBBVbjLsIf04Gbop9TE0
lN2mdTeUIS4Uh+CwmhULTSKdAWPXqIFie9L47Fo87QzHA4+AM69y/ZO9yy6ARhk4
7KMIdBmhZk0U2x4U5hC4d2f8Gv4V8jakG8X2bNfCF3LuCiwlL/Qizl8rIO59/H+r
FHzSBauSXR/wgtjxGEZgv/xW79E+QktbImaPfnfqzAqBzYbTKLyScCZ7QjDN+cqe
lAEpZVzKrysgd480WhpLMRBcyeY/3DtRmi+pldMAKA33CGKq02L3leoJVG8kW30i
EmIzD1XP6Y2e+PaRZ9n6LwwM9Wg3GHNnkKfDkluu5qbh9FL/frBXlprfzw9TOvgu
4MBsu/2btDbcMhPFJ7Ohum2Ty6x6cTpC0jtT/20MaQggtWyeti5E8AguCphbdFLA
aAyyGy8M3MKgQsd/nSEHHs3kB0rzJ/kuSg9b56NgmTQEw829zwUkAMPVfNL69UH6
z+LfpgzYpf/ezOMx2MITtNrdPrbcp9sH5ufqk9u9gWSfvyb0bgsng1a/LLYaMeH7
Y5PvjuqZLL56yYgpapXilw==
`protect END_PROTECTED
