library verilog;
use verilog.vl_types.all;
entity main_fsm_vlg_vec_tst is
end main_fsm_vlg_vec_tst;
