`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uJDsSm+sdmcYeaqQVL4YUFPR7ltOccBViKr+T8/ydxnjAoeyAK7jw6KbneIizmEn
nkQnWhGfdHuSLVsQzKJHv9w7A2zCEglK12JyMAqvQKpi0TbZfXf/b92Qv7XtSSPO
gn0iyvkkOVLcUUPV/XWkdZh8ff3M57V5Eg8Y9xbOSOmUXwv2z4NxdbIgu+4eKyBV
/i3UFdhGoa5ZOfkURxHw11q5yKly7iAOtUAbVKGDs7ImITsauKOxPZPxc8VdYNYo
0X/niw4NUvCWDc50HIE4/PIq6tnjWrhP41403bANs7k2LvUeoDl0KGgrDnbhcwuE
OZHwddVNhQb9Rins+sdJ7V41XfGdQ7Av38oNVy/wf5P3ZBUDwRQmEqcKhoJ71c/L
9inb2njOI3MupU2TjHT9sdmwvOtrkBKtEKirN+XDn5aGTDGpdQNT3GMEmxwtswMT
22wb0olyHvNNGRG4Gw+w7XU0ws948wbVW/vu+O+JslLFDQQFqTEKny843P5hJieR
1Q14NMLUiku0tz9B4FZmEyL7Df2XOFxcgQOTXEqdgFEmslbA3mS2mxjueQO38aBm
wSCSSJKsdXbba9kyhFabsEKHRFMACe79vAUQEzh51cCsp1FaSZCmNm34VDvdUZv0
oU7cWqJw+2/5TF9HOpMGuLUsS9IXfXKrHzc9PJuyjCo+NQxFiCJ1b7vhS4Nuym6T
aGdyxBFoI1Y+YGbdraPM6jWKdBkdszmB5xK9TzX0lbGdP8dPzT0DimmcP9BGzFgf
NPNG6hS90LD1OGSXqxX2ip2lTO4TeHceK5SxEzBKrPy8wMWA6hw+U5Ny98yPfVmQ
tAEZ3fpT5xHp9M0jT41Ooxt9XRms4KBGCqJ6uMtrz8ufXmHs/h14QSR8Vk4WE1eU
m28G7LXAyZhx4wLAdF8fjvL8G5s1nn+zCP/B3sKMCuwH/Avco5IyU0VUBtwX5mFF
FBD88Nn0V3AbznGoG8td1Dt6wti1KKp241Bzi+rG0TVy4HdGwTReeol5FM8HZZrG
fX+NR7zwh62Hj3pRBN5a0bV+q+cfr75fQC1VrzDqmTsW3WNHr2sDtbsJO+hBe86p
biobXPWpFbxiHeIaotx5LP1nR+s9i0FH+Z5ReIRjF/gZcB7FslQuccu8K9tTW9fS
0knm62ixU26tzmhqOEP5u3nQZBHoyRaxrQSiQT3O4sfoUrQTtueXNc4RqRYZkxRp
iJ4f7T5X8Z1yn2Dwbsz2vf/rPGQUy3Bo5GwvjXzr0ZUyPW6rPv6jRts0JWMum3Oz
b6ruFBwwOIPUJuoeEZLXChXQh6v9vbjsJxUzF7Upmy97rd2/5xlhBbXXX5n8SZm0
0iXSQkSRUO386S8hJDrzy2GcRJtiEwPrHjYtFwjLm31Ug3lTaG/HqjKHtMGbcKUG
mMb8r2MY+3U04CR0XN91TnK4Hvaz/G5JTag9EJnBf1gzcu62hpek2OzRhTJhO55R
EGydmtdGnF3I+AxQlFp8JcciKOBR+BSi0UqNjG5i6WV/WZnOY+P9ncU2DgeVhL7U
8alQwR7SCn98QyQNGXLuQV38zE8n5xo6xB2nz7GwcQ0EiRQ0VIKdsLvBCZgofzBu
Y8S+GSKbXoR/iweYoQHm4Ew8LXLx6II0fhuuiwK9H5/R1SRFixi4dBAXKU9A9rfD
8MLC0gW/TpokvEwm619mOTqSg3og1pnndpAVjd672DA5s1dJudBN2yimnhZnKQ+m
+3a1Kcl73bHPwZoqllqN083k+JZegqRLHAgqR0V+uweIwj+uL1VbGsse47nkzIYd
GvxGPeffmJdwSf2juqh6V//D3wCiCByOcbYDYBFMBbkMIwyVq4HO8VHtlOu6AACj
si7fIhLJPLsA9HnY4QGzsQYnGTBIhxRvJzhw/0mjjsYoWmYtGbio3WjePLziiP2q
WtIItzMMi5NqbodVbFLafvl/miAj9T0I5/rQE03mDNZsd3WbqyLsP5TBOuOyNir7
5Tb+vNLu6nrGzbCUpWfx2gKuESHIj702mqt3Ds+TuP206fU9B9o9tIk6oN3g2MmL
JQ7omeDTC3HYxmDN99JzzuTxs5onbd15KMpSXEzHRVq1xbtLSVb+jN4++YStwV1g
YsoNBEGRkpLEK8DCq6YB3yi7SwyXYv5i3+0Aln53MCO+v+F0DQ5R9gZ5e7Ipj1NA
sIr/2Gb5MTCafP1ZXeqx0mjoXN709xkVd1bkwG8HffaYU6HZbTL8zqhpp8KGXS8l
UPS4GiwcwBGJ5npWJIMFDe8o+WNi7uYW4HvNIy31Vi9uiy3S78OfwmvKU9lOfOD3
S+3n9sNpIC5mr6c6V5N5Grow7xo6vLgeogLMCRomhV/A3kod+P8iwBFATrjE4ynh
KvP2Wzc5qVqEJLhng/FR5en1ZFVxuwsGkPYPugviQWyYCSWV2z2ofazCKLw/70/1
9f2NY0Er1vfn19hFf/fQiXrMCducjIUnxJtKvx+WM/guKnXnI8SRCL8+1TnZ3mNx
xrisb7uV+qya6fFTGm4E10OYE1e64G+lot9yRKOtCbizxG2OcERBD0FAJmMHidWt
p1/tIrle+xqM0YQB3jKvipzaM8tSShCz8CjeOGrfBX8hdbYdoFfKc4OdhjUgNkWQ
2i1/xzgmf4M8FJztGzsM9WM9q/l3+lu+4H2DDAjIRuqEDcF53s2/17cOt6FA4R4M
WBM67/u6goWiLGvzqSx1hToJScITLSCaAUAD+mpllJ6Rd8eOigR2seSbx4KKLhF+
O9HIVAiHdcV5eV/Fd8npHhYGVbK2NFUxV8pAtcIasI47VDmmBjUDhDsWnDk5x7Ws
RzNSC52mseiYV1tw8MxlsuiJxr33ucPLeWZlPbpqci0=
`protect END_PROTECTED
