`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AWJKar0SJcbQ7ClqMyVhMMTuidnsFsR9vFdIcEqn9XHrDs1dfn+1IN47xgSqLr54
ne3jlqHwEJMDMnmrkEDs24Xf+ZZ6/pWpYYofYV8uTdOYRLHNQWG/RiDyFaWOmxDf
KDKWRObTUNeY1HrO0vefdgolfj58WeYtvAGKRyiGSey70fGV1GPxgxTu7PgSOxeV
z+ohqoF+bvpyPns/lHnC/3ZyELl+FdQX4UT1ezGn01S9EbSgQog2oxCrC2RTICl2
17JKB+hpH4VfwSMs1FPBdiEt4wOpELHKkLptiCO2NPJ1CM7UsJTXgToULAz5MlGd
AqySMzmjFmKT7jEkPulC7lWAATgwpD2hBfzhJ2/IHxIGolvFDispQpvrHWINMEI8
`protect END_PROTECTED
