`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
l/gsT40oskLn6Uv/Et8cKKsVTY7NBPAnOAN2oxGvw2CVhb+cMsdrToEEuRsfacne
W1DdSSzxi/03pJI7u2R//K7e0HevQTAB3RF9KClE/EwZs1xbYBgG9/ltduhIaeP4
KDUU62ayqSDxjjBrMYYypyDAgEIJQ2rgmhihmiAwDfubPq22s++8wN/PO3fXfz1s
2FqoLSFg7Sy7DTOcsaM+eACJJn3ITC59CELG0jJTuXJfhtwMC7F4DWR7X1tdnrBa
95nDpV+ZeazZe+i30XvFB9ROYEOYv70mfzy5GwoA/4w8gLAedHPUkZ56pb61cBdY
n3pX+rvF3k7d5f+JBvL0dgaI29Q9LZmhKtfBrNNLtmdhDcNCqRqck2WxWxCEA0Ip
hSCiY1pcU8/KjzyTr8PzsU/VT4Wlfeg+XzPfu7ENP/jeBO5zDGW+3OBuIb6RzwwD
NWEykx6tsgWVSh6uS4Tj9A8K0HYg7D1Scq1FCZpDQuaMoN21xOnPD2SmFm8AKxtj
xolp/Y3bzYTAtDA3opaxmckKxIhsySvVovWReSK1ubUcKo34bIJMeNp7yRbxJK7V
b5TiZ6wcMizOl97gyqpGjr0Y1vi+lTgCk3fcc6G/CoTbNo/319S7GE0Q5hcxfLZl
dgtHmkGF9OcI6twM4V+iF1j7IpY63MIRvYh1COC1yPzdf1aiA1vZsKoxY/wl7kjE
TtfKKIWYqekg9BVtNN578vmHBeRnf7TSzs5hO0iR0rTJTIYwVesnL0s+lYA2mLa5
UGQFaDxi9fYMqFSRBE8pTA6kXR/742GZ0oXT5WCelx/2LxsLG12DIEl0ZdhAFGyz
69gIVig9KI4VMhVJrn2HXqyVsEUypf5xUzTEnID+B2fc4QYlvKZv2ZksOrhMk3xs
YOsPSbESWhz/MPh2Azi07XLxOmaJ3Prei2biDgAhkriH3JkNenA60vmyko+3QXvM
M/6p1/BY6yN9pFtlP8bkQfz0fHCRUPEA95/WEclaPaF6GKWn4yOLNfSGX4EIq20q
FyiIXYqIlObcdzaVcu99KXiWP8AzGDgfe6rqkDZNc8vso1c6qhwriZfEWsuM8Qpj
O7j7RjofXgGvDX9/GqwgLMIy+hJPfYqQpSp+tzBYdk4nYrLdI15BVYbnlaBNTu5e
gU9gSLaLFHzlNj60yLGWmYrsI2ZJ/wVGSrhpnXFE8CkoRpKoY3ADH0djQm3sQbQO
3lY2hf9RfSB1nPMMl21Ix6pXgUSBZ0+RHhua/KAcxZEVc8n3nICJTYgpqjhxogiW
EO2P1fAT9IpktTsSLORbPBOQZPXBcsWp7Kk5kEB+Is3bhdS9biIaTvTKlhrpHFpO
XcByH/nSpjFU6ekF0uTaQMbI1rdACB/RpWTRTQVp4VjKF0SNSAejGZN/EOwCA1JM
JCoilnCUBOy+/tZ9MaGBmvzjvdbSc7Oc1Upjg2+fyJ8oC18uabhSHlrtsj1oQUTS
ARxqgwEvCAHISnkvLoePJleQlU35cPQ3fZyg+LuKFH1PM03FH8jPiina6FcWTMeE
tpFKixhX1w9lfnjbpA2+WhI40Z8agDhEg2qKLx82ykxI0SCNCO8Ll/rHd473BfHJ
R6d4VtzSNH1xozqpnA/j2X0JLiWSkYIGCaRxkUvCXEEGv5OgPij3x4JXU44bWE9Y
CvV/augjRV0HiRWogDzzYdsFW5doNkVzgX0k+2nmCnT1AzpEP5FJ0o23wk43Mk0m
pl0vn2bymrChUrCV/NXMPoF+ETJ8G11gp/baCmINAtsXFJhtOQETDrjzL+W68qom
hZm6lPngh403IbbtYq2ZpqnE09S+31+8adnpgnfArfRsDm9wykpd+uZulO4G2yd8
zFVI9r0MC9V80tGN2O8RjHEfXRTg9VZGNYiUQw170rcKpylTOcf9KHQGu4yapHKx
yPZi3FXGWrDsVfNmk8GPP6JAEdMLVCT71V2q7jJPE1UI8IP6sOhC3lXCCW0nU1n4
of6yDGOj/sVxRO+fIuj3EWAGGv2rx3UOnaXb1bQMTFiBIP6NUY8+Vk+/9Dz42UqT
/hk1aSWJah1w09CpNBklCpfkEaUceMy81PnKo+moifARBS2CRsZHY5eYzfmecn5D
9+JR9ny2dL5yNw52FpN6Br0TNIvl9YKgm2H9ApOGPi4378LR9/ka0PmJbKUZ7TaM
3h/0KmQhEu4eEVhWoL6GZwMa1NP5NxkKmBssT1qeYzT8H8X2X517r04/77dfBkL6
7vXU7oqwzIdfSROoKrbMLV6w9RrkS2Vdskn4v0knM2Hqsr3kWVoNhpQM3YC3KpAP
iztdU4ZUDHGwJQVub4PwCnqwtxYicitDXXvqMQHMDpbq0ZOBf2aqvfWQqaxHHWyb
8ksr6z++dJ3VyDI0HlnPGSr7i8vcGIMVLHjjw5dHNQnAHIOqT/N/fuPiAHrzCH7A
yZAvD5z2oQOIrELys+g7NgGYHonWjDmqV3u18d0E3Us2buVv5n2i2827mI+mW2lA
s20NrtZmg667ZrhVYY19Qzqr32PTLOfmCXmAtfA8BXbbtEI72zJNkxsf2ZCbVhah
yToiNDlFAveBlZZTx9NKKQB3cUrJjS/oqPbSWWZIQNLJp5ULBXTCXwhk0D/D3xPz
UO0uH7Zk7MSLXG2y0/WrmSHlIXlyQre1jBV8QnDWCLL5dhP8V15erlUzE3SccNjl
7JvAxM8DaOn+Yh/hxDgcsHT7IGh1Qn8Nd9P2QI5XfKkpsb/49e2FxswXp9lY+dU7
koPYHs78A1IvGqC4dM9ibCVAZze6YpO14LUnib/Tx8ZauLorOmA7e2VVXV30JsLY
2+L6AjYI+ajwqbALghnNCiy7nXsfcpf+lSec7BTpcKLN/ngVi4TxsmCECZGOF7wb
o6+cXG4XuBtEzQy4hxM9RQiFyARSIGuz5mYFg9c4U4WxKsvMHF0EeZRl4jXqA+CY
4A1wzpEdtaRoRFOxHWIc2vCd3gJsRVxP6Uoe+Fu6bwqyQJvDcazW183X3kzsr7rK
9pEJsqjQju617q031vpOu82061677OLyPzZz1veU4PLo6TExGL9SIz/IM8HCtYkv
/mUsha57IymwMYj9wE0Oh/Kx923015MkiUSRvZIOtEN28tM/sSEcJ+eNOG3FJU4W
jry0rN8209ZVtF0dWz02ud60wcJEyTBLJTXAZi/1k+omH4cg5oBJjoWosD1/StSB
9/Th7I3dxI/2zVdgBDx2Yw==
`protect END_PROTECTED
