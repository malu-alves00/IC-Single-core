`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tjvvNnM7Cf0zMLKuno76jlXLVGGZwNYYVj2Ypz+UB/ggQnYOAItbmR4LRPXI9Z7j
31s779XKXuDWNXsNfBL0/pcAjjHDUeLiowhnxSYU7X/oTngzZTvY2DS8N1INW5B8
Gc2ZK/6zqePp642HCvpKD+f/Yoa3qpdTzcF4aRghgQZ27MDCuDxipzaN4/F35IEq
bPuE1ztDRPpRBbtyZH+sJzzJNx6ovsqFFFHQ48ETiMPC8iVPvhQGoGOJXU3tbYVX
k6TTis1D3UaE9VBc5pZ9sCM085iVfPy9u8CxotwOZ7QEbtzTPTa1dLLA6w9XV1Rf
o7tKg83Hgq8GhikKB1bmfaXJ5THeTejP9fC4PX6jOfEaMQ9vOjUBUQTlYBb77P4J
HvYbwiPsG6kP7hxMfyLj7/2M30RDRREw2bN9D6APXnXW1fP6uXkDaEkRovCqdSZR
2CXO+Ah5ePSiBZZK4dkQVYGVyWKfUkElifIoMWjt1YNUyIi8Lk/mqF225XkkjRlB
O2mK7XVa/3YSzkFTYOrgZDqnkb6g5eNdKD3qCz7V7UKFGZoSlz+rSr6fF/OZoDcm
p9EdBlrBcbsWy7WMVbk5Z6V+F/Tl/gURg0XY+Rw6iuDDAxZfP1bFsgiPA+nAoyJT
sDnuCJQUA8/yCyMgyxtd5yQy8nKjK9WzQ/Nq3rsXkCVZKVQxq2kb83V/D89VIAXd
KncLLdr/5My5Gff6aj0jEPdxOc1dGVNaYbXJmuxPbkVCJlM6Koun4dpBfYCxTN55
QGClYloJmBqS5GDu1+r+mfJH2HJ+vn0ExFOKV4T36Ekh9FLZITOeoBIww+LCk+ly
3PLaYskXmp6kS3x8UTB/3ZPOyNouGyzF8zOueEikpVoPd1wFELuVB2J/iakwgUVx
R6dwb8Say0w41fV364K84N1Oe3rP0EnY2yRxnVwtegCoIXUpHBdXuBK/ng8nWJL4
Ebq1eZBgw5aQD31RV/jET65HiXTd8qjbjpoipaRUFWHvO72uSjE8VRMafYeYhEys
Fc9w0kidgOpFwwsv+8BWGkcGedoh0Ro0hRexl7U1SsWPNvfqB94T5lb0//z38Xt5
iCf8tcGZsmdXuV2wv3IowqaXpUyc64t3sdlCuFCeYdoMVijuQfNhkRPANr0DC9As
EezekiMcqaAZQcQJu16qJ+s5Rs05NjWY2Rir7x53X+GeuvMGeJzsK15ByPhU/ETy
LggCY27u4U96InYzaQBhfcD5lKfiDpMN5Gw14KDsGx39KwAX9UpZvAq8oNJn2cqL
puEHnBMhSUSit++prRpCHXhhBfXiFH2pAeA7z5fdE6RJM/aVqshHRBKbcixUc8Lk
l8cPHxj7cYOue2rM8ZPgdsPq3FFMLfDQdz2RF9LCdm6j5qwN1asWJ6N1MFboq/ed
75mONLqOP0W7eGB3tAiRqpH0wV/8XlYcYsiRAIvZygLEw6smgPS1fa2bi8G21txH
5R3Xlx3HNRzOO77OnSkE7hhq2txbmukzhWuluGCv6PPOAxSezgBz5Gkh4JGLi/pW
6aSkuhaUWwzi1y5gNBhP4e01fDrZnITpnAxJWwttmm477Z28OqR7/4TA+3EcSN3r
YUt/lmh9tsQ894lQYpt5xHsIJG5jnGnLFyJc2gHW5zoAuXJGHFzrpXbxSYyKEqjP
RmA41DQ2UwKXTQurqB2GnJaijVEpuvyZEHOXunpV2tJPWHq/ckHG7ZWfusL4u3Ar
2mbS1kjVlEM1MLMY2NzdIy92JdWw8SK25c0C6mNeKlh+YucT+Du5gTU06GtHM2sE
h/oeEwyRJ8hDKphjQnrTuz5wsbtV4pwAQ84EwhiyDiBrZf1LJx29e3xhNlrSbvGb
dbSYrfPrJsg2j7P0YIu+z+jwJojL3LnNBGj77wZu2hw6XMzeg8YjSfHqLA9I2Hp7
XrbW1u8kxOcgBLP5k5Lz55URKVz6LD3NVnak830Au6V//UjEIc37qoEVojtQGnQD
x6eifVZRTgslbbQOg0Erv8O2h6K0rjkWGWwAN2MdxRlHEPT178/w7zxc7M2RVyfS
Uo21gb/75Nw1cGxxje4jU6jCAuCodLZpluBI1O2/Hg2aXQmT2xoADgKnJpPbsRJk
c1PVLffVjHHlp5EYCPvPkDnUg1D3OVkKNGf4ysvmiUp+efodH38GNbBFwzMyZAYr
2S9rh850tE7n6uHpmGLUEQkly4QiMLHIa+rSpKMyp8Qz1SEYJvA4AP39+qfnhCDK
BjlBJjGRITPcvtUoUSVyBpiVzXBewlNtfYqoKaNoNUgxXW4v9RNhmrqrQF3Mi6Xs
xNnQCJueLfKV41TSFphqKPsXy6ZXekbt1tTbE/guMR84qZFYZCPUIHWEtrrtdchu
VaBu/nLf6y1mI1SxSwG1CgGvO/vhvyTXz1bVQhmy5+11S+VVg7eGwcEkKMTysuxW
hy4O9wcI0qDkQdBQMsjkiFgy0PH4FAY4lzuGeoZ8UOXDHRYRFr3X5+xXFbxJrNrQ
WTrSGrHypr6IHLI4r1WXOuwPJO5ze810m928+0Hhzfugfh7a1RjI0HuADfncAlpi
BioMKT2IoOeFo6eM8SiPIArITSSiZEU+uS9oXt0VSk+tsUg2FWxnjYOjQJpAtHlm
XQuLY3uR1Xam1xpjCUYikJnEddvq3votyp3ZXmiFGrbQjDS3YCiV13reY1lOeZqs
6e3mxPGQyjInEy5te0NdLBUtIo6sv7rpZyYvXGKTIpNAOipN+zp6kd8p82U+tUXy
zF/YJyNHEF1UW3VXPb2FH0rBkh01WAWkSQMdweqSMwWcVQCPneHzqyniVECYQXRq
lzcUlBmtwjanT1BfZUrwR0yyNlrOhgggjn5jo8Xh9ZK+3hXxt/bBpGUiiesMPlC6
FFxOwn80+rJkeY0bSd0rP+XlD6av2jhlIlrYvcE1Wk5ri7Nx2G1caPp2ozJfEUJs
WYM1cX8e2cnd6bh2wAmvTqaEJ8PSoIBQ+QRYCpC3fouA18jDaeKFV15jgrwMGmRK
3DL68Gmr6hACx4WEWa0rK5dw8fGeXVcSkZkzTCE+fHQvJJxcpzmj5HdtYqP3sYEL
z9hEnpANqdQWTiATSmGbKvavCsczg5mYpkpT87NuKbHLGBw7Vi2XNdvoL8w5F2Dh
ocYuryalo/PEz2Y8vFkRj75JxWpeX57rYSHT9/TqHK+FVYF27dKs1psY3UeTQv3v
zFtS1tc6Ea0leJJMJ1dqW+W8e/79A4O4/oL6/ELI7P/aLqY8B/Rft8enUCASvcZi
KMmBFJRXaY4E+H5bwKPQNgbBAAkn72QYg/E05w6nygKxY6MgQvE1I5zIB3aizDcg
bxBo2oYXgwbi4fakkaG/TbYjpvIKthHvxWFTrNP719qGV8DKjuuHc7j/Zc5DLwi5
gOVYkfP8s/uj7HUpfIrP2IpxDnFaJfmUUoT0sSfOYPzGFVfqz3pYdf52dx+rkrXm
spxhLxAV/xt3eEv6J98QY8lUCj7SejWv31xOvVfqfdmq6X65rlb+Pggr3uMKNU4Y
URMlIeYHxpTESouWtbzVdsXvsRxqRpnr2ir2WDIWKVdXukgXGUvSZ5UG3+f3foYl
VnXn3gP/PONdYopnjKzr5Fl3tnQba1fxJB+nGb5aFZcPvs/32yWisqjKN9cSiPBP
yohpmbeMit14d1ZANs+3wumG9HP4T8UVsHsMudqtH7D6B/BDTBDBiYd2LmqcdPXm
Zc0oRG5Y4Yy0wYKDQ/VsmFWRu6nvO/nb93OErJVrTo1J21Q9d2DpQ2K7nYFXHsXr
pIh6i5AnnqSoCxCJcCqU6Kj5VvD+lSvnqbvglafTWNQfYrunxOlAKPy3PInlrYHH
00g1ZK1wkZxrPuSQPjzm0MYBE94Xurc/p5utqc2Zibo7/gskGB4OCvhwHnTvqgSy
V5+NzQfk41/KObFQrGzhSDrfbFfwLx/RrzlL0tR7AYPB9QTynetoKE9afzZMXfIV
NgxNfD1qbCnyfIBncJaRIS+/6NVkEtRY12UTGdDFRS40SuT7NODBcFUUzf++ULMm
ayeRG+qlrDJIZ/F6hKdfHQSE4+wE2rl0ui3UBiqw/5BD95WauDPQHSAGu7TWkomo
pb0kGq7GNcsrjnS4F04tpqEZ/18qJjqXrYREbF8yYDWRoacQoaNYdgwuBapCiKpT
ejXPhJxYfHU7qDScyhQxT+l71QkUOED0ROIAU3zT9Gh3gnMX1g+z3DDcRme8x6Zz
SbxDRDWHQkW++44ls8HaI8hmKHV/C7u2JrSjMImsSRivH/5r6+KfX7FnNmDZpbgb
fANaDP1WEYXJjrfeSF5ZsiKSZt/WtIyFUFLpEz5nvN5s7vlt3kGVlvRS2xwVTBRt
YgMH/AcJZavV9VVc0t9RNSq1omrJGi7eesDxwLYkXLIWI6kDQ6VLboqGagx17C5A
IFUDTB86RuXxLgu2dVYKAwnUVvWOAivUJoL3pi6xmbYkwPzekM69eTXCtXpexFye
uYKzoze6rCH0aocbdGDa2AXs0xI2WdHIxoVB1d27pruClDD/nQrO/hVKRYaTWp32
3SV3YoJoDUOfdpsARV9u21XYzRKy/6EFKHdZJ0xc3arLCb9zRBqlK3b/wqXiTJXH
BkGLjSdPXhS32GYmroaKRTAAhObyMLxyTDazmp4VcAfO2op0fcAsuHSPvUyxPo3L
CBw495rMYv5Cxd0u0W/jIQWgF7TBjY3pirNHpGF5hP/S0Fi+lDoGFbAxLyZXGc2V
ZWzhifAYxLewdlCHo1Dxfi4bTmDpugLs/1xJM7aicFRRIZSe94Ovshc1KO04I8JH
5mPZJd7NlS+mppwaPF0adLN0whhBCxSylT3XbDsro6a96j+yWw6Up3HrXo7kt1IJ
Yy07/zNjZd+RTWxvd67q97FvPPaAA7HRqLoQUK7culaxMcDuoH74drJkBHCQ4wxm
/FEPodjKxYGCtp+bAhhwj5hraJelGrSfSMSlohdu/K4a/3/c0HsjeQOGo0d1jSht
05o6r4h1drD+RqsamC/kIjvd6xkuykbdc+H5IKD8N6HGvst3miHyIYWiS0EQGEX3
SBihHkOmuVNboaP4bjaRVVR/4K3gxZaJXwmzU5lwNrRMKCl3iAPi7gMVWLqIDkMP
EF8yAVZGpyRY1xxxaw75guSRSIp4XFDnDDsAA8TQiiKg+tc8CCpAVZdmg4ckTzvP
vpzIQapYcy4bPCXrlUFbJB3bM9VTs14jU1afWH10HNTRcEYZorAeZ5LbtN/LAuu/
c/bMo+iE+jkkoy65ZxuupP3WPY8p319nd6uiB4MSqgvRsUv8LURphR1YonUoXA2w
04pJ6iArI2DPTxp7BZJAWiCqjGyf2kbLFrhH+9galEE1wHKXwK4t/tH414ruqc+0
Vn5WG3QLV8d9kR5eitg7w6KV3r1NQFhANLZjFUn2IjocgihDsSjhwM0sv4IXch3I
z6bXTrKUIKuHbv2R7noV+cEqTyE+b+Dh/+VQpHw9Wb4Na+8LaELzmfErzrZTu4Kx
/uKvOxCDImT4pKgrN8VF4Lq1txNEL3b6KIts9MpIz1T4pUaToEU3jkKzgKExMkqm
E/8zR6DRjEYuuY0XJXDarJBqoxkG2Zo8j3KioEWp7yCvW0ecPsN5d5keN+2BTKfw
VwURL4CwmyoAVfflDhfQHo4qFFnawqoDnXV1o8y6Mj8H04yXqzCHVPHtMlBF540L
FdBjTzf3CBODaNoop/wWO4XXd77sQ01C6D7+QkT2PO9Yanf3hQOzRl9hWOsJ8X+3
vxej1yKAYRUSj4YGA+6QMLjnhuy+CgDVQpdp/07sqqPd1mMTt2NCvKGoN15MaSpA
GFCwjSYRawQGLSeq8fGncQc0FAQ4d0d5vO3LN5Cqct3ImXqC2uTOtWb9iN4UpHww
8C6PwRZCRauxXCu9sn+6CMA9/KecCBCaDSH8CcR+2PqGxE40UnXCk8PaWQsEFSCN
55s+N+o/wDFnqr0O9VNM3zmHIci3BM+059Diftb/yJv0Nd5AYvDwhDdk/4r9HAsO
EJmpucZgtwMZRhYADfn2wEwED9Mlvg7+3jsl0nHq3ZTUtYBR59Tt39R+Vjv0pC43
qsOMwrWHDqjm2X9w/VoCLcrzVfjOlE8wawlUu1YBxuAUY5+4/2w2D/uBp9b+fLuy
fCuzzKXgh5FYj3szurXvqLKw58kZ0JnX7YPoaQGW0+Zbf9l/QK8Cb24vs6SVQQkP
xnaVR6s1EXo2T2g2w+g39Xk46BwUfd4wsphfVlct1qp/qcsNa3o5kPwtQTV+8Kp+
gsOVVQ3zvEobMnmbTyaKYCz8eL2ddraYoCWJNKkIQ25NGEH4Goyy8pJ2xxR87Pbh
Lygc+a+siaMAuFBb8npCjH4L3FFkTlJpxn6LT4Fhs8jCK3nJ+2djw8IJ6mjwelW/
2edXv0CzRPN32hHrbhHoGK+t62sViP7Q+HC74gCM7bKpvUU4oxW1H4BuaJY5/jLC
5dvj/6y2f0SSkSavbbFlTM3yn/0C4KbFsoQPUwh0Iube5RI96cDXqSvtSs7XL1vR
BqN14BcjzAB1bQb0JMnc6OocQPetHyHXEO08xxNLxSW1xpHzemU25vC/qn4TQiwZ
RDJGRiNLqzVa/9mUI91fUZGgeSw67ux2KXyjjvqJ7/4oG+0eo3IfpFxrRjAWbVaG
/47yW1fGIsC1ZtSQNDvwS6lrebN3A2I7btASUmTouwkS0E+mM41Rx1tojNLaf3y5
h6fXa/ZuRXUzSYnC0f3AUIZxcENubQ7KhT5yCuBRtobSWHMKVWdcCfnkU4Zd/5fS
f0YdIBTW4QLjbDE701Yw73VhV+kxO0lGLXL6SHmo5p8gLUnfWMPUTTxp3SY0v5fU
qj2IdDdhuZQQaynp1WKzSzuVHlAJY43v4tZooxDicuKckRILfRKT15CvbpG31lA1
HbXRdiIzD6+etzUp5OLCmepAPdvT+BUuzYqoCp8zWM6SwkjP2aoBesAvIC7JLitZ
QGWd0qMnBZMI/50GB61WxswiOR5QBUz6D3a5a+zslzCIiS8RxYeEBEQ/orliaJ7x
I+6mC6VCX3BxtW8hNF9SUB8S5qVQVCBcwr3XJS4Ki6mxUfhcAPBHrV+XCSd8ff2j
u/FonNW3cgKakRUsI14jm3fsi7WGJ7/U5AOidMdefoU9pjHWddJxOnxoNQ25r/n2
pkQzX7IA2M3OTZOeUXKT0jcWjaaDQKND8g8/9qTS4krtNtc0uRE8FeeOcnDICEDY
BHFM7ORv5Nv5k2HvwzOKXKrq5m6zyHrRAeFt/9ccK9LHU4CaRuyHq4wEWlSMshDX
eQxx8HeaJDZa7VznZFeFNVxtn8Qc+6eCMn6AAW14kewB4SpQeUB+c9f/YDJAc3Rp
urMF7R9Ac71JftRo2wX8gJiggt+uz04BuVk+4PyIppLyV6SEzzA4eGDdG2V0IZpH
44AwfNjvPMcLdqlUm6BErKfIrUwLHRFh7upRMyn8GVAN31UW3SpqjW9kDFuWY5oq
yFyA5BxSmSvg8Kpj1EHgLq9mZmngPIcZE1oJzGKQIwAS2gB+Ii0z7DFcPEcqBXu5
jbmKp76eFvHpImhSXnTJH0O/4GnjTHO8K5HIyz/1qc4+g5RRUTBLkf0DB0SskBPL
IofHWzVUCc+n3puJSL7/s3LukGk7ma6/GFuaoUIU9NxiQJFj9bcjmlNsmVdyveCw
NH+22tV7d2b6+cNCc6EegLRidOoOnLBH26IOIKVk/JEVPGlUb/1HtTn+KZUYPL+n
2fW/8pWQkzAFzo490OGpSmEeh5fjYmzbpTqjXCsS1CZ/9ibls/Qw4RQLXq+KgkiL
jGcR8Tknsp75XWAqDG6xG6kIoJVjskYgBCCknSXAcp0+4BNqPzYdgGR2N4S2yqki
WBMJj/hZsAr2iV6rJNiOnQjC8dILiXEnWl25JXbodJDMJAkJX1/p6//lJae25c8d
XLC+rPl2dlT5Y8heS14ltTBgw3q9ATAyrisDEjWStnqF9QgHqDfGv8rJzKTAAnlp
VhdFVmmEQsIBgv2Gy6qYrilMz0Sm4zzXpWoGd7dWc70CPGyxafJsOyH5hZkAjkar
4i9mV40n+VyUOQI2es78N/k1VHuAjQCXoEBQGZG/XXCpTKv7WZCtZdnKit2b1m99
CX00xvh7OqdkpHtZwYx9znB/xKEKpNHcwEK+sJlSxIgSQ7OvsUWuO2t5jELOE6Kh
IQ6sR/jz5QmamC3cezP3cZ23YzRkGcOdOtABqcjsjASTrsXx8Rr6Bh136pP+hxJO
jf3j9Hvdhwal//dwkqltlz78xsdJECYUwbmb/UFIC5I2Ee9dQmDx7c07SruKigHO
X1vnig+PIIMKTRAZUV2a79HzeAM0lTaDM1OjbRZe0gk6Ro2SgwFDegMyZnHE50n/
MojhkbQPUSbK5LUFRY3f3dgwkLajl+zCmIl0XhDbJHpWDv8MXa8oYB3AxsgIOyXd
XEkJOpy5vaeMY5alMwv6oiVLyzqZbjqPGLgufH2nB1hJtjn1fgLhUQ4Bq4JhWmOT
otyhNduIeCU0Svryq2h3mQprleFwvE2sTd4Niq2jyL80ALkkmMjKh0wOgj/GZy7w
xfeCfZ7FqYgrhpszc+Md6r/cS5APqtn4Z/DrGAroqfAQ2p1LPuKq0Vr5rHYA9Nbe
Z+rgczMg4nEnVUUA0u223TufRXnPQvj8P4LIMH7C9EIBG9OMaGXzme4y3TV5KvJd
TKkpzrLJZrj5kn9IAEzyinqGeZBQ3rJVW5zNC8K5N1PebzjE85p6zE3q5cp57iB+
5pqOnPUZkOnIKCQ954fK5OYHWARfUuRyrE62xoo3V3WoxFl72QMK4cWeVD2EVM/6
K8dAPFsGwAtfbln2HDI3USWMNLh9rXsZM4xr869mHNipkK1L3e/+2bcQpbr/5QGh
hLOFY+FbTK6UGDN7ZRMWOMgEL1lUVRqxN2qgCBwXDn8ESjJ38vBwOUd1YF40G551
b5GTiBG+b3X6OfLgyFCzPdHs9rhK+ccME7BSh8nnWxU/0cxZf8lbJnBPAcDJCGUF
Y9u3AMQ98xA5XFDxdQBd9j9jEjbpxSAXGoL4jZ8RoGC5zS9F0UzBjPIQuM00Bcw2
tuBeseqOrwhCHsEjzwkSX1eMSSS3/DblLJWzKUziOJDbL6gSvaqA5k9GAgd2HFof
86Av0AC0NDmd0eQFSycHp9oW7/lPAu79ToQFD7nDM4nm7FgpCVXtt6Z4Nyu7v3Fj
7eHDV5CwbJ7ub5EPbDT46MRtIEMftCtVMw292gzpfmTWGKyE6c3jRTDzrTBo09bv
5MV+IeAJfQcJa92pqska9iZTbZ/TfptttjumcOSwiw5I0ddkrCayxHjRaSYEFcRX
lQscLe3e69I6MSt1nXgX23EAJ2i6iIB7zmyK9uSGR+buvlkJuzp2CLPhXvjIr7b+
7MJrxXwZHHRK1+K3i5SNTM6WxCLT+sNVkouUYjh85RHoW0n1/8Dp0jXntlG894op
1ec3dKjO7BnfIHVO2o1q8ndW4h+2Eaz2uAUutzT1v9mpaC/5Ikud4PzVX8NgmQBk
DMkZwNtVuMTcvEKVRDSKmA0QlbLJhpa3yTS6Tu5Ik/8+UFaF+DEOvr5RJ8fUhY1B
lX/0+Gloybo3RWROnGriCt+1AqZbafJRwkePaRiLcJFoSbOSNj9PEf1WChKBLU7w
JXNwsPAuR/RZnL5MwgiC3Gi+5tIW5F4hLWxgnB5MtE0c1oBvE7X/ryMyXTieqvtb
6E5hqQV/7W9B1egi5f7+Qlk5kWKsXYbAWaEyM/oQ1Gu2xiGaM+fNnJLhyHShSGMT
SxtZv1lRhv1Lo5M1TLxRVgAWjEZr08InL4AraXxWiq6Q5xg5J1pr6n1keKeRn5xD
2R2QQcjFh5WX47qAyq3yI6gNIlTJu3CwxHNlkxpBUw4xSSMuXyL2fCcGqxjHd6vq
skHnBEih5R7Kq8yyEGp6x/rnlt+x8ZET6UR+4DVXseaNTsulJpPZbazmdeOo9A7/
ZkIfDxztHAO2e7sKZFH/1f/PPjhGrI5MYPb6zxfe8s33QtvzDQnhYNrDbjNyL6ed
N8Os6EFlL2zzc9xgxdaYr104CU6zsnZvzwuRESC515pzJwpCLwPTWBpCzqJfxrB1
dk5uMb9s/RpnAP73qaVy/tPTmlW0LF8uhXnHdVWz3NqFqbkra2wSAimLE8nsVjA9
BXfIZrqGvBq9UQErEySz2iHvYB4EPE3ep+6iAN3zdmWTdeYBdQB3W/7i10byI7fq
c5dUQxkapMFCBg2gzR4M3+I3nWnZUnUUC4qCDciMBRui/WXvUBu82aMo2VyKP+Pi
o9ees/jw5uUrfih+j/3jM7nrYJJ9/B6zEoPOou8IoCq1RVlvVzRPr3xvvr954j/b
3e4sC5ta5lGNooA4ZQQJ/GDKKPrXSy1U5y7p4k5msW3IpRhhSwYvjalht/Cig5fP
yvU9+CPpO3c5fu7EdZQ1Ce/wX3qd3/tgET9qtv2DELIsDh6Qi8lynapChAqWm8vp
qIH2MccMX5pX2EkWjo+MeyzEVgbQoABRm0NQ11Qd6mFQtpw0Up9AtfmZ8S3OImux
HqZWv6av9JQQUNjGfKafJkH7l0u0BCTPMlX8G0robsY0JB8QD5xW88sy55PsHojE
CIPtXXuFYSyg+xVEXPuJb+AiHBYxEgBgtAn0i1GjRxyMDUfuPSne7AvUuf++YVJG
7GkMbVWSdjYwSczeRh/r0v4ZkX0taqZEqWivXYqvecwrFYUJ9x6jlCW/wUlBhGz6
40CF83+0dIUh+10Jf0mlNEkedVuj/loaWlIgmDDN8eLKJral2rFRWcIQTOR5hBRz
maiKL/Tpntyq/fZpioah/2motxPmCJwW4K5Z0LiqZQSF/Txf2W4gwkiuRsOMjjp7
x5ZzvHnLkKYHQMpFosecYW7hXhWto9ENSzIrOyZ3/P9PSkhHQzySfSJluDiqO6XN
Lho/STpdnafkI0Vd7Pc63kcylQehLZeSIqs0AKu1NLGvGOJxLFCwXSZ8CQrtlLfi
TZkxPPNWu1VrgDVHr78kuGtioeLaQ20FO0wcHqlnGTuCv5yaLY96V2wnJbD1um+l
elvaoDMR+7EesxabbaZtnlbEQfE8qmRxoQj7sHCfN4dsadFlXIq1M44G5TAu3Gfq
P3yRsmbguznm7BndOhblA04dnrcMgDRqImbnyNmo/YIfH6TcMRqUVUdF0+DCG69+
+hEWKlGFNl3sOFWOguxicueoioFNDHMM9A3789ZUrL31pPVpXmDvS+HiPLgv5m/O
Qtk5zoMCAS2di8o2RNCtKBL2Q5w/vuVBLTMjoG+mshgJxR4ipU1MHXt6oFoN1PGA
LP20hbAOPd/8mYkTk6+uCeME6RKSeWyyw8t/o+aWX4mJpV1i2iOuTmdM1r+olLKS
47BmJGP67GQCxadPSqlZ+Hz9g+BJRfDkt8iseBsfByJ6Ka7VCXtGlChFIpckZ90B
Xxp3N3c6AY8wDAh/NIfzh4sL5n7rIAEVf6WOqBPCRUexsIamsXWaJiA0zW/6fAVh
6fSH1CCsuovO2HwxyZn2Fc8FxUV4xvAjflgNijUwva6xBDXBwXUzN5mi41GDx3fG
+47a38tVeakXCCMvIYJNr62bsjYXFdiDOb/wJijS4/ejUcLuqo6uVpaqWBbiUmJ8
lZ2hSElCqBvnQov73t14wTtEv1/GQILz0j7/8RX3qtYjMbbY/Y53BjjAuL1kQR/F
7zhc2Gg99IHbMcveHHFLCiDaDmaHVNpFd7Ir/RrajcmfRwJukcOP8poLfhfBg316
pOHINKkMspb7iD2g1Y2STJYjIigXurWtMHLyqnBlFVEipm1BQE+Cq6Pz92BLdLfb
PUjSzKUIGn6WfVj3F6VkUl+8gLiuCxgIqACfgrKN+fr14virBUSyKDkN8nBqkejq
6/HJNrFu7c5H1UXIc533R8+Ug+YCPXSB1DTiPnjG18xbmz/0G0Gc5YlQbkZYDDtH
wKklrUA8+capKax6eTQoUaQBD5fup1R//ldAuSXuvLkEK+UlWg+ZeCnLHO06ky9L
ndPUnVPoj2YU+4njg0AEr+g4/kTPIPjaRU2O491gf5R3W98lPoZ2hLTHAWqH1icA
1L/GpGCDHrEJOJjeg6ykDRKs5TdDI0eIgEQFT78jbsqV8KUhNl2B5fV6gSqW8dEk
q4EUjUx61T0UEqDKlLSbDilEF6SLkIcoAhm5E98J54VJL+04r1X0Y0gulKZUYUXW
k+3vVEglnmv9cuabgr2OaJTwYuUNbOBNcCB3I3v+VyUnIlOGeCVXBTyfve1KRWWU
9SPilX0Z4VOJtC+KCv442r09CnyPZhbgzBt4Lb0S7nLLLv2cXb7h3ke1u0xujW1S
CXQYcI9dV6oyRThDZ29i9A4lL3TUN3Ojb1LGpcq49lpg6PzfCRnGu57C+8urUBY0
7kgasQrdaQthc5/7ZVd4kRmIDMOydL7GrTnj1FKL+XV2PnnNkLj3+r6IRC6WuZOP
lUuPiB85tsLY8Tb/zxOPbQpafDKDKR23J/1pUHM4nIJbfkr7zhsYkGy3PEroOM+t
z1Z8wNYrhTI0RUVaSkVpXOl9TVeHnBOngiVkctHlDNJXyCw541w5U2LKiQXDwuWO
QnVZWtV5zQRUpcP7ggrSDdhV6tCR6Q8gPB0tXVc9aufjhTXxHozIG/JMBGMsqk8I
+OnO7fMt4q8ARi1Kg1jBqPCjcsBWn3vm3fDHpYI2wojE3LCYKYRvu/YkGZ7MxzmF
SEzBV99wGQvVFOBM5ri5tqaRBZwuCLExDPDrHkXRFtN8BFw5YqdYtxToz/EKiy7o
3uHMLA2QOa7fuhKDJz+YynVNj/Gw0wnXzuy0b1NkjDwVa9AH7FydaR3987mKsEoH
k9Hg/Q7oF04Yf51ccAX5aUXNc8/TKrZ9s3dmsgyq2DPieKNnTxtsxdkS6BXMJHO9
`protect END_PROTECTED
