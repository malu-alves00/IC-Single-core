`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZV0h8ZSr9+iwsqmzHXXD8d/SgwlOXLfquTQV4OoY8CBcfqQGDsTG3nQTSUuqZQnZ
yMMsBCuhykhGhapwB8iYOPigIwYR7NGnNn3dx9K9coRvaEAtobQTLHDXyNvSeVRk
0ELCvT5iEpTYr+PG79aB3Dc+8iCJ32de78aRxRHm/r3f1mucVtyVh1tXx9WXHKGM
ZJCZo1JPM7i9PtJomPgIofLpNfwKtSOyMsbt30sWM4XhQEj+Sc+XYNbhKglweQyJ
lDTuc882oTUplbx3CkQ9eaE2ry9Q4INJ8O2rWV4Q9bqpoJ5ViCYWi97bHwkniQmU
MtCf+mbuw4XjVQzWc+LZGWFuNHAT9DL0Hzi3+nfQvTOp/kBGFMRNbVa1yynRHpqG
6LH0b8u5mk1ynYNrP0d3XPjoAAlIdFX0IlDADLrQUtmmu83z4em8Ub6Bnv/YOcK0
nZX/dFqSbCxOmc6iTum4xvJCLsYmrRI2wlM48z1NZesfSO8ZbyLJ6s55DjyJ/VDA
QuGz4Qu8EEq4yzT6vnc9HuMZV4GcA8JS6aYfko5vyjFRbIVP/cTIrfoNpAM8jBN9
2wJ8nscARVd1RrntCJ7fyurELBiR/dZ+7UI26tjoca1CGuvrSJEwRu3fseetSTuo
cjMtyujTDxaOiVkhrnw+lWm7rmDNVtPOzC55pClaTRgdb/VpACHfpt9QX764+Cf+
2xripUqjbebc9XFNbO87KkgH0/lSOiKOUq9/ZwNPOYuql/QP6HhSZfRk/E8IWxtL
a+wuwbBjT9GVriAhWu6zNnvSUfu1U3vDORo2Hc+cv7H+qK++GJAsH/fga/pfL5a8
wIvwwzLyiZqG6C3gabyIjqAFSTUjkdpqweVAWFKRBSnM2ZjSL8lq2S7ZYF7gkMbf
SthwLFLug/NkNRpnDhlJMNHRs7AOWyXNZ+36aN9B7f8rw1kIRRIRqFaFu6BG3CD3
owPe2GION0W5WUbeVGDXS6P2xFlpVOx4AK73OJUOwErarJtSEY8fKAD9D+UNxiLd
qkohf2+1Ko6611MJcGHhGROuuxtCB4iw7qe1SgJzoL7i2IQlFYhMH/ZlWH29f9Fp
Qu/v7mOo1ILQ+bYcWkAQMerK/8Sq2iJpxRSMsVwPJMZJ/nfdrPzlOcsZR+UDALms
3tLNu0VoJyT/gzqurEOljUz9Oh4dkYS9awv8VIy5S69uQKruP/FQSqKunv2xb7/J
03CM2KjCV5dkneCOEkT/HYPZf8FmBCXrwaMqvyjFWnxmdQ0Sr/ekLPqL7PiGgPU6
Ad3YO8CPXvJlRyZVG/ksiH5FTKdjCjvqqJMiQrV0mJmcvgMGo7VwhjhAbegUCtrg
YJGPMKvsnj2fwnYwOiHUvRW7h59dnZuvNnW7tTV/X2Hvxu/H6uZsSN+IuafyM36Q
HkjCcNwmAa3sYu/QvW4k1Za9NX6CcRdgo5gMg4IxSTUYm8aheBnn1WrYHOCis4KJ
C8Nms/OTSZj85bLOgS5j538+L0SvK/sQmYHT6jszz1PnMM82ZGf6a9dVNSWIxVtO
i6dIhQAs9jVL3ZZuwyvBq8tF/X6Ok1dXNnU60uemH8ba1bvYJhTvd9TM/H78r/Wn
UiyYhoOqgiIz/mb7iz/28++93szJax8GBCik0oAH9YTZkfcgaM4+gFk2llpe1/1y
zv7OzBUB7oGw56GiFoQgc0/Ovp/hGLbeLKG0L3N8HNUV5rCOsmV1gsyKTcCbznLd
fdG3o+/G+J2rVcLIV3WokcUhGaZeLJVg+291AzB7a3kVrtJSJ/4ahmBmvcFb38hn
E1tQYSm7QBhtTBJ5jkzawcgtTttwlMnOBwTlDJUJXvRYvc2BjVSdYzCBopzbrnPa
1BswoUazlwaZPwYE7Cfky3Z5NI3u7r0jv+qaeYjxXwvC3y+1Oe7Y9odoW2BFOsvh
JlLr0mf3nQglSpEZcOrBo8lL1Zb/yBqDobbcJwdXwZVLnBuZ1Z0fMTkV7FGkfh84
pzK7/HdA5zsYZBiRZwNC26Cc7otieMTllY0OH0LxVqqF6Kz5ZvbRtWwiTCinQLu9
IEL02wjzorJN3nWIlT7pBQ==
`protect END_PROTECTED
