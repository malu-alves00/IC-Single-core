`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QtzFsKFMIEYgAklNOKHw7gYqrZE7mglPqHsV/YymhJ2Q30WYECBPFng+PBqHo28R
x/WSUt9bzZq5fHQXpS95fy+HiRKyIlxJ/fc1lxJh6RuyAp/ssHg13RsIs31IiJj1
c7tD4sc0PaxkknUSEn4Ll6bLhEdoMpdiJ2igTpzyK89qijefIUNgLJ9nIpot/kll
/cpYwss8+uI9na+ftBzx/s1r2AjqwOA14A9m/70Bz/2xiefVoW3r0p2xzRGEX9s9
kWr/T7nNVfGiZjwbD7gNaO5+lR/3335V8f5k7SkBaG9kZBdug8Uk8V/KpO4dKiXA
0EVWFI8mu0PfEGveFCMON7LnKPix05CBlmqSuL0VqlIOF50NY0IxjYOmVL3JoISN
Det7RxWrHmyzMAipCDmlYKlvtEFBtACwMaSCxp7EIB4L/s5urzllZ52Ml7s2G1Ta
XVm1XjCpK+mEsEP1dcTTUqDtgoxn77wKSL922N3yUWIlHBLP29RFiG8sU4CfYExb
8FZcO0Vk9FnvjXLeWIePBmtkU6A47ycs1b4IcqNZlNHihI+BiIaYQs/zetDdToLF
WJig/wwuDaiVsGgboUTN6VtBtDsUHYapO13Cgi+fY+mA5FePGaG9rE1sOj0u56BX
3+THJ0A0mmys7snVQd5ZUw22F7W53X7IbA+WLZHxIbWXJjv8q9FktG3rh0F9Unxv
KiZPPlXMbc3o7MAO+HNwVnioKmXUWBc47W5H2evczFoWt/DNElR3QA4ISQIaCtvh
2DeHbrW5Z6m2SaEhb62KnwooUhD+w4ZVTU1BdvfD/lkjU8GCOSQI3ps237ZyN/G7
uQBPes8J50H9cNpnpBoeVnzRx68xRcqSA/zoHHERyuFtu3NSbFYJrrT53MelvYOX
KyaPQdB6f7uH8uV38LtTCx93zUj21LznK5foCzISPhE=
`protect END_PROTECTED
