`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NUE6eamTonfCjapjeEldGPMDIGKMrZvKC7LE4iUK9KGhZozPZEb7epkQa1sIb9+z
iysoJ908LApln//GCb4u786d2FEGCmZBN0GlzXpiFfL2fxF3mONNrJ4SEOZc/B/k
D7BcMIDB1UjCC8Tcti/bQ9h1y1rfgiyqEf+dwHBdqg7GsRdZ1SXma4RBQtMIXFRM
bWeoSMEPoKn+WilHIR9RstcjNH1SY86thQGXVJhyG7frZ2dl4zrXMsY73JB1iauj
JjLmMFndI0mdYwvQ0oGuaixUmFv4/fMIOnGHut1UgtEKd0PRDq4L7Fb8H0hh+0wt
t3pcQIoO2MBZuF9QZWFYXSHk7ri4Kzj0eRxOTN74x/peVa95qhWxrt5PDPOfukZ+
zt7oQJoyDnvX4aCCaod8+7eW83ZPrG/BTVp2w9wSSbcONXOh9ne/y2zhiU42KaKU
NtHvMJPSjRWiU3HjDxgsVFDL3M/QowY+uZJDtb+sOXASXp6zwlYg5oAxGy8ahmvU
ICCPiAdIaVthY9w/YPJctQ5cjcvstBRWEzmev3CU2qxzjCNlh0ZkmI/LjZKwMany
+S2dnVOKh+hEk6d/k/vAev4xeztFuZSDOW/EGjRGSdz9OQWE4GEeJkldulUCZL7j
M+9sEaoqIoaLBfAXRz71HjpJCAj+OTpUeUDWB8ssIv+Qdr9AtGbgSfCs3iOGtzC6
9ksAMULnVfOPAS0d9cDZhXat62fgbQfjJrCaey99jw2UI1hU2WVoMXguXrlJ2iNU
+o3KeYKxIWh7m55zc1b/bcu/NCvO/nC7/Epl4YUvAcXyDKlQfDYZEOh0nW98+qi/
Jt+4kzXA1nJso722xWEu6z4T4rQ1V2IdwlTLIyYmfTcon3ObvS1aQTx+TNVZYR62
/xHDXnKHoLw+QQ7AM3FA8vXNF/E4XfvP0bV4toMfpnNHIzGEaF5s11JvVKEsjTuO
Fcdc0VSWp7CQ6/lcMwbVJWpzrNbbRYgs/VlQ43WvPaBKB5NlaiNxXdPIoYCxdiVg
bYWSRQwOmbZdhwdSMaIIwzWYaZjWmdEA5Jbw4mU5bDDiaBZ0x4JEkNirzgUO/vwQ
e+kP78n7o2BqnEsrKepRO9iMoOdjtxBCVM/jHkZ4J4Z1c53gRHDteI9Xx7bSdYCU
7oayvUW8xc1rT7173JHyekWy6+u+DHNy1VMozFkGkDAf6NdCAwaIiH0sCmOm3jeP
K83bQu1nqcRRljWZewxe8nw/EGkViQYA68Bk2vCfAP6MrrIVykSlRHotR+CH+/QG
W7+PYTYqJ+i2mtMdWACyK8SFrc5tluyTmsmNRZIsYfEq0aqreJrRBPd3UbVHpSOG
zZt8w18RN5vlqzGTtebj5ePPRhUNriaiQbeH35UJPItDz1fvcQQ2kvpnCuL2tnIo
Z9Dk7yvddtSGyZF+pCWJELF828MFzIeqbAQL1c1tbBw3Tc/smwd+8CSLmLjl25Wr
AXTxyNk72QPYdAji5kkRjD9TRwOatmaaQpGp4Wp3OscYApuwCwJW/cI92hmMYwid
cyuQ/xpaCjJzCRNGCrjGFJ8dS9Pm80nfTS04exFh4c/ilBd+67Z3IpXnFD71Jzbp
17HV4fFTY6FEM+FTAc6J4vwJc4+1HhCiCSJ3tw983Vzl/vNzrbjVyiGNpx1QXNfR
QJVhWbSLiG9tH20ONHhqNlq3/aQwsUGVBSaQk5EaGZTSI7sghsaSGH8pIQBsk6sL
mmTDnxH3kSS+wjbktZ3yQJObBKQ8+Jtb1+FIRAaN/8s88o1qXy+PfwgauQByp/Y8
icj7AO4M+DbtObFYtsAVyXrDAej+Fn1yVdh1aprBfwXyJ8AHvOlCAx9TRqOZydt3
kK4rMulTfOZ8POzbzzB05jv3tuLMozCre2w18bjCj/MvhMKlK/WAM0rT4AEuyGFy
dbzmio2qDA3hCOufb0+q+GCmczBl9Z96OVggvQUNXEm1f9VskcHXVkrW0dc3nUzI
zqQmEQWGcKGvyrtgHvsDf9aG2alxLvHwEC9rdD4l23bge5bEAqKTZrE9xN7H22Q9
p0UKkNif7aS/YCnLcc+hlaCa7GQ936enYKnH0Yc1870psPlgzQk7jxTkNnKKjIJb
Li/N9CBqMTsSgLEAD3hm5TbupQoFI6wBmC3i0Aanzgu3ogmehS6XpmJpge0/M72D
4QYZzG1nblyD3v7NL22Od854xMu7QOOQtw1k/ZL1XD0uxOnSZj4C8MGsww+zA+Ey
cy5D5EQGOOyxZ6azWVrfP/pVD4jogZPZ3gyPHvzuarBxZx0K5tp4TpBtBcV2ZhQZ
pJ5Ot2tVNg/WIQew+3kxM+MBXXPQJ+LaFzyyOGXGZyXCRH4zYw5V6vcH+13K/ivU
XtL4dqKWKzlEskgYPJKYsUsDzFcU2FWRBmGyOYKtbECHR/Rp7zqZe97Fl6kUj8zb
vQYXkgaicUGEyXSpIsT0YuLuTZRkCGLBtZ8fhOwLCJD59CiWa5BfhqwZLm5THm4I
lz6OC4JfGuVpSinoipbdeBueDLo40ONik1bkM/lgHWIzO3+mmi9mCanIS3mlk1H2
iZecVsraPKMJM56hAu7oaZ8pBUGhn9cNzUWgxSKxeqn6s80IPMO/mBLuISqKpoPD
GDfXTtP2uGiAuK+t9JHOR/ihA1pECfSSgshNo8cixD+qTRZ9oo2kBtM0BrKSC5d5
7EV7Ctai9cQ2X7suJtqVExeg9DAljQ4+wsYMDy3f0CxftvF0Z3+CCIxjqq+lcmei
A+gb5kkmowSpTRQSlf313LrsnUeTvTa48rd4fmAhjw38bp+KWk+3EG/VlBL22j6Y
RHL7+2+kC2I3agF1852UU7XXUTegCDMt6o3b37noZ+50z7n+k6N3Bw7P97vPfOFc
GhyOeJFJipi0z/pV0YPDL34Qf+/g+YrYo1piVRdEhEhj4OmPuZl9FkLt2VsM/udJ
yi/0VGHYym7I2rrhyvxv0UgeJqld/NzQ40MXoAzjTWXZcRDV4HpzrAN2TgJBcZ/t
mayvzhGRNAfXhrhKhv8V1pGrGFb/r/IqJqPuOlWEgk3FiRb1CJIwTCZy1jN3Bomv
qJhMQq59yL3Yt4A/qIYd32te/7MiEmy9xvhDkWtLWs7f4jWYjKBCvBDpNH/Q8Pqv
eBJAeOTaqgLmscLI/1bzfnnrc+glsjdsHNLB0bfZYzORIhbi8NL+tRa8igY0QtXr
Y26NWIohJvHUWo8k4kwAsE8dwuDaesxrVsZdNa4vWqq6nefmKnv7x00YXUSHzTUR
MGvd3TwY/N5ZMOtkxtnYNbBvmCcFYFL5V7sqLe4fEQyELdYr6Qxh+76xdcK8hGPT
CVj+/EQad87nvTtHXaGYG/Sj9bpd4PBYTr0IEvJllvPzwk3g9K2TxFZUd4KXSdCc
bcU0Y2j2QJN7UtPzNpgS3mdlNvx21rzGU+60BPtvUQ4NDTSYdyVt3tCB92S376eR
`protect END_PROTECTED
