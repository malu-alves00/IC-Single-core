`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
g4QNmiR3i0VTwAlzmWOn9oC9KRf1NxIyQncLSZwWEm0vtFW1Nyajhaq7l6qmc/Q2
8xZxhQacbukU8P5LFeSMx0itPnhSdJkRnBlz8YbxMbFhoc5G9QN7fzOVVZBAsA3j
/60oHtoAlokeBUjpGYfUwT/Z4siphPQDGPW/TXIrWvTQ2h7nJCNqPDQanyZsiSgD
DBeJmCN8YJXkAd4eHcJZexwSJO9poEm1xzqVatn3hQJrznuH9ZT/6G4o4eJCZALW
BTTXPb2ppVo9mslaZp0WDTTWN1N/FYJLgCeFdXfAvzt2RaCLnLbttUKh0mF5l/mz
1jxrQI0UtEn2w5u+iUosRt5DRYBgYvMYElkyzOskF9NVRK7mdcsoRxzcXTpk7YIJ
64Ybv/IWHjtyePmyu5Th0k0Yl0dnC4XtAVvh5inP3glsL8hTQukc6B39hJZJjOf7
9Ie0Rlr65bEVZzP0C3VPq/y2W9oJdKGjywUYdK/hWowkEXadspkT6ONfD+ASWmqC
72X3UPZFTaijlwKxzZxqKtm2sM5R8O3hizRX6gqjZwcqPySw80gGqOz5k8OOeql/
d5xhZVaymuBPkVeLVvwbYtGiaLIkkhOGw+TV1U8j8l+qZtN8+FiP1K9UqK9FR+dy
40KLWJGDEWz84aa7M9b3zRI2yDlx8Atsu6/oubAzIbPrtqX9qy+ycsHmNqPi00Kj
x0tgivGKVjPpqgfdo99ttLyWasLPVYj203DzcGmX+7tVd/63We/bT3kPUQs+WU7C
iQC43ifDqaAZWDkqz0ZvXdzPzOuvRKJKYYz1t72qrP2rXbALE6KNm7eVDWr0hD0K
B+LjOEA8hN67iIw3QqY75dttCkbazELhI8uF5gVx9InWVh6sDCtn+Hag8cTR9N1n
JiqkY7Rb0EJiAe25Nw27AW99XZlwkdl8txXM5FJmEpL+8elkP61CnrVTbD4moNiQ
UXDsoQu35MItV3a2JH0a/9iih7ccrqLFuXuRxBbsbmRZJGCoCJ7Fnf1noQ1rQ/t5
k+oKS9SfZOf5l9qIOUc3qL6VZQ7ZAQGAHKBm/gu4qIdXgWm6s70v+X58sAq6JFvu
K/Zwv08cH3KOHJoD8nVuLhpJROMhIvcS+AWlpDTi9QtMSS0YvQv/51Fd5dEW/7Tr
8FhlNCyrIe2dQ7KE1E6b211anwvvYko2JydjTcTto7FUccAyOD2LbTmDnn7M+G2C
6vbq6vsEfL1UnvOVe5TMzKSFn9PZY1Mh1QW2Z9PhxepMvDYd67xG3THCLl1Q/VH7
xoVpYu7EmSXfdVUaZrh+fb4q55E/v2tINGJ/G4sGlsJVer+Mpb7ihyWl3yFZ/4+T
vXqP4POHiIbDTyHKiz65JEPsZIg7+nPugJi1wt444Zcx5gQPQcmwMBmajSwK+mKH
QBiv1x8ubFUF26qkzmh+FFLPL1Ir18vwmE28xFTfgS9zZ+LwGGBqKEZM5G1NBAmZ
N+vJ2Je9oHBMNp8GZnOVs6wgdlSO7O2iswb0N0CLyoelpW2wdrmZRmn1Xvh2JlTS
JrGfIa1RpS1s9pune2ZB1VpjxOCOyB0xg59Ren6G0i3+gLJfpP8j9q35GBgg1IPv
Sx1GDi/smUlzOjZukJ3b2Mk8LECHC42EJvot1ZuC9tYYHOIL3sTCbSQhCBXsILS0
kz4Savg1Uasrl9SBcgR5NZmns2fbKSxWYNQZXFR1fsRfm/k6kOcWUwvCYZ0n1Wo7
J/UG9A43aGhzOTcJavYK/gBQJXJ4eiL9M1jP0J/Sw+0ZkVOCw1M/uZRCvpOrh6B5
BnXxkSLFmW1/+boC1ZMPAzeANqRLQ4hOf4rywHFDEeCNbwqn9DwQjhgOr++PfBHi
D/kVDi5M4GbeW3DrXmtAfN930gpvEtmC7w2fCjG/A26mSV4lOw+/RWpujY0EVoPJ
JRIXcB/YP4541PxjHs4gHYG1JEcr9fIUuhd8bWzDzXeI6cacQOTKFF/DDcpDnYw0
SKGpisMvUHJ5lwx6s7pa/HMQf+E/6fu1xBULip8nEbOOIo0c6VKbnaT4Y6U0o4Du
0LkWiS291oydfAhTcR5Isj9Bm9qlx+HXJEg5jmKBG3TbptZE1B5kaYDMml7mskpR
GYrq909sneTUL1KeN2KlBFggYRL6QGyN9mrf2gIGXrXFFdrG7iOk57H3ebd9m+2/
d2PE1NAES0a5xG0AevNoK7GKhQTSW0LaDM1OLqzJ3yXWBGsK2gKhhWTF3cggZcoQ
rrN6RdVsutSR4dmQorSKFXDn7rxwv1xCi3gtHxxBdvoUaIQzTvP4aoivUK7/aakj
0nfgziUrG1EcXB5I3AQ2D8k2Hy5NBmaLu4YkdEOBwIZlrye5latVmzZQ4CJq2a4z
2HmuaUChIiOAUiORAmJMmCOOJklfm904nJNrLogCs88B0L5QQ0LiFFA3ZP0Ft97u
g/EKAg9xWxLk3hBBGzc9EM6j6HyDYlS72fl4MJCWB9Zg+/ImoFYRxZWeYlytHsYW
VI2eGjEqejHw2yr/CKf0+TjXVXNFkSf33mihDGCphZLl5ne0e6ROf/6wlxf+BkaJ
oMpF67itpJWJ6K3qZ1+FsDuaZrPTwrZajEAQ+Zj9ZzrKKiBQo/X9sGbbf7Q31c4D
K3kA8ovEgdi7gkJcFYsdl4BYDeNpCmxCUMCQILcTVoywi4uMqrHsE272ng5xSirF
Rb4v7f/qqg7uUnuQCwUaKRp13Zy0S5ZR2Eewwz2t6o8Iveib0ubErBslwkFV79RQ
Mt6YOrmNrNMtlnL8dkVWHWeU5bWQYLaXpKSKvZjFqvjprUHBlCKnyAPsBgN+NyZC
G5YaT62NGgou/AheoSg7RxTid4/9QkXP4aEmchSOotYSycLor1FLHjxe58eGKOF8
xiIEG6sprMVn23vz/fCM0sRsfTJdKJMkeSU3c2FS8MtJoaWaV0USZFZ6oiveF9JS
vbcsdKBq9Q21GRYEUPT1hCGay4e9gXhqGkzTPhVgtkH9Z+94gweVC/SnYqHvt1Cn
bFREBbIs6Tvn4/N+C2V0r+6hpVouGJhoXpl9IRlMeNujiNfb/BlVFt+/WwZgGFDn
Bqe8ihCu7jScULEBHAGOoA0QstnD+MoK7E7AH+kQstj+CD0WelshLZnBRWGh+7f5
dpv186iMih9Uy3BATbFPxrLtTwt13UU8hs8zfWHIh2OK3DPvC0hcMn0hepRJTaNh
cn8+CpuCDbDoIESXLtPbAzI75urpU6RBRjtSBoCmdBYeZ9dSq5NZq5upl/MW9Buv
q52zAzezl8m525pOZxExYQpddjN9/RFyuGD9QC1ivqiiQ2PVXhyd/2ShQX3Yep8T
UcloIm7yqTGR4eihWJ/qLR9FG0QS9QoArR1VkWlf8fJLiAHVMZP7G/mEEUr4pBxq
WaLL1LVr/YfdbMrJBILj625Uh3naQ0SCFITDTZuEKnPOcftcO4mXupMdaSAUbfMt
FErTgeRG+Hv8HJpwC1YZl8jjC9okmBMqVmlveDsfeRau1T/srxEmWIQq8OxIkxSx
0PJQyConyBqI99q6QqRFewNK6FH3wg+V+jfWWwaQOGy9rnvYuYpAwpGrYyd3fTdN
E5j01YpK01MdrXDIntzXkTSG1Tg3qxUtjT0i0XWfnb6ZHAhLyJjjRSSauX2KcM/f
awO/tTvOaFeqDif8hBu7dd2yJLQ2woDG1sNtwFp+Od4TNCSVjuWe2DJh2IDDPQD6
bXAn48EvWNhloTmh7o3wQ7iSRO1XjCKX+K25bRDTbN21xJd3lXdpKOk+LT52CMOw
BetfOB9CcdIeYuu26EuB0jIb1dFMIdelJDJoWqUNK6agDKEYlC4Rm2DAgMBpZVYx
SqidDcRfAwgFnGwZZUknOrjdKh1qAura2u/1ZJauUbTx8ke4aDbmJPA0XNnJaBQS
shQtZ+/H5UxSK9CMbw8oYVWWDk8pwrPPOYvWfjyEZyeGTdIuEicnToFhzgYXuOlK
Bdc8jN/ogyH/Pexd8RYSXUwBJC/FFel6U4cIDWuKRm7pf81Ie+g+ZL5b2bFy9Iqk
zy3pphqptjNiK420lSfdBu723WeB6OZ2vPfpm3v4p9iIN39RGOWrbCmaSCrGWhwi
5eLpsQ+GXKGlO0riWT2UDzPtJqN4QiUxgy5IHsVxmoysjVqxjHkp9zwN6ZuSy7QR
6q37ZwucOxD7xhKFzIp8dGQdOk9t5V5NspzPjz5iLiWI5Zae3nUNjXnGGTW9EJcs
w5CwCUgX5vTQbbDlVPYDnLvjtPlWQ89cBEZPGoU8DX7YPO1OgjjMXlMvg2x7Sa+R
a4LX1IVcdOcQmrmNpdv1UwspPUJKShuk9l4gDjR70lZuDTs1c7IgOyB019pfZpR5
4juXkMAVlm4L9+bp1fbRSogcaF12pSqxn8zFwBR6T3kb2Jk3rR8+Y2ddYZ+dt+Py
rbO+18wtj5PIoU8rsWx9Yrt556INhMRTAM3nl0Www2NlYEzYSWiTWttBp+F+bBFY
uKzr7Wyo2cGkHIUFcaWopig9wBCVMe/C0c+pn/fJjBS0pBIE9chI3J7FfEsKNf0J
oBNjTeHRIHTjic9IBoxB+V0n2oZ6FtBC0s+5fl+FP7usGrK2iHAu90uskwN9lgxT
FVX/zLfiMTk8rCcXG3fEqoPM4MrY6AXGasRlaoKVblJWbmB7JGvuRum5CncURQNi
utnTVu1KW0eF4JSvQW6UMU6ZqXsi72NHoWv4WbWESdqcLx6IeUxex+k4Mktlk/E1
Q5AhDjc1y8A+1af5HFwDdvjgtTsrZAk8f+vtHq1KDJjo7l3MUKUemDLN2APDL0hV
nS4WURRdx/QEA0v12t0D3Te3HwBm77WncSLOukuOeEYMn0LE65BjI8DD0B9VWVTk
1pj4sEjRE7XXrBuPOOuCsdZd4/8cvnxuITe930C7XXDghoZTQP+4AO1gi/ZH0DHb
kVWKZhfP2cJ7HlRK/a5aoRccRUxnMLD+oVROsjgsf9Ud4yehFIZnmqPHXNMVEN+u
uwWGEUae0KD+fLyLsW4JzP7gJ2FhaCQ3g95iBXVN5X9diQMYjTFJaXKYdNEm5Gu4
UTCyxIbQdgku9/ZF3PUhQ/CXUx/9Udude4P/vF28mDQesidp2KIdEWckMj9CjV/s
MefbZmUXPTS+Gpi6opW+pS/dDUtHc+rrfMIeQ4Xd6S+0pI73KgorSHwOQ+IYI1OR
5y6Xvd6C9nXGsBWhQG92+huPr6IB04tS6PewIUyBWAjEmbNAfdQh+YJgEeYckKDe
7L5HtBuSyB3rxr7bM8FpKT/tUckRYPGjrOulYsxalC6xV0OJL8/6LM3k1jWe3oi7
PCQ+xAZht+4dUwhEsBf4THjmOINky6sBVHi5btGoMm5HZT3c/4Eo9ksae/PNndqD
Duc/94oSmDCy8DNYQT5946ttm9GOnvOIPiKjQS1JazsSxTyRD7+8uVdzFcHqVXlT
iOOjQs8xvkwE9/Dg+7V7Poco3XNkgIZRVDunYm0uQieviqhaQCOOKkTcjC7BzzTL
2QC1dl3W2iI5auZPZzyBMDt5Hk2USgNOmou44sGXu4af/Shk7vRQBbwPRiwp1a2f
3DptdYZkvgNBfiuAVDg2iQimo0PcEBShi0yIDv28/Cv8OVese8yBnSXK9HcdWnoe
RCwp0a2luYlTf4K2rFN52vtqUQJcK6P/2LewAX8h6jTo03ozMz40yyj4xVcjcfJ+
BA7ScUtBImQe8l9mWzO2RQdV7AdNt1uj9vgc7hTZqqXQIWNtyyrEKJYkRMlaAeOl
xuWRWCl/X4GJReZ9OQ1Y+jgORWxp8YW146Nx1xrHQNruqfY8UifXBl1QGSlKViLB
ldIWwva+33LDTop6+Jbtmwpvl1gWwMmg1+rsr1Tfk5td7x5xVVLFyZHXOswLdUES
DSZHDmLQoA8zaqTuwTGExBx2g0AF6DEx2+qaH0VNDa3BsbIVhM2MXDhecu6IlnwE
ElL0mF6OXk2PU9sOh81eO4AaEY1CvopfRi40dAkkpTnEYfmAq7mZ0+cqsRp0HOTa
CfCpN+cNr4UjROLhaZ7u/DRQXtc/+Ubec/V8drov7qm5q6sp4O731kXMMlIAcGku
8hbTFuPYzwunJs4jAmQteDV4xC7UmiAzDYGgCOYcGU/GBi+36+NoQLNhSjvwCF9k
IZRwS7V1isJXAEheWyPgRDQlx+mDguY/MtduUaZbKkBmU2vRJ25EUwtCEGPesuxB
mAirZ4QRKtGRf9PkcHjkHwU0VhGlzbFpSuNsvA/cxdaC5cm81UU7owLcQe9wmsio
ueQ6xROOUyAUoXEJ8PWQviBHfy5e72f7YnibhqO9RP30JFZV+Nph55Uq8JoxPVJJ
TIXSO545DdXNMVW7wT4Wgm1b5/6dIQdiQNArFyDoINZpWm5nXsqH738qe+DBBGmA
vqn1RFBaKe18ifNEsQ5MkKeU9ma3wtwlhVq2ozlmR4opBqLDIxQxB7LyL+FlerdQ
SfXD4lz+DLob3a2R42PdK9QhcMblVUN/uLIRb5UI8bfefueN2w0+w97RpIEm2312
V5f99WWM4d2ITP8QE8KfEmtS+DQEisxXZ4mioKx31PfOGMuXQCPiqD8Qg6xEkbQH
7U0wIkdk/b6ZhEPJl3bPw/35VULy1UWBvyVKoVEVex0SHW7zuM1U1xAJjXcao2j9
pR0eI9+zMSatLpZXa/2NNpC/PB0zGKLWjm/A/gcTgBDo45FdBu7Eb74+zJuNLhyx
didyuVYs/qMk9O7WFJ1rY5gWhIHVYjYrw0Iyt6RcNM6szB0Bj1wNBsnLPshv5Lu5
jSTtoBl9mLU/PFfwG8r+zE4kMCl+JhqlsLcqbgbHkTw87GMfjh2cI1a7t1inreTY
R5cbVse58nNpqJ8zW+LM8TfpENdtfDMs2v3iY7DXoiytLyqyWasAlysOG5G8wYtp
Dp3Xa09MO6LE2xrDaowne/fmqssbOk9C0nn1wi0hQELun4rbRmiCTWOtVQcrprHQ
RdLhoapnNSuUgorFnP4v+WRKGGoT2/oCJsMYkaGawxZedvVOwNuMjlS0203eNJuQ
31GY+MfSHBxIj2Vg+Q+47WZqRK7Yf4yvnCjluA/6Z0ESNGOka9GRHYJgtw7TB2jm
/VvYFeu45GCgWycSPx+Hr36Z3P/03h7elU56x7iS8c0saWmPsqPkK9CamaIRBlz2
v64/shsUN95h7BDpyilsUFL6Brm7YSa81zjxLfs9JX3/K8uTybO46JIU4KYLn1J4
6r/QtdVTm6RNmz58wuONKB7BTd+Loi2YcFGmK1lccqWKMrXG+lsHQm3lqSlyHYxj
CEPE9IoBqLpDiL1kejxxOz27wR+ag7C3RFF7JG/2YJzutYo6xSuKPBt1h/W/Zt/X
weLy/kryIJo+hVbDQPZpK6aQTP57R3dZ+kKoUp5R+UOXOTQlMTNHft0vCXw7SzKw
mCamB9PaeGhH6+Q12Mv6A+Yc7Q4zSuW34l/obI+MNfESp1O9+gstIDnlREhfFsix
szmWzW/2CxoLjitlK4S4zWMl7m00vjA1rQ8EpRz445Nlik5K5q3pqJ+v9qAtqBh3
DqtMM57K1gp9vwqiJeib2rJB18E/53sE5lidXIFKLn/I4safHKfjv6HaX+xZDciK
a72DWBW8y8dLvw2QrZaGBGLqz3ZqZyixDamhZUzLtyWOggqoeCfpltI8euHrICve
ZBN9QnNLVJctER8oyzQdPA4MTueUupWG6vjcSnKZJcKkrbT456WOgQtVA1EE39Qc
WB2yTajn0nlQxJftPccYcki59FzwmxlJ1PbCmttRlRhKTpQnllWtR8lCYoRV/hnb
iVDPR3ZtGzsvRIdFdObFw1O4fsSxbbxs+4Cz50bbUhY1K0s41mkK2DFPdkRNvabs
sOnSgiuVUJBx0nHumxdMdzF50FBT/hr7XswbtvgYzdLJLDyfGwDnrxLEbyRIPuGB
i+I1D/6m+xkMJH8dzmS7DenyHrDWtByJaMlOG8H3ya1RcLtd9J5SokRMSHknWCF4
qlPvAeKt3mB6gXR5ARywDlLKOOp+Hbw/Dwh9Ww1DMoxKd3BULXyDbEeVlgkQKQLW
nExRJkh51CxxjJQKVAb8LUkAyGC9tsJNco+HTjzt6vkS6VPJG4EiQoQ7F7laYkJw
dcQO/aTB3sZfi1TP+OEIe7vAP8SGTMH4DuG1RUfXV79bFoPmuO/TuHHOVg8IvvOB
/qRTqTZcAc1n9xYJNp7YTpF4rv1SPBaiIvL6f65FmOgTxXZyFMW/a+qBX+7t6ZBt
RCTNwgvO3Z5iYIzMUlngUrKmO5iD+itGTNTDc7qP8Q9qhQwMhOHQENlKjA2riCjN
sLwQWPctVn6SJAmRPr2Y7vfZzAKjh90RTWMhyuttlxoZa/vxIv4k9bak9d7asjs+
7XgBtqNjoaEOEv4Xa4umtG1aXEFnN0q/zvq0btdwvSMs3Mm/C2/YlP9C4ORbU9Ji
vJ+y9/shvOpvOFn6fmvzsQ/JbTxfmLFNj1CBcjSxbiFA+qOGGVvgq0zVQvEaYz7e
FcENSLPcPspYolHo5geVRLCj4ajETUzwDn2b9jkoo7AJ7q70/mv4HZESL1Q3EEz2
zW8IvVwQkAtsA+RYS+zOu5nkeq535/rpxGgYFzQrV1IDojacnCBj/izCfL5OPyGc
ByjQDvjp/W2zzo56jSWlq2uUN3rrUOWb/cgFW2e8FEENiRVSXyY8uMKHIjD7oiCD
jDk0140wXj+3oavcn2D1K/ErPH9E5gwikTPQu6bx5G9RVygCGGlvcTG4KpEj+QOO
V7Z3FxIZlBNoDOTiEhQEB0LV1XEhHdOUROav8a+EpTRLMSs4QG3wBGVSj7Q52zyH
Tl+/SIDxJ5Fy6xh/zzfrjQBNLoWlW/NLhNJoPteKwO0tN3jw7nWUgpzvGfXQALVg
0hycL0RSIO4jgpfh5ITpw10rbRYFZ9vaf/FTK+WwTMZ9mmZG4a/3mXAcL4UC6Uoo
BOgU6+bySwURPMRDAUKxtxuwmU2oAsrAeWs71fzCh/w8OASjRp5Sx/4eYuYvY+Io
iAsJO5m6TBFqfNOyDg/DlCvCK7AMhwtYBAy8smrykv640C0P3rE1WAx7V5ZY34pJ
L/38TQJCH3oVWKisDOzDuegmNyT1FJZJoRJ85uI4m2QRNXFUMa1r7XyKYEcfhSYw
d/0KhbGHWg64/5YYEj4HA7atdGoprOyvLO2ZUuG4CUlWCxSbNoaKPxxLbr12iOZh
NBvRrFLZQkZEQqKFriOVu69XYbZ1S3wK2rlvTWJOV+MBffsNQG7zwZBm/8C3J08b
DaXT+vO0zGlVgttD+Xp25WNF2DHyHOeQVnjhiLeNPv01ZcrDyKiAYLW/R52BwS9D
B9WKuFnS0I1vEvIIX18piPVcb/iDQzEdYFx6bjYZ2dJUZGsZX0MlU5HPjy2i/iAA
zlsXjqZlG4sptNkAJvJ4D+hjrrRLkW8VCm2TknpOtWTswNPYZTtZ/gPoJdwPWkYQ
hEbYKPmol02ttYZTZdVs0+hSn2Qx46UI+2WKENUDlUAKsvdaUPbmVb+JtsFHl3pW
rwWp/DQFRB4eesJ2I1/9+1pANNb3XAe3eeHmo7NWYr16ziQs9cRikzXwL5LT2ndg
yPYdEfC1KjYlv7wlgGZtWIQGkoGtBBWWS5PJcBS+IVLQtD6HkV3nVP2f/81W3abh
n6P+DiCXCwVM3G4YDw68g5xDBuy3el1FV9es9jXiEoIoiBXTIYY52UUQHQvpM+WN
yEbSZKbHXi2YsNtiUt5hDHT9weUCXUkTNOkRd+S5B575fzWvIElU2GbJ69rE5xMa
a0U0Ea5HfUQyKq3uOEJ02bU1zM68nGI0kRDbu/8WGH1BIO4tWMimxOxPLTirtisq
+hAlm3nfL5X9bH+bk3wdJCj+0FIcSodkroeF3JGN0DsipalGAOa+LQkd4JI6lavb
T34KZiITXpiHTv46i5O/w1MSv9j5B1Vh3IZxSlzabAmv8JT//REqPQiFo5Y0wr9l
U7uF2mXmfFcn3KmoxdLA5KqITTALrfOwhqmrGj3Sj3cUAOBsHQWeQobC5V7tT4xg
S1kGgUcV9E28hatzrbh25KhMSDtKyBFrutnjfFxVFitO4dZpqlm0d/EP8ufLcJdW
DsXzWwStL6VVeRtXFmnSsIFk1Q3tqWHffRVFjaUfrx/X+v8wHmt3DYW+wlfHqqLR
xgw1kBdvdjwxZTxo1mLxLXHdUNFGc4reWNUjiKqt3NnMIg6ZLKyw9b9NSa1ZR1WP
5eeNLbCAYdjWZy0wNWCXrMydZ/KOenmrrBffRiO7Ph7KFNECdZ/6RtufnG2TWM2b
Jd9cxDxPsgpXoOfFM9PB8d1jy6SWYuyQaB/6r9BrNdoirb8Oy6q5AGK0eNOazsmr
48CFe9MozGvCAk9te5HquAhA5bwgVwjQ6Oby/Bq46XrEKmV0Zfq2YmVuebIwGaow
pLv68eGAHio2d8+jv35MsleBivrVuNIsCci3ujDSnEh/iCovt44SdPcHncM7k1fI
FEeHfpqQd5k8NMNf5S4dsgQQJl6jTb14f9K9++PMoVcomw88A3HFmk5vrXYAZxU/
+6rfKq/pzLNixKAz2slHpkGLQdqFYTULcR+6Ne1Jj59gr/CirOBayqJpc6itcmLA
YUWRCwaORPqE2JEiKekzh89DURVHatEbznLetcpqv37/OqfOhHnuCTtQtGA9djf9
IQW+iFm/AekAh0J4F31aHgoR9xAmbRiwoxpnJy9sN+64z31RmbwhFTjmLyhlLBZF
nScEtq3JJbcKD3V+9CPgLTH8CzHH8JcEAIZHNFqck8PZrxVAUHTeuQWd2zhpz1EW
vb7XAcpEQMdMp9MtB7ZzMdSjGpQdVQIeH1qHp7SM4kGNa8nWEE/FQch4cTVlSbwj
XjZ+/Y5gLHf7XX4cb0Qh0if8c3KnGw03qNe+8ub6FLn6HU/YU6fHUHBI4ueu1eZl
x78NoaPT1QAMI0tTh8b/3xx+qj5iJ5s/QxN+W8SY0nCuoO5rvezuPscGzL6QgnZy
EwHaCzwLX2JcpU8lzmO742CI5PxMslAoKodd3BBSyAAD7y8bd6HQ7iWhpGdntBt6
eFDGBFsMtjWlJVK/HvC5/Gr7/J4e1TB9K0dIMfDvQrS89OSitxiHDXKX4IO1c/R6
A1vPOqXFzqIKx+2LI5q/+xgLjvq7JuZtMY3bT3eAdkm6bnKsXh1X6TETmITCVd1j
5dxsnmOHYHOaUVAnydhWdgxasim2NB1uPhFcwCitZSN0QMO7LTiYl4ZVKhDRaaeN
fXZqTqijm/3ERL8PGOUXnlae2O5hQ1ClVuI+5pCIC8YUCej9RzWoga6E/oWemxmo
sE8AjhkASTJnYcCl9+GesAG99VFuHdMWvy74WBFCwRyyAU/VtD4W/Wu7UKwWfGHT
k5A2i8aM8iSZsDwK969I7T3AIeKjfN7ji+TmgeXiZeOMdZ3mm0xHLqOyMByJw5fB
0RAHPMzpS1x1cmblZQoYRKo4r6GSCKPwAEC9xKs3CiAmTnmjWCF/TMJ8kzoX1MWr
8DqoP3HII53uPoaKWKVwxTEIxL4WvwWw63wH2ExWS0pHpX0JRkO8ll/ocEx8U5+x
1pwkSJ+3gCxPLIUSI8I4vClfnTlTRGPD/JUvDxk8E4AjvutNn6qbcyRsZn8CbbUs
xy569csAw7J52Hb3vmM0itVDioqsrx5F0rMIycz648AFvPVVd3WGxnhohpU6lncP
0SJrrNIxgqRbN4wNDuwQSzJKKtGJczHUSSUKmQNQwRLn0e0JFUXXu2aFE9LwRROy
hapbQ+LWegIfLGdR8l7MpCT6kz5ViJuLjpCYMFRLmyiUBptSHxIu2ALKi13hGPV2
KFe9hD6rYuXoe3XmftwOnC8lfsY4Do/SOXp55erRwhm+bBlgc/VpjBRaPRS7r0cB
CcWg/d/sBln7EAnyu47oV/DAOVfJ95xWigzm0+FAk+oYW/3NgyQ7NG6msBeMTxCn
TZSyarUo2emwjlz+sFbsWWtCmFQg+PSh0NTpyOB34QzJnj7YtOT6YSyMh/0nPokN
4NlpqcDpAMx6ydZFbF42efNofP8owYbCoUeZ7sR1jucpqYqOHA6Won1+uB0WEbn2
p84O+AROCz4wl9kIjvwttjKO2++mAbwvD/m930vjnHD1BybH4ZSmJO6ncbcGd5j+
vC9wQmGiaym3X/UUiaFI9LlF9khVuVsbj1zZU75WipStWMBheIHxeSjX0p2hOSMv
ETGK4qToZ2RQrjLBxWta6LdMLSMM1H+B6dp2myT2AuT+VQvGrlElQvWGyEFuAWiF
0nphCjuYwd6ZhTLl8F9W5ZSo8yVlzJnkDnWgx91R2K5zP7w2W4JsAbX9HB4BN7Zs
2dJuiYD+W+XXop8q73p7K1VWHPCA3VciH1Xq+p48h4+eisW4ui1LdLxxXAXzfINm
kK0tMTG7YIPAz2FkkAm6+jksawKdFkfbVJarCONipac7NofQpCHe9H/qeIRAfdhF
X/a4aHjIx4vc8dqw0CJ5/tq+31a9shVDQx0pjfrNE3rokTkEW7fg6K08J4i/voEg
o14Tf+uRZNAxKKHVXuvRHdHWgivDmxwhwPC5jeHyuk4oqCXfkA6J1xclMmQR3vwV
fqG7i8QvwWEibtxUuaml94jXGmT4uCvvelG+UONj772sAJOFbkH2JzODcuO2SapE
oxnlF0bQKML5gfGika13epASUPIsnN+Noi16WK1t+axdX7JM7+4IuLAVaYnSaG9g
JeRZUWxY5C9Ul2QTmkVr9C/S16UdhYFx41qu19qoxJNZwPc93bGKCajbaj6rCuZr
GYx6s9MMjjum/tM5Kd5S4sbCHmLUTJ5iyibE7UAOf9OhUwLY50cBZsoabZztf8Vz
qvTYp5biY302T9Mv53hp853BR9w2obvot3jXdm7u7HYseGHuNXb0Zs3g02gCuhtD
zunGCB8IR5jTIeXOWoeSB7wPEfsN/VoQ8eQl0GdUmKZ4AkBRQmmzdU7+rLQNBt5v
cmLUXrbBsSO3o5Rcw2utGjK0ZFrQvUt9O5LQS3m9D2LQIcgAnn/Bgik9TSpmlu07
B63uRZyvwGWGZRudLSvsu1ovVazl+Qy1DV8RQ2CA2uZ7CREEE9EMrovhQdZEhp6X
Li2YIazoVyk4D4LEuRdsCHCmc8IPmKQAl2ZzrrkHNv8yOJu8bgRfOFzcPTdQli13
93fZYm/hQki7rTx3beY8dJXNgVnSi/qn8/7V4BTuWVr0EhJhSgRV0UJ3UyfvRRl9
4NM5vaVZSgt2wKdqhhP7ecwaAfNJN93AcpF4/7VJhjpRaDbtmYyfeMzUuAyIyMnO
`protect END_PROTECTED
