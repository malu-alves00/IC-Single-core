`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
r6ByS1agO+jgXy1napL3Y28seH+9pRRjFpnGdbgtkBYHLyZlE/8boNqfKKdsE3Lx
ZlCnFl3rHtASfxybaBdIH/YdFCovoEmerVzFQE/T/q60oamQ0vE+8N3RFbVi02gz
u/gOs1ItyekKY8eEkBkdTJ5GcpMrGEDptYfIsp6tdCfRdl1qMxouZo34cZRrtx/0
YH3HoIBLCPjC1M4UvDZF6LVZrQkclnk/XucCLPUv88d0sxXyQynqzA5UXDVSiTnl
4gNm0jSaKGx4DttVnDSMjjr3zrVk73a103m9id2MQvHEJfLIF9aq9joxbDQ0jpql
i/7maPAv47mMBVBvXHZC+FHAseAWPW+d4EouXb7Q4hdkCnLaE/SE4gmFgTbjGShg
v96G31hTyuNHlflL6NuZ7ipRzyhIVhcBshUZZ+o+Yh8plNK6+oeXg/8OzBJ3qovk
Ex0zSIr6HMZpBGe4h34I/isCmso+3uljiuVwD2w5LOO1WJ6j/Hv528oV1Sco2fMJ
so9YbVeYRKdIVXO0bNuKMEmUNFbX4V5r8Vy8UitTEzeR7JsivcT7OOEsGTjINijj
2qz+EvvOHmxciGeErmpVS8MID1HO6+VGb5aJW1GNC/JR7XF0x6ZOZ7iSl8ecWQjf
PHO33wy+9kr64MdHOu8vLSIaE2xo8AJ/y86o3NMrTnUVl/liCP7aSiqJbQ2v7cYD
FVXYGP2SQg92/IiEPXeoJ5/sfF8vBvV0z7jKzj0Kd+Z0dyEeWJRQaXED8Jcfb1yy
esivQMkL8Mvr85tXy2jcX5Et7IlFcOTvpiMKM8elWNlXpHR86S9Yo+uIMOp5rojv
4bFRO5Qg3c9iFglw0svvelmf2tp+vHnRKP24SwKtbSQUVmzdP5Wbkq+5GrN9tXTE
GE8xhQk1t6lUbv2prmFjh2ZPQ55M5B1a3qnrgAEHjuEQSDS3s27fKrnSzmhMteLw
gbdkimTNGfiRWRxMxytQiWyYN0aPICT5f9FDNhedFqMHUTvEsoxc5rsHefedb+2k
jvkZmowmLqchcJr1McnEgQw+UhnSfPy/RiiQtrEfFIv4CkwJKZysUXuF15+f+c7f
hjC+yJATslXBOoahgixMGMJh8tdqBYpcQ8suYd1ocUHwuA45BelBNynRPTwTiYhY
ck8euEickDgkXFdIC5JovkWke7+5uGXJYsbdFHIzftiDXuPi7ZyiT8/1bZ+tnm1Y
C1bBA3UMe7lgNCw6Y+aShh8JHpuP8kvB/DfsPgn4LkQ=
`protect END_PROTECTED
