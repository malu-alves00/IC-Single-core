`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
N0IrbnhjJSbI2iQXPvX3a3NKa+uUwghHO1w37BnV+dLo0UkvmRGmjxvM6shmJcvy
ji7RS+xZmSKk0CmBwcJGPrdQdZApM8L5ajKXC3RdMiyPj1G8WIXHf8lA2Uu5743o
OTlXCe2UtXcLZ3yoHI+XsZL2iRyDEJWSnmqwAqYDqlm6FtO9AxGE6BAMS3bsODWQ
gbRIsEvXPAEbofOTW9p9yW4E0+RLr2xprVIgz6g1/IaHKbtlxO58S5hIjkbHjR+H
kRLSRVt8gsSEXTvejgGfWGTWBtGsWbQsarnvdHN4XZkY0QIaGmjRA2CvQNfILHjN
wTAY9ybcXd7esryEW4AxK5ShpFVvg+jPV6NHU1oru8KbwnO2VcYvmGSUpWluLvCb
tlS/kxWw5kM+cOD1c2eA2DECPz5Sry2Q7JkfXYEmM2zw2AUNjmr+ZLd0baIWBUCD
YTgBmII2HMTUgczShm8dH1uCUEsylx870oCPtYeVjM47Q/HgHSOSG6nMf4l88x/c
O236aPhDkbredaMJrmvkwNX7Nff7Jhre55Kun54CPzYD4x3pTesb16B0bCHI08//
vhcUMiDKhBaGzRFXGntYbpciJiSa0nQuFWCCfWHmTI5EuWYnoFvFEnq49Nv6YmOl
QtL4k7pu+SkAvSuoYuxtg1pVYMh8gXohvSifnUYBA+pM9VQidRsfmxPfQVOysucr
NoZwFvxGkJYTJ/RaTgzVWB35cgc9cCV7NnhvxNr/1DE2HXZCUrN5+rQlQz2ikwTJ
SBONV4LELYTp5ml/FWPZx8q6TuZvH+Eiyl5mIMXX6USeOwUKjyNMHQvfKTBQ62hN
gv0AphsaV+k4eUuYZ1Wrx1cyiqlr4zVXwLRAIlWVpIJmYOVzA33LQLsez/VmhtB4
mgA28abXf2HUAMIsWQNPZylzQe0ZVvw+qmy2Ks4uy1jeuHuHn8+sijuting5lP49
POEaMJkWto0Q22a7rintmM0HHoTjg5SyWEOQJpQ0yXA=
`protect END_PROTECTED
