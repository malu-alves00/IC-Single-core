`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6XiBuP6ojaXZbTY+03sMbPSyjX/MicoyL0hCMY8LZrVM6L2GBox5VnIPkjnfeyix
39WNPCV59ISCnEId7PVRM3c9YWHxN3yXCwLMOJ7vMKw9+72FZhxCNjZfLqq1qLMA
pqdm4S2OkQPHmjCB5eAFj5EAsd2IUZ4JcHs9ig2iffcABLx+WOw/GP1Grwrj7rpN
vi9NDtxYEyBlhy/sP2q5P40L8d+6gMe1+y+NlfaGtmDvIsWGZGUnbrnoJ6e2uqbG
b31A2UhTNOQayY0tShGVeme7UkI6VVqdxz19YjTf3cmImf17kn4nB9/19uJsiOEt
EkZcfoYgO5kYktQt5gISYfV3CB5upZYQDlI61UFFlLWCZ3rC3Dpq84NzemlkgcHP
1DrTO/ghfyHBYncmyhzQcQgMOklCcU08HBdvF8JTQ4bNXSPZ3FldzdrO76IZkY9V
6Y6nnET7uCJsnbRkYZZSM3cczU3C2wXMlE3Z5cpLqYsyMvDQc2MSvm4YH45ZMVgW
zXNHsLjUIrEAYIkVxx2kn4xQ+qe8DphifR9RAgiK6xdtHGZZTvtAUDjdcU1n65Lc
00Z53uT7RNeCj3jcdEGkON9f7Umb5rJjwqWytuo9sxhBtDnDXitq4vn1eewyRZcr
nwpf2gyIM5p5M8rhaIxwKXcHwxaTSvbpsNKnKNjvE29BWowu6HPszjKAAocHZTUr
G5NA6bUQYv7US9NlWPnib/gzUebmfLKCmFhcT4j+o7c0P6lb7+Pg8/0JMaEylzyV
FTSeLaHflHtvQGOV+629Zg==
`protect END_PROTECTED
