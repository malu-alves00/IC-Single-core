`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uYEzXRI1KSbv1+Cm0149MrCHt0pgJRwlAF2D3EwuOV8PQMjUMpVEvtLjnCp0hOYV
l3ARqYZZXqkAzFYN97pmvs1gvP9kespKT3hbTNvSZi1Fx171UOSQP9iDZMlJKLLn
u+TXfwyo2N50+EQSvIZo+mGRygBEbzO/AbwibNMXYJE/sk4EEhQmWyejD8Ihyvly
UWWizZM7aubv+dyn77oIf7zNJTwR18EQ2n9Pn03lGEJypvh2MEX4JYakX1X5gmI3
9ZKMpQkvK2EdwlQwggYMFX/Vn5LsejpV3vrJLxoQU4dFNd8k9OroQk1AQYBXdY28
fhwNKWN37GhWM63oF3sMtrraFGG0emXf4ftcq8G7VqtOIVt51W4Ci0f7NwmqGH+C
39Koqw/vqYG8zgTGiSrkjBnTqT/koNXdAOsUi8q7VvubnQpZzWDUd38CPJeiKR6x
7vWB2HWs+a5PW6jc1RjQe0d5V97IlUbcFqaVjOmOhObt1P7EZHBl2cgWI1c3B0fz
gxWgb8W6oK3v3rif0TZIWEALaoJv+D6rIeRHP3mK31tXbsKF+jnequ9/uFj2WpJ4
b/AFFygkZ7T+zb1aY43P/G1nqTPxTmcCvcrd3cYSBclg7769RrPtgdMBotdOotbw
PAXOu4lB3ma4IxN2REn82iwUAin8s/JnGpxz83JPl/tM2SVrwmTLw64jADQ6fPq/
/3HLH/YwUwXdaJ2yKcluJKjmsbjNcppWF1j8C69LiM5+O1pE5oQDIQsET+/Geqac
ROQTfViLPcATaJ0brGebQnREt4SRJ9nURHQ0DYjxK756XadK4+DM0AwRd9959NHa
THOALjOi0rxVr9T7WJGLzFhSuwcW8Uo5SDLTIu07ipgE5Uk2Ql5NiDRuQ4wcs7Ru
uNjwpzs/9qfNWhobKY9OqM53IFFEiR6KcyTuVQLHYGv+Cwg4mmCbfnhIqwK/fxnU
QAmoej95h+6GQNzVdsvw6SRH7UuhkU1yTkT/WNrbr/5+CCFQUXy1EPOHTSQE5I+s
W238CEfc2eP6l26vpkefVjOYEjglqJDXCP/iudnv4yvCGUlPzCoMG4lacduyggEk
SY8IZRHNJ/MjOV0e1dRGR7gFG5WMNoEBOR/xRYtP5zDopg6rSsZhpbTOKxOH7dks
0M5PA0XbaOJ4atxcMkQUUEGRGGMt5fz0mUtHi9YbaAamhUrzzrVmsi37/c5T8Fx2
vV9A3fDHKTOquZ/f8L3sKJq9jJp/RqWm1WEuOj05vx/9oN2sResQb4SvoeGGgcsA
/QraVrFhh8ey0k9zHMrG420A3dyiAsrVxSAbesfM86DOFPJhpWZbxfgsZC/QHZVE
ry7TdkykCBD3zkAFBQy+CCl+VYNYKediYrzy1KEbfeckdAAfkhIdV+Y3FCvXw7BA
q4WWmhSRZPhM1DoXsHlkYPqN5Hs1znYkK9K+9TKOiCYpGuXtpGeP/6jc8u7D4szl
Xm9UUS7kRUMMHWXenkV6uA==
`protect END_PROTECTED
