`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JackzEDOaz4F6/dobHDrJ25Ym+1tK5TgkgQsysUBQgcu+dhIMPfYeipR22TKgXxi
MzjcXmCOxKR9R493wQw8AQS/1uLZO02UbHtM2JrPVx3mPJiY0TOWQFOHY9hzFJOW
uBq2aTcp95NrMs/2NXuiktlWcz4hv34ZobIT2sbkzZIBzH/XCWUALt94/mbIW2TI
wIUaOjT13rAVZHjieECm9nCMzyRTTZF035CJU0KVuNRlOfWUgTWz0lzXLJBs5QEh
MY+zSamCGLORCmBFReElgmNMP27gVNpBYVMl2OUX2PLz1rRAJdLPSn+Or/+awht5
KzeDif3wqKj40Cc7CpEisZyun/j6uK1zVvYBMZ13nbB4MmxzyPMMpRKRdnb5dsER
9QLGzmHVwaw/P+rzfCqulqFWStYXVuCT32x/0CnsRAhU0yR6qpNs/AiCiBN7tnt+
a17nFkgha7ziMoH7ziWWI2xe8c5VjyfUwaGa1Gwqpys4NRg0Qzqgrsixc3NIb8UZ
LYfufS5G9Zcz5KGQeDoVVBC1Hj0a2cX8tmKMHW091lbyUbtodiZKueE3uI67F/RS
F2NuUMrGEQtNNsois9ymsLoN5EiWky8YnWGHwdQx5AcNXamEdYwKRe82KbiMdDHD
slHOzQDGjPBCnCatVdC/6kA7IipmxMoUJmUkQ+wr3GtdLyaddDMptVLGRuMKgjvt
kfdICfdnQZgBlwH38E0rt8haKBbT1lE19agFEeHu2z9sHRicuxWODeAHezQbpPBC
U82GIeuocbIcWS58AS/ETbAI/WaZq9UmPSqPYOYnEIilnlngxSnNSxO+LPtB1SF0
ETiTYN5unM/BN3prUdO1KEQnAhPW9aT5q9AsC6xId4u3Ck1KBwEIg3voPpzcpo2g
uXPDxF/dzWRrV2GEjQp4bp/yeyWUtIQTU/QrFEGQ4d0pUhlHNUMuJZJfoWT4n6ZS
c+o6BYPWao4sInUZ1DtZamCCx9Vzu6AIqfL2Ko4dl5jvCpY007iQAtRUPwI1+GpA
Xr4Aw9HxrYbx63z8UYTqD3IEeGe+ajfW3G6QeHSj7y+6k/Bo8S3VPAeFFdOrQO2t
fALEsrtfxJCjAkAqmuwXMSj/NHQYYMZ+TLwAe/L7cPsB9pSMj617evQoPMfYOJ2h
36xeE1/mG9CxDCIlHLNZVgOZrKkDWk1ln4GKNd+R/98D0NVeghq42kJ09nME6Ig/
N7RRNGDLDpaiOuvYIQf2rU3e75aAlGKr62JnkNLK1ABeAVpkfqhlbdb1sAkIUGaM
GwyUqi8ElOv1n2za0aMPuScgAqFeoW2oQIhYV6rqFhm/YCT20MwitM4sEOtYWQOk
6SmurYlSTl3dbDiSNDIt0AOrg/jeKLXwSREBYZGU0sqPS/NZWd7HsHlf/EaPa8/W
9CHlvMyRbA0PBwZoo0A+t9HJgCXZmGutbV+rxQJCWsyKBz/zrhVephHDFS8IT6Nr
e25tKbn74ftNHW+nnBx+90My7ZhVECxRHXyVq23FjsU59Jrz9eCZFyTfU7nJC5cn
DAJJtJYNDYAcX5a1z2yxO8BXevqt36JeY8jDTt9IkqxodzwUFWG97xEmI3JCjYH5
RtEfDuQp/wVceLz2D/O/L1vAn9a7cY8PMMHXKeT3mx3opqknaMGnYkwvyCDUpyTI
Q8x63L7X6LVY2fhnFm8hJUmpP++hPUhN9eO/lUufK7DtCtLTEEk64ZG2xLY5lsBW
ApHRMLNyoh6nV/uqqX5ma9GfSolExWKo3DvjUuxEfF+qljDffQQwrwt/msBAVjP0
IFtuxJl6aUMyti0iGeUpzH60FJFoJxC5wc5tLZ/cc79UImV4oIbNJlCnmkZmcJC+
yz24dxctgftQXYluVkijXUXArSpxwQRV2Pdjr+RGsY8hSbp+TAQXDnO4/1CLj0sX
bidoEAbJ+OEXCFJeOu6C7SfXVKzMkmoW74DRPYYbv4NSaBtJqPDVpaqejEbA1+mU
8DE2T00dH1naQJCcOfn6z+pnR+bd0MRRmOwg6r5QQ0ZlQ6zHGgJCtE87Hk0BwDDo
5h2Bn51q9dvXYv1c4dJ9Bx2mqgv+4XEqA3T6Gzd/8nIEZsuxPNqZf/9mjF+esSWM
vRO05UlJa4hDCCiVKhBuVc0P+hOO3+N8E4uT8lkHBSwctqAN2Zn1oVuEpQ1F/DXY
YsXch/KiPEAi6KvgBz5Lo0dcLUPkysnHYL7vq7cMxC/J72RvsyzvVlo+lcZ2vjPQ
zi+6n7ehJG0hxmgsUYBA7VGoi20/QBWattzPRgm589DVXXAiCFrZ5P6m4VYXgLFw
mXeeu14E9vddgiMpXCowTIHEVvHYJjFuukHGpEalhMw=
`protect END_PROTECTED
