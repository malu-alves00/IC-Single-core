`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bqZMjWHt+WU0cm6tWpGfYDEO7LaZ19Aoxr+7JTCBG1KHVLiAED42mJScpFlZyJr8
E5QttxPPUhVzVOKmYuVyMrBA6llUHRj8VmsOxWXBHGtsZnysJju7Yy34zivcm/By
jEd9ojdEW6lW4H4Gu2U1BqTN+XWIjevULZEmavUYIc3DIDT6ANF2wup8Wyd7Ejzy
VqtM7uDvUU24b0fnklw+gupduv1VoTvryV3UBjxR4BoocdpzuVajkG4wqzc70k83
eKjrEpK37x2dBNXCTh3jqbDJ5FvaM0/87WOoA9lnshY6PDyjqtr9RuDXa2g9tOgE
+c8s30wLz3yp3xe9wPKIsMk4A5limftMFVBAN9kbn2KTKod3dficCyOGIiMXoZDG
XdfV3PaTnLBZu0T8g0S0ObjUIFPx1AmeAQ3UIlA7IHSQMbpf6/JNKDJjpRWQM6JS
KOJ2R6pNr+/uR0JJDoCqJs2DWkhjOFTXus1tB+y+R3ZJ3eEvAbtSJYS1fyws47Jc
q7q+8qSfYaS7U5A7aYJ3ZOWOeJOwExicQ0YuD8FJsGaLJ0AqpjpIuEFAv5Pn3ZT/
V2o3dYwdPAJqkM2OqWLYESlZ+RUuOLQmOwUofk9lhSadLEqn8BNE3Lc3iB3jXlhM
6V69Gg5SL+r3NW/c4lYtX5S2qELrAFvy4m983vlva4DwIyfXjWOGZ15/Z50bBd03
Fmq9lgFt4L2j1IGzt2uRIXP4hBLlgYTtnTgpmJZsc8yRieu0Tj0+wkvZd5dC7y/N
I8gHb40d8h3bjFqc8Oca2N2eBs6X0YvHjbFjgP5esj3tR2I/pieBi5XFFNubcDth
q2LPcxfNhN1OS4LKu9iyqOoqFL16SwfyfeWcqjOFGvoFTqsdsJ5vX5yFHRiMknzK
XWwFJkJH8bWt9jSnAJIesHzRu78VVGXAohl6l9whgAc0zC4e5B7dMFy0V5TQDaZQ
VQ1s4vpKABhQ3quL0XV6LGCuEPpRr98FphDx1q3BDz5mkAc17JCsjOISspmBBu06
Fcvuh1Uqe7XSf+nY4NLCkBzNC5qinDdDS1rI2fCmx5P2VL/mXNGb5rvqffvq5UIB
KJ0Izi4fuSfRwfYk1mUTPVKImYOfqRXUxf7Q5kgIKsBVrpSKL3Y+uDxLkjg448bs
EdK608QimV+6B1yfnLfaSoKOWwuYF3pfu1hbXQ+2LZTfX94b5HEXxLsU4sMsuONT
SzJR8PbAVfta/XZwF2LmXDAneCI2ODd3hgaN1Lnl3yuMNkRisECqeJGhg8x261tJ
6qcBkl+eKuQr7pOvZn9UK3rC0U/P55pV7116dAg12sGMVV+NKuIWmqSwzvx2BflN
v5/6xsnG6KyngXBKTntLonXK57Ge/VoPa32gPkitykVYrdm9aMd7IrxcZEM6CzvV
pUtrktMko4JlRP3vSh1Xxmjqh9TubJuHMMusdmWxEUrdWCJOaWhQMxPMIzmtohoK
x5URIWMZVPQPliNtmjDnpB+j9dqPcOhYdJaQ5zWAVLGyeTT9d7hw+L8bggPU0OCg
ijRWBPe5TL1N+IIHLurP4DW1yoOMbVLqbMLU8xkZz16EvyEax4VLm6/cWfBHm9m7
0V+gUC9JOLI8OqdvaUxXYfzhXKY6CsMqiMrjPIwTAhjCVIWIxzRZqMkNkjzA1MlA
2pBbKxBn41zjSiAhBVTXleVuieESiQ0kQkO5P2/LG0ADasg7dqx7Y+JPO53MbUPY
kAJZEK6wVCfron5l4wAC4UCpRa5vapVQ8q5bhI+8bSp0Xce7dSMKqKuzKqwQf3CA
1CtGS2AuERLT1YC4T/1NSDEvc0f2zSXwQjlfukYj5wQS4Tq9hWpkxChR6SmW0RTw
DMiodFyXo1mBNG/gg6M0eD2iTSV3M5jRFpKHn3RmDEFy4ljc4xLVmPWVgQ552ybX
mvfQfzo6G1rmlHjkDiMz2t/PBQeluoFZse6lt6KdAI0L85BvWvEGovkThCRfeX8q
fcRgbMudPj3+Wh892J4RysMSvg7D2vEBYn8TOQUAi2imClplVFnrVjX8rrYbJpSt
16R/V71EVrM+L75Qd6DfXQTSGzVB4/mXZHrVBLLh22GGtsSkNxL84s87BnjSKmus
OefPp8JIyv6VoS7KuvjmRVtbIvGy3Dddpou8xyFsFJugxivvRE1RUNi7ov1uUnyk
SwWHlQ9Lj9/XsVGaGWfbEHEki9CJeYsnkviGXEC1BpsdZ0oT1jkJ9ajdLR6MyDwZ
DGV1oRlABXkdsJEOSZSFvjKOqfEwA8DZLCn4hUU9OToy99SD2te8jJiQAsQCNKbp
eSfVPOfsx86owDFFVpBw2DqaR4vnfQpg+6mabGQGuZGW5E2lhRnC8YeNx9XjWt2Y
p82ns9so2SdtcXoIY7dTQQ==
`protect END_PROTECTED
