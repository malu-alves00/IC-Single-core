`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ufIEbV1bf1wPWLItuIJq8HUgXmyBpObkM7mGfce6WFjZiUO2BEvBOPIJMVJn+JYX
pY1fnzYBoPDkHJkgwbukbRgbG0fEyx/C8mnt/NKsK5O6vnKxij6er5d79cJt787c
UNXh3ZX+GoJWtgfQk6yDDivBonKsaFhWzqCXGzzphEBdZnyDDjJ+I/S0BX2e5XG4
vmY8jdJ9oWkMuct1MoD78qwcI/XDcVUUqWppzGqDTq6a0zSaODC0RrB0VxA8QDiX
0nDaXUBR1O7ANG+GLoS9MIZaWsQ+54jop60nkOpKXSOYa2Qfrd7t0RHKddsi2c8C
scwCXP5v6/rBMwNcaW6dqPJqhQAFvTtJFf3pr4CNZqoUx0l0H3JhL76TenaLj2R/
jmIT/JwzMhvrv2yLeAVNNX8kc2/GwLbcFpyp4s6Nd0yqzp4729sMU2c37HH3p30J
FvmgtZE58PdlmlMh64lLeJOyMAQi2ZgLjtGjsObSmSLgMk1fT4R+qMC4mlqiTE1e
8g44PP1kORrWJPa+J/EO1vhLxbUUaT3iwZbuVMRGq1pLCbSUOVYkMqL4pSqN/04p
/sFTk0dhP8TX5/LOQ91pbpxFdH+xYH98bwzzyF6WGS9JQaEaTcgC44vOY+9toyn4
Vh2372PmiHHkZz+gYlxGogbbsuP7Zm+K2meNuZiWWYEjxtvKkJeORKdTQBTGkogS
sDn8uepZo1QhV1VhSsk4/MGzORh4oz4h6BEHsGv0pQeQ9Svbu1ic/n3hmqLrZerG
KLMnX48F4RQ4quHBCr6vk9nmz0tQvmBdfWu+mUJLigDbiVXxlkX6vXwEbKisP5Qk
ZS0A+UQO2A8OOFjnyu4H+EiDQsXnUT428DAxKXHoGdHQozjlEo+ZdwwHL5WxXETb
cxe7GqG0ZfnwuvvKeRlzw7de+5hutrp3ryIco8Sli63A5+Va3ft6QvhNwKTUNAig
oCj0uoo9a4yCnx1lrMiL6to3le0QDb7nzEircg+sItfnPP4iX6emEczKw4eU7c7D
v88PqAuSS4PGoULanV9TTUgBten+NrkXzGUaZU24pq8ztctbmFJk7WgYyWyE3SVJ
iYZYLDeBKDhlIEsF9006YQT2JUOUU91/B6yMKiShDXMn+MXLNavl1COUkcXSNtRn
i/SvZMfB3OYgbDa05B8eMjup0X5Ena9tyJmPspEQJsLJfKVZlPyU8bvR+C3VZUxi
Q+2Aqj/3OOvTE/PbgamKz1z9U1Np1mlWzFAtslRjY51Kp5qqomuRvYnI+XmiDR7y
4GcWbxjbLFpDZ7z5rJV83/yX1mBX8D80dRXcFvpn91TPz0WC9IqyHaW17IVvC1P8
XYvBTGsX5rC6T4t8ub97TY525E70/to2GogyjGkfizwsi5N2U0WHpR9JPwnyS+Jm
L5y9ACObHdJ6z527Bw+ysOSoHnW2s4DwDepC/XhQjkr2cjFJgKi93C6t5FTmVFNa
Awz/mz4Af3rBAg//iYYu/KS0okHEvRjBFN5nGcbqq4jQi+ldil4Bxj4a2CbliTgx
`protect END_PROTECTED
