`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zFOs96ailejWQK3cgB2sgM1Hp1fgRGPniJtbdBijpQy/Oo7wkAoshUXM3IxBUjyk
iQS8LHSTccrv8qljh6D5EvZjOApmZjZhZgMi0g/JgmQfyj1bFLSTeB51su5aDB8L
fr9d7dzF653FQog9VMRUxqDpkGkEnkHIXGImBf5uDhGutzDRMHo8jq3zh0p2Zhg3
sPhMsAtLjo5NneOFXxBcdcHc4wZdOj0I5CWkIAE/dOG0OHYKfEoO7xZxSgnLmP2D
ik4+uZ5O5LlC49KHMzltwGbi7ZzXfrzeX1PTnelo2r2BxnKFc1GWO7bnaW709wVY
EM8P9U0y/74IFc81qNV7JZoIhG4k7HQJvXQLiKe25qDUaAcyg1+Dsd+KBQ+EiQBF
PN3GwwI8I1GPV27AlIM9a1rZdISnuO95pBkgCknUvrIGW4vczUoXcfuNwNwhEvsb
NWJ7DUk/qChMtewkRRczD7QJs/CO3CrwJMltGOhT8Dhw0sQ0l5hJqdBktn1gjTAI
6TKNWZDahgPtkhXlzXGewuatXmcAGT7rO5AQwB9oWI+xNS8Z5jv/Hi1qCOYd4QxT
U6u0TZGzbuaaZ9PxTW4I7gbck+QRmzm770LKJoRpy7g/4WBDC3TE3R58aHFGe+us
FY/I2A5wkqkiyFxyEUhLg6CPKoG8UgHiiswes4NEm/OhNnEHxWy0I5GaL6EKePhf
y9wrTJR7ZxnQiTBrb8G8eVaEXE87X4a+4CrKLFzPWl8oC9pO1dYh13GzFSD66xrd
KEx2C5C9SuQqewQiyEIDXCiOd5t5WOlRwVpXGO753aEEaSvaQwU1uItD2nvnYIFn
68RYCn+ypqUESc2CVBXu+eoENdmSKpV/ZWdk1UrDi0uTWJuJfgXMwp48xxzfzDar
mQ29wctBtpgujuZAro9hhUleL/HwTgHf/2HAhOGbpn78CNH59yS9cM2KHzkK4n2T
WdgfRQCFY3+u25Qtnxf90PLpPhranG+Vz491d2ljqmbkkq3MS9LFd7JDy4vzAVuW
YpPc5aP/uBZ6SIeA820EZZxNvJ2VOrbC0Xn3ec+m/CPt3AplF1sskghrp8wzKPlJ
R+B40p/5NOUCbUXKreZgaEJMrDFBjqqF967ydyoGLxriWXktI1scXXukZJoc9Ls/
R4Xo27dqq7vq+xXoqk9ph0V/tmOVSJQTWLwdnEsZc7iCl1aw0C/KVnIe5K1LNUA+
bdG6V8+pbWIWzAwpQp/Tk58kHXUW+IeXxu53P4lycngdWm5X+WU8ikz2uMj+dt+L
y35N9h02lVNwhGzlX1ZkXvVg2RdhnriWFgySY9E8zBFRDj7iHSwHksvFs9IgLBGU
RGwVn3A1/FaCdTKiiEPyDOTIn+G6Nm1nj8eZhVZmkI81nNM9IThcCxSiy34N3ji2
ZIWIbNqEtz7Hz7aJkcFfrZFr9UGr+W5shMn5rNkPYSGv5LnlW3b4iZTkvxy4uns6
XtJe3/s38xrr0DHS6trGZG3azv3f3H6ddb9523qUda+4Gqu4BEKu01bTfrwov7JW
LXjRDz7ISEDbQD8qjsbA9RhdaCmyU+TMoRN43J9IfMxChbRi858LbkYHejnTSvGb
Vkmi6XVJ3ptEpDQLrGIBxM1FlacraGvzekOCUEzqlBTif3XogBszapTn2VeB1Tyh
a7BfZVPkwUMaZeQLf1fzpWQCzVk+PGvFD1YrJzszHi1t3VCh3AzQrIQeQcQwGbe5
GIFnS4uX7LXVq2ypEkqE3cfV6sMOkwE1YuXSIeY4twSj1UEZLgBEP4Udb79ibKl9
vf/+WEu57SrYd+Wk0eRyaTU1yAmp/BnF9cbE1EDVbIJjV451zQ+UrOn/hYLJh540
tTCNWZWwcq9cYLOKWZU/Z7IypRw37li2luWw5aNinqFBWQechMDPPpqRAv2E4/wB
fN7oyDdf4ulSGVijmiX1SapI2JPgEZcmV3uUVqgWK/XGmy4OiBPNnmgR2ddwmcpa
InxGfkdFxZqbyEUawvj0uxiu/JATMPM65sEf60NdD7RJ6lyvenoGVa56RrRLh8jN
10+8FmJ9mJwIIAmDZZbvQLoe+xOYQcqeduse9ZMJaIPqNtRpMd8XLCW3JNWHUkve
34q1nOAYxPN1HTamYRJakwgHFxippLTrxo4/p65MKFgsK/0OAeK/1Wkpviro4349
b6Vc6QVdxoqwQjavyxb7RnDBCL6IrLMSnkTghskl4DcZ3S0ABXsIOeYSxmcqIDnK
rKGnsUKlgq9mB53VubNZFSbFIuJkswi0TwNbu6HvDOOcWQu1tM7zGzljjnRz8FN6
Go+pxBHbKoy1kKBnFfTw4lWoRzydPeLno+SE1CcDiFHsobx1BKbclRJFJaBdq8fW
E1UQMH+ePzX6S0y6Cq+UPsoxULs+HbfdH9hOmPDxWUXp6VS+R21cQ6WpVKMhfJHU
C+IQf4GoninciE8KyxW7dtwjN3lJjyPySG99NQlpzyGX3sdgTW4o6MBQ/WNwE3EB
mSQjVLdd6/0el9zNcX5hluMMrDNvhTNLzwFC5esle5iF6VYzTazTSXK3ba0vdNNu
sk6NzKa3b1lMe9TG0WbdmhfS2MjAHx4u4t/qqH7xSm+CBE+bDtCi/pqqT8LGr1pg
gLpwD/w+HZ8ZSPxIgikE1yXL8bgSo11NBZeW/9RxBYL1reDr0Ie0Ojqfm7NcTAVh
zK12Mg5nFHheqjKk8CsC1uVsMwqoPM6vd21VRDk4GWh1dx2pMrvPo+7ZAobTTyLW
qQdCRrRuMJGswglvxVKlpeIX4RlwnavyLsKRGYil9IAD0RQvtuwGMazDsaswUMJa
wPbp1/3HjKmhZA8GXAUt9Pu7HpGxTFudqbt6k0SiO1NtBks7hAYHsrfMqqHJc0fy
76Hn3dbaE3CdsEV2Ca3wJ+yZKBdbrkdYijTV5I/getkjtuQK+NS2bF5aHcoO6zqK
NpHs0tRnufPxDd+Jy3YkoL7x9FQYizMm+jKzg17QN6m80Gd3cb2sfXZo67JWkMR6
Irff7bdam4+TUZ9gzMhGoQJy3IugEtBMtiaIpEGG45qKz/9WvZt/3AxL0h/y48fE
Z6uV8aVMBR9OzL/tm1FjppRTzMsgzeGtXPp0K8ECzSg0NGZ164jTbi8afH62le7x
f+nqlBCyxK74XUEG4VX4keYUxzL2Htl9dgb2XyvTVsc6PTk6TSEgKoWeFFbTQQJq
Tdc+0+r0CVhtXLINPH9zozDCIHcc6mm9T5hoSPjdjkel4OKKbksOvvh4CvXzm+e5
6A1J7ri+QZ/JCdqpfChlW972lS0ckNcDwIMi3h0H43XV+gzocgIZSL3o30ETkaSP
2Muw98Bq6cfbDJ8BJDVIOM6bb6oaOKxPNaDe1XollGXgtwnQOOw64rq8OeecyDuR
6xR5MhAj5N0SoZ6A7bvb44Kyzc77UASjwg+36r3tdoGeaN+colkHxSVPoKhBZ8LM
0K8AjzRLcLj+N7Gd89O5BybFhE1rAyeCYOWWQx+aC66+ZN+ZAalKWpqYB73R9fZ8
hRYqFudinuJsU91oALOo6GiOn5UIfBsT/5vPuvQoiZ6xFr5twF03XdI2Vnxv19sK
wlBBM6y8G197qDdJplhv9pmdIEsdUXMCdl5guOf6x9HgWhOeFRXMWr1hSJLQZaHO
i70mbTyDOl+wjFbjwgDCPZXPkrE+MM4kI6W9pje+CNrwZCgx4IAeNWs3Ld/VAjHl
UfTtvYfCkfSm+Wp76T7hZV+5p8Pn6EKr64OV5lr+pO0WKdmsnuwEU7e13egj3g7X
npp2wfy7BYuurB4FpqJGwrva4BgpZRWDtuNgvsq8mdNkeOaNQylUMeTVzyVfv12u
xvUz+TrPqSn/2PbsYnD9hQknWu49Sp3MNQs5S/1jtEjD+RKmxLGT4vInk8/D4P18
GIpVsDnIR0c2p2eORp4AagGlkAAHYMAVwe1B/Vu223bdxNJPaKRXB6qWYR+2jBCJ
jMaYo77jE47tkRx2+OXgKEm6DQ0dyjMokuBQTdHwhQJDDPcCqFwkz8jhKW8JzOqy
weiKLeUlaSZv3+qYgV564D2mGPYbcybHBZDj5F37CgTb721eST1T2FDU7rfDS6Qm
OeJaxbHV+qFN1vt51Ghgttr6Dx1aG8UtGg2hS2CBOHer2dJAhb7ezr+S6lY5p0Vt
6eYhemRrcRi4XaPewPf9EEft1T0/83qdJMqk5XeRjMbnzvHe8bGGGFYo3OwBi81R
8uoPGmUM1824D4lAnL8V/A42JV8RClFB8Bm18G2XlnBhttmGGoTX4jajXRhW5hJo
HI0Kqw8qe7fUiZd0ihM9XOl9wPZM553mkOzILsvZRVxucEWL10MEGD77I4jMnhgM
UgT25NUDRRLKsLLP670UkMhapyc5r+XI3lhPAovUqU+4w4LJ1toxBiJXlyQIMELl
dOb7fyZqer84tPRMmZjVIJqyfK771bBJdGsAwiUoSklz0oGkJ5XgnvehB+l4UzIH
RWSux2bcVICiM0aTkDh6vxaDDkYLhhdZUzlix2mSPAhGJDPLLUaHY93BEx4b7cC0
ye9VCKdCK3O279OXVImv+DH96cJJ+oiHK22MOSMY/5FasM3MgyAzJpfbJLmzv2QY
p0c/w120EM0nXf+t7pW80IvgSTOXstyMrpHFaVjpF7idxYXL7U8TfLfNrtXcqQxG
YBdQUicCQsShSR7h98iH6mI9LJBIxQSi6MlZE3Nl7ulV1Iqcp2uCKAsFho7ge+Ix
DAZjkdKzPe//Nt8A1NMqRipSfPeormgdpiS4CCCOmBsol5+KHTt7j/IZQKjB2Ud3
iBhj8+F+5XbN74ky9KST5Sjh7y1JUZNCVQvodp6npeygDtebYtUnh6BuxFmgej/u
F1GqQGQY0/G0+aVHpwkD1Ykn4b58WTOkb57XP8Qt31xsl/OKmeGx9QJ0cLMwjVBu
rl9CxYmEWuwTskDL6Woy43spBx7zC8SrleTPdEKbogichpj/GLzKQfLJmD8I169e
1h8n72qUmkbIQRSngzEQk+ys1jNrbmtG7ZU7d3jrJCCfSWvJ0xH+u/MNivQ6WIm/
MUwRIE95LfTbibbOQ+hVFBS183TVEMcH9fey0ZLJAQts11jrO7IhJ6n38raLt9T7
ZPvAW+BJLJ1/wjCQOyvf3emI9ecZKHAuwBnnIdPxoZssyB7bDs2+eKBPocjLZHRG
YnHNi05tTZ7sSjUfBEokSzNP4UdzFRfUqomlp9rZCUSwNGTO2ULAZCVWsMJG6kdM
7bTppi0qdQv5B+Neq+JRPfaJcAilfkKA5AwTsHBHPxNjFpTO1+D5+SQZJgbFZBPw
kKMNe2XPPpvDS9vQWhk0Xmz/N/XGP13pvDm0kp3KpDjDdVsNrZ2GaLq7QroyUq4g
eY9V55RLT8Gbbp/6mJFIFUT4q8uTJiwDbAKQsZlp+PpYzRTsw8z5ZKiCvFOZ07H1
H15q0GSkVVIlb2L2NbDTlVpqX6l2hmkw5dh58eptNA4EyL/7sP6VGrMLvre6bLg4
0dvLy8rvV+s3GnNeSltIJsrHdMLU3yptZ+tYUuZFc3S7tGXGkK+Vkqi5HywzmOMy
2xkIat/U3gFSUl7UvMP7YQbL0wws6X6/LUJ42FsRvCn8+nSwkiOFRmV51MJxlbdK
DksRYc0khG30figIim21cGpLNjKzarC3cKyikiJ6KPuWXOdt37cmfbxMp1besOdg
UnHhsuL2SzBHLD0Iv992uZ0bBiSmweflolA5hwFSwOtzEKdnMv++E1CBM5uYQ0Fg
CI09R9JQKlC58p5YpYXtxFJPfNbvkOfJDUSulY+2oPfbQu1HhdBRlwR+ASt87EDs
iPdYBByRYqexSc+OPtbZ+j4XlKNikgqT449CsPNQlCcBA7AJ6fQuVb6ywjl5t9Yg
/mNKXk4p83b0PdUzbtwK7HUVP8NEvjBZ00jcAC2ZEwGKeO4gr5t02dNPRlJKRnZu
4uhihmppvvCFlEm24U/tkTXOghnFok8egj2YbVy3AQt8bRUHIBmHW0XEM5TE3PzH
H90VUG64jV+1LI/TIVbfBrVOJzSWHVfLtjpQ5nxMgKUEEHl/rRVeWY4N59fCjqEr
FHPR1kAvYir81NAz+kCJGHab1C57zzR+X08n5sEAMeuA1NK16qR6XHV5zl2ofQuz
ERX/1Y96E7oOvPV8NI//W9y8we2Rv3pNC1LTyHp7OlV5Zjrmh0zilrZ3x1PQqJFZ
0su/IgSkaxFmd2biVAGeX80Ji58WHRYTC4afei+jCvpePdJkRaWLnSKSwSoNf1H2
+YxjuCSitkVLivf3vxTgbupTxnNnN1+eUxhctn5YBUnP3X3pS7Zy4z/vzYOwpqMx
NZJ845sbnnxpyb/VwRyHvBL6MISNkEv7uTxM4mpzIq6MSoHqkqv375vm5d4n7sc6
gKe59QtvJ7u8v9YKHGYx1gSZZOP0w9Y3Nl46/M+tEMqFhWKXL1sgKb4pw3Ys19WV
Vls+bEI3tXq+NG1SVYiiRtG0TpTYT9mcQVnHst/cVlotVYOkkb+P5Buv5TW9pJtp
V2QkjiknNBIArAvEM++THz1P7VUkTwvNcpVYsOc79Q2VWAvJLBVOiUyUfWMQXX3S
E1IwwrxnN6ItyYdWrcnJgA4KoiZ0qfI/n9CtDhTB/yWuF8ahGGulATPfQFeQ/aDB
dxfeB8RANLlsgY1CdMCpDckuox0g3UUfYjuW1rMRl3X5u3dw8ihgkG4ob4wfFKKt
1bsPR06autRYrWl+PoHgdPCfn4IHDf0mx+7KRiT4WYLFu6ZpjZ0AFTR0ZmoVQW1T
Lsu1ob45AGo68a8rvWAoKsRcordGwoZb+qOQEdAsAKP4edZSoy+SDvC2yC+wHFng
gNrRTeWbwCucf4iTSi+/VXV1LJs9LKKbCuBD+XM7eKaD2HBoWpgqtwBArnfYRrAv
v7oyrtSd7b+tts2ZF1P4CSwWV1e9PCGV7cmyKJk9KH0WJ5M2+u2DE1Jr83UXZVw3
U0DHJd+vzcv3gsQV2Temi5w0J9L5ZUJUcu4MxjChKAddQz0sRwE2ucdsnoe/h9Mt
B7Ph5YzT+VMT7xJOhtk4olf7K83f7mOufmop8tjGsw/l73aBUZT8JyFLq/g/rs04
oQ/jMQD89395AWmD9YyjxCkYmO9e8geroHyyaei29NpvOV3K41YhxFhOv3w1/+JC
g8y0a98aZnck7/0uod2LeOCS4N775nJJZklch1ssWGi5Tt7Xf/9wfq3cT4cZqasm
Fs+S+aQmXfPq6QC0W1/SLEkJ3vt9AiPUhmaZvhsQrn91bUxlcBu9xz8hAHRYRJmw
hTRH/thW3JZ3jacgiQEqLY1gBs9BcPIat6yf32vnEFsDv7V0XWRmBmrCLTZLT8uv
H8F90GtKmMBnN68VF1wI8PvQo+Ja+jqHp47u1XQXZmx/bDDxqzRkLEc7yvGlsJ+G
hJeAxQbnK6Xg8o3kSt+wvxCuu5WY/DtR9Wrm/UIoOdYdWrZIrVHoyAhXKzgziIiV
J4kp1kAiq+E0FrpgxBRg3y3x7/C3ywtI24vmX8MwY7MRuaOHjHel5OY/dh/0ZUAD
cEB5KLVQvC6hZ7Z5YngUpGCn3di0uj4ntP7ffOe6OmVsX7KakJ0NOlWmsiLVW5Az
0v8c0LrqFYzrPuFcbCZVccgvRwSDmgOnicetFzjRzOHoRchkLPX43aDe+cB7Y2Az
u5XltS2a9riolJdH3FV3uy3wU0W9mvRxSk96QyY7xdSUqxUW0hsPo6UgvSb3gTzg
efmHB5v+OzplySOEvGftY9doIm2bDj6btcPYz2wXmffw70WqPWNetoayh41WHe9p
yKRLzQdC2LrfCxw4cNmQUVBG4AOQS9av/oQ7X4K5egJDrKAo+mbpcanNU8/73Q/N
VOezI7zy83naVx52bRo8W9799NQ4ArzdJ2C3eKw70JfpQK2kNrICMMaBV9pwN89h
qdA3Tx8cPtYL/SDjepIXXB+XOazGG2CXYO74AGrTRGhLFEbRXnLvyGNenAm3gTNx
2D5gbu+mdNaPP7h4zRGyMmmafyM8uaV84Gu8s11rTHMdtVeB+5RjsEg8Zc9bcrAe
npZc312/LcRZhRw9fOAMFuIjN8f/roxgnrNQrQBS+2nA/CX/RCvALH8Peyd1vOJO
fpJeaBMONqrt/zHApAA3jaIoi4zxNvodaCh0LEba0bBOWYN62jctH/PwPm9uaBpy
YcKb7DoTvI0AQNwpFpwh02GdunyBYHmj4HmKfDqzCQWAmDrpD6mk5UBAdGtBMF9Z
5PitFHVVxYKulbw3hn7DSF+stoecQL7ondAwITNrD8Z8a03PA25v+xdnPXnPqkM2
a402nCBZuGkeR0xk/OvldJzE3aCFkdqviMuXFg/gWyj7OohP53vBFV7OxICeI7i1
RE7IbcBcY5qv8Y5IxIse3oPSHIvAprJwtRztZi/7Z8yua4T81MYDo1kqEV+dHJFh
hJzTczIEGlp/vALkoHRraoUB5WjVCE6FxX647WTpTW12R77bl9HmkwdKZpIqMMSR
/D9tn2cnAWLj5BiDpKbbfTU/eopA1L5HAI6TZ6fY8Pk/4ct+9oXwp3SHBCcCMJtz
7qF5MzAGx55nncsX/Gi80FTs3T3mxGXmH+LhFIXNXl9G73pIPUn6po+/0Zwk/0bj
AaxahlSSKkRddwlA24GeAhW1qVHR3pAJc3cvB+hVfQv4ocmZBlkEJuw/jwJ4I647
oequUTUnBqvoSu33IsRWluPUX47iOHtZOK0vkrckE3dmzRdfravRL8BNLDuYE2xa
bofrsWeBreWvlKgCIzyvp223UR8srHJVB73IgoKUPnUjRbqnWjqtU2hlQJiSpaHj
nPen0LeMik/fxFOk8lUX6kbof3woeuKjVZTO1FH62GsnW5WrI3Jfs6ZAzxWMhaN3
BRZX9y+oA3h4epF168YCQqrLOdjHKFREmyAG68nb3TM6nPeMh9whunKn1Swqq6XO
mmGf5m1DWwcBQu4BER8h5z/cSi2l9fsabpOY+xU7qKejO94qHLTksPSL6FXR5evn
ZGy1Yro+8sHtSKFRam/RzoGmmhCeMCNvnimLs3NLNfpr6Z72KgNNGosZSvZO0uTz
OAdW936fwYjLTKOwsPJOOVtkU1I3N0NPr9V9xCwX8s3lYEb2cYSIJKvxdPSPCpOq
rZ4vqDgV1TUIdaelrtyaA0VKGAorOEtNJ9vRzEuOrLVyXSayhtBggbyBpopiSDeQ
tQSTJ8oIETSLzyrOxEKR5xX8DqLnHaS3i1eu7JUeS96yeoUYtuvZiGBsgZqXL9du
EKfzQNv1E4Cq4UnPsRyEB4mfjs0013qVAXKl7ZqaNBt39UqUEolkbyhqFvk0tEsU
+HWqnU7eYWZo8YyyYAp0KDo8TGd7DI7WhHejGDc+isMBQfg6LXxOG3BluVOIIiCS
zKhzHNCk/VG9KOC94zguLRb78ysd+lX4e7Ss1WFyZwxVpk55olittQCMQhZT6ex7
h/uHhC3zXtcBC60fIg2oYarJ/5tEEHhR0osmXS/KKFJ+PlVMphxW0Ap7iX5oYR8V
tXF2bX4icS+yvXldjE1dKcUJeKDTlgJJzSPe6ddu0xYg9Xpwpj7gHbMcOkjJN96O
57kQlf6mc1LAXiS8RfyNEK05XgJjFxTu8odnrOfpLD7ZgDR5+1UAv6GRTIqXl1re
VNFWCNSmDcpoVDgPCI8hMBReMCHy8GbKTPvWBie2FCEDE9EwXDVlBjGxkutlte//
hdUy8kFiEXZYlV6ipDi9ndJ4NlMUrrl0Je7tUcmcHD2augGPY8sn0/4Nb29pedHB
uD0wivlSNMwwKgUQuZj+j76jhEsKbh6vaQIJ02OSZcXVXL0jPFVoiUmJJ1zTxHQX
cUXNfqFjK1C2Y8MGvP09c4UIOoPijUAf5OwaxTx9+hwuh9/CwBpkfgvBgpguZ5pw
Ci/ylQyTPR8oZyUMPVT24S2Zo8yyoF1NlU+Veci64JyEee4j6ROTbVl74fENKeTR
4ULGl8z3zO/FvkfolxjdZS8qwZO0B7kX/AcW2t/SlnRetFOvnsnC2BaGoFa0dgTy
GubHdpteto10G88erBLxvAoE8AJyW70Uj2H4Pl7/8E/1NmkmIPf2ijhs1eOQWWIk
l7abNzMe47h8dq6mJOTMIl4zl6qBKcRIiFeFMJ/2sLbOZmGcAIyQCL9rIORpOmFm
O7hFpygvSP5rzfONKzg3kqrlno18Md4XyhJqSULmigGIZStAAmJ2bnuX3lfYkSzv
sDJayfRyasazRfkbfS/iPfyY9g5i2lyL9WEgoNk94e9/PTOvaUzR8nZbmTMMDL0L
oTvLZaJOnzLAj9jq/35aEPDHiYFhc0saPPKelRfjLjQ+pczVEL4lxUrftfFdNF1b
5XpOu/h4GYZNnnOhg9DIEgIkyuq9TUzPcOSQdpFnq/Ma5kLlPwVvj4XmZd9ODAOT
hhelxIuloonJ989ZQ7jOrvYyALgeBv7ITHKQxpsyvKmkaVVjilcYNzKLl5RicfBr
EykVDLNYnstLwx4Q6srt6hozLgTpKAUJJlMO83qeSoKZjm/kWOOljhPWwaK2ip3l
cEImtiuUei+velJ3BwRI+P96+P2JVR+wX+AeGX5DU5XWSCVRnCAq0XNeXbIj5xyN
4qSB3WwyhL7UJPeip2hf5bfg2mytLW0NedbMAWFrKVNbHqdXdpwOOXFSLhXzaTXW
LqrlRp1BlMcFP7PLQTg8I+z7K7MPQ8L2IhqrfQUIGA+ZhPwjeDqqzvlJx7oMjIIe
KzivgLmSme82sQQONCNef0tOsjR+nJ/C6kNaJ9G0IOFTU0qkkDXroETqCsgh10e/
uHNz1GbT3S9voHd9ptOezFfHZ+wkzW5JSE2v2EGSsn2RKmOjcvf8WyRSvvKlrAWJ
fl+e15jIGa9PLGJLIdMqVlgajpE3T4JyF+M277dQQDNz/g1fz2TJFtM6EFIji+EF
TXxST/ppPK7wTdtj6Awy5srd9EeJ4ZL9+RzekyYB5XbWTSXTx9c7KbMu4v2Lvfdx
LYiFYv/npT7U+xP1/E+z3PEUgaQbcE8h3/sDGB4LyNpobcTEyavqnxYt8hD7XvY+
36rOJVCTrRaxVESIaabTtqUYqPELt/JHFRO94P4EULIcvCxPmujJ8FA6GwixDRNg
JLZjRIRhquPhqLhAxYhZq26MWj1VtwruEHPQQPk/WPSyDXM5zLeF7HjbEUSy3LME
K0v1HW9DePYJAURVv4CIRm8JhZQPL0os5Cf3/Q+LJDp2E5VmbHVBkXjywOU0i1HZ
L+fE+XIVBKGaW3G+nUg+OVTW2AKW7hKfU/fo1kFMMl2pMXSExjmY3VOmQFuY8y49
Tukvmx9k+Y6rbmyXZUbD9tOCe/M3fQ6tpU15qTy2mLZQwiH/0EVkRzl7bF7Bs6MR
cSee9/QawR/NJyzupkzkrqs4l257tdFR24v8VMOdDb0Kmknmy8mQJs+EbLpkSsY9
6RQP9ao9mcMngb07ettdKJ4k5oE4N38WvAZfxLL0BByomQhIAL5KwvruJ2tx/prh
Ba/4hW4Qm+DunLpyUy/231L9Rih6Rtu6lt8EcIsDWRHjMWhtnJNJWujBcihouR3Z
of6qsYtJN5/n0Ul3khAq7tScHO6TFSLFvnwGK0anq0OYqzMQp8pcZijAv7j7RyoP
Yc6raZx8vDe2ZgWrIDhJl6cZmxYlf/wQWD1VvfmNLN2Ry6c365z4tsuETpELf1ei
LDXFhC209YHA5rtibk3Kzf71fn8fq7CB6J+mOGrqJ4ocSqzQYgwMZAK6DG5k7yA6
lIuEGGPscaB9ky1qHqc6F8qs0TUPZKQMEKWEafsRea3FlnvsCkfpx7CiK3C6+Hqg
V57+ApJElPdJcW61icZmrtRkweq0KYZAwjE829aZBn3yM2/J7oNiBADkUPgCCO2Y
FZg9Gu37AleGowleqJ6+Iq5XJHdbODgcO0pkMXXLHpKmS3pQrIldkAFx19Bp5cFz
0CUKmzt50uat6GBX4e4XOT08Y9mCT1PcQoVbHwFd9EPiqftnRLr8NvC5rphPihyq
4OiJ6ij1ylNESRxq1x8Cs0uRii3A4fOu/of6x3RM2rPg8phcr2GgXUvClgS3INnh
u6FTlYoZJZ++TK4AIJMyKHVM/30PDYgtvWHV9TFl2xi10L/a2nGdKJ3rujxuQLyE
mGt+IjNAoZ5tWRV6O/6xDMr51pspVr8mtei8V39iHkwp06eKQbAaKTvIHVAThpYE
gRLjKtUb3W9HqXX3Ro2S0yABnq94EaziAZBgMet1dSoABT2JtkYqxQTzvfUrSpmu
7UiwiwmcWp9eVSz5DYW/fz+iz1KRAds3htFTDmXRyUdXIdTkbIA6IxPk47rdEAf6
upCpFUQ1bXvr5u8meegisEhHQu98kGvBVRGs8FOeT4athSlhqUoYcTe36KXfgtK+
XizvbND6SUOwtGND/xgi5L8GKuRnzjssswlrv0RkPlIHQ8OD5PruWoS972rEgaDC
bBrqQnnQ30puJouAs+BpwcHvPoEMDTGQnBJsy6wB9f1wM1Q4CJWh3bY1X2AlBNL2
ZeJ8Gre5vLphLoMbYeqNSrgre14K8goQzqRQ9gk9C6DxMElNXlO+OiONDi9Hz+vT
U1YTVWVkAVlyDGW2tVwyBZIbVRJQjCu5RslbcoWsjRcZmCI4NYif6ElZ5Zy1LQY6
I9N5iVxDJFD9Qv24Ll1/nT8AZ8h1GJ3dVr6vyBKlQUqoUz02RYbzWuxacIyZPGDI
ichpl5AXH5gJiAMwdanL3N5Q032c68vDpgu1UoHXaJP6zhtnhXA2HNNOsiivnNIB
BdEW6iuuC+x0o5vtsh/wQOKm1Jl8iHH9JqHPXUlsLAa1rjtJgA6hTip9Tr0iwovH
gbvALjULkCvLypkMw/J95OMLaA7rlDaM6+M6EyT89r7K4yWeZqG10bI5Q29pNabp
Z5M6R/M2OBNvMUPvZlJRav4MuYGUfYY5Wdg4DwkK34Dh8+5gOMntoHv4SilmpHag
5AP/cU1kI4q85+Oxs1Q+BTHiFJ1eT3TtWzjLMIbqT2xf+RrVqxw5HWg0sMjYE1UY
sHBrfZjh2N2sGwT/MKPR3Gqajzha3+QTb6V+0Rw8eDRfzjCxt2M/NWp1IWmG6WUI
5LnpIDTkSXGVCVyq9kTbMH7SzrbXP+hg/PTjDJFljlCewTiCGuvUog/NIkThmM7M
UklbE4GcGlEz4HDaNQyM3SmLrIkUicY30Rr0BtrKj8xdILbFMOkIs2Ig7iZFiLEj
7fwzjOs7rpnxt+FS5lQma4p7LEovJMhHQOjvn3stmxLSCxXFZhdAnlQudHIIPV5z
aal2DGoXMTMJpfZfwZM5LUg4cK5HvVP4lYRPo4RT4Y9RMVsgr0GyyZlILZUfD9j7
T70/SnaN0w2veKStuT9yUQf8d+CmURCtYGIDTH9UuiO1la9ON1Hg69PrcxAa2Sik
2ndBX8tcO1givt7EDeOtLVaIYTEFOaBUBa3l2tmlf+U4kKlUoW/BlOgDe0KiqGO1
ZG+7fx30TDcOHeC+lR9UkXlEA37gF4BSqZFoGG39xs1qhAn24QGrzrIE6O1X7iVF
7ZgYs5Bj3/DZDgA7Xfioim/d+x2X/oD3d3Gcb7SSySINmfoq0TWGlMdw9RZ4Ns/B
9lwvcjLnyamIDh8KG4r2oEJRMhSsxT0/wr7RqxJma12CE5mAzHKOdZ2OwCe/iiJN
5xp90LS8hL9lpMo6qql0qE3w0ggCkyhIPhLWd9osQuo25hUiL60hkpChi8gRaU2G
3Md25NXZExJK+F+mZYalV8/nBXuiJgr6zj09yuGy04Em2H3wiBz1fJGTaL+iNe8i
xeq6NTfZS4pjMgyBZi1OVG8ADac8weNrV6d7IecFP5T10Dpdh8RPCeiiC/8AJioC
VRAwV19VSopQwYbCuRe9tZEH0SIfqvhpx08Ls+zGctFCOp6RVu/umG8p0iZRM4kR
U4+yqj61ButmkSnIbbzhYYqtZ+nQHtMcZPcZaChj68H5Fbg5Saz4Ms8AMLgOIF/O
fp0w82xupTWzi++rLUNxWqvX59xd1Io/VYfaW7mCIicIv7Y97dPOdgFKZZ8ZMf64
DSyR9grPy6CZ0lqpzrgJFpCBnKzauF3xikALjp679aZnkmItkTeXIwq8ijMz/jXo
FuitQgtMXmGtuZrHOZ3QCCtncNLYLfZVRhI7c/fdqOY0GlKuFT3ZZJ9XHU4EFNg9
Z1ksfr34FC8SqVDHbo8nTGOUu2bYRlJ7bPJmOce+pofNt6BF72tDcwv/eJwVr1f/
BSbzM15sjPQxCNAPejhYGKuLsg1y4P7pAvzhTT2kySxZSDaOcYGunJxKa0UpqCmN
/iDpbJaFQITpcclTAqJW3lKVAZOQS7h1Q7UBpSx0JRjzdZ1sJXIvNKMk163tmzNi
VO1OTe/imUJQx4IoYbtefoL1hpJRkLoGTIDRBsS8AuKixtrRG2zpvwQ+gh2hIskD
20JE026wKNrTNoR2jUXqTGzN8Z+N15YDgJYaac7peh8MTTfm2OPt/nuJYGoNCVQm
kGXhFutEsWRQQwRdTcLRe0WVhH6/QP4KwGEXO1HFRfQE2XD45LqCVgHgXI9YS3tu
zKsw1DzrUnPuz5+vJj2ryJ3/rlc0QRhRM44lOPFQz+gGGq+VmK2xGLQ3WAonPfzu
BePT94brG/f/bOpdL5Fm8o/sbF2HLkyVktuyn02AXyiBQFWOKrMSR6k5KW5z4SG4
9xxZTbjTci+cLoxP0g0Szt46u7bDUWkLxtindjnKLTlYH+VVeFEB++sNufGUWcfc
MB3ntsfssjCRzmBgFwvvuQAosPTu1FCu1q2VQ1STBG6LxTunPjSPxIMhrhX0T/ob
jt0RGB/Wh/beaZytlRnSYDxoM+kFjBz1mD3E86O9qVY6lM6C0v8NeM907ZiDThQf
STIuVBKXXPjzG6rakZeR2N1NSwkoO4o9KfT4wimtnaVFvGBlNIvFpobAjb1SIt/H
wkpii0KsB8DOgIrfA+gUrbHKkYYOWA/fz5U7ow0fNRnj7Z3SCqPVLGmT2OL15RNy
CA3UNpDMEJiCIWLgXYBYmciazfgXldPcIBk1loRf3hdwoz0auWqoEilvLjwc+76l
fkriiDJsc/YfQf9Ti3f7LSzOd2+gPcCNwsk6Sg3ThFlQ0kDg5tcLBh5FgqH5z+8s
AkQqKVsdLE2mcY52S657a1jjfbJHwvvliV09d4U9zHaZHqUpbqWCwCSbBZ6saUPI
kG1WHJHGv1rQkfMbKwwJufq3G1oEhe+OUmWZlL2DELz7cwhgU7x+uQLcatQSXYyS
ftR5+6I8bYt+k6BDYIMBcVyRJ9u8s6TYkoHOc2zzpZ9l2fcCO0wRhVoCSpenlvDi
+MBB+tiwMWDKucPsiiNiuozaUQzMDsHXUENsmRu1lp2UpSnVbg6HVTj2nhzVL+RN
i8DRigsl82VLV74reNkZfD9xpDy1q8q6ESL1Flh44E7uNkpklOklkCjdcKByS0No
wMNJ9GWY05VJhdBHpRCrfkArCqTogXMbBSRBf5ft/UemD091F/XifiJoX7Us5W9e
6s9kbtqDDnpKaea9qp461DdbAemPACN6gbScfeO24v3RBvrXeWSp1LFoE18Y5AYu
+V891bChs9GTwKcflBYQwzuokM9GWgp7pVcCEH0Hxl+62xpEor7pb33rVNs3xKou
YQTBA92oHhSb/bng0naEi9ztDsIN9T0xc8zEZnAeDb09YMWyQcl8H/TKK5ttadng
SzeDSalXnoYDjWkFHf6xzFSRrIUe2pTkpyyaouYzca3OnYWeNNt5lhiTGkjFJz6P
7epwEEXO+9nQnN9tCNv2hYxdKqNS7+2vjTLoXn4tZtkW7Pnq/9D8MX3L9afmTsS4
AOZ3d1ZpaWsjvd8CxBOAOSc7ZlDMIzt5/3wZbMgaJP5FTX2/1Ux8U+/sY2ZzrEH9
GPGpYWh01IsMQKWu0oWIDluH/9yScPjJr/xIC30zkrhYA+/urHetNaLPFhBzhIwo
yHEb9WQ7Huwywrt6OTclibsAjRtjRsbz9V6oGin7FYQ+Y6P7oJoab10zkaymx57F
Tt0Wz/GqGvV7k3gAldXvpsRfqJ3Wp0jq869ghP8aLb4fYgMgkSvL2BcpEep/3m4c
DVt5zzXmoBT398IypJJoaTvmwodD/P3SMWHOKUB9QE2RziICsNVwzl8eWhrQtoV1
kUtLkM81vNApnHfISu77qPwdr2vkJBMUag5OsZo9Y6M2TsszRqX/uLfEk6maRD9y
+mAkRyhbp4o1iz4BMYpjwiBi4QfshUOwTnfzaaNEAQ8I2Hm/kbPpob0xpsLvCnlB
/zEazjkdWCRxh/yoN9sJf0Jknt1ZcMjpcYBS+IJfdEOtwWTNapvwM3enuz6yYuWd
zldZqTlNfc0rNmn3GZ7QDx9cv1hCaFZ0bRVOCOIWV3VKDy334Psd3g0LK434Uiw/
WO1Fi7iQwujXi/JC9RW9A4PTHOtwGMrAah2dLRvD0I0KRkD4c4me1DnTqD96FPMS
5JVmzfxOtXOcDLzjkBzAAone/pw/OLI1r/k2b4V+a8YABoP7WByq04WLEkoI3ymz
XneU09JZqWwA+Dq1MY8uf1R41YmFI9D+9PJLZVg45vBAnmuGlrRY7sHVw0MA4nZ8
zjy4axwE0JYTzTlpLJptktPpfRyKrGLHLdrMbd+rI6HTjKz4pU1zLOUGK1COQje3
JqbBj6xVdx5nhxjPhA0VwlcWz5jYd3kmMWtJMmXktTnS1h+HmkaM6kn4vZcYvSEW
d9yfc2x0r9OjOcwdkXTkT/50/ELS34MnohJseowXXNEYw2CEl8aXtbvqe1OMBAu9
HdWCI3zNUGvarPk/kAOtEqJdpb5q7ru8U9bwYqf5jsn4W9oYnJsCpwi37Us+i69w
++fWrr9ofbGG3gehheFdePkSrByuefDiU5gNWMMkpCy5gdLC9PGzMTNdAx0xdYN+
3doVlkokF/5k/KcqWcuXXvQV2lWHHpjpqC3G+VA5BCjXaIVJ/mPcFJ30p1ZLgcEX
4BjNFpYgyHoUu/FY7vccn5uDJ3t2nwY2PQn0uysZohcy+91HpWfxXNvTmEj5iArz
0gual3K0Om0vWjp5d7UYDqmYIHQKqostrzG/H5FDaeCsxeaCeOQOj97NCx2j7K+z
VQgO0jleULIJwu3Lj2Zy6lWySsyC5GTM92sDnl3ct4tQB9RggMOTP70q+N9NDUGL
fnjkmJJv6JugkK2BwKsPVT2XW4XLVb1ldaHek/ql9yEECbpr8jiwv7Y3bMcMPOgN
fiasvDmV4z2WsJAoylXn5WkU3lMbjpODGemIPAPiFS+x4e2DDkMVm1fPH9nXHfWi
JYxdLQWCVgTU8cLsGQa2v8TviUR0o920QVlRR2nFM8BJvrcMk3siSaaxWt3h5ita
75JEY3GC9nVQpFbfVDWId+MggxLbefdZiEsgWoEgWXzimcIVBQ+R4Ooyh9SoF8v0
ftK4NSFfD+59KvCzVPZKAcN8DXus8zhFUslPguAamK7aHldcAYs6+Gh+NcGa6ENT
yhmD5kPfUilN3DM+/HD2MkkBx7bP3FRV0zkZrztIaOfrfvs20tum/sJTCkKipC5k
GFquS7d3nxUZxCsVab6jAcFUJSRauxb1umPtjOqM1K+i+tI8NbaH+2uhV620z2T9
338tXc1+C8FZogWZ2fGN5F36+b2mu6bVcbxaaHQm3cpZQfhsiKTj80PhXy5+uJj8
aiZ1cohY89KMYuURUf5VfXOPs7fdS7+83KHbkPgmQYssoNJ+qEG/0bjJzwsSc/Vi
zSFmWWECMSHJy0jMFO6Qsu6CXNCHyNCRvukN2AeI+1f/0zm9gaDByX5HC9AIhAVd
pStvhTLZSbfrGTb58c6NFOD14EpcWsmbSh4i2Q/JaOGABkxFQlnoQY3SMNmWwv1P
nFu2J19ebkgzXYm8uqADb9ya1yrsI2z6b9bW3tMukaSX+Wlw1dO6jHNXIgQO7cnu
gG8Ptsig6gg+dlA6ak6XqR4q82J8foJB27IxjKTouf5vhLJME5A3ieLE787kzNOO
zXesFqmgXNyPWKfQobLaPCX1xKlKCmori347yQ0zesyy+bFvgeQQunKQ3A4Uk5PE
xLLO841iuXD5D0hkncAX7vAVKlxmrciJ0WrIvfvnfqAFTYLKJl1yB6MhYyjpUSj9
mUaNAs7bRfVp1Xe9kQ2Y5bqw57vWhQzKw3B2ptLNV6WGQ1JiWCisJtMUiiVWShFL
+9XelSx8iuejmtoPD02oflJPwlRjwZ8zRCT1+Bs3p4JyIXbOjBnU4vsbTEV13c2t
nZkefltV68KEV5nuShp+cdeWxEiS/KPAJLQsc4gPAoG/hnULeqhWHe660oS8muRg
GtJJnH3IK+6X75Lm3KmAzfE6gxrWC8vtqXsUhrrMoWgyco3iMkwWA6V/cBGyKmJ0
rYwEIeDB2a0Apj0Uf4gKr64sFSWz9IVmKarMeMPiYLGKDLIdgqvjOUMV4jsTg+Yv
CZOk4amHEgCoM9kHmrGdNcXaetbcsH/sB2psOz4XmWSHfC84BC0tVrSvtqld8s9t
mCX35t/6sNkfGXMgrr0gMZuiiaJ9kRPcU4q8+N1Nk5yV6OYAKAJD+UjwF8LHM3gU
PTORWWBR40cxKzINacHsU8MxfCv6+QlucQirztEV3B38dRqzm03iam6oR1a8IgT0
ds0K5ylEYC1sb7iPlnjZ/S5Po7s66rcrRSnfbbaKm4WhfkHyyJRlHVqV8bAXfqh8
30I553E7A/afs55djF+s1KBSwV8xUdxqJ86CkpbVBvxsFAfYu/Vmg99HZjk/1nIX
QxA4o7tzCyDwJrAeAKdKp4cVzo6uV4cJoTqtSeqTQQzu0etuyTGxW+qkNTLu7ttp
bB8at5z2h9uDZR0Emg4z9RcQWe4LGZnY0WhCVF4pihbgLcHZcPwKjbjb45jd9Y2o
Xpi6Hv9BgI03cK8AsoBb1H4QKZgcWb1+SM49bTVEW0YRJNG2rWmA+Dokr0JK2EHu
Cn3HtQvQR7QIfPTrVQDhNWiGvYIIoVWZKLaj00lBg7vl3KsrTMA1jFhZXCr18LRB
+TuLarPqEx6iJu2iJu5QVbnWYiZVzMNGEkPRbwpls5A0TyMGC+sPRbcVcMMUuBBL
KWzQ9J3/OlQPsnlJLhkLI2U+3Qi83FSld8mdQTHBwmKuVOfJRYgmUJtyK04038GA
K4yWrCsqin3d7ZYSdv4+dkVQDsJOb6ncUCwxkfUgo2dfdUyKed0w7QYt60pjBrEX
hxceUXTT3cc/2pJn2APiC2oqlRBKfHbkDMk7pVU0uQKlwhOXYdqiHmJXtLxZd8tS
tGdROjg1TLsWHoADK28reEsQwIzeAh1AUqdzsmRGZYAaztDgseQUh3j8KvvJRXWo
S23QsOx2CzHvu3zvWJkiDHKKLFmTc5GnW7t/1lYjjWcel55ICJ3lSPeiuI0pTYfO
7XA/4son1HZ7S6cH8lzxcVrx2u7G74PTKDOXLOrZDV/AAvPRuIjZ5bBA6sXT22Wu
a9Uf0AWhMmC6Ak6ks28cf/RlRF5azDx0dIOhsYTa8tlF6QdNO6lTLc4RMGYN19JC
VBaA7WZ5koTUvzB0F2mDz+PALlWc0mzspVP49tTKOe67VZqBkKB/B/PLvQjmyneO
Dr+ZnEIHO2Ia7QfbPpm6q3gk6cwIeX2KzG0eeGyHq13xB9foL6dwCGamBduVIGIi
zBezKV2/p1uMeKPcedILTJejhia12Ox5EceDaV4uygrhl5Zw2DxEI4k1+gZDVdhF
idlgGANNCamD59IuWdabGV29YPf3yXq/9JeKT3IVn9TTCZFG3V5RY9f2IHBPfhVT
UV+D2O9suBv2UGoCNo1tF0HHUWbzPeHwPQBoDuXYL1kw7ug5tGgE61knqx8AMf4j
P8sD/0Xy+01yjcqx9Kfdq7BNrKW8XYlmmwyuN3lZyV8RG6YG5a/Z/t3SVbL7ICbJ
9k/67Dn8pXf75Lh652GZZ4IzkUYnsobL0UOaBdq/+zDACiZF6hwQDo6ZJk8iDZAA
9cGGc1MtZUIPnUj5jUdfPyu9G/Zv8ZdwPXmsUrtm9x0kTFSN5V8Cvq4qQyJ7EATV
Xt/Ukucz5+32PsApLfHrbEVBmZIRFHuSoe+i6NOWRcjxuvUgmyVaE3+d56lPijiX
ZH+nEBVcmMZ150riK3DopkIhJDDhmPaL9p5JN15Y1scrlypxX+QC1xqi1BKEjs6c
otR+HQGbDqX98xmgG71NCWskveB+n+xG3dZiuZFL56aD4O01jIOCk01lmsuVhtnj
ehO/yktnBnxZcnyVLnnWJyDRhkQFYm3hnCT+BHhmI3COj5o8Dgpk/xIo/g/xlI7Y
CTXbmqxlUVP6SbYgloPQR8M1eRO5hhGOU3NIi94MfBYd1B2L6JKtlR4RtTMaXwhw
1DBXVuXFS1wgW6QgBUn9gY3UCcuBzfMW7DwWY1PXv0Ixr7L9PJTz8KW5w09j1eNV
lyYVdNn6h3AY33eJQt55+BzANIXoSTbARj85RDwly92v/iYwobYrJF5qA4SnZUj4
0z0yGTNPdXXCNRbrM1eEBy6Ti5UEiB1M/pfbeazr4f24+Fwv8uUaqdl0zEm+2IWE
25lQkLc0saEDiYPdjZjSXnV9N2RqrPv/0H1h6AD5vDQ3TzYx9adPf/XWlW5tDbvD
75U8AN++iWdMM/C5mRnY36FeYeAOUFQmZeWqUGgW8boQvfgsVhByEejdOttB7k9r
ZSkFtK8EXTZf6Ulfwf2nPQLgLNrYNQGNs5+FrCcpo6TYNWx+pa4Eg83uS6WeHtfU
Tv1ZMDLHF/C4afoUoH2WyGX5MdxYcH9mnB0C8EZW34JBtkiqt1/c5BdUH/TfkFMQ
147lhm+ANKIfbQLmJA5K/U6DFkHEkfb1NZf6pSpJy93l/TR0hDj2Ch94VILQPJ93
X9OudEzspZ7TDTzUKXvar2M+lCSWKrMv1WiWBn4tnKsCFPc4GTSfy6f6zq7M41gh
NqlGC36MVMusBSYMDwKgMSFJfWk1roo5vgCkuekDJj15a5sc7V83UflLqmS1Y+ob
XrLqLFTbl08/b6jl/wJKZDuN60GOfpw6Yb7BX4+zCqFUAgXdMe72JKSeA9nJbx3d
2KSAr3luQeNbgKyIBRWnYWXahEDmlZRlpqnziIIJ8ZL+1WkVz5Y67AjCBW5CTU2q
E32epMPiAVZ9bGjMEfs3PyH1hOXDARQ9ZBhuObLQ9Sfq4Mp0Os6ecNCv8amIo3YL
q6U7orMdvVtM5IdqXKT5xBqJqCJQDl6Z8eRIqPtDlFSkaGLFQOXeb+TstNyfmlM3
MngbARXt+Sl4fAaJFFxC8/shnAVJJMDFDR12xVweGXVu+O9EYJ459TsZeoMj0Vjm
B/aRPGtJUpLK32lB70jJxyR34mgfzQHO87MJsdHV53KEe3rCx7O4sZexplt1daF5
Jt9Ww/DBhNyeLobHbxXIZbbvA/tTbtowWb+4NTRnURvbgL27H8qjHlt48gEbdDDH
VccYg2QkCA72SzmuzYZ626AoEggFitdBlphQKAJb0e3jPlEhC9gV1qXjp7eD6Q+l
zUc/7uqgKlWiZDGPww1Bar1HaAoa04Eu3xOh5Y5EuMK764x3ksJubZyVsMg1tJUo
n29R8mj8rV8njbgL3Dzu2XnGRxrGMAzqiYcoa0HH4bs1EpqAmQNrbWzTfI21c5jE
5+gECCNL3YD7SPcb+onVrZ5f3qcpRRkL1CQKhXR8B3gmgxJg4OHs8+2X5lYbdDi7
OmzBGWq0uGgUMMraZ5ISklWNgXJz8CmKVyR2X25TOczpoA67gkzkiAwkoy8fhEVj
pF4J9m4eTDa9nZdnOUuCgDfr2hgGqV9sTEvUBw6fP3wEkRZoAhermZQleud0xh4c
A1llQpbVDVxcPPVLypFXXWK2yvRz72BFoGuseopZF55TehwwxqPO1YncJnbcZ2xn
vLSB7ePq2Vr+V1kURPjrg/8UVJQZgXqR/3NEZK2ZnzOu898bv+bS2XzRwTqc7vT3
cue1McMdtsfSbAYuFNStrVDgMN9+puF5SG41gDuC5g7/ge4VXWJco4AjbGEkQVxK
PB1iYxAL9gJMCVXxk5sbrdKq/KCb1Iixefh+pvSi7EkwKQhI7FDtWTTRKXXZsKzP
ZBj04/rAaFTG9ZrmbO/pWAJMH9K0G1UAcyGhtKTLHwpGF3+rm+8aRgsKGZ9qNSRK
rUwEddu8PpPf4kphnmLGmL14r1NwZe0UajViipS+l0/ppOkIdB9FxYyWdM7qUN0M
2H74/llBQt53gqsYShy52CGF0bt62sf2Nfh7+8eUCIrWfQVwqDZk3RKWU+nSvjkf
9LiFyWygv5nXGaR75CNydXWxTuiAX+y8SseE4AY6spgGq0lijfbydo/WBJninmXy
AJo5lOiuyTtIOJZqkXN9x2Z15R3a2FQNiVkQx30iaOWFW7wxS1i5A3qzbqqXxmkV
s097yjoEnJPx8fjWgPSnDKj7aTEB9PzhgbNiex6EJuoSFhHQuDNJ5gAYqSPbBQwT
NklIhJxNUV4MSDRM0IhnN0V5eo4jXHQQGqx+Z9INU9qH5ajr/gTWgYCKxDThngpB
UM8Xff4DOhGDPqSzzA6G3yuK60vxLL7mpLkosp+qGwWKciHrY7a+HkFL2RlCSgf4
RNhHSPvisbjnUGRrYO8AVPZFbW0pXDtw385DO3ogTTZrhk+c7kCVakxEdFjTXMqp
AKXHylaQdoKCHbWTWubhn4wloms3Swk0QPVW7WXOKRJqW8oiZ8u4rYxIRJNeSxwu
swzvVCKtduKKI9F69ppw9yCuv9Emnwvtu2xvy383NZBNEShMwLI6LvrEQw44fvFw
xE7YZb7hUQF6dj5np5bkpGuPqpDS9tbl6TkVBsVVXOinrbNdSwjf4o6v+xvjFMre
t0KZwSevW7JGai/ahhyAWE/6fAGHlzXUv+otxGLfsElpUQT8Rchk+xUycWQIPJn6
uK8e1ttoHaCHDbTyLR5cp/jbAsaZmX8gvNsMc5mlQCJ3ni24z6A+c+/kDBZ3p669
mfCiR4iTyfH0ad9MkaCdjiT/e1w2mH1iwtm/MGDDYHkiOHBKNPTNXVuobDQOW1V4
DlvAar9+0giY+aol9/RBtuYmxSYsNoqauAsz6cGrunLWLPplCfQMoM+QQOidARRV
OU6CZuKPDo+nxkFJnl/ywNq96dleomeuHFxPmocOs25TuJ+AQyiSztFqrHNV9CPy
mR+YEwdVM85U4DmhLy6xy9yQM7dLivlgDfbbB9w+a7ioaJaaEp8aTtPQ0nTQRrLp
a8E+8SkejVz8g22GSwubFlePNPvS+Z1Y+fwvMuqqiynRUFZEFWy4DhltvpEoDyQc
ypo529y/EsKIqicLzAJiW0jI4BGXpxwL80XKAbJiMP2Tblsp0H4gg+4Gk6tyjHK2
dyajuHE6hfYUeiv52Ab2pEEVpPn3XWZsb3myrIEHyMh+nsdWL8LeKUfKxaaZI5xx
VIhvDy1LofDZ03kAE34lRFypnmeo+g4eHD4czO6mhqZ7zgPEYJ5Rx3k1JeL/pdRS
n58b33DLg22jxI4WAD1gZYydVWwCgWDIWcsAzorUDN6VoURk6DK7/tBjM4zgLOHt
hov0yl4b+g0/uKX6qeGfLuHfCpCJ+/08Mf/Ln06yedZqf7iA9gytqeTbq1UuUotP
lGCxancfZ80XoZXxZjBcnQRph217MTJzhvQ/WttfJHkeCLAMWzpjr2ywdCRc7cKi
ak9HpaiZ9WmLx2pNIOXWaWezQIoLOLWM7d/pzZbDMrqwD+Zxq5a8KiBQDtOukeIG
HrpAofG4dG5tA/9ElY4DnC7Nd/URz+jWk1V3BgaYw4LwVf6DLyFkuMGByJrR4xcb
bEkQhXAj6YDJan6Ywm7sB4rdY6aDMO8zSnLegm6kXsieLAsz6drs0aNcWrz7XTc+
wBpSokyk6mTAiUYP8eu6a3k9ItiANXQazEFYmemX0nM3JhdsXxWthLQVyAK8Ed7r
Q/JCFbNW7t3YSky2/Exx/2tQLD4RtErsICbpDVCilnqYpRJ6Zd37xT/M45WKVW+Y
IauQijew02/n/urGX30BVC4V19F3Ee6HInjDUM+ipvc6NvEKB+Dt43QO7pdBWhlm
QVYcIt4MBReaTw+9cEuTTeUzghfXLaolCszRkhUzikAAnosb9rO110QPnhIy5fOT
F7B+XlxT9/dXcCyr6ZXUJU5SF5EMest6RIrr0UStUimIEzKWu7g1YydsbBzus48Q
ETB3OX2i7MXw2uk7tyUqmBwQKT0NhOJ/x6cIDKsCNk51NJuxoyY5ta/CQ5dZd5rk
F9aGc2q+urcxN4N74JTFT7wNKaPRTXCzaueMHm1GJfhZj1I3EIs7W8A/TrVOmwUp
L45UO1ZSEt5B89b04Mr3sxAoxCatcb0wTzoQrKsvEMnvhACJegiGbisRkJbF8MWT
yEQoAFfsN1QGrWlXAbPHCQ7EgSoRS/XNicLsJAQOsCSQMhK+xi4ExPuIbrqY9yry
DYQ8qWICu5VOiu2Ta8mbK2XFGinZJfo1Ta4X7O5WbH9IL/iJc/WornIpneyTVah9
+L1nhTX0XTpqv6j4HZdgKv96nyOpJgCILY4KmL63OBp0Tr4523eVzjL4DP7fQkzC
vZ2YoBw++GrcgHhf9mw5awOK/EajGe6frgGII8eMP4INV4K8nD1zBi7HT7b2uYBg
ll71EMoj41t0p/mNadMcHmUEfYlspO+T41t8J6jRIKCK49FaDv02H02aWRMRuqM7
eH6F3cQvccqiBm1wxsnh8WRELAZgdx5s1r5LBqfeCajxut/4yCucbnbvIGjd6vx3
oIBzBZ9CDh8m3obBuDYUV1Zg76EYK35a/3ukAnvFbW3C5LVAAtqsktvgFWE8sB7G
+7PTJKgnRQKusuGMOTzLB5GCLM8S7kz02LEacoCIqvPFdC8Rg+BgRfatyaN1/b4l
uLMY80Zn+N71BhYh2GwLqQBe55R5RBaNslYqXmPFYJwA5KEzhY0tDu3zUiIYJCvh
BeojDAkR93UUjSSaV2wE5bMnIWbaf2rHutsIgT2EfthUBrbeLqzoSL/XgQtbsvlP
vBGRwWKU3LK6yXcaCaCO93ZV7/2S9bY59zMq3sFNZhRsUTGDgvI6eXtgZOixdeIf
jxIKTHtjz72+8CijM+oP7R838OKoTchVZxKtbiOchOJShONoIOqkwuWwcD0JJLDb
9wk/ALGTB7zQpVLlOY2BNo2W2VQIUnHvbxUbwPM27zR4GBBzWVKIFsyNqv9pOtVQ
z9g3C8fA9B6HW1CV02AB12/6CVegLgM3WaUoiNeH6sfFG9tYruxcuzPMM8lv28+s
1qcgG7wXaTSvIE/t2WVVC7RxtqWOggsROEcHRV5NNQ3G5x4r3ov7fz1yFC4OzmFI
1sJSB77mjely+G8fHah8eLmHp5BvfeNIbmGbF87OcfDAN/eNGO4ocRmBwd41v4vM
g/DM8AJGykSKCm1E9xk2tFdEmfQfoyJl4jfJUqdW7ITuf/P3rkARmGMg6oehTC+7
RwD9PxbOFXmPCh1dqEM8jqp8zOVG4LBz7XWXpfOYhduuhelGjonVr36NU//YLw5y
fL7SNzHxCn56Gzu2lLUae28J3hmNTlQnP8eIvDYKWUi6mQ98kM778ZbVdR0mC9/F
iWRf0mcIZM7Xl5cyytCBZN7y351siKIfPEdpSVqi1+BKAT6T/jsUQQh9Ut3z498W
4Toya13kB5oYQZyAtPXHfOk165nwjA4AGKUG82oL4qiI+FPdD0xV3m7/FgYLcRLE
+FxxW81fo86aDoshPNzoOQ0pmr+0yMsBDuJUQVVOW0B8fCkoKLJ7dUyeDxNVf6vr
fBBruyY4nv7YBL0xTle6vfIhxRkKa/ltZQ7rjgaMKgcA5pjHnJEOiFeEwCTrwVBY
IuDBefkC1APqK2HS2eJpSQmpzeIPbFIWiNv3BfK7PjGx3+lODj6F/mE9edPLUt79
OLLByP86/UL06zorRO5Swa4h3L32UQTbd4Ka+wQfMvNL6JZabozX2lv6Zqc54bd/
u7JS48a+DaxRvtFRuLfHEiFJGHehKZIyuqeWK2J/E/rv/gaulAwJ/o4PR4B9KkrI
k0AECepQTgHzJmNsagEgXl1PRKXrz9XHcpBE0DjVgBKeYNaCCTo5jmdRhzU+pfYn
Oo2wX7FnHTrmEGVyS77SL5Q4TxDE4Q5ZiL/QZt+1aGwKANqbiOd0VHEOPHL8xoXy
sPwlyCbGFKcvhVbT2cstj3iJla6luQegcDZA4GrHlHI54JQ5fIG4rUDN9w2oboXs
JZOU7e3IfURwY8f3klpRqnjww2idj5VhE81XEsKLYXO2vQEUgSo/h9BlE2figs74
pwU7XbHCLy7ADI3GHh7MtjqjIKC+5wDupShCfntjQX93kRIAHIr6N3qHnBKu7dDC
jswRzdxDTZ7/9/5oaFw7YIGM3tVeN3Xx+46AnzaEkI2nNaDGs6ppoP2dR0UIRySX
9fGumazT9+NpoxGzu5jEF6rKP3FoXU5jjOS9GtRyrBJ4MGUSC75o/FKCmBxKWteT
iNhUGVeUnv/jIIaZGRdB/LiSN8RamQg3tI2uxmkA5TcP6rxv295V3lYv4Sifeufl
RjUYn8Pehd3uHQmedcKXdw==
`protect END_PROTECTED
