`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DbjP36E5U2weHVDfN/kZRvpO+knp8ULr7GjI2yy1R59+1he8EngUK0tGB3gnVv7I
xwgo+fWPHOEx1pjVjPciPHsUH7zREvyBNJ/FuJkwzdJJDX5JZcN8ZR7RnwU+GHAs
MzdKLGKte744BaXM29kwdpplLyJaQrqtXcvUNwIyEaDf2YY/Ob7LtHZYeZ+oVSuk
e7c0ZBxSjEsdsLo9r0rlGPFCnh0fIaodTKQMcHTI6fb3i189aHd2corll+yYOB41
Wh1Qzdw59ufxT1qYAHy5bs6aPDgEy1ZoqyEywhOEj1hJ4/h6SFnl/1nxG0X35pts
OrtHIxjhAJW/lIOV0jA3qu3RA8CMGBQAjIpsTvOVDdc=
`protect END_PROTECTED
