`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FxMMW5my3QjZA28UyhSzgSTLp91l6k1dm5RFoxhI3R7xDYUHwt8EZB7Xt8oH0YE9
Ar22/ZRmWF0GxL+6c8U/LqpB7zVDEUIHl1BfLaIu4N8ZOS07BENokDIOK6b+lpR5
oziBfKzWSg1VBbHl5y00RgMe9rmA556fP2MSU3Njn+w6EQfrmTmJbt/Scx/sOAEg
/VWz8NYX7p8XPf+bLed9+2bIvfw9ucOko7V1x8fsVozhNIDbcyyjnCjZNYG7nHQz
Weg78wD2zxHWB/shOd4C64tbb8xuvRk+H6DeBNiXQ7QBzL46s40SV1iEX8IqK+yp
lzTzpXpI/2CcYJ4QgfB656wd/1ocAAMJpSlqUG0+3wh7EPL5NnAOXQvOUbZ6p7wX
7CCj1wNMePqywy/lKRFu62+Rc4e62fry8y27y3dMZjM4Bla5LXXsgs5QJRx88vi6
9Ix7hA59TxYoKD55hDY6iN5/Nj8APh8nOlab464SJBc80o97C9agiJoE/JBuO0ei
Fuh9lHDOzkVclEo8bNWDSrqqYwsffYpIN+VPF22Dc7uwlIbgthG9EcHIZEqSlm6x
`protect END_PROTECTED
