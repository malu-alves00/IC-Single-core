`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DzRFWMALMrPvgYeOAg2PJTepAsfoOpzCnDtOoEMDw2ll04PtX5xeL/XYGg9qKerM
PDbro6p67fzK78asX2TRUA3EagE6ZWSINa5PN+2by3N4ZwBO1Z6+98/6FoeI9NqF
zJ1RDt9z3ciLX43QCswPSi6SPPNQdkJpCcWHIRpLsAj81mM91rIaYJyT9rkXWKB2
Ai6OztpiEoeQO5e/OFgDoMa9FxGRTiuepLUy+MDec7VZM78w8tr/DjnRy14CIc3W
jsTzY0yWcFOSCMMnZliHh1LZZP74upqP74EIyL/gCgLE0AyaiGod2+Y9AeduFFKE
Rp0axMzy+SCeHUy4XfcZufGBNSD4yCMPU1EqMo3YmFyZALolMZtG091KdPswUzTZ
tPXvIFQHisv/DSETSWg7lgCTJzioeg4Ls8HUJUIPZdeyU4k70UZDYJ6mC9lDH3EJ
wOr8JAqjND/Cmn2dAJoXDMNw3IP5MQDyw5DKCLxUyqH6yud+M9LNvsNx4FKf472z
m4lr7EET2p30CI90E45lM0vskSxlyYHtwGzdgLQEv/3GGE6jM6zByLYjkw1pEmmB
s1qB/UKl1rLELX2UxUuWU60j+VymJ2LX5Dj5bdpy2hXXQXVqyBlxVSoXzTtncdVy
We8bx3sf50v8mwgg3tz2LqfMo0OyIdxTv4HLzZvDh4LicYOAA9bI09B+0p8FHvb3
J9KMiTK1nbdbAfyeccJbHabdNkJnFyGj7y6GzoB18mrRdGtQv3KBI6OsM+d2r4PJ
08dhUxhAp+cre5I94m/LE9HIoiwLABozwrDw13viwFzY3d8+IMQ571NNHTNhljGy
RigCI1IZ62ayFmDFNTYyFPy65G/ka/PR4x42EDFzk85WdaBt0hOZmb9DOi8PvAHJ
3ISEES12E8667MG0mtA99OIcImT647kXOuWUUWKmN4sAN1Q1MwgIRk77MStS37JM
AarGKarp04IhCqYvjB3gnWMMsumILWzo4QoNiY8/Evc6rgJfufG3umC41iCUQgEO
/x+pLoM6Twh5l94fNCyZm4FUNOFvrjRSVe22puvWJxsTvRbEp2Cx3VA1FHdaQCQE
lUdlnqVkkj9hBxwr4EdA0rO/6nUeOeqHPXaLGAVSLTcC3bhZJNPVflnshbjYPIec
5ZnY6fo6REVF4Te0j3J6kyfFMmcsOyWl39tR2zPWxe0qjt2Qy+0hi6AdNM4u5A67
l81BYW7snDQIUVAKB0NkC7shrbybZJhAzNziHIl48YB9bB36CZ6po0qDNC7r/H4e
fz9gMAE2tkKcjooJySnwWykVRgyZqxJX4qlqiXd53ztO6Q0r5adi3O/+GgnHc3jK
qbV0EstBoeJDGT+VYWeHwhp322nURO2a6JzcE1LAyDHKx5Epq+HVH+8IgjWCk8H4
IMczzagIE0WyDeuZWbDzi2zyNGfsXnh8KQ/9Al/tfLhYOeQcMTseZq7a21nCnhFg
9agR57T70lbgKfH6p7NBS5fqctP5OIb7m/GzP52QhFtjdqHSaFIysCA2dqwN15YA
uDkn2qtGdUy0P1sb5gvpBmE9kG3aiJFf+BBKOdkP3nn8duHl6UT0vOSjD9Sr6vKD
GhwBQcE9u7YQLOfIuA15yWSmbe/GAj//eL0u3LTfjXnzgDIdj5mOVUECneQpPyZz
z2dyJAN3P7J8YPlEIE4kNDPnZra8ptAMwipJqSw5rsMD4KiqtQ7yT6dmk9Ts0h5V
JXORIKvYIMKU+brQ6xLN9EnUZkMJinrjRdNb5Qupw7hUTnmE/Q2qLO2i5G/i/6r9
BRegWTdI2farANOr4J5CF6PQvepQWjcvTkhXx3TdteO3bjNVqWkL91nAQzeqUrRr
YYlBeH/yww/2yeyBFqgzpg1dqoqIs8gVeaBXNq03d8eVVlGqKOKi1XAfu/7ITML8
5fjetq3DqjIszNaSiwR6/d++L0g8yJkAqT6hGHmO7HL0psGa246x+tXWhDaSsWVP
x1QVaU0x+KbV2y+2DBA86eWD2pMLJfIWjILRGNt3kTLZbzVLJ79a9xBNIuUIpHeB
a5qj+58TGUYY9o3G97mjScNUYKfol+hueqjZ2WwIyQBw6snjy2hzsq44OlkwS771
Rpq/muK3K993kWSCgCoWho26huj8OCtOf0OwL9XofV5laB7eiizEZgEZzFOmWrcO
kkitbIgvWYSvc8qawkYy6FPStRpveTwFXFtuAjBBVnHMhYKdiylp5iayJY9855Cm
HGbLJLHsC98mJKQV3E4CWioh1bG/pj2uRVRBL5WFG0p15busB7G/WRqJxN3iJO62
td/gWCE8r/Qq8QWwFL3fmYh/3Y81jZtxBfKqO6DKdaDKj1ia8Zfhv0CVRkXZwhI7
HbggvV9J4fU81E9alpwITcG4Jyzd3MQv2IOge13tCmA5sHEuN1oZJRa4ivfd+Ivu
rHZJ4TjOtqA32yLEomqgfpJ+KGi/7/TXJ3FBC2hwOsLU/ZBS+nDDbnsA5duEuGeE
eUM+tre48l/sB7SP6Y7h5K5s+s4jsUM9UN5gOQlhoKgsmPc+aBkaNpjYbmeqlmfl
UIPJOEvkeSy9yF6433/IyGmDqUiH4XF9qPOXiYJlnTgn+eSo4KsMCW2TPcejr448
1qrvjMM77HEQPYLIv8Snu989zLkevuix49A1ullO99HJFy++7+MMulgerFvQojj0
RnXF5O5ttiurBZ5rH2T8hrPNTXVz7s6ZTpNyxqiF/oo3B0+PUpbRtR2U3FDjQ0PP
ayFuXHP1I60L2NALtDjg0NgmgelPzqlk7N5wcf12lwRd3gPhEF+nGGkuqnneA47l
Nu/f7KrUBBx84wAHAQAGa34krSvjEUiY4Gpl/YEY0uY=
`protect END_PROTECTED
