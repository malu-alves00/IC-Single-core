`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DZuGtdwcU982FajpsUzzey601tP47OUlrreEAWyAaGp519Ah014QLVUZqPjocTvy
FCPs6zxfoW9ghpX2PdHH7TXwjviKm65P1sHAqjZ++622SqKQ2+XJuJ4SADaA9F8J
sTJpvExB6ry8V1PdGaKk16m5nIxn6awHFqbStrTv/AcC+RvToi5xfSkj05bzkB4j
1w8NqSf+U7U1wq8FRoHZu5Ol97Q/R+UVhv7HBadNYbVFN+RUGiloWxX/qkBIcZD+
s8nya2nfO7TZ3J0u7eRXfvhV6g0Uo3L3uKMe6LyQuYQW2DRIlsdZrs/ySVLJOT5A
i1mUHSXbP9UFarDx/sfKCfEz7VEXM0MQB3yDqoTGdOrK3p4aJgfWfTeckYG2092A
3vIty63aEvG2019ykFNUbWKEAL+UOI3wjYSwDSrEQuksEZeqFJjKmP3mWGRWaRXY
Lvqz8rgWFVXgsDqxJFpYL/b9V8xb5dBvDzKnX3MF8yaZJg+T3OYWyprrGyXpPuS1
i/EOyc9+r9fGSw2Rkj4oMb2JczrJPQKpnOUy5b7Upiga6L3WSetqe71nVe10oSLS
xkTxnmoPIFBbrcjrKXgEQ9O0AHe2tCpRqdlvJyo/+0hFD+sICI7yq2Cv1VhEx/l6
gPSCuSGgwIHon0y7gqHuhW+MWH6z4TFfznavx2/gsg8DYmbFjULKWzEsWIk249WR
d/80vsa92xrC5/dlZ8UR+q8EZxxIDg7GaXfTq2xyNgmoR1jcA9sK8nO16v3Y2VbP
NAPn9ju2Z40lwnzMVp4vJonBPZhKPpuPPyRMDmoQP/rhVDU3ck08z/gsluWEPZ5n
OBqrd95cK/c+epLYMz1+8cfoQKWW6lUy+YWqggy2hRqDOJ6T6lHZOR7dNohRO4HE
`protect END_PROTECTED
