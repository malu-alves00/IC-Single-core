`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OS2BwPbvguk+PfNX4vp0fFLSiPeNPCqvQ7Hk2FzqkGEpZZ4qDoGkJ9KFwrSolTJE
vw3S5ft28/erA3edkTtoP/oQtx7LBakQdo1z4y0VzsmI3LWMjkS/eUON+QGNNMV1
XRy8VclZktQNQ8dej1rIy+5Nh5Ac28zFiOd+80FKdIP54n9kLXqDY+EixPGAH6Eq
ejpckYpi2rJkgPqsyo8YezqZuvwzT1h8d1oo+imtm31Z4NSFav2E8WqbP+tqJpas
lHhQlhLj9EGEp1MuQQIAAulBS73j12WCRwpEpJ4wZRWaByRYWkCiCCBaKwGTy+yx
Y9s2Ch3tAI9QJ22pUq58S7wwoXkWHYKBKWKznzDZPaj5AN5GRqciODlakstrJ0sR
CfG1R85FOA6B2AS73bFV+bbIP38XflBGx2BfVhDZaDHbQMbXNzcXUh8FIn94YEqS
DPn3ZAOvsfsFjKX7a4h8q9BrZmA3fVc4S2KZ6nNR4zTxlUtD3TDcdql44fulXXyl
SAohQ1bUBskFjY4aKXVKoT89dHjxzngcphiPwd2YQO/PxIJjeuTv7ZMjZqf4jrVh
tGaOksEiht79DOv0Ih/lXYnnWogc94aQbYuc8dSqD2nqEKwapNBRnZiWGQjY3Ap7
dTT2aowxOOCAXx8Yx3eLRgujJAG1cfubmgengCJFtBdMI2uxgr+HeWntPKVeP+W4
N09qSYsPtbJ5vOH91T7WEWgDwdf0KPy1hjUgASNmBFFtsxvzvSVpoAuCtIW4LURx
lKaSF4SyZl/hO1B21ujqzL/zAFzBdN9ZQEmDcE0+/Tl53j7nUf1NA4W17+PFsOCS
LNkvuxWsB2cYGN2bhOFbkdA/5j5Qi3uYKNidfyKKw+Zu/WTQmRN/QSPULwQnzbcs
imFqJv8kdgbBLjC5QqwCtdXpQis0ijmDnuhWflszoGY=
`protect END_PROTECTED
