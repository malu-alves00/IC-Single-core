`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AUBHyvYCeLgQh3Y14toNWnh+yAo6X2qEPVEoVt46lSW206zUHPbnQxr3A97gJFZo
TSG5QEcCTlz2NeUYlaAyzYAFjQWKTDjGDfYVy8b6oweTM5gxuaskNCrEdFG8/5DN
m7X6ICt719jBANec67jpyLyOu/BglarwVDoLRELECyMvPzBSLIlKMuh88wHivi3t
PgQY0lGYzG4rpN2P5mScrqpexhtUpCey0gkoGq8pSAb9M82To09lT/3x8Rlk5pPT
v/koyxXdYWJtgO+iKc1BZH/quFIc3OPGgmNHijQ7CCwom4VoFrGrE6wQbQImJAAp
gKZ44z9LIfdu/cqNyopTO5cy5LDNy4o7pugz1UkvNQv5Q7nnkEevgT4tmYIGbCgl
ab45m8tiPaQKcs9ur4Muh9NrWoiiOaY8/4ciqVTvCKX/Dnd1slAR6ntAdyhVrRJN
lpyOZDQuuv76mA0nU/2SYFXrnRBl2Uq6YI0HzwYrb34JDFPyBTLgLvO12VsjPsRL
citIt11u6qvTv03W4M5rgBdyBDGD/L9yoOuAZm0oHLHZo0i69Vfy61Q4QdCa182n
FS67WPEqP0ubmYIPBWk1fijQmStZnWutVz9A350dqfJjhbJCCnY6amFh+HMARF5r
Ku2lt4weOtALGRoaXPqnkIjQ2mkVPCilQCM9+3eNHOrASzYGEMBMmsjnSQvmDI+s
d37THGPakZG2ns/q0jS7tPnZrd2UxRaYwt33BYGvo7z12xa90ZONx3TMI1rp0rAQ
Bl+E0nMOoZNOnkcxtdyw5Oh0qKZqkBgTk9kX4LRLTQISJCw7qMFavdmWo1g7EqDo
FhMEcTF1u6cQtp9BHS3o0gX4YL9yW81So7H4a/xtHeSFbNhlUf8uGYSLPbsSK6p+
Z21OuLTEI/u3MpXw29xLtNoMBIAFVRDBxoosxuOP9ICTiYUh5L8dMoRzFdqnO8QD
HgxO4CAQoe5NZKyido3e6ybUGmXk/1f9h6bxMjKurb0=
`protect END_PROTECTED
