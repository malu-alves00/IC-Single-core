`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6JbGsIOBuo6I9pbs5DJa15eH9l45yXzB3NGy4RCDg/Ri9iGvP3hFnVr5o3yh0sry
UGJMvH8Wqthc93QuaJ/7Cmau0bgBxw6FoLgqHytwUxcjkyWwOUsGRRNE9KdtXWIC
C8GnDQ/H0+6XDeb7acIS3w78zBBOmp+PLIhvTZ8Rg9Ts+cmyJJiUI+DuHyCLVhJ+
CZrVdurl3NSDrdgAyZft5kzdTyh9bcEQmFfSyyYhh5kxVS4HAKJPNmAm7ztloyM/
6cz4a4DwptbWFd0Fi3CHpOPm1ylLe2QiW9i91KuswkQbRuzLPz1A5505/9u9PAfA
TsoUKqvuc/U/ASGfLsOz/+DuX+GUVuLADz3eWPTIv9kgIXYzlLsgeWbhP0TAFtEK
J9aqUzLCTvQZEWLW3P3dsGeBoOM3U7yG+WLXMrWfrQRagqGF3waI6l94gIbvniqb
qANtaLCFs/PQ02uFlabFOXXN8moIdj+Jpsm/j/chYDNCuyLiK7+5sS8SBGYu+w7j
tmmO0NT+CBV9sO6p2ehjwPmAAEHOaE0PT4mkOtAXKaHfz0K7Bd4F1t5zJMt/meYk
x5gcbk9WzF3sEvWxASvnKioQPt9TxrO8wL/XH1wQM88dLNdr3AA01tJaV8iq2Afe
FAZu5qE8ikf3qE2vU0RzL2IlRS/UDx9G7Qg7H4ndqlZVWBz/XK93f+HkrlH0TbwE
vdYkVxm/vjbfvsEB8XZZTK/uVs8I4AdUngUzBMrvSMoprI0pjDICtvHdiDWuJUBe
lxgob9PI///tAicae8Mmkk1MK578gVjvvW8bK1oTb8xs5gcrv8Jagd7fNmUZGDvS
UnVJk2jyxDHPcogFbSK36ckc/KXya7iQ67003Hw7WSHMEcEDEoWn2wUHeU+1Dx61
qVj9P62n2mdEbaedxFZFPv0y+cNOKJ59ERFFFvHwEIgxDZgLMSWqfIUtb+APpvAX
Yyp4Mey0k3MVQ2STmveJaPUxq6dcVWY4DZwBdn/eM1oxB8yjYL+9JFvGfJCRAUPx
REJDKVt6L7ns9iTxBKK6Z1dMD/3OtZ1wKZXzXiYcUN1OTS95NyaY305lWejH7b/v
/m1b9mWK5VczOXVwa/1OXGlFD0oxrW1cTAk6gtpPDkX2/Wb9rqF+3As3RYdltBDB
V+rr2QEN2PldztQCaRtDQ4VWK2mAQ7l6OYORyd2689vezA7LfIG8P6HoRhrSck96
0nf+pEW1QBpRWAZpNUNc4DPN0zbDpLrtUWuoyljk3fZsMXOWp1N77dwjSkZ/lMIR
CScsZ9DhZwzwl9Ib/ElBn6gjkuYSWv7KISI75p5aSUCkbA+jZwP27ir/u6Cp35It
RNJsx1A8auLmbGd5QVrQebEe6BxSmpc6PNJgzCnvy5fI60rsoFordpHXti+qvlPE
Yp/Ad6Q7cOxxbyzUTZOGC2rcozqKY2PNleUbbi6O2qSCnN1tprqNvpTTmIRFmIIZ
uu3oZSNora2hKbbHc3BilzSnrU2lio2fbTKWBJiZqZ8MJPDtE5fN3QtWM+EvIFUp
3jo5JDXsU2APZsszlQPr4Gp6LsRg3fpwYxzyFyYbb7IK+n8y1VHTXYAQ9PHaGyvD
htiUVhCtBYpmY2Gi8tww4ycJGR48X9azJtCXkolXQ6A=
`protect END_PROTECTED
