`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ls5ywzCkfG0yUjvPrrsP5VKWHHxGrdp9LkU/34GRLT5/yw4TmkKre/8lN/KOMuIY
Aw6P6VvDIuEgU5Duzrd1yxi9+pb6PqDzdBEmZ2V4aaoOEwdsOtxvcZcvVUSessVv
Ws6q+/LTtk+EvXFyzeRFq7WF77JUgjzt0PUnilkocbo7oMwuGVvt7KCCJHWKHBtC
F80/fHwvWmbdB556eAGLXI4DMHqKELE2x/D7krFx6G16DoAkYzMDXWQaExzYGUqm
epvS472N3X24EDvKx42TsnNJu2zfZTMOKTL0hxtdz5w8IrXwId+H/UB3D+LJMnvg
LWT6h4VabX03wW5a+T0pGXIL6VkTFP51ri15P3VV+wQM3G6tVKL+DK10+es9O6m8
lx87SSILWuHMCJ7JDulvu31ZIfhZzwJNLqQBM9HTOeNkqYqdUWvBLQpHdwD4yGX6
0klY1INpGCjVHoTq7qeSG4S3CIvXF6ARPeSzyGLHolUV6gjzpxFyorKXVZbFrg6k
VZzRiSpUYnEDMtRKfn9jZqKuw3MOggcAHmCqghrVCXpi3NwRucQafGq6AK6yAMIn
p1CtSFWpsqLD0GXph0jx4bUn4isJuR6kOmWfg6YL4opaxZiFKrQEkj0oKm7UGFPM
HQGX4E9W/n8a2jprbRpAA5hkCaQPv4bBOLBOjq7sJyYTPtBRS12DIQ6ERzgAdlI6
WKBEmG0K3HYIRegJxhC0dTRXVvAeKQySmbH8XmFfe4lJb73bDn+GDncE/ENF3RdF
rOSu9e2pfUKg3pzIphdH+g==
`protect END_PROTECTED
