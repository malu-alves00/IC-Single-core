`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1bJumcPGk+z9q29DYJcRdcRfrcym0Ve5EK8NtU3ArGQgNtN2leWW7WsLo4pb4+cg
M8CywDgtsP3eEjvh926jLTp220z+37E4gzRROJ3hml6UeAQR1GpOmdJlXQCpH2Ml
d5LrC0+qxt5pKuSiAHVIRBb+bi2UmMgI4Ral/U93cte7F38B9W4N4ZYc7apqFqgH
TPGBI0f7IMbYCf+bSOuirge8GAGv/pNwDA4aco2eDf8bLHFr3+vRwQgEDciQ6NaM
UHrRu04lu0qDeX6ECOaHJSHJJ4jBmCE44amUlKkkVXxAe8cIYiQt2ssVKPuKzlC2
/aCk5pYUug+IVdePRJbMuVhnh9AMtHWTCLbiplHzdkXaoEb4bZ5kZ5LATSopAPPv
CFwGHpMpxV+uZm/7A/PF78gy9VilGSvQ8NXSyMz0fDaIvSNVqa5Byl7UGrQxhsVM
9OSUxdXlGG+IujxSX+Qtr2Gob3hoBxBjHG5Izdp4XQf/M6ivJMdjG6Iw7BLVn+gk
0J42iK7unu6hMmMf35Y+ywl0oMHRZHJYu9KIoSQwyf0=
`protect END_PROTECTED
