`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iiNW8GATcOVq2t+NfR89haFDhIdR064HIh68cb6rkPEBuhMtBTYYPSfwH9KgTx48
IEkKoXwPDrr8fVheIdXccI9qtbUJ4wWiG0QJeNBg/cu1jxNYqaVXxUm17dQebezW
QG1r5DuUpMBA8cD3PDMU5IAOR7npxM4jseyF/k3Ou+3pZa2OfseGGjBsS52fVDLm
VILVbImp0M8XHI0NtzaGYC69K4au1erV3IoDI9BJB2+ZsA/4UWptkc9L7F7gqgpN
JVncqnv3J8/mN8qG4O6VR04AqbdSS5S2OwYMTKUwnd1w6W9tYP+gP/unAimZXuRq
qoFNhVsjbNRu8h8e2zq8uzTj7rsSw4H/zpFK7PCXgP+R8z55gt29zkbOVob9o9hr
xqiwfZF73PgIMrf48m9IXaCIHL5gqjhqCcmRIhL+Zu1zKwUCnUFgJeWdfZBLEbMm
/wXwgnBOeQj3xcKBbKtQyA==
`protect END_PROTECTED
