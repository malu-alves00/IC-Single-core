`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XHsA6EiuyWtWO622qZBPP/bqD7qVaPsk8VumnuFonqIku3SqGy863e7dAliNaLNq
j8z2L/KkqL32FnR+/3Fq391sOOsRQja4d+iqvYS4qKhDV9Pb78yYndyesnfuqEMu
cHZN7GCGcpYdxsWcUCGU+ec8BCMB/548siackslLHyuw3pBe+00c0d2lvFbDn3FK
9+9aSpxdLijshIK1dKKo7n24fbt5abbN4jF41hhtvWvrRqg11djy5PDgIp7z/UPj
TLQuTj1WWbxSpLWxzawmu5MdQCSu3XRgOcRPrbvxI9V9mFOJPnrSPNE7pWYX6nG9
hIMTN1dGeBlz4LR9AABhVTQamIuhabSmKp0L50HuaNJaUWzohkd36mT6FJE3syQy
+E7mo+P6+hjMIqAUwdhhGKC/0/pQi+/ZHbas3RFEYVWcnOiTimZ+wkOhGaqrY6/3
8NsPjecS3V0Rif6sgAwAmzZHc1KseJM9JLDDWC4dMaifFjvvRIUPKMcfjfeFMPfk
taPUh0alLoBapnCoYyOiOlOYpMMLaji3C0idwxJKIiW51NtDKFWQkXblseli2ngU
woK9oVA80qm4IZX9Tj+ei0v5IKZOIVZzS2iRnkrA0adF9qYR6OxJVgSEZFmZnPY/
GiEJmCahEm3Qw6w5M/t9bw4BGC4hO2HmBxyIVjzSElfkTFMvDvGFOfPTOWHZRBbs
fdzA4uT9h2NYzq8oX9DfPcP5yGsozism7KkxwsDsFXWiaXqpwTsVqqu/ukGf5MQS
3XAtx1v3GwY6qT+Hsqi6OZMASMHULrK8u+zJ4VqLS6nLjNz0Dhb+a5s6X/PlrKKu
OcVgiYH/e7OXHLZrhKIMc0xY4qv9NwnuN8tZygRnAYKB7zlUVi9MD0A7MMu92tt1
XUQKQ9+I2dKRgiT2NgtkH1ZXrvWHudbY9VnJoshqwcANvDzGRD3D0EtdkkAyJkiB
dc4mW8Is1Qs94PHK7Nbb6MMOQDbmJN2e23cti2LRi9yupD9eI3BbGgnmYRLNqfwp
THCu/XfE3Lcth3TNpWzloiqfg3BoVw22NIwwyjGBHPxlbUWCl8i3mhquXVlpSjtP
zfnTY1apF39iXgLQruMPtfeYtOAqoVtEiGpNUy00kX6VQIw27c4IL9gGjALWnWsp
vMW9dtm0MjnDsKUrU04WaxsVkGe89jk0lM55pSrBZr8eu6ngYGxHAGvzjJkJGZ4Z
Y3ADawyqnfK6mEgIEW6/Jvr+khIOkd6xEftLZnS27ANsxyiqk+DtVzOZdHIG3c7p
Ltk2/u6sHv8W0SGYryZPYKjunPP027HjGebd3DRe8i0ZgC8Q/+Q0jNUurVwzvnYl
prxd5p5Kf9A8Y82DszeOs09x4/tlyGoeH+qlEWIQ+eK9YTarV+k1FogC064GwBob
Na7Jj5XqYeWlJfChQBNbLZ/7ZyrMiINZqiB8GG2iffoV5qXs94Y+cjhct53giVOH
2t35BDflN0PwoCzqlzRXWEZ4773g2D3UpR7GrjJ4y5bIlcnCV5kpJj1CjCdfstDr
IlD6T2wfuvwNxyrq95pjfILvfEnT4njzVOqc3XuB1t7VQ9uZtF6cU1uiwPKnrN0p
zXgvpRgHJwdv2K8SVbKbVEzetPF1PL7IDFxXLqnnJ47FNgCyMcCj9PWp+0oDIuLY
eAnIjKwQUi9nUKw9AHxk8i0D5qmDrtCyhEFpiPrIMYKo9ZghGK7mSY5FtxlqhCK3
Y5lVek2xAYKhgj6ZwQ6bBmBV7s5pLRZaD3v6lQcYMqI/3bdGkLVlsrpElO3smPsP
J3F4kM1jxbbEfjrOJo1MOoN3gTskAmdA1IqrJDrjDs7bdU958rdOr5gLu6WUGKD8
1eVYD4MmaochQtzIJHw2azL7VpLKjumju05KH6zBKH81Lcv+/iCsWFdJh6ARRfTF
p6rPsrfFiLICRdDUzybn7rnb5lmp8OdWi99y38tufRq9RB+eCKADMSH9L4t8Ebvy
lhH3qMVJ7Hb+0E7niBzVaHPls78XUbjVusF14hS8YNizKtI5xcGVEHc0DkohYcNK
PAKZbbM2RGym7pHb7/hYTK0b20+Zpm2oDB5yEo1kJb32zyesPG/syGFpz5s0yiJ2
DDEwr33XyOKnlBGI8HlWElPKf3RDpFEsScKwup1IEWHBc53DgvC41gdAlkt3eQhG
fMs8r2hiyqlPPgOCI1521eQ+reBebO7aLff9SbRKi0ttdYpQfk1ze6ZGMrxr/nak
WV8otWQ/UXnk/ZKj3FpVtzSh6q6VnEhqog/zNriCxumMOEBdIowgpfz/dSwkg3AN
wCgHaGSEOXAn1+FVb5qNacxIphxE/P7N0HMg7bUJ9IJTTQ6bLHXy0Ax1Ri3+TADa
0l0C6/c3GoNlyr7w293lozoYxBspJidbKJO6a0bPtvKkwm7v9E22KWgjq4aLNMQn
Mhokjxbd4JoRosiIbNErUvhiVPe6MaAsRKi4RmYnoToxwUCI7cHLUXkrV9SRrhBX
/qXoVWSFCe/tLeKQ/VNYPDibRUynvvxTxQyqY1NRQV1FXNk04gVN9Z+ALGQaLtKo
Aa73GNF1hp26wVIaD44AUWfeJlToXr/D2m8S+oD/pi4p8i2LQ5lRpqwbAfBXz5Ki
grjsaJClb5vuD020AcMD7rD8BzV6bFhciMbch0OOaCDtWJ52+eXgxjjfiperMHM+
o5dWTbQyMunkmQ94VSBbMd0FxYNlx6Oiiy5JdWFjeHU6j47GB5jbr7Zx49N/8Ksx
gcfD2KyStPTNWwQ/v+RY3iSWN+sY6JJU/5GiCPA3t3re14AfWXNopVVuRqqESurk
FqwKTej5Cc9sS4pahEPDryCgTQ1pp5zzC1X+vOSVvoAtUhi/1NQ8Il2sIIoOwtjH
`protect END_PROTECTED
