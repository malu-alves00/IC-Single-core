`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YPWqf0la0OOWdC049/qNE6OzzNtQaMUVf0RCTpnojqn7CDot2OONzBJIvywBNJ/E
32pNsdmhSSQrCRuYqf+N/CRBz4OyHK55MnQvVcX8iM1Ihm62NAxtL/+dsHLu3p59
847lWzJM0HfgeO280Vetntm88/L2YlX98/jjMqYMNSinimmVg0lQ1Z0YHlcsPRVw
nA//6TScIVoPpiwdgfgTsnkSd9lD/bKlDWrheCHmJbQph+Vk6E6BZHBcYxpuA6BO
leVacqbGoZU0k8pXOUqu/ktaY9xzgqvOcvjXL1CErLNWjxT8CZA0g0fJGwnHh27W
pNIhhS0MR4aGGFMh2E8m5zHC40sWbfIr8OSeNk/1bPOUJ8vr5eGLz9zW0hF1oRO5
4+MIue33lgaIQhA6NEzHXzqokdH3hUs6HB3/5ata9d9NTU9fS7Q9J+J6GbyVPA0K
Ty+qllXpEjHTEYGYkpQW+dPUcYtm+66mGrsS/gdi7uLE/SNfpPJj0wPyUqCe0o/V
yi2fZlEQMY0Ghxkkse7tv0HGAditJVStk19SJEitpRHo5O3PPYMjVRBDXoXg8KQs
ix6Z6duuNynfrSA3J2TQxVb5QmDJySoPONB5Ebc+cT6Mvk5YZsNKMyDGJRi9BYWo
M0jeMsPuMyQA3hmxrx7LuwDWZ+PXZFfLbxfubA2W0yWZj3QqcC8hzbF2qXUcZYjE
KRt+jhsZNkS0IU/QjH4AMD8wuO6r+7RZdZ76l7Oc5nAGeZRAznsCLaAnSj1fOW/z
dKWBal1Zx1WFzRGICV4ODyN/KgVryJ2X6ztD4lFpm8pEzZUT6ymwnzXnKALqxWkk
boAdMclMVsp86buH5fcjP7Ofu5oVbQFB9mKRejy005IKFWdOulqwg3ThkmlNe8TI
Xkb29X2sqeHplOYpVdHf1syWlMbp2NGjnu/j9mR+STYsd5Et5c5XoVb7SCM+GOQY
/fHtp8YenAni122j5ojft3r5D8JnwlAKLgBefwdHy8QJzKFE1Cj8MhmgeTcsHgEZ
oJThRR65kpLltqgBgwUI9C+3xzRmdeZCNNXv2jJ9ek9sRkPJoxyFFPCEeaIkZyDZ
1qmbFs6sqBG/jKf/YDTqpdWOs3EpsMyXpQEpGlpf5TGaCuDyfGtWRpQ9ZUCl2giW
PI71LlDKbYB9lnoR2t84LB0xEOZ+1/3wFBJrfUFtWuIaVZu5Fwsu8GXG7P/wbRFd
W9XvcA/z4vAPO0+UeJoTrUwguB6+X6H4c5fxFlA+Orcszn5CH83m5vV0ZMoaBC6y
n+Vxrht1wL2Bg6eOKsXSjfM0tQN/sBeQ10LK3gk4vpbsXNZLu1xYyhyaZd76RZpw
OhzP5X1fHiXfHBIks1hu3//eA1loE9usKUjorbN5rpk+kzJb+6hgxY4qiBEzFDEt
MIlWxcSArEMq2bAHLWVRI53ma2UzvFTGniMrxoY9lUGQtWAjn9em7QroWBZvEII6
G1I5kYGSdBH1o7mVUyartPB3Kfc5WhCsXAAypeGxvfe50qgTYiHMsCg1A392dQ4M
bvZBEiHVMOSexnhxelPbDW3wAtXk5ar0fUWNo1mfN9A96cbHuO5/9dEpC/bfaoGp
HS4EcfYMaz7RlIkqNDxlC6p3EWeBBV1ztMYROmZPXc1hWY0/sXBXXBeuj4U7BkTk
erx4uTtsk0cWK7YMNg0372sZeCWhYVMXY+qJzwWpEoweJpVs6cYzvyMFLmK38R21
qjJfnRjZVG7S8ZMjONE9zlJEwFq05NBWj8kPASd9C5DPt3vPReVm5YGUE6jHGLn4
I274u2/o0ozgmBT4zvzLx54qWjqEf9KUBqVF6bKk6d2EpAcnfSdLMF4w95CmDpeA
7OnJWMO3OmPtetDoeCz6iT0LzQ6SjfmmqhtgDMyV1SIvEjUClOywsayRMjQ9eeXs
2nqSa/7mpy0+d0FSHNgecQcsGy1PD1Pk8O6h2KI8kPr1fXMVBDi6xlnF14f6m0N7
n7bsr3+0CZGv/IMWJeuXqC3UHmzbgksIk0I2QE/3zlU/03BiPv+9tDPY6Nqz39ag
cRRjggD5YIKJarG1T4Ut7TqgRdvpmme16RiQ7vs8GHO2/ZEVc9xaLeCWNWQUuUiB
2XL7fjV2X023gApubvI6jzsCoupBK5lt7e4TTUPzMrxgQ2czxhHCBag5auSD8ZrM
fwVAaXokmeG90r4kDqbkshanZcZBlJwM3RQEBM8c9rrG/cCZVhGwvNZl6Rn8aTwp
5QS7NY72fW083fUKQmom4lsrRyuET6S5QOaojGRn98FNWPlF53a21J2Gjez7fP7h
dF5qKWBs0lphRjcf8c0tPLtG7EIDUknaCqA+xQumVG236trLibvIkwp8Dxv+AVL+
JaluZMxtoEcHXc9pQWZbrOyjmhSs+nZXksp4Wru6LSfiqenJNGSXu18ck9Kz6Hld
s2LbfY/6lYKyL9iGLwxpW0ZRnlZ2UnARfI7UuDkGxJSoM7y/qGLHBR2oez0HftVZ
c97N6Gr67RSF8oPHeSlS4qRxwcFLsk87tl4PaoBdsGeI6ZXs/YE+Jda9cHYeNw6u
D5/BE0aHO0QK7jRSV+MWgMdafwdpZNCnoNI9uSGsBHCDTxThgGfcXvdQ55rY3/KE
nlaH8zMhHLDACtmuLpEcdmRDof/4bR7wPzty8mzHlx6gI3qklnvguGB85NA+zsUH
CfIxcdCI46zbA7yQRYDx0gqIIcBMhFGvDrw18lXvrdVz13+5+hRr20W1MIwM21dn
xIozf7Ejxh2OguoNpFddGhXm9eFVMUnLFgZF4nMmOIGr7VjPgXUwF17WAoOdFOPl
oEsW/TDySAveejOC3YGfdKVYSsN6eNGMBZ7MaFy3L6b6jYEXWn/eFzvKOlpXYAZj
hrtVwElZbgrmuJrECCuKcGbNfRpGWHvuHrsLjudtrT9fKm4mg5A61jaaQJBkmZf7
GoUojHEv+NOlNIw7BBH5HGwkbY03vpp8zhxX/BiM6ZDggnoRawjC+vntrk7fdYrp
B0Uhhqo6jnnrzxkad7HZg1D6DNXHu6FHLoSOo4vXPNliZ6F7+XqHmtPP1bUSaGwq
J38k0GC3+LIbpBIEsZC/8BkC4P52dtpZiLolwe7qBieqc7vXkyDIa1qV6z4bTT3R
C8aXMXqHHRCDdCcWHEpuqOHdQagC4j55zrRUIKHdVhpUHBdCZWE/J0S4HoSZ2XDL
/tfFL4CmxiLgxENqjJ/2ySmXLqCFJMErkYcXojiyXO/JbRK33RyhDGCb1uRVKq0z
1C2uwF6Og9RQ2JL/uvgqQdPq8V+mbjV85svJ2y4T0DvvTVRb2PcoHIMFprbopEpX
2ubVksPSG+OgR2/hDFVEyw21FngfqSTJrXT9C/9yBElXPQ1DrZQN4hAKb0O/POWV
CT74MU4mGIF0BUcFiHryv1u1NqdnoMg1z6EpluPp76Q0Bm57iMxgf1XkjyLxoZ2E
59bUClB/qlFN+dogylqcb+/aUFxps8fOcnjcYoIKt2Xm8c1we+oCF05SW/ogpuJE
ZdVJN8nkhdXcZwX7+z+oCb3sPh9M0ODeDWDquQGmv+iIvmlO3r6omzjsOywBe8WW
7cUS5cHckhj0uBC/CFDD26bpYJ1UJ5N/nrwUDJmhOUo4JkqeXdQPALny37sNXWs6
/jp5MA325Cy2oknXexM9EpFEJGFQ9vSmC4T8wRh6U3xlzl61z08XKE1n5z8BoYck
U0eUOQGM7M20dOBptHD52jD4quePMOM0fZKxNX4ZUwj2Lyp62NWkgn/3c4KGshN/
9FoOI5bu5jaidJNeGfe06dUQfM+kAOjkunCEtJB4/XdYYYPnFX4uFe/94xtsiAqm
bnRmQ51u8hufCQWiw0RYl/DSG/xpSnwtBQTqeOs4JlWysscXqJr+lh12oBg89arV
/WUAKJoRNZcvxKwGiN7fc8fh/3TFnUzuegGJWfjv1Ay+502OPEwrAawS7qrBDr5p
Ropc1kx54c+IcVplDwHaWET9ShBvsh2z1iqLopEVb/YM+DZC/Q9LsCNjJhvusPY6
/VnkJC1GU0F1TuU+NJURWwNMIC1yVv75KP3gY/kNCoU7wSPQ3MiRdvnkRl7RiHxx
iIiAPjgoooniRZQbkhJwfKoRb1D93oSLnLNtSCe4yPnaGWUrCvnJhjG0jt+w2LEL
buIj2rqDJ0bg6QXnHH0pyKBTRU2iMhTrGuJweCyT40aWYKRBX43GtlnR9rMmhBrl
xU2EYHAOyIwlDjLYtx3Wl/WsGCu5YGk8x8ZJT/3in+KHDBpPrLPYPB+NDJPz7qkU
wne8wuc26YwIV1GPqCyrktVdKLGwb4aMCJN5YPo5yvWVfgJ0WocqWAwJ8aYUg/I7
lrphoxqY+lnyAjis7K8H61XNd36tlckrZFQ85BIxsOCzEwmCLR2d+78L1W5muzy1
N52/tq3Yz/kIKNtdicWyKvbwDpLkYuT3SQYPpaPhCTLOo1+vdafE2Kb2S9P1Z6c2
IHWQ/XPWStTs7LiHBIZ+gey0iJZumLHIpKiXNmsW2aTO+w6p5m4s/DDdQrmJQ1Od
n0VwKEfB29JPABBioMGIJgVypIwZbkXopreAfIOK3jFcO7EaxTtWZ3NWd0jOjMFD
JrFE1nZd7jYW2OvDAhecwbUC7GjwC700zujWdq6KrPWcEDojEdwrFTrnm8tayk7O
ofICLN9hTVFdC0/wUV/DErEdua8NQ80+6ZOISmmH+7+7jhstzUb9wFu6+OiYXpBO
BROk3HCyH0yeaSbI5BU1ruwYQoDvYrS5E9a1Q9dVT90QojoTUPlCBBqDjcz+akwi
Xf1OyiKXgjX7gW5/laepBAHsQFKhzrXfc+tJd/0zoMZ3w82d+GgveARstHmrjQQ7
Wmy+p6nt4d9wyQCMe/mTfEkq5NKJQ6vk1uZrSGYwl3ek/dbE+zl5rjiJt7PejfA9
YeOXqap4gm1fnffFxcVTdUo4A/gXIaXst29yZ0eOdlwCHpPraiv+HemG+XoZVb7z
dktPwQuy4G3s+wlhHE15MxLf17Bm0Kg30mFwelswEnIX7wv7zd/5724DVaJuTh7k
6ePlplixBaNmo2q2buhZ5SOYk2Oq4Ml5ySRtERN6FYF+/41infe+5ynJ3IRj83eK
YdpOiVhJ9uQnYzIfK7ZIrazL6eYIb6BBamAXkDLDOvVpY4WDdyFSgrELtoAlDJyc
Ge5MroKRdZcgA3txHsKlpa3f7QIx/n0dGUalEHEbjHGG2eF6TyiYRjgFNaivUHbQ
iOSHUSCdT5C+4qVJk8C4pmwIaQiuSuYSdW1ALYT/QnVZMo3KGAarzibol/7pgeYo
9ipjNqa+O5Mngnpc90aR7cwCfQD4bkvlrD4MBoYiRDdRxR+lb6ft1gKv2rarOH7h
SkxO4sTqhjIkexS61Pfk9Dn+TYSRZ1/d0i3XRDZh7sq5AArhuYMTIvCNAFMg1fwr
akWW3eA0W54K22oBrKmbEz8GUW5w47IcgYxJCrCsw7hVn3XbWM50IZGx+QCCN7G0
JxejalldohpDEVdT2rYMzUGats5cONMQhvzG1JJ7yBQdlSIXzhbIiWLRNll8z0Fh
MMbLGtHxo16Q1J9MkzinOj65EVvSoGGEdKtDl/BVXLZ+0Vt3tHQRdhp8Hb3B6TVn
jXlI2Ehbglwjn6DtMBPSDuKUJhBj5FOIvuXCamhzf+sdytwuUQr6cpYGoenJtFev
zerr6p8V5B3LS8QeJKbAt5Ub1sJPTsKoPyEk9Va1I14GXDhg0zUD0UnS0avAfXvX
vwaHMIsyuOHi3S/+n+z2+kCvUwWjENTKvemR2d8+Yn6g/o2PM0DJ20qnVLWXAMg/
hAf8Y9Cp4IcN2KHX8eXoepjUc73nx0M+/B0FGZbm36wwzz06fZi6NnX6nS721vC2
7QmTk5+wZEGVehoMUcZHxVIgHRj+/PpiUF9Kzc4tag4TL1eX/QnqrqFVkyN4sE11
rAoi+S9+ikabUD5p/utZ98jX2tt2blZY/6seE8fCu2tjVzL4e4SMx0VMesiAjiPM
4/x/02ZahROR3nHEpqjcpSBu85eqI1v9jriQfwppWkRTuzNyK1wqHRMWVUJZTC8t
vEIHR3fcMpfu4WPam5X919j/ZoH+Xdz1RuQl6HQz97YO7r7WMbC6pimEV5ovXQrY
31Odi/N/6pftsS/9OHq86+GuXe3WVF7brMldAPUkF2kKoNj+r0JaRdWktnAROGpb
cIHK2gWEMa/imxbwrCMRGd0hBGgDt7RfPFQfhdiGBCWaSyxK9Sn9YYoh9MnKESUz
v9IuEUfWLLO5i5XK2PWu9XPGk3Wtd1t3MVqk3ZPFyHu4mm8JRVBdIiOfSm4F2TJn
hqTeiRA8WnAsDUugwZvp1ZGWgIzPAb1O4/giKZzPaLUIgEo8Q0FTUjordEQL7q7o
JbBwjknLTuSACbgMjHRoQOKIxfqCFYCfiO8otrSrz9mYNp+brsk/GV5bmBOxUVrh
ocz+JcBEY/WoVpdco7rKS5MM97jIyjr44ARzgaN+tFW7PYYlQardAAMWJlmJ2bII
o2jSJEO/GxHB366+a0Ecn+aq+c8cY3S8Q7h26TBolzwzcpOBw40GH3j0pK7BTVBL
94Yu+S3bUR0Q0ZpcmWAu9Jzc9zS9l4QL5ZJPcPq6+lyfvq8QSqVv2Hh9OGXJ412r
EK6ldF/gBzQsG3ClbV71dt08+t7lqaqiguYp2mzpI36fvKq7aK6ghaZJFVIPvzm0
CIQ7ZPBp+8ZzY1FHwz2DLVQ+7b/HtA7t+X9CiJ8kqxTE0NGrd0x+4mQ35pcdrz8o
lIf5cHSf04IA1aoGUcX6xlFO1QFb0cz76Iy5vjPTMhZaErJw5Ssh3YiAI2LCeq0n
/aCO9B7WsKV5zW/5Jmx7aNypf7bvNYeP5kY1x5wrXr3vK7ZpXZSqVFXj6ZD/01X7
RPb9ucIcSWtnXT5ZBXN1/za5bJis29EAM/HbBmzch3hV3CUsMFIhfAA5YS94n2Rk
NwLpHKtsibH7qGE+R599hWYKTXh2QqHKInAgT7GbAqQ5uhcwgKa24yZzAF8xRvpc
L1PjF9BFXgyslC4adGz7QnY/xJ9kZ4jv3chxNZV+XZjL9iiW1JQC4NJkBdtu/12I
aeddYrEQ2/HIINzli/VFpODkgaepbZAL6G0kH4dKofrU9kRIPm5F+T4cYhiT9lTF
eo7mKB3ob+HBSWTy3tE/mQKI3Fh6hwPfCoMODJ3o1hrvk//pQ3Bzt2m0JY9ar4vu
jQQ2tEMHg/3xFKB2N+WyhklImzqdVpdlgtlS9Bm2VVubGeuR5G8F3N4BstshUXsC
0aDPSbAjNR9hQaptQSyz7SKys53pizsabzEYRk5cwLAzdHuhPg81o/EYBbp3YTvp
lL0DDtnGavZSh3Ysv/MmYdS8dv2MHMPTCJ9JrbJPxpOm1sVuMRkMaVFaCEKshZVG
xV5VZjdYtedzxyk0j6IjmsDEoAoftVLA3n1b72aLpLFsQZEcV0jvJ6JGLJYk0ynK
NWhXWi/5riZNDdByu2HLX7hrxrobo/KWLi4JvyF4QeYsvHrvvCScxAavwz2PB1xn
0yZn/ysWSX4Lm5WxnMvugRm4uSRN2PYPQqw4kv3QAF8JXfd72IoQWbAYfPadilg9
VQOxZeJvI7jdMCpMBrwUrztijBJYIb+mg8jOvg1ncfHxYNEyEhkMwC33XuA61UHd
WaKicEH0RAW+3hCo7JOPCUQjvc2sr8phUrMbr9V6prGlNZcvXAOxCBXJYHNGok+Z
yquiqRSp9c/8cqWqMBwYmAIV7F3JpUOLVtdM8oda1M1a0TF0/5kp6PnTkfwVPjYx
JZe2OSTu5VfEaGZz6kEisKzGwnTia2O43LlObA8XxoWrrN7RiHU5pk6rO/V3nyd9
a8hpcFqan3MdqAWgvo0/z6tnMvV3+9zWqMukBz52T/wyADl6qjtPEmKaL/+gwRo1
qu/nB1s9FM+40RFtEt6q+S0tCnwb253ePMmgeExKke5zO6aB1U65XK6RMk4Ti/jC
GGSvW8Tu3seU94/t4lrqI3JHltiZ8c8pBi8seoLZtlUy8qy5dn24B+sNNkXpQ1I+
yxAqFt1kucMoHszqejBDSulRwhybL/H9I86K1jUcy3T0IiTn4b8GiWQLSrrdOMxa
kHtsDPoqXEEQ8C9fiUYE9j662jUYdulA6BveqW2wTx1M98qw1GNgER6H+CrP1Fx8
iX8iZmFpggJmKgsKTgOdtYyqtx1QIPqEWemuynaogZRELTPI9onOAUkTjhW4EYGq
Ji/LABxhcwRpzYM9O/d7rPa3VAiK/p7xA9ai6qsHELrnZtKn2JKLH0e27G/2aV/O
nSWfUKLWqeljyzlYnkSKQDy/KQB3fH6FnGaMM4zJeAJwM7kQBilyKgWHG/H2AT0F
0stwgqHDdmcpAmlXl06lorLNDuKEM1i/dzOXI46hAFDXhKMvK+fNB0jvpDSk0VRR
1ohAlggHx+61luOv4seVu82qY/+FL7u8irUN/g+h1gMyX/qDGzIUvuH10mHsvtai
3qTv/fhmvklROaSzFALMMxo4eS9XqYXxp5ug6lAEuCGUv6XE53u+3tE2ViAwtlRy
UJyrmMhvWdjKgxqNLYWHbmINNhZzaOdT3MdMczJ6KEf8zlYAcN5Lfdh5+wXcaOUB
zb5pRX1zIXJH3hqemItC0jlpsgBuV4rM629o+Ziu77UTbwGr9wzzQToIAguGNw/U
HenU0D/pP7Sx0hYBun0g/N4S+mT+2/KYOQDi8er/ozStwx7lJ7BotGXue6a8uxoU
abhAyUizDDzrO9kEt8BiYrHS+xc0JecyE2D7FDFZtly0IcQCo2c4WCUNbUBinIQY
RGXJxVsJYB8j/uFCrfGXBXuzYqMgU1Z316ibLCqv2qJtT1QrmKJPYzSfjZJETBji
tMWPzJFx5oceGDfj1bboxNCp5MPB9VrkDLBI5BDaTvLHnf6bQhVLhaLeV49dRCjb
QyqDzPbUToIGVny+sqkWqyGo2mw6UzatBbSR01WPgpJsDGeshKGGSmFUUfy+f7St
bje3M8TC3hniZRQWoQ27jmyovIrexohiwVgilNN322L1JlgYSMtji05QX1UN38j2
7dOjvcYS5MIfJzCIZAssGT0Nr3EUtLqkOkaJ8WrBXEkx9Q8olFnzhkmJ67SkdS1B
A7BQgSMioqil5NL8fOJU8wKKWvOvyb0NuVEsvnGt3JtabKZ/GR8hKdAeu0OMSQp0
ZzjSfDjOn2hE3FwMbLBPiym3WBaCxQeSGbDWj0AJQW+HYJz3tSLHi+i/08WBoF8L
2kBnqzUS/GJORZrqzWTMDtMhL4+ysMYJ4yQT2N/VZk/9xl5rQqAgv7PMxXLly/3v
KK/veEtqHP1BMHgz2FXfhcKkV+TA5G4uI63XH3b4307eDs1+k74IFoav6M/SztAq
OthWf95T3wJNOK2Af6RiZdcp8jShHn0M2cmUZBnFUldzJXfX66PyhCVfTqOOaYll
qkVEcUWhLtxSfsJEX/SJcVTHHShJV5Bgf45vbZZbWMnyyvTJx0nuWz4c7RxXN/b+
1H12lDg/zQf481qARg3qqRvIUzGHSm6L7PTtGpOIOy3Fm4xgv1qckbhD20lssjao
qYmFKrvP3HWeZygCkJdj3fpbctZBfm3ckibwfSQ63BnQX7GruaFQHlSivmuL4WuC
OKVQ3+mNOArx2J2QklWHbsH/wd4JyswtBli3Nh4j2p6pxlIT4roPlS1c4jBQTexf
X85/eVOPAAcamjXK5rL8Syj5qyWgwwNq2pAw+E8I3Y9+RwDBT6X/8ij5LdRGJFXL
zvkenVnmW8XkE0vnNODaILHpgM1CoZYd5n9fKN6Wm8jTgFFcGTtZ5GceFmjNiAeO
nGQIMQW/ppNm5nhhVNgGqfRRtQqjAQRBvrbWCRN2WDLpGAfPq4OoUsVQ4/LCST7p
KkBGHCQAPgcSsxxjv4z2XlGpGbGuZJ/ohYvazUzK5MchywdY6wRRRBQuKFpxBKfr
XP5xVEllHATRxoyY5MsBWy4TFWhLRBvlfHq/bRPExAj9eer50+J3Gy2pDOMD+Pl1
nul1IBBwH7vqnyVZxAD/0Stpp0BrXMZeVdipid5tquuGIFQypzDXGoxR9iCbh+0v
v0oZhGq3eUMgXOTbs7EES16HhdASLNon3FH7p7fCZ7z4pe6Qqk7uHPA8EO9FJb49
vbSjQoSTKU4FKDRIg3Ht9SfyFHDxHyQYAo/ouRyksfUyg47GnEk1LQ9y4EuNTnJD
3/wUnlQ4aGJxFnPBHoFXZKz923tp9Sej/0bUxFBVEfgUCmxanz+MGpFMV5gx5cTK
rD3Loc1mVyVtarw0tIPG5fxoezNpzHFWLFbaSTMFZ1uXnZJNB8cYCYp2ev6qrzsS
v5mqwC1WxppONVPq0diBrJuHDVFELKj/Dt8bzNpgujBJH1vqDssLVKngBzaMOyFa
3W6dzzdKhpvmdVJUgN4vJbbQvUjxQQYyLSJ0mm27lBUBgnMQ6VkTRTK9Lg5AdWOl
rsbmzzhLXxi9U01I8EDUd3hNSFnpdaWul4ng02K3E7sXOVFYioZZcTQOUk+hwXCv
PxEuoxoI8FGZrTPQvA+/PFHo+DFij3Kd0MleVZnCk3lu+yuS1XPLWJkQZRTKRiNR
mvDNYeK/C0mUYKdt2wLpvE6X37VkntoTdcS2xkkZ7St5nRf7uNo2R9LZ5IWIYvDe
QtqTgKB4LOS/xMHRjPND8Yzy2HDdO1enjCWQV45mtuHg7UBSTPlRjjG87HUaBr8z
2f/4MBnowhQ+4GJNR0kUxA5yRhOrHD+3rhRJ0156NGHJwWiSQmNFLwoCOy2NR8/e
nx5sHPYDVFBAZg8ML0suO7MxJM8E9rodh7UQiiw4kMaguR5lul12BkXFetc+UDun
/WuNEzlI0UiTHdidV0IAOZEPwsnOLi4cQf5xJow8WUctHDb35cMMDYKpVvU3UERw
+WCOndsd3AMZKkMMBjf5PSUtpbCH8se/Qfp/Yth8l3Iaj010r/GZIY32KaTjPvm7
/8UVXWzTwY5c7pqMuQncL1V68EEt5eMDn/0bbad9GmYWrGBvfgJvPc2FbMk01Bg4
SSXGWRWljMI6qkrUEq8pVX7PmVtoGj4cpYwtfgF18vpzf0yLtAmxhaP+9xytd/Tp
63l2xaQ+AAmTe1g6iK5GNE/6BoQ6NQOtflJDJIYyEpBPP9SIdWR1m3gqfgJQXLeY
Ulg9xOy+eJ+9JEfAfU1h3AgHXzrz06efbHHpgb9cXt4vqjZLEfYrIuI+grvTG8p7
j9bgvL3Ei0bJKEXH8YLEL84C+HgrC3Wq6XgR1n3k/OLiCygP6kFACtJCpzeFt7fy
QXFjzFQawvDX3E1f1t09vWBdrOFpCnXdjvVAHkHFzQeiEtCHZwb1mlq1DlpknMfM
yWGA0zQFdvBqBvHXUDKpmTwgoMYrShER5I+brMpIzss/ukSRW8UQ75FkA32JCQy7
Uz3qy0dVt70NOI8CS6pOs7yKMYJ6cR/D7uTSNlRGlN2V8QwH1AYeeEVZ85DCiZ0N
zXJzUmqXZmc3FfSRK934JJEO0gajWeNDgPgUWFcO22EfkQ6Cu34UN549qRZHAKVu
0dOEs0wVo+yfwvZJr2EvDFYswhylQeD5mEsywCj32iOzoLObCIgiFDIvpVlLhDGB
TS4as5ofV/5AWu4Pctj/AFx7U4oFEnVV+neH2nCgzIBTLOYXKtZyRbEIYW739dai
lUNL/RiENGfxNmRMCl1YVI6t3LUhQ7wvzj6xN22M826CY4EknNKmtogco6Hvgt8o
kwrGsKowhXVq5GAWiA1bQqnM4GRunnqURmQR8EkPCdNkq5gQJ+HwpY3yt6WtZnKC
VIR/AcHh9aGsSA46x0NinNWSWI1KpCe/9Mlv9P7BMDpTL7R6OBPHW/70OMZ8Uidj
D2HksTEZwgojikD/m4oaYvWXEhp16zn56IR2l6uqYyOIN1i+iOWrrxbdjuWmomc2
44DFkgfszR4bNNRFA10kKKse82Zpyj8jtyLkV0iHGJTaHmBXbX2s8vymwIXOkx9E
ZaryCx2+bYEArIRuJiCzQL6/9jXuwsXxeZpPnHt6EG75vq/K302epxZmn4Wa7xLY
OxwcCUTM51zG0e8Wlt889A7xPtCSOnnK2wIMgchnITf36+rf83lqw8aU4S4yxXfj
ZUVruFEYDjaVwa7I7R0mcPPmVvTf9DYpWDdg5+SLo1mfRwd3RsQsJRVWqZmtwmf1
bXLBaFZKhfbBEU5nZ0tQOtzytzIK0i5j620gpqC43+TF1lisi7XwslI5nmtQODMN
F0dAsmCFUHbHCOu9HJKbJtY0eYsU1Iq1ShwDsj9BnJNmi21uMi6dje9m7JMvcAN/
r1EIY6uZFYAnpgZqKPOQTKQU22UIufatPWSGvggzCh2tNgBwxeLl1aXA1XoUsVay
SRGwBDLlI4ZfvV4tCPx0YxJE01pvVAHtbTnmevzuFw0Pqh6foxfmAT+7hDOAOJ3k
IxZREiVuHE+elGFQ8bBgUpljvs9lgOg+YhftQpVPVl/C+wzEVYymclJ8d/+a74PA
xiqgtUd9NrUN5lYmkGRVxUW3ALlaDcVW67eWus0CDpR0IZcv29yHdTCp1syCKGkp
DlXsxaY4kOLS59OkxBYdkFiC0h0OIXFbVK/PUbT7BZyiF+BCKfic3J5dj5EW1KF/
ibhR+UBFhVXjOJbcyUcFmpsvemd/4PKY27MNcll1SqSJ30uYJTAfyY4+z3gcdbNo
uuy7yjHsxUL3m4lg1NWrdl9mMsVbU4Y0U7VBl+w/R2CBYThbZn0ql6lq14hCd8RB
hepsDcN8SvdcYrBY9hAKzfQjda5/Ef3YdUOcc+kFgL9pN/D1lqAnF3qtTl11sXIs
4uiSl6VuLLzv9Ar3XNMeucvIH7/06L0+MBrfU9Ka36Iqy+gideJmLtHX+4vHKGii
YesRb46Yl5mkT2bCdALVKAV10OnWSmGhictZTI1g7UIy1q/iV0ut4KISdtSANYQc
d96D/Yay4x+jCVLtEPi2gTgDpNK2j2c9yaUI/FqkzKzMNpSeuMHG/a5CiULhwFj1
5OhIW6qyHsqs4Tf0yAh+2BjXQe+rvP8Q7PgIe8ZiyWdkHHEtS+xNOdLxrgiSwtTL
T1mr7nTvCQgHkp1jCv4024RQJ327VoCvgT14qgMSxL49MTlXH+naJKFDvV09+sXv
38bsx+HSkO8vofJRqIxcxHq/vZV/PrhP9Mt2tBaRyvSZX0Zb1tzpH2NWBX9hiKxA
vrWWwWv6BsKN5HXKsi8iv/itE21wSYiIrwEOxSVtZUNqHAK5DBthQSFdddchsdwc
POeQGU9GM3I6oqCXXVP4sS6l584RtBcwV4FjOgCt+l2SOb5sCHsJBSeN2AHm1yNJ
BerjK2BLzoyi/xiu8vMsTsu3Ydm2cK8INiOAP/HXjSZrJE0dNwXqctkqMlxUJK5I
AS4qCFCFhevH95LLjxWTWMGV4LYu0MprOd87ryQYpB9xZIv9APpqd7V3Kk/vZ/Yd
Ft4mz3ienc195oSGZEJoE1IvnmEXqTDTRlrv2rpbz5PQWgG3bgHlmtsYfX3yMFIx
z2VZE/iRIEql18kAAxjbbScBgbYUwTl/IFb/pQgYeOl1Ardd+yNKzf+Tmebtik/g
y3ETmIWCuZzsUBDfqhoLgA5L0Z2aE2mP7idKuPn+tm0m8S5tKx+5Jq8SumMwWSgQ
wElrFd6a8lAaCULYa7JZpRrknWVdssvhGDtW1d//Lr3O5HSDV2g7+CNBolOOhj1k
7xWWpiwjUu2M31rXKBNc/7kVl/j+YIVs2GXGVuVD96R8/nxYtREnOtYBAfzwDXX/
PyzLg70Wnii5cDYcvafvqaMJthlrKxcdFi2IKdQnGz3fhLgRqx2Ny+UWYmM7uPpT
jbPfSztUVUu1v6fTajumBxdOtAQ5Uef3RgK3pgUpg4FPhLb9m7jmgce4BZ/ckhAx
oqw17zCcqHX9tXiGLKZAEHRa2Ud48XTFsGrEGk/FuY8Afo8xqVjbD79dGuBqtaUV
lUloUixJpqexsWR3o6ERRtrO/wpJ8Z8RfGEW/yM9yY/bXjGLPe/EXOC0g5hdem3P
vSKImJPJmH+990Q8fzEAwrm8wmMEca6IslnVo+BDg6HgvOoPvDbdU4KsodXzrb75
hg202cVogeSUM6up/C5AbFV5kXL6GiwNcNawMx/rjjDvLp2tLhIKdFHzUUN003em
mKeqgM404+fQl8YdqDgpwJ1Ngg2P/G6nxd5OuDrbgviBT+VQRyHqRzUMF2mKYPVk
E0HIsAonH19U0E17Ufx1VCWQ93R2vH5QxRaRIzoUvXu3XySohiMsNkAShidEzeIj
ACevZHVg3G84nPKnyBCCw7QBQFQ+WtYFn4xA4hSHuWK9u3YziWjzCx4CID2ug0Vg
QpZM+6TFJCUG9qgACzX5KFAYrBIVHYC+UY/zH7zHxC/k8YD6NqkYWtOaj9EgTChv
SoeIqXsNxLbDReNsnqQ7taLQmEF5KsR+gDE7jnVgebqFgaijYBPH/4XSzw6VH0et
gz+UsRC+kW7nAUi57zoPnlws9zm/Q58TGnPszc+AfjWyHeVNUqYmezzw8Rj4N2sj
aQ/JvX+5BGCqUH+HZX7GirjEOAhI436VclFGp9qk88cfmfDrJufgeugxNfFctA5D
OuwPSBCesx5bvy50O29vKAV85bdfefYoGUu4rv1KjWF/qCK1o/NQFCs2xGDP3bph
KR9siYIphwKSuaxAA1r/h+PaQQnlRycpEDolmM6iNRoLr7iHOFSFwgFhTwBO84bx
LxTyzfcJ36QzPxHhswEXeY5grrvdgkYoe2sn3Ds5O0Vdu6/cEzixAcnNdbv8Th/u
/HXilVHedf7MVMhJObDtWn1NkCRk7phbYaJj1TDZik429CF6ahlgRjRUVz1dDDJN
yoCRBajMoRWDAn7067F3bt94K+v8xOkvLp/X1YPA7wjLwOit7395m6cauSinLci0
nXG7JYd+IOfIf+VTNq0X9mpIT6a0vJysBHrtE+LHiBGzHVOX0OOynxTItcnMKXgA
p7H/D3kmVzBUDQO0OPdjvnkYO3G3g3P/hYjRqnfzfNSal8LP2GpdLBpfo1d+XkIy
p4Kl6Sf1MbiDTaKcu/2M0uVGRYmTKxFUUHtc9L7JdBgFkWFhF7Lqm07EsmLxBd7H
g7SfCeBx0jnLau/4dcrn7gXur5MWkZ2lDlKOabjIRI/0RDqRuX540JJkzl6BD6nW
ujUTNOXvNechwLvHogjsgYEtawBgNQqXACuJTIBt9WXAMEdcHNaY0GGpBcxNG7Ec
sSpJ2Xe7m8gIY3xPKJAvCZcB/NcYuOhd1KUtqacU41t72d4cGg1XJx9jNc70PdBs
SJa5sDQpcB9QNA4xlAy+Zps23O0AKhiJWtrndHlv9Vgc8f0On9O+d6l+uYL+zD+q
cbX++AfJ5oF7NOxEMi/yEfkfmPEiQybDy1Wbx7z3GMxIXwKpmEupueuYX1SrzZP4
A5w0jLGeJ446Q4rhKnzZxvJIhaugy+3k85P4/1TbYL3tnEycoOLK8VgFolANhFdn
t5+a/OsSI7pgrVtrkqqcs9Z7lXeeCmDEocK+0rsJ6164MGboOmW6HXfaGXo5mQiz
nfZC4L47GEBUSMCOz293/GmWHqs5dGqJ/h6H6V36VvyeeEYONZwIVb5xLuXPEYSQ
3x0MguNUiUe3RXzBcB7IBETmDySPlwon/EVAfeXGMGJtJeT69jXkTY1zIEr8t3wi
JTPX2AxVQJQ/KMblt14bPcmq/YeGnVwj/CtMeG9gaAJ2V9gQ0GY/tQ3j43fFp5g0
zV2vfeVT6gQjNy2wRpXBhC/zvHEaUJ6jGStXFcNi6AGvfmKYDmbfjRDj5FTzzAUc
8Ee4Q943gRmChFleBf7jZh57r+QRtYOotr9DGe8WPJv7GFwasVIGkXnKljBFTAKw
4dZssIi+GUk4eUYr0bX8pBBOHSqaveWyV8gTXOL6HUNeOdZjB7jQLqCJIsoS6lV/
GVVmEqCfjTUlZ/g/DmeDGSypYQ+lGLkj/X3BjoCG33VJZc1Xe+9NONFlT3gH+hj8
/Z/mVeSWQ0g4bkI7deONsAGxqIujetZtgqmYHmAA9+lmjvpakjEcTBfNdRsq5/v7
fs9mFY8p7493dV86KwnBZ9JjQhASzCI6xMmkH7m3srKlBJME1xRhGWtuLk+ioV/E
BN9maSNAvxvoCLdEGrhSS3BOHyUOnAoUjUwuaF1bN2QYNTXfRi7ojEdJBzgUFH+4
AOJKWQItZqmtZEnb4sxaBZHpNMXd4z2f8r4K5G3Fu0sArZ9Q4SZ2jsDSV6mfnn2U
ZQz4T5cFCxqNBdpeY4JYzlygoEdNQuSyR/xulKVrbdioxZ4GksGoTm/RmpqTDHmK
rxOZb4+AgEfdsyD8krASJdMnNJyTbqtZm5g2zw7zX7FOb/o7w9RSnlYsc1ErugQc
0NlnXHqICrX+ZGqIWGn9cZZfmtBBAhIR+2MX85EOCjNCrS/1bEIDPcrooZ7KG5Km
83rIpf5dc/Z2BLonw8Nblnk/gTPvGqI5380w4/slKlSY+815oAOP7Gfe+QVNenj/
SmFZvALUt8WzQvRBMhfQ7tk8pJWYTNo3GQbd8AomArNC+tL46a8J4yMCVtgbudP3
LoWz+KifNAcKGoo4sDMPzshOkhnWLMcLdCxBM2G9eHWYstIS6sin3tq2UmRGx+wn
QsA5HbaO3UlBcLNhlpkACWMPczOwTOS4k7xTon5fjc9k/iB3PoXDXZlTT0Vr4NhT
qf02TevNFIUAIvRjGrLQiTkkjuCpU2/mqIPXdMJhnm892YLW1XkJwvCaOoxX3Kc7
C8Zx//UW6RM2eRqpLitTuC4Vzu/dojicLnKSwMS1EpaW1Qyt7h1GDyQ7YVZKr5cs
tQ++xNTSyWfjukg9it8mBFGkdfWRlGBi88ds+sp7pk8zDm8qEz4+SiHegLYQhLSo
10YQEDSS2Rxn5qDdfAS3HhPqy+xLUkjuopQ448meljlft9ILisjCLsSain2NIWx+
TmlrRHwpi3iis3gR4Xr3Drw7nnYRandj0BIE/Cj3gMRVKmS1V1IM//6FVK3dAfLW
PRYL/Fb3R7P2pjvi6IwIHk65bKGAISSj0vNySKyDc0Y2m0oOS85EomLRAZe0hpNw
4P7bRyj+kblIt64Oe3OS3r6+USyRgW8gGjD9FiAmVZcT+wIh9M8t9b2oIzOBza14
uRCIzjxwK9C/f3WIz9sbodPaqUGTORdAqpKoH6t/EkAVNvfaVojbjKGj97EJpPgF
IoJhf4Hm1D9uCBNr3hVDBUaQ3PL16aSYZi29GloiirVdvyZVGJIeptc1e5LCACDu
p7FXCp1tPnm7UPrxDhXznQ0rEYhdf0Y9LBb/s5xUhjKH3fUJPaB9ebGmvW2R+H5Q
+WqfDaKjH2qnO2IpTwqjLK6gemG3GEt1Mu5WGQnxzOByfDZxALlvoTXNNqYhxME2
6fldi4Ef+Ufk+06Zg8PLtFvUuvbuzii4wllfMsHtrKoKNn1NnSIrsBYWLqoTXblz
gkicOURrt1gFoTsMhK4RAd7kjUT1XoJxc0NCIrpvlFCNtg5XxB6D5BWxbz08relY
FWrSOgyLeEqfgWc//5CqceLXjd8WlrdW+4qmnAngVh0A9SbxUwNsFbN7RsCVxI5r
G0Ua1qFZjjv/kvqqjC5XITlMf1monWCBtFJXVD88o5BtC2ybQfidjH1Ic7ZcMsCJ
kUBfJ+0m6eTSuhidYzhaXUMpSnx6tHDtdifN8R8buwFHUGEhqyq+FliDh6iQHIZu
SaYeZv/PmbRX8pY3CPT7tsaPOpXnnEbn6SJV/xRxMTz0bDqT72HHCsYmO7vEYxOs
zxB4UWe5B4bdvn9WFR8EPY4m+eXyl4c+RYQzcBzx3J6uObpkmrT1BJJNjoKXduIN
YYNniDe9DzB+wnYqG1TyGk03DOLBHkyIbHgbat7uowaPQPaxwviSWgHoF13NLhAq
0vCnYsO55ERPVqiSJnCRlkBYLWH8S1sKk4NvoEHRxItSLInvD86/MizeKZyIVz6y
vR2opZ1+pSC8bUTGezWSDY3cjddT0gJmf3NIP1fZow2bToCkxTxzQluWNO9xOqbU
71tdc9+ik+CICKC0rj/EkHHdAGp9NYQeOFbT80OsMpa1AW5jFXZOQZX3nVXzatkm
9PB61lX1FhgbWVZu9frg9Vnf9RnTCHcBWs6XHhrU8bYnqGILeDXBARQwkvXMyTNI
hoBSRWNaP5M0+I9Vyzb+EQ21Beo8btkZIYjk7olgGsT/oJnKWUwYg5C2cOh3ymIz
QHGzBxt36DqtdE6Gv7U0hTTykgvGch45iHNmwWdoVAbSoVt9VvtcK6p1zJyQVThd
j4ilkF5wICOe37tkjk8nXQ64xJBxkaXgQWr9yx400vinNcJGVJyO+pewIY4iLNww
ye47LuU+aAguI/t78W3l4G9W0PhOmHgi8+iauK3kkIj52XuEI22G3fa6yElZbcFc
uvZ6jaucFw8xbJC8nxL9vt7fdszFpXGPZ9pPowtuDedpK328q2IzgKwEF73wbpXr
QHxw2ofti/KvfNA2nc3fAtyqoNbDGWA+d60h58HLFktPrOXh78d0576491L1PxT4
Eozam48ckwApLR5GfaZ/NhEaFM4tBp1EgaCe/INuhaQmL1m4befTJal6FmzI2rMs
3D41dr5tpoIBvDxRWiU0/KtG3kAzXGY2IiUCKRKBd8HC7pYTYPB5zBKnAUJYUINM
QR4+U+3PB/k1xz84jhSZ9tqYKGL+K6293A/nzxfYYdfR1vRP7rKlsxHQQ7H0DV80
XlwbNtkuTJytEy9lfYep9okUIlt284HKG/BUoAta9PB003DYTlz/WBZEhZ7VTFxq
e5gCewTiAv9zUwFklyxEpVW6DQG5rfRROqB1zHArb8aqnfU+QfWuL5m+0WkzBAon
B/hokFeNm99tsmxEnQki/P1IgjYo165U4QJ2czsyGick0ARh18fXi0IfdwTaIxVr
NZqoepMVMHMG6pzZ/KNBy6TpCIgWOds+dQSoQK3pF26blVR8oEZ0Hb/9w91E6Ek9
kZGv59+SrnH99p6cAaJdYDWf+it4pTiLgx/P6UDINvOjqrXuSrRoDsPGZcFnhipA
lIjuHZNdd3yrOAugOFPd2INRhh3O5jiryPUwXmIZabFnwmE09ITdnGB99BIKFLPj
HgA6ioNJUG+oZKeqJti7bPurntLillmReZmVs9BPWZ43dBOSvAh8OOjiWA7D1b28
HUu/eSWmyz7Q9Dfbm5a29K38YTqejBQvAP+9hb5Yk1UYk38Fh5+XxJOZeT46m24m
thvj6Sr0wUVz0BQ2ukWOs6/RcuxSyyaVYf7bcjeojFepIgDaDGKARtBgzTV27ZBr
TwPJ2LPP2UcaxwNb8Ws7mrTjBTkXsbHNTIu5yUlwtD4o+k/ObT4McddKbJiuxPJ6
jnjS4tauIB6yyoPsp7rtILp9JzLXbBNBVNXKuD35YVPTRXKf75YeJQ2M1pSrwKV6
YNCbEX+c2vg1E4lhLlpG1xztdqINMhQJKG90XmvUz8OL50QEQkTcZiaSqPeVjyhP
LPS1LqReWROGoAiD7GRTC7rYzDC1AQivwdM5rGdWmsb4stynpYSz2mTrRE4Rc7jG
ftbThwOPEAGAZKBHfXnl2AeA/uB+gpvyuwW6WQ6IWTlryxgiczOrDx7M3szzjvUY
9jx8AOy0i1Q/aYvNfrQt8rZu9AOQgtTg0JvrlJEmnqBgQBGEKt0i8tGUEqCPJAK6
dF7+5o4KNtzGKs06ohbIP9cYQBrYoLLdgWt7aLO8tVvwdgBqvHXUjvDSrqLpfo8a
qvZjl0bYUn2QeIDzTyR+HgsAFqCuoUU52gdI73lb4xvCdfwO38rt+J3yfpp5G8ij
+wgt/9WZnACn9Un+S57nRFfcTLFlHVPb1d8oJyeal0jVXyv7Ts+TsEeHaV0/2ND9
TNSqA+P71kTrSx/jRWZszVlQPujv+eeMpLqeAb8x7FGbIDuMQjQQT/OYfYSOWVON
nWwwfKVViZacGPR+XUvuxMKNmaOI3+3qvqtFuM0IIvN2HwAOVxjN2ldWmEjhu6L8
kOJmJ0bQ1fwOoZo8ViPL6N5P6HP6JDOIEPmAgKFV+CYAtiFQ1vMd5IthJoID7yTh
naRiNDteooBouCrdaLkiXv8fkigCH7JKYg0sHk8gM3XZhZ2Mn34QR2XPXKUlXsT4
0KADbIQQi8nLcpi7plkaIvzxYdD1tk2WTdql7QBMRMOtbTdwzqGI9+RrOC1AOTjZ
qTLItsqhoTV4+VaTT6gjhfk2hKvPKDP92QaA8QKQrgNTqhS/A+03fT6DfmntYY2S
6Y+JZCyZhKOqBLjOBVypSg49VLxcEqAc+N/CZ7y4/tfJ4ffLiyrn7KpWbA5qG+dz
lfm2Bi/VQP2SYAdOwT8v53xeBfC0Wptmyfd5+Nq5AOQamq7EQu8SwoQ+1QkvzHQ/
H99YoDShyHFd5Fwx/Aehj40/fwyMWtSvAv6tzdCgd8AlZGdKP5LyF4oZ/VyX72h7
4HlFAM3AeDkcAQ9Nkr0y7mmrMCf/G2u2Uoa4776ulGv0EgjaZ3bF1uTuQzh3lv0m
J2J1hHcfAjtneyKy/NyYnDiC+QSXSF2Q9sMZXl3Wv5cs78JzaB7t+9hgKxXTW/ju
8vnu27OpjqyOyXmss+DGbUvRasPXy+3/76q2utQ0VlvGoGLz2WllydvjDkTKOsXr
ks9E85Xih9dz0o+fjwk2dmxqYtdLdVOCF5I6I/lj1GmElE8AdCTRPQJoTPno0euu
koHg/FUeQbgSTbXnsS6C65LBQzNSphSY3Ji9lJ9fetCOJScl6zZBzLu9rWwhFzMd
AXIuUk4WxVBlmlK3IaLRYcJEmvtgvBuf+IC1/GGEdz2wFOQa2TAfgJATPvJbX3Nm
JpFL1PuAHPq3/gzrVSEYA7CwpS3M2ek2d6LDeLsCqRzKcR+C/Wtnc5xfRSE0H3LZ
afrXiGuwbWeobPiJ1d+CT3gGEAvpCsUDxF5vhpC4RfHDUHMY7IXxIq9sZZWjhloJ
0XoVt87tmWhAO3lgcLNrfaNGRISV4l43TlzwVT0eDAkYe7HbJu17gC7takb+Pwat
St+BS92aSBhetCDtNGsN0+cEs51MfzMe+K2hlrXC75nEqPDSVYM1wPd0bUpxOA4Q
Kwk/sLgkS6+SbIow+afwof4JNdnw1AV/UGo+IbhMnAv0EX3VzrHCcJ/MHq5lyI73
TBTgfZMAvArWIN/2xaLHM6/lsYHMkw9iSzPJL8i5HQU3oI40PxxmHhOTbTK4zdOg
WBmSXS0f93dLNnPJsZ+DoC231eF3f/9eO6dUWVI5x33CbkzO1dFHCcjjNYmX88p8
ylWEwPQw/zw7f/bIbGrWtIbdtBbfdGJGbteIkS5cAqeX1iBq82jw6L0BgEjb0+fm
itGhEBcpKf0Eo27iIVIXwjJpJbDLgd27GTuf4dE0D+BRbdYJuar+moVxD1X/jfPE
obujeaFaQ72VJCBo6/+aYnnkyaKtvvxWqj9wF5zowCHW5BbCp8U9CEs0fOtyjohM
QBDdRL/bxRLc8untUwmQqmbE3efc7FuiLERYCpkvNw/95B0aKcHTKrbJjGWZLZNx
xjiijcg6DJZTqPv3tBDmNjUS4ajyAC9Suf2VWlemnirrDiYnaUzgL61Tj8QSE7It
dubv1v0Lli6fXDfyMezWZA0Z1awc+2tdjOHndp6wpRB1E1zbI4QMUG88sjLIK1DV
KpU5+4vUDBYOSmxObwBKefsWY4/KXN3bViWHhOZXIwNdOy9GXIaWgLq837DvRB66
bb1l9C8NM2eI7/v0OOgsCNaU+CEcuyTlGfu1VO2C/zHNsh/hkYOnfPyDwqWsf1QD
5+0qDgAJNYpW0qGtcSFHeASPLv35+jFxDzcvT4FrkGdWtUWwKl7+qFcpWElbgMo7
2HuGFgXZNm0O9LTxdki5UGAPQU6ykort05+ceDwR75IM20TKORK91l349ZBjPIzT
YxzxXvKRFsJy/y4aWZxfCO+0a7tQc5lSmPpZzNZSdEnrL4tBm+8e22W6k/WAIzvn
JbTl7Y0a24rRf80rUo3TRxyM6IvBk+nzj1m3TJROoVuth4GLU9qibkZc+1Apfpjo
hBNjqp3iewHRAGnHBlqyP9WjrkekOoC9S3f8K4V5vyyCXpdBnQaFVVK9Hzw4PRn+
SXOGYkE97JFBidtffGoAFbS3V/z3x/4lBYUugKyRZna6A17D7pWOH33boIsp4V9z
vIzTPae4EPAFBv5LlkFflcDEODfICFb3aTGOyk4Z/qsIX+osFh8d5ii2h5wtSfiH
vQuWilYUoAHb4T2agQCFBRV7IsARTH4ySN3sZJeKBwe0gzFYSGHgr8KDHkRt+2Z2
cumo3HZzKYHTCavj7ZdoMPTYd4umCcY3jCQsx9a/KZ3wCE9vZj/ty9vQUGiq4Fr/
gZMZ2KFMYPqIZmnt19phYm8CZDnlG87W3pZS1GLidfjCEbQH3y7aHHGEFPD+IS1t
OI1cX4yb0oq5V3MSNtvJa8+cgfrLqUvF5Mqn6Dvh8CuUlcPFU+ldrGPC80mZOVDJ
Rv8mcRTn6m0BFntpU9vY31OHn+PE9uwCVejRsYFfCqRUC6kp4sDp+dpPA0Et+5n1
bxi/6q7mzaJBODJwBDeSPOfXuq0vmXATtOVGk6VASO7xJfb0F/N9o8FGMChXkx7j
WXhSAPNaQ69XBHBIHsNbWZCnyrIRa8M9EcPxPyB5fAwtdCKFKKGUn9DNhV6+nXXU
HKZO1xaOjA5lvr6NC40bG1ogYFdPFl8es/4EGmBxwp08cOF67nnNHvPtHqFHsBai
MHY8Yf/YsPsCYd1LX7RFg26PSo4C36F4TdjeYtfgcGHSX4tMdvurMLKoVSvalCEn
3Pb+mNhha7GqnZj3VqfWLDTuijXFTKwyt18I4AGkK7Io6Z6kFwnqQewG7EEgTy77
Llt71av6y9cm/BX4X2txqCkVxZtUKibkDRovdaIkJrM/B0NjVJ02V57EfZ8vBQKl
fG0zxjga8maL002M7JeWFP0/4MzFEeiLm92iarOcElVvN+UWkiDGniVyU3jBgfMN
KqF3SxoGaANSLplKDYCasgW1gqZ1g7ZX/LfWeveDRvB/J+OmjoVOCDz7/Cqsmwl4
fz+PFv+KcxMgEFzl5njZ/4gY5APuRhT/3B0VKw0Ks5ftvWPE6VKvAhBr2gv0vqu4
PfR3n9lFmFWng7P0NtlixiHBdxqXIfxxaAO30MOp/jvVYNqAUJE5CX1i0ZoyIqlv
GHS3etHNzHn7z99aKatd40y2pao4hYcmpMcrgiTvKUN2HOsMMOzoGhA3zDjh+jtd
QHTOBNa56uI1fN3gTOttz2bu2ij2jIg7aDPqKD/ha0fCHHoTvsJ6vtfJ+I967cl7
ySdp6vxKnTiNpEvlsOGgCAKw07xbTUxFG7wA2hua8WSIbWw/+GPlmo0VzDUGQ3kt
wcRg9Vogn/GH0n5Q8xuzbVfv0tZrwBBVS0KQ/qj829oKPgPdRIZlgnk0Z33kacCc
g/6KPouhPHutffDd/LGpUCdZHwNUyVBmONzIhbOVxONFP/XVuKVu8oCuXXuncx/u
GzszysX1RexEF8rZ1XCnMG3ln1owXTjVnVmH7joGMz39JINZ+Xg7dIWMbkPAqmzO
cj40wu0Y0R3M8uuNj0I6nqc06SifFKnY8Gkxaz/i7HOAh/gz34CCtzycYcXMPlGw
py84W3rj66AfswUCvI3aE7scvp9lsFH+JZ86yVRzTc8OWfeIqvLzbD23ZA0/Bkyn
Lpg+NEPDifAP8134T7yfRPwCRAj+spqfH3ILnu0EXigMTUVHWTpnkCBlBNsbI3jE
NR9YUD7VINRapwmlaCGuJ3sJ4rnIYDZo4svgQMl3EdwFrwh2awB7jGj7/1PLFaZ3
PA6ShukD78VfIXsLZ04OOgfqGGNHNqhYqaslSasVhDWhOHFe1ff0kCzp213Iznus
u1+etVDzxidPvEgsvPnjHlw+awYgpIs8SUulWMTGIC5OSpIjUj8snaV2GfdHC9vv
scv63xFZgXANfQLs8xJ58RdXWsWU4PWXau25nWNn0KKJHKskuUXBwr9HdIr6Zgud
JRVtqlPYEZNX7N0iDZgpJDoSJnTmhR6SlJBH4cKt5dxxbPoDkxOKD96/gnYfk99f
EHQV+l0FyW+ZQ3ZbprL76s6dnymhT3y4gXIC3o2+BEkWyJottERQ0Z0c48Z6FsA7
xTJbYBlQdAtj/XyPX6e/oANnl1xVaSlOrTf/UPE5ZaZ6ogFcAce+s/hKvrwfNne9
mQ2SMghfVz3NJqxDr2yr5GuhHqPqO4OjmYwp8rN+RsseFz/uI22bt4ISXufHV4fV
aefiBvDNMmjWzUbGRl09Fo+ZaDwHYYEdWhV3HeGfiHG0rLsnEiOO5naxudE9BHUt
jD+jR6nX6d8JHQlj+2dIhV6uQerd+PNIdj9zwLDThB8xfALO2ami2qx3CyvXXlgb
KhiwL4WavR0tJ6zp9zBWIRG0Q/JxXYRLfJIK98z4723xu7K+p14aF6SvHPUaoElf
L1LkMs3j3wLPz2buuUpanh3QWAfoVaNdgweSXzolGTHMThSV+cm0fIPXPzea4Vrp
t7Gpeh2BIlNDMq7UWkpIcGc5HOTa/jZI9t6FnnvijjyJzp5xl/lK9JislrN7Wv5k
W9HbmWz9qXawTWpqiuoo46WGrMk5ibkSrm5YBWqZgaRB0SjhSXnc0Ql8wh6eO8gx
mkt0aCUR2vzpDRX9qgnVgD5L67+tqmX67skoJlN300h/pU4NuALBAS3/VQt4NHGS
GFL3zJbM+JqL8zpTORQiznt2f/PN/2b0imcRGx1aeend5J8Z76ei0h8YKzkRAVZa
j1ZjayE1fAxpySmcZy5AKJEILqQbI3W2cqWxT2NRRcEUqsJ15VEf44ty4Wc3j74F
oUats+0Wuq1LjPjfUAy5LVpaZIQfGEWfluRn+UvrQgdIRa4hp6nRV6aUf5RXuWtR
75F8H82aT+49uA+xx3jkP35ggBVZTCTEbIJ0FO55UO2KFJO0orVrjjKKMknnbJQg
LgY78nyezQF6mSZglOOxzIg7TAnVy7yI5It52Y63/iyLKFzepubV3ZnRKggdm5Jp
/4n6vXn1Vd760s4BKZbSOJFvXgZlXLMHrcEIwtCX4CbeUl8lKhJPebI137HagYUr
4Ih7T/ySN1xSvwLFOrDQdommFsyZ2nZ77j3QjKq2gdmy9TPqHOco/el4elt2tns8
ynDFTWNzBF1dld0Szc2+C6/CyuAUfL8jajRFfmPrBW0G/mqmvK0pIdDaCJ6ULNhh
HXHjvvKajqUjyheqbkfYxHFxhszbTlb0SqD9rubHqf+e+5ZsNmV6GvU2SAcP96F0
rPEZxrMfFGr0O3L4fcOVUesO4YqF+hnZlM8S6wt93AfjEh9NAd3ZR7dxTGBVOFlG
fwT8lmtT/ituUyK3UfF3taoxeAInz8cYDE6sNuyv9PBcGzKmAO2lSehJkm+jLjvB
ZcpPRUCGav/X0Y3XnRtT476HKjljb/JCCvQB3CIxd5juK38GTMXUcOApXhfJ5dX0
6/11JkxRo+quID5awqF7JdBLV9/OSfPdC/Yk4H392XGOPAk4GWvod3oRf9UNOoSY
PjfZmi5RpMkF30UhAX9+TrOYUWQQ5QAcxl4F66ACmRaixcEEqQiwfSLZV6o4dnzD
RBMKshxEUeUEcHgZxxxP/kZ71vUIkCY4+zGJkIBnWhLsbro7/moGiMIIxxQ6AP/W
a5yS2QBalnwmB1kxUPaeMjido2Xkvrwg1ZKwYjcAAmUW+HFkClPHfIda7bveTA35
Y6Ra8Lia8DH9xXj24iIBQHWTeuKUWEb5pQ+lAeWEL1svxYJp412xuohiIYd2suHU
voK6xdZ2PYK52DSl6ybFPDU5csQZQILfCN7yMdiIEoGHq8+MPvqFQMs0d44dfunt
phmfHjOzVIDYsge2NecxMJK1wqqeTVpC1bB4QG7wJpR4N5s1/mpaiVZLG0sXrAQs
uH6dYcPVXIzs9YZLS6G6lfrqXwSjyTPR1FjUFpPQ4BjaCNo7sWBixXNwG6y5z/vA
M7QT2UgcgbzY+A0ykD73tCFb7z/GiYaxE/TwSWIo2sIaLnHyGmi1ceMq9HchQnzR
AO7aH0dIHrUtJb/NVF5LWc0bLHRrfDBoEXiGYNUWFb1fBrDEAdmV715HYCHo/hGI
13wTfnXWrsglQnq4UzqjqlifG78FKQ1vMXuTQMYtUpkzwsAmqtaQ5GanAzbpz5CS
h5rBXxsJtq0aGA0uwjxMJ5lrRulZmVV0r5HRKzk/DjiXoVzfPijYCktcQ6faDwNu
WGrhDR6XklS3xxamEgdhlv9dkUacpoD1jLFM770S3k/g11gHbzJuAtrwMVdj4Xc+
YDkCHZ976D59GazB21fcYnl080d/PsOZxnRahI8gVuy0xnDB3b4vROUM6ytX3dUj
3dIDUfKeuXS/h+GoUpqy5hHbT7/Qq1S5Xnl947DncStnt+F7tSYK6o31f5PdLNKk
1uUMuqpiniuLKErAuA9knBxiFPd3dMc1EEifF+qyBG05ZOMNog8PQn5XUU7awB+f
bJKoleFeHZtd2t5/3VcIUp3oVpDQdQLuQ1tzNwF1pdfqcC8HvikFEKrIXGBCmcpq
T2xssPVjacHTlrzNENn6GrY+7eFZRiBjZ24slfKWy1eCqO1UUhAbWQ0N+MpGLRUK
NG25hVS213G/bccENluzyjhODX9g3lhvDfYZ7sGYqcUHxh5ySZvVquByhZttp9I4
zg5g006g7CQtGfW/+xnVQfBSgCdkRX++8NQF/r2icbf9/Aus1fYAVC6CbV9+vE9W
jxRaVTEUa9628qf6D9J532+hfVbzN0OHqNUIpJF/j634KG54kRL8dRjFDWJvxxVa
lsMo83iFF6oq/NfHUP5z1i72dDPMieVaTAVYm8uDvGHQRyTs9ifaiU6KOwd+4aBt
E6hs2BATAaVWv3Bzv1pboghhlIMG+HdjCwh+Vz/enyYCq1e04LTTB5MBwzvyfwxy
fr3D1ipjyNJCybugmatNg4/BSxdUJ4dhg9TFljBpyHWUmOi+6hJsCmzyG/azR+Q5
CztwtpXI3gR0KDBt8XGamRF1vSyraEld8QmFQoITsbB5XXG8DuAbQ8DWrrGgAJo3
g093ymUgBd/eyYF7S2XkYcNKwDAHwd7/c466b6KeXk29cSPIhvTGZwAJDnXmX687
eXZk5XGbb3oKKRlsNUZhkCCi/8C+I8G5sDwj6WMy4VWS09izRPL73syWvXkp+FDe
GxCgZdCEq2W5w29CQHAKM1tI8G8aFKi82hELF06MeqnTft2MqFNaOZY2uZp0IfRW
ZvIl2TXeYXr97DAIlqdMso2YdUAVbCJPEGDXthU96WCbzPPC6tJu0A12JkdbdPHl
U2ZnstF2dBgSyfuxBnyDBqUIMtZgF+bjKzVOW0G+k7Pi2WG1X/et4HgPgf9RWoFm
oI993qhQfnoBM/aas9pHeC4XXxg41RlHy9/1IBX3951M8DoI61OabzqcrnKs1iiB
wKRyWMhde5ICdtxM9jY47hMvBaILc9pQZAUSyHDJdH1ApD/fYQBETBBcReHNeo9t
MdIBaMFJIAND+R/hGjuHW4Q/QW12wSGXSXGecZj6ExxkJQZBQ/bfZeY0lKG0RBQo
0CbyJRvYS7wnU6BOIcVc9qKByYYP+4V4XJE34FXykNj5fq4YpI+2IbjCEGjfVDu+
YU8t3L5si0inam30KkNA7ZHN1rZou5lrYhH5qNiEUA/Uk3mP9c0YRsHlnmfQCdUU
EvraXRPbWAIL06n0baY4l4qAcHa8zU+QpwAC20FfJn+3lQqIeLUcxAqKvYAPszxh
il08QnOO8wuO3TYz0RWYrxzEUe+HAHYyJ0c6/ygTcdkmYuJlYWGfxW/sladHCmB1
O9+fvwnH2FNEfMkPvWLqmtVD0wTrPfZumLmMnJ6wr/HVcYutUE40brGQHosDfZfj
3RnEbKM0N2H6faT0qyfcD6Onh3Dy41MPUUmLlBjCJ6Js0bJGmKrUuxxbnJZEEhAB
H5qnPkS1gsPWBXYlTrK3tOFRQgLnDmmVr0cZ1qwWqLMbK/Hiu/t7qADEltIA0wQu
Ppd163kvAEgRLTOx50nJCEclCKcDEbqDBPG6KuL2as9nfJRWup75sSnDgbIYKJ/4
M9Es3dzG7aCNLCvaLXQ/Wd0WP0yCN+WroMhVlSn8YkUQcTsRxQ28hq4bVm8nj9Tp
6rceu7OrCb5e/cGYcoRYf0UTTeR5eqUxb5QMQjX3cXUMozXSfFi0up35kXJ7FK5D
J4wKFN4+NzsDDAtxNxoq6f5M9fpFgqz+68nThpdkBGN4kRhuQ1fesxsKBKdJnzxY
s6oNBpqY5bnWAaxK1QcndMnNfX1Wyy3TSPEgWIHr+gfzHp/g0JDTXe5V9olz1sBc
ceoovnLxpTo0hU9P6VVvyDqBp8uokafMzv9lJnDkyrrxwmjZBczFiQ2Eqf9nCMua
R88Ko3G9bdqUgnmgmNYLWcuBnO9O46ag7PSVeopOkcmLg8r2MdqmDhJGxDar+tcX
xWzYUD9pkXRJvI70sUANtJd/f5yupBpNOn3BSSPSpxt/i3HvkoBiim+d4oXflPSL
U8BGSKV1ZF7OLlYWPrZInRNVDZeUV3JA9DB5B1oCTw18c3V8+ZW8mdwSeQsuKXQZ
wjIzmMvPaFtEDHMu/hSMLKVGwNxwLrr0s+FW93EPFlfxywW8dQ0hcJJw2NVrB4+X
8Cz52rXQpvnzs5jtZQEo9QrKMTqpFeM9mR0c15kGcFAofGksxBNJw6Az/nVi2IX6
VvMe0RdLQNOJ+1vcwO3vZHFGLVi4evFQral7o48JDmBeqQNYzWUxkT/rMggNLgYr
dbZlUAgGpADRXb0Cej7TyWqGlOGiEaUPXfA3czy/RMc5HspmJML0T7fSmIE6rSbz
c9JpdaHT+ln24ML+k0+GCwRnEY1L7Y0LacBbLztpaJR2wkM2Lgh6X1/fP/t2dL9Q
y+lUsuNZsEp41+LUBxsfgoGombPxzCjAaR6yu5Ug/p5P0eZQ1kdwEmeIA19DBqEv
N4jJzbv1c1deDn4+BhpGLAyaJloa+qvZMZflx+dDusjaPDhGOKIX3leyJ3IeqowB
o9vr5fw+6orJmUc06v93+rselDLKUm43PWBUJC18O0Ef8vyuPVI01iRghr4YGT/p
eqYkDCtzr3zs3enPgiBcOjHZePmSm7seNBEglNj5bb2/qFL96+zVXlNB0u04Vjdb
bQqMJX8+3aiX0kg0oyHHdNov0Hdd1ZxN3wyi9pI16Qvueyx0VThvEMgDnM3R8HSG
78674fONOsgXVncB7RghrK+qxx4DVpbXnVuyXeAM4ZRV8WMuiTgjOYhQ6gGD9AI9
UD1NMts1HPese+Kb1eH/CfGAmzAQFy2Xde5NR+vRbScGDDVVgU49nkJGHdHobPtP
kwS2NX+dkBMwtBsNZqBrB7kJphYOxm05O/S9WLfx78EETxLoCkYH5U20RBF3RNS8
LGW6YsQf4QssPoUWrTIkcGYKO0a90Bflq9SzOvaF6v8SIWGCJvoGQEbh5haFfTHo
5wczENAYi+dLR8PM/b8hKqufPGSUE3BoxAvIrOwZj4/jBAiT+VkHO8FDtsZzvmyE
p8bMxo6uazQ+4tJi/4ltMelq5zaqx3tzfr594PZdLkkCKn92GNDsxYWSHDFfw1Ne
R40a+Z2fycdmfEZvVdLfpc+vOdaFjjbo+WcfLr2Mnnh9lXH2KMpb/rHd6eLDhul1
q9/Eb6aySpHdabnbDp2PPvHheysny/yhr3692hGDYikem7vCKalP8VEfgwHlrF/F
GQUZCMhFmeTJisLDPkGcsbFE/nMamRjLfTJVPvXRawV2NC3mWhci2bQnArXQeaDB
EhH8Io9FS/ZzB+wqfoJUy0GBh/cIlP2PEwNR6iD0It+d681BcsQ2PfsmlzveUWDJ
+rFeV4LvwfMemB3vKnx+VsB9udflnV0yuLeNeqHn8VVumg6XRV4LDxr/tBTNBzko
sKPrPlQs7gdYDjtUhgvWLjHp+J/aMrN28tNkhn3oZ3f00MkxVWnpJJ575YGoQwAn
bCf/OvlnzPvyEoN1no+lbc7QUMpPenjN5lORtxrX1X3triKZKz0a9DRMXNpyh4ob
b2vqNVga3N01By6MHFsSn+hd24vgwoKaj0UeIUZDwEcVIzeld4iXDRml57rQ5JRP
SzLp6LIkc5qrr1DOSmKPldFIa6crs0K9w3dbNFcTg8mi58/hfPpPtYVP68PRLh7n
AxLmYMTSA/U3clY71/YCN8etZgceeYoyp0JjyUCdbxJH9v3w9h/uOFrWNjnwkfP0
UKQ56TBy177ez+A5LtGWxUnnJ268IELtm3gSm2Nj5KdQivRC1wZtctsRlZzqO/Zb
Yyu7lA4ioyz/0jf75UI62v93lXbnwAVEUfB9ySi9nXBUYYYkgeVJbfi+GqWtE5OX
0VIUh+exBfgw4D/Twrn6h+7zqTN/w8QhDBH/xTGdpODPMXfSmjfx1rya8tKRHs+R
1oECeQDBwUiV001mCC6JwPsn/SeCEjvv+kdWWyfcteRbBHD2/5xOGY+3VU6Z20EP
cvzP/uPO9whG02zIRBR0YSvMx+MPtIvIP/1A+JVTXJjqUFUj5Zis2TjLZljyIBT2
acD55k5O3sQTJAyzoB7kf1YF+hRt8sutBW2JlRhgL9zDB2PAO4+6QVZ/cLPXeG6S
+HkrI152YEzc3/vg9Z8aUIWoNHL07igaYmd8BncGOvTHManigpqn1Xo6+jMKE+JJ
zibyJVYIq7vVawYe+nH+Y5r8PrvyslytiKt2roDEEQbmY9St5XMvjuvF/qKF12Pf
GEinC4LKKidVfCyXDgYZvGp/l4XYOo0mi1Qk93CA9SNvuUWrW4x2s7q4DOQZYmgc
ujJ1MulL5DEs3e2ZaAK4xao/RrKSrFL7oMEyJsZMD+OjmQ3XkfQCDLEtlnIK00ud
zpmFA4R/qAsTAEnSu90lNhYqx5sN68DurIUsN3ekDekJ1YwRfeD8yWPRPtuEtCwd
DMHdJBDXNneyKfKxcglX+oHQqFsaW/LM5fQKeJ33Hv4d9oqR7kP1RwaeUPkcgNKu
vFeDhETsHCRGR0dip4k6tgdelmS7vFOe4l27Vd+xvojD6y7jOgFMVG/s/u8LQbEg
k7H+Km9gpzlZr3VUou4SflmplH3lDHU+eD4B1aM0dI1ty2Jx9OTkQjgI8TrWH74q
+l4ObFjuM4ipX5jM+xp/dUjnUXTxYQUhN1C6ZCRRHJhe1fm+8pnpu2UyvcWZuij+
miVzdRIfT9W0kK9rvd58WnzE/QF/W/Y5TT6d/OFKs1BzPQB3rgz8I2gFn/MafyQm
yRBKebqebNk6RMYjVYNvzLTaaxXct+pK3efpRMzGSa/vGlOQJMK8mT6SE4lc5H6N
LTFQiIClx+nxV2Ywz3tVBsMVyO7lhmpoB3t32gdfXRFZ+1K4RXpbrVvaT0eEq+Jp
PgNnfZeRXn0JpC4oDswC8e+twdTYvMhTZulOwJVlC6qYRRofQGOmJt7dGLJsVWba
W1P9D8BjgclNlHhoNTE+NK9hzoPaSqvce1lCSnnSp+kvhobPApQYQRv0Q4TmhJCB
2CTebzGIMtcI2SrOrlt0fXucIzI3GkYeGCU1el6l8NAgrn4zZ02CFPk+xqOLydop
Dg47/eKsEREEPhBWcSuZLgcer9q1U8L9lj9LxcXIgM8XHOljqKVpW0fYzwcBT3Kc
FKJMFpf7d/IA7bIgh6QTC3KoaJh1IeFL24H12WMLSzmmWDTwIZK6NQvIUDpQ4gMm
KFTCnuGbMe9wcBB+4IT++W4o/2KOnkKeZcdwXTJaJ418EqMGmAV+dFCAawW7i5To
ZjR3U68YhwosuVFVw/x/dUjFeT/6XR/bFOI0IaRzfZ6wqkL41ltfzIm0qz4p3b8M
80PbXE2j91TCycSnAJrJV/fkbzSe4gYg5LXqqwAw7tBNgzPi1Y7zzOGKIVf/sx6p
XEP6Px/KCVleSxwXNneAp9A4PA8RM+Mv3fPVPTYx4hYkTfal5NaZvOWIyLchkv//
0JLjOkjnDGpZOGPhcYVkbI3h79BcKRa24sqvPbvXqTDoJ7G+Ei0Opzmm0+5iKqNI
vvYYUkJHpZkKrq4DHMFVpPrAohWW9FirleYlrvTbI3+Kx6hiTgq1rFLUkmkxs+lR
ZRmq6p3elLfbg4fvg9w7GRzYtJs34wkpbGVYJQgEioH26YumfJxYfzVRT6ccMyYK
jsfa/4Rxos1zsVis3jkJ0bhkzCIPFpW1pAhsZB3zVBiW9d7DjDLsFQOEMqkVWu+j
LEOtCnF7e17Ry/BnAdtfiDAHGersvFWE7omk8T3d9zIEYwSbxicy3gYVHLLhytmm
xcMFc4ljWa6fsXRcW3HUzSCsRoLcBWOxRds0pn07KX0zaMi3AXfz4U5iUz4wCwwB
nM5mdOOUezAPHS9kbso6eldNSmgYcwRXQxhpSHBDjj2QQRj915PkmB3gHAK7MJUR
+RMlhr/DA96nVpsDGr9Z9T4+mBLYbZrnqQlkXUQVeTVTFdOX001fYb+Z8/DFfced
I7UAFGtEk2xGYUYq/McmxtTuqykZK0fLVagFr58sfCUJGfPK2AWm0bv96X6YtEbU
Gc6c90hovcg0e62GpEKLlZgVHhmDGCVr1deHTCMdlvGkTm+Iq6NAKv/wjOdGgRHw
XVJDRV52by95OQb9WGzE8/Flpl8nCBSWPsQksGTsrlY6VryWaBQ/t/YPzG6bJ9MJ
2iID0FQiI1XfH/W4pjVcfxjvR5vw5zUwv0brOeFggKykGuB/MwGSb4aE5xK4MNrq
f7Fw4ZfxrOj3lveI3ojAco1N8RlDhuY7vRLEULbYJRd4t6H9oS59BjmuNlBc/m9s
3zTtnQdWPaoV8kuDEfTYXWiwxszulCMos+yKnui0xYp/VvB7bUOEtpBINJJnxASQ
ayygJnCkyUbol2jm9foARsHs4FkDQnek6bNWOUQvxm8d3s4jS9NzLkEkw5qvDsRd
+gHdr+NcB2Z2qYRIc0RXQyhSdhZ6rzayriqE67WKxGMgVVy5zBEesDT6oGhV1c6d
9ypdTu6zoebWTMQvtaKqZs6bWPTkXregcwOaqhqZa2znpT8PL+Zht253peJzK7C2
FXhz4jPl5Aj1vrNnAl5gSwAxkASkN4+bL/FAEUrNx0tZvIb435uZOn7AW4teiqQv
GXU6qQI69VHOhNANWSX3OwPp2W9itGXmlGItCwwE+ZIETYGWyz7Nx0YGeWMRrdym
bnFbq62L2BaLPE/kpLo13wuXSSkpmIe0zk4Cx4KPm9Q4BwqBp+C9EGrhBEQvh5ZE
8Q70+9HYxDYvV7mMsTJlld3sQYMSdYRk2c7YsqbEh4kggU9yPgNymw6ZOxj3xUOi
yFbb2ACmz/wHUPutLpSMCwHJTWV4AzyKM8GFUgOZn3hPukizYPNaRV4emIiu3oAu
y/GvgD278CxFB5eVY2QU00A0kZvojDmrjkLaHoyBwJXb0aYD4bwkdD2/6Lw7604l
CMXByLNyELP58fhmZwQmCCDqUe+GBKg0z+lZR7kcCLyn1Zl1gcv5VPxl9VGWTmkC
+enfYUQowKxoUoVZd3qtzNlyg6uDoqxqiXh468seeQikftdVWBJwZXN1xk0YJ4Sh
bfNOqjv/b30n6TyUoLtiVNErgD0dkzFOKBKEBETRrIiubQ4afzKoGVuzzVkx0ueA
MJuAzvyBkeeA6M7OiiU+waOzIXSEPeqpPFocFA7eIygFHjtv2Q8K22ODqvNNI7LJ
tTjn4ke7HA5UXlxXjKSJhzU7zLjlOV0HigZhe0qLCdAjqZsFkTRkK0FQMp+CU5vd
cC6rYvSNgYxHG/u3c/egDkyGUb9EaEO95Y135quEAKKaQCsGO7ceuXJ/fXHTkv1S
R90p+uLd9ZX+S47GPAs5+5nT1EAkzOk7Ez6YMB5SDdRkP/raF7NSLHkuCIHag2Pi
C/1DEo0E6uf20SnWEmuUbQcKsvBPRMbb0VFI1vViSbNvTCR4xOQyeKm8pzJPyoEZ
qakIvAhkGXbpdI+mhXTuZEg90r0V4N4+TDlpIM94bunihlQN6tYoDVL5v0fFSSPL
u1vPBK30KLR++qls4cZUQiHhKRK+41oaXaQjBOUXOFWYB6Bj21Chh6b1ZKXeTV4Y
FcoLefBMJztgxO3jUlTbbl8mnhEYn8f049t+P1eQkjgbum5c3tH2VofOZwa3q4AO
P0qUKQIQhhfnlB95C8hKREeFwD9rhYQa64fbk/6brkvlXoZ2Bs8E83VEupCyDDYo
Ou8YwPNH9zyYn++/OR/q57hv+N24edG2SCeF7udGBVuSihs7S7jvew2P/11rfa8w
Q/ZCqw1nBK5R2KQBwANA//wmQrJ0vms8GHveVjLSQuII2w/ZxZ42fUmp9MyGKsCt
cFZkXrhcDp+vcCAny5ZphvJHxPY9xt8F15NxWWSEGYotY+M2sZtDMpJ+Arlu3fWx
bF6UGsRe15e7fxl5LUN4ZOcGpYf2CXsJmec7GOAvRfBhRlaifI6Dcqhb+tbyQY5m
esBZSuwYReXVq4loLhPksFk9pRCyWxui/htnDs2i6N3G1+MMwr6dLcXXY1QJaS5G
Rv7CrDUdJrhRPkK1Br+QsdZfGIBVWLetXfMVobSWGxFs8lCj9XxByE6I/AexVGs2
YhkSDftFq+9Mn+51dqPFD9+0MpA1lcJVLVoQwnpirVbJmfeiWiOBEYgmwgBEO8Ea
XlMq3BLc9RwFB7A6t4WVpdCxCEzH/XiUi5OutpgNItxizD5GXSDpGHeRmpawGGPO
Z63zLMjyIrmGwF7PeSDwFPFrn448O+D2mJNKg+AdAfTLpzrjM22UWq1AvyQkpISe
9JSd7IpxbINbvgWHiD/Jgyw3cGgTvT4xn171HsXNXG5Gro6auyo/CGZXxAtzkXjG
ZMO0CYbUHlAW9fotIKctLBGYqkSxERikYkG8gz/QSzGx9XpwLqCPNaPW8gAl5tLA
hLb8ES6kRROJjj3koGJVKoOobbxOt8pszBz5cCmKtAn/NXCPE6LJ8mhWCIN/hnp3
sEdUVHzjfnRmeXk6yy08kcxrBBcLk9gu31bFqIIYJ2ijjyqguNhDXgsJrlcyviuv
qPiIk78r0HB+1jiWJ+kALtxXlTonRKEIAz0gW3cI1ixSBLfgCb5mquCipAVBklaw
ic9GdCCzwm0kniZQ5GqJ3O9hSCIUHe4cJKegmnOn/LGxq0DiCD+w3IoxvaR0qTnB
ijmITfOWG3+zCEe0teM9uU3UfbiBNTaS3w7jnvxhJ/KPghlf3Cgp1OmY/tv16JV3
H0wcnoIqwJn12b39CdJuaex3EBjU0Ax9/5peTN43oLRJNsXlkFdYV2ODDEb3N8rX
8LxB1Qfh/yqsfVBn8sYz/nGIVgHd5ADjpTz0zkBR5kmGnqWs8QFXwmo60XPaker+
hgH4kP4ZIFTiXu3Y3Tu3z4P+AqUQ8/0VemgW95iPxUQgs857bEIaz5/53v3o7qIo
SmsgiT5YDEilp2nWp7z3EyAO5UXQvQ/GDb7MC325MUK4F4dKNtNr5KIF/YStEDYF
rszPiI1AxnJMcMiyroaVIbk+F9TnJRaaAUD51j+neaGFpiC6JbM5GFGu23Zdp6j1
glez4kQ/WzWJhan86SS6qX6a6mxUsOaNhyPIJ1dllR+Wz6cwspv9nalDtmYQ9fjR
rgCxgLQsnb7R6sjAu9qeON+A8eZ4a8frzYTwYp7wTqJyRexIEQCIvqoRvpBzVIfL
fWPZHRr74KXJ4ecNTuh4FY/2WTvasndJX56oyl+eKDzGctfEsPiLnwmMZpAAfER6
ioJsJHQ6ZKR+/fNC6bx6gEAMWzp0xQ9ky+llJ2x1jBYl05zNib4h9EvPgw6MKW7i
N6P/f9VBHGOoT3Xn7cjFVO0/YF81sTAVkadNH6EokqHpT/YaVGCGThzDehgFU2fe
m2whRC+qZlZSptr+exuvdVygWi4tqwXxfXOKNxjD59a8+HqexTXoD8+OlLHd1Etx
vpBp7NpaYKki9jW4T1mtAR4xASdfWU45cI42ch6TODVWr71Fc9fZnb59BoczusR6
0JPNkgaV2ggbduH378eiJ7GHvgiIPQZu+8hzybN4x4u05Yc5jY3mapDCLmPlMRws
Y4kCfzJ5MPtSgAOP4rsIxynxRuHWXVF4kV1o5gzFp/tEiPSEyB9nbzg4k16Yc29T
JV4/aYiTXYcgbsswDg8kc1pWJhw0ENTXZ5liaeu/eXpT3imgg0mctLY+7ejKCvZd
6pQ2eTftlm5eviNwUuaAJuQM+SFbsjkh97bzJkA6qpwI8Uzvo7CQsa7IRIf+RT7i
AyMhIZgMNZy6tF9ryaZL9dxE3V/lFgayQUQAf/5i9e/0oMndWY5bnWkXiE2C6nY6
EbtBz2lTqbwjeTGD0YRLpjMPEfMx+FayRjyq9O24yIpI7aUmCtKZpTIJXyXEp0X1
KNq35KxlU6W1OvN8+afVjzmSITBuENx/KpjE9pg8n3oiDRhTlo/X+9xuQ4XQw433
gWasY+CBDLEceJZRYHA9M9SJ7aTqcn9z7E+WGFH4sIVmED+1MZkLcXYSwHSrkFPl
dDPSqBmiDxpqzfLSsMvKDpXLehnH14asRPsM98ym0WTcFvqwWb0WscGcoFxuKh01
Gvhl1MXDMOzpqJykI+KSgT/yMmyWYqSxWSXG7na5z7K8GyyRABVTOnZlAfuKkzM8
rVJx8xnQ9cG2U9P2NE2Y+8A2bL4MGItgj3z3LvxI5otMv49/E7x778f1uKSCHeZ9
2R+bGeVi4hdc5pFFyBKK7JJDaJrgWuS2aypdTOHnDPA1XmqMVMNFXsdgc6Uk0Ovq
2IbkdRNI1gmDVpVfEtsK1s5+54NYjOaUGGbQ46a2LACgHloz5vBargwXSr5izK7c
2iROGbLYmn80+F2x0ryUcsPv4L729S4WblMTflX0h52QB8EmxgHvEm40WjMtq6Fm
CARPPPE6ryTbsmzIpWQ4pTAt8WhvwrZbI3Tt3FB9UUeoBqw9I5IAGu54uoiCx7C7
DsOGJQVHYYxWEj84e5yWxBLmJSSJgI1agQQ//1vIgZ43QDVn4Yg4Y5/02KE/wF7G
dUPhiEUGR0XWNpjAQZE80ozEonXUNicrGjYH/TjN3jU1zh/H3PamYwEq1phUoaad
F1okiiJBBz2nFyoE+5pdy069EDUCh4n/jRfRIJ+8d/sHpETYzChg26J7EHXzlXIx
DiQ1uZouAGXwagspPjAM+aWxBvj31N5vrmqMTj+B+ly0/YxmbL2RlNeebCRrfVh2
YThXVkZdtp/GhVaK4LmbzT+PhrwqhF6lpt7sR8S3iSF5t4OvI9jjhV/0lniZoFLI
ZAV5716VWxI7+6AivHZDshC6DwK4ZoF0HEHDxA0CR/EdWIxSkWPr8uf5Kbjz6kcf
1QdXxEorw73IwarC61kQfZIfhk42jh4U0uR/EJK5MCuGPde89A2XelkPkKS1veV9
Z60MYZAPzklM5IE7+Qy7b+IIdllkQIUMlUSi/1ecvpeA3yfZk3Iic9dVnskAdlpe
jtWF47SMtpvPYv714IMUWtZhVrqCzpzMAtVJN604UsweSFceFnhDQmLzBKecUol7
yN1vF94G96PNfNQ5E6NYon4/+nG99cLl37UxaqdK5pLYZJPwmY0FTYGxaFyrQlBE
o8H5rNYw2KVUFbOdC6b66vy8sfaklXom4lUvQXadItDJvmLsSyeUSuf0puY8J4Hg
dhXYq3NNFsIvLybDXnUH64+LY6Z5rIyWjVghEDPrpQ5w62zSlVkjVAF0E18NM/Wb
hDJ2JJNzk6o3bmn+6jXgO+ltXhr4E1ib/hJMLZ1oy2aXE1+42cr1+Zou4PseQj/S
rKu8/usP7ZQOfMxzPnw/yEPuVordCEF//7LnN9rVg8jwKRZN+RH+VW6LZCphzMao
RkDaZ0J95ihUcU5xNuiy7wFbiPf9JCe78aDRc+D5IZplPJbDfP5XHdIJhZ3zw60R
535ptdVz7tqoeA2lNRd2y0rER5wmKmeOa7WPODCmmY6iH1pU3spZERFg0Q+NG3Yw
WCj0ICs6G9wuh5XST7X1xjjQke2oQDwAEzvnW9v22UAIwETA09Wy+d0bK3ipTNGb
9URDoNn9UzzRCPoiqiNRuojnrAO7a8TKN2QyOgYNSPtAXqxCw+gU5HRuYEzK1ZbY
YFA6/jTH/XvC5M+DR0zO4MoxoueRrf2EZmUHXhmJJ2b446KzCerJUF3VV5Z57tEM
vDzVNSBUtqpROqR7HlHJodwmQ2/zG1P37pa2Th/gIXUujLFPKDvuf3QXxjA4nu+J
EoDQwZdSP2O5T9oj7dscQxtRO+Hvo3fKDOfRm7VwwPNWdnYhOaYhO7zWlR3M24mR
srAj4pHQnpmcWNSiAhVaWAaaqJ/inusGsu0Ya8rlsLhHrC5ZYBMBCzRLhzujYoCb
cCsuEt96GZS2NNNzDTluRijO46dlfb1PefPFnvcuV5NBvSuuROrmirOEYNf2ydmP
bd8OFzxHE2DB5BQeiqC/+ID7JXdIwfOKFEH5NCs73Xxvid7B22IFZpPQ+Pu8VRIp
StYu0Qo3DNqBLH3fTA01yIoSI19/CLepqdxAcIvnW061qaHJCd/a2xjUJYkTgi06
UlkPMigsF++aFigyvgi6uBH/0g1HHTUhgTOv6soeEs9UAOUOFsNQyFQh6DJHOur2
lb6tltekjERPGdAZBk/iO4LuzYHS/imwzajBiHtUcINyNZiGFSdXrDUr9kC0oXtW
p6ftv2PPTVL0TlNWPpWsytF4oTvFWhGpnZSDX62JWgheUxb/vfW16qcSG7Mz4uJl
uXUapqBZQ6+CZxmjq4oCPnBWp1GyoD8UILWHo2xyn4fO4Jnf2wDNQjAq16tG8Wr1
ezgeTdkdJJCd5VsDf5bIWgjQz1rHpJUKXJyGlb9laxsVtlaDxU/A85W/kLGXgVnV
bY3JYf839lXOtdTL8Wiajla3MF2evoeEQ8WkXNE3Wt4XPWjhlRbW1jyy2xpzz0Ju
CFseDEDbS+PvvYFQs8kuXaKKACI6id/jJ2BMouY4p00T0k89nBerDn0NRdwm17jo
k0Dq0ot8kLZXbdqSKCysQTHMgX3V2vDhcNs1zrbv1v7r5QnvVl6tn9sY2nlkZzeY
d4o7Ru479U93vHWQz+4XXz+1jdMJ8lwlxWnDCm08EAsfrsh2oeAF2fXX4HQGtbfZ
TMX+Mo8N1aQg5SBwk84nYuNBIptBDwJUrUOBlp1qLqJY2NLyiUJlpT4bYaOjhWBr
AtJEmuWv9CRBHPxqqOiDCcBV5XYBdkGuMpofUfo0c68azQeb2mOGFUHTmLIkH1fY
ZeB5QRJ9mDg6ze0csKqEdV6ZQoI906Bvaj0h4OMvY6Ra7cDP7uvxR+ypp3SBU57k
dHKuIn1RV9u9LbwzM2Y6yxmnskyKW+zwIHjokDhkZ3JEGzfXj0wNk/Bdi2a7K/OP
SgvmhTsaWrrHfC+UhSadKDWETkbj7Zvg1vPUV+mX0hKj4E9mz8+1bL7s7SF8C1k8
Mq3DgZ21oarjSJ5GDG6ofazdTj1qub47XsmxH+OKwSZUe6UMY0+uFxiXHRZGPbsv
0JjrQHyERsYM8Kn7rnWAEgLPsK1i+6pN9lwok1i0EN7EoMW99yuCyiccclla1/1p
7NiCHz+Hs4TG0ScJUGK522tBPvydva57Uy4Sm/E8oKv3MNajUp8W/EiTeE1fO70F
ShLD1ApcUSBlZ2VyWl0etHr+wmlmIoDw4wmuTMRNrcnYRmmBq/KUR4Dk3VHDkZ5m
/yKHCHbKABraivthd9QPnUEsUHfLZYKv2hHRSGcHdoJL3AVGVgXBe/cW/Knrfao1
emrsJvrgbnTfvEC1Qwyv+26MEUXWdY1rg5IGa5s3ksNX5XWAopZG//1yHENZsshE
QnGk/SaZ3P6xQjXBsFaAEjJQjfikrEAlJQMUi5aL6eHXaEa4DYJVpQB6toVY7xIi
5xqAi1OWMc3eG9D7j6CtSe4XgKMRET7lBu0+4boHABT3H08A1+eKJZssF/veu3S+
pdZOgXa81SKFUxpJPwAj7sq9Rr5kZXhy4a5xoq4l9IZwFe6N8TvLFks9CSH6YBUT
1K/bZUo5dc+fPOysigGVXYHhUWVU7SIlpPRNEWy/oHy7m6Z9zDjmv4AaPAxC6V6Y
F0BsrOywZI8wQbj85owT8kgtncD5sMzec9PkdW3SzCflPfNXMdKB/W7trpwu1Nko
gfTy2p+KC7AThKAFS3ZO1OxzzHIPj+skgdUMnDybV/46+AQ0wpAsXRhMe5eJdcgn
xvnekpK6FYiIcqEeMDPlKd5KIw07+Q82+sdJQzJeV2umBD67VV2MmcGYGCOZfMsm
Z7KszeRZ7F9HUB2kKeRmJOaYpDQMqGIURcx1yCN7KlKj9HyPvqtl9nWTlC4OW5ua
PSauUEF1j/vwz7COZupIsi8IPOeDxcZEt/dAWLz1C2LmuNVClYgA/9EUbBs+mijQ
RwM4USQYfoT8ZqEzFs7d/ven9jotkkrOHA4ydZiEaR4G6uh8auzWE5ruMnZ7gJM3
OcPvZ7eBg/RqUS2h4FaXPkgJyyI3UVTiI7TBiXlnBBTxMm7DnvB2RNzJCk9BImjX
Z1wg4/Subk2OkekxgG4dbBOKGKVqnBt56ePWAhgnQyMWEEYXXOmp1v9EhGNpItBT
MhlYeROTtgYASfIpWAFpcTZjzng/kyOtlcLOtV+k8pB0DnjZYclaUM6K/uGIHLpI
rby3AUVpdIJMMABOBCHBSl9pb2IIN0pLcnEyx+/31UDi/dx/OTV7NhHpfvIazPvU
Fi5DJ1Oga5iaZZJsLBvTfNq5jwXFYNIdGLrVveFe6eFJwrLQ+7u4kUkQqqUr6IqQ
iCyW+AhUnJzJxH0/KAWP0FfhuW0GKQtzm31yVFo57N1COvnh9qhVR/xMmEtP3d2U
EG0LmhFSUbgUJuxKbMqj1YXvN1V1+il/jgNmPvuaoVmbicPuQj5o1aowBEnxvial
XC/yhvt9I3961/a06oOYmn9CVEp+rNU2zy5KylHkGuQwrHDXvF69cQZi77YHE0+s
ecUqUtAApIswUuzOSXRpQ+oyvw7y3ruEZuCApsRG6+AC0dOLfJ7QbQMHXk745OG9
be0VdsLf72uJvtpFGFED3WbvtfOi8w/30AI7j0XNHx5o5yOUw/IzG6nXAwE8r4JQ
LEtuC7YyOmq0iELDvg9ET/nHv4+BzmQmHSEf378Hola7YxkOEWutO24jqXMoypy7
rlSwQNT0HLD+a2HoLsndcCxM62LaGUplYedZJrUUXbdFD4S5a8OsgTOsom8dWvde
woCo8/UoP+xPhA09b2jGB9NsxRWNn8cXjWJXvbD4049iHfvjIIVNpjmDuv4/vi2y
JouspdLdDX2GqML/wlOcpmJmXfIX94bCHrjIdnryWZvPwszmEARIpXWHsFRVhcVB
anvQlB317rpaMcl+nUOClzLqZ3J2FxO/UYyQ1btQRaqre2cs0WNx2JRSM4R6yisX
bObzgnYFW8A1uHFAVugDAnYuIqBZ2jCPtsPolmqDMlyOUAI97tDX9vaoZevPR6Me
h4Xza/pwzosZWf+ySfQZItLkntm9D2giaHj5slh+RwPN26tA0f32wAViY8SeY7Ds
F3drQGsOoxsN1RjHaJeMhap0+qlVFq+xx8DC/NbemJP8Ea58oBfdJdvGNiNPSTXA
U55lHAeVc+HOjJTXBTdvl2+TJnJVxvymMEPh9M8pN41ck+mBb5d6+JHvjxgsoyvN
XrLJMSjRQIzeJfErHrvs5mHmHZPJqNRr4cNzwp4ZqhSTnSYhnUzNd7p3WdPMvGs+
kW74v4dR2vj6tldBSa52XhizmWeKlUYSihZQT3HezftqY9GV6hOcrurUopYcdjnI
NiMGKcjkKuoafa+dm0HFahWnmD3PVX2MMhUK9F5MMUGeh0bfFKohgb8RfHBOXoVe
b5JP5I3tfSnJGcrEo13dso5FVGsFEndOcByeCcToExHLX8tVDQI12uG6o+1KRmtQ
W+Q+84+yuqt7qxsim9qsqOO6HGq6CvNFHZcldC6IStvGsPXGgGvOE/FzcIw4FfJh
uie46OC9fzAxjbH0Ao2/F8jun0UiD3OlkieYSqnUyQKeJ+fdHMAiMxUrIdOTmx0k
zyCBQbobcHMhqG5iksB4mMm0/a8z7aWoBFGRXOZdW5P5E+JKg1Ufrd6o+XKYjNR3
SxADNCAKB98od94SCujJZv5vcz2IzQBXjqKLESiC15M3Sdj9V6zn68bh2kub28VL
0tfYgq6CZu9lNCTHn5Qz3X4wCEcfmRXO9nA8OL3YBXltbn5R3LPWtjtWrF+2p82h
aiqkNB5CLx8EZsp7RQbjQgPvB92emSkcl/7c0c7ZllmayERox3anz3lBGG4TbTIZ
iaxS1C2DHoG3pJv6LDFVvJwZyXFLjC8BifxtCFTBZFjngcaJ/ZQkkk78NIMYfEqG
5DgDpw3VX+by/Ld4D8Y6wqz/MPkG+PelkPnDcibfeHmZKfxFaJtQE+QXYmG0QhuA
poAfL+qDXmDMI0ZTQZSNJIbwJ2uE1CgEPJ5iJdxBjToSOsnF3Zw28KONjsicJFBS
UPrJ3FTSmVNa95jbGqWiZRdpu8W9KoV3Yhi826DhqherC2tdNYz8gFxuK4njnE5+
2VkNaS4Rdughaf1T3bZJyuFg65dlR/9tl6wthhHmraVFqp2QOj33Q9+YWd0Hi2AY
E7B9Wn2WBc6ykN4LRZUwX36UbqbBlcht4QIOi5qJtIJChPMqbx2mGulOfyyngCH9
/bgoPiYjvztbbVaomollwrSGTgIx5aDGkUWkHKBKTLo04Nk72PkZSTdKGWgs1/zX
YolT82xdK9WX3fqwwvbkdj/G1wsUvEm43YUqgwuEAH6Jl/Sqg9Ne0j+hrqMqdhGp
fScobHfd1x+Ayuz2lHHhRoLiWB20VrVTCc5Iy/IwzBeVId8HPnI0MMFWM4YNVVXD
cZitja587S+dU9BE2BPZ+k4xGMb7SYFJbIveiru44XNwPh7oOStvmpWGWGruQNDA
mJSFzr+4fDjzvt+iFp1kWxsmlGFB7aAiSp6MlhjWycV3zdxNUrVfYzV73Yhw1HHw
pnFO6ZuSO2mgWbaGUyBRw4EjmUm6ArjA13XeebvM+XyBcgN9iDjdHJFvAsuGfXyt
NvKSjkiZU7+upBFRjeA9x+A13d9MABBl2y9WByuobsIKHr3ccTPRKt47ubSbM4JJ
HJv9bJ4Pxt0ny+Vs0eZKfRcxJX6kAqFXpIFKXJWLMRSdURVsttTuqqbvKLBHHJiP
8RqVywi9o2RQBjJIXfFbq19q8As+CziYTFfTqJkOJxwNT5uDbfsky9mcg1v4fOpN
a7k3/MXXu9nKKs15qVTreYKzYVPxV0P19JQQcc8zcX87xjzShoiZo0K86zSY6Een
jhPj3PBEf5XzymsptxMsUxzXdMV+A1RJs03+l5p/RnycfyCblFODusUeWF6Tonct
ayV+TiIr1QPwS/by2Q7+j5gRBwiBYHrqxycffYRIAAJNJS1KN5s9qk8BpNjyVINm
HoCAzfDEngt9l+zPzLgO7REenA9MTjYm/nW9DOHwQ8q+ZwLi/pPXuKDnSdYJhlLP
EjXNuR7kqyOQCILORAJB1QSTEG2HKPPE8KPeZfkhKswmMoU2MPBl6eAEgfRWuL+4
7G66KhIKmegWk8vLsLz6X2M0L/RPot05lk6K/8VFfCbMrhte6bxza+K09VoMa+oM
/2AjXGYwDllj0h/XQ+srdXEixmIpffZ7WW7keNXz8QPkSt8ncQgrZT+yooFPftPm
YOJj1B6R/nnc5Z9hyOXogGfc+RMm0zZ7NYw0gj98bqMTLaCESOFTS4ax6xXwkN7p
fmPGlpoYRXFXfpUVR7qjVTpa9RjJi73kscXfC2WSm25Ny8KDZlGWaJShSlLh1Dkg
UQIt9vTxVf4k1tV21JnylOoqKrzYJFsGb0akUp0Ohu7vanYzUbQ6ZaVotYAGTDn8
+iYX90+mAxvFcm99m+UzILnOXeaESBrjJJ8hPRJCWC7wVqeJDDz52WonPw1Pl6Tg
yTCR3+ZCQ43TINfLSbLEARybBOa1NUzNIJMpptvPrcibOP/JYhT4yUDrhaHEdIqz
YFK3SPwx7zoQNTcOSKTBaIyekIkg1SOfRc5RGIwhbHAVwy1/NFns7s14miuoEuRd
TovlY5EgQWMAMaZg4+nwtr7McWDYr1Czq2tNWrQ6SbfWBibwG0dFxXihrngBivDW
1xDakxoBGguRVP0l285niyCpnOr6UGwHRKI2CqL/JPxPvkHWAn0yv6uhwb4+gLnt
SvDxSTWAvvZJ01ofuwqPJQ0FvbgiQElrGF5oEkIQ9qsgH5wlnyNOCZ8yif+0GiNh
1Z53Yh6NljBlVIapqtfa8LTRdCRc0iW7uhTVHHItfZqufWOnFUYlMEe+MJWzCgtM
25Bnptc24+1XLPddDrXDHf1KNzGbbkIiXa5hlOsjpFS2Hoj6NpwGbgBte5XJShfL
8C0Lo0vhRS+Kz4X39BMH7qGOYRz9BoeRcDZP65Yh73o8fys0Blu67sCbNPDCYB1J
/gSyAVEFpp+KfM0nLIeGAkmUI8ICvaDlqvSncq7dLVZW+KjYT3EMHtc0oWdo9KOO
BRAX0Mx0j4w17251tI2OE7pmYSfnemzhJsTJg6XkZeydbN6tmCOr2Z7jS+ktA//N
ZyHHO8aXG2+Xu/ELJZsSLi/DG+UJ3lk5lqi3V4H/MDJqQb+QCf2PT6pzU93hGqPV
7uuQstsMVHNbuvl+822Amrve9q2MbG49nh7cElAtXhBUSJSghAvyuBcuIoilvOF4
mh+PkyQ7gGkDq8NDKT0rmMre7YqGpVdfbJ+BA7AV0JQwvEJrDuMF831QiUwITTds
n547jEF1HxgyQ+j2dAOp2WYzCoJXNSvogTtPY0gY9A9Mx4xOFuCB8RlZ7mSmdIRf
WohnpkRECjHdgcJlQRpXWT33NIEp8CtZ/oo8jgjxi5PDDqd+UNhrNDTlunHnHWfG
WC2U0YD81/900SL5I+eIOFymszXTARJWIslOouS1QNi70JwJIWGSmvRIlWWIxQQD
h/u5C/fLrsyf3iM1EQwgM4odYgqQ8maooG9cW2S7khHWzNGejDePz00LMhScnGMF
D8I/9f8SRJZg1syG5ZQb72AoezoN/2+EixUJq1YvZGRFobYVPtlBHRJkQWNqSLdr
iXn5SgUBgwJjI7XRJXUa0NKpuYgYKrApFtFZZDevBxk7yC6VgIMjcSzLuH7sualO
ImKkec+oUNrBixcKhlCkGUyPcw81DyGAujQGIiwf50g8mCFvDKsIaS/GJvcv/0Fd
tGmr4ewXVp8cFtHsOvLzm6fs7lz+coOMeGwRuMlMKXRfdAcuwFwHYxCWohZFLsJD
0vMm3VrMziubW9zYGb+Q8WpkUXfttH23RSCMDq/DwHdookYL4Qkl5TfW6DtLm5UP
x6n21aIpQmKcYUtc76Jxa5tb2vI/dpTbbplU8eoJ51/UAPCidlXyhM995QoV51ef
WiwtLga40JIEXZQGAZwGM0iIhLk/PCWtaVQm3ntChsaYBkHvW2nstD98YFDnXIWu
+1WRaO/QUUjwafqMWPDoX/DsIc61ZOdkDkbX2udkhkx7ZNgKawbbmm5uKeGzvsEq
k660fYE/2NukxLWkqhShmT5SdkILS55pq2AsQY5h/pJuC+dYWanD0vnXZ8nzdT21
fK5H4xH1pIfx96zWL31Gq/b22bn8RHEAeKk0bkbUs4GFLtYXVRapKFOioBlNq2yO
/pyZwQaX1mZCrG/h9O8D3YYxts3YHCy65h7jJxMNN4jvTgwPxRU4QOLFUwPWC3FL
fRt6UMZ2KpWz8u3NaWda2IyBSlWiCi2sztgcgbV7GoV90Z6PCPot2gQQzuVUFINy
v1JVnIU1RnrWe+lDVJX22Up/MV1QqMNNsIKBBlwnpCe/pTC8SoHuaidsTnZmIXTe
p6H8JAxT0gIVE8aSHbWSAmx6nnEp3UdM0TQnb75zJsa15Pl1hxV6Q2vVAmof+unJ
Ub01Zdp+USTsnAAogLpPjfsJhBwYX7Buiq0kMfzMzxhST2QZQ62SQmqMOvYOtCil
4lRth6sU0DOjy+VrTVCiv375fzPLIpcy9tNCWa5locLHvMXI2tdgsC5RXEkG9eVD
gXbZyH6BuhUYIvgv0t5x3suId4sVMdFD3Gek8xqvUuLuANuuvY5NJX6uTqG7b99I
MVzTIfnHMFHZtCS5SRG2mGqgcfSYDDBPhiiKhjlEN58SPMtoJCczOX+MUOptPIs6
eXvVvIiyZz8b+rIDb7DMUPd4tiVU+IENh+Yrl/Frh6kth7pRZnBimcK2q8iCTQVd
yGTmV7H/uV1HmUqcxuQyDL5gycIg7obdtPzuhlg3sN0LDULlXxccC0KKlLSHTxUu
EHP4dg6KSJRFp8lSuKiMHw8AE+YTbDvq13btPi0K7k2842s1Lpa12w2Bt0ony5ia
MiCN5Pd5lDlR951UXLybHFkqB8rHCOmkIikBiQt9Og6BbMyiJccjwV84hsJqJQFa
L0kN4UbYD2h+NkmXZweedG60rxEEbG/lc+E6HQKi/zhGmLrNsox0XPZF/T/phN3H
pr3M+ctL5/iXDPjTZXLUozFUs/hCIRBih/jSXhymVIYtiGlGilIhhCV5huKa+rLC
pJKjXCp9/nlVOtL9HmPoip5azwsO+7IuQcEgeszBFMcR/UCe0uMpkeVBiCVYb6d0
KZEX8Bxc+VdZ0glbv3oeomyosuNjdAEBG8L8ysbTTo2c8Gyqnx9mdqtVJLIa0xDb
zuSAHs8bzDMtobN0z+LBa6HHc7u3ANyF71I/f+vWxp9MbUaoaqalMEiX3j41FseO
ZzbYzr8tEUHBbRaQUKj5wNNmS7+4CtSqF0UsLmHponYH+VjIJNI1jw3mBrIB4UM2
Q4AIrOEe3xypqLwmlTSADgkGoaX7kSS7HIYN8w7M4HGVqwxIe1tGxE6WoMsST/eP
cNVQcS2HKp8HYn0441Ypk3CpdicudATAhKz5WCRlzZA7yx1UXXGD/8DFGljK/+MN
Ty/m+UAFOCMav+KsNUxWUuAY2SAXAv676HhCiCF+VaFatH2gS6xFpK36r7H6t5E4
gk4NH7Ez0QH7BoZsjF366gN+MPb74Z5DkcvD5nSfqUFaHytvkGUy11/qDG93qe6g
x6LJOtsb7S6ua/7m4TvC0VMC7/k8U0dSdQvVuBgSRig8WUbDCjA+P10SQsVsFxF6
3iTo06o3YwOdguc+JPtVpih0vpIAsCbuZrXPDeYYG0wu7Bp0Evxw78eZ/BfX0QWK
R/MW2iePhAltjCfT+YD+CxtDgrnXa0TGr1cppQWlbRdx+4+ikg2+2r0aPNTUkwud
pO8rjoULQRbW7nrJhqnZc/VfUiqmCe0E1Lx3DnaLh89HrkHzXDPrEConFh+ze18x
fQRW96jxr4yo01e8eYWPQolG+1GheRtPOTV9ZWOUR5dPcNasxFhYm+Js5gz8cFaK
Me+7Bw8nq/DXzUrRVvIJpfoJvstBGzBtQws6uAOpCa/7M4WCE4T2EL5KDHyQF2pl
uKuywAd/qI0V0XdcXS1bAnUg11fV4Sf99w8uP+EF9YUdjlk9CzLwv78DEQF+nrkL
nboSmZBaZSCWc0Ipi+3VPUHnp9nmYceuiIixuxTK5yY03EW9WHIEdICnPuocKqB4
UwPFmmvuR+Wg5J+ItRD2zCLhpdev7dwnNeBe5IXmmCWJ9EgW8m3iH4R14avUmlUj
x2jtTaJG0ExYkgNbAsWA0lf/erz9PDT+cgugYsj+QrUeJrm97FQmNVKoYGC6wLzT
bUb8mU7dWtJedtza29y8cHa5O3emctGjr3TdURWImg3LAt4Ol9UC7DHrNkXc1Ahb
Fq5fDqOmphnokkJf/o0bGuaPBOabQR7mH2jHmHzZ/vWIgV9qbJbbE7Le1E82ywCk
M5ryB8DwiU5cSUSM1YU1SGOVmRxiWd2HfJpcWaPXrDQ=
`protect END_PROTECTED
