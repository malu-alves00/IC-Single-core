`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xHEfmMfFnSXPqjMTvA9+QKIUGRugrA+QOH9Rs7HggD5AKMNY0pJcMis8OKF3HRC4
dxYacZuGfYTjtnpYKhDyT9A0MoiGDz5whrXidAwxAi2i4eahGdGLPvMIVKmcHLcz
l4yuSGY7JQc9MvEkbw3F5C9p1+ZbUMZheLAjc5k1/1fvYMmebjKttryeAj6wt8iP
1S5qTu8HtldPCR7ILhdWKR4JFhP7f3CuFPdrJ3I1IyjkgVbPDx9JMl48RehCjelD
XzNEDtc2isp9TUKYcMgsAjm2YXCzoyIvQJ9PvUDEUkaMLHjqkd82gJ9Yh43iC5aP
rQuWRaWdiC3A4OUwQSNldKh3fOHpV/HLNX8kkGcXiWHjsxOY2uMQlO+kbC6V7Ezb
Q88S+zPQYqICubHLKuwKmHWV1FPUgdQ5S7VgMzdw8X9lAO2rTVbYs376+Lc6TMWM
7KkNMbbZtNrTEau/3+VNEiIUycDx6Pqx5bftVV0RqtQx9IVujS0QSnfObQ9DgZ8Y
8vBuOgAq+EBpjAKPvoRpESEeCL/IaD63LG1XApH6InOc8UlE1GPjkMQr/rLjRuo7
XWsR9VhjezESTswaeXomE84CsZnr5YMTNTmjdH+n7h0QGYS9C3/hVgdnJl50nDi4
9CAfPcTIkqtpRqxDaNBTngCud6k1VAh5Qiglt+akZjrt0JZ+Vlee1176V/Vg8fzN
S/4NKAxWayhHjgLfpcdbpb0BSUEeXTYQvheS6zLlm+SoJrWjjGp/Wsds3DKwbbVY
jMBLAQIzEx3G0XdElVu12Ly0AV+xJo5GilCEvs6hZOL97T2P2bHyfQ9AXM1XFE+Z
LHbzy1/liR84UgXvmX09ZMV5oTRbJkAWqZACkzvJRNdZ283e4PXEgFYghbDHuizf
zXLmF3CJ6Ie4T9KhDjaDzR5UhFLS+CuxMXmir1e099L0SkEB7q4eGXnvIKP3ukTZ
TEaC+88yF7pDOVELH916jt70ib0gzNEdi1Xy0oxTp3PQDbZwv6dVE7I7IElx5sXw
mQzu4CgyQzD6VLNVsvx9CmBkcpyL3jmZ0NNfsisiGZUE25Ct1HGsCMxs9pkHI6cj
9RdVf4HnYDM7us0dZdiBrSQsWf1hHXF5875Sved8ReSebv9fuRqEg5wjzEA4Tmjg
6/Noifzcunm5yiiEinENDYS6VupKaNrRJxGLDM2KHo+fCj107/DrXfw8b76iZ5od
vCpO9QN0w17gMwsLnFbA3FEsXwpER61Uo8KYm6IdD47xkIHaDhXaRfUFg0LmMUQ6
cEGVpQe2/Crt6GME25ETZHoTmDAmJPzcR4zVT7B4ICV3mxPGIuvWUZ5LfgZn5sNc
d084ILwwFzIMHRF5/TR2x3Om/4qak38fDxZ56kguDk4Q5kWkEjFItg55RnkU2yfc
xPX32Mwzga6psxruBeGuwDOxshCUM1g18Gs8gKKYfNWH1+Uzre7YJbCxGHw/WBHd
LxQSD/Wf/DkSPYPvkYRSV5V6psM9CuxRYZtWLxwNr+DKhzaroLGyGfw/6K+cePHT
TVecuk3Yj0DXAcJ/4DwASrHnwiPXvlKyA/Tt6BUlPbhvbv2snEE7I1X5I8Ime3XP
W+3NMLXvS1h+C9yJb77/4uN0vTRq6O2qf4H0VDRA81e0BmneWjb08WxyMOBjrqgr
YZ3Pzew9IacX1qXLxYCA7Om80xjN4v2Z80XMOcuvT4RHe6OEaAXvsXl8LvpTwPKB
GBDsNpdlIWLyT6qxL0ksmcbT1gZS7pZK29ohRuP0TsrM6F1tIoZMEIbkYWu7/BSR
NmWOlbikp57iqSdBw7FKQZiALr2GfkgiSBMgipeq2FuGuX6ITeMi1+V272a+cdi4
FTnBP7pZ4PEPimp0aR+Tg2vir3gBYiC5Q4Sfvlug+vLbDLbODlhVwAtUb0Sh/dnC
9oJb3A+aXEo4Lq6kNYiiw2JM1X3tQrdHR2Qb/oLcwraZ+4mxqobkruk4BRR3fTxH
f+L9/H6Hv6zmlYtazsafiJKagpuJ3WFGSDb43lWwBkhKMjFHqJF3oce8WCAD8ztC
SaUNO2ZxO/QV8l0USy1p743mhSSXsOPOlZ0n7A/KrogkRvpgKar4JeE0tq2Xzd6N
ZiMbLwUEZAdcP/p30CxZwn15MOL7NrfLTdu+s0Uz5KVSRrPcqIHOIYhsLSBXXQWk
UPKUTTOtxN0WIHNGqK6WhVvI149Hl6awrsy7qDDs4+sqjYOs1ba829n6l9NO3oMc
65GhtrmOcpMB99w3LFt0W6F6Ldet374Pw/ebyj7OaRAPOmfrIJi9Dt02RPgz8nKr
C1wFIrJOM86PCTcB3evmzIJrrigBd/FJLA26/j4Oj3Q0zQK3h8jDyS3+bNnOhnxt
UYapSr6PpYIDtm9SylfUIH4ukHBYh7qQGTTzc9URNTuJTqAoWGLqIvdyheyfE8k+
IkgsuNziWjL6dOifrivo5Vi3Sq/JkLe3NjzxPt3SxASKXzwFbU8NV3J+21U1f7XF
dR0zXR9TJ5x+wv50SWXKuR/WPi0/Jrtxd/C3jRlRm4LO3w4GCF6+vsOeYIT+8Q1j
JwfKxyEQ+n56ZjkTdKnSUdxCzTVPx0aUqlvYhw/8ufWr+msQZ3wAUF0BnM8eXkZI
1lGzBmM/1+5LVTrII1OIn8ffDSEHD1LF7lSQCvJaye+tqa67OpenbNbw01A5+0qT
gLxDOptp858Td+zgkHDeRZIsEgRLGAEEG12UAgtjIToQ1qS8k43sldXJrVFs6toO
paDtzRcQDE0JEMJDEBKB8w4i5MPlFgqFOnZb//BAbNMRJn4BfU0MG7/dgRL4YRLF
cw6Z3p2YdKqFdtdW6sv86cIrNec1tISyszr+dGcs2Dh8P95A39A+SHCzq4kcR816
LCECeZ13CRKccReqLxriQmGYKMDZWb7JWWkCakPXrcCMg3OsmVtDgd4hxtI+X05v
3f+FXQ8ROrGYjXoIomhd6x7ZxzFw55MakGDwH8OJDgCzv7gMI/ZHlqW09yGc1ePR
piywZgIr2Tc+F4PjyV4rbMcaSMDGhdROwkYbzL6qWeB98RQG+KuFB7HGgJanLpkc
mDRf+5mEgji6GtDY0RuhaPYyQO81olylrsOiMa4teqAhwpe/AbUkx7OnFaJrp/Xn
R5W5DgLbyn6OI0MYkFqJ72A7p7sGvdvAUuom582qkgB69tKEmZNoChQs0xQzcF4Z
GzniodxlDGlOVHQI+iFLpMlz3Nxfqd8+/E7lflluhmDGKUY52lkjfna1Jow9DqX7
QomUheHOAhC/Z5jJimGDVISTQ1USqUekbQSFQOucBBp62QwpIVE0sNaeW9mDXwjW
skNrlAA/w0o6Ts94Dp/FCkexfKkRdRHCbS6nIFiGSxgqA8TKwBrinCIzEwDbTMlR
mT8+BIhuAQCHsRcZH2ZMBD48orxnSFbDOKjtOlZmWO6dE7mmCZHCICGfg8gNfO2S
LCqqWlWqdUZpBa1XsfZb8N9PL8i3qFpobEE9zzR4W/MrWqq4c3ocakiYfboLg4qj
skQRtvYRwT+jw9YoObEt/Tep6sd2N0sFPhMzqBQpbULNbDkvmKyc7nZvd8hKlgh9
SR3Aouw8ud9K//wKeiR+86bXpcLpWKK7kryYbdyJE6wSqbucV0SMltiN+VBjIuSb
peZcF+Nt0y54GQOrP71wSfhB6LC7vi0lB49Xl6miZtR0fUwEcuoqIAs9S6dJzt+Y
I0SLtQ+7jC2o8i980PGLVsnVXgEkSGNmnwTUKS2Inu95CkK7YujJQSbHKnmJ1BmY
sG58PYZq1aeddBKECfSWu83OVOZs46Mqztv+Pu9E2l6BnwuYmnBIB/8QfDd+AwUm
Pa2yBzfPu1An314yNTf4+B+1n6brh51OPq1xxHYEAQcfls/Z7kdy1ZpYZ3fi3+IY
mlj0nebH6ZMPiyUVbLDtt4GS7mIWrhLlAsMN6gG49Cg71YGASCLsofndxuASqXBc
42c4pwNpX/oB8UoD4QmfsPGTMW+v9/K/9sJrxrjjgqUSNNgKHflw2iMKpWKOPTJ1
EDKh/eCPscKhuPyxb9Z8NdLCimO3LtjkmJNWjDACDwSPWCT+BFmeFKG0Kt3B210d
`protect END_PROTECTED
