`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1g9LZjRgSsEwrZBc+EFXjUd6ZrVAUqYZqI1Tl5ag3Nu/yP4ZHwla+6rvJ1tnGh0f
wFWSigHxUgZvkGLPiWijlmMQcakLHkssMVfhz658oFrCTBeGGHRtGlOZj7TLoPkB
qS16NcSwR3YRxiHG8D8MMG1SM0k1Z/myroaT1PanUeCDdct8cwaS2azJdcZQyD4p
bLogzK7d3y2luEsA/YFtnObGnP4gCm2FsetWmql3Kno/SFMAbPX7X6JwJIFfcgX3
lhdL5htc0YyEZF+AsytKAx8cgmtWQc6p/CGPrvs9APpT3tuxPWOHHE04l36MY8pa
SW6Ptuw1uOQKknNDecvmhWWxhlwWA6pk3H2RFCeO/qpBMOBw1mrmRdaJiLWvCoYH
+gXkBx43T8tH+MLbloMFVMe1PbggR827epZx0skfis+czYqrdygDe3GzI5zjig6N
RQttJO8nT/wh1Q5FmryUgtm46ted8e5775+oBsFsgy4=
`protect END_PROTECTED
