`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3LUuWcBmjMP0zPq/ujixA+nixv5uilGHGao0hZfAHVcY1vGfhzX5NVK5G/GoS6xw
4/FZs9yaGNFBxeBRvR0osnaJR/+//AqdtKH70pYaZNdp1tqW72UMstqxbSTLOwYZ
+Uy6YDTrkEAGkPlkQc5sJXQZ6RmAN8RUS4/7j3+K+jnSn+ou4tAO5BXbMwqQPGxi
zZrGaKNOa3rJrDoWnikCe+mw/AD9BzbYmRfHtg1o0oyLC7Z9Op5PxN6fJO7COfVO
0zfXyqrwipqzxJRjOOuQC7Rnlv+TPhQCVt4Zgg6dmc1C/q6qzbT/XcuQYKwqDxbd
+2sWlQ+gvZMMv4tQamlUx1Zi9/ZZTVWfSk/yYm8kwHUuQN5uvSTp8NveLcHN+POt
Vh5gMdjb+mLhfp9ZzuweCcdsJcDC20re+QNCXIl0zwbNu9jn/C3d+D9i3vsdg2IU
pC5xyZIOKRLtNC9qYEhSIOep5Usr94Baj7B3GA2yFvucAcFDxIn3e8gERltv9nn0
gnbfiI/1pKMUac10919bfkuCHXgoH06dD4Um2FF9rj52SpsR0aYdF195FaSYeNf1
FjmxVSdrekkDBahky34mfndHaQuaXQtUJ2tng8PjCJSzfUqobC0vBgdpivhcaAiH
3+mWOVA09/z7ZjcNkCIfu16Z+tdHCeJfV/i0xJlPp/3AO/XXrXZcM5WwUD933r2/
ROEJTJnKKb3m3qJe+nCIgaxKz6VAIE7egiscnps7qjPSmMnnBWE2oMSkrVhNpfv+
wlGam8vvPTbkmnZLje1kBeole785P8Aydd3+J5KC6SZw25aU2rOpGW3jKW4ed6r/
Ji1BLKNvJvCGC5j+k9x0gDvIVDO6zGJcA3WvnI0wHBFKlbUKC71Lrs2qGzX4U9tv
kU8d1pm0TYV62keOlJQS14gF8bG0R78ja3A2Ho32zIpoDgYYsnOg1D5huVmEer/4
onpTn/yXjoqqeWYXW13gpUMHZUTp7+MDGhRrz6LwNqCwHiDWcz+c2XTvXZu0L9JA
0xUqtmKE945AYbYt0ku6uI9ouAWmygQyIPFZaTJqL4ibIxLH2v01zGhrbcOsP2xn
NlKVJ4OuYpbsD9DhIhz2a14laiHCoGQgbg0OyBGQXuUeWdjbOqGrBwvildGLXLXt
YbtfhCoG1Ac2l4N6GkpSRc0E8mDV4nITreMzGjwrFO5nTRkJeJ/g3otb94q+tM6d
bYJre+8bY8+AuGb5Y2AZjjPUlSyEeA0Bg/P2Of938iAYYXYWHPzVqxvpDKtNct91
oH6YvuqlWzgBzdez4mPDzxJefhGIzUl+4dK7MWgWS1ewkVtICgU55iNeuKD7w0o/
7O29KtKnnWKpQj5TzzwtkrSKKlifXW27pbqUgZThXXeT+hsVK15ob25M+6UVwVkZ
dvMZ5RnP2+1vx0Kfhx1qB2HfrrKd5PLYjQZme1f9Uh2BCOKSY1GZlPkzJy+zNh5/
7w5h9dpzLGVpwKG5aDg5zMNSorinBp5S4vatpslSs712AnoK/rUO8+bNVPQMedTY
TCWl2hlsYo+K+0K1/aUmLXbzquZGqoC9jXiUk3J5I9tEizT3Q2lee/MvEBra/aWQ
AihTzQsVR4sSxipuuR4jgmFcJIclZKkQvpg1moPbUPw=
`protect END_PROTECTED
