`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/u2YHbXDnsIh6QQJ8a1KMqm4wQQtl181yabA41qJP9mm5pQcxzF2+NO/Uh9b4499
sLRUXpQeE3GDBRS3g137FHpEjAQUXWh+2y7TqAVE/8Jl/sRwpuT2ctmlLv9NBLyJ
+zIGB/B6bGIxIKYwfn/5iD7UUgjj5GDs8MXKGW1BOuroRkq+FS9ZfZzYXvxTT9rg
P2kbhyFYKDBB9ga7f9/3qMuCvk5R1MFNd6reSmYrOkL8TcDaC5VAzbetc2TxHrAV
iPpXV8uZoeuSMK6gs+NbYWZmQa2pOQMktmL0yC8EkbhRfUw1xwbcxJV3BZcPgiN0
9nGL7dTvnr+rf1Mhd0Phj1iSltRI/wx5GoovdUnJOPJz76jAV5knHViP+GVKhrcd
V9+gX9F9siMUOg3BgnS7XNNFq4/nT4H87N7iF57P/oH0nqz5VAcXzsH8BsOjKKWu
N/5+MV6igJ5a8jEEqUsbG/NJf3iXSwtVS2qvVTuAUqvPuPyUt5lffhGguMg1x0CY
WsOO/PrPYlLCPWsO49gAjEtrkPd2LOcUB/md7mV8vCb8ouE63Hvff0ivpGja01f5
qnTPh8YMWjmuoo1oWUfY2FCsIarixFFpGR3+kZ5O8kIgEeaicvxfwGV76rC54QsF
cqMpZAQJmL45HLxhz4IAsXvyImQ575JkmoVSmwgm4eQyANvGz4Zzf3jGitzAO1nU
5Mk1iGlJzS00y6FAnJqhLmh6fhxjiewnv5Xe/jKMYaGeGbW1NbksIKgLe39IXtRb
yfNlw6DJV1tZLQEEpDUAT7UirqvAKtBn+Xwt4/RwYQjUM8VHwPODZi57Mduy6PNg
uJkeVaqY17+HxvUuOD5J43QKC0C1eysaMFGiQ1F/c8ZiJo8kSWlwdN6JAqiMZLIF
6T/tFkeavuPa86SyI/yauRSkMtGV9IhLV/5DJnbHKX727oALUEtGfjfBe/NDeGxi
lJTMWUN9tPRs4tlJ8vobc16us1Vst9anriJuybHD4FqKJnGzESXwgpXZqwJexc4Z
bkveJ0wpU5afNg8q9HveBMIHkx+5ZwtmsuKocmQb+T0DvqDHKO5Gid7phYd0OrTo
kB4FaRZQacpcLexZ8qEVA6BpoOTxXVIpqpHTywCAloXrVaAJUsBT85F0ky1gQmEJ
j6DxyQI9qa5ELovSlFRSsz5BoEeO3Kt2tx5A6KexI+iJ9//ctS49lGESbiVVAZBM
b0GVfZXZUj+j7y2fyVMBV2VqnfR30q5woRYj9Fn7i2SoEiSu0yZG5WkGXoMAgJUH
rkzS2Dq0EG+m4KfvfwjSqCwpHHokP8Y2TzGMN8SOjF73F5IoilZkjj3Z9PYHwPsb
nGqP05LMlShmiIQXa6AOmkIneNlNPzONxUCcec6gbE8BaGMK8F61PcSjXzIrCs/T
ZZ5mC22A/fvD/KhDZ5I/EDiH+LPttHx8GSWViHM/NeDeGLeyIkEq5vSDRBWc82wa
im7eXd46hr7TqnoY6R90OQYXVqUetpdvrOxssb09pQEzfkaFYyClna0Gde5/Ck3E
uWcSAghv2w7kNfcrH+zVCGt6vRdSF7pcEqKVjNz13eBvf1+6Sc8Up+u/3U/2KtI+
C3fAZLv5TjgBqGRT0jLDDQDeJkoMAyuo2sGyq5HhOS5xwEQWohVTKtncwmBSbRvv
pnwUw6RSFWHn4E6Mx7xG2udQGVgHyNu0uRzjeSsHj0B/OAxB6Fay09FydG69mQzY
2ymEU24ENzDP2GEVa0ztNSbCt7koe0PgUy13CgQpOt5ihj46sVe6plu1sonVdN01
rBdNSmXxFxo4YDfCHtErnEr8kqW7i8Xtogs+sh8blJPsnEQXOiFPrvpvac3L4CtW
HVIEcb8fP0mEIHWldQHEkFMnisveEFK9xiIkjRAsG8mEZxC5Da3MuUMtE+K7/Bor
f87T3qdWXi+1dj6cz+UKIVIspFhZsGZYiIzTQmjrGLkx1VPqpZsbPma2Cit9QYLH
sxofSDb3siD3UtMxbfNl23JOQZdesxtSnBZ2aNHYECiwMLBT87Bl+8B2HmD2YXLM
eJj6PZJpoDzGJWUAuhr9eQXA0ue9jmUPINMEPnBOT5L57RVjX/OfWkpAOGvanJK7
ZjfpS8EYLcRrnZJGk0UGyrZlkimH6hcJlu7xAv75VeE/HpIhxphyeXb8KGupuqQe
cIvJwTXdk7hmj22aL3wOloB69KyzkJwjJFZ/GnJy/rNDVFJJRrY37AnxlUqidxv+
zlbG15pv12SIH9PLiftkKR7XLTRCBdxsGIqu1AzhPi72i90EwCJgql06PQH3yGym
P1zSG4PUloc6CHfagQO4PHsIfAWwY4X1fDRtQSJU5Lubyzn4Zbo+K28NLfY1iVcB
tXmqRyHNV3Dn5sI6qH6XEQ5d8g4+lBlo8q4XLV6qnKSTCymkKqtR0woiqAR56E/s
ukuOr8tZMq5DKOj2OPGZkRB+uzE/r3Z7HPqWYK9XTappObilQ4q2JxUIVPzozBcI
ELzEpaKsFAb3SFTdRtFEg0/M295IUOC09uHaPb325ch8Gn9BWSK6bGIrU8KUG5qK
Gfi+Ts3nkKwkhopqoOc4RAFjkAow1KcHtvyg6jhmnGyxSKqXchhe9usTZwOPnVvW
8Nu2ncL4KVBEyKoLVv+dMcIfzL2rDNf5HJtB5BoGm/QzEf8ewgDic25Q2PWk8cQW
G5UV9HJ+NHIRwAvctp596W/2SkJhk3WrqA/QkKeHDk4HAb/BpFyQBreFP5JMPG6i
wqEAbIV0/rxGan5tI+Fkv0VnMKFnqp65pXhB7tqL6Cl6dV2BQOnB+nQYEoTpqgsX
aIXaUJhVqIKQk5KWllDb2mW6qmFYMpu1hh+/Ou6RTCQBB3ZnXMg9NAfOXm5F9AUB
i0yyhmGICQV/FsOcptDatqELsjwoTcMhi/3imxI6wNlq3bPby0kZ4cF3gpYgnh+U
+sPnEAA+nGhYuoaQI1fa7HH8qftFbdsbRlJ7Cq4nuWIj1h1GHCusawbpHRNawmLr
yYG16lp85yR71LHBWaVqI4kykrBpijbOFLQ93kquPiMj3ryErYnWXARPokbQ0YF+
g8GHhYhlqDVa0d29K77cTaYujqtMLbquW3ostjNwG5oyXiRwL1o8p/Yn2DmISXso
xRasgng82bX0EQl/u6SzuM7MBoKUFMe9+K7nIOS6HfpkWUK3xrxGs9Hz/G+vMCp7
yxThG4MphynwLe2il49K24R5UtL1yG89dW/w+ImxFlUGhuf0XZn9OxnHcd7qgSBK
WPLOZs+qExFteUEWnujJPQpsvgLagoMrw1M6BfLLpkXLlc4ks0G9PXxQKFuyvN1Q
PcV7NWBrDWgVF0pMzdQ2YM7S7certeJ/r81jAGemx6Rh6rFBZM/Bwckyrsoa/+ey
vb6UfdikR+hBcd5scAlRq2q7gE8zf3b+O9bd+CUmGWksZ9F3J/8u/M5clP1mG2yh
BpOzraSVbbPDeo8MeCJDAJLx9M9n/4xuPGcsuOyYFKq0r5gedCaDVFYtdcSFCNJO
`protect END_PROTECTED
