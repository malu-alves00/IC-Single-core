`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tC8lN0nQ75fs9ZJo7zIpKcm4HdPVkFsDKAXQqOFvKzbZY/kpSRa2Qg2wxZzUyGcw
IGRYUt3gS1ryO1Z9W8LgYitLZtm6dbraEcvcRXzmHd0cGV9dxD9Ay42IOWY/Cpe1
OmcQsBmoRhg3PQPwT7rEFJ9qIXpX0Cf/DVlF9/+e0ugm+rM5rQW+8uY2ziDNpMxn
lrLfiqnedPadGkTTzibd3GoOX4+SxahIF4loOeABwL5/P+bjFgiVeHyKxGsvGosw
wTuVD4wcRkhivIXvy2877vE3sMkb57wJ6sZGuGgq2pUUpF5cUC38UCKEgQPNCNie
XwKHEF0LoU808P2+vJdMt0Uj7/tHkc/iDf7qWElYxXPvqGNwXlVxyWYty2aqCEgQ
necFtZK5zoFF/Kh2q9jNdZ7W/clqeBVcAZDapMIDQJH0j6aS7DvgNTN8A3irfLQs
DGjwPvTrcdw9sR57XW3gvYFRj0Q5zNrJVp7JMpE6ajQBH3cU02+rJhUFr2fYsLWZ
nHyxSyMM5Ns5Fun64ofJY8qIg/Z+38fsQOWLRgszPM/CndNb7XK9FsWSMCca9nZW
KNQAG9TNm0azKkmhIs68nuFD2WJ2EiIS0CmqqcSkQPvg+n2voz4fRjyCr+1fqQC1
dcaOPT0ZNN56jT6rV/Wcbsa6PjDuC3jjzvi+aZ6aNnJUYmWozWYhPeQzq1uEf3X7
35EM0a815f7xEuEzMGjemDJQW2l70uUNaxuOu5qSuKdkrm+S22mRMipCA7m4Y0/l
MHvfYzb0p2tH9PU12/6649NUfM7JbfL5MMw3kGd7O1S+uWnr39vLq2rlYHy9N7+A
1LcdZNaRlmjHtO3MZQkPeYsXXrmkXPvr9k/vF6NABShSaOyNnGhqnQ+cpVEAoRrI
3idB+GlqYyjAOejOh8XEwtaxjpctIUBm5PkzwmfCRNpkK9SFXSkZebjLowqcUJyl
XSL9TdwKsqwMzlAfV1/Jy+3d/j0D/2nXpvvbzeaN+3DI++L0dsFfdVzMG5r4i1FO
ZNMYisiehVKgIphVdfzQ9LTyUIBvy/dzKV2Qbku9rkGoYakuErYUJRsoV2xBiwB5
PJmF+Zz7zLDCJmLbiXNtWA==
`protect END_PROTECTED
