`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yueJgpEMhkVshp8h7P4bjsP76nkVpu1hWedNutKBtcCTI/H8Vq+Ryh4tw8egDAg+
vv7y4SmGHrS5+a0ZzLKkRyeMnIKnwLgzMM2l2hazckBK38zhIaLLbmobpLV4sl2m
CBT9sOv8BEQkIzIzzzr2uydOHQbdHCSn335G6Y66zSVZgCJUW4USIqjt6OTX5+Jz
oiLsGaa54bKVUXYJlAsh108wOqSCEVIh0ngzMn0BpDIn4mpiOjI1TRdps+wnnzki
He24hRsJ680MuCJ3iG/xJtBJAxiyqIURnMoNTFSU411vjpNQiKzzTEVcZpFh/TB4
Oa6TeYvLQwy6EIBnBvf0rDCh/SHgntQtLqlyI8xkR2Aqj0JHYQrEgL4bwq2OTn7y
Bmz06LwpCEhEcxx80YyvpmyLCZK2H2PB4jULglOdFN757uesfPfb82sLWMcUBBd7
ftKZdoBFHtrfFdIFGkN71oFcsu3i/kML6+eCPwRQBx2vkBTL4qeHiBOaVgxVQsqA
zk2dHrra/FEi8AdCHhEb9imAG2w488QUE5g/nhPLbw3smT9+LkUsEewAA4X0tnoy
/WVyiRjyq+8emKuVQwhFSR8RQTsnOonQDP+bGLkMY97N2X2l9rquTa2P9IBiZi7A
hJ0Ih63Engx+SPm7BvrQWqRgs27uc9sf+a/TtOPiJ8XkSeA5IgWl3bMoQc9gGW5O
pagBb7IV6dqf/ehpLf67NSF22uEZDCF2kIalB8P5MYFri3ww9687AUPp2Ioy3xRM
jZe1xtTSvw7SfQPNZYxrLdot5WDB66rohPzSaqU9by/Ld0ZKsBDl1jshXi/DHAVR
i8nF5/7v1DdHXBa05AaxiET2e25XxGkzDzscJGJDxqpE2/odAVpycaUnR4p4RqqA
07RB29Bpbr3dp1bfYRTjI02DBJFHJu04IwRI1Ia/Y7db+6+Kn0rhmanDq2qmBflP
dZIUpyX8Nv7/JkwhiSCiCCdk55F5yf91I1yBwkVla3Y75lSBsgiQeCGaTd2yr7Is
VuPFMgdfHae4sTKsV41yE1JBsEpkLnQ4D1s8hloaCbxh+JVqDyCni9uUYmrzZPrA
NGLnbYnXFDwYKM1I1n/Fz+y2OD1GMEp7hk2jfzAKlQYORBYqqQNa8uRFLJsbRgCf
UfpreaKUBSVqQS6pzOrOzhYZY1Ds/Ho/gUpg6mtZF+w3gNCm7cLHzjicUEnnc4Gp
B2s8ao/JxXxuqfyHXEpKB6dJl1hwPvk6yATIANv0q39uQo/+mPAn5Bh2V678E5YO
rJlElzH+VrAdd2AZPgszxQ==
`protect END_PROTECTED
