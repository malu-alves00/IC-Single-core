`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RGmFE77+zO70AjkQBnkZmwsCB4LSFFpiR1L8qu+VX11DA5pTeYf+lKnty2rFobWO
Hvb7tPrEGIflthUvbPi6x+OQ5UGyZt6adqL4YGhiDxh5idLQvW8rXXWAxuzeGgBw
OwpxQTCdWwA9uHv1YwIibSiG+4tO/D0DZZV8wh2JBrTG+xFI3YtCZd5gKAcpgtqy
jUl2nU3xXb9dKHRp140aACzTC9d3AT3LAoQHBCRFJLyri3lsVQJyFEO4A/Skk29l
V1t0c2ZROWzrnQJk+is+GSfruVXMfJc8n0Kvm53VXeuvzlkZzmREUg1kygHAKy4f
eLvh+5Cp08C12QrZOgdXSSwYt0vKl05hDYUcr5xMDVXHwKOjnXPwKz4s5UrYp4RK
bNC68C9TvbHGg99qS08/woJbPcpDtcuGBrPVC8KgPP/y2qTiD+GD1dn9hzMGAuuY
Zf0U+e2S1eBd9zZvzbkFlfr1ADcW9mtU14uVUAIiF4Hu0/kruMiO3oEtvl0sloW5
ZXEBpC4wpUofDZVfuTBSgefh0l16sffIJ0zbC9HfYM4ZsRaLO4sKXbMzSaSwAXrU
nugwMqD6nvDqWnUihb9uDN+1EOh1bpPJcdvE/UydyAf2sW/62lw44rGu+1BSsrnS
uQ3A4kiGUGdKt1DIGL4MlVpNjrIxSM8vZiz44CPwiSL0z0J4L/Q7gBhko+aE69Ii
uFv0nD/ZWcJE0LLA/3ewbQmHSSo8jqhGltI1GnjSpb5ZBL7j9GJpWKoHLALU4XkT
Rwx0lxMUC2TFk4shPT9t+1mrK3SYwB3GD1I42QEa3VAIzEBEBJIaY6G9h1rzVpou
qa6xRNFagM8EsV2YCwtYweLJ45h634rZ8zCsFZH1qSMPSvhUHrX0orZ9iFgEWdks
B/IKcEpAuRGIIX+sVei/3uYV/3S3QRJ3M1hequvqwxuluCm3NWfoaWyldpHdztEr
T5B3pShS2iyLNs51fEwY6282sFOsY1n2QuV8B9P9XboIneKW1ECnko0cbb1kLw34
SQvb971kD0WEGOV8elLp3RdmOKN0/XW42ThmfgVyiWTEScllebOQbqlXcz/7qm4C
tVUZtmbkU/a9n81ehoBINT5rLv8FG3KR6Y107g/2Zn5Q3RYIXiq9HvQrV79lOKTP
9Zcm0IpbDmONXbtb6O81UhGRBBKcpLPiSiBHVklxUkSrjt41CzWffD3q8IghDTCL
DkqD68Ys/DbJPCIka66KEa/6u54+W40dRqtGnnbr7Pk7xp94F4qsjU372noOA5Wp
F0574HkVyDmbKkn+dRnVukkIN5OFvgdUE8LTtZar5Di4+q6Yyh4XvAwkP8PzI7GO
Pj+Nl/yiXDRzWf6CsCjsLRbtSVH74MdSzz2hO+eqGUccfhamz+ZgF3s8iMDfE8ol
EEA5UAgKZzFYlq2O7C3n7Bo8aVW8520zmkTe9eWZOj9ZfVdrHDETr1+RVHTMG83o
g7b2SzCtLAn4Un4Q2QKxOuyGkmKXgR1n1wJ8jn4hhMnO68WxNT+0M1pp6s6hinEQ
qDrUM8E+7GLjPgpvR61UaLAJICF9P7iWpAoO+mqQ2Jdzp9+Y+GYoyMLDzM9ywDL5
fbwbI+/R4LU2nsmH6sT//3kR4D1Hyj6EW0IDHXGsrtED630GxL9PO4YXIT5IStr1
PmD/1NKC4MjP/5K+OndAKlqJFL2Pzo8gw08nSyiH6qJYke6N1ZiRvThNuUoAZI5/
+PlVL7EZ6rD3ZxDcBaJokmsJTRZE9ehHKafLkdvv9v3dXgpFN31cBIYtsjfse80U
srNm2CTpzukdT5TjBSlOn6nxwwsRooPvI+3oKlsdRoKrUFewu0Ya7zDkv9GPMKKD
B2i6sNuwTYXcjDXwOKLXETa5nruh3DSwTUSS1sUQ8jmqggcpHp8ugPsJCqIBIByM
UHwBV25dG+m9rOp88q/IIHeSVXit7wHkBLdFc/L4Gic5tqOEYrGYiJY/jdoXD6Es
wQMHqmGk5Eot9H36Gidq9Qo415fMHwILp0JCzRE/lTB2jblBZmV9By2xWe2KkdhF
aqTHEPEb+TsrJfHEVNDsIZ5z3+H8I/MZkwZxQ3ct5Y1Fjkj45yEnX6seG8X8B1Yf
kE8QPXQ6s/l0jKDFrDYRwP//wE5GVt2i0Ydba6LUhqVOE1R9QJVwa06+EU7973/i
DK15Z1I9xFX8uH+IPtBDA2tnihdxdkxl5q45pPsmc5c8RnOy1dTxcv3yi61bj8p1
NqWZR7rtSWN2S0yf+m6apw2BtaZiZtSTv5s+HAMevZ/jGSVBNVpE7xXzxrskzHKD
RjKNny6K++f8rJ7z6ObbkEJ62dDXfNsCSMIKK1L3EYhf3AJkQ+FBy2pzGhdnptfX
5RV1PDIZVpjjymPFx2I6iZ5gJGSmeLRjgHtLz6ifE2L5s6z1iml8tRRHdiwZ3/sS
kZNyPVySlePQrtleU1RazS1MzJbre17D0iavoQAPtglDN0sVCbaioBHctzAGzEVO
0rH8LZoovMlZrptRDn8GiFaFUr/+KCqYO1WLUqjAc1x86akPSeM8wiyszq6RSDso
FI4gFIwHdLKA5WW8Oz2QoYga+HxPkZG8F8tEyXk8z2BXVAHEseGYByOD1jSEd+er
47Br9kqdKXmOciSjm2hLETM3QyhSsR3geAy8102Gc8y92ZtdcJCt77k1iWPRcqi1
bsUp68uQOas+rps4GvfJJADyahYIcWYQUJy+3z4w/vUztnXnNtbHtuIN6nm/X+WT
XKy/PWnNjdjnLF16NbAiugUR+cRsTtM7oJvz4PUyf8JNPqXrkzyunwq2OgKO/mn2
URhFOFpUVvUpk5EM3nM0hjLtoi9/AqgGDQp5JsSgibzMYI8WOcszEFUe7G1MNoTK
0QAzN2vy2lDxYZd7nw/Fv1mEMDzDtIgG+Rg336mkVo9T290Upff98ldVIRPiOxDO
RoYtrCkDOzvrb26jLQmTHJ5Q9RRn86c1XaYrHj1QHFVjH7rTZBpuBQiUGKQYwVqz
1OR7OCt1B5SkI4ec2HFZ71bPzfbOrz7Pn/LVuloDEj7hd+ukmQdNjVikg8yfyh9/
bSAZeDiER/zLdkW2aNK2/KAEVMa/+EIEx1Ygci940h/cKYH5snKdCbg6QEvCe1mG
07uCnVPwEH759opXuT5Bi7axyx9zVxf9ZDLQLEB8wjbma16qEUTevAC35W2Ce5r2
UFyBFc+CPQKJ4AXxa9Ys/VRwDIBbfdrp24wYw6jxs4EjEr+812uX8nup5C6g7rP8
79KVyBN0lv7VZ5xvseYRlKZvAAcDLZT0L0zuNBYOsdLg5QFXNJ3+naAJ4QUdItat
bFdkleOrq8g4oHmMG8adMa8One8EOm6u2DfCJYChisjvZaTZYBYmhq+ZqkXKv5wR
BOW5MES1mWPsaOoH4q9Bqz7G5zA0hTaa1R472gO4tF+MT5jkBLicF2WO0hMtVJpJ
7m04LHt719hVSxPzBOuQnrWlptWU/deGUTHcqTm6eAdou+MFM9wrOnp4Utfva8cK
p3T2Q/A547d4PMr8DcRvvAlWmWxH76sGzXD3u9WEvH8DeElY/WK4dPxM/+f2F1mW
Pz7AcJkLwjG3ax004FnlW+6yekmzIIu55LhRPB1VbygTexSNmIf03uWbashsK0+D
xsl+6fHxfBzIumNS5wYE3b2VwXZKtsfxcDzkBht9Wjc4KvO1nneCF9EMCQbQhJEB
Bu52okLZVfIOmuccwhpDsWPboua/eNdOLCYtdtDmcbBzGMm41RuwqKGK99ayy3oo
HmMw4zG5cyeQ+6Vnr0woP8AW8+FYasXYohoLbx8Je+TfE6gaBa5XAn7MhDJhXSLi
Gzj2BmynipF3CTahv+NsaJ4NP3ZbiMFYLAo0gq1/EMoP3fYR0Rzmalfjgqujffe/
FdFKd1wWqK2TG8L55RVLjSCKGHMlNOpSyZjpgBtUfQklMwy4sOptFLQDDorhR9Jk
dli+ZHTxizJyObdh5+hoHkzlOZa6yETJwjPz7aZT78iLtq2zrBFutGAIhTjcUNcc
abs/6Xt/gBJckHOn0sSYFQ3T0CPk6a4j+Ysjrz+OU7YUvA8BYPgpGMEHsXj7wZET
akdPC//Bb4g64wmiwVaXVoMZ0besYQfK14zI6Q9Kd0Vc/P6BsbeYRcw3VaGmKcr2
oIyjiouWL9bUqGWtf6SHHxU4YG89YGTOuig1xYOaBuRGqyF+m8MITjJBXeM+ebi8
c2WDzn8m0LrSzMIEbZgpgkrc7TkHUEOOcjn43Ymjqarurf7PbKARkDt8ntXYEsA6
xJo9KEfJq/nYLGV7IjJnYSHEHOqY0NaExFdwq+rFpAGsULbRuZmRFqq19GwTOwl3
xV9Nr+ed+hrcK2Cf1/K4r+uxrYAqNR2U3J7D2r1u+2HYAiY4Mdna2eos2n6v3nye
KcELJcV7ZgPIcYYLrPYVdv6oM6nmXkD2wzvy8JfPEd5clBuO/2P4wurSiVL8tgLW
3QuLOGS7YINtJh5HANaocBQ48gKuDAxF67h3ICFYBL95WGa18HTrg+2nGeHbe0op
+m7QHBLK0kx5bLmVYcr81zHx8XVeJeMV640ZLeImhzeMcjPMTRPqornQ04MI7mrL
6bAwsLZ3Y6BN009TD2oSl66iQKEqUZkYtXCi3D2shK+c67sWksHJSdnoXgXm/5IM
33cO6+kob75SM6kPg+qCr/OPkaS2Say58GoF1a7SOvl7DvMXb+ciAXuRLQv1uzbP
6jXdTnSvqUNQ7mlAXbBRHn2fnwK6l8FphgVvZFI7wgEGcgF3C6q7XGwUGwZ8Mwiv
2cgoeDSKLYBJrEZnAQj47ZiSqNgnJ5IlGOJDAL8maKciQm/A10Gmi7Obrn6JAfjH
w5ozsP/rwAFktXYLvc0ACn4fTvSs5oat8FNLyJwd6Qx64X07aLKG4oFqJEZDpPMT
9B2384hKIN0KeL0sbtmOiLw/rHejwGLP+6osMXaiiaXweOuf1VVW3hKQk4Y7i8D1
L51w0WvORC0q/U8+OSB+7qS/OVmRsIxNYPw5iR/7+DolBLDz6VPIspSl/F9wJS2D
PJST2q9a/UoomfxZ2FN5L4zndbJMTEmAD80VYYSYtuAju4YH35SSAE4GmWgeDt50
lZUTnjVWFihs1c/Cr4xBiG5T3s296O4Er7wSIzCEQ0bgC5pFgnaCb+Gm3Hml8Dfi
SlHChawS+h9TOdkCSznAxqMe+9lLLFQwLNX1DAhNGBWJNTeZU0gKEEoCkcSkj6d1
gMK9d+aa8sGti2DSey4n1BHSOW+tgW4Kt4MVvSlg4LX2x5kzyg4Zh2h8sv9NGhBR
Dt6kQh5kZjWvF96L6xkyN6eg1EEmvTB4b1UAdueXvc5EgdrQQ7iIkOuAT1Vg7DRl
lxJEGQK+X5ayIJtfF7EIWXwas7FPpkNk0SpfRSvqhidFiqiwIVVgx0BBhNqo4+f8
V49XBFxAAR5vgEXm7DaaF7bhx9Y8eHH14AUSjEyj/GriOsMcNe2rzP8jJJi0JBPY
5a6rGAP040Fuosa3sJQHyDQeU9CYHgxIIcqQZXRTy9aKLwKvQe2DiBMZquVMeaAr
i1sIkVn63BCx1F5GaX3F0E1sgAGtdnb3tFrFdoG5eeOnvUhkETrKfjjFT7+wI7MO
8eydIZWRgm4d+KMsU+Bj9VIffHKLjdS3yvpDd3MaJ+ZNIaQCw12kAKyeDv+CqzBp
zIkBFCsXAARtXE6PlsOG+jjnk6DS/RRcjqtJx6h9YQPjpmER1WHnXeXKAva+p1Ks
/IbfKxvjOxHBqVwAsNPpZ+8m5kZEeIG3q2X/+/uo6uF43l3SghvsQkIt4o0teRd5
eaPLeACnQdY1DT+5XrVEn4eSLSnCQbXi/O1dYU4a6bjznI4sohdrkRZ1hP5m2X8R
/v7qPBTJr/vggBPLt7EOddIRpClrVRuWYl2WmrSe0iO9Nk5WVNBt9epxZK/R5vhH
71qkjHGxfFEczG8zjGpDzLs78QwDBPi3AkEPw+JMsaqj1ZhJPkVlralj0LT6AmzH
XXYCJrhzQb57G2vXgWeczfE74eQkRZitK6wVk+Xc4f4EgkNVMbIBY02LVuhPDryz
aaSAivAnIFp1ccFxmiCbBTBVkL3n3za814S62UeZ0RGubcDVB/TPmMUlUzDJ1A08
FIoCYn2xVHY7YjfMt17px4oP73IiFiMakPVnwtCcFVIbF7hR4/PK1rYVwN1Oj+Lf
QbQzYxTzkXpeJQvHc3TaCNlFrGSuMI6EiXLRhST3hcJVR0XA+ckbFY1Y20+csp3O
VNconlSPEYEsP+9lR9BjcOC3QZnnagzVSuMHRIWwrVrdZF/E45qQXfxfv+0Eba6z
kYC81TvX2wum+de4y/+lGfap7DCtjGxMdPzVUnXev7z5chx32h5CrkdxNPoo0WO1
Hj8VgRuuJSbPDc+/MYH/JAc3gvu1BufgRgOnsVRVIH26TvQUEDw22SNRI8vbtsnR
ZIa4jfUBRlVZbY3pGQmPPaqd/WJcooF/9Rzw4U0EKI387AryScO0XuEgIO77ZNzm
GNKCRy7ihf5WDMyek0mw9UYvlG9UBflLkHtLATWfaXfyn/xDRWfXj3hizy4KXvzi
Poxrm+whx1Ru/A261HAC4TxDoKe5m0QsPbHPUD62auG9HYvO9qHlOBIUvzHSLYp0
KmsvPW+DClTzv6Ka7DtLaVvLfUBuXNuGMQDff+hCb70vd+noEsS1RSsq9GsbWKi1
+S+/2zNChOfhQBLS8p/tTy/FICoXIcbiJgjj5LoLL/aVhRq462cj6c82H7QPOpim
9zQ4dG9lYYynZXrQaHND2WoWKtTUupqYrsD3yObMIbYJxXfZN0kJPQAVDpJHat3l
AK3PU1NmqJxkkwkU1g8QTAl8Z559RPB7FzbfhoB/HgfUfAP7BwANrAoVP82I/Woa
uqRPGYx3CbRG70Vd75/fFv0BIGfhRuFHZ5atAXzqRkdp/dOWu1QPJSmIZj/MGmbl
shjbu3jwK0gNy19g4ThlK7SeO8rqViNMPthGemYYsIqvWMJqNqQdFUHlroplQSRG
shY8WI42IodDxfut17RzhLrU6sTPd73lJc/yfqKLaR+yKFeI/l3FQvUYArMpnMeL
uFYhVZH3MkH/p8dI7sQY3FDl9HUz2EVz/LgF7hq5VqdopRvEHpZuyMThGFT6RMVd
YeaCAirdXjrXfj5yY3Gsg9argJMvGzQc4mzj+GgnV42Tsh3gxRfhHgWHYMrivQSK
0JkdYGJr3jG6cwHierYYEzfmN+ZkmMdrI9sryHb8NzJr5r9uHFuqDQjB+0t+wdm2
aSqMYZ7+MPn/ZY97CsmKBG/cs2OkpOTqoaJMPD58YsDisowUgRoJnou3M6MqCpqI
xmpRV4ix4530RvClDKITjUSq0IIToA7UEZLDwzWd8sotMCWwTxzD4wQkkwgLmrPU
hK31P48dfRPKZ9cQqzWhflZ3mAsxuUXJLNkQ6O6Gs7lFHGM3CdbvYQyloIo4HjOI
WCg5cr7aXIUQNLTmJ3WjwB0K2zD1us2gpvJTmzbREY3VzgjMvwWX5GE5I6QOwKC2
94fGmvryoHky8ioQZIVSLDG/GsZvHNApyuUQbxjD/l6NnPDX5uhW7yLSkwh1KI6C
9gO9q3Ox1z530JmWZrEGBzYzdZ7P5seYregO+5B8xLM2L8boNZwIKpN2BzgxaCQo
PuHG0w9qrExoBpJFxMTsP2J7teR0uYcM05nZUusCyi4ICBoTRW3kaOtNKeVrPHiN
GHKKiYCR6Px+XlyQIDMg/NFEDVaNJavcKmWrumkuJz5bXFm+3uKhqKp/LtjCx0IE
VQhQsN572PZ0qRwTPR6StkkTP3EMhfSSrMH2NV6fxhWY/E72hsDCxayDAuQRz1+m
MgRoUNLlscYpVJOzr2iSe365hGijBeQ7EelLJppYDvv8tPMgr8jDfWziEnvYVtyK
LNV4Y+slR1p8CAFCdpgZmmAry8M7LCDRxEZUwtIYdwSxN12xPr/5kyxeCRkkSOij
TImkGuBLaH+yYG5lhz89qpoU+ALORy6gbsHwSNsBBTjnafjtXn101cE75Y0YOLUU
0/b9O2DShRrSsksvyhCrbeL5K4/aQHeTT+uZyg0LETkVTrYA8SGVf+Ch71GkApy/
SG+VJVRPvRHC/7cz9ayJxsT/mQWQX4lhhsq6CYkt1nr67vCL8PGBNdMGDF/uUojC
Ew0Gmg4ezMa2umJrCMsplhOYwRWQ8U62EYw/kOim+kzxUThWDxvFtnTwV7HjWenC
KU24m+LyJ7PyPy3G6b8w/AyFYqM1JfdLoIpOBChtfI0KUE7XeGGusDbsmrGywTyT
2d7WDlt1hoNvH7egChCaLdZ3hBRlsj+P6fWX40dV8y0ircmfkyhGZHDP8VjfbJvr
StIFOg7uM1C51mmjtmGGynbEoGQsQGpfD4Yphc0ndWFiF3pq9TvqvGmwr16RGB9m
/PuRsgL1YxplS67FD1jShezmls4hRicRVDTtEO0+E5NPqwXXhBDgdrDrvVQ+BzzW
2FGKjg2Ca+o5gM1tn3Dqr1As+MEJH4Fo7sdJmAZzT8mxfJ5u1bt5LlJT7gR5wn4p
m8FOzJTWYpE3f3SBWnXLk3lyXb+wjxcezkJqNO8je+nhdsM3iE3gIUqSr+/wOjMR
ly/YIk7Yt5B1FWWrZBTgc3ZCbsMfcw8lt8Zp8RboR+fi2J02nTKl4vY6hDA690MZ
3wGLnsaiXaJnQEjWXD9VwN5CWzziHwjABvoitN4TSyGNHNOOpGktAweOqVVRgUAk
DjLHQMGh1nrznh9OmRZRSxOEvY4aW9cOZu7StGVSMuIFhKxAhuzFagf/H/1e9vL/
9B5OqPOGc1cakTrfLVwHtcOx4WD2B4nj36FFxSwhrje3WMc12HvGKFpSpeVsdJmh
wlZXMTUlzwdYuOBZGshm7R2yjgbf7hgYMANQqgYKRwjq/YxyjVCewBDpfvb5l/oQ
+1kXMiYW7XbGBQtNTGZjAfWOEsrFT2wyBlbonuWCyscFHMJl6Vy5pgnV5649iGse
834t7FHmaGD4ihIb9+nA+LuXGWNjRhbyycCOfV/EYQoTWlYX26kRcbiBq1m8iV99
e2ywT0K/TetAmoZHzV9rFm8I1WU8+VcrZ8VICq9rdY9E17C3WCRmEZ+b/Fb/nyEE
M31KX2yNrhdp3DFrzoTxyO5WAjWe6emnGyy88qM7x6o/i9HfrVCPrv5lxZqHxtRa
BvDqunHzyTnswSGmogSl8PK4iW5qSg8Y1olPvgaUzdyK47wNEpJAE+wPJwxtNATH
XxQqWB6w8FoyESiLL3/Y+5ewqLvxB5KbwpvvIwIU0rKDiR/fAOeoMTyFJt/RieDF
mVa8TiMsOa5cbhFRPCiBc9fWkelYG4txlaPAVuftJdtj795vEOIqy4nEtwf8InS5
y4jBFSw9r9C7mHtpLZIAlPKydfeq83sGCPNyT4dJI/ARaTpfB9514jYKJnBKgGdL
W+/Ng3gXJKtn8Nc1nwYuvXU9ArK478pHR6S3yIi9OdAglLlkod8RztjIJxfoU/6b
CeLEJcfzXK2mOy3QGWD5j8gV95lBYOP+RS5a9FLyBX/5fOvvIvZKqLg4aR9P1Lyz
cIQPR/Rd0AJd4KVHUwcUCp6TxK1+zzBSmUrG45fyBBCIE4A/fSBeKerBvKa5fAOu
`protect END_PROTECTED
