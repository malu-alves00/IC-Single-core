`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gVaobiwbu19ImcdgI3z33PuNQoCzzZCcyhCvp219JsdDChyX1ZDCUO7gAFkVKSzj
CB+VcgV5UGzcA7DCJUmFdBCuEHLq/dh5uUQHCwzeJCwR2H+0OWX9YWAqm6DL9MO9
6Up919JBfvF5o4ApQJQkNL8gZU+dTXQ1v5u2/HGIH6aE3eTrvweTA2FwmGWi8vm2
TZmCS69yoq34sGzxwY6H+TycBTswhRwZA7WWd09g0rSI0zXwcKvGFSdSxnDyzjQf
65HJR8Kh8K2bex5nxvdZZSHwnj6K8QNZuU0zbvPgEjcyzqr9bTLYe+yvztLeqp6I
Z8Y18gE7r5gtKWNjBmZ5qjp+1xgfJxxncgcuggRlF+qq7BaYwTFmRC54+E8Ggapg
MeKzt24GDoTKmuP3BSigg0HrUkudLszSnYlBnj6KgkpgtxCVWH2CsnJ8xXLyHKBH
q/Q+nrgY8KK/E9E8Wjv2kmASlwPU8UScF1wDPf2Et1M+QMzFRMdUigJVisVx/2Mq
E0Ypiz1LcaouNtXw2kItoeIj6qbCxr+ZBIknljPMproJ7BijQ3oUldDFjvM9sy0l
BqVSHfV+epZgSCMBXetqNqAjQd9aC/APImXHONipCAmWEpy5p5MoO9TpoEMrOgVe
1kWYxsqYMyNvXBPaTsEEuhHLlu0GLMeKaQAPmH2xrVCGZ6YztAvJO1iE521XrGy0
a/xibqMY5AdxZoWb7QmmCEloVuxmkY/TSnJfS1zXvf2CKIVKueveRdZ1Oco/Um75
7YtGt5JxsssKUf+D5kKtvWiOc2VSMyO1yvKEyt6Sj0EeaAzRd6sBRYZ3az5Sqxck
6e/swvw4WqxuWMqGhL8cmomPQt8fdsgz+h3P1wf9wrAL8Ei7D91IrGh1N1gZtMVZ
F0wsAdztzEHdSUpSP9Y0UmnXVikqhgpQPglkJH2VphZRxYA38ihWXE2D8YHIQTvV
VURMOgmwfLS1Ohw+FE/6Z1pR1zY8ro9PTHwNlc8MhQ/msrEbX0gPmAxI6TtULyPB
z9s8+ZPwAMB/WcBSqP+IW/Cw3sS7F5PpVn4XZZCH3AilXO2DXenMZ6nbWr7RifZx
/T+xO/nTznInIZ+S9vpO51FgMTwU+Rm18ZiRm8QAgm216fOt+vQDmwoW9ECJ4sgd
UD2+gZoX4X9U9iO8S1v2Uy0zd1I7wwrlgtR8UtMGW8euRBicda63F4OhSvAi/uxV
noAwG8cqIQy/lf07TQpQ0yEl2s+Ydyji3jqTx+CBQDt9xJ0b1+vOb7Uef7ZisecH
2EM9HlgqbHBuQ1ovaWFTHBAmsFabJ9ly3QpZ4Mli2TX6kRk+f3lvskstwqIC0dUY
a4IYwrMTRmmf7QNN4pWxruITUHLzy4Q7Nws1tiKzRM24ilOCBSneRkxJOzz8UqcR
SplrsL6imJx1x7H4K+tRJvJGYWrCQnOVS4PPkBOW2IivqeIj+XFrSe1YRITNsb95
qx6tf3MJB4w1M5ZMKFuZLSIBRn+9ai5DfJwNjNt6rltrr71Wp6Ki5fDX8Gq1s9kK
iI/y1VGTDnFPCfr6xPH5afjvIBwPD7yUM6GHZ6snyKfSupTDG9ZVC3aKjulj8RXW
WC3UzlcIvXSJrNJfkvi8aH790DxpseP2mcCdLftjdv8dtpQ0oCA/57k0x6ktTrBl
gipREWy515FTU6T4THVqEt13KKieYOeil+4umh6KHP+Ra61m+syWy4qIHQxiKjK7
GrR4dijw3NAJEIiGmrU+lBrfyAp0CCqle8hf1t7XlaUX1yhGVAB9o9vemf3HKeia
myCyF7rG+4oWCvP0tNkAKu6vpdOSUHtOz8jRtow7pW/4kIuEFpcBVlwmTy4VpOb0
RXyLK31xZq3WqYwGbXnYfqWpwT+yU+1wWGGG3va1h2KzuPSGdD0HsFOpBSANhh2j
ehsKn1gYozqrPrgSc8qYEKbE7XFtwGsSJf823BhAiPF0Gl2wsAKhcoE8Gbyd/Pmc
a6V6rcno86zFpLz8wL+gQKbW4soND2nP1BeSzUoA4MY6FSMNqmE4SqdHJrld1aUv
AiC1ZDi9HVcJEknB6tTf4vX5QqYW9GBPfObMSyosOzFQEdAFczIZzRbLO7hVMzWT
I22/fOI89jhVshvFCyHO9wQb9eziJWV9p+eqsyymkQvWPICsJ+iFav3KQrPp8l0F
mC2UKkxf1wVrrYGnvoAV3zgeacsNs3G3WrrlJc159tKS8YVodHLi3jN35UX8QTe2
k6WCMWUpJuYdBiSMoYQ3KideftlDyLm9s0UY2+e184DyyIl3cs8tHHh/OxStZAmm
uWXsdaMT9gdvBEtjJOGoqw5+cwFzSc2a8VOtprl4yAg4ZRyKJbJULSe5r+0yQbPq
PrLLva21BTXLXtWfGiDANeP8IZefarbrN7JrV2CjS4ggg/KQLMdbcwoe5843pvA5
`protect END_PROTECTED
