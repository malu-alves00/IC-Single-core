`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JhyFLSlbi2BRWgIIlmLIAIQIwGZ5jKcu4aG8C/KcOql0PUBGhB2Z2AK4X+tRQoT7
flpxP5nocdXjov21nsu+ceSEV+5ORmLtYn9LKRpJUnetwip8xcQ5E8R/yT/tTU3x
PVo6o5jQj/xI+ZdQE1Hdm6aW91LvgIT5SsOUxwBlKnLtG3vcAJja3MZGVs/NJ/di
jmLF8qVHQHgIL5FPVTD3WX+LJ9Zez1W9GFYnY75VaQyYancv5SKZxFp/Af1BSLum
ZsPo6MDtEIgmzV0oUomYPp/yNp4b6slBTavvLbTS8QI4We3omrSi8rOdfXXy9gZR
+BmpEhhzZw7ZiwWnQVUPZ2FDaktlgPjNpiezXFYonuDlZbekNXSZpin1ben37oOu
xjHw4Y2/xloRAqrVUbS44QFkR6owzaMejIpnPeFJuSju362j43D7cL1seZFlMKbV
ZRckMkSBhwCdZiuSTmsMwo3a3Amla3vsSjVsOx+KY9MDyO5Byu56E/Q9EhduFIjL
juh+qf1wvpA/T//QziYHK/7XjW7A/GI/M/PWpGcVj3b1NYd8MLduvv1EbvG9rwvu
CDL3GCWeR6Q3FtZ7cnOYtTaTE1LSIKUcZnZVhWyqOvtJ2lXXtj2Pba5tzl8SM4RC
pyHWJ4Mx6zxsAya+vZUd+wiUjN5Qy/xzADU3vb2y+RCWUGcXHP4zTVEnfFvBXHzy
nZ5FgawAM8Gn8S00WAinrcbx+H+/4/ETG5Vui7Bdaq4aEc9JBvPsGei1PnyaFTo6
iRBxXcBL62w12gIndbdbsn5LAnVS5o6A9qN+mgffkpF4Y0msKOxNw3K4mW+aImQc
PpB5EdVhk8p5PVSY3tzWmzS12z9G+7aSsJpH8X6u1DMpE6rZcFAXeaLX69w7cbmC
DUjsJKvOC/YTSkgWUMErLXqzxciIWfaS8b3TWPc/nChxB4KtsbjPqpUYZURr3ZgQ
HDCLxJQhiAu9LJ0ltcgwaUyS4sMuJp264zCIhZmtC6ZwfFAU4CdOlcga/+vK4bRA
AGzpND/XcL1lkEBR7wAcojamJTKQFHyLsyCmoBuQdGi0Sjm36jRd902SDutmOGRo
CH0aJSChNNjY2Zda52yMk9VGbD+yHyvyqngRZ9T5RD0QRHlsrimy1Zf8pOaME6p3
/dEQsAHWXZFwpY1zmrucoY0etbIDmiTrbbMDDpqTUS7MvduRUCfbKb7BC0eUpy+R
Y9vRhfSuxfVN+9/C13S+fVFDKH7Oun+zAMOI5G++NvH66VjTZ1v6R7ZxvSFDOYFE
ZYSTCBmRi9NNeEnfzV5+QBNL08lX4qMp6e1ScT+zvTBXRdpD2725kjF24d7n15Hj
yPNaYWWoLvrBIs+uuO9r0/ZdIy6hoECQbDPXTeC9ingj4i12hPMGBHIV1UZNE5UK
LMJkFMRhZezmjp3cOGUwuiz5xEpt6SRmrRDjxeQaul7vnMVcZJtdyOfk+9TBCzZf
GW/GLYFLD3hZ4GnpAgOnrGi7JFeRhwPEln1R+cEVT7hgc2i3V1M72tXaqic4Juxi
1zkaFuBnDqqRdiV+LPcw4ExAnFaFBmqQZ3nkXEd0tdN+SuCbO2KZ+OsXO90iHOJy
YzD053b368GeZ14HjPYnooPkkyc1auTCz61IEQ9hitvvHBlqczSbVCVP0auOEc7U
BLeOrLNCtrsiIWJm9xeonjppIEg/KST5E+qOW6FcyhB79Z+ltKo8SjRvrMV13EqL
OFHlsJTzoOCXLYxUtNSuYwiTZfM1yMvcgoFNJU5A7lLrpjUn5VHVM9V4PMdkvHvE
qFDowqyeAMofvzgSl6I5UKri9YioCU+2VOhtZFn6LbJpAKcAUJLVkSsIqvaftnla
cIbNwDcYNlkwZz0IAhxexQmKqNLDH+pQ3uDVurtjkwmouO2UONg71tTfWlIWmuzp
hlJPByHqlu7v41Ob5e5kR9eruMhZrRzdsTViAZRsjJapnajIPaPE6nJ+C8V19C0D
2V9YXJLgqTQw8oC7jqnvjNuUpOr5uCNYooP7VziC2X6HYekG+3ONZd08ZtrvNjlM
QKmbY7Oa0i/G/uo0FcbilOvZD4hqnkYw5DNXCDAwyj1CupJYkMK76FLknprUBLvl
zatkDsYoxtLVwy8O7aRniD7ju4NB/eROJlgv2ENv9QrXHDCz3W5zwBfy7nVQ8ywl
WA20aGmHJHyax8frRwjY1mmiMYuzSwrPEs98DHBe/MTtJtalgZtqetdnN7Sx5Uu6
+ohxN1/HP0z2NEE4kn3REsX9zIEKdK0lrmCMqE6slgnRsSQ5awqwHQ9DHFaXe0aV
YT0a68dYl71Jr0Qmzi+Z4bv+H3ckvPcArEtA+W+Vgvo7Ggtg3pynxancV6ZfK4ln
YQonNfhpUuTXHPheQuDf6xCjOBCHduLoe537GKe5+TOtI2VOaPMWeBWaD2cu52hq
IaDTkCn8oERapfuJ2UK5JGsEktogdCdnXylG8VjYXv8DQfwlz0zlP8yU2VK0O0Qc
U+Hdzp86p0hayvWBdAIJGNyBXmTwiMh7h+Nrv1FzrJngJB0O6EZ0ZOWmkOQpIzw5
3VxFZK31Q9HV4vzgEXNEj8ZUlfmfX/EX5uVtn4SMh9AL/tnXpeWz/l1eeecEbbRG
cJCT/AkVYHax9SfYvduvcggknYqPiVAhpiC2FJ/wmXnsakNJbjZw+bWRduX3X37W
MpIVAhjHSbsuk4x8c4kazwoUR8qecwGpNr3vaPzc9N5+wV4KaHAejEZXfVyVbS0B
LxEhIcBoehoUmiKPfMF2AOjQeTpM1S2bTI063yDcDTp/lS3JoHKd3MT8rG1shUrB
8f9Tsy9Glcpgt/vbrPehl69AjD7ZtggicNi7f7vm7q2u4qheo0siw98XgqYlHk3G
t5ASBfqFPNxjasxnx3uOXNVKogIJ5n4SvE+1IMHFZGh2uNpytuyzmgexh6pZW9dH
YwzrrYdbnTNSaojvwC92OFKidLlKv280K5sd1FnnDuVfmNPKRUpAJhWN4LOcLNmN
OdMm9ZNGA0DUqo7Mv/UcWpdUPRasEpz6epxYQHLEOLu3LO8RAK8zxN5DIoBWK1v1
8sZSDQ8YbTWXbdTwoqtE8xo56xBdEFg98GIPhqIYlNw0dYdrWVyQZPpAQ+icA0+i
SvdgwoIiGUoIZvYmUDJ2KDNQr6suQc0nFWJvc+Bj3VS46VoOanJev79S6SVH1Kmh
bRbTu0Gs5reMMzDaPw2Nn3v8QQVVA10PORmSn9BLJ96gGJkvlY77Fgzko9NJh0RL
2QSPEcgXD9/bvP8+WE1YNMnvCu0Hyw9iHINAkPUuGd6LlTIQczsVKtF623K3bPgo
WSTuyjwPEsRyfuLnbsQZMOeyQZE4IdZqhU42EJbgpius4clYjmK4uQT9TwvT6nXl
oO3QFlpENT4gmiaWXAwlaw0Nd9KILOlRVXB0DXkWialIYThVndqftUCB2o4+Poof
Zsi9GyFfxuHAFYErqC6F1qzSyK5cDK8E05vWmkkBiuB7i7tQIgi82YKluIt8KbMF
ZvDNrIlf1HJmA/e7ucr2rL1uKWZrvHTBtfbxrMzOqZSWMlM8F8J6CANCi5LpoNez
3sTI5Yy0t+4BhM9zGhLFV446Y+WFIDyeKv2/PlMv0SbcMRCdIeuD9JVTCbv58P/l
J0whBTJDsefBPeCU8ArHVao+f1Y1dPG7k5bY2vZ7XoXO8lBbW/6YwEsjifpGjV2T
KPxTK1+qZEWb3MWpgFJCU3/KzegR5KaXzRD0gqwFLD8gfwQP9pAbC0MMMg7iQdmr
EaUZcSFk1IbdBEdXDvttp8+t16hy9zgFMOUBemf2cqoncMsRKee9NcObnqdb5q6k
SpGxB+sp4CWJgHTegPASd1gR7Az93ehfDQtsjfC0q+GI8F3fOYhJ85mdVDt3v1uK
VzRhqAf+VXyA9E83iApcUk9eNxjsYxbZ8AQ8z+/EXOyizH5LNqlVW+CNygM6Bqf9
/j7rgXlH3np+UskPvdi16Tk+dFF7I16PCX6CvXUAwpSWonhaXWxYZB8z/spPTuNS
QcjDnVsbvoO6DQE/gxkCAUjIWcok5uhj/SOHq0DTGKtVZoWOStxpBdwexxpOqAn/
CFFyw89O7fWhQWIrAH7KwNq0APX7z13YEmYG8QfxqXN+0TLL5OSPguQe8Ekg4zjK
uEEQm/eS3RZ4HWv2XiodwvTKU7YCu4CFSdRXiXJiCVjvsvMskVLHuT/l5Sm0Aelv
bto9rWlWVrtukSQTRMfhG9/+8s/RSjSVXlwcN/oWFToY7FVGHZ8U1FsVUzhEvD8e
kfzER5mVMZqA8m+38jTSl81y+2fDoeTzTNorJocBqHLFDhmMo7MdI76LQxjpb4Xq
T+ox2E8Tx5Vmv2dADlNq1KPAE53ja4qoE8lvmiAL5D4B84kcqUduls3vW0dfZ++e
AUebT79G18qbBaFd3xzdkFyW6T2Gi8nVkxeY32Ky7+6w99AZvCQVfQgjtADnwhSo
0OaArQ2APeAnKVDAgPvr+dArBnnWC+Bc6uHgI7aP4M6pdZvEaPN3qLocc//YYLpn
P9dvSk+Cpgc87R/uzkvoCMqS1YKgUj/IBh5KjBjO6zFot8qHH4lKiCgxadNM/tqG
VDpg4ePlv22XeocwEZq4Bg5w+iCsC3cMrrv2gtMcx11uRShtvDoxfdLJeJ2Vhl6f
MnE7r/geWpaiFAvEk9YuobpAjkXeBfOI6koWJzt+OhlheSJlURQ477pDSGjVn3L/
KvKVOCj8fwqhTcanppKikkv0wuTu/Pd82zTJl8rqsvREUgDvDvQGCPvyAfQxw4IU
cDk1irY4YMe0uf9jUqzkH9LOh6MDxN2y0RAWFhLoH1EcuyQK+bcEqa+KXzmNyv2q
U3LwaoE4aq7ET9cmN9e5QqrseZtKyqt5qoRq7Dvl39piLdIzVbU3VTqBcA5d7bjz
PW+3Vofm7qSCO1EIV2bj5gvNUkHzdXBAtuiOaaFNk5Vkc7KvV6sxCGF+lbPG3njZ
S0vXrYByg6AVOdo108ofNjrfZS66RvbqtAxmGLu4P094vOLBrGjXumIsxTs5ozzd
N3foDd1DCeyFOjGkkoEKChiUuXDMCpwS4R/w7rOuLnsDRLB9c9D1t5vSWF+4+zJs
MjYjYYOb/ppS2Ns19EyezeWx+4isxkzBUCafW4w9l4vzKvctjzfzIwc96yoNSnBC
UgnP8pqHfVo62ChRKrkW0Fsgu1slRruDhq1Cc6XVIW4JDuoqDiMf1e/nsQir/v6N
50JNVPrHrF2o8+mtrVTL28HU+fP1SbEIdL2Yi/9oQZ5VGoBXeCA+Taj1DfM0tnaJ
kbfu+c3d5+/U5UeuqWFje+WjeWaiy6Qzxvw/GtSgakrv4dA/Po1qe1JQl6A/B+sa
UC967XcbwPfcPDq2UsJD0R2VtK0VFkl2qDuyhyg5F7zbd/l+BVP3KqsZZ2/tL12X
WZ/zmgah+wO3vYV5mij8fY1zzxTjxh+8pgy+QF0GAtCHAzyYk9X9GGbylnxNDruY
PUNuaIqGgOJegR8ndRmF4U74YB5bG5VhlFtZHXye2bsEVmhT/5B7XXV0DfmDyzvL
5+hJhuehhCYe/5BxSscniqQuO5uphu2jISy2hZrK7SMMCkDSyBrLuuMC+6YBz6U+
3DV4X3KT8Il1lfszaq8YHu+WA/M+7UFo/biBGYRgwwDXvBvaAPUcU7ite3uuLVgv
q5gCzyBMMFmldWO18L4CUGfnZXdj3gQ6A0nlY2M/ymO1zlt1D9juRQtp2RD+bn9N
aXz8HuGcwy5PdBvuRN1bsHu5gOxg8IOPkG7TbghdnTFwwIXFPGS/CpWRIDcnnW5V
CRb20NoYoto6f05Pp0gEDz/vPXflQ7kneINEEBbbGn/Qs+Kw9X3rhzkS9/dd/oFA
3KNlY8I/W3ByzRPyMvlrZ2nkw5i9QBrSpCQX2n18h8yOfLb0cPhATawXovW6SMgM
55e4u8Iq+XEAsUpc6g5WM1yAxBIaOYVx5Fw7Ahyq+ADQb+S82BxUVqmV0kBoPDV7
8aqRUVQ85gASQFQqvycoJfIHogFFLKeaX/sY72ikt3f7ToiOicl88XC9UNJ+7W9F
cLzXFMp6NaZy/Qk/kKOpPNhHMEPcclJq1FJkbUnoqpMUuT+OpIQUEX4u0ypf3gHQ
L5VYW7YlO5Avqzl/U3To4FG/nhAgksjkfIMOgtEsi+U16HHr67PU5XtURnWmErAN
8KpP3ZKn4AH2R9BN2J6Dxx6IS/mt5d2+pkaKAGFJTrv4OehFVBOO0I1P6qSQdhU3
ehvFMSnhJebdy5L7E5XQnt2JxkT/lbpzKx3Eg4h8YMGWvXyIQA/R9AJvOpv3eXYG
HZGnWukR85Xv6HRlzpf3F3CXXQS7E5R5YbTG2lGLvYuG576Opobxoy6k/H+W8zc0
tSZ8yVKfhi2iSH/WRWYgnLY1LGzCPVMqKxeo4YiPtlIKhDH0zT4jkm00zF/EeN8g
ymiNsIIWlmzqzll2yJYbKMJnZVrMWMXxkEsPWXxbYmPswiBcryvtLU1BwAFrSlcI
vOj0dYQKBj/DWeawAt08azyXHyW5yGxts+l7f2uq4ATpinVBJfyt1jNI2eCNuDlu
oFvf5yUfoklgbmXVk9De3ZpTcbsrRr2qM7UEMOwy5dG+xoyxIhYZ6O7lOqxXVi6R
vz3z6EsTldVWPZrj12tJcQCt08iEO1bDjhdZT4dfnV96vsVeDer+zuMpjpGfpoiW
Tbz+sDqKZtTMb+69osOeJ/LC+VVyXvE1g+0eSy5v0ma1e920Graqszq1UI6swzu6
QnpAIUVOOwRqoZ+MldmIjzjgLAWFx2rib9ajXCeVS2VuzpCyNZ63e5uMK10U0dZG
SLsthMQraCe276zJ0Ncg7gC9Bbv8Vyp86vKOYRrzlSw/YxfTkX15LEXQcXgintDa
0x83w5ShjWwsc7GdT4+oQkr9h+a7Cz/PjSUWpyI/rfF9MpMa0o6jYzbFamNya5hq
LQ1n+Tzhf4gU9f0GPIK+V3vZ/64fMhKIZwCQ88tbaA9WFxKFWP4TQpn+ldAfuVwv
PNYRB72zsNE+sPxsInoC4W0FPjWRMvPCjgsSP4AqMjYnw57qYkU9ZRHOwulnYe5G
xQNgs9FDMaeCYgW3g+HL4l2ZW9jiO1Y8iAJsiGpowwyxZCIrneggPqWDkoOox71h
fuR+rM6S9qo90ohMafG2UXUeGCk50UjPAzBtwH+Q1ADi1Rh+6m4TmSlEgXxNgq57
b0sPP4RXiH11IJSGG4/8edipiuKJMGGaFQ6y+aESYapwX5pXGpwP/O6+OgD0ml8G
9vmjk/a585NecV/wJeqHmneaHiQJdSH9h5oL9eQQx4m3a679nLW21zMArEDThU76
ktg7dgRk8IqtUrCqYBItNhtiULJ1jr7GKekGhNIIwoNsniGWlpj7P+bN5oeFYydr
U4aQDDWtMZbgEOuy9UX2eghJZkU34rRA6M0DVKwW4NPICObSWH592xDkY9PDnpXC
Z8eBjvpZRUHVOWxB9WnlVpyLZ85O/81KYYTr2Y5ZtXT3LGO08yTdZCzwImIEXWNY
UTKn2ugIS18sgsWOjVXQHHHH4QqWyqa/C3XbrQ7FZ1yrFU/TqP3trqfnO8U3sC4P
Z58V8UmMduqISxkygtCXfjdkzvSxuqfhDezUYFTWHlWAVI9zu2Nr+agAa1ozBwuO
2WtccHULLLcsHcu6uJuV+wOwbTj/J4+SNeNIjQi24bJB6jjQXvz2TQiuolkm2YG0
MCMafVVw0FWoc3CBan96kC9TED+xRTdx4egNeLBSQMk1XVI1ucRCBcC+ugERJm7s
Xl6w+wlny+xowVgbBvoUJD7FcXx/l6jxFGjydjfl3W+8GO+6Gu3ReaR33/Tyuzxe
EeXcjV/K901O1fpx2rkmkOdJRxT1zRHcqSul1EE7/aEBI9qYtGDqaWamQ1r8GlyB
nxQBc5VElUgjKoF4ILensmyJRdvJAnWKrXgs6irDA8FwyMA4Dwn82RKHt2vBCziH
SdK61DMts4USY3Cyr/0A1csHXckFfxc5Ayud325eKw/JFk31Pdv2U3xo67gLhYcT
sPupxIpJybdYluFIZA2F2FLFgrKdUMNUSxegyp5ZCc2VPbgrQzN18JazCGFXb28m
5RJrVKyYJgQnMsIG2tzYoGNavVXPVqUlsOz7H7AOtksB57IAjGEu2oehAtG1J466
jn0pxKJAegpKAs6gbzJ1+s/mb9mko3tDdI0E9By3/VDIgbiaVFW/J2iEofhXe5qn
oOljPc7iViRuQGo8gXuSRaQbzlloGVSciGYj3VtoqDU5aM+V9hgAChnppWVuEz2b
AtaXVCgwHUAJbpuNQcnXcHikTMloqO1alUJS+WlbRtrBOqbrhskDBiNHlLxEig59
DMlc6zZ+tJWUXoMvAIQ+YtYfHplsT1/FCU482UxFoC2XyS/DAPo5cytH1i1Tc+a6
OSjHYmJoPtqADF+FtvBe3XTOMbrmcwTr4vcmz84pX04hx33ZkuLF5vD3k7YBSTag
s6g5GS4wJHPJ7oAd1O9ySxQMLtKb+gOC+RLflBYlOfofqp4g6OVWdLTvjAjpCiYf
m4aj47wh+FdQfNgXQJDmJT2sT9vQvfq7vYfwf5enWJGpPix0pNl2p/hu6OfOfd1j
oHj8tR3oKc5UVQGkSGpUT+LALuU1vXdfmCNAbyeH2qkpE7LVx63Fl335YfDD286S
CQrcYyUXwUWv2sdfIKAHlikdYQM3GoCnBI4bGv7Qdy/mygHzyCjC8RBibHH9DRft
Yd0puGaT+zw6slflhdrn8K/ZK5TyOUsMWNF7igk0llNVh876VCODoL5blOlZ+5Ay
WTrL+wwtgb/B5g1hho8+Psj6GdFt5pskoIlkUFSJgG4GPpz9yVV9MDcHroeBSypa
yVoKXDgZ4CGzRUQ3Zfw21JgKE7F7P+3SK3qIY9oIzk9oAQHAGp8rv/2GHeWwZoaG
ThEGIEPAVA9CMSSc0gGgKtuSVToeonGZ1gh7lYk7ztr/qy044x2rtm6x2YgPB/X5
ZlA4lmFVBlgaQMt7cGXI+c5OyXUH33dBWRiF45AlHQhgd0B7Eti1KHxxgHLRL7GB
LOeLn3IWx++Do/QnTCqeDxbX1wIkdWC7sneGqxJ04YikLs4acjwms46/U+Tm810m
tpgKmt/dqG0IjglEARWrBEyMNtR+SGGL7sERcQrEN9vEnhtF3BHnMff+1lGGlM9m
sY+BrAgu91/eOMviSUIpg78BGX8u5gzuPbvDC6dCSm3m8u2QuTVaZ9gBuTxzxntK
zVSRQD4kIFFx3deBfyF4QgfGtg7xwH79nCa65SC+Ml4znLvulBnoljpEHKi7u1ym
P23X23304DOqWOTH+l5WxrXFp6p29RC1a3XTB5oTztJfJZnyFv0k6WEC8PqbAg/y
DT3lyaxZ3oQwyndFTGq00R5dfboipiD4z5UPt0hraMPUVn/0xKr0IeDobcIRtKol
RxOn4a887LbVYIi2dwwYyyMMkT52qUXziFRX9DluvOyvLdcc5ELkvvpI3scCVj4H
4pkW7BAgrXQkPf/0leU/0vOpfsKbFiHj9P6M9plZe/rj3yfOIQG7Jx8ezjPc/csJ
shJv/9AHe6Bg0EjKCsMfRwBPLoPD87K7fcpr73lt57JS4BG6VFULGb8BAQeKIVFD
WFqePhnW4VuWq9545H5KBgEXw23NRhglmH2VC1owNQ6ixtqkfw3aIatKccnKwqCV
VCQaC/hJWdKHysNn+Sjz1aQR0Y+wXOdT04SKUq7FWQBYAiGhSD+p6EAQT2rjBlUP
yJxcf4VqMFEoqa9ehnaXWNCj1WszasEbcWtLPltwnHBkNYbXe/UVvkpbWBQothw3
zs9eFjNwkkNctusvKBjNQFI9+H/v7qAMaDGxzPqnsIkyfpPeT2XSCFEaxGQA1kdw
Gy27OGwKV2yA3YpLv0eUYR1qOjLKuX5HW0uADzwzCIIhdRYLHFBqbxZAbSgxg8E/
U8qlqnq9Fe/lGCkMidAudmTD83eYa+W/Qktep50T86wq30B/ZCUJxxhVCXdPcWlm
yYgqFXilFAH7jJKxPIQ534EiSwPDzqnwVrdn+6iW7p3SSOAJSYTuEk0wTpjwDA/t
rrvEkYQIj59LvEdyDbRYmRKfuXYj2cCYf5WDqkZRAATnd5HWT2Mig7e4aahrhrzP
JIfruDcHMhUMf3DgNdgcNY98mLdZojklOs76Lxxg8a1KaylokltupQqm4uWWj98Y
XdbwVfjr2yCZ7aGLyrS+kH4E6jeKmBjKy/75YWnaO1qsYS2OOR2abXhc2X+Z5ekU
K3AS5ZHlaJTKbY10Z74qty69Bbn2MFWm5l5hIK5xYGd9d0a2sEOv6XlEp+LUyqfW
i0LgJb+xv7c0OXpktjEOGIPQSHyGij65rsm00T7mFP/RbuiQaeLjKKg2aczdP/5h
p4JYn1Vvb3dgn47rCCdqCal1kWhrsDvgxcro4KlLmz1m23uBC8280LsgUrKfpvxE
pj62faRE43ZdANhPkAzI27LaizR9lvHfl4LPjCaf213nWvfnWV7Qvc/+Jp59u79W
jXw31zaj3d7sMk6aauBoNPMT1b2ruEOyVnQ2YYZpMuCReaLBgiuqrEeYdflGUF4o
3wHrl5cVFpqS2Nz4cQnH69hhqePEGHOe17G2yMKLemrCgYPnT2jGty5KAUqWF3Wi
BTANpfogmWIGdY0ewdticv5ZbsU4hnjUIxuoyvgYBi5CnxqtIeRM+SaNdn5+mOO7
PmJ8tqFx8bQ0X0b95UT9h6XQyaCnvdyRE1C1wvQP1F0+gCjkN6E4XDqlpMfbibbK
eRrqVrdt7f1vet1PI545spezQZBFNK0O3hmR9V0+jGmwod4X+mt1ehayGqUy/FoM
MIJuR9CkW6d1NznY8XeI0daswKAT9tPZgl68QLSJjLSM6EMkxPKMMqEV4xLHAbxY
/K8uXwa5pmL7hM8nlNFYqVeCSFHS+SwNhSkRg7DyDHMu0KlcBMQXRM0kpNLScH2y
UYWDbV9nv5d3AFrk50vyuf8ZRK9IXTJtZGYU/m7UpGby0LlOjQtuO/bdLc8TVgHL
TIMXDZAmsv+ThsL4wL3QmkSEFPMrr/3tHTTGekWbDYCZnoOIysabvIwOxGndX8T/
FalCtcqzVJGJLxU9yVIJB3yTTFEQukMEyM097HTl0StdHxR8V8BbNdDSrnRVvO1J
aWEWmU888Dlq3M9p3iyM76DK3DFJNcO2gEbhG0w7wOvFQPx/U2vYetgibRl/bX6X
8iEsA8B0KE9QnZuh/Hr6aqmOAbmsIrMyueZCbYDos8TAj9ozUlIG0G2h0TPtqKdA
Hbu8OUeIrtHSg92CjM1z3ctcVJCKDkSpYGShc649LvI2/ulIrTUkmq/f38D7aL11
n0Z8OVcVC+L/1/xzAHeLMcpmfV2m6v9HYkBUuH4nlIE49vbkNluwWuuODcB5ZsN9
EBiwL7utrIcrIVFA2w5Q+fdtXvu/CMEn+0a6aImYSejRLJCfc9qlp44lZ+e42fj/
PGxKZyiN/DJElGDKHuENoLp9qreoWX/T6jc2peic9md2Qt7wnO9Q/3zLBPrMymOf
LvN6j6qB286Rp9+L4c9DtISS+GpDJaG01wfGOE6xB9ECqXWTSR2A2YJCNqGbHSac
HbE2BsLY6XsVny+Gb9qLhKZ8AtVPB9mRw/XxqA8pk98S+lX/FTLPIu5SDdvoxWJe
h4jyfsy5JvsgDX/cJrGyx4hSl7cXJm8k0tv3GxQGZJTuMPSybqXUqW8/uzHMkV8U
jWR9sMzy62841w7pHETSp8t1KeMF0EEtkwKVwT3lzqtqQ/zIlSZ9tfSgbMsShZxQ
nSvCb1cLub8bpyKBbQP6i8oKzXaYF6m6hWzaCUl1LVhM2g7g9cPTqPLp+f6ewRzW
a9PTCLAYNDuNTEx7akGskmECVPN3HYnhUbeUD4xoiI+Ymz9M1yU8e6T5uQ7YgLw9
SdwXWJxqYpsR+BhFsSUV1Lq2zy+8PXzhVPfPiC4SYanD/mpCZw1Jc6HxB4nAbm0l
3f2KAVaOsdAXz2JhFuCf+6C8OFrkohig6faEd8hRfWlqhAh8jYksb3ksdo1NUOy6
BtWvxvMqCY9BgbMDZB67aktrB8ZvyPDoyVLXirjdB9VfPpJLo4R6UsZz04qRSq1M
TeGr/AVRdDkCZqrAZ87C5pdfXT6GtJ1u6/qEpuIxG3ie5c4OBiBKK26/6/xyaIOu
P1SnhLJoY6LHDbD6N3wlWu9puuQlUSLalS4hVZfi44hiGS5wZe0wIjQXYWZq92yG
kf1fWmTFOokEYRZDZvmHlImc3ks9lOc1ZcLFmGzN151XgO7vX4VFf0OL2wQ0D+xt
5FZOe8OOyYuumf62nysaiPfj2CLfUSm3zZspj2fn4YTvHflk/3fpKy6OYiItxs8y
soIof9v8AvQ2OOmuYK6a8HGIxtC8I0raGBGrqFPzHtnjLJ06VIyaipQLVAsyFZtR
`protect END_PROTECTED
