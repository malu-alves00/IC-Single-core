`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
h02J2x72sEex/hFPVyh+RByqQDEUkOmqg0FWafBuCfiXnrbg0XQ5JQUvPxFM2DNv
ABP5RxRkXYB87CMgjBlVM5Qk1Stx3UjD+UeAMszo/RjrRYltxVzv/1UpIMUHLc+c
9S8rFI1D7AU83EtEVjLE1J0hKH9ngYCKyJduaLJj4HBmir4qY6U7UHAAh4swT9QF
yuU4I+4bb+gV9sTiaJK1AkJtjlYmsqorh7RndE8rRllda5JbEk/2fFi4gHoWI819
T7hLbO2ncpV7QanL8spOf6dyfjMOXmdpf2YqUppv8STx1ajxdZPTsXLPEml7lDFV
t4Nn/6ADMkj2Bi3KfMx4QtsnSyuDyZkLg/gSYPECNv/QtWdJJNt/Um0OsYhOnmkS
LSsvAY10y0DOdB3YNYw+k4M++s40MaeTLWZX1hMnmchEjz802Ap446pVPCFR5TJV
9+ujLtJRFfWILe+sbfY4E77ine1YeomXFSaMYYDNY6RPRcUUEtm6EttOTCnepNyh
1far8y32fxg9ECaPmNa+5ZptOP0NZCPb2yRSOhXVvt9PMJ8C+slBk5LIfFJYpZYg
RLks//o7QEFZh4AQK+2QkJ/7MzGSeYZhjGv32HJH916GzzoSLykek3SgbegCQ1Cb
XmYlDK2MZ+foB3vkAf7XfnCz9JMWDv5v5C/6gQ9q5jajGN+uTidxyPbqWKspHTsU
154efXKybvpmAp1aBCzYug1jF2NI8ceD63D6b6etHRrv0aXQypDIaecBRZyAL5VW
TIXME4Ik+TpZSlL1IF3N/M64B4YxGpji4FxOYW2n3YdVilEcA2ryy52k9QMmdIHl
8A9vjfv28LOK+8nV0JSVtqMVs6YG2++sqpos8NCM3u34Y6DKfUtDS+csTjSeuAxY
1+gOly3KLfWDrdN/C/GaIAZjIF4Wy6fTbOzcHITXlFCQXd5tZsGUWJoN6YJ/UjwB
X9npAJ193D19zkNgDlqx8bGN+zv5/T1eltxYF3ePm12RQmY1/XacxZFt+Jg1N/zD
qx+uhVVZDFyxsgkWhFMYw5J46Oy8aO+TiHuXu+WQJh+ku+x5jZVWUu/uTultLRv/
emp2EgylhyECFEIZ4P7hScGP/CxiSQ7W0JTje75vvvu7nsNWaJpPtx0f+Q/DErwy
Nli8NeJKlCRh4dCRgLKjzbL/PQyTYE/AmOtGGemZuL1mc6udYBnNRgREAkMVG5MZ
QZ+AHqUOZ9ygF1NffBUbnxOUX96vuT65b2q6jsChtDAIhhQvH0rEYttyMErvyral
ZC1f3O6uBbjcZKyE1Xz43a4nzF1B7ZVAxrtZ3jPsttSbM6d5EuZFZ1i+k9jQDQEK
UC9H3FOoUNv2ySw5GrwLYybtKcJNteFTN8gDTSxA8X3sYVfGP38ddLsDiiCuuJll
HEZYjWq2tGiCOhn0hWB/sDp5oqoVAlA3yxKVvuj6QcO9kw2XB1ggXrzED1au+dk9
v7qzzOn7/8vJx0FrmC1XT42WcQkIxM3g7r6jiJr6xELmoGfsnM/sLbUFvjZAaOWA
1xvNBiDMvNEWtha/32Opaec74PJoMH6Bq7G90K4BofWIC/cvMo2p8N4NjdPvvRcl
TN4Rxt4k/aOAG/jnkZpfMBiAyolMk2J9FDJs8MbfJcUpREb5cygp5bQoOIK/tDlg
7NyZPPO9uXqydROUd3ehlBJWxF86XkxgrS8qs9jOiJ1KzKnk+v3+rCeiBl+uKf+y
aVomO59tQAda1ecUq7YhVL2W8YlOKFrauW5YTk7IexKA7hj1ssnUbDJRuICj3j58
CNbwGqr7vMZklR0jZh3Muex9yZGBlEh++OdJzk5tlkIGGYagkjoxeA7tL7FumgfZ
/TGwmoKpjGkwjd3BkHvMt6fbm/oZJNnJFpCtMaog3CL/MGqdLSJrA79tONzDbbhT
6wUmc43hQ3kFPFLuMaRo3oB2Cs0Nhrt6FIIy25VcfViZ2eT4oAv5gbRf4/A5Ww3M
XKke/ljnZcy+NmWoKh0OBbIR1PVBmypGddrCLyNe7tyr8nZ62s4jWEg5tz7VQLOo
wzPba2hlxSL9G4Vc0Cujk35pyYOWkFPQYjE9PDZl5V3Bj6UdLPBvqnZotnYOSCkY
iX3AxQ/2+lhxDOqEKien4ixTq2AOPxuY5YAVl30q8Soqzitb97BalJ4StPhskPVf
vZQ/nhQd6g5eE3mYFKdNMjvtF4BRz9kXU2ZX/jYNCJYlF6x5+HAPjbalLJb0sBaX
c9EVelaUOxo1nNz2/c9jK2BGAFDot8k36jMQYjkBFFi4XYxv0fHvWlr41H9MOTpI
EI1v0YCZsz7l1lfGWlZhjiZoWidPXf0y899+XJ/VWnJGSwYe7yh9IzoVsamV3/ox
tVYrdIYl90Tzqy9tNDbiSw9CYIZoI6offTUEZ4pN/rKRmnfU9nQqocPBhNHZN17t
`protect END_PROTECTED
