`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
93ltoXHfk8piBsjucMBCjJadSKKKUDyP9l59pdeLxs7xVIQljGzbHKhEPRdyv70e
T8oFMy7woQDa5wiujbZRweC1R8WKT9G/pqaGNZ9h3FA+4xTkrNHLRLDxfOiAVzEm
uVMBGlEwHErEgIZ1l5SPVPaq9N6KPhEKmOMKvc3fz5pIi54ioR1fDTPPFkXOY23I
aWoUKjpTaDgUaSrPIUtR23SFj4weTUzpIXHOqs//LnaNKrRF/3Dzt5ptxeFEWk4n
G//ENODIbd2Ru2DV3DKDywYnhf4Vm4YewlUioZj/FcBrZIJPTi/odiWkOZ+5B9me
3ZJQRyb7sw+/UvyxvUhYvxPGkkXlPvgqGpLQ6aobNLRF/F/MsffrVaxU9vKtnWsi
ju6NhusBiizEFSmKz9XfifY0KmigFuM+1eg61DcY6PwVELXqA5zbKOuyz+Iw4KuD
SvoTRjdEHaDVehNpmc97TkM25qIMM+oOTO0VxiiFs5Infb3NHMRAaWddi4fIlem5
X9aKNf5q1v4OxNvkfzfWuySOwKZbSsjJyN4yPIff6gGyjglynTXsN+jhQvSrBbYP
LdtLEePB1PWEKpQqG2awsfbPzGx/IeGYBJOlZPrrQ80rqlB6/gLb/baj4k16AfPM
920jvHZjXkzz4KADfI6v0/F4QQJ3cxdhhs1U+ISEXkl9wzrXnW/mpMqAqHfDSw0p
7Lf7UggUv1GeWU/rEhrqq1DgMummhldsz6eAKbHL+BXp7chDe+irILjYwj3IHiG7
`protect END_PROTECTED
