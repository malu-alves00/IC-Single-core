`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ifSd6qVmX1tSCVUMryFACkhWB47SFrkYVuMVecrRy5PONW0Qy08KrIPwdyz5jbxL
EGk1MRAag1sJTc31+YM5JtRBjjzjmV3uAT2Sq+c+LU7qObT/9e9LJ0nYPJUeBOgm
IYy5qZ24+p8FAn3m8E7E8CX4YNELnCNYbhfYtCQMvz8SG49u1iW9Xh+AMMsyrRuA
qzD0ybcWd0vg9LaUVH75SU5kQ4cxLN5ioXpEQW0K8DL9nH/SOrka1vOQdcv4rz2L
oSDLmJdidePI5bXTHrXfPXiPMkMsMgmN4H+cERGdqKup/oMbjLRnZUwaSuk7JBGA
8HMW2RC5vDQciyBRKHGCp/AWwNqLDMI8AWiLJINyceieqMJwDb69g3bMN+nizKoi
X7Kmd/S+RFyo7DkBhYjmDeyPhX2cpyIs8TQzRMkqJvug2m92nMnohniQmGvUVj1Z
5rVOhASem1635wFrM5oJrrDxUIsAiJVUhe6zh4wvPvKHAWZu6M78uK4YEsVo4lEv
lBxYeiwzvKm3nEhsdtrTgNAmfqPguyoel9g4j8en4rWdaqf+hxtlYAzQeDPe7r8E
iYhW1vY8IvE7jkZdvlAZq3L9LzsX63otlGwg2IK52OqZfBbwL/BfvHjpumCYupge
D0ClfTpv125TgR5QOdCnqNCBU0jxVaqI35JOunvsL26PNYDAbWnoIyuQQoB1VF6U
bIL9NZCKfJ5PkJExcSOnn/dodi7xbK5M3lCSqMjuqqxZbnmFnaze2YjpJ7HC4pgJ
wkOjWCZMUGwrRdEg+nYBMn3Mx9Kyfg1Tw2oquYFDBlP1PjPWegETSTfChHpT6VZJ
EMb3/ANX0abQMDT8aDJpDsqUhLovD+YzNHzGSLA5RGbb3U+7c3bOod6748pRbEVC
Edm3jEXFwskJVDki0j8/VZ5IgsgpYbAf84GjkH6ZYVr7KW7kUhrvsyNIGhxGPaS8
S9JV4FK0HbPCaPGNMGx53VHSxRHZBe88cjwleP7gf5yeQMJa0piPy2T3JIamTSgK
Y+LjzosclS/MKQWSY75Zf7fn7KFSkprVt66WGc9TO86w5j9hK5zHSExRqxr4djTc
P82cvRop5W+nkdbOzGJBNPw7GD1GZ5UxgUZqt/k8VG75cdAab26JyTFSO4HaSQep
kqJyvIHHgksky/ErLSY9nOk16DiQkr2OVrNOF7eHWR4sN3a1I9rPnHp0kRLg+wCO
3jGxkBM86Fvm2SNhDsv9/eNEE+HE7NGDYYPMtVLmOXU+n5bsdLIx0Bx95lv/nR/h
W9Kjw6AivHJSIy8T5b6HRdGHb8PAXrPQj4tytimhEmGJSUVSs7WG6ndtcmoXjAna
bcBYmU+UF2zJq9Y3BRX9CUE7RcYIqggiahiOfRSfGbtpvg0Hkiz9SUiV9RRBZFQv
MXAMYh/AQIH8ZWzmyXhEa8k64MqxBis6GIIQtJUjTsA=
`protect END_PROTECTED
