`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
krrkuMHr5ClzEyXeKb4hk6hrV2Zz/khfQgk9pFRg/wtFzt89ufQnQ8GrbdhbausD
DrvPBMzIwklMBPUlvbfxiyycZeGenhVCcj2bVV/RM3YxaaWHG7hhdHe4RUVx1oNQ
lynVUvE5xr7FZGyWVYoAA6s9ndmGY8NaJ9DyR5p82j1asT+G4ydItB6J7CRYb9ha
CJJXCCHykmNvgRh52ieUyIKWWK0Kr/wR1/Bao0Sq/CAWFNAm3BBq4od2UapeVZg7
xlvo7Hfw7NCyE+OqUj9CWUuVOd4NaCVkEmbLtx2eE05zeORgNMtsp8ur16JQfEOt
fS+9WXnG1Xk1CFjzKm6h1zFHGnUBvUlZQs3HyDYZcgECiLV8nTLH4i5NYgT86iQ7
Qr/vqd1xsFRno++4iFbbqg6WV5uNwGjZ+HYTgU9NozFucyasj+L4uIfXs9MELL4Z
4ogFNUzwC2PxChF5si6g81MBrfsAXId9wxYpKbBgNh5zD/vFgtlxsRSP9u6Hrf7S
fwhb5cQ+TUkVY073iwPUBNSeY+/NyXwRPdKs4nX6emNkolBs3DoT90y2pV+Q0Mig
YFN3EAFTc1oeM9WVp9dDdg5nO1fjofYO+A1bVM1/wJPzi0HxCK+ULhV7eXdr4jSA
vfeGMn+ET0jOblsCDTjPwA7jqUBxjPrjIIUj4gjbdso8btBtcM7DsxQC0Ll503c6
jN/4jy5jznw9mU10mROcBsDLxorturxdwpAJHCNR2YjfyJafsfaNFUJvv5m715yB
YH6ouQNQYNJ3+S9JNpCSJPyNBQ3c+sbaSm6yKnKHhF25QPw6V71RksxFtjkTVvGZ
VB/gV9mWcuuy8eyt47bwvNjflUWLmUA/m0tjlcDlzO8narx8aQC+kmTpIXMvBVbg
luJC9LexVRiIFD32Xv2XGlWJCqLcvwicQa81qzK9qYAVqQxptSUqMjJR83qHQ3PR
wLGq6v00YAav6fQeh6VhKW8UdpbTxmrxB9Xgm/6Goly6sVjWgQGpJPpDrxR//dj9
FjSkfs/MMEVsYqkMTiS0cEX7ncK4KPn3+kTmY+cwMWEvR9DwNMGVRaFl2vxDOey/
+Rldu0T4hsaUS2AzM4FLxmSmT0tj0LerztIjDNi/ybfNog2g38SNLfACGBnJCgkK
KUoz+5aHkLx3thPylBBJl2AMkpMUG+y5aS/9T4B07YfNpWx79tfSwSlgP6TrsTwV
15FOhA5TG30nam/gyud7ah6sSko1JCZEGTHJZE3IMxyMeQ9n/xbkt3K0eMV+Zdsp
ARPcOd/7eOqqKXMDnBDxHfJH+w7ntCRL8lX7rpcwTTqu4rNeBPMlwoClHypHhtEi
FK4AKXMrk0+KecQKMsFm9p7jE02A8TxiI6VIMembjSlvZ11z3WEQRVg4RncfFYyW
4HVgRdDFrXRDJPXGHC2sFOJSB4UU7M35YGWdY7xPKiFKA8jnlTtSn+LqAr/z12FW
GRf8sUFdhXW3zBVemGRlQSYNUHLI8vKDHuF9PDsjYneQ5Ni7JTv750N3xIhI8VEH
+QrP8uSRzr+2c+TTbI0Be6XYgJmtzrwCQQkVOqTdyTh4KN82UzObXwyKDWqrxWY4
MSCpZPikgHvdnMmB0jeZqpI2bx2/ulaJ0MZfFJuRq/d7Bd2Td1ULwoz2OEYf7wz0
f4qu07zVlWAzLXQThXNfLfD1Fq47NtE+z0lLi6mQTq6+C7imHzoJnR1g9OYg4CCg
ZsTA4+pLCdmWMBzkog4Ur86bLxE/YzCGx9EoF6WcLR7O4yMhZ2dpjd0WgonxQa/u
vm/CySRiQgPQXRHGWIuwdcOWqgchyMEgub2aaJ8XSmzyctCND4qRDT176Cg+I/Sk
dp7atl5qE8laCBrcz/94rFY045jqIEvh8b+vguOCOqpGeBT7bWvW0jyEpOPBCJF8
ujzaVvurrzZvrO2+eScLhlS3bQdMFeYVXOz2MpNLAcQFI0j2G1Rc6athFtFMwK/L
YlBv7J1vLH8Lfh3almh/UjoIOhiHRKpa3+cAuGVXmGKF9wEZQzcJMrw7HNK9xDVP
ubHAem4oxSQeAKdt0byuKhcjjqV4hoFSABeQ/qESxMxYstIzIA8s+83zFX02rzWN
cuDQQffM4oV8FGah+KJauWCzV3UqwGW2yP/QgbqVpOCRIBwY4psrBTRFH3u6duzV
08/D6a/G3cwd394xaefi+9v457O9uQbnASeoRqprJ0KZWd2ZCUBJA99ibPed43tW
PCxgdDszx8QHAndMmrbleaWqRWFgXwTr/Tz6WsjPvrOxTGqy27nxjZJpoDjEl2Iq
b4pE9VkPlv9SBUd9jyh1cASek8DT8B+My7aOTw47bYR2eu9+azcGyqGBhmMEzx8m
qidBuNfp68W/aPBCgW7IMcc6zlfz0UVzIAtA9itx0JuvmXi2UXFAC2OH2jDR4QeS
5jRsbobbxvnmZKknVJnHGoVC9QqOUqrxnYoUav9FSn6pzl3TW8EpqRCD4b+xzIxg
bMHgabutR7RhiXFp6iJKp8l0h1sE8q1cVK79q1ocYUSUdW7pR9ye7xe+oXe2KkCE
6YmjvPkbLukWuG3MQbT2HFDAHr7ElbR68Ge6LzhYeX4r0DoGbzyclBao+9vEzwUw
e5u7qOCbdckprnsJAPfd+uebsHiEE1hMe8BvGU+Q/0o1fRckw/eQpwlmc7bAQJMg
pXaKHYwfawNciTGBsedd7QLatWl0FdQqxMy6xWl66wKKWbjld3eiNOlcY+qVbF9l
87XnLfAiPmbLZ7RYVWAGqjib+0uzXvtnhj4fVCSeFLf2l7qqHSsf4FoqOj8UrGER
aZZYzrAKlBoukJTJ+C8sqvDAoUq2GZWrR+91uEKave1IdVOk8vCOgXqkn4BGhmfM
DR6BUY15RCXMiWMgHYA/vVMq1FmaIk95l9vdIfYp+ewAyCzlbZQnql+CTeIZEKFP
OphGWUFCQvt5qhRVvKJj86RYVgZbtLhmQmRoin53s2cYrwi/ZqeuC3k2bzAK48jw
I4gJyYvzr0aqIpGSgFNWhBXliFcxNJFwFPbe22C/qU+eUW7Ima7VcIHF4UY3bmNE
XA1R85zUhmc98aSDx+Y1xpRNMrRv4/3QJ1iPpqZWy4p60OLJfw2Z393aFg2u8Vz1
4qFc0V9CiVwX9036MXzNth7Dk96iEG0goz62am6z6ekH/A3Zhu0JWIjvgclEF3Jr
oB7jG1h2Orv7ho2NFl24sc8hcwTsgAgDhoj8GF13pFIQOqdORN7flhwhSalRUXOU
38R5fmH39VsFXbWWzsvFttNek1q2E2KQ1eagKXFF0NchoM72EGEk/6toZYVLEpfi
StA8OaQMqZSVts+jsNDFKb//7USgSS6MIg8lSbwv6qCnRheqgfiA7X8BRmH81afD
NRkUTBL1RkHF5aUxsAc2kgugiXuxYanaVv0YkaNKM+Ru9ujzrrCdKWO9l65d43Op
HgJtTfOB2VTC1SCZMexfTFwKZHLhF3wgsRcxvwQQYZIv/sE1JOXx1/2Fvm0FlDZ1
`protect END_PROTECTED
