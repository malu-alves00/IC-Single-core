`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GSOmmo5nbdzA4YjTAD8L7si6Y9Ty8E/yB58cXBH7iBU9+6hLpXlz0xVBy6UhTinX
wIAm31HNCh1WI2zBuZwgEjSvD4X768MTHm2siB7DVM8MVYHrSVp3SkV35epyExeM
z1AeBDINQ3qvc5q2jBy/bwGygMfRqlzWhKdo1eLxmP8wr/NNGj1u2brEqTlz0hgA
Hp1wPesyf/JeNNwoEoFTYyt9JEM6AtUWZY/S+3rMkQXJimr/5Yb8MZ1IgnWwz98g
pcc5cLaqTvWz3Omm72uE8m/BE8Huo+nkj06+TCe52GkouFqDp7JYO2PBK+e4u8qG
WxEQWHEOVUo9w/G9LcK9lGwWz49glWVF1Y0zbHAoAhE9A2ZKRKq1rJBEauJbhNrz
a24+UvN0X06mSOJbF7mWpsgKndugRxKLY+WIajxd0IQG2tURKu6b48HNwWYpfXrR
g2z1f1QldUQvDFvtyBB9Lg==
`protect END_PROTECTED
