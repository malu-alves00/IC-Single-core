`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Zv9eRd4GT3BhL3IYMq2phOeZh+u5BDdhtIIf+Vw7t2pH2UENs8m3Ogku5+nAadxK
gWxx9LGyDYfN1ykHX+dD2Qw/FIsaY+J0/geKPeS7eZkquwH7S8Ji8g9elzzZuM/g
PiCA+STj7tqiLNQMbjUBYnvG2+dAWAW472couo+V2WwA+UriBH6D/E7gp7YyqH/n
ttdVJhtIPgDy6mgsEhL0BUZ1ynaa4+bztq3UTZ4uKM9W0/fkgC6kOcZyGL4FdZLM
woOjhD2ljV3bAXJwKMysbxhw17j4DMz1iCJBz5epMDWxdDWe++sU/xlXBouLB4Mx
PPi0RLMfSDQL674eHq/CYzt8/MX1xSHhMvKZFDp+MKIPpsECcrn3aorcBf/CwFWl
HK10DcBwtvU8AXPjPCmzpLgFjZrIoDl7nT6gJ4UUMg+zaSz+hFmeHcofbWEHljNe
zbRgPbDsph5RMu0hlAJwG9HbisUBW+KDG0yVkX8LiRG7Pv4PJeJL8UYeKFUAXcSE
VygsWM1Abe9pAZ5aumeOOuVNm0s0+KzfPdetLd7eCOfaFUnk8BOQVFUhACRo5B1f
FZrNtCfPX5TOl64xoRzrFrxPtpuaVVT4X55O98pYu4tpBXQUPSZe1S/HYRoYfAOy
7JRnkpiPAnJvIS9L1yQ5/F8CL4hLAioO20a76GICH500MHcM7u1EyYTPzb1x5qb9
WWoKJl0k5ZsH1vlE6YI69eUvp4qYRTt2pTdUOb8qXq8=
`protect END_PROTECTED
