`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ff5rGK41yUVn09WPARjmvcgpS0TxVZ5bmgWpXEw8dl123Y/LYWbhQPx3DPoJVhWO
XdqCXJlIWikA8F0u39fWraQnINf2qfe2w8fiQs/WA9tQLd9Ib4r+7CtNH4u5wUld
BY/z/Q/ZP9GizhkmLp61e18vJr7/csK6FNU6DUsHBmhl6/9nZPSg7S1gmjBqeTtZ
XOMx1FeZ+F2E9AIYNdh67yaj4j4jQEyP6sV8jsA/WDhlYdgxOudTJm21z7sEuJwu
KaMBpHETRGKoUWgFxDNFiuAOAhhkV3juP6f+cOGSEpcMX7C3pcSeD2IA9rENLsCj
2v0lz99qF39vWf03GH8aggJjGf3Z4YW47y+YeJEV6Zp2WnT/gDhXpr+ddWorXwen
Ojda6XvQePxLB4UkUA04/Uuhf7FhT4J/QqmGAbKwl40lyPL1obS2GMhCNjBAfJJd
Jqz9UMmpQ/UtccGmAVVqr9Zmm6bYcqytr0b+lwWRZLhHszwu0ISCI0RcZo9gJlcv
KrTRYXP3myW6xDYy0DfcCoUa8hbC40qvAuse91Is645SAjVKtMOCiaq82aQn6qsI
d+5HYyKK+U9vhHYO+9Ud5vYqzl5slbQ5JT0NRMn8GwGWIbtTLA5gAxQ1bMzaP6AE
Izg8CnFs2OtKBRhjKZiNid5giAQmji/uq6nWpO0+j90qyd3m/tNofqev1C6XMijp
q5AHxDHmHVKtDLsd93FtLxEZ40BZ1yhe2r0IYdw7KS7va1novkTXjhmtyFEvMhuK
WjfBDLttmeYSiOYzPapWmr6ztaBYAC69tiPn6K6U6mbWOCsEzMxBG2xeow67oVvP
kzLeXI23EFlN9CALqDcJrBP6kVMA/NDJB3gPnNt+O8FPKQ9/LfuKSezuZm2BZdZm
wO3Bk8OAwW79NjDxoF9+CETch4dxm7VnnM6pKcepLHJbre3bDlgFf2fVIQ6EgIUU
`protect END_PROTECTED
