`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
E75PW02itwUrBbXcP/NYojdQIQCMEPWO/gheH1/X0VrhA9NMjS/pWKtnqDcXA7FE
+/NcKJK+TKMPnhTPjGoOFylFt9jwk7XEMTlTlmdMFM70QPq5Bceff+bvNC8or3BN
jpLlZMssuoKKLYBj9mmsbSBBTyYn7ORVWgstR8DCvgsbp7jjx8zf6PO+fzhnfkDz
9beNIteUjJcCsftT3Vr1BOX9Xhj7zR+4cLGIAFjicT3JvyiNw2ozIMHXrx0xxeYr
k0QMb8ICA0V7DKKdX2gcboGgj0YzVitnvWDKirwY8OkV2eSX6E6iMmddWT1AG1wG
efm4W2bC6On/GmIz3Jlc4J+KLZtrHj2zBrteFM7dkRBV8GAlVqdrHJgRNeXenDMz
DVLPJB9jWzM2X+Yi0VYPVE6bZemA0fRVQvVzqdlUZjO4fz/udSUmGxQwPbf71cgY
3e/NuQowCEU4Ii+i0AlRiJ/lTJu+YETylyQ/FZceisQYFjQdIg2WR4534YQfqqFm
/IQZNQKxSdnAMxsqOJ4OuY3LvQ8Xi0XNbRyK/JDeHjpCWYSE8f06sju6LCvIOOcD
unh+837ln92uq/gDOFBVfsdxlr5GFhmfHA56EBm653Kzvvd9cLtQ4C3cDtuemt6A
OcBNrSF1O46tEMyQmus3IRdAVJdpqlEiPsibaBF/p0gTtcsCuAOjnHlj9t6qzEsT
fDkJdAPF7v6UHi0Yc8RF2DQRRJzDUuy5u5biifUILcWMs9B6VIx0QXhYFppFnML4
AgKK38mfxbtYlA6jGLQuyToAIIXVx2KXb+YHnBUuSYeUqQQo1TX61I3Hd5om1xjj
ijc5OqzV8H69SqRf75ahlWyKjaackYnMAT+aUczQNM9EKpxYBqr/EeeQD/eBO6Nb
7E9WW72OElo+aFVdlb2pglUT7BKK+dnpzpirJ0/lY7JwbOCXT0k0SPPC+ggOfU9M
AJpEzJu58RSfC29qb7wqvf4mHgdpvgdzmvNXf8FdUsQX1EJxfPHhgTJPivqjmjr5
rSghqLlG1rKq2DNnZ/pzNlt+N4+609TCrue/DYs9YIvFLip8PcKqEc/K8mMREWrm
H/V32R6FuRwOwB9MxKPOFjez3djk7yOm4BCphclFmr6Y/DBSdzMT5kbkzF0usqFB
NLDZooA+1/TOGqUPeiK2Z+8ALb+AdyffcBG28pWjcxBYoNgJi7Hj3uHqoOolUze0
GfsMeGVFHp5KGDHyW30b0xZFmItP0qLbmvOb90A9xDl/w800FVefiqZ8UPMjTEAP
bFmWL7ZgOZ2sxBNKaep70hDTsryAUoc4EQbRaCAlEZJPeulzD9om5K7cU6uUiGkd
QrsJHMKQYkpwPFSuDVoR/Ky7lV2Eg+6sBBEmDdeneyhXFjPuBjpxs9Xi82agkmni
tvmTs5QQCysGTmD6PhrKM/Bv+4QKAj40C71le0yrS+r+EVqgWzQPNiiqfw/o4ehG
9Np3L03L7V0ea+nM6NI1zH/xfGR/uzV+mPurF6mHWs4dHeLsahkaogHkYzrJrveG
qfFWqrhNjjZwbWNZbBh4ZmypL9GzqNV8Ctesgz94I5uhmw9u1G3Zf/xEEQiAi/Rm
25q4/O3Dawlc06jFTjoBhgmHbwbUQf3FCtYq2KQBFd9lsHrvCcaBgWeDHDZHIhKS
gXOfMGIwwrDUdDmmpkelYZljJFSrBsD5DUrQzQESV2IX59pD1XSQ4ArWKzB+EZOS
/OH3bdTOKwDgqbct6/Ee2RaJNTLTzE6xRdzx6CVnkS1hj13I9TY2ai+llI0H3eNK
0iZyCRMLzsVgfWmLj3hQKb8+9rE7TCtTlszgblgfZh5eC2pqhwv1C4lRzIrSh5sF
WcbRa1f7A58dDDQz2fBgpZ8FpCuaOpbYdKW5OCzITRIaMnwSTFvtbb48m1fXZkFr
/o83lt4Wv2E4j+hI+gCp06F9rKkPYM3q0viDmGiamCo=
`protect END_PROTECTED
