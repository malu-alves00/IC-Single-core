`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OEod71jRWSdha91IQcLYeE5heA9z5f2OtIv+GBMqpO+yKL39P+un1FUsvDVLoha7
/daxDZL8feVEH0szQDlnZa48axpBrY9s52knSxkxL+TwXwvLzbXamOQ+Kk2dGFDo
DQtApq9IhNdr98OLKxqGo0u3XCUtcSyuHUhdcHVS1ZsYRKj3JnwLTJxfHBT+lBPu
P4JTx40e1gs1P5OoWjFZS5a0HG2mj+OvwH8FEaN0FL+DlO3W2tnyICs5J79KmRWn
tja7SvMeqFTuDoeWTg22yHB8/u7B6ED1SfdVybVEPwLjH35D6iDnsfnrxmnxUSA9
EIvNVqGnEfZFokZwGeF19wPprXFCOmrNTzM10Y9FFHTfKU8rXwjuNlnOed6Op4vd
kT76imX0A/mLPYxh35dVQoYA8b8BUSfwlW7DbIy+OhFDxaWx7d4Wwl8vw0L2twVY
ZgmwP2JANvhjlKy+3agjzwO6qof4o6kCRc7LrXbq9LccbC7fckX8UnsFOb2Uh0nj
p+xrev0Em2+3DuTDLTE+Zu3A1hpotl6LAlaadDF85EZ9qNx1+ZC/mjNUZ6fK5dkr
YycujLZ1D6yhGtvm9k0in12A+sVH89jEtgjXKlwj3vi+yx/kx/TG0I1N0JZTLAle
XWtNVXe8w6NDwjqMYkNchQ9GiRhBx5gbEHfB4BxSdgQ8254TNDvsc4vvBwhIDbp+
yQ/+ffFe8g3YKNS7LSE3dqeHXylNsU+pDga1NjDHEz+6nwPjYLOtRVF4kImhf2B+
lg8MGLuqPi6tr0yJubsqHZwE+F3rjSPZ1RSyz+k29iUugSj4RI46QsAeIBM/UPso
CBm4syd2DbjPGHsSvzL47nyS2cuhn9G8LtbznuykAsJoAyo1lyu1+JK9vLXgr7YD
4CjkzNtqwmzuV6SyPI6TwJgZqZcYVOUmVmhBHmRmJtc2hZMeJqL4Udm9Q3g55/+7
MnQbI2DhnjJjy60zEpJbgIqisA2iMV2OCZbiNrG8o1GYb9DkNpRZTPu/jlYb6iY4
VyOwrM2+ZWpA6G2Smf84h6tOzmAwA66bXpizDaGdnL+jMe3hMK5ZDn03O62eDxvE
UvRClhBeY7UYvC8msJq1MYilDxRsUk8ujHKImSAca2wk208Q/P2JrZlOb3sU5Y94
glLnKU3mYwTq3q1/PXbkw9XouvdK1Vu19FHyHuk/eWafkvX4wLfaXFdJvTNWmFhM
Rpqd4KIUPy+/ydwbrsIXBVhgVgVP9vBYdiNaAzdZue0+6Vte8XRz98Whw5LlDV1y
914k8lv9Sr9OPzUiyO8VQU88aXpmiyoa+2nRfrhtklXZT0Vr4F2huqBBFYrIEgLl
Y63xb4SNq872QXTS1VtTxPwG+uCbdfLGl/cyTjuTEa5X1Q03vKewo7xHMfB+ah3N
e+dFFrerXAuBjNd0UNDlMRgDAUAcPIo89mFsKr3TWdI66otO2QyMX6RJdKU0cfDA
WvCp/uBuevyf4N8X9h3TfxBzVvr+6esWB9rPTAvExhMp1FFSaVjVuNzYWlemC/tL
pJ/3vXRJk4LnbCeJ/X0RirXXhDU91rmXebopFtYB+ikdwpK+9sZb6D+23hXopRDb
UyBIKzaqcpCv6aCL7lB24qwfpnjjdZTIZg9vVPbg81YX46lA40kwDvTNYLmQvBbc
YnyHyKuhEFuhMKTyqRcF9VfAdl7FexWiVpiC1/wN7Xfv+kjd49ZPGNXyEUIaVxwh
Z2Y20iWxwjKXCjqlFIIqv59FcNTIYZfRs3pLy6xISve8FiZwDlySQiq33GseEzxR
Es0t8dONw9W91xcGaYj/nJVdGnj7N6749Z4JSBpZ3a07+5NShdfHU7k3P97aJiTr
u4dGbf8JTDhWx110tMn5QbbhSBvDSX0qzi/g6n1oE24DkaunCUw7+Gr34t5QIw5r
/28u+UEDxCrPv1KkbqsuU79tpfCeWoURi1WG+yPQ/3pDGKG9vE082kgEBFSSeYVe
FwX+E94juxuv/nrN5mvX9/qsSSrDyo1Jr2FpCxn9yfOSJRwbsLKmmAQK6P4/hJhs
h7PJDr91CXRIWBh5c/Z5mXctRoqoVX65nMhLxj0IZb4rGMJc4EAlo8fdOHlmSwYZ
qcYG/p09IVHJI6UswGwfI0UpzI5a92ILVtnCRz1/suIK3g1YsIKA+Yi3n+l0zN8t
lJOK4LqjVEIMikac4dYQUesWhU5FP3rx1a1mxm6HiWJZjGthdGpqyA/pEOYo+L+r
ffIuYJ/WpkoJpwz0uNVPrBtO433YoPpqhq/nIehqv+4w2Gkcp0HpMVQuDvLIvYOB
cApW7ClpKJs4FsTjots5VUg/bt+dXRbohO2HEDwEUBtFxxkt1yNb4foiMluoQfbq
G5bnaj3y5lYbhcAfVFfbRIo6QlCxWlbKkl56UmxOkkBxoBtK0R1502kS+67FglEn
jQu5MMF5bYo5NAvQB64aVA==
`protect END_PROTECTED
