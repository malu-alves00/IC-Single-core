`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pbcXk4mHZdo93jwvjEC7WYv8NxswYvJQjZwD0WFaXCFOoompyL5T68P3pqXCzL67
qsp/IME32TMrWFYb32Vd5wU8fxxL9z6ejBeN35bDqQ/J/K+xGPNL9NjaYOm1hOra
RB8X4Y/76a009dnaaFl+HnmHOz9moMopWI4V0Cc3NfB81TrH+AIv7ai6M8xB93Pu
cRRVlvlXODK5/1ADtX3FbmNvDe/XrE7J5+H6ZtcLwH6RjiHA8UkXdXcFWPf7aAa/
fIkHQHuBMXY6uyGQbZ0YKES8gKrhnkWQhfEX+z+7kYvF7I4WJzGxDNBhNhieA9Xh
6S8kxRTvuBbbPdrjgQ7CEWr35yWU8DjJEF6C7cy+Hted/3qdKJgUaqgMV++gm81l
UIwJrgPS6RsMyh4vju41S0gM428yKFagP2VSQOMcNdofTmeeZfkSlS9Nvq1yo4ly
hG/tDq1ARcEZVwWgl3qe8RYkyNz+7xDY6ieM36/wJ+XaGtRGKfFoF294Ni+pny8o
EivBJWzwZuE8TNNil0uY7Axqzb2l6/I7gqgR27s+1PxICAPCcieAgy29PInqsIIH
HLEUyJ5AP4uAPAh5cCq635D00CVZhTeEUT9uSKgQHUkv2DHUcpJsMO09Pd0BbX0o
PJCTbNqeVkiN5JxMFYHEuQVxVLCzCmYdacLl4CcfzkNvhPmgUPjLxi0Bm0iCYkP/
MDdsY5Qgng8pY9/+GdAwWatQAqJW6VIGZuSdrF5uz2KkXzYXSjN9Zqp9B61gph/q
XxzI601oQAZYDK1xHP/wluaB4YQjD1R13C41G2Sm6k01CLrzL0xA38dTLZlG+2+H
l2Nddxvelo3+Nc9cdoiBdgIIF8visSkU71kJ+NZaQJ2vJOMh4FvIzQtcw34bcEbV
nOUZ3EwVssjODrLyH6jO4ApH2DLqUdVXQpX6RtuzcfjZKxh4TYkeF1a+yf7jomSq
/7/aKHuOCko9qYt7nupky4I/4wfEnzdPV6APjDwTflgOzggGYMKfPY8PaMLfDGnF
YkuRQnHYgOE0FsK9bqgxv/BfsOC+8mDwg7aEk/wv60Ah1PiGjbpzaJVlF+d9qrJw
ckhe2iCzWcoIsDSgBI0UQ22OfN2x3XTMdW2PL6faYnDC/dTBJ8abOt0gZ2oDreT2
tsTJGPS6zah1Gegx5g9aexnO9eHBP6bF6qd0QnToEwts162MSFYJtTskGBtA9ccv
Wo90KrxLPg+zJ0oZp6FBuQqiEOPeGy3uOlAf9fvXYxNjEFWNkzpwVsEY4YSZk0Ut
`protect END_PROTECTED
