`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+HOgNkz+g39Upyg99j3h3BGfHXDKOQ5Stt/P1kb3dUO8GXGUezSrRs5rOxKAOzi3
xEZXeIfOeYaWdywAUdAmsNnxZIA6l9ej5SBs658lOdMzfjS8fJSm9pLUDaoItHP3
IV545dZzYRDI7Z1WI+wqex5QDVFGFj1VxuR3Q2TdvET+4uYvpsD8MQPOROVvDoSO
cqAH5zkeHZlMgleBBu9jKbu3MB7yrjNPPVI56XiZkCDDswnjnQ2smV5+2fKD0dGw
WOOgSd4fZlJWbhdftUZGEXEd63r/GeE9pm377Ui96YTzwV0I7BWu/frH9LZAEHRl
62XMoeRQ6+A+/rpeSbnO5VFHZuM0rj0DhUiRIjICIdQG8w2yGGNc2ogVO8Tpt8rm
P9n5H2zkR2LomiJ4iWAwGCwBJyF9DadrtIv50VhuzmWTgAB3MQZcWelKBgGC7R98
0TJDBxs8qGLK/x5bdDQu60vO7Mi0fnXBtRvqE2zps2gNFUxcKN4IAqwMxowZSZmO
dpE6hJWl7ciuwdMUHZHXTD4a6QOqHtPOgdDYsM2SHJWMV2YZ5DXf3jMxn6KGrZcZ
TxmDkCioNvmRfctKDj7KbFRqL9zC5q5rEOVLRG13Wy4nQTRitTUu0/qQR67RWpcO
qxtbxUpPM34/Ut7k4yLlI5j2RhFhkO9SNzDkZSw34LBl0D5bK2w6+atmR5Ob8PDN
8aOSRI3tqi2dHy1LN0TmKMLGCtQZoB3/UkrD3LWsBmBueEr05XdPaxrdMbAJvLne
MLLrgERSjNwmpsa2ZIyX4fYEB46oLgg3FsbNtmJ4yUf57+e3dcJqKYQuoWf0Q3Fi
0cEfJKbeL1LhaXvldlux3SN9og7wnG7nQOI7Fc1Ocesfngjfw7hOT0x0mG1IDI81
jJ4x8kGEaJNo3Nqtldsd9y3wyYfipYCRAzLWbk0inqh7Clmu5eoQVVfjnh540Wwc
HlxHvW8/DHeIO9cTWPZX8bukaApEjK78K6RrvB1wJOz0aZ+G0C+WQry5U9o3tSPf
2QEcAESPs6KIA8AxiDmSEMjxbRPvb+imhVe6/E+NxrL7I65ldltMFqpyrOvm3h7h
3WX1DI/R/ZoBt2c5Wm4vIZ8VQTs5oyfC0eNJZ89nreS9QWvNfbI44HL5LKse55d/
LkS7ensCEkukyFjNGKYsRD1q0G2Q8ag30wIjs536cBLeduXinck8snJWeJwy+5WI
T10VvUSbpGpwnEgYav6K1GS5Rpcrbn1D9wYAqVlw5wPd9q7xjS0u9dqHeyeZ6f2k
V9gVvG/6XECRPi6n97q1YEtWBlr02y1n/z1mQ3Pvc+N8g7XwQN7W1MEHcz9GhfPH
3nqGXy380KzMmnpMWae1rf9+ZdbBieSwj7xIQYgAwkIIJ+erZj+/ObhYq/b6P1ki
lhqPc0gYbL2q1q188oopwDiTNjpbYmAufWBeLUPyB0gY42EwaB9td24X61ZwF+/N
zFX6mpR0+6v7nOqXKM4cJJUTDv/2NRXqKtHuTIEQuFI7LjcHjVXX02+B3YM/S4Xt
8Lm6O+tADQSMD9X+CiHIq35aoU7Et8dax0tV11dG+tNJVPJv9t7/vjq0bax6UcPw
UzH8HICEA1RcFR/qzuXxw7+QYEEsZ0mqRJ1h/4dTr3LUy/WVzqtE9najblhp5E0+
aGROxG1TZirlAPstFlTtIMvU7opEOSHY8S8vObOBbNReqOR9zlrdEq+pmuCJOamb
+gjqeJ7dqacRzo/LN2zZRy+Qb+31b+LLIEuu9Wq1Tv0=
`protect END_PROTECTED
