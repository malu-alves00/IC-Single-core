`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8clT0QdW5Z5SmiNHOHcFYjSxGyOxiE7xufF3TyDr+VjXnVoUkvfVogcCCMsvrk93
u4uUHHMhAUEA4DkXZ9KvDk8bQdEdUB2s07E6r50jxPnllACgBqMCBbaJpBrZU2Vc
2tXWg5wXfiN6zS58jMZKiZDTazsyYm1qLJam1TOI1qkWcisJNA2cAxeUrEf/Cum2
16xrIhe2be2aaPlv9uqi9AoE3rXaEuOncUSCMJUCKU3aWwfM8OEFhKQI3hkbtiT5
15oCkv3ND4/FFQa2C+ahO1SxVR7rGBPjXjDD5HBmEM7ivdHUzUBstPD71dc2pCOR
1jAfUxtXzmEFhyAaJqAhWIdVCoFWIQeTEfW6+WHcQXF0Mj4CdHIIzCKOmwE76Nkv
VO0uKk48rC228EjAO02vo5vCxXF6vAq3jYmGbO4Wu8tIiIRUE/PzIfZ+6mCy02ib
2gouHKSvVeX3qlTjQ/43jpolG/vIZHQOj8kHwASBFkBE+5glqXRK52EVwoEb5LCK
fK61mZB4fOlfpgck2SEhK2nHKUZRsomi+jO/jz/dIFo1o9PIRHo00I780VeSAXt2
1asvqs5pduKFf11AGqRHKY/LfmpzCVny1zEVJAP8p2ovsPhwNJyMRKG2DGaU41db
RoMarxMmHLAGKM/RFh/Z22grxSKFOd9RJYlR5y0oyeX7aeB+YV2AJBwHT+oVNTFJ
X4fWHGvEVrnswAyF5XUFkoa8b3CaGetTK+0Y1bVPAD5Pxgak9abJUy3pKvzGotym
FxGTeaEQTaHkOXRS4XgapTJ6mC66+ms4hGXRKL4dPwN03zHen1Hb3vCKej5pbM43
ERK01PbwaeTC4Mg3sGsUCNIEunuXXD1G2r946neL9d3K4xYivunnYolTo5+wQohE
Cx1aMpy4t0PrdXhb0GmvAOlUKzmpV80xQ603/k4sKghXe1uMW8p5/aMHO8QklNpB
sfJZHrhD6nlozzqGQ9JgBfJ6+ZsrqC9OFEVGB5nzaokBYgxPR5EdYnCBEQH5+0kz
bcmESSMb1nwHLR+0LG5RPdeELmxDf0pfZyibwinJ5djWfLKVcaUQtDmS+tL1ierz
1/S3roXidaKVJ24FAGxI78SX72GTmPy6RDJi2rDEysJNetd8VX8LG3ldjTAGQbot
LbGnaxNt6I2afk4+STsF4G66GqpYWuc8PvHI+Y8qOZTnPfp+fqLOrsmJw3vHAI4W
m5iBF2KGR3tV0tbcvgz8ocMUFJuXZghIrCajwSQK7P0=
`protect END_PROTECTED
