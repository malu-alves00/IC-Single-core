`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
su3vdbKcpzbDbS+GFUynCubK2QFVogCcx9IGkd/u1t8NvgJBbRUY4Xsk5amGgNeC
kxXLTiiUF5OnOaxp01rDms+MDYzuZQ9x0C6TSQyulwFLfJsUclH5ObG8U2bBuBG4
jb7KdjBHxzwFCDd4aUfJqaeJAtXIWCrQYWL8qZLVPN68w7ukuX89c3YegRDSrFVJ
WQROCyXgcT4umEA+tsY40rJraderLu5sTS72YH3r7oQTn50JkQz306VMpd8dZnRe
80RJHeyLAvlSSrCFZoJ15GxUu3ZIOkUaPq72/0suVf+Xm72DOsvJY50yxMH7CRnv
f5l+YEBFjECIdc0rWAoT7D6S4vDArIivrB8dlHL0NsdQOJoj6K1m69xIeJ16vhbg
b3ctQzo5nqA1x9kpmB0ty97pTM83vay3vFmI3v+tDfoo8fwhl2u6d2c6Re407VRa
5GYF6cRGC7S2yCyPs+jLVKPDJUrgN3WraLyeOuv3yFhQPrVnwipgO+kRi4fmBNVQ
G2r8kXuqqQTj1+X0Id5yRnOFcF+d/iIIMbsM2HSGi1wHTnfmO+puGKY+aV7yz+fB
KmMYEU4LS6D+kybVlmtao5Sqj/lBz9PRU3sYnBoXgkr7z1XmbrU52cIa+mYaEcoC
bdbhGjmq0hC/E9Z3ATqo5mLNacTvJ64sG7YVWGIXg/vtfMXl6o5CI8oLNp9PNu2Y
wo6PJsKRv99K5L+E6LusKAK25b1hvH0qQi9Q9LWKmOCNwnkaVE/BLkQH/wWWGK8h
ViZtrHYOm1dmPSipfLsyA3MZx0XQ1yYafaPDCfVz24aL937tPGFd7fi8mSH4TH3U
QY8HwsOdIVryuCuwKult426ogTvwNQ21kVDzMfFfRMLv6S9dHVMAYHLkhMWyLj/E
D9TXqK/3z1K97JZcy8tq4DewQfs+19dT4GtCCsbNn3B3tFDBYfsj2NtmTaAc3gkN
2h/Vi4hKI6TEnjtCNGpY57T+hKDhm95OX8cp0jKESv9WXE42FZE0tsMgzaqU+JbF
ydsDtprfXg3b0ruJqm0TJvA+nbfJTwPTadZvDtNfZaEh9OuEsgwZs5eHMSbXmdsP
rnWbkyQkmbEzgBJk42fTC3VNecI+gi+xR4HdOTbd3+VnBUjrkiZFMgqqy/gipCv1
01/T9ovJiKgzy1BtWBWfm7GZRkznIme2mrpNLDkQxH5AC3nn7e2XYXMwfqwznrGI
QsjW5UylRaheLP+zELtQHikLa6k9JMJ20K+RdXSAkKts309g/VysJOFiEveVw9JE
`protect END_PROTECTED
