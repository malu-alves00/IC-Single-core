`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ICGLxNwYA2mjpIPWBpsJ+/kd4InDO+oqkLtF83ijTdtDcS9sDWbNfsaTy/3DbtZ8
7btEaTvKeNhgk3QbFKl9O4UMRKZynf62wXJka3V8/Nfp1QB47K25joPqGjhgbDd2
BBC3iyi+lNAmhKaix73qljTZOccrDUP+PFwNujrfhiNhyIqSHYugh5WVRF6pKZpx
yWCgS9cUyn5lanYeJ/ZHHVR0bGxyqYwP0obzX5lSIqZurUky9ruqEqZ1uYr4UC1t
8I/MiAD11KthBhtUG6dtQtwiXBXiA3emACbAXo6sLWqEyJoKLwPemO3RseKQIRbF
H2IUk/Xkii9cdINUk/+eNBgkaghxt9tysoI15ixQycZS9jbIWCw5n64x1Wneue/f
6ZpZnQhhOQcWSUd7N+XXxYAJE+QfS5apoETJH7KyCE89iAWk6WGE+KThRlGQ/Dxo
OcOjOTBH0qoGnkAnwV6BmY5XybEakPYWVb+UHEPdJFhFHjiR8ri5LkzZ5im8dyPT
B7DEhJU+AgobdE4HDtZc1m/4qHNqcx21WBtJZzVWccuvm8yWXhN5lUIfZNcwTWXs
NRyYo21Z92Hu7doyEEZN61X777d4HO7gKfK3q6dltgX2qvqD3+bDufkf3lfoQt7r
x+pVzer8HkPPJbLrzcwSLS2OGJSiiAbfkP3pPrSRbpiREKMK6+gEfyITqP0MaF/s
dYbs7Udf+Uhn/z7BqetDZUz6kKr7mcO7yb6GVDE/GuDhTvL/LO9TsQ8aYhsFq24E
Jaw7OAxw06+Fiy2d/NMlIlfbVcPg9/qn0XDCQ3wsNnX26PyOYRy78pZw8k5PxxR9
izUOQXT32tKl/Fn0j7RK926Mg3mHZHX+liZIexWrQBCbo7Pe3XIXke9otCxVG91K
4bqA67EkvRGZe3VoXET0xHMnnOX3IHmu6a0rSZzu109Qf/t8AcmBNINxudxrxrNd
+b3yTssGCqEY70T6hd5qvzVKoPES1XpELobC9LjjsPe7JXkAtKQA4un3qMJysdj3
bdK1jUxMU/ZTnE+w+S8OnqcEL7dU+fACVclEdlfyqChoIdrmcWtMb+g6ULS/Xidp
jAUvKLh+SNob7vEktVzvcqoGO6JSdXHWIpqmTYMdUNGlVzzFRSFI91nQiHmDZA/e
JH0BUxxTlLqj2hYoWbAnvNKqCsyhCBBQbj1qysE/ZRB4IT9zHHAzoyTMvVArDUjw
3xFlr7JOMTTlyeFtPQiFXMRaTDO4ni+g2/dIk7fEA4ZceFARfG6MZcFkc68NFaO+
2GPgTW47ju2sm62IpJM4q/CxvNCg669YV5ADe8fVIOWQ/UEwtONuDjdkMZclLmLC
BnJ7WD9Sy8x4yN5pA+aAyNeZnc/j11i8k6/aX/L20e2zaXz9z6QUV7RUPiDwmFSJ
qsokdSt1y3Avh7pNQp9TPvtRPJfiRcp3uDIdkxbtGvvIlykkPBP6PRJgHXdLe257
rqwYtYNWh3v+54pdHs9+DH24EHDcf6QyLYqKrhzr8nk9m8X18FmefY8ebphj2P3N
Ul7nN3pLkv5se2h83REnB7hhhgW3iYMbIuXeqINMT18C87rdH87c1vgkE5cEyWW/
fHKk99RP9QBhVxjJIDHjPQxmxGk1U1qVa5ZdZsjXsLWoUYbtui8af5JbSGDduCOn
OkTznqCfqDoU5yhXbQ2sPoITz3A9I/1XmaGB8aknfhkbO0z9bPV50zoYhMhqJn8X
TijDOcFIBfPNSrZjP2kbVKdy9DnKhmzdqlNFf8EVVwlyBLtPqNkL7iPnFvKBvsF4
NeU3FTJ5ESZiNdx+rHTdPmhJnyRG4UVjAqFPAL291MHpLFVenDlN4IW20/7prS/e
UBkVMwXdnRM87chAKfT3Mh8p39Iwi3+oiRD1QZ7FAUZUfjPwXRV6V6c2ELGG5DxO
ASR5Brhj+BHQft1tHa87JA7fmqOB7jezQQvUMQTPdcwpYhviw437e2BYH4x3B0GQ
HgE3PSLGGZePys69LaEcQg3xwwMwiB96hMeWEAthJKWRuD16UDVTzX241zTbnueN
Nk5mw0UQab4N8WNUu7zO3yQ93wcG/WVNyJdAbXdTJUNdGKVGB02xot4RIELC6hnF
pWHmdbt9+ELeHjVHCRlxW8BzEw46VbnolwGmvYT0Hv6sDYXuxqzgbUBFKPnC/syJ
0LDlXeBxVupA0iQyBRAEX9o3zhdnwZkUlxX4PIv0HYeDXA9k6dJ2fflyGv/NqtIG
BrErGWaelwMhn8g4DImqzpzFOMfbqEwqS+oqR4MJI4ygWbjep3kNMqNvzsDvuYB+
TauaRwa/iFL9cIYBO6Mwot4NLfJcT2FwgZVXbC2UEHvX2dDAV0cIs4WZWbjOVL8J
PKdmi7Ly8eFxZ6Pp3ZLC1Ubqg7JNQMTol9fLliuQGqgiEkd/eS7Ds16GO0tl/+gO
55l4ibgFRCmApTOuulTD/0FE8pZfdViZGlWwi6D73gRGNyf5xZmjf0/LNck2ku++
LAAOSY0tOw48RqkDEqYOSCIH1G5xAGJVnVLmgFGLtQuYjbMhXSidPgEOJB5Dk3HW
S97uiqbioksZvp1ZYZrUKvSdgArP07Z9METR55G0ntbzXHLdSIIU42Ul8JCjxVk/
IBVjmqIU/lpC38IKUN+aNnSaVgN6Vy1ixvoY+2MPcAmrbBapYltFJRmpmwkksJ7Y
e9/mhIVbL8HSHllV8iXW4ejncxiznPXZ/f/apXE+p8+JuL1wJb80rD42ShFEJ8dG
devfLQDP2+u4LOwIZpQIAJJsrd4Q3hkNFxoIHVXBvZyE+jpPH9iOYry3ZDGnseHR
Uf1t4v03qMYoutafpZq957BcAY9zZX4wEAQYo03vZu5TxF9usqwZ1fz8WHDzYlfa
oiNEs2aR4g0cWKjO3bQ7F+ZdO2AeENfEjnR37Caz3Pt2c5qZaamku8FFR6+RGtYj
PQx2bXaFJJ0fZTZmcu95sGXx44Bn2YhcjrMWgDKbEXg0TxafTVmAL2c7rDU6dnQT
lkFVl1HJ9EMe1Kpj8yfyol4aP2GVpBgkefwV/CKWMfCbewm3wS1YHoDQ5Avn/rnQ
w67KAUz893YoTjkDH1lZmYBDGCpoSumUyRyXYKHea582ewmdl7MmsFeGX6m+IMok
qjyEQqd79tiD1xpas1Y2aad287OIt295wz0qeJ4tJVz3SXNDRPCTh1msYNtP/xuX
pvTjKSKjKwdAnmosDT7AOpvAMDyxvx3BxanlQ3WzGYTbSysnEWJLTQMfc2w5a46a
u+g+kRW3pHyzUrXz33LU4b7U1txYYB4ZUmIcrCKqXMACzNxd6mxdF19oiyO6gxTz
nXyvP09eKvtyd0hKyps0omIP7w6fF9XdxXw5KLJm9IVfVCWreoYtI4+7ZvxKgKtW
yLkULCZKFBWz9Nah6NlbEBQ67/I0tcH54vhuiCti4dFVo1FANfh/IBsnMANNaboB
9tCzltAEKbn3UCuzLeptBS1CzRo40pm6nhtbd371zAgrTQRpPvP2/TrQ2Ln8juFv
hR8dtSKYBCdlyD5dBI+uWZn87W/GX0ellK6zcXizRZs663en7FzqtzXJgHIEh1el
V1fm85tfjmciZCDEUWFE6jO1MOz9ZXHVsZlKRSqLCoIsyNqkPBWiiwGzl7V9psq8
5Jqiu/Yrru/n+pQuJEewO1t0CdaP9mFSVlIT439txxSPqPZS8D8pNjBCWe+WD6Cp
H8uTMSN/h94xDpszK+/+Y84i9Q3KvFqX6xoCNyA2e3Too5fpWE+77YKHCOYSlpWa
hPM3Q662S0u3kQHXvwmp7cf+hIx7ssfUnTHqAbQnbkMn0MWykyneW7nlNsco8Jn6
zJJ/VnvmnjMhoZ4CVJEbCS76tJZBdVB/0iYXhSyLu5kI/MeTFrJz1NEHV070TZng
zXI1Xhng6U7maUgRc3+eajdrTu6VwhU7t3AaErof/0aB5KSkVqEzDNwmfhOG3B/K
AA/oGL3nxfHee0XPHMjhSOIrqv2ER4tZi1igAugck+vLIwpDorXekr8PSfygG9uy
CE2NdpvBUZx6Xk+k7VNSFpZWZBgfAgX7+h0+KLBB+l5lYiauk0Ga8qPg6PCU/1VN
`protect END_PROTECTED
