`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
q1SQUvmwZDcv0L3jSDGdG81Gh2yZKqUSwqA9HfTTlg0BNofZntchDqn9G7kvIXUF
5VPSr9Ot6b8phmsJIrNbH6uXx7dCK7iPpek9KdyAMQar/W9WcnscEhueCgLGuIjM
wRORZebmhv9yQNGCerq2aOS8eZ47hSafOJkTn9p9+EGPsSunQsOoWdrql0j8Pf5b
xDhOl6yrJn3JenAh9CIg76DdiKF6S2dJ2dw7vpwqcewtRdqXZETq3XWpxsIXrzc0
IycRKkg3wwmXgnTgxJvrIyi+Iv0+jPvkAOR+ONHYiMJMJfPsd7umS7vUcMZpQLYZ
pi/yn+cg0DHqx7GcWS9k/QWJWYLMRKVgoo+R3szJNoUiB5Sdjp+jzYvCo5VZkMKx
155TPDjQUybscMCzP9G7NSPYgMHdqyu0Guh3Gx7X4W/DYNWWtOhapFzgL5z8Wzs9
R3ajaB3f7adVJZzmgdpIPN1Ujdi6sO5gnnGaiTJGJemTuxbtcFuPE5t4MPUFywjF
hGDA8VGOHWlSV2BmsHyk9gvR89JsHdn4yH+mVMM8r3vDlUy9Ba7DRdqV8cxE5zup
nc2Qw/DwMFCwXbY92Krfa8l/Sy6BoQziWKtshsWfC9zYO+XlSnsMfJeaNOyr7Qff
Rlmjy1YYN/2yegDm1ft2RCwdhFUZx2OwKSsUA6FvrRjjffob7J1/wLM36WU5VjKU
uOXhEEdVJn62wGO8h50LAvqeWrcZsQ4V5UtGlOuQlgETSJefVOqPb2fMOb4cU8aL
Ol/yl/WZqoeBKuqYAncHWL9b9gvsZ7GTpACqBK9vbYbFJdqkAAyZ3/lB2i3Exs42
qy7eTns3lAOmYVnOmdV7noWl0KjAakn3iRnR1Q9RyAIF65gYu7P8vEaEB7Qf0F85
fXKmrQDZaxWBI9+7s5+0nL4CS+pGdWXrPssy4MYnM+rvyi78lAx0HCTtHyuIOkIQ
w14wKicoBg5BVcfA11dYg+H4SX+MTqongOjCZxXQIUveX1zTChOhYiAog79aJJZA
+VFd/DkncqSowEd+n81etNl9Wb96sMTJ1w/1od8oARomRqdzUYfLmzDaBIqoln2u
UvZ6hCHD0VI9XE1OgDspCTuBFP7AIyp+JV+yW6/LNXwqmD/zCr1r0MxR0busRXBa
eAsdtfSALOxxYs3D/fz/q+kKknooagE+C+jM5gZFFyybGOqW24TLAIdCtDB5ANUF
sJ5qbOEYJ+2fthsRLyn5YwmQc5Eikcp0eOKvbsi3+5JVwX6cW5MhItGFj0YIAiKJ
WjIhPdJEe9DjNVclj0Pvt2WRQX+dmlENxEjXan+0C/I2lIqjujawsTILpCSOOS0S
POXLIadAcF0L0AQZrJZc354eKmotxB35GURx2JBvupaISI/G8bH4v6FvzGWE+RL7
au5U5LkvuG1NGgbE472BZxMu2+pah2/wZADz7SVbMoHFD2NQO0oVqz57gW8PNOZs
ImdcHiC0+8AFMBioOtFJCpHxLoTHn8tZBjHZ6ud1Kp9vdYZ5f3tOXQJJ9NC2lLvK
tOC2klj9c9MR8BKBYb1RIx8WXOV+outacmFAeLdjL5uWO5JA8zCRshh13PvBFvJm
5xACppT+GAlxXN4fBz1aWj9an6syfYlNr9Fx1aIIx0fbr8j+ew8fHLSUUtolKV0v
5RoB1C+/BGNNW/QE0lzRrBwFPVyAnmAg9xe+Q6v5oUMTAMxYqQBjzbpb/ilkfPnt
/ck7fCMUsudfz23zhWuRzwD37CeoaMjGlF/bj4H+Wm9Stp7IpZ/KLkW0SLhDoTm7
pDloV1IGZ1j+jDMhGr5U8EFu3zOIR971Csvz730RrTol4yxHJH44U2Jc5kzNSXlx
wzYCXfbxjfjUo9K+FjCUYn7pdpJzvGbwOTOAh3RlIXTAtN6rPm8aOirhrMhfL11z
gXt7NPvzixRRVhG/PNcltq3DeZPOXKbmemYjZNgxpM7vPt6ceezqkIYfskeXcvWl
6GTGJD3ZlVSKJKc2I0epa6CwDBbN4sg0rGyCaOgp5xOZsP+8fBHIGULx75RMoEP4
6JXRpdrVyMvZAKuPvF14xDJEXq7LR2UunSTPg6F7lZqAjzXvPX7QnTbyBINT/V3W
65Y0XlrSubhR0jcNG2nud0KoMnjz8JnILOjZWBQC0Bk3UGo1Uy6wCmvcMweP53uZ
j6eb3D5lTWuRpJ2kuiTGw97gOuc0OLMVgzgZM7AGFrn1EhN2kYeNWYDGbMZdgOvN
DQKrbpnMD8m2ApSIuS06xjgczMU9RkUGSIN3yhFl3z8zN1WnyTDbzPeA4w2zzsjo
3dAe0edtaV9IvdqtCfl55qVFrtPdtmQDsRQnoCyoQUaN6Dlu5sa6X1xF9LhlRC0Q
UXvrBWTmugN6kqci1H+2jwiWyW/HSn6ddoKqrgq6mHpe5PHdqI0PSly2KxBNluCz
BxguDR/sN9tmqdjpOVyurxnlxxwycNrBmnvHE7lxjADxQSiXMBKW3ikjghy7FwUn
wGdI7UsibeKXbnJyYcogY63Q7uUYw/78ebaJgdqK7RIpt/cAgRKXft42rB8qNJxm
ceclRvSucfLGoHvdA0PKH/PXf3xI+2IIMlimTMO+d6kKbLEMu0NlqHU723Hn2xsJ
qXvm0yWOpzUGCQ4JrPXW1pu4qOf/ZB30LHiImfvxvkCdI3lXqGIQDk2CZa/q+OgI
+qDDNo/s+dq9c8TufERxVolfMJ25uFVhQ9xCdy4Uz7KW12lLoTPLhGZ7aDF1sQ03
5YWYQ1NHJhOJWKfP5uomMnu4Zw+YC8YVIb3NmFUm/ClvD0VwmN7ROVCkR/9Qp4S6
aDymcdIhXDu9qkEUuJqx5zXvQ0QoWNJ3wRQKkNELAH5q6WRnvD/MtWtjpHPX5DA0
oZjYOidqvDKNr/LBcVL/idNMpMv4Xr1/pr202WPuJUmtZMhUlLCEBRp5roLIZh5p
uVzpuQ9LGstFxllW0y6jV1ZeDdAsfc2et9oeWXVDnC3HgXm/gnlEhdxX13F5+N9s
taB7PVfSV+PrSNqEHQOnwV33kKRBixosriILUJvMEIRHi8Cv7if56FocbeHwhSFx
kX86pVMbOYZuQ/3ydYqoEU0IWpQCX0XkIfgsvKIOGP1WNJd/qwR25cMm/CteVd13
ZBf4euIUqlzYqAkqYhgu/UXkZWzMO7ZhgFmrE2EUMKsTzeLL82PTQinabvqZEfwB
pm0NDHs1Vn19Z1L4e9AHWaBXsvCs4WB2NubLudP3owGZ9KHqMq4TVWV0hMJAbQki
J9+RSWFvp8LrUIMN8WqMXAnLFn55RQnCC3HvVUvFZY5QsW7hyrIfdfLFW1FFUnQz
`protect END_PROTECTED
