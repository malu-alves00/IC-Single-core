`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hx0EWF+l5t6977hfEzSIdceCuv5PMIqke9yhxQpuZTvVgRzjAr2JMNMcTCPaq5Wj
XY/D5jMCrBxwRcXJHY/BrKxcDB1CW7W3DFHg+TwnR8D+jFZjpHvuvT2AgijmRu9U
qAS+RDBq4F4I1qOdQanGnd4LhuRg0HXLiM4XZt7HywlGh0JhziLJQlSZMoBY4ObV
5DmS0cKku3m7c3+FdxlRFlM9/PnO1y5JqHXDas0qLlpvqC2Pf3FsIg2jgiOPGtn3
xz7WyySgERPRJXx5AuCnz3yg8HXKuVuh/w8ctMhFYVEeZK3pPyfnEozVzbEL0V9/
r4J+IiDIA+KY7kRgHI3ZYjUX9SGERZY0rFr/rWM4/nchN0KFghe3E3Lt31pCk4Gb
WLqMbKZGfeOLDCxq5JoanY7MdJb21ISekNSeRH1KiX0Z1q9M1XiPMYUhheXRxqOj
jt2VB6yIl4Zha2/in4IiQY/RIALlTIuCa1nhHvvKkQCsMS6qCmXMXpHRXH3srCvs
AavElkuIZoO5rXnFAjlRGSiYXIyo7Pu+usgaC0ZfHCLZDDspxf6uqdyL+y4Xs2vZ
2igfK7M1Fub0545BQlsryHsKlut1/ZkwEb5nbzUyC+c1Nn4tyuI90waGVux1slbu
7Va2kTFfyevhWA8N20eRXUYtRm3uQtod2DMUw2Ds9XHYemuKIkRqlOZEHm/owLgF
EPLBq6WA6Fk4gGeITiv7ZcV7f9vHGxE3e+ftccjJdv3xXFKHG0iP/CYCO4nVogwW
Ww6hrdc9uAR3Pz8hTHYorw9HunmWy8UuAF435juFMSBDFvLEBut8knZZwTjrGnsZ
B+6Rcp0lkS9CjWrEStm9/S3VvwjgN9MYzQXyQzzUqq9TuKUvML9WHiyVlC82pUUU
ysa980zcRa/Hhc3vxDURh2QdX+5CrBw/RI5qa/FJppbE3LgooHeiIm5Qs0BhSZST
2qOam3zHMCFOPzvN99C+qDOET1+5+ZkCK/vHUtDg+cNAQHl4PlpqecCq0qBBdwFu
xixrlPfB/k5DwmkJryoavqPi5ANzkEEETsGsn4SgQ6NaUj9rWHnLQtlFOyQlBc/U
D+uair6c1mcE5/OHverPhopjO75p6UQAwIFe4j45pBpQ8ApehYEYVBId2ubtIQI6
ltHPzEYWKTLnRWYg7kqZiLJwiJVygIXcpTYovQsY2UtbV1czgPIGY6rQq003lYqd
t8jMse9AapYVjMGv7IfzcbzcbyZN7vRNJSmnmsnunPLMJTK6D5i6ezV+GtQDYmuZ
RQIyi667xAhSvzn5t+LcFe2Ku/HJeXrBNuyGa5p0f19mjNAEaLE6RZ80YXSgmw6v
RtC+9bRhWQU0KAhzDF0dpGugRaxjzGgI5XSt6bQjRwZrYNZxTMOFfRU/YiFZpQLE
Y7DzF2ZfrhfJiZHHj9SGNN1UAT92Vm0W24+opM2iDicXzxb4UKsIc9YBY1az6W69
hyf3Fp1OACinpQWPpwCezpZbeykwhHqNHzF7z9KPhK7fT5YLYD0KyyH+vaapOQxK
X36ZdMI2yN01QRKQhmBX+pA3n0jYL4DxmRg6V8L7cXp/TnbZq/I7CnU2gho8j8ZQ
WefE4p/5DbpQezINUNxhKkMbaeM6DEXS7coLB4TAk9VUoaJ9UcRPopjQpP9IT2TH
lQpy3rXCS+acVHKa2tM3ABop8J7R9FweyAeLg+iHlcFjeJ+iJq95vsi7Tlrm0O1h
kbz0/R+K7aF2sE687iqktKHRtz5hIkDhsq+zxyPeUL9gIU2I02mcWn8AklQqQhKO
tIVtFjbIkNDDAKyfDMclhcvcSPBVNB+KUZxtB4Eh/ZI3BtOnPLq664646zz0a1p2
GfGXcApuGYDBgGyMjSFMD3Bdojzknf696s5EZnVJfWrWfM1DvHMfrerxgglALNRL
YWciRHwDsnb7lKAHbCPfxhYKbgvXroBQW+/OVRSzuojfgTuDNimPtIgqaHz2mZXD
aKPoAu3GoWBfb+5C4aad9rgvGtI9xwrz9pBsmwRdfcMUUAsL6vHnsdYjuOUCT/tZ
I0TX27kyXTCPnh+fMo+PC9txw0aIe/mXBR606diWgzG6fJfpNHFgJaIQl4JiYcS1
r9hVkxXvF9+pJDZBgH46G92DP2tWP5fsl/V91GqI7Ws=
`protect END_PROTECTED
