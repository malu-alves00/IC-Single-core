`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZpDVojg29sXa1zARPqo5SaL3zEQDGipy51ZU9yS0kJIY/hHUtuIgJ0ghUVaN1I6M
fZeY6CdRZE538uNov+Tuyc3tnQ0p8egi2MEROwWWIe/Y+e+qeaSVhuapHixm2URO
Y56eTNGBVHj3g0GxblgfUwEJo1MtPvOgF5PrDEHkgPpT8ruI34OozkRGHj9zjNFK
Fe1OEoDadSAjmQYmz1WPvFIBwt6PmOxhfl9TlIEKV5oDvpXS53lkaGyiWPZroMxf
TqfRuiVvfSE8HK3Cwr1MoukssvQWWKOSJdFNAXd70rIGmNmv9OB1neljKtmijGJ0
ePW07sZu2ydfuCgd6y7beVPnHLMFj5fpwoCzw34yP8lob3UdMipq4vQXQwvYtOm7
nul3JFWKb2ahDt5OB3QAs0yDfAVkuOn2bsT/SJxhDFoBb/Z4z/Pe3qksC3vkTkMV
VqhH73DEDnKQSPO5kiAuQiGE2cEmaFWlpoqcQ4/hJyYnMKC3guRGnl0f8zXDDQuy
eoKSTWriNcNU8i5Zfgc+8pPqjiyTvUnlNRbAP8Fac78/FNrDH2ubW9OD7Ug9fyEf
iISJXhAP3lSsN1XBW/ylwwOwA2GwX+DpeALuadOsX9zhjTgrrzvBadh8tC19iHe4
wzaolG2r8YVI0aCFw0N0t07howzXliSCL+v9Njd+hl/STU+ACQmdADifTYju/Ghm
n54RFuexny42u/UTcFGAJ98oGQdqdaxRY6/IPeHSHaCGZufCd2p5ttkO8BlG8LBa
2Pfon/RzBD0IQj7omSz+UOmVNZiBpZ1wjEtxcLUde+Uz93UeGpm7H5kGFoxUCFRS
vtJMYoF5YN6/QjO9DrGQNypaXttdyyzmK8jjj3R0bBDJZCNu49iKQ6K2jL8+H+iR
`protect END_PROTECTED
