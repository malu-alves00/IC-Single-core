`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bvhYguRg3cXRsH9OyjIOlQCTW5jOBErHiz9nqfvTDyPMTM/bRynj2kwXRVt1++r1
ehhlSs5WsC54CHbwPlJujmy4DDiiDWIZWueSgH7sdKxBCmy1LISY3+gp1YH7jf2O
bznsb0PZAcFG/RAzhmjJenz8EaAuXi1bI1D+ztPPcM2vHm1htdy/xlJOHNf/SA16
S7zyxhGFR11lc/onoYQR2VgFMoWDXFfymLg39TwiGa+YjM+zJdJsaXEEqdMHTLCr
lg8P+Oeh518WtY53a23ZclnTyvvp1Ubr/k6z9RYwOdKlD5HNY96Uk+jOJuRL8jsB
5GJd5YiSKpRdqHMKTq66zSnU0OlXp8vWChHJhdpKHJvDlQqVJgxxNOsNKoqOFP/S
aXaImDULSjOJ+NfA2y69fjSUf0MP1i4hnogI/3Hh1zqfNaetiH5uPq3ygVpQTgdY
qpst3BYYSWCWOyKwS4A6+qhHSpNUrXkemfwsFMsWBCUO27AMUjtMC+c6KFZJl6qT
l7Opc4FKUMjQUHgokesEpZV4gir4QblWv/sIhAYGIfPvvvVg2ilWzbce0xy8UdZF
xd+LjYNqdNa/Skivq0rhWn5tLEtcjputO1dDs8jmkLgwOsUC+K4ZMQwkbzMRvVyv
nuoRqSyvSeVwjmX6jZ7w/anh3wV334FHn+y/FGV2cC99tDYrZfzyR+UWKA1qjF/n
P0oFZacqlQeBPMbBQHkvmFDOm23q6XIMPGMvSX/cVQz+/VIfFEAGSdKiUMNis0Ng
g72KA3PIhFSVIlhI8VWaPTVlrmRPsveym3fAdYp4pIZfUn1E8phH7T7oCM3Rc76p
HtEVAh2pkpWcXz9gnzUPOK+qBJ7OD1VRaLC0MOCbxnO27GuZ37I7Xe3x8oZGSBZG
udkNYuWHfDceyTow/MGimnE+086zG/AnB77WBW171tXZZbNUeqxgbx79vyd74R0X
CPXKD26phQnq9d+Mh22hpj3cnrsoymwRwS79FownVyVfNPyig8GRCpuugsym+eOV
Mha81l/lFafSN2vGe0l1KZCSW9nnhAyohpUUPeBOJIijwJgQQpDGtmPpFEmD2gUj
Is+FtY+XonfZ5d3/mvxGfMM+eyFck/G2FdiCVdQG6d+ip42FSYN0Mex1EOTzZMcR
yHia5Lx8Sh7XSlmj/55pNaxHbssu8aQtxfbOObbwiY+J2Q3YYPXDpA3gvbPFDfpk
FEqGdVU/rkcs2qPa+t2qrXRBQh28n3qedrwZ2xIzueKZe9PqFWDCr+y+kGjOgj2P
zyD2rNLTGJ2uRLl8GLhYjBjMrcSCQAjwGA+onZGbPD69MmmVSfhoqDw6pm8E8nhg
5Mg2i7nV/Ho/L0Ow2QsFqjug6jbq7OzPshbHE5fAE049pY7wo0yBNRvvWcNqUabb
8EWz03VYjMLHZ2s8pk/p0WrNh5qCupu8C3akiB5dWjMqP8xewcdKp/NLSgkmWg8/
x0Bn+J3YWg2ZVgLiTlLi+4nYgGQVMMfq4QkASrRnurYXxaL+5MYbpWqlkpdfJSxY
ToZAMvnIkc+ayVilYVkRymQ6vi9Hg2XzPtmxedDldQa+KynhOLgMKkpFD2eZWSyz
kiH+iHTdxtBShk5Rfg1LhINBh1meNnfUhkF104VLx2oBALGaaKYQM2GqxiYFrg8B
1+nnf7YEzmrjQ0QV6J2MbnClmgJVkzXtJf/Gg1CJdWdpL/hha09rIipYaM3NP2t9
5nbp+cKcaDpKgssrIHTwuahDJWNZ6MpsXTzGd1Y+ZS4/iaV3sSDPVgFSYLAvlIxQ
I1etUSU0EO8p0GfjFMzt1ObbD0wpeFiMnr369zCWPMzUI/haSVPGg8yw/rCvk3/N
r4T3ZnOo8uWI8k9+t4c644+GD9kHhEMuvvahuv+cXXeH2DjjTrsuE4NTtEVPksyy
Zm8ydp+mDw4Tb6B17Vg0SZhocWaC9M9uvxlswHV11djElNhCN8Lqdfn24T4jAVd0
t3To6e4HnEaBqbZHKDRz7n0rqqIHsan6gN1WX0Vz7iDtDYiEu5Sc/KJLpwMqjQXH
WS9ey4thIxozdHqkZwnDHLtnuQ+C6bC4cTO7EWQwtijPsJ4VSBwQupU2ezYUR2bT
S1PIwjII35eEAMaehwJaMxqlxuAREYBF9/2uSJxjr+Z7bsrzTq/8/RfpLmKGs9Fc
RoK1aZOhLoyukVlJEBm8mu2m/1RRdjGXEbihGr3sTwEPW5n/KrCLw6VQK77Zbkau
LjUpYSVNYYtHTQHuxhouYheHhJprm/73QF12Bb6CCmbyB1l4UjFLL+6/q3yEPSHX
6fnJjBQrphPoDtFoJ9T9W/697ZXoyyNSLC80arZRNmErNVXndZV1+eAPvOCliXq/
Sz9LwFO3hqq/S/d/HmM/IbqB/4vtENTDej8YH/cImeX0tGx3dopwNXXhGjz3XReA
Igj4vOffMbAHEhKIiD3Jf9dK/le2oD9cjA2TUm3J2faT+Vfwpuo13H0rVBoEGSPl
fS5gf94MqHrxynzNou4k2M9o0MKA1go9+wyGMsgeQztFNJPhruxA65aR1YKt04b4
bAtUXgF0T+avkNpMmoisFeaTjBecz/w7wHDPvbPu1LvTXUadOLqd5kSn1RUn753b
YlwuJOSxJhYeGoW29ku8Wn+jxRPikUHqYzxQfyFZAiTwgMIYQ5MDQzgbylsKlw+4
3foJwpjUMe4KLBLeTOfTlT1FDn5aNCpeR5nCtVE/JVoJ4Ch4ZZUTeDaqlX8Uiv5y
lReR17cco5g+q3e6g2Tok58xRb4pwyFIqutnFGXsIcEEJjIr34WjPUVz9Xzh95nU
5Oiq8NqPXX2zyBgFDeT39LaLyA0Wm9UwirRXlCX8e1N/HqOA43RNr0A4P7bhZ6u6
U2M19Z2wz/FKa8sz4qH8ymZdTMsX/HrjbN+GwrxTBO1Qju5GiXwbMecan2rqh4yP
oJJTgXlWM+v6TWzpBYz0qxTadTMSYp/YSLoyGIJIRFG1TtnI9ZWYXxDap+HJmYO1
wZCWa7H0toom8ewX+Q8WDTc4QdC5d6OB6sbFZxkCF2qUx8vRhZvcRWHrD80DW56q
ty4XGFrER5cvps26/Sloq6O14bdYghklfMfvSYLCibLriHyNdQ34ne93HPdm/gWS
TCwCS+SI82/r/B/yYYu3m+MNPEit/RdP82uGlShwa9NurcxObFpzZmCD2Ifau33J
Dy0EuNfN1lT9Y164v/8vlQ==
`protect END_PROTECTED
