`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vCV0Lkke4937xN3wRzbFbuL6Uh46rrUmhuQnTRR2R9ZOcV2WdGjoW1YC3ENzHyYC
hecDtJCVgwBYqIxvV0/vFgKIzO+tw4wY81Uf6EfNGuycWeqsuCM5B8gYvzhflMfA
uCv8YfPIihgomHXqx/OFballMrcCDPMcgGtk1aN+OFRCWu8PT7z2C2SUWX6l79aF
AMVhjGPQ/Xuin7dl29EuAYLABgdFPPd5ahZX80LZ9rjkuHz2mBR3KlAKNQc2AoZK
SSYsLJ1R04jbXk69/iKW3g3muWO0AxZzZA3OC+uCUdpGplb7wsRI+VwuWrWfrOQM
UN7hSRZrpFALh3TeVjHObDj4QWmuati3DqD9Yo1K5mLaVgomC4uNLg8mGhSdhUHF
tHNPrRdYyJ0rjohZ/QHqsJF86eik5ASIs53t/rlZxsGvwnijcSCaFQmw0OIui11+
Zl/o27nIZE/rJOMXKimh3y5mV//RxiQqLjeuM4dhUjuPBpSbfT56Q7DwHfOMwKFR
CWFhuEagFNugtacCrbVGjj40eM7VU2czM7klHxoW3fugueRBgVS7SlXn30gb0xWD
17vbTATYRdKyTrmB5idpGCaYf8J8N4MfpFYT/RuPHW9y2VUBDovo6EWttdY8XeXA
iSbVB2aA0gQiEL6ufs5AhZ1ZwGxKlWXJ5xn0lIM8qRk=
`protect END_PROTECTED
