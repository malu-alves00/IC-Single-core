`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NqoRddCzea2tORN5wSOw60vReNjWHdfbEE7+a3thmcjfRNGS/cJZHVnkaR9WFvpH
eyW0zw8oDl4a9R2QNOtyRQ7Ori2nAfWOLmxLtpnMkbQMVZdCiOsM0wtEnQWVEand
HFGsaX7o1mlXfRlVG3RGKiBZ6mCRJ2z8VvrT64bZRusmASo+W/4lMWBSYgGPX9gN
f+m7Xkwx1nHUXijqBiYjUJrOnXnLmyl63nw97v8mxO96ugoCYK5K1yc/8wvoSjSv
3cOQX4J0Kv7Hv2JTZSe0gGZP3vTsdXBKsZO8lHLYnrYG/SARTzCWsl+Lx76lBpYQ
T7XzTZxgi7l9vevcDkoDYHXqKZpUjSGBHuZzs9x/qO0v8qATxWusDL357RYj5/xE
i2hzCiZX9rXfK3rlJL2hNP6LVsX387oWqtyFEVWRtriFuWNqmVuBb7vMB37Yz5Ng
tiqhkVuF4ENmxI5o3yKjZHHZdjXd+HRgwP2BCboTr9y0JVFenezetCdOTHf1nc3D
T5pmNjnTm8PQoWazAKZs2otZ+YX7rhGkQJZX3nQ0HDompvpyx0mIH1CjFtK17bN4
gJlNNP/rvpXwfYTBO5suImFnTdDppi0ZSUxGqJJ0TddI2nrIYp/lj3BZKPODre+n
Zl6fPQYqXnhGQPTK2M9HtKNN/8RROSGHTXJkR9M/EzLrEGeKP1PLsCAgiGpfBWlx
jMEowOVho2bgl3FBofGnWckvCeYPCuNL1/Al4GzeLnb6qiFKqs/PSCbpfPyuBzZp
yOPpnA73ljW6UeTG5McwHx1+UIx37DudPxo1iJH4pzh08ii7ves5yG0VUOSMytCA
z1l5mv2xdeszyNx1VPiHZFbkTMZjjR2h9Mg1r9aihNW8bOegcm2a8iT1bq7h1qA7
cSHmh6yxIFm/MqFteTWXHRffjhqhSHTNh4XDdxjKTIgeC/wAQOl6hCgHV8upNhEH
kTDyzf/SKCc1uB12dAMw4JJiaY7qVHTbUQzfH7CnVUZqU0YHiCASpRJ3S9ZtIopQ
+8tVxhEKhZkk5ozLz0fJ6B04qwRbDVV7OYW8w5YqH6qt4eI4Ds/FBKSwzp/bdgin
b5x/QovnjqSJgq8udwjyyn5l7IMVD1D9aMTCi2QeJgWMz2P+h+/T3phc4zBMTrN5
7yMQHO+I37tDdvFU0qwqkQeecpD+1izma+i7kzmKSJxqXcIcktq05RXW7ml19DVH
J3yZ617b7+hhX4VBVFTdyL+zNhIv8vMJcd0FDF8/OBwxk0JSjMABr7TGIkXH9ouV
EiSetsZ2KzIiivi9u/0uq26jHIp689FhKb/XNT9aiFJAtqg4lBVGwKUaa4kP40ds
tOu7WwKklEwVWcTykkeprW1k4W0Tmsj1nN93kxKLn2Sh0wIiBTVdwcc5abA7h5Xn
PB9996tbrcgYVsdPVZE2WbRHR+csgAez/077LhPdulVLE/IWhfqoZHWdi5GKKnWp
IGLKvWQzkrpHmRmTboEUII1eClmKzEr4tR5BJ+LRtRZeLd8khat8laF0Weddk7Md
dLgtabq9gNj1EgxqM6iaCVI6Ub4iC1Q985UZvCWtytpHUSpWI5vzunZwNAvXCzQq
SvZ4vzUHMoPPixin1BpbR41mAo0cLQ63SpxfvyEQ/WIjeNc/ZdVBEdze6JnXrYXI
fUcweivTJpn9/WzEJJCBusR5JTgBe55bF6nKrzainrLabiQw9MMiJi6fEG3lhsbO
oMtf69PtTMElNBzsvgHb1VtEvoH48/4xM8ug1seav9yuuMIr7dkR0PFZOxO9RTsE
eLXWl4IEQ+x10SNpBxVYtUGIl70wy1ZmEeeD9+/ldHLiO7IVazLhrfh1C4WE2NHT
4K693po1rhqjU7F3BL6WgrntcK1ooOYdMKMr3MAxFferqI8Y7lbZmrI+RS/BEv2F
oETdIGeteeSbPFcZ/EPwZzPCmVnlmAxkS1mnWXqzBLAUd6GiEA0EYObvOvgE/ivc
/iMCIC6XGnHWhz5c0sZeVsqOuNb+R2sJZPNOOkcqMY1aCy6B8fn5BYi3ymyEExhR
vB5YwFHwOAezRu6mswqOzN8RbrDZ6WdwzJObsKSZ/P2XMDu9Uw76npbXhN1IahG7
9yeRJAxTsR5W0S8FMVUHkvmy6sxMEToXpbsbl9ADhB5FGh4T+Ux0oO8NEan1DPvI
cfr5oyRMepfba3aa7Js1TvThygPmaGWLU0DPYUZTMvmqsVtPQQs7cmI9KYcWrxwd
Gz5gwss43TMBnhbH4TFMn/HxEsObYMLrIEhq5W7e2tpo22f2nxJ4EDOFSxPbRSet
mB1aP8uaTl4/dc+EWyVoQfWlLbLVbQPVm9GdlSmu11ggmwm4pfnisbD+g2p4jMFt
++/wbi/mCty4h4JWI5Y6dc8423Tjq2BKgpIapT1KCsLwuTPJt7QUqX1h9c70Atif
+7sAJtQxX8mMfCDzY2WWb/ijQ+o7FEXXjq3UK1Pkbz0WRJSZd/PMK8fK3WcmLccs
S198e0tNZXGdZ1FMyPsdCOTdEOQ4wFlZcyLOgsavOCbHkS0VrauVlRRi0GEp/eh6
OmoRuAkDKoL7OgMLBT1mHG8Qqj6gAVwskuh40n+MiHZAiQVO5UqVDHNjdT3n1mTB
9V1s9Bjwkhee2vLmTD8+TXmXR4acsT1ZeX/6bCqSQHySkmPIwU/nJbGUEjzDtwcF
F4eaeRUYPqBt9756FpOzE96PSEBjPinUilXcRbhVQn/MkB2WI2E5Wvw7pKeXe9/8
HeiwdMu+riNvC+IM6xbbY7pgN+WWPAZZixdCwGVLP4uUUDCYKEdRrdnegsU9+MGM
aQU+1W6A1oIe+aBk78kCZK8FSBeYY+UPFMUNJNe3kk5OjdUF4yHwJ32LMzw524nx
wVOu+5KR/rAO3Kc/00tDhwup7gLhQUqgi9uPoA7Ib8x+EKbdIsZYhsDIWdkuoa9P
15v5AodScOte//siRnJ3f5XhXHk6SmOoc5T3wLhwUQ67OETvYiK9Y4ypL1wIKQtN
tPlBksrJdsSXgENj151jym0gc/pdzaRsS5TdYd4lxNtU917A8/s/x0Pt4VPpOyJI
RtYLtvPKP4Wn6cCdSUwyDG6NjYRoTW0OCb+FrcR8d7pJiOBQMBdIjHLVPWHjNgee
TAWRwtdnL5zxg4V+/qq2sOzOe0lD0eQWwnhjCGEWD4XL+Ol/MB5w9LXvMaVw3QN/
MdMOMmjOQRcR36mQz6bdqdY9Yt+MwUmN/503e09Qt5hXjyUQBMKXdGQTTiBi1U5S
VeTKCYIPL1kNTqS1Xp+TLkGS2nuZdZo7U1bWc8v76SRKDI8zn2oZOKZ9riPtG+2S
PNJDG9fQxx2D7td02SBsZ7swBU7WZyHAmXHsifY104lalPNepwcbV43UNyu8OHvs
ra8dGcrzK/vC6wqYDUqPT4DFmZfYhIIMryk2//oVMgg3MTGC/0smpxM0mnIBDm7W
/bpJz1B5fGfLP/bfkksDngEQ2/UKwiZtaCUE+6NUgnGAs94bcmqwjEthrZ6WRLEv
zX/VwydP5410O+obRVUbZ/8jbdleZBWe3R4p+Bed+x9rBM2Av8GNgz8yxYH/ISAy
oJruI2LS5s+WnMkogULOCcAp6QW9U9R+zrs4LOfTCBhqOxLZUBb7eh0DTBhMtTE2
Y4+8xSErvNqODqfhD843/Ut5hGsRLeR7HCVc8X28cqn3oesNXmAQoZH+vmP+bZIc
w72gfZAecyvaATHMueX7gFtnAWAfPtvANqbHIYhMkRev2hGOWxl1+ujaH2pa4cnx
BBmWiz+LNc7a0skuQ7ZV+7zbhjcw7DBI8IDc7idBZe8eccE9p42Oj2+9D0fA3wpw
MY5L3Anbl8MfrtR5eaRV9YXmJmIMoCE4ohzI6LgJ+24FsSEc4ryi8DWAnqEvHORW
Gx4D/kNrm1+QLYmELutTe91QpCNPAAyN5OS9nqvyAuQJzMUdyQ8OLVVi5A7WllMs
aH6uFVFTUStpfrU3VI7482SaZKFUIlFWIBTStnhaY8N3QQSuF2dHhA1+BRN3F4yE
NBCvkD1l/ljmUzaxol9xFoOt8ZEB8wLEd2rJvoJI0nfXj0G3E+MCgoqP6LXB3vQ3
0gXeAJeUMUJ4SFVWwdGJvTzI0d/P9BQmkawkbHmeP/gee8gSH9gNsTNCYS9UIp5+
Zx0BHAx+pRyy62a0agA7GOH2PJjr1DdMABY7URMXFnoze5UnGvg755CudaL71uRd
VvkYEsGIkmq0BPc703uvL7V1ByvCQL12LYy3Udu7f4kiNpwgorAb3Je+w2Na+R6g
HUxXlwguHQ7NTtreRNXDxL3qfphd44gYH69Hu6Y5+gUXZyx5mNqZOcTfgzTRazwn
U/3KsGvfuuqyzXiqWMowjWlDpyZcxHxRXA6cTYbjPECnYt2B5B6cwjNEoXoD4+wF
0FHSgmkGyfDnxO8eP8bxaW+Owe2TIqXnQ5lG4N0fidjf6zf2pIs2UaygZNbyvU+n
2YtBRTRim2by6VIOz0p9a/QgK9URCCMf7Uyzt0A8RZrQJmUmUKA14xuPvmt3JdLI
BnIHkpISVBj3my3LsMf7ahI2juYEOlxXlS3uttjLofyZI3PXWedmZGUXrxqlEi3Q
rWYd6ACkQY7kzko80cii54aBynqjwyC1OxzhMWLgceGXnuxsgjzuAHv7eNTmGVhS
b3HVojJ02TAE50LZtsvTwo9Fh5Fs3ij3272uNRO43kCGjasyAhD9RU9I2X1qXUp6
B7Dicff7qvgEdKOhFcRgR/PLPKWLIsbu61NH/FV6v6OVXl7OstOBFJLsvoTBGiGk
H3F1SGnryE+LaAs49WmO4qKWpBtXkjR3cIyyAbmBaCWX61UOhotHVJsTblubD6XG
XUVRXNoe1bfTuXLhSc9dpX/bFVkKOwaKM9dKn8+f7kwN+w+oC40j75jHF71y+JWC
SkB+K8Sa9BGwbIvBN9oYNRRcVbkFIcj+A7dnd6cTEJlpA9jLT4y5SYBSJBWMOPku
N8BRrt0gyC/2yq8FwaHDBBH/eASPpq3+TyXibcXbp+LvpKyZYN32R+PzKEnMv9IE
OAdEzNLOdWEakuAMaqUpUDUiFqw3Hwl9TQT79R1NFf8J/X0glgpiyCdwoNgd2r3G
JXQOhpW0yQOSNKlv78i0YrzJiA1oFrPgDu2UkPjOdlOUk2g4zc3m8ObEbxSqQblK
i/Nj42PfI6nsm0aLhxXE2GdaiYUkIXkHDVsEO4K4bkaOOCCPaVrytV6zUlKhBJry
tow8LD7BtiNW8sUNapEVbetz86Nmqtsri8Jrv3Z/R9lR8k8W/zTXAqm/vyc846+J
SnhEzDreXo82nmNLLiVbEgXXNzrL+RiTGi/YE18pPMm09UOEhYp9EpbncCPs/WQQ
9VtkNk74+WLIw0g4uxEzxc8Ydy3MRGW6piXp1QEDCIpy816H6VrgXT1UKa05vPoa
xVVEhYYe4WF6useHHxthWl35dTStrIqwM4YbNbJqJOXzPwzPPUOKpjnUXZY0Thph
5pSs52nD9kfc5m/39IruxJt0+ju2Ca//LPZ+JTpXpyvhvggcbbj5T2Sh5IxBQJRQ
vVGKSSmog9WOjDqqCyMhNIzYpcyjHx8GytLJulHqPHY0NVhx4Md5XgLzOXlI6UgK
yi6FtSTduTdu9WuZE7zHUIX6E71O+16dCDoZjrRdYHH8Foq2u1RJheoUmpwlLDoA
snG8bMgVIZFunRvcAwwNau2zt7LdH8NkQ/antPLyP/7/1pyeo6eCfOm33vkpkqOF
fyAv6SNOGlXnFHzfyyCHQT/NKspJhSXL3ZuJjd7VBiiMfjU1EOt5EkKjxvQ4raxQ
zGa3/NVvqRldQEVF9nlV+F7yVc6FW0OGFYGjkCNg5bS/C96cm99+K6GwkEiE/l3Q
IcupWeji5fwGDabpFu4u71i5Yj7mimEQs2qqjIUfrENG9B9mRQCkhn6XuKkiCHRG
ZmxSPwkU6wVcbKuPUWoYMMZyqPfTCPTeBY5x2fBiZy+dXSDW10YJFjA2j0inDAF2
iwD6Tn/5w6OlXRTln3wCnqJCvEz08ErC7OIDsyQqXOPq2aVDrIioO3+FT3tdLE7u
NDmBC6tvMk+9ACTDtcOwwfzuv6fVwaigIReDAyuD5TeXAUOaEG3FnWb7Ne638aEM
6DA6TF+u8zVQ149v+muPBuAXGNTTbrLoN2oXI5ABdr6n95u/G09I7NhNj0uo0pwP
fsERf2sWIOSL/Ai5GLb6OJkqWd3NQm9q4oMBd/a5hJRCrRSu4xJob/47tOu4HWSy
+gEoYYDCgE34DYep03CVQmOr8mZe+o1AfK/OF5engx1u6/Ygz40d8K2HCINsLhe0
WYt+fFQ3Q7yMZPjB+7UDrcVtMBkdAC7Esrf7NckoX5spXnGTO2mzg59PoC3MfE+/
xvr7epua8HsrVaRZE2yEcQqFBmA4QtmFVSx3IAjN/vkh5vTv08lz5bpBZ8b4nCCc
9lMrOVWVbPlqx4hSn8t8vbM0gWvU6/Bb13N1yGR1APAWFQgyF0/FtZojia7QhFef
qAet3JR1zmEGod4sNbwNMvUbgD+l+Qs1zAhi09e/+Koyqqq0jlchxUAG8bse+d0a
Lh28KUb+I0hC6Um9I2rQ7pDpJ6u0QxzuEtDcL60VFN1LBPR/2QIi4qarK3nH8j/B
0F1IrW0WXNE+O6Q9ab/9aPIPtnyz07na1h4qB/9bzNjy/qQeY9RiwKp7PeyiNFIM
+CH8Bu7nCA92mEjxVV2OqwJVGkdP+P4EAEqjZRxmpqP0upRqco36uXbHQd8KAtn0
ZtcUNYimfbbL6YNWslAFODD2fvbf7jcmRU6o0c8LYDK6Oput6X4Rdz0psMXFKH2d
x4Vke2a9WVGu4ZbvhtXMhLI/MUemXDzf2Va4/I8qsjBrhgyVeepS9cEBa2F8s27G
zujBK6Eo11TqaDyWozuHGazC9Ue4QCTLjCpa7Mm79hasO6ADfgD19YVmSpdtlBoU
e8KBY2mgqT28beTl/MrkCqNt/5lH+nvIWLhHl0lNQPp36tAP0/iKDSkOiyoPwziz
4apUHfLTIT++1A4Xd9N1WtkqBoY0ZBTuD0IsYWxLWNHhQCtJk0/BCpIUIzpUH4G/
e47KVUuLMJkBr6q9bMLAySnIOBSdtMy7cR0wI/CmHAZ+nXYsTUX9Wlo8ySpefyIG
mY3YCbiNeSGzIL205J1UwcAVGEESq05ak3x2ErYV36CpEpVK1euPazEaL/hWJE4D
ZHWfLEEuClxuEPs1i6OLeau6uy829Zo0/3WI29tkK9Z8dho8kY52ZYUEO0vrjVEw
4VmnnHG7ubbyBoRexUthtN1OcLdeJMm0zZnDukj2f4SJfHYIlG0Br+fK3mXk/hpm
8FVpzuv0jPNW2FsnGy4c3Tqf6MYJkIgb2+QpAhtUU6Q0rZsMpFRfFM60G0tl/1Bs
vMXchOGPHyrGUnmyxJGcLslqxaza1j3EDHNci59vsMBjX9XdGrgtL49qytxtdSsj
HM6zs5dUqxJjSnHcYqco9cEzv/mt4uPzmIhGmAKFLmSlfh5awlcPWtsQBxiCey5I
KT0OeBclmgSjn0cRQlfKExcl4qkC8zo+CtI0jXw+NNF0EsZzqPjPTffj8l8XzBbA
foHeFvGHMYCbKyFMdgjCyYYPAtVfEkNlCnKRuz8L+6NCqJ626FoFhyf/VMzufW8p
M5Uq29MvLRjX19wQyljM/2yFPranF5cEocC+wChXU35ulAqX8yF9YI2Y9HVDKzg3
p8513boNWR2/sD2Zlwr9sY7HyAAn32/rhXlRXSmAJD9kWVCYRMTO/ZmQrdmpvg+8
AsLTR0swXzkA15QU5Dq0U9XbsZbPprWL9spjvv9M61TdbbgOLah4xJf1w5qE5YWo
lc9EmfNAV9TwXDROizsRC2hf50eI7eyFdRmeE0zYutt2lHtvFrrn2FGiEgmEEJJD
wrmqmlZtJOxemlfAHp8JVJ/aJdjzzz8890TWUCeQknvsRC5rSvb6ClxpQzA1Nw78
Vst2tEyOR5kj+zXQG1JT/R7ucYZcR4qUd3OzC4H+Teae2w+WvTvfvIXO7Mx7OX2L
3cD9e1jQtAhUSzIsn3+fEVapxDOd3LS4IQ73tK1lKpGe3iNFFw1Iwt/wLAac34SZ
MGQ81Sy2KWTLDx+gMlYtjYNFcmHNLdLx1Ppo1CiX1TQyaHwsRa2HMo48tj75gCRm
84beXJEcrObvu/EfsSh5GOIPpA/+O++1nt7NRad1z/jlvPkw3d+E+xdO289qwOsl
CbCkPmdQpd7Q0vTq2iqtUqMWacHw75li9pKM8cpD60wWNZRPWMPUG7wCK5hQpOMz
+E2N5GWSFl4jQbSBLw6JtvaQy1srEB8s3ODIJ/+RpBpBUYlkBP4bhhdpBko96/HL
Jh9Wjzohqg++xDFAzRlEygan5kngCVVthN5N+qMHpcwVMyargftGPvmJtXAzAYVx
nuGT/5TZ2WD1tSrU4QTT9IkclzPZyzpC2FtA6GuOiPEjHB+1vcBY4GtZJmt8/fNE
4P/bFWMfd4tjKDKTswJDsVu0YIvKKM7OuxJW4bXwTlZVtUwQGwnPZo5Z6iaAfxrn
bG4mV4P33RM+55YFuZqPh42wzLIlnnGElfu2gjL8zbLuBsht4nl6L+oS4Xb1hb1V
yv9FoWFsGYnLeckegRYjJSRD9jCQm/f209kumEA24Bm9EW0pG5rKXck+7+KtUUTs
QDabIWCluCGHKV2pNefsyOjVERBullpfUgqHajtBXcO8KJMW73tkyk1N4qbXWYmC
70hji2vLcm2WZm7o5Kk93oGc14LlOWUcEPXSlyMOzyD65PyeBPsCsQpS6WOdp9JE
mKyJMRVSHsKe5KmXy6w+ENBMw2DuFKc1koT2qdt4l+1tW36Esc7OXCs6CONX9Y47
Pqe2oz3nI3YgoYNPjgO/CvOr7X+tut5YSpZDZ9HMrx/XMjv8y9aQYPmkos+5ZL4Z
Cr0vCTpk6GE+j88K036yBNd/gsMhpewWNYcmWxwHfDSMZa1aHHFUDZ920/SEV5j6
z/URh3r9t25I/HwXqUKC6ORD1Js1LLvC7pN2GX6+wp0BHjkadm+TvmoHRHGM67Ts
UyX1JKq178fU5MfDscUDI4czXleQONwS3rn6HGSPcykhtjLDpjgFBF61YQnL2Aoz
8V5max4M3fnZRs04GQTiYYCSfF3SlkEO6uIXxBzrI3cfsHoqhOeHfr0++fClpwe0
sGyz716WJ70UkPRFZ7a8mpLjzyCqU4P9OTWcq8ZEQ50V4c/p9KZxAdIWThDeJbpE
4cVfQvDMywAuH7Q0twd3ZE2OA6+FNA9zI896T1DMJv8UUlFobe12It205EcD4tTW
ujb750H1EWdj/WBJA1xHfYXqppYq7ZHz7zIbRDPu+WvAdRZ++oVj/1qayjVQ9sOm
Egz+4aO87ZGb0E6YpJYFHL3tc+o8P1X2B9wquihGJezdUdycO1uTmfceBb5plENo
omPdrHmy67U3HRrduQTegsizpspUH8AsB/LM1G+2wQH8s8LKPH0WKCPHowQ47oSE
68GHVUwvAn2+1KmEF3mzCBEsBZVnol1qZ73AceyNNtlgXqmzxyc+hoZ2ruKsFI0G
bOfNWln+LWGCLzjUoKA2AUF82UthgADaTeA4iKITYm186MSAALSmcLccERa3/XAr
KfZ2mTqLAnwgtI442KZl+gMdZlCnWEkBlIAlxAGtsh+1I7bJbH2EfwZ7V1dheCmO
Vj58lU0nWsNK6bMg0JTIolISaVHCUs4DJEXm2hXv4eq4gchIMq+QOIF59sbj2wl4
kRFl4Or58LtBKawChlJsKjrqM2VDzJtlZnDDO9GfJshHMh3uD0vIfnG7e1fnQ/9j
c32+exIUHQmRUHAWJ0uZEqHd6sGl1sfIPG0p+tEich1iQlgpQl6dXK3WqjVxnWuq
oF1sAkr7z8qQh8U6QwXN6Zg7sMgMFvKtB0bCMCE1hZV1LiXQ9hYwkp1D1EoEoksF
p86QuIa32ooh2NQqbJmZhgJo48U2BJwRr+v3p0ddUT9lgelji/lp5K+2W0ek4vgF
m2wRewMvmfcxK4JYtAGCyZWN8XXvlM2d1SxnwMHroI8LuJUepnCd4Iz3dT6bVM0G
XUyfzQDHD9Y0hYI8iI0dON+frxajtOMcD2r/Tl6o1u5lQpgO9riF403n+kyeUnUK
SquLDDsKNNeJb3I63N+CBNXXdKKJBiNxovxuBJ6j6kzUNnMNjaK/DhxiGgZqpLJW
ekvN8JZ8RL5GNDVhWieKEVc5bK7UeMo9tI06AJHvNqMw9DoIJj/E248aXn4G0ORf
DamD7KqRv2OgNxv6LgqsY2eUi+oIE7dw1kWPpo8izPhxgeJYmCWAOrmQuXMTIVO7
/n0rhw9Ul3T3de5CYuIPKjkOkmAKMsvVA4cO2wGNAxmkbOgSdX5HdISABcdCrFkl
o5I8Co0Isf0fR3pFs+tprjXiblWXLw3ILfvJirPHrTuT1oWEm13j1BYIGa097S3n
wYnLgVn8v4UGu7E22XW1HR4NjPIYcCQfWPXaSLNvHnfWDMJl3yeBJXBrjk4NaRCY
dGdHn8jVhpk/vohNyuzp2R+URwjx3pTTWYBws1QBoTdAmhBStFVnsXSPnMbb/8FO
7uCQPQf1cX39IF4scOl3eQ7gP9ZnmObpAzz3pBaKqyaxFoQIjP2R8QSbrXWHh05+
JnkFEojABEYZwrAPLOr59AyhdijvbqFEZpa3+4F6G+UO2VODGJMvzaUiJfOrlB8j
njbkdXrDNz+c9G0iFJDa314Dee454FqfR96bmziwkj8bziMZN6X89GkhPamaD2R+
Y2u6nUZXP8YlbimXZcSsUVkQIqpGO4OdPB8dh8jGdjdJCtyCNQX7SudjL2ws92Fl
BJV5bUAMlho727lx91vT9lvgi3WGYw/6wRzk4OTPwBx5C003bNuK2fyHkV4vzHIr
R6/FI4111+esW9atbYWD4zFNtL+g0RyFD4nts69BdNsRes2ICmmTZESFfv59fUIC
WzwcRM3VIVMLFWda3/uhq+vz2MlmDQp2Dpwpdj2IGPjl5/4HJfiRwZKmojR6APTo
VNP6FajwmVnqs+1e809cPmYbzn9sS2+2uC6AQpHSxBZjip308AnrLymS3wq33j0Y
XxFlXEAxJzjAb8OwUpqQgRxWI7FahtahMIDVEGvBGySbctOwN1Hr72qT+r7khikj
jaf0r6vZ3dJzwEqx8plObNAVw2l6qQ16OTQlo0FABCN+IpeM7t50klRdPC+/EgiT
SZwLjpTsWkMb8syrRj376eB3/dB/eEdJ2AYnrJ778C2y8UYlZmrAtxFhXp/1WB4q
PQZDNwzsqktW5t0vkvom+zkSHPaRTBoajLlhUcKdGDi6DjIYtfzmzLo2glxuNAO5
tF19WHhwCtLlqD6SgLTtDaApGGDvnOnMJddrGO/abj5vk22ggEY+Aql4sp+qXZ3K
RN78e5DA/Ihxq2Z8TrbU3idMmZQCObbWfQnOu2fI2C6D1sNomimqlavIjKqabrI/
si+bnR5IleqQbq6Wir1gxNqxhvohj33vkN+jlCzBbX5nOQcOzz4+9fNQKjxGo0u5
670RR8LXhEWU+o0kzgNwvzMsWhvvZ6EiRHsKsJf27Mdt4J1gNFTzpJmn4z4nZwmi
uipkyJ2KNMPPGIlqKWxee+Teip51PcNrePhCBdQk+pVHcD6hi562f30KN+lQsUvg
0bx5YGC1LwRV5rZdKIzuLgoXXD2ML0CCwngIPgkv+gHrKq7bINiCPH56CcNQvPx+
vr9ETbjkVEnPSCXlhTekkcg/jtk2KdSpx3WuRl6tc5+yiqVGDUElRaL7xkwovW7M
g9PiyVpxzP0TFClcMMfwx8wxFmVe5bDpGOTMIp4WlZMwQksCuFtPI1tWR7b/8bJW
lV57SNfO+aXoyvMaBZbmIsk6MgYiMvalhKwFw+GGQDIeJr09nn/HBjkcWa8Ul2os
VOJaYuVguqYiiOz7Vfd9JlPoGbLar7A4+TENytFc32PhaqMtCnA5qFx8ASguoSbY
+fhjfFs9UxKwAuXAOiTq7uzKPua0eEO4U1GgEYrXLRhWkObmSd/Po06ON7xqPpgR
ey395Pp3/INiGjzHFN5uNApqNykW5SafnHlphOLSbrrI1k1GOGFYoob8njAWD4O2
2CQs3LxEGRylsYE9AhHk0vaSCEfU8rRQsa99odzF1UF5WwkawpOVVD8A16H53KSY
RFHXU2AlRw3TPCdp4N9NV6iiPskxvy/cSz3uHkVcHmEM4KcHMWBwc9PwpHWsUfgC
dmWnITGtMKWV47TjnaHUnLsnXfwCyaAgKoS9gIPtDSSU4Z24TvPMV4vKejqY2n6r
VK8l2hYwd2D6mW1ZhI7ImfkD1S8Waj2p9Wrr7yW9eyCEEfx4+C/BwmgUkDu8cBj2
a88CFW1IEAVDS0mlLgYinqtL2DwL9b90yjPbNly6ihqOsAT5vfLbjEvM4mFH0p/K
CBjZcCGx0uJZ4DVBN59Q1eYt9ohOoVUunCPI/DJ7liC7YDVcbkFp44SJxb7Rb+90
KMVf+2fNB0aLVoRzf466QQKdWgmnyDftbsswgVWeKUGGlGc3yVbG7rdAYG27zevc
3ihmyNqZBL6cRX/Khe0jNTjE4KOmJgs900e+ukRpmtwMfAH8d3NZSfQguj5VRnMD
bc5ZrxUqFO/xHfnSsNuJIolesW2qtKH/zAahUzjafVXNqHQU/ka7mj5mIg675ShE
LlifvvRb/HrJS3823M2cbahzpZfx2p0xX0GqMuZ3qfzcm4ex1Ge3xfxZyQm0WzPD
6t61KV3B8J9genfhew4nq8IyrpWVoDiaJdMVUaTePJjTWpFaqo1hEJ4F2or/rnOS
6jixwS7btpYQSafZm1nDcIeWprf4l5mLzI1EkO4eNvxBeL4fOHC0mKdXqucQuggU
p+Qn5n0w7IznLWCM1KFyozHGs6fnzEuSxvSfrJM4jsrQDoNQUgbSGwR9iS/+A5f9
P/4IoQZTgxv86nYP2DG1+WbP/XwWm5Ol+fVggkrnt01pqYQA/fYEJBj55qyJJ0hj
OKSvz9FpXdGpca259ubZtYayb0nBF7XPTzOcEfnTyvii/EnwqFEOBbd5Vo1nolTY
qUkfY31Zgn53irAmlLG7n+/N07+lqBHbJHPk/EfXBUHCZmAITG09K5CIWfd3lpdV
jsjmAWCqcaNGGF3YrEwGAPlNujXvRAGgBdC3CDqmVW2S98n9/3yowUfr3L8ORt+3
afXeHwh62GycHURYsSa9wowpwMGcOj2Kirs2RtkZZ3UsbkPpb4BketvTTjy1VLim
FnT+OVs+BF40tcqMcMvq1tHfdxny9S2Kx8g1ceM4TM9OVciZ1C+6Yzb4pdVeTE16
xqoTLDXp9TR/S9OlEAMeAMW6PFjHIT0xQVdYRPMy3QyjWHnUdl9aSkl+dqbhxm2l
kl3EPjqAPFD8P3UagBGzxBmVbBiMH6dCt/uDAEqNtvLtgZaCjR1c/dP+OSyzJXeE
TpgJ3HBpQ9VODRMoG5dsBc95Pp+/sA3MdaMHocxpAL/kDh+TJl1jerYc6FXhYAqy
1XYq5mmBoWqQmhTxyrsEADludKv8pNgiu1awPjq+0rxryKJ48Z8MY7ITyarSA+Fp
lin8OTor4UEYRGXkv7Zr0SvLhkb/u5ze2uADxksAK1XvotwS2Jh90fxX13Qmy0bH
zVN45e+USOuyRSLEI8L3/ggHHRAVYpSlo4Ljg3fQpqZLlkcLLi3eCH6aaIfDq9uP
PeU95U15OL7KJgX7ddzKyZTAFG9OwlUqOvTKQY69MxE6mc7Mm6qh/xxwftaaGzvQ
+J7KKg2CiNVmAejFJ3WC+FCnK8oE3uJS68zX39y0iMPO9Bt46LzEwCHxB4I2Ah+A
kYYInLCxbUKFmk0A0wC0XTmyip9L2+t2l9nKwfIAe80yleN7w/iZwCwUH5z9ac/P
3xxtDBOgvn46W8zUFOmrUnFsazCIU36g/GxPlot+iMVkKZ76vUqUyPRyro6vrUaM
MwmXJKzO145GNjP7VvlsSCAuX1tWOeyFnV9Acsh+nMaHX5KAUlIqMuiT5NgJa7ro
V+3Hgs4xE9eADW/AFHeebUV5SEW5FoWy42TPkJ2je2WrHXGVigEVLwwym3zSJRrx
Obb9PtO1MBOpPnJLSdOwBbAKKhHhxt22Q0IT84E6XcrjoUAivwuO2gySCxSfc10O
/XrGg6SaO0mJmmau1IBGfG/WuAl5R0J+4TSLGGu0VF8VfHW9bb6vQpW2F6Fqx9ZU
aBI2jT0yhpV/aID6ddjmQ9HPBLAUuIdql8LmCwIs7ncukbyTRULX3rLfOflTDi/m
BU+HuIZ1zpfBdpQVyB6h9Jq/9R4GmBDJQJukz89weCFz/rS2UWReI/OePvszLuKX
pA6lppUin5eX8bgiN+ui2qs3B5WRXm6qitefqH3XvpM9f72s6665kO8Nt8A2/RUv
biBEQKbJcW+QcMrer7PenqTRLi1Z6BWBzsC2NAoCnXe9aaEIzEZ2mnK0ZmARtXFa
7vIXsYWHS8nL75uINN4tEOd7OawGUtaFkoRWEUHxiicrMC2i18brJk3CXxgV7NlZ
tRhmJLTjdy4I+tE0jyvUm+nQApRBAzqCySRjo4kM5hIRnqPJUzW4UZ7//oGt2AT2
DWRADWDLOAd2U4yAE3LYwaCE/BcF4YL0O+JqjlbY+DiBPMCJhsqY16v5lZx3gppH
pYQNwglDTN1Shuk2sZzrMkXfN7XLiMruFxUCr1QMWvcvOgt6vGNymfcqFcY8CdoX
4+OaoDTqkYkNhszwxAQJVg1926Re2WW9rbxff0TR3hbTdWNQaJWWIt0Npc+hBMAK
0Y3QVCLZRLJJiU3ouUdEH9hNM3P9vagxutefpJPeHI4daSaLqFai9yznO103Ehla
tQ95UoU2MLULgctDaXCTwFfL7uX2fkQkfLa4+J4xi9rkpYGg28yJVR/+ZosPP8Hg
rPsq8/aEUsJ9mLuD+CeKMnDpx3VepapQXRRjE5xRcQRDe7tWsAGQgTmIbVpXYkjb
d9cQIvcj4WA++G5j4kSKbh5kCxrkmeVWw0CWME9hooXYwU8mf+rXpqGoDS14xYC+
W5kWevZ+veFW8IvCR/aYhrHaqB0lsSHc5gs/K/2/jgWGnZ/s4mROUc1ce0Pe1dO5
NGkZZ6npxg2sLyiG5Zq84ftLF/K3S2DICshmgd3IWpHQorRkrnvvZXlOAp/sOeRi
/flSMU7LyiQZwGVmAGJQVnnq/qoG1a9/JEm2J80ZwB+ChUDunwQkKlBCrweGZwWE
bE7w6NvQXNjPBdZblVQhvhctbeE+IkXOLOFc4G7rnf9XgcY9SnNGQ+CV6Umm+ekQ
21hAfdiSqH5u9GnbZDMmJbDJD2Zr2sDqodDetbH5Bbx9I0DJY8M/dEyg/xSDop3Q
FmCga+dmnwVjwt0rynTCz4gML09Qn4My5O6wcMeYktQy8iBfc0XDcYiZqDwPpbPR
fwcMZP7GbhDEtpthlDGJdJpmh5wVqSrohvou6VN6NaL2e4rrPujlxcsuPYSXCE+Y
RiM6lhn3hZ0IHL0fb8WYj2PAKCfqR9IfLBL11Wy8j9l2ffwkp6T6v5ue4yT0t75p
hxIjVkWxZJl3bIDIGMiqRTGauL8DJxhNTDPhyDAkiY6h1uS6ZKa9G2tJMCZBYgbw
jtyFjOGxdnfZjXKCfWkLJlmQpadktII/kTY5OnWtVkWolIqGe8hwXgVflOLV54+d
6K5fHYHFHdo0lVeXsyzLbyszDjd+CJcnjESDjcklgwO0Zla6rPuY0oR8eVW17mnK
HPQNJRbkWTYd6eGZvMKjUqwF3yw71bFVrMC8k9UBpNB5niFDG4bO3VKRoFmj5l1z
q+8tG42dL8AldvAe0qj+KP4ZarJ6PaoTyeLytDQI2dKNMzuNlKPnhAD6vN07RUbr
7xIjO0F2pLKNgNK03lZSYM82+qIJ21xiARSMb/0gyIKOX0tIxrCAHt7Zu1kbYWwV
WQx9XcH01VsbDP2QjkHnpqi+bMIp0CZY8/TLU/7w1mTEA9Hp1IV2xYvjWC15CRdk
Rb1aLyDcxyrxcveXDT6BBk8tOiwtZs8R2KiU0UQ3r1fwCkfmVT3ywiyF3kzO4o2z
Y5MGQyZDeRhYzPSIZZgbNn7tHtXDiriS5+koBqMXGpIEbVfeFgaQQuJP5Pobx/+n
DBbbMb0K9Vz18mCZpKXoLW2d+23rhD7v1WDwpAHfA6qt7E+wuaNdNi7FZvUGYBOP
S4/k1KEgjwlHkquogQ8cV7JqX7Rze/1oBilekfav/gXV3esRMCxCIVMJ+n22wREH
QZyEorbl+n3gK7ior3YqoW4vrhG4TyU7OqANZbiO5fyE7TVTIi6tAZFTFZiRyCTN
6shJyTbZjWZ/urO/fM4dt445IIcF/BOd0VTkbF1cWCoxU9K0VrOXX8Qj8cb6vUYp
9IX2j99YPcOVLOT5it2b4GuC+XtJ+10mFGieR3jueyaWDeDNoOz3gddYjggyPexY
GEpo7pre2VzPuQBjUT8T7BbDnJAQu3PTV2+axW6eYfR5jnlQ9IP5awst+9/GDIFi
F7lzY+T6DXUGf+ZxKDMDInlQp6WdOXVTvwBD7DbG2e2dF5rMqGAN2CcTOA41XOS1
nyG5Uy32IQSEcZNb4p1K8zCeNMeNj3+gCKAdNolJSiSlNvESc8OmF346dQk+0/aK
YN881O6bZ1mmZL4+FbsOHRwai6lyPc0EUwewEK3tZ5eLw+F4fjFTdq04sJFFl+an
qmQSmS6f67mRBabyF2k4oIQj0SDMpMmxCarWXIVDVDkf9cNqll7r3bL7NsioWBzj
5FLQgvxn/IaH2ByVmaVFNcWTuUlwOXLTNH+RUNSsXoSPTigfFsqv4effaGnDYb4s
U3hixHpe/3lL9V5Y2cMphhIUuBvB5Bn6FNt4fdSFJ/2yb6+RW96VOmzFNaHuRnmd
Wk7MRvQolSwjRN80kR/Newz8SLo53kYMDlK08XcNhwlq7mLBqtLO8DWAyUC7+aBE
f6YvfY930+0lHF+Lk6m6XQJqb9RbcBi/b46NiGekeskTdXuewvQuzE4mvQn8K8mU
BslnsKFQrGkU75gtk+2o81tLxIsrPKVpGw7AihIl1SRMRP4noOfFZ+jnpwdJzvii
3/mcBX9wJJSaS7w6OLFaS9do+IGo3xCl9WXbivf8cYHAjkFUWOPkjnLwyVSofifF
qd/ObJTTExzYshvHueh9AIULL6/6LeonVtslwO503W/Lcd/ilDqy+JVBC0o+OPJa
yeU/ku4g0fNMa8b5QSTYeQY2+NGu2Z132O3A4+bLC2tEf9MhYsNCcluL2IA9Z1mD
Set9/jiIj8a7Pp7v2pXYMTkGliR1Z6H8HRn3E+nSStR6WV49ZGZ4oKVvMT2bOaXL
uGr8O8EXT26xCO82XoAKn+TJDc8N+D5Ny/ZdJ7zWlKMqQ9q+kSPt1FM6a/dpHXNM
F9dfNHzET6xtzt2f0t+FuN7SjmMxrL+ixIIWDUTaSdEJQfW/be1vL9SyyBq9QNGz
LIsjpcXijYlEKZS1pePacxUqOizN7v7rnNFqudomlhvrKZDkb6o7bHFOzRRN7qFY
PCIZFBVk09ycMRs8YizPI0KUFwXCRqbBFtOp9aD+BAyHJyRmuYcKe4S47qoeAJdR
KSWh+TNi78Yw3RuZJQ07D9RY4wP7cgjy0xyJz4pY7vpQgHHNesIhzXaKD+a4cauO
tRuj42D5atVzYbRgPVzK3EBYsX0CDHtM09zVjImUgAFmOTPeIbOndbZ/5ampZcGS
xrm6+sV7yFvf+UwyRdCq8lZpaALUZMBYxfdg9tuqi5/B4xEIKfF1yIlsrJ68IPnx
KJYr5IglQYKJA5D61FdIMDznnovvS06LRXzDXZyCvpQmYVMBmTI9gREd0+NgoEla
IcibTIm0eKnmYprXkNBsBoKrhftmOIOtowBHrcMQeNv18zhiz+XlE0AEdI4KCBd4
RR5Ogr3zeQpXrJKOy/N1FQwd80YT9l3kqrsD7zi79t4m2rCX3f8w4v+5PUWnCUtm
5WRpsQ+vNIkrizJxVR04qIoZxjxbjwB/Vm4jKwcIyRjCmaiWVWeQa7BkgtzKg7E7
TiUcwcWqP8dpeziKYPFQlTViFIfYLc6bay/hCRc5WwbLNNKdx52jQhfrXongzeBn
XQ3g3bfhZ77S/Z8pzPKBUTWhOgsyKgdFx0yn6ekMvan+C0QpP0pmbNZpWN+BebD7
2wRUpSZA5JghEi2AS8UL+tISGTZHa78gvmlBeGHumng+2K3P4kJ0S6lTJUyP3PfL
C4PUbtoKAjPL120EWNj+x7Z73ajwjrUBsjHTDP7CIzd/F7Oan+v8nBCH49qmQiIJ
gFXWH2F/8ZK3xf35UaUW7wdlRWlgmqtLJBsM35M/xAgONHQAX5TsliE4uhUIMNYL
kgkTi6hQu//mHncAzhx3r9gSevwmdtNvLwf9LzNEHIkebXsrablI1izBZJnsP8kU
oda5j4t5okmAa8UNtRciJYjll1XzA1ueG354g2mYCnY4ta8s/lSGG8QPOZUByPlP
EfUdsr3h/PJWW4n7Y7reEXT+aDuE3vF3QXffDg286+Dp8WLbIsoPQlLxP2PccMms
a/8+5aCaYrP3mkrHuZhKO5/FzaQz79xh6Y7a1U78Pa2oJivfFLMrYE4sCGXyRDb6
C7l/EMcN4uI0cmr2XIP9OyPPxvW+vHkMAMYtgRcFfsMqc+a6mZ574ftlRNYJ+DI0
cMCRmklecTkNDkbl/hRKcSClsJrAm4nwE8tLt+Sp54d86RB+ntdE/R9/vh7q3UBD
gwM8hjVdpvkwO8p8S/sJqO/pwvFqeuj0CYMwbbUAzt+AbRFZsR7Tn7baW2FStBgy
HBiB2iRJjzix1VjsseeWQORg0Xyhc8WKt06LjxJ0ySYAHTGIjptmyLOk7J1P+dKk
vohyzjXMeMKjFpxQlO/12aDsGRAd9419opuOXCwAfIxByH6Swb90Zsg79eoijpI0
7z//VcCOQoRO8Phl8ITLDBD1ZGdxZl00TTq3KNx5Orq3LcD9EMM4p/JxCPSRAPUx
JexZiXsNSX0TutZRZ98IpUX7wyvbL22Z8+Z8be7LbLdgsjfvFX+1HWMYRqmb62MO
u/y5WIqjkGLebmVhTFcmR0+eEzBUqMwoD0PULPPpU/cwIwKwLoc2mzjeYPa2o3CT
LLwsfp1hm4302r8UA5MlMPKjPcwDUkAbQ9SNEcNIxDxnlG4wxO5+BxbRXW4PX8P1
e2r3Mt6huMEr/eGGgHE049SeCQeNgKT1sVfHu3/4DeWI9dLaFndhJyp+Pgzc7Md0
h268MmQAZzE4crfDSWBmcS1ZCOqAutx7ex3iE5rtv34tgwQvkzJt6R3OWEduR+fc
tz7vQ47o9S99OGieZMx40HSS6Puna5tFOPNy0wPsdaIbODKhIy7ozArxQE/6LES5
Dy+wxFHJNTQ4uHE5CbAHOXp7lBnyp9lrnjEcyq75otbS6d5i3waLl2eJKcpfQdA1
0GDJGay6EmFwoeEqzJcIkFfdKk2G8TckmG3LglRThFBfVxGpEbMwxb7S0qiW09YV
ploWfkWy4Il8S154OAnbRsUyPHluSNacDZz5oea+86XQ8IIZ2lsoa7knX2F5mIxZ
GB+cWZW7IEAY6IRAYpspG//EpNw0Xkwz9CK08ucLmtUJIzTkVKUbVBYb25Ad1tOe
/XzBeNfERTxiSOrACzeWXbTGa8EEciAcHG5MT2SqJyMtWKUIEpUhl9I6tuEH6Ypp
zU1ABfA7tMW3opAfem47Ui6W3tjTQsjvi0KubhRmHFY60erd3onSrivqETFkAryI
fw4OvQu1j+FYRIqWUukoGJD8+7Z7aXhc/z5KtYzzzn0adCk8JMkmJQ4lD05AaxE/
q36AQHMvP46ZJp3EqVYvZZlFykXKO9RYK4Nb6vwkeT2Eg5va84MAsh8VeawuCvlV
bFGljOlHfPfqKBdtGOPG3kRdvpGZz0QfJ8kNjtMlHsrZbokbz1z7Hhr415Pd0n6l
/5PtgVJOCQgNlkVFJKV/rDDfvYJfxdvG3YgjCoQmMp83NT5bQWNcSkAzw4GgOG1N
noryXPZepo9cdzvjKPQ/Bef2cPiHBvw/RxBLC9sphWnp4QJwIvxitINHcpfg+xku
GwL1gO1LXotedkxvOdGxwn+k421t/fL5Rz/dE6XlcSze7qfLLkjgTS3YKAkpyORp
DUjbBY4HLgb+ksSF3EQof7XXiUY2WO1SiBT8FAytHiKdc1Hh7AWCLD5yui1TuffV
XEDlsUIQ722ZDCpkVBpcGpDPUr7TzOSbg2uq8Hr0BCj4THUuWGPsmZ4JZmOqOXBu
bqH6KIjBNF+kkfeoXaLiMTMplq267HxdakCepMa3Vtm26cbkqsUnVTruRHTpnwQg
9v5mTHY1338IgRR5Nb+2fY4irQxnbPiiEgT+jINmQzhkoxqcIebcKotnsmeQbzzq
KJwvQ8RsePg/qHP8C/ggF/pT2P4NCeadTctbgKBqrKTSTNefEqm++tBiORi8ejw1
ypdCPDM+TkRfUAUuk3BECLnzoPRsLIj950khq5QHa8qGer6xMNwTo1e9x4Uvx/M+
wX9PgbU7Do4zPbALnnamnp4pG8MJQYzrXeoNrulEq70dDoy4V7Y8cSzUS8LtKt1S
2egGwL7XkKMEJKWp3tvKfdfvRTO6Xl8FjJW5s0q4leLsrRzWXLEpRPaYmOSGpW5M
5K9xYln20BhMxyr8VVhFwCX89/r8buZC89dKRy7LNbXT6SX0s7WJWZa2FtwIV5jE
Cx5LCLyDcuBqhSSgouiRmhkPHbz2LakMxkS1uDBAcotKKcXfH4+WO4S0ymsIo8/2
Rj/kxZG2qPlxaxRo7E53pOyc4airFAfSbBxmRM/25sPqkpbWcGYktybkQI9k9Y21
m8hDj4oK5C4F67pcWjB9Ogox2oolCo9C7KdacgJR0qyPkrQSmZkbPCVb4buyKG1u
rF33UupYq1G5i30KQ1t48m8+2aqrRpzBGqHdynZGShFMFbDhpWoZbmPHpMENhkdL
n4jQwLPvn7BaZ3w0S5Jtpw4959eWGG74CRtlciRarYfy6QFeJMVu/mVPrDs1UCQr
kQ08Qn4avswYZBVaHY1W+SMpA2WK2+WmLmEApt/0ekHTmp+uEUIRYDxhgquumHHQ
XVK8Ki5GeSvC0hyZdFEuAk0ObwMNLL35KLOhMGvFhcf526zhhvoTG/rWyqXimcVd
79uaE7WdWzO3+atbeRAMaa43WLwRqLGrrRCBWyEN8X86WKRp6V2+8hGkzdQgfRXO
kzxK92KhP7QIptb28ijWz6pS2WHabWJdQneVtmWyRzoWf0UsCocxx4asxZXG+ewx
oQXwnFM3TfJrVXWAs0Jc2y+Vb1DdQQkyTelOFlPQ1cWVXJ/B39sXdDTowTE93+XR
huxfPJ3CeVszCFFq73ke8TSqVe6/MiUNxQw783nu8ADdUPW+V6QC8mt2uhNv2IFq
yGoDKICmD3IwZo2DaycbH+EoZQVkIjwsUlQPao5AhogJXM+oUgqtGjm826B7H9CW
66jHpmw6XoYYnu+xbfpXzUfE14NW7tmao1Vz0YQMnDANy8/UwfU8f696BFNlbLyT
2Z5AeHtwcywMbxtKBZhehEES8RCFYl0Aom9hh+7zxjEgDHdiUupNHvtn0J6v70EK
sy5hzFS57kPEjI0YJWSjZc351qHexF3pe+gQKgbgeigYq/VvwMNhiWc/dFOVB6ba
vxdq11kVvkjH3ADe0A7zzRD5nxhzSplOS32zAfDapZo0GFB7IPhpPNUefwolAe/p
UK4fotiz3k/Xw841PxDe2WPytRbSASBLjCc+25RUhLYAXxI6u2Ydc2yBRbV2CzHv
SVuV58rj52tytqIsR3+W/RYZhhkdWvFa/+RLt+SJGrQyoiusuh7wrebwqwIURggW
Sr2mSMKy1hjjJuLHVBstcGrlwszwpI/t5wcEfA+0qzaE8hUccwzwc97rDBnEAAVY
eThvkg328scPQmKr/rXAG/4FUy+cJqc4r8aijCA2IjlKAT8L8yeBPn4/+OsVyw+C
2r/cPld683ze0M+yWVmpj5Ddpg47aFPgI+ig/6eObTdoDtzocAlmTujK/2REfhC6
kFG/PxPYBUt8PdlyFqBH5QivQvo7KXqe8eEX4j+QqIX+ov0DV5b8kVHc4hcT1aXC
Ny1U2Ha3n+Z+IUTnnSo5BbFmSm89gXq914DI4wLjmSXdS6wXZEIeDbgcN7l5DuIP
mB3VQFv7mGC8kYq2HWqJDgoRk/YI77p0RatYIAruOWKn9WxZbBMHIrm7i7c/47R3
YxaSh4B2QFA0cWzIjdQ7oaku/4S3keikwFNjmOIVzRIZXO3IKv/WEuZB/fpih5Fv
HBWoBgCaE/b75728M6V0M+gX1mxGDrunBJ5YBGIDVF6rBFR+uzR3pyMmhLNGXWU1
LEbEpkz3yffjuzXhEBShee5PG5FsmwsIqK6fKNR3eAhw8kI4IPY3UHQpEa5h9dGm
HkYjVx1aWUe3L6ugHTFvO78KRxroy/kcZtHjCRMjpSQFaIWArBh64r6bGICK7pSo
p2iFyDjwaTO2A95uATyv8U4tS77777wrerwEfrhMd721Z+NrPHxG58Cc+INJGvHt
OQrY1CdYBOov65n+VkPFAp8A4Q0SUlcrjcBvYt5y5/GUiRihcW5Si1MBiTEWZ1yI
ygTEtl6F2kovqJTsPx/MK6Vr3lwOlE6QPjK14Hm9alH75qs1KECUYEWTi4qE59+L
HoLiTC+oxa1sycMYCSeLS8nkwDZmhMBcGfppab09C/60H6oiiJH94FfVgpxaUrxh
yRA2hZOiQbr2VQHoYQj858xKtXxU36A+wJxRXqHZRGEuwY3ZziWUbjUDC6ofG8BT
XWmctlI7k61/K0wyb0h7DERytkvKMPKQmwAOeZKakITr2T29YEsL7u9wD+L8EuJL
y0fbVPRU9qQqhczir9DkgCpEodCpdKEl/PShc3vD4L0Y+jsQp/UuzDtRHq+22BOp
/xx3SnAqjE/ZWsLyrldEL2EMT8MyjXbn7/xlvmZWLzPeZwDx/9/gYY2ZWkJW11BW
Twg3Z53cbo4QUh0wp1QVASvDrOPc96X7tVlAhxmnmqt3HVD4ifpMFX3AwJYWyNLH
MGYU5Swk5qgiP/ZIGW0ENE0oQpmUQuHQxHJi4DTLKvGaW0bkXQbGdak/uGtCWgUQ
b09i8p6R6NmqzVnGA/b/sXTu1E44J86bw1GxWvN+lNoP8HgDuIuG85NQm4F+zSyV
rAsk/9guk93dvCTxttiIaVVHtQ9z0KuF9Ca/Ntc6lU8gGGn6cT3fzjqtYuWYj2J4
HmMp7ggs2rfvHHDNucOfkaD95JM0G+xnmXKlJ/cWpatIMEA16hRHaMo5/O1OrGmQ
N0zT+InhZPMX1NAnsEJKLDtq589XTvkpIYkQ9OPJ6QshdlSzOWi5krkVjl9Iv7vA
lU28m6oGJmK78iR8+JcI1jdLCAVWKzx6sSsWT35SvkwPDpsk5QxZbX45Nkqui2HQ
1GGEJQgY7hny1Tcmk5unROfI76BQb0NGvtvk4j0DxWzgV8byUhblkwlfo93nUFvR
RooPMg2kncAxAUEGSoifcmAAjOULZ2pSDZKuOA9ASbDLik9qR8wcNhigKid2zsnW
3CMWF434qtv6lACG4qTRxAzub0cJcJF7fR1X++qxSxLAM5lxaKjtMUr9RC/6XSoi
KdepirQPmv8jLWBfUCDmPCIM95+C/d/5DNo9er+NZ6T+hhtIJPOB56PDK1GbdP8+
eoD8i2jGkyDuq1CC3EVUUbC6fC8bWDbGtdkf+umcDkrGsLlSiI3Luy/nOAHaQHrs
ehZI/Kq/TZbusud5XM2I8MfT2Aym9tO33DUEFxv9CQmZGslf6sW/jSEjGKwb5KOk
ulhuYMjwmHk5dU1MNGMswEYI2J5aKdNAzF2Ct9R+XfJkv+R5skVitok6gt18ti6P
ya3Yv3HCT1HEW0zDp5wKUboCKsScGXyiTXR8A1FjeHyT/NMo3otL8SUAtrcrePNp
pY2kgkF45GrFJi7onvrFMA0nsCSFoyd2WFXwj2KBD/Rqe4b6t+PlldAukR++f5dV
eR+7ozWGZs44AU3PUOIuaeMGA9L9uo9sJkq9D07T3atwX6V/16RS/rTTIuRtthFm
lIVupdZjCvBiFuHvDyVUmXZ/xv245AMkOfKNrwQAp80FP3ntoEg30PJNEPyTIfMz
VAkWqnMGispf+gDJH3RvxGYh4IC9Yom8CjcLoR5lCQFwT9xG9DQrQr6mMf8uS+dk
LZW8yC5WYp5TJXzQy8O63cUWLW5Vrrw9XBe4ZiLCu/5swy1wxBsRUaI4+KJLTMj+
LdWihUqpiqHnlZLVAfuuCUuwVI5+RadSk2wwWQGBKFXw7kQjfuMJHYexbHzIX+5h
4il4QfHgF6dvvFsfilzotUPHQJGy0JihKv7D1lqqazJ8B1L6+pPHXMulj0yCr/yC
o4pst9C4ieSqw+288NpsmAl5bfBcrTxIKMPu4LdfVWWvsFHrUvFD74lvWO0Yh7MU
MrRkKwde6NAnVdk6bkW/uDjziGCyN4GoZmFThpekgdD8zz0Q9R3DVgZhle4+UeYA
fzuEj5v4rSlCeJFqjC2M3Uq/FVupvXh3jKIIitHiQiSZ9ZwJXDqLYzzuv2RwKcuj
5CSSYaf5EslRvQt+lx0AJP9KA1dguJB7Vtfbuh1W7lXZ8QD9dA0+CK2iaY4WaVba
J6U5QqjTRDq5dno3tt6cKjHcyDKAiIY7e3fBG8t4Xhkj/ShhnXJ+mfIROx64HrA1
64sJzd7XhG2TZZTPAQHXnVX7/MQliyYZXgkdfp+n+GEC4Td+ynjqzp6qri73a75e
7BV2baJ5FisrTqhNJBa4TQr7iVgBxVRj8gNXAYRPsdnT2BokwXIt+lKGX5k2pzfC
S4/C47OTqvJnnhhdVmITUmP5SWb3QzIBtkR4RS7smrHQqL5gwu8Xxg3tYWR+9miu
+ShY9yGeJfzqpMEiD13W8DCsPLL0lKjB/ph2BjfcLtcT0VpRNyzG1j67b2YwB5RC
e3/6s5oJaGk3AkGi9cMSQhUKQoKkLSF0tALvZz+iLDJmsmb7zpO1GCIm/9vYYPZt
MIE6mX97/q0A3B+Ebj9cxwxKAxTXppTYrxPxuiVMbwlorm7SPae80MbrxDHfmJ6Y
DyGZ4rZMFQJUlDF9K2NR8CSO6VmvJG3TBVuxH/sH6ot4PH1FmPF9NfwVXRuBLOql
H9q+82syJfEQaPE0Gj9ylniIylsozn0IfmlqrpvFQxP0zlXuTdBhdBwvSZ6l5enB
aqfgMxnZCc1pGILMGr3S7GDrrflTcoptUN5uIF0mpVGQVTv+AiLlFcBxCQL5je2I
JeQTFfXDBO0AXKsC/P9Nn7Jyo4zcBnJWkizuzawbPPNNB0XIKupk8W4d4nnacSra
3yTqIP47RUTjLnsYHHYW7K3zW3ADOvTmcGnupM+WuHlsHPDqAXJL+ZtWwZ9UEKMZ
vCuWq8ts+6dQ3c/T7f1Qx0Syr7WO2hqAfv8rehLpnrZRfvSsLetqz3Mg+1gYLNxh
g+kDneVwN4wXxTKcsKNnk1BaqlcNBFIAEydggsldy60tL081s/Ra3ga/u3fzV31v
+V/DCEtrRiMr8hDKJ4AnVJ6+SITeykFO62tLCaE/87wJzh/gxjNVYdPajTuEQXUN
VTblngzBJ3n3OBHfcaTqxwbNdp2gp6z5iUfzRCz1EA8PP942CqOEZg3HFze53kMu
eSLF8KNx3ASsFUihk7dDa/8ifGviC+TFTpycERUL80opD0dG0ttkLM3+An7M1cSr
pX7UydpVVJuPH4SPbqDwokznR55KldCWJoQRTIJcDrxD2PKWenIcB6UrrPFsdkDf
XmhSe/SDe8Wo3E+E0b/lZfPgcJqVLWxKOiAdeSA3n8DIfkfhuBlYsnP46WTiBngK
EJd5UlQTRemhn3rFehSLMBcuwitoWOvV84Efaog8zS4vygxe6rPbFhtxT//osjIS
AEmwLgxSaLS7j+IifJgAshMSH0umSegpW4YXqXpwu1SmRqApYqXBOBtFU5nUaiCC
tUbkt5I8cm69OGmoRpL1BFD2XjpfN4Lcu9j3zsALu3j52yGjizZ+S2ZgZqNC1Zr5
6TYr9Xe4eLIfmCKZhpwquPalH1qEBMwWxxCh5rEr4QIIeR4pWur+k7MZDQpJd55L
h6GsDAKDpZR+fIBV0rmXkczRiSyDdI+l0Z4ISQX/u+Ydrwcy18UUxQIhW2fGkSn7
oRRMJpktWSE7obT4ksKzv7sotf/hUug69Xk34eYhxbLLwxWrI5yRV5wGir5W6Ro/
8d08jsOA4JzEbmznOoiSWlMGO7lRQ5BowrNYrxeQrEChQf+kVwMFHOEya7IpviO4
rxt+N1OODrBERZ/jhgwJzo64t2NWy9TIJGkPF0uCCiUS71yXJBhXhuTJoUn9OIdd
coUk1HHIT3Yl/Ke6QWH7TsDaCG846gVSso5LjsfM1N99FKt6IUQnvTrn/lKfrtD7
fX8w7xRTsWisB0LBX1tFgEaS68AAtwAuDNYCwniDN+XJRVHZ6ScKy07txMKMHiQv
Accy7/bfnuUdWsqFAy0nd+TY14+lY3Sphi2qvrQfoZ93xGi/YDUapVuFWNc2YRBC
B58RYWKhoWFsfohdPtfszRPakHYm421mBqCOWME36ZMtWaOCI4MB66nQYglu7N8t
Wuvh5yloBVz6iOrB6MEgIem6M/PWm0gGuYV/5VEemtNhvzzrbqBbv6kEzRgm0def
+xC94VmerjuFax2ljCkJtLLBlRfFqsExlGJDX+CnN14mg74VlDXFYx0xyvNEhPer
HtMV2cpQd2GvH62D4pkjLE3sezCh446gM2wYVnLq2SGtY8lEOXT5ts/Gdyr0H8SF
M9QsxVji8s463EXdPofEks5ZM30BfYmObstluTdRlDBVzFC1GfLP66XoNpvAnrLm
KzLG+uMIHL4mmDXDe5682A0whQ34NEQFlh+Oc4A0XSKLvP2wZalXeCLBhx5shHg6
fo3MxnFRfEHkKwtGd1xc61o5PJV25fZUjcdK84IaF7GbUUkGzNM6R9NdCpuzkDsj
FfNlKqVuXzTU/Ify95xW5Wsh7ei2s38InZ2DNEqn98QHEZ4Qe8fVSf5TLn4PXjpd
2mFpC8vJapwiFjm1EwVyosSd/SkgIavUfqMHwNTBE7LxKFz3tLcH58i+t7rcQOtK
pLQtaUAuKQHIAkLCBBoyNFi7kHJwi9TYGj0VEeLdr/iMpSVmgfw7ku/DDVRRwJM0
Qp0oW/ETOYpsDLFAn0uBWxzoFxATuNovr4cD4bBzNWTehESVFYLnzh1MO2BhB3l1
qs070Ayj7THNAj8cJu7LkMSzng5W9f7ZaQ+q3igQrioIripE4iULo0c/4R8ZgZPS
Vkc48D6vL6Aa4LBbfWIB54/BhYrmP3oPefVTjHRvjVKjeEr9jedqxmYf5QRmvNIS
Vb4YshyMG25gxKPhPdoQMswhpZC2HM7Kx0SRJhHruF8L/Srg1ZeY+sBK6YFzR/H1
RGS9samvtrLO230qUT5HUb9T9Yn05/gZO//gnAWuYcUdTM6nUKcbiPnqYdgCMiAB
++HkNCHgNnQIA4S9z3t/8ySB+7AP37i5OhrznhZnVIjNad+ORt/PPXFa0YRruCsh
MAi2EmuoSlJzBVKRr9iFe2BYs1NMbC7Y9CJh58IjKmsCMegPQFmW+bw3PoQRjQ4E
MdaYbpOcnuC2LVcqTfG/1IZj7WstlFqGkuROElCnF+2mEGda3xg0npk6RkQsyqK5
29ujAtLAVzcoi9tbv9E6qf8MYwepcUmH10nZvLUm+TFX9Uv1G2tdojgZ0YLHgqA5
XYy3LXLa/v4gKDIVrxCg+Q+E3etwYAC5Hvk1u+OgPUH9kDu14hGtO/VCJ0mKrsOk
Iu4/dA0cUyjtghcmfsddTs5PUwSBxrWzRWNOSCDllv1/ENfQS79vnQw+9kFEMkYW
kxYpKqePSxaZm4Lhra+D60hs1jn7H7A1LTsHmwHXeSQ1KJ6GEHP/VYjctkzaFqxU
wAoE6LupfMZD8HOOap/pUgoTCeedCpYdT1eGu/lF9+ZZcOC3mpCMjLpJDqBc+jcn
t1a9t91YM1qQDEyyTBezrcurPIdd8I+sWo5TbouRVOX1w+CyCxi+lEbjZHEh5IE2
lYxxTYTmcxk1djakGMDYw70rEU3OzGA8sEsNcOZ77TI2A58YjO+qF7c0VfjzG5/S
g58DVoXSMMLg8EN9t5QwN52WZjsKF5YgVGub2RuE8vnpd7TRtcsRHuHGW0+Da/JI
HsqTssSwOF22Zzr0HWuWnfWmgAF9EKKN65SIOEJwp6DIHk2LmWegp1uCip71W4p9
98sysTMaInd3g+SsY4TJjNC9waf8k/zvmle1yKWL0ZSQRTEeX7tMzh4h49wchgl5
vver9FVTVrr93LKnQP1Oei8iAOxBnaFwpoZcArfnDBuxcfeBdFzXf986vc+rTFUi
8E7kn+3Z/YENVDvRXiuE71pJVXS5CCze8BsRfYNAqVf+KxKmKKfaZYhwsv6my2kt
omAhzTX3NwMFwljXvYl+Hbw0UGt794yn0owSlXshxRd8Lu0HOyB2eI1vunOuiSes
Tp76chuC8cZ5Vbat5brVxxb2eeC2ADuNvwcau+LxFoDeDoXRW2heRCHVNoAgYIEK
Xus5w2siUjbKha3kkG9nJY43W3t3SJ2InPp1n3N86a20o4qXFqcDPDKGxJCTynug
Svy+SQSiRKrxxFWsYdlHA2jKC0E8wNVbuW9e7sN+zuxRA+B8ET06QhHQ8wlX194n
hUNDgTsKvOFQmwTQvGLndHO1LQlSAEHz/m7hjxAjUf6QaBREnYkbWMraRNgut00S
cdupcpCn+hkp8Wzq221Tu6p6CXqS6GZvZvDhPdUf+KCkemKwXuknUe/vgOeecn3c
rglzILbrDWutt/i7jvMqxE2hILmLy9x2wKlyOKmneSqwSWioixmxwFU/okl/BzYl
TGHh9BrBECH3vi+WJLa5nWSgU7oGOByTjUWlLsYKWcsC8sbESrnnOXyrBe+bHv/a
YGd0rlUyj3DfK0BlOe11p0LeSnX0muZFZNd9VMR75LjOsJRNPL0OT1gYuyLEKlwB
+tFSwAkB489RmX40ESkBeXlVbBVvQVFB0a6GWZ4YrOa+/nPa6GXz3zIBuq9//Lrq
fOcli0r1R6U6tY/8321F67z0lzB5rUJY65FdgFi8SeoJArhw8ARK9xHB5qILA2ra
2B24sAu/fgTlujMadQ0NGvoFzt8IcnLrlGdqwvW2Ozm9BTTQJ/ctAKS+SzeitN3G
GoJkP/PXyQMSxGLxQHmsix+zvZqjHhrK3tEky7fXvYCVE/vu7TEtThEzL6Dq8X2r
w95N/U4aPFZGpE5M5kgAlL8QeVnYR4Yh6CRDZTqR24nR7ay1x27nwBiTCAsdpML0
yicctlS/ylpZE7KoyxSp4qOzbhz9AOj2ySdFIxUcf1CTKMOU2P5AK523tJ5blhP4
XPqRdUPswQhKnOE3eZZlf4WmNHAyphR/biRpmCQdwKbilbtmuwuqCTawRxllhplg
Sx5CAPSRig4dhfaGUCW70Gt1tltX4im33vkmm5ZfuWdOtTmrZ0DjHvpyvUSgPuGg
WdTR2kqWhzm8fWV2wAhzd8/cgAwEUr2cw9S66Tg2Q8bLJDJpRsbJMewgbWjt8w4K
Lhjk0VmzvmxvRTHipk4y2UUnZvbla4wpjz3xLQZ+1SjzJItzq+ssJ92BkA84a5p9
EcRde4osLv2N+gs6xs9T2RHyv9PMHNy8nR0n0rxOqE5XNpxMHAjRst9k+JifLrIc
jfDUOrQG7nnzAsFlzE8AS7zPhzyQKJHTj0EXmVM5zAIDfPiZ4ASdFjhgsVHulRpo
TFLM2sgOohOFPbh/mYRBvhe55b/1guDW07/BVGvuUid1f1xA3CgNX4MnrSCqO9Tt
KjdppGF/QsR8PkFvDqaPGFeT8ei/UL0CXDtMCQgciyGPN34WyejNiD7OotFuQEuj
+3TRSTg322362IPyjJusiSblDaTyCuBLjEXwqGym5tsrVYd+LRraVuhWx/TYzHpV
/ftfssjpxFu2kG1TC5M1Un34z3S9QbKRn59gXnAn1Q0OKGzJZPu26e5KyQYf93Jp
fRMi4BhdldQrhWja8ENzV8U3+ifVJecVbSVMtrqUYtQOQoPp5QjbAqPS0wa1YeMv
1AdAzytsbksbo1v63rax8r40geEI7q11ScGFaMfPt+zFwNyHhV5z8twl+NlYBqw7
JSh4umU+qtVEqd4/M0MPU9utvCYvZA6xCJgIxwRsvohA8BTRhjC+bcNUVm4wu57y
6/ti1E1N9Pz1baeNP+HCWsHMMf/KNzxzjR466W/0+r1aInvpEHMVxGrCPpHr58Bj
jiC6gOatkwpM4thSfrf+OzLn2612Q2wiVuyETYxQM5NR6PKs4amonTt3e2u9n4/2
rp/il0/kn0UHrFRnK0GWxgEDrnaXH1viFO+agF+7LNR/PnMfWLtFao1PzBUJa0Gn
zOFdv5sOhEiT0OomYlv+DcqLZSsB8Vy3a3Eouw982/qAAcF52R9wC3x2tq+m56ql
9GSgjcNPmI3YcKQO0U9bksXFlhElyWsKoDYlLVcNUOLKFMdwFChHndUgqxgHYXLo
Sp6dHWIFH7Sq5Vf5C5J2ZT//onvQjJn9+Y297ykYwHVcQ0uc0mvs/cUcUzuQoJXn
wGn0kRlXqd88258vesphqZ2E+mxCxK52mL0+PriiuAiwG44ntiU3I5U1eZUOywA2
Fbk9nOsErEG2SFidNQCSB0GbZxBKqwD1wo50vdp/W1r5VpxvolBodvlzU7hViCXZ
r/YpBUywjQAxRrjK8EArihoEqpXS6Txpa1NfoMgwzoa6w480z9ABx52ft6lHPBz5
BUJOKI87RYeixqMLxjvuZbw0I7lCjN7sc9ZkI5EwvrgX6S9gw82PoooewDJpdSgU
lxexjapeDJq8sWdxP0Ts7c5OmsZY9nVAhI+yWiPNMrvKo+O8Cy+HQLj15OVG2sAE
8u8a3EImO7w9//A5k2ncRUl0DShlMt4feQl2v8NbYmTzNIn4wvbzgFE6riSc1hew
0y8WpXK5qvzS5muAVhQAlbLyOcba1uZd/rA3C7wEQG03TIKbmUjLFTiQnHDPJEB8
wb0cMsHH6Wa5ctLpRZLyPLxhJ7ISIQFPGFOta3d3RmPvObKwIvFkpmvQA8VjkhUu
BMp8ooG6tFCti1vIJ+f0fTMH/1Rhe2Y0j+7nWBXrk2lvbN6+3KAD5uoohrVvGIwf
PMGFXdRdt2UHFe312/5grTkR4uaol3cwriz70YP5caR13sDxfG8kU/xldc+M1iGx
AlXdgt9dvdMgJaEvpMbynSytRfHG8yBOa991VqJa5MbwYanK/0JiDxUiHj/cggKn
taqxDW/YiJ45z6pk+KZGFmd6ol14+GkfQ1V+1P4oSYkJzxw4z/5Oobi4B1xrgLG0
mZ0t+LS6Ao2Xe7Za/eIrZp8+BhQd+kAKKnV9SlBQScJGGXW/4IHXThj3jOhAUDgr
lvG0n3gaj5dBfDeyG8OE9zEe/Ha+R53iv2RELpKTDx7C4svDWL7nUUswVwV5QgM+
hzJSlr37E5LcmPbS5KG4rovzLiqOY5HRoPl09lYUxIn0JmQwsG/FYSa7TKQMxRHE
YLTg0EJ9xok/r6gp5B6KJQJuk3XWb9DsPk34wsVFL8Uo8krDjqP3ghQ8KvvKlb4N
CFkhHMq+XTXic9HIu2zZYoc1j8guvKq/64EsUbXA/Tl04VIPWOA9hGFHS5G19sY5
Qsp7cE2aeN/3cHqo1tK7ZPX8ZyesyHo5UTdPZF+DXuNcd1uraL6NmA7JyXeskVDw
yBkTBTvE/DLvPSDnJ432nqcNM7G8fZpoQn4fWUwGiq8FIqUt5vd8MpF8F+bYCSbx
nNcCn7YJY66TWPhXc9pI6JV0A4dmDF7k47tAs2D7wfAI7rxa9EOJdlfmxfefouBB
fUbt6WXPfBfAda6Sx3iQPtKqeP6OOtKOiH+72lSCmEi6FEoHHh4fdU7I5+XGyjV1
4uIt/ceJ8m8rJv0ZjNqNn4n7XdceOyDG/DGRjQuQfXO1qKmSXOZCF5miS3+gF7ZP
uXiQ97U7vXKGg4WYYCB3uXMbqh4txhnNTRV6EFRqIx2VYsV8N60nifD5OQZJQQ3E
B4hMY51DQbeR9fiO5tb5VU4+BgdNjQuPB+0SOai8itb6ORwB7FkS7iGZ+AWsgRYH
5y2IaU4CUalsUwQ5LpnmU3cENVTCrEpWEWSQx3lInOchmmg35scQ7pr782N3JqFq
dmrmoyG5cgceOUVFnnvN7NbzPQUO/NbDD8idS5+V93pXEsAb7mTPPSG32nLLWzEz
rqh/G6L6GkmzL4A/dpErfdXhSETiJ3SGzyj7tDJjw0QWHNb/67P16vN8SABVj+lp
hr1yM+3Stp6ev4Zqlkx5V6EfetL1ecVE8DDlDAC6TvR+VzK2kk8J1RLUGXLFcmz8
EeXR2jkYcHCqKwb99S2M/dwGAlu16MI4LCJLjCPKk+lot+aHc1yqylDeCX3fdasj
+TUPK/GOd+OReqKZseJKa1ACvCvk0sMEmYraCEyHx3jdjxqFb/OM43XwFFaKvJ1G
us58fTTYG6LouDcPD9kl5yXzGwnWpZog+Lbg+lX5wsUUTgQ31YiyJ0dOOt8y7G4J
ulylwdPfLP+KfHTuSHd8m0y7Ha7HoHTSXovDRMO4xWgv842Xhq3phXhOEnBi0N6X
ZnaIQSVRA6QfvEp9V50csMCk8OJtAwqMw7Skp8HIGxsEVFNJmBE/ys3Y0KTqfLbM
/m+7qIote4id6ifzF99bxS6R5ZUJDEIEE/bGWSbYK7FfwZ3PO/vR7unUBO1SqZuX
yKCqTfPMiaILPTLOPyTJFZ25z84S1ozb+Z3V1MkBdcQoJpTbDicWupeZPOtnTa9U
l/hc74MUyyqNkb75fERZq27hqE+OLWtv/xexE7ENI63nDoHOBY6+4M4gzKMEixah
EKIN76Vzf550yBf2KST7WzAT5WYNNbYLns1UK3EjQxdquXozEjPPKRGqAXf2cl0z
QnA0w5zTqVrvagWBt9k7RJT0LaVCmzu8tdIme0W/x2GbCMDQrUT1vFXrJjZmJN/0
3xJJ0CaXwkaP078/lnkP4Wzq43moI4ty0PoVkkS/thJ2jFXIkVSn+aen6pNlpBiu
oHSvXwg4TYytAv9g4Xo9AqcxmXoD/vsp9/2JP51BW7FrWHxnp6md2OtG2HYYhHqz
CRLN0DQp5E6jm5DuVnm2K4wGEZ51pN/P3DEyegii9/aMuHAhsKUxV7ebQq00J6fU
Kj83Q5jWzTgiPpLuGAQGGRQ71FgJyLT1MDBTmmLj9BhlDCZSpo4HG+ZoGbilURpF
eFsD2V2iLqWTwncmB8gAvlkQwuLjQTauL3oacw1QUG5iy5Iu/JmmngqCc1KYcLoU
m7ISAEaR33bvXRnmC6BdS8qZPK0Ws6bp/o1ttY2bjCDpPgV2rch5bdu8MvjglgJm
FpQ6540W820LHIFtAZuGLh+4gkytalefk5a54YklD/6hRUzyjUx62msYi9FA//29
IPvj/pc4Um4B0A+CtW09BaTd5qi0mY7m5n8okrXXkYX34tUo+xnF4nGJNfHKJzXO
57F73EsFsfb4ToNWiZs3hRqDvP3i+FBOkx6hEjsv+hMkdvZM2BOiFFAwCnvAnb32
nW04SVYm0ojOJVsulNUQGuyAIdx85iMP2n9AyUl87FYccvrsjjTsPtfVA8eDvK1Z
CQ+eQi5aELB/6AcgtqOXER7IGqQIHx6lUlTbtVuJq/P38Or2SC+Vf/FREJ20QZCo
5B/W3u2snMOz1g7fxgpN/M6Iv5CVB81VjAyHYB4cHp1dAedTj1ZQp+lZ4kWczLfR
syRj3pE86/6NEMCSYBoE8Mt90vltMX35E36vmN3o/UD+e2WbXkbzGDvvzXtbh4ts
oYA0dvwTtKj5Mt/YdDYRrGnPGHH1XojEAxgyP2VCJE6s03IhkTc73GMIEWTkXyms
6ME9uUdqKqM4W2XXzStgNBk2pmQi2mGB2LvsLqvDaMwFpkNL7W2YL6itoOyRsYJr
9lh9+VZWNyvb9rjjSk0TDIAyBRUD52nZ8wVl18V3jDDGt/PKeQIQ3IIpJZBZyc3Z
8HpJb7QvTJCCMfPm2A09JZW6ZdRYgWm0D+J/0cNPrA1Y4SJFTqyOBPK1r/AMiaDv
KU6bnr0a/JFIcNl1ML0S1/LWNOydsFTlBRGytWc19WJ+rQqtcgiACaYZ4rqx9gWT
gSXixIQjt6PAXry/xjp/hbfGKDkBbKzW/VlJtO5pOpOMoSnOxZFJkar/7llfagWE
ovZT5JBEC2tmU2CMKANUyemNoBxchfM92W0WfVLfulTxMDENtK0Oy3RvIeXL+MBx
+AM0v4Kf21rbroWKBNb0GGHCTrPFbQ7Hxm9HrvvDhm3e14VYS4PwTDrmlmu91WPW
/YXg+toMU7FXDIrQpmRTlZigSffVAHiJQLwW+5bMxpV5S8GZn7qga4jUQhsxlg68
Q1+Ut0JJnuufY2GP3Z1W8q/8O7LGAFnYH6F+2m9E7v+GbmUpOoOON5BsNI3Wg7kn
2OMYILNMtnHFAEl0ynfwNtzv/nBcmOORIQBzyWJDCSp2uiVLbVYvsdGgLyVo7J4l
DBmHztcEOMtjQaWEphE58OOek1z83LJoGjUI4oAu8rgWO5q6IjrCnEURsTumDKW8
OQ/Op6Q/Q6EnqC03JSvKErX7nX+jkV2HQgAW6wG1UYf7eVl4m8i1HPAcRJvAUinN
COzEIT/947zevpX2JwAQl1oLGDNgZKeW6RSmBLmCBbfmi+JX4JPVfjspNqm9j6My
vRY+9KGaEmiL1HqhjIP9S1I/3k/AlQvRUrSMcp6c6RLW6c6pPL1nU3C8QchlGm6I
SSPDVHr2Z9VfT6MokOcUq2t+AhKNJ9s6WaLBXGeUubuqainCuSxYI0GfMrK1xu+/
qaNo1Th1fonVg+nFAhamGOOsP7USlpL83HSUdOayCBGsvPIVo2ssf6WFqxvCvbts
Xfya+t+BoQxgw/W00YRc7N66QN+XYXwiniZAPgcJxO+0Sn6hhZL1ibJbliVz8Pvv
2XqPZMP7ktibWCjBsBE0b0Nl+GqL5pQKzkaBSwPgv881VHNRMgQFySlumfa+505I
o3OQWmyzbBxqxD3wNF3VKQrV75WHVfNvFwkCZoSUN9AKpBQAPR4eTtwyKpGI7Z1k
IF7FtG9e1ZYU7WQR6DbRss464tVPvj/v2vOmLak+WEDmRtc/dGdPPT0khH8CkidY
dD9gw8izOMStwHM448DK1y6ibX4ETMCtKbytnaWblTW2AHwcpY0Q/g04Jj0nWpSR
aKQz2eLK5bLhMGTI5fBcLrrDcrthkjT0RWYdDj+FL9aHb2I56X3ZlFX+XZBEP+xx
GyC9i1jzc7vTMnFOuTBTPX2E5mKxfJAR7SzySSI7b18wtI6NTso8SrfUQRV3HK9/
RqQFyYgZVgKV+F4s9e7xqPy6r8VFq8Er3b5ueWplRE9Jia054IqLpsvjvNc3rbzK
qYiTTbirKkGm1hVOrsEcMWdNO/dqCpbaJZ8nJfWU8T3t1xKBlILjTy5KC4IMdwAU
/WX+DhfQhNABKq9oPFF3T71pouakYwR6vC0ck8j6WwprBRWxydvTVUuf7PtSvy6D
y3O941ExG3ICKxSqrNWQ0a+Ihn+ykZtJSrCUTywhC2D13w+orCelAMPnNA002A8v
b/aZ5gngbOqIaNqWgIcKJyNuY1NZ6U1jkI0MzHOuHK77JYNGrY4qVG4iTvLaxh7e
NR8K081wZhnXPaosI0AN9i3JS2f7nz51ksbn9O2rPL18Ymx48eXZrciSE4NQWgfn
ETy9k09eYTKTPNzEjvg+DmAc0scPhzQIX4T9FwjU8VrGolMcd+1z3vo4cZFL8FJ5
k+/u/5+6EsgeTKtyxuE0qtewFNXVen8QrKRCGkmCU6DKvBaT1JDDW5/WgWKi7P9D
P/t5vgYOT1zW65Oup+ZD1bShbZyoFb1ff7Vj92BweF31eIDGEJkLZYflIeycinWF
2roPzsJDDNZNeGLuKanQWwfL4bQSDTDEaswYO+JvI7K7UcoUsVL5wuUeT+gerH6i
s8WT4K9wUBmQXzXUUmIs0ZS08AFPOyWIJ3duyboddstGTHnkuYkvmoaVcHIytb1C
lBPSOK9RvegOEcFsxRQNRe3cmBD6c1MCf7tZFxueXnoqjF9lLzTaiLP2DHWpyXn1
5jXRAn4b15FsUxz/sR0QlaGJ3FEWFEyg97+twafeUapfjkAjjPAVyfYzeSo8LoEC
HlerDsISPQ6vVAxKLDzpekNL0i74Xl0XsHQcIbg9xu8XFecQU66SlGtzrQpb9hvK
uTOIAKSFd9CkxNJSmGRUQNEl5aL1Z0rm4dRJ9qkxE1sqJ/DOd8Fh7Eifo1TjlmS/
ZGFfhgqBNGc4HtsBJyMPvdE2BI89jQ9vZaQH6sDxjGAoIIUwfTmEdpjEXZl1pm6s
1hFyYTwCddmmOFzXDfhaPIEmOnaCk5eBMyH1quqAsdEERurNdAHSlMirOF4keo9l
kUtipeVchURFWfruv7YcdBNhDcbVymC15GObDi/3nOmjtLNT+N8OATdEciSXZdGH
mpE9lBtaVHkD/euV/Do9+A1nhxyl/kqgP0sQCS3gZHm3WKZJ06rXqDq+7xwYcgPd
VZa5rYGfo58EtCamViqabh6fDoQqDFzGlokGUKSzWLmp78XImZMQwIOA98MR5FGJ
7GvVkE1ARE0Nx2ObE4R0zYeDLDag06++jS9NjHRxCaeltrwZxCHTqpIhy8BHL2CR
9SLbj0PtQcm83dJvoZFrdUeZonlTDAtezf5ojGOrx8Sk9XHpQDVNTQ9fpBEtwqBu
pJo9HFFlweqRfEoFmQHLpg9t27KV3X91BKDGWnuDkZ5YU/f6x3QqECDOpG3ZD3sp
sxjg8/PtJbjkgtDDzghnoYBZm7nSkfVSCyAOn94CkrUlefMy43Z7JCjyjr6py6Vc
3gktqs3H8dWZTWi7dojUXcmFq6ieKuz8N5ExRay24y4tjhlIR5KH3QtP0uHa9ngg
iHZ3xTIDvJBIDQhzLYrDIBfsyzdlS6MRe1xs+t0Xho29PPnkACqm9bnZI15zRBVq
1rXxaKjPsc4JMBmrRLOeQlIqel1RFSgzAFlo+dvXMiZVF2zI/7aDmW8sNQlKjwAx
EDyxGazrq5847z+4g5nJ+Py4XJpcBo7fVFS+udQoxqECzjpJCGi7lc2hZAEtCm1p
LfyuQr/hFYn+XH491qnvIVK0Oj6hmzpBTjla3m0WNqEromdGij7UiHcHxF2tYoQy
kGR+aN01qN6BsHgf9teo1euEvVFja7KddGGWd5VQ5TUWxFae1yVJVTOIeSDCoxdI
F7ApWcq8DyBdcpvIEJcmJXAxDC5rUSIEd6/cF1A3oEfxrteMYm6gimhgGWS9nW7U
3rrXgp1HHR0TuS1Emu2CktXJSvlHd0XA7iXRipLr23R9GgHM6+az7sfa48ZMZw19
I3iipotldKZy466apMPJo1d7/rgQVweclwT6i1lWUihHFlJHXmiFgK71mhs5ETZ3
qLMdZ5f8k5SoYzDdWD6OyTLKMVVRPD1Mc+FBt+L2v9RKToYLNAPVscA8JR88T1wb
DwQjSaJ93JhWO9EgkXOKth4kZG2Hyxgtnk4FM0JS+umzfcZn+5ugjPTxB48PdTPs
DX4K3tOnkKw4LbGNT6Zc9t+HSlbCdq/yGEJgJExYciZhvCQZxuCyEupB/ECkJZ90
QoEuPmCB/Uf/T91KyI9c0Y4HEk6FW29Sx9KPT+SMzRYZgV25rBN0SPaxu3nWu8G5
eluqs1P8IEOdCcaUZ09ziOuvz9uihxhmEgDFIyZbuUqYhAPhduCN421+iOsm7Esq
4CAZSBMa0ktU3+lMUv9iCRUHnJrd1HRJ0gvpe0n/MCvLUWIi8tCN77dnUVKyHbD5
npGB23gSKgFbOslYcy2e4ACXTIIyz0IQ4q0Qj43fxH5ztIxmORHfaElr91AU/Gl/
7ycMzHVm+vF6cBEG73W05MBVHxu8lFmXliUnr1/R/kGpO9U2rES3WyphtDRgP9ub
lenH+chKBVwiZggaqLyrbzL1oPbKyrpKSzpLZkC5RNPdTbMnJfEeJtVJrPBK6KvN
Ece19NuGoSI1JJbzi978IIK22s/X3OMprSR5OkJyxlrK6vjm6ViX2dmG0bbTULDW
g5C39A8ZBnuIAZUnNKGGPjtDBdlcrDkNtlGno2XQ47bDrqQcrBbwOPhbc2JK7wpY
X6WbFNKAsK87LbIaIEeUETFVzQc6Oa5K02IHBcMRsXSk18jgn/MRCD0WTBgdfx7e
qKlHcYcUixHQu+rABmqj673xBqCAkYL4suYQNiu9szcOiSdx/xvRAS4NRpHJYTI0
9d4GgAi/UrOIqIffxT033NN9opXJBINJT/ywZ/0gK2Rv3lRwucHEo7SNWd6Ge50U
ygdqNNTXNbcemTzAV8qRaXxySJrMZTNF9UE9jHa/Ehez0AvVJBqscqx0dJxNdXdn
0rXCbxt4FgCKklXUQtIGKZ3WWubhdnDTafUnZrL0OYSR32qtdylnMljOqzrYeK6d
jBbeRyNFy/OfPqKcnXYZ/QKw2iFMmIOlqy5smnEXEjr28zylYzGAeMPcxdKYTVdB
J8To+g9rVH/54+DnWfzrjVN3LQbIrjtCdxkRelLZQRz/ajw1kr1FCardWhYgaYQS
zAYuBTSZbzk3oFeSqCNhqnugPiPEzciMJ1iR45GnBpMHArTG8xfEkw5SJ1csEj3Z
4znFFM3uutpgU8XdY87zn9DI973ykjEnRpfKfeOaxvdb6pS1E3NQt6X13vUj2Pvz
VAOeIN+qRk/DN8dU/2+AW89wYhWCCmmDXiMJ3o82uz+3JStFjgNLcX0wf/poRFPT
QjVNZUD4vE8c8tIzqiD5L3MBczDeCuSNntDXPGP3q7a/vdBYzB5Ym34MLJehK6xW
SNHdLKdCiEG2HxxeEOIhYweUVSOn0fiG9bcXcx2eNSfixcyRCAoNqyzfnF6ypWxk
6LUlf4pzdxCiLl4abVV0tIw+2QA22LhMwvT6arHeES/+JBq705E8TihqpslzNZic
Or4v9tQhs55G7R2IvfMg1zqDG/AwVQUE7Ca3dDLimUGi37iRpuS9/gavFDq82qPq
qWLL7BANjx4tHAr0nKqDPRpX4CCg9yATnlvSyrKDe2YbDPR6x/xrRpWZrHz+bnbv
HUnNQO/PF9MqkGZNiNQwHbQ/IWg4df5dPZudflq7vfoSJFqK4qRkkAyvHk+jze+L
TBCGDTaxgWKqOxdPIojYcZymYQ8yTBVWWJYnpYmco4zI2qxSUqZP1fNrkvTOv71Y
BIW5eX5zd2iAjiKforxwOOjdYGGYDdw3Dbk7rAxtSiDjnt4uNjjBa7BBD1SLXaRU
Lg8/sY8AhtbW7/ocf0ikTc8ZSkKDMCjr7sQqEaCE7MXWUKvkAcyxneoDyxyproD3
G8HoRuAUKsAB4WcjI5n/UoWXsWsOlGhfrp0KZeWenSFKpyP8sKPXVz3zgsJpYwy2
HpFqTB1+iAm0dYoZal/yXoX3wZxIiznsJzyVyC3XkYOf8T7IkJJsk1u3+zqvq2Aj
Cudw3t/oyxofSXB0DrGpl49nl9r/Qe4Wr/7EjZQnJsugKwzZQ2kWcgcfoWDoTdua
v4j1/usQ+gF5cRruM/7QXU0SHq04Zlco+QDDUQCD4KQgZUr/PO9B/4SfBagXt/yt
vIr6lLvTQNUTDfelylucx87a9VpxwBA3gKokUxfhe464CwPqfB52uF35g4yNnu+m
Js3kX2fxANjoFKyq2B8JSFOQZc2lU4JA41qAk5EIrF50uT8wWNZrHxsJ98B4rmYu
S7CTA678ws5BH6o/7i26fnuGn7qfk2doswaqgmXLnis6QnIYZ1ZVCPHjp+nZLleS
hga2iNTwEuPuZl3SNQFddU8ukZLd8fOZBT32Y8mAOkCw2kMeSBORUgZzoymQw+sT
i71mcBlFelRmLyjErrdWbiJp067f6VA08EBhRbqD3Cd343XRnDMghhoG+BjDnQ+G
+L5b9+vmmbX6+Wut2X2nsPFF+/a71BluGXmT/GLw5zxBz0Jm7QGwLj9gNjkC2wJM
Fo3scZqg3VPB2QMfcsGXHGJjt/UHLw+YG7nJQQInNqDER4YSG14XOnzhmzc4NOLB
Mm7fyYYaa/1hcMb9uqn/9fy7AnsNp4WqkRINxPwvjOvXBOkghcdLG097d9PRef2B
uUY2NKdX135RJoCUHNJfgHIrAVCdjwSiU8rmLqsGhpXKqrfqwtZf3c0no9+Gd7WI
rrMYS+qc4BZRxDDnx7+7a9r/fs29hFG95n7IDOeUl0H+YsKq6QaREiKTOs16a8fL
70S/4zEDB1aiApLmwH8aozKbsBoKexrGNxgYnm9esL0ixKhIomCE++wJuNMwX1Gr
45CBk2cmqhecwKn5Qk4TEm9to9Js0rBn81M0oVDYbmBvt8yOrIOZKfpjAtAHsbtG
iwvSP8L+NuPLVbH9VMFQeOWFL+g4JWc5xlOnuzzOGOfglIA/B3LMFqUhEyVAFf6I
oe9FHZ8RLU2b5My0C1KAZ5z1Xk1t32FTwUwi+xWJ9aS2JAvHG/1dn/nLFvLvrw4A
CPqOhLHBGkICjK1joTfXPxr0RtKzbzN3cRxoOhfB9y3VmlQjprOpVU07L6a4/HPm
XqwTcdN1O88WPzZ8RmyZ3eMnno5Q9kN2Pc4atYtdg+6Sj5D36B29SYCAXNo/TL4a
2YmPzCU1dLs9Gcm1FAkWajhsf2YAsL3AoxXdwfYhHC61jNke8asKYr0APQKIu7vY
pQ50LcenVe47pBdD8UfR1Ip3AYVkyCFnyk/ViNbBI6tDGSg1JnsQivHt2kSXcNrY
Sfy42n7nESyjBZOdModlbxq+RGqKsHl4sEeOW0tKTSnlQbKbJs7Zla+Bea1g4aZB
uijwgse9EetU1a2cLolwUm7oUQrJQq4Bq8Wbo4qRI7DJp2Ye8RRpMY3Xr/POJJn+
nwQCLoEyqIaiqMlF05xJl7txXemwEjSxcW1kl4ia0rp9Wzxo3uoeqhkt2A4JOiXQ
3hYh2TxflPdbVcB47KC3AF1gAFg/jSsriz7P6/0xNIQp56cTbCKbIdP4RgDzu8Ng
0jjmI94dlkU5thh1hnigsbOXqCeWIa/GpDr/X2/KLIoPSP4tNoZHVRP8yvoldg4Y
Ul/VarGeF1vOATiAtqB9pAkmr8HwRRnV2W8sFr6r6i7gKv8SAgRbxThc3q7he/Xs
WusQWHBDGZ103WDqOBlSm2BtwyyVo3P4sTs/95nTKPyZW2x4E3YqCWQjyDxZov5U
2ynR8y0LWEXAwhs8JhnyZh6ehy4rRP6gpaRIz7itax0OEvuw17HdheYA+vGuJ2s+
gyD4SOTeE9EgGgIC3uz9i9kGgwsHgJ74JQho8Hzfspr0rjbzjzcgpua6UR0cJfba
VTqbipFa5xwEEXKu1JE0PaIbSL5nLGJLMM1Yp4mcukqw+ThYzQmAsHs4iT7cDhid
df3NmFXcL1Te+Sf9y/YvLWkbJmyqBnQJHqoggn7hBdl77XJ07YIxa/8/BVjryq9k
WNoLwkXGtj6zAS+89tNyi8EF+u1TAFI0zXLqFM0Ls4RXIWOwPkR7pGcW0g08AklH
aFsMy387M/VeZAKYEaL4MNJ0eDo+jRd6pqTRh3d/n82FhdVuore7OZf4dMC/H/YA
7aqd9dFGzUm89qOi2ik7SRCA7QqAVSuTNHuEHrvbMIZMj1wLGy5gn3J38B+sllFl
eDpSqG2ZIBI4MQL2eTB1qWu+DMsPF4sXaJpZ1JWIk2ZNtmDOsBXa+HCJTc80AqTl
kXXffUoYalSqr2Uu9rN3legsI4G2jq8Q8JZQeXbk7Xk3XkCXjBjvi5ieQWxYZUW4
ifCY8j7PHdwLhSar/bNGlN4Z22MjJhilfbSioSK6y0R9190ZSm6dfe7tlB7MlbUt
acspbLDdcSlQ9tLOmAVYipdwQ3FhI5cxcEwD9JuDqvI9K+IOzxJ3hlqCZCl7tVVf
9X7s/ZjtYB+m20B3jK1h+vfHd76fmDnam27B6BAL+Uoh1RGDud5dFNbzHv+IU3xL
dFjxANQTkE4g1MtVSxvGZlB4UWLb7Hbbs7pxXdqnKHN8nqyF76x0d8YeLhEly+fJ
Tzr27QLiE+8wBzgta08rsZIeC7FYKqhZUSN5Gh2N4Y4vxxKAHmVh8xjQGknwmV8g
QELqy90u3D0c39xGzrI0ICW5KoUMtWHjoaGcK/x1jn0ksdp7NzyNoNvWiLwhS2Vg
zQ2w1XGap+C2GtD/0F/b0dSE3wEsUJALzE1B+5BlFEQ7TJvILXGbzIFFYmvnEA1k
U9Si5BDxm9TasOdmzR6J+sYIzFuZs9ng/zuFimbQLgoerew0OVVBWa9l11n38vjY
FD1hAVklH8/t9nlyQb+sjQAjU1cSHuX1W0IJ0BRq5QOupV5NPtJHYKfa8j9R9cWF
z20cXQMCOtCvuSUBdScBUZTn2ABCqCUvOhvOwdQMIOrUppJwPqruqNgiGLYTeScE
ghj9ADMQ2RSjT4pG41tBvrMcFlge1Ot4RrDLnE1WMEezJXsqzqyG2bgJbxsp9VpU
DRCq1cn4pMxmQaWraZ3Gq3HPr2WQqhUu7ODyW1mpCY/uRkCRaF+zfcbpcKcwCsMq
IDyFkP5JGHuRC24F77JqOEL8/4WJpJZn5Lo9rhY8PMUmp3aOTk0+70p08JxkwCKx
Z0FVkwU7sHEDOh9yvduCLqaEr0wBUXL+kq3FJAQfGrjlt1l7oZaXGnGVU13+y15a
VaM5HhkWYPyliM1KG4dfjwYoRIM2Lo0w/BEwbptiD06tLH5JRnBAY/gNKMqlHd+0
AmH/oMW0CQi+FjwBfcGaCSt/jWM1YoV0VfNleKN8SsOYpxBRY6cutVxX/s6lH9oD
KyQ2NUqD2CwlbRcpoDODDQDK9nSE1lsx15rGB10zAZ9PBNUL4Gn2EiqEytspEpmx
fYEcpkzvclm2pAkyUEtC9ApXFnDifHczjxMORYDzY7SGi3whMcTjdMN63NLQoOgu
ILvqsUvSKbrY7L03cTky6WsBnjus04uFtBt10T2ng5fTq250J8KRsDvVHLsiPNMl
fDCLXjk2buK49jxwSStD58UIq0j0ButqINc5gXw7XE3q0aLDa7K04qmCwZNDBiVo
06Q2Wslr5Dpsm/NHvk6RkN3l9JuQBBgF6JZnySxSjYUgQF6x/6KAJiDqlsQoGmsI
JgQXLhOMbdD7rI9piuOkSiq5xP9mRo5/GW7GSoC0Dur8hN9vSK/6+ynrUjW0ZaM8
IwZn9t31QJXm2jsGelxpgdOQZ8/9W7eHrUUkUBCEPFVS/v8KylSlF05uOgsEaa0C
DyF7UMX/BsUFphxEZGTfmjwHDR60xxxC9yw8MuHIB2/cx5aalLWALzH+5hDhzKAI
r/QHpIDEL/hHFJQPPjX2SVODUt53H+1zVjuByaXBhlxFoCfrH1yMZFkYieNMZoYr
syvfDjdj0PJ71Z2aETi0nPZ4yH2/yCxOgRjXFMKmdx4Ff0FNTd4Go0LHe0p6C4QG
I25cT2sEORx9HnOvYYS8+kCPk5Kxy6RIHh683ecykV+VO7k+ga1fGhOa0uQNo/F0
DCgO+lE2hWzxywTXMhiU6AGtv5C7BFYKs+UmQ34H++7qRHLFdv1KlgMEmmUD0rt/
fag6k6sgSu9jPcIgWWf98XjO/eIEEDuVmjy+fGbcUQUsXXyv6zKzOCc6te4mPU8R
sSyhEXTzT4D3FcjyLreTSQSQfgwNQrv16tLMR/wMeP38GfE8l9KhG/oM+62pzR+h
t+pyzSh6807uId/7VdqqSa4WJFYnibyMypb34bNi7hJrwRjeeobdtazKpbCuQ2jC
gOfVQdEuA1YiPe5P+ybg89MbH7OLkH+br5NRi+RbCWZWgFA6w7JWBvpmaAChCF7+
/Jxy6TyS1n+v+JthbYNO4KpXLXgrUiUROHcsID2szNxaZbjEUT5dnJuHm30ZKcpg
KM8QF4/9Jj5dvAeKxJ4MOFoT1xO0sj0sRMaFB7BGZ/GE7TwLxTG7F7efuG/KzNWf
diFc9Mbxi26Ay+XyY+M6vZKgr2ILSe6rZXlTDcLeZRQwhm+1mvwnhijtKnHemx+V
Q+K6ojtfFHAS2G8FqNfrQNQetTgbppH+2rpshWy9gBhOpE28q95NADJVGI/Cgg9D
E30gNL49nCpe3v5b3643hyGkT5KWLZmYrU3SZ9Vgow2v0ap2OJrhT/C6xAlRI2kL
voWaac9cbcaTFdjOuCAhk/T6wVjKHoa60GKrTx9XJqj1uqU0Wn6y8x6MnokvlE4p
v0f0MhBq6vOi9Ui1dFgj1b0Vne2OwxllO0oZLxKTZVQTgAKbFSxMcUdHkuhiYnYf
auzjlMHY3EmkWD6sIx4AjQh08mJVOcdiL24Do0LXjYoAE9I91Fe8K6UpSLRwcYrw
eSOyjlpQnFFpB8qRf6bO7PCGt8jDveY7bqd62gUXImQfxy67iI9Kdhmfwxw0fqsX
6D44zqFT0cPChOjX8nhcmXeds7DHI2xdFM1azAE/VA8d5JITfmuBf4Yb0N73pJeV
LIGiWl/JhmVvRJVkoWIxHML8IVg4WJS8Y8RIQbKjE1V9WrR+hr//3yrp8/WLXshT
FFrwQuUmHaHoDMiT8ehd/GRtRjBmY7rHsRDqFUqM2cS89azkQmhJxtHPaS9QBNiP
/Xtvtz8kN2wvzLPWB++oIQ0BG1G2y+UAflupGyJiSiaAWWtbaBcq6Xrfcaxlh2w4
EsIB3v6bvmRiPLOeA8SElKkqZY9ZVoVJ3O5SA7mL/IYhXUuYpbfsVxyksypbcY8V
GEuX8N69D93s+J2Tq9qGnRWrVCp+3D9zf4V/56MKOn4k/2Xz6M8ySJeK4ZsnUIa6
yYjTvcpdMC02M4ea5FIMPozKOpSSUMD/DnNIirQTS9QPLiUvn0M3fQYIlC7LvILs
08QNCzL4kvxYQpzDopQmsDjGtpuGeecmU5ojfrRQKSo0ikx+QuFMIbWPAXrlPLHZ
Z7LJstXJd7YmPZuJg+y/NFAER3hKR38qN30Pp0C4uHvm0y2Mu8qBxteM+dzXxAuU
zy4VZR6P368aOpG/4h5R9swgMDQi4OIjqUQJK0RVDcTia3Ra1lDsDDXhl7y/04Dn
CtTH90Uvs2WdsGZSeBMigTkvz89fpp52PwSo0T59kWW/X1x9Jpw6zfAeLdWPE6uV
lfIVizIIpCs5FojWRMqYvVkc7egeY7dL9jtWTd7nxMlhdvvnkmnjRkf1ZP16saxI
Wvt2cmrMH3IjegfDYEwemkrJkcK+jMvJjQcORrlHmrDjgyGfndCI2eYEQEl+13mv
Q87wEojAYP8Z73DhLXYNBuln6XUE6q5OF5o7pI9yJF+KdGsDIJKa06RffKTPLhV+
+wb2zY1XGiubbAHmGoxIWY1CU8SQPARGVWFrthWqcubUEPvIfwfprAwcNs+1PPf9
4UFbIL2EKntXbqEqo6AmfPAbZn24K7d9oTdocAOwirCvjaLEKEWkzoFZPhEyn4EJ
cKN43gENy1zsvVM7jLZjmNtmXFXBOhXuvx5Mcr3sde2S8ESg+l5fAZBmIOiBtFEX
4S1z/3CEmHMkCoy22p62xGEu1PPjEL9HVTNZEHxt0D1WJLNTVIBglCs4xTL2u5+Q
SgcTcuw4zmF7VTOGtO3zuOjJWftvyWmVTsNl45vj6Lm4uS/Po/UjZJ0f06SjuwC7
G4jVYWsqzisisU5437BZdsPPPNKwDRcgyYyWajvCxzAQtt1uvEuchcUajC+Xl/SJ
oxeDSQTqjsjKoQZpV9DpudVx/e4QRAMHHSNgelzsjkyGwvymNfuD3otvu56Fg7b2
NDbGRfE42nVRl/1vn1/AURT6+ANWThB4FOhLz40xdE6MONEKOjTn2vwZxtCNerF7
wMqxNBOMhA/MpQkIOGXPJ7QjWz9l1YvAgWYOfO9Mmt5meTIgFbz2Ue2kHSd0nQfC
xy13mw5iOQHsZpnRVIrw1ilYg+8cmqbW0p0/nagrwHIazV7/f7INwiso7ayJN8pT
7C4nMyTRO79AvdXowwQmB0LOcoc52v4jVRsN7uwm2Yuvs+UsGhkfbQ26Z1axgZUC
cIAQT/ghU1SdGBBospOz1+QAR5x2kNu9E5fVgvM/btkOzQcbEhXEyupjUAOxYcDJ
XWhSLWMdBcVTNA2zCslIkFzmCXyhn/Oz7dcaxvBFuNWjvvYJ1b4oMLhsX3HaS+TT
1XvL0uFJf+XNRJnXfK3432AUc9uSZTPYvmPbd3wj5ptyQHbr64rHETgtVkSrrTq8
tQ6cdrtL6Sjw7WOqL5tvoKJRL1/v8b2/QdnA6FoAAW2luHm4QmzqZAfZkvK3nhQ/
uYN8nHAvdKOx2zrIVbMY9kgIPIHV3WzkTa9vSeS9JIXJnau7riHoVYwv/emfA0Jl
DLlSCNoEuKBgOt+QdgAoSOxL6G8InGniGDTWcSjQy5cnNHSqWwFHOa85ONlqoO/H
KLWIXt8seAEXny8rDCNag+A4Ly2mUfckB3lEWSm6LVQyS/d5NHQFbN6tMh4BJgcI
odScAEzrkDryuYUSb9ZgIlbhPxjaSWrV2UxHnAwdLNe6m5ql7gPkCVQymUNpOdbJ
ouG2hDfxeZsP1BeQx73OqfhrMy84gtggRYo5ARSr6r5A8DaTQf2QF7B8tdx4RbTj
U2RWCXwD4Hcrg+zT0evhYuPXe+iIWJZZtwzMoGtegN4n9XEKwBki3BDIciyXdrZP
jP0lRrUnQY8KTFAax8Y8/n5FvN3uWeB3f8F5r1H+BZHEEe63gVqNVi1OLGKDHgBX
jHw2+nozxUzf8j/x50yU/elcV9UqEHRrKZEn82LXdmvHxWB6PqWNucjUMXCNTMDs
ZckcGy76LN77enZ7KaSwyt1b6ORNHiqQv+K2JjJZrPuFjtMCB4uuAKebMYRPI4GA
pufPXwB7jgKnG+Tbs5kjNE2+hrQqcSni8GBjJZetmj1VzWY9YbI61j1tZq2OBIx+
pB7P+sO1tLrxSSkV4PxK6U/jYSJciiYSQlyUw15YP5NBKD7JJwi/FO6+tUMzMHWL
hEPcITIPfoMlkH7WFkFV9F2Bi3eC/SMLFNsfQYiS4qCnxhsG+X7HxbzONK1oQtWJ
oRj3uBD09tYWfxUMyzFF8rU7oKlsLQJkR71MxXh4IXJPMWQTINzVAmSrXd26TwfG
zGbf+xgbggi6LMnrvN8QPL0Hix3IHhsKPKM3h5Qe+eacoE+qejQpVSwuTYB3kWFK
4F6Pwqg/k1o2dQaelfYU9WT7A4Lefy0Hb+TEHgzteiXLRTQaOPau5Yv1KDYCUciS
VtkfR4f2TYNTUz4Z0TGa7m2HhEFRTZDjn70uORte57s88QcsK5oxjzxQwrLXcQou
yJilnzSqM86pb5afbhEHWHlOrAIGxg//MvtMvRu/DV2jJEbmNjTgMJ5hGtNcMQll
efY7TSFLaddl/PTo11+gmpwJaOa4DutAZ9/bOy06AkV3r6O4CcWyIHQn5dqtUsAz
cWtHtae3NaTBiBYb8IBAPRAJMVmy9IUl01unfdNlU/xmrW9p+mt0epP+ZDcVK53+
KTWP3EDXGmhJUOzRqRY1OMCC7RciCqhM5WrwDdRZYZ7qfA3Tyjqk9aJOZVi0xRzu
z6YUd5YMxifxMW4UVKxDPLMXBVtBJyUf3CVxbXVDQIJSUwKkiTS/5awd6tv8ZRy/
0BOrlsRjCqjcymZPNuNt4nauhsmOysCcWnjgm6/FVsIXBuo3/Ke81Vv8+NYQldrd
eclq7whFRLpZ/ZqxvGXvxL4F9mmNlmSzzW6nqr5CXGFAVqW9u8rzpEnDJxIY46AB
NE+lzcOYuRU+WQjCfUByh43l7bdZtLxh4yaLFq7EB8yDWNPNY2AaNZhEwWl5EGXz
eHV+yy3KvP/jXBcIQ/juuObejdhu+tNzZnXAPmLDQQeJ9K4jZv/tEfpJ+Bb2RnPg
KxoWyKw5aYmSCgMW2vhvX1yUv2ipGolEkt00xvKq2NZXRr3PQAolpIUdGvC9Ohfl
grsoygKHPa9gDSwzh5FPx7L2yGP5kHIV+bFI4rSM56/o8h2vzIeyi1RKvY0MY6Sq
O6+WmsZlKC0kFlxotzGTKnDV++ScJu5S8IrR9HtJILvE0aw0GWpGt7lZxX55THoS
OocOcZpg8kxRAMTrK7KpYWFoyFUWA8v2XxFLfCnWgCxqlqSbvoNa9UCgV+7vSJ+0
Cp4tVVTpzPOjtc4oajl1IzhVSzV27LPHPWXSmvduZBWi+uKloTRzlmIVumQzX9xP
NEFNPujeP6+peIy/c5YBMGORstubl0crb8yqi1KibyHxgBmitfW4MFPA7MK4SuTV
26PzIGEHOnHl5JVffsMlyFtkNU6hAuW7p5O4op3S5QEcjOZuVdsjKJoiJoPkBOQJ
1ONr8tHxffU5Np6KIIN8DCPTYuStG6UmvIpzifmuNcd1+0ORW7FGNXSgJpfEaAr8
m6/6n+PbQS4CJzSavFwu88sElErDiOny9C+lEigQ+/0cMbPmDJ1Bji/hk9mU03PH
auM6NLDaguCLc3xApOlU/3jQPALe7WsHHQ363R/ynAfm6JY6VCfYFIAK3DSc1AOJ
00xNTdWvsftDM7NpTMDiN33NOV6IAPwZcz7NyFpbh+rWe5SoDd67biVE+KNI9lVp
U4/++uM7yZGGiof6rC3Xa3rOkyLHtBdWo/vW71LQqEyrXyNyS8fVVa1fdhqZ4h3T
EGhnzFPIsGPDeQizS7OlZCqZDk+fWdctUJ8G/zMjIUURhMp/qtc0j7Jsxj7Uw38p
suMnK14srAdkx5wEOT0Miu93gIAzUed0sxU/YzpFG29IjONScew2B2YrV2p7kkNz
ncIzMsHIXdOHQ96iAPiQbEz1rPObfLPCp3vA7sNXZNLbTywTU8TSAqbThuE0oGAW
Ukn461BHb/LJ+5ozHEqjMkSk4c1CLG3y1Es5fP+4X6sAm2YU/Syq6g+pSlPd1K4j
u5bhMPOcs08GHjH8XkMkJZTi23e34oHQzHf04nYvhqLrf6rI/XMo3WZa9zrB1xsM
cusj4JGvILZpjGulam83diGHWxquR1A11kS2CGHE0lpAwPbHrgrmMKR6L9t0rI5w
2Nw3VMD7NdpkhljK2/EKwQejVnScuWd4a6iK0NFgowqQqk1LISE/jOtIRa+Uiy67
4L8FsUGEuyf/X31JZ8C8Nbrs1pgDA3wk9whU/+EWgDBlT6Uk5LrllgjD50p+p+8u
mJGBRTIB/aVHgsdDLzLLxBwexvhwGOaENZ9OhJ1CSYZ2ibQsMcDROaNOZELSc6KQ
zcgE7CUhrOIr1vVNGHqgaa5yFVElyOwI3IzseZ5/T+AxQ17n+U7gNd30PRl30iBz
oV0nSaiP4xTMgnjw0x3uWT+aXlCEPyfBCR2SiMgRkQr5Nu/XlA9UC43h2nZq8aMc
CNX9xcfjx88X6WzT56P/wGuHsvmmajPsAmOhvBhgF4vBSlXphf6g4vcBfuKisI7r
Md5uHvgrYEoZwiM6OMQP5gkoSfqyudMh36WhC0Gp3qYcPtcGary/y5DRNEKm+VIQ
xRfncO0oPd5Pnz/2NespoSy6CVU+8xv39WiVqNmkafv+N1NR/l0r/omLuEy91gso
c+WQ+n6wnW/qUrrXXPpqpw+XZbNQdPkbQBreTI+YRpJtCxgCGCjQgWHPoUNCp0oo
or5qMNn76N//unsYKAzpkv2d5QnWyES8q20AmcowHRofOaPt8xF+1BHgIKhvjCZQ
HN5NwMv5t/TkKxjxpjhGiJuazABj+zvojnA7cvkFe2rWGH2nq5+YdTDhevlGfBgY
+QekCdTB5gUzTc5W4EN/DSjsJav5HRRjK2sCj6VVn6iQ5iARr9VhoZpkXcKEgTas
pPpZ0rd6ZiGrgldSeHboTi5IqfMv1mI7ddmTY4yZ2YenH2GtjnPtIC1s/U6QtKkq
ZG+g1ncg73tdjyofa4bUBmyAw0w0ZOHjAv4PqhsFR3BWh9dzkR2X/+j3g4+pAHCj
FKiBwpmGVuM+xYU8WepxnMCk9E1t8bZ3J6aDwjUwDcudf7ISuj/dD2KYie2S0TWT
2LeUuZbrCYVxfX2psnjhgZKrMpQVwTECl/jsv0I14vM0zd33DJqLpyRPoNZAgHIy
iZTkaL3+wOlcNyb3OwN8oLBg6GP36CSqepq7AkH0FKJOUJyeH7kOnoz/L3Viydvp
ZSyh72fdpe6oFEzSDeMQruolYaL435uTca+nUUR8M0pk/YCjmJoMzXvlHjL9puzZ
4AIu+EjT7MeT3+P03J+lf4AYg3Y8GLo3VjR9uc3nnFzs7qXA2uxm7PerocaUGA9k
h/z5LzTwcF7o9/d1PI3T2oxzsPgBPEJoeFS8We07lExVXfYAkfGsH5veqMROldt7
MR+NDGq1k/swr30fNK7zh6+N6jwKYfb5xvzhaTG1P2ZrqxyowBP+ZWtpcebv7TU+
DX55EiC2YLgKwrYn2FCKmmdXg+9AxoPNV9PCoZz8JcHQEkfK81qCZ0L3UrKurGoG
Ho4Bkbwygw3+EucnR5Jt3InUG9+MfcWBIXcnYIlHcMhLQeZcoBWs3eJO+aAO3UeO
OJ+f3luezoWAtJo4LCR69GeJlb0CfjVgmYNdpwpJKMEfFOPsduq1Avf1G7QdjOma
Yiq06l76R7ApgtMomYkoc62PrrKb0UnNtIYutHSKCoYDKMYMIccZnXpw3DkdeJ1f
Cg/LbkpF/shn43VQnBtHMoBzAKkXFHjw32yIhXjFphcdG7UPxAYb4Wo1b7AXxszs
QW0AUwjn1Wu+vow8awmaOwIDQowJfRSSArOAg9ebvmuJHUWsDsziAga+JDmRwLYH
fu/KaqUqoK6+oojsd4kStgIzMlK62Uk6BxsOekdapmdRHMnzqgf6ZUJyz+1+J49f
CfNQqyP8YM1cKTwRNB8iBHYq/7MKxGoqJ7+Yryq5bfjij2tLLuGy3FtCnaTMYIZ4
/dBWUYtkMzmHKz7CvrPjI0VaM3eIudK67UOXNcg+1tUro8siWdGrtSk5JLsUOK4g
2tgfu8WNw9uX2mDIDsAc4I8mIR1J78Irn4KpEBTG2pyeE0ysQgRMujXfn5rkjNba
wvudRJp5BALbFt5MAi3kQyQx4GQxVNT5gZ2cG7FzD7a5hL3042QZ1+pNLXhhqkPt
BAxgM8Wf3OBqg2Fo31HPNVI8T3QXsa2JznhvJOmJdY8AvObgEYPG6YIMd/wnl9xr
eSwRk8GF+Ec+q9KSGDr5KG8CU57Ko+jdWT4/5ObsXzD9EjdglL3qF7lneG4wj6vn
27pyggziWnHtBSaEgwxeU2fXtlBtAqTrFD9dl0McJBIis3YFGNb5RPV/6lg3DEQX
a9DBAzF9ENouAe+KbHhOGiJZWfpcOpGTGaQZ+x/++sebtumUUb/JK1BGiwFqEx4T
cmSGfBniGU+s45zrlVim9Fcvl2Iv8M216EljcQlLMbV6yxtASCsGMpSAEIyTDKiH
YaiaoC1b2JZY7muBRoFLFv27jynPZW0wRVXXOsI/sztrYDcC5YcmEP4iIP9QdnTx
X1PjmF8MRaBS0NDxQ/K2E1ycMvjX5wAQhlGJtuag9uYSKIIsV/tgx7TTt/TJAb9N
ciIi6IHxxhLHrifN0DInnzlZnbFFk367hXRAWWcwT1nLwXk7oF7tbrfXWa8RlYei
SKP0xjIEpRmylTeYS4YQQN5lfN2AjQpruLEvsWRPf96NqdMCUB7vXVQjan30m4H8
WPJOAlbm3IPPHEPEBO+2goiKjxXvGnUqRn8ca8MyHykr43wgHCA1gbAQyRjz/HbL
NJk0cyKbzrcgUDRm+ybqKmRyo5SPAaspqCtTiuTvO94Vv4oOSK2dfUAFn7bNZdzK
RkD5JRTbRy9f4aoS1CMzj9dtuXW4la7e3FAUGL4zm8VqD4CJG4J4sKmvzM00z7M3
kw16iSR5Hp5JvUQdk1Q2F26Q6oY2ynS2l9kuqdylDjQ+qVKLXBhs3pIfIrj/CHLo
ZOjHZu2DCFg9IG1yx++gX7La/PRKMiGXFVb4tDxVkKq43YBTEBaSWsODeePUN+Xt
ZKPTLBnEN7hsuefyUmYkNzIYjhZrFsszj6xpYJraM86H+106rM5lUPaeNmdJ/WEu
0FxwtdbeINcwvdvc1mHeMgwsu+fD+oZ18YZ1v4GdNuthGdASwU/+4da9ztBEzxUi
NM6jMNoNaa1IwxlkUjcNlmfopNobjOJBxJzjUcqAMlUJ9UstMa877RdJ5FkVuts+
CPQWrJd/A/Jpd41yOvNv2d7/MlvjN0V2+NPcMS9wrWvN6bxOAK+j2SnADPsQelqS
eXiBtv1KC3JA1SBZwkMmgHBUH1ApKS8T9EXRtDkJKLiim//CEO1sNuhLLvgfCkwe
cToo09p2jFvxFKW2UKPPpx0pkvh/RWN9qujvM92piVoiBMVpsU8waYWJ4r3VJaLO
oV5cxH9uPHddUwlXBCzYzsGoK8BSGDZ8FKWXj4BDTOO0tH9EbOo2mqiGZ4vRPqDD
TSpxhbsYTCgs3oGDQZZxwkA90nVAy5Fuqj2gXPnHkx+RHjrHUSYPB6w51ORboskn
bvW3eAN2bWXR9eCK8lxPZeD2RreDVL33Rhwzas9kQ+LUvom/RLMGpMJvH3YHLtLf
sK5/UlVjiMz4EDt1MdFC7rs2wmAyM6xNl9XC3z2Rk7BkhM7NRNjuXvMFfFbluKXu
TUAOimAhkp3gL/JSVjBI8VPYEMIPw2IUz7fbTmuvEi87qPEh8VbMM0tbdWbDKcSH
/gfsuwBg/mIaJDbrAMqwTYR4nxi4y3fVmKGNO9WYcpNrXZAElH3NiDb9kZ6J2nVI
NlXaI/FXFC449wlnSyEM/fRWnUteta4hGelgtJdm6NX4jg1InLCcTBA6uocj5SgW
D8GacKiFYh06y/Vj3BOZM8aBJpLI+GSN2gY7KdNmwZdeHvnrfgEN6/NUgzQXsyqi
j4u1ytcwUUHi2Ozzgzhk/vAhMogsYKdgSnL+R2XRjDPhXN0q9yuo9H4hZLhHLJd7
PLgEu0qpvuqHCXRfPTerPgeP6RGP883MkbyH8M/5r956dGG2U1+7AMXWmmbMzk3h
JPlWB+/vDnx0T6GUKsBM4nlezK7lczo4BwiCl6GalPWuIx7mD9XSA1lsNVwARbjU
qxNMqzBn3x52gUmvDYktZO9y0RejQZGmbHDaZXu9D2sG8z3/Jwnvn7yFEVGGFMuQ
EwHsWld2UhQPUzXLxVtqkZiJXDCOrVo0FbELBPq6G2uIlPvIlPj37ORV9rkB/+Nr
bW5gudgC1I6k5mBeA3lSuRXAOoUYk2ZVTU69xFXBcNABNHqQ0Toxaofl+vJSnSas
ssC2IC8oT6m83191rwguZ1bKRzUwXYBRap8/P1/TlQ/ydyLe2NGQsbt0DV18i++e
S1vt43MQ08vAGJUI8UT2aPNprQz6RIFiPUhxep9vePLrx/3XzJhYLDj7H+kA383s
Blp4A3seFLF1kjmDC8qKmbqWHw3Oh7H52rsRgeHVSAubn6mpqBoq/R97U4FmooAB
bhxzGXgwEGPiaWFo+7AJjsQePz1YaYPkYy7Y2qxGQX8ubTgoBldovZkHJRoEUn2a
URkiDPpzA0R1jLhqxb9isQpbp1AbUGM1X/cTZJbUMgrT0zmYrwvHZp+qbMwiAtzR
yzL4DNDMOws8PfmoHqwnk27TTxV7yfba38PW6EjMSOq+ctUUD55GHtmaO/5edtGS
NytlLHoQ7PVZ7y8hONYqFjWfMXWnk3C3tVb4UcdlhSUDXTTIj2x0xJdK8g40iM6p
55QIuKISZZqZKdWBskWXMycCqOzSaskXuUo5EZCqu+xjd2pctVKWF7fjmOYzW04A
YEakJ7A1+MF4MLXs4I2HMgz4er/rfjlDthFKJE7e2/lMmjhxqEtls6/hlTf7tcKs
1e94rWRcdWfdPeNbucLgLlWPvNT02cqOi9vezoA3zdTvwGGGgdh/FoPtEIC9yoqI
wIUDgQyh4hV7sCPxGhyAGxGIpRTWy4V/DwEnJVHMWwTuaMvBh7aq64aPOSU37pJb
Swxjry5p55IjwjHClraBBl8HgUY2JBZIox4JA7AmaE58ZPgwOejavfMXwWVTbDEn
SGunUJVaWHBj0C7j9NEJVz9xnqqsYl97Of5Z42E6bqUC4YxjvxHaIuRY2+wF9PrW
rVd5QdUwy0DU0TNR/phAr5K2e58DiDhtC8k+YAp1bZhZoPL3q/VstuybtFzFjI+E
RqS1q9st8Mv6L/lEByeLs4Ypj1/qif7fGEgnNeE2aElyvqA82Av+OIvvj8SQczCo
ahn3BNj7IBocrc9/YXXlh3b8wyJ+inIZ0OHPXglAPTJlrt/xDyz5LYZtxVr/QLiv
UhEmAgm4BftofT4pfT/RE5Pa0/CWFoAW258yzxghivnafLwv93OaAmsa/ukWdfgn
7gRu+aq6fuSAe9+YkTMPgah3me+btrhMO+v28aTORc4xDZjBK2eUDamc69Jy3I/J
KuRaCVRE+hdTRUJSQ6RY82japry88nBZrYly9g1STk5tnlNvLfdYWl12L0HA04Qz
6tvVI5hOCxZ4r/XtSAwijSNQppVwauNOQtWuYdNFotRM0U/aJzCz0AEjN+OM1vTY
EqaMxOMlLM2/FXCyGPbU/UfuXNPbL4XD9KjFt7SOr+MwXp06Hix1mh3xWUZv78cf
9E976rPUm5mbTvWYx0D5n7vspUAIuLM6yOQ3W9RWYjFzswrjGdxvHzaghz3GaUMT
uBoW3DnmQK5REg5b8Ffb/O0Xk1ItDUO8acK4qavYzqK06DeBgrS0A88zB+X0uf+j
knh6hkZ8MfeZYmoAieht13Wjej9jl7rXe03ECXzFxSsBzaM5Juxd/D70ROh4VhWG
YPFCB1fIMpXFx/BVIUxkt8pBCQJwm8o2+u8hjTMhb4uvAj+cee2YT4PZVHeDLd8r
NXHEn3HfM6VtBDcfffXc9sc04TXFLsKMQ6kPfuAWmIhBs5SD+5PmM+7L7g+B1o84
bM6KoF1GzVCzv614PewaL4BJtAYN4TRfbZT7Sg/n6ZVeWrzorv4PxdBYo/JMQWg1
mDiqZMzDyAbX7hMOYs3bhkMNhOPibv4KYsK1GLBnq2U0s7+QMQfGKdjQ6OrpPBp+
TGeET/wpNTb4SLBhqSXZCEPNRYLs6ijxWJE5pnp6p0UWTuR3cSFT7lkOxlzRreCL
bMzYi9j0sn6NvqDoG/V9yEQSxetbxoZF6BvxcKs9pXPLDvpwy9qYzcOBUqSkgZ+P
yEKsxKyc0AjIC1TSi6/qhrtiuS7MdWi31etbi6bm0cwhMPygILHzNe86P86GXxyf
n/ggk98J8V5q76d42EKxjK+9ROK++EqrUChqNr9XT2QH7q90f/NDFIgoZwbmw+Bj
oBvs4KP5M132/nr7gt+imjIdWqyf9yABR/3I9duKKtAa0lTkBxyt4FyHLTMSELWR
TkmgxRewMgCJTqdvwJfYS0HG0HMhCYcnml836ZztT33YAKGLtS5T0MQ9yjOF9eJ1
6C/ZbA708RIUMTpJVt2pJn79R15BUOjv4Rddg25icqvXhplATkMyeWGU7D98Ku12
2qijFcj0qGLAsVIENs1xMjGi06sHL+80gnPAVOjSh/UDE2pArOKhB0FcxgoKfNYW
fSUNr4blVbA5BIbFaOsXOC50VKF0oUNiECQURnExpariuZTWn0o7UWGMedN16KUr
24HSt3dAljzhvDpZZrsKtbZ2R6JLApcxvnWNkJ5NPYy8aC0pS7qEEj6HvfKvR4Hu
Ka8Ud//okHC4vO4nt3ZI3qnC2zLQKrv2S3gAG6iLO3b0xstJsZtXj2DmdCrxUzq5
56oYo8rc/fKT2wfWTjZulKIwpsTpJXDq8lpEpmkA6uHsRJ5sAhMDNed+oIxcrbZ3
mboObh5TX6ed1LyEIVnqGIk76gzVJc8Ia2FEnVGGR6qJqvRPg/qj5dUoZAlmZxsA
H7k40an7C8gOCZHf3U/w87tfMPqEwMLzWH19q5ImkaSDA6VHrE+Ma/RaWZvdN1EA
e+YtsOejBVda1zs6QERW03Dd44/8iE+V/ry5kVk33wjjPBxGbczRrwBPG0MjEkGo
h2J6wzItgsor/k9TgNECVpwvyVfc257qXywn1d7X2/2RssdG/lVpCzrDFEXtv9Dk
HshwSKlQOT5roWv4R3DtbgnyR8bdIbbxavPyRcg9o3UDOXnUVHlJTwbfgddBrFZl
yheWszkIBwDb+HR+gm5Qhf9UfgliFArqpMyLwTSPRt/F91a9ATxqrxsMoiAnba/P
CApjwdKejB5NAQFgMXlObNXC46LWvAIvBj9I4Edja0trmBjBMEeu8sUi1UuBDw/W
fVVO77907YRXTWGUihP8GuJyLaAwUbm65QPN8B6AeQ5lqgZUb0HzU4w3e0xIwBV1
4NLY60l0EDgpwEQXOYmJkwn830pWUKBq4WKeyZb4vd/AHMkcmeyT4tbgGahhgLF4
NaiHx0A43988U3Al4iXFaVl4E19bgnzficH+JZ7bDZvc7Ii0lob8VwrFOhJQzU4n
h8rpS63TSA7J7HU9GNfwtOrk6KqGPP+hDo7Pz7RC1N/PxsWXKIIFPGFB3koL2skG
18GTlbE5bSiIcIDRGXLSncPEd1XRMbZx5iPVZyrsoj7WWGdITyacYbkVAWevoiZ4
8aDSrgfE19THuUVHgvfT4ISaFaSj1NpfqcCbM3uQRXBweRI+tu5fgsWmu+vWBpN3
UohD7kkC9osy83OpZWfjlqEtodML1QWI7ZpKZahuznjVD039l9SUywOTEy9i6aE8
G+qp35jFHhtU4VmQicCU9fdKiKvr2WWotlTT/ZG/NTqy80mx8Ymd83zFNl4Md13O
vm6UBx6T5ft2y+z3s+I2ciUNOEIm3lle5ATPJbW9TQG3I4tX8vjIm32cE2yGx5SY
HynsnsVvslBQICRbhYbuYQ5DfJb/d5P1eLQdZsDH0IrQRVIFkPQJ51uvbIOFmvJ4
chOzPNntmt6r4XGN9UVPYWQ2EOEF79y/Lwxav22nCjZXI4hJwSx7bpRq7jescalc
Kwb+leSxNwy9QdaMipT66HjRctc0QjHXgV8mOjWsZbm7+oFhag/sAJ8EGAf7DVNA
lZnPteoMjKld/88vMz1oKKjSbbyglsfqORo41EmrmZFf6TkekxqjvPDyECZ+ocrH
aY7Gi9cOrc8qJCAUrVCMFNyntWpINkulGQx4rrNdh4HOe7U61dD9uxTv/mO2Gveh
hV0FjE+5UxJTcA6tFtUnc5EElEfRBGZC1VCUh4IytZgqUDiBxUJMUP65QL46nRBI
N1/5oHJTDLnLmnpW53HogXlke8X4OsGnQOBdEoHqwLPY/uFimWzHWQe40Xa/Mqd5
afdx/TTSIRGANYtnXoFrPvNxGmP55de7dS5RdpBR5lh3J/2kXYWN8nqxTt53r6cy
NLDGVjuvUXkpb7AprfiILxPPIyke3jtlao0y71S3acqsHAQ4aK+dt+r9s2MlcOBV
67muu99ybYTQdqvs/NrW+4sMHqo3HsdwczB/KpB9H8WkzCnXcc2yJ8o+VwyzkkSy
rDYk6+o3XIM5zjjoEg4dwgCzGmjiWCiaHrN9eco67O3OkA4cFPMufO2eIrMysCp7
F2N/D+VR4F6vR68Nis1B0VlbbHEw0Sl+AmLCAxuVh/Rpyo2ENzQInyfL3cuwomxq
t7ifNARYhqxG3a5eOtNVMxZeimZ4kiF9ByFeldeMfgLVyb4QiLJKDHhGKDv4fAyP
NbF4Kw70cbd640/fDdil58TGjYzRO7MYKburPVG/iA14K36g465LmY0tIj8AlbJn
c8Le0WglUvFHdTVW4dnCL0n/juhAEDF5MvIU0rRkOqn+itPwMF4w+1MK+vHBCimS
BGOrsXCnL1JWpCNz9MxbKRG+gZEOUFbzImEWhofZXJTIXgmvew7TeKoZ9oLmzOaO
UgCaOnWTcPynJRHw1S2EB2Tq6OQzS3yeihKWFV4xwecAo6Qi81ZWLCfwIGmXMnwq
tnqL86ixlGu5U7wZZsVJxHUW0FGiIV5o9ajWk7ttUH1hivnMUzuhV2WeNZbyPuH5
SzZJ1ZVXa+Gg4jJ8btCUrnoM1eZQqZ5K/dp3bIlIGKCIwKmNEXHd7PAE5RnHLCpD
fDn6oJ4JXIYZ1cuw5ehSn0+IM4dXZM91TAmIbxEvVVqr4qZT/ld2UdnOfhnivoNr
538eBwIyMa6Fryca0lmxbThhcifaeyq9rquUprggSEr4Q0gtpihaG54bXJLTGirj
ns0n9501fzLknVG98BrgbTTZKuFjywWHU4YgbOzpgGxpHISycvXhuVCu9t7wwQOr
TaCr+9kSX5trrB6YkJ8JMCDm+nzLL1ghoFubZQevYId//astHctLVRX6ZQuey0gP
TJUhg02oS3o6DXzgR38eOvFHo1n70PBaRPByTggYYhP4X/qdes9z7m8ZcsxZR0MC
IFHkbfmC9gOl9+PX2QxbV6sxdZJdqcMWDIltvhimWnfne24YdyLa7Q8jBKXtFjOu
ruuNUCEXtHShlfltnvO9ibjf5WhfrRMDOUWJIanlu8ZeZt/hFuASS+yT4839+CdM
14cSVIOtiQ2TJuTOB3ELX+DkyxsKUbqZ01b8I5HYZkBoy3AhdDGlJuSmb4s8cb0i
1kg4782QVkDzYAgMZiqSxJgcFRwragplMMvwutme+dT0vLph5Wy8XewBVK3kel0Q
6a+IC+ovK560F6t9B+P7Ci1XuBG9HVj7jmodN31dR04Taa+lJulITIyeqN+VBshm
lv3m1KB6TuMvb7PpNC97owm+S/T0beVkVKmvRHvx9Wim56CYZ34exOPea4tslXjf
Z3y8O4RZM3vjmtUxkooUYjd7ThgFLII1+GDDYcPZcyO6ZZAI8gCLCUFMn8p3o0jX
vxajqIjvlbnQ67s74/Tr5hVJOGZJzxQJG5f5CGGeympEDUcGPKod5PMfHPWWqTDV
ciifSBp6OuKdIH4VvxisS3IOs66WJvB8w9fXulxcDtbxnbDsm5dluImzg9ma2M40
/4ZexBUCpQEo/Jo5adm5NXpLWi71+fLcn3N51SOQa50EQ8Ymr9D5EyrAIZBmQ7w5
GNe0ErUhCzxVC6GhE+/WEcsybuHXExOPODwE20yxCC1YmvvHMFBBKvIwoPo2eMvC
MWWoUsF224zqby531TUKO/Fxyff4RO/9mueb6oWJ4Mkv8asxQRknaFXNeiwousf0
6HbJ1Gr2woStfPL64s4XA717PD27oUFnuUQ4H8dGaE9Nkf3aDkGm9fFTfy9sXQD4
SZwYLDKf9wa1JLSuT7Q/Y4rDIBBR2L0GrDV9kkkcrYyJndDum6esovbRq9cpLwEE
T7c/j4NG1wV1PpINcupS75vi+knlDqH6oJ+QJkrasBcLoigfJkmD+b1pfjir5v1H
NpM8nNzAYYkX/Lj3LCQQKG/6APS5fPI5DOmC67+iDvfWoE+ezZNRw8psVC1uc1VL
/nQcjWnFJ6LmmRpQ3VVHhPeoT0umrZe3lcjpgZL/i1b2h9hOTs0HnqURkNJR+ntD
JhxZkkvr7F/zA7JrLoVb5OgZ4nPZnXU+HE1wfPHpT9eds+ATG6Xi3JPI8ipOdsDt
dEwfpysOcaoukU3injHKGQs/nvp0Wur2mWa6LlfMaMdhjH7YGnvBHK5lS5zmIfQE
qbuIAPdSyX71Iu6IYwTeaJMbbFskAekQThWcuCQBje4J1WgiJ5NIXPXJlRs4Yyc/
RxydpXwRDcu9JNhBJbljOPjwu7YTOVDq7uC9UsXYLjK0ZpmJK56lU0H71AMM0OE2
RxxSS+DCOhL423iB47Ulef6jKQMOrk9hN810TqmhKxt6csDHrxKqD+Hb8pQUzGeY
XRxqP7fIoGGXJW0wHhdwGxlEt0xCgbXcr1MwS1fhT/8gfU1DOl467tI/V7NQ+E6y
Oldd7Cml9qKqrSU7UMena5MONibrb0slu2b+kcrB1hl05ORv/ahGyqPuUDTC+Y/N
DvFu5dtq2DVWnZd1TaMlBRL/NgyMh0UkvbZMG3vnmZVTHiBG4Jyd1VnelXBSsTNM
da+LY4dSfsOAsiypIJ6AWIZO6rnmpSOmAtX9zaQr3FK+t7hs/iGmHtL58WgDQIcc
5weKHVlPb7LCquCxXpsDW9O1sw6HXpEsUQnJnMD0FxQX2Udy9GIqzavbt/epiIeq
bkCQwXGW3/KwQnYwOnmcGmAUCeNmQW6UBw7q19yZ8txzWKoiKhvlKusG0isyGorh
5DmY9uy0IK77QN9IRkPFUedJYaf6FFcrC4oS6ZhZjVTuuStUxCQtucwkSiPXAI10
ZkkjDyQRoiEAYSZudP1BgIX2v7pJmWUGyweqS/WZPJH+M2aUPhzyQ/6Th3W5NqyK
DUlus5jMlbx4jicC6IrwBJqYMOpFNGz3T0UnMBJ6JdRkBYf/9J066Ztb43kvp5Is
sE6kxGIUP/9/R/J881nmqD/U8Nd5baZpwJFYBvRos1xcIzhTLxFnOFT5Vk2hScpX
41AOiA6l6djgj6T1W39W2m2oemhaEFZFDIEzZf0pleSWmupsfDpW1ok1sfskhJPI
HlKMuNoF50jbhVpkdRlmYlpceVTyyb0VYCqHJ9VFHr7T08N+M1TXTaA4kPlKXEK2
ZXwwCc7PQrWW9tGwUeY2Wc45B2oL13asLhlH9z5f+TrRh+fjGsA2QsiA7BMVL1EM
tgWYvrIY2QEnd5Jvd5s6qnr4R4ZKElf77jGNNxSI5BGkzkHXmkat1c8KZV/FNtV3
eho52dnWGfCN5856w4awR/Xn+SbQet5a4wvz6O7BPOSQasSGi5lg/rGS2FUVZCOO
Ef9+tpoxszbsbavV0gBBL4AMQM/ZrErQJFz/DZssmKHn/oMIPY1en2lDg8aPJID+
7NSWOX6i4+6zNgTwN+5Zv5p9PUd7BQp0FGJRH7Ez3QKabGwVXUdaYypLkl0N3trs
jt8XFe9s/Vr1pYLNhB2yiRNKEMgWxMFEjjsidSrDm57yUL9QIoUrZPcuX4nJCMF7
vPnTVSCYNRWWURGq2V9xxyXhBAEm5JWfoYfnXdL7P0+4/HfV9eVk0668VP1LT1ad
39B3nFDA22LaFnYw9XhXKiAxtacJ1yYgZI76dYDPwyeMsMVgjEw3zSPWgGLq2syJ
KuMiXUrkSlKPSWV68DurkybYKBvz+7EO7xyrWanyxhS6yehnE9ib3oMKSymTuYAP
/kn099JzEB+V3200rTeI1CTOEGrHn1uVzacbJa7B3/+7TXly5ApxhS4p/S3tib+z
GzBXeShmpRM1eXVa1nQxO5ZFqo4Tvhdm7WYvaBTtnJqAGcla5FUgV6VdcccomZcv
/61EqaXV5UpWsjpa+Z99B7QZ7Ziuk8CXPZKKEjFpPHeXdu7eXVe2gugHmW3ACkn2
dgRUWWQQ/e8okcqVpWWdNQnikS3Lzc3Ief7BKzzUJOw8/j/lnq5fni+67pGbjGlT
X4GGs9OEFN9xzY9pJ0eKN5gtj44Vc14sLyDAxeM42vsMqlPUAzBkV3763jZZK4ok
tbsEdqwKBdjV6E3J3ZVixNp3hoEvv+5F6Nc8bOhxFk4Cmkr7shnbqCg3codlI/w2
8cTHlqk5Z9TtTjDpPZR8nkJmNvV7xSVjGOAvzUbF/EVP07EMHvyBmWvNtC8ckkrr
kxHASewdAWDbhlZT1ugnLeYfrXsYt74djdahh4IasuHDp8ApEUgm+jY5s5WWrNtJ
sNX9LFZuFF8rvaLTMe9K9wM8F/fscWvZ/nHGGprxIk2lfFbHL8X7yHZ6DO6LTeZq
RB+1QUsPO8OCAPGmyLEeL738YjjNrprQtTh8LhO8NqY5Q790yiZJuRnrVsrN1VA3
wwhlIp/asK8PcPoee/SXjQ60L/9XoUSzAnhDKOC98m54L+3kHBaE20IXfAMDM/+Q
XwAa5uDROwNKPtyUcRSNyLAZV70Nt2QWgvfTw1xS895UwGxuq/3TQOD3Rgjk6lSo
6XQNEppOuLW769Cjc/vYOoIPcMtwNFqe0DUYGv5z18xfJHeg4qo4Pb2CHWvkhxsj
sqdGt5BJY+dlJwdzNPqVTIs9vDmfHR1l0mwho07uf+af94fXDrpq0vGJXUPYv1W4
VJC0X7/XHdlz/5MqA6cIQsIO3fdpzI/T5AegfCCtu/3CK/a6x4+sqyqHBYsDyrsQ
LWPvQ72gPpdXvWha/u/uCRrqbgxd3TC/vfjHoGuj+9hS5J+YpJSOmrentOd2CMUZ
LihDqKB4a4lFKfJOOsnUrmecZcIlwy6A6mpu67L6zdz70YWsId1LdrFIUlJwMfSq
Cd6BKnFG1bFSRpLAlinHR+A0TlUjFoYb3+ukQYN6TGlGbJ8qqWGlRtGoKfdE9bo0
NFHnjk8nlAMdG5OJpTqTXcEJd4Ppcchz7Q8FJEhU/TgEAnWlrDc1F7WjaoArYtfd
+8+F/j7byypApIVzdufrBOZiKyH31aYpBN8anBS13b342k41vcs3YseR9uD5CmSJ
e6MYB3MbzFLlwRCB4oJP7FqIw+2VbzaCWxLK7MwZSxqp4RdGYn1ixJRbmtOKrR1p
iJ1fFbV7ebejkHFcGINVdXw77iP96tHZTRQ8nhSC2GBxhCUL5tFpDMBiBOFhv9/R
41vISMPbrKg10A2SmH8vPbXtzzsqopwHX5fPhmOlrtbPHwh43osCv00Ey3SaL+YR
jWaB2kdfD1A8O7du/2S4L6lk0y4BeIag6rz4S68QESzLMdOCgHy8Mpq459sJ5sI3
46N6gOEWhTTKdgGlYIBLRq6L3CoM0MvvjsL+wHCVdBPKlBmBbRw4be3bjnLzuRoa
ykFS/HBPEgiLN7ro+P6PYZwHlE7rJf2L2e7bmdjQ/6KCAyugyFoSQWMYYeskvO2r
UngLIZGtiqiXHXt3gXkff4lMJFraqUkC7mxdYnXvBJjEgzMjh7wQzlGqM2slZfik
EZoAiflvuxuc/ANy9WJa62gdsLd9KaFOf9eCb7JTrC947o+6eEDQv1l37tQp4sfO
vmd5aVx03SvrEVmhlb9kOnOKLuekDvrWlEmhn+lJIGegCf0O9UNk4KovxR+ztNK7
QLH6vIoBVsDdIoQRNou4OiCpAT8XoLE3V32Dd9+LW9PnJQOFQeUYloVDV7gA38XH
qBlrP32cxBqhUqlIO3EKJKCNag/Ex9bYKN0/Urch17n0X2XyCjqJBndLGBB4mYfW
lW1VrbWHfGZiu/AS5mxgjlboX8336ikEuNyU8ic7gZILdd77BpsdETrBdOj5teKa
6pMPeIUne446Nbrxi+nDh1hLx7dJ2qcftXs3rUrDj7oPU2y4mxX1LvKYYqHim+bC
+NGHGpNUke+jw6o2gBDPU9AVYGW7RWcb6PffZXaQaCZBEU8IGKHqhOT2Y8lTNSXg
TVXlYVARfLjvv91/qJryzYQaLFHlZdRTnNJpCyLD9aXMQhk/L38UtCyDwDLo3QK5
1nWEwOmjL5ECgRrY+wfx1gMLllTYh5MRL3lxbYuKCous/B/7Wa/nKnM3Wmo0cqD8
HQ/u+tuiykqTvqymlw9+mocM4bWBhtX7e6mVWmJWWq2nFHYSAOVGh6ww2eojBh6w
ip3va7d0wt3Sn4QA7IYcfJIqs8UCMyvu+ky/2RBWxy5ePofX546QXWJw3vF8CsWa
Tq0JVRZKq/MAaqArkRLfDRML+DePgPggRY5dPFuVb6XawlO4CkAXAzP4RNlE5701
hVGLrlSnXxdo2dfp53aIx5UOjgszeKW2bXptaxAi12sv2vSfalzQ8N/vhmxXYede
iV9b+t3C/nuZzEKw2Q8JM3N4Habf/T7NtYH0cNt/QfOKByD3kbw4o+zIttsqWJE6
Z2zvX09Cg/73Ul8jb1WeXzLE55tcx5eFBhPfacWrOAu+/vEtGl0qcZKxeXTTwmRf
/Z0EuuNRQEzxhQ24TPJ11Z39dI0arOa+kgPbHVWcMJmSKbGEolF1oByPcH7HwfBm
Qw68v/vVItklji73IQk4MsvcRVf1alI4YgyYh2rxrDuwH2BOrzNhCttfP3qQR+f/
VpHJ/AcfKCatpI166P26haVHvo/vbRE6mag0IJdsnZD/fBNcpNhAF0aSuCGQ/e5z
QOk7x7KduwtORn9avXXhdeqXAU7q40Jsknpjfm9OpJaFtg915PPgOrfsql+RCEm4
9Jb7Jvd60mKehVpI4G+MJCsX54uXgIoeOyyHDvVwUEWyexsJ9A4e1sCjIN8cmuwv
+9d5H5OmZbT3qPJTLAnunqnQDTkP/YWpc98tojjYYhD9jNedC5Zs+mRiL72atRSv
vTfYlXSFaafrvzFu8Js1HBWPv8EViFx6cbjpbyWe/d7zhfj21z8L4ze2UGrAb6NQ
9T+02UzmsP/L5P2ieWYJan04NyPI/qaDed6rKMU8373z/B9M1iquUKY9x6W8Dnf3
6nuf2mSVBbyA36FQb4MbLFqFzM8a7u1oAdK0h0jjjw2bHSaH+13dXT5XtB9wkpOE
ZasU4+7qpyKzSH0uoCAdFZsVjK5MUJ+5vM2cqWIpf9hqqcSMmoe8Qjb5fA8MNMp9
5FmdnCW2/eS8GB7sjvI29klA3PVDI+jKaQoRX75q7q+yl+owVtRV9usYkkz9pHB9
EdJkwwLdHM6hTmfBwlhnF/u5ugutchD6vzm7unz2W/EIFuW+wBGYQLc0T4a3Kud8
sc70kUYIDg4AYRdlrKZjxKX5hQTa2jZeyeUtv/z2GGQNWjwCCm5qJLrLSDnFNMMr
n8+yrlPfqtA+O6OdoaAwxKl7IQP29fEQeBwZHJUZHs9fcw9fibYo/1FmKD+6yluh
HqXLrRZyWgXmws+2aSoj4AiQYfp+Xmim7pcdn/llN22lvLRFIK2gz9frqeO5FSGv
JzRTjli5GORars9sQ0tgKAJDVAS0OQK5YXCxq/5/CzlzXRLfxnqMoLFWW2ib/q8w
rzBAGMjAHks8QxwxuF7pEkfAAEYaqg809F+8BtfJAnvi4YvoRxs8mAUX7LlsSNPn
4EYywdxlWqESH9FsnZ3R/u9Lz++ST+4+cuzpUgLUZIaVy2TT0x+dRVdmEdEc/s1z
p00A/vMkVdRx8XjHGbqYrv06gmtGaNNSbs+Nm7ibrRzvoXgbj7f8puIm0W6nsdh7
lKPaksbJ2mt/im9DUjLXBEDkJbFHOnRP/9ior2sN691Y09AAkrSTTJ57exyJY6OP
C0MfqjWVhMTxJdOjUYBjdG3+atwLiD68bs6EPMMEGlLTwegnfzglS6YK7aPj8bMk
7v64MV2ADjAkSlw+vsb9EMUzzPgfcwqVkZ3itE8U/3DzwIyp665M1WDy1ZKVm513
xcuPRHFrW8YfLOSTxNwjET/gfh6pAeyaUnJLWfVJT5l9HN8pueb1dLydK25IebM8
RC1ea91Yd+/Db8bTZgcKFoZTnTdZGJk7PB0NqXLm1osX51NftSE/t8eDBl0/DsTH
u5ld95n4XOjJOVAhDuE767GuflK0VpxYlhnN808uy6v+LWkkZLXMJA+kGiArcgQT
rzbT4m0hgnhiXi+KMhd1fzWJlOdo9r9OLwFi+DdZVUQCkx9tV31K7zJod5SQ7pRD
GZuxMeKZVm1QIrN+TBdnjfQ9crCwOCtq9HOYDYADWoZIGK07fxwPRUIZfNiw7EAk
AkOEkJPkuTYWZF/it7ZIPhRkq9py8NsZU74UxDitI08BSFpiRkCaI4Sx7DjCs6M0
uesGDwQGM0dP/ETmMHU5W4sYHEct7rE2pZJKGhu44a7Z/sbw9uZZeMyc+hC+xlQC
Mp+PTimyEAv3Nx7sghsXEQv/Ib/8ElI5nEwyodaA8MvQIFHH2aSzVSHlujsTD9PT
2RXeCO8L3yBjq+chG6oR1cGIbs4IaH9y9Nn0d20gRT650d0mJTYpp4veLdo6JQ4X
HNEK43zhGOPUd8EDj6syss06Um98jAgoTy8wqiB/KU4Xhx8LgYNCx+ri+bNnh65g
wkDQJp0NAhBNguZ7URt+VLGGVCLa14SsUdcpvnBIqgzQ9mie3ZyV/APlROS816Qu
FT62AIph+R9CSuBKwYItajqMCP80sp/UNWV/N1hnVXuLqOdUexnsRksfPsySaDCB
XZ4h71dGVRdoIjBD4/WHiUESimyilwc4knnpqy1W1xUvaws8bbmMkdlbSP7TV6tD
OC7QcLxSqYXxveasHPcCOVDZomm5Z+p3KDk2HxWC68nFWDfIiZ8c2XbaUC7uSmJy
an0O5CyBsW9nFymGwSoZTQN6GzQk1C/mMDrSzPbB+7Q79u0NGPf8v9sVItIYbyah
CRg7D+hFF9m3lyv30we6EYe8Mzby6Js76SurE5IDon5dvOEPnV2RhoTlf9pN0MG9
X7AiOtrLT4zr0zj3SyaD5lsZtcCVqkHwWdusoBltn87mL5NiW1mGGLNtpfhuUewP
lTAlUjwa6sGI4eFHdWqHZ8KnX1L0p2aci50adz5atJFlmNskVikPuuhOrg2IHt/A
z9j+4A838zGYGTbh8AQtbf0+DocdjtN2YcKvI5ahPZfxeI/Hka/t/fAtnxQ4BxJG
1UX1sqS6XQcWNA6K6TvrYWGP6wi5slRYSYUiW9FbOcTJl5yHcXARiLdrVTMX3//n
98kKdj78pT+C8iJbzm4+Iz/F2pk4GGkW6kQmDPc0Up3L3HJ4YuG0y1VuH5CukJmz
bafmk/4yxelQlwFLZHHve1rw7ZYg23fhAb/5SbBGzifuA+T91RlK66NknPtuMLgN
03j8xMuNEA9ih6N1YSNFZb6cTFGBnxPVNPcqFKgwyFkBes3NgcHjNaqfZ7DHOfOW
MhKnQBNB8e5Q8zdFctBz4LjcalXGXOFOgvkfrfUq4yblT2RH+PgM4T4lUjs+kH2q
muRCxs5rvorL6/3u4qzdQhtreB+/qw2o5tDpOSnVGpZ0NL/Wpz7wUD5LFjBAqkuW
bJQZYTqhfiF3WXTvcGlhmk3K3FJObEmIpMEDPci98sfw5ffOpgyGZnhBbUN2wPFt
BRu18eiXtU9I4UcqoQHu+8zjspVl5w0JEicZLqH8LBmXGS1V+HSPjWIiE9VTC/Wb
QckN+lIpKCf7gaVwbfCbC/1rzxGnEiS2SzEQYBAR3d/rcTT64JVBExMDX4QXC5u8
eayJtenLkPZ2kZjA7kvdupws/Fhu8YzRFLqf2wk24HC1lDWTcVL0YwM9lw6FRA6h
e/uL+jrY2W9u9zWj9Phu0lQ4f7VZ+kIfZ53miErIIuwK7eNC0zfSvxALTPU/uj3n
4356jIyyGMDodZ767ndQQMfc7FuGLbJZMfVOBcsJxbzUho3dbLGuMus/hlUmsQzj
IpB3ECIvj/YsFBgCc9CgwMapvt1rKH/TDTaSoXqyebpU7HLpgKTK8hia1/F5yVeG
ls11yil6I3XE50yc65Rbcz+BHnb49akvKf8qVtiEMUFD/6EfVgSh7yXBOgmZF9In
5V9SpdGKEku7MyWDU7x6JW8lSDaSyzLyneCA4ibPrNwbMJRdxwLYSI9iz8RgbM3+
aLGOPC+ULWUKSe7wzklbSokgom8k+M+D0fYvrFFNumpwbd6AeIobIaTb01agnZX/
B2YBf6i0XepKJOawdonsF5U1vP8YVNQhif3sx2IseMfaCYTJFnhCHj+M8cNbfO20
i5k8ztezOfsDsnnEgWinPpsSxv4D2QW+QlQFv9Tf0SC8qQlQgr1uGNkGSeIagwmz
WqHtKep+sR7PPaWoWoCogZ1tUrZEVvX6nZgoAbtROPPS5f0bj4Uw9wCjjlBwEoJw
D3fYkL/47B6Qg0SJJf4ujIZSWzEIxIpnj1CRk2yGkgGLyKBY5C2yXPlmJoDviKQ+
Ewfq4Ocl96teT44ELlkx1OEjuV5ysDywSqNjK9xjx894nFgFnFw0dtSKT+IdhBe+
LZUVOqolAF0CPoE/JPN+iU0XlabpQSrNVAyTmi+LVSJfg87PtV32TQOdNc1nLWV5
TpWGLRMrqjcLB2kT5txKtvv8M6GGrF1TSVcMriFcGnOzw8M3TKWdPZDP4m1+1sDs
gYesnWpWgXnAaZMuxvw5HvWVmTH+wuT+3oNYl59J0sQYaNdKrtU6s+IZ5YLmfnSi
uscfMlzRdCSYhMS3RExD1OORWRpTpnRW58vCTFi61I/0wA9SgQHFwPhdtY39pah7
OGjt6jOnRj0pRW1lN0GVKGO49YsHbFVxnKs4zCiVD51E8RJecUC8zlTUHS+Gb8/6
W1G8Z3aFA671nj36FLB6hoIHdaH2RGNtjdCp89wummow7N1105ZuPUaofVbBOlKV
TfiKnvil/nG+zqhJ8x0E2rg4JfVH9OfUJugDDxuOSTfRu9qOTlHqLt3oWbQX6DDY
YChk1lXNBmsdv4XYAPT4p2eBv4yCQmwGaNJn0gxZS5a1t750q8BiZlqDqGvZJSO9
Lkve717wxs6iklE38ks20mOeUgnydl15qNH+ve4kD3/z3BHzIBZtqoh952eXbXHs
RkBdQH2KLHNmMG6FeYZTFWRJRvMqGk+yV35G1BpmsSNXK9V23PD+Tf2S2138ksUk
I859vmSRMwIDSvXsIuuU8t510G8ZwZ+I6q+EzGKSmNaGHi6Wpb/z7xvPy+Qetjq0
enrgL8SqEv/tb3bKyhpPpGI/mbWPHeyxdddWT6U5W7zRJk86g1bC5TX+8osn9/BM
Sw14zeAJomKe2Z+1BbGi1xc8xHNSAJKjzmDCncz0t93aq3hosbpc1+idc38JFn+R
+hfaX2DN7Z8fjCLLGNmUfDytoqUlRIktEn0rV3vc+rHzJMT0Q3dX9KvcZWFfiXU3
2YcBp/QZ/fekRJgSO0CFt5fUMDOZY4GuHP/huGzIQ3Ncmo6TKHoROLIXCcmMwdl1
jsudH24Ldie2YXlIJ6tNEmDnPCDmEcaG4i8GF/msrFoZMyAl45LCY8211ibv+dCs
GRtBPhoAQoesp9eDFWM5bd4WccSB8rV6VsvXv+R0gJsbRxLwaHeMLjGlBDnKEFEX
3IfwxgKHf1nazu0Eeg/xaOCVdHG847UUF5zFEzj/ecN9Ij3nTBSHZPe+wisl4cWy
ni9GudnDyD7VOfznsAIXRL+Ld1/7mH2fkWXa/LrGeo82uIKl6F0BHk2TOwPW61Bx
oYSUARxZKHzP8xIhg4ld2rXasXLN1lCLOm/wcnRCZvpbelxRhvi3SVLuFE7dQydZ
tK4KajRAmAk2GGg9dvdTPPodidU58hfParGoMbpQk1e4/ZmJz+ocigleCZdNPgzH
PWx422IgOvo45VaTWphSXouCMDwZ+0RDCh3hvvyrAVsB8YIwus3QzaHCV6hE9N9i
fHpg0VoGAaYsoPYvhktiIjN1/jSVy35htFe4D/ua2+bUW09B8x+7KRJNFVl6tHXP
yrS0tMF7tCQ7RpLAVpOJYuISMGIOaqTAHPW6IzhSl4bPU4kS4tOMMgjk43Ga1E5H
bK0zkGrKRN/AE9OXcfVjQBWJ/DjdTfrt2VfiXlcNggzTmZj/28Trl1ohGwfnPwTj
P5DbHfn7y/Z4s7DdGYJyUFkEK4HHrv/Di2DM96UzZSvTvZVJPm3Y0T/V9Qe+3j7L
Zv9gb/vQpWHBzXDsWQtbRGTAQwe4AHSb0cdXnGo6xDwqhlNj9tqylBGQlw9accbd
8Oafo1h/ISw2lEYOgup4BTmxjuC42ItXFDPIn9Uz3TjjV37xBFq4zjSiSdrDTfcB
E0siyxG4LGwJ48SPWtWmHaVIMYat/adHgGh07NneKn9jD/vxsLqKGCACUP1r9lKY
vhHIFfsiR5v1CYJgTtS2GMX3zb2pb4ymwjKOfG9KhwAqlMvsOqy2kx372OqQg0+O
2Lz3v4fugJwRS9igJjvnbK5Nc2IiOoSFoIUPvFighL2A6M3nkBdQ7kGbPxPMjB3i
W39rSdJBK3m4SgOOUPhT+R1wSDv8k3psbVBHwxGkYov/XNya1VT7QTa4sni5P1JU
4u5aYa69weG/BpfgDi18bT+bPJFc3jWmVx2o0brJHT4pU5CIFOkIYGN/wwJqDhTq
C+3dJQVPTetbcEDa/8BSSK0n4eWiNGZueL9h/CS6GKSkWcwwPXd4uz5PEFungy6Z
hIo/Df4HIFmrv22pXFAsRZEC7zdoLcQ8Wt7Ka179f4lbL6CsrobQS3TQudCGSwE8
zZ8QKB7NsjzmhnMZkDa+IKBwPYRkUvLfBKqfbiWZ2wgZ1vLgcejrS6Jxo0H+SMKK
wHfZ2h1rgEThHRuQvcwCv2Jq5pXbZ/9wwThO8N6umSAnXWPkH1rcuPfIFoNkQzth
MEaxLV+XE8kwE1y+NPtAgb9HT4ZbscWRqnDbQz04O9rT6anPQAF1aFwlPdnu6UG+
prW3E+3yX0lwJWCgm4OtZRAJelEuPTfv0W7XYKF4344eXFHluXA5OxZXhDNXUX4D
sWc37ItEhiQP6hLXj4Zk7ZBGjYO/tfRU+JxHnwlMzHLGpzpckGbWsv3yrKMhRvgC
A1wcSyWLGnP/kljcwwzhac/SR7HkNvcxc7C5tb0h58l8UplDw01nQRDFvCe5IqIZ
H/sOfFTemltTEcrKq719ps4F2W91UhnuYdXu1AjsDXz7XCJ6I0wsmaU4+4yvis8E
NqXuThCHsIPw6bF+XUxHujOCec5gCAFJKj9Pvik8ocuKlFpWFcNSE60Qn5JVULvP
2x+/bZ7hPMPP2pYQgNnQHnToywHbRln13l1PySwKeaY02/2j4ZSHtTXWHlyqdx5X
TX1gxQ/PQnVdsom+y8CQrIpLrVqSwKMfhpwHo7TrB52ZwjDog0+pk3o/U3XwU/59
kTndIpc+OHAeEK0HaWtZNNUovMr5Dy9j76o3YNJllYhq53QRQC6Mh2UJvs5KNUGc
H/RRK7JD+hSotGykuv2daVeec39Hl9o04m7STH+miqYbGtmjxc2mTx4i/uyG/p3t
48Y8Gap+rOrEVLvUdM6VEZA+jUYti/8oZdjD1vZjvxikc9S8c9UJ/IqG8WTvdKSS
eOjZMs9vCm/3GUQG37tpTlLLmbnfjYzRBbE4f0yz3xY3hpccs++8rlKH7SSjBEv3
z1eNzOzmLF+CXB/mxRvwFF9tPJdTLDuduCyVdTTx0u01oOZYxW1KCLo512cxhWe+
YexmT8+dbuQhlEK4c7IC4tLmJIW7GUiQDV/o3J8D0TUiHgOwjpLkTlF0sgl5SuLV
CQsoc2zqFYkxms/gnjSdMhEaLSu/HxTG4rZ9NeGKlhw9XaCIllDESvIx3mWRDBXq
G9nGO6atZU5Te5lGk/5HT6TxNBG2xNuZtsn1+6A0J1OityF1rtPsQh6PbWjAt8d+
2G2YGEn6LYluCx4HGi/SUmFEIAK0lwVIdTHMUctFVHbKUITBuTTdOca+qy7T9LKz
rknMgMQ/j4P6OgzWzrKQQaXsTSa5wue5aQdFyOmLsHQu7jYzFlYQ92kx1khq5W6P
/RS/p21LVS72FBUsE4zhUU3Wl3aZ7NgHYNhYSbTbrYewLeHDnqxLefvvCq/rVnPj
k1AOdaTbx3vtzQLFtAMgADU71bD6INcUPXf6nT0q9woSGhIVqwPYJUSGVpTwI19D
1Ii+Lch7UYmM2yNtEBUMLNZ8Qvplug/Jrj9TYXdjDgvCi5fxOAfzBMt5ipkX6e1F
MR331wQK1iKXZQtU4fv0eOYCZ8AdwYcgAlocPh3I8DZwzvVg6RlniQgbpyxVhYaL
TnO9082Ot9advh91HgbQGqDWgCVgHT73RaNeBdEkOZP2FyhkLyCIFZy0gXhxL6db
cGNDMxAU2V1Do42CDGBQ1ZV3VQsvQxYB/tA9nW55ULztXW4sgpnJd8mRnIG0tcFW
GiWmSLGqxKHCD+aYRhmCdEOk4xVisGuIKZzZtZPKUCphJ0YelIBK4ELf8b3WZvfw
tpXKEg5W3BpZHRNM3zkba7ZP/YpGu3oF1ipj8Vl2czOc5BfkH5zb7au7GdiX+H/Y
0JnXG/3X+HeYbjy/hVFVkPNvRUeo87Hmw7XDQW4gr949RVwKXq/DrBFOGRz/qpOJ
5rK0JtycKTDHEl3aaGgA+wJmJ+hIN6wvHQSiyNhr6OgY0J3F/euWxDPc3DFxVnLb
YG2WEwLtbOKqkIysh+g+ME17GvltYer23IWB03lExy72CJgoQAuZELrfh7S5L4cp
tN3Dcb29bv8uVRkbqdC2cvmGaKhhoImlc1wnno61ySzeh/ao2qWZpkj2NNqFRO3j
yNspHABt9uZsUT/G3psqEdAU/+JVqDltDF1QfZt00TfgypOxTKPTv7u/9rPxiRwZ
WxSN2BGfGpWvuGTtHwrmRrlSWOHfL5EkI/A3eOcWwQTtpK2ai/49X7rTxqF2VlJp
ViFs3dcPiCBPDk68JKJt3PwsnOgrAvpSqezXYPz40qntHFzbxE4D5SnBULTIvDjk
Kqu7ZAXpgFhUOi9Tbnksur6sNBQjTQpvHxrjTAQTIXuMx2qSRNfwR3n2ri37dKRO
CJTzvkIH0/5lztHb2iOaL9mwZtG44yEQp6rNrLntth5rz5H/GD1dC5hYyIxh9YPp
y9OV/sZ3pALyK4hdfL4Vg6QSu8NMIMoXd5nj3Z2vwddGz8byh8DGn1HMKtX1pb87
LXRcG+wu2hA724DjT/EusYoz7KyHaOoc2l8rvE5nEYMbCX1yVjJT3gTxrltCQqsp
wclIyLtFcD1HJ7Potlrld4mwvSS7JRLWsTfpMFFbxdjlweER7/jH2LYvVAZqhaFk
oK3T2D4UnZC77C1qnbdmPN1syIROy+JHHSnmhxGlXt12i11ArS7E6B6inXwMxutD
Ckft6bIqlhvyYZXkMfAA26QDrGQBYFWOYzUFhd68khlAUp3cgtf826Qw4VsMnR6f
Kb9KpTY2wMhDdJcX3qcn01GhkY+Ga2iPSsFzWKADOOB/FSpLzG4uIv1PJGr7YM7k
2WfiepCzpeCUCpaL4A02qkaP4HYUTglcgZhTu1O6h+emCdEtsTnIalGBFM/j75rt
1E4NS7YHh2FP5Uf30t9+9R/i7zY0ALNQzP/hGm6xwbStutYZWIk4maBdQsgmURGY
+H7GHoqA8OwRSGHus9vnlYoRXFqfc+1xtPJxT6GjdPkBv6zxVshQz60B2VJIQuuh
BRbaUf3XUnyorwYbMjOIZMb7w63oFnNe2NUuyn33CRcS6c8brr4O9bl66tz4G/pb
PnBWixniBo4jUvcsVPVuxBWvt8yJ3ydMUTHyVagMUbTo8fasY2RZqRT8yB+4os5B
uHUuRjft+PsDymaAkTraOqBEVCop0CsUXw/llCxZ+UL+I7s3MbmUSDXWGWuO/+3E
vD8Hl2eYddqbqVE2s3aOHV2E1jwsCXZW9hj7bUMLXljmjHUtV2FJCk/0ruzN2qWv
peUstsQnm9dtORsUeW+akmxUJB+3oWIumCPzcw/EDvvG0TyLy9uitDLGXhSDsa2M
2S1rWr7DEyev/AVR7kC3hdhfd0pnFVGrPkDSnRciQkwR567ZY5jgjNALyCQ/0Ggt
S0sb8aityRevg4QpCXE1cNa9rAaKGpmIni3mHJ+sjH9iEYKtVVx6xMYC0uiASt6j
4JH2b6CfT/b6+7B2c0p4fixcjP32ytsHXoeRB1TNXPQAea3DoLsY2X67KCIWrFzx
XG2KDh1figFvk3PNGtsBe8mmYzG/ZNhlZGw6sDDMBmWQIR5zELw4hVcrZWN3auCN
M9mNibcEvc+HxV03pW1I4Fo3J4JQPNjxR1PJfu8FcecjJ6oKN0JY81yUTPNBCQZG
9TFGWeG/PY3S6F1ByQyJ4xjED11XFCuzfeO9INsCsrYnRoXZJENpwEapyb1eGBq5
zEsPMSsLc5xqeiq0z52Ryi+4hI3eivdo1XQl2+OzvtS6tf5/J6/6mjHwAlGbQhoc
+abNIi5dvEtwaWd9mJEGHSveVQs0091asOHZ2xUV3y6BGaoyefFz7AIff+v33fV8
3BZGDxfuUeatg9IJvVgqMsNnh5y9pOJoCz2vm+Cg7+IbPZNeMRvDIAZ9PGtwb454
cXv8hJsvyEKFNVC4rRi8ljtB+IM7/DnSRsxavq4f8SJv0VXsX9hdO3h9SY2ieV2O
re2Aqt2QXNseQNXrkc6B1boXr8fbuXwWr7t2nHqSlyb2hJlMOJCXike2xbwWPmf2
tk5NhUAbwr/wJ2u6krcco3VNmDC/UfuJiiU57MJ8PM9yuewq7UwoepUyQlRevfok
SPTQfJmXT+Ch9i+xr1kCxtqwBPEpl28YchBnTXs0CA9azGosGxYzLxdWP/NMXYrG
lEjVDfhR7DRxL+ywnPx0MBd86pN/bm0bjEmuNuoke3A6kp0rKT9q8Vj/5TLXSYA/
bM4XkgPxBGCbHkRbVfVV/6D/i5O7HbBy01uipGt516EIQUBhVKt4b6Dtt5dHttgw
+d2RXNZraSdmfMXSC0YG0O0TsOnfvB7aSvtXJNWG+emScnMU5mZ9F3bmCjjZNUD1
GrVZ0Hh2wVoHIO7ff4WddEbAh0eH/sdh1Pw8YEDlFhdmnWmuh4GRejkj1+gNAgdO
z88WRBIY8WPnpoew/CKlOU13Py4BC8CfsENzjWcsRrBCLPTMfqlfvu20R82dnAbj
oDzZD2hJfCkIfIym9GTDB/IX9D55VsKh57yGPT3RdeAA73GhRoaX1ZWp9ElR3oSV
VZOmTDLqt5oxzLXykyWdPGLuzOk9IezGyZzbqgMYX8DM9KAvGmtexeyYcDrUN9NZ
L7R2OXAeK2S1wnKKlLe9pj9jEM/oXpBhUchNTC1BgrRTYJnPQJ+OxCNMUZcGF+7B
/zDnQV2D3l++lWHd4vUUHX2kiTZEaLl8xDC3Bie1WAmtG7XCee1YvbZQsuFq+Dqu
p6ts6+CZhsPmHW+5fg8MRi4BdUtdJR1TB7/JBqCFQJrivB2OYwefm1xbm0OLxXeS
8t7bLViA6gVsOSBHMrPG7DEvMpN33AO9kx9A/ixg2CBOS1M1thUdP219rZlTX1pU
V12tpx0s+cZHlNjc9p8RE4rQP6moTeWG5fcStmMxA2upcwbMPrbbnimDpSL0AcUd
rdqli3Rs1CagfzMVC5Z0mZerlXMKMdBwjcevH3fKWtLiY1qpwdIGCsWq/zgGInR+
4u5RmPcW3Z+GbqgFAoXIZTEGmpVSDsKCsP/dwYAe3Vp3obfanTiYK/FnhuNok6RW
5suAL/80SbDsEZZQFyqM8pPLu/Y0AbEt4MlVVZAmVG0zJJeO2Q+Hj9YaRGN3AbR2
PX6msGMqGhyOMFpdrtz18SIQHu7qXmDnc1STLb7qRrh0IBZrC4bDsNlUwu+FVsxg
R/W1s4qtA8a3ZJ1t5euAsctrypOY4hOYNke5JM3xFz4TnWPGqygKNz8y15sfsVew
8h5D+agdj43J4MBoy7p087ssJrzUcqHjpmABBPTs1PAr05LlblTMdDt3o5jzMWWB
By2bshoWFer7PZZFS0N+703xMdHK8Xg7TUr734CjMURyL1vjEDR1mFt6623QXsxx
fIrrK9fWHgbzVDDhNO+C4GjC2Fv3HHal9sQ1E6AYHwniTM7GLr7WIZewDXYuQtb5
E9vw9FygN7xM6RUy/3usUgBUoY2ygOI0XLRiDrPh5INvH8Kfw4EVSCjnp2Y83bgV
lVg9yRSJa3GOboUYtZ/QPh2XHWYvu11i3PLN5EHbMUiHBIVnyVu8X5NqSDclrp2e
yPbmT1MDNbjidjIB+K+T6Z8BT7/veeT9RVQ+76HmCDWQbxjfYSJ6OVPXZudNEJXJ
1r6/t6O3XWCAjBDxWND55vX8Y0q6WFCzZxteNIXlmxHJGKB6SaWqXP30WZU9kQ4p
wBpRl3s6pC4Tm6ePQ7+NGZaQ3dAGAGxLduDbcoD3RE+cL9gLzFWcysI3m+NR3E4M
e3pszU3cdr8HNjtBiEPsSYMKCOZV7D2wB6Pq7qDPCUYvXAE4tMV0eG+FRakVo4e2
hS0sdQl0y1lqHzGkYx3OXKUftZcgCI1v/V9jJogFdhnD75d1NEq/0ISIcmKJPgLJ
z6ZGBX+MKJ/bUAVDqXnRwIDtMwd29hWQB2VqUDL7XPZxGuR2basksT6GWybtSHd4
lhZW3p35TamWLIqpKvEwJPwIKyC+AtknADLq4mkBCtRh+Tqt3zRJYb0+EuB2Mops
yNjnVYPaL27j5alwGJj32zB8mBxmg9vpaoG+pV1jyX5G8wNkVamPFtyYHehnOC8H
APbtFI7rrpSnkRJnPuGNuGfrQxt43hzZ0p3GaR76GeCr3dEmXFLI2o83rYVMVVl7
qDzoasaPKjau6JmGgkk4DaQYPyxSITDie5zE35u6Cy1KRI4CJ246d4Jla/RYAzld
wm03B7f9p1VPZlycHSdhoOn5lsYad2tvOpSrxubV8cqfqULJgu5FpUnnN6rSMrX0
mP6bDFLB1g41GEccqokjXpMwxdLs6u9jDM4AcpKQThDPh+lffIbFGYxqp2UoB5cU
5/BULP05GQBxYHHBgcb1xFHlGWrV6Rs4qk5FXVRmTpSe/qg8/WY6/lqgJjSSSTLD
PMJQErPEJRyTtZKyNaxS/np9wUcY4KeS3gX8nf+ho//FJAf83GhHCQPveDx2rwK7
fOyIv24rilsVnLjV00BjOL6+WknlWICdyDB1mfsBPD13qO1eay9Lguus+UkaO33S
GP3DJgiaco4Iz6/SwjIE5WZqNaZ49oLQuK+4OX7JqMeGPiVdCsSEQVBb+pAtUuPo
Zsey4ZdmRMtz5lJZd4fzX6UTfLYDz8QYUR1My9lMr6NBdIC+gMcZvRBF57aTvJe+
nAFtx3W7UFtN4HIzWz4Glz7/To1/H1MH0AzcaCu5+vWUjz45yDm9FtB+XBH0DH5s
o2XamdsEUiLs0grfWppHsolFP8eZZ37u9X8n0pTV3MClsMTNlch8GiUPzEYdE/Xi
Fy/2vpwCyD5lOO15OCB9ifBJA0n6NLD1kGy7L6IyRK5zWemXPUEUhRaKLD3+wAYz
j9+fuamkhHvVlaUAXXBarV9iRvlQKD0lS5SEj1Yw9qYvrhIdqJn+jZQzJ0JdCp/j
thYQaThAk4ICyX+AlcBP2MUmBIt9ALLm8KnbjYVV2xpWGOUPVEzCfg0+oPEUJ+qu
SfvC0J0XQGv+wkKYQicOB8ulow4uQnrNBVqqEYzRE6RMQq/A6I0V0WCPMsx9ve5m
z8dueb30C1uk2ylOx+Xe2jdCPFDdXtUAVKuXT7Qe9Dgu4RQA7Il7wSvt7ADoRBML
Iw5nFUcMDVEW/B4/KPsorzXLP4Ut+/Lp9yAVwvGAX3AqnjQem/dpCNzbbPNUap4S
dW+JL8q8GY6cHym794zoumc1HFpHBDtCKzOMT4pNbWs+Jp8zFztgl9Staa9u26ID
bFB1uUCn1QTiW8nnCtyUNLVRBk4C5kdkldA4wt8A/Alh1LM+Ea/0LTJn4vu7Oc9S
hdeCevTlvgG2w+LRB54/7zpjEjMURR0rRHSLjMvHVe9+P1dP+fUB6Zo5G7Fr5XPK
Z0cU+d0OWF2EtWmyRHDG9gfIMJo/h+WO54zxfOVbZuIiRBvEnrmSBaP0eQ8HsvPj
0HFJOrxgPWGEeha2JHPdeWMxpoNW9vdsWR4cbmnfZJcYlxQPOUDkqtA95mVLu5sU
stZv+QdYY/QCGaHftM8uuDt1y95TiOFppyssc+LICE+jEQeyb9CjIrjg1yGa7XZb
49qSZFbTKpSSi4mqnPTjj77Sfx34Imc2lANxB538m0rGi4ylz49b5Zx1/HnH7rsq
6+qkOhqVSD55f8kI5GxNFk03NCzKLLg2EdYGIdeSsyhUggnOlkwA47A+uhHK50oq
YPRaHHGXFvsEhyFhKBZKetx4r0tMN2dU/gHr4S/O4CFj8ueITz3KAgKn7hIWuGeI
hBiksjBf2IU/KA0D+6uyMg/yqnqS+wgDCulrqHzwoc8ce+tiDjSe+g+7TXtya42Q
UcBa6+vlBNPxC0Sn4kMTqsbYpv9e226+JB1xVn0IZz0R+fpUS+zLj65bHek1lNQL
IaZ6La2gHA+mwOF5HJrOPlIzz1qOefF4DJ4IBt7waNCBMexddMttbClA2svxj08O
pPZ0A3mnwGpK7N3td9JvmuICcNyJE0rxdURb8HLwK2ydmz7ZJpjUlCIuH/o9Ubgq
T7yViW9juDtIyFKJeHUml7vFoMa9JnQbfWswtS5jnjcIh50LqJp+F6lkAZRNLtZL
t+F8QSZwDn6vsk5BTCj8TrEojOK74u/H1jPK+5xfkD3yu3P8A8/KfFIkGGHJMcML
Bnqq8/BVkBftf7aAhDaEUJHW4oKIoKmP5ExtCSj75HzA1HIQmtQADh7ivYxqIFdv
YSMiTrI3p2MJwT3B6n/WzBvZmfOlAm9HEFNYYrogxZb3qu43+HQe4Y9DaULv/6px
Xmb8Svgs8aIGrEujgN92jv1G50sTCCXxHIw2/vFofqGxCy0L1Ci8rW1ymoJWmeX7
3lO1rOMha2LuOqywGXgK6kg91vuVzyeBAwU8ZlMXD5yZD0PjJ9wobAsj1F5fKp7I
/1ulf0VU6vwWRwbAEOw187JC3uX3r9dRqbUhnr/5lIecHXfX9gA+zo2QGK0QHd/Q
56RzTkNAzDFOMppskztUM90j9UomlFpn33vJ+6LT9kKE3C8B3gJjWdwPbm2dx2K/
N9wc2qUKJPRmVH0G97sAvCc8u7T64HqRzTOc6nQbEtEAdklJw+2CZXE0By/csG8n
6tnwnR+Fj6TXSsuqkcPXOX5ZnJKecMtF9XVx8NA9jdU4ETufROd4/MRqp9GIf+/N
D8YOTOLJxIiVJ91l10IPw9fFQE82fQQVncx6+1PvNF8k2pk2raBwsbvqTsCjwT8X
m/YT4YzWEAkCr1IYbyW7s1IWJi5v8TY3JgFiS9NafgldbRJFBj6HdXTNPrx48xkP
VnqOZMOkilaWXCc2jpxTw184rFglqXiZiKP8kLGdHLuMtBiNmzrpmP1/5QDeWnR5
+H5NVlkLU1RgDRRYZWhUc/5oem7Jy2dd4YT0GkNIEeEV4Wsy/nLmgCAjwFMEgePH
qg5pwHVhm4w34pdelBVjmnxumPtk6cAfZEncP2hYyIaigworefWLOcUPgUxuMako
/SosBK/Zt8LDg+tw6EhAq0x/ra+c12byOmoamx+WsIvIvs35Q1EOuy9t3cFOYfbK
oZCVi1JyUX33UBE2mcaRTCaIBS6btWpyLgM1Jjj/sNfmWr8vNlvnIYQs+aoMlUmd
uUXDLR3nEBNcrTJGPvYn2YF8vf6P/YJvD6FzV1bQqbJdykSNKJBbuwD1n/Lvs+iw
rPNlIU4Qa7vkaosGuwFrbGT/Byu5MQKjIn3/QII21uymlrACI7facYndyWMbeqTV
5LXYYmaw7W0MJmie2N6kJqXmNvHDhL+7adRT66fVJCJzgO0ZEwFaa5/hWp3F+t/I
MfbjhceiixOPxuogQ3I0HSfEX5R3ipiA3l6/s7o0+nqRLtvR7eFNlcFdEnv2eb1G
yo4txAk13PgqIgdUCE09TWfvOxW59dOExn92+gd+6swXrOTySpFw3unOJhzmrpJk
E/oWbS2iC4OCUbtCX5zinvRz9Wr6t8HXRkfzgNlaCCc13NNOBmiX+oAFN1YpHxhu
hbkuSO+/VzhuxillLoZyiJhRQixD71ZWAYms1ibpmbyx0eJmPXALu4lZEp58DsZA
LVVUGz8T7bGoqBHo6YQTAZXMAnuJv02E2BSTiivXYjGluEtywp8/eExXJILOxT+g
CwQnccvtYWqGvZwxI/ZLyksJCRacxwt4RvLkYexq77vys4MUCxDQcYoekpxtwAfO
Xvmp/e9AqPkmqA/RyzwT3lL8+fm5k0r/RU5MpFp7+tH4WsXUuRbdCyYM0tVQekuR
xnhkI4ARjOh+2MR99uQQyRGgzS0bCjBzXul+J3ZOXfdfa/bpWfFTyLSOcX3CcPwb
OwdoZGs0HG3n8glcoxF/0Tknx/YLBRc4F247FuztWiyVcR5pYP0W6YGhinXEG17R
KWXpMHtK0yfvzupv3iBWluYtQVf0vFJ05ZRhcvOou9t6XBjyg6ZYgHUEtBlhkWJh
ZOjJCmrT8hcn2ZuEsUbiymSU1fl3Uu1JvA5RrKcT3sKjybtNXnhPtVq+h+VcEMIg
NwmJQTld+xJydI6cf22NJBk+4v2qiBc2mq2A17/8tB/Iccq2G1Fu5TuwaD772JRc
rT35AGj+xLIod2qnKNgT30Citib93LFGSIKZL/EUEMk8G6gZPsr1TGKK1PZd2FI5
VWVMeZE3+I6+uP3NX0PQgx+koHe7ibb68GDZrlrvTM+6ZwXu3XDT5hiCMBhu3K6K
KOb9dV4sTX7QokRT5r8S+GqfSLVaO1g2XZPIu/SerI6mmKKfWwTUViLAYPtKsdyc
7bkQEbdjl1Ghw7xCqA48JTGdhRLFHabBycMRiTSKG7HRmnUh2onSvwMUw/JqnWew
u4+jsw7YtlBRg5xm191LNAR0BZPqxBtNEiu8CvMg5n9ZWV+rNQHkSE0r3LTjeC25
zhQvWA/kV1CIk+nC/5uyqcQSl3maLDM6LHsWn7GOCNrDI/dvi6qsNLp5xc5LepmM
jbbBG/BQmdYKVq+n5WCHgRrPtviWq7R+2omFZLeV5/PFkNZcwIycZeOzI1wNzK8G
VP8ZAS7opUoK7uRRcCelBFtVRkjbnRB2yPbIccNNpMSVcHniEGNhcF4q5rrI6hl2
j7lKjzc8mNRgAL161Dk+LdikESCerWZNA8vbPcx4VeBnge3FbrWe/dN+zS8P92yZ
OMdM9hQJL+Z2XTfxa98HMWy0RrQP4U7wkTn64t6O+6L2Nxfpr7vxzg6ycmuZCS9w
LChEiRmB6Td23CCvUwJ4ca9mgtkH5DcsQ6uSaiCKFHJ7NCG8B4fFiRxCzgAvxsm0
moHHAmuBDDrqJcAL62A+iYmSGethZ2Lu/hvHZwMl7Z0+fbT6cEbZ7rzC7ws1V1vL
hwqtbJuV1LJxffuVqlz3u1NTAKTfbYOM0d/W2394h+iRVJPuwwkMJTapsJmprXL9
bQurCZTiF0b09qO1hG2wTA6BjnouMv0BJ2xYb0rMSluIbBPIB8mv8G1auyOV10NY
vmBN5FMSHa/3deyq7gR58uYnTRwOr+e3Zqx5/QqNOc2WRO9c8eDK/3dVP9Sjsafv
plsOoseIr03kkncoOE+L6VitZf4JvSltCExs169OrCNl6+AEdW45dGV7uQ0L0gbt
w0rqXcdSpb7pfCc5gkHIRd74e/gS8X/+H636S/lHXR3ONA8sOOf8n4/FH8L2/sJo
Ag0jPAGvMp0qP4Xc7j0EEJX0rtKBXGmuaP65AfKMIblhkhCFmQxpZu/PTYTe5oEi
77sHe1RUJHcN7+t1iPvyNBwyGf5Wz9sz2j2ZcUveC+HPDmztqmew9gUODzLhMsyI
OwrOqUEhASajHoC6klAHLH0r+7mTktoTOVWBj8MEmeqRDs/lH1hPWWAsFPiI1Qf7
RfrScLNT9CADAWaA70Eotb7EUkTRdpg4JAK6tY9lZrAo+HcipN2gZRICN5edQP4v
UXJTrYu93g5qNJK7FzVhX2ZidUB6DjlBGBx55hE87HFlSJC04uyax3/5fTotMT5N
hSONhvVX89zgyoX8Zg8oNzwNmkYDgOSI+hofGpy3C26SRnL2E4GA3AV9OPRCAUhW
hZ7AZLtnlkqnbe4IquITMTM+CAy3qn92kz7UvlTMde+va34o+TM5RCNSmZPOrh7S
pe3bOz5h3nazO8fVoQJ5nh140cl5//W8gpevQ0mC8yY2GqFqgImUewKVxZqu5Nra
GHze4hK2oEOPs2MtsLDBYRB7Sih8+NDerdIuKDdTWLgyNuNodsbFgiR/hYvgPBjS
O3yMbFrC15hHrnIdf+NrparpprB5xTA5po6z1bbIkfZ9zuqniepGIPOAhBo5Rocu
A/o4carRu1MaAzIWkIIKBCJVBSDRMTkUC/mcR05lidVggoSwgl0oh+EuzdtUxkjq
rPrrfY0apio8CutTcMxPBImJf5F7QKDPLMMR3XKVtwPOtpUmGVSQdf+yMB18wZtx
5BNKFCBbzeD+63+uo5iXx7FdHgOPyo3v7C4ze/BeQhQjOncTAzYbCkfiaey4WEFR
jPpA4Y54R6oHE0sX678QmnqxKQJXHC0S6eHGFjZOh6mO8YAFXxtrgU0lQFdNuy2E
qZiVvHlhmnQ7EM24vez0LiWu2j0HYVmlfnaQDky7RBecaeTNJZYD9dz2I06rJFH3
yTWYACJiNCNnjfNzEOxhfc42g5DB7IzcVjpdwhB0moQziOrpVmhi2kozkKFtS8xE
54RVXiHrZOB7/ZZa2q4v4+3YANrLlEUJFHYYFjZWp9sviLpqSMfpaLtNqYXkxqwn
uLLObKDMRdc+0rZUViegdT5NXEqE4CKVnfqeCIvSsyEyNjTYhICLRm49QVQhbCpa
0jNlvqIJxmSjvSusmdyBlz5SFY2Rxh7LoqJnXKuhS4wsuikBvSQsh0EoFo7PeS0q
0whfisrg+/xA/2gzIcdVyb4UdLf66O27QgNxixvAgQFo/C4LfIklY0/dQjfaLvv8
Gj678TIn38nocVNdIk+kFqNmQm2KBaTES1Kitvx6G2bqWIth9b7t13c/cjdxE8h+
N2g+m4uvQ2pm7AUkA/ePWL8ENmfefj/1mgIEVxEk0sV8G5P4SL1sLzETJdZPdGJq
09Tpkr//tTQOfrh1RSC2TvJgatYWEsCmLqK/Rp4JMWieR/qL4nEgToRrmXx9XMrW
VIHU/41Tb9frdAJ8g4HSr6UsAUGODpK4oc4MUHi+QxKoHXRyzP5v5EKrQksVMlIZ
HMzr+mPRW5f4rnDYLZ6EE/0yp816FhD7NYpCi6WRXO/lhd1om28WFaygO1aP9yYy
NFTuMcw7fc85i9zw68YJA6yNHaaxXFaiSIz1zdvVFXArAJR3hYZXba9Ad5q5U+OK
1Xn3kFYftG2MZ3CDmlDKRWTv/Exwp06zFY26Wguo4i2S9iraBsuYAUgB2dwVEy2e
7OPU7DV+FgOozut0/0iip4Nhe8KtLo8WVIKP0nVw9RZOZjt2XEUmerwDuwYs2gCd
tkW+hzHKjX6kLhMwqPhRv2ZBClQ5+pnBkA2zlXBcKI3t3ZGWIFLWPPQUGIu1lFfD
uJwmIodVbHfbY7R4i3B7/VnkNaaMhuIYynsz8P/Q9i8+z9bxKv28TEiT9CdmS04B
gugMFv1/hxPfnIW59C0Imtd+JGMFfN0g1Nlp4xqjXUEygGZlx2B1Yt9rkQ02t9kk
TIGQjDPsu19bgBpLgs4RMZTyCaU+YWPhrmHSer2528meXEVSMics4gnlYgPIDrGA
MHMG2apLWqzKDhPzCqNiJgWZlA2eEVihFQ5K4xJypmY3Ne5oy8d2P9gRjdTLPQy5
o02wuiMo7NsKfBKLLolLAdKecP2j52BRFYipul2+Ah7ET5OKAT08xmZ4k9DHCL79
azdmFDF+VIn+O+N9kAcxdurt0m3nyE+hhFuL04Tko3ye0srd4FAiUuGTCHBR0Q/q
Rc/9IZ2hj0N5GCdy2JHK4aPSqyTxMiVZguzuEFXwQ8IEb+3qMtCaIEgc+gCWyYZI
SBol3t+Ql1QJlxV14kFqrYZ2eS/6ynwAiNDswmxT0eVj9iGB1nFm0gWUKDv1nulb
l0k0oSK6CuGBaj5jtjjXyt4iSpWJ4k3FhLfOvv0xHgOiSqMXoGg/9wUuWyoys1Yy
8CglTw1/A7XyXwAyExTkinApAD16Uk0p5LoksxOuLouH6zAyWrciH+pR+9dPaXKX
UxGbuDthu78NYFAmA0PEP8XsVJojCBHGA7qUm10MpE42DVMFkt5qRQnGE+RAbhb0
HApRRtce7h3aHi4kYpjTNTUXm1fNSE+lLyeAM+C+ctfQ2DpAwaAOEj69bJdYfjzb
3ancSZGfwQnKWela9JT6COoHR/ziDrhtGTkTldIfMlhOLzwNpqB3WTGK45ohgT3o
OXpxe2bS95p1LLz5uoErWNnw7Yjo3JA/TjRI+B8YbnG8Geet7qi8im4/aERwlAp/
I3yg2lschTEiZzWalcjeiQ8Z+K5h6/la04y3tG01IUT5QoCHoi9ucL/lY85V/3Yg
TnGah8xBd1/jDtHEMxiI6aCb/JyvCj/NCIKH9L0oCDwpWxqIgPKo4Xk08KU1CXKY
Q0KN/V5iqS+ZnQv9cJ4mShrHSKTbEQeabZ/orgDWrW7YY6Us1wHhHDKXbRJzhiP0
Y5NbtxSjTDUl7RHHM0HMfpxtPjtcbFTqT53j36RIghFXFn/7wL1buS06MYiFK7Se
HA2eK14NZusnQ3lhypmuHuANInmIef+rfNSeeva3X4b0s9TsjJqcD4Eq2r/QXD4k
c2OX4Cg4IV58U6jdCqF3n4CrhJZKhlOrmnepg9xfCo8jOHjPrSx3Ko+8SJy0XIFS
JKcp6WUQOuyxbMOW3769nGNnbCddaZqTrURVZ+UHiKDT/vF61kBSNAtH9H25Gc+P
YzNKKuoZKpo5KQbZxlXMJQzxTXTJxZ407vkqChfNxM/94ajsdPt19fvhnK4Sd8rv
KEnnuAg0xwnYu9OWaWP68maybLxBW4BLc9bTR/U0hgexPu9oB5LrUcKCA+wHJO0X
I3TDBzQRdpbmCpVCubOi/vm5rxL4LRucyGqb4G0UJcL1MfE+FHpaoeXT541do4IL
EiZMirkj+/KCNi3U6ckiloqBTwDBMlvIzFceZMF4jGC3VvwWgZxpKDnMlXZJ9ceT
BVqN660WkWB4DUiFNl+PcnJJ0zFT3ECfyKKNr2nAagWMFdtfU+z7zen+2g2vFaCn
JwfSg4UTMZ95wahu1dS+ywsHg+h685pjRHscze5tQI4uU1/Xw8Xx66UsI0TNVIRi
fCSLe2HfIn5Uy9C4gXwDNxbjJbHodJLR9HnmWBXPQtOoUEBjUp8Gb//zYL01h8yj
IX5H3zcvViYqvzIlr+H0zqnSffxbuJz8S0WIxOqo4BbLpRf+bhyQ16PFkONUARPO
uVzFc3G5jQsSz3A/RQBLDjty1nQzJ9HYShbXSsYTI25qHpYU4R4EQDdhdF8AfX6K
3jOJMFxLp/I2Ioi4bjueTfJJ6PY6K2JIeeabUCBs50oQ3fzHJdOV8bIU9jFlve5g
9PMQGctM73+5FdBFRGiTw89990WufRw2eevoUi4HSebtby8pInRp12LnPYns2ZP0
xw1HFQdoP20Y74RdtqUnDSJiFDKShQweNDU3jZMKJFzZ//Afrv9AtnahubUBUWc8
DFGDPUjxs39+fws/SMzisbrFY3E95lROAhqRBrHIB6aJBgMjvV014WeveYip1Sgk
qzCJNE9KOyRafPOFtMF6S/JC96glyLmK+FjupxaepZXVNgxqwtkuerXXaeeJ7Vn6
dQxa28dEFXfSpvWS6kcs0ySbSKWsyDYrHZ7lznyiJ/aGjaRv0sasU++42Ba9jR1t
f7Fb2j6sU44ohkXe5aFUWhp0nh4E53qfZqQq4G359ewtOCLmBlSDWl5utCjt8G3s
FkJijRM0lDIUl27HFJLcCkDTGUGIebNz6g90aGsAkzs8xMijED9sWSfoGuLP8R8b
eXo8WIzirVOkm9SzlzsP4D3g5Zz65yaXG3xf3zson0UAG0fuJHc5ELX999gtUYln
+UtNPwC6RTRPzMMb9WbXYK6G6Nk4wIPXk25B+Gk74kn4CVW5g4TIVQFQaiUqTXZ/
4qHYT8GlbRbKDAUACOwMzl7Es9NTDp5FRh9Fj80Y+O8VTAcY3pUNNyWnrosoukvC
Rww4iBJ+xW0KC1TQxwEwyZbzckezxk74jzw455DOADerHoFgBgTVVu07zYGtUjKi
YcHIW2eDpMPh0W+lj+B53LxxGbdyN1FBulysNs024G5IydsaqinxauBRrHIy0sdv
xzhJBmsx8RISP4NfoHLkG9C2J2PpBfaebwEwXZvaNH9u6OzKoBvkPanWXSZVJdWf
bFbjz0e3u4aNmCUwAct0aHfoxnev2Gfbl8FQ/gYIv7u9dSo08Vt/93Mc1sJ764VA
kmOS1LnpvyzWobGPTOueGxg4UqXa5wRWgFOF3Hvesk4RGor909eRMCCAnuuJm1l1
4hJ3zuOw7iVSdbsjhNwaqnY0DglOGr91+H0dqL+13HijuCsPLmcaZXRTmoMxvLN7
Dcu6QWkYOUDyKCzNMuQ8cq9cc4KYl5bWH02rEeOBg3OLcUWgDjss6YzNdmqEou6N
kqLlARYCLnGTgFpppCz5UKQWSzv+btVcGtMaDZls3FLPpeMiPWMqEdvprx5uzLFS
3Y9KxdRKKPJq3UZlKrrtYPcFxFRXYI1L+vefG20eyFKTx7HO32B304hOKZKPazCP
SVqtsD66dqguCvjEghdbPhfLvg/jxB6Odvfk88hNTSQqZR+T5Nl2LccXqRLFvPkr
CMpmnuM9cIkUWNLB245asDrk7YW98RPFxtv3ejHb4ucN18R8xv60tc0+6+hOsJPC
Lzy19pKkwtL5FNsaq/wOsUBdbk7Ru3cVzXNc4YqVuDxTGmqKx0ifUeY8+F9rmKTF
GIKN9k/WtUVaTYFuxdyyZGJXekoWq5cSVL3jztxMSmKmzrU7eMvIpqHs69gbM8/x
jX682lHpP5AYQ7pn8QvvQD8+f07ETk/KKIl7bIL6Y3sfkfQ+nweXvTM31RBjiUJQ
eQ8dw5q7WjlxO2MTkhfSXzLuWwYLrVwcB+QBIdS7h9wAA1fuW436xk1rDbJMlpQq
rtuoLyFcoVxj9Xy6Y/IutMLo4TiFEQxPXscT6Ra9XfeRSgfHkn+HdRH90wDd2eCW
EcbfT8PQHP0bS5irfL58E86IPUgUUGzklHTEkItb5hdw/oOFeZK4NTKEIG8nKo+B
hfK/EKasyFP6awe28r5Jds6iTQD9n9L1bPjxbQ7exwMCF8C3ue36ohzzIpDZz/eb
7DD1xHAHTxQkjjdWMuzFnnYlyY2DhWbiK07VeD4UZccGSUAlN4E+z+ztWslJUcVu
g+x1baJAtsBb7d0mZZMyMpd5AFiAJnfZYH0GMCq4suoJSo1tQLri/r4P0qugYrOK
t7F+MBX86MNLNiUso56VjcRhM5y65+qewES5qxWFhS1LuYEL/P1P7JuOGvcF0faT
2DutYE1U+g8r3mPlSO9BfonXMiMrp32J9w2ETPxqIZZiZorWmJfdC6MmT1qqodE2
dLO2tWXcPs7SEW7UhobEpuAGafrof9gQbtn4tBNLfdsBnoKWyb/W0fBaMwYu/mK9
kGYc0HvLg1w1AvsaIBmjYxG28wXC0qKnXZ024DqAu23nVg2bo61WdEcs/zLXuQan
AOH2EQcQrMAd+KimwBPNGaVvr4IKyyeL3f9lMjenS63FINDIpfLTxgrv8hy8qyOD
XphOpWoaCRQvANb3msYDj8/aX6NA8uwf88o0b5ZCqt5zplj9iqqswJuvvBQW9F8h
Hgxc53IVayIZrXMv2BbGL4dzzx3Ln/SeEVZ4ZcgvwUNXvQPtALez6iSg/h2piWx9
gyjxbuX8qTS4VL3yj5P/XP7cSqOa/XlZAG1G7xQxnapMfsalbTidD3bYq6pubMec
y0kFpb3vVVq5aCzYLv0nCzA+FX9+U6UuKJqscY+gJmnO/m86uoQuoX7oBaUWq73A
e9FSpF3kgxEsl2Xov0xXqT3r6yzGHRlHtzpqY+Q24E21BOlBmdWH80DyxzjoBLS1
Q7taxcpcMQKN9ki6iFmjnYTAY6vT0qgalFeJ72jyQpVUToKTuSkTh+HwOkMFgufW
z6io/5BOuQl/Y9Kadnn0I2L6ZY9uKcuXivxir+Y9oRXHjLmLSg71XEpsvwaAOOr0
IbAvqgFhIzqzB4p85ZQ1kkHik8Jya77ZnZeWuKcTvktNxaIicvklkruoyT5z3ADY
fUtbDTK1EDOCrkDeVsNRob2hAOXA9KPPi8IDn7Ck9fWRXQJu3UmmcoauVF6oI7Zf
t8Wf4Ni4Xa4RPAb0fWMQmn9KQPiTnmnQs7O1D/oOrFxeb73mswwpOAw/7bP2oKFo
E8Qkaaj3/bGmq2/VJiTmzpMJV2Q8/Y7IPkU3BwgLHvAA3iYxu1w9pDR2J0lwBLjf
pN11UzJODRBX2fRMsVj3pZp6Uu5ndH7Ztq7Nkt+Yc/NUtDZdD1DcBQtqcycVsU8e
2KuWmdOR6IPwSZnrN+isAmMamStZa8QIiaUsEOWOriqXlW78z6UrCFpqbvlfRHV4
xuGcXUm/ZfKOYxZXmpHlU2CZ8zWe5pey/ZeTClPNEeTHkLFcbMt1YsiVHKqfjVUh
wnkJ6kI/qy4/GyOtbW1n98K+Z6CrMypY0iTmZfb03rfSNB5RvVY5HkpHx+H9iwme
axRB1UxmayIfv8oKxI2iqJ1rNDdoJp2LsY5tmBB75GC5OMW9rRzWPU5FrWuYJaNr
MKjK2kXBbOqEG0AQULHOYWPDy0eFoKT9FGDfh7vzTaDcgonILAo9lYt+p+L2c5Dh
4ewjN9vB2Li7yn2fkjg3uy6czQsQSdAr2MXNb7Q2FaATDdictzfB0HpYuO592KYM
f9R+SvnaIX0uHLuSlZDX1bEh2gvK1grX8ll6V9onuPNXfEPBgGkXyNaIT403c22P
uNIUKKo94eLK7E98e/vodTVV/Ahcrw8B4TqnHQixNkH1GCj4HwBr1w27YoXUl5Yq
zmA4OqMuzX76c5szO7O0k11DdB/e8DkpgRSXKWSx8TlFMw5PnFZAR2ckgIPo9aie
oPrwGE7CDjiuXZ3/VbJHeB5b9EQEfVtBE8njrpljOe++X1IkQu4ZLCg6mI15Ih8v
rIXTSlCIHVsuxxT7JZiksFBxYxmAcqCHdJpgClFlOE4fMvk7CoxOAAnW30epe61C
KaMeBUFIYwPQfuqh4OXxK3DSPCYuQtjNXVQszqJMM6z+/BYe9f6ABPjj4lii+pTV
ZrI7UaC4aVqdvfHXuRgVFS+XIloebpvHTJwnaBA/3uKvaHpJaf538e0KspIKGa3O
Ur13gCddhhLiqfAGJtIFBDKAFGANfrpob5krLn5mb1oV53xMsa5PjgkqNx03fvli
F7xx1bSENliowCD+Vxkfp2LuGJWvIsDhQeCgk/E80i6dUjP3IkmhRvgUy7Jw1MNx
8AfU6SQrhejUHAaouLFvvl3FcLKjG9RMjrwXY+BZZprXcwVgpLjkr+2Wi81e4dDx
mi2xJ7L5t8eH+v66VOS6i4rZWk1HAIMNO3Ct9p7Lgnx87qst/qpKX8zzTB8/1v8J
v4FEqBjyfBAK7YeLlAQTvIM4pT4OT6wP/FP9NY3A4qUOUPrn2GAAc6jpYD2TwddF
uDACS58ie1UWOK0+xIYDjkf3mgNniyvnBO1QTDZbrdKiXpO65qTCy9yUvHr7Pjad
/ZaySkzTxT2dnQiIEn+CL4pqA5Y6wRB008cB5eTnGnmfdLpJXJufE0Tvd4yTjX/J
EKmAQmDEVSOG3c7nT4yuzfRGIlAF3ND1P4Ny3sJK1VoykuEpxV7aHmF+Z24KCG4S
m6OxuYeQO7Q3OuLEdbq9dENSlsyLB4GLneFcpRgF22HRnJNvmsPVzmlcWa7Gkn3A
uOZlW8W5i/NrBMQyb2VByf+EzOiPDJB/PxZIQuMpJbYnfXYYjOb1RNdrDDaMK502
OIrkjOFsEvgQs/2YzoXNEJZPSkoNOe7xOC4sGSUaLcDTjSRkGOHajB8ZtTRz2WOY
M88Goyey58gG6ZUhN777EmK+EGF/qsyXonpkOxA5mRdZhd9BDVeHYBeeBQgM9gsm
NB7wH5dqrZu20DBID0JfwS10tNUBrc7+uufcPv2fLfGbvW0kFeZbXRmcRfS5O+7C
h1p0wltFY/tuSNukzvVzUrHy8VkGmHAvK+MaOw6KwTkYY8tzCrvFgeNyVyO/UIYX
e5k2W8BwQsva1f4u6t5dHWtZjsh8qqBJI7LL4E/hmup3QfLL6N94Ai5n7XyFUNAd
476lupL4nRoiNCAlvu2VGtuUMJh8Envkt7krHtahCfNCXzSQrhj0ao0YL4Y8qgtO
kmSM7yTfiXMJivq4+NQIhTO1v6kQao9Z0H6RmmEH6xFj7vlcw73S110aWIWtS2aB
n4vfqrDCmsIzKH1YQ4L49vqDCXslu+vSYFoN66knOhvpgGuYWYjDqJAXBSGNNjej
hv2h6dx6SgxkP09EQCK+mM6T57AHsswQ8aPx3LUUjDtXnbBw5gK82XKp8jDNUb82
4hJgVdh0RlOtmcBjE5/LDy1k+368edkYX+WiPMIlwfwXQ4g5PrxqWeeZCEQZUB7F
qVwpb5RnrZxxp50nmGGrpRPELgvOcvVollIpVTUqgjZlcu6wKsn3WEiPzWq3oKAl
gc1i2ZTJY7cUb7CEp1M5sqHfzOneWd4jXCnzNlhhkhzGpYcZf15v2R3O8PrM8uD+
P69/6ldHBdalf9e+D5MVX46bYawBxYnNJNIJxJEqezs/Cj1vz3tmGrLkCIaLLqNI
BKMs1pKkhhyHzpPGmXQrM5qtbUx+QC3tPqroDwupkgupRadHqb6kSyE/A7JoGQa9
jDxd55xOxLzqjEhkWQeNkqjQTvYBrAtwiON1rS4A98xrgfaE83GwRlw35qST7+RA
Wy8ccTIAuYgJvD12KhBB8tFkIoOl2sybJPueVkTWk/bN/Kl/VDfUCoDQsfUBQrHt
MDq1tJ+2Lf0K/hzxXR0G7L9H4q9rYQz/LQkQ9mPjACWHjDuT+fduMMoOX1wFRZzK
YZCgz+YXWXG/29zl4ykjg+UgP7/hTfuVyFjRnyq1ODBwNEFCG7JebDlStKs1brQ6
TOrEW9AWvHpk02Ybn5lruOkVnDNYHYdOO8mMGPxVHINIsFFiHh2JuDbDzHvwqEnb
sG+S2cMdLc0BzmQVDDSNYQDC2Jomm79k28ucswe3B2rgFXDMuVpAmtGuXtD5REI5
8N3+FyIou0W5BC7vjZVqDbGy8yVLplVhJUuc2Axqsjd7XdMeC3PNA+8wm8Lm/fQM
FLrzLP84IDWuUgvbP96qItkvVbwHZe0jMwQirXMGbzQzuNpwGLDhNl4NbR4U8Sbc
jc1auH4axKY4Hl4LGYDmsP20bD0520eQ5UcBwTYonCKuS/S8JUSNIDR+I0jDsHYh
q2Tk7vd0fPV4jISV1NrZrcYfX955n87RMd20M9SolJKQHxb5SNtzF/Z2DXz/ImsI
wT1qnglMCuiYF8kvJiA2/iighb0+GVhfK++bDzEdN/wpzag6eHoj4UkhqzLvJxF8
Xv/Pi5K2fP+LUE6d3MF2bNWegJJup0B/e+xBJ2bDTmJuGmgw2f2FedS2b9bS4cgH
UaR/y2u5iKGxI4Vj15esKAw4kagBmExnXA1/kd6xUqLiXPulhGc7WZJTdNTLPQDd
wJtRKk0PHf7MQrzJWwzWHgjrCdygjbKXR/tFTemJR4e1mfRBl3IdLC8EzriHjLO0
dac8IAMj20hVIaxapJmbAQfPgJQSJe6SrD4C4X8sdKtcK3Fub/rjW/4Z0JT1FbIA
9KiDBUUnc6ajWDS74i0UR+PQIjMvfZGHtPR3E/QJCRErSOScw9fo09WeZrdyZ/9g
MdrCMqIIUaVWK8JBIMt3fOXiKZYdB4F16Y4kNyN8y9YIZzxMg/qKgvfzeTw8hB0B
n/oJsvP/JdV805Q9Yj2FP458/NQMIf8u0uceF2/+GoXdOG8NpueXNOJKYYFRmdOw
/0nHCFZUQ2tveAVJemv4XDUgJwUMR86ZHCIpMW6rBugXTYdOsDT6cET5Rj4TKiIH
eCyzr6M3dNT7JBqrxfCSVZgLPhG4HPt8zVc2BZAXiPUvmick5TIixuQvMYO/u6ZH
VPm9KWCmq4MVgOUMh2gR1cJFYc/oK+TtT9AStboQ8wIAGPoDr6aok+PVhcXcNHyT
MMQ/TUzKZXjVZPjmjWJvnvKej3FpVa5HA4DfOSGjf8CinSYqLSt1O27V3Zh67Of6
Uu54r9PQaRYb74jnMy8xPGm0Z9RQEbfE78cAHv663nY6gsU6wkwsEaO2oFEsEIP1
yf/mp5TbxqqsLm2FC9ZPYRt4vquJR5y0nWN129SYywf4f0P2YYNTFqL6V2q+Axyv
X5qh8+066Ikeo84cWq08WOItXT1URn6JvtSss4SwSBb0jn1YG8wJ17B0+cnvsUdN
t1UkHfqmEeNVsXO4SOeZLnYV7JW/IRH+UWsspZMHdHlQ055dIeDAxetVIZFcpYa7
dU/EiUZLPooQvIAHdrDo3I3xf1j+Z6ckQsa/DdQGT3nmqrGuUbT/dx5WVi6Sye95
6aPf75n7YKtc5dO/ufC70XyJODamv5TLjjloSmEqfH4fx8sxLvr/++8MKdUcl+ip
UB2jlIe0mSGaJgzUkWumf6GjpnXuI3HRJp4Lhh0Ze0LxqN0csP5s3YIAik7HLYUi
P+UrLgWmEi55L5oJDlUvyLFr+nwfVYcgkkd0IIBFoKFZu3smM/T+MgxRtyRQO192
jhJ1uxR3Ru9DgIMREFj6XKCRgnXj2ndjhHivI85thfaxHDTinVvheZJtycbjypqy
lOg1jWL1q0NolU+0jA1TrxYIwQge6ZSBt29bUtkyiGNLiz17K9v5RihyglH80ZdA
pWqW3lG2vDP9vVUPhdtMNrZ3CepPGeLdVCOSB3ju6lOriXGOumkydtorVfuh1uOv
5s7rYhJwy0fYmeioSnwuLK6S9WfRR0NP2GS/Y/43w7j4c9+l/dF8+CPYBcALX5d1
/aqK/a5DaYGOGxdMNgUieK/JvSc3wAQJA9wkki5PKQK5XJ+xAn78/pgdFyAqIvC4
Hvs96IYYf53+O9Mx4rK4RtpTx2J0NooyWZQ+Bcrcpnlav9gqCoT9Fn5DDq4yBHp2
2ZwzF22w9c2VgRzahTxAGN88KOU+fpugsqLSjmlFD2JJ1+G0pZaKtIZBlAngr5h1
+RfVsygGDUPBvuKomN6MTbJSrPleKEcBGrdoJ0FAVGAcZ7qqSmX8dH6pmNG5LjrI
rXjaTSPjWm7I6RcxPGEpr/JnevF4WHHUQAczGdq6NR67GXVIwuJ2r2Ecr7tOuX2f
OdIz4J0VNdRGQ+VCWR1UlNY8qzZ+vxakshg67xZ7n93VLMRAMxoNfBwnzVFfJLZ6
9kXAi1G+vqogczEOjwXOsFPFYeDLJ/m0T4cs5Wv5mXTfj76qWeijp7ajHBGvdVQw
pmQPsdnd4fiowmculyqAifM9UgB2xbw7xMrT/B35ZG3qftFX8hPqYFOkjYkGr3D/
BrP/XPUCQSzM6L7c03jU2MhnXjgrLVAEu1jXcoPh+HS94KZLqtCdRbHIDirWl7eJ
gHW0lzFO8K5zVf5hNctSWk/btqrSyb25k9CU6XxWZSFZl0z+GjtdOalN9XVAyyuL
kboXbSSCNX4TRA879OyfiSKmA3i8ft7WlKyPx8tr79cqNwG98t768yN8Lbm879RM
cM85KlIQ9VLzcHuLrKLsozL1aBhIAxJWPuRuCif00uT9X9w7J+AmgsOry/Smofb1
uSNEF6fWadYzljrDmssjIY2O6egewfwUkSp9AzEXk7K4JcwxHQ082sARcg0T3UzY
ZO/4WWRnTUivDv/EoSOgpS0Rx20iiX9rcmlEpgnaPF5J8R8ooM1Gc0sLoZ0hUxOG
0PQsF/um2cQt00hO529D1M8ptB2t1ipUEk7SpYBZn9yHZ0hC8+k8mJ7YLXefMEge
DVTOkNCY9l7D0nkILF0DPhRLpbqZ6R0cirMN2gSKwBV76xpjhmJQg2j8bLMgsU7H
HTw8foD5rcHcQHy1U3laGWQNETi1Ny5VTHEn/KelXAwwTpK56PMa2WhGctw6fRRP
5oDfuwwO3gyCBmXR1y5s6bkx5LVh9xPBUVYiT6tifX4yyD5vnZp7J296HAM1i2fL
ZYmmnmfzDcrCOVy7qBUOjZBKU8Q++yZWI15ZDgiUgZySMTVO0PMA/rhPxIN+vm1O
zMVbHdI3rrDlhSnkTI/sGZ/tFqRA9n2r3n4UOWSdYvAn8P7hsSAscJ62BkZhLh5O
EQzAan+OjYbhqf0hTy8g7lDM/dITqnWkR9j18yHWNDGPm5pjVqghBk39psZrbBIk
UzIoffZhfuWPfqJaDWWCtG2tO6khnDJ5MHlB403Ym4QjCFsS7tX/oZPz0O7eLLU7
63b0RF0T6MmQGqpgJ0Gnoar4uCzi15+1P6FAkvTWiAgy1GTnhNHqfdUaDgKLgVW7
4IlVYEkj+UoUM5kAQO6zXAElsCLzSomqq+if5mEE7gYGoLzL1jO/n+KvZXOyxkfa
rJKFcLewsSZaCh9iYQAv6H6LmfTQjOmZPnXcw5OqF3G4JGhJ0grIFNhH6MttEdef
WU8CT24E/PUTJxXoMhubd2ygVefF1h3I0GKhfTBZHDN0YBtYvC0Ft4G2Xc31WCKH
L1qiQtXh0gbupYX/IGMsB0w/wUBQFV/V8uUUva8NHdeKr0QQd+ZhuXfdu/JVjF86
AEGHI4oT8Fd7FnqtZYOjbbIwyfMarqtdbTT8PaGExPxoGBpgJEOLFzOVIx1RM6bt
19W4I8OIsk3//mbFQbpBQGdD6qX4dorG0iGcuSGrtfEyoHBKqiwsJu4F5fVg0wd0
AAoA+35K1WbzBtKZpnnkNPZkHq0GF4on00W0KT/GU9MIaG8xvrSyWqsru9xIFqOr
YqFyeCBIiKlCVErNAJ1LxKf7E5LANK6eci9vO+PLQYiqt/eBzwETTcTyaWRpkt9I
cOg6zC38SviaaUms6nTPedP69E71eJDfx23pOwcUAeYEABswQ6drs+hNkugjRyxz
8idBm3L0LFQaWNEyXEgL9jhK387HL988igIMOf7RwGrSMEULYfiRImhNXssg/bts
4uleKEXQw4VsRs5eITlE4Xz/dJNphjqvuT+2T+7WmTGaTeW6EI1E2jd/Gdc6cYFf
uBtt4W6PGZxs0gEJXzit56DgQbgHf2HMdGPqNYVKHRaaxuX8SgY6pLqLXr1nL/Wy
4hTOCvlTU7jcV6zO7AUAB+IFMQVttOc7dH4LKBoaPBiQLyyJLWWN13YpAD1RYzTs
NPnSL8iIbYg9wI7GfS1MGOkn9goWJd8lJLfGsPR4w2wMaK4q7/VIGkfUqmpAw+4D
9PlVrXN93QjHuRPof5QOlnFU2Hj00qynGNqgfYwmNCQH8ShlkVm/QG0ExY0N2FW6
uhrJKACl7lPk0f8itJ3VQKrV/O948ZBIaDY6LuSTyABr7gvxFYex0YmcY4pbwCJn
gKIWAl/+gkf1qEtCrUVQ4Ih1FIQjQ5Ds3T7TyiFWVg0YCZb45D2NuNTND5CORQhg
xGimH1mRAXN8wnFhK8lqO+7WWn2Z6ob6ej6r4j/82sCz5nPU/r2acjNaATp3oayL
KLjP1r9eBCdSq+joqGtjJ6q8+SWF2o7/uEoGVOzPEegG+j1qePjXFT3TLFdAXd9V
lYi9SK2m/4ryB+JEDfY/EIoyze2SZYoWaQ1SUA3ej60tCuvrNybgBt0XkAcJXWSb
gC3fdKcjPqLS1vGnnqUgAdWmXjuteBCW5BQ5jyVTazAuIGeRkmWd2b4eQih7Ukaf
dw9lvqjZqs7V45GzLjrvGEQKW1vF8jaWk/g4FMTrtktZQM8F/vmP4/fy8wpE3UTl
ciCRqSgWg2nTmK1sGKGSCGJd/quDynnDNKrWIzeKDe/r+Cd9DJSlXSvEXGXHi+xj
ndGOS8qyWq8Ki7RrEerfLUBVHa8zNzsV2gO9jRdcIYqGvpGGTqwDKGnRvhJBU3K8
NAGIwDjNC9iYmffJBOikaRLe1YSFs0fOaKHOk87rRkgLCXxefGevm2xWMtFiEfo4
RA2jMekWyeLIGKFht04S8k3/u/73hF3slbjNUJGAgbRAVhZ7KlLp+F1PeTwrZ6rY
HyxJOuErlzhBzAVmtsTUBs5Yx9QmFVoWjQx72fvUch3GZtz/9JmTxT3uzs74Ttjm
PFNojEGzYe8OmTmXlTwEWzzCVJ9pLlSv1GtbTYoJmXPyJEUmYtdtC26tkdqrCTGS
EdWsrK9ALauuxmfXxTqW8u2zTBhTiwme60oof3lwEaboAVDyZFVm1dtRfEpYAeV9
AoYm0Hzs6Kop2Gyleu/5+0Zy6rEjh1r0iZo5v3ThhI2VLOPqhRudir6XX4Gybzpw
8DusWnguiUZ9yVUT+JvPrHvwNoXAJfoGLoX/zm0DmRaNJZAVlukvraQ32hR6N9DY
I56rQbJTx1rCJOj5Rt2ApMWip/lncnvIcp0kKYHcLGuxgQkB19jk1hYjIzH7KQqg
w6TWxdV4ZYIQBCVqVKxbeCLBl+//vKxnHP/mUnSMyHRSzAN6/Bmp7wWfXsqXHUvU
XBzdJDo58GhKyQy9cs+7ar+egwro+sWD+jLK8b+IPO+Vzqtd0ycngUrt+cREYzWK
fuXAX2ts1KwwAkdnfqiCLLdvq32TSF6C21iV/4UaR6yGfR9kP4QhnhVKqdcsO44G
Wh1UpAhKJv2UjR8IXEYJoRGVcp+DA/k/HFaa336ixIwFnauOR1OacAZqpnJIqJZ8
1+JKXOMlgyFMqOcZBbL57eVVnKPFy224TNsSG3cmpeyo4z59YWQCQeapXGH3Nzeh
gJupaqvjEGePbqQ2viOJYeLmcd+V+KwFW/yIx0tXJ2FheKjL2ceUKQ1XivurHMyF
a39JR3n1U7MqS+pwJ9YXarhB7MFeA5n8AKIQ2w9EYFRzJbgUcGpF4DyO/BMH4Hw+
NcwMk7rFLXfHXzNhFosdL4kVlDzhpxrY5/b/dwA8w4IXaTBjQLVER8nzTt3fm/0k
P2M/HQhFwlOwlOTypkTv+pgRnA9ek037qKtgK5f1IKe499xZf/AZXdxY9cHKFVjE
Dz7HMV0z14dTTZkoXN2IeNP7XMQEEqwwssCcM31MkiCmk/GiDdJ4sGqJSoLfel/s
9ZGSzzLZxxetLohG8rnv5d17N3lGu06sia9Vc+9aDU09Axi9kNb381TiTKKjS1LE
5f/KfDVfDRlz+fxi/pSqKFgIqkkp79pRC/SacjAzkSt+T26quW4Pjmh1ZpbdQAmc
R3H3opfTH2CNlJT0groJZV/uULA/tJZQhuHVqP1CGLGEcyA44wFs0w1ouBM3B7kt
3ku1P0gtHd39SdyaFdKeB/5SRnStnmo0VIJaPKOTAxGDcH4elknCwtpzwyQN1fH2
grB2jaK8R+914lB53s5ao5kweBnFGph9ayaeNYLfKadOVfbh3x6CqHgeZL7M5LY7
isdxS4Us7KVqYazCCM2YcbqCIsTlF0xhv2tc0G6QotsIziQm0xg09MsYKZ+ZEqv0
36bTVXzeBTZFVCvQxLseJhclwyUMMtJvG8ZZnXqwEpqvcLUgUvt6cecLwe87xIdh
QZWC8DlgfBr3NJVJg5E/6r525cfcdUDCbxKPivWUdmgLZPCMwuLPcB2de4ONt1hT
9p7uMb6Al6ADRRrwFeTTYKBEqADJTuhQh3bz/ffdZazUAhhxE7WDdgBAQdgMQAYT
efsBMwJa2C4sLERkuBN5TjtXRHYx+qwJJ8Ob8Y3fdKt/JNF6V3qHPLuEX9cxBzOF
I3oHVFmL+O3XAir6HrFiVbmCm9MlE0j0xnIMl1bKEJQIUxfQdXxDGS29jxRYVJLy
Ols+qilEBY1gl2nahzBELFL/xdrRJh/umJqdHokFkerbXVnsNvEKMll9u3NSN2mn
j1gvUkY/ULVSy2izm7EOCO+GqjHR93dPRfArSVW0LkvsOg2tmTjLB2TW7IIaE7je
A2QDZezYhAJ6mkruBRGxp9Ga2QxI9tblxqieRFkZJsYnhgjdwV8Q3TzadlWi1pqI
hvrHQZlB+/NnHkyP18jpxdutjDZkUUqKUohCXQxOSnWLGRhIWtXVmuueYKP6tsId
akTzsln8oxHRwaTPcf2tyTLy10nhMF37qVGGc7BvMhFuyNHe5eCku1zhbqz/WMDO
K5LUrUFrGmSrHjt+MDLXjdnXyyAIhRCsP/zVnMImopMqSdL5OnSsihqEbq3Avofh
2RRa522l+3virHaZjtLnUs6xWmTS09Bl7LLbrCkdaE0o3xoM4m39QB9AhLyB7pQd
jWHRzlZxIQIPB/pMN6B1Hursuf6BPZp7nWTp6bcMa62NBYm2S2OCdvNtKm8NHkjH
4q1vyBNjvDYQZWhsE78CS9JZlHeTXyReMlV9Zm2lNOY/XgbEAZOnTP17cXTgGmzu
M1DVnnLCn1z1cDpdoR63hne3f5SfMhNK47C1lvriNcBs0fOpfWEXeVTRSkNzi4Np
JulIG7O0YN+RF1lDTMlC6zquLZgVX7dy2GWz8w0lMSRWY41wfLNoHys4H7x6WODx
8x1CSPsdsuooahhWxepheRY7zINFumBfeY1OxJF6G95WqvM+BSh0qpk+yYOForYo
aEh624Sequ3E4/vkXnKBFUE4KoWrPjor16T7X6T0S+MzM4P3F3myiCD1GuhlwfR3
TKxXw9JULG4eVmmP7dJtsHU6Nc3Jk0Eef/WgG0Axhx/EnSIbBFSZc37W9wpn5Cyy
h5Kajc8WXMSOqTKvsNMhlJWxgd35HEdPSiItuJ3ro8S+MTjnwEVKUcCAyMh6OBXk
GkGWonazXH8NflEF3PFLYGCYJ7nAwgzpXaNsXhCr+/6UstVXNGUsTLwxI71DKgWr
wOaftcfJiuSxBzj9B4EWzApSVaFT+AUvTdEg1skhYufq+iccStUfV69w416L/Grv
kYcP3+rbhaJ8+Qemzj/OoDjbVESXfHh4iDGFGBO3SjuwHJLnZwAtlMKNQY3oskVm
PF7y7atydtyfPMRY+geA5s20czymAcXiAN/3g+pzWoK01Ut6nj9RXhT1/ShhtXyg
GERS2q4FWWnUkSEqrfMVg5U4YBiM7R1dWAsuguKzukPKizgx1lkhA4FsX+Sn0lE7
IvVnRN9UDYhf4eFq0KSHuzt0OasCUOZFwgDNYl9Q6PROTip9tfhulAJ3pdYU9sOE
+70CCXOWvSpdmNDarEPqXPBGXRKeJmHnZxD0OsI11+M/jaRGmqn7mUPNFy0Aw0y9
ljC3Uhy+dvfwy5r8GoKQbveWjwtmPMHWTx4x8Wl1Sy90TNp2tZN3cK+C+UnQ3qDi
whCeyco2RcndnVY6WmMPKiWoPTpQ65AecJBYOfMi1D7lXXLqOfvojTM060OLgRU2
DX2ClB2ROSdXPow0TtVQ4sT0/dcDaFh5gMn/2WRCmjlzG3wtOC5xf2WdgsdDCLnm
Y0ixsd4flTq0fkla0TAGGtqGQk94lYR9je8Zu4J8kU+xpF1f8uxAzmeuDL/PGyV2
b9t0SnsFcLbijOAV9IspcCgEJzZ1FV3DwuCjGIAE6OEU68ctZVlbt9uKCr7iWXdd
X+IevttlarSy1KUZ5nmzZBh35EWJne0xEkzZzebOjxRHSJPFDdvOU+UKrqPTvbpv
eXq6Ti+AcIRTI+GjlXhN+iXMyJSuKhXRMkl06gF5tJe+Nlarf32z+ncX/4qdWQoa
QjA9hXeKGOoxQItIJTPr0Fg4u7e99HAjrVHTVQKZI/r5V3+EdvvPteNIr0nqCoum
bKxdJfPAzebZS7rbdD14zsNOMQI7D8qt5clTy41Ea2rrXcdReSVuNMl8iltksS2A
ysoMNXGEjB80wMlIlkwwxWNAO7zCkpGnFcqkIT7cSkVoKL69NmDZHhjwQ1wp3Vwp
+vIjyGEo0+TkKvBq7AKGTlOQc+H8GZsEIbPT8odRyiiJs+YynY8Fac9oknJLi8N5
q4yj0QCEOMWmN2AV82h0gS60z1EcQwth5wH49oH/BdLBoRYS6sulld2nUV7a4qE+
8k2jtkr9qxtmXn/3G3CdOOUPidhqjS/Wjh6YC+1GpZAO9RMEToTYShNEgXYOR0jk
dp6/garKsrMdwXofXVZ4JzEFw5J2M7iYniu3qFu886jg7vbPoY4kZFwSNDGaRewz
G1VMK6p9bJuHYQUG3VeIsRS2pWT1PzlVClHt8gKezqP4Jb6dsFn3+aEJAygoMZOt
N5PSMrzCFSklCrl9c42OGQk3x6AqQKo4wZoMDOAaN7onGwLWySflq8yodCtJASHc
4+aZ0xt/K5aS8XVSSDomNGylreKGRCu026piHBap+m5g26KZOjKReZt79M5msFeE
3mk/6z9UCdwGoCdnNnBS0VZqu7rYMI7CGdXTeACQ0Ga0cOkVobWRguciKwO5M5qi
CY26xI93Olz+qEkgqjdUpetLgypk838IXb+0THKfmzZ5ky6VBQX8f22evAPo0D/L
AdXp1azpibXMvf2u4wrCeCPtv4tAmxjIfL75lFrteksyU2cIN3lLEQuUSim5KSFw
j75HmEyYQJmqux9qehmUoNq7qNZg6EHFdOGCcA7MrjNlL9qlfYLf8fxMt/g/WjCr
05qy3hU+wydleNNOlInrpedXBEUV/JUCTwrM++qflozkKYapSXG/NoiyDkcEaKkl
ZAd4SOkGoXAiVIwEIEZIIlo5h5gdIfKTVf7z4T1WBv84jbG+TFVZ9E9uuon5t5fl
2+xlUTcfKQIa/Z47JYK8389OUyXYJc1E6Q4mJ+ErMjJdPX5S8f3hMwUkc/X9roZO
HBOe3AG6vKwCqBJ73btD9KQq9ESJ84IZJYEHvtSlUVz/XhtTfQ20s3WWqyelNMtY
4uPBkSwAwNs0QJSck0Ub2YdMHSTvuib3aIKLC6T07Uoi/jnVHo/54lB6CNh2usZd
cdDEF4sItbchTRuGhaNpvj8ncevr/8I1OHyrMfI+glo7kztw1huLjMfLRacm/SC8
eKFmIGFC5N+bLT8vvBpWNwhdOBXcnGqfrzVoi6UycPpQT+eEFo89x1S2X+nQbRdl
9QPiJZyBYpHuhcljQEdCMAvekNd1r268smW0hUno/uor2qrkjm88jgW9T0yfAZB8
SIF2rr5pKFlyKXpad4fqmznb7t/BEO7mPGrSg/41T7HUMKR8w6A8NLqTU3xO2Ftv
D1mcEQ4dXgoSGzXsoTn/3m9oA6EIeWLW4rRrQh6V7g5/TkJBSM7Rn1+8WSVpm0L0
SBfSMPUYcdA+BlvKPaR1YvHeAWKBsvBeSa6XV9UqEkCdqf+ul+Cmm8QRj+0lu0r4
YfJuezdg1V4a7EAAtgfcJRoj6krc1gz+Fygzf3t6MqCRjjkXRaJk8zoOCjAXynGv
RGLG8a6UYgdnpP/boDxl1Z7aqS9esdqxVcQ2BRXNeHx7Xkl5b69vHK7N/iw9+ozz
0RsjxLXKfVmYeQy3TB3zpcNr1B1Brv1W4iqcIhletLROe72oDh2TTi7rTM1+Jboi
3iimHzD1DjzlZAjNLA75KEKDZTbD7FPmEV4sClDOutSeapqH3mlj3O7QrHs5tA2h
Djlc61E5Pk9tv5x0P5p9nWBbW83s177PezJ+aZJ4vtPuKG8uenTQ9/3wIIoau+9U
46s+aeGmMVDSyh6xA9j5ymz1E1q1p9VxhX03C9QHQfBuVxdZrQGsltyL2O4ihv5+
kfA2ANwUVxEgdZ5HLGG6jlOAHc34I7vMC8mxUiis600E/dpnKVR8VJriZrcktwOw
s+Ka4L8OtGRHRZC+KRbYUcf+bXq6Yz2D285TcLPRPmCX6/wDibkDA/60BJjzb69R
AGhMm+4hyEcAb0JJNy72nIzl/szALJhkyyv0NKnegm0In45T1mVj4PUBr11p7+zr
cPIFMGjRZ7GOsOgLWU/f8Wun+SZig00OIct4clGiueVV/WDWwS/ygf/hKc0Stgmn
7omgOij09cutdHs+1MEUZmW9/K2K23B+iGI2k8BiCizbMaYtfo2t+HW1sdns1Fla
X4S7D4XyKFpLQh7AGjWqlwoacx3vCnX7/UkN8mOrz+yoo/ai4IP8yd4nCeb7Fbmw
6XlcSzAllzctBFHgC0VsaanEZ5+/SSMUQSeY2K9APdUjOt4XTFl9e8E2zbwIklfc
MCoYfF+2+//veboQoQ6+WFr6bhtMpnDslZSvvqRnF18HxKPjdsS9Wymdx3XdyK+K
IsbvLCNfrvte68JCQx5A5rBPsdncyLAXGrkG2fnBVt4ejmJ4WNAdwpP921+N7PVQ
CT5UgLVjgOjLo1PIrTa6jRQAe8o1b0U7U0lwKu0eWhfcbaDe/Pbf09dFX3nZVI+K
sqX+5tF7YoXsQo3VqisxQl7kPCX+TBd6CXZu5zEBUViHKv5XxfpZHBXPSz9Uh8T2
CmxzZF3mRaRVR52Sr5qL4p4eIz2jYGVwjHQ+Qob6l7HIV0bPkRCeU1+211rxXxxu
91naW+lTObMyED00WEZD/sVydYZL4m0Wq+7hRI0l9zun22LwTXA/Jpb4iujqeutu
1X2UHctZlx0FxRIkUxjC19DcjATiheMjyWLjkLq/V8B+7E1QpH3TENH0/Eu5xkiU
5tIX1+/MOSCT28KuIrlmd1tLbD9yuk1M/KV8vex7FDqqYsJGEb7qXqV6iCVC4iq7
GP3H/VkR4eua99LYUGuJARAfLrVLClja4isbqIXFUlY2CH7tLgq/lHHznOxiSsrt
TG6NwLKrYS9YOd7L4fICMlLELqgowrFyfjM5HIhPt8aR/jQ5J0kRtdzW19ZUjvN+
yEwDmLwlMp8/zxl6nATJjHxv7wrXKBi/JTr9Kz+7Q7IinzFnHOXCuxINQltIS8Qy
ZtvsMopvKhm/ZfNUdfbQIYIbzUdZHU+wUbJ31A0KD8TNmI1Z+JLRRa02hdc1x8JS
zFRRfDLMNO9gOwXYRW3whn2b+UZfRBF1qp9wlEWboEGkLijX3tNgmUgUbqGUFouc
q4yOwbalvWdB2+lvkuqqm07/pe/k7Pk4QqV4gaOneeTDJ+bhYIjHQqPaEUl56+HG
/C/4crJ+YLaQCtCAMfPYmrXYpZ/NsPoSTVsvJMfdD6VhhO075nlBw6Dd6CVa2KFY
POoj0mKaCUcHaYcn720T0T6bhx3n3UUt9l2AgbYNpcetraKQ6pObtq3b9rm823nL
KpofxT6r/S6PlbmJjTrhq69NkUtX5XX6djEsKSAA2G5zdT2ToowWsrb5XBB3TqhH
oqlIuU2mZ9pLZtwprYcDQ6HgnG51bE4VeNIO4igyg9B2rMl8jq7G8XhECTF8wPnS
DttXchMaQe37CUlVV79MWy/uZneHli/Sa+9v1WBYYqIuRKVnq/GCEoZaPtbCVGlB
7/OZGLHFd759Qtd7RHkHgHDDXHo8J/WSx0Zwlu+Yyiwyl4LdAKW+AOTsPAgT2thu
sUuY5+K0QJ0cU5NCL4jazhBH2joWVgVXwNX4DBwzKhAOzW+e6jPAWv6WlcVUOHej
f68cUrR/lr3mhf9JB1L7LJBsnBwlU2e9dvp5XnDZ5lSdmFgi0wZDqbZ0UI31Qs3l
kMcOe2TBAXJXl20n6KjzlsAaarOG5DrE16NFY07yJVeaaJgKSCp+RGIggBwUOyMK
kEfyVl6iqQZveTSuwEYsIKrXns0LK0O8FPmY/dgLKq1r4BMguKcFrQ47VMozaUle
rIIL55IDej5FTEoS49+ej2rI6J77SOBAW0CVTFmd6ABuEVdy5Wv+jpMLRNxvYTxO
HgMXA0zri26q17Oakt5iAsvCQHW5A4XibxkhOrQzeApl/vSg91byopvgop7QR02D
/p9ga9UDKdrZHT9U662ddaEX+ED1Cp0RtYKhI37iNDa20QpuSEAj5BUbcLejkLIy
K1f+hUFtuxnSF4Hi1t5NOQN7vHgVimb6GiXvhgmr7PFIewrlzOvQN35UW/wKvotI
PXIqhIo/QoR23NauYroXeAnhxyAWQGPlDqXTM9G8Xil9HcKfvOunSn5NvN/8dDeJ
T/1IkCjjxdmQZj/PpavpZLOOYhikU2ObcyJJGbyK4+inB4ckM45PcX7TJ/C46y4d
wIXixCTWXWRTA25WlgaIi14S9grETqF8fuvcdYqYo8hCxucx21A/jKnVYTTMjo2y
p46L6wyZOIjC1CsFusyzvDrtmDIQBA4jFE9L8sEsivjpimrvTaBem+0SiQqIvfGH
7dx5A6PpGGFePfrMypvV1s1Tbs3FgEbPYmexq/bqxuZ1L95qrF40bM08N21eUhWo
DIk0vxnOhxpuic1LVNy1fD3Ami7PASFKR+3Hf25XjTtwEqpFRfist9O5ODi0KO58
rXArX3j9kTi5xv4moiwgbmznl3ZnxCDDE5TVSBJr8+MJ80IO/G7R68snmhdDpgvq
pcXc4+U4lb3yNc8fGPqG0AZN3lpP9fHPT0c9xwJtHKZNi4SPj+YEJ63AzeLsQpa8
Z916eeRN32jrvDWPqF0K+nR/k5R5uo1qBGXEuDhMcYmhQom7z1WqQyYfQ4lkP22v
pqjV1MBkpIjGE9BdDkYQN6K04u+7ZcqTd5GVU3VlU8AkdRezUJaonAECz+PSpjiA
7uL9yQrkd4amHOJ8lZKuPIgrpkQSQTBx6v5rFRi1jPvY8y3sWkPWCWgR0iKQFGmg
gQ7njWRGiaT+hG+6I/2ZVHGsFN0VuOmcpPh48TCDqZPQ0WAd3+uDCI+u9QMen3mG
617fbZH4H7MW2dgOz+7C8sZNRW40AhCW4TCnvvVhDXTF0k7kOFA3RK9vA6qy4YxG
RcSOs2BoBC1DW0hIXseuqRuIhYc7btJeDNPOSnA0X4WNHOWiYX4Yyxum6NqpBF7D
xARGtPBfHt+zCo9myyk7kqHFMQzaDcFvtmbHqsE0EauSSA1RtSV6CIJlVVEEU8MZ
OR0jjzRaVejmtaZgDi7SvFuFHda7xsjNIWMXunvgr0aeYnAvIstZfzSL1W3Wf4Sl
5aXOg1w6yJeFwn1bVjn4PkqKbicG8Mq3ZxU+ASPuFtiCEpi8EMl/0zD7u6WZE7ei
fEXFB7Bhc4Iq8hEf1CA+FWTOemFeTdZtjdFwggX0/gCKRv+WO3E7yxOvH5CwQPH3
P572JQKxMhuh5oMQZgmPQpYAIA3BoRy9TxAWa7H6MLq5Dq5Y7EXWlgexm8fbnQPm
H89Ph+riKZK1pJck3Cj8AC2y/RnhkPaQvKDQ0kLZfoyq12LMT7nQ65LsZlY43bPq
EhpJI41Oev72sDjYFRK/IroxcfVkxtVhgk2eWsWnc9/N7V1WJPqB69m76muMCiMy
y19E+o7nHdFfcWA9mWOO9blVJ5g79EaT3AhPdwobtK3ZkEBhOdYPZjV1N+tBM4JW
R/Tdnp0pFjc15KVCXpPjhpoBya76mUQ60P9S1+A+ZilufNov7QFpTPR2LEEC+vmL
xiFAjX+t58ZL/ts+bRspWzQcPtFHLTGMJQsNwbyUr6A2Hc0UlaHhlGLgnW8uQW8U
QD/yFHQW3jBHTTAv54APFNwiHtMpZG3UzahCh9kHQTODCK4BHt9xqAhLz3S1pCMR
vjEIwVfI4EqUX8CMgzzb5Y5rmJmPJAYISO78uHHi6yh+YRf7O+cAHhCMwxiWWGQ2
UURd8/yNPwCyZdVuicHwgYsTFKG8BUJKQFvUXpu6RxEXt5ity6j5WY3qWw4jbsd0
nJOaYeYvDvTMFJQqCIu6L9wAVUuJc0o1hwP9araVOFkT8o10GQv1vu1mKPfSE3Qo
VX89tNt1XzfuC0y8+6BNeNI8AzARnr71FpDqo1LIliBz5EtmGWE1bM4JbrM4xfkC
UAImfhYBgDpzhL5FLA303H0m4yzW1Ee380jqU/5wfvd+SrLtqu9EXq9BYf3qXQVo
FR4YlIJuNspKoZVfU/SopJUhZIQGsbRVKW7k79qYyy/vc6yY5iYo6sd/80IP2a8M
7RKa3Z59L/ACNdJXpaRV5DCZyQkfag8h+hYDIdIvWHOU/MzkyRB1OCqI+xABBmAJ
7wkITOhNxiJ+ujoH0RBPNkgmCvbP9qNDeb60h+uEj0DYQ2JjRA7PonOKWEEWFnKs
56xFCX/MPcFV0eQWsoopED33pzGqeEqNjE+AiOD0cJDgoioTIT1EhCrS66g/tgDw
i87w37rZM9xEyD2wQSnvyyQd/ZWtQUa/PE8kE6PiKrlVSowLlhj9dcRneTicum6R
XEoJwzl+1o8L50AWUIaqSnirGUo+Sf363KHOmEBqNnzzykBU9mAuxDpTl3cDlIMP
h6b1M5SpGyhfcrmkZ1E4nbGPlfKu39fuTfcFVSEJDOYBtER3fv0BiJM+ooPoquhI
yQ6gPlo3k8oQTNbUgdOSj/M/4GZe9V40sW95eoRc2rYnxYEg7GfxtVJmtX175FaV
PY+E/p2yq/L2kk4HVjbmh5c8hIyaQ1j78ZGmMQCqNyl8SLgQecoqUti2TORmRcnC
y4yxI559NLGzbw+OU0BlFJ38VVS/KtI6IRaGRKna9tcTmMesETLRd6KbGJAKUXO8
Lug8jfBNIMWAdBPze2bjStRlpjrWznFCMeH07lp82NHDKdftWksszN+pr+pJJj63
wbRHpF+TCgxgNmKWgSGldiuHRBBRzW8UBXh1vAAPBLqnIsK6FgNOjeOmSiD40iOK
sN/ePfgjIShNMC78R9QII2gkgUEgkcU7CtnQnhIm0DP5xMLURGx2FfkLCnLO+fCM
wkR89kyt9iIdlOeJgnSAb1TCGwheGUOdfu4ZnHCKoSGgdPqXlnkq0MuwrcSAU7nY
QEYDXERuH1d8bdabu5OYnzw0Lg6igaX4slgtoOCp0KfFi6l7KKyDM+b5efvbWc5S
VtkfYRXP2l91OpaEHSqm1LRj06yHUqD4d8lqj2Rp7Q9x2mY/kI01RXyaOVdCGdsc
Jm+JFJITfKohmab64CxrivlWo31OgjWYHT4wKka6OL3h7nIM6RuaHwrCAYfSy0rO
T8DnhXouAnnquPqgCnfiGUT0Mf/GwiLCsA4rTMC1DftRSFr27DQwrUmCLBb3giL+
AzZ9kS3Jdei/jPoQVgjc+ZVRR0PhbxjZ27q1RmgT+3IXXSh3aFKxgYuIwRDTdW60
/nFLpFziIAVzp77/6e26qyqASvUrKzxo58XzRorDCMwYyw3oI107TOu7F5TJdMm7
M5HwcKQ7TrCXxv6lHQd+d7z1Mtya2oe2aYfZDjkGbt5q4pCIVhSOL/fgrKFIYiR2
3412847DnukOl8vpDroo8DMRvVujrT/4hfzgkSjNp0/sM/gRmcpzS+isXNlrIHnM
qhPFMyUMY/gINcbhjRcacdf3x3tEbp+JH2fhGy3KFO62IqYkeSGPOidZS7vDhLW3
ExkvXP6hlOGdK3pLaE5OwxcWztMch/QGDKfN9rMWV88WhHohCTFCUR7WMflPGc9F
hBjxgsJ3WWFcgu/7S/5pFAI1e2xg3ap9H6l7SHP88ZAUAognkyzmymub85AiUpDx
1vm7sNfQBFYnWlpWBVwQjAuIwr18Q5MJWdEKztBL01j29jD/rhI8porA3PuLc9pu
Y/AQzhInFx+Zk/jcUsp9qg5f6WzhMFJMldVquRxYZs6w2yINndoK9GmTeWmlQszL
K5PvtkdKsy3z7xmWJM5AWYxfsal57IPqq/tquPn8ydoQUVHPfl9eFFiCJAz9H1E5
Z/HgoVPdrd2MNxqO6SOiSkPRePjJEOLwCidA1lgXxZXi2pB9qFyiMZTkkZtlt4DF
QubLltc+Pm+fF9a0NrLLSyNF5nFzAqYcCV1P15o8w/Rf/Bvr3YeXLUiyJSoDcbS/
z9d/p5PTGhfeZDjbgjkzrh1NQtG4qXMf4krzSCiXx3NPeYUfqCAHEfmhkl9zMmq/
xP4Gz0gFe+PsfDLFZpvqO48DvgoYW8zQi96fJpKz+NHj+vuyFLFRHVov4211aBw5
FZLs9ga8opPa2FoQwWfBKtuKep+2vGSf9Ynf68CO+Gm/5SLoMcRzSLjCV5k1K4Xt
er1/s0QExfsSS7bFeudOWMOKy5r9o8OS32y9rWf+djCQJUryApgiXfaiOMYI5z/B
FLsOItg2QSiHdb0q/iHFTFYXMm6KJmlwJLUjAkUtd2UC2lIJquen1iZnhLNqHGDh
ExRdqa7R4bj//GMoTfGHISweceUNf/OitLrEiqxPFBghzVbBQ1q8xJC7TbKxO2Dr
N6SGmV2/up1EvrqNudPbRoQ+FASG8rHBT2kQj4124uK6/5riYR2F15k6bw4L3BCY
rF7IXqLt+YglxLgvKKFIwPjocNL0FGtS+BwaQ7C1WVkruoaZD+U83V6xwiAGs9lX
MOrUP02paWXOB6HYWX3Fn2MnqOBOWQVPUq6X4rJAHhls1WWtTLsCFPsfTjWhmx9p
OmQLB1H+Ee4UWp3gxtOLy+gpAttxn4Cyem9CXx+CHqfszRNN3xdCw40B0GLMG7/3
FgmqWBkoGyPpT1Ln7tiFVYJ4M22wdB4L3eYN4gjedc0fUIHTFQAhGX5MLFDTAOdz
MqSBBgfw59euh59aI4S+/hag+XArp31HrX2c6E2EPHCynP4bXwQrcDpOgyOx9bij
KEGbl5eDEjgF5uMf6mgQ4laZf1oBaeOFF18J2jayvxIIwYUI7a1fllC0KuHzVoEa
Je+6s7vQH3/BuxvRrEd52sBDhXvpZonr7T1jcNbPvWR6XvwmCZbos6q8MvRXrKHw
PthXyPKagUE6YUIYfgYmtuY4tvF7FjMmkCYrWjTxDq1fQid1lyuiOh/yyirbp2Iv
Z0L/ZXYtoqc5z2Hsz/kJK+24n3w+y4e6qrr7u63IG8CdVOz0pVXKCZcY2dyTucT8
oCExlZCo0W/5YClBSMC1MFLXQdVMzrOHzteURtxyRBHPF3lyiK6d3HGruvTptUeE
Rspw37gBUVz8OSwGLstCW9BREgGXleE+xMdzJhUciSeSX9BGpPzbV+rrUqTd9rXo
0oix15cfUN2YxlCinfFtkg0iB/A18vC5cQcZN9sJtVxfbNl9jeOll2wxsIieaP+Q
sbLpLMLVZMc204oPty3fKmWiWT29OyuVetQMw5XIL/M96VThQyt0lYtCR4Bb4lqs
gwOQb1xrYAh3viVynzgWaKLyQ532S46PwyKW8+nolrmVsQB7zggiqTMs0zYAMAxs
DXu2A5u+k01mmG1JEwLjHJpjOM8vWSQ92Y+EyE4RdULaLZB8Xg2XUTxxncQfsJ0x
k77gjQRdFc38ZAdER4aWGk2pVg4+sG2f+oy5XosaSv165t42bS3FAJvubqHaMR/P
mvaMTuWjnBUldNCt96eANfrIGzECXUtql3pTBvgjkGuK/Y9bsP/T5xlcOmc2rY35
Q/s498uWL4sucS0FR0ZYNGlmwD3rpwbHNd0NnieNwxyFJF4/9mSib8FXvJyVDusa
1ZDPdZOV9X1vhSGE93Tp2jHaPHSA3cafsAEGLhVzlkeKbPzXUwFV83TSjq/xM9C2
4FlJfR5L75ZbZAIlJXWrm6UzXqSMcnLGHntEcfQDKiPe4mTC3cwIi3dqhz0zfwfB
muBZJ+AjV0Dty1yi0Hox5OfjwlTkpUwYxCykfnjzMo01/iJhKlzoOVSxsFDnG7z9
sqj066PLXKwzeWnAlXB6Fx6QI/+7heNGLkoSwKseSHYQMhivTVZKoPZMqSw0DvkF
DAEblAAOmXn2RNSeYVZqCNE6T5y1You9oNJ6uYbv/Kc+9jnui7xxl7Dwc0nmTTBH
mSTrnGLeg5ms6vCuTtHgk1OG+VUKXXIrz6lfNfPBaFh4ac1Y+egqRtzocknW//EC
RtT3bn8ZRyvTthHt+Xa72iM9MCyRHx4tfc6Vequ2J2xR8fPDU2q/QbqGQ3tqofIK
buaskWSUF4iH6lUqPmQSzwwg85A3ggPQJq7XSRf5tSlc5IhrkuxBk340kGnA231J
HuPs2qhXrF9kxdUFXclwAcaRM3btWghQJoFTha/3jAgxbDc46+eAz2vJNTAlJ2FN
gHag9nEyMW42TwKNuxVGeclCKs8iY5pxbhDvtldJb3V+3Ero0NJrVi67wKFhE/n9
/uIiVfmAbCbxeIH4P4zTQz29mUcTuFMMLpL9+xBOzQ3CLKhWzG3eaNhrGMx7Ot08
6mb686bzCJAeKjIeaYSqukTPSEc1P/IgOFQOEEZbZXv9pDccU4aFbSUkBpHV/o6F
qFOKbATuHeJpsuWjF8I5Hn1h/+6QmjaYsCtMk4ChohCdAZXtSUO3kHRS2R5nvkOq
phBBDhXUmNdrvaR4Gf9lK8FRyrQSqSzIS2lNE0JlFJatnCkb+ARZ4+BGJtlDX0p3
2aCAWdFWpqC2VcewXe9iJp0hMXNGmxKUS1izo6HwEo957/cloyrY/YtPdERDJhxA
QmfDga85U5gCY0RmsFihrgrB/ylX72YE5uPsZ05FTmwT9UZluPiNbRHGNy/7N/gS
VyNhCKxVpqKUQCUPQ3WTt4B/HPGBMmw5kMcBhLRMsYfCnavi17gKP1oFWzedxc7/
tNxgw9JOpqAX+8PGWgq/knHZuQFxcaG/CjEYLrlH9/bOquo9ZQIGb4BYlVy9Rwfa
dcUl1KAFOMt4E+lgd1c17DV4iHwiFaDdXydhsZCe9ILsAhZ8tvvlHwb32T/4bs9O
3om/iUCPjghB1sUeO1sWG5n4z69lflbgwLJ+WnPckirtYpjxYskEaiEWvhFmSxW/
8kwW7YP+4rIhRSVPbdj6d8E9yKAKDE6LE/sCwjEuAk/vbDI7+wa6lU1XzA2GT4yo
QTLZZ4fxitA7XQEo/HP0VZERnISmYYGZrbvKgFa/S8UQIEidOsuoMgr4oUmFykFe
qTdqmgbDBTQGwj7MemnpbqDxO1TdnbfJMaRKT8h3HzDtfQFaW41VLydt12XTkY6n
WMhsgNdoONJhz4f6SazbGGG8HSv4qxbcpQh8HZ1a6wZjs9CTAasyvJ3igq3cFetg
NoH0MjJ3rMavBUpeb0AHSK3z8v4k5zM1s/BstsaLLuYkokYyq7bMZMObTHWxX5zN
wcHD8DQoTtZHV3vg/T8TEqbWdyVJnI0rN7G0asXk9IFpUIjfiyDZoGxMf4Gu2RCV
Yasq4Aecds0WB6vnyhH6XwTspoGKA6VuSKkWAydzQrX3xADsXAOLQNqzdTITnCUU
+SQnj5yIizfpZsza/2ke86W3F0asTTXHXbTNoGGdLFgOwlo8cRYoUpFruztyT2VP
wGZjDv9OP7xV84kAXjWn4tsTp8de0lqe/xv3j3khtzaKJ0YV7hpPGOoAbR5GAJDA
cIhBEnFKqhEj8l9777r0RjlZPJRYtkhoKyoQf+foaVJh5UpBkCEbOmGGKwcSfiUu
kc0OJGGS+TKpN0wUNZ9Koe+zAoSeCdYxdPkIa1yo1xAIM+jbfF3cCNt/3Fc3PgqX
qLUc10TDcAGQKv+6RMbYfDV7c5I0zeDVMCyCoRnQ/miHbR4k17heW+hi+wk+rRly
6VNE2JoTecx66k4qJsDjYt+Pt24lLETjsJNcF5tGwv8jYxi/ZO6ckwnwAxEwts+x
fM3GRPPNJJOZGJhpMw9XPvsT38XsJGIC6X2dVPrsvKqnudOcfeNyLyKImL6EubAR
/IdmKfaxVqOuMQbfEEdr11ohOuIwBKYKEwKX/+aphDTLXFCWriESVsXHzjKKSUjm
X9faEf62E7WpHbVvxfinY/K5XqJjtnYj+jq/09XGSVZ1dyUfE8JMRg3sig4etZAm
q8YCJf3ZiSqWIwEu038M+bHi7BJiWVZNNfLM5u7r8u1gp+udY1pGDANsoOfjo6jk
PUpXlSyAO6ZPlXMwsClEkDkIvaWwor73RUeGhlECVK3OcYgyAX394tMS/hUy+Qur
dYiLDgQT1ZD0CxrdR80GKe/+UgRZc67VhVdxxVbbnz3Mz6BCVnvpylzm1TcuCmB0
FuI63IV2tveiIDJm8/EaapkmyDeDgq7L4jvhbEh2+kU0cKnbqb9xRAyhi819sVti
qKFfA+vRgx66aL2PMHIFIuW3O+Tan4syZlZmjKKY8o5XLn6WL3Ejfxjxf2g5U5Dk
eAHJbIXnl/PqRymC5zP0f4XYsG+1VtKXOeBx90nqOnBPa73esqjmLyvTA/7LkJ/s
mTwW672m18AUHpUFOe9jCzR21+TQCkgFVFZ+FZBFaIEzAqUeOwMSliFLIXVX8E0M
XngRPBMoC6Nm4CYDNL0YrJa6MTFY8sN32l09Q9/JdeR/RpoJrdcZY/0kPCqY/s9R
QM7izVdPTTj6oylGU9E1wXdpYlsgF3kMTnfvngXCEEZF+lXWwWh29IqXf/FJKxB6
QDpTTaNzjM0z8k23hefPDFzuUmC/joKwd7tIm14LBl00KvJd8l3xcTECxAZU3bZi
d//jRXrxSA1b0zOhKwF5ntNfTM5SvmuJ8aiv06Md2pstDVyYL/AvLmXklTsQEG2N
4N/ezg+EQ5r6u+t8zEPU8iDYI6M5r8qnSAuBVnCkRBnInyxzqvThqj9vnI1bIoQs
dqunAEGrq++PmDpDMgSAPVYPTvBnr+06EnKseitTv5hdJAtP4In15NyoSToHX5NI
I/tLOZTYlPDY85ymK9x/tLLMBzTD6vHHvjGGyTLOyQDbnlBm4/PxDddGPnug5BJT
I0pepLiZ8gKaZCMOYpLv2tI+3nyWdcBt0zBB0cH//xjaz4Q+EaQsFVbbAKl7WDYH
xRSuhiRpFrWQ5uJafa0bT26pakVq2bAARaGrKuyby0BfSjM+hS+qcS48tb0NVcxJ
I0rGfxc5UHXc6uuQ/1PaKIfqdt9wnA61j9ByfrI93vXhTrzFwfn1lmGdlElLzqaQ
xuPnWo4eZA8REd1w7j2C8ZCqo0zpJ3yRAuTWM4Je0VBTLPa1mjhGN18AcgAm9O6/
IrLLA7WUK3N2EhDldWAC0VRq+gp0R/wdtHMAFcKK0ko1djTZWx7fxE4ZwLLtj/Vy
SkG/Ul4pWPSuZnDLTv9cB4SRgQzasDpD9/nxqmoCkzPd/ETxC1AE7ZHOf+KhayHx
bNr2lg4mUdZMYmSlhx6ZcpfJHvjTHyRkpPcxSETe/acJym57uffhUnbRsuoIDjCj
l7aFIxGs882ibfdUDV4kOqAlRg9PFSHsR5D1/LPTDM4eLMcKXJwQ/SaRt7t2WTdp
X5UeTGcb0eSMxnN5Z9hGt9NQdoIft3WmoO7TdbE0uV+Mr1CogcrFFIlDEv4S5HNF
AtpxbJm7fEcxam0A6oI368zldd/AdPWyMKgOaNuPY6G+9Kb1b1XJ0a/VElS+mz3S
0QeMZGtvLGaGUL7rHx60woQcOpqPJ48X3Gpr10OOh8QHiGRVUIlWy/Jcu5dY+X9n
XMR/SgzKd95VwIs0yYJcnm9ZgrjWfE48hsrLrhjkL/LNDDWXxEo+9vKrCpCX3fMT
/c8yviZTwaWIUPlyHFaPMuPoe/UuWuh6o7P1qpDTIAEr9DCXO9yjNUkEHDhV23Lc
G8JA4N3uhtfoT+WNZAhjzaHTzTjo/B9F8ywyH4yJhL+imcpfEbbEy1qcO23aHcgT
+QMS01WMb+e+83wcJ6Obt+5PYHIiiwew5/PBVCP+y5WPU0dheOELpmY+0FHzO81M
CFO6ut3bkxn5d+Zz0vtwWwteACOyopXa3eQzbjuK2ShpPoeOS4S035SDMgwU9PTp
nvHL+mIqlgIrA7wma5aZv282MTfWmBmrn6Rv1ypE/I4T2BOcbqmg5DSMc3PjQvZK
/9YTFjQAHA9IlQz4L4cTth1H05xTTNuW4fSS7O/W01p20Uc0eXGbn1wLdlGqT02z
FcNP33cR7hhFOohGnyt0QN5Ws1TJ63s0coHx22Tb8EQ5j6kRZAMZli3eBfh0fIB8
T9pm1+Ou3m6a+4DzNab+T2NZe1WOUGc3FdU1W+zb8li7CFZI64B+xTCJrInWg3Fs
uo4WWlc9hfQQFiY002RSeIZuuufaDRiEn9XtBt13IDP2JOLgF/m79evsyrYAw47d
/kFTT/zoq+OI2kzgnLaeHEC3t92Ke7FJnGgpsVE1z30/q+xvd4FqY2BCXoB+LoWz
4tqYvugecuwrdttKBk6jXxm4wcpeF9bwpMfrLMBEbyLIwmbhrfsMn4CfUVlEbzz2
6YtlL5q+OfEKbvg/TvtbZvaxXvcYmrPFfIbgPQgtWJPuuNAA9zifpY6DhXt35pSj
vm2Uj51Zik39ZOMDVTp1mCS56f/DUlIa7xiiNYB8pD8HBrb96b2JaNc3+KIvxUem
JPNKmojeFmgQTiejL93i/Jh8rx1SehzKlTW0NAmr6Wb2sZjoqPsY25W/SB5mszij
EjOsx/FmMYUPI6R5zmF3hPWtL8LJ9O7LIw2h8nZiWADFuaBsfSOghPKsGsK/6Uh4
UmTlSHIAtwjpaETsT41QT6kaJMlBnXcGe1PLcW1Xg7HpZrwNGAInCjwmPDTc3slr
CkW0ymIg3NnZHk8neaxYeh4Z+KWslG+L2hUtySTKW2uJLJuuA3p3Vav6rCuhk+dK
gHFb7iIt8X4Cf6B6M1eti36z1HqIIoeogv7rvudZTQ7LLiOJOVGyJZbZdICt2dBd
qngYTnL9TBmI86VvNo7XAXxLPAZygdphAu0DRX1HsYNlpkVrLXRLIhiZDtXAQi0E
m+PfF24EmWQmrZvSFnZXEUTQvXOF7OWc99F1CByYvY72lVTC08tPbg/0f/hLsQ3p
pTxXq2eeaYo8b0PDqTeWK/jHawMwTB29y8fS5QRfzzT+h06a9X3GBXDbg9OQdXVq
NleCrmUKrhAAWMVbSuiYiZ+0tiNxCeXTToiS2GgaUzDJCJMnKyCssArX/mJZE33o
VmYmfNmuhkA+TDF/BnwbpHIINt6SAdRgeArOkng4YLyLJuoJxb0PTlbKmoPpKsDd
o6lA/etF+DrB/mvOElBQlO4/f7ysy/bD90YL7MLrbDbqJAjiz0PEod4OOvNtrC6R
uCWOrHgZ3IaxNc0bxVnY6kBjewm9Cz/QR9YSy55te1Zq4BYd+OPo0QzuzwsFQS2i
WTEUhuRxPEtdKpAde2wwhpfDgooH9DVjRFs/6MKkkY+bOzaI7LCMivn/a2yr4R5p
IHLUDelYdHpll5UkhFgP4nHmVhgN3TZGp1EKDpMV4LiJ98HligrfDnee1XTewUkn
33bkLPZf7tx9dGTSh2segV+DNqRdYLA7Xlcfvzeo3qTcd5L2cyC4GACPAsxT3Jtq
Sc8yjMCspkxVhf0OKQXdMxHCU86ld+yWbn8qARtJ9me7mfszZmJtO7Niotgh0kOR
MjVQ4eeVclLlpWV1bGJlFSnWooY/7BJa01OUp2G5hSMbbSv5g6Djb9oTaAzol3BX
aFM5ZnnMjviT1H88ReFAtCFIzDKA+ENOpV1sMKIoNfg93QvkVA8tPSTDF5Aq7AnU
Sob17cFHejYkQ4H/fdMj3ugY9E1Md3A/6V/LEZcpH7EeDnib7MYUJCngL1CfmNbU
RdPXypcfEsoFBQ5gSU5PaEU/nCsd0mJy+l49sxrHWyx/gkUQTmQ4v5YSfZMQhoNo
oXuqGStLNVNiEWf+uny3U9RxJZ1db5aLZyojrztHRMU9nI+jb2Ee/2l9J++Yfw7T
PT7sxBUJeLY77HjS6iqkuXkXXU8RXyOQFbk3XDLvQHGbNABWa6/HSf6du5cn5/3z
0pXTL+3JE8TNmQRATPaF9AT6fqX+LYBx35GsS8jXB14ZM0TZkRt4NfKNdqbv9rrK
Gmh9tD0Ks89/DLn7tHh71nI7C1ABYL0H2oeDglABXRLvOd2MlH2QerS5IVLi4Nnu
q+TkkisqsTk5ZpNEHL8EmCm9xY4ioSrUGlp/cm8QaqlSgsgt4WalvZ0DL4id6B7O
4fKPH7XZ3vSuHscEgM4e5vVtNQN2TnhDazmYSpdxD+oB7lnnS1sEbcsiNNvoDNbZ
MxWrzeHImuuhnl3HHAjEnTMPNu/89QVNWgZ1/qt6QSK6sje4pBClb19NTO+cwnAL
FIbICA6cnWKB6APWpcsms2aiUC7wFiS9SNrSGCHA2KsmhmrOUnFRb6L+2bD5jRsS
UYGAZ6l9bSBIqvulBFN7SpXFtFm1TIBnTij+ztVbUDAvXilo7V+f4xRMw5AD/Jiq
4TrT85livILGVXmXZycJevcnBLdoWyCXW302aL9SsefPiUaxsPiT/5L6OFbz+b1i
0JBjRSAifkb7h5YLdofQwOFjjho2ZHNgN3V/yKxXz7i3GNLB1bW+xqXwAI0/h4KB
blA9PByivFkfjD/YhExcawveWHo9amAVbqMgICpdkRV5s7jFMle0NBKdc32SvGnj
R6pscxstnT/zqYxW2ircwdACqU2I24Xj3LFEnExak7xqOfw7nc7kTuW9xejtPLOf
Rj+4/NZa+U/eKdDsWj6qvuQAyJ8aU0rHNXbfTDhyB6CN19ukBvxs088PVgjqvS4c
XqpXbajM9PSEHOf/bBpaOfCmwHaVCnWfdTCDzgGPh7pG7s9j04CjZrSmGqiExzln
CoukK+CDlX1dD5zdbd3onbFw6W35WCODk1pZdtynwZ4MeuqtTJ5SNE+Z8RGrVoCY
IVMpKTzX6InFd6gOuzggbFN3G7hGHFEoRrI+2G0ItdsYpxF+xO/E9zOWq0T1zYxe
/78I9XaTyEzqxAgMHlIzZ8bBlgFEXjDOuBKEPTtwvPmoyPR5cX4wgHMWbsh4FLtw
HYtoxONKj+9apIDqb2yXnETN2frVRPZOr4oO/jmZx9K3yWq5PFddAQPbB5mgfZ2f
WTUbDInTHvmGn7tvpwz7UbQOe0Gd/8FZcaMe6dKiGgxL4LTIijmbxEcomIEIoG0M
8Ql7phd89ofXe9ytzJhRYGpWUjd5Ajwj2g54+E5Xn2qVkb25Bk/abnyVO4Q2bgGd
QxuzHZ1xPMhsnUsvz3gIqViKrWVs3Ttxe2qOei6fBzIEXDskF649EC9zbGImgkrE
M0Swc0SXiLke58pPjy1cRl14NWrNhCvTwofrWbyht5f3lry0Qf17malqAr1DY0Io
6GsGPrB7oAjO7+gP46ag1Pg9KGaa6uMjc5Vj7rdR90PloCblOGnNRbExy5OmDvVo
dk31qnGTXbG5HzxL31IioQ7J8o/drJJ4aamb6Pgfx6bbwUJ0XV5O5H4nJWr5NnUO
DO/Plx1RdbJprvMyHCtyV1DcucC2K3FKAl6orafBnI7ElxxXwP342tU0B6+F54cS
ueYQhW5qN9LGaw8N3fULOqHIbMR2kv59Ke46OaT2vf/aZZlqZD0ifiU3zIIDLoQL
WnNQoxxmtvAI+CsFgx6dotnfRkLYfiDob2zeIlYOefKOMctZel1hwSIhawt0v5C/
Qe7xDJUpx5AwgLmZNW+scIazo0cD6q+DyPnmQvvvRYMXhTYXdd44GhPGldWr6FHq
HSOhfWuY9UY2mcnbyZyP7TthCdo0DqCpIULcaPe4q/XJBux5PoZRFE86GvFx0wIG
WWn36KzPLeKmF3IHeXX4Rqm2IKoeVKc7RtA673QnVTX2XOs7xcfQhTQeeiY5cMFQ
hFV2PB8lAvUOSwo3pqdBeO4oJ0Wk+9heDHR7xnOx4kEPBqSIPicJTMVOOrRn7zGB
vaVHU+CcfuJ9OCVM/KRaUgXL1lr5Atap83AazajUtHYqN3JX7BVbPQ34Dz01Mx9t
A7BQk+rgyN0r4XElbM8pfkkl4/D7Fbyp56bxYTabDLcyv73OEQuKr6d+0qVaY73m
opGcU41bEn9i7mMgxltCzo5fqpRkVRWoIi6xHBqmUvk3SmF10yxhcMYgFVvif9ew
HUVjG9BzMKTkr9B9O4QWIFECSDhgPzTOG0qT2bbm8ePhnVTDXsIbw9TbLH4gOtPY
HmMdcY8JlqmW5mZ3LgJWAjufQmyDhc/+69RoIekUB5JtmKZi6d34OR3eFKyiCCTz
YsW6DgibWb6pxef+moO21bYeSFVBumeS9uOly41hn+LFZxWQf+B5eaFzhQ/C3eqs
4WDRQBezLdDDPS2Ieuy46PIvbKQ7ewF5RGw6BNXtF4dG+Gdol343cP0X9bN16kU9
6Gub6ZWghbRzVuFOzqvjyJKn4FvUuTdYsZTqdnX/Y7kpS+LcV+/yH3q6SM5f6oD6
Hm0E73ovQmO3Z7aFwP5NHS4aYFTHN7gADAY9D1F7llOFvnjo5QZMm2UUbk9PnrUf
+t/B75cNQgB3dVkbB44h/Mb6+lJP0AkAsA1Sakuc+EFMUJqhjvkMITrVmde6A0IN
O7fTf9gSLRB02fZl8HkRaCD70iGn8nzn74tcSyapyodOpVQmsQvilctCmjQaQ2cR
qQZqkCEEQSMbHx0RkCG53fks+BBBijoAOvBBTfHPGx7ZenPkPqtmrsjU8fGSPxvM
dlDCv0jN+JqnQ0M37JAu5V2I06O86Z5zMlHtY0KrxFJCMYEhiqYH9ZqL74u4fgpX
kh18dVvxYj80dmRB6PNe6yn/QZAVxk75/dV/HVkkEacuptZUvgyTT4lUGVYQWGjf
R7Qq1//tYBMxgqWcKihhTuxI0FwtUWeMEx0d6Jx2WtodweyLHJjpZxrWWNM27Ah8
WGX2/KrDQuYSiLf/+lRqUttAFrWW/AkW3DatSB+7sONQKkrEUJmR7uBR6RAq1q5A
Un+3Ixi2wZG0DIWYcvAg5kAtSDARrhSeSAfwBuFNs654NJOkbDn3bHvI/u7oJJUJ
rwabyD2MtcDlBr2WNwlnXSnIOAfAz6qiGsjX5g0n0z/kQHFrnR+BPRcwnciSbjWn
QPrO913MkQ5zm9jS9z+LYGDeJpHInnNjnzN2uCkXBoJejc/TSxaDq7O5u8YpO4i7
WwjvuNnII3YET4pLRpJKBWX+mdzGzvPvP20o1sCADcNr7W7KFRROPUyxWhqlOpUy
ffIETNTNQZM55skh1CjVCQhce825V8leKkogCFgb0J5xaR2SURcrul/Fku8Pxqac
GJ7Hi8tyrVTQVKuQrOMGrmNVnT5mS373UM1Bl7LVyjO+tRh40/Ve2YMCFQ974VuU
VqRzQCkZK+iG62n9hOUtIHUvyw5zR3c/6/AXuQMNHkzsjvjNQl7twKAzIed9/xTS
C66KM5OnBkBO9tonvDtjFSfE3Qw3Wd1+FD5vvZ31Jz1K8y1OubcGsEzLpDArm1i0
ix0aMLE4+8/5MFNwBAV08b2KfBJnTs5F4IJ+o5v9yjnDiuDOYSTx6kiPpktoPPc/
eg0bqYwdjEL3pEgN3SgdApR3x656MENwCpzys23FH6r9o3sYCH3Nfu76amj7kqBN
irbtKpfJapmzj5IdIw0idxJpqfjaj/dTRVj8IuYQ+B6V7BE5Pxmpn9Uh0uvMlXOX
u1mBtXu04eZs/w6BwsK6HB9kin4Z19B1gQO+ELvko15t9C7S0tBX6J5xdVJWW2Xj
MpF1Qll3c03Z6+6Lx5DvuRqYhuuhPVS86pIx4RN7nB+Nel5wTOc2EtLrmPKEzIFy
1KtsRmKa1ktuPnfnBX593vl/dUFMOKfmsF6Ip5kp+G+9Ng3R8Hb6DlpTOV4eFGJv
u/fyPLsQyyeludgBUbGi68gB7I7ZU/oXCgtdbJHvLVPcYjnn5lkmwyNfpwYJJEbs
F7Lt8KqSBdWCA56w5OcVJxd0HfGkR8nb2Z5hUY6HRJJBuKQ/+dIK3QhdFo4ddFCz
QBIIvqsX50B0bsh5Rmidvb0A03Q54JZqH4Q42CVd+p91enUbxfkVPMkxQk5L5CBP
cP9AALjBtR9lamjrmBcfTWOGrIgYLuBOuj0aOo0z0B6lPDLYkKAuihlaDZfkPSNa
1ppjjgbIcwrAj8OFz8QweyAbj5lZn6+oPWeJ/aeUnAcIaYf0cdzHJCWT73eKCGUK
v5g8ssnyn4S1tr7/2Y/BOpX+lo3XTIY9I1hWtEj/S0YPfnes4MaOAkENT8AGgPVC
NsWtdteN6rtU7bLn2/aL0YGqG60TwKORNQqIvjRxrnZKccPpzLaLK65ljLAAB9ZB
jk+aEK/w3nMDFyYIkY2kEOcUlJVpz9GESHsoPZOjVl6VoU8/5r80z7UFHB2Q2Thl
5zWqMpw8PyRnuW+7DKwHovoIuhCanP2+6kslorNrdi9Znor7PBca+7K9R/G7txKA
t1C7ygxdoywMpeSCCuN+CU5pdpVC9gZpTDNUGZ69bHtQFiYS3cGGaOEzRvC3k07Z
1RahmK3SZJ2CFR245Qv3E8Jqk3oL3GkTKAPn7ayi+CcHz+jKe3PiOLUtGA+a7d4H
4n8C4eGaFqcH3LAlXn/0pNWxE9qKq0PgXU8PLg0+pc1FN8Utt9gynS6Ac/oWoprG
dJPDfGfa6sSwt/iJkEwlbdp7RoHWm0kSiZzaSQo8JBKhZ3SqtEzGK9+TTWXXjvN6
yXAwupqeWchxzCPHAKpumhNAqK3h7Zw6/vu9rINBBtq5CosieDUYx6Wf6nwKfA3a
EYDeHIGyZZHydwWwDv5wck7+vWBgtsXRJwXuvlJEfTDMQTKEMQ92nK4OfK9uT0Ji
Perl5dt5oH7+YOb03jV1unTMxfgrs5kxleAtKGhD1OuMO6tEBIzt62vKc/My02lV
clALT/TBtN54egyqV6XZwFfCv58YB5SL916C3rx62JPU7YEGuUL25aEW1uV5Uk74
PjnYpR82HVctQPy3GCe+xvlZtt7KSPArtIlPwK0qkufakOpYkMhqq+AAVBmY4LAg
nVzyKpTYK+HGQNsL6NUbpGRp2AmBax4LNPZR9dZS/h0iv+izNTikAx8cypSbAxDw
42sTZiDa4ph2At8fTx1jFvssWUm2QWSgB0U/zxQdWfIL2+Gq/S6Yr1RfkBUyUU3I
rQRwpFosQL6FG6UAHQUvOJPVKpOoFP0hRzrnHw+RqdEfA0SzTl6ArFm6dAW797fx
QdK90gXFQUsMEQCSgR+CFWfuMX98K1+hF5cBJsrvpc8Pqi5BnZ18fmKuJ2ynbVle
7ShrfaB+VnPIQWzgF6LENcM3L66isHJyCjVs1Ct/jmna9lgKPQl7Tv9Vag42Rz52
CUBQntl3a/OyqcyGj5VHksWXur70OUQa+YfUobQcVD97lSyBO1gpfZvmW+0awbjJ
apNa/5ZxpdvPXaGHFRaylLinmScnwxeTpq8HM8LOg0/lqpU1JqY055BR+aawfZsW
r3+rRzqDj7CkhGmmvMC4z4raI0HIEZ77UKYJlozXQGpi+/4L4it9UpBtjfb+UUAM
QDUuaYz59eZzOcHMCzMs+jxBfg2NvDxUtZaD9ofcAd8ym52Gdzgck5BiI86qfdF/
ECUZFwnCbWjcQBorGAqEU0EPXq3PeDoPt1MXLX4LSGtG7PLoRJIsrwWZiPqMt2wY
QUjmMwgPQ8Aj3eDU13oTdRhwo3ZunTahVJswXP61aayl34t2Mnz9H6GnbpnnPkm/
2F/mceNfhT6iO/pVMq1iecnfFSiYgmPWYd68deIjsb2PvegyevWRg+jSFarw604E
rZ0jAUjD6VDg8OMQAz4QetBKbwLifDtxeKQetoYEM8n9OlxdkV3YnHrdY1KxehwL
p9PdS1PWyN0cu8pJIit91ctXBgz597SzvMxmixJwluMYW2PGZEjDCbI/bbE0wQeZ
2X+8ipK8ldXSq0IoRmDXEIye9TvHxE47RGMuZ9S/toMtgoc24PiuGI55XRHsaZM6
Fd8Qjhi20G+ayVnWC5XDpvVc2TdEXFcTNO5Jbo2Qqoyi5AFqcsaICANirPLty6ax
6FW4ZwWq6LwM2ZR92NHy4g+QQTaB0y1gRHqW99riT+omritfhisT7WHeVwH7CGsZ
yJEuFrczPjdveu/2oocj7umoOka6lkJOVWfcMwaTWnYDROVyCiEtrKQESPrS4Kbe
DQzN7vyS+Se5gUjaK5r2xClH6pcLdVBopjAH9xtygLCrfhTLn6ISQnRucHyf+Afp
zqMgEYOnYwwuWBXFhIF634t6jVEdOVs7Ghte95ShAYM/9XSb6lCRuUbeRRgRA6uj
XqVfnqk68NULxAzt9wF2v3CR08L6NtW43xhv2dVXv45lNXripjNA/ops/e+eP8cQ
8r0bTSDeG5pGh+zLD7EUp94lLJDhD57SC3IZtqZDZBwidZRE/t6tnNkF3dA+xhoH
OzkgzPO5ECUHA8+pf8kQpoSz6JJ6pHb1Z2N5tyxbFIwqZJGEygoigWe03qRJvQkY
yGvx7+uupcvoKo73tTc5r63cfYCbNUhwT0/nc7ghE0aQXg3bvf578FVy5f2k3/2C
npiK7gMDuetmRGqhmwSZc77JD7JGH4qxAfBTGpJJOtgJg7dcq9zXdcC4vhosOsXq
fE6zWW7y6hQEVqMOMP40SmQBkIYphWf1mBIKoSVoIHExNZ2/9oF5jRw8cfKGfncg
CrFxCtlSmbkK1V1EUE39S8Nlrw0bdmbKmz9yR4Y0G7YlleW9t/F4ISa+PAiPw4OR
YJTaElE2RDIuvfezR1w2hikq07MKwksywkDHGxDnDU/Sfvu7kkh/trMvvSabzRqX
zeIUEVoAAJKWwGOWZiJLNuzToH0qksYe8qrhhkurMUQmrfJyHCR46AoqgNOmvlgz
dLlregciJJ4H1gG2xUz7EusK7kNiEGdzaUiWGZqcIWQymhD1m71x9/Dq+cMqizCj
/0/y1oVOl6+TmlsG91gejFE1F4noFVlVJoHaPSgcoPnCYHUOhdjgOUIt+xpmrEJ/
tmO5LI44GcMgJdF+NOLgRDLIi/pvrbDInKs1YVwAZE610vVa4x+sCo8pP0H6dvA2
L+xRtRsb3fw6FfzwyCnQlaXT+D48CX6XOo2d9grwEWI4ghKOTy+mDb452f/QC4ux
W++ObjnL4cQJxH7Jd2M119wgiyhia7YVYdaIvpF+WAnVql0O0LSVroX2GEuEW5bX
Jbh+FIS+7hqyJFj1P2b/ZZuIyVbBxjymLNjVHPO2wyJ+MKw1NXBVmaWHoLqxSNLU
nYB5WpaBHIq6JL4YyybsdiFOOoXBsKF0Ad9WLVli5HGQdP7UGsFYfKTu5Gt7rLRB
4Nn5/FtRNUwdgbEuHV2G+2aINsFxJblVxNr8JNe6Hw3/wH1hLf9wgAAw87CSUDLm
fkO/pvalwQglOUpiSGkXtCEZbrbpLEyBvQ3xsF2EclFaVnfLVFzw7WsyA113wcor
W8strYPYcDm8HC/AiFO68p5TBQUmnLdd1+E2lobSlMkZK+4K560yQTu3Uro/dG6S
4FqAIPNj8Vykns4p4+3DQQEoqhkSQzUTFFwDHMsIlNNVxoNSqGieBIeRmRbQqm7b
L+ulwpZAg6xc0MneKU86fAFEtHD7bIZDK9aQxtl4Qp/nGPIZkK5CZ47sg1LZ/Otc
CoyIvWEGyUs4E0pzdUflZaMfKi24yUPJJ3hBrdICJn38U4rFRveQhrhbcAa5G47E
vhH/fs938nY0si2qWr15VLV/ztoUQxRqsQ/NH57IFPyi+1OItPqE1zkQtUc5WorG
6kMNP2jqFliYIkvOctFekYr3rBS05cL3kFyI304ZiBrF6DH1OLtL5xxl0XR0aFB2
UK9yYdt98nzMb6du6L9gI9m3ErHWiQeowhG5w4euCnt3OZxdEEBo47XaKVPYpqrD
iZ97Gw+g+j7GZarfKPQTisDgdiY+wvCU8EZ+o/CquKpZrGjBapxBEkqXeShBvfR4
wh8J+DRF1ELf5/10gRd2oKbnSCNeg26HTpfmkhX5mxsDL9stWBs8VxBUXJAFzXsX
K+axUOYuvHwA5l5zQmlKZzwQXb2oIbXNGyNP5Ma5EkAMfTE65vG+OWVdnO3fPra+
3aWm7yUT9vJcmbZbCfhZ4YDHT4hxHGdku2ZCGSrjGuJQZ09LWan+bE083p10JRtR
4jt4iyoiHGzz7d7rFxakw3TZtsmSWdUXmoTt8LtLWlGAl765RJyu9qGR7rDsb7va
gBVmvckQmbQifF/RfjEik9NwteVdl2HXENQGTq3Ilp/JC/0skxkLh3MP13w5B5rd
miC0WMmz7lRwMsbuNfWVuJlcyk6rpXdpGlhvICmDktOxjvWhLjV5juZyhaEXSTHB
7Xdh2F0ech9eH0E/x1umqR22lkxt/oMgvOpvl1XVmw0yM2+86lFY/GmBz9kBoFJr
b4luDwlmNl1XMph1FmhJAnV2D/LRik3Y1yf/Bnu9cqHFblrX/HY2JIKIIQTAO8eY
gWru1jY1kdJqOxzEn4xQ2t1NKrN3UkamqlstZv79AALuQozDvmWNKfk3Yho8vRhF
SYk+d4gyfrsZV4J9Fxr4HH0r4ia9uZriAXlsvx0wGzO9K2W57JmMF1tZIWuls+mZ
fjuhwfqDuXTjxFDn6Tj+/fu1M52a0XtKyW1t57K+NSnoL0X9XhBzf0MZiOPzZfJ6
Wxl4Jle9VyqbtE2QQ4CNE6h0o9/KQRfN+v2Gqnkky5eJc0H/UMBxuW9JvzP/fwD/
zMTXG6cZiMWsa0y1zEzqNpNnz2Rk51PmHR0iuSFSI4/5DY+j/bEWogSv+Pp4Qu/+
78+ZB6rDWFBZ+2sbf41utgzQnWqZ7U4t/T5o6X4q0B0PJQ721XgecuAEENgv7ni1
wpKiRNfr/5Fr77faeDTpfWMaq+HnNcBaieMe9gqljsGMEJUSFQmIV/hMoR8IDLZO
1Dfn/RnickRBEiWMOZf4qkSx3wxjysNy1SoxM+V+A8HEfA8KaGd55WEDKv0ysRgN
yh6U03miWgYxRLXb0Dv/RtF+LlP4Q0ueU1saAVsZcjpZA+d0ZuKxRxR9qKT35umO
I0xrBXCYHLqzctzYAfydATTQnqguYssxYcV6Bjp4YpfVEKLCzVe/z90ijl25SRe2
TGGWDOgvqN05+kpxPn710q5qUIluz+uAu175su9SLpt6ZdeD5HsoC08EwXq8rOaF
bHCnGCuRVmIzdlFxA7oOsRmpS3jWmvRNSeuYd74U40hJloPMjzEPbHEEZ5Au0jXk
2vpEQ5GG6QxsuZLpfDp7tIIu76aFU16ndwtDdN3SKgx9OLJVSlcfKhRcpqLwMvKA
CxQNi92veEbvjEIiNs8x9QePxdoeWjPvL+CslxLLR6J2xnrapBKNdXrUHNke67JD
4+raxOnrOlb2wF79RFEievR4Mnp/UgPnTpQcAXbAzGT8UeqPmVHMEoI1vJTrmEXB
2hZEv7LSeJk6wuj9Mq0NlgkbLZzNXjBKHuC/4ce6HzP+xjXvfd5XHKEE+vyT1n8F
AQ72RVCM+nywy3CLXOnW6kR1uzRsN8tg/WauSZWuqhJYUHlBlSkP+Q0MqtTI99CG
sIWAhI4LXP3TSMoQ8hsfKxDnZwpkyUdyOC3NchR2NbhO3wZvjz1USgktGoduDrhq
FKduVdoQ5KIDNljqXayH5FydBo46e5Uxb2lYz2RDt/ofXa9Stq6b2DBr+ulBIxRl
APLZfo74tRrvuVEjb6pmwpQpgzZpyZoLYHvL8dFf/vVV2R4EdKtekdkQSZvGfnxf
lUWOieHjhbxlxcLeG4grq7vBZsQl1aSnpbKVO7OWRvPrmxeV2+KxTdsxwIY7x5VO
LQFVM2ihwoeC4BgKM/UrlIv2TMaweqducsGuW8uBsVmz6P3g+X/OZtnOrfZcj1N0
tv40XNMpD6OG4zzZNGqOtaSdtn+sYK1U98N7ZNVSg1B8kKWUkv/sUUmNEQyHsL0J
U3hQUpaFFC6v04PVg2X+OZgX3Xqib48i50Ap+K9SUbB/JHFebqxosY4LixqnsHkT
OFWEyIfeG2T9AAzX+8zgMF3Aja3XFN7PqvJCvoXdo5wKM9zrWLPr7uEHhExmcd5F
7PUSKNdJGOI2uo5JxTV+VSTLGeepKIko4lPW4Cwmxb2NylAcoAmnTh7koQRrgg53
e2xBCdYcIugO7fxuMjThVU1RFxR4jliwDHQIRGQ2rbTJg5b6C92MoYpCpBw+tSnD
cpQrHkTyj63OHyKGRLb57BCMvWE0jYvGiwEPsq8yOlY3MktWAqzJedmrb/KOJpV7
w5i5iALnkDhi0KVLtlsRBR7Gh+l9L9ix5S0XtagdMek8xpEdMb1Wa5WOsrp1F/6t
bNFiIxsxLI/+EXnribARtDkmb398h/gH7vv7ZkIEwSUHF2jBa4Ao17sis0QPOwd5
BpRJM2br42GXRTUHNDXJclLCFouyFvwzEZqbHwV8zwVx6RmopErG2rZf92I3VGTS
AY3D1m9uGkA8061LImhdXbOEVIE9bWJnulFdb1qqtCQrhbex8+RmOqkCJBVAHCSv
di/O9fp+hmRAKQvJH76uHu3BNSYFTChyxiyOVTsqB8CB7iJcDHv+TfhOwy3aLrAt
PdO6WAUwo0ThNjOhc8Nc+0+eTHia5SEs0T5EgJGDvDoy4VbdqvbnlJGDl3o0adPn
7uh9eyoXGPkqL/HGhIiKg5HRwTiksICyHLURxQowtKcWyAc8GEqdiJKM4aIkYI0o
6JWpADKDziBgJmCs20VEmhXaKz5a6hUpabpR7O0ovLwbyitWb0Ir95lfusxtr+1J
AtbHBQ35aXPnztke7Pil/I/OrAyMk4Ob6SqV+0EL5oPzYbXqXyKcC7RtWSpqEK1Z
yKkUOLq5Czg5jr00n1cCsa05/wW8HLBZD0mFP0Ltm5wYCWCQfcu9APIiJ6hWp1No
nIPixZ/KuFMLm4iolJCAAzfuXi0T5Ur4MNvxx5lWuvEWmonWxVVWlZ36SkM3dEpZ
tCXYKEdIBF6RqZFsPIQYLWZfxrXTL1WkxuhUjdEPUSHN3MZ+/bixw8fSmu3b6D36
nRnSZy1RRlRfLj8k7Ze7KzHywBghugsNH0r8zcH57YuSAFlWPbzrBJCliViNDKx5
zBlFBgKq3jO4U+p/E+6XqbWqeHtVClel/mB6pPvyX1zbTNgrnwD5IIpmtNiudeZa
TE7mbAeBA6UXQE3NbWdn529odqka/UL27GVFG2snLJZYmJyFfeJ7oi6Zz10OY+ok
NiJ1h8Gtzforc35GpORhumbSpIuii5hMv+nl36ktIvhB1NNx5djcr40jF7UdcdkF
es8cLWRrUFACBU2K0WJIlpNjD0gA/DR48cZiSgbxEIOI0dZBpdxPS34wfNyAuiz0
ikPRPF+S5PXi/Ivf0RbvichezMwVAq7ycZ4i+0m64t2RTbztxNwcEJbogDEzP70+
uXoDLZ8xzCR9MiK6JCUTDp9CM+q4ws6Zw5A0QE77BRC26GFrPXZMhFcJ0BVx9CSl
D1OuCzv4pK3F4GEjI1foA3fnYxjV/laH2Qof2ErRQaUd3zX0Yan5XNTZvzIfKtHv
eTqfg8FCFpZ3TUArju5sRYGtaQVMb4xujWH3ETFnv9GzfyIOKSN8W3tjGrszTKhr
l+foySUZ1RMF2wfcy076L/KHxSBka7IhPgON5LWqdoKSMRNZceqTJg7n17jZzr1d
Udfn1cVnLBV6efdq0MrW7xRx9mDzlvq7n9Qp8WUSVhaqh4HHgMLDTVuTYRNnrkHo
NPE+A/0ykXMlUSR/A2ZH3cZjkanMRfPIA4Is65gjXhrNy7Cc1Psh+rxdfJCbYk1O
CC1opG+1u72sEKqwL3Ak+Xt01Oo4eZaZhNw4uA0sTUUUJJry0AeH/ieUjB9Zh6zt
Y08/Mgx3CaelMjf4AxylF1FM2EkD+XvFRLrvSma45vW8pnYNdK48OvArZo15COPG
GzdWnnDul/QMgDJi3ZaaKU4zm0o8k2hFESVN+aZPRzzNTgGmVtPq+tVce8dnhpa7
QfI1kLpodZcGu31U/iPIQqUxqz56CixG5Bh6Ue7u0DOkFhRK9DChQaZXuPVom2X+
ZvnzlnOq9SwxwKrs23OYQvZlTyxJ5ktIVCqucwdNiNXJGihOrVfIoMiYYhg9EtWf
OtBwwuBlsV2RWR+V7AIv3xH8iQDU2P3SuW/Vb0ydhbELdHqC8N2hO4Mvbjk445nK
GLZxH7jbr5mLh+xJuAcT9p1+fQ+O843RF1XLFvPo3uu17WWHUtcCFvIJG3BvQxCI
a3JxgUcYC30xg1Dm8rInLX7pAqoOP4PFipSlYnrUHxVocKuoFmeT41Kb7IKyrsai
Iwjsum9RTldHfRUB4p9NmPMFzsZuM9bN+UpY791DCxx2AH2er8BtfwajgUdmfyB8
iydtqyJp3gMfThN+276CLlOTl9oN/9vSfA9/zeMcKqv+8z78HwEtfvYJZ7E2l8Vx
yM0G3Khvxk0dMsl7YmI7H+/iP803D65ykAxri0F/TRn0UVYSyYn+j00E2wcXRqaw
XJrf5ZyWk0yHxGLAssasufGdg939uZ6hsQw+iq6R6rMb+hEV4I9OVf85yba2RI2T
EAE1TeQD3FuRnr1RyJLL+lKaGD8lbYRd/Amtf9xcSRcE29WX3Rt398gC9856zwBG
XO+5SIoDY2mcDaEN44PFEjMvdiJ/brS+PfqnsrOY/zzfaAahGCbLQkiSgTsTJq7k
TCyWpUCUEDeKDNY1s8o9Git99H2qaXMj2Ooj8jvOLWLRGT+062auSH3ykoRPgu2B
dXzsrwQ2Dh9AVuEEEzLI8gs4NnI75UjHHW4uKmr74xChQd5F1TCtOC0x+RfMTBTa
dkEqxmI/AQysZx7FCY4u7kBfp2ugswzNpcrOXlA2gdnN5aULR+F8BPepCEwvjJ6U
M4UYb2NyL/LU4iogqMnL59Gyo0HMIUOzoxP+72lZvQfMti211K7kU/ZBqWDuNQOj
XBP2TUpYbxIT+FVs8dS3aDSO19zXFnHXf+k085+czjjT0oY6rzB04CXKscIS9Z/J
BYSPkfDSKGo05qzrmHj7uwW+0ZT/dXqpHVmRu5eRQKM2PQHytRhj5YOfotYGzCiE
hOZ8IQC5nY8LPX9COaF5oFEbDuZkNJqn/1OMX4xQcwBW6MptFwfkW+HoF7qR/eLZ
+PyY5z+Nn4vgUDNd2OP1gVXBANrxP3RYKZRehHpZ5DqvbLLTr0Iv8DFMSz89wUW0
FbUiXNnVLFoT6y3h0v2dOnIjDo+c7ajFnUHoZyJRV4mBv4j4OdTG18Tm+lVVVa2e
T+GYEFGlI4nkTwJ2iCoGzsP+E0pYxCdMtECKynNVjWTIEtO++99ebiDKQL7zoO4h
jRaTmK0Sx3+zunO7l4RipQf4dCT97hKMGCfhA5CnII1JQKOuos6uF0hD/PadGxBp
8tuj+0tJxvc7fM5vRUfW+Ok7IV299gCCIemDjQiB5QPI+Zs5DQqV1E6W8GtFjN1c
J2pe+MNkB/JkZJaTySjvfHdM7bEReEYLTUwqp7glY2HpdjTM33z2EjwTrhNZ6VWD
eeJ60HUA122OAEAZrrWZkurUTrgjbJDpgaCNMY6DL4RT/s4qURYF7xuoNxMbdCF1
NcfIKVOEpuNPleZOOw2czIgeWknEBuLs69G3dNWupOe4aijv7lsOxHJm2D/Tu8yA
synAbL+bPeWxweLJzCPphMuTi1t9QZrMGgASs7eVtZDew9lQCSt/BOLrOvjwaypH
xWBsdbwNVknbKH5b8Xi+HkskvjHP/+Eio0RwIlomJESv6gVZKdSrsGlvdIBNbkTs
fGw0a09xf1ilfX131+kuE8gzySrL8mASN3jX4vsE5mcrHNdQAiI8hknzhJeBkmGu
D3ZwpK5XTj196vK6jhFy66lkudgkHtJgJ5UgmiaqSctkJNRFfHiOWNoDRjgb6G8I
j4aa3Lyj3Qap7PcFLREMSObAuiR3pHY1JyLTGmttBxn2ko/FADTWALvutqcIn9oo
8wmixnWoBQ/gxP64OxuH4mgJmUX9Y546QpOnOKK32/lHBnJxgbEOwr19fYVUw5yO
Rkrv0KhapTDXL3JaYYtrM0d5FVW4DZzAqefHKZCxjRfuoyQxQTUkmcOzpfKhZDz/
q5gCTr+fuqcUKOG1h3qnOB949eqi/9v+9AF0QSDa9BpE+b0CTSwqDThzx0sGCvNt
yMeyXIMXD0T85SNA9vheTL9+qx0GbgpI70X1U2pDG00apLluUpruwgMnh8To91br
HpB7RpCOag4kHMOA2puynnB7E/6+abjbxn7NATpsSeqEZIFhi48JJzgCYfPjSNma
uiVh0L00mt7ZmDgla142BFRY1FJ+qPoUyO5642Pn+aRSUp9CYEx+A95y0VJMCJlf
X1aeGqJvlQJIynVQP0j7927hzReIzXHSj+npRKzSVLSw/1o/MjjkAwLVkRdETlL/
GkLl34D6hOI80vnzesQjW97GB/2XZwJCNR5SeVODP23w9cMELFUP6FQ/F2P/7uSK
CppryA3TWW8/UTw7a3L9fgS0SM1wy3PhiD8hwdKOX7xVSSaVgsyR5tLN5qDvmClO
KopJjQUyw4eo3TllWGJ34AQFPrLFuFjOYVU/ATLCO0ZfcoU/QaXNY1ykB5Sgbumb
Xi3YCVeChqE5Rp3u9AkusTP6rUqG40uXgjzfcLC5uLvGkmNrbge099Nm7nQjMHRq
91nQY05YQ5F/vD/J++GFc0dvmQg7yIKyeU2/sq3hQh86uuosPftBaU56sIS8YmQO
YLBSciZX+up7hxqNGVqUAePL/2V1u8KAC6xOUPoZncPPDXKK0Nd8XVVMq9Z32w+d
USOCf86/5u2vx3X3jWb1NxZpYcSYYQqBd++kvATBdTEQSKj3nzIXedQTDV4mDnZ5
Z59QscBnKAHspM1YXy79J0TdbCzIDqNOk7vyNCa9zsiRGIzOF+v4vAsVOepHiA5w
d+we4kcz/1uJlOW4OkO3eaS4UtiCe+JaXorUm+8Czr68+iuDuVrWEhL7dth6DGDj
GtjkxjINO9/iAnICAypt/fYkL5qjG//+Q6yS2zFWsdaa+OgCP23UDefeV5UxPb9j
MJ7icoguV+PDcBvdzFcEvooMmhSW53g+tzVg9omNshSfzAelMTCGAPb/ZS9BpjDu
DSOlRUiVMalR+Qo1f7+zgpEQM7SXjptKlcsdNG3gUPbPhQpVII5VeOw+S4PqN6Oi
/eNYfVK+0SzHtRcSjcpgYvPMnHSDIQKz4lqov3ZAd7AyTEU86Yycq93BcAKHmufv
7rDxZJyk6yb2pfZsZVtUgj1U1Y7DXT+jY4ldeO81NJKgWlbcRALynCMMnq81uhjh
Sb3re8/jGVcnQfV1fmfLvyUW0K2UUZFmTM9asO9Av1g3MZVRPV/WqufvS0c0PWLe
Tl46qiufqBndIs2y75gJr7Gu5IjCdjpOmaBWP4qxeqkypbK6Ec8AVtTtfukqeajz
eU4Cyu3kfOlm2sD41oebZulesquMv6yoIooeqW4uY/jklu/hzjmFKivN9tmD0W2I
k0YZpD+/w7WqLkRihIlGl9LbLftUXh4S0pFm0HhrFCz4IPHVpBY1tYc9T1ZnDE5a
sJjOMxOoRazuSUVeU42+OCct0S7H3yN2/DYE6Pjozl3NHxaOwPlyQqZFrgnVBSt6
SQ8hVZWLbIY/HQUmhpx7pIdjImWRDM/TII9YhbKEFJklZJ9wJhqVmFbFwDrkwoGA
cEWbvH6O80C5mUG2FiW2leXM9XBsFktEzJDVxq/CHKd8ym9Km7Hl+Khv9vFnkKV6
//NVfzJUGU+wAwdm8tCqRx0OwUhf/ZV6lXXo4jLwdJxkqM/NFZ30SgVxT40/WxNP
O2y/V+3CHmXF0Yf3xlvkV4zBzvseB3zbrL+XUTzzlzk2Q8D2V3jFxnIE3Urg7IN8
4OMMNvhVHZ82ZCdQBlz5M6kKOjqj1Xdp/VQT/XS4C3F7Coov7y8ChZam/DnNfZ0y
7kfyRx18/7le4UsceILzcqlNMkQuBuNjB8/z4ZQn5WRblDPCRrVC8d5Lw/DzsBJa
zNjjFUZd0g59q1UG+d8DbxQ3ItlfdTnWhHsVapl8tzeG/UNsMqeIlr4gXb9PqXDi
tUnPzcnoX/vsaJ7y7Z29DUxB7HgzQVQfcXaJWS5YniHKoarEeM94HH3W4hDMZeC8
rBa1Fp1VOS/5eyqlwW/HXyImXTVKlaKg6ftHAapbsMsSlDTWhhiSr+PVTIJ7wbtX
mwtxTEmrunLE15+N+2XXStKtfIVSiKMsxbxCItBwhU76NgWHhNRQlKjozSIpd20V
kmKibwfIeAVVEWWRUy7+G7tBCofmGgzPnBXCl/ycwUM0on0AAkB7xDI4qXCQgkRi
l0mPW6zRNJ/h/OX12BGhzxfsLbKtXFLyc4uPjgAxEhimWd1tcCFEhAAcT+ic4Xv3
aKWXr5FyOULvMzzIdc5pS8ymBqfJJHRJtrb+KdmgQ6SK0Jgcc3UyYkBk+4DBfFDY
sjwt7AHEvJwSYfHM+6j5Y0lhdmyxzl7TtZc2aK86UCpEuHsh2dbZdVZ52yfCYoGX
e1zsakb7kxROnW0B6bGIa6b2oKy58EPeIO60QREYMFpS0PNgRyFPy6ssrybcuTyh
GFsCBIwaPsT7ikafO9vFjYVUNPlI8HFpDxOn2saIP9HNW4huz5Zm/5HWa5bu3hyH
x9nWZZs2cusNZlBDoI9BKcBn2XhoSB0GM0vy7YniVRJ0kHO+Rjq1NKsdLhRBQjJR
A3A1pxL+NBGllUHk5Se2wuGVqZdkcoVHCnQpOSYEIy/SdCo3dPAjvYKk99nWIXXD
PI2nGcW0aZeX6dVCkWIjGOSI7owGIXObUQ94ePg49Q040LIfhGPfnBkjiERoZCJy
1nBbGjbmUgvfW5KU6rLY/cgdjJC/LV6q5cHrPIx51E4yiyDoXggA/KHDh/LAATd1
TmPlqWbo1Ys97zGj5KlzRAZje9SMe6mv2TAbAt7eZjSFvKa6OVkFLDhWyF6a+wiQ
Jv/Hu7JfW0Z1pUl0Vy27ImgREk6w+MTzWKx6GipdKWa5u13cfTxmF2MstTeR7Cmj
44KQSDDTVfqxFY368myBRXbyZQaXffrw9A4nsC1AECivUoe6t2Rz1/J3Ww7zlm+0
R4xy6kBVbVK9XpDCh7u04I02cJN93l/nkYVJw7WH4D6Z2PxvEqqvmmjVksSeHgz2
NZGBT3ossxoH65sUZe67v4TnqqnCh24cMQSiIUkPXxZr/EquMBY07XfsWg2yAOFo
3uQwZaHQDw5juA8VGdVVr4fdReZhtonVrQ/Jubb6O9+VDGr1Vde521BSWtO5nBGN
RpAKVm0N3y4Nqm7TcOkWXMnE49oyrgmNIEjDYmrCC/ggdseDi82hDuN4KejTa8pl
U6blZmbZZCYbC6b58Vo/WtcKZK3UGgdJ6TGqn9FmoKGC/5pu7UD9H+GfxmI42Gu5
gzOdHo273hGn08O04BvKP7Ns8o3wusYua8cn5IS+qySw5FZ9uouMW7zMZqJ41Qst
i89eHOvC8qww3FxKAutnGbQbYWGqM+H4VWzCyp+b7+PyjRMZyxtN003ptf5XK9sg
Q/N+j5dvZfq2kjFrw827Z4moZCGSKzJbn1HZGI8dvn97GjHNUEXlHWFqiW5/kTrj
HoDwcpxmRi8itms9Rk8Y4pFrOQte0PExXjL3JNrA5AAz+vF7x1ZarXwA6T304e4r
W29auVsZ2zAlxSH0bI3J4OBvEcduRG97IP6N7sBbxei94KK07mplSQRFpm9wOAeQ
w7nRYcA6KIXwqo2q4kbSN/Aj5A7ym3d1oURI7FyPHp06vANibQvsQIsvfbARd8Ji
mTTk+PUfrdyCDV0WG/luOKOI+74p2H+WNvueVYt1bs43DvInvUiAYAY0MraCwcI5
mCJA54h8DK94v/3EPmeGeMUJWvW2qt9NUCaLfhWoRFfiZz2fPoXZkPP5Vv1pJBA8
Q7Lqo2xFekiW5WHgmnDXmRBwLfT8DjIxpTD+tdCWyjP9L8B4D5G6qwlF4c5tEuaS
Te7BLxRoc2iPwB2nHxIGwqcQVg6MKHyKq8S4b+YYByxozrtNvQPVdCbwlYFyPM7t
2GRmbGBqsw4+Vv13Qb+XOJyEWOQvjH8+hadjRMR+Cs9zbAG59JsKIQW/6zL2ENzK
DA1eKYJEXjjhI30+1KA3dQh0kQ0YT745iCRJFApATSBesOyfNWWbxbHwkLqXHUZm
0HwvBolrzwkSvsbnhllOxDuC2b08quKgkdJu3lYhFdhx1VTgcMBcSfYEZel7VyD9
CqhA6cNJm95L7BFBE2A9N5gbfhzYKXHliKVUmN5TC/oeg0mEnRiIMWzMU9dyNBOX
43ICivNdMJW9ab5BA7Ud9Q0lBCBsOKELVlrDvToTZMyNLpVGD60LAWhRpiT+1uzI
2Q6URbN6O3pH1Pj1uTPigfBoVczesNdSKsagbUIuFye7wUT7dlL47qoIG4fUKBRl
TEVvO6D2+ij2CJzDLWUXMgrdOxsXJaJ4BpIPx2SK1vGz0R9NnMpd7HewZaZeQ3VI
c/jBn2d7bkKZwIO/cSMf2CrAb+24dSKdYiu48IIDr3I/zN/EZLj0ghyy8DnjZ0i1
XfCT3fcDYYqRoWUuesb+6c2luvNx7zKKhdR09jJUZDsNLAanyJ+OaVN1iuBd9z8f
bAU8NvgHvlBx6CLj0BgoyA07dH8xcB6QSOLb1imgbY2tcyh5grADnqZ3vmFYsz7n
nV6HocneHpMBURTL1gifqGGVTzU9MhIEDlIGb1dQOqPBDWmrK9ANOY9z3TQYANzC
lp3KRnJC5EEIGp8mwh4WvtsgEL+UFPFuTgkaDzscppfjstMZHDZVX5YldtZVKSWZ
Xfs3I14YveR2tKq/J3+gGiLJ+pQBzoQmRbIQgAXXfoQaBP2AB9uCpQEZ7apj/xeV
CvTAB7aRP5cpupb2BxN1YN9sRGGvK3DKUR6a5P7jwfoqqPyR07GKsaSpNULikc+F
Ow4wfxjffMtOg4x8+52QMD327KyjrlIrVy/g8AsBWfiv7YWe6wpZTYjALbMLJtmN
L3v6RyGsFKxR9XijST4bOhOTPwahsDdGJSgq5EmeZsrkl6ETSwDiTnKccZbk0fiV
MmL5U3cCjk02vVFFVRqwUojJ20c2shtWNMuiynmtW5Llm3VGNM0YP24O3sWupo3O
wuJK+tIJJ+hr/bm9QCksW3imCiHnJW8MAqf7ofsAg9ha0q2gmbIZvOzpmvLm+D9s
L9Kj4kV8Oa21w5/K9LzzyPMycB3yvf96q7EV/oSCqGQgKxb7CQ639Asm1F/ljLku
0MiZ1oV2Eh96Q/qnIc/5jbHJIrWzqyU0IQIF0h4Jw5e9uTXTIY808Kna/uauilhg
Msoie/wHAjSrIlSgt+wyEzKaxpdIOeodVllLLNqE2wActTBmthjzOwhJbrfOFNG/
AUp1I4TVac+LjHWajgxHK6G8ygxBE/QoDQin1W0Ewkw6Jf7NTD3pSwUZa132YoRH
w+BGNrprPq8Lj/sadIBClmGAH0uYyyqIvEHptHQUkm4sY1dmo81H7SIDJU0XVJcz
ahiAXSyXtx5pJ5YqkcI/hDiVt9WFQABErr3JlwjfPjrj5t3mkYyIIBSNfp/PvsE9
B2l6xEiJVy48YI4b1eTcirwrWynLP2F+CU68DhaILQrJyRfR5F8tEVgxtjkQSdw6
71usobFGLGvYH/WzLvuv/FbpMI4qSiS6fzOVRtHoOdkmBVr9WO/GadMJ+GWXYcxF
Pah6I+RAO7Qs7zA0Zs8zgLLgBttWf/uwj+qlKHvOqWRiSGuNF8rTKRP/yd+jydQP
T5fMgFkc+4vniFui/N0qQk7kZL+UCzk6cufInmgz1NGUN8e/Ai/cIq2SfNgCHGnO
tgnPAQ/zdb7CRZFmgJUPvNf6TIN7pJ7ADlrswDtwE6HAjBbMtv9pt6f8ffN4e9SU
Sqt8qs5jOHIa9LX/l4U9+xPyFIM3sFQ3D/h5VKkSqbJDTRRP/Js6mQ0nITtP5CYS
26TA2nml4ydIufmhcx1vV9a0Uf4wjUrkENmhpINVTqQ+ApSp86hky0bwL2YQlYz1
EHYzkFRqDBhZEfpIss8sv6HOI4xWqMt69zihsl6bACkyB7c0OMbYQ2wq4ZA86vsc
Mv9/OMO0pTXYHjAqgqO5m57rUkiPlFgSBaMmVtisn83h1spiNbOIchTHlaYEXBY9
kdjvlqYzJdQgG1cIE8Nu8LAoaIcEHI/bYhUvYWNHNo/tN/zKGPXCFDVWvws9XpJq
5FlSR/Sn8djew7Gj/VPCae2ZyEoctB16ye/UHkTUd/cHue1B/X071CqoBauqHF0F
B6aMPDQkNrby4fxYEd1eVfx1YW7xfFvuwS9et4D5e9Snjsh7+4LZais5+JbWycna
1K3F7A8KJfoCqQrEkZc8b8kH8mA/gZ6TMe/c/Ro1C2r4PxNEphGipwfBMXjmWH5R
TBSs/q/9oGzzEfOMZTSQZzePEVCi2TUX4mO1SsS5Z9qjS+Ytjx3va+Sui92n3+wY
kzE6lsZ2Q99RMPMYe2vi3Hhc/LyBvlUGSj/ZIFF4keMDsTtm3mmT1vbLcLck6h1u
fV02245jJKihhuIP+Hkl/+utX0XZj1VUaHERwZDewcBFZGkHiJTnc1v7xZUiCbB7
VTB7+iLTYdTXW8pMIo5pV5YQZnFRp7aKVeDapA9Rq+4LMd4LthmOYUzL/moBJptH
tPkw42Ke1j9JF361tkihVLKS9BphFLYtTEP2aYriWumD3c6JLnyhVufizLSaB2/1
gBb17lN+fWBqnH/b3+AeQAAiWORBmZcf5Rcl6zlJUZ7KhkbEzub0BrT2Z0rhTvJo
IuP/ZSravikD3RoSlP25cm9/GgZ+16XhydJw9fL5PDxJ4J/HUvL3grVy3orLtWdk
WAMDni0g9zuD5xOVwrvjGCD5UVhaC6n4jY8wfoZREu0mzDgjTYzQQ+dEXvIMrtAo
DUtjorlAu+X5GeTTUNI/zmkqqS3/GJSjjnLxSd92bEGhuI/iafhAfgGUAy+RzKZJ
L00mtVjK9aha8DeBdz5e7BYMkuV29S8uYWGK6TB/PrmNTCEzp+O4vmKJjNn80zGD
0chNE8CSRgpLPOwFTIdwTPkIgt++QIihb4BHffFrb/0qxUpRAXDUJapWUciRG4hx
wB8xcZiskMEhOmv0rXUicDTsSOVxGoJEMYYainqD+qcmaFvlv7Yi037j9kb9dfaA
VNnXXSCMADFBLlrtHbphl5sl7nHFeifvwzAbi43iVUJRxgtf/MsHmhYE36nx0U74
KYyrb1L0Lx/5x1abn8V6x8/iIAgRkxJr1NWqJLjvTB0q6Zx3YO3lEt0swACnxyaH
3dUJNokVR1fqlurxgorqRZMCMFoGdRZsT4rLfs8c9VCd5IbunFKWfPeNyCk4UrGK
E52DzVncKBA1Huoip92+4YxMoyQMtHWqrcUNmrIGHdc1wS7PwcrInMRyyRqGa3mW
sqJFpFQXnQxAtFV9IkKPLBK4MIuK8XcuSUb95iDitAGpcsBObJ09ggjca0CrU6tV
EGQoI2lYwgTBAyD9M33OgZKy7L0ZbGqJdnSXtS/iTWnE1uT/oTyP3Cn5qAOHWwUZ
WC3EMIErVoU7LY+0JtMCNXaKEwRcPBlN/ZwkjUdjrccEYnGuJQwJ+M56pFw8Tre6
RfqPsOxs73GjP2FuhYQdAv13Da8OkvWHl9o4sHE/87HyW+v48fH8GrJ8TMHI9TqH
ffXdz6I6zJ3KmV2x0iQkfcvk0YVjiePS8OqWeqgYYR9hyaTRIHmGAaUdrk7GAdKm
50Vin6L6My/e94nneUDJ5Z7YuDRf/DgybxapuLhwQwjlIm+cpy7eO2Y6C40WYwg8
139EA7aoty5WypQfe+/UAOlFE4BXiSqoVpRrQ5JOEOh94xF0kWmsMxz4QAhW0Cxh
XF8Wlfqqm3WR7PpydHhqExr19NsYg7VLVChV9BohKQjLMuz0VCCua6LXZXm1tCE8
AT0pIzcG6U09kQXtx8yPfAV12J4l0aNfeqUQNEy87KHFNLwqDgc63/yrfsP+0iYb
TdBP9rMpeMBEj9ZX91RHjWLDMJnlKJEDOAjvid7Mb0V9pOuU8JW93j9iRZXvI3t4
7faJcNgFEFGov1+sl09xhjEClInnERB4St7MK6HqwjuxLWg1i81k0XwGEV0CVsRO
LN+sZLJL2QG6CW118zHyEMGIZnxv/nH1g2kZXeZxypfMH1PKmORiJIsW1eDR6Zmy
JhzG6kScR7DynCeGtyVzYRyDg4ITyJfAlWf7dQs0IQExaO1/Yiwdnn+sc8g5DbXK
irKsfcw9nhAwdy49Twu6/Ad2JaEbTt1OvFeyIfofMGL7BeELKmYf7fer8zhlfLQB
TUDwP9g3PFDHjkuY8K7bWZ5a+y/xDDXKOucr5tO94qDM91puQ7Ez6ek3BK1/EVNc
0VMMRX3dQap2QYffd4YUuOfsBzcb1Li6wiHaPqUG/2bBgZWvC1FDiDSvI0nmRqHZ
Jr+Bd8HXA11XBIRyVhu703UAgGMzdzT1QICkrAn1wZoGIEqxw9WIqw0LIDzYGDs4
r07gvEpZiRNfJvr6t/RvG81EunGEPUsVt1tgrstmx1S2oG3wLFkJRljpF4x4GmXa
rWqwbQu+/ZaU00R1YlgP7tySbvtbyRV6ufxymV5LokC5haFFgvNsTvnjhNJu8d5z
jp4xYFo2OghCpYAiTQoC/v6q8ZWUTvJRMVy8fJZeHHxVff3WcrW35cVOO3773Yag
VTKJiaeNWySjwX05PhmQd5elPRISjaJ1qbaUyKk7UZKge9RwfIte2Mqb3ZH2I/ag
HqYj23dIY99gJTB/l4B5UKE38XG60gSJGRxrh5XzxwEu91dzFv3PJVbhuJHMVMBF
oGOoWNZS5O3qnGlMT7hz1z/XxWOzEO3zOcyWEanGqWBFOyC8LEcvSpkuYUNZXkVr
C0x5UKigPdsDgGbjYv+fa9mrjUARWMF9HKw68SjuDa+14UcEGpV0Li97YvywugpF
GzAsYcGWgrgQfQBACLj/MqQk25HINi3RWBbLYS0aiqJQzW/zR4d19wupFbA3YSoe
Xb5yL0GNtOO2Rl3+8eJOI3tpu5r8qGd40DwfHLHeoKjBoulSfCoEdj9/5c+4EOjH
jEAWIrnY8vYJ/M15qE/70BcoCViYaBnxgb4ud5NJ5fl5u0AmYMriP1/Igd40BELN
5Q0oqUK2Esk9xZcaiefw8uTWRiTPJIcwSkNKIB7elQgKekHXUJbOCYtwpY4WwsGl
iu/Z7lt5j3pgK13L+Za2D9DR3J00TDUkURWOWSg9Ct0Jp7L2QVuxEOQ1JEFsL3dq
rvrwGr6+uKlChWt+dmmKSjG7NCetP9IJChfQBWRL5GDNFlQGP8TXrJGxp3TODrAX
HMJ+yrAfXFxq00YBQVuHLghki2dEPuipYq+CwiPNTmJo8pWUEIO1KhMZe85AE/D4
3hMg4930GU/f8JFbzqF1ZEyPuTjqHGkuExmHjQLWskq0sNcctbKWtCAYH/ATDocD
/WhYKvUkWEqL7GM4nWbEtVKuRhrFwblujkh+dewY7OyHOwRNIp+A5d+8bl9kfx59
aHWZc2sRd8Zegn5Yx37Nqw07tv8kod2LmGEAv16dhGzJeP0THMwK2fjJ2XZ3z3JT
Tnf0Qg/U0zUdO65/BCArzYkzKmUlyCwt2zSvn5nRh8i82qV8DJ7jc4ZgSHY4H/Dg
GHBKiZawkiL6qWvZ3J7C75iBU36EXwFMbdX0iIHoXyBQmMi3ZIcK/B6/p/2JYppe
dTDxjRL2HrvUV89JlqeesOwakYhSeb0TjXMs3QWIgFz32QjjMr2Mqqx0rgi0AswH
J4Lg4y2ISS54JKemxhYvQ9LSXDr46hR0Jtka/Uj7s3qlePTpXd65M28EDmPeCR9Q
5TF28EOU1mKS+RvHt8x2u7C7o2EKpbmq6V7aME6PEKUvm0yFbTolF0nneWmun8JH
FIXrBg7R9jVV2aul3jMjSk7lak5wAX8aijVAeUgwoPYSBwsqxRbe0SGItBkCi28v
vtpT22ZSbZ/7tYFR0j6AzGQDFJYvje/hbqq/svXHPXYquH1Xu7+PnfDGeuELRc34
vf5H34eu149L5OI0WNqQZZAH/kcYBrYtgyIfTgxWtjY/0wUBlM1nbnJlGc2SmSpQ
lDXLGQjILvl9pPbyK+FtW3fjPhlLs3n9tuiT09uD8NmvkVz8QqyxTwyErXmTS7nO
C/oV87FNGgknkmRLB66WMmaGdSSxg/v0qQzEMl7XXepJW8zMWZDfLUnmZWmuI/Q6
jbuv7UfoGQ0wn0Uou6yMBb+fkSchviTk/aQcnUH2qXof5VUA+OsMye5wJ0pMeIZg
t2gIbDByavCjv6y6Jv8riPBNM+o1yN3HyNk0FHAEe6KSlhhp+39rjyvohuW8wiaY
g0O8v0QA6enhWAEawEjdWm9vXhBPCK6db/XBVvdjvqCudkPMQyOQ2I9qZv3uqo2n
IPJR9rhSWEWPTX4aHmuB54B0LXvhVBPsiHHQInfIDcRpOdvxsZlU9AI6ORYHf2dS
lVEZtit//oPwRJBMREntodIw1pSteM/akeLeguggROwuQtAyvMb+00/5duPMRyFU
tebrb0qKsTb8NQdvs6DmmbW3YdMxwVxfJgJnEqD3+P6zGcu3cPjEwDaNf2xv3so2
j2pmDnsfIUhIVxJz8OQoc472hE8aTIej4MkqHY2jsWVv7SKf7CM2rNhgWsjBNx1d
qYG48IWkxtOAMaQf5dL6U36ymsYLuRqCA7DacYk6xn8iAFb96GcUdxnq0+lxtB5r
V/C2Pn49n/1e2nAsNxx6FvNZqlNZPpWNXmbEz9gNgCD+2wA9Y8YdBA5s0zFeS4a3
eVwg4C8lbqxfElS++cbUP7DOS1SWM/RHqQ1FfseEqDwMmwEh2LzS5IFkVZeCDbiQ
Mb5mk5SQ6FVaFFNErFxEt4GqtkvrNOVZRZ3PQ5hPrbxtOi+sO9NuEldMfrMMda9i
920QjoGXxFjttXwz3UcyedrIeFxvMXCPiZtsVoTBEAlgA9CQExSR9h7vt3CjPKGZ
ziMzDXkd++45+saYjfRVeqavl6axfL5tMZGWLP09KQMlaIgJjnIL4yu4IeAL1p0I
9HU9A+iLC5Dk2fqdjU3BeQnkBOj9OVZSOmBATeMAbRXEysOGvOVISCVve77GUoGZ
he/bCWUopFTwZj3joCukIVZZQVd+Xw9BZaZ4I5gPwBswkup1Xa9jCJBlz9kqqyS8
5Eggn7z1xOkiedAoTII0pl3Q3kcGXSKu1Be2X1HAI7Wx8FI1pG0aDyrTCYDjfGKF
Z+KxvI1yjhfCCYoeGWvBLIKJRFrnapsAe4A2zE9DzGwQicyjDFxQgjz4Jeql4jja
O+hM+XE0e8TRXcG6JqL3pyAnoU0B4lN/D70dMptbRk9QYK9/ux6LQBdFNy7uxsv3
WwnBmGlWCFzYjk0PuATVdtuA4TZ7KRf5G6OI4a9+VYQ7mDl26Iy2NuaMk5sUlKnM
YSxvPo301cbssG4B1Ge9h1igeWuMH1ddtjBnT4EBKAxE2ImzJYUSye+1QDL5DEIF
iRskg50u4U0rnoEXoYpIIR39EJMAR37fdOzep3ORlI3ut5v/TIS0SadcYlNDopMw
L24nDQwe+tKzehipsacq7D/CkOYN+bsUsvx/7hcHcYIGOMw1pheGAUUZ8Y333iPH
QhqdMQ371SdB+0wS5Kzuoh2boh+xw8odgPhFhq+y27YLo6KfiuklG+Cpc5dVc5yg
y/H0RMELathZqSRDZTwdHEiBLCHNvBOnxdtPqEu/n5p3QhWJT7/ow+OOkvJVuRJO
Nw8xL5u1LsZP3kdKzUYO+SgyCOvwuR1ClfbxRI/PF8WHcmHJshemJbvu3CJfSkcD
FG46lQEjI/Y1fVUby40chPoUWKJu8Zu9l+WhPDFNry7pb/ly4dlobAvAB5qYj9qT
RgCkJmccr1+97I6XS1CuxS7QJIIGAEXlHAXBI3U13omJ8UWA8KCteWs8MLUG/8hQ
MV3Fk5Aszf6HJ1jj6YlaWDfMLhEyqyMhhS6GArSLty57WMOrl63Yh4UYM1FvnBXP
KDVxlOMgeRql+6ldvxoDfUa1XnR0lA0il4/U1bry6E3gB8bkRs6xIVZ/2NrZnBKU
5RE2fhb/sBBUK6CAXH4BSt7gZnwdTt9yhvlCEaFeCuaCLEmMEjoV+jhetNXZtMd4
HTUK+gRqni/CtLVhb0k5ZfQj22JcYjIqCulxd9svh+V4XMDjg6LVpb6x8VXZiobn
RfuImQ6/VWN2uKSjKFRoYTpXsoXtxIVzuppKWc/n+4VqWkSo8IfmujTIVvkn4jIk
rqZdyWP/9ewnz6f21cbzlCCDcOsy3+QdC4lNVaDldfFtdqsVnW7xEdX2ClqjHfyr
UYue6I7d9X9DYMCbSXfrmPIgsJbL5qNPGnM9vtZi4ab39rf+HXyjSR5CgbkVebTU
ergcGs/PqcTDcJtauwvNC8BzCrVcOSMzBY1Q7cuqND2ngZNvCG7PcCTYYLaYLQOL
E6ZA1/OmW4eVbKcuN3tFQqTY6c6YxUuZ65K7j47c+MNuXleZLaCyflEwYGO23B29
CVjYcRu7sYvL5dtUxhrcnpPQOeMDlaTiw0p0fgMY+fYANTfJYE+LDnDgK4XgIMSv
lglu9foi9mT0RWLuEWUC1SKMmuJNnTQJljDP8JnziqTXwlLLiAcmj7TBQMScfK+n
NAVLsH0E7aWenUNTTuiM+T8geaVGJePa/Kig9jGHi8PTH3mlYq/4quH3K+giFv29
wKLV2XYgiR86lkSGIpTdu6imWokontEviZH6jXu15FLP8pQzDH/7yMykhEYdhKHh
8C5a8dwQyoAuF9WSBucxYmeO9J+jodjjjgsWicKaBMVARpoSlxyQ7cJ0XPEhIWEt
rnxsJ4cHItk7bSsdjTFlzG/JeZTWXN162D6PG3TIYZ81gjYQvBRS13X7UmmvjbFW
gIng1C6eVoG50yS9lgOHSdLtvXW4ZUYrNVdOmb/ZntxVjM+Mymdh199bkW5thoX/
VODA+RTssQFxdUyy84TSe8FFryzwgsXx5EaOF4RF2jl0DW4qxq4K8i1kHPNgYVnU
w3rzgVi5wUuGIWcHIpGolKeQ9ahc1iwsJxPFjhW68VOFEbfkKh6psT/i4ygTms2y
D7eH/QuUnETNe2W8TRLL7zGQb+5TlecvNHEVP1UMMNMlSpWV12SI6m6JC4i2RwlW
pb/yPqn9gQgvFHoZZWg/i1+70AL1EV3FgTBhz9YXOxoX/HN0oUyMB/QjwkF7povs
wTaRufip454HZhV/SDqK7o093ho8bRYacbWAYzuXxMshm6IvFpwjTOzbpO+nxzbO
N9qsOCU7uzHYtJ4adBDZPHH0emx22FDuZVNqOUBj2AVnZXBczDlSbSag7VZuOsL3
yVsRrq+vcOfmZ/EKi9ltiaKkxlC2UHcgsgeCfDIWn+iC8P8q8I8blV6UDzIuvMvH
zvuNiYyo4JEb1hJpIJN7kmDZdib7DdWgnkc2ClGctclgIgj266OEV0G+o6+597PK
1fD7SXRxmW73rnFD+mhntzfZzsrg2RuV0w7sAhu6/sBmLV04KM7OEJ9++Elx+9rm
PD6Q31cVYB8P7hCn03RtJHPDmAlP8xRYCtmuqzF1LXsqsoQmv21IpbRQNboZ4pMp
uE2nRfZv02i+1d5dPaBXLLYncjAWFM/ioL5HHOVuKZIZyIFt1Rj9Assi/9xnJbDy
buDc7xjW/ShWZcMV1mCPyoiCDLgYaUVmXpXRYiNqfzD0o7Gc1awX4Rj52eddABTw
AnFSUam5EpvVZ/0CKveBGol2GcfJ61vcLaSGBgPrsGZ9pP6ILhQXF6Jw/Tm50PyU
mkuze6qC3BJXXkisb4ULGDH1I54xf7D6YGkjIhya4WsqlC2ogmpJ3ZXKZWeBbFpA
/ArbmdgMolkF6Drz2SA7S78VJOasNhLU93DzvDBaVUlFCnWEHCa294GuowfKAPfA
o3FYOPl5Txq4McWmJFebOaRN2LEKpAtgzm/FWn/GGEVHz/2tnLCHIrugcpV0HjbX
AG4xEEuVdqYT0i8LZ86qIXDpJM7oKJMOhD6VwM+bxUVsvpmNDTpGKCC1nxAayyAw
xiQbZAKIHEA9D+WA+1+spxBvT5Mu7YurJH/KN5xIK+8wlP5NJNMX7OFJ68NSpMC/
6csejTpNwzVXZLBaG4pa1FsywxXSHMyX4JFgIUgs7n/FBFVf430BqsWgCUNNw6tb
V19AJLA3vuNRqnORXE4vbI9l0Nskk5+DjuIyHtt5owLQufi9zuUDvc6UNxmp1Sqg
amRRuBAOqNQRKUCGYkWahiu015diapPoDmIQXX44VGwYbZZCl4q+kr/nVQSzUa/G
XNwCY8jsxgCmSuzsgrR15n/Att8CfbwPcsmiPToAEB6tu2WBD7W4SkmVgWlzJQY+
lUg9rh+2fnChqg77HSK4thElEoFjM7kA2eXvPwyp92qitCacGY1o0eso5duHUq17
jRtLN6N4A44cCvku9oyT4jZT+/k6QdQtYp1dXoi+VtLLkZXe/Hibr7OVjh/XhPeA
uQPeh5cvu/1s4bbTheUyr7M/KyBMbAAYhgWFMwhNgOkkYjKBez4glDId0bHO4i7u
4iGVbOdbSKrmRndHXPoQT+ZMuEIIIVCnkSF/MpTsIwtrNy5tFDcGW11qowy8ppXp
G4LvsXKymHKSfPSoetOtoic3BZmChck1rg/Ju4vsMLFoT2b+nYGz6/I+VE7PgxFV
fjB5FcsTztAwdD/i+Y8VisFCf5voE4whWJ9LrCZfBt5UN/HSpUtoKFRfxdga8f7r
5PHBp0JVukA+r2IThyWMSKpMS1xEb/neNHY+7pa754eHvsYfigz5SMT+iUn2L1Fp
4slbG3d1YAzdDeLLuCjpJvNaRmjULWAjIQlGotavcbAzUKQB6iZRDV2G8vRNqV4T
l58D6VSnUywHWhydUDCg2CcJuXpTDNNU2tHSUIJskjWeovF5saNzqcwGTuMdcPAN
BjuZhWvRQhbIo6GX2EJhWHMoTztxrtVCy9fG4zOvzDo/h6RJPYKk6DIUkaRwHxFM
36AAB6o+T3mrf5DzuZ+nVqfSZPllWpE6iEPu3ktB/NdAk1ml292nMksp1miBcb6J
A/EcxerGB8yWB+iIpoKdda8ntVrO1YPRZ0V2xrYlUPxgPYaOb8ZMqgkUnTYsCFOU
5QIJ++ziZkW6HZGv3DP8Dv39zEddvBfHNZx88ZiW4jLxMLzJC26Krb39WqG2HAdy
dcKAOYtAOoLzFd/VWg0BIXGL1tNc+Sk0hTQsTDVi712uGDNr6+RE5j4WBgitaSQ8
nHl4RIuV0lPrgSno8snB5iEVLRfStwyGhKGRneUwMs+as19bSsccOteEr9Gzis0d
SY8YbGfa788oFKbvvAVrkdocqj3AhNMdcOvjoyEUizazyi8LvNK0yVBpd57blm1m
bQ7SkutJXYl2zNPWez3fGIsg8bt7gQxSxy4+17zjJe+sDcf4u2vdKO1fp1/Ajmhj
2H3ZG6pJnS/Xq+a2J7XE+AzG5UPZlNi2TyFbVMeNhkiM/XkAk5CaDWcKDENGcmU8
CW2KjxmzRBgSFEp9BediaZTbGfvYMretfaPRXHro13ccyJvQNzgoheI2ingW/TFV
ZdRPjf9AiYrkwzTykTilNGtHf7XS12LUKXuG3e1R0XH/N2VdpVmjP9eYEQaTYOcp
ZQqJrDEl4PPJw/FuF3gftnKP+6vh/iLXrEWRiIMWjNzlJzNRqRczeMB4HD/eUvo6
cuC2uAiqHRZrr3PiEWD6B1BK7q/HdtHSZrPXU4A8icBfpQ7G8TxmTpRZ5XY7uQNN
3s55xBC57Ssgh1VGPOVIjH0xj/o18n8LFDc/hJr+s1vYjzW/XupP7uo3V4d/A8oW
48eRJpTYtVM6vwPnm3OF9yh0ecXLGhIS2jw+nLeLEPY9AagG8sdTrkppED7AEwEo
ui9+IWZFbpf6eea2arATMAoMIRUCABwuMN6UaYK1je8Q/8b+HusVb+vpvl8+7uda
015ofSwn0NkLyNsrKGaXxbb8f71MjaOBxLSi24NbhhgJO7+0uhzNj5Mm0tYDJiJY
72Z0ykJrrKtj3o4MmRJNIq9joerRgW9U44QtpcAFgmy/j0UFS3wgunoZCRG4y9qW
6ZFwr6P6Pr7WP5QavIYwbClsMZXCPr1TVPVcgydYgXYk0FZp4CSEJY0JG/E4khoQ
NORmtRAuDKPBDxi0NwGF7pmu8JcHM401fAMQVmisNgV4TXefywFXErJfqyyjawKF
UsOB2cd7zlBCAATyQbvqV0ej0FSLfoJfLHAyH/Ok0WjJRR3J52S6uAbQ8t7cwNlr
V9wEJV7LIdeRwjbMVzTd6SqHSGZyNYGjrZUTh6u9SEZvvm8LXctWG++H2oXJQNWG
XTWjtfLWKSYzKWDnIorAXOUDyf4XaZnyUkrBExpvVojct5UInpQzFMbjeYWo5mbT
8zVHaYrR039nh6kIlin7Zwo9i74ELRe8TPGbAsrBdKZUXKhca8NFqe2tB84Y0rL5
JKbQrhPeA5CwAOH6dxLpY0jTITufMLHgIaddfwkxGjFSn7BhhbzN0c28doJzsRmt
oiYq9obsdgawvoN1LkODZA2xXE5p3eNRUGHZgQCM0dBFp9grmVE0/Y/DOUmTjpqr
PuQDqBwL261h4w+unZZ+DB8RbdcbXSmCI1ingCRwHcWHn1wL+YtAKACDqsypk0vO
R8Q+i3tK3LgKr+lEznLTadKtDFzk6M1VOvRIyDlkFlpG+uhfR06dOSDIq80mpIT3
ay/nTnJGsBQg/2osiJMOarjGB/zID5gJbQ7cvKNDismbmb9NhHy5FETJqytlPiQI
WYCivXwWB5yeO8kwK3lSMPpFzPdP114oC9xvffAsmuELatuDmV9SM9bC17+tF9rH
q2drlSMqjjmU1fHS9tlPZsr8TenB4W9u3Sd5pfMSXtJxhCVpK5k/mwP5kvRA5Fra
Mu4Wc/+wWoCOyCYlhylYerRRvtVaHiCMIsvzDFcZ56TvdL9ufnmqN6fLzMNM7L21
ztI8Xj3dGKDlXUhsQGDZVw0BTLN+A9RvzQJI48/nzhPWy6/U/nLuPR2GJG6B8a01
lyMtVleLp323k5qdijRgaMwUo/Zn3TLBwTFl43MI4gf2j54DpL2khlzuzijX3WHR
6m88iWxIr5CZnoFFr1pDHzN9yFJVToQRZ917tQG24n1hmt2VbrJedr92VGuWC+Sp
Eha2epK1MpAmb8TK9IccqJAPjusxMgUwsTIPrS6F3myDSAseF+pfLG7dTGeV3+tq
3xSUjArkhsruDUVMxGREnhznoxZkYE3OaWA9Cn7dcwVjbfqr/pgWehEN6jDZlGMz
EAvZsJ+y3ECt6Y/0azp9fT7bvYrZbiJlEEd8hb0nHKaLUZr+RMhLeFxkRNatUlHy
wO//F2HP3as4xwBzFHUEBrEPD/pyNtSiXhcW8o2QqAEn9bY6fS13GSAQITWTfu5r
y/u6oP/ozHib7iVC6MLu/ZSsn0m8N8Tg6enBISw0kyNnidt21AERXsxFYKsTVMOC
+RzQLLGGaKWX0fSdxoN+SFdLSMVZxHtSNkzaX2th5bhtsqkYE5zXLa8j3OgRDByE
sfA+7/hrQZTwm6EGRT+Q+IgyaO2vNio3SjhKZsiDmifeTEOxyBOiWTY/VIPlAOvJ
Hx3XeZ4yReNM6c1zq8yExeKg4eFdekV+X8seLc8yfgg1WiXqadbuKWOG06nKZ4pM
6a/PQ3Y+M25/S+8gg1iPuO8BIfvDa3GAg2VLpLRzCYVdhyqkgcew0AdKNbtXoQip
PFfFYhXqvuRS5slOZpUJQ6rnFQNUBim7sACDmIgEWPH0+dKkI/hX+hp1UUGghinv
3n68N3jGnPsHyzKC+PoppJR5rnjJZZ726wMds5tb7jkb4YLEmJJIOLRyXKX41u9A
UHzsqQs5Dha+7YsrUvMiNdp3KxZSgbfuJ4r9TlfKwqztLmodgqjGEgCH1RiNpnsx
N7EeRRskpu1Or2CFVZIygo+k8f0IsJRzgDCE+EKqYTyUjkNhf9juC9jqU5BIm70S
DJSVr+W4uZFJ0swvlks0SZVPr35ApSMS39LjTd6VUXdhP5ggT35i1OT/QIi2sqRG
NAE4oTjW/Kdu6OPknuVj0TWeklebw1xbsnMO60fot3PeBC61/VnJ9D9ZQsXxtmzt
ABAKxXnZ0bHdjJlA8jhxYbuih99wFbv0Hetm++Zi5RPbDpFVDa96Onad/TC3m+x1
E4KiRTjdHi4vttKAbeJZX8Jq2MTIFxoVFrOVOzEbsb6WEzEhA/pb8IJcqVv/CNpt
EFh5GcxTtCnIOGaHbWK/MBCFP2gMaX5Kj0AQ7sSmvtTOETRO357uJB/qMnDRsaC6
db3YIy0PPP9NcAvNYqylxKRVZ5WG22hw8QPqFVqo0RQ4fCaMlEL83i0chhUXGcjS
xnnLJ/0QkpISPAsPz6ahZXM4pTKvFSP22kQ1+I0gVtopGSBUbw+r4FY+KQBFBMch
YmO72WqarmsS4Xdqg8RO4zyVWjNSt+OcKO3eVrB1njvt0TZkIb8+CGB1rV/ELFdJ
P30WynFF1prfFV3p25MTBL0cl/qzjZoqcrTZqHYoqxWUZtXZ1VoVnTV0nRToiU1T
WLwMC10Q4yq8J4ZKyL0Afx5rBQDblbqtcyi03TiebSchUf/Pe03eUwGJnHot4gjN
MV1Tapr0d5Y3OVpuEPIC7HJ2mREa6OfmlLD6+YxxD+IT9Vyldnuprv4m1lh6Qv27
S9KCVZP09R4+a3AYIxLJObwuHqA7bCpcHkeqGFHA0AOk0B4fCiUDvJHzMOrocL+s
pJ6anJhdQSL6aIPnzi1WIOyZUhoVbE5BGsmiAtqw+khuyjd/6zV+C5fSNzxubSaG
hbYpzACyfdCNbUJEWNv4ST4avXddpP9RhwfgXQZ5nDKQh+E5LhpYAT3vHoIjRJAL
D1OILRP+YBFZfrcmjSbGYJcDd40EQlhqRmBRm6t+fZi/dksrY6rLyM4VS9+GewOc
a1gjvl/2SDNsj5W+Btcpaiw4ACf0IFattmsuIrX+Y8v4uXRvNbXomjC8Fad+mslR
PFaXf2YgIOZZoQQwRGz3OIcH3AN7eI/fJ5PS44p0YVJUUFZPhGBf6ulJOAbixrO5
WJqIGOldWi9oLYT+Ad7RdOguBMUllFhDBHaYUMBvwaxeL/RDXB+dnc5//UQOf83j
e5u5uPo8UePRs/qeUlKs2L3ZOrhBDa0Z/zsdXsFdvRMVr4cX7ZlVWIqODF1JNwjD
i8ymk1hjZTHHYXkAubGiULMs6W27d1HEJl2cyUQau5wn3ssqAIAwOeAhBANaTJDZ
ItUOh1YXjrDdhnZdcGZ22vTosvLYprItFnNhEYbkmcPpuTTd2u+nTXdz+81Q4raz
xCpjt2qhRKRwB1g8Jx/DDo+km/OJ9THKibYUr2YGSerBSQkmRrpATpzUA95BSFsZ
crQmqVyKA7NoPmJB/GuhIUV+SRpBfzfnW8EVbuTOQgbqjM2u7GLb37OFVAXb1zSV
BkumsMxzLVqL4IHkHRsCY0r0VZfeKmyik2j0XNAvObDUJc3iNiHrh2Y3Cjv+eldP
GhzQhRP3n3egz3GP4KKlUfhjBIhksZosCdIfd/HYltG76re/3dKAobHcyuWJS/55
TzBD4YaYHu8a+uwEWTRbYFz5J/cszRgM8b3yoMT/l9JVAIxfEUNjB8tYpQMy3jhM
YCridhQoOcgRnvHwq7DPW6Lf4h17eKzPajBOKeMmS9R9TzZ76sFejnIN6XVF2qS5
oZ9q8l0oSjeKpoj+uY/AWDdBgsLdbmVHRVo5oLiyXlJWB028z/W7foF89I5gHMNh
9E/a6mn1cenzC7IDAb/wMLWQpQSCMo7edX7FmP2J64OrWCUIHq13Pt489FdlOmP/
k6bfSgcMsovTIEcoPKdOOdtvRsul3zeXlUVQ74WnYG2gIWKPTpBGASkR9TJm6CTi
aQrS6F0nsyPYJQCBK3NYvY20464nX9tbDypOJeTfz3ktgo8GseMl0Tm2Ft5jR5TH
H1qZKNgXtFJSmeufYV/KZs527BvsvY20kc5huh5EifnYHc49eYc3NXpEe89nbhrz
nFYs/BkviguZOyWelf+IO5hNKTF/gB7fGCxyo11Nrl96CwkSrCIAUWLWcEkqHC0q
P17lM9WqkJeuhE7cgInsOom8H/6V+C+xaO8V56m0ZJrFOh9hWXqa3bFZu9w/cg8a
zXOSaGEOOGvwGQ7NLP1DP66IIKONTgSNsMH0dSPO/v/giYC1a/lZe4b3g60JoxFE
uF9ejFrrucL0YB8PZfECz+ZCdKpRxm+DvLZTMYmscG39jZnDIU64rdXPg4wv0NDW
rlQHzqSJpi1pJ/0H8x2H7F5uAq6qRT+yR80Nos5zZc3O4p3a2OKvDbivXMBrwTCV
9zWDAJOyFBTFWlZf0X5iIJ37+ajFzeufM1XTn0+yhe9jXV4XT7AWKuQ4wHwN3qd3
0liMTB6ac2gOjLOgimCV9z8bZm0EOpHdweLhzQS8J07xUWtrItX1FXOTpcdo7ezP
Et15DsVPAX9d5nvFWxyrFuUAq6h+hLCHKozwGa0zBOiE50fGVIxzFswmr98DNwzR
o/1YyZxBljcQm4ChrZ+GU/+Kf4DQ2wKXVVC7pHDOXJfWxU3QSI3SReDlVOptnPwe
/wLQBK4IwKtwO1gqWut4g/XI0i/PXMX8ZOVm0PUKP5ej7J1yQF4SG3HM12payL6L
iovBmI5vMsCTUhmHZYR+JzKLD7Qq+9ELk0veSd7E2GVxBWibJC5W4WMYtIVCi6RH
H1w1405sGJdizbUVUBwBAiERPsb9eWuePpIepAq3CRKrHUXp93Otkc6UUU6iBo3D
3oZzrvlo88ng8NVvfffFpZVojcmJ8NdrlXNeKhha5htdrtxHDt+RVFIrCERoRZdX
4f9oRHFNA2esL6vrbGzdQhJ1p/QqdbvzjnGMoNi8snibjbwzNB7Qqj9FJaHhY4vn
Bce8JbjG+UlmGGYQ5YMf4cQIoCsaSef9/5brBq7lTrg+UDL6lwkHETMFJ0/eIGld
3KfGkDMOL+6wxciWjHeZEgclPlrC6fj9KOGz/D8VOuwXb7sbMQZ8pFXVDOjnfb/m
GaJrvEOrsKyCiAMetZLOSxH7xa410sFWBvKjDgOTVoL9lOSu1Yz0r9wF+35ohAVt
zYu2zGdQ2YtxgcvA2ISXU1dbtO/Uc24Htbk2SUnJfT41MiYws655S10WR/pTpTV7
dYcHcu+mJjcQrC5OlVwQho0sYNHY0hE/b4RP1J/Z8ThjKdXK79wcHeroB/UmgaUZ
6NNtN2H0LupDJTN7wz40hroS4QFL3S88UvBphA7vwdDsfhVfVHIe06Omf1PZ8Cud
ihQeCqcSrph5I8UFzqwiGD6EQWY1Cw4NeNjoabq8srpGs342IB+Hj3JiW1roEEf+
Yw9FxO8QirJUDjHAmzfybeNzjhpTKDHIzuXGLkd4Zv8w79LpdzwaLe8T2dN7LbHa
CeNd3aAuf3RMO1A/z7njIEfqhSdAHUP8hZvjg/G7IwrDTZuP29ikkZikEy70hmXI
4FWVjS16TEKuNHDL94yYQDSbUviQGj0vrIE3xzoAeTvg0tQg6HSZtrF9thGSIack
3I6ZRtuuS/CeP1wPBZkkf63HvDGiyQfVOzS5xUXlmmnuijs92vpxvm1wkgvrWWMV
w6vibAx/IJosXldaatFcgbjBn00C1E6JfAmG2jOrc3ki0z+3TQatEKTmw5bUWbtx
S/9ELuUmVQQ/upYOV832LZ9v7pwW6y1ddHkUiUGR6ubJwHKjlcVwm/29/LLsx0B9
16V8Ig6neGNd1JWTYpG0g3fc18N6hy0pqJDaFS0QHvK/hXP5GKXhl+RRDpswfmON
5nx4ccf4uDn9Vjiwr317L7alstJK8ZOw5i32PZYAUSL0SEO4vYk/8bxJW0t6GJ+Q
7kUtmuxFRwX5hKPI+w+LsdcKm7jQyyCql9MC+OKQ0gblz6mjvXft/8OAzQlTpeu2
0OxTcvDcQAAX3Z4kpFt9Sxu8buQpy24gMsNzrnO2p/38f3iNbTxM8YvyzSMqT/2V
XSJYAn3Gaq4L4SUV0mFzqN/C3T31+R47cPTm0Kfty8iJZART7qzO2G6jkZOou3C2
tFGyY81n4qNnIGaz0HSxxLqcyr2nkQKdWI1z9h8WyBiLlcCJoLq60kY4EEZoBoHw
MsJTii/ITmWFVpSGR/i7Df7HGViJ7KUxwkpDpBGQLgjUUsY4O+IU+hb6svPoUWXJ
wVhOPwjWYGZfTAEOQv1Khx/WyKqscbB60HE5LNa4EzW2nmvLu/+WV0F2UeU2RZSp
Hgk20O/Of428mK970mlx9Utdn4ut5mAholcLQ4Oy0ELeqMc07wwzdJGrnYYoNvsA
jEeIUVZPjSPf1bVHVSXYDtqanxqJpwRTMgm9cR2CIYvpRkJUsa3eSd2SNEgEWyzF
Y3sEnC8NN7nQgYmVwynGKGdRYbTLly14UgRrlhdp6GQvarjdn0jE0UbJr8NzR/4l
QvmR6OWToPUMu+KdRVVDLj+YkQ/YGXbL27ymhJbCNuyXadmQPRrH1Oe7o3M8f7Zk
hYU32KE++WtabPcmCu8Vt1aC8IIRj5vdWd5HseWGZ0oRxdgGmHT6Zm4lyynwXao1
NZScg/YYQiO1kLqqqjIX82/yFxsorVTOktih7o+2tD3ovGeOXh8pRPFvIC0WccW4
tBUF73YZvKSqAP0zrEAGUOfml6X8zaztsZU6tAFXReBYHHEBvphGcm5/9gBV0VcJ
GdUqY3v6xT5MR0cWDFUVJGkGy7Hz7ZeLoBbSyu74FyMC+eORBZnLo02Tv0jlkUmg
VvJzToXpGms2ffLjJbf3moOsD+yxZzJxmQ5N3MhjbciJymdBFz81kooGSghs+e+W
rdCx3sU47moyx+EZ0F9wahLL5qGpF4g33wG7Mk/9HpNukLSfeRPX7rQM+2ooBK9O
zRevT0pThEn28XklTgN57E8K50a1DWAsVx2sOOUpyL8EDXycdIXOIpKU52CwyBGa
zwpSXoeBa6SvewdGTm5cnZemYVkjuIc/nApJ71xNhCSWqSQNsN6eZ2arMVMIvoo6
B4ByPpIFLvMazfxT+df6dCZKi86qZ6xDhn0IbGY7QzwSZtMkbHPDt68+fzFWwZ4L
PN3K4Nv7zDhxsLTWsK4RQsiYACqrLpdj6P/wDKpn4XIv6OXsJvnKNbNBGlTcvFQS
+cQSXOGD8U4jG527pGi8mEmJpurKlbk4f98flON8fPibPpUW5D8pBUPGbbY7/IQK
u7C+7hrwKHikFhnahPBxujsSHUw89Y5jmMtJyCTj73d/oTEU4WUj04vFlcAXI5r7
8GSHrkeNNah977pn0CLU6O8L2GzhbLKfeYYsoA3hQCKAUyNeVVniCIYsbeooXsdC
uNs3ftuyXSaqNdzaEORK+iguO9cBX13JdgANY7kFWbohgbUWarn8CTPxFWb9cgwT
XpdZy4jUS2ei3MAwS+RAcyrafNQY/wdhiZy7eLMbwRVDTqqv34JligBolSBYWzjc
tzvUhk6OXMinvmEd8Eyo4rvaLxdqG3KoKh/DIZlrtGCxukwfPbtOnZR7MFmO1IhK
JDFcDVCk9WtiIQGG+++Lx5ZlecuIz3cjKs3pS1a7y2agdILO/FJX5sReMQ/8ByVO
VWNEFp5DYZL+UyOseyrTcTwt6pvp693zlQOjKR1pzKgCmNP2MojJDWFHwhrD1fkr
Gj52GI+WYg8s+yzyNGi3foUIvuiWYIPf4ks956kcoozuG96oQ6y3GftxFX7cyiW6
djiLOjJhPqUi7XBNZPvTcGonZJgeES/8bkxTUYT6YagbbqaKzJayaIA51BnzrCsV
NNifM2s4oUDbiZsgmJ6By/gHuWBFFiufrXccwowGVNuTMmnvdQgPcuoIHdXEIzbU
15Jce61gArcKttFETVhmiW/8hiJbr54Bm469mr1xKsqogWROhXBnqeYZxSGF4rna
OD9rFbSjcroNVSo/NriuDVA0Pj1jFMz4c+J1eVkIbAKaCLMhnRRgQxZchA62YWMM
79UvS7IpV8frc9fx+KDB3jkJq656QvdH/pmXh8vskDe3hW1NhQKdjHxsaICbiVAz
Ir36lSSqtTalheEJ9fPN9ypsMVvhZIQahCHFus0SJBQnAxWFOksCQFRR1xkSTeM9
DN9kIVQEWHYKisHh6zGclRrsu9zb2V46xISlZEG4fJXc2jvCb3WtgxZfNj/lDnpM
+Bg8+itQ+ACO98yovQrT9V2DAjKB7p3eUKrLQTvfWw9JprJwrtZYMxnhtUIwbQLX
wqq0hb7CAuz7espwsMkzcow9JAKaUZJc1l0FTZc+/3+sGO7mf8T708Z9b2GbkP9O
+2GJrr88+B4xDqEeQE3lMdNyl7ylIGg0aGtRIr4rTeU/qodGg3/0MlgbIdIC14PC
hSR4TufuvZaZU9h6k9CvY6vF8rNjtlDyEkVEEsVfLv7nYmHo7MwYxGYj9wvYG9kB
52ZIScvdr86UBGVC83umHzsaYhMs/g20GESrezLM8tC6dPXJNdxdZKPxY3cu6++r
670L44tvqqAtpT0ITZmcq+imnmdZrlVWaxbfxB8aNdTjmx+zIcaujRB68D+drBIc
i4sGTssX+fkckU/qyrZghkpoGP5uAbU/hAWkm7ItmqpWqbv8Wa3aRkau+2AVW0/X
OefweejLk9b8ekcFPoK6KMekeSUQSv06/OrXPXJ85przskXKUmHC8rxY852Nw7TP
FuOhyFkVenZbpys3XtalgX6ElVmdQEk2go1WyXvK3NElEXgzCK0WBQsf2t46Bub7
XfKh0/u3IF/7b2YsefUn4yA0H2DG3DsaOyQvsVtvcjSB2HSdiBo8QGiaav3DtIT/
rXC8Q5iZGENRQaRlQbRN9ZzMYjBKPii2rfCi/9j9PIBkDJz6TlxaAg8XPn8Fon85
I0EQY9bSEwnambmnYULNKX71vzWNTVPJU6+FZTsMjBbP6y9PDz/wSJ9Cp2c1V0OP
hDKCIaCeZdFsZ3nIqJbYgizdJ2h71yVDwXC9AGEpO+bv+g9CUaV6XBAKXUCwVvs8
zP1V/QzR3ph045RDzuK8/TVSViBUWrQAmcMTgNJlXBcxkJ1Pt0v/WBSvqt+xxWSz
SKye6vGDUMMAIcOek0bs/g3KueM3GMUSHYFu6MizkZf9A/JuxjbcN/tVBbYvWqgE
VS6GWoJiAw2CqAeKJsQgesvKCBhlkbErJj8e2AtzOG69862sYvNCvNmmAv1I0xEy
lwhVlDpY1KsdfmrE+yTdhX0M98lh6inoSaX/5hClQDsRa5xGsFFLHXCmmSCrxoq7
uTUaoiHcKeUtunOCmAcbJRXKcFfVSM9O7j814Ng0BMvZZDcbwI/cxjsz7zq/Kyvi
E1bUA6S3xxiZE+i1E0lCec/IkmngZizTfjq8vsSeuCVhv3jbtCaspBOBkdx5nWIP
YZjydGZ1DaQ6ay++++CBkq4AInKx1MEgPH9k4IVMKL+FJ6qmRZxG4iW4tS3RvZ43
VPAumILGtgFONeWLgl+3sGMhoUjbRfXzJXsA8ytK7/WPMe5FTkl8o6fxqhec/Rk2
/OA/8CbKcLTelUVcFalFlJoopd7ZNcB1lKT7xIif4sH7ofr5ZXnDbU1mcFVANhgV
2brywglngxxy4JCGdEytMQtubSRfbUjdLf0GGok0VhlurCwdQGnFkuXPeo7YRR4r
n0a3KslHnDAE/FOQq20lIr7v+rtvJCOIb78nWZlnYhBVDNLz7m0Kof/lI4evbym+
oNc4qGs0n+LqQ3uGdRYbXsd43z7GeDjMbTZkJoqQHK3FFUeH4zpeMwICftTVgAWk
Pv9YdVLq6tjr8/FOzUlWcOpdXX7JJ4ac45/I+7eltcihpVLAgROBuM0fLb6sRi+i
Ee1Iuiy9ZVpXmisacQARtebwRtQBQX5UDgimU/mneZolga/zmasoyxNGSyFv7rP5
o5EbkMUKet0PdrHmj0e5QqA3OWOiVKbC+WYUTh2TBf3c3xlRmO+IQSXpKXpm88Ux
/MeybsEec+v2cpMIWDaCRW7FNoZGhcsuRZLXR6Fv7mxPWQtJNeupmD7w2GBwaZiW
UU8mY05A3berGX46lNhJ9eHi9FVhfotzHLCW1Fh+DbEzZslFNiUbrC+eFAqWfjlv
xkeIlBfcPaczwowYZffxYCGUeKuC2K28722slozLS/vm397ubUPX6dZIgtC88hGo
NKQAUlum0bQSdofLkBWfWNVadnPAKfvMvltceoNGMPg1sxfP/5g6eIhgpiW7pveB
77Dj+KyANlCjW4qvedlHUoQN1IwxmEfRQrtIJwBPa8OtF75qB3N+ayeMv5CK+D58
wpSH3zn8HlwGJMftlqphuLFeJ4qxzbw4V51NbOxo+VS8BU612uLzTUts2Gz5P4rJ
cR4TMDL4t2Uh9Vc/5ZVs/lrufPBn/y24jW7S0M9kwmtHL00Z0XcAa3pLpFgwAHuI
tolZtyQqnsLJsASqSrvZTlCzIreOwC6c1/B81izfh6zCyV+Ee4ADR68trXeQpaX+
Vc8v/uf0kHnxyaLwXJq1E83AKFywp1Wy7Joisq9JDJh1miGuHwIuM4Rici4H18NQ
MsgNKc0Xis1qDlhlhf91E3rss1XAVAAb4zN1cV2cI5ubYQ09kR/7r51pf4NyDwDH
sTBigbfnzUJ3hLgZizXcKXBmhQ/dg2UU1rd+u1ClJ5AAOAPHe6goJ4TaQELG7mwT
MHUMBM7Sh/DZ+sxcmoDXHTVqlxhhZGASV1nuXQN2JJzMWzYEWxD9VMnAJB0uEapu
zxMJXnSaIRR1mHi780sXXgTcJOenPzt+UEPGcofEe5JJJHMmKMdDLl4GyZOiRFe3
nC5IFPYegG/2sO16uAeBRQK/4PDBT8eKc5sROe3FI27dSaqOvdN4KhcV+V2pEhKP
E+aMAwfvtAg6Z8h3CnqPxSRiBiq4aGMYbLCuwIpLwDL51/s9Ob4k3JXX8MrscVMe
f79To0C9I1rCCpa875fPSSypSggCrmpwNzvB1UXjBfygDmIIwkjFGV8p9fzppIKv
eSNkRi+E5miSJBYRh0Mjj5b+JtriznqT+ioAj8ua0efV7ZDamepnlrDDk0S03Eaq
iNX9nS516aX/2w5RdRCkmiFNNKBQgHpgncHwZwXzvzuHJ7zkRaMpqRweXbeSosTG
zRE4fh7ATTh55OYv5saSAqnbS+m7hzI5WD+ufIYD2VlPoc2Swpc1YMzbkmKjo4X/
ilep3MTxS9t54DpMitvUaqx3TNPakaQx/JXG86Jl3vm7pPXiirzTbcBO9frKsCMp
3z83C7+6F79LAX7JQGKmy5Lek9IFdx/ECPlC7XlLzlcRuKDQXx/6RRBhakyDEVks
lhNPj4zR9vbXeTGxQaCOEXLBtWBOVFhNGRIU0MeXGrMkVzm89Gl/UuxvRl4jNeEs
izA9zOP76mGxxSy5Oj3TFaU3cyRJGiGtJs8lvjTJVzp3FBCU5BkFfOrpo0IKWY+L
JpLLr2TSSz1mFCwwaPJ+m9pN6T0HGMUFcFdpuLMIHdx6QoKNjdk3u4fHQI0+j/Fi
ol6Pveg06T2MaoPAnf8pgxcTCJ4dksHa3nYNAIVZF0lIXOGoXm7eWST/XNjXMTgx
Jdgxp5JroxYFa87ds+7POT4ZfkCB6Vmb+TvhMUVBEYQVs/mzhMmH+Du7DI/zFCfx
JRZInZONqlNJ6YitbsjkIDBY2/7XoGKywoDS+BdivOxiEh7a2O5GjAx5wd4xE/M6
IWC7X0muFYuuaY4XMDkGRecBVgK3SHWBMZt4nfHsz/JOqaPvES3MrSGMEA15YXEP
t1W97gZsaNlGoWZ0we9VvozFVr7AEZl59c25ViyWr6uA5na6C9iTztswoKx0Q1Ta
IXPQnjqyvrH0pQd91RhUcNati18pUCnLCG24+Qzt0dvJ1+ditSaOjotBooES4zBg
dUWMIXNsJ5/ffOE7UQX7OsuP3x0rwzX3zMqAGNzhDT/ylSdjSCC7uplrHs6farmJ
ICGdRBCxL34liVRxIp0yNWqeBr3TeTt2qR8I0rlKhP8CJOd/PkYLJU3aT9++XEvj
AVYuMj+8KvRlUKYiwMMzWfrxnFKiOKpjlE94rEgv313Js2kqASmQ547+9bG25Glf
x+gqg1m1didViJ7fgWE5C9+343x/G4+u9Soko7FkHbA+ZEA2a64wGcMUpJ9VHeTw
yHkSf47UPrxVkkwfJQ5kNavuVPMfRBaLJ/z/OczViGI9r7dm8y/sZNTnUPGMOdS9
etZNWghFBOXCs7meQtTKmAyWH1bhFh5dvDGuEfEZ+MYHGPr9STWhbyR9+LkAMNuy
MYwkB0CPvKunNJA0UNUMCmJ1tlRMrTrP3LXqfWLf5WhTOusLv7ozWDwokmnaF6qQ
CPuJOyvpLLmifSXibUTGOLiTsQaLzeRg7aED7IMaKzLn1y1peRasNQj7qSZi3HTV
dft7+TUvOnFOphsgnaxTTcycVm8WT9o8N//Ajjb3dN90wzJc+DKQzDulVa4PGmhT
3T/bk9oBzcypIWpHJEA7q/Etkmm550NzScTTkxrmleHbj+KATnJxmppvmfpM+BSE
Dq9+bWZNymPuc742ccUfX+BWPSZZfqpQBDCa94VwQ5f10UGdIOJUc9ttc//NDuAt
HbXjDymt5pMV174IMcL5YEL+cObDGUCgcS5Ac5cMCf4GH2OwGiviM6qcEgDj4cvM
c3AY3Y0m5/NTJBwi6SRW6OqoaqClTYOGZSjS80XCjVN2AKImTLdWtg2BK9x6XFHo
aPTa/CcSGJ/47CmkWVVEvhach3IZOIYFQ+wEiXNzrRwQVnSaSSiNJ3Y4rJZNgW/7
kBtXuKxDUdvvhUvWCWRMwZgfDf0QZGJm1F03d1oyLgfgsFO+Mq+rBQMwd6/F9EkK
ROn0aUpRy5Tiz6ZnXXsdRISCNqTSvgUXW3gBpFFqngQkGcFPI/x/VgmLbQbuzUnF
yTGWC4bn2PSOTa7z8Lv5AecqqRFBrHJbE1NeCsef9gRV5c05zvdU1wcDi1xjk53p
DBcG5Qhb/tnjHcKPyzNJ2sH7hYmdLqlelt3BZZXb9dPA1/nf8HyRiE9qZDA4+4gZ
k897eSX6/IV4zMwsW2xhxIK78yE70siNjFpxAPzaBhQbwv7qUsItPHIpsYKEQae1
F3kz0Ujkz3LB7Z6mYqTsWOvuETA566uE8olg3DhVp/SUaKRJfVRP8BllxSAyaVrj
rE8AbFQzwFrXQ65DVbx1ISKdWKZWlmd5epKebZN0CTiO3w8bV6GTFaJvxJyX4xOh
k46cYS0jqSutIVKVKR1YQMDkXv3s9zVENeYasQggIcePP4+5A3VHaV8wxHrha+lZ
59HTpgRKyiXOcxyLacM6BC7SHurnDL2lGK1DJ/0TIwFq2PfF9ePnFTdS/f/59Rv7
6x1Nji6klFscYWuK70vTm4T/j68iMMULjhXvLM5reK6Irmj0FxT9ygLmh2C2NOro
P7e4/mQQUFysvAtVOlXJWEYAenbArTA2xvlnkEuGqaZB6HLIMMU1lqrpayWcIcpm
qoPxmw0bn23KxbeX1ZHnoQy7m0NLEUVbLPqfQfOt7CROmzGK8g7oH0pJfnUYwK3G
zM+JbBGuLft6HO/xdNkAvurxjmfoOko+HM/+5LI7pu1W/OcehgIohplcJoTVIHKt
ymlOGdJyqiPJkDLpIgPNtPGhRQr8ePpQAfAMSvyIQNQsmaIldDpHHXABfiM+IenF
aRMuXKyE5R8b+XDb8Nc6rEwhTwqVcyW9bRtFAGaTpWDi40aFfpJknGf3PvLP6MFs
lKDgYuDU8Rlty9KXQ3deIyz18d1chSuzH6xj8aVa9GJ3ycXpG3JhyTfazcTMCNA1
n9Z/kUYN1qqj84ZGABIzjBo7FDpdQ3hc8Pt8aK5Q85KAovZ3NsAGbJ0QqNF9eJkN
CAT2rSRa8IitMHuCW2dXsV7g034WtiW7u5PN/NDC3TjLEhU1mImiZoukukuisTq1
flk8CshTdZplV8LP5AI6Kn15Ha7snGGnridM9ifayME/dSROOqKKrfJMyUGI/WSI
rGGt5/cdMOdOnaHG1FBel1IF4nUfhIiRNRKQcij5zk73OiiNCnVAX92s/8lqf1zG
9MGvSgyqwDyn7HsI+Icspt1fmGL8jIPU+jEWmI6zOr0QplixXfKt8NUzEILATjeW
xdolfluweEeLzNqaoVx2sVSalBr6D+VBycbwku9E9z0R647fg0VHEIwYvObOHCQL
QWExKJgmSerfI4a0rneopCpS7BT3kCm1IQf6Vqb0THZhadwMqdxM21W8N8l8FMgu
NuJ539FeYX1hwKWf7F/mGG9iOg/PITlhJr3LYSDafwx38m1OAUpnKJlYKNYGkw7r
m16csBRv055vKkPptPkUPoooZcNGwy9oQ/DmhJA82F4YAOSCm2byc6xuFT0IApMg
/iVv4RcGXYOWi9iUsW0tK+2xu2hLibxbPQi8eqx2o7D5GbWUWiFWKNCkOTuVbbBO
NrsATAbF+CB3EJ10a9xvvh/qrYpc6v4KkEpFsaylraFkiLiYd4iiyInT4A2QhiTR
Tq7tJ/snnoaGQwUhI9nVpQUrs9UXPZ3RnBeVuF5kmEsUfnw2j3wBmb/H7N8EqPmt
D7OG3+5Er9bQW5gEo+nmahh+vNxHh02e9Lz2Mz0kKSvGgpmmpZu64L+XrAW7kgHh
vyk+atIIprmFU5voAy+6c0aXL46PfRfop8kxdZfnKdIWmJ/rf8gcLle55i+d6HKx
qnI6dVx3kJ9OIHJaXXTpfQsiUdfKdy0mcYK86G/0UzRrWMYDFcZaWwMx8ZuMBR/5
BECIxSETuhWRBJEHHZgW77O0EzezGYxAAlnqTXnqeakpncI8+JGX2/t50FEBc6UK
KqvoqK2Ll0zXPs3JLVAmw1uRsETMkLBrWKp8d0Affb+qc6SYowpRTXYLXt8wwfWE
+1g0WUNHMKN2hu2lpSmAt4N4k5OcOVR85zjdoTDMNUycdE2oh/ry6Wovcq0WjJrV
itgH0VJVPgB2gqaaZsXUi3X/E0PiJq0mMoy+xPnRR9AULmjlA58JZUOVTefQSikW
+/8lxc9tO+7gTywZMLWV4vXiwnD/PT/f8nsWurWtWjk+mnd81585ML4x9s4xRPwI
cscfz7RDOlOv5tdxvptL1L7vrW4pXsbsfFTLA7e7/eUbcZsbkEONvPE/YAASCjDE
1OIKfaOx1CSqZXG2Pqi/t5nkN4/ZoPCVHZzbpE8gloChocRsTa9iO+HhqJRCKEEb
5gw01hWrV9u7ohXGIHPrio+7EpLF+l3oxSUXkNxNGTb5JFj0kPFAGfTazlL4GsP0
dz9csaRQ+WUMGWFrkOu6n7pzl7Y+GbNctHW2VanBfENSVgPzyNLTgdDlmexV06df
4xnk3pgX8QXQhOYDnseqFBvrrrlGGP+COwo47Ojk7QcxvAPEl31gXPB1e/jUob3E
WoKiPblIbLPzQzI5+6WEsgIuZzQU9wLJR3X/L3INkLy7Bg4lpYLKZ1iK+XE0SMhb
6TJuLwWbb/c05Whk8d73dYE3C82xOdYImOpwyymXnn3oE60Cp2ARCHe1IFvfGeM8
7m/CXz2Q9VYag9vtuCOORNwoum2dmOpPbSNfPJm71OrTJNXE1UhSu8PGV/1F4Kmw
kv+Ynle6bSonN4160V7kfl6YLnKJ+yxADTjkwl2iUzEThZQKCR/GLRekMQDni7zX
W/cN3tSgMi7ZgXRltfAY0VpRl99qtOEhWnxjcuoqMS0zyYEQ7LT7HoLqcI+SUnNt
tGjnCYaxU1DLaDubdbNi/t/xJt2y11L9qG/WMGp4R50IUGCkPrCTEYtdiEHDw9/b
gdt2p/BcTboSNBB2jJ01tlFrnVQevilIIIoFvDsO1g6tY1BJGae8iUiXcTK7WS29
in+He9JxFXVGfCQYHUaW07/BB1OTK+22/PTJ5naGrSKzHE34g6uclpXHN6Furc3t
GtlnXDj/aEZxrXEJzs5gsbemCETLVZBgKjMgSIx9Z1IBMcIpcPrxymFxNdfB/Hei
kswmCZnJtThSrAqRK+sM3LcEVW4mlbfjFLCt7ZI8zaovxIZFS6gtCFhSWglyO7EI
tsjwYiq69C/RgOVIQhAufeAJwlM3CIQHTYMDQ/D2Jk5ompzO2R82o1gnwCotOpse
gZPHsAlAeFiY23FuHq9R2I4N7pqXisW2RPYgG/v9Yv+zPeqEEB7pKQ5pcuO+dPbU
vqJJvWnAsLY93x0qjEk/YMlykiXb1e0AwDnVYVjTt8FbbaxxbV+jbPuOv4aaHbDm
KSgg2Ap9fMWfOMCZ/m2GfnhW7MQ9XxU6woMGyUWIA38F5H68Bb5uXMvL0v4AMMeL
R+94eMNFvVtOpvuQnkwBtQLQ3CKe0D7/WyJKW3BNiiLhvP8Rbq5vVkkt5xQLsDRL
GegJiYOMn+1TalKHHKKD6dJcAdRU3caeCHq+rSOJb8FPY/XveJhnMYtucnrk247N
CgcCeLO8Ifo8MKNdLy2HASWDGco57ZehYFcdPPKTh+7nRvBlhKDTPTQfcyr+Oe+k
o5b6Gw840EfqyjTU30S2Q+iHPKLVDwq9TTN8YMFyUXHeH2vNXKT1Ako3N4DLULlN
rEdTYVZJ0coOTqvVjr9OeSnyeEwvgvYaLn6YXh3ybhHqbKgvBVpuFV3VKgeTNsIC
tQfFZlBNzn9dGCjYfHvj3Azbm8gXwU8u/nNHNVtCt2N212BDwE4U0VbthYxCkudx
PFKSOM6mbN92BqvO52X1R58jV9idmIdmGIfck4ZJdn+JWKgtHCOGr3gi9l2NihST
5sj9Mdbqm38qIJDpa3Nz7uj6AXkbqEWs3GSdvaVjyI5Rrw33qguwNaPM28harpqI
zYW9rFwET30tKh1jOASL8AX+0BkAuDGtxz2ayRodcJb1tr7wLAW4Kb3PjOvaUz5S
IKwW4/aAI5rHeH6ULZcb/HzhiraKQn0yE1DPjfKBbw4BHi/ZyN+wcTLwpe70iLQf
QonKij80HpWqYnNyf3fkuZQUMlAcvEYsnCm6nr5gt86QSOrPXZBG8rY/qbXKMRHo
xjjQor/ND/nTJrKeE8bqGgfuncZai3I1gdkn3/GRgqfKIzE9zDWSpF7cc/1fkNpJ
74k7lcF9y5Uw+wCcyaaNhmxUiT6qlKtF+zUuY2C7UChcWnDD/TImyIOXnRYcRIDg
5B3O3E9uh2yTCY7yJQeOlSa9U6Icmnx943vNwr150hqWqSC/OtlLZ6exkiALTt3T
CBOasGolz51wDrCfpMwRzktDvvEqY1VoZ8uyEmLts4ZhPTE1FqGTLekzXBRbujGB
puE85zn23Ym+G5tnLcUX1rn5S/7BMo3q8ApuJNtm4HzF66YmrSVYvrdEHpjMwMfr
1q0BNE8rn/ujfx43vJBbs9vDYkyGQH0FLlzT36eYfzSW8PiBNUsEWA9m9mvGPnqY
2lSfgKRXwnnVGatAM1q7hekwqL6hc/xPXe1fuzoX67ELN1IF4x5cW4P/mQ8B9u3g
HvFy3ge4n3uErYQNy047q6yXTjtrpSlstB0kJlkNFzpJWc6NI5XaAVXCBtrgRrSE
etcbRCBDTyxwjMZXwdMN+KRnB09uVyiIyFULRMmofF8Tdd6YACMBmzBQXeaObo58
alPed2aHWjSIeXPMZP//eU96/pIww0EGk5gVys/TgdxW7IyhlzEXYDJXrLgkpVyR
+FIGmCkq5WmokXVpUq2WOgYp8LClSvrnfp5s2ypAmP2Z5H8xXQb073KH0OfZ2NvS
1PH1LKYLjrRLlnCpbHrAs9A80TFwFVJiMXYiqcRfo/uNfcpmqZ8Ligm/dgGRUtrv
0v/YZQiw7UtkPCziQGIR9m+ivKGiMrPWswlbq2Q71tRpsL1V5+XCYYQpPed/9e1p
0wMAvH/T+FGsml9BNfn41zbqLYpOAJ6vY13e8ksixXZwjpjX6y7YmcnZw46HUCCT
M2LjDZS1kao0cDdAp59yvND/vGjiUxzL08icH+UYoSiW5ipd+v42fOw4W3gOrpBp
3Gkr7/JUMJPAREvW0OQEau0KqlwqmOOHcbryXTbr1054x7EQGu6Nl0zrW1/do6h3
cFZm0ZdjL7SL6hcsToCv1H+KjaH+3s3mAabvLMV4JvwVq6sR8ZMp0flvdKg2+Ian
iwrJRwXo2TsV7Tu54ruvCmVILqQyVaYeOLJ4wkznOXkO3JnA/l/JECC8jf4kKLtg
zh9XH5OTKDI4TNrscIVUHogdIGWCKPX3iDk404MnP9pDuvs0saR8C6inpCd6xie0
dyBzpietyGbuFU+xmBFHqnri3ckTIdMCOqZ2MCDYdzzMZex+6tCVeWa9wH2dHtGQ
DbmVXt1qINziUMzgUDer8k1g7ngCEsL5kBeEpTtJY1cBD6g24Eo+EtscS6/i/WL5
7iu3SZ5C80JtRuPvW6OQX968Or60OZi5FFMbFEojo7vgggKzZqDrxCkHhUZ+QizX
82D67NYkGiQkKm0qUbo8u/rmbY6ke5Y6r0M9XyqwuHfo2rCtuT5f+4LBfSpDBfaq
8ObQfodO0w4JR8czS0je07TY8kPDBWJS0vDrPI5QSLDDw2z7FVRay+L+ecvkKrTn
AhkGj5Ww5gjj7VIZOQZbYU+5+4O6CmVs0H3saq5Jl5XZ2imAAWGThrldRVKbK5fF
qcP96n34Y/HHW4a1AxELgwIXPuC+9QdyBTEy16RP0ZuMlDACve2J/596iIkruUar
3EJCkUv1oKMns5emXBmmMIbzKFpXEK309GRTjaEsanTMln1KVYjwegdT/wvz52t4
qzFvTkYyPh3tdmFQlgLwA3ve+Yws+DkGsoXPGD6+cYg5THVl4ZBqCAbCrSv9aFNf
iHv9DR4jDoFcQdl5Z3p0lCqWl5EN1H1S6ERofGtTxEZZachoc+V2jrI11dnp/I7s
s+z7iUd1Buvp3a6Wi8R38g0EQBEUZ1MYuOF1MJG3iCVPWhvsQW98AKyO6kcRDiVt
COs/vDI18OtybmcVNSwAW2Y4JXdUf8bp2Lpqpo1V7xw8NFqBAH5eyyooEzrm//Y9
SafHLdOmIC9iU/lPuvXt6oGJ470tY6DawyJbNL4humKMYvmLnAzOkKiPEjOxR8ZG
DmgoY7qchoeplJC3bVM2rN+bVcNkX04UTd0sQvqt48D5JS9Fs8Itu21E8bIcR6RH
ekrpqrjnXy/zK41gG/o/iJDCNpea7HNG9mcs8MgIMelXAm9j/n70uI4OWNCzQFyU
sbGmqVM88EGvlCcPQU7Fwl09AnrbJ2uY2Jnyp+Ju5okbMgz7Pi9YaYcU+CanthYQ
Q7y3a4MTNdli37+edaKGUGSLhzSZI0wqkDLecC0tb8h9U3D4DcRQodJpa1jqnqBQ
gbsRwm8ntWI5gL4hRxETfKFz7YytEyDzXhPAERlPt1dgFa8zdNU/uXjSv11hkjca
oND9ZYQa57NcfouqKT5A5wqHDI/MFYWWoSnWpeNow0mi4cCvkDQlXuQNxh+grDqp
U9QOkgcqvhkrl4AeqRMuB1VvSOM37U16xVaSRT1lPbUMMLgEyb7cnTEDemxU+ECO
KQ2JPCbT5T6vxBIOBtN0Xw76z6RtDBmLy/zTaaU+N46bq1SmdZweHGrzeMRzFEr8
wd/LiRVZrvEgI707WWib0vMOtG5nFWYuaYgVzY3+OwIGjYTr5i0cLzxRRK+7v/1H
VQq4iU3o6I/y9/Ay8/8+ZLFlTsgjkWVs8jf0siz+lyRSXxpcZHCeMHVUaKb5B6FE
CT+0TAWNZgWC+7T3m1c6rn3QgdeoPBdZC8YXMU9EjnqvgJ7hBtXf8QJPQzPGegb6
aSmF8unnM63hXO188lFy1S+ZRvO/zS/KVkSmBjLtPZ1zpbUfvNrxH+jBVm9g1rJ8
i5DmIvmh9u4cAyRZhWkDa6GiXn+H2LS/9PfsjDZHl7lanN0IYz6/hcAs5UjCqe0E
1ou9ZoERnxZveaOO/5D8Sj4ji30ddIWn3ALKCF2RBseKtRZfoZg+9z0CKypspqte
/RvJs248+zvXDp7GoHQbm65X03/PykpUZSiSojeIrn375wkgN3uDPmudYScdXJd8
QMBSpNaHyGjEyTJVX/FE6+rBLKD3G9FrIXGNd5VnAzlUf4zotJGJN0zfTQho2Y9b
IqmlrGthGs1/5OERmPuzsk8Q/umcJpzvbRgDCV3XVIHx56ZQcgXRZKikiNxAWo4B
a/ydV+e0mrUPaxH6XXfpwoFB7tCDABtqLc7g90rqQW8LfB3SJfHP+Vl5XBrJYpN1
8XhuQBA+QmjlSumja3XEKx9JAXU5OizBhLGlYtmRR1YiNpO3VTnhyN+kSHqFMFQ4
ruteUE0YMDps3DBOk4oBfFBKk7Hq448cPLxJFrVk3rrVC/JPI2acXhH6/kowc3RN
z++wW0vudeYon7sNKTxpvXyEBugztgqr3E9aSBEvypSjaD1wbN7vbQaHLXBQSzwZ
RLOqPDTC+LnnplkCZdUyLILnll331YdMq2zOTurTxQRVTkSV7V7GZCvnEaiwfMDV
miuNVEFqvDG651kNgTZkXP6uWw2Sa+eEOkFRrWlceILtInFTztuSvCSj7tEYyNJR
PzKVfCnylwXfuNdSLIrYjqdE6yr7lXJlQzjN2NxDaQqA7o909nQA+sVvyKVYjJwS
A3VjfR7Kui3nLeYNQvp6kqfNIdfV96vyv7+hS7Q+e9i+c8YfQFOy2Pu1zl0o3lGl
+f4il+NDPJ94bsFNMtr1F9eW3nYPzItADRTGq9jokB7yoPJZ50h89E6elbXuQ/R5
vTr01Nsla8R/KatD4IeNHfiSAHe0Deu1urDZv45o7HROpDT0V3UGQLmf8rujd9OA
GOBWPe/OW3iA489vVPEq3glBHcSWymLEbX12K9MQxbz7Z8sqZQVpo0DXo74eVqhg
xvxKjYWh5hoQEUv5hpuZAHzTnY2KBMcV8HLwXg6Q9Qgj39I/+4kcxFGsUfKkGK20
yM+xvDSVr3duwOEa+8C0FwgN2yUhGsL0cnNKmHuYIkttpq8ey1PSrmdOzhsWeVGY
zR5o5wLdpoeT++UXEEft5e1oKXqvpmkNikoiNYE7LU2XwyVCwzO6+Abuuj8shX1y
g8ePC+7qLAAxY3B42cMiMh3eovUVCKsQQr/baI2fvydGHDzttcovmQnIStluU3Cr
PmKwE6OGq8l0qoIB0nE+JGL0NVnVXQSqVtJjlfpqXAxZi+pmUWiD+MgGvdf2fUp6
zYg2+1COWsBsfeiY9lkj8CSeHeJGm+zte0QwKAXUVVx5QXwSoiTWjqbS0hsdPblr
Rb3v2NAm+rHlCO+6dKq0yP6GgbWsie23CNtPta7jU7KO5F0EWPPIWpF+E87cL6ke
0bKzHqBBTuMFPUaeLzzUbqsALdeeKEFO7d3CppdXxqAC4ofqiJLbKoqcf1a7UTCO
iBPu/lyt4EuWTSTQ+CeaDlgR21pfZ/OJPCPyNUegnTTipyG5j8ZA62nC7IYjULCO
ky/11c2oPSDnurXBYS4nIEklC84XeyMi6TiYIfDqa9M1yPfDAJ6gkrdX6fEM7s4Z
ihJjchOmOczwfV6Uwo1jB5HREXkoX8VbX29FMVWh4jXWxX1ejbNpVOPi5lBCKrAw
xBxOt20ybUQyZTyB3bDgFNQUY0Q9XfVmnfJn2JiLzkiAoMHlgk5o5YPKE1l49iYF
xIlfdDPv+/zNStQ8KhYdRHmgJ4f1xvTCdgn0ed7k7EvPgoDEmD8epTQPGv/vE3Ns
WTkWt79rAXW1Tw/+RHKTVMwrFSNr6eDAca3Y9BoJDn/4b+7fHYxoipwXNaNiAlqV
2XjkrqBNlgceMmH1mEK/I9NhraO6KXyM48kwG042xn/7CYrSLc/Upf5v8IumorWi
mxcvnj1K0BAxjSzcNnW24j8fvBBoHbpS3sOESZlRWqw+i55Q0KzjH2BFj6sJ+CbP
W/zCKwqqoikKqYBz+EXqG0GamQ/79ldAg4dBhH0th1AzkNpQregXpPf40ul6+V/Z
5otayEwJPYv/ccfLgoGbqJ9pZIHIh9Ty9s3x2h3+I/cU6wiRNPmZxM9tyAosoE6i
+oQUcD8hTYpC/UvK80lzId13LGtfE804I2kxvhYIi6oWMXRbH/bDyaOgOR2itKi6
uqDaDKz5IEPgR5w8ew9UdOl4uL7Cz4F7PQR5nBa8XEg/JTu5kyWFq+wpm0wY0ijZ
Gny8kDBRS5JjWb3PQbZwk24NvBCZeyyFjaJGQ87YJIn3m/lS3yRAT9nZVGWC4N5X
UPIheqXBTVJo0LK6sihtHtWSNCPNeEnRrs4qyPvJhXUePmyU0XeFNpqsrZTaAaGC
RNIXMuuAg4Lcd32JTye+bDNP0DrOBF0RnNd+/p+RlmIJFnHgzTndlIBaEuXd8Qc3
fn9DWsEm5/olxi2IuqDQSSVVdMgqScpSPBIGJ+kYFkmA6m6C1581z+CahS0niU4R
66Em7zTBb7CvnHW0hhUHAMfhRw8LSr5X/1WYzHX4OLiDEy28XlEOEHjRFcAAzPOm
jLkaasO5go31mWamNI9Vy4TwHJJ/se3uadVni9+GPoUdCGgGgTkq5VMlSzuLldxb
rcOfGQEeQnTQKGVfFADap0kW/hNjJ2Jt3d52Ly+ck65WaPwVq1YC0Mh2r2Zv0Uuu
ALE2ArxAGZdMGOTClJPNuiEBkrzvkezqWFOFvvCZz24sRARhwL3N4lPPSLaOqATJ
VV46vewwBaFzp1cIDhH3qxbL7aT4sNripjmBX/fmeH0RiuJle9Kf0uJWS11NYCy/
knpXlQnEpcd0Wy2c59LgFWuHoxpOJV2PYPsGIr8aJtJFE+DvwjuWDObqnJFkbR+/
DJ7ibhNXgvA1Lkp7ZXCWapz9oIG2B6bGEJDesKRw0sIa7qm6HXlJrcjFYQ3SfPjg
5c8qjnoOKhUvHgzYC14kPSISuie+vpjkfOHVZ/nmyXZm5UtU+mV5kI+Qgi5/NYDY
Rmf3hu653QQe3HcV8p3pVL9OaK4NdAYKzKO7NQsS9SBhk6rrCQjP82W36+d7xS1u
zEf16KUklqFMmyNzBLwPNhAtyJ8uyOefw3UFSXer1m4w6vJVAa9XcAVryqhCRvT8
49xsqibSbLWTmajtEZIbgY0H+1p0BAmv8K8mLFi0gBbZcCLDWGnc/XqkHtW3TvuS
fq27liHBzOOTItrqURByDtX2ZQbxlnqqE/ms5Q9qcYmyVnWIc9jnt5ym48lgLHmV
m11emrsA0TEC+rkPaQd4/N/OIV8zIY+sSTQV0K32hb0dudlRfa+A4nVBXLdXlk9p
WKZ8ZA4+OQbQn5xETOeN/PO/ZU9QhEx5/n7Drgr9N/fOxirJWndEfCjbCgRsjNp/
vxTy5gr9/s1aZgEjcPPfn1S4Am5Kz3sCuUdFkcHp/6CDe51xtBUzL0rolKd6pBMT
X+FY//Ar3FWRtldpAxgZWM7uAji/7g3syieuP+BjrZ4SmxMEy/+zVfYgH6u5zGMG
kD2pXBVpmVDGXDpXMvhJ6WrxaF7VI42CeAw0JvSleCB9L8+I5zrStheg+h6FHSkg
KiYEzQ6GvYP24tNSj8DROJ8DCwHAdYJltu71POsV6yJoquMo7JXnejaHlnjpucdw
EiH6b9xkwkDXMA6Cz/wQ+EQo6QgVFaPoFMoYh5+X/QSDdIPy7Cpv3EZjrx5oXhVO
XkJJJ2tIUEUFmxZ37FvFoOmk6Bod08mFOIMyiRQKh7Lt6Gowj0IvCYFFJVNzjtfC
N9x7Q4pfJRs5vU2F+Ccu75vKH3JU+pVu+a5kgC9sDYP2uBdIB6F4cFgXI68xWUjn
rc0zqMCwIyzYhamBg+YSjg3pJmMWwsEztin+KvUNjA2t3NeNjuJQmTNGDK7xllcf
eL4APaVDi+SnwZdYhMkGBJXh4Fvt4324ivaqY/ghoiUA2O+gT3bB3BHoW58mCg2K
5+exusY07We20hjLKAIyaNoN+fo4FNApDr4A+nbKFQrbFTQJh4fgRIs9cPkRxHDZ
uNuwLdmv6VtVgX6Dj6uZAkYtF/eKt2fym5TQ2OQhLU1q0NksNLkGVziflWFu/vaW
tGU4as03nwogegjaCW0dlyqYq5nCClvUWBRKT8xNUDfKndJxh80mrZ+5r9rIsGr/
XT8t8xQavXewstT15c5+gSMe2G4TSKMLz0TbADp9/pOaf0GkuLuNekVBLq3b7Apm
1/dkCIr9VDAmOD8OEtKTrnPUU+AUUkN4fuFB/Tap5sJzlLX9c2z8Bd5grcG/oqq8
yQ8M/0wiX6FZRz2bJiFCy7z1O19RpVk6+LpNKNl/tKvcmsDSQ+4noWJvNa4lZhRC
NKOm1Mv7rra7t/9kQ+6I8Dxx0sWoCcTcmo9zMiPuIDLoajLGycznmWhgsEiO4bOx
f1vCLutzliwuFQBPNWYM+cKHEr302cr7evvvUq0qLqxWfxGiKWVHQSyp/yc2lL/r
jsTdd3k6GLj5lVfJvFr/FWg+G8AXB22Jk7YC9QKo065YW0QsWmE6Ej2DWoqLnJxV
aw+4pbCuDJ9XjnyTgQjLofkqHB8zSC4o2/zAcOVtw+49nwdGPKsy7Th+8sBgC7LC
C+mKkrKXybbbgXVHx5LuCiKhDqWuKtqpiDpwuWL7Z1nlFRmFMCNjb5Al9FW0djvW
IyBG8xCwoK5eZFsvxAnHuxH/Dhwd//jrKOioig2XZMQnszpDh6oIsoPMgwza0m6K
lDV7BUBO51TJX12jcwzeka92Pyh5XOBXmxXTqvAWPPTUNBjnD1MVFdh2OYAuCzL5
IJaWfLXTDL5NXjs/feJeDF+sIYJE1z111TEUMTmTSCRBWoSMmhQhORtBeepEzjvb
YuYcC6ZxwVTuWV3NXMYuupoVWzq7koahmgGKXYJIeRLRBH13E+XkualI6pFiNaCV
EFHggTBFGsCoQwtRNL7c/3CeUX+c+aFEHuPKokTm7WO0TVLWhixYqO+t7tIoJaaw
xYesLqXHsUom8m25rtL4UbVuH+KpeK63yRBZh3jKbqNwOyeHcnmahfOQRXjD33lk
qfo6uABvSV6VbBIE/3TPgNMqn/WGno1JAZ1K8ik5qroe+M4se+p367DDRaC1QkOV
L7ZwMeDrJ4D+USM/cn6JTB7j+9SSOQ0/r8+HiEITsE7RJby2A/48Jo+sJVN+CLH7
OBymeiaWaz6DGp14DVMq8iLUkjll0ztx12sWNXAAeCnOkU3gSGhmqEzbe/OIxepy
UbBRtqLK/Gqd6wc1sPWEfaAJ8VUYcWDBAbFexbI0QlY8TJ3LoCZZs6+6b4vKzR4G
t9LAQXvkEsfRtyX5C8CXyDZKlikBWUrzMo2xEiUftSWAPKPo/IcZob1MmksVEaTY
WBEnCLNxttbLkKF2SSL1zzXdOC/GM0ycVsgtEuoG/U/EODJ3VtHve6C6MyiRp3dv
CL1qyRPP8D3V53wvMDx2CKS3sqn5LpJyO7w0pynF/VN8NNodnMuEvf6xXdqTsZD/
yrmsHBJ9qcAk+P4uwFgG1EGl5Hxuej0MRnI2y7kHPThY7ti281281YYEewSF6u2q
v09tSIIoCy5g+z5TWJbhxOV0hE2EbOlx2Wj/D7UTqj6oT9dvQIb6/FqCWTPpBtTU
9dbC0GYnAnaA9KmZxNGtZRJWwOU+/+gFw3ZwWm98LD+pUjP+saywl14FEKA8FtoW
EpJcSeSmqTw0ac6nYAlWAmjpEb+ZNqr8+0kZNY3y0RjF0aRCNz7RarOdLoGKxiqh
8kGdUxNSAdK0czNMMdhDtO4R1AOAaqInRaqF+XSUuQ7H2J0hQpp3pnORZjRmIINH
wj73D9IfazSFQlgUXBfTp32BAmk1VUh8xfgB2WwhhCj1tHfqeCTbGeki7I2bOLkK
GNIS57PrwvJ5OMZQmZSM16RbQWp0ZJkfN8d9TVCLZ5zfX7TmgVo9xkXHP1iuD1+y
hmWdzHOh3dlnR3DoLl92PJO2RnTp865YclN1ncXma9Wb5l5uYdebtW8IXtjy+Yyf
2bhpuqhFc3u5nKEUivgMzeZ1j9d0g6lEMu/L6Jt+4zVThCnoPP0NFFr5EIk59cLE
h+Ra/ge/I2zYQ3X6X3ScG9IKVWRqBdNherj8e23Y4zDSa55BjlDJWfZDnhxsVh0r
kfbBr5ZOVsF6Va2tb7ru9COJBb/5MBKJQHe3zPgcjIIr4072BJyo7YKShjmxP1my
r0oGKo3bhLMWsqt4VF8CkvekA0NGjqbAf1UhbRMt4tEYPpUxEegig41/bTRM3kMZ
WlTOqWqcmhqNudn2Nxmj4azyI1T97Ke3cga066aFQxghgA1Aaypa0tO4avLbVcri
sDDVsXr7iqLuO+Cv2jNgP1i144PcPJjVZyxch+R98QLralfvc6aoygXPoGwoKlGd
8mdlPARglOYwiTBfHKkDAOrB/a/ZsdoKPAloGP7GpUuOqg+Lbvrz3FFwQS9e78/v
Ws8dr0jkCOR2a4kGwEqlhyyPKs6pIdIHwZgfAB5ChLFq8NNW+pj8+N663TfO13KY
Is4zQAUFfyokZOAl6DtRzl0sT82AUAUnOq2BS9Gjh+9y+tLBbohXX1puVQvtr0Qk
yfaLt5hTvNGLjtIzPC39wy5Lwzjbbvryev9RP2GTaOBV5L2ZrelgLSCWtXwBqQWr
hYktqUzNSwb6N3GzxQ9iZMm8MCB8IomQmg5ZXtkKl3GHphUX1/KynsFgRAyP5ErI
c+Z3gibiM50eMrI2+MIdtrQrajjRfxyoftdhxWC+8lqvtkOFPHhNpz0lIxwVAWf6
d7dMfwEG1en1LpyHPzAnsw0LZE2tDJlGlWvKegbcBqQCHKzmcMFG9H/9AwqMsaHt
vJMLObJYaYI7cEvSpRKKaqoyaoHmcA6J35LyNzU7Uj12WmBT7Yyzy+IdtIJfFLzm
PO3mXxte8aozHJj0wjvtgyn7ReWWVKMn/J5UuRxEK3C2Kfe7BYZW2FxS50TjPIcV
leTnfI1HmzRFrliUli3i7ne81kdL+RO8rqV4sJdkwqVSIlciltHG3BON3DV7oB/k
5/Tr6LxtFknK2xjVJvlyKjFQTEEGz1x/rTdbRAOGhBmq1nyrlI8cv3+dX+tV1dLJ
b5pJ0DyozKQ3/DV2fyzKuV/jIeobG6gk2dBAFH6FHn+WITcPZa4zcT0hgkJEoJlV
kyfsL3zhQR+n2dWFAm3rtk+HNGASxADJMtm1CjM5ofI/8DsP0VttNh2GahtNt4yx
lFvUVa26aLEyPVY1+tb2UgUbXZW1DyEFVfSrSvhiVOpIkLZk6wHKCmF/pusbQyIQ
UB9Lu6yGvCG7diZqgcKZBG9iO/vzWjM1vHzmu/aECQCOn2fpK3j2v2n+KuuQk9qS
uYU4YluEqRVVWt1bpc4pnTmycQOg8y8n2LM7quvwBU9ki0FKGTQ9ASl4/o0Vub06
qwI5zOVjt0YG+fPyYEP0+KAwfIAyJ3o0MkHcfpM6iI8jGsWnMbSSVqeQh2ruqUOg
1CLj14G1FHw0TjYE7pAppFvUpBj+mUNN0H9vieExq0+Foy/X1v/O67owT+UEvmMo
AjigiGen9TZM3jJjisq3ZLQ7HTzFo1LS4qsgHVuMhfWITVcH8tgb79KMS9inkQ6U
Gv5GVJ6oJSHr0HDSdhjEGGs2qfa20rr+akEc7F14umIxNeGRA/v04Q8xZWDnrFCl
BxWkF340bkizEIGWBifwhWmbXm1vdg8dVDQwb8IGbgG8tr9sbdl/cCtiSEJjKq3P
0GLfZRkHytxkhiQK3rbFgy/50VJb7K2+6rL9t7ZoHLKJtyeEt9QGUdOy813r6Zfw
AwY2h0i2II/ilqq4x6fpdH/Y7ldtDNebOQ07wshKdtnPJ/WdT7ILmq9PxfcjULI8
4D44JeP0jktncwGtyCvYc8XNAZiZy4PqWgjwUFTYEKzsvYebTmLXkGo5y/HhwsPF
osAiwYAjmRY9JS+XYO3KvBuxEC3s0dOvCVkF0n3kUjljhx+ZgvDjtYMpH1j+bPVV
s+30tGVqLaok88SYpH+elL/UfFagmnspoFjDcVv3i+aDnFcuWJB90NlT8mZjxWTT
lMvcwSHJxpu7igbO0MWcGu58Eb2eQCuhb9WDzhhIWh3MNptCKlvXe07YMMEugxQt
u2qF2YUo4kFRYurxSrigX2hS3bsJrgXZIqe1+px1tfUYb6b4lBItHbnsZzAjsL/i
1Xu7JlSbL0PxzclTVQ+pxXqG2HB6M7k3S3ua3F85ulps0rP5P6PCeUmq5NgswLQQ
jl/BqoEsXZ9BoCWx7xXS3k0QtMuy0AlJ8/g7pFX+DVPY7D86lGYENGyMY7Mr28eC
1i5rdf2Hnz7mJtzU/v2yha9kNWaAMLelMdZSILuDx3/JaU8wkLjrrOxedEOW/njL
Uh6CumO7alY1RzqqRQPTuBtJyl3lpAkld8p9Y49yP6gCruJaOM6KdA6Cy2JHJy2G
bRVeF4f1UmPPbFjRxZu/nMI7l0U29wyUNm1Cw5mmZeSaLFAzNMmbISqSQu9ggwFX
dxasfvU3HVceVZ/0ym5Tx79V3CowJuI8gKdZVpaFwtsr3GSJWK0ozjJRzNOhoK8y
8UHxy5wjaI25gxNY4DI1DycAPaXkyOznJd8/A0c4SWzqwTl4QKgnyB5LAL6960UN
p8aRstrFSJs6sTk8hKU9xHf9jd2nYDJj6Bi22yRKOW8QRCm4bXys99FGJLJPpzOn
+YQqsKyucInpdfRtDdUBOmNqtWZ4Gmp0g8Rvox2XrxnLACYHAaL5B3BAzkR/N4aW
R+CvDK3rlWikxfnu2+11IL4rm7wncDka2pM+6rZp7J/TWxU2ufgK3fq18gxq+ZHG
3tESXzJLW3waJdnytMeBzVrKyhI65ntZBObI0wQ3wL3wescQzuFaH7Pz8B86NNQh
FXqTsZAqLGCPzFzRxx3eO6NlFhwiBt3Pukh/0bct3rOFFK4UtnYOc+cDBnQEiEzI
wIBBgrFV943yXTsB4GL4NB9bOC+Th5OY+aDRXCkBNxfZQSuqMtjzcYFf2lK8bqAk
nEGRbIjurdHn55APJCGgYDWk2juROJEEa8mIWb+EJePhJExFNI4G0FPfMYpTy6Ub
Lp7NPBWJf7OQda6+jTGIzEl0/rIOgj1bKy6KpwIq1DNHrf1tU2OuZd+96yIOudUg
8SKU7scn+DpdvgC4umlWIUCT5qZwibS40z0fQh5WC/Gvcl8oK/0picVmUG4j4htY
1Y6sLfWJw0U0+Z7oYYWGBs5xkMO4hvMsKCxwMg6atD+HmW8G8e8gVocELFAcYB/+
9lpicTp6ziHzjcisH3oDCl40zOu2bQbI+mw8EN2fyjqilr0f5KlrVW2z2I937GQE
KRSGb2tnDPvPPTPInWofq/C+gMIn9IGijfdhEKTq/Eg+5MXcttjpBxOQTzWNUS2y
rq/43hTodxzuIHXJFy3bs2DbIp9qzS2ws77/cVTi6voudnixUiz59+l5vTZ3xLEt
TkQ3xQIzCxwUP9/suia/qRotiUFjlMZKPj4DCoeBm8Dg8tYYPSsw6cqmD0y3XIO/
i2st4CEnIqvlkJxnyNAOOIxEyhD/4rQugqbiJKKorzjx0i/whrf1zYcOCdpEv7hz
nyrc9s2SBgyAB10zVQlZMEPJyo+5M9p1eKgOdxStm3MKe5oiDFm2M2dORJ2PolRp
0yAjR5KI5vwATjQe+KW+8bvWXWJA52c6GRVqC7LevwOcuMs0RY2FqQcRwKfxVzNj
/rwvzZe07+CMMALuoSfes+0kfgsqYTROo3t2u6yjIWCCvCAJK6yb4rmy5PAEq82r
fftXoyVXecFu6evxUgBvWK4CXIzX5mC5PBRBc/3ckt3XmATwbnevOFSjp81cgmRp
vC+/Phx8HccGWUAiKqSaYL/1fLaf/iZIPY72xH6N6HJAw2pxrygWOj1yQFoj7Bk5
ff5sxNZwQuH8RKR9aFBRzFdh3iQI3uDM++4MrkomuwbTnD5GTBVGJE4lAFpX/f5x
JHggPCHuXEy9SfH7hAtsSui+Rh9eeAk80qX8Vh/D8fmOb3t+VVeyE6eB4KfGYphZ
u9iwlQ9EN3x0X55aLh5Xn21Wc+GtFfw0S495GKRZFALCDRYmvWB3TS8GY3qX3Ykz
GVsDJ4Kadn2QZid3wsyVbHR/4UwZWygS0pHPApzPWcgvVJiP6AqJbmt7N7RPnHeg
C6t+7hQn2vpBHjppLyN4ies0Sz2k2YUy9lJwIkcLFXslapgWl2yvyhpQvBRvtaER
+E/yIYASqNdiaCBTdyOUcNfLyV2bSpMgaI8w3JedWOZKUUf8n6U+0RSAhXldOwdF
B9i3qQsI1+xx6J9smabBV5VDbzieb45LvvLCFs7ux1gDLKiNuo2B9VhIdVNsJmi5
6Z54B9p/Ozu4z4N2RS02kSqR/H3d5xH7SXIjRl5+zMu+O9rjoU3uGgeCw3/bkyQ0
pqYi+b9mkuPnWtcjSePaez3ScOkqijR5MKWVTmHspzaQK/tXzLa699yJsOU7V6xL
pvsZ79aPC3d3Z3LAa7KYsyn/pGgapxI4lMyGuEsixmjKR1ok4xiwONb3Ek+YtzJl
4HyhndLuYfTTzbk9tDOE61g2p5Do5GxgfNn8RPejrbD0nLzaC79LAVyXrI8cIWkO
o6GQMwmourzY7Fs3EZwor1nMwMi0d32Ilpvh4m1BGdQV/y5ut1G0BNFBLoAFCmb5
CEi4vHgy+vfAPgfXpBhygzzOG+5rf0BbzW6Gx0zqN/xOvZQyvb8uZSG1h8mpw25R
FZBf2CGXT0X8TCmhSS0PbpySkwhbrryVR1QyYkpMFOVtQYoyEaEQyp77hoKmpj1W
cUrGAOpdxDQvJFGKPvrZ3H2Pb0J19uPo7uTAcZfHtEV8lOM0ERHCxUR3FQ7hdxEc
QW6eSqi/U4iQybJ2Fb4Cj1aPvpUK1szotwLM0GHi4XSQc1hiFFs3oA5rb70ciPuP
16v78PIB+2E+LqLNjJ3NUie7qF88JSvyi3N+r0Ta+RdfGCxyXoBeNaLVP0SlEkIY
aBgVYDrpxsRb2JR1dh3LoodoyLxLzGm/UdgwVR7a5g2uZAh5m/Of8svI46TEu1yM
uII7YNEZnpHAl+IeX5icNF7fgnJs98ZAKWtg4tlq6sBzDVAr0E8oX5WXJWOU/CEJ
Gv+aOxHYV/pS2ZEko5G6/9Pti25j0PVf4ISm7SkivBFRuh8cHYe210KmE+jYY1+C
xzlh3XP7rwzEuJ+KMQZYRY7OupAWBF7i/JiHqSQgzo3sCV/IOlycaGOB+W6kJ/H3
9nkueuoEAIYosj7AJ4R3LHEBOUEQZJYQxyaAOFfyANu3zaF9Wy5FXmmro/h0+7o+
F+8N3q5nVUHMslrcd7sy0jyPzEGLUc1Xlwg9wlb7z4LpaDFpxOuV9sfduQgGCrmY
fyR7eBCYMzFoYJmOfT4SneatFnDObfdFfnK5/y/2t/GQ5s+ShFhFTdzTPkLQeT+i
OOGcykHP/SM1DhTKWTvfbUjKUUKkyPIscGon3igdTdh20bw8zM620iPTcSarz8bg
jOvt6n1WaQw4vOrYN2PAXzGrjXLELExIMJDPJl/WZ25YtPpw9OxJdwVmqqny4kJi
ObYzwJlV/ZxaFqE/LjBZ+HSrs4MqVsvrqoGWBNNjkQ/+yNPYhTrvoILs4ZEJ8EGV
9mqeCK0Dzi7QJ/FA8roDkhXtBE65oE/FHzXzA6MIkZ1fL1auTniiLt0OLSxE8ewY
hAgNN+QDCp1hY++ckAWGTU+G6HwYAblJRSX7AhZmi1CoLvqIEJwS8qjkBLa1pRoA
b0Ecr3Gf1RXKh4FKKCEtTrS3I3b01ffg0kI/AdOcdp/VxcXEmhU4nslgmecjNqul
SXzAVIYHGevBmPpL5c1vQVNC2evYrM5zUmWT5eXmKKfwWWh3S9IiCz+Psxn5pUBB
uWIFtP1CtTw6ruLu7tGSF3f//iRYETpdwnJNIlahUJ9T3fb2LUB5fqGAQNWFebGE
Kl/+cRz14m2+xqRz90cvJbBrGHZvq2BK6OkWs1plvit5GjN9wH3tcpHwKJabdRAa
TnudCUV91MCLyE13rRKPmFjWXQuw1MQ12UAo1cetRdxT+3QgUi1h80+NgTjJGPWi
vcFXof45sHyGk0nK1konbEoiQGrwG+8u7OXXpPcIsc268ZHvZJ8tZnMZ+pspaUVE
MkoDww5x1sRQGfbTahcXV2b1UOO2vlvfwIgbAzyrsVeh+NvJZ6asFueBlemVY1me
Pil6IxAqK+Bo8CZ4cXTKZ+cm3TjRGcM8scL9IYKrX1v7HWnZFOXus25RI4uajXNo
n4RoKzJl6KWVI0jYMg6nWWxERtOqE2BiHRtANksXEAiwUuAnkqAItOW0U3QDXIMa
BNRyp75Odl1sRZUguqqPxkgu1TdHo+cQdBsH+2/jzc1WQQTphdBbqViIbOPkc1JR
lYI/vLXsj6yLjJvEftdg/VnnabJXF7+VTmt1WuhjXEfdDL1+nHY7h/SCOqhRkaPO
u6phHnS4b7mOjtwb0GYGIFfY78+b11gSv7RibJqDlNKm//MYr7GUY1I7hdgP0GSL
pmKnyQXkN9B67XK7bfWKhjtO+3HW4c+vRs2lJ9vxV2IkDcdTvOH2tVPHPGtvYZ4u
dDrjPufU2ArCm5y2OnVaF2F1yyofbrrG4K/JSp8HlP9jUtjwiWICiR2rezZOHTdB
vcR4UoN4g1U2m9u4j5I9vTGntne0TU5Qz4RVWW/lSXvfVP8Tw7CujNnq4z+An1FQ
lM1AfS6NEdWsG8u8o81qgTLAyRmenI2s9v5GDYhxTdUsAP56f0UwTNvPizkZS5IG
3IlTVuBfpO3mfX3VDe68C1Jq6AcFhexm3qI0rikTQWdtxl0chCUTxQXQMwbZctEM
ZSqXWTqbbtQHY2dts+OlNhM9pP8FFgq8nO5sW86dNf689uZb4hirzU4AMy0AqpAE
hJagl7XFeb0HP3zQlvwRN57AKsTGXurdkhrZq+g5OQKQ+Gz+Q7I2z855rSA2sxU8
HCASH4awRd09USha4eiGDrZbOqomMo3ytYFveOS9CGSe0A3k5CtmmlB07Jjp8QDV
hpThB4CLisAfLCJwHZWF9bOL07dPuo5/4ndFsCFBXndwsJrw0FGmYrfL69C+dvgd
eK38mskq19ANX+5C+GpMby1bbWa5cqZK+aa+s7BSIMCDt3MPykaTZnEI84V8ioqn
u4cuLPhN/Fqe6Uim1WSSqgF9CVjF7cPsALw7odOMIlXUwKAf6HF8h/1gUeDQ5Ab1
gqAU7BDuk9411RUTtcFJG+Za2waazue87IqcptKP+bw8Hon0tDu2GnzqfpdSPD/+
oblkXelAT8v9VCfJEAxJe5heFKPbIVNlwHMtGQO3abZqcRMTeYxIzbQzhKwSmbrm
r60MDTiN+F+87LC3yyI8cTesupnce2YztnNzMyZAuZdTeb/KUSYgi+KYdIBUL0eH
lPEt7mJz5BzOjACTrrpk9cGNxLTZMjYYNK0hARv2Jyv8Vgs+VYvLIg0XYFH/2I1K
87ItKDLbZ8TyZKJPlaezaH/RscINx1s0qy9+tMVjNFKouZ5plnXuP/1OckCEKT1q
8fG1vmjgYisBASwHNr4TSvsY1oChX1rLdDFXlc84ufdZ3970rqaD5Ttb3W6CzZeP
CnqNObvExUR4/tkfOrEu2LTOrkjVttZfXazM8PeVaN3Um8QZ0DloHHlAUqks4NoF
7Hr4UNPytHABtU/y6A5ezSb7ern2ZRrcqgX6fH0Cxrmmp2iqNPvBtQJUhUAgPUlg
F+KuGfKfhItl2NoyB5dDjyOqAY047JTfu027xgsw+qITpPlYLW2ILVzHPSpyyAdJ
dr+KCYjNx6j6wt4NaTQmkG5X7LY4JOWRLdJXFKWfMhqjyOArodGh0bi8C6LaeoBh
hJCN4cyEAKg4fA8DbQontP6uAZTeOBe9SZETBqE+hUvHOUcpXWaS2ZEMhPqmaZOV
nkJBdEzqv167Hc56H+YzswQZ1FKLmXmt9qAePCedtFRVnjguL7guXImOCveIziXh
B44ltzIrN+2gLYYNCvYC5G4A1oJQBXlZEIC3jxqAAn1DV8xktViz1i1YqMbFZVjQ
9zMC0jT1zk6CmCfj5tmQSmdHUHBWBDzz3YPdOeLGs4g5YuDfExReNMohTbb2jAOl
8P1bwsmEkXqrHsAJPJWFCRdBjIgUrR6+8HFDxQG1K55XuKz1z/TOH8xiBodnq9ln
d1oNRh/ZN0jEDjv+OXL5fITldLWV4YU/A56uvdWPOumA7EEgoHtcOfp5X4oif0aC
eUK3a6LdgwqhwzSfdDHk5Nb77NSl7VEi+3j/S4bm6LBbKMSEMJIdUOg6gIf9Fy1e
DJP6Mms7m46sSeYj1H3N2RH2ZM5ETCC03LQ7NZeLqb85qeB/bLflHyRVlQpxxuU4
bG+yb5pUF34HD/nFemp4Sg4BydaosOZ3kGV292axDetag91dwO8iRk4NZx6iDRPz
QdyvOt/kkeZTtXSIBYJoDkr0h4exGlu3CRtVpkpgaUrBHkvpbxOvEMp6dWQwblFr
Uy9/Dxt5hWyQ46dW9LwgXfwueqkJUOtNtKUYZL0oUYD3/d5Lj+/Lv0O3KaXLrUxI
PLQ90u0Z48d0P8fjexVEkxjTXJk/CdFfiD4JlSarMZYbTy5kbeDYSaMiFGz5otAY
K3Q9XMkyeqL79S/VWCTNvj/l11M7P8J79UcRA8umtx2zOaUkjfi1F/2DgxmPZqlP
1mbi1AHN71UH+kcjw75hKR4zwQTmZVLDeJjF/+XQkcUM+avhlBG1GOKVb3OY1q8U
uDQCTGQyYetzhZDOs8k79RB7S4+luHjjqWcXRTgMfPVs4WODILZVi5t38J3UAik5
9ZkWC9J3sbxNbLfHiLydoH6rKY62cZoUK/4lKi7yCAN+MSwKkpEXs0H0fRxlHsdE
/qJjvAxFGVuvft1hyfmNb9ihK1s0fJ/D/ZQbQVCNa5UzyrrziAFvZh3I9wZsmRqL
MosGGbSFcX3hdtXJOeDvYzw/eKjXkSNBs5IoIH+ZUUt25DTepWhXlbKoXhM+Grgk
Lh/An9VECSDORpHpppO2tQN5uRmXFCv9xS9tv3NAXhUxuW4Lymninoi54AkSRSb9
pSIOuqXuVqznVWgI61ChS26A2lGnhWxweCuOkOrT2+gDYY0dRqZfKqO4Ue3QlEfk
prv9q1vCUlk7X/N/V6rbfah02t3aipBNlEW76oJXgcpxUcBW27viG4IWu8g4dDMF
PpH3HxgGN88xS42693xoMg70gCywce3kLMnvzSV5N4rpS4bU7yrOvmkWmbZjHGdO
mwbfczkzcZoOwl8abz6F27XsPkWwoXYc6/O+9VNJ1woEJ+hE9o7BXwEw6X/YmhSM
PaOEUPTOUQAy07CI5oEZ1azVokfd12c145BxqKyPsQ+a7k6t3s6+W8g/dgliF3Ml
FUrpFqqQ5Sx10g/Nc34+bj0Cr8eoMaNYVdXPOOwzz+6iZD4+L5AEM0wm27l+mdYn
Gd9HOGLlfX0Aw/XAHTbvDAPpFq9HdxjWw/bFgp7VlCesS9hgC5Lk8AL8Tbuo/SGQ
JrUaTbyiFNW0wMstsww5HworFDD2+//6euOyjvUiL/Cyz19GWv5MMAI3e5NdfGu2
ecLmyjzh4gwsKnF1GHPlNtXTfLpSiPKZKuxDkii8dHd5aWuStOX1j1CJGolOyQh2
k6H2M8bD4vSbOwMR0KqYnZwqCE7wqZ6CukbFpYO9PQQY3knN6XJHOApQkAebyvk0
GLDnxEmSyfaiCwNYYoKQD6rSIv04odW+1oky0BjVm09ppy0VqDPFkYDwy7iGA8LD
q5wrcDA7VTz9phgbg89U47w388y0kA+39gI2p2BInvA3URIemkq5KLQlaB+jzIht
k+NdhyWYlykUMrPIo7zVLkfGsvnPh3VtJ33r+d4LQqckMGLnmg9OLJSZsl93qC4K
f1FpbJYeW6sCsxDp9Qn9Zi0+G9npNHwwAU3T6N8ceOSUpSzIFP7lKLjCeb8wiPiR
P9lGAy8zDNlT22kcNnfMNNTyqxY6jl2rBnFdQjRFku4G/c0oeV9DcfFJcF2CAwc3
qNWofmN+oaSS2VXvnJ+wKCKQu8Y3PtP5w3C3BhRW/L/0JI4M1xYwVIVBfpALS2hg
iIT5qgVkz0FGQRj5HSDemSodRSTjCpt1Wy93FU98nxyeqXQPL+lRjDydUBlKl1uj
ZrMKrgNbE/GlD3zrqR7yiB2RiNlXr8wdpPyVxskuixtnnpAIPQGsceUFcHOHtUwI
BIGwSvR5z4ZODGd8YOFgKJRDx65HSv4n7OqMeW+PptmaDhwazFE5MkUg5Up5h0Lj
iIZKVd6vvIlWoVOIz4kwAk/7qtGIeipIJxg7Uk8d9I79pxcu2O31aJd0dFMyLdx0
BEQ9lXkgB+uq+J2mTHiy2qzkCyUOdfpC+jUhFBoDQhtrTzZQdWQYfNzbyJU4JGQC
nB/uq1C6N/dTEIpAt9CVDVmOeb9ZiYgHpG+wRH0O6/OIgh1C9uyB091rTSg3Z/cb
5xkHkTtX6VKQAN7BBQuR/al+sHYeFSlGq/W+FtEfRNK02QuMQovBtd9j7KzwaXva
b6VYNTr8KpCrUkPbspL6RMMMecVGSYRFUQaRBrkFc3TkWPShJOiPul3VDm/lxFRv
QCcwhn05qgG1omvOQI68dpRAnV8d+IceK0tCaOemicQ9HcO+VdqRwsY4PkBezIo1
7rrKF3t0XpYGYW5OHkR/rEe5OGcR6kzlDWKcErwBSZU+rpsB5PhVXmsoRQ/ZfWje
GhPAVKke5O3CJFdTUf7SnY3GVGNX2vYZErsIDzw90YqO8MBVuXGeqIWLHZ4kpXwE
s8Q9ktlR/0SW0NMfQSfQZueEbV2Ddsrcdya7Fe/6BBUtWG39VDt9+jwZWxlyFQmr
gtFOyl6aGnijD+ubpjFcTC8v+8VPk3Q0p9ZpbmkZUB/N+QZcQ5s6oOTY2Ig0lirZ
5J4i/QblaSccjcs2MUS/7EfAcQE6s/LapmVg2VE6sxsERgcpZrBwvlvnttipBHad
vheiaOpemGYoABSzCzAkInRg6ZfGvigxKnYKR3Z4C3QnAP4+23fnjuR77qdU1IWN
zy0sp9zQ2BW8yvcHMFrlXPHIlIAZgyzPMIwCIMSSWyOhJY5Boa7YQDUk8qnu1Jc2
K9oJhEjxT5VOAUEi9riEDELcn+M47CKhq3JqFEvkApmbiXHcI6h3WhQszzMaAYXf
y+lBoJWA7NdT9+vIKQ2zGAIytwbY3a4Ysn8HgwxekCb57LvMQi2Y6h4sV68AHi0N
743HCwF8CdrqgL2SysvSd8w17pMwHqT0+OY//5I5/ZjMVYnQPXlmFrGGs4kcfm+l
uMCouTii3/k/bR9fd2J1KDca5amwnBDG6piP+p3NJmPTDgPt6XEDn39I3GJKn+GY
HM/bTbhnc6UwWeOSubruCb8xjwSn7/YK9UcrZiH6BVp9+yeG45ubwGpm6vqzaH5O
qzJK0DgWqynDu24E2us+fqrKp0yOGbOamuEAX12/LfMRFHq+yLcvCOO5T5MnquDa
dAiad2FKh23yf5U+VVUFUKuwkHjRoW4L5/BVw2mDjBpz0xOXPzxaCLQtOYRQCgDj
nAQEwBoCjawEJLz63w+tvzmDRJIFxpjkVcoV1PztQEI7j9OEF+N6pYQbVhscY7Tg
+5j1m0OY7O6MpmOnAB96ShJLOedoqq9NWDM8Tt2e7N+lWIfAojV7mHRUjErE1yiA
W+kQyyPnXogO8VPQMCfOim5aTSXUol5Tbwc7FKQCp0l1SfmrlVo58XoZ0iP5goAA
zbbLZY5nrTrlKinHbIOSqotU0vsaQt2xTKXBvte0pE4Zwh5PkXW72VmUiGkacuH5
aE9Hw02anaLK7Cs8IvanjG5z9LuNkpgRVNZe9WirbfhHgciabKu+9Er3HHj5Bs1s
56TazhgPoWIAPAXHZ/Fugj8RtTM0ZlhWK1v7i53rnMyUmCBaM70GryhzLv6EmGQk
X2TqPHzYj/9u5CvLUCf2Qqf1Jb0Cw1NvFDaJlEidDAcYvTsL1zFNqI84LMuSFC4M
vrV/okSyfRu670ljlEUA2BQHDhnRzaAgb3w42nLoGKTTMzpcJywyApjUqCx1KUXF
Z+Eo/sdvn0hwCoaIOLuOYWYeNT2uhNQLWmVqLhiL07Si1PH9CTQKaNGdzPlReTXh
U/CacsRZZuyHWnsUVT1zVFZuaV5qtJrjMniRodsQdFxzgXkfJH+tQc5y+Hb8eirX
/0YP009ajsvL9TQqLh5PyDCt1CFVzE0bTv2AUKJ4rFJLIQYAKEgk3kcSAkvt67a2
tbc0fcfDDplotqPzrEKAzNnTqEJenIRzJjzzfjkbcMJOEFhaWaB/XNTeedPGPJov
TJoRHgb/+g4wEJMAun0XqBRrrdbESld8veExVg5d8DQ8SUYlbl3/U4j0H3N2phk+
KC5THDQFvwrPlPfPb3ejDH2O7XV35meFyoQCi7gYery5cl3JQwbGPc2DcMl9O6Yc
rW+aLaQoSZVJaURjLCrNeYcTa77kC43q9xjYlKqQPGCyHOr30rjl1dlc9UaAO0p2
XSo78r3XtGCNDLRi6aWeBxVmYYxQiOZ5xRM5ydPp90yuVQquIjvODQPvcBtaDw4p
afYYnJV0eN9uPOiOrqIel+K8w/s+KqxGW+wx+OV30OQuGs/EuTB1xge5uDLRHRYj
mKpq7vWq1vsLPNbzBz9MQpd4lyKcWvib6ZoPK+qC5S6oZ35WFBAN66yxu3qOUO2Z
hC674Zob8YMjc6FPeyLmg6m+zem8GLEawMzM8cWoEavLpy3rYFlm0IiJIteder46
XFsaqIsje5Pbod8BHFslWEaTM3+sJSGbvPeoI/B7VqMZ/3bqYxCDHE/8moUDR6bY
6sLxyfh1db6V+IoVS6f6s5Ee8jO+E0wNCejbGgWZ2sUnvjE2yaeeootws7JyufSq
QfugDlzUyNzpMUK/yYaKz8HMcypIWfbEXxfCvHqQbrJpw680ReP6Eqki9tYbxHG0
Oqmg6x9wLso/118y+M17oBPYi7NcxnexyqB9oaTPxxOWkwTDALn0hDa15BudUa2y
Eh/RowftQxl2oZ7RT0z4TJ0xhL/Hp+oL1ssmXDVVBZJ6l79Jjj5pcSfsScuq8wtp
7X71QnsuD5ITRJK8B/WzxkJpcnpZqhkJNBC0v6zQHwOwHwKxyajG+z0DvqvbWkGp
OOV4c5+lvP1EdSFXYJ4rQHWQNhdCo2GPOjfj0MrNcR7ER+18ROK5e1SK5Z8B6MFR
oo2t3hmPINafUwrIZ5Z6MW9yxY1p3e1UEUAFDeVsVj84i2vzH0zvQz0+8N/T7vhp
aJpMq07RFJWvyckusqzG/BonmZUjLLzg39RYdv29V5XyLezLhTr1ulk5zqbJe8iD
e4bfeGYqw8ILws3mEYSbLxAu3i2zLih/Z6sChZPregq9iZ2ugC/tXMYMsOKjWf+T
Infcw5LqkvmC/lc7tU5BVJ6vXavhdbjP4n2bYhKYKleYnHQzGQOc/vzaoszqmCaw
8Hp/WgcPv6TH+XhBgudnDnl2pUiGppWhnn66fNMGXvMbdinnGewqb6puAIxjLsbN
M0R3eKzwi9vko3cEMIuCwp4expRvU2uaetiEJ3qOl5SxVtWiSXn89SG/L/EWmINY
6l9xjG+iCW6RWUmbWk+8OJEbiHUQs6dFqwUjb/6Rbr8YrH06LOhZgYXV9amS9sSx
HBTz+j8Jjp1OIKfASeKV21pHVpRdFVAHsgr9KT1O8aI73l9UjqxhL9TfXRs/U091
lzYKeCAfrFZXWurcUmpsARunhZgiGALn5yitFIr938JI5vojX8/aIP2tLs7syQfg
PILDKMd3UqBSMu5tSYDAB6jOW5Dr0BBAL/IVSdOotq5J3K9MhOG+JwzgTOlYKbZL
bxupUSnsIQzL/z0mRjKu6bDZzV6YFWjKd/5oL29Ew6AeDHEw6ie607jPisXLKdax
c25a8TVP1uishnePBgYzsnSqpCA57lxFZmCegS0yyw8Y6Jgda8B6JdgLYy9x5uNJ
SSIsJybdby67IhUTYqcevmd9jlSkdUvNcmvoaSuwSa8q5VKPpHSqOvvisgQQPAQr
vvSR9I/RnwDJGQRth8WJ/6z94ZJa8MWoYLDHI80aByUjE47Jk87stLOTOfwn+i1N
xeRjeNfwixqXt7pfoEYUy4CI+aZD6l2NLX2WjL8IW9ZvBxsfpYSomevU2TAMF+mP
ze/8K2XdSJElkqHeimv4fj9s3kIBBCpxltrrCX+Qen7dE5XRFkJQBhM8LgXhfu0/
8xYUnDF7dfT1aaTLEmeeDv6SsbgNaEcq6/XoUu0cnUcJpb7SBrktYzTlWJZlfd/S
FLW39W+0vU31wfLjZyikdd4mLkNsWxNH3aWuF931rXagz8JkVbl3gbaZbiV1qxca
k6nCkDWNVFOc5iQrRZ5mp69QB+Ni//vXtjC2H0R1UM6XI4303PhP6z13xSFL0kAs
mPXTXLkzOTTiGfUk6uveuV1yY+VIWGllZMf0bCRbEMNRtvTDIIkTVqGMesnrFORS
hr+KZ8z2cSXBsDZA93uh8ayg5hz76kSwSP+ltu1kCHwJO9BIZuSfHQGZ9LRi9n6l
/XDnkfIpjzotOW0ejflGmHkufvrLuyvzhYbm/SDr1Zpm3mDeDPRSdfX2b1vP94Az
NUfMJfUjHsbzKzjoO445h5U+eaecSTb7P8Uo/GrtaNQ5+Ad/IwgpaQQwpldfD23B
YAgl+5AKTS27pH3ZY+ONTt7MBpVEPogY0wFQzVwZq2nGBBvE6s1s67LibW9JQ4zZ
zUEl2Ug7cINmLh0DjXoVbxEFxxMeKEtJ2Hu+702veFctfdsXpkyh+dYAFwGegO1s
pO1HTKcaJt4c/ypI2k7zpq9wNkcVtZsuceXOBbZSET3JaYdkWyUxuzOGpV6JRaAY
h1Aa0yMhcT/NqUaknb40/TUz56VW9EuxSyrigENVtMUPtxyk1CVEZdR68kgby/s9
jfFNZZiELNsk1Q9kiPWna4PvRIDqQXolqBzfscfdyJo=
`protect END_PROTECTED
