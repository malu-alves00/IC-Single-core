`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xf5oePakyFPZKFzBpMZOD0gLYoHc9aTWypd67j5w3Qho+TkGSkOb2IV8vBOxnGs6
wzXtlEOlDZf71E+f1n0W+tP7NBU9je/RbkhzKqrEdAzun6GFpRGbT0u+j1yHM4IQ
S/jMMLXn3z7eqah9I7OZU4oy3KuN7vFpd5sN3Qr7vzq/TX2Rmgwl6E6cyVKtRSml
aX7eMFXAyQPQPDbtCjxGgzUmbCD9eIFTxU0lRjfNjl+Sho6YdcqoXG9xxRP8yDH7
FOcVA5nkgDfZIeWCiRfIMK9k+2b/IZGTsMpnaAN+Ox3mA+hFLGYLF3NICTFjrl6a
NGXlc8wNLKrqncaNriAvia+veSwiMoVtIK/NzSeQUo/xAcHn/Yz6/5ppLGPnT1/O
5AnODPlcfo3c8ITvqhfw2jZS1PT1GtWwG107oDkrweoC2XATC5N7uktjsSlv1fY4
UCg7Ki9ZOBpZOQyCda9N964tjXvN24zMZzQQnD/9LM+/q/aCFExku2whT8oxkVWQ
JiBa1stNNxAGjt7/yvOKEWu7GJReTaJ1ulxjo4PkTWMLP+PVl17G7ymre3nY2Uow
IgUd+YMg2dGxbdFf4DNR9PL6CJOEH+MlHLyIbEmbTBO39WvRXYkZv+ZFGbLgaQy8
Gbj8A3IaHjZpC4GcAYvOdT7WRPSnGmpXlW5EzsiJmtSF7gqeNxnOkuDqaNVaiHm5
sm3lAfhZYVFOC2s4O1LR/IzOLTV2HUV8mRjpfyvb8unHuH11sd5mpV5m3//Y+seV
8/z8YKXEWNrRiee19igEo1+nVWCK8zc1SPOsfrMpraduCUvNwfrjiC3WGrM91WnF
RHVldoW4zhWs+Q9iFJ8JY8Vme9lAystKE/jbwGg/VJC4ZzQHseyRItEXMA5EXFgv
sRPLy1ACK3ACKKnUtXe+h+/MOrLLywq15cmE0IJD4KqlwYnp7n/hECUo5iXyFOHp
ga+73VCL8FQdr9i5LGIJFMDA/mFMi6Q/QiRd/UfTG6/YxuRMm/zh6Et+J1Euih8u
ecVnSIELs73lcgns5HqAGfBz7PQ+IVXhuZHyTA3hnGouq/ZO67zYkSUiKJf6Q7Af
EvaWoQkwo49Ee5Ev7AzhUvweCkY/+aI+HHZes1Bs0MxFrEiPJU98z0z0Q3lrNdAt
w9ioQjshJmQFfBuWNf8DdMlSQgt3nlrat2L6PbyI0al+rsWdi0m/XmPuFB0XRlaD
c0T9Ms4QaeNvqb+ZG9b9/KOTR00eCf6AsAI8v1D53tVTNUMFnBTc8vHWjtdzyAyR
7OcBRaa5ERKh7jM7galvi7mZ8Ztg0EGSQt5VaxSCrHje1jPdOgmGLbU6mIre2ZKL
WiFS4CFRIw9HkheDV+g6KNdUGzC0V+mKM4f+RejBaRvVp2S0IkfZIcFyRk0ApPuw
8+CIVRLXRfEmzRMaBFk4EmtbjeABLUTnycdLUzBT7mrufpPRHOIEofl9bfVtdBIh
8Is5msoojxej4FibFwP5wS7EGLl8DcFhI6YP1BPMRuEX1ARyo7lt7aT9QYQAouy2
sZJFxy/tIQXg4VDf9Zms1lqG+PaiGK60+vKScBg9rKhtQxn++wbaR790wQFjkRks
SZ1zM/D0fjjFMo5H7amnJwVR4XIYLzCKEDUi1f5lOZXIwKD7kev3Yer2vchxxjSL
Sn8FIMl98DkQz8xDElwvslXXJzUGFRWcX53lEf/Py2xinZCiwVtyy0UuN2tgNdBF
nRl6eddaZZPsl3RNBGvv7jCXRjbeznuVeDhhUiSXhmM3wU0urnCj4ekaMl51jqeQ
yYAK6tdbIFGlvCxEQt8KMVG6kuMIG8UC72liOmzDWLCa/vG2OtHdlqhn9tpPjCCL
O6GgWCeSCFZs1ZnOe6RBd8i/pdscR3IcA8FsdJyEdUjATdJOZACPyLFD+F8aishe
nonhQV9enVQB3Z90RNHZsQ==
`protect END_PROTECTED
