`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QBX8HFE017X7wGlyOracjNVENhM8lkIcSflJVmJ7TVYYtWwVXb3no+oCR1fBkg1L
QJxRDu4/HSl0szw8z09Mu2JOMG8MXSC+qHBKBPtIefJ8W978L2WgCGyk8C97VOvH
pJ95P/MWUFGuOnVzRZrcmHsDZMcg5rm4p/cYfoFk8b1eUSoGNdVYpWHV2bC4RzDu
A48VQEjpw7ljntkKBgmOPRh1rlSoeVveNJdBWb7ELVxivksZZKKCTfygQ0vD8+sx
FEwmZrJffQJy+dp1zy0J51P5/i7kbdB38gG2siOlmJnbOq3QEtFUsu4MK7Vq3eAU
m0UaB1o74kAcEP1o8keQM4qIhL58b5Z8koTlbXqK6wf3JAj5+NCoaWMWykmBNI6P
IrsyyF4PIOpbV7CI5u+YiIBWcgfd6sWz47uvSK9YE9av5vFp/D7AcxaZAuJsxQrX
g91CadLNiI9itoCrmNQZLx2l/zkTiusW7erTZY0pZLhE4Kwa/9Q0806OzaaxEZ6T
/oSI12kYx7ibj8/e3PJx9PrJ1g73rejamyJh0U6sMtPeGJCPtEt/LSE+/1vKFlJZ
dMMXJlkdf7Owahp4yLCZEMmyaiuuIueUXAT35CNgf0IU2Zm8UjW8JF+lJfxiAD5f
Jo8cvSGeA6juct9UNL8Sk74npwPcQZ62MobDDdSAbHeFEQ3NxrIqz1thTdyzjbvY
5l0O4IGQsY0rKvAzUysC1xSuFvoS/O1tdOzrIVJFg84vyeXj0pIoOFKy/OACqWBe
REVePMIcveSVgsOdahIMErTBjm9uzQOJ2y9W+alDr9vYsrbafo3T/20vBMoNsvaL
hoiwhCsA/aW2iDOEqRz9W0LCYsUmh2hbfIqwPzXIyzROi3wwWlnR7tEhIrCZsfZU
xAQeE/uc9pWHMdjof+Tus17JW+i9X0Om8SqXP4D3gjB+UlXM8L/b1g/WRKzhxxB3
Ibl2KGIIQ8OjSri49OZq22AeUiOuZFiXa4CwETNvzx+qksotjP8K976y+e1sIkVB
/r40yMVrfvSxPVpi1PcKE2oQI9GYsAj3QwCLodmA4W09lfoNbsDh10elza1y6gxv
95ITGfec0GDqB/qJ1w8sBm1KQUmSIrXcFlAdfBSAeMsvm5VtA7y8itt8RkvWeOIk
jVipUEziOKCVChjJL8tmudtMakDlwPKilMy1g9/bAvyvXp/jpYbEi7jb6AWCgBEy
sYjmrEs5kNHN3ZVTd/7mfFunWV9KpTIDMZSttnBaRkWGlkNNip5vO3DRT5zYbjWr
EBU3zPRdNMPhA9M0LyoTzMxML34/YDSiFE8ELVBJaF+iNQ+lCoFVC0ylyxus/A5p
5lpTZ9oPe1F1ix2wWegIvC5o0VqBlrvW9FRYmV5i3Uiqmbq5xMVMaQCKQZ66DWbR
HkqecRwFxSUB0b1fomV2fNyH4N+RuItmdo5BfqWKJg443aMZiVUJ45LRSpQxijD4
stHrxPl/q0iITHt0ZCIxOoEVYHZijN8lM20G8HFsQXY7zYF+bErp/se70lfGyNU+
OP2FQsuZ1ws3NvwtJF/0TSH966vMET3QTP5T7MhNe7sVxxB6XSVEYuRe1E1kcIHj
r9A64rtUPInoUY4EX9JgEVjeW04CBvORjbbIyIFlhSlPxQROGDaLDg7HruMOrrt/
f6Xii9qayGy/YisQUkTIDtmkmdn9ACKhO40CbvWGPMsEIioSmo5yxipOifwz8s8S
PPuRHY178iA2YnVs45O8mc/xCVhWTBHiAkIYQr85eY8Tr7yYPO6ZqbikBD2oHR2x
T4saDkwl+UnCnbOkQku1KX+QOP5gA4bQZ9aMcD2hMB+jpWSCR9y/OYe2zjs8enag
oTKBY47k7dWK9xn0xdBPLQwJ8fOCewGEKoYX+DrvHHVxU0ULQEaGH5T7x7/Y2BBz
wzl+tMQ4nvLsCUx2enaifT7NW1Iizww13AylMZA5jPaCgiQhrUDaWJrvHjjT/Upx
JiTYX2UxQ3u7L/doz0+HOkYig473BWCK0vGGAQSqcwoC9CPtrn2zGFZ02n/c5qaZ
m6OPOQpZh3Y5EBdFM5aCFLGVkz4DD6cS3kSOwIWqLOGU/K1cvE/+KbsNStQjvmG0
RcdA95+Z8e77aco922hT5UOKjHQyjmTCJOpBGo6wbh9CI8Iw13xzi0yU9/yFtKNs
NGufMy6nlUGPeBV/iDNij1a7tzFxRguyKYF4bupMA76K4eWfcxVy1wh3vk73uY7t
DTy1sBMRP3eyIBE1duMvUzMN7Njim1naes0xNHjaKZbHibK1Y28ZDYgRk+SQQaRJ
c9o19WYnzy6JstQu+CBAnIGTYJJ9vHEQ6kyX0YLdqNbvdtZvt+gCwnnM2oPaJ8Zc
IezxK5x+m5KEU1l7QQ+B9xKlQIX+eJQu3IdjTcSSrSdHfhoFjrc0v21/fa6BEmRX
Pt7O5m86sdlNizhn1Rk7LyBljd29Ehfi2y6nZyTRHBynhrYBY7ZX8SP3cHZ928jS
vSPFi9Lg8EpHqMoFYCFapHNtXp26tErXouLq97WT9mLOX4hrTL1+93r2Byc3CTKC
PPZND+2rET4NlRoqAgzFFmy84rxpScA4Ab3VDc12mvF+/gls7LmKmKed6/q317/G
5p0ST4jONjTi1HJZm7t9hVhCBtPNNj7ircHTph1WUVDTZHCzL4RAHXCN1AmRs6+W
0EBAac1e7SBL18zhKowhBY4nqt+ctHw/TfD1UsmOmEVqGaWlwpmM5awuIv2TPThT
+Sio3JPUd16wJGnnzQRSjufcti9CqWsKzGpGgf+Fvu3SXuWbgeeeUz/ESuspOYDQ
J6DxrTLJVX9/1Dfh/bxPEfh32Ejg2bJeVgMOOpvCCqahJVoHbOSs/vlrh1XWNG6H
h5uOi4toCq1Mw65hgZ1La984hxiVwNrtd73/wBKnt6JzRGJRxbtI/41DeVhMwP+D
rs3777Ty/sn4L61+UWEaVziMQg2rIPYMDUbbxT9yTXwmKAdcPu38UJm9ZS7BXQii
q0UNrLzdKSlTQuvM6XyY8anBMh45etrud9yXwU/PSIFzRzGyEojjgtNjlnO4fEiR
yuQFbHZTBtwjCMOu+/1YUp6uVil3V3JxkDlPn+COIwTcHjjmUcoCQqXH76QAsXns
oroZ3qE1SPaTx14eOVBU+qMaahznBWN2kkIDGZZ82W2KoFt84pukYIkdUU48wM2w
lwKGZdOiC39zuMDGaWRr3rr7/zETsj2ski/sziwfJ+b82jI4zxIcG7NFDUb6rBz4
eMkfAmwEmU9Fx6w45wyx4XZ0AOKbt6cpTSopFTBQHDGdljg3RTe9V4DvwVKiztYk
7/3yGIeFfMV/Dd0g4ORD/D/vm2cPmHVWdACW35gcI5axJ+qHQupDDQ2tY6EujcMQ
+UvYyh6pJkrZoZrIqh7DSCvszULlCxTuvCxXPHUagzLrbxkFSaCtyPwaCOQuR5lh
lyhjQRVtQYxnV8vbtEaX1SOM0zN0fPBTqgpC2NTrjZbIMNjoChU9asZbFirmRPHL
1r5OTYUE7iGOQkSmp5+HCGuLnWD5mW7WdwxP1zzCJw/is0wMMz3kXedKB1iJaBth
BJXx9sEujKVvyPH5wOUS5OCcUVUtaVDfMxXhKN0nYCwdTm48LgYpFFRWXqmGdC8+
bm1REvlGf98JQBkBwLWwK5Snm99jhnKD5ZGoT/PWc5BAYV0MBvAhvLymKv6fplFa
fjhUYr1Hv1VLm/B7YP/g6KE+gywKCZyxcdSQlDwWbrXuJeGMKMhKksecz4r3HSuG
o7R/wY/dkh9noL3lnT92V/lLDMwUEQo+zk5FICYi2t3G8RZpJThThOq/7h5fo1KB
MuriU+EquyGrFmcE6f7NWodddENeQXZJOuXx/B1ATgsuOWpercJVg9a58gspZXC/
HAIG7IldOKgFMkZRw3XFpFjH6RXWDbkJq7gAFdjPPEX6JdO0mGUohFE1PFtKfD4+
nclX23n89iGYc4GCrqNn09FhYfdyQzdsY8apxUPeV4Qy6BO96XI/5MUJxTVhLNkx
8Lmcbo51fyXNh/Pn22Adja89uxffDdzb7HEzXs1CcuWzTp4OP6Oj1RHwwzCnnRpH
LSn3xhFTYNMrUanuwwMviPmPbS3O7ra2kiopD0+cG52Mua798wwnJX3Xkfebqxul
+INVrBPz61ZKyp+/5f1F8NHeF0K37TDAEvkwFZMUZg8kNDhqejT7CVC6btsjQaoz
br+zhfv3kMX9JNqxdE22kbCQxJXUX/krJosnMrkdv3qCK+kkosTikcBPN1NjMDeQ
Pk+RobEdmuRr8ksmgLBHbaWK2u5GAxbPFS9ufS5CCtb5eg3cR8HLm/GCz/jpZTer
j9YSnuJHdm4MUrSDTbciPnurr6RMrAfxivPo9KScOBzd7V0h4DX2n4JBkCwIzrf3
aoLm/a4Jm+FdQMFvdmip3oy+swFlr2Z8oQpl4TQKOhngLGWEV8mqmKFs7y0zev89
XjltehNYBod1kSOWVl2kTCnCfq4aZEbDD9dbzRyBL2l6KU0hW5lTH4mRNsu9esJN
pe0ocjdYXltdg/zBnoHqvMXsvEf5uB4JNAQrLXhzTTSACJJm8vsBxoWVoPbnyj54
iKpz6WlE9+WzTwyT+OC9CA3FZU8ge5FNXiDfQNKrKi/f/bqqTqX/wyLniJ2K3pez
kppD1lM5Z9v79TbWG6M8hvChNbC63kMRgzC9fPNxMuCRumDgTv9wM1MgVwCl+or6
xwB9Lm7+sGhY0jhcmxcMoyj1ofGpgTbjgywWueQTtjuWdnAg8cLFyhaji2ASq7xa
JEZ5R8bE06E653EKliQY8faREhB2zr0HZmDKVse4LTs/3d3kXjVF/5uWmYeT8snc
VCVeJiFvqYiDkMChBBFM2wbV5I1/7+9kbpXUyyVgLCr32FXgSZYfTkddrTQDe6YX
iAnES+o0F36+GghbVRWRnZBsHcK0T2ORYP2/yyoqfBAzom+U2taBhjvUspJvCIXb
HYOatW8LsgjYKmkbUw1kI6/Tx3BbDFHJkeTbaNvgd9aBFTUbzkg8qiHsnkkA2USC
i3HUJJpW7ZubRxct/htnT25VoX0ZL5xXm7wt/RvQHt0omUxdVcfZ53yAWDCpCPG9
bjujXYCYX0LL7PYOqOWDtWLOrXos1DyGy3KLMA1MbP4Das2ntZHm8VQFnzOSceHZ
c8XDB3hGRyX1scfwD80kfF/n9D3Bd+R1GSFX4qyn1LR7Ip3fmLYp9ufZdVtZUzpy
1jl/UwHz6C2hBSnxvVQxrTfWd++ZILbCQi8hWQ3JcYJI1SiEf9U7lGXvfTFQpdON
5JCMLDmGcG5ORWv4x+6kLQYNKo7bC+pai/+H96QvmDYFxI3R7cTF7mxLU0XQw0Lh
Bgn0OPypr4XZe7f7166hulNUEGUEaDQbYn+ElY0QXgQk9RE+Hw0aoYRRSGphGpNd
K/SIRUenJ5SA13bxSXD3kLEErYrD3SSQqGnfywcTvOl4vbWulrE9L8duEOoEqgjT
TdZzWCBil76MteesfLmZ68Cv61+aseORcIMpiWA/AwjjlTBAuNt/z52N7Tr2v63m
A/3XuqWBQjsoIzGpaSMMCTcVu5UB4yRc0qR83E/gWMMwlx78V0QqzJ4aXzO7jDu+
QYzGDG8Iu8k1jyno44Drw34GZONp5MdCFe5+7fX/ZZZu7UNm73psK+G52CucURfy
qWUnWF2eBv/dD+YSDhmfwDB/cFQN34qZcdyaO6zNBXoSSILLOct/R5oaeYZSvWvK
4cEaKy5a5YMoj79S80hTZKWtQI5i+Eir+oCzzzoi32dYdlDMTelpVJp/FGoY4KgO
fRlYYvazltUWVfA6HuNtYVu00kM/DpDT9Y9/3qDmghYW9ChtxydBqeon8FxnAemL
woEeFHGKtysd0Gl/DasL/AG3ds1L77DLc49jvJ3FnaCrzRJ/tW4OoPE8EWA87luP
/U8hMguP1OLM695yHvcw2zAwlZZnmLEgLBnnV5mps/TxRPUg1MD+akBDZ11qOXbO
s1snJp800JJiuKnpg6i22irrGda8stEygW18INPfduhqzoT9f5G2SFPRbUD0uQnc
E5rdR8WKUkgDpZIgIDfr8ghSzK0NMFtlLt+UIEy/TrMFsIqkSQJhMbq5DFVd65pU
7uPcrPbPzy+sJDkW0hdfQnw0Fs6gtpew3do5OYexVpBNNOUmw+oEbu2Ax944HXuf
2CvwYODtRIzVn2kVIoIRXpPzybJKE+Qz3RKn20CpkesZvKlIGWCyKSEiiU9t83kR
aTQ6cfCazVA6ZjUmctRsJGe1ozU6Zh1vSWC3wtJX9CBqX1Yz7wK0YipKoeKb3WZF
AmxynC1Xj/A3b+BlWNLqJgEL2aLjnWI3dL2djTJOC4Es2R5mE0SA7YOfemQBldYm
jMQkat58/OiJWSQ0Ct1ILRYvaWqWvj00gzKxR/k9S0nlV4UKlO/lbGDALSdeasUS
rqcAcBXxKHS4HG4/XCPytu20T0Eq4dNHxFeXOAz6ZSc6LU9RKLHYB6bYXbLxOXjL
+Pju3xe2FX4GtGEKLsKvP3FcPb6mABBg0gzc7UEY7d06uiYKyWYBHH445skUpiw6
+Rb21SzWdpOeWEUlaobiM6oGkjWtEDmLmoSxwla96glOSbQrFYzngpo3UjRxZd9D
Ry1RF0zJ5d8Bnc9hk9xzaW7KblYCx6/7r8teJqLv4ZCeKNLK7FRG1RIezMeXrV0w
k0caB7zUoLjwS5otaqUabZJF3J+uG2KdRJNuntVuXExgA9uOpIhMd6p1u0koNDUR
PQ4BI/DWYeXeqJptdlsVSSDSyhgZRwxcKLrzKjD214MJCujqEHvTY0tnHTGvTddF
4/DweMALSGliYo2I1/dtc6grLz/9HzMBWWyZTtMvJdK9X8J23O+9dUVhP/Ms3F2k
idOQO9cx/OoWazMUIS5hU8DelV+/3D5HgtrrS6wyq84nvjdNbCX4uGdl/dUPS54g
pVoJTboRQEFkTIJ6s4ot9t6zY/EaRc72delje/PAjLCoi8YWZzpY6pQgXpsgccsU
qT/VCzLJdWjmBA0A260PW+bc8+jJVdZXAtvmQ9H5XShyab7jZmwzvsbd47dMeQzI
30jBc/M5Q1fp3X5Xin2xKAuM6z6YfeNCQSI/oLr+OeVKzC33KTLlw7ws5PrysMHR
uIb33B0Yg9PhRbubs0CF2sYnwRSXVlYlTvioYmkDP9EUWu1a6svf481it3Hd84aO
7k8B/HapsUrW3dqmPGiSQylMD0BPnVgNiGDCZ0LC5QYT2G7bOFfs2L820V4m3LD2
Oz00CH2s3w5wE6u1M3CVznOSFyhVT6vvKmD086mXpTL8bPen+A7tc01dINak9KNh
rKzIhUoIBOZIacsZkZV4h0rx0lq8tR3IRo5L3JD6tL3RQyeUelO9+zcZBOVChA/3
NRVCpYcwH2ySR6rSW1QUWk86ga3XI4Mmt81LNn8BLqPZWZtM6pMHpLfVNZInrhcI
cwrKRDuuw95Mm1F4BPalvK3cvnHf1w5oY2DWwBRXlx93IzyowyL2kPYD0JFjk7d7
QtEM1Z4En3u+Vv84mLYna55sYtEqpouGQapEOz8RN8+NKq6lr/5Mi9/F0zx/oXXK
bc63EYsPwcqncdVkDcvRqjKNXW55776m9X+3P8FrZi6hWwF1ohsLfWA4RgRa4R9L
yf2ZZRNt9xnBj631NpP03PTdyI7Ortvsp5li9SWk2uXduUcMCJYl4ENE0AHqdime
SrHGWwxmee9yKeSLWELhOvOqlIgthGszqutxzrqn2q2dKmz2SewsyrDapbqOSy71
faJmCVvORAxYxBYC4BZYwN0LqJKFerAM9Lr1TTCyjK9N9ZmMcjEdrgmggtIHO6ei
JcSgSqTIX1Nf7OWejGrxpIPUZ2rsrgJrLEV45ruWlftCtpXviSENvAWlYRJYn2pg
h/Ww6Ufmqfj1hGe9eg+xuBHiU2H+dDlBC7KNw2guAtwhuI8yEaJSbECk6jaNOvyA
g1SHB1zbMPRDXSirg5Uf65cL4xFIShxkuzO7pawdz5paBLcUDV9z1frV7xxpvyBL
nWgrkyYfV7WmeGDOEjc5YngzOkr0u80SRJemP/X5C0bxTGxImrbAEc1I2z9idRDs
JvSWFS95BtxPrGak18uATueyQZYQUDP6YBvrnf+dh71tQWIkhgz3c0wfH0zIJeQU
NxkWo8AMR2ZA8qjuXQbT6qHnbRnIEIgKlzqfVV6S6DECHN1fnidi+pPFTciTf1w+
Ds6npnITyxQ8Je4assqM7A3nCAGqKpnSlXmILCCLw9L3NgRSOY7zlQQCr4cDiJ0o
YJQFe98Oy60h7h2B0VlPgnXkG5Xah09CswSrd0vuPxyTE1IneO2wIntsqPtaNqe3
TM0MCu/+AEt+FVAS5wsoiYi1A2c6LsU5XCevGkPARzg2tRqDirkVSfEYPpptcorj
PvhFOYa42owCb6CBTlnkcpDfaBrU8MxAK2JyUQEbrTH3Koh/3pdSc3GD4cY/8b+L
kWxMJ81U90cxztd8QKweXI1kA//7iLpZ3/DARzbrz+ESjb+2GRBXYt4cZMcflH2X
v2g7e5INrN9F02zp4iEwEPaNivSum+oRKCQBFnJdUcuqjl/tBfIkwWx7kSbvk9gi
ckUbUK5YzUq7s4eJUIbz4xfdAOXPnTGJSlm/ziDDCvk5X7sgF6voeCfgb5VNSUi6
1wjfjRY09OkNU/r3lKIgwdeHf1xxZidZgDyWjtlPtrV/Su2onut5OnfqNUzHNIsi
X2rgziLHyKFtb8DUJs2cwL/ekoWeRPB9W4le0HpbsdyzjJAr5UTDnD/z0odw0dck
tY0QQyGFfOBRk4rFvhf0jkzUWD9/Rq7Sz5zdtOQpq7rRxut9whOJgCb6Njeo4K58
Trz+NMHB8vZyhmj7hrwuYsqxbAPx0irxuM91j7A67A30UnprKTaITCbEx5jkisOo
yScEMd7j6+NgAWXiN20Wa+3A4VDHqEZDS5UNTfhsTGy7cl7nWe9gmy8Yc55dWT18
cYA8zo/M85nb65/bonFDMxCiU+jhzCmwbgJwbGiNQmuRMU4iOP/KeSX/2Gc80Qow
u2XWb8SHkKAcsHYwpaWdtpMlenRKmXIei7YZ/jH5kQSxEqJyHNqdVE1CPrSSPRG8
0Z8Qpr3Kmhcpy5LxFNYrmXBkdGXA2iAXIbgi5zvyR947D2x962lG9a0tZf+sWvlc
7LNJOT3wtTraqqpe612NFcgg9zfDYCFjgDjgz3HYfJC9Cm3mv64B8v16eBnihsCo
YDZvtvBfP+C0y0csvdqD28MCca/FqFKmeyt2r3GNrJnSAMdSZR4Nk0f1iFuEu0iC
p4NDXoaqwmwo0e3BG40GmZoPoiN3PRj+E2ZL+LLPq+cU7YacRU0aNK2MNvliDwbV
0m47yV9f8Dd/nwoOBQ61Am1NIBtIECz/PAAWUMZl2bkDZcVGQsJq3u/NHdaBy1h3
S1GHjgId69JuAfgnu/KTdbrv0zE1IzGFJ2eShaJcCI9q88YXl1AVQRAYMHzKB5tp
05NeSAew+wbmdw4XtlONA4SxBJU51dC1wrHt/Kgm/tHquV4W5UW5EaiRD353Bo0J
Jh3FGZmLZj1U50pgaWjqYPDZDTGPTbJyz/81/BgHllfyIZKcOhKtqCE3H4/m1xaS
RBrvhkVmeqffsr4jUs/uMk3edamomy/xgAiIVf2x27R5dhe7mKRqv6UtBqA9TEd0
JO7WtlIT2abcED2oWl8lqjVpdTiXhCtjzapBPfvDIfKt6fahXwamFsOhxp7BS+AZ
nj//FrYOYNzlTMPtd5lN0vLRCxdSQo9gBXUokWN8Bl/yZm3ED3q++nq4CWsECACe
6EBf3mQYnbt2hV1zkvQ5okLVyQdsWALzuby3mXsLmhTHsHZ1dm70GPvNK3hZSjz6
m36CFcqLU1UbOIShvfQ/Oc4Res/1NX1XFGVNm3SsQeXJIf4UtMZKwxndF5/H3v+r
9Z2/XaF6L8hvFaZhzHSrzYwa147zKSRwKSMoUof0NfapgT0KXjKDJOWv3s06O13l
CInoRQxkZZZ3OCYtu74I8IeHArE3SqGIIRD8uz9owegxCWev9BQq7FKp9TwE6p3O
tmhdIcUh7kBcwN9hYC6KspfoN+T07MippqWyB7H3CvucqBHaq4tvpyxm9sCglgmz
SHaL7LpgixekiXPuEmc5IeD3GCPAHr9txg2mFjfVGWZeT8tsSO3expiCkGR1e7Oe
oR4sNeh6IGQGsDHoH4oSJ9ZXM3guBw1oMeOVlM0VRGkmbf62A/m8bwvcJs9GoGxl
W3cNevgxrxQcwovOkT2MqL+xwus8VUIcRr3cOKYlfJmnttU6o7cFOQwFW7/HGBmm
tNCEPb6TVK0t15T685MXmR4DRUsbuj5MxVlQL7e0vR6+ibn4B1CkGO5d3c5ubuAU
B41sH5xy0tJBe1nCKLZAH278XDZYTMzUoghBkq9j6qNV9J3dbrvjUDpgH9AybjwJ
ikydcxgZumR7GJuuSGvg8ApGQF17yaeINE+vA/mIUCjv3ecOUU/mYWqwQhwIqYcq
J9VtfO4RCXbaEGP2csKc9AuxdKhJ7s0T/K869G8oE9W5kUhFdFGMvwQbv4rELG03
8XSP35vo0+P/bS8S4wN4iflMDrte0MOjBtmp1OdDbxKFODJpwpk8voCEik1IJ1JG
NYMa0lWFreW7LJTYKEAB1iRs3w9ZZ7dYVA/CT0sh+XJBT98QBsi3k4LBqUp3hoGx
hWJpDMnvUWgextUOTLNuDopSd9K19hSueOfNQxH5Wx7FBwffirWQSmiKXsRc2lsP
zmqREiJ647yK5X9Uerw78HSWi/FcSa00lXVX8cwKFx6nRAKcZ5QxyjXUzjCn/Af+
+iV5jjXCTZIgBrLTkxwj5PHuwcQAkOJRxgEeLoQvfZhG4+jlC5W/hoNZpmpKRBhd
TgHCkQsKRKChLRg14kOnOPM3l6Dc/zJeqJqC/Usl9T6KLNiMZ7lOEvdeOkwZlwUe
o5twkXrrtGFF164Z1yQyViaoGWZye/CUMu/IpvUiaz5ZAI87vk9bWi03JTUYlYVw
O8jUKHYgSHm/8lV6HMxiDuMQUUrYH1iD7HrGPqPDBEDu25v6dTAal/PtKfAG+0yw
TJTjMpxAk7QtIsSusCFL03na9R3kSLrsN1V4tiA62CDpwpr68lQSi9cTdFWOQqD7
5XrPZ89A0Z/fOu38anO5evCDn+9vJcZqdh6Yf7yFLNFWCU43+ePWcTUI4vnABTeu
yau5+rTXHNbs9ahxFL+vef4ZiSwysM6IiZetu9RtVid6bhCln9A4j+Hj/hwIQ4mx
iWVj6t+pHMm+OsyI0JvGVonKcp5UJjm4od0s4Fi8dVFFV+Y57DnpemVKUP8/Z/0j
jsBwh9cpr5LK3jpdEYcQrtSiBFHKT8X6QoKWzx0r01C472G6ipAs2Z+kxhspxyWW
TygtJ6oN2t3nWXGONOrZFF1hD2aLwbZUPycmZwn2tf3ZBK120W6jqxgBWTtmEKjr
ugL6UogMkMyl6Vt4wCDxH9ckDkbA13+jLrLeBWvDv89HWT+YIvrUXm+VTvqkyLm3
75q/PvIX5w8IJaIvsejGObeZh9e9ppkJkT8LlvBOgmeWa3xSunQ0QZieXB3a9bf+
4ypjNOqZGM3nd7mSUrJ2KWNwyqSfeZRpzVaEDng/bu7S/ERHbW7Q7YA8cTSEFvrW
PgpGBtVypt1cWLVA7PRMmFLpu+lMh7x59Pp7xdmgsd4Co+nq4Mp8U08xu5/vgocC
sPKy/lyu8cbRH/TTbJc8Sps6Fv98m07My7sy6c/zr8mQNjfoEi2wKFn+47a42ogR
2ndP3cnbqlpm1xRb5LdxxoVseV5BqJ9ouTRCjNA5AkCG+ggJRu05FKkscVFE5fAH
w5opgBFNG1iqIGhuec9D+u8semcIUKQaXKBhayFqjBiqXPHBENEDu5/OrrTyYKhl
BJVC+z/XPBpA2HNVa8UJ5nJ76tG4sg11kU2+RRBuTqwHDt+TFhm+XLkl7ixmlwb6
lXYyQfxeijj8ns8ll+sUiuZBQVwun+ShqoKAYESEHApfx41vPr1jtOQdLhHlCaft
4N3u8MpG7L+0NfdfksTwxW+pV+MP2FyJTJr7brIsZGWTcKdXKxT4lDjs+WAOEzKc
1oh8l7silf4+cldKJRs4h1YXddh6T0wZVnT+berhZm1ejG4n0hHtZ4qmSbmUXzQY
0wWM934mzpx/sgegd3avI+sL0VJtDyyYwdzGd7LdIOcOzr87jUWs1cCzGEe7l1ZC
Xr+nQILDSDKFPrg/H2IjVbEm18CRGiysGi7/mCmK9x+BibKrTexKybbKcy5yg8I3
n1dP8614OU8qjERcsHkbyzrzBWpPTmSzxVibzs8w0PyULK35a3XdlrIJLxbecgAo
hZ1seNPMLXrbZVVhZ673FAeK1AEn2BdVHAnKiU8jILpj5vs/wFSAFQ/zkCAITEYB
/LOCwY++74P/6Tklpi2igCnr1wcHrHg8+mNRghMHnUqTA6Txnci+gpb5xqid6nj1
85Ica5sL+rrZ2simeyUKluUB3+Fmp8qTLQFYqfN7j8VteQ3F5c6cYb6WAGFUGJFN
zce7bVv7JzDE9FkcX96m5jcO5h0X2Rfht7QZMlKtPPN8WRY4Zh6pFx1UEQk4aS7K
4fxZHFOMURDzNN8Kf8Jwu8W2wbNB0KJYFwLQUpwoakr6TQz3QCbgBpIf+xQ+5BfI
ClcnQcEt5d/CWpyecJ3hCOw5cgoGxV0dUbvP0OoV3LHCL0WM1tq2DSSAZf2steIF
aklKPDeJQY4CdBgvQokNnMAScJ7ALSiWr+uziwM0U/kmpUrfHdZgOknDgbThiYlR
eJZ/k63Qu5LaNqPscIatEMFPL9LwLQJImSwHQFJCDzZ+x0NN8mGWT40URPtLE+mU
pb/p+e2QvrlLmz95ODr1VPB3wGPPah/ZLlH/0SpiHZmMVivkFtrf4S8+7LZZc4Wh
/e09fQx5biwngUIzrMrfr1vkSMk79/zKZqBnZW24qKTFF1HADFGTEZsXtkJz/Rob
oGkC3iOG6dyUmycAGdXuMTx6T4e3UyKJmuEThGYz2mSq+I60cQnMMfIGEiwEjFFm
N8p2QLeDIPLgANTGXsBG/qHq5gIWMDwOAR4SewtJA5RwCxT1YKIw6lw12a1KrQLp
Dq5AcWNm6NYiGqjP5p7PSfiS1OziLUUuAMTqaG4ZBw43x0i9aIyVS+CLufYKCgfq
ZLGnKpTsUp615RC8FdIOfNBgSrWY5h/qBPhyrfIewYF696oCCP3BHvHh5sK4a9OE
0QFl4t/ImGrhExBD4Vaz5ErdTsJnTq3mujodAbUFyOIS166r7JI7RrEmCa/OUTfK
61l12YQIXbB5qdtQGqx5aGrmKjfAdB2yKFCnJVRVb+4D0BOG0CiIdCiSgShPODwH
rt4IBAy0HIQHnTfUq1Fq98KEZM4w6MLvsruDTY9/JKgJeJ9e8jCQ3RbXZbOiK3Vj
afnS07aFzfc8Za6Vipt7mKM6Kyipm1z4Sws9SnsRhabndmIBSaHkuWS5u/+CPWmg
tjdP/gLXevQjEnqCtaWmzFTHZkDMd+AfG+csIebUie/DDWbh3UIzn6H0ADyDfGsB
+JaWU0T//SAxNucXZ93SBldgokq6DZ4yc+j9pATvl2fTKtRtu2J1N2Jl9enfGI8b
we6j2aPmMOEw6XNRQjyD0XyWbKvpbmFKtN9baG+lJTA3eAm/twiVIPbXfQZDGQOG
nr42XUpAqC1qot3fr7ZVSqnhSRihmc16lfGwu8XRe5dB7DeioiFAiL44FCsDLMLf
Yin0kA6N2qmtEcNsGD94Rb+/UJlq8Utm6iqrde9n4/9boKcpmvBI0gLiQndsOD57
rQKIc3YJm/oD+qnhfpNQoRgZIYBISwgMFGXBvT4LoUx3IZyf3xPPbeZEPBrIgQDD
JLW7oWwzdH08f1Btk+TqcRiuHSXCx6Q+9eCWNCafbYuhZAWr7LDo/418dO7UVAZG
JxWCAWEhycYga679EObmG9FoRaGfMKXo49ypLUMp1JKM62wsA8PBKH+wwKHs7oTQ
e7q3Ef04rP7akC9pvCn0wWqnCOcpf61YWWCD1DDsg1PEYUUWAyWKorFglv728DwP
unRl/CpafYpVUvXBSBu4gTZ9E6dc5QcbMn3SZE41EsoQR86ynK8ZpRfeuICyfEG8
1lHM/UOO2PS1gPT68CsyFFzgCECWp5+pQ/HTQjCGciFfU6PzBsmn81NSylXWMjj4
UxEsImTtgXuIxl4K15hLPJwzzESRsb5CoDlB5FJm3o++EnGX2Z7GOaJr1zdmeDva
P2knwuirHJyTpg2pUc8NeniHi5wlt43N2XKyQPUdDxOZ4nV74WaQZ5HTqrfQ0xfn
XlE+HU1cniasWVtrJ65CLn3uKhwv2/eNroNGGJVO2/FgFSuqRst8Fs1/BlTZUKfZ
Rir1/o+6/3Du6qcXzy+c1mvMZbfHTWzJqSAZaFC9OF1PXO0U+sVyKpbkB/6z2JVq
zhG7yNuJTo2ILvtzK57n9Q+UIDD7qi+KRY/hI8RvWlHTC/+GXI6AGm7a31fubiPv
31EKyInLjTRwMSd1p1PgRU2wbeEI15oOvh0xkcrn1T3L2D1iG2WzMGuE8nMTXM/p
ABkVyh8p4aobm1AP7I3n2wNIViUTADcIOVS1YJY2hvpWDEv70lWdCpaDurm+NsJq
GgW+49FGl4cLsmv5yYsSHsjGX79uGIaNFcMPiOYG6wM3DKygURw9qblhI247AXu3
HbdmLzerVMVYz9+z7qG9JVxYCYoihNLX+isEGTOOSUA5jYOAfsTfepA66Wukws1L
rYY0Ds8wqB66cFLK3utIkU668ayhLeegX9fO834FuAFRB6PzclgiwM/n/OBKRHXN
fgCWxdsTc4Yyk5ubW4VAly6h0sh1NasN1ZAbra6UBDqettvvSMbca1dDUBcgmyRP
gE2ZhO9tZMlxRDaIrc8RzMmmKLj3GpUXEnNGD+BHYde30EYwKvQTt06O/2rYSHe7
2ApRYQlC8+HtRnetpLZ6+q2er6E10Ag3dn1KkRV9s/z1Web/SwnnjdqKGSMyxXT5
1gykfYxhuuXx9lVngG1wL4zeC0gsv/8oIrAecpbgqXmXzqXO7BcubjNPPHUrirCE
RqNQ+22ED3pC9M/QUqiooVjd9MfA8GIvHpb/14W/06wmt1d+bRXhdsscu8OLAoZA
c+5um/IxRRvIer/RAHBU+6RXFEmygNY/e2v0BwXhGun6WjRN56qtlO3RobTEzfDW
YRtY6zlhKfsnB+0zdUGpKwbxlfPzv6g9JQzOZWFXRd/Hw5tD1tOp2qsCps03hCaQ
RqlGAOuBPH5YWzNyDcIUvAqdpTpf+6eHWci8aVu95ei70Kwj1BRK0PXWLtqCG51B
6IQa/CUZcna8+qlt1BxoJN3uGvHhJpKCbq8czd+3+DZ0CB7K28MmWVvAbmAfdvVl
dnXP+ljNTfim9PgoeUDuaY15Lcj4qyOQaSY9CHdoZ2p8X91h6JnSoUye51OsSreW
jzCHUdnrk7COAHqwFYHgx3mJ80LszD5CpdqiPjVkuqpucQJm7mfr7AndbHw+bihX
2Zq10LjpXGnpaaEEouZ0Et7P1KF/J1pYp6rlWkAUB/gV3F3qUcG70vz0AnzLRTkG
QS2IgrG+tf1DHDCDOgQbcJmEvMGVhRKfYbA7h8iVpgMHYyNw+WcB23fguCgYLUjL
Bs6R7+0eh+NjaAVAzMjQcrdujx0rzUxfYIGB1dFa41yDGM2e2a5oZ/Js3RPMjyDl
aCYqeWpmtzlD+EeuhrOzt7k5jtHNgNxA27mLwITskHOO8gqB5ek6Cnq96mooZAi9
469pai/2R9v+43VCF/M3uPsCrqMSLpCeyEojRhD95+HgaG8qPXdxmKLByQzAzowu
1ecbcTgmVZ301AgyS+IV1VkK/sWyX28e73kCs/Xkf55d0Y6/krLjHiYwCisLjYmW
wXaQG5COtZD/cDKaEkAFxilTm34Lds80alt60D9m8CEe6sdEVDD5PPzEX8DYVXfj
ZeCvT5bgvBvqX0bCyYjFTDhcZBudpagAZFVmNwk42aOMTYSU6IgKYvovf79XhA80
7pYzdENQqJ51utCypSrBXzSMysydzW+Nu9M8Z3C/DgcLjLvJtdDPRhdpnGb8jX7/
nIvJn/uCFHutAcIzWtvLu9sxxj4cLlxkFaWsKjWJpnFup6LL7SeUAOKe5hfid2hY
xPgzwsHsZtUba9XGIhOCpZI2LSUPdqqCPvA0RAl2PdCI3pr0JbI6IP9FT+vFDxMm
nOpjCh9yrCi5XMEf5z5nKGGMyhse4DQU1ISuokvAPWUW8lWRrdw113/+ObspsbNy
kS1DstOCOBQ1KkQ66Rv4/tMKq9yrxFxCxJCVCt88dWFUE03M0lyYYHCkPwv8PONF
HDWGxZGY4WeiWNy/S8rvt/gdhwd+Xb/Z7+mWptqed1eq9VyOADwR0O0gKFwO7U/a
+PayBpVrWgtAzf6pymKOUDqUTdeaJE4/pxG54KIT6KiqvWrzHvxnVkO2vENGl809
+DBhhOqeAWN8ZDOzX4FOKPpJIPAcpWp0Rw2tKwKe3ryKcp48gIX8ir4Dm0lpAm2X
mspJb+3272/E7FF0r5fVTHbroZPV9+6/35uCmwCMBBeO9Ga5cl/MZVTuNaPpNTHs
RobDByDmr2OzD71WpEyM1v72+xbl2+oC5K7zyzhgSNfp1+XrpEE53DaBgGugLGp4
zV/ETyIv2ny1hIKIpjx/McdLOlPUZVPa21M3dwq7br2tktnR1IrPAGvXg6r4sjuA
TwgXrHsYAdEKemCX27P/LPelWXjwRq53iEUkJcnP59/sSDf+MqiUAA9guXswEe+T
4Ms073C8oRkSblQ0W5aVWi5Y/ZZ8weNWJANlDcduN5Y93bBDFxjKSTnVgdoZIGRF
pjHjVWh49bstKYjG9+54Xnc0v1vp+tlp7LgJc/48PRqdiQqlQfcJVEDR+i3WkVJi
CijkWog7A0Ej+rVWlhrmCKqBaqitx3Z6bkQnegxK/XbmKbowjZtJ/gfQKMmQOuZA
UUk4hmU+GVMW6JEPCawfUhNjjZ33u9ygRq3ogvOGyQlPUk1et5fz3tlFCltQMEv8
JXGnyiGwWRsDAA4btDXL0dI1rH0D4EpyBc+C/1DbcijPwnnCynaDUWawsty/7mOA
GgC+gXUqq8kkhHxj+7hXO1/DzwPpdzunlHCFjCcuqhvB1vlu7YbdqsPwByeqExb2
QskDrGD+kRiVBsb40CWnC9/6CE12mVahPl7kYn871cRUKLt7/6NTeYLMlKCpmBLp
OIVmap1GF1l2PdXZvHF34hX4czNx/lqXDdtOwEEj13QRS9/oY/DutG7ppluUoHFG
nn/7warQeHZBcbSyfX7rFwdqvo/G5ZEsLL4Pb8bi266zwm4CanFqDcKan9T9IeAS
MLdd2fpWNsk7M3I1sAHRhWhctPBnf17c5roH0f3mxZ0HEe3Kly3q2eeGYRxi1yhN
h0uLEweSggo8E6fDOupxC9z5glWSRSIb62hTr+Tb1R6Ji+Qy6PjaUi/wStB1t78H
o/t7uGGCap3r6Lvmx8IC9E98+zSoRB4MHIRIQRV43asE/Yt8mJf2pxnXLZNVRSs/
jPMz2bV9/j3K6voSh/77Zr6uf3AXD/w5R1zKyVUtuO+QszuYKniX07qZ6MUif/8L
afBdtRlXqyH8zn/u35/01/7byn+pwNhasjO3xpKsuAFkMLS8UWxLTUEsRzHkuCIR
uv++9oIVUkJXn83d7woSPi0Oaev/crQgE6CkDD9l5Vn8N5KmqNMC9FvCN11q3fe4
2gw++Oe6dprq85X8YxhCvtBv2A+gDMslrbBq1LX7N4klBPcJeeSOdEvEncpgMAoZ
hTDhBnEn6a6PAAfaKVj+w7XX20FaWhgeY3Yw0YjgJy2+ZNDdy1Iex62oX9iD2c/n
iVdSRtl8Usvh8HUTd45X37qLNacxTD7XSvwjJ7Jhp6Eo0sIopTSHtTsyq3iWhZSv
dgSXx4e+/abYt2+aznDmt5G9K4g8FaN99cZC6YLKcq2BUiqrUxgMkbggWOldWixM
cmIafxLpCOV7aulM02zf8YAvL3pZsK+H0Hjdut0zjE3SzNdU9NXgNvdsjruyvo65
iutAVAqIT0+MobC3B5NUxL6VdXQr8ZoKrJigbeyR3zp3o91wsEuucGf1rxLvk+hz
eh49irlC2iis1WXwqQUSGVovoYdTnjELPBNFYI+bT/tA9onttc5t3ryakA4y5nDD
DZTv/k50qaCav4Ih9Mv6aVqAcntH/uTy2EnNSeZCsM1Tb0udYPomoD8oJRkXpuUg
94RaJrdZdshK8IXEdhHxB2tfcAQvlWaLO1swojYd06Kp3uAiwyfC78b7d+jb7b0k
sS/iuucwrPmgqO8kNTeyZ3YDMW9Y91mpadKMPCCaDEz/ULnIGjeEUWRhWzyKgdwA
ZurjuD/DDtsy15UNih542EZ51Jpa0GnrikhVXGh9KNaESIqEtK/+DJR//U7okEm+
Y2mpCagziNKxmxo4efAV96sW9q9wlysYv9pvITrLtM2ov58pzHDFSAmcb/R1OFS2
dwgDKALYXMz5K34tp2RMwcx0gYojTkJ2k5c+Z+vG4MLoAGA/5BIX+qusUYK8md5o
6FhjB1POva9QS4tIgXabIZk5ON8MaHKcf5yJuUDy+Dt55gXBCiJKo7loZoVek6eY
40xYJQE3qF6+i8FewsQWSLnaKfVxFbayDZ2EGQbtOhXLcfqspxXgRkqC8wUeX/30
AZ403V9uIvKfkYT4xTcU/h3dKRXOufLISVixS5CMBbnkObM5XrLWpZALSQTbui9N
yfBBicv/4Y/nRIMaREXDMvhXakI3x5hYfyUxkFxPjcTz3nAzoZDNy62q+n7vCTxm
8FG/yBjlBTh/nS5yGztqwXBLyYtjuNYhQwltoFjJKmBuMNL0rsBmcy2eM5UVtz1l
vMVIqc0sM7ZdvJTEw+dqxcqBeq8WWlaplxkeDRHbKaIlq1bfFiCYN1lxV7cVl6IM
dJ7rnwG+Wv2jUgPtrq8cKUNGVSlaWxDvlua2fGaGNekxCxecKV8Sh4x4FSOcBquy
1mjfdQya/PGrNJ/pmJy1EHhhPKcEQOE/lL+UKNdmZNWQhnHMlK9QY3eDxrmZAd1E
bogvl6U7+b0Nk3M7zp2EDTAfFGpRnIkPRME0oBzi3iJClf16DODtbeuapta8rpXX
AuA6R60Z+uiVXPVEB127ViauATpLSxdpnDcACn0FVq+3ZT24yPYVnWRGqQrV2//Y
yWNQD9xnboF+KudV98nX38urrZaIfUCK5XulbkZ51fUZr5G8K7rDy2qCFNIjHEOM
LxqF3bJwwNNRCRtYlE/r0wR6wakHKB0PSCsLUUrLCZAaQVz3aru8IFUoAOjYSi3K
N2404ZoS6UzkqfvdvFizzg3A60TWuwuHzkN11fKqN95eThemE0ieojspbIXQY1Wg
ree8td9gkKfJeiwRTJ+dHmOAFZa+okLMXRnCC39iTKetRQAJa1qnAhkn6kysFRoP
k1wvgZtocQnCpZpiqqt5zfxB3RaABsJbKKZf6jW/jOiiOD/wZaaBzV+ipKeKsMxo
oE+5vPAR3I5cP1fAUIJRCWvhPc/C87aVOOpodqfrRelJ29XqvS5LCrkAvQ2Jtfl2
xDgBij/FIXl2j8TNpEz3p8Jmra0iPmoIx6TZLQlF2zXPMW1rCLg84/1TtRdkFr9z
N9ikAqr/e1mKnoA0L9+W6X9vqtWejK1SRixO0JwRQzhKcylObMGJnLMtjXSePdpi
TEeMJKBWVWC6bXd53IpnCw==
`protect END_PROTECTED
