`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
237TwMV28Km4IZEVxcguC3ro6gxYPktqvD1PNU3jZI4O+tspDnTjIT8X1IsLE//c
A+yVxAUGKZFNdyvsLp7AIP2Ful8103Li3iXVDTinpJWbcBtLDstBjPrW0fzg2pAt
s5F5xFx/LkI1Lkgl0MKYr1v5KdcWK0TM5ziyhWgLajeMREoTvsh6GeLomzlvgH0W
Lu8GoKFCpRuR6W3fSIXEAluls1gR12CQBVfPTJQ0YBby7nSq5EcH8hVkorRfi0Af
pJ4+IDx8sKVCVfbkC6X2TGjkuUngVSt5McKFQjE7EoOzuwncVYHga0HQ1eAbyIYV
5UHEetkevM9KRTnthmtwQoi4HH38VU3wXFc0ppU96fZaTEo6Ft1Uw9WLLDc2ptOy
vLsNYT03959GH/0UUH2kE4TODG5/xjsx/SJXbQz/XB4uUReaR2CYEngnPclXamQ+
EYfX3YEK1YMj8umqPUHfp6OHuY9M7fnoQmuahOJSHlYK1qqTRZLkCMSF1Cd+xp0s
6RrA8NiiR/lXsX3VFz9Mb+vP6wMxwr1zhdYJahuxww8fPdKtZomsZvviQQMBpRdb
Tfwmm+NH4lOZ5fL8X9DjvPOdSV1yOts04bbVURgv9M/j7Qz7R9xHdDCslSrXE/Wx
eRTf3PsME53JmGtLh/UGGWuZDcNPpWxCkTBpzyS6idjwcucky4dTXePJo1tc2a7e
yYi89we6NRR8bU+xbeqf+p5HVU5IdxWrIVTgKBrVJxD1UGgVT8Y8bIgQMy5mrLcH
qy5cbJrUbCbF8yIZLzfFzywty1UEd1O2411340YBjxvB62lhUQdHPL8IjgD0tJp+
vSSl9avSc7U5UKFvTw/fOx7V4z78FIqg4gznM+dJLbB3pzQhbg6ROWuP9J7M5Oii
HD9n9Asb0HLdcvxX3lAh/0NVX47Yh9uN3sr2UMIWHeMV6+po4/HjkRWlU3gqyj4Q
lP2HvEBASe/if1X8xWjAra9+x17+KPLxYkQyLq901ScVzttDpWPv0Y0ew9HgK7jo
onWrx2dVpPygQ7Y0Ea0gWiJCERjd9idwYviZsNY5hBfT4fMnEbe/BveffRbsQHyF
0pATOfdtev76TDF02IWu+Hc30gPuim4EX9V4AEt71ZHeqZG0q1X0AK6ZcS8y1DVG
76N4Kl/akG+ZmYpTSQ0PdDB9VVgK/YormaKVA/fPlA2PVb1gZwvBiKmHVG0U2INu
JszGuiD04jqKNmNYJaFiSFX3bTlQOGneEvxQBw9jcbCcANX2Cdzl3Y5hon9PmSDP
DbrVEgaL8UDDSUwjVuBfLGrvs/Vgce5bcfd2lpWfxK2aLL1HgXcH5IieYnr54vC9
oinwvbV94S1uaheOPi67blWKFfyk47/0Rw0MgD2Ma7OwGEuK0vVRYtJygFTWeIu9
Mp5kIANfs8csM+ql2RIPBuz0WcsmY9smnLewBTMUlQEQo1FQBnEbBPz6pPsoNocm
mkJNS+hnBc0cF4o1X/f9K6xP97wNTzxrvvB9oZRhpUct1ysJD2Aj6t9X7FQXKaB5
Ue9x6LLeO4oms5rmQOwiWFLi/FDS/o6WAN+NkWm/Ag59FGP6ZNiAsLRGHu3s9OMW
GHMsCELG5tfAhtMbpxXs2VpStFYRNHPm1X3UETbxR8XxqZc98+B1Hxky9rHsTljX
6Nvh5vtEM+M1IDYjEiFZhugBP0+OBL2KP5iga52tZeqf4nSSb3S+J4AZeo6TZw/d
/QWiAW8DfiuvDo0zcPmZhvwnHOy/neyu4NuoRy2Uxj/TmvUbWgZ8RFk7dFOwRe5X
6tHdZqIqRa5ackXG8c4xUQ9pFY8dNx2QaF6yMztGgN+y5jaHjzFlaiw+u8iQBOk8
qQf19qoSCfCtYxLPJbMVM0sfgauqkw4z1hqK3/qNiNs=
`protect END_PROTECTED
