`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kL24iFOi5VOoCLqPKSXnwhB9iW8LW55MDjS7Mbwpu1gNVljrTav3gnRYDwYr+u+m
sZyA/wgcvBz9/74BH6rFaedHj/e576k3sKA5jSkV01w7BA2bHTdzQqKZI/878jnp
bJX7gx4NqiuyV1R7csJG9IQC9qBcYztvCfLUtqkEwEdjglQy+6OrEvEOf9/JlAg9
muFjpnhBxWA5RZQdOaus7xG+HszQcsVERpD+EI1PVxW4fxN54/a/AB0Pxig1R46a
Bl1nTnHxEYG+MB+4XZhC1O99W1dQYjyi+xGuoGr+gF63yWaDfB11CMMRiegeuE/e
BONAjB/hzFrMUoIBQJO24gAnCkan3qhVEOlFb9Ay2qwEyeI8qrN1XI9l3SZXM7+e
Gb/nbp+eTEXomeOEhCgUIpkOJmu7A6l9ZpNZSVL2IsY=
`protect END_PROTECTED
