`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vHI88wHCd5oYW8Hlmkf8vFNtkpTU/NBW2Kv0UyuPv8YevGQxwugceg79tR0kxi/1
siZFrPRt2nHghvSjjlOCthiitu6Mviw/mDNe7XWp4nqBw9t+j5wO3Olf9UCDVs5q
rbxcBkuPr8OP1kcIgqRK9f21VOmk4gjTnqguXPja6TyTcCNEA/km1a47+31YuO9j
YlmJpV51f92FdQkqVew+Yha30nnfoJXnnWT3GSLZp1Cis1CNzVWQ7Bu4SD7TTBvM
j7bASpP5DC0H20dcTaHgU5JDj0NLng/udLvG1MlJ4typjzdLiJkzkTGyNQBhqNL8
pjZPR1ApTIfuVYsUtHDHuP90t6ykibC6iTLu9pq3+KyphQmrzL7rcbIIYxSnwS4w
eBVyMjdDKSrpRyt5lgHTwEQpebo/dTgR7g51tu3W4apeg2ohHcT7fpH7nMCwLsFR
X3kpT3wOm+X7c/FArkoSe6JOO0hKl/CqyNIz80S2pmh8QJGAWvex37cWuvxrvNfm
PpAofxgR2eG2latSyAi4t4sPA3XjQd2rJKOEAvutGbl/6PkjlUZW8LHbekFFpDIi
zgG0y8jaEwhMfTEt3It8J25WnXIpdU62Wydpj0qXUzP3xFGnsNtutcqKaJ6tPoyg
ax+Drfy/TW/M+nq5AjLRMfou3r+cBnKnpBL0Q+6jjPc3SwHYLki11Xo+CGzRAuQI
fYCDOzzzcLOVmM/4GQuUkTy/ajUShzLp+d1JRfWGt7M7DYjDAUOG0o/xQDhKDgod
a945+KOXNrtkPnINyfdNYdAiyq0KNzdtyLWLdlyXLjOwTv/QgstNJsABW+ioqUEd
JEp66wg3lZjTXVg2oepuVAhPkpZAg2mJBkA58rVYmjsK/4inmk7zfq3INlxaQpRz
J64N9i3U7fOcbdRGBV9OPM1dsWY4aTbcUQLHMxlFqP71hOz6+7133ytzsmPnpQI7
LljgsXbET7mv+b2OJO7g5TiBMnmSeDupitbPFuNRDIYtMWjHk+PiiZrypE4Q8y2r
EoVxJwx7MLuw6SjC3McPR6TUXQQ/Ns/sxdr20K0vpp93hNsni+o2h7A+H65rYQx9
gVLUtksgWS7FTRsfznTmmDEUQLK6ecKG2zqwh0e1MEY=
`protect END_PROTECTED
