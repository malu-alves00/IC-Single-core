`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WlhrZE0O0GRxNij7fUcf+tpLFMDyMkH1T/p51Oyj3MkVLvWhHvlLA0gVv410OuBT
LwmqQWOECPNVdnG/S5rsiTQfSR23EHzUar2Mye5y8rxN7W0o5OEGALa1Np9uUf+G
CfHkHJ8pTiTh9hhz/TDZgY3U7WD7nn+H8WNT/AdJSF1S5XdvXb38GsxlHL/KSm5s
RCQf+mcaWupwIKBpC+n3D2I8Fyzv6UuRhUPyV8Tg4AtVTgTy6V2jWE+1UWUvvd3z
SW3hdREWz9YiOLWB5CLHVmu9Vk5CoCWZh35lOFFcje7wVM0g8NzAg1xaTf05gZqn
9QX6v3ylbIdnGA4KHWGXhtlwXV4X0w6C0y8GKY3z9/Pc0FuuthZxlRtV/fturLdU
j9kz9oU97fm3+z/loBSi4wCqwyClxsUABQUBh7VjrMrgfTcu7iNplCXsAGdEoKy+
VucYbQIJNbUumTMNP25fKiQNzLy/z2flQ+emNR3s3Dfe9DlZPnrzvk48syRH2vOg
zM6MwQLzkITgu6sU/rfqmtOHCo1WwdK/DQz2sSBteYY=
`protect END_PROTECTED
