`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GQyLB2lakMLwYTaQ2tVTQ52fCNNc+953qTX0jZqMMl/NwK119CVHkORqQ6/BMH2s
ODllz/lCJMsOJ2M6wIJAc9139h2kEeQUkA/t4VFkWar0TH3Z7zLFDGlEyR9ZXY5d
fUIZprxGx6yco/qkoZBjlv7htK5TcpW4PHrkSDsAQCaJfHSw9vIvlYwEe3ZPksko
nxRmz27gsYuVk+DHjByZUTYmJ+fbDx9mBgwtbVkhQhoRACkc1nToH2145ZxdaiJ8
YWMJCjl/wqtVnh05mlELF8C7tzHgeUoUfaRuEtEign2yD/YzTik4vzvkg9Xhbtgp
cPxDY4QQ9DoHeon+96t1ndRxbHyEbKaX4dG0uzrXZ7kHLtLVfTytkxUWvrXQJOMm
RW75MR2WlJH9Ilsp2UL4UP9XL/EM7VE248MbpPZAks5gIllIteOQs0SwUwfuIUmQ
20vkZg10a2kBgeqlUGPvx9jOi/F7MdKn+tTjRmol8z3AUxARvZlPndGcLgM88koJ
clRyNod0HXxxKHWd8FXd3IUAJX44O+yb2Jf5GoB8AqjUEDluagPpoRy/socItElm
2/e8Le1udAjnJSFe6q7mVddzrQNA3eHC4V71GAkGM9QabsGOGhK9olAIXwJlSkyj
oz3lkY2AWgB/CDgvwxgNvM1lgCw5UoOSvEOZST9IfBKPEFiQPN0E8ISFwx4tZNFX
CW0cpymd+RaYTXhBsYoAn9xnMxYGFaWaKeczd/iIA/EB5A0vQQteXvtyhhtSpW7z
oPiQlx2dmpVsydt/Xsj74B5UI6op8VCm2QVBRiludbKpzESt0FMWqIf0yr9JBHee
hznDbvU2XxM+I4nWe3MrkAJpCKHgUCvla6QeZjLNoWFlVv85YbQU6fkxYhPvmYLo
HtpnJxlDbnZo+eiyv30DMbKucRAWTTPpAWgbzT0x35VaxgmB1KW4pZPF4wHfIxsY
9IfhqCAUo/TPTMAv9XllD+prBfLXb6q7r3Jy5zXFLC+rhvApTohd4oosZSBwcUis
`protect END_PROTECTED
