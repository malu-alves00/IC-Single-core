`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GLJU+CJlmLy10MfMX5R+BcL4fBlQFCrHd6im/tetmUN0rrum5ZJqep6OH+OifHoa
5ygodl4QIoVxYSnnxUMeBwxKrc85Q3f6Jhn3Wc+B4jhYg08jW96glleupLFYy5HZ
OMMEzlGExSYgxTwRin1RVmhyWXPC+EHA+c7fQzpF9t6N56krkJZlwsCe8hAlCO62
jWGCQoFktaDTO67tQJNOJB6rDj90lwzk1z2MCR81077RR0+7Bw7sIyJ0vIcaPcTg
PJhkvXHSvv8f+ShEaJG54ZdWQlc833CO7gtoGOr7IayLermUIc+ei5zxKX6a54ov
184eEQ1dCQLzO5DVYXUCdVG6xi/jRLp5FBWv6vNQBbiaqu4qXZbI9lA3jjHWv3jq
5EUl/+MOk6SCRs4ki7gUxk2Fv5tyvMXeDXbSDK7gYf5DI9gftM+ZLqgVIEO0bXIX
udosz9IsxW9Pu5RgEes80WcxRGuULVgXweIwAUhoMmyLkeXf1+4JttAu8HHBF6ZN
2wr4Bg1J9b+mRjTa3j3XEAmqvjbhuimGZ3wx5zwH5+G1Mt9LLztjmp/oF5Fqtkun
wR+KfenxC3UJ4FrqURLTRrPWWT2Jp16XdsIpV6q2wcNbAJqDJ9U10NTlhDGGmeIZ
QNCUdNX+FSjUhZXibyPk3Waz3B9veA8UHYWDYbYGWGvzXIF/7IlJiS44UQ4Qoftk
1CnQR9r65c1XjWSw3XOqjW8/Nul8uHiZCqwdMuHw8H7eAW8GxObQxyA43EBPylPr
BoXWDuttJJHFMcEHjXnjp2rfM9/jqSAWecqn+oFMmCROYLIWmsYH26EqZC7VDBma
pQhEagh4zDO6gwKHHS0JZFUUX8CaM3DAiM7CQ4BdDaXTZyUpyO+lrqO21GmsK5YF
l4/uEhIuaqFMnsn6bwKkwbwgBy7f2VnRtYTOKCvEIHVXAc3MudvZC8R6gNGFLc6x
anfOIKx1yBR581hvq/3JUOxRICgIIVdK3Vmaxq/peEoilfHK1yE9Z5E1kAmUihme
gSdrG+cCMk8sqMLKMDt1CNG6pn+7qC72gCFS3dc2itQeE3X4VXTTYxTwa3twlZc3
DqlAsKclHXpwZZePJmy65mT3APURhWOIkXgYkLljbKO/wGgFEu0ZxMSvc+AchdS6
0ixnxwDozCbAeh7WHDSZYWOq5qBCQ1gD4mwA5xW2xiOqTVaZheNhfrT+AjkShzqp
KdIT9MSXP738IOSw4Nwi/VfR5dzEWwsE1k4uMjd3PZyXh+a/0eTh1trJVf3l1GC9
N4bN5odttIEyh9/7a8Ml+xPcH97+3LIG0E96pgGon9+PLAYxgdVLq/ZFpe1SeuOf
TXOleRTCVmwmSMr7BcWm0o3KVySD9zB5w6ti71Us5b11F8IH6X5XgV2YlbFHK5ga
t7GiucsTmXe91XV0YX/W8cU107iew1zaNV618kq6WfjkzMI/DzOUDnmKvKfwejRA
jsJDKWri57F3w3+VNYYL2Fo6msq3RJ0/UKkSAA1u9Xajf/BZwXUIstLLaOVPCoyS
9n7uslpEaSlnygCJ3qoujsyfO/M2ATH9nn4Ut70W0+53AjEJTfI0JuJTyQENxkZ5
mYHSOaWA58Z//XWU4xw94wbrfhYMDAvdpoJzafSuelW+yD5D1sbQuLsffGkPVouu
jtnSBPiZ+Vbkg36bRv7vmep1Wpl5Kis5tcwI61ytwHXiY5FaR7Pybo1TNm1PdMdE
82v95sPVlKLU6hzLRJZjVwprBYBTIgUZ8UKsFzoyxRnJvV7J80UgopK4DH9oHCYB
/31CRF6Zvn6r5tecf8I4Mh2CwZXBlu+bFyc/b5Azmm263XHZCYb5YTjExAEqa19i
Me+uua4/+aVr0ta0eliPF6UkWcq2/EZnIL6LewOp/My0a93Dn50LwPdjXBSyudoW
FI8Li91/4J6hwbzllIdCbu/frobiAhhpHY6xQ43KTviY21nI2V1QbM1KQSHrkT5Y
BMYSTc+LUZxj11hkFagDP939p5ePgEQgjtQuoh/NApCJXGg4R061xOZjYQjF9Bdn
QQUv41mq9BUT97rwYgdDrNJtIwOaQxnablaJB5bTIsS8G74JkA+oCC9QeMOSWz5n
OrOFioVWQJAMBQLovqf68PjBpPQkcphpMU4QXc5c1pcqMs6v8yl9djHhn9HvZk+d
L9f8+md5jlIPMHbY/aF+LmgjAcFijGhRb31kIqfTyY6RI74aWnLFDDiEy3h7OsbJ
Z5dER8eqmEWn2R4qi9pvnfNyDKmCguQgUDo7rxCwXSkhZv7eNDuU4ERP0GqPFxCL
64s6kPqOnyZLsx2L8Y4Z4+EzQVniMGkhA2G6A4+QqaDhJL2FeKvVeFjybouvMH/f
XXSrlHknosV82tKAqJ0Lq7xG3O9HKqw4OBO+ZfUl+GGqKNut2F0RDay9Y/GEpbNT
BtSbaLvs+XnZa6Zq98swO8WRBE0iXjAiMM9apRAF4Ffdy3oLORFNCiA4Cb3r2D5L
9yHNMZ+z22XV1MaK7GoozrmCsiGz14fTBOwWwLTTlmRX5UbJ4S1cQUrnWilm6VUJ
afEs5SziqGxbd5iZYWHzHbQCpEnbBgJmb9YIN7iW8OxXAqv64TI5gsUIP2siwrhQ
KdF4LEbQzdXwDLHj8UfYEa6H9IlzwMEdWRK4K6elapNnr5toTo+o3H5hG7i5AK39
R+3QEVU4lGnNBQHBoPMIqYEFXyCQ+S2aet37lzgSSuctI6J4w7S1WcUOOkUGI+h6
r7Ke1d/SdnxhUyraMUkqpklR9XVs374/DANqi/QbbHqZVaw3sXB8YEFIZHFKzEMO
pwjuj6eWWI42dFJY/3ar5RpMcvYy+svm3CJMNG3a/JW7m13a8dWkP797oD4hE1C+
xtm68vCElZe0Gc91a7UIHoUdWANrTLsZBwCuFD86bt3e+kPHxuKDbi1zfMR/jYm9
5lNyc5u/m8EBGZCOaGuyPsWfRNIsnXpa8LqbuhGS9950cC+0MWQlst0ulxBuvxR/
99JE3sm5XbcnzPNv9JMcwnZBJgcdhPvb7fsDf2IYDvMRebaYVILywuqn64aSwZKm
Gdn5QYszcEJTAen+iQiE/nLodpwjTQG2C6SKBjshO9usotYz4OHpdYu+R3c7DNSK
TbJBzpgWJCq23AU30yBwQXqxJlBAPJkmTJ2DJrOuznq/z7m7+KPBzHfpiNO5ZWPV
4KYKTk18P17MzvlXVOi3zNPW2C//RSyzyxCRozEnuFNB/4yAQ7cB840wN0p7f3kB
vBLHpJuXL7R/BgU1LOhXtXI/hT5TqzbKaH+x01/PQnKBP9e+7tNA84enGl7Sf3Z3
q3G8EsK16REfmMr/HoclElmSTGCbmz3CB7DnY8g4T+rPuEPdm7/qGQqC9SNy7mwZ
9jNaGsbLuLltj0W8wAvvE6SnlHBL+vjTDaBeajkmHZ3U8AoylSUURNPZJxX1bKcP
YW2bfeaGmRRg8LbrgaJXn5vvU6RE8jtisLijxO6pR1wym37eWjBx5Y1Aj6kSSfOO
XregIRUuJKy+29bm//NhtMXNJ5mSdiq3LhATVzKsNr1F2SPMjLzTMHWkSyfpeFQ4
qawm2Z0iTKucVawEvCTLeMSjK1y+zxIjHq8KryfN/FVN6AI/FalUaFwptFJtmqGc
wuWLaxAHYcJLRInPaZYN8XOh5SJ311RMWeEOWbCAIzyDfLsIoya/fjDAkC3txajf
MoBglBQO0YsFybWkyewuEtvjPclOw4rEYf4IJNz6LDHL9KHoh5nptzcGeM0/uJGt
mDojPOJoovLwtSM374wL6nKarMJvCCHI8jBhKHSuP9uX9JGP5K4uvH0YbSt76ock
FHLVFPxhJdeZ/kK8dJMeDy7CXM1FW4t5C4foAsRdFHLbV91GhoJBbRMcCv7NJK8/
9QK9NeBrkB8d127gXFn9DOaWDalB2BceuOhmPKZMYayHTT2am4HUfJuHuek+bFco
EK56JP2xbdAgnMDuC6RLqCJ5VPZ1+zyQ02ciiNq9r70vF6y4P2eArKnbz6JmRcE0
hJDxuOrWvfkOl9dhySH+Hyj6SLjnBoknpMiH3aomIYf5o13toWiPjsSm7JzmJo0k
pdoGwIhfRNv+EY/vc09tUtuwFRFTtgfxV7qmyU4+D09FviG+ORMgaubVsevLGKj1
Sd8xGqaRiLdI+gSLqrn+dtfY2SiSkt00mB/Ypi1DZXYSeES7C34U5OIz5TuL1+FR
V04Pi7Gj128G4PzN8hyKBvaQ12Se3GDaxShJwrQuW9SBv5WZbT1IXeHwWuxfwwHD
LOThrlioXIsD4N9jcTJusvPMl+JxYuApLSqnTUUCpvauJ+OEV3+mPeTE86WW09mR
h/AHmJD+kumc76hCIG++feCt5oxcFrlKa1+2CWDYtZ6V6E+6NTCzLucYV0pkMrle
8MGWjxzdd8oCdqd8AXo4PJasZwRo8VJWt164YUrIp1b7eegJzpiBrni0Ub9Ti2LB
qf8ADFCQxowB+rFv8/k9svH31OxAnDfqGV37ihFWEN10id7hWrHh2uqHjm6Lh01c
8XRqeVCK29wBD9iKlhW6+wHm6Ya3+UnmtkplrLDhPlZQ9QcKclkx4k2Q9N354E+N
ofEa99X0O7z2O2AMV9otQ//vEwbN0HzUsNB2CTddpUT63bWuQV994b8fHRxWcBa5
jp4C+1+dVz9rIVBJnR+M/WeqSkftajswSSVQrWe+ZZ4QZ2JiU4K6Ass0PJN9175N
0uJPiy21AxmNVwiYGt/vs4qSFMj5lSSjfZ6hk0KkTWwZVz4CYBuQU3uE+Nf2SgU2
EiiMM3msW/zsrA7blhmp7Fm1Vy1AyMKsPuNz94VyIpGOpvO64YC6UcPUHt3brQZO
VzygKSbgZKQu6R5wcNNXUXC0sS4cfUqFmKiJXWljXS/WdqafF03OrG77ZZxEYtTZ
VrSeOljQSBfa1h8TIa9aW6Oqt8Dw4BpAzYU94kKrRIzuIlJnXKy6MY3FFMhPn9mE
PL33wO01AWh8pVeHPnIaFVRSCwypZBpMctiAMb370xYMfYuDUELRXF8hJbk7qhEE
OqrtR3AdEwyLkLHxngX2YqcQuO20zllSgbod7u5Iqj99M+oMC8+4UxlA/9M0dbwB
iV+5BoiZzIvgBntM88MkaHQLiuZQvVtA6aHMyOEFnznMQ8ga0g/3mzwEE8e10g3w
MA1cXmW77nyFRNiyhuWl5AxgAUYAzfdcMGRPRLH4xNJgM3J/bDWSMwk9lTRNXDYa
cdnWQdQSKD8yJ6oxtQWkzu97UZGwO+L94a8DesjHVLsZ10IpIWRGZKFBQdl7T8Nl
SFnF4J43ySJhamnZE6CBvuE5+Tq6rd5+vK6Y6PAvDq2eIFW6ZS9al1moAe/0fKma
QHxj+aGf2hHbnrFNCQVqcXGwd0i/9yLUm+nr2UqpPwM1P9+20riIqB80hrT1/ox9
uPq4p0lyyh4lIqqQZ35ul4Hu1LJnttBB2I5xQVp8E98h6bxY4gddJeOsio317u37
YtroUEjmKL+iMQ762iW1en/LBNhUlp0R3OQ8KpEEZcNEv5WCMqDFETE4RQCmmLtF
ojQ0AhX3TaUyAH7iMGS+9RKESVc7vXaiE4Jm+MDIXwD38tOJK2yfXws7c3paIUUK
QyUX7GpJ4B935cCmNbgVwq7+M8Ob9+xteQCjALdzsh85xL3t7m24ArFEoh3qBuVQ
agHWeX1gBC0KNs2gxL+V4FDzP7X46GetM64aFa7RLEiX5Z98R7ZAumO/bSs59icQ
phb0jdpDIZfFjOVW7CU1Sz54iUpjFqzG4BB7XZJcvo1uH5HiWiERadh6Q23Zbgf6
S0u9xCjLM9o1v30/hQCMHnHm3c+LuiHCEMr74nYjDO3sEfGjyZzy9JfSjLU0+ZKd
nejj1cWc2q/LvdZK53aCQj5+Rl7eoJSNb4JgVSzDkAaz6lk/lZxIXB1PKUK0I5qq
XjQJEpOwc/cjOWFoLHPX79NUbysuAsbpfbYbeXbvHhMcX3vsAz/c2PgF28t6QcQT
kkdU6C3V3PBI8SP/tXLOIVOBjQABJPHdLWybFuYA9elpw4a5sj5fVpEIx4iAraqS
6cqkecmGY2vffdlHzhwBZJc2hU6hv7x+tefIrdMXPiObGnuFRq0WqhN44AfMHDYC
UYqy/h4+6y5RGoWHvTpv4cGTnn3x4vu0woDyFNZCup5anGHu7BQe+GtyCtWMzU7W
CAhjApSyDwMfRqPUZFq+/QurYW1Y3MPZjVPmgBNaK/w=
`protect END_PROTECTED
