`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0sLBkH2xBbDX+jskQ+z8cUFbombeyI8Qd3bZeKZitzltTQ6YzaOchUst4HP5A3xt
KmNYyRwRVqqRKJW+vNZYscehJyH1V2STidpKPYdodwAqp/Icubu3v/ut8hlvo2MU
dTqiTdtCGYFHLO6tKZYOAvuGou2oBAv1gMriddYkeUiVDiVQLkzrqPC3vD3gENzU
wY9mNxC8zovZP6uNsWza8OEnRG3HMjuZGtxHxAGAwShnLsK+gb3RRuK2kChnRjb4
mXSrztDm21T7Yaiad6EzcFGDJgMAgTweIzhL3TOI5GSZ8nJMdwM/KFgqJHpL7w/3
LJ1M7yEDbIeS19amuYqOaq2VgFwOjlhyuqwpPeExpCFNe16zF+szSpDH3jSYF0Mv
WguLbhUvAwI73YkFNGuo3I1d84i61jAD+l+jA6Jt61XA6M1sCzgVSCZzsck1wtZ+
t36ONCBP8N64K51lmx4I76OOHS8X4KSSnYXeDxMvTdc23+N3GegRHbdv2Dtg7/8R
kKhwTjca8Bc5CspBoiPsAyeN9SNiCU2iWs8JT5z1hUg7RhlxF0EfXlTZ5BVFHEF+
1TLnzT/9jtSyEZgYOGq7MTTMnHCsB4vqoIBn5vSOwVEaUYzGZozg8ov9VNZNPRA9
C8Nwf4yfjy7RzC3Fyuktwe862kCcpxmwuJrCwPE0+rt6V8A7oD9oddM4qt3uGuSo
3GqnqBtWzDKPnij81oEWJHNPWUoG5K8EDhFw+ik7Rec1aXZ2bHxPNL2Uo1abY+gw
w/2n0PM2a8ITSAewxH7T6qtgOf/px/wPFg9ZvoNJpSCXkX2/fhLJl2fZKq+ojebD
M3kpAg7eBbFm05EdNcln+qIfzIlCawfdD3/YzVYMAhgXK+ny+R3FZpUFTTcNyOqv
MXInNMG3L7XMGRPMmWlqWlIVzUBNP/UnIr/ARV348kqmxv1ufQn6dRck0HDtJjLr
DKcZ/ZcGOX3lEukRY0vV1mPruGmTz1itmCFUgCD4E24Mt1upe4rGdUvsEORCefdw
0ACPre6zOgjCAL0SywIJsQTv5yOIneVAXodW/0F8c6Ze/Kr3QUUpcRdTUK2cw2p+
9Wku+4nPq0W0By2KSXH7lkmYtyN4q60wHErKjFd8GSPxbpwKvZwOcLBW+rMKw8OK
ygGotrJAv28BzEftMY9IyUOHez7vaxYs0h8/OOQ+DLT3jTYpU49fQsxWiz9AgBm8
lSLXaTrXm0uP7s2hWGFVf8xBo8T5fSVe/b0LDm9OOP8AuXqnaTyYC5YKfyO44p6Z
Z7TrZdJNYnYhvEzgzr36xFcTQt02pQD+c44ZWddQ2Mlj/RrsAVIluDAQT0m+UOAT
jC5M3EwjLr73U6NeiVLys2kXw+MnOJ0dujOZzLEGp6xdJLhjWvomRW/hA1sz1U7s
Ggg27uZZDmlSDE1cDrR9aL2OK/6e3qXWlRE6XB3bHeEQov2fPQAzxb9APNMsTMP1
s6/jYqZD+BQUGGGHMGkPzWiwcxQ1iFvwYPaPdrydwXQbSErAcd91+VK1ismA2x0c
TclMz1z6t0CZs0DyPoMrVZ8RMf4eo14itQTHE4gWm929R9MEs3TzgybxMQuIp8OW
QUZGhXT/tWo9fqQ6ckxqZo1CZ7GvD0r7NWeoN4N2U2/Br+FFovdo0jRYXrtvt6UB
6pmh6QR1L+nJXL3nugucQm+NA5O+PcJ+dk/yiGOCBIMW2T3SE8SpIZ5Zde+t8rrp
mZSsL6W/DbhwQ0DOnOdWWyUlhGemcZIa0BU9oU+Zv0jKOFCECzBkE8GoJ7yYg7hA
jvm05/46w7KYWz4E9EqraV2su7OseYbJBh7903zhonSsS0nuxN5cvUg7/e5Xbk9N
+s0WILwG8Ho9iRVTiVoJqvrnqC/+wN4tq8Q2zAKgkJSuXzgGSvU6Y6lx+asYVFfm
DFCe5x3e4BTS4oOsQ2r0I4L1hUSH6nhCLU39NZYAN6O4mQmlKU4wTkkscn2gffUE
mNC5yHGQHhzt/CpjrR8xZKlLVCrtCNOLqvwjlcgll19sLTK0R3wTjgAApVr2o0sr
6hMYd15krchhW+XOS8bA9ijrLsfnjfspOUtHNfSsL2wSDoPLQf4qwygn6llUnfrM
8wri1W28PycVbLFhmdRvQxZ8BTd7QwWtwnVphh9ylnJ/HNhpWgpTB2u+3xlGKdle
5MUpflUn9DsrTVrhmztl5rBpYBORJ7tfjkr6IxSKpnQ7n07iZ5ai+6j9ZR3q4aHA
Y1CTsx/YpFmVw59vWN50MKz0lOeQs8xbzKEC0ewXYFFEzu7xAybnqyJeZG4nWmP3
y+0dE3aCleyEqJBTJsBnvmS3exbMSJq6o16TgRp/08r2HHKL9A/wP0PcyxDWHJfI
LEtykWInZ/AVXyIeNx6O1RPiPHMiA3lVVpwks7thBZuL2E0/vyqlvzt9jqQF0eBG
WtHxxhDdWJaJqdpwgTQJRptiEpwhoSuuku8lDuFNESzjO8oFincxguRU9OL9Kc6E
x0tvG6SxNxUJD508bbmrUBGJnIjpVdrg9zpCXurvXnk=
`protect END_PROTECTED
