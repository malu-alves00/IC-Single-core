`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fixE7V+OZq87LmqPcsitCj+ZXa8bu+hVwbx1W8jcQXEgZfUi4y/v7DU4NgznKmYw
obfh47tHpMNqTkZp4sdN8TGpBGKU0q9xhnvkd8tDrOASgwFyMunNIzdwyiN1jU5F
3sPG6dGVvXWt8cqvy33R3SYnu5LNZdSk15o2VpE899Hq2hJJc+AVcaISWWrrMCjj
V9S/pjG6OrudYYi5XkNo6jaAXeba/SOJ1sixJ5sIq68PXbOwblwEg/qYingZPR9x
YVlcg4/wDVsAzH53wbg3yqkphqmnhZl08wYYOgDojb1jX32DAYNNlm9MzeRdPOMj
wDRpHPp1QiWYswCHCVnpkuBc02LD6HMoKvhdg/zSaCCDBLelMiUGL+LST6YNT0pZ
8X0nv5c/GbCbsupcIgr+bqz686IKgjuFPZabIyJvtAPOATs5EjKIo36d05cVZV7p
hC2SHx4ysRR/emS/GHQjyXqHk/w5BZdyXkgNX5bxrcNe0TKFfFQbPcevPxrqipUG
gOnqBvAeu5AFLKxSu+sNExnNaht5QzAAGZjm7p8+nJMj5yba7pyPIb/0ELK5gY3e
2jynQfnQPtHCq99ht7l0TvZTJj/ueIGkQyyddjjyGRvTLHJmFlN2RHZiGsONNbCq
EmDPhVenLpk/9iKd9SBy/BnibSFdOAoyFmmFwIp38qa4ENU3lZzSP6QtMt+wcmAz
4urWfmDB/AJkJA2hexIU87czi6JrOv1A/pcNViy/S2hBscABBCwZvBR+PMojDu7O
B9LJLWgxyBveWh88hmbydXNYDamqEgrFsqZAgUf86YTNd/sISJYxlsW9pA/YsoNG
3HuTEQpdYl8zNi7+DUAxMNwGIaqD+gWUiBKhdkKCPRNIBJI0/KkI5f4D2eFLMqkO
oQiV0i6gy2gPK0HA5r1J+6UtUStWwBmhE84R1G+bARv+eZsqtPBEeKo+Bnio8GfE
2VUPcraobVD1R5LuQVOtSJD7YEJj6Ja9e8Q0+zlLijhEiCpyH8ZMk5pjvbPhM/+Q
rVAq9PlvBpHihPWDRpbI75lwM9V2SEmtsWWty72ZiaY006o04mbNteDmTFUJpgZa
DJhwIdRKqtQ/38eEISx0kxsytJU2W/bFCRrUy3ckbTlxu5leg2S4cLY5c2L7Hz3v
TbyyfTYglnIH3sTWnUPtwdmgeuoMLqdWZrfHZHHrNlAO51rXPMpBwKYyAmv8VAjp
og4ndpaiEFlWcojzlz/GYyGIiHIrqn3tzDb2rZWPKo3uCBmUvQHxyXlWcfOBJYx+
eBHM+6+SP7QTmRHEDCZx0jl4reaRmYO3/1Sb4zeSR9ctackrk4U1RJQukTV2B9xK
ufUNEj4+W4S6zXeZHNMhW2DtuKBplFoGvOGHQYoiNqQy8AA3YZMm/1KC+IhP+Fza
ITDKybK67d+PF7209W5J+aqvE67QxAlvgteXsxdPB2Fw6RhhOkmSh996CAi22NZz
BEuvf+1kSac60VsTSvhxxl2UNrJLe20XBk/gEwAmNIJ1kzlTiQm40G79b0ytfWSl
ipMxshzanYRmCQ6Eh9gATbfXy01O/X7wvHwE4v8a0s7/jJ1bd6N4rrOPVhaBn0iU
EhYd0y9kxQtMn7ypBmSv9M2iTEVfruwgFbQyiqRxuXWHJxxB0jhaz82s57HH214A
riLp94tGf02w1FIabg1lYiGHCl8TPiiu7F1c15WnEOVGUu79YNjsrCLGV36w2V3x
/ja6H0HKmU8JRzlkR/h6zSyNfbNvy7xqr2x2tI+GH84tXcpX81AqPXd8PX0otfMt
wpuNMQPvZLoY6ccJ2gOfPfwrI1eTQuB7wxJBiiFFkhVGkyieRIRFA3SEj9+D7ABD
su8Bca5bt3cxDvhgeUUHYqZb8V16K9cTJuG+C36Zk69Tvx2jG7BLKiiuQf3cOG3/
61crcLPBwh8vHH4GI5RTFrKX7r1MOO3vIDovq/VvTcPQwzowLvxf7p/Eug7n6HNI
VTuF0jg78UQOtC+649hzrqGsWHDaL3BTLVaSOmZ2DTov6yA+JWUtm9AXf8VTMP7U
MrxX53lswQbCN/uTk+ClaaEujkie1sfKrp6dAwJ3JptxKLUNSy2EHHrTGc1l/tvL
9ahBYXrBfTFJ3A0nWUG6JQIT9QIWyWrid5D8wJbx5mtO2dgPy0CszET18a3CpC+r
H/rWIkRZk3/JD8sl0FfDlWRf9P+p7OhXQ/PjhTNKo1+YYbN4tSHUkvl/pGt8TFEm
o9v1v/QS8oodoAjoSz+XXcJ1bS2JDEBsvzK8bDl6FfpV9nUu7kcXYxIXnKLOO6hi
rMTInfKAe0n8nqhK6/DMqZhGICubCfsZlxc0LG6848TWSYzSWkhpmFWCX8HDqP59
nnsDP8den+brxyxQNjx9cpu+4INbjUVzSyAosJD+l4m7Td2uaJom69pR7wS0mvqo
tjIVBgrZ69LoLHPxunWt8Ec9dOWJyHNJKnld5xun4DObcFZ5XSyHHF6nz4QXOnXN
e9i0JZJEPIZ4PaYbL6dJ6wANkxWWQ8fZqv1KoDeKhQ4SJ9RJWqTFakbJ/5Y00+Bh
WPJG1xkm7iAtLENeSDfGpjIwdqN0Gb+gBRfuZg8K+ovFSu82V0vETf/UyoUdiLT1
TX2jvKsXHPNTNmswJxpFoDaYxwhyHjmuz5nskjFn+C3OFZes6O1/uWj4jWdqP0HP
MDqYeqRW5BLXkMrSO2jfh5hpq8655LfkkgrU4WeVZmH0IQ1uenmGyiCzoJ+N9VG8
emluyymQ4sNQW7WnZDDpMUeYCjayQRXud4vyIuLgwkGI57hG3N7uHrpa+Kkiejyr
JYkpNIs4IeZz61mJX+oriwalRMtFVx6DxDhTqNfKVXDEpYSMEHYNMao7DmCc4gl/
bvfVTvRvttCsOSUElP9P4Munxw+xL/c1LVxCuGK8dYlmH4MTLNnpYLhSpcegVgIo
cPSSX13UWMB4H7dNNvzHf+6DcCq1ziGPs2eOIoWk6UCEJtw0Y83M3KSjI+Nm7rx4
EYW9WjiO2pvFykSTkCSYauWp6yIWXwBwDOLKCAQCnluiAl8tLUpfJntWFEAu+EST
IPHnbCQlFiwDqCs/IeC6StKZ/sKlky8PcpVtSKcIUBcmulWbE2qEez1F2nF+6u9q
elSGqvMT96UUzMWzjCJ/3lJrJMqSEzYoAyLcO2lt5SeplTPLYtl+cCLUtQJheNO3
aSfNWjtPY3547dotqdlPfAeGK0bavTyVL6ioPXTUoZNwfhnp75pdbTbZTs7flztD
Uno0qgkIkMlbXJXZBNn6V4wou7/fRHSS4hfXILmPkDosTg1qKibcIeRwuKJE4Dd4
XvJjy7A8+r+ILdy/aqmjBstQUerTsZPOr6AlGZieorJwl/fGJDgSiTCfBnDaaTV2
HTAFLoGNGc/0MfEJ1rd4swpgzIMRfrKqOOvs5w1kS+05+BKeru2fMEzs0zmREFzu
b0olSUySJrrCKgr+65eVGbCBMN1a4e3t0oRJzsPp2eWLMrBQ3n5VaB1+yJRW8XqW
6cVAPVpFLv5FyNb622k6uvINvmual16P4gb+4jXPs+XxVirQI0rj1WCxCMQxzwYU
trhMU7J9egmbGkTsmV4t7MsVZDXjOqDk3UBa36INhzhOLjakeUO3l4pkMniPFgPn
dRfUh1H/AeCJe/8uBmELRcNX6XureA/8FV5AgrppSW4JQyWjy7ERt9J2HmTOTF/x
7obF7nBES5MCTDUu8sL4Axqt7SXk9RJs+vV+Q96lQhxG2lsGu2KHULJ/forB6qkL
NZ0NQVNuWoZPdemE3QTH9nlseiSCJmBRjwvrJeCogm30kV3Nl3w3JinKZpVxyvJo
7lAaKFbiH0sX17MzOA7Px6Iffk/RVyU5hm+NbDl5IUU0p2pmSAIslYXIHjx+biWp
pPPp06XnqPOExmuBlv0VaZbjtZovbdJFfsi/pHRobh+uANiTvc1/EWkmAimCWcA+
EqackBZG5boGWdXKa9Z7rOsxXCAv8aENgRr60GbEsYLNhLDxD39MiqXjKyZjsHjR
fuEfWYj6UPkE7hbBAuc7dxwJ66CY7CFltBQUlyJ0i9EXZ56IaE9aI+pes0t/6H+X
8CCOjTb00vwDYMUyX82/UEnHAb4AlXmxShV8uA/6KA7kCvGeOdkpIknvsV43YUvH
J0GHTzIOh5F9V94rzEUxZCRxbTXbll+lizTQObA/pfgzDQGHoaq+XHiCYH8ussjF
h9wgVYm1jBDFkw7N4xB0FVbrrmyM6kgUj+OeGhogMxU1aiAmv8C4WYHJKmI32k4t
0Q6ydSJS2n+CVmJRB7Te7eo8F5wtzl8eR43bVSah2Dt+IKkKHjbd+AE60Gc2ZDXx
C8yEf9RIVQWaElNlHxeIUafotY3adtnpyj00Ib1JB7v6WiHaqOarul++CuDGLSUD
g/6ct2FVVS3Jh+mSkCzB40SJRjJg5IQtcWL2C/fzvrON1EYka5yxK0zDxrFfK7cy
1R6xUW+Jkyr89DVAiQ2ro77oCrtZcjCaybelZW2+10SWo91TIXffo+LRLvYTbMue
JuLFDudS+v8PA6NdQu0+SepUsXTpSqWkOG/HRr8dxnSKj0e4WTlX6urPEZzJh8oK
+LZGLEN61jdhpVVeUUwjxmYNtm9k/5rvrInoZXgAxaU6Bd/1PxhkYMkvbRZCLhoS
9X+Sthn+yEwjcSuVQu0ckqlfbjcUPFX4CfwrUiR7VJ6IPoljw1DSVGAynrwWEOaa
WDeM7O+8TewZgdbIkkPCZuw9lBf/u3S0FTOGpy3IxZbbyoc6loRC7/EzckonLHhS
jRH+YnHbVSj+Ukw0oaBxi63mJBWcwhR03aiJybtnDyRhcbzOv9CTofEi313iHJZE
vaQPF+dA7YEDQKa3zXvzrvsNsx9aBz+bKlOjaKkUOTEX/6WejcAOmoBzTKORLzau
B1fuyNDTOVxoxlhT5Va+YHlfPYqrITW899kCYj3PW9uiKnvkUhkgHOqUV/m5sI+x
Ca9MhTuGt37TngC1+9ZdmIhWzf/aNImvl0/cIaGpAW8B6yF3qEj+UUa4OrTaz2KE
vACK2y3Pl+ljMWgh0637cznRf3CYxswKoTozxhYu8kYTqBhN5DIulBAsH5HcTBUl
SYKcoSz3111JDJnaqccPacS2IiPuAX9jd8tAfWUsVzqAT2vFofCNP23QCxWMViPd
UhtU8ugE40/vOsVuQ+iBUYU99wd9Y4d3qun1X/z+CvoTdacA8CtaRN2hwl+6g7Ad
m4xpHKvy6DAEE3nZfv/0GK4SHbL4NrE41nJ30FbQJn9h2IDxLWjMAR/nD5sOOl9k
mki0VfbaM1FjsokKh7eBQvrbyfRCK2YUUY+OJxitiDk6d36I1DA64A03aiFOwlk8
IilFHw6dyc/xEVFJI9Ny88uL1AKITwGHIzlTs70Wv0J1iU8IUAKqCcWoR1bOc4xg
X/jlv6UbUXWFK81NGuIX1hbs/2mqhpkXBRn640xdjTKecx4VgaD1HWT+OC3odXon
0WHErJUkdiCbjk72m3iWU2O+hAQAp4Hr94raMsyAOc0/W4d2qiEQNW8ZbZbEmaCB
tQFVcLAGZdNHSQSqy5nDE1oDDPmsvZHduMy0OhaiFXAXo+9JRegLu3MlOpYvuwBf
QSLgQG58jXhHa2K9z3vpl1NoZKwuPpsdBcSmIthwobKKqoCwMKwAXIPuIYBgrIov
DsJvz95rBSaoeYLPr0kzVG4qCn7RE7iihP+taUvcaFEKizearlqb+WgvReaxJMPd
iLSxPIH+KsxQWj494iu/ogBo64+b3Nmt/J05p91vlSe94WjzsuIhR3Svdg0tSx/G
sRNkAFanLxwh6yyDK9/Gle6f7rvRwf91GGvB2d9XKc77CftHrjDCiiMjhmZn54+v
jkiJr+27zwhJDQ0P1k/spveLrpeLz2rfDsajxTW5tcN2GrPxPNrsz1dOBqn7pL1J
LyaAUDKxGX4CBbQPhM+zUahnsUuHZ4q5A/OQER0j7BTC10Z019c/6qH2LI9Q4JEK
xRgEr+cUXZG7holav3tN75SZQgF/DIlGc1fZFspbx8xh5kEgKCFDBTn0hjLDu8om
3/tMBd7e8WxXs6cdPgPiDG2YsKcMD7+fF/4TFVCEkpfV3SwBOeUNx1AE200zz4Ka
1lx5oOAi0TOmKKPeRxQ6lbqtBQfnGOxCYVJUUXYD8l+Ps+OC9VfOb0AlCz/ua1OJ
/hgJg0JX2ioR3lK1QxjnhDoUiAueF2r6JSrNzeoZwaH7VgyjZHXJ5KTPMGZxmEV3
rEmd5j23ykmkbq9XHlHlhmYqRCKg3UyfwiQrkBjn+crw3qPE/HpUNSurCTMF7wTt
V/kKXIHL2UEDMeK+s/tdxfaumP9byGtLDdtGEeDOTwbIYSqzwtqnwN62EvGtmyIO
dMfZYy0VuHgRfc2AigvEolXlJ4l1eKKosvtU+K99t6mV/jadnjUm1P8Dpc1EAUCO
OQXxHR5L5z4pC0x5Hyi25ECD2Ok5g4ysR2sRX+NS+P4BojuMyhrtjvNuuDh4fBLw
GvchtEv6ILb614H5ImkQ6TcD4FH+JIPB51dzm/py03vjvhFEXiFnRBaXofgpgak0
6juXl4KsscUOaTSuplJEHag0F/38440qNKq2nonTLXTbC8MKp6UUmdQyarjeppfM
oMUopJMJkqq0uGwTOXvlT9E/2D/AZ3hmd2HRk8DFoMtrK+EDkgRS2DbCYXUN+fhv
rgY065A4LVRjxovLLTwZXz6OFijQgGYh7tkuXRTdIXVjv3WeLFBmfKFOU0DwgwF1
1DVrBoqhDAjTxmJRLRjSlBWTPMUR0TaE8B5OEirPh5bYu7ztUwKpVPxIetRJ43Ua
+lSyfO268xe/mt6G4Giu7jYth8xiMlSUE2Cr7UsX3rrT9RxjkcUkYGON5HH3bul4
mzRBFcJZHT+7D4tTERya6PnlZub1ha8qqolKlcTpYJUEvXrTMApTpYFrxd6bMzlE
h2e1tpOmPC/32a6Hqt6S3zG2fHHQ/UUDdmkcMErhtRrgma6iuEt4DVyzooScUnEY
hrCoTN5d4wvVf/tvTIlXjUnrMFmD1gTcqXSTJQPjTFhJfu2SkiXK0eJxFqUjxVTi
Rx+/zPA11XJqfxugyDlec+VENZ+YIMngvvVW/kHm52GsgunXqOggMTVocE+9yRIX
sOq6WEEEOnS8H+8dkO3bGA1U91MNdk7uI87dOqQX2wuXUUuaCNFgki8509JUFzYb
PvBhJLJDJz4RRkoG8xToIai9DBYgk2FEvuS3GzHlll36vRUoKnn19ytYcpBdCeup
hcjqXfGZT6telgwL4jnEejUlkyT3lLv4GvGfugNKdi6NYh1cWxnR8skB8tt32J7Z
0rtPG21Nl71M2HqZ/ugtXy//75E+e7gLpUZzKuNDriouOJGFKg8w1ciLKJCJYrSz
b+E5Cha5YVHLk/O3XJ5ialSYsEB7qVdcT4NjTFYV6MSOgnuEKX9SVdNM2Yt/uIdd
TV6qW9MCaI6ateAT7Tsi1Idz9Yi9WAHpK31BzGMJaxsEySY1YZ+gXAC26c/hlOpT
IAvuGvADgxfuBVJmmrknXidXPRdlkawHJX4k0jFNBagb/mha/1tV/vDdyX9NxJPu
yxcOAQBJFzvXTzDV2SoiWXaShxX7pCbIol35yz7sQdLiI0PYoMCXnMBs1IHQB4e3
CSi5okGOFMTIfvaS+xUdfhB5ohOIXaTJ00T1CuAXSBu62WVlI76g6KkjFcOj4m1e
XShVnxhK8gMLB9xAipVZMVMvpdDEqKBLt/wUPoqctvCnOAJhDsRM+4aPUIKgAK3V
+ib3lUA8NZPh8SsQfxyA2/KfjDPOiIFuZYEAQNlOsDbfHCMyL1OoN4LV/4wqgk/H
dTO6FdlVn/xFlPtcG4TlvexdjucJlp1FZ740hBRilJ76U4YUEXpa+8S6wrjt3Qw9
Ev77Bxt1XkDY08PKAww3fbCHxV6we6hrP1RsQWnHd3jzAAHVEFZylanN1nRJQqlO
hQO+iLT69pJaXpO4PdZnqXdjGcXvAKjSOUNRI1FlHMJLYylWYF1afkoVzpe/MIzH
ZZNmdQ50YRspI9S6lOMpWbR6FQBR31RTWvuaW/MM1y/2/ap1bIwPqfxNq6Km0Jjv
SKktsZgdTcLRcAG+Xgz1PO4wnOjztarWI7R7y3ypP1+I6E751YdRHMIGb7zRGQkk
juUa1oWSwEwBDWeZre8aIF4a9STwHeN+Pmw7tLY1nW59k9gDIwtbMuj1uLJlyntm
G078goMkCOcW0oLv4xYkM6aq9EmS0VJycC7eQ8WTvH81chAhK6NfYpC2JkF1/QjV
D9oJYuji+YsOd0UjwTuKFY+L4wDjUj6WObeewrCFF1w0UPPyMMme+hGUI1YquNnN
PsDQXKCvNQlvc3WyL4esw5KvbmrVyUmpqwCJXbDJj4bYbVQNueYZVSi+KOEjZjwN
zvNUTqHTTgmfQe2aXJvy0S2BItY7VHJO18SNQ5dOq4/KaCH8/7ItpHzlHvRJJT/N
4RuFGdbKdwjBntAJHUU17dLr3Ha3K7KG9sxbwfRXE1lzzA8C6KFbrC8Xg4b78QEe
ELbf9WL78mduRlbQiBBiBeTEgIcyN9zeK/rpt2bFmt4hGr9scSuKmF4GIYohstYU
MF5h20wZ9rU1++GvXWpkPPiX+lw9X5PV8IJHKmAY20GL8yTz54p+HcXxLuk4M5er
HPB9RbJBOnYiXOCEILyFI2FPbJJojxnevsWi8Ab6uBDZHaMmLSiRodWlm9jLK0KM
4FXtHL3ap6x97cDXz+h8+oSE1uk1NZHfzDanRLr6aTGWLdFPTxZZs4Oiw+NCQGi6
3/ZyOkXzFxzo7pzpG5nL1dBlGmCJsVc3mw/evgbguLEBTntBKzeRwq1eaCa4T6/+
KYny4K9SUs61KVWbV2uGQabTYru0rRQbDQ3fDbbGo6zqfEWuXXvKV65fo8Cgf6nq
WrmpfPZuswlWcxXV/sQishzdKKmCgu2B5ceVkbjPAWYf/+eFcpwMcy8vDb0J086V
GGS4E6I4doH+Xm/w0pgXruUA5cndCziA4aN6rSPcd8q2UTjzM6GBqDnbs+vj5SzO
sD++bBR5Oo+wXEvXZnUfVn4Oi1Gja1vlvHBmdPHr7LTwXhceE16vGbRZ3VijlPqt
ufkFtPpWv8qrFtEZlh4gz2Jc16ufja78+vXVldnbFqauHjIMcafAIUk7rKFrj+B1
Uk86TS8HohUPft1lnow/tIQ0NLqicbvZy38u4usB9sMSzQLTj7nkA+I5OIZl/6Ll
fnbO+cNgRyrelBWiiCF6wQT1/BjCXHOqWJjVpe1M+cpkimcqm8Qxr0ReO6gnGrIw
S4CzXqcNF21V2N8blLtToGLP2zvYW8/yVcqaGGR6cVkX7e+rBgDjR35fnsIGqUoA
HcI7IlELroNoMNxX6GxsWhVlbOymtmQIE0A1O4K2GSbQ4RZZSp27FUavObcshfiC
K4+wTjZe37FY9x+3w/oug8zINmodFDKVlPK451V1uExplkr8L4+J8rq8XWbFMRYQ
vsjvhrcpIXx21fs4YBkRFniySvShOBVilX8+01ruXqUdU4riqKGTsBnModNuNA9Z
QY7+qcLt1ivGFCVSGEoJgX5Jqo50mFdunY2GbSmolmAOIYeJWxE/8zZVLWq7PNiM
CZ7NwtQq4yqtxjENsmqRPQQN4D/8o0QBkEDqERiUn1ImdA3SF61kIGM8tPxEf8kt
ryekXHdCs/5Gh7ihOLQe7gibRAWow1iHdlDaNcAZh7LCauTTHUrBlsAq0gG7nM9i
qCWGMfc8mmAfmEps0jAj8vZN6MYF7Xd/DAFO9vvT/GDYjLmlk7qx0I+B/au2MSGE
i3Yj2XIn/8GtfdAIRQTtcPJOXWH1776ts8vhuBnPmZsWGtMO6b4db+jQUupomtpF
hieGpdcexlwH6NWzd/wTuSrkdcGCwNG4ygjyjoXRXYf4VBmTBmzLw0d28foHKQVs
DOtbRsMTEYDI8gnNd725hNov29//I4NSBi0JFTM2lS1N712H7m4dTqYzu65utc4m
1JwIJIk7mrQyHZtxeIXmnbAyZCpOb/1UWkJAHaVp/WIn4t/U/aXPWginjvXZTGnJ
/YVmo//ebH4FYhGj0pwNPzT+Al2J1DATc6/QcQbPo7xbH9Mc4Weh5sUNlmuHyvBS
/gLqWYT9qyUhAtt9c2c42CIeHip8xw/XEFg5YaH34VDn4B+070OCZmXRibNm4y6C
aWdGfrhN3T9Ke1l8P0beNMfYVVmtXNPyi23hS20veW5w7rNX1UPnksqKsYVJzGGZ
//XcmbAiYwx0IY5Kp/29v+Anx/TDfPi1whnfQuSIQHKbMEm7ttl7gkrlYGLpZkpP
4Mk8risRXOlGXXUoyVXMrt9ND8NuS2q4GBqQMRvZRDBBp87Yc6Gojh8gSq+XotS1
JOyOT8g6VHTeCNMM3V06oJZtUlh20v+vH9N5rQkTvuzvsCyFtuTEs1Uk7rnNWa5r
8gFUsSuVYxKGNq+QwlzL1eWd8NTdwKEuxirLyLVMml4e8D6x32H0uQnDvmNsyWkS
61a3+eeEovk4jJCxaUo5Kjvy5aXLEa3hpEBMrPQ/Mtk/WrC8nxG5OZAkPl0MZZ7I
L07WV9sgQmZ8hv0t88VPCjgVjAb7oPJ9UVdbrWZIgFqJDtk3HNp4cq5WaIMw9D8o
S04rs2vJnNLPgMsIo8axiCM24SRNqLCxO4njbxOksrkhSCVP8m7qHWczQ3IizBbj
Q4Y0Su0wQCiLa4RWI3LtZcuShyMEcA6YnPWx23OjpCdt/NGT2n3kOATaZBJVzf8x
/BS5X58ermvhHSqLFU8fyz4xsH7C38jXA2hL3TsQt27HuAC+XNm4z62+UPVnHRjW
2oEkYtZsWfiy8zdES4P+ouM5z7yc/IQklNWaG/ifJC/Y++alwQS/80ErgRwwQ+7r
2iIoLAUyblvtAZSY9FBREEAmmkcbnKm5bE0r5tOPqnalk7Z4KV8gME7/9HLTqVHx
quX/PIZL0KluqFoBzVRYbF8184FBPleVLdACeGldVexqpoRlrb6/4vcg7XokI6Op
B16lsgaghHCd6YPex5G5aPfrM2NYGMNxpaNHWvtzRfB8pS1owaCazwhR8VNYZndU
ji8wdftEiCrXgnoTP8Z0nyfyKOJTlSfTof6esvj7jclrLf6RXAJ0qRnw3sdvuDJt
6DcW90vDEmOvYvDersIIoH1Ibx1HaHYPmJQ02QfhPl/HVPB2qhFjhToI6uUKUYzd
peeBxCxV92cgOGyesnXYYIf1NUFBlUmxn7zmYPxqsEUhosFUZFEd/eRU6dI1zzvV
f4EPXhKzq5cEGsuOALxzOeu8tCHX8Wm5rZL9PF1UDdjeBX9NqGUs8e07Kjx3o21o
CiJBJk1hgDgUvHUlAX0Mxlad3pledXHxUROtfM8J7CHDnjMMToUeTp0CMZzQKezh
mLVmNAW2yyfq/qT/qevmUrZhGjmKF3WhjPOn3eRHHr2/8076rhvqO2VpjDW7K7mh
mYo1zo5VTYyjhe8o/ULbqg56EPGP7vbQutMT+MQMCRdAh9c3+86SRwoVhVmzZE1p
drgcbHGP+7v57ijZz/XgoDpq4mCjty7Baz+8PPAVBK/VF43LZkobn+wRssciFu5S
DoVGMfotSQoCl3tzB2lzK6RT0AYMftype7m88Y8ZJA8rkNrHAzaDVkXqEc5fPdCH
trnUAr0fQ5A8QoNV8mVZNJtNJDy6qdPLICFGkm5P/GYdZ74mbvPDim/OTm7YxCEq
I3xBw9TgzK8Kcxmy+OW4LM4xVszy4i1HhRCKtp8JktKVmn0N8prpqa3630gIveRH
PkYDlVRjj0d5KvJgVSHJtG43NhvqA3vIBFoizJF1u8yqKbnjnAL5khshC3eHW2Ju
3QYsz9DeRwWCmC7dXFinUj6i49i+QwHoYn3wxUu1LOlLcNVj6H1xxTRmdpd2pLsj
8Cxg3JdtRIQ/HX6u7LOAWdwmphqD8gQNniQEWU2Xw4Fv4FCrD1ChMdDslAjRFd8+
Yh6lKn0AuDK6oSMM0s2r6f4t4a5oOxjQrvreLNbJDmaeoz/8dWCUjokFGQ1XJlv7
lJpaDGzOOozTDge3DE4AAsIERJj1AqL1rXYQd6E95jvsDes/VHeFD57ld++7xIJY
YrTm6VBHy5fbqEQZ8s6wUI1hPcW/h50ZKJogDXVJEh/ls9kb/KoGBd47Vejp65sQ
Kv88rNTSCe3dfGeVXdCs9+s/yjtFx1oJYFSeS1aUxVlEJPCiUUtATg7gAAA5kXCT
XThxQRqv/VYl/3WH4LuY2sA/CinZDm/9Vas7k6tneiiCg8AvytAXigMPY9HlcXu3
CDOz/bMqLK7URra86cHeAzhga4yQqNJ55XGzBaL6WfiY5c7VmohkAM31B2nCU9ly
BgunsDd3i1g419QB4zgDkXIFW+xHlfuHKCa3Mt6wsq8nf5Uj9pxU8Y776yWCCxE8
1atc+eYIi81TFyKr1yHZ3UzG639umj8iem83c0SQ9pVfBU3jpes3T1+lqGJqIv+P
7PdY4vVZQoRqZDoULi/DwRx4UX5GjvkAWh5YZYk+RGTV2acMujmXS6znVWw+Tkry
zLhSCDGFVm+IHtwnagT1CSt2MMOf8U0PPW9oNNuiU6tYx1ZrXulCuOBxREWWdrpz
6OOunfO7EiaKb2VW7HGN5TB87J/f3gRzpml5kq3UnpJ9hbLOe9vu/mHcsE9gN3PC
FFzMgowf78W9tyG5VByodwhEaHccqvvrH89pXbWXjyThuTpJjWvS4KfCYNB6y0VP
Hh4qw5jaegfSiRCBSrPHBc0isxubZBSJ+D0Udssl0DPe111/Hy+rZ7uIHtwKRprz
qnoIhkrVcKRiqhsZ8OawE5WQGZ4hoWuS7QC61u3s6YPdH0/+zsCLh+7TCbqguULj
OFXVN1KtjOYONuyS1FjpkJn7i/2i0ngbXMUEf11Bn24aw8JiQL2jSuYVewUN1z+9
PRrixABJp7GIqfRHPrhC+ZKQqI44WsBxy/dULmLNPYw8tGCKBsAFXRuEJsnZcOxQ
g/NBzztkcDWSuPLKpLaF4joSIu7+pM4vSDzXkpK/2JgHC7MdGeXj5SJQwObORMOl
P/4SsMcmnbbhNzIXkA9urEfcIkJjANMrD2DPF5VeRNgcPOkI6Ijs92f9/er++oaG
f8H6k0FzhrZxWOYILe42A8T0NPNT5oYkiSsPa2vPLlUGkNNaYvsP8UgEL+si+/3n
Enl/n+qwiCUVdFsGeGYvNdnqNu5Ak4M8DTXGJdvP8HIqx019mVxOTRzie5nXUjaM
MhyveijyTVBaJYaqo68MfeVp0KIrRiWkywZVjzjya7ET8vN3FDousna7dT0Q4sRJ
oOkuWQDIWx2qNlRle5Cz6JMvLw2jGAaXJscDA62OClxnBGlb5dmWE8XW5IaqkTIj
sja+kQz5udIYAdHBpjstEVwcOlD8PEftFI63n6XqR+nqU7GULtuUuNKzOKw2ze/g
bgOfz1BOw+knDsUbYfpUjRP9R7CAhEpZS2fq5KnTTcOa+HE/lOlhuWQMnjFvWcLv
RqsxOFpEjWgM1T9+8iee7j08mz7n4XhR36UJq3A1wY0LPD815R+cGjdlSg2DXTpd
cWmldizIQa1Yblx+dw2c4j7xt2jjSNUF1HNxdAIvUzMJdcrSqYRoaxGHZj9k5bIZ
svyJ/QaRNTFGQ0sqZmpGloRsahAlqf2+7B3SptbfBS7JYf+POo5gSL0A7b/d1lF6
kJ37wG2NaCF/8A4HenlgBbUGRtVf3rUnAaxYu7Vif90GdBNJFglsIyRcXqKOTYQN
zlFMyO4SIJtXTHqNdXpJcJOzNvQcJlmqZwRDdiffNghWOf0w4nlNBI6hshvnqykC
Pmok44eRQGAcZzeEK/GOuHXvau/ltq5xF2jcVqyT+MB9NIl3fIJHCS9N+vLAcYoF
s98rjIjjV/JmKdGifdrE0EjQDkWArIvsL/aK3lrWmpSVsc7KF46J6mCCuVA9B760
xD05dUFbwweyviR6wFlutLo2gBcwnk/br6Ov+G7uSnJaPGjYblxadvX7RZhzEg++
Twlsp7FajV2HxMRJKM/2m6W6K60sH0lfJuitFSrDJ4L/vbL/fhHjvBHNY1c+23Jr
gwJ2zluqKdtvNOj2aHFEIY4kmyY8nq+vruO/HzvUgWdaQ4zIwiQwy5NxKpwpGL3c
/+WovkUGhtFp91nAt2/3S/GPbdvRjxjyUMg2GxOWBsy+8NqwD9vDeCXhPZ4qDGB4
`protect END_PROTECTED
