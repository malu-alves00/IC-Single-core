`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0DfmhMTNfFNv+U7Y6VWsAZhsmrow3ACOaVHUi087Ujw33NtN/pyUw450D8tTJA/3
uUPYa5DKvgMmMha+g57XolffQpg/DVCoNBnGI4meKFsfiBa6KbTjd1NQZvOX8PKA
yaIT6xLDCdoV5cEkYiY6/NZ15vjPYy2qU+ZpT9251BP0N7SoGPrTR9Zfd6w8Jw4s
dccxUew65MeufsxF+MiTFX3sAa3Jy/j7Wt1AKoAr9KxPBsRuvR2r3FYbqZyBDcK5
8Se0Cqa+7AhWi49EpGZJ1+yL2nADxYrzEYwdQwtTFsuKhESPLvUf08xKPPO+FSkA
gxtdAfReeFMpbfQDEJMXjhg4vM0ozv6R4wH8RqKOfQUsgz0nrS2aMGh8ex3dn3sw
C9yN7IxS2P20n2fruss2xNJHE2wiH71lGs50X5lB6Am3zVjGGdkdwvyhJYOPNsoY
p1Uf/YmYtmyKkGKFygfpcdaZLPEHWAUcOgcx5Y0N9E/JzrsFjkj/sWY5+kG6QsqN
aFsGKjhqViwKTw8HXPDdTpaESsdBoMLlREeyy4R19aGDlJ1VNcG9RYe3KDOuBVc+
BGU2BgJ6uzj0pCXgZQKkZNB8VFmlQT4GiAzQ9B9sPEbwX0ImNAvyMJKNbAYd5tpN
IEbMgGThZRIFop7bwKg6LN4ewCZEPPu4sOVq79hQZWW4PFgmx0lShuWkL5xmn4OS
3qlVfTj1jSvOhSJgXRIlXlvEqGz5wbF4I06AesR1WkZPEs7NLJ7dRP2krjLBQvis
Rk270uD452uP8zE5T1zQeg35IAU/cwys0G+hZARsNKJ9w6t8bnhJtUQaRfRioqgs
SgMWXejMR4JVCw7ehkFEc2s6LKALJj2p3K6Ofb7DwdOhoWUtWMkvxf5oXlXYL7JU
lka3v5yRbkZWHh+Jend+L1sYmT1hFl3HzbIwObgpbwveZdER8wgRX/Ub0yl94j2u
eQ8rxD65FrMmYWElGxpJScle9dLjj+HzM5+RNjqSUciCtLt9VVPQukJAI/ukXBJQ
NzapZpYeeoQpRSov8bTYmkgtRunLW8+qDjEB20QSBtKzceE6QYAvePlKhDNZBSJ1
RlNxMgeE7R3IajVpFcQQ4EY3VbBoJuvCabUY2P8lDSgpgXZy9azNQXD6crrIevSI
Jp4lnHxGQTUTJlD2utGbFyLl1wT7RumyFf1OyABFcDkru0xm1Qd1CYPb6WdLLHil
7EppjPxG7iveD9rCevqi4bw91c4VX8wH1XGwtPiyief428a7640rFhOIiZhF3qDh
7EV1w0duizh4eCS1KEJBXpis5qZ8u5rcqtin8MRSqcqky8bstDW3aFSU+MAvE8+q
hJJgHjKubRBIfxOGqCgkBH12Tgu9E0oJxw5+cvp+yjwndByK0k5ppecIksScWLxv
Kf2Q3lRxMDnRtibq1H09h/nqrblfv35COHegQFtauf8SyINK4jOB98Ixf6TkKk1a
kbyI4/PNFAOMhYKp8rtk5K2YlXHphX2Za60rqd0uMnJ+8mwO1EW1xWEKiLO+89nN
Uq38jZvTdjOkdEKSHnnwikumbaxix3n35QJAlcED6/1o1fJRItMi7PRDH7p9wYqK
9i2iJZTdQfb3Hb94WTrKHUMeBXh3x8EXbmeAeLkUQMIzZfOF+qNdAWlQcQiHJfFt
5vTBlAxz5QEK3YKs6oPDXg==
`protect END_PROTECTED
