`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mPy6w7+w/jjQR1RwAOxkWvaj6VRapF3MBDJCi2+6dh04k0HXEE9rTrkYRq74nNE2
yhHdS58O89juJc5XuWbPMiEB9NQx3IHElAmGS9auY/4LiLfc2zOSNS1lVv3kclCB
rRuSHdTaZr9KlpH3xe4u0TGGPIcu1a2FTqbpKU0b6pLoucTOFXFW6sNmh2zBIc5+
Njhp2Phf2EcjlxbIJoYr8s3uj0WuVWULzccPR+qQUZLvJN7dHdyHUuF0K1Wu59Y8
mUY65FtQoigNHnMXSRKhaD2vh/hxdLq0chrcabcHZ/uOp7kB/NPGuTYbop/puhPb
muFgZWZNxWiw7wDjgZcSuLhDnujrio8IH/xbEQuPxavdvx6Mi6ouESlw3z+gL/G1
IUD1m/U1t3h5Imw1IjxcVHJnwQ402Pi+mQqg8p5WXPnL0+cZN23CntPb6fTauI4p
aoEevDzPOTY8c4QMYthJqByMMgf6ugeuEKBG6Zw79wJ5mD0d4HM4YKzW5Zfg7css
E5+IKQTRtFiiHk9niU22R+Aj1xnw60JxdoZtWeKkzCzaR2gSYuXRft90q6P6eDLQ
8GOf3j0+SUhKXRm4JcUl662JuI95GDWjX32wcBw/hZxj6xbOpGamXrxUbliNnHHn
qkwgJghozRvrS+2HnH1xcQHiMZgSLMwKyBBpttMKYZdyuN2yVC+5ByDjQw2o/tY8
LOAXtUQZTJzNG0GOSPeZ7PWgm6VTmER4Xl3uRd6gJtyRMQeygGaCqRUpL9wH5m4n
DILmLO1CJvT31Sgn28WjKMd1IhxOYCjXJIN1rx21zntPtTt31aGYY3UPOrlFdWhb
Qo6NZeUethEL37OxaDZ4DMB1f48w08+IF8+KPtMPoVk+Kq9Ayk6/qyQjg2lQOu22
VvBJAh92BY1I9CYxNqq0ZfSZoNgyGhKkM3USfU4QCMdofQ2umtOFOTmUxpfM1IDM
KWdAj2uIiZKuksv/NA3f9gmqs16rANyD7GJg5qesF02DOyZqPfI4fISeaFJd4OnT
stGjLwX+KOODEuCAvoYWHVvr3NdeSXLPGeBAmxqJOnpue+9CuzwoVnUhn6Y+9Fy7
Y0KKjg98DCX0/S0GgzMOCvFdq0LjBaCh679lkkAamTN4BYGWnDxgWLTANlIvh5EX
EuNFTz75rLrt9gTGGHpbmC9u0JacJgy13izT/cTL7r3lH2ulEsvwsOzBZnY9KlcS
NTokPlMqlnNLnF59Gp4l2jdS3uZSZl0bSnsvL2a0akd48WnVHvISBbS4najVQoC7
X/NBrUmpso/R7kd+MXLhmkgSgEGU6VYBiyjedGcteTTNqINal/liwcO0Degu5FKh
JBVrpUB5OI6ZAGaxEHsNwM/aQo8wlhgjbUztS26kHBn7onDDYtcTKjFdGulPUzoX
FZdwU3x1GE0QeHe397M29p2eSE2Ba9QBcBcwmjLTnBNHEXZioz5dpktJjx4USxnW
GI3NrCOZ6yWbbQFap6SzhexJebq1AkjYX2GDXX5I2PeMvMlgcq7fbFMGUbiyGgSi
3+wj/4SGsDnK6+CtbrO2SQ46Fp2hg7gqLUtaQuaC4nFw6aoBN6uQJIVDTDxyU94A
cSmZhfvq2JO9kfNmFW009/VCtN9nf1r2rU31FjPGAeAjmNPum7GHRTUTGfp3QR2b
rTy0SgwahfBkcg7yXym5z1Gh+o6AC84/ogU0njc1iiJCgUPRGMPi5FgrXz0FyPew
VdVnydKUQW5gpvFgmevQKg5wJo3s73iL+ID3jENhrXAy8AxydsdKq7bkU/j9/8Ew
DkfdghU2L52EhI4XOV0rNFQtvvmSYnoFFHdKPdQPxNr0k22qCJ2UtSv2jOjFG+gG
CBOY8Y/NeHw95CbeqfNmfEHOnjwdpVHvxrjImgNObRpu8AYDZDUf9kIlOGdgsEeJ
g5iNbta7ey8uZOBgFGfSbnmKziY/jeK3/o7crZAPt2sosR2+/jm9zPoDhEg+wCAE
plHQxXZUMFhd+BsttHG851Bl1xaPvs6is9Kc+9a6apFkqPka8aAv5do07Ha5Ibaa
hRE3I2o+KYjhck1As2nUEDq8uB30K4erwKWoLc+iAHHUtRsZHP8NBBhBzpeLSWN9
`protect END_PROTECTED
