`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CZddHAKpEFKBSDbvNA2eFVzhSdv8+7r9uGX5TlXvZgeodL3NkY6CFlvR359w736i
dOsWCwQllXty4oL+Ivv52oaA5QJX0Cb3noZ0jAXlAjJV6mOR4qE4/2UIRGLCq6Jg
Xmil0yoFFMu2tDdk4VrAlYlEG0OpcL/T8pA9V+wL3UEQSUbmT4VkaXY5dXQs+oW4
uTqlJJvvWBNdwOPha2Un33uNUhITdlZqXH5y/E6ThrxR/obfXyh2LqTYMQemCbdz
NL5BzTAWwIfbQmDYHsLbtgapkl1+s5uAjkyW45cmpeVULDetNO2hZ1wqDZSddZGJ
A7od0a7Qg7QFcXlmAsrQI4pDfb4IQ+pESSrKsK1odSFUf1YJHIqq9MciMI/hkk9O
MrKT7ZKTuyRofB8bxauf73IN5Y3IBPa0fjuar/GGGVezhZsIb+dTC52uFd9++Zc1
plZq3kHGGbczWow9HFxxNKwexcualnWvPGZNYGVz6kPa0LlGfh4sInxSaszsRh+w
1MMK52A+C98X+v6RAD95KnF2DEi+cQRy13DOi8+sL3LQWJ8QaaaHp3NMXmyPQ1H2
r+Dl0uBIudfLusrXag7uEg==
`protect END_PROTECTED
