`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LPJKjb5YUY6+3gL17qxQ+g1ffYQN2yT4WfgzGdMEycLBJljt2goS6eUvmhSNs8eh
x9NclE28Vy6Nk/xNMedt9RCiS71vGG40bArFKTwFizfedIjBiZDtEgpGLjRxG2F/
zPe8Gs0+0fiot7d6gUnTh2iy2rhDyGwJI7trNy6+GNypEZslFyEb6eVF8CiPju8B
nI16Xj37on6mRkUe6AlhenFZmRqXyCfeNvefeHJ24OvCw4b5P81bNWA7vxSD/QqG
VblY621PDMLqho56chO1ev1eDd3u9FrUCIyJnp3DD+RW8kBACN9TurnlhwClgAeT
doJi+k23Ym8aMZKB25FLVG13D1WEgZOboxhnbJND0DPBaTw0Z+CrtvEHINObeYJl
mKQuZ04Qet0+9S4kk7M/XeD6JqbFfiFrbGZpN/oyo7M2UDzzVLiA4qR3Ia7NZRlG
ltCqLo++paOb6Y1mxg6qcj6C0A23Wreus7URfhLhhh/+nQXIJ1iDzsflD+8tkS4y
swAr7pypmkre7MwCEt6aeNMbzblnYFQSt4AP3SrZh+Cqzg4QL82waQ08TfSXTMW3
6pP2u+kvMWi8+uDHWPmR92dC+rTotIIVI7TqNHdn5yuJyLjTObd6P2OrRKtvStIW
JO4HjYdiN1ddNTMSoJcs939BNPmDan5le1m/yNf0phU2rFPxVe8IuAv5w1ropk/9
a+Bbm1s0g1TFE/pk6ItL9QP/ND1S+7BboQm2PCWL8e8+hzb6MjPO+5H6Bd56udCu
FGY6mEC9hm/KKjEsQDHgmachqzIcCkVKtnzT/K16eVIt5F5MtdrQJZsafIfTZLi3
dN7uYhH2+qojUuhg3htVFV0JYU50R+dkutyAGVByO0PvL9WMoTY5WrVFDGOCk3hx
pv5818mji/+TW4TaTKyUsEBp6UBMCJPuR5ldobQetVvPLRmfhI3n3Mc8jaMqFT/s
EyMwaCoY6QmXTT1JLApcFuDRoJfqeVRVZWc7q5lpp7VlRndIUBxZ4RIJD+Guzp6y
70YW/OnSJ+F0ky3PdqUfj79h9pOz34DaTFuN2InlZ2KjF6AlGuIIjkrKJZgxBKI+
ESuzNoJu9MGjgkcFsyUcrkKKq6t7wXW5QXeBrBC7hR5U9bfcXrpmmZBsfkYq2CSn
PAdFUc41hV2N90T260CGiu3Wjg6IKrnFXLWhpJuASNH7Y/71Ali96wNQv+wQjt/c
34KXW+csRE+0MZLv+Ao9DyBelHJRaYDaPAxn01V+BW9XurgvaEDxqY4+803laart
8oRbg/++PDbg12iVBDohkoYClyk4P5OW3ZFJnnwj/90O4zSYwuV7De1umZGmTjJP
CklJbTfPsiRlWXEtdSLo1WuTi5MgtSaTO7XEzx3JyvKF4k7xYpJd/l2fAkXCB0pH
f7tFIQGzjbwlc+zCIDdsqSALVuwnUwkh3ilRGAiy49D4Wqx41PVARQEAx7SLT2m+
UkP67bC+XbMJ+zDCkgQEWGHpJwhQnZYdGZd6oTjcmb9TSPq5VDuhYGgjCwU09Wag
5KRg6a4+Zs4tOz4Aa2zLt6uluEGUbXTkMxSo9XEl2Z6/LjsWixjUCCdhs4DvrwZ6
URKzlodiFo9V+kWK+kyZPXmlSlg0XQ7Yjd+CiSXLOZHc5YX76YU+1zKvkJnNUYb1
XjI0WD8HaqORQXMjH+LQji5EViPbcskSHKobSIG+4IUUe+nHW7v3IWrjW1T1oyCm
mTUWQoi8op//Lu8pekeESx2h9kpSlYs3rLdeWi1wxzFlzUhcNf6fW+yV5Ih24RJ7
Y2iRC+ABYoEUe4QSqXe8UcWZ0ud14rV2OI9Nt15id88d8QozpWNiZJeFv+F1rIz/
P4Xbl110V16jCOmtK7jBLRVN8QWcFTPo+daMCAoUIfDZcHCXzrQoJTT/u0QkbheO
3Djf1BIe9asMw0YVnmvk80sY9CZLXaWohRMCmxe+WoXSzK2m5dtjmpRqKU/sBeRT
wKOLLTGfOg6DumPz8DtmtMa5So+qjNBat8ogj+0vvavfN7qKxdWq+/8KMu/emEdf
5k9T1zjowdwPaaEQ3tc9QfcR42suVxiie5Yj6QTq0ahOOHBCjbgWwHJ3Tui+y+/u
aGouTSscgWgWmuglyruuS1rV+mUv/ipxdt1BWqh1nwZgvZri0wINI52W7oYL1NOC
/7yTc704RirgX2vET3argrmsi7EgCNFG+ovq0g4koiHwi1JiqT3egkHW2zS3CH3W
N6szsvIjqU4EM8Hc5B4VP60U0VJJgYeZj5WHrf1VLubn6Bx8ZR53fX9Fojp+jW32
v54+E3g/4E7x2Hjn5wdYJ0LbG4TJ/VJxRJeqTCp1FAcH574zLwOeXPNqOJKOwBDF
kVjCKrhEN0iuQX736N/D0A==
`protect END_PROTECTED
