`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
H1VRLx6yZYS0E/9NCouaIQB7cxuipmS8sntjBMkacPLpXgHxj0bE9IS0H1A3+8m8
THQVDQAksPXtOR+wPR1MRIOhvBHmclGwfWje9sZhjK4NICaqaKwZZmJ/niiyq7jF
BSjGk/EekAOYMaC8We/k9FRnAmcNn5uwvTkYr/GmVnfnk97eiJ5ZpWGTUgJODz+s
rI81hAS3BDMJeZ+k+4SPXITYofVGSfB+OeneB+bEkVmjH3kTYURq5aBguUMMi3w4
Nl878nrysh3f4OCDJ7ACtoJNGy2BArj16TxB9/aTaNeoo8S6g2++GQYLI4tzYdLr
iZs0P6u+rzu4xfsaGtTfY3KAqKxmMJ/6bOSk4dxYtFkbRfJGtzR3+jOUHcc+3JfI
pdUw+5QFPpWNPFZifaRMU9r/I2++nbDKYY3B51LVrK05iY5cXdNaMeh3Nd7WPo6t
cjVDp6bLwKNakVl5iADOgOxmDpKA6rljrM7YLZsABIc259i80XLhZPE13xezxRmw
Swg4/cyaEAh2YgtYaOIs2VteNnQBTwRGLSJxqJcjs/jIEZKY/q09aTL05wmU4iPI
dWqxQtFZFnuEz/+3NmXKWUkvsUP50mxVxxr3m5nwUNeqL3m5wHSm5SL8iZhiddLi
k07FYJIwzOZC66V7wfgfgqU1V/kHVjKBotaYIZHNBgQ3wErhFuPV5z1GxLD7vhdO
SchEZsGgIOQY29I2IcdvKqQj5AW8Kjrr1f8NC0N4ZLS1sQfpLvklKpCqfp8+lZPb
iYl7C/mMsUJDjJTZtLHiAA7/oHIGsyuRf2wMEnYF2RBhA+GKlXezI0U43pdfAKKQ
Eb6GNY5axkKVHth/1CWtbfh4+bOY7gGeC6IxqEKda/fkcptGdItxNkxhW/ffZOxl
DBTx+57Cc/US9sOTk7/LgRsoAHwCKEs6LQFQwqnUMcGWo0f8+TunvxQ5mX+UeNqQ
OisI463p2XmV/YYmcO24qqsglb/rVcIPRIkKTESVD3OmULZy/oX8kPmxZbkP85/2
ga/WIPvx5kyGVSUDTBkvZIx/SESPw+bIaumUdkyNRTUyxrK5xsVMJGuL39KsyIWZ
CtGFQZiXF+zWe1qJrDEhUpHzq/WpvO/vOFseHpeG43t5lR8oFwL/hj6p2Zo7K0j6
MCdLoOLhXOXwEOtvSmoTxVPJ6dfiH/WPt7OEhdlhOTrl3rtUntDL1jqEG03yhbsH
VGdH375lNg7/xBTFsW5Nt/UIn2RqigEppmMvH7TX1Zx8k/NLxay0xSGCpoQtxJN+
YiO4K1eaz3cxCJN3IoL9R++KZjM+m1y9k9zJsdGuCdrJSGco19Mcc9pbcCWhR84p
ls0BZWamEUs63fdiEk4B8LReVt8oP+km0qby3zLsiUh/N5p6r0wFiSjecGNkBYi8
MXPn+X2YNGRboFdAiAcBRkrZut9yhUjZ92l9urwbJ3m0UGaiJS8Lx+BJD0jtnpvA
/bDtr1RvRFXZkNz3B6pt3TG+WmRTMyuD4Vcn8bLVP3BDKnSoGxrPZGrxODO6roZP
oDdva92pHP0jgGQ93A4nroUGw6wzyEkTWpjwifU2K/hbTxjwjc6y/kxvD5kHDico
h3MwIc/+vH/ku+ePuXDErqYveToPgzlKs64ymo/LBMX93lWWyLarqqsok/z8NYf8
oEv49WIr+dS6OXfMiG4I5/77sTt4c7HRrCQdfnZeEMjRM6IMAb7Ced9iWjcO+oGS
CGqTt5EadWg7Rw894MQEIBvrm3EYfWt3UOyWImMxoQ9TYubkyX2s9TXY5eaVRSsQ
VtRZfuuvlcXIXuM7e1z4iTxlNEP2U2hhKWYUjaWN/C8xfuqG5CM85pZa4iemVSLH
89SzNvyBG0EsHxgUP9ZnWeKXvAOuo6+SBNBAq+6p/L8kAPsF5MFN5AgDV2VVvJkd
S0UPGH1ea8YHSyh967x5qEEGZMis/rU7dgVf0xI2FYjkmKsHKMVd8IyDs50A9yDa
Lrp6EczKzo3NVRz4HQ23BuExaqIFxrZ6+7zLrkSDKUhshWzzx2PPaiGImqf93Wqw
Mk4Ge20OdZ27qvb1ukKO8GZmEAHH1gd5eb504q5VTn/+5U46KCKc/nIPPzMDu7Zq
JVlf/+IXSfnBL+OdMRfIO/8BTP3k52wWc61nEHlkX3AS+3OstG2MoEu56xywXB7w
jsBd/JGHrUbrOBVT732tt2BrkWDzjGzpaU5FRi5LiaHU2HAGo5ExozLNUqlPyaIe
UUqDn0Mc2KTA9IUzf+mpcpuACdLGZP+kJNFSc2T6zdk1LPXMTmRItTk9cIs2v+43
BtDdUEA3L73JbbTTkDv9Zuu0esxVybz4961u+nooJbJsvB4h+fDiOcva4f4vxBgu
1LT2CGE4ErWZyuYqBed4cwwwuA9Dsljp8LA8fNkxEogT/UpkpvB0SJHwxP9etwje
4BMuEfLr2vI1aO0FrfY/pkRywQGvE+YI3cUSZa7oEmXVG1tN5Sp3DywZ/3xJvbXn
82ZFnOfKLX8AX5dhj/XOk/fNFOv/7KoA2h01Dt7oJL0xNajXjERrESMTzEqwkZrM
icDtM/5vPvZGx4MYdUzaA2o/oZPWOAXAUvcOEYaJ/bzf64S4Ko8NERxWS+9qTJ8j
ebtRwAjmOfKhQPsilVldLnoNCnkxJ2ZLP5jvZ0+VY5AqxHQ/y0eIaE/hND8KgAuW
im5feLtk0xpdkBrTTpfSPmddeuNvNGUWu527chbAKjuyZeyXV3qK2lU4iU8Wfj2w
X5PJ+jJoXsWMz5p/0FcE59uWzagmHhWdRw02AJKY2DuPqXa6XXJGZu8xvDKB7W1T
ZHbvf3CoaYDjgF7cgyV+5+PAlvGdRMJJErjX6GEawSzev6LFEaw5WJzZLlxMGjYG
zyBhVR7E6p2AhcL+W7JK0FHolY5oY2oBBOEj5e+8OUKZKX56tPUtvoFFyZyCv+OX
pl++crVR6zUnI5hYevz/I1NadWkGUTL9DGXHuPTjUWWxDBOnkggCv7o7n7D7gZFe
Eo9c2mqmm7JnFkuy7BIgmkmFLiOzevEGHayB2dkto3d1jVzJQOVPMM8HcEI2TGVV
N0hmQWgCxz5a++kP/WJeG6WNNx55KhR/I4XJPNoIhrd8Pmyv5J3FjHT4hIMWjVa0
Jjb3uXAzAhYfVWvhprz/bpIvg7bJyXEkXvryuuFz4MmCBtTyKXrk2aMgB3jEC4ZM
AAnLmEzEWehB7PgWgT6q489eWwD0bCtDKxosLFnl0byiV8hz0TW9+4Z8qvI64mlk
AOrExFiCG+Yrdb8/xigv/hqcNdbdbj6rYoc2bS/cvotgN1VhkottOX2CKZ+LSF8m
auObASIf0cPN860WVI+CvBoykmdA3h6VGEOnaXNR7vldRadHsIaDQnstvaQ044RH
sRRyOwEvnsCFMq3I8uDY8mL5X66IMgjV5vpTzv6kh+lubVTeKee0m93X/pj/dves
6Ib/iA2B9rcl6zsb2T02ozMtpToSRvw9Ln5jptAvt/F1Jd0hgRXaWeg7aN5pdDeo
TCFIARsyk4MnkCUqSHeOb2O6z0R0W2r43Z/poCWOnpyAHT9eeNbIQBnDZng+IBR8
N1deH5lULf9sUwEg3j20QoDnPYt/KSU9bVnw3vOd9qmiL5V0rwlctkGxhpAepdUW
e6TgIh7v1dyosXo9nSsOzWMwWgcQtluJ1+GtQreeNpK7YkdtvdHxpsOGNA1642oc
h3Pm/LopJEXBePDJzZ/ix7no/YBX7RCpL+ictuyuIo4FcjYKhXs6fxmnAIRiVzvq
GkWUeDJuh3hdO7bMcXJR7zvYKtXVyah7JU1JYrjk9VTBIbDAvDDaT1ymMzGacffQ
OTHC8fuayPua9i4ax0jGWTwfbxJwazQGGLaMyh9WJxy6J5QE3L4ewXZaThjve1nt
jm0HDwbuYVUifOQmjjd+PAZF/jmSa5iZ61EV1MApoSFIE6woxKi3P2WPXMr0udbC
3U21Indokp0N7HBaFlffOSgl96suaC7Gem+ZFbzNnPYfVHy+fh06FphTaReIcl13
qQjGMrn4fEwtNOyjq5NiQbkcKi08tZcBLmXwvU5J1y5Vkdx2AKTZarvrEs9RzRtp
uthsBGxjoNfsLLkSy9n71AYEgjdtjJhFrAzS8lss1ozaev1R4ccFZO6Aml67M0nV
q5EGQHRvehiL6FqFqZuqrgYhfOHYhKd0k5UcBMztMZo0+Urmz3oa71dKCQAaBeI4
G/QfoDxjDhpiJrvQRNFOjwWm8SBtqoeJW/pFX7r/IY0y6KPAeuOMEpolCNeZtBIE
0TkbK8WY8psAOcl7wtn3BFdjjIfs0QTVqAWpIXFJ2idiHa3R4YeMJ9REta1l5H5X
Spd5lRqt/kpP6JtANytBhVwnO3zh7XsJsFw8tBjs2OwzZmEXAlrSB2gSiXXAKBhk
RWQZsHscJpDBtd6FER0/jfKKJE400wOpVo3YXjYT6AwB7Bxlz+B2lOfHY9ay6fdO
ZIFMm3K7dWIgWC1CwCqUQOen+pIQoEPMmGV+wsG+/RGciT3rm5ohUiEaBMGzkbcO
2LUutpA3LxvUe5fmiOFpzIwbXEPOtnwbRENweyilOv2oIlLu8Xx8MCaLtWZt+6OV
O9UIV8DtrBgVfYCroJ2qsCm4bHDc2lxMOkfGEiGc4pntSX82Xjrpgihjz95kDIEb
m72iznXQb3kKDs9AzFcQG4kjP0d9f0W9BfxcDPhVKdcbJiE0FusiZOej7Gr1P2VI
Zgs55mAPgRQHlLz7k1qyZYCAgGoc/X736MkLeuVipN7RDOnOVyLYANLt/1gkb4st
tehIpyd1QYbcW9/VMfB+Ybbr6Ot/jqtjMaCjxZMyFf+bYezTeE5YjfO8ih08fIKu
mlGPUyCe3PIm8he5JI6HN5ResnyrrBAlhVFta9s8TxvGQSjHoPVo62+057L9dQPH
OESTwBdKSmM4+ADA3yRQBVMRDq5JG0W2020syRbsAFlpN8ThUpxTJSajd+63ytpb
kjf9X8AIxVNv1yW+dIs3zQFosb4W535BpJqvDWXAb5WRIoXdOUsOlqRM0aviwJo2
LvR57tuo/79vbgNBqCpQ9T7St9iek53/VQKIujA4rmf2eQm9nKsQubABkLspW0nq
fpCvmB2xDsgAo89TsRGDaG3xqTCsPF8JZ8NFdtq91SqFdkFoVepPQhC5tChinzVz
Ta5BN46qcNdRhOPSRe+r6K3+WJmPl47Jg2PXPUQZ0f9fX8n6/qEaycHiWESFSbJE
ynqx0nfdTTCp6j8/3k+pOuuR+mLjMfrzXw/M+zSmb9tRZlL72CIfTlIVYKzgIREi
jowRvOnEIF8Fm0u7DJugUEw2kNVRHqPF14fr/pi4QsMoz5RBqWNlJimU+yxBVUWd
jGmvziV3Rbts3WxXAR91MXdmgawvdYhj+XkzgAQFromBk9Vj09w0uRlVvM/gIeSQ
Cc9HJ9RTaShGfJnR3Lhr+cmUG9nQYUaYh/GRk9PHSUegYwwHGhGamLbqDuSTl1by
Cw5mRNzkc3AdDL3d3FtE/8bnUW2fSEepxh+REdGltYPgTw6MmoqHl5b8mv/lFEYb
d3FZSxRqa3wLY6x8tKpDKKOBdAWcdgEFUqUCSikYtn7E/fKEIMZSilYv7BgZd/i2
Cyr21C6eLBXDQ5i3hyKPRZRIaBigt44ozhDn3bwFuwNE3qZPyN7AfHrT+jQZQgdN
51j1L44CTvzXt/OQCiNxh6r0Xd+TD/Y4DYcuS0mB98UcV4D5xyW5Pq/QlGpHfl3F
2pQVD2arKAdmjUsYQHiEA2TI5bh4ULDfFJ2SEXgkFsDjY4YtihP+zb8WUJ8TqnU/
9kk95vhTx4LUsKcp2kUJeVPDQwuIMLPr0ClOZSUfCElxOG2ypzZM4/XAkzSZbEf1
rcF/8xNn2mKLc+6rxPwLO4+hx3j8wVp1jXE432Xi8K0XSDvKFn/d4bxuDDPqX6NB
WmBi8n81vsTapFYPP9+OP8v+sxDuXed1hXwcSQR9Xxdqul+W3xyQtJ1MUA5pdjiV
0ErjXk9tIl4ik5AoXpitzYEje4p+jKulS+wnQ5Y+Zj9ES5nxtHcpoKlLOxNvgwGj
+KHcCctKXAmTp0ApeZ7V4OQ9ZL14gU0Tn5t0ahK6CdHNy+BFiFiMRu8Rn9oaUq7L
gVR5S+POo3MYiFz+gnRXMT3n17v2uLGQUm8x5PSuC/SAEWjqtOkV9yfb2f2OTQaR
RMb9jHgNzXflULKcyejlL0aEHSZ6n+slUVd0xxn0dmqDaWNgGBCAMdnyW5zXZoIL
03F3groQfTfrgFKMSxJ1o4SHwApoFBynjZJ0aCbR5+Dpt3KWJgVrCgidN38mdXIh
1uB2cR4PFBgoyec8LtfpcPp4ZIrgmfLyFZZ/ZfvMscA=
`protect END_PROTECTED
