`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WaL4P7huPmU0OIW/K/naWaVln+rS+DC6k/r0Tx4AZ/vBFvUapgP1wHfZocZAf4j4
ThM/toRhGFxrD7incePZQ694NEuu5LOEGUn7XYAFeHcKpVM1dAFfshT5n2FVWoXD
t/yD5ZDnN59RArSWgZcjHSS9MuW3Vf7Wbwg9LtvOqxEgGFyMyBlHmgQ+kt9rrLV8
jpXVEJW3AzXPxaARm5IvRJTFaxy8lq2yiwxdRlT6SHOo8G79xk0gJHv29rO6blxi
ucn72Igr9XThtvonH936X9HNWkHum+XL/qUU6ZJIHh4Y709a3+y2JScBqKxemln+
0Tah/wZhbsjAR9QN8BiShB+t71M4vd+1MBHQaCEX4Ev02g7RVVQ57WLNzmjzc/RH
4J6zzIDXKzx6pKc5f1d63g72JiNa+YMiMpnAldZUBbJGzydfT5Np8csFtfP1t6JE
3e9Gz0dcgYaXpl4enkMIZ16l0zvmodPmOAC2VhV5g+7o5juxylHg/fh7XFeq42PG
NwZgXkAbDTzdb/CyZR8qVtU62b6qCeMs3cztknC7j/8MUSdgji99x0Cojs1G6zIb
Y4GrPc8iaK/lDnBctYtkuezhXaDSGHNl4gvg8bKxzwaV/6/SPnsVmMVmF18Ej+yj
vZZ87DfjB8bY4zPLoIqVS7lJBGFjrDrrUHAhLkYF/8C/evCtXCgzQiomFYWGzLI5
paOn0S54+JETxUywr/lubcPHKtumbfSusH5VYguu38g9Z56uIy+8HI7bHaLayzXi
9xJ3y7nDWIINmgudsplBWYRxCp7GmH9gPC8jOJjgUCPlNInI+FKOhTYLTx46CaCz
kXM/eBJsH6GUN7+DNxzRQJ6MVVl1HglH6Q5+rg23jIhktkTmwC2csT2JKSGVeXCf
KnuKdZc1cuVBPIwzQMV4ezMIzralutE7amtcw17ivp7phxtYxnJTQUzS/E5WXblS
3+s2J4sAhAcQ1ZdrGgbv5NUvKqWvdDhd/lgT9FoZ3pS2zBUyHPXuozHoDfJrMOZQ
OjYwjDxUPcOfzUjtV/93ltOgt9s7V5jJdSPJNc8Icse86QiTx50YLpHwQ8desLol
QabEcz1Y9WJsDGV/HPgtbkmVVx3j13ecgc7qKCxme5iqi1MU4acTnB5sICDjlJeO
h8exWBaUthgiEByg2UJ7zBsB1CrowdAcAN6o4htYQatvKuVcHvuKM8QVsCBQ+LEw
4owwsX9qM/kHxhrIEJaT6IFbqPNaHZcvp2LM7BFXyLB0l6Z2OWQdt87GW1oMKCjW
AnmS7ZP6IqWXkAQJBa8q1b9FFXN2gxEPWuLQHL2mG7Qnq4mUvnt1klixD2VbZpfW
F84k+q+UTFKlgjTFLaPgFQWS4Tl6a13QCeLoYDuMidbWNLWLKi6IS4N6zxzjbNe6
fHOG1PstGAa2AYR1ZVx0+4dLjXDF9UoEDYX1CSv7ATuUZFlhh72aocbiUg9uh7pk
ddgXjI8VLHwALprJAKIeDUJtaYlaO+EQ0MRjeEsWNHWTEwIbjecEV4yU5en4wOPl
NQduAOHpevWNIu7L99T+rRxFEhv0oIKH43LDlVOLyjx2NOp3lG/3TcnAwEQMxeSy
UFGxDEdnRN5z2ZHYvKf0AJxqY6r3CNOclr66OqJ+S63fLDn8tS1uzoP2ewGnWS2J
+6o6dHQn4uyDLNVGvuv1xV0958llgrRgO1cZPKGEWjpvliSRkiU9K8GL8OZ4ixbO
5F2fTR4UI7VAGeOv3+YiOP2X+LE3SVWOfVxeq0qqnqfRj5rJ4v7B2HbY+t1GbK30
QdgqGDH9bQ4k9Ef74WXBp0Dwsx+rC4CtDSRYQLGXxU6i/rj7M3NIktqrv4baaa0f
nU9urNZwDY1ELQ+5Cit18OrL845DE2w7fd6I49IULpOrB6e7q1GKPOcFDNFb3Nyb
RECce/g+ZO7DuM1LEvC7y8LHfHN6qaBKahybQX1DtEqvXl7Nn0SHHeATi1DlUUKQ
pmcBOTdeAXKd61H17h0fWOKxPBf38MTIDxNUJM2EhVS/EEVmSBakUEdkbSMycK2G
+ikcNoPh6L+QwfHx5KTILWQC/U5JKDS9HZ4Q/hBFAMs+XbjoAr0N/9GKko0peFbc
buxJsVNilDj3dsW7TM7jBUifQ2tMkQgUMHhNq3OPaenqTQhC4otFAHFuVz+q/xP8
fFOj0YT8WdKVpEM9AvuSCwousfS/KCW7A+nqJZVJ9RMHRFB5zeZ01L5UHfotCR9M
FUzIM+ZMfIhBBY4JzG4ygV+JICoGmxdMxVsjlqMZN4VU/O0BjHxqMhq4l4+vvDbd
7rXEQUbVVbBrfl/af8SsQtPTsSfs1X+LS5R06r8JtJ5h4RK0YXu7Np3/3aQSpnai
g+4kpBj8gxtOZgqIOWyOb9AsTxzilIw0PCE5o7UJ1CM7OTvX7nA785uk7uZd7j0K
B5Au5/LAs5vwAjzAC7jXKmlzT9bQU0J2fid+RCRIIWbtkD59U3Ztd6DpdpMS1xjc
AszTRe13aVVMh1orMADEzrbsTQlkqqYwDOC/o8/YV1ioZHv8T8Q/6RVDsS9UaoAd
fQglvHVrId/BfyUxhd01TrqLGco7Q/H91uLyDtQxpc/AZnr4eVAdY7griNYKghsT
P+mnun1bGMuftlEihJ3LZgsFpUyl/J1/iMxCd8sL/CPsRvvtSyiR3rYzdCkEOGeo
49gn5eS5muBBwRjW7fR0u2dGKGZTsBKaYQTgubhKkrKAOhe+OeOacuzBUNenWJtP
yizWzmlEvliNka7awRHjUZRfyC9NNJH+qa0ngxHpcCQ7Rm8ok9IyWbztma2VQPP/
+csgxh8rg1epjQCSYQpHWzuDxDqhelo4bstZjBwmKojJUF3kPBZfRSL8JhVrGbvs
9rzOMt2XDf+a9YgPFchd7oxUgXpGlmmt8QMS7cWWXOZc6pnRJeaUgWv0jOmSe/Eh
vfhvKebmVuS8HIgULz+t3vs7SbFO+a018uTdfblJkCqXs0o78BmIMMRQbPNqYNRg
0L8Upyg0o2QyRxeUfReauT1Y8qJ4+YMh5+ZiMfnFQLatkk7sPKFVABpR8jhkl7Gc
kZ2TGkYh4yYj6s86JPjpQ/YPVZic2s48FFzgebd/piadFfMWmn3+hr5VG3QBbCI1
Klw2KDIFAVlkoTaT4Tl4c/ZBw62b0d6OITvq73SivLgcvLbEp1Md5dSc7jswMCKK
DmcnSqUXG2+6vcAr9VKMxgx5TdcP9Bo5SsaeNBlG8AAGSacBiMCJTV3MHTfCKXA/
7fsOuAV8Tgn4aaQ8VpcQS7F3HfNK92x16rjlEdSkmU1Nsyyny+wKfhAS2xbvqcQ4
liw21nQtO0AHHEgGSaMr+2nVtmoH5tGwOs8sde9FdPB1Jq9hra5tooHQKAV9u5ov
nV98hapOakiSn7LoWcD/4hnc1yx686Y7ttcjk/VjavcyxlEx+DN32XVsOmoE6Arp
VFlpOyFEAGdiAEy/r/re7PKFpm+DMIp+Yg6FhyGMZqRYZWt0ZjS97eIjbvYwbrcH
8XjPcW2f50mv/QHA4wIHEkSohufSYSG51ngABVKihcB90D/7fHXiAXcLr4WPwBn+
60bTdPHT1lgr1FX4wRMdhptf51nUKeSwCz4R3DoobVbC5uLIpUR0005FTErHc4S9
4kxwMutANJWxQIMlVhse7A1Bir6sNvQwrtHjvF4W3jlK5OM3paUmk3CvtrFyfnvP
YBqI3WEwIqJzVCJBubheS5D3gQSLw4Re+W/Mr5/aO57SfF1Fea19kuiSh6vkr9RG
Oxk+95RnPQoD5UPqDqPwuf99nWpLhRt4xy+UcqY53z97S0hpm8q7WxyRnfz/8PCt
n377XA0jpFGHyglF6nyEmnrdXEGEFkRuxmfmmhxCV3KDL1+ASwGQnn+a4NHuGmxn
1BnTenMHZy4MNfU6W+tbWZD7BdGp4XnKnezkHD8Tws8qDUfp1eWGo7ireZnJZuje
k9iwfgJgsIK3U1FI1oNjTZECzW7tx84c8QKAleGCkdoK/IsLUseyku8f/jOwHnol
Ycx2uGyLZaykvjikY3zyFmA6iGUNAloJYIkXQAv3fIVa1oWKJ1YibUsKtwiMPvQ9
FN3bPWg0mHw1yAnDhOGbjLvzFCvEQ1DRzHE2aiVOzyFLZChZz5c5plUErgAOvZx8
7XGQEstB2m0+24wUonlYXjosZsiIdoO7yWrxhxwGtZvFjyhbPQ/0/m5gfODbufPt
5G7k/syw5pu9A0Xwm+fkvfPprU6gYsOqaxmtkCbQrs20mJvbOGoF8nT+RsfBP3f3
3mnPvwkUYdnIPIAt6uiGh7/Eqsg2PPe9c7R6Qcn5WjlbqZ8dJL2WSbW7cLJ/gIyJ
coPvxGtbvEqsISKvmtDNPGH3Gz6zHaB5upvgkC9/mwWM2BqkxwxXd7HerbQE7COQ
QrnVmqbM5BcURmQYof9fgN7F0L9C6eB0sGhGRRI6zeZDKg86KUsY/v8lgA3C0Eeu
RiLjr2BWoV+/87JnTUzLIleN73gtPU2p2eJJbhZf09RWyjewJyoldWSX+qdsGaSB
ZDKuI8sPThy9M5X7zlGVqeu2AqPk8acX7BSy5bLkCsULxgy+LSmx5T4c0RiGpaix
o1rqQxwT8LzCJKhmhDX9D8g/iaOGJ9XuRKD5lcwesYlh6dXwGGFmTSLisvftVQoy
+xi4vS7FBR2+5PqP9c9AikFapXo39Zc2od5HBnGModBVhNcYx1QOPgHGXf50Gc4X
lRx6numdAR3Z3iuWUe0ZdnnxuW+QLcQBckG/8Priw8QOzFpq7wv6faE++0qbiQby
DA7xZ4S9ZQ1da8DeHLPN25W1R3T9C8FOataPasxv91yOV5uCiGcTm3mRLNLbkw7d
ACvmKHfLV+UoB/nhJtNtiTrSiJypvSjwQOHp+VbBCZtpf79k3xSyjZFv0IQqbKLZ
Pkcd1Xj3o0EsBQeKw8shkp03VcvpVDAq2Kbpo48VHu4A/rTJCQYJ9I5uPfTD8bBw
IS1t/mPSTr2074/XpOLzKzUY3L04LrtaRpP8x6VZlLUVUejRZi/TF0Zpby8gLqE1
+1M6p1Rvaas74fjxbl52J0AZ6i7BsWvgYuTorGLOmG9oXq9zlj6yeNZEsJDU6qZi
CoQS+J+MPdgZ3Px09m5gUQkSmWQ8koFAZMAFQeNfR6F8GnOjPTN7M8H41iKE2MmE
cWH668FuSVOQT1mHYHvdrg9LRlJQSgRYm0nuBPy5Eq1fzgzsi7azVrtAbQ7pNKmg
sLG5G4A9rI/cugUyYfWBrhfvzg/2kAN02P4XStn7e0OH0o9GTiQ8O2oKfDFt3Ypy
XjhliZW6EMmPFK+zSdOjHEfngPx3+NYVM/4iRbqNHEhpcbFwbnetCfezoJcE3kH2
emDJJaFdwWMNFCdKZqMFjztPM2+iHMCpI2k570fOfOrdggO135lFqckJCgYHSMom
+rZNBBGCCVJdz21yw0zzphA/MbrYwmRS8ksoBVIfFUGOkJfPe/GhB1RyBpOfpl8/
vO7hWUKVRQFTMGqWkqjEQ7v/JyQ5WrrSPfvDsDn+SLWFd7G8LIixPCiLZ/v2h8q/
jj3D8Q4P/TAx33ubaRKxQ/cTgNvW4s2NzZ7tNpr/N4zYGIcMit7o9+OxTiGZRF8Q
LvxaopbOtsi3YVRfMA1MQYgkl20dQcPBthnVLZ0YYaqkYEv9smLx9jFS0JJDsBuf
KB8/dE4mVW4n2QPsPenMXL7vk8TQzzGwpy7sshNJZ+GItPQ3uirhsRmCZC6iF8K9
UM/faFKcSnlxtoOEVOUR7i2JK+uu6tvIqZ8GVuwhtewHdCKDo0BIAOrpSpF5BQdY
88IFJXSpPnLHJnzoo4/sK8Px9m816XpTkcTlLohpir8/XvnfxcA7irOoLFfzxU0F
N0DIctaF23Z4ZaNfRWqE/tzs7Rn6FjL/GKhvjTm4vIFzFRU0YjrK3pm0E9EfXXtP
cCoyusoiCTSoOnGEDNGyblROmbfRQhIvAuFPiUoHrt40yy6p7IhtBuQcShUaXOBj
hfn9PcFwylEXhXzlmKM+9whv8q5RwmVp2NFUfRq7fC18qyP0X78TnTGwmsnB6lYf
O+KKX7WvtS3onUonqB/tgtED5ZikIuYXKrdul4K1ig1KLE/h/4nlMyr9NTiwiBPP
yVajkrztj93VOXQNt8bikb3qCEDMMRypcnLhxZcQd4q3ksQoLKu3s4b+GuzpV9/P
oH3McsaQJMpTGbhmKwG8OheMXj9NHQUxwMNYEO+7bLnDFHAEcdXJVOJYhv6RlqCf
PatbJvpbk93PeRFpkuSSRGToiDEe6Iephas0oAl8wdi3s8/pm5bct1yNskYDnIhb
TAVOS+2nrsyTJ0mad/HS7rn0wl58Fm9k+r0DDMtGIAoIWcINB9xcAKfVUiIKyrlc
r93Ms/GPF7Fb4yV4HMA7Cikoom9fv+G5x2Aq4lVWFPjCspCXLIKD/wkutnJV+Ea8
XXtJFU5v5E6+GOxDhJUVW+SDW7ClWn6A+WfCfcb0jxtkn8nT3ISZ7hycKlMOAL6s
Fg5h0ztq5uLPEUaqM+OTectuyJpe6vVLVsEx8ZMWb8ROTm14dUzTdINw56/LrT+N
gOcdoavYvQZrT1GJzhMJ+ym7JRbzpZOGWBbt4zRZ8FFErG/VjbEexicFifP3k2Yr
lpUL1H7aT206GEannoZ/DVIgz3aagcC1JSlcJDi6652CxeoEPs/QaInWEHt42cya
ZLNpxU77KX9e939ArtuHTe0P/Zbbr3hVQGnW2MhBL4tqNMFkQTlpxAh0aSxb6e54
dvNQaRmeMSBk6u/rL7OjQpOdsDRCa9einwx8gsEEnU3vOXMuES267ltu+/IMZiRu
gkQnrAx/J8ERumhHo6JaEc19o281SKhHz4gqHT80K0/jJdz9lmru0ym1CYV4diiF
Bcsn41dVIXd70OSHQsc/UakEKmPOptvdYLFWUco8g/qIthVjYiAhOeTZPEzViGki
2fLbpTogyzn5y61oVclLpNAsKcrgz5J8xi3nNCLmlob2UG+dbgNNt9MZmjk55Q6m
eVQqqEABEuoX1e2K4ddLNMWjHH20q30/GqaQ4DsDhIg/5/mxJW+9U1lDbLclH/0i
6fs32VdYEN2U/bEEJJKf1bpn5/ypSWsSdvg8fkTMhTHf97l+8UW6mYW1xLntIeDI
5QvsxtuFZ/wOZWzl84up6EcwE25JissFTzuiMxQog7OEmn/0DslQ7s3mkk3DoWOY
OuhQZip9aLhkyUB89Zz5VO249YzcNaOzwdwQamo7ax6STZq7CzcCQYgForeM9Gc3
bfBXrfN88MYa6UaCnSQeiGH64Zu2TrxP1PavzRIXX2p/GD58kNjw7viJGJGNbuDr
98vDiwVg+wmVSFCzvWLiuJ36kwAiJxUw2axiinDBID2x1E/CW+MPGYtf6cqgqTy+
1+q+F0j1qI0kjREDwYAGDFdTQ5Rubt5HaOR2WvE2g45jNZmrXZTo/n62MZ++ySZG
cRGLsG9BqumY4A81vqsM88ViPEULV/uGEjsgs+Xo9DXCCJy09BCOChWnLHXg23nb
xBwFvDb5dTJg0qmQPWztjeoZKPfPzEqQJ4Kpl/LnQ7V/HFZzLrnyLVDlYWT8U6rj
aWy4MNXhLxT7QeutoKPIIXOuZrLpVzCZPzM710GLhEhCJIjf4KLUmYlFbc2FKwvW
vaAg0y7azG0to10/MAsTxB0i6JDLyc+tcUHz5Ugt9XtepRqdGHhwfC9u040hOc9f
oR1RAgPysac9pruxZih+W8iHm+IfH4cXErZHrLzVydvQWnmYCfGaWYs1ICaB6ffg
4YquOtYfJIQ3s0005o2q8K4JFaJs7tGEBQiVJub3YWl0MSdm+V64r86gzIIZRUu4
0PJnHgPbleBvhP6b8SmvFrWxJk3PhLp26NmhdS5LKvgJz1pS3iUleOEscejeAl/C
mb0i5/yBEfDwIoW42F5kLlvWnQyvhzNInG3HiqRHCvFED3kImaq57SPG38H0rx0z
i88+WUB3pj3TKd3x8bLpSDE0G/kXm6BZ6x2vRnEC4lI1zpNfL6hxfJ1brE1AUiVv
8nSnsEMGaK5+YvEPN8Y4IJMeN/eg9eNZ8O2znjThFl+agOgosdI/c3fHpK7ZtLNS
Qkh4e7PU/FydShyu8IdKXD7ouKBzuD4zdCNSXxnEh978RWUWvT7P4pwyi5lQ5GVR
ULdb2FmW3AZIptaKy6pG+gHfklYcYS92ucYYJym5xF4=
`protect END_PROTECTED
