`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
w1mRkCfDp3mqCwgcUikKYw196z80iH//eYtkJBrEUrWB9zX8RaUrtAPo9F0Kx2nc
X/eiFziS+MpoDyrBvFfBoEatrXCZ2F6EDjUQIqCJ6U61+ecOmANLX04eyX+H4+CV
7P/KcARJZ96UfeBbM3tZXlSAUGXzcIWajqS1Pgt9CM9jn1tMSI62sNdvrSnNzPNL
6R51R6Q7Ydu78q93RtYrIQjoUEVycRFZHxbcdlFro4yd7ybvq6Ea/vFO5QHJtRoA
AHMepWPdsXMLBsNuiHWaECq10d0i9yBu8QITKUDj83vK7hbx5IJbhIck47iPJGDM
1zNy1MiQ3KlRcdDphW6KK2bDW4AkK/O2lXMPSu5H8Idy99e8NIewwYCVeesnwb8O
sXf4ETOqjVEqReZ2VbYdguwxDtXD6ySoXezJVZ22cMO4bU9ovzVZurtzELksFI74
Uu0h53dV9HmC6g3oXgWkcorZ/HwTk2mc/50EPQj3PQm7a+IMIWCTdArJotLbAKtf
0/G3td353xcynpByTYbOmUY35Xr89ROkUgbgqMzEuXwckzXPK9xBy3/CnECHgqOv
PjgehD5Ht6yXFyrPQTFZHHvZY//U13F/26bgmmiIW+uxdbwUEPM4PqCbLXZUcOwJ
`protect END_PROTECTED
