`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GTj6QHnsjawgp3QfHomQ02WpWH4VeBrO9fOTaPhPCeSenM5sdZJkAG52EeAvaNPn
n3/fSZByz7BUtPu6CiopZDzUtebKjvTgtsyhLyWO9JuSS+IdWg7K3KTe03khYxwp
x9kfJRNMVdSpGCunOw4ISyXmttjW4qj7BcVv72oqpL3rrT3nLpSrdgaGbBlBXWw6
PF2Ndi+llqmP7LexkvE52DWDW3G495g0/tH81vZzlh7c8pthCvRTEQiay+5B9QEA
t8NZIc06g2SMHeiycaOi0sbWh2poBpzSnLze8STn4udfSLsCENRiSezLo10Hmqd1
6X8EEDx22Un0FjjlDC4gaqwDCAm+D+Edk7gwsVWfhW8wAjcBp+cTLh1gShjxyKlm
`protect END_PROTECTED
