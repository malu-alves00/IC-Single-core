`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fK9Mo0bNv9NRllna3C3wEt5J+ekIcsTY7nLZ5nyW4GLSqUQv/gCH6JFcK3qRtGNg
MKBnvLtV/IO03mlXCSANfgbyT3pwJKUhB/Cq1g4eCI4KPHuAXdKOPT4mGM3SpW9t
FHqiCFQHs0q0Z3GmaIziBxar9zugjEv5Si2+wV4KlGWTGxnUwy4Dn/ZCHl+M86as
aG7gZ2x+tM1ysIHAf90Gh/THjunbpEAdT8y5aY5Y/9nJY+6DV8hS47e9Qo/1K09H
3agTPA78DK4QA/AvPhgIGhOTNL9w/PBR8UBankivXlm1bvE7NH0+VdRDZRnM3jcH
BARHA7l5HqBygqzniEnU4EFw0t2YXUe5vkITM/B2zORaApZgFpdIfnOPXEH0rl9l
S/OdlVqGdIfuY9LOQF/DZnNDIks0aU3LnNZJ95DmduNo7GVGhNMHEdv7hixc35Wp
qz1ycrj0sFssUbH8W7Ntvzf4LP+PtokXyJjV2zbve3qpmqgrYnNoaIDTr7c8wEwC
2lkZ5ZJSh1JjzkwD+0YWA+lf4Z+SnIDtLe5cKqctX2kbyaJS5AO0IUGx3+ENKLe/
qUwCfPIsmqQBk0D/1Wks9sWJR6bnOLCjAySurX1YLfDO5Wb+ym/AYMfN3HMmYAcP
iCDtoQgVPvRSdBNTSQEaWdtKVVRVxH2Xdx6qdkGIa1XZPcGXJcofIquvgxOyk2ts
4U9Oj3FToISj57e+s4cXBO8yjBFNdW20z1R3ybwS9NDS73PhQbfgBt3Jql1R8eKL
wvm8OEosonsDaOpzwXHLel5aZY6+lOWZpeVFlZW9fhUtpxrZKdBsek9Ss8K5fJRy
VflZr1o4FXsJ9qHYfckqdQ==
`protect END_PROTECTED
