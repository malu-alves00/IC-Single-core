`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dqQeyMefoOSb5sOVidSMQiy38qIyI5M1lqbh7FrqUZtUd/tP7SeuMBt8iMTourj+
cX7Zy6kx8fvMxZvOmTLDuo7WOMSMJn1uEi3JLmSZcbx44gX45gJFAoAcRzLoQjLl
JOzn52JW4dD3yXDt4zghll/mTcLlqG78DW73Y7b4nX/KuYwsvjR43mtO0qYtnRKr
7nKdw8L4DFz9FrCSJTN+DAC7bUJC6KG898mkKQHSE9+QNAjEzuBxTTxG4Ui1aj/M
+MByd3Bl15VRbduujDAx/AOadUiyy+cljXl6AkJMoOaMw3VjEJuJGiMw/7ZkEaqV
rJ7giwyWQe73lduudLAa1l01M+99q+9gD1+jRrBtYvD1nh6xw+YLj2FRRczB2Hbm
kqrtp2jHKNktESmxJOzlc6KbwYTsWQstS0BzKZFdpsVR+6RiNEfo3+164U3ykQhj
hzXHvt6tNJ+5ERW9GYo2Dj2+VSqZx4GqKJdvRgXyytioze3HpDncwTNWoiNKbIIY
K2/EL5/hNuod9iEGR96gD2z7j4LWwVCg4Yc7VIeSFlKT7MV8L0jswI957ahVZPbF
bS4QSG2ssTndQNiLlSgCwM1GjxlOKF9XMzjgiBDFEy5cLd9bWZzwCz3TiwubN4rK
sk6gdZ8dYPppy/epHQXvij123HeNw6Cb5DDwn6VE1P7D/KpBJPE49pUI74Q3HSWX
UpmtDsV9RxVGyWKVOfSo6osnCv26G96O8y3gb+oNj/Njy4ME2lR2yRH8hK8NkzIy
TMr7hLoCpV/tU2r89YDm71oh3EP7NywRtBlOlrUaNeSNluvlTH0fFu8uGf68vZ1y
8KfAcQhv0Rs7kJrY4nCiraJiKhuDe69dZVL6UkuNwcKfzKHrtgo3LmEeSevDpnaG
Rvjq/iRdNWWgvdVlj6pO4NemsC63khNUzxVoWF0ErFEMi1PPkFIsklPzWxjRRmOB
wbQo+gVj4PuZBZ8R8cZs+bTSe8OfOLEPWSsf9Tm+/RWmKkhNphVl0h0HCERyKb+u
u4ONWIIdj44zv15IVY/gnJi7C7YgdjSUpN1Ny/fml50Wvx3oADujBLh7FUFXO7RJ
TUlFJVnt3yQ27BfFGxPAlp45essHVvaVzM5kHHUie23Tp7pHkUPa4FeUjq2e+z3Q
ezhXp1GfdaNsYt3Va3awbyJa1Xs0ZngPYMRnPO6o4/C+l5N0dA/VkAhw26d7pq91
cr0E3Y3iHGER6UT8COqhTiecIk42lyzGQUO1o0hwIWNwgNZXXk6KEd77iwwhv6JH
Xu6T4N/ysyhglIyCUl3hGNOq5KtM9GxtdnOLGR5Tb/NjUGzTSJoTAdRhkV3W79PK
MSnITfgjwE7GLv1jyqrYQ5umacIO4NsX4J4uPbDWKLu1Q68S95DzX1mCFMN/Vm7/
5a3mNReyG2ra8iFNBXu0GI79fY6GR28s1lUuD2ZvluD1Qiv+66seN7ccr2AhPlwH
LtbCR7PwVxYa4yitgltUg8Gs8R1CQecdA/i2JkG6yDmZJ3DCoW/GF1GT5PjP3wxm
TvmiUaChELkI4lu2D2hKBPnjdSDj3Zz/0n2Bx1Z7HlKTIDbPqPoez0sqF+u2okh8
t9t2sUesE2vWb6Cs0gVVMlTB47bI5IahlstHYkuSdGvHk0h3J9LcU4DejSpDQ+rZ
ZWvWttGmUIizvcFEEZK/jiSFVGwJqLP3eZeg+SD15rIn0OxUJdSiltlLeniJE3En
xJLwdlM+usmZhDFK6U0lt1HxtjAdZO/l7okJyP3Xa4pNysBsdCXkuKfk9uVb7/DB
EQs41P6ZQxomtfQOVQLmArJ2Yn5DnCn1GT1Gt71Qpic7LW4DX2tBWghiD2K0i7tN
xMNUxdWmPOFEe4JZ0gy2Oo/pZx9RdyvlvgDjf578Bd8v7LY97kxpcpmW1hYnAPTr
oSqKGOGOpzMSzxODKuhphsbxtX7Z72rSIbpo8dzrQQYYnEOcvSecFoiYl44FQNRV
YeeuwLazIM6a9ykrFoHLJWXoplFOJZsdNZDK42LBpOSb37zI8UMTJIXBgRJv2F47
kacDQF+oKbqEH/x3TAvuWv+1EN/HUR+dt3baihfOor/MzRcfUZC0QlTweWL8UPU2
WDX1gY+nhqhPM9p2rT85SLwg5t1nuP6jCPX+2mWy1aiH3r8tJmEAmnbDd+LEwVZM
zyQYOXbvL4WQBMTuvlJYAFM68EL1xEJ3BjW3w7TbiqgiYdFgrDyKNhDa9jlSu0zF
vqw0sV+4wSXxu2raR1JexMZ2CtVW+CXrmpekVTbhY39wLn6atblr0ue3lp8hJygd
3fJLCTXGCDy41wCII/3MyJeswTCLMz5QruG5IHXLvFnJpOj6BWjPoxoodaN2Xjbk
OUsB0/Vo0RUiSiiquJ0NT9VIWik9DnDAZ+UlcuPge4543x1q+HW/QDg9ne16+by/
jToWNt4Qc8znRxyOpWwqC6Mw/+ejf3LscJYEooSriE5IxDCjtarqUM/GRsY/TTjl
YrKVwIIV/OEiqXMwsAFbtonQqdQ44WcMAiH+fU3S4zkhjF22YcFXKxrYZjgW8VR8
f8qg9SHOLWH9+J9aagSy2YcSeOhlCBNDaQaS7K6+Gb3hD/sA7MePQ/mWg46/NlHm
EWtwL9qfYzhQZZ2chGRosnzTTlu9mgLwp568X9prNAopoGoW5WoiBxqfNTA3pgph
L0LhzE24tPW9bhYKhh6NgHcxR7Q8fGPCgpcDErvRFd/qlxWoTA0eB3sV6MdnWljg
EWQXLg+I1CvWMqwR/qo9y6ryns+tx1s2c1wRcn1i8DUomuYBbQKVhJFg8T3Xa0Xr
krVQVG6PoM7/zGV+B4xEewK7L3XicBvUvTUXxoQsd0FMr6dVzKjZJ4S1tuFXBOnC
+QjpWKQ9usUVEHY+HUWnETtl3dkXSNlLFSJ/CFqc/22gP/2uv7bxQXZD2jIoOcn4
9ApxytFGmBVm1a5NUtYUbCl1PXtM/B+h/YGIZnu3nyeuawIwP7Nh8zqeT0CE3ATG
DuOI8w8GQqIRzFhOtGB86otXFWI8hKwamgsWM7C8tJcsZmm7Drc5u2yy+ohJLyx5
Nb/bcw6KFtnxJg/2z28mIX6hWJ8fyPJAdc/ZrU14YmIB5bPBsY4RquoXtGaUgQsn
/AY77DU6klhiRh3QIfk8l0RVBi1bRfpgrqexEuvZu4g94CRWX8bZTHpKW0nZi3hd
szvKKlktObpXaAa+XprmkJwkg+P0nP4sAiK23HkwZQ97SiRpTrHZYjG3nDzUqvbx
Hr/7fnhsuByevOv2zX9kNVR2SUOUijfdG1sAMzKamg3d8gwpc3lIwRK57Wnj5hwt
WiIbdUonMDucj6bkHwr5KpW0/G1Ypl47ldrgfaq7O1Qi+hLvBDo77IBucvrf+trR
C6ttBS2RUlmGBffixJuItRqCSbI2V7HVtSB0hyg4HTly3eDQO6kO/AWkbpma26eu
IscOT4xk6CfOENz7NNPO881RXE9SuL294O7t9lRmnyllfKKRO/piK57V61+vyWE7
9gcielf/l4NucdCqBi7fbt0Asg9K0Zy+rNDsJa6lRkRApBQN5/OorEEe5SF1laZ7
l1U+ZIXdfm/ruypxNO+DX1BIRBkBFjrD4WQqrYzQb1YS75/Ey9NRtyAxb/tYp9qm
hwChsNOoqMeijJf65NLz6hgFbxlU1CeKvJx7mVFCtXLxZiECTpsIKiJtvhl0JQpc
DWFt6El37zijB6ShmN81yzkq5FB4ZLkn4gbmd4xs8kokqzll8vuAmt8K7LOo2AAn
iJFpkileBL0LJknZuoFbAkOFWurk+qohX5Xsl2frrO1xUblGbWjlXZ58tQOimFt3
gDlnzzYP5gJSVMIJkvO6pLnlmwWuiSqYUtWV0Jxun2IBYJmZi6yDxPggY3AjYK3Z
XV301UrPBCSblHNotIsFCirxNEL2swSWwKd7nYfvy6iF329t8hcj0hAGe1LLEamG
c2FHqFvCNbxejBKtRUd6tCoYAKyFZmcIQL9NjCQj00cZNBeldn9RH/mLR7xJMGvY
19iyW47SJ00pl30M+Kpv+flZZJbVtUczt1Exba4RvRFQTDjWov5fb/oxMoH3GqTX
YoQIVh200MDY7LOfNmGJb/2KY2pdaiYu4k6sX+MOpKZCIcicKdAuaiUEJo001Oik
F9RicIB+ZtriPTYhRH7BTEr8HrkwwMU2OalnUJXYHtCt7VqPAQZxRUlTi3w70iGo
6kiR60jI81Zj8V/T9z5clCbfILULPWp8p+rh+JFMFE49t4gu0hPg2pwAuCP7W/ty
keBzVnU/8USaDyzYuMjDExVHfz3yICFwJ+NJth2fI/U2TeHcbLW2QuNWQa9jGtxX
dQDu8F8dy52oiqj35UJtmpmmPgpuso4p/EuRR7luBYHczwwghvgQVX8a9+JuCIWt
qR1UqukqH2fcdfvQc3Y0Amj/6AyDkbpRUgJby0ddDdyWQfSxt+hddcbiY84e+lkV
/nNlB3fKxhnQAXFT9HipBAw3fWMtv/cgxFzl0gWPdxP54ifoLRUvJKA2ghVRAqMU
e9XCYs794hpC715IM+tVlddc9i0M+5yaUmNivfvF1woy1B5hDqzvqacHutpKFtOu
ivvpv6H4riV8+M63qnOnE8wPB1Vc/PsQqrL/2pcynlV/MIByaIVzZwAXSHsZrfYO
AbkbEXlXOv6lBZqRZgGqksnAC1+kh5bjAATcghVont6msw3v045lCKF9FUBCaG6I
GhOMUht56QQ00oOazBnUzro7mnD2KOCGUAQI2DkHyS39wnvNxMaUWghF4cPb2jVF
pZVglJWc9AfHrGN+u2LenvOldixUAz3mPFRutf9HT0V+5H3a8ewuJpPTrXtb+ply
53F3A8fU0MWM2THNhYvtgxKDrML6e6AWsyueZpy7922FFw7uHqoAqFtkO1cvbq9O
JanR7fJHpfVmLzYMidBAlKB6/ZqhKpvAK0A2qm4XMqK9g9w10l4e2qdvVoQAFrGu
XaJFM/zkI9wZ7jD5M6LuHONjmOd5r19X3hsR8AYgRFAJQW6TBQO6dzRdXpBOPMNr
30Nr1Cy0+R/lLm9k18QMlgQxa877RcxUkK9u6mRO01q29APIHhFKzgCogKwnMazl
5XVJ+8DIAq1BBJJwc0h/3X4B+lZfrviy+20Xs/tJ0B2BUqPbO+uRd2aeE0KZpZxZ
aQ8qkbHeZi7I+YSgfyMTNz9W8a6aSoPaehFm6ZBK6cCHdYzLs1YxoIoO99o4ihrX
BnSe/3Ls0R7aJOyCzrhDZdCRvehETbVmunSlm14IWpd1WJ9QztOOFitbJ0RwXNlc
P+ACQQKWzmSEqiqHL4oY9ImweHrEqoa0XD6D6vqIhV8NxaOOa9mduYUoQsNXrvv1
nGaBG35bfRY4jQeb2jATIWqiJ6fig5e/O83906UW84Zz36PVd3YsPv8HAikSwu3d
ozmLseutWdNi9c2Dr5ZVybralReY6sYhZwdFEb52M6uxAKyk8oSjwbNVrI//lqZ4
KkXbpPF4pQRBrlvUA8MFI7yl4NI8iukr3iKxWlpr+V4NaNjVDvUcou8EgxG6R3Jx
CJvO972q4iJbFXtScocODESumy+QGy7wSdnWO1Ndqw1DXh2x6Wwhh3Fsbvu/QLvx
knjlRAV31uPVAk+zYC4FumVeE6ClW2Tj6l4BBHvKpohZFMex4FJ2Sks5lGIRBzBF
BNlJm29A2qC58WWPd8d80pXXRlRy5EshBH4u6c6+chGNCtmTRoa3NI08LuCc/5He
z4ffeoTljKWYyggfxAWMevIkC8yL5dVc5OvEZhngSIegH0RjQcbL74SqzkDF4MT8
deeywucNN+LqoNKGJJ/Vf/dBle85Yg92yr5l8HpwIsMYgv1FkLaa8vUwdM+G52hu
l94aPx5L4UdSqxbSlO4WUJ4KDTOKOwUGQgFEhndq0G6HhJCjeYeO+JAD7Q4So92f
jmxy7BS8e+WAYYrOqb2UDBW+JY2KZPtthl1uPuxpbAk5f8fNG/l5rP9AZn0ZRKpX
RTSovRjr3HY94M21p7RU/dccK2eo7P9j/o/rhF2FXHq8ni+5+5JOwK/rFMs6KOJO
wHFaEtc/0R6FIFeE/gwUVqD2Ug6E+5Srq703ZgBfUjLeL5AZwzUVcuZvPxyihCN1
06nIsRPpxfHv53MlhTpe5Dzg4ViGy8XJx4RxAw+XC+WAEd69IEi9IwzCTXKin/+E
nvGLB8Lg1boigELDz8W2JhtyKbalSnFAPsEEL59I5VIJHXRSLBqqe86SASHGf+Mw
NwYgEikMNlrmK4Zimd5xy3B7LYqgA6CK0dJZb2dFYPuwtxTlamNMhU3QmYuzAbvD
Xlka1xeUxbmnV/zc0tsM+0LmuaFbmgCxiLk5s1cr0x/Ev9/69EkaVmLQuOAlKrHN
YleBZ403bA0zDa88qtHTVTwzOjmLFCBT75YKWvNy4X9URCQ3In4rjQtepOBFs9f9
rNgR65431oxsXtDuEasoSH/yZ61MXYa1BEAkmwfPxGsGp65koGFENHMA+baHIFpA
l2qfae1ww80TF+/O7UFIBIWlFCvwp8b0JrGvfpbPPH1ApPGTqbe8BYuzwa20ZzSc
dfUlc/LmxOoDjg0IgyxEPz/x/gJyAmfuse1lzFi90eJdTu+D3WuX6TBzSXRcenrG
LOPAXLOrPw4Nf70Cdlo6vLQH8s43rLlFInUKGzaHRi5oFjuNkC+HitOf6finzIr5
NfJxbGUm72gGGQhHpU9zgRhXvV5Vy7CiKxFHyxrsb3/FICj4Jtxh7Xvt/iLp4SxV
eLKn8H7mq4qKJCG++FuRDRnL+0IikeedesEP4PGRK/lSCUE+5hfgEEh4AJ5rt+Sh
sLzSyWHRxtifGrzpBXZ95Lhfq/BFZF1IVSMcN2/nC0l5At5WGdqTwKPEocLO7yh9
qctrSEwa2gUHwO0I3ITmldSZzJY0pxTYijYNKaPTDpARSvPlITMwhfcps0PPJRRj
`protect END_PROTECTED
