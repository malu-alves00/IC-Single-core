`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+ASKralzHAegGjycJ0yC96fX2ufCxSDcAU+PTCeKzXWPqp+5yEgKumKck+yDA9Ti
STxUQVdCaYRZyUC9Z05mapnYK3/N3xdG2GQCAHhiv9JGDFW/spNaoyAQ9qn/pu2j
DDmawfH4X+NKNJK5OXStvlTEEqGKel3OE7lghv6WpquI4oGyXF2224Hn9rVs9zbD
3nQXx8brYRLIx5Kh5xklI5R09uwT52LH5ceE7bxnO0wv/X4M+KhXDvHv0U7vy8Ok
g9CsKTZC/ePQiJu0UnMkLLXqGMEaO1HTlod7hVRrOIIE75rwO0bBZDiwb7lvm43w
hIHIb1cDdHTDwqVNfOWTUlnBSPUDnAd4l/uiT2gF71Eh10uF9Zwct0ymIz8MzrnF
eEKeQESRhXOfUWJJSviuN+0cHKvEOA4V2IYW/ZIpMYDB7yocgSX/FHjP1+LW0Q6T
bMZgLERN19zHGG5zTfgrLpaRJ24hDxltUGJofNhVWTe4F8+S2LsOgGv2NjuRKueg
GJXYe9US3UBGsw4vo99yTqXUB29I/O27eRW3d2xnTAMlMeKT0WOfAmJ0Qf6GcZg+
Ebia/PG4dYWWZ+yY6c4oJv9Ghd8lqc9lMHFCvO7IuK1xbW7QDKB7cMTxALPtsuVM
VoVgeQvYj8vAw5ZYTejvua6elH8I0Ll0+rZE7p/xE6ocUEfCUL/8nkkNQpr7L0qk
z81+Y+Us2cUc0xEwcE4yPLFzDNW0fzpJYZqTIieO3j/M6+hW4gOzbbOEJ/jvmsfA
zAWNfdoZkhI5oh1BWwE8m0LuYvlELdbzXDVdhhEr2Nc/+c830+eqOm+iYn6/BJSb
6oTkxRrY0jMt8WTtpeqnXA==
`protect END_PROTECTED
