`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6qUd7Y1BXhRm6dFy2vdPRdxhlCeuNP+RGRtWswWD+TDisgBovhgbgrpuNOpYdkQi
p94gmgY2QDUfrSWvSdw6rQkWQbg+ColghyFiDl4BsTMb30Zw0xzn9hZ9M4EP5jNe
dcnwvrlTJlIJghgyq6lGLSYrFELA4RpN7XqZssvy794Sx1g++fLzRYPu3TFGr7A3
0ed65+T1FpxZeHrebEMZy7xXik+pIhkAT6PG0Q38irPGmDCv1Am/NEQA4ixrW2jS
h5ZyFV7iV5/uMfAqcKv6KAIt8lhWmS3TSvA0b56GsYaLR6Ydi8xoXM1tNb/5RTQ5
EXKZ2JxDyO1Fx7QKahdkLarcXoHxMHOgNo5gJkCi7uIXmz3hOEsB+z/ibPd47m+D
aO0z6Hq+2IXMuurs8HLbRZfA7Of5/59/G4y++1T66LY/fdxYezCbkdFYIkpUbLmU
S6NC8tZrXVZ8ASaFTPYhO14pCJMJ1gzhHLvY41QMqH61H2ilWLsWhFlUTLFOMMoR
uk0rMVWgD6xtcy+c4oMc6E8+hWNjIIEa9PuusqtbNbQa13CZLgSDZbzDIk1YUHyz
9i/tw2ml2Lz49+JQE9L3Vy3dzFJSTCRwVJeKeIRqspYWalDdAlWmMT+DATNZ4j4H
BAeBsW4kH9AxHmBrfThvxahShlCKYcgmm5Og2nxFr3Y1WSiCVoQdunHUnKCf6pzA
ByrQ2Dn950t1ZYfQehX/oaf9wCAMdwI1TP3Ukhet4EpWbDMsAwIZ9mvRkDW1NPgA
JfOa9oUfoFqzPJyY8aCqPVCDy13PAkpsQrGCgCGnvM8TEcmttHFDMgfKrzXr+u/k
e7ANqDl6fr1JctyGXhgM6yEE/hwPiVvqX2l30mhMxasdIb4f6ATxBpqEBU7SCEfP
ur+6FmG0mi4mpnfBt8AjGy6pP1R/2vO+l/B+bBM6rbwpwPkzHjUaU3THLLYnke95
bG3DPXKzUTMVS2AxgdQNOz5QLsCnKHUJZdA6M8BnEZRSNh7aG3aBmrrwIVAUKFCU
b9fE7FXQM7uG0LObNsji8Nd3wbGZt0bJ5PJE2/8e4nVWLJM4go1bprL1tH574A4j
dyIm9x4dZ4XC+y3rfIhF3e9+prNUGgPCFualj0juwesnLo9KlReOEUOPofgkSbto
AiOGSakxpdC8/3mWjcXHym5hrgLmfvZi9PxxAIfCkrbQRSt4jjIGObI6CoN6w1mZ
YNw8PXV6tuTq9ig6huejWoXI0Ua4Gvp/SVg/HhwaaQ49d+L0DqyqrLdyx588YcM/
0ioZ9oowJ4Gl9a2Mw/utUxLpaFbC+G0J072aNzEV8LVHQ+Ypkx9sMYZaW9EC8QuS
R6s09Ax8HeaUyBVo5j3oeQA4u0nDR42LMMEyz2OQ1NzAz6SYISUpjByP2eG5Dx2/
BbcNHbZd6defnwZupFQJ6iUpF9WGXIpbDGMdXARDIddD4pR2020JJ1U4Cq/xWrRo
dMOCHOgjk7nTkmGQJUZO5CAqIColaI8nNPoFUWGQlC18iELPkSTJ+sYhis0m/4It
oAlrfJuZCdcE0GR3at91SxurkCOAo6o0meV0s6QTNgFN8LPWZGkXaChxJ3jghTof
MNIxQT7x9JkWTido7vXzZQDOopqEICns6AcjvqDcRABCx16EYkNFapUpXl4M2COP
XXV9A+949TIROa0/9yKXYQp7ixVvdPOnpZTY+x/eU0VAett9dx4Bvb2WnZuIeEDO
/koCtF1/13sWGtSSs59or6sHcSIbJFt0uxldqzivmNa6N3HSA2xd2gN8uDAQZOYW
DvorVBRPNTVoglCTOv0L6VhRFwD4Ye2ZhgCh0JkM4UlIC4XerXO9vJT69e3tZZPi
WNVVs7ypw3zrVe9OnTBwnkJ9jeFFBhbxTDLpZBYoAVLscqeYPpaOISYW6RRhf43y
mlQ+13n9VQkEMdzxMJdJJzNwduLnJLw3jt+iduXMysFWhsubmmwxueQZ1mpUPH4j
fBfxZbzpG5Pw1DukyogZmc7YOVUrT+IcXdm2E4dGzlFV5JEXp66MHYfbNbR16o4i
vbZ9W8evygqCSGaM4sh/G3OfJPG2aA1sXoDSCTmBa52r6FYpH7tz/fjnC0i16q4R
/P8g/eSZlLLXqJ14XPq9L/29TfKYUfyEypxzPCmJR5VYqPLJt5GjoF2m61tK0FKQ
5aPa3neT4kT86pf3YnBLNt4thLLsGh3lyxjW5rwR9Y8fBzM6Igj8yduoV5gO1ADA
RaO1pDBQvmNqAaRJWrQb7/zPUWzsEbY9wt9+O8zYJ18RVnY+FeXEWCzBhriC6EkD
2scsJZ2KB0C9FGureTBFsho27dvkRlHJy8xs/4WXkMQDyRcOOHUdi2LGQZm68KRg
ZMw0flD73CsMV4hhzMySnKI9R5N0KCCWfrc/c5qUl7skj54f3fg+o+oG1UziARzF
fNRZyzVKUXU2uuUX0ieCX9EVoZ0CdXQeLTqrs1ztPNEfH7Kkr0HB+lIHQidvMLM1
qG8+ntmXbuxtZYs2TpUsCHDrgLJUO4JYFzgUs4snePkrQpyyc+WynLq8hb5kvlWv
+ZlymTbcmpbr69wmFX8s9AA7Y6T6KvKzaso3f2gScGPdiOAMlv/5VhCEZsT2kEmA
F3G/A8ZCTSiXSjkVqFyl1i9PwxNMOnKX3DdwMWRgfPOFjEtiy68nVeLddeJEsuHZ
TCP1wu073u0Y+Fh9Hr+7fzSIwng0JMBign+rzVJx//kFXUDRtUC35DvPAubNB/7p
8aUwpSbAiRcD3iD2AnpyWjadSplFNZza+jyic/62JAwMsQAhO9xbbA6lACevc5jY
Xk3jiPOcmiSdQBUwfZgPxuty7o/s9haYXlkmTrycDXc7RRPJBAv8S/4CrCVtDZ5e
zCID4CttULiIGMngJJbGwGeTP8HSxX2R6f2rexTRA39iZRMoOQ9poc+S6Tazr7iV
4LKacNZLQfebzkoCQbCrFV5T+/tgR5oWXywfyivRM7p1U7SFIrUqlX05jgq2ZjuM
gHror/gyUphPjfD5KvoEisE/pRnTRewGua6yxzB7kmAQRHg9wr7CCNpgZYbTdrPZ
VPSLU9HfogUwFcmUAf0MP4KKJaej04Mk0RWW/gbEzch16YND0MjZXo53On/KDPou
YgRQNvSKxKig2mUOAoYERU0iJ77K++q6QR2iQ2mjMlegJeLYDsQ/rEHWm6G3BIIL
qldJqwprz6DewlhTWX3nRbtu1VOcBUDP0n02NLHWZ4f0vo2JjqejkN0Z7QlwaO3W
fig1M/p0Yaivz7FlS7tel0hF/tMDOfnJBsuDxKT9MjA9MCtOYmV887TxeRz/3fAj
vK2lP0Rl+OnU4gp8no8kAorrIGoF4mKbvJ5vln8nP65T8H9FycqZiYT4ZUcG22XZ
n+pkM8nIGtT0LhL1B2DVUCWN3QVlLzBBRYR7aDZ8PdN8XnBCYLdBPyZmja9MCnAa
mjliOPaOydlHlcpciKcoYqADiCqyJVd/wk1S02sclxK07uRXo5lPlYXXCHI5sdLy
UKRSYx9GJLKeFTcMfkOb8xeVEzRz4PCcM4EUn0DmvDCRHN5UhAasn4dvvy4znrRi
rL7qUbUEBD5xyJgBtljSvPadHbv8zZLAG9z8HIa/3zfzGbfyA+r81TwKshnld2sb
IJtBkj3l7ACzSYgAqj17JZD6iJfuYMCpJUc92UagMNLRaRLR6Um9OfACgkc+dwls
/Kvn9ij2f5bBKbZb7AhJqVIbmNmnAKbDTGORDK02O8nvJ1xIHtKJRSSCstr1AVHb
EMwDRFU8gt7askKPMhnAb6zAPw8gUl+7ZmLNlvO43LaTMKvaydCC3s3l7z3oHaej
XrQZ0HOth6483mUK7FnASdQiLaSa2L128GKE6Viz1B+wsV2Rusrcnz/HMobhbict
wlwAFw31AtBm3rdaQoi0Ja2YUBBlgn+l7/v8MjDmzW+xqoOY/zhzDAuSvlRJM09T
gSNZu6Bbnih7HWn63aOHoKd4soK3b+/uDLGm7u5oegHymdhz8zo2/2c/1j7HMiG4
8GvKbHjyEioulTr0L8DS9ndat70cznpljIwabZZUrpMmgyzBxVjoHq4X8lL1iW3d
IxDLSlCvva9dYGYKf/qFh27FDCXa97LT7Ecah+jd0cROOhBHpeKFfOYjyDz5Drhd
xY38rF8cHSkmAdSEPb9yRjV/AZTtqH8ZDmD834GwVN0eokFXlfJplAQHXBfK2NNG
BrIb9qwxaO+TKMralAO0ZbeOO6Yn2yHz6YXcHOdBreFL570Z/umgCuW9j/DzOEjc
C7HwV+kxV58SvWCTF0V5isRklRLUvWDmwKHR1APpjrnAvzIWSjyZWGjGMQFbVfQl
PmPkjUn2tYVMjgBZPxismJyRIhRfaClO6q9KapaO1+0Txrdj7g3mOQspl3nmySyd
Y3T/tWRUsDQ2WbPXzCymROkrvp6XmS+HKMF9Umh9LNeGXgECqqYXJs24WOJJrejs
1zakEQnyTHQtQvY0orrtevlprpjJChXDJVl4f2fHcavaFTZsdZYXBqMKK8GYiJsh
LVR2Yv0uLO853zmJF0z1PoflYgwKFGNxP1Yhc8UBfYKDUvew1Cip6jn08NqIf+m+
JAxq9ELLHF9mA+DYjbNluhQG49TstX6iRkJkDM1ktEsxZoncxG9alXGNCPf+aGoy
NjeWl+Vf26KTBUThuJ40KvyPNHSSms7YqNAxZ0I9U1DesEZ9vq29MhBurcSVm/HF
inTwurGACvuYx2sDXkSIgFHzpU+aLiRi2B0P1LzoMOnyiMYP4nVxHhl0ecrGYYAP
2GSQ+6iTHQTNoqfpln6aho/zJ/f2/Cd7n2UPEfeipddlZKyOS/P1jNdFnjh66rg/
znof4uMGo0vCsLGCNCDT0/wkaj0MVS4fPUcqoRImwPo5gGlCNwpcqsn7zjcEo9Aj
lGM0va/ObFHIVfTyqAsG6E/uTkNwTnuGF/8uVmnSSB5JrC7fbhWfyBjbebAW9Zdh
DMf+m8SPL7Ab7VbkwJ5w2m2CKQEBjmHSS+ul2NZNWrQ/hqVYEyKRwFEe+Qc5GOd4
sMV5JCeNu11FLTRy1ePKzIy64uvMxHNuT1W7oSUx/gVal0Z1CJi23+2YWdUJOHaH
cMuG1eptcx3B9dM2jYDTwsASJsUpUiO2EfLWZDNUEOOOZxu8RgpPz1wgAe91SicT
Gjmnro979VFegSIRWrIK+k1QmgDWM3IXdHC7h719AIs3y205EO+bNsZvzzRiCcpo
3ru6E0B7jl//h6V2cFxbRWrVzPg9VK4WMsVRUgnv5VeaQp8Hpd88rOxAXwnS/m2/
Vu6CAsy3mEY8mU4hCvDlCD32ct0GhTrMO2r6iPnofsaQfeVGna4qzTHfDbGiZbyL
IZ8MWBrE3pPt1dffwMWWChGovxytmQaHPeDnWj39DN7hbi6Uqy8THjBEndBmP528
LJu9IYknFM8JSeHqZM4T16rq2+vDNQtT5Wlo8J0DH5G9nQOqJDdSL10mjfir3uV2
B3npsvNM3GjhTzTn2TSL1Ky2PGB19cN+lF+riv50tlktb1Ns7bFNgaRgXe87L28E
tiCA3bVc9WQVHoY9TwGkEUV5/KcGYn2Vbbk4BMTVqRvaMAPL2RvUSaBmx1zjl+nF
Wp7bzAE/pgc3g1kPoJCPGc9W9wbUGhvnYN2hXF2pNmYZpUXpjGK2bCYMGiD/6Pt+
GfjnATljIcTGthAnS5tup81/bgkSlb++PI9Ada4ztDQ8zaZC6l0wrCcDV7b7n6pc
besU3u6wK5GH5tIj5uOyLWVdAzXhgfCuCapGWvqf+3A3HBD9qYLMWvn24GeGHZ6U
gbGG2xKI8f6b9gagG/5TkMpzfKMCE1yU+Fj3rmlqPqrAi7ECjoFsp9lYV/WJBUpD
v0u5fNFuo4XaaTnQNBAQlTQFGgdrwVGzfbvTHU2AvTBWWnDyuHezxqneIAMcQfFk
zdP8z6uHFJY670EEw6TW90yAMqZmxoZdo/vXXU1tlSM=
`protect END_PROTECTED
