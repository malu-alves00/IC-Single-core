`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sMldT9o6R+2RjElfwQEFLHLhdJeyVsEJcI0uAATlbzHRWs8/RryFfKo6VTXRwZV/
/pu1r2q1xB6ftAXr07Curgdi2kr2/Wm2sc2X/oH/0M4HsP+XhXv4/lLF6Xiq7Prx
qn90m/PP+urIKJZKPEOQg4jHH7h99Mk3WIZTUXMN/GxCnt8jjInDBdYH1TFbxg5E
Ya2HQOvh3kAPnmn4/7Zh1qZGE/idyP9SsqDOw//xVGGFdy53ugeD5X94hIcl2SxC
jN8d5OKPFrhlJlfbr0ya1nD82zBs7kNlF3WbR02Gbt/rX1iHo9gxPkCjhk8ARaoK
BPeWrcA4Y/JTN915joXXpWUjQSiOL94QA6TD/h8nsEusy2SerDxCrnEfcHEc+p5K
BcSo/OuynT8ib/HURDH+lWlSaaMNcfZuA5nrV8jJkgjNR+8HKvvCV+c6riqdQmkn
eo0FAPgr3ZJutxegWnKWRlD3PwsyTo6QlrvESaWuKSql8IfxpEAF9EIBvUZWRPQ5
gzEgiUCizCqBpU5+kY7bQSrJXbjg0NisM1BTfZaDO/hYHSEIFenN93Nfxp0wo0S9
PP1s20UtsHk1UNeovt9q6yJChTQ9E3CvJFQBOf3SONyzUQNyO+9tEGDxesJ3SMB8
yFEHQzVUj4Kyr+30TEjGfjwxQvNbhgSAj3YkE9CQclKyRi4BUBkYZnZbmIQaSftx
E8DwhxmDFeeqvUc9kqcGsTqSAbjywKIKQU5AroNFWv+Zv62UtJRMED2+t080+Qey
gQQbl9OVIP2s7VwOu05maFUTrTECkrUaI49v6XqNd9lDvZfC6lCInL0HdX1968y1
BTfg/vDLN/16xL4QhXmJ2K0Ykvxy4CoU9KVcakU9q+1sdaSYOsOuMjtpUcUzWYIO
c+F1ZrCvocaua/4WqLfacoKip4JVhwrXhP6mlNBPijg3Lg7Lcw8EDdelvPcPJr5L
E/AzGZ0PEFO07ueogYtbulYHIcepCjMhaicMjNKTdso2vV6VX1tKhASjE245Z2KL
TZcajfHlTW25ct+8E2rUCxqyywTN4519PchGz3OIRaoeKGzKZlgEyiZFNi8vUH3w
0GcLKEO0d5i4WJJqxBvDc34GdSipSatC3GYdxvckQjPc8defsIiCTp1EbVgv+75G
ZhUUZeQ8M/ZI1gNd1/2cE9Tq2L0u3SJOz/XlgOie94w4GPbH6El4d7N1RWEL0aSc
pWKGqEgr+Ke6BIxyl/7G6A==
`protect END_PROTECTED
