`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
y4B/HCeMWzu6VbiYpU/37LVua2Zd8kWcpcFbQEMMp3bBDLcFXv+bh9C8gd5GmvZ9
aruwLqnL80My2k0Q0anvYu30HZrziIny7pHEbWMJEfZqRa3uJeQuWecI2BClzZvE
gLGlY1mALdSXXNAcVlkHFspCtupFpI0J8Fx003+1jNIyHQQkiCfmIPkQAVUaffMY
O0ywbEeXkswrJ61Wdh7gyRkfuDCzRC/IlLpQ6BVOIcURjCI70XLR+E45eCLkuXBG
pEbuRg/EFbHnLNV6cpCzjtWYHNhABPcIjQqaEZXCmcirk+bOEhSOr4IHFLdTqGsX
dfIR3W8BCrlvzVSU/cNV5CA34CVtUSZKYHrPSJSNw9zTp6fQv2O3fVBsK2NfNTk5
Fo5b9xwL+rNqy4PyGjHbC60qF7hwh//WcVlDUcUhJPqlMRxSlaIVmC1bFKfF+j3/
dV+0bqtP3ZRqT7KCED1kFQ==
`protect END_PROTECTED
