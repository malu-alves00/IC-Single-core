`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SD14QVlThclxCRI1hsYNZhHpmq0LgUfSCDQ0fS0nYMOiGD3qZKFs2UBUShXWhMiN
oqspO0nqYBEqXH5lu/QKExAN7morr76n2fpoFZPHY0V7W8GpVy7cKxgToD5yTaqM
4pqpHaDMGbzpW5Vg9QQck3fTy/g9yTg4orEnLZ8YZYuysztZfPQzDhHy4FUAHT7V
sgeGXFNQGUocyyKop+F2HfWLjdBGtSZaztFQv96pltjLYQg4uJjivwny3xuArVpJ
LGT559zOpCxD9Rfqblc0tYezbqklTHUpC7tG0rQABXBY6cAEUq3hAn8SLRvWirUq
+FTblSTlx9i+CI8x58CVcGqlq2dJ9IkRI3tgLrRxGfdEz7J4IZHJsd7C+hyMCDzO
nwMcOYS32Ii/C3TXyjywQ1eC8mOM8zUZRvvGUcFIBGTLKtc53iDYUyd+HeMbY4cm
KOPwP2xXM4Aswt/X1FCIHytqJE7G3jdom8CLzDqitfXd92wIueSbWKEMjdBAMl1l
Drt2ZI8NooIjuR0OzARh9m5QR8t4t/MNenIJGgHasdgHL7ldFppawTGhIbADoQEw
JdHXnYljXsXmjc/wZkCGU2Eoxaic+ViIXnbYDDSFNnH2yvO+Ct+4jf9oNlo+Wv9q
Q8ArADV2VrXp8kwnOblCXlI3X714s15P4bRVek/W3ykBQf4LUnP+KFHQfGF8b+Tz
AuRTps5y/JDYanmR0RqJdl/wWoWD4x07VktLDzBr3lujXxbwDGid33U1WwSU1VHr
idQKngV/Ezvhi6utuSc6LXFZpXVsxgrmtbRQftDCPDZyNaJ9ZVS+VHApDsR14z7m
z2SxO+8CIUPv9gGgTW2NXo4SUNrJWum10peOBMbIwpk+IoHjmadOTI1nq7ZyKklD
MqzpOjU4gdrnUhZ7WaTgmJ1YW6HEunTeZKvrDk+QfrTQQt+CetXvnrmLkS5quKNF
L4DLWSAH6BkMH1YB0PVMGs7mwcEZVze4rEYkVfrwb/bZ8UwjnsGUtFk6xtv/0Pka
0UvkG2fePi2GrMhItYkZeOkvTCbSfQOHVokW8VKLW0pH49Q6d7HlkADefa8X5kfj
CluqzKcW5Kp1X9UfyLiSRKF2M/CQCxiEpAHmq+it3Nz0m59fMz6Vv9+R0w2d3M+3
8xdAyyXBYJ0yljbiE3oZ+BL6TOe9OaSb25QXgjv4YxovC8U2ujy8cOsDbPPYAvxs
G2f84mYY/pVViVX+ejPBBnWA1LLI63iPDqVx6g4rmaXH204ccmxrcM6o+dBO1IWz
IetWPXDvdTJ4bWC1gVpzLYiV1exJ/M/1JJkis3uyjzMf4zK4ujFUaiPEzgRmGz18
C9jndwIl2HMI5nsbWgHChcvGlnBzsSpWlmEYlqZaZh8Meb0bf0PWW15cG8Da/xWd
nrk5pz/TM6UUOTqq+qj3Mfc/NwKyPxhRJ2gUUMbUPiZ2yHrl+xMTO6v8vwOL4K+P
RL0k//xtnnj0boEOmtEWcBJi5E1OiZCESPEAItlfa5AQEmQZZNEfkGEjEtQJuu8e
p05MrQ8n6JB+F5Ss7k1tspwtwurB9OodSSpKlfVO6/dQm3MPIcgKDaVx2DA5OkBu
CyjF2vP3CivNQlRY0OvBAyUbTCz5zmcCUet11/kyrBNrKXF34e14xxxDnnBYdTCH
g4epCvbzJs5lWsJ1K8RtfXvqExm4plxIdFHm8qsyyPtQpdh3vrFFjg7wErtK3Q2j
LnJuR4D1vrGfpyU2b1E7Cmqtwd9IXDeRt/shj34h62Av52eA/CX3wq9+8gaNGylf
I+9IAfC8DUTu6WQP1xD+ghQbVwxexf5Ak3LqmbX+t4Ad1fCs/DZo/J9U025dhIup
8+negsS3uM0LmUMzfCi3w5oYKEDelzo/4MNU61jaXNa9mtl0zAPEVidIOh6oRHws
kKwOahAS/wp3VWmd/z4j9brN/qeocxNPlgFAR7Nou5s3d4CWIodMbW8MajV0ZA5r
/r/OI7172NcBGlWJ9pBOH8mn3wxSbY7OLHhEHRpwoRvKcv05PQWKv6O/1Ii8iK/Y
YC87n0S4oJdcpJGjqZk6zJEeSscwkVFUhsNjKf9oxQCGzOLRmWjgzfasLahH/y0z
UjWPmh+Fs6Xi6BqVg1eR0ujXCRmi6wJhnqiih4dJmdREAww+0lmj2FeK7R3b97qO
EiA0IcEYNMC/FlTi8WjizHsJ5gL504CAaVkzJdsgVPyqxqd7mynPapNVfLNAEu3l
hXUL69jcUrzGOhN6kSTARzecu8GhCzet4eYDTX1gC9KQrapyI8/9tUq+oIxC6zP0
yft87N4sR4axlnQ0z7FAKyYXhRTviB4IRFT8N/PIA4V4qIhofrDhKenaUlpPa1cb
aEkbnyBjhkZEpdQoCshWmErnJyeeBvNnitPBkBxKnTP64kYwk56Rkx5XApKGIDZR
Hor3LrQbI0RQkJlGA3QKFj/pqFicdAE5MefRrqCX8qy8L8SEPwaNVnjCfsWfqhVH
AtU+SR1Mj6aQj+9iVEu+sVF1YpKAN1eplqyglskCv7rvh8Z5+4PyagKm+TzWYOp7
XvTJyh6Z1qwFextjo4BN+IWiZe0yWAdr+oS6WUD/vF/NIsE2SCQCLGk0kISPR+KS
1QFkqxhKz0mhvC/zAGCX/j17+7bRPhSOSbuzYlm+wJICfGW9QwezM7cHKQ5n4OQl
s3m8+1oI+u+j3rf2sG/BcbcaE6prtT6aa662tEjoA3PSx2kd4Buiy26mb2+3PU6p
ageWVOHazKYFsdP/Uzm6HK6uMEEzldQpOcr+KvDlYUFzJf2oFPKBKzx3R0Pg9PZP
pOE3ZwqUt1Yh9dMJ2eoIjCLoCP84vy1+6rhKc/xbxijL4MEv1n5/r+iUy1Y1e3We
Ewz9SdO7NsRsbqpFmOyyxK6TbX42IW94QQD9HEE5+MZN8H95Ufw3A77Rb5EvOfRV
YrjV5T3m7xYpVQhuiUgkHhZTubPTRhJSZG/E6MSoU3FcmnlAuaPBTnyTcNeJS7YU
kVRDLrt812h9vVa+cQjfilLKaTIx32OLQQdDs+17aoSu/d4K+sTVEoVpa5CRI2gS
lhFD2dWx7jL6RZrfPZ7SoBTi0dg8kRmrMQlzlq/FOprbR4iqiai0il1Jt/Iv3c9k
nn2mvEj43UVH3Fmw7QW/cLMPvXj0vQU1bzKrtLsi1jmPE6T5gXH/5j6kzw8JJVzq
1sR2fGWm/R/zWPnE2zIeJeMXnx5eXmoDuXhCChD+Dqlha3zktOtKpgwy9tCo3kJz
+ytgsNMU+rtz3iZIuhoVBJBrm8Pg0t8jOt/4K7v/nzLmvY6AfyIWKfyjFW8WQoFp
Bmf0yWz7Bz5ixhjCIM6zymNwm5og2rTDawLGFoRFDpvG9Uvh08TSWTF9bYcQfo/9
xJOc5knQGwy8ZhhAfDMh9iHCxwAigr9x6ffwlQhirM8wyOeQJbqDb8IJwr2WdK3h
3ZtvRB3drFsgzIw6S6bIufAcL2+0gFHNPmzXIvYmgVJ285SaeqozK1icEy0fZRGf
nCmOftdqStfaMCYEGkb3gxvmFDyqovxCn9/s7+5bPAxY8R5BLaihNJKbHvk3URbM
Jx+CyXzKA3JPC8TEAOCDvOaPm9VesAr9h9nk4xDEctWjC8HsQ2vlh6OwfnS8Vqu0
dQN+a6TGe/wiWDfuKyftn5UA+/bL/WuxBeDwL53LksVNIr7NruCOhViXPzAHYn0H
QXS/iFyzkQ2arMZ4Rf3lEEY8jtSq2R2aNFV0m9VCWSLKxf4ynIAxlWLIR1itgTsa
kJM3Qg7dHmwCZCv0+NRcOm8FoNo82hsiQ9vxsDYch/eBIR3QF4JVEnn3EIPBBj+N
dGPOwPNogNYuV2jD8l61w+FcIm4BPRDa+cq32L0m9lcNxyxyVaRVFb1p7pJeG+9y
vq/FoUPc0uRlL2/C+avO21id3ZngjY++Ni6TjxZSDdDFmNGWz49gUYKRyFkKEQJY
L0va+gYSFVKbl27jrexxz2V/r1Wb44+FOHisjShmpjIFpc1+uCMJEX9zWd4Fn5/o
m0G3+lw0/vjT75d50afOOQVIi3IO3i7Em46OeGeCSzwC88cDKqWWUcOjyQD0+GSY
maf/zMHvaxcRjNrW0eev56sNrj0ISqLBFVDBTks7kKmjicn0rLAmJ5cIxAOaLKx6
GFH1pRdq1oJzAEa2iYLs6Xo2zHKi62Z4cxPq2kLSX4ES+oh8fHG5i34+oaFs6PFj
z+84bFwgRHmFtPh12At/H0l7ejCC61u+9JQz576mV/GGVdFQsgUJWa2iGwsUV3ZE
vM23aUJCPML03TbgCadIn0qGteliCY0iGRqiRQSu+yhUz1TmAkWsIYTxGOOF4Y4S
5hOI1OmADvl3V25Lum0sX1RUzy+dYC+KKKW+ailjfbeFW9fYOdS9snGnBmw8PEnB
jcqYZsINey1JPKB8wonjmJwlTKL1V5xxwakyCLbMWWfLXGaHlO8O0sQCQ1EWrQmS
p0/a61U51ntN+Q11xqJyYdiqZzm7Jql67NXpvaP3EhbXJoGQ+dECM4KeDVwKdsKH
eA5TmCvX24UhEkuLws0yPRwIXOxZxbQwn3wFp84SgxXVZR9w9gUTINBCOIP4GN8I
SGYiasd8Aqu4pfhTM+5ovi/R12/4/kQCVRLpxZy+XP9kBFIiNmnsMmmWi0AnzDdD
eewd4DrF32GMOpCCjpGBGMBVO6Qpx9+GAVaRrsVNTo+UNPTnlqDWHpO1CRnUnUo1
G4QRky9bLbYuOOJs1AtCgBXBDsWZrzRsV44oHNnZgY3EKpBumKRJXt0z/LIREG8a
UAvSR0V97slO44dCz8hCPbkIZu7SCLC4WY0tfDnUoI3dU+i0QWd+g3nJgt4+yxw7
11y56dQ30xqXdPHZabnsCV/7FhEAf0DGlCU6JOMoBATR1xEjoPEotYXj7YXBFPeu
WDphFfk2KBQH1gfddd14mcoblRBjXNSi/OlK70vuCgTZNhHhG6nR+s/JiGrdQeAp
HTfxc3YmuSm7VouTQVKTeJA+PojbiZw3bHa2NZyP/tDClTjQNlKLigCslc36bpSS
TZr1p8Oxlg96uXYRgbfC2BYmErwPYANgfaU5QeZZ9iT0Ki3nYq6C29JkGfglv7cH
zcq8lnUKzh4ZT/eJCXs8nijISK1Fi63wy0Iq17dGvYbJ0XaSLepG7c0pGGZPMHzQ
LTXgw0aP/cBh/RZ8tPGRc6mMOT0h1vvNr7w99xGkurkfp0/PJr421j+0e/snyt9p
qRnvns64FCyRdJYuW+93ApiO/H5xDLiukXti2kftISoivJQ6DFb3IHGq6yU6lBFt
K6eKFRCey/O7g2pKe4bJdehsl1dqNWmFlh9NU+d49AW5dmO6nZT3yFenBgCg+6Gs
UKp+EmtiiWSh+gT0kIWVLnmJl/W7s+jarcHoR55ch4xeEQWPKB5p/A/SfHx/qZmb
VUyy7sO/Fc++HA1rJBiXWdAZElpxxE5mb2++LZD079jCgbS1PV4oLRDWizc5RZay
y+pnViVm8fiS7/tK0jA1As1gHeVK62r0h9phe6WOwvjGOnTdLTVapk1yqO9K8jjo
8TrAQoAyHFm0AKioWhSIBygpiyWSz8hOUIaiAcRgoJ7P81NYibfXX97b8TO90nV7
CNgxFviLDNmSccsmavl7uWAYBO/0v8SbnJ+1sG8hH8wL81/886Rx7c0QXh2vn2qL
eoz5YIYhw5SyfDCD1QgeNpTjoKPM79KvCJ0R0b9wLLWQpXNaoh+wMq7a2MYuSoO+
lycIC+/CAk1xYMLZPZl3EzR4Bs72eHzutOEvrU6TkuE=
`protect END_PROTECTED
