`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tlQKJRNM3pBKjbLD75D/t4VoGJ1pgqZ6WeSOHTY5KDxkYMGSOilMCwSPGKN8Idx/
RQdK+578ElYCQtl5NGa700/c5ggP5UAXlnRBDaNCgFSyKWA0ZtUr2n+kgzD6kikc
XgwcYPoUC6m8ZBXKtkY09KwZ/4Hoyz+vawohhB8xAUvS0+0WtzVncQ7HBFToG4oL
0t4lXDrRLemoM+NNvwjh/14OFMebGopXdsn4NnUc8NjdYIhtTGxu9EUPtel52iYi
xPfhHU46Tc0WcUrT4/v+pPCgGEmnstmUJOxMypBzB4nozYkP3ip+GixUSOlpGTTF
MgRJF56e09/YyXx33im3pAmhMb40EzGvw3glirSIxrIgN/VyiIH3n8nJ5RI3zrEb
fZ0+5qItDFLBI9c8Yrz/nNhDgg+GQ/qBWPZc7shlITd0pNtnw5/7XkJ0+lpTpeKF
QUOqSG4iKprugEb9Tnf1zNjngHTcNZKKsei4GUI0KrCXDJzoyFkL0P4vrXfvrSLy
2RVgxnnD0mPy87f/U4zLjr8a2GifXPUXfWwp8JjcH8bPveqsnugipLDQaI8RU/wp
JuWAqzAi+f7h5f6+MX/B2bhFoufZU7ooq84riUl+pP6d8abIsZNJFg4OWri7LbDn
KCdSHYJM2qlHAPM/NU89zsT5ulrOtG8HyT4E9j1ypG6lUuYirkaMuuI03TxeJG0S
LvyupSd2t7w9BnCR/Uwm4cGujKxdxfz+uYTcXa/C4diH3kF9vmKQ1I3FQwValr5t
c1sMFqQSLpGHSSWcnOPCSKCfNp5QAv2uYJluLEeIvC+q08X8KXklWu1x68kLVTLg
gO1YkBCJZT7jwXrXHy2FSKHcAo9nZcqDwceeiPTEJARH8asUpuvm4VZwh+m1bZGn
FQp4MhDUmYKo2XnTEj1ukAHnIgebidqZtx3KAlyl+gIiF5ZuRYBaUR/DL3hplmlj
zIVTTd7eL6/SdwGf97RG+2GkJ2T+dk/ZygwM05k/mg2cap51S1iWyqATwZQRVZQl
Hr11zynER9dnqEN5G5w7VHiAy5uNcy4d29nmWr/TfPCZRWvewPm99/JGHmKW0M4w
M0laAzUPe9XOBIU9qk2m/0aFJA2y3sEcTVBe9ehWvnbeDCz3cw3ZenED0jRUFLW/
sqU8vtnHXtASMQrXmv1Wj8etCjYHVLGRZoXuISKCdreLu9fHmQK6O28mb5jBaCYm
fbNC4K0BaX6zibpnHLJOlyvrKzK2JKLj5q6+4kOFzGNazOXxbUzH/v5bA/dI4/c5
UHM9HG6Miny3ujGqQWecFH2sMNMQ0/PxY8GLSuAnsTsD2N6YA5ZbKAqfd1lExkSo
NgrA26YPvpOjTf2ZcYXUfTOPV6GkR6mmo3KBGc+TrXwFCdJQ0jeJJrTCZDNqAH+A
cgmB2Y0JKmYaUHERYGZ2vZrlu9OX1zcmn6zScBUxz/BQvgAdrBcIoE/46XSUuIk2
FzJZOy3saX3BK8cY3/y75AU5q8V14Eivo5x7iYzA9AJezkswKL6xmxsIn5/9f10Y
3dMaJ1EIESZNoJjEgaLVGRmk+MngH4FFX4V9IP52BK47EPLEp8Oro0Q8khC211Yz
BAoipMeehNBytURX7ZgAz0kdSTopvCJFp3xYB37SvaMWKIp8VyKcht3s7oEuyRI3
nTyb54UfBL1lGGZCcasinJNVpyw/Y73AEot8p5JPAaboihc1UVok8TLm7Z64KKtC
QMGsTTAXOCH2kLXC0t/vs3Zi4bNesVKGg6aCtzBwwiCVzHNP/XpEgPg4dJM03ED6
OlIMf1qLiVJYV6at+92rueXvCyYjg0IXJvPNNDDEctTVdYXHaL2hWVNceNkGxprN
0TdwaSDOEUy+vKtfPONTHmvXnvN/vB/9gGWp78AJ4S8FQRwlODF2q2ZoLT1hvLPq
NXre2imByvIyOmuYXeWqiAy1rJh9aQAkRcDZyvJ50Vx5NYNGApqrta7hbm+/VjQI
9Fh0NsWppf+HS+81gjkCdsOLJgBkslBNpDdZzvrJfxP3HnrVb8D9xBW3qTJIfDxH
8hbmpaRDmwVYFd62iJgup7Hgodn96pxBFu9oc145PzfAM8hEqrnGcZ0LS7Ny4w3C
b6rIAovas/B5O+6bodMFBB+8BjeV+3j7WEpC6c6B+3358SOoAluRj70xu3z8eZby
xaka1UtOL+PcXQQJA6kxoVtRZszMoj/ZvbBlnOSiAPzlss8UrjZWqfsTNfi+iUAC
G55ozsnrGlE5mpYQPTH3ouD8j9tF1w9EM39IZTvnK+VdipzvHpjUf4jPfvYa3oK/
Kg4sZpEQRja7nus6I7PwRQEQ0RR98+gmR8zlToV3yYpZU6iiQY2FawXsZ2X0nTGz
nZyCnoFo7YuNeFE7Jx86EYp6JAkQxRsHa4pMEs21uvS2fmBI90mDMjC0CLb+k3od
uwaz4xeEPHExD2irzgI2olnSUyyjpWLRSC9GkZEWvuBuQki2t9ztBBZMYDVPiKxn
Ev7hn41WKjsZqIODIALWxNXPcmV7zjvVY5h7ltji9RPFecOUZImbzHh5mpOK+fnU
CVyOyxg2/hjHvaDXq67lx3y13693VoHsOy66JIrKvJq/fGfJodShzdaLlWJ4civL
5e4YEkB1ymo5kDoR13PfOo+pKOshopgcYvT3YUnUvim4cm0TETpF/Q0+PBz6m/oE
tjFDkGgwX3ukzmOzVXr3jOH476tNdckp35Znl/ze1IfMGMLvTA/0J3XyINPH1GlI
z0Wh4ZSgaVbmUlg/uwEmqKld8KjwbVN6wEzQ3RQO23Ps2QQeY17PBZIV5ETOu29C
udfwuv1b/BBuVomKcdHZy9S3+Vk8GPJo3uZ5/gvy0EdJ6PPf7axfoeVWhoYFNtzO
EjcUa4HlgMGk7/1kzdP6JjPsuARphqWfy7eDuVU91Ke4GbVGRK1APLMswQ6hfk5m
VVTzkwkNCXC/lYISYQO+ePQojFsrxJc0bidGJG1lGl0G7ExSWYNVLEbXjl5eR/fz
8F5l9/EXu0GsInennPOQY6KdnkhFBstypB0K+mUHLpKqV8PJtTEeUaDAgDsfGSgE
q3Wzm4QhCbEXYzHhQ04dw6CyUgY/IQ3f69akk2x1Xv+MIaglZbo+iAaf1rJtnaYy
i1S6jvche1dYuyWj8kpB9tsMX49jigJT7K5NE85U7seCuvdFvkIAqHWVGK4znzr+
u2kY7yZUi/+OOECDnlC9kMUzseL6tD6Cg1LrJxXrTd2MNsEMEwnpP6U7DrOvswTl
lf0Nb7gtGGO7uNZ4I0tOpebjyXsqsaKd5uCscqZehSPh5OouWaIAsD7D6nmtNyTg
91VjDiOt5cc61CuZLVQpm5nDKJ3ewEGmPu2IhQFkoLesD6q/FaUssNJqPhsMOH0X
yCcPxIlCyWsj0ituwUwdvtfdkoIWsLiScWual0Ca2OUzfmRYyvzAFIIvuFRk54rN
YuchIagJHipNS88H+jt0m1p0gpdre7qzDj66sgdVspz5VY+BvRmnEMejylM6lJBT
Bz5PjrSFZfxIBNUJTdMvrGS+7CsNWB7KH1ST+QrgRfsZ2CsFvzbAue9mJN3GNbO9
ZPp5ZWHQNhdUFHb9eD+/FxFuInNihAOCC7bX92wsJlgN631Jk43DyNTI9RK19Ed0
bWkfR4HtDqsnmxAp4nCoNty2AnF6AkekvmV6T8Cj+kuF6fhYZGWOhlgCwN0aj+k5
ev9i9QuqtR6eCTLyi3tW9xZ8/f/HxrBI9pvk1rufnJrn9717uQFdyk85exu/zw0s
/Zcl7MzZCIUBKw7F5OWUUwELRqqg+gDNg0d25VfLdUqNpzdntAPl1y6R9ktQUYBN
WUqp1nL9bdIKYW9PmXUeIKXPrqLb2hTLPamchjOCADQEX+kFi9lKJjt51vm3/dl3
VCqfi2cfGKhRqBECFdHKsIahYssB21S6UWL1oMuSWEr0R1nFzKok9BbHSYnWGkVt
Vi4VYvDRj8kRhYKg54gH5GlOzpsXyS+kab12aF0/P7Qevq4OYxGLZvWfr4V6jVty
KO0ZNCd2dJ/NTiFJMzAAZ34mzgLz/L6H58uk4SxGgzhB1n/u77SrMPwr4V6QfQuE
x4wOo38Gd2Rbna42C5kebQn0FZ7mn/v8xXxQblFdiPrNk3hYlvIUB5sltVh5heJP
u0cJ32rKEySHwz1KWQepAEigWm4CX9sUTH33p2WWrNlbmYy5jJRQjpgrYCz63zYQ
LKzaRtlT4s9V6gwlxTX/hHKIQx5PIKOmdk1ci+vsZ7wKWb/8Gg5gFGWazgfLg6GA
8NjLxYoTcOVNJqQ1/SMPak+XLr50duqTbvblpqGMIaw+g95Qk+O7wL/fLNsRcE3k
dOL/nmiPxGm+9RWqrbpg7gKpK1o+8B81cRym/sZ/f/ZYTBNn9jbYaYUDk6Y8J/Lc
gwL+iLatp6VuIHLxFWFz+fsoEUDcSo8h1qcaE19Y65SdtXb6bbHiZ5wVM5v1noWu
NihjugF8+aOYS0SQHK+iKx0aZBjIQwR7kQfibSjm8n/SHj/Jbz1oCPr13BnBirer
MlLmUTH22zHOdtJSsOTpCC7wQID6J2Fo5CfiPjilhdTyAPlpB53VDrUX4apQwWqW
dtZRL0Ka0ir/y4PlN+5Ol6Fz6I75xRLCG5T/ToixUUj6i050CTaX1/yJqpQtEij1
jTS1YpZ1apTpf8xyBtE1huH3TpNR0iOm78oSRby97fnYZDMaI9+3q0X7J12rSMls
O2h9q7vD/oXhka+ubJPURkhxryJka4hIbAQCotlgrkdKtxB+FqncTiYY3+IcuHLt
FpRwsYU8IwULLJc6G+752rQK2hyyGZseGugv8+9kI9O3wfV3jCeA51EYhw4iS297
k2fdbGInipbWA6LjijLxf5/m+VpNUz2NjK/2hMJoga9ro+D6IlP4/URh+3LXhFK5
P697CGVvbZrUdVVsathDwiQjHnyG/C7u/aXh/UOPoHyz7m5gZZUT7W8wNZyKPd9h
78PqjqmZSzi+6QswBMD18armEHXBEokcP/XrBpuPzANf91shhh9++rd6GVOY648g
6bkNSYfesPoJpOKMUMDgDHin9F0IPBD1z+JzgU7p3LyhtSStHb9SPZ+kQzQT0WW6
6j6qfpvAtEILKr4mHQPZoYbgPoN6cU4eMEF5w0ff2ujS8/RQ9RlFJJTWBz2aEy09
F7Fv8ETmHLhoyUqUblZqFTr4ynDO+HmfT9d6VPavauyjK55F4ZYvsICsa4wa1kz5
+bVdtA73gpcgF7QTeQoEVm5s7i9fEnMu09tsitH5gSVI2ioSeA6ArKfiHPAOApqx
qttvTnkZLMV0CO0KCgUc3FgDq2XSoVus8oYyC1YYAhpHs1ajnBtVV/5g/tbbIHjO
c/Pu1bPhIZ8fZ0FzMLYXtBmohlKyrWMlTV/sLJKcI4uR9qngBEeawaAcabHeiPJ4
0ZklOCp9Q3t0acjJlvwaESm0o93lB0WlJPvs7EbYy6zKaP7N/LtJ/zf3WnfcRHqP
SzSWAed/74TCRMbdQ5IdeybSd2jd9uWNukSWdPhiyud31R4p3RPY0TFMR+epQwQE
9N8hhO4B3b8+cAL6G/pvtrfOKqyShOtshQhKm/fPvi6JMFpbPrDZu0uO90UoCvxl
2YdXYvFCrNkDHBEZlU+oxysO/Y8pqbP739+xWKYGIjrtkM33kOkwzbmCn0uubIB0
71UfLd/i9BRwIf0xGL+4NKiDS7p9bq2PP7luO486TucEBQtAXKaCWnNjLuytRwsn
Qysk6EjPm2RXvTVK24pHP+XA6iswRIpE4e+6O+4fZXScdd/7XXpJNE5EEMHwAJny
39hCfHi1+KiwYQXqT+oVVNxs5Kkly0EFh02CUCCTtonovVoAH6hI5se3dZB72tfs
icqv/gSnkEmij/bwQF72QPaXrLWXCSf77FZztganAEX0q7VJYrfwqXb2EAViKWXs
kWEt9uGjSoeEndwsqGSaAokW3G+P2s/liFeV8l2Bzt6dBd/di9o6O/S9usnJjzWS
cqjngENwCSk7DDGV018vnqEjrf9qHhfeKRCyPozCgi9cF3KqbIXpTzIiTymIA4+U
EyqOjoQwJtD1ei5NQkK85x2XP9Pp6VKvIn4wLoQPiXeq8s6MjzYPjmYg2Ua1z9No
89HXfpJyEgpql508iDYMH8CKU0hEf+eR3xpXniVS5ItLi799eofWxok5UBvXHMbZ
XDIkVjQNT7mUCOspwVxGUVno3rOqUm5dzQmqWKDEUXQTdqlgUe4gEZlnT3u+W4Xv
9jbH/RfpcTDvlaQo8aKA8TMB12JAsW3SC0c97x0JK15WKT6EPnJYgHpYg3cYPxgh
+jP8sPyA5tzk+U3YIn0j1D+5vZ2mnt37H/AtNPpubj/ycmZ/5p0N0mza57Y5RqUW
gG5+F457u/bnrQtdhNsGtoAUHFfcUXm6TRdab6s8EJ1nUCXf/NZEsP+2hEoXHrlO
NDpo0BNmna7LaVKGoKgs0GAvLZo/Rs/+TBVsl30OrrFc3j1AxPGN3Jth3nmYYjyW
jCXb/mTv0s1Ere8kknIBw90t+UaB/ZXb4ttutLyhbYC62CFpGvbQAMiOn824NSwv
tx70qOJNOigxukflg5EPb/ntvs5nEgp1LTLAsCDYgPsXzEQlXQSIrO8idHpu4KCM
fI08wyCBXhNTMmdS2FdCuhY0h/qllgLl+TpZA/DXLKgu9HTu+ez9s/2UQYAwzDNH
yTrcXJ8CF+eYn/SpEptssZ4zdJaEMef1jjJsmGP5OF6eL15/8Ohs3piagBICaFE2
XEWOlCvD84TJCYZD028eReo/YGpDoj+2MJvBXmdIk+n182/MOoI7AtJIlggLOpS2
ogZbyUgZXZcTDuMRp302I7MBeBKrur3L1oD1NiCL77moYXMQVl77uPQTCXOct76+
OxMHo8F2wtX2p/1LKCSZZolzoDUku/vY0NKgi7XPhEEDramONUNPckDfAKtMfNhY
DWqInimUAU2g4i7EnTpT+GP5fY74smYgdGuHJNoewvwpAcY1XNd3IBqwRMywW3dw
RGksifMHv6uz/swlu8Qtsr1YWxLwrMrhZVAP//LVnzRwCt7NeKbKRFY/oDKNii5O
sCAmqKpwFrx4s7vxX+Kl4CgmxyCK74yWkL3zcdr8otJvu3x77kWW5T7ccEP2a2kv
ZDh1n9u0VxaIhzVhcANq1yjyIqmNXz9JWsYTkpnmHY1v8OHM5xoJONvjO3bolWCl
pqOe38A1FOdngAGdx6EFp6K/ge3yXFvixFXr1fq+0cNg2Z70qwZPeNqKfFfaZctT
7LV8938JevZN+x+6pG54PKPxoP5xI5fRXUMJt2BA862oO2n2TerETLDljizHE6E4
0kBmo+iG3Kj/VI/ajfYr+0A9bWkY5z32LW0/Tu8xohIcf3VbO4rWhxVwjaQSYxBa
a9dt+kvmtPhgrTcrNa3d+hLikJ10Obd32tN+uDTlBa1B4jRiM/bchCuySitgMznr
G/b0yRoMESkoLCuaQAFMCw9zGkuEJNbcZc1Yit/euPgQcqwruScrS+vbB+bcv/UR
thBzn8YWz211DeJ1+P/mHlhImN5UQmT1poEXm53AtIbtmFfoUDmmObLEKlQIxYFT
d2LQv4HSxdKLvxLUAlz2kDHlFo6VfN4AhR8c0hsHNO1srXP/AIZ6jrSdM0T5vAug
hsJ8noS8fTYWY0mBO2+txo/VRnViXKy0udrnlw2eSZsbYLoGurkaVQlnPS4vqkfA
kuYf8OGe8k1MBXmm2MzPfR6Sg/LlwEs3NKX9v+6J+mT/u1PK//qdOca/B6L/Fl8z
caH2prYsAdwqBmjkYfgaOIk1uTr1LFsFBizw5VcAPTBIddakfABzgTtIyGs194oH
9vvkfwFar6qbT6s4sNNklCZWfYdUntQwCrpMPw3oPqcL3aUk8vIHoz4bDq7UEzBD
8/DEirPnIGxfxxcM4zVVUq0l/bx6oFWHXcSjSH4rf+enjAXM5+A7TWgnInNMIhxO
+EXyttFXRkPJHlbipYALRBPKEVjxaglqsIn7FCL5h64p1MyP7UoS2UpJtSSweU6w
BSi1GO3jvbiFU1nrxdqF9P4lQTQaRNgmsOCvRmxrXaHjdC3ngjMhWncR+GBp5HXR
IdiNCg+a5jcvIsrRpUXa1S6NkYhdBZvFgNJF/3E3Zm8QhtGfYvsuOi4BNPRp1ABI
8bZ4hHAwLnfniJJ+1xCY2VKZy0bNeLJp6kpdZSEzK056tJTYCEqbWZ9Cif0bsHW9
yqzoCdQ2LHMrfhTYjJ7d5wN3iHtVNIyVWXyLtpVL6guFlcPcR9gvEyyJR07GbFrk
67yQ5JVndQhr4kovjELtnJKSqiz4Mpxn0XFMEzd9czNtoLHz6cwU7EThiAC6+rxn
yedKyjEEnSF0Ox3Gu5FCLCLiWzfwTFTvf73HRGC4kkj+jKGF920A8UnEKHug8kxj
pN49y+8zdmoaAi23YDshEp0yZ2jWH7+KPyCVgeh7VvlhEuBxoc8BDqP9eHLBkmlE
EtsqmvtmXl0+3CxmSDrApXORKy1TuheukTSN1myClBc=
`protect END_PROTECTED
