`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
THJ6v86GNb6otmyP9CsFR/tDwc5wmWJzmYMbt085nOSUNwzuQFXOzg/JuIn5w1Or
vUv3d1roT6aFyRJoLpZORROtJXPT7+o0BcOgUR4OSPbVkCecKFRrKsikVMo2lgLP
BFyxD6bcU1YldpAO1rnCSZC04H3waqqeovpo6ouy5coSVWX6mySyEZE0oxaNk6OU
Ze2cR7ZCnk8r/zjvmr+N5ovI9Q9m3hxFx99VpIkQersQhL8IZgHOMPW9hfMAk+J7
D4ZFdasivdvigmPpTruf/sYi42Lhr/YOazeLB58MZILYh1BtblZFmAiBDWDExtqO
+9PHeOolai4FQKXed7+9tF4pVUwNaLSMqnxCbo/hJrK+XFG3+x3U1GSKxgF0+Fqc
E3bAU7ctAZWA0o+ymjTYjYCVIF5VdWwGIfMXczzGriU=
`protect END_PROTECTED
