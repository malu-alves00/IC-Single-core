`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lqMKh931lEOdRYYTWQAPSZvK37WogLF0UG/3D0sXGwriWbw8N+Kf+7N2VQ2/chqU
JbkZmtuq7HfNPuZ8j9TLhuhtTIWTpyPUfAKDK0+VWOqH+f9fTxwEjivaA5aIUpEx
YOW5Z2TKCiFB/jIaLc7oh5/ZuojP1NF9yTHjIXD4NcxtLZHHVbl92cUlR3MlvFaZ
LXIVHDpOv7HI9xjib2+Qxm+90xkyrRxWKeEWnUljlpC0kVhe28nUirTjw7BOn8n+
WaYxY4vaCwHdhZkIX56rhE4Ey2qzacbkcmzqssUuxW6/7XeW74GIPfee/o0usws+
Dy25nIWo6K6IchyUrBWsu96IgacXMFz+7z0DC467hYkfL6Bc79QWMNftZ8N9bD4P
djQ4a8G5ciw3luUlDssmra6U/mEnITkUV3yxNrBEhe1GWWV7Srksl1+5cSkIXJeC
06uPLEb6d8HlWk3X0BZYiSTO36PCFWpD3jBVG2qDw/L8XuYaOGgBp3XETr5KYs8H
LkCVdUZWefp6qD7oKpk9fqIxPxgaeY0P6l8EjcSK8T1P8MyE6B5nqwiXhaRJO+w4
rGlz3BEaLhLUx8Vo+LhEskDTT4tBYqnyMnIFRMuUK7rDESwe1vVvAqTLaSZBZxEu
/oCrh1SpbBuqLhKf/VkTtKryYehMs8UIW2yYzTsyjI7TvSaE93a6rxAN1yzX9ybc
bQ1R4gC+qc8ZlueyLFY9fH8HkbJjeDD90C4S413H18H6wv7hJn1+HGVWvN1nwrCG
0QV8w++Mef3PBxkOlUtPMCMT+rakATFq31I+hQ6wm/oRsR0mX52D3uSEFemBBoU+
UU3kUE7cT6Df4beYe/RApRCNqVhAys4S5nPgMx/dwp9AHfyUoVKn6ragcq7k9ota
ThkqDrqWVFys4M7VqFf8vAKXST1wn4jNobv9XQvpMj5VkgoNKDD6c02EFL3zKqsI
FtylZdTffz8I2C3H5vY8IL/J4LmURW4d57tih4HNQkUkOtwT9fC9GjdANr94FarL
1nkTjIN3EMaSLH//CDIwhx6EmPLUpwLgGNVFVtSpQB0DOBofX+pT7A+xdB54tnXX
jCCgCp9CO7oPA47MtAPbnvLyMuXZeP4BCEAUjfWnhEvxX0d8jN+neQDFGVtKh/j7
tcMMLhpHp1p+Oi6mI1h51KhY+qIICSv15VMu0m2rhO3xXPXALekRcmDic3Eg5HJk
iovJs3WfzLDzRmtvLw+EKpKZ0fPbiToKN2WKJGvqk8ETjlnBbYXWBho8OzUUyW8X
G794vJBcrhkwVRCaq6+WmR/itviPCxYiHRCXbOpV+EOru4+TvpIXfGx7hSoRe06g
USitilcTkZcckgEC4YcojqmowjcSDWBM5M9Suuj8V+lA+grXXEoKrAYXQmTc9chi
4R2i9AiNb48BFO3oVzcKUyYJi63ia5cOWG5QoxKLjoyRbY8H6eOYs7flPqvqVUIm
qqa1v0lhitBK4xSzXWtOKg1jG7hMdW2Nf+fn/ShYaq5K5tl9hn56dB+CON2jhWQ+
BwsZYCgbgwDotM6mPphFgXbB8/g8fCwU7NShSeK2F902qkTx+lPpRrdgSjoWDQP3
rMB/ldv7Z1yD2JfVnDdgnBF+de53tCVyVPjQEV2lpxs0Pt6arpxBX0Ngf7lW0vCG
s/k4IjKixlB6l5SIxW6TbXCH1dErkRM7Vm+0WsUoPAuipjUGHfFF3CvYaA2z4RQB
fp2XUufQlkgbvlPX0bVDwHMH78l7TzGJWpmUVWLQPUVFp2ZEj6Zbzttco02Oht2z
nxOyQUNs0L0YrndDhVLx1mLLqn9AVnBzXGxvstKJxDzm6brYk3/m2R29WUR9p2IY
NLPxmg3aGDFhT4t2LS5s/TPBtECXSfbGrmgUTAbGslsLlvAHl2XWHfRIZQ5E/pGl
ABjaqs9IyWVbaHHSZMNZs5VF480CtS9SI0elGARCN4Zao2da3zAbI1TtgoGGOoLu
duEvOCjMTsqBxXFcpLs0tjR9caiBn+7yXtSMLDAinGgSSPTqC3806J7zYWreXLx8
+6MYj6GSePO7n2RS+wJnTdqytweCaCEg89S9W60sHYqhU59Fkzq5NT1Hn0jSkVc8
zCKjrdheFDih76lzGJZvyQ+l/lQjYJOpo4nrk6aDYBjkMrruF0zTamxTpCeT/7cx
koGpDHrczZ24O7v9fPBJhc94Q8Gm1Br5dAuBWNcbP+Zwx/AKQ7fLs9mNWD7jWmug
3OoOgpjWJ18rkT/F/eatcU0ao5+bGVdkQhpmpVLgBvROkvbFd/OcGxirLUI3I5kY
OpWkOIFNE9K6T6lZnNzmEyIrpw2sKvb2Arizagds/zY+Y6ZjAC31xN3ACqiT9EY+
4sYJFuKOo6Sy8NYlOUBE0XtwBrW30E9Oxon6ODUHHyVSFmcpIa3JvzRSKjWR4j01
z9ufHIHmGcipT2dzHUqJYvbQXBvihOPWtLzW8zAuE/vfSPg2kOa+Yo05282cVaLS
Tco/ZTkATFMiEN3wVZ8RAYB8MoC10nWTnwe0pxEvAgA8ka7bZ1flFC8QjHNBN0YZ
y0KZgzh2Bb7qpVAnS7i4mN7jJh+J6bLPsHBPhkjXjBMdoqIJ/AhrO/GRVHLmWyIY
1q5k99ZcMTBSU7cZnS5Y2qcjjaH9tmT+4FfAUraNveKYg0N7cz8Wax/m192pNJva
SZc8ETqwEWMF2cUp3h3gSjLqv8jVPH0Nc+Aco/sKlGP5SolTRK0TOF2oaKN4d7OH
PjyrMDsdf9XsAt5e6tkPHllNgodD1rTfdrLtzwG/lLuXnpcu4jto4N05W9GTsvEJ
6FWizJPAO23F3TBazjQSBO0bVVmgAmxYALA/3fwa756swIYP7CT1T3Jf+km0Z71Q
lK/UnbpOrj2d/O16SapeZ9s3JHh/MVgnfAtdu6zYW2K3DEXGujFZC5nU1BBmyTK5
IviteCQjPcqa4Qk8oqssvNWSPre82zD4mybtekDDNL7YG+NhGwpRvU2/K3vWIbmQ
tYjrozSwA+m9Dzv1QGjubMARBP1gOC40Wi3LgrZ2MBwZ4cQD/1Bn2n6zj7rZ4WtN
ZnGYXfMBLjir6uLHx1L4JnYkcOhl2vcHYU351m0V3ajiEHQoeXLacIElbwsUhSP8
5Jj5ShFwLcJ+ZALkdFheeXQc9Ov25mzrQHD0zAJfMWVnxZKihcBCEaFR+WoIPmOW
2FJqfuWvK+N5kE14FkV0iW41+vx/0vQW0sV6fiuD3CaGFlIzJq1c6UB/yZuf3Uvk
u3h2GthJ7+Y7N+cfd9Em0cTFABzT8ec0jK27XtPXLTorGWan4RqmMD5f2cKlZ6RR
AlNKzm9YlQRWpU9isbwAIz9hc6pJVOAjLJ5zry6T+dzalX2MQj7q8F899Cocyh4W
Lc0YpkPuf0qRPRJdV0IsjVlHHsWUMmorqu59vTISWEdqOLXLpS6Lyb1t63EKVNlD
1nQxGY7dAsBOLXEI9FrXm2GQeN9TR6e++U2piJK9C7ACIqhWXOSCFwCUUXOhBONY
u1W2+eLw8MXGkZHjNg16YPb0luUzCAMBSnabDiQOzm4zXsot7z1HaMafcefT0za9
T4Q5qZ1pX+GTnJFGp/eQ9glypwfUuuvRNs5ZsHfGA8fDZvd2UufVn4TEbRc7XAIF
GQkMueksNRjZD4lWWZnuIwPo67/reepb8cvnIGR47IfM00YZpzp9/oRwE4Wg+TiM
nPpKf/PUrrWd6KV6FGN1YHVxkCUcx/vrcMAnFXCoKs2vljrBD1g5ylNkHld9sXrs
lSX3vmZ9Bxxc7fs6O0L0OA==
`protect END_PROTECTED
