`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Qu2Ua/siDcnBW7/bpmBtd+zQIRDlOCJgoSzRLRe+1Z+HxA2nBfMyvotVH2+5EMMS
8yGdkyJAoU7EC7ikpNP47azAwXzi7wCdGDqyMPo0lLmFgAGPxSQ26sLzBIqS+lDe
sVeiZe3CNKw9aakdOAbluTEka0yFHqDbXbU93w15HJUs/ZWaQ4LlUo/O3mMasaWs
w4Da5Yi5QyiTIkb95AHjovv+AdBmc4WW4rn18iuDNE1X+YAgJcZUafWrpoApAjia
8vrdju6ksvgdEIaWUrLZ6qSCwld4BfyWhqA2BTK2IvgR1Y+0/POl0CiivONfGuYv
I+QIk7rOTgBUX4Ohh4lz6ErtODRfUxF37fV/qORgcrLs5qpwWLfrQU1FyZewE3jm
Z2zdn52xTwrOVGKOQ87b1sIymNtZpAkKBbeSdSyR3EyFNLxSjSbHmQb8yiPQXenR
FmSVTd9e9R8AmszCXy/djamViW3oeXm5wXbbeR+NValwTy+SVNF/abZzvcTVOKZW
vTDSH6Wdz+NVo5kT/LHiux1i9iZn1pXzYC2XBm13nm87aJQRYUZ0R5rl1QTs2Vo/
UPM7p5SNWxc7OUdCXa19gNW8g+jK873voQU9A8PUVhCleVvbvAGnzXE2S3JWfsjY
7oRoj7NbBgsfvMnu3bW6vaZVHBy9/HxbLfrqzdvifIWA9BbNgDrt9kL5Awf7AFw+
Q/3kVNXrYphn6s0X22r8r8QReQNq1jtp9OvTeWl8F7Z2ANYcszq/cFGq3uf4ISY/
gMIJA0IIq2B/h/4uwjEe5Q==
`protect END_PROTECTED
