`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fVIPwaeYOSRCw51R+rP1VYKBS268u15hqQdiZ91JLtHcqQsOVv0YYse6OSC9TghP
o8qQzdFuTu9h93sFPRiu23tfZ65rq5KTsOL2jxl0HL+4A23/X2enANG42kvo+jMK
HzmuSH97eLUyN5D5SPT8lHKwh3E1AaxD87rMbEKv0EWRLXqSonVm+Yj3icn/StSc
c48uXGzvHuybJboyB8xToWEOsEwuKYKzKzpmBffxa/QqlEBtqofOKfZZCuSdeOQn
DoeYMxbXP+m/vmBQvoHoYbDed8cSLp+6ItMkn7Vzh3utOjjJuRWtV6SE1BmN49eV
uoynxe8EhR2kRcCIv7ltSpsZw1w2X/gObQZCA03qsgJclIvbeB1V5PHAJ1Jddzoh
ZkWoe8v4Q5pkpiG/U4EgZykkcUwAhhvtstelKwrS1WCZmn7TM/Anf+K0XTYyLCfB
iHlJGhSw38p+pPU8DEyQmR1fdhBvx/slxbaJA1hHHZQ=
`protect END_PROTECTED
