`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZIaM5NIvIurBgK9ntSPDg1zAobVp1O0nuHYrZ8cqWHSzUb6UpuU54XmgYPJh3H7s
ornjDFqLhxIQeeGku6myn5FIVYqhXO96ZfUMTQdnQUVpi1aGKCKJwdPNwbdO+S5j
10nCucJ7ckRn4S1ZhiyEpcv+LAKVshxz5uCbpXWZ68REGfTvHNx8g4istz8zSvMD
izuKDrL+4zGtbrvXasRAHgovTSGJVh1KYOCi5R3WN2xWqx685DET9TIHUG4cZYYD
dBlVB1UdeNXhPPsMpbmgQVzUqSzu29ZUkS7Siib+4lgoGS763o1ZtKXqzKLbGLBm
G/3QaQifVfvpcPHR3qB1eNshX53Xwe8EMQTXMbrcp/IQZK0P2baNT7ctJWXStXVM
u6NIiXXYwIQOnmg4en7WOa77Hseah0H3ybLl2HDSO0zii5DTj9FhMlR9Sh+pvg7W
w40/Pvy7uYbB1m20kwC6+Z/qhtUWCdbNcNNnUdywiP7KpEQI7eF1UvFwW92PXw+G
wr0nn8xBNnJu4KlhxuwnJanf0okX136TLL25AnnN7lV3JHsjGyKRtZ0LUiHE47Ep
9QgxsZvchy8rvt2hF1ZCGzpT2iu3IzcsDGUxlwiS+bBqwacZVq8n+U88/BgVqvhQ
Y3aMx152Hdd93YCXrL1l4p2xccV2B7yX9ySFWff7jmjQLLRPc367PMQgM3skpqsU
`protect END_PROTECTED
