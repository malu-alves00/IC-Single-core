`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
i7wFYETB+DRe0/ql0n3vqDYkhsBpwyCjFzrevo86+NZkwHhFnX9+qnPm7K7mHopR
rVxInAx0uTaD8tcKWSYE6fDrFIL8qYJqjusus4sidZRVYH2ipGmQzE8YWxFJ7W1u
FPOZ5Rx8PcoXyZi9KOKZfkjv05VCetV5ImyHpYRPmwsgkSIN+fh5Ba+JkRiicr0+
wxnR1KypHN99nvvstqF8InPQZfoCLKjy/EMHlcCnLWVal/sYK+W74+hqlSO0mo/Y
a2k+iOu+3vq15bxASyRHFxf1BAEEO00m6E7lGspCPBCIuT7nRD9PvviGsAUZ+Vdj
crvfeNjz6yLEBlbT89VbgC59uTdX4E3xweGGrw/3JjjIXAJMf02d8VbbJ3VzuwT4
C/Cb9PrMPCv7IEsY1nmoBad09LsAGrTrXu6uab2Ti0phpCQPr8g97DsgS3zyOf5J
6jIeaodchHQriDfv2Av1H3vGgnmCwdcV/x3NxABYFB3u8VEsChPeKS//pNyhkM8R
XRzGsFfIkufqEAmB4aScIoYKtWu70WPg3MZXTsJBL7Kj3IXFEYUwuXc8sZYdo++H
ceKfsGnKz1Te8e18C0Sv/K8aO7oIFE6X4UnNNsl2zNnMNKMOw7KEGH6/LM21RiS9
z7rZ3A+2DE0FaPDR7Schm94wkSi9jjQhMjRCyToqg7rAi1TLkJG+jr+W1Hj+Oltq
sw+LOUkncc3p2OL/6FKmfJM0C3qed91uvP+5RA6LZgahzr/3XNSwpPRxlL2m418b
rucQMx4T0gdeTTihxcJstAgxcAREJKrWRRe1Nlhgr/YLt8nShD9EkOkdLgYjkbdr
/QcOrjGlrWkNkZHcEviOAuo8X8i9uoUdXxfmLDexT52ggBBg8P2zUBV06bR7mF+C
OPcd5OMVWlmxXAhqPoJQisYy6oGUl0PG5Of9G5AxIKszxE3rsgMpi2R45XlWvLh5
b4xSBItVdE2oGG9b8iE2DATov4yymIP1cJj6+gOLPBToYbt4kxmWz78h0yAnvDZS
yhl5dgqISh6pdY4CBNyDLQQP8mJCi7n19OP2X9GzTRUPBM50xJYwO8Xywl3Z6xar
b2Tj8LWNS6BDpwRLfBu+LhBGPQihxCVbp8VNcoROB5epKGs+mecagrSp34ifM3Ig
wUoJ0/u0HIKajJEcV/Ikig25TfbcZCS6kIZYuAsJsFEUlowcjLxcXossYwhWC4SZ
RjwY/jFJT6xjTnCRbhc7cPkVEtgi7fx4ACyKJAgsWnYNioacuHsYAFSAtmmxcEEc
lnk1pNsAntWIEnmIBxSRW1NqXz0Gyq7b1rjlYdy1ADiTuRKP/PbG4Qw7Ry5Zas6C
MHZM4a1AkWEW3j3aV7BPaLC6aRX43jMDJFT1M9onvC57aOgiDkbFZ/YMknb3nonS
4N2SS6SvAtXSkFVs4f6kb61Mg2NdPNnrexaAtfPJJqAMkHR0keuAwUpDRf77dIUb
ss+kcwOxPYgR3SSri3WkodpzUO8sGPp0nKWyfXXOEUtHAXRSKU8MkQNu6mzK8nag
y5qLyrpNeVag7px72O4ddmIRzbA5B+UIewoS4TF7xW9o7FsT5/Xb9RkTBnwxlivN
xtrXWiKhNKY/8+3AifIxCBIgdpRsaNeqnLLLIo6urB7gucqFjupODIs6rAZXXNTz
vpWjzrNKynCnlCKSKttcFYfum8lvYWD5IFLi0f6WKELzhH7e/sTPrtgmkBB1wT1f
igp5UIWk8P2xj7ITSpKtec2o24PmI4DG1FvH6JFJ8ilDc6F1ZNRXpygOgFuHEOp7
JXzPYzpUMkhjBQj3Y3jnyRqvracR74QI7/aCI+vseY5vUfHPL+cnnEGyJPnMylT2
T2Fj/1VEngc1SpYSR+fAyPr9W0D7UhFzhni4GDhjvI1KAgoJVvlwuUBrRbOJk65j
qeYUHyQAzUHfj2jSQVMggTNnZFqQKjS3QLZg2at7g23f7+0f2H6VR766uaZiNLNU
2i4V4RyPP3EuEeBTyRuwfLlMXEly8+ie7nXSM+zhDMRXV4vqoXArAUZ+JcpjIffL
WRCerBZkp21wt+h/QuPWEGtqyA4S/7yCGYbIUUS4Yv80yVKO/I8NtZieBVU50eBv
6DaFR8sebUxhURyRiq0gnoBjjsQ5XBO+XdY4a7y8GKsGPBeJkiDBG7ZCOSHngRhN
SW6ItYH9wt6UR/mGN4iGqMBLvBF1hKbD5y1ibVDCRY0oRXyrye6zdN79wHxiSE40
gXVN4/K1zvLzxyayJayVsKaESDbxOB6/qMHnYDUL7nCvJklHID0RRnxkRGWPmV+B
CCnjhyZPpMmMIKwRV4OHVqUZy0A3xktps8VplaqEY6iX5bz3JLSixuQF2GCG4oFL
IvsL4X6K4EZxA3DfsZkZSuc10fwAtIv4lTEyBKWRXmZGiVevZ563rTHzCIhjGkmu
623FriO2EV3K2LZTHbLhr7ymlaLapVUwrl3Qhdz/YukShqJL4arPm0Nt+x6NKZwp
M2uiSqRsdmCGvGJWNpNSENiiD9BLP68i38d6MHw7tnaA35NXo4J5JfF3TXH5CyC/
zj2b8WHAtpMgDsmjQg+u9F99oKceKknxEj1paGg21ytsj10R1CezdZBcnvLtzWZS
ahr7b/6ctuRhzlXFj6K4xwL3vOLfA0diI0EPZhSU6ttPq/qod0D0JtUlRF1kdlbL
ecCm9pADPbkusweI6TDDj86PIg1ft0/tCjrO9sLhP1KIqi1hAHgjNBy/dapE5+iE
TtdmcDTN17TPhCSvM7lBSIhnQ8PvD0ZaX8WX2L+DIm+zGKOy+/6M976CxpfSSW4D
tfjQ84wo+3qDPhFafPPtn6+L6oSf1CQ5ZcAfR8NihiU1sh284TnnQIc7FdckxvC+
z42nk8I6dHMNsjn/L7VcqAF7uVQOxCTssp6Ygq16o5jvnVaIv5To8M6ptf8AJshJ
rKAUfup2A0zVEgI7mq98YfnJNQqJtdqdlHXTHfkeJbPWAbtNY5/ICti0QwLhJ/7F
5yNhflMItk5edQUdeWpuCN+Eqq5IJhw/RhDctRP2sBWJQWKp+8p35UTSvxC7oykb
bnQnrFL5X4b/ElrG1Q/s9s0q5meQj6ObV30yFws47Z19I6U+DYjZvCreN0LgcxLg
9U/XFBe2R9zfiTGXLluYw9Cji+iZOr5yTmv9MD9P6rUOf3rXdxT5OHkbWBeh3F9+
9/QMHIx7ngSv01ff8mCl/TIaPsYJlW5NVl4UUWxspHU2KhH+XWgM9qKsXT0f56zJ
HgdvM9MVCQc0VT8PCqr6CVVU1Xdud1hP/lSKCoX4HfsMjyFW4TTMxiltoqrReDJT
SuWAIin7hB1mP+amwWH9uRHlNXYW0GzzFLuSQUlG3Cn9N7sbjhFn6+cIC3P7sXEw
4SLHmArT+yXpc4q/1eC+nC8Fl0Bx5UOeTlymwpmyX7LkyfZWfBZwPl9CqKQdqKgI
BHPZ8d9SvYbPueRjWkPJG9OtKaZMy8CyG2k9IOhz7i93cdRKWWh35HJLQOR/BsQC
1EiRqRB8PKc9AOWxK79fljVhsMx0nYtSOwNKSelKz4q4ByjO092fOcCrjzJrNf9X
RXmW++We7hp8nlct5WAFkeYFxGq7LofyuzU5IjdxgkVerCCoZlMbKHR2uZpjGKgH
+XbYS+mlsPJJZSxmCvmd4NtICd/kKc2OODBJxeqjs/RR6P2dVQRdV/8QHbOpxC5Y
9pRIEW6ZSMDme5SF87xuWYJa8nxpwRS0iejzWMP/SDOg2Voty56eW+/ymJU0+RS1
rIAc+/Ad/fm4p3NHO+KinV//EBZqQvGeTIZV9ZuGmPGQBXjm12+q7eLWYu/+niks
0/LcoZyov3N6+JYkLNBr3Wp6Lx6pMRrgi7LELz/aMeg5kNu+RxnWf7keY/grAvF3
CXZWY4MySbYiayesiS0pAgwth2YZClEkaH1Cqn6PlokRugODy0M7DN+Tdw0AX5xP
eHGKsr0gzCilgRX8OqiYL4lJJlBmRr0BReJ09BbzxGdz129Npi6Z1pZA/4YPneQI
RgNI1UF+0Wxsp2OOHVwF9nUwQK6AOygR3XdlG2TeiNIC+NirqYtowBGK6uAAn7uV
I/ntaDEbYHUOX1cNRCdq2OfrCSL+6A2xQHUyCwHcIb4LsbHtxmfMrpG9rByjJCgw
VIkwbbBZe22T7lP36OFuzs1GNkxF8PXGyZ1A3sM0WOHk7ePEeaoGJ7xv+fnvToAa
pdDFrwJARE8ZW5BImHze7p56YK/lRWYIUKnPEssLtRp2KvZ/e1gdX5/1QHs+SaQ/
Aslr8bd7K8wq4GtekP52JXqf3AZ2loQClMiJ5usQCaIipsQlThMaUMg1d8wrmDaA
3qPwdS78C3kA3IOCrCsDkAb4CldofdgLvjZQaw96lLq4xPqEqJWcnjyC64AgUwmu
f4qknnUn/Ic3ebmzWzlgBXnaj9MludoFE2s1on1Jk/C+eoAEpIxmBp0uDrbN9Z6m
PKGCk07OGBufqitDjJ212xCVtOPl5CLXK7fBYlN/2joEZDWK4AnPtCelMVQw2juB
WJDpUaOptmsE6F9n8bf7X4prFgZayqWKB+DUTwU2tTEAshbKzAZU0ISHyqovK/uf
ynhWn4roCODnkBxZxvnESQbsTxv6NEoUOh4gu8yBQoAk7wvEez0LLzCYYzWr4Xne
xvrWAy6Zb+SrbfT9cR2dJZECHxV3eDuATTReqOyyrpRA2w9Y8dTnoN9xYUcdrs9P
P2HTmS4w//i1pLckg7+an2O0iPhJDJ8ePSiVH1hgJCIeX0X7LIcC9LP2CIJ1y5vI
UwG2aeK11CzbIsCaustRdaRxUKkKWuI4l5j5OSwxuEA5A2X+RqRJ2OM/Nkgycq4g
K48oIJmEHMAXmSZFJosqPwFoctN3589h9Agee9yvuzE6sLD7U3cXGq2eaYG5ghL4
zkRXm0DYFC4wuuApy9UjaEqvThRwhPhhBojJHKoG2C9LkK4/E42v81G6zDcQv5r8
cCmErZeP6aIIsimLCrFA+z8QIVjtdUzbe9JxKQBBGX2lvEu5eXvvZ6ep0oWzbH9j
vajKQMiOE9ALfHZ2gg8Nppbw5gXjBhwsuQXQHszCEVnAIVNzqPKtRt5Bf98p+kNU
GjgNaGdQTc3WLuA107tVnAs1FBdr4zrSeFhObVaNJafB2ghgQWdfM98cwsySlxBJ
2jBXpGb6ETVY5odHudq36rkz1P2flgVh3pYA0cRZ8ohwwYwy8zL6Hsi7k/y+apdb
iDuFiYFdFIoV9/CchZduWEwAuiUidKmSXwv8ENxW+CEYGZ3AdqMaXAzY7bsArzwx
osRtkmHfEEyXvRiw2PZpPeok7S5zYyAf7jAY/+kNWhChS70xW06QjKCgStDQlLIp
W7xl5GumBDd2GFTsgAd9EOXJIhDJkBR5JJAqDm+AFO9+Tw+iY6Q/bKlPW87sPGJh
2URNiUtysPPF8qJvpYl2nrVww7BVAsFSWadWuJCWTcSFADMKR926rdHJNbTodSfG
uexzHsw7M8gZ1uXuF7FTLDhxogZfBSOh6g/AobIQvCDHjw2CH4cnDIEhNkWbaMcl
j4q5CT3wXd/GQ/5HF96F6XAoe2RtKwAEhUBI/9WkSKcL9t8zYjz3l2e+WZx+gWMt
iQobe2C7Uzrkx6pk2maq0HRzxMD9qE7e1TdHZyuvO9Zju8UyZfwc9qnWGUfnM95U
i1TX+9igh6u90FQMiWo9GetasNbEdwN01JC9fc5cx65DtFQwkyghnmYVmOMJV1d/
3/2VVIUVjrvFrksEaxkInvOd1SITKKp9Yr6/4GOYMPd0Qn0jUUG6SMnfbeCtQ4bo
U55v1Eqf7ZvjZQObhBrsvHVHkZpKSWp6dcrOAnHpidu7Vnr0tIaC2eAL1mltbbp5
NZAFJrG376H2Xm+3nVy1rTnSRV1RI9fwm6apjvV3+yz/3Wxjm1PK/y6LH1aCmQ/Y
RukRXbiF80sA72iAXoo717F23U3LXlUGXX/1gTNoBNHzuOphsxFODpG9TWfpyQjD
rJoDAZp2Lh1YMe9HQkU055oBhlB5dHV+vBxKXNfxqzw+CxCm10A47ZuqOsORmuR8
ob7R0UMO17bgnlhBTIf8p67QugCRtJrO7FXwYGhA6V31wKn/bfhrIzkkOipKP9Pe
SSh//n/jxgN9x7A9M99gkurnF69bzmhlQZ7TvLw/mJS1ANBcSonV84APpiHSdvW3
xx5nU2jufUXxX2AnJ0ZhhIeFF4OAlFUahJyk9TMoLB/oTUINtR+QL89axI3HqqIJ
2zjnIErbnb1ANXyF4Jh2xOGikmGOL/xS6PeFR5DibsW5uuAJQDKc1EGG6JtSJ777
QxwUd61xOocKGneAO3k64VohfoFdQIKlFeZz4CpaZZF7hC8t26oNVWIcpp1SERfV
E88P3p74V19OU9at1sFtnv4aPweFP4HpxZvSEE+EnnjcsODrlUxY/AYklT+tQL2j
eW7vCHwVNsnS/L7BjyGTsrlTyQjgz9YQ4+T3HPif+N1wj1BgTu6qnAGxGQkWV0rK
AV5sjoY1Uc62XpyFdVzVUkJea/qXJhFyuHIXQBuJcrsvUZsobnHvTj/eEagZRfvv
HomlHTIuImqkBILEEtus4Mow6mFgstmi2TNGT37m7tMC7/uBpCEpw6Oov8aMyj1O
YhvefTAG8bqOZY2/OH9WW3J3j/KMqgxFSkrsS9JOybteDExb+wknHq9Ia1gPVHmQ
2JyQ1Q90R+OtLqb311ZFqKmxwVFEtVP5ZNg9avEnEFzm/fnV8esXQQIUe/HN5xaS
oiPPDKwq2HVJTR/Syvfkl9Ksb1ADvKbuYpg15HvV2sbYF0iBJUjCed7wzG+4g5Nj
Lvj0vGsG/n3ZshmcwWdErle+zu6/+/LMI+tFGkq+40FRXksRWOTRbpoe83XX79ja
/xEJ5u5H3gd1WeYYw+4e35jpl82TzmaMWo16uYewMXWgJcDP7ZKqZE/TmitNGfhl
Mcqp2DWvl1arfbXIHqxQxSoWvU/v6pWzXwfpb2f2FrHJ1LEVzNsHvEBHYNrJAuEQ
vGSddEEf3qagrxgDAG2LQ+aabwr1QWQZRWcfExspAwbgtNFwl9pMC4TRoKD+NwcS
zFu9tkotPgYYpp37pud3zF5V5yviK4ki47Wz78BBbn0mF524+nHqCDfCydKfUTQu
nqHrDNff91HiWzPPjS8ROe2DTLIXOkBoAd0pSKkaxZGCNx/OFbQ586AkoqRTwKQw
4tRU12DKKux7KWMTEJHzcYOiZKxidczK3WodfakC78Va+7oqF0ysW3XG2aTRBHhT
+g3wspw6d/fYvppigpRIH1nX6oHcKMShgCaSsRfR6OCI8fIGKeuHZj6IC0RerVHZ
cRnKXQVdX5KdlMgFFjfzHGrWIiUzzXGJZsPPaqr+ocAIDHv0gZQybh6/01xjo+Rr
5I62bJRjQsE6kFmeIBualDM86QA5qM7kLjPNxr4eAzPaRr1o0FNoF/Qi6Cmk3A96
IA2J2dAWl1QD1LFsKiwnx6M6F9vJcTJ4Ff/FFVO8kRuq+PZ/re/vgQg49WwX5YRN
pPq/DzPA5Za3f0K+0fRR5RyaFWiYrHFgiHXgpUG6i9gqUJJjaQCP5Rb8O/zg3iRy
86H+m1omLqm/R8q0oWWUkMpKZaYB0O1lA6iHzibp1CmKeExz1UpcaV1cdBrm+yvZ
Ui6h3YMqBvhwmy7dgdSQZ1LhXwMfwGjgra9HcxLzfTYFCAkXT1Swd77/J28Lgd44
EK4nr4oGW53UPgu2/ln3hm6e8tPNo/5GuPZKt1YdbPCgUNL11TLyJFR1Qt7scYlE
tXrQRmRnQvIqCDwFdk59+UUXExv8AxdFGhARSOk9CGUk+Gl6dm8IdoxmPZqVbCFp
14di6haDgo1A2cnM6KS9bFXfQUG56WUOHVTmWp8f/E2flxdiQQiY2p8ke0vHkmlr
x7/rcFe7k2qlL56/BZbmUQh9vf3ldkRVJeyaqrXDRS8wLMNc2pQYIcNaPV6mmczA
UaE0PYVX3pq3mNoEUOv/pbdkGKIxEGMPcpUtmVvCvNK9pjh0eCTTrIr7/UwUfK1Q
Kyd6+3Hmqpz0JgG2jYcEGQp09pXBxV3JkaNHlbUl6+a1+xpq6X+xOGGbRZRYugnx
KpMCDX5QmxKf5q97Tyb4wb6sEwtjW58Czuht7iudD30f8OrCNvDugwXs9rEQHfJI
uAVH9G3cuqdgSbXmyyeIro7mKbuZme5Tq5K1cCi09couydcpIIwt1PoFua5j6GRq
BaCyTaTskrvJ4S35ybc+zSBo5VP29UNdPNBinvHu652U5ZiOQdCOQl1X+sxABUvK
DpRsVO+m/22IvR2D5yUa8Mg4OAkeNPztv6U/0LuMGrjfBJUpGPgc/Wf4YtA3CSFB
ZzT1Ri+nkQfgBIGFimr9u36ak7NgfesTXojYRawRE3Q/pREoI/jFGEryWg4Hrozu
sbQtCakRGjXGI+61Z+vxQMyTp69r1eq5wASMtMMTveuqyGuwUlYvJ62/lXAjGyoy
A5liO34WUyfExEbFX3dmOgG2pKANa2eboG7AmP/574jpWn/u4SHKTgTjgjAp/Trk
h20QIIEFXgUXw//krwAbDsEQJmPb7z5cg6kLcdUuGDrgs6hzWpvsXPYbHHG2KASx
eB5QneNbe5Z/97bIT+10mkyWyeghJXwkVEeSp5zbjxhtLzj8+zHa9ronTymNy9kd
Yl+EHiQh+Zk7DHWPkBH6FUHLSCL1zqn59I0I9Bt3AuSsmFhaI/r3JoysrcaQp6Ic
5AdoyY3oNmJiXKMqeopstXmB8ESugIPNW/2MBB83BmP3QlQIq1ru0loy2gLPD7SQ
cdc2gmpxFvNjiBZvg6vMjDAzbSz5wK4Z7+LhW1X9Rgt4bHQGyQ0PBrE7tMWEZNPQ
jhJt2+3mZZeyxjpewnHebWALfjwnZ0y6TerFpkeBc5JzxYP1yJwRLv/2yL3Lxj9u
PlqlWRPYAiRwQGCRJS77YC5TUPYhCzRNDACxxCwfyJkAkIXi+g/JMdubdNrOq99M
tXdhzTaebYeMgwXxJ5wfcgvN9lREKcIMMt0F7NrJxhopN8+cgFDb44mbc6m8mxS6
mZf1pmSjm21+ZkB74Quvl8hdzmH7hQ3odPNtYOTDvJhp34ncEe/KSuIW3TYgxajN
hKCS/UGPkitAXzVutokQG7bY/rrFwGx440V1ZJTRIF/fI0SAcsOpc86dUiSKqo6f
LzJl+nSlHtTS1j+3SJJluFFahHPgNQQyNBHPZ116zjGP/1UMFmlx30IXe3NJq3D5
3T4ENA9zDfUzabJhUzJ4fDCY6PsehpAIg+ulgBVEuE/VSL4Tb1zmbOn6OBrHRvbj
6VJ5MjxnI+PVk5dRTzephDqGVkJ1nZbkHOB1JGoetV8m9NSyd9ozOwGbxHJ25n0v
DC0Nx7ttw9gTzGdd3IOHoiAnpTAua9VxwoO/+e96y2jZYkWob3rJEFPybc2+zkR2
9K8PjssMqG/2Ds540iYNwr5GNurs89Y80jEw/1sll9Xs1frtS5Ol/9t3Ow8JxTLH
RcMqBIMmVZ4QrrGnzoR51BqUiOrz+z6nRiNEi9rr84aWQsqkT3S4rKvWFh3GkH18
9MY93Rgcxl8EWSWoJKhqRVSpRPP3+NAzByKoRDkVk6Yoo+sV9BdDX4wjhJW3SV9j
r96OxUWjxNal/1/bW2QS0RV1fEnZqj1AyB7+0yTbneWPNbmbiZPeftqc2RwmEFZF
M7T1Z9KLjMvzx16MLBIqCy66Jw4RSrnXP9NHxnnbP4wz5F2V8PkGJgewaJlrKAWl
fHXJTGYHLbKe1/Af4j69i/eUJZuFdEuxVvzprvor4RI=
`protect END_PROTECTED
