`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oZQIiCnS9jXRAKZ40i6GqyMIvmCEc6oPNVVw2y+lYHNu+XCVwTBvk1jBcA6ekl6Y
nggmSv537zQrNdcCOuDqDQw2JFkANmH0fwX8laULc9iJg87KqZHcecoWWHUaivs+
udUYHlc0GHUDJ0nulEOe+PC63ChL9zvBhpfK2CJcCYXlOWj3HkH2wdkjOopJyHh6
7suiYin5F/Zyi2aRIC5W+zJcIst6URrKyQaYurfjwPNAiN7y5rGvJJzIBL92UllS
f5AF6ZY4ZRs873tpr0ipO1a6uMGRbfhOVML5SnEQOwmDZH0iLMc1o66rGQ9UxeDH
sSs2v1HfPXd4K8ArR71V4efd/pL7/93Q6Y1/quuqLMgNpd9WGX2CvwSiDy+kp3S+
Lex1oQ2+Pl4YJWU2rAijY8S5VnGWEBet7pxjB2fPuHkTvdq1Oz+CurTh7Nb/jPX8
GNWmUQt7Rv/npxT0x9UmaKJlfeDdARqvxpbfsZINfkg0tO+TMsETL3heoa+h9BwH
bBNPX8b7dSUyQBOKSU9X8rTjVW1vOkNehboMcMDbvSWDSMpstcxFQ44TUGXia0UN
N3D/Oy6y4tzoRARbLps0W6eA/b1waI0rL1jGfxOf0Z/ucndnFIiBgcBdk0RW1mE1
ueb2HnlWj/ddeNMzMqv/3dVPZYDvH7nNNMelUQH6esvzv0FDzRqpB5ARDMFCpegL
fctIdCGtDg99UFsENWV87wK1s2kvCzeqI7b/hCRkKJgL/VFkeoQZh8EGNc4XOQP2
iKsAVAVBKkcn6nUJLJCdDLy22uSaKrlsRDyZ6EmW3tJxNImDyQXhlP1fDFDYjZBz
Glk9e37w4rE7UhtxWDB+cRYvAS5tioEOPpQ7jGnY/dNpYEaJUnIJG/nIjQ81Roj4
3KMw3KH1nlhJby0uN0LTZXgugqZeXoz/KmOQughmQYA+rw8Iucitpq9wuzAn7eKu
VkSjFKE7Yc69vIYK6AYoeJVNGrSYsD1yKAnbilCRvrIVKcY4uV8sjmkOsjUCca+d
bIgGqQuggd1+5oh4zDPZAHCPY3S298oCtIwuZneHO+W7At6tDsA/bdIHnnI/oDW1
ZXUiG6mwMSv8gRiZKRU1e7xG97k4fIqBicROYJoivqyKJg1k9EgDj11qLs4Zw5DP
0V5/ksAi4X8GT7sRDxgZeKk0OqmhiZiV13UBuD0Y40IHzaj7v88JGXVy/e5vq9hr
z6E3oLNlsG5ygSzX3stZw2v8zvlr6gHGC026tVYt1GFiX7nEcjK5rnIdhDeZ2L0L
trQ7UKZtRM9yItbubHxjXwjLOJowvG8Ynll+EsfMAxvEzIHefIaptHbBpStUslXg
ee/JFVhJ/g09T2fO4qDfM+EtALaoC0umRZfRfHH23WGjgZSWVVEuBZObxoFUipjv
26+ay2gbUNtECgaGAbYjgpPzUhi2AIE5J9hMQBBwzL0C2/26E2BSAKnZ804VICTo
sWaLosUOB7AZnLyDsHUIYIbGGZsifbsIBMEOU2et6Oxssa1hIU/xbLgJR0Zx7DI8
Ud0FvwscL0FTLL7hpCjxPF1ml612fxYNdXjWXaWioArLZtbHWIscLVwyDaQL0TYT
jqMfQ0hxZai/QU0G4rSNtBl+maIJ4c6b5QCHcWUrfBIolO71KqJPg5L4vjpI9LXo
RUduD7agckJkeyU/i3O1fVXXGYjbUUjf4e/65aP2HbBm38fe+AIZlXjCjlWoomX6
B9L2MFqwUxKcr0fXVSuh3nI8/rDs462v6opI1ucEc8Isd4xSKyazu8jzn46/dwVZ
W6ckzxMGtInNT67ZwvjJ1h5PBl/1oZEfXcsy/btP0JoiSxWRTM9tEHX8L+PbtVxT
l74JnEScnfsOPdBQnseQJD7jdBLUdLlBJmIZqxt9VzY4XpCxkOcbsgVcPtXiIaPk
NgjOCm1LZ0eUxjCIdtxHgTwaz7soT3SZsp3ptM0r2KtNkeXiPFbnJhO3R9ps5LJT
pO1Lnl4gToNHOMkFjNiMEuS5ibzjSlBE8lWRJZ05UAHY+qXM+bBF/bsXWWkFHNds
z/2CJUG822mmKM4uAdv5XkAnNeXL6sYXOYKT1Rdj3uWjcRGKYhb2bGXX0wijgDeZ
JbEX6swmlJfQVednRBRZ4Ga7/D4NfJd8rAwtMel3OBvss+fGKdv0UBTBO35kkep1
n9HKsmWLJcd25h6SmUM66GZip8XSV/NfiyGMbECi22M8IVinvIsLLORpclSReeXQ
+VkRuG73+Vnx+yWlCJmWpTAVcGYWcUkETPMluNOr02HbcHrINGmw1NLqixUWmsdX
6FPR8lzc0WoRzCrCMI6OnX+LplcUDOLjuCQ+vPMVQ1yNi8XE27AtIHcV73CYm90R
IGE00OWmCsRtJYhA7Bw/9PEtG9dxm5gCoYFE/sGrHQ5WH151yBRcC9crNUzF++zm
unSZg8fS4qDP4/j4xiic8KtZL/4KguWHeV4jeqYuBoV44Rq1wUfBLrr1A95y7iH3
IPA9qQLodGGwTwnf0JFh+ddvWNMeQLqwgBr0JAG/aK8TUc9NB5f0TYjKVjso58J4
BY9FzE2Zssk8OXJW98Rb8VtM8qnzE3kT4DgsBAGVtrrChd3h1kaK/xUcfz/Hjv1G
CjGVAaKL0Sk3ZyU/4vKSINyBlJ7XCS8R54IGX7IjX9+dEwokrPxmqXy7QWw8nBqz
+QFRci5aeqSIboeDfVSzfbsOB3l7o+KcotnXSCY9sWPZCybbqqHovmRaiUuFLOvp
Pez+TTO6eYuERIxEYlHM+boYZeOycDLGYdX2wHFQMKubDhzKqXlRq1RoKd1lIbUY
fNdCGPfD8TIi4PSUf7Nv56iUK9XDtLBfxSRtkSFInV8=
`protect END_PROTECTED
