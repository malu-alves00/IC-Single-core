`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7JxtH6YztT6het4MUK+EIVr8tSmq+Ti0obmRM3IYg73hkCgMfbgzRv6L1jjU1XUG
k/Q+d04ABmYi9sRwfJTplEx6autlGeQYig0iR4kh2y52ADDCcJGrOvGsgfUc6lmb
TtyJFC9k41BP1BjQnYhd0Qe90Ym+LUoGFG5+wfZYTOmVE/wxVzlVCf2yiDyFRNk5
+rj5AmbKSUsK+pToNIQdW96YX5RdOjchYi08BoSpBkGEKrKoyWYmpxFA8GoSgH08
TD4Z+SVl5qY5caJf8wVbXIDWWoVTHa+wgLGC7LetQ/ilSzvnIGFRKzoKEtdWcGPF
6C8mbK+pZ8tskQM8p1FYU+cDyK+eiv0XH8vVuL1vQrZbMjXw2de73aVw+3n7CzGL
16u4I8s8vUyQz2Lz2XLzRQBO2LcdSJFW84bj0FjCvRR94m5EMQ3SWQfIXiXfQI2x
UdNcAM5GF4x9HlWDffs5G9lmc5Sc0wePYU5ClSxtcOLbYjWsdA8mdw4NyvTj4pEB
oNtGuVxkcf2+2NsEuS6q5Qme2hjT5sAym0YTdje20GB9P9it1WtB+ROfQgQEyxCR
1gi2rx4JVOha3dltw3cxbda2PZ3frGMFKzHteCAeLkqL8FT7i5xsauk8FVKYBsfW
SCrIKpePYoN+/g0Z1spTfEpGqtullsPRf67rtuLJf7jlENegdhzFQyJf6/n8YcBB
JiAi0saqdGTQUGwlDxdkNnVNHmvMY2vmCaUFoihvTTd1ECbKTwhEHZvg37M0n6oY
tF1qPI5sLI3MPDUrVS7rQsF+5ZtDnZzevBDJAMjDGhEyVD5bUrzC5MGibrRg8Ajo
DmY20gLb2GGAqbJQ/infgLHW1CfBPtw6/necVnoq8ChXK70lzhxwwq5sI2sA/vLt
xQQRSJdUySDZDAc64EWHh1yan8isj4LMEaUwatD5hikiU+qMhesOYYhm3CCYidRW
WTk7QPyfYXVFUIh++YRIFLNKjOgsQV002I0IomSjcXbfOxsh+CUX3TCy/Fudxytz
6ffPac6/VPWNWt8fpz7M89AFV65OQQZgshdHMdJMtNiibcXFUx8R89UMvi0v8ZuG
rmxn3kQ3nUg9jMIesw1AhjiOcxG8Ej/3D7oVBF047wfQGPCMFi/Tb4yq82JlXxYa
6pLI9MI5HmK216pOjFUI/9OX06pSL8qmLtQcXPfpFNfJ8pQNyAQwj2z/xut9yQU9
LLukp4EOficxDCwclTuxq/goOVD/0+1rPHV3tlhPKUDRCDIo3hMno18gmfEsLo3l
kyfk3I6j1dy1K3E8yZtvRRW03W63pimCFZX1w1VNjgtU3YjIGgpukB7gOeb8DpHa
gWNuOPdVSwf3/mo/I7BnHcjljXCuhmEjP1CCbheL0oeugvlcNtxZJdIYSsHn/7Rm
klpTgUkglEaDtFfx6GQnPg==
`protect END_PROTECTED
