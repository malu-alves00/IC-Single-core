`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gS0hOH7zwlrwLS667vBhEcg6ZlG988LBDhMc7UTZavBeA6G1Ne7w6oXDErA/BjVW
/oeh4jJhv/wgsJfPpr0nHFkcAgHvViPYqI6362SBP8z6ADCvScOMfsT2lnRHNM+p
yBLDMsuXjygII7uMDF4ujEFNNvpNAPhIR5n+qD/hvhu6sfY4NQwNjNW7exgsduKD
DuJqcVwzzDme0h6jka+rE7qLu3fYdp8GBgrtMwpXPBwRNZAuzlJhqutFif+Tp/vA
ZifLYrAUEtLp8OyBo5LaVM+k1s20YIDzpTyx8KknVd95MgGN/x3+mtBt7/gLVwFc
N9DV/DjT8cKP95xj3VV05jkxV8glaBdeyuVj2pMze/La4qantU2gC1kV3Mf63xD1
iy/iFGYoJgE45yEi25nFoWf+gEBLdgfTk/YpAydqFDrKnwhMOGccohc+bT2294B6
9DzFGVcit55JPG65f9bW8/8re9ZZESOEjTnGfD0sB0ez9n7aXkq9mJr40qnqcPoV
eh0EONbMsyxCS+oFgRc8CjjnFPqS0+HcQ6Ksff/TN6Em4dA9Mi+xFt1G7+cKA4Za
abS0DqA8uPEoO94ewNcQ8v9RHrtu5xibW6xdCMobVlo0IsmsO179iLTShmHwZsIV
sfh7h7UX1x1iK0+yjHTmnQjjg/Iel36nh6WfZQgMIXRt2r80h6GUl7pcp1Sl/0Zp
CjIlgI7KBTvCISZYhQNKL5ChAFxsli7GTvRoRPHNiaL5UxexZKJ4Y4A1UM607xER
n1TXRikHg97jcPk0rwheWqvmFnnZBa2FZ7iMTAvtRmN+yCU8ICYMpTzUEpjd+hsp
xrHF5+JGLPyGS8wrpRlnuxcjH0FTDyxznFo6xIRx+uQmpeKycn6lX4k4n/oFw9Pl
/mNYBSvPRU++TRPY+bj++QBNiuAinZOileWv2R2wrPjgAAoHQE/8AXalXywHBpvQ
QZVKSSp0qglpAvIlAob0WIf84PENJFvj9BUiUMTvDZLza3R/lSB29Jz5jqh9yrmT
+5SoN9RRiiZOsqMHgtZt1YcCzi4Qs+83j1vfhPtn7gZ7zssekDK4ZDfTTP7ZINO/
LIHPhWoiooAYQgF++i/MrlJBLkH7ALQ2vMBO8QnAhwUr9/7Ww/aZm6dWGLbje1HP
2z5hTXhzQQ6A54GkQtBeyIaBji0eBCzlkD9ENKpKe4bBhncdxOqnyMQPujSihCnH
FweR9cOfXicHBxlq6OFH5DXz480ap2caFBJVvmLtJTyW8FpA87fZC5+JPKxLlxkH
Cn9SxzdQL6Fa2FDnrkfLUZRuk0iSYdCrmHCyfY+6xtsxSZi++MixajeIDXYPixC9
S6ucx1QBRPXgZnF7bjJpIXpHhLO3T4UWW9fk4Tg1yndo4hr+jqH0sJa4spVMM2Wj
BWSt4kjTZdY0vSCS4V+PxqKnnyY9k06vP1p3DjWgC7HxI+mDvPX5qDlkmww974IE
7FvI6aY7gYQ10z7kw/4BJwA3OynzWXeaXmxfl2UFWOCSJBLhN3GYNYSl2cr40wYf
ZlCHErJKlJmwPQqkdiytnoVxdMrp06hkCYzbx4b0juQ62FgGLMJ81mNcFFS3N7IP
gtQqltxQXZ0UTcsfCVwCMvWx+LTZ4Uy0mpgfdBtzM2anQwz+JvgX3LIRUJCnAUrS
WfOgcoY7abaJPtUen8NiVHsjhBqgKVFJElHF2N7mlQTjRSuG80rf18XIctroDDBU
`protect END_PROTECTED
