`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MTD+KVSp+K0Dy2WI6bkCF+z01uC291q9jrUMzqnlZIqtVzJXapCKUKf6X35N/DVX
zA9qJqkzHJB/VeHrIM0VGIZFHvk9ORPRolm64I8HM/9pH+QUlF1IQlJalkiYbrm/
6tvQX37jcov+EtMf2Ji9eHKVXlof4ueu33J823+19NBCAm0dbVun+PgS45jCM2Au
jA8SWMA0sd8s94zl79gqztEfExXrL8vyCtWzSzJ9X+pyfQfmFxVVRFum9Ax3/XjM
cRUWQB/6d4t//uw9LVn4Kyc6Gj0vvZ9n/4ITj/2AQpvo0y1+2poOAomiHhog95BQ
bbj62CJurIcaVL+aaMYYteNYTCQ+Tf8EPBP+lB8LP4TExmFH7nQXVZt6tmLOBrx6
Ka2AM7pDNbI+2VOWSbCR/K79K+GukJY4qcrk9SwaBtlb6knpQkQB+sPBxenD6UJh
3fLw5TlE3jI/0Fo0IVL77W6DyciL3A+1bW7Oozezbs+YIc11DbWLcJbTTpeAJlwO
CVusM3w1WySutjKUUU+52PJpGiRpIKuzoKj4iObdikZfdmydGfF+fMUbTeYSo/qe
cS/URFa55vTEtljNdpNBQP8o9b1rfgUKM2uf43IlxI/QK0vJk05W7vMAhzjReCLR
t054UvD2WmUiftSj6wdNvPqgOnyLMbLyNpq1O/UwyE1bBlQRxKsaq0gwL+9eiI0k
WOel3SoeGURXABWQ4CQO5hqn5yZenynpxEpBhgqOLWZmufzKQqXedVu4Tks2/XZs
Jus2r62eobXnarPPEZIs4NvMit34M77G/hD9GgzJ4GOcRLkaMcTQqkgCr25YKe4s
9Z6aGZTwlnrsGoUfZl+LRkTg0G7ofNv+yMez6k3TTzUWmvLj1Cw6xu6RK17XfwfB
LrB0B7B16VWc3yMX7fQ7e2An/RbBVEQjGUPB66nE0YR9GHfsPLLRd8jC1WLj0AzQ
giEdCy3d1o6NHnVz+YavMaZxI1F4ez6NufsoatN47EgOYXPWVXkWi1sBKuz/ScS5
qwfeOirNxgIxdS5EkyFeM8Y9WFqqM+wOVxej0qovKDUVzVxmEQZMojZgLWmQmtID
Mfiqubtq2HghFia3MUl9aVWVN5gW/zHCB4szNVq4Vt0BYfrpl6ooaLYWBnlJn346
MWU+aeZzVXPnRIoDGBHycnvv+WwPBmVEiDow/pbBBVCnvkmY9Q4P+WaMLGYIsV+6
c0UaMeOOKsLIFs9vMNsqaAmqm5424hOW4vOIptjjb63vSDVzIx0GnzizFZ6L/2F1
BlBQruHStRzcRu4kvwmwzcS5IwPPjdz/cPxDp4nVW9inpYHsgAeNT9TUfaUzfNdE
VaehpZ97r7/6GDgEKrw/rJdDd7B6WWxVQuKPURcDuoML/zEDUKQs0u01gE/PMIFn
/d5U+XLmh9zhSlsq/fYkDxDNmaqGHsDFWS9PIgv7+YCx/ZriSv6wl/Y0Yoy2djFH
pK9tACsKqF4mSAJHWIE8SihA/nVjB7WB9r59sOFx9BAAAhyFR0on1dcdm6K2Wg7a
r8Y2YFGp0iLz+qXo1ko5aTgagOQxUyUIfW1bXAILjxFCx9SJp6iYKPKJHXz7hZwG
wISvdqWa6/wTmZZf/HlsNg6lIYWzK6tr9++LfifjwmJQBkIdYOF+c8n8ELMUsBNc
u9lsr7agtaTpXUY7xR6itRnODmyQwT2+WqdwXdMfooHLLuG2AxR1vHikBDOLLmYN
Cq70BYEZ15BTDfasmBivGVcFT3whF0cD9c4VqzLZOgEiGMZMYIsINztWhEX+j2Of
IWTQFwLQWs9fEpfgVESu8BGKGEF4n3CgShQYCK5aGUczFI5cwdz8PkKzf+67u6K5
nSwVjH9xO8+54GejAcCLC4ovMZ5rslLjV52nikSKnuu3uSzLtM+ft9jbsd8nJkqG
j7F68noaete3jVswtGoROS5LR388NJzqYvN4yv24QDnQUNiJe5vt7AWHde2EGUpX
r8WRvxiWtqs19ot4bgk2pkR1P4rkBFOMjOx8NypzsVG5d0jzXVfzTTvcU+QRr1eU
WuZefMaapw0/tQBsqWzlH/mQNeslCQgl6Xpr9Jm3KCO3L+q0Ny41rYBtFBi3LOxh
m0ymYjZPr4K7qy4LFOJ5QcoZDDnpqLFbabDhzaEn9aW/SASD9cHi4y4jKN1g7Rud
qspkG5kWIRpLYDxvc6Ho9kwe05TcTX9k6ybHw/PvTjkfMCAMTkVaUlrPMQzp8MM+
YDlh8DrKTg1DhWy00impL7ctdHqojQGRU5hRR+HORJ4x4gJ4MeVh6T2X7bWdY9O2
f9a/JUTF1iBL7oYlCq+EUTKSrsn/sdZB04OygwsNLWE9laQ3i4w23ruQJn1KyH4Y
NnPTDb19wkEXIKPrwHY8MNmfek/Edph9dRTt9uLfqxJLJLzj7RL/XEKMPpvwgif/
cDQGSk53Tq3BCcxoPBQw0wIAgaHPBq8hYTMFuMX3WVLQaVj1HZLISkiugBQYdZFE
Y+bZ0icI+VIqQqgp5UpBR3bBmxGYpc8eNbrpn0ZAm+3kG0P+xT6IXwPQTzhJboVd
Oeq78VOT2sK1hOg1jruu+oslVnoaoEM+5PEbIsLhYfQ5ra9U/e15vZ/+zbo10cnA
zzTfl4y+/J+JkXj93/eSQrq0VckiTwup3C/rx1FVqkT3ldo4eLcy+esfxMgbBG5h
HffUoovpQ1lcrqgNaPesVaMAr9UHsaxCz49oBPqehxb6468/6adEfncLEYTEMCm4
i7wf5Cu1/Pf+cphPrKEE7iUtBmliN7rNEpJRZhnwU0YbhsT+zZr5y4GA4IwTQ+G+
8eiEL+xtB4G89pyVXbgyuxABaYRTBrg/HNURUwppm8Ez3IBbDGiqZWzM5gObz8Xk
vh0RfN8IJ0eiIRBKVG0aoaXMEYXzs+e0tmZt4Uv63GTPTKRaa7HlyMqRlfDbhzVQ
BP5LZvrDu/YAO9X5l0sz7Rf5etN2vcBy3pKqSv8SXf12uwuZfaEps26hu8us4tzd
KdjoSv0TSw83RiPraNYBU9V1p1IfE2x5E4u6WlTU6I6sKoXE8+OQGauYPteeE5wZ
Iu5hB5dD4bnNuSZwmLmdwfBI5BYM53tbPzHVE7VlA3OrtIk/ta/drW5BkPOEeTn3
fkZfVnEZA+yYN/pFlWuhaeKhMAmT8047wIBM76yjyR4JxSP/a/JlxEONUvQO1p4G
ymwWHWbvsT/P1LluPYkkyWYaBCfPBeOnyuPX3Y4+ES+X8mO2OxBamLoYuJxhtcw3
LBdviph+FHT48Geqcc7kjvS/A3eh8SxLSGLt+B/U5NIvBJXHStX2BndJgo9gzZmh
+TH5pNtCZwIZ1uAIFYSHMZGb8IzZvN1DZaiQmV9S9UrDbM1H1BrrcRO6kZ9bXVQD
Jefthcp1z7uUAFiCfxnb7OFp7V3DLKpn7DdK/5IfEJuKZ7zBn7aSXd8rtl9Go/iq
U8dWofJx/BIUhF+7enK74tbeuD5s6ia1gVeSUsDAZdVdnf0gpqHlnSVvH+sHf5FJ
u9a6YNKj0nZsckXyybGvnijY6ptLUZEpsNv8QNBAMxLo46CHEc0zeJQzSAfTtDHL
A/j5MmBqVY6nbPajlAT2nW1i8j0rGFKCwNVobTmCtoIPQXJqmElbvkVVQ6Y8pqjO
K0G1Qc1mFifIAo+hT5lB7Y7R+7HzZI7KNIxOa4+VCe7M3xLT/7+33ShNhF4OTBmM
nkA1XH8HL+tvUxuk4IYGJ4aPEoDpcp/c1boHwawYaFmQlaZQAyBctZ38dLWdU4T9
69sOwy2huhYDQrCMhkTVViGvuNl/liNroimR1LOBeWq7Kk4MbM7bP5VBMeucjiS3
lABzt/Wl+qkEwjcBv88Q8xWrYOWEOajv4dePfA41UDlIcHZyEzPQOnbFQQiP/IIL
wwCxDf5k6RM4uVkVL7Sn/+WpdztKXqNDumWCehRkB9mWfd1gFjv62bTDx4nga0Gw
mJP0/PILoKPjvUTmPddAzlh+mrcPA6xHGju/7ck4hIiEUlzZvxbuwJOdZAROtk+7
qRDUuTNt+ENj5i0HrMi0+DTdzyNTZm7EUeZRp+MM62Gk8oKLXVE/Izwm5QtNxwB2
XhTMoYD4xg7yn+0YnPxsWZpyael4MDTolr2dwL4+BOlbz6CZ8FaOtr97bXz91CmE
ZCUcXW7eWvXok8ciliORIKcWjTp//I712kGgdDoKlzWsNzVeoUh3m3kHu7/USzBy
v4HBXb1MkkXm4JM7ksC8xTA8CYyPgE/831qjnJBwwrX6JqfRCxnqmJUo+G0CIFFK
FucwCnhxAD3xV5eXlHU1Vq4XGb7bEmNQCVf/zZm2NsbTOc6/zO82DLMs92Mc6zrG
EDhxFcLkLSFsB0CNx77WMmcU+sJ8pTVpeJFfSLlaDpdRHgRQwV1djRlYZytOMlRp
ZWg9tgETkK6YxYHJ27mBAwajmT8LxWgNaTNlTy6t6ZCevffM6OzSe5BmMJHUCsnL
aqSMmvUKkgEZtTIx5xG2z4koYiCuqDbEvNtKr4zHg7faN+f7uyq0pmlkKDQyJvtI
mLeuiOyuJOygZfKY4RbJjTsVCHZhaA5i75QSNkRHI4Q/l965ndYJ9jaiSzdPhEG3
AtmIdwLKmMJk1lX2c/SQDbFY5AUz/y8E1WrRCfXcnTA4fQNxfTVOLBalprkIwNxk
pAFoP46fJ9lUdjNIMc949HTXNCT/JsleaBVBW2P3jlCMGS61Ti+4BeYJhnKxNbEZ
bsJ/1BOl1ZpRdHNQJ+qVXhwShweURyVFw+zzqsvI1qgQL5WGAuFkRJNHuhpOJj/G
RQ19FQ9jyClwpxmAFAtx6Rziav8agWHqz7GZw04Cx82XwLGT/36qtcZ76Iv7xJ8t
ghIjxKw2leusRs/3af2K0ltee4ABXutMK1giGZS+BXxtXjOK+Tx1I7i0Rzj9oS+I
8VuMe+G12kS2CInsCjotcDFvFOj7afT1n+ByrAq9VFc=
`protect END_PROTECTED
