`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IGYiYcvhRubWPNE5W2BY7CYZA1jd1BFmR7jfl3ArJoUzYBAG5gXQaqrGGRE7oViH
FuHjjNZfsppMWKENm1lnmRjEJw5B6/XMcTEIGdrT9Vw/Toye1wLzbIFk96OcXiXW
mdUzZTk70eGvHvzOmzubxgpO9mezLZBYrhYI+46FloMwfY7Jr1CWfA0r7a+agBUx
bHhE9WyvtozIiDtP1+fPvlKoFoOQmAmvVMWQVwkJ8glzdFXgGmSR7jyy3oKXXvyI
UfwEPAD55rxPsnbDq2jSP9RsaiOQV7EX2YumAZRXpFSiR2lVVvt9RGhQltm4E1zE
T3Cwra/DiGD1FNiftg2/oRlD4UojVnve16kI63+woXs14HQ2xac+JsyJJ9MlJkEp
Yd9Gita5lx6spv/Zfqq6rxppU1oAZrnGe0yLjqS4YEbOCYKTybos/bS3g563Q6k4
BMxVFv3PY0kk2Ue2Ov4QrEjEIKkQ9yxifuD3LOWqrqjaaIi+++7rSBM0OE8IG83L
vtpqQ/HuxcLhBmvvwLy1oFZW603t/HjuBjFkYTik4cTDYj0gV9qd/BizpesWE6em
SaglplNRdvHcCzOHaLfBJJmhqqqEkG1OIgDiT13BoyWrhH7Efia/z4zcjiDBfp+a
vmxWc+9db+HOVR1RoGyCNCFYYZthwNCsJGa6AqbDkZ+Og9CZRz+W2k4AsNNQ4I6L
HHU+7aY2bnCS21g7gFtytKdU2LZOi39tpNjBMw/13L9K4UHPJ6xUDHUiZQBB6c7W
GyO2IT1mBt3BnzmvKZ280TFie9+H6yNXbFw6zzRB8+Cnb/UZNMVqkcShAFGJ3U6q
a0wtAYIFEFXLnbYge6kHSw==
`protect END_PROTECTED
