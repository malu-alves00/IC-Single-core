`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GEezn+oCW0ls7uI+yj5j5K+XTbiSPt/k4aBPBS/GBMz+5P8KmVhF1DmYSEYqITs+
KdbiHawjBq3TGfjDM5TEoS29z37rpfZ2dsWjMsfduIaV2A+6GmhwGmcSt5nbkOO6
FF9lIPotTL1hWN/caejPEwniRRysVZuXaIEzeXHkiz2m9YPIerAZ/WY67T2dsQeg
n8zREPz/VIgfcIzyJXTJ/MCxPCXe+pnjWbacDNQ87RsuPVnpZW0o+ke2zr+pYC6z
+sHva3/6VCHrw2MsT7k6TuV52OmlgpzC4mBFy+xhZvBOdmGz+U4NmaE2Tb5B+AXM
/ytfnPM4dKxCVqq/EfFq0t7l1TVWzIz5gNP7EUHHqUSAap7Mt19nYgvei32beDC0
LOf3XIsL33n3klre+ZWPew==
`protect END_PROTECTED
