`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fhmQOaKb2Z7MsZJfCrTg1vvOKzahc6rplfJ74kfUwm3ozDt4JOm+y77TXMB4rcrl
XUguqOpXpStoE7rkNKSs8yVXSuVvrm9Ah2DR4RfH+JJAUsjdCbkWF2SoWEJiz/Vt
Ka4PHgxH+qINAXWwIZno2Ac82wtBkRz6m0ri4KXtChKGpXo2TEfVSVycHQCz7dUz
cIqd4pYwmJlMnEhbRpoHHi8YlpiehvmP/kYQZLMB41zQ0dSDCYx2B8LfC5q+kU46
z0OQISmEcpzjsOcJlJcyC8kwPklwW1lXz7gmeneRdLfrTG/vqUN83veJ0PwL3uny
xV7juggCvTjD8ttFqta5yb5uWmT4jhKVNTCJKAbo9SdDBPXoK1UT/Uwf1MJW2SAP
TIZO8yUxpxKsSIahFmvoFA==
`protect END_PROTECTED
