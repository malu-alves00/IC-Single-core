`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
b4RKiNWUIpP7oV6ztUGqN15m+gSEP44fPpt3dmKrFAhPU5L9vyhktdOYiNkoCQZ6
tGJcwe61X6JL41pqVB1qj39hdA0CiMcZT25aozK+1q72qEJGEYaWRyu2HekAm9co
EkRX3iMvMl/ZPBh8myEiilDjjjLRS9EEqdZ2e+bpAte/qJEMsEhUegrC2mkUYWTP
S3DEDzUtdJzGkyxWCkgWFop6mn7qb4011CMOffzFSMoZkGWnWS3h0J3/Q3Bk3Yb1
OpsBMDe9tS1B2LYjAcZ1dXAj06d3ZluZ+G8VohNoXGKRGfMZL3AuDjDKjJqrzFMz
vHox7LSr7+YBqRq49I4hIPfihXiLBiKUf8fFGOXjKyXinGjBznEO4KQyhQZbtrZM
JvDyN4l/W1vID8Vy6tPbPl0Mr3LUACpQPB/BA01sdwBwkeLnDOpO0cQs21p7u3i2
9JseyfM51CBONzTrbg2zqThxEJQWi7Nbtk6SDCd265TPQisLro0fHVClabFgSIFv
StH7lhKlqTCCOuu/6EZxteyFfUBdYyBf0koaEctJG9PjlUL0zxjHGoNGFv0kGZVF
vPckkN4YY6OEs3YZZv/2+h5yIYixVQi+SkO2qB8ZVMmklQvNwtohuv5ZT/kIkSpb
BxKzNJyMa6tQrBvA4wDa68Ow8F49xKSJheP5j0KHuDu2p3TAt8VT6w76YXSuM5bI
VUz7cVKCpJbvxwGVKKY7EUF9PglDcnVtwRgcYx7B/MOvxCSdCrHSPNbDC7LwE2Zw
d1pvW35SO0rTRNAj1HGk7d+qW4N4gz3rqbIu6liQRKargcfVXP/7hopgmnZnd7eZ
j6M5zMprzelAD01q83JoQu3HKHkDVqHkT22fIUBFZ8D3YlYbKZuiDVUX3oO/6DE8
va53pPeaNeIqwQrnH5/Qmcg01QxuYcnra84KANC0r6G5zAjt0AQwB4blC34YjEdm
QxE9pXfFvJIJRP28lgp28QrS9jOq11zv4i+gtO3r65EtStDRsqXjep+srqsCcZYE
9ZOl1A07siTZbKFZ2uw8qRN3UgzOliYaMfCq74zKy6DrMKua7C7C2kFFz4kLp+3K
0hmjDISIwJ9d2eIaLOF6WipyY77l10B7UGbtFjTGBtlZUcqeI4X3iFsdgwCZbh1v
hImOsbfa/L9H6z1JQh1QcuYpto1KVQupadUL7qa2ejOtRBOebB/IfC66c0A/Gkl9
Dw9paC/EtXHSHNOwslcDQm5vEhKZXmOZadau+iI1mMRme3llAL3oZ1sytboOXKf/
0jXioXSom8YKRzi91MJ30VM5fzm2QQBsPWQZ+iyTSjFA/QOp5pIxA4T5Ud2gG+xK
uYQRtkRKN+vkq4dG4N7zr/kjb0QZaK+zTvQipJa+SfaBvF5sfy1P3eUk8vDfPKqt
R1LxDJaNt9eGhmZ10uh7OUdQHb5qf1jnP8M0HtO+IEHquzTm1vTQXKcqJ42KRec5
yeO5EKiAzI9HY/h2gk16tqPzMRqp6VVl7JDqo24my0FSKfPUyt4p6MQGAyPuxCtQ
leYd0P0NpyfWlRuPU3npwepM+IHLA7F+ykA6Zq7uvOhrALMfIPmauE1wawg76iAC
8huvOk1/cT2Q+qs5BbSMGtM9gxr7OEIaV03xWLAAXfTKxaP7pjvyo5Jl1y5OGbEo
2HH+9aP8S8ftBmNWv1LGyWJJo+5QsXzD2HoQj56F0zPIKt4PASgxt3iLgBrFVI1V
MzBDwzT57yF9rtWXw4uxd35uq7JIE/bPLs6ngg5dcZPv97T3I5JjpDa/GBUI9Awp
cp1Nq5KNw2SDzL6a6bqQQ3NS4ySvlV/xTRRW67nA+2+PMx2GljGvVUKzmx2v4BqC
LhczOk/lMNJ+1EJCwPZJ8AWJkIFQfDTw9PzPp4ItYZLE3ZkdI8ilbhDevCwLxEd7
LtpxnfvegD7s7EICkTx3AQ==
`protect END_PROTECTED
