`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Rj2JaZdrdrTVlGJBFtwrbZ66kG7c2kWz46z1ZRn5r3JjKjq2fpY0PgGs0+rOl1FB
jj4a1J7IkIFPx8o8/wBd1RbfbVYPfi8D6ItrWINGeuTCrEYjp5qD4r2RbJDYKxRf
DNQTijoD6zFRz6DDH/AH1Y4+SgDDwwdSdZE8B5lnbzCgJZ1D1UfH6hKcR7Iq7BU3
uaYf11OSDEpMCBxIOXK28TkwTJLUeEz54qOfD9h9sw51jI3okWybz8NNpAQGWHov
pdz/8MS/IYfYFsMxAIpe0AAiZDS7yEoLA9GXPochhqZUXJdgNmjadOJUBr0NDYMJ
U7m9wxyCypXrg39C5+oXxMb7sOLPDuCKV9bwnBcm5LiRcZSMaixIoFDod2mMC4Dl
Tq+tgHJ8rNFasfARg3VGaeiRvXA2XpPcfAdK2ju5VMgtu4+A0l4+geX3gbeaJMVD
t0EfYkNv0Zs/HP524V8FjebC/bAryUATfW3xKNeLT8LecuLuB9p97677bR9v61ZH
FxVufUayWgnufUmEA3u+GQ==
`protect END_PROTECTED
