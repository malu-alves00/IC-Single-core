`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gOzJO5mzPp5v1hoNyi/pt5T7OXS2D/oqsP7MNfY0uMRZPE8gxRukkrZXQPB8BVWq
qwRcq0ZDPHL2A+M94xmfgI71ULMAgtwGb0jZFX7giW2ci42WZOkL1vt5zMwItlHy
xckvW3QctMG+478MpRDBUugP8R7U++xWXEpgEsKNwEj2QxctHfzELLx2Es9sG6hA
TLunv7tGP2R+MF3BUha8l+NtgBOxuNh766+Jv/3oKHrcqsHwDyPzyOZKrQoWbip8
fvg5aDO5BNeXDhxXkF6hrK150A4WlALa02Fb6rozb6zVQ9NGkQssHDicZW4aZ6t3
BOcNrRpUoqiJzFhcgm/6fxr2+NcgY1WhX64ulVJj2+CHLgPia/0oqcUHzri7FT1M
BZgizqRiyxCFDbdu8nOABBVH3Xfz+fo5BcyRBC03IAFHpwS5B5i1P1pR23cbNY8u
D+Fe0EnQGod0rpL/O5BLQuk6P8SFNJgfm06ZQXwUMLicMP0fmxKYari5nS34zTbo
WO0BWU9/MM3BsSK78Y6PQEv1aN2VlHZrqI+zKTiMDFtJs3Lt1H/N+HQs7AKGoBpX
q85n/e52ToEBtxYbvjs65TAjWE3wedvUldJsUj8bWusFlbpB6JC0nUILhZ4OIQzQ
bMZOHHEFYt+46aVBIX/n5zCHg2BMFbEZANbX/YjjYabk4F21GghTWI1fqwbyg8Dt
oT/3QM3SV8pXfmqWB1B31+fGS/2Ynh+Tcmw/SeHtrYcaRzcMyixcqLeZS5j3fZVg
eQBl+EMR0jeBXttnZhBI1vC3UHqHU3q1x4SHCmZQyaqDpiF4PFMIYmISccO/7u3i
Qbdr/hhUr3uO1uq58JGO41e5u803o31kEnVUJPs9XTurGZt6i5gNT+164jQzVp3+
EsTISmtPgllvSCEhxJxkT55Jds9fEZKlYVlCAwazU9opIwKmwtixxli8vC+b/EHX
MuYXdlmxv0k+dEsBlh9rGE0Tqgt5dFEj5bVFQJ+8fIOt2vlT2PDHiC8NgSyHqxaI
lvh08WGJnBY4dtzaFkFS/EMF+uqggrBiIAtR+kEzPsNMV9g2ioancaa64MKMX9B+
W6egPvmqnRC7GakAWXw3qFlPkLAELendmDkmzkqLAL8HqbiovTQyZtE7B9pceES/
APd/+/jpZ/fLejM8sDyRVUnk0BWtc3gIIx8YP73vF2zhRUgtJ2E2YWkF3qbYKJSf
YEg0WCqEUOya9uLAwL0dWtTlVF17j9RN7Hf9reDekQJ70AcXqLuW6Y9D2PM674Pl
Wgzk3SmJsOZkOYXFMmz0pFxiZcZTBnVEy5cjfbGkKKUvKcn+CDb6IhQmQHewoU0p
wgCuH5HeKObZVaJSpwHOl8QFxQlZmcBNRq0W7faUGhRf/n8B/xx6dMnUyzs2d4yo
0uDOJmconduu8CGguBaMQGpv5/KV6YgVTV8YF8dhD0qSqhaqA0i+ER6s8i9Mkdl8
6zgtKsEZnQ/YOMlN0aenEZxRFCcMF9sR/Ff4aYC36NjIf1A+LNAjO9T4JbF9lUtQ
WAqyYTTomK9d9SYAHA1ASxXJUtaMPBNH4NU4cDEr4BfMIT/kYJheIZ4VWoGQmiXM
Bj4fYGrO3mnOPhkWKkOFDNrYHe8aCXctJNeeiwAZrCEBcofXDLZPImmQw68AaD53
5zpjq0nhVkrFPnebCMw+LxVGaG1WBdcxn2rbOXXAF45IphR5EL/X5otT5znCqLLb
PVoW7Nd6/KTbEo5BStKc4w7gTAxhNKHtwCX4TvnR0tk8WX8kf46SOstxuA8kLjE9
5Q0e+ek8s3kxF5iY2uU6DG831oTMGa22sZeIagelOQQIYw17QlFygdtH8g6f+QLW
kUmsmgz1cUxMypcea7Qu9wOFwYroy3FQ0VECMdfw89f5cqkQ9k42uPuQkFyWpiRn
GFwiGV6Fig0wuEKoeNtBLbj1LbPB3okTh57rbsL6J5CQfztCnbLFkHt8J6o/BUtt
r3jAUg07XOj4RJl8rAwszxp+SxFgKjhZJ80yJbzVvj2ERqW/d4HRyIPgj1gso7y1
J7YNBZmX7D60eegVGGWFKeG1iIqtx1ZbAzvKQuI/qutPHUo/sMiibvfoq3di+lot
3etysh5TKrtNP7jwpw+t5jXkWV6Ke6WR6YAftCblNOCd/UTVqt7uBWzCIkRlIPRh
NTROL405+fzDxA023tKejp6Mv5E2IOGwd3T8r7ImMsMTeTbeWAmCGZCAMkL5raS9
W3BAGybzK4/U8i5w/udQHSFgBvCtfys9LzmP4M5FR2JOtsI2dwWJnytRHL6rVMN1
a2WUTN1H/DOG13Vl0RaCcj34+fV5UD4uSnybXbV6WWcbAePKsqRf9/Vu4MM0YlEE
AXuU8CPhcP5HurPtTjoWMC3g0JMFSh+7F41xNDzOtQzy3/Rnvxp0uuBod1BFYrwH
nmqxdZH6bANXeKcvCLSp7gnXEJfN70AHGwhO5cl7CEDzP7k+AZ3f+YfQP3MbevEv
TP3OpUuuqz9rOstgfreQzSZJt2jMicEB1ms91/8wfeJm5K/KXqIQx9vvrruPDKGK
w7c5mecrhujTkzsjSDMtp/A1bQBtWYeU2z2rD8bhT3aSPW/pk+vFdHwCDD7vcqa0
SVcPl2B3CLtde+UV4DRkjG5/cPvHRY5dnbNu/oUed2UxKVBOLjAOpYv/4PciSzGs
taQEIBRizaBJ0XEESnCcRdZcPKe9VI9qNT+S/pRq8oSoWvQI0Nfy9OTs/ZYfTmy7
ExdA6/k7gp7OVZ+wpCf2BFLhbULG78AQ3R7Fich/eRHNyr2ZN6wfPgYJt5RqgCvc
7kZ6hEi2FkcaNQ1mlH6gkx7Bl6eiHcFutAVENkNlzwMbbOzZNLdId8GzZZ9D4VQj
4YqKPwltwjljH4mf+AJagMhL0Mth6WPAraPA8+EdA+IV94453wJ7wWTq0Y+XWhca
K0X/o0rPNoc2MKOLwieuecunpf91JYIaTclPx+PLUNFKs59F8Luy8+KWd3YS5w1W
yEC8ckKfLoy/jCBPpD0nIOo8AaB8I58hRpytyxskz7hlqSLciVaSJlIMvevDhy+m
NGNp0DmiLqkZrHjTXh9DMwXgRY8uYYm1CL9bhu+FzHbsz+wpg2+aGoowCS2+7nJS
KKUx/SYhoyydmSt1kG+GcUIn1Pz3m1XRt2KDmfpBdaCXnVm5gcKRML1TZGWFXvUB
b+RpoIgrlKlvwyONXNpuFyRJSU3hGE7UGugnmA65cS8LcmV7rF3UpGAw0AkaZDET
vgxrx6S3njFGJT3JkUYFzu2yDFP41txTjaEke0mlE4pO0u05cCjzULdIWsG47Ep9
9V4F5pVgHl+3/N54YmEJ1juhv5lDHsdJx4AAE3eWvaduwdGS0IrEsl3y1MYN9cPy
QE75T/QgHZgMxRGkiKl6AolV1QxcklCZDZhcnCIPPKWzL/WWFIpKGa67E3x4vOSZ
EjPZCDG/Rj9kPktuBBaUsk3nhyxTIfLHoBUlWXv7TlGE/Fm86nHNnUbEdhJ4RtJA
rzwm13QaATtBq6kvlbgiZ8+/ufI17V7YGROJ/CKYbGJLezqHDxQfObwaeinURizz
4ojbCQxn/bkMGqLxdmgbfdLRe2X1nmF46e+MMdCyFr921xw4miakOh98V6/Mdscy
m51WCK6hoSE/GKi3kWlkFTZnc+hQFulelcEgApwn4XWTeIciduedf4fGi6bFSNWg
6afxp36NcbJxrIbVpUNbieSXYeBMjVzC8K2C8TeBU73LiLFan0Vx7xZgxwDE+gj1
17cUR06kztod2irKG6xFb+3d8bVrYVJRw6TQ4kRdVpH2HLicpWsvXOekkDprrTMG
tlQ3ySVKpoTuD6zEGg/0qZ1n3lVzfhNubbX8TwWDwyTT8mVKoXI40lL7jwDm+3f8
58tApMud+ziJw7as6raYkDMdFV48RvMTmrJ774c+OFpmgeRjFDPNMtOFV3HWzQHN
0wf9qAydr/f/K9u+xt4gViM3xUaVFSbHYkVDeR1nmLwQRqGv/ZXDqvxQR3crzOnY
jFDyjn21fxUJEP5jrWS3iW+tiJ6z9o/eCj8zKzZLChQKBbxBjpscb7WVH1aSq0rn
1zQ15nvPmfrxvATlOLOT5GYwXUjdg73pf74t2n7bDL3DH4kcFEWsliHiFYm510QU
PAIovJ2nJ1QCzt7ykqEdhcYOSEfwKoS9zUUwS08dfFBoUAKquEuh1C0SQ0kFUrA7
zalM2/ApPgZky0feiYozn3A69E+7d6bOYrmIgcejm5gwaUe/hm4L9+RI0kl12pXl
rr7yifH/iQ9TGXtl99Sq6EVmsfl7GxRDj8xKIwME+9T9imVsfYf8Y6+2H/D+lzkX
CQ6o2XXd3NTKk3IoVIklKbWS4nY68FbrT85IL7fgjuKg9FAyyRbUF/FfGYRO5Zek
zPcrg9FkibNy6jIE/JwTOl9B35zJ4hyurXEei96iY9z/qA8TUVqbKtgmsG8ccGdf
VKyrW1Ovp+oaGtm9EacCRin3yeKzThkDD7KcZ2d1HnfnirkA2tCatUPzmumiani+
wqL8y8XUY2RG4C9YxlNqX0CKGzX8JrKJ01l6SYpEhaV1Qdse5EdYySpt7IhUGBeG
m8JPEMFGj5DxkIPJZxagf0FsVOBISJJjuRBQLJWsko6peiVAmo9wCdJEYSL7j797
SPwRkN4x6dayFrwIlhl7HEiaHVMrxAta1nh6lQyZAV7fY9hOUx8hHTS2eZsQI9A8
JjwBqudv61nILCSBwZoJ8etF8huroJ8bzWYPrbQVRLHobDSKOMylgSreJzW3GvNv
qgTcY2u6KE3Ov3LwKzi52x9giivLeoTEUPzO3uvzQyo2uJz10k+wD8koq3kBCbw2
fEBZZZmRl7tXRZFsgSk4YFAjUm9wBx/BQ153IrJq3UCl7vFegpJV4VP5wycFMOR7
VqCHJOPw6bw6fR+ubaVfkAZmBVpAhaW+03VyevcRGXXTuDQywDEej+IR1XiwVfaf
PbKdhhUVikjN0E84z9qcXhgNGHA6byaXMaW8WxaYtVMfEz7czC/q6bt3jv4GrqrM
QaUQ7RLClcbwd9pWYWZfFCOmMj2SCJ3PWtscbImMA7WxmnJp77xx3L44qe4i+HU3
IzFRPCQV+eC9hkonhFlE5uUlfi+ucipG5rDmZOMoGvmFA+eTkpbm411XfaMWh99N
NhMolJL9GcpOeeS3uYkBaGCLzwXmvdU9NCZdPNG3HgxPsSX/qYnPlfiT/3l42BPe
7SCfa2F2ydNi/PSAk6dLdndrzpoGdCQT41j+Z3boqI08sf+eIHv+5bV5gsWf1kWL
jBkiOLn2aDe5G0KtjeL8iVQVkJ4FIw773xccyo0sqvKJn964S5qI2+HBnkgFffpt
ECrNh/UR3F1bV367zAPLEOHRmR7OXp8KWXfnP+KJOHaqoea+fXd4SplxKu0gFdoI
W3GZpK0Zg8QOBTUqnENvKR7+CJGIC8a0DcIr3l0Vrp6HE3SqErctUpqqS4Vuot3o
ZXB2+ifdEmJcHsMay2jOQYz8PANwzPmF/972AAWP4fhTruHstPao157jMo/Zpueg
NGtMDR1lWAEen59GQkpBdI+jlk8rXluShHm2m8y2zi4lHvksI4mMdQr2togINmH/
rFZqW0z3dYgm4C5+HRCk0XbMAc8pEgj3OiorrLFCrlQmC146XxMbTkJrZ7u9bNyb
wy1RwPBVmhgR73duQNJh4b1eAyGgxZjkF2NEEqsJ0SSylq7A5aGhxIjQgHLgwoIB
pPMC5s6zZDEdeZ9WogHP6TG/FyJs5usAiLe22itTa6v2qBO4bW62FuliVlLP4X4o
iTUghxwTWBvNnnJ2eOT3v2lW/tgxaGp8FOjuieaFn3IuYDeFKgUORJIrfX+wmbWQ
le0PKDQ02c+i0zKJ9l7d28D/RRw8a81CUdeyI+dwLhgINEwAmTcrRmZ/YrRrFUD/
YuxaH26DcHlsb1yWsPwRpce7ewwQ2+HSKdm60ssb7MslgiCK3Op/sxksApIYvA3I
0XZB5s9qyZ14vt/jQdYygA2h3qUc6JpHt/j3CGsTFXvPW9USj/c0M6is2xy7HRPl
f3lXvLrdPIdYVLQSaAr4bKozkE2cFSymnmuNNdlpSJnpzPmWUFWF6/K+E80ByUEL
cqZdE5TCTt8E30YT2kCxeu6g80NFKLUesKKSLFk/1OsCEcbqdUk+KXSixb7SUZcF
TpE2LgHfXZsSCA6ccEdfcHHDgXEtFihaD7+Xpd3m79zQkSFm35/I9AtzvnYA9Svy
Xaok+Euudc2WeTgr/6Rh+0mN9L3DF9Rno5gurO2CwtyxxKQTqEpyvliuRu+W2S3A
UB5xVTOF6ywGzUEhYaK843fp3S0MloJZC7ORYMHKbFc5AbINRRkuKTR9ZWIVfHpU
j3ASZZZvbrVQlEjaDZGcN4EuwOmrjmYvsGxnB7Q6sPFMoqS9o30NB/CNpOLKJCpU
38I189H+/JeuWZOuS4HqPjB7GqfgfAl2QGzW3SvzVw5ifUTVImYUnk9Pm1mJQyzb
P5b3HSX6ljeRcfsgdpYC8C3wPxHc+vI3BW1qd9lo0HGu76Su3Wz4lvJguv3uea8T
6ZX7tRiQqUnodpTSLruyF9BmEvlavzkji4OAgba15LZxfXmfgwN7N0bXcTs+DjSR
wlvGjtsaVWWgvbE+1jTLSNW4tTFLUcnWjZRUIxHM5QAaShl4Z77h+4CEa30hdf+B
mYb1j1aE1Jggen33yQA3HV/YKT6ELg6osAzkYbccCXNonZqSoHe0WmhYrF5AgY2J
CmS9c/GvwW3bkMvqYGFLpePIMJGZj6YYl8mjeUjG5sHsEKwH5txVKQxR74HcBTA7
5aO/KADBnTPCr0h02TzIhcD+wpJOwS1+I30MW0AuuMoJbH4ujmOL0E1skmTEodT+
TYDP3kP79xtEtfRu7W2HMnqpXJHKUgP3am99WKcBG9U5qhuZrf7Ra9IS9h849U4P
jyLgBQnlUCCkM8eJWeNSzgFLDVnpoCtb1Ecj4S9M69OI4u+q8B7cV6Lsaws8lAiW
w9ZxeahN/3CRR1gwnRh+E1kGYlMw1ONAJu6InrHeQ7ALkvXKE12zgv34ejDFiZv7
07gXcpm0rF7JYAeaAujjGcBkr+z8U4XQ9bBn2yB0xyq858q/5b//bWy/T6DK8lBd
ofyM1+lPdoD53EN/CPSAczJONZ34MrFyv8yIHBXe+vyNmKtx5GpZb3IJ37XmstnF
P8P2X1XPXCzQlq/IEHzxlUucMNmBv4bf9fyocP6v4XT0of+90GOUG9528X64cmUD
vbeWokRdEid7Zm7r93AAjsqZjIaPqJ6CdtG1ghjxgMtTCtwQinEf2yrDs5iJgvDe
OmtB1QxVTxSNl83XqPd8R6/4r7mM4rZWtoWujkwWJA/WdWUIM47GcDqv7ZyKFDym
OxMP3I8YnFF9UlA3UjCv5NiBCZ6p5dQ7kBYhq6mhbW8WmdxjiNOrLtZ6Pu6ibJoT
5MnD4eLann6AVH2sZHRw69HE2K6ndn9TS74LIeva8ErqV8zNxp64TSI/bnt1r8Jl
6ElcJRsdfhWEBpsxXexRc+y8NiyA64HgWeiWlDT0fumcoFI5YoJV8GOzM9ne7ENW
YuWjBrMz+QyfC9ljsfLexBwG1nIL+wW8+wxvUlavksg/blPC2/CtZ5arkC8c1Ckb
TdxRW7tAHRgqWnIIbN+LFcgMjWmnXe2/e1yIl3+tOKdgM8MUO9Sgw8CaKicP4A7x
a3pHQewSRkKe61zL9XcD1faJrdHDHxhbY7+DOfvk1GoaWON7azxYesdrdyZTp5bF
E+u75e7Q+rKav/gPjeG3eG25bclOHy3VBxyBo37fS9Lf7HE7TcEECuXhn0nio7Ao
1AXZ5eqpSRUnwKUH24JQpNAg6I6qDVy21i/RS4mmf0INOeM9PsaihC5k++8CvPKM
v3LDfQpe9CQadwRs6hIAm0EF6BaiNv1dIEbvZKJAl796DRqzP8ixR75fy6qPx+Nl
DXayd1nR6Sg6jvlVwmYJkAY+bvsClrkxWXpWP9oxBZbNwNBL6UmC65jtFLWHfZZJ
s3EfHTNFsIQu9F0TQD1bhhWoGGn5MY4gTVSp2h0TT/NsMO0JtPmcZO5tGNjsV7G3
UDKhb5OjBmbxtNM6MgryI6qmU3vHNcb97ipyd6wwQUeBg5bs6i/BlOwGMUwCKMxN
sD+SYwG3anJz4b8X/7WA7Np8cs0lh2RRTOwEuStaF4bqN2iw5WFZ6jZpwej5pwNE
kwsg5MxUbVFYFA4S79C/tmaTQXOLo6DfjhEiZltKAmNNkdp80SLdksQXdT9VccHj
nQ49uSiixKUZleqQpZx50rJwfc1ATD7gL5GZ5oLVY4eTMlzTpkdtNRXIcElPNsmc
niXnteszt69kaZj6Sv+otjg1UxaD2Rhe3RBkVKd+t5jQhF12kpR5LqAaZ2v43DhW
S5nNUr3B2Ds3l98uwh2Ro+xxGh+Rad7wQJBcXex1WkzWQD40pN9MoO4n1lSn092T
WDgVAOmS0+ltmjin2fBWDGiw8QDL5GtEbGVNaurh3UFDSyyfaSYZqxYPAxviOeky
7vd1HYPsljAfQDNyC0uK2PeAl1SL2cDiJ8iXmJuq9wUF9P2DQXlGVRpaCD28Ysa4
0d6yBaQbbNFHBDMN5zBXJXZjpBqTgLb1N7CCT+P46++Te/C0mL/dH2b6LhkN+f7m
yptx26voXbc1OfyQstxVqz7vaYUAah0s80vbXi0Wc77M3BtfEYnvioXff/9f+LuB
YIRf3sDVvuMaxDVNIGzmkVi5YNKalNKYHgYSyCTuv6nOFxtR11gB0I4QxqEyLvTY
pDt/uNa3btgsqef3b3Pw7W3hPDMLHu7syPZGDUysH7qn1XE0fpacsYrmtnt0rpi7
JmyDztbIJ422Nhz+79FLyVW/4tqYH1/Z13jQduPj5fHyiW+M3l5yTShF/MbvNPVY
xOWaDb0eW8IvuvZq+qPRTShbuCgax+Uo23sOrr8u7rv7HSU/dgIrvzdGfu67mm6G
CV+8JzSmJsyfUs7BmzJCA+vCnX36GJi3n3lB3p/XB90UlwmgJAf4/ka0dvvom3tp
gIWeicz4gF7g7130lNk1FZierBAbKGhAQ/4rvV4pnAscA7fEl2irx9lQ5Cx0fTHe
DBbs2ChOZqjFUqD6FJGwQxY3CYU1KQHxHiBMtfI2Eus7dkUzNkHi0zmU1QXM8HG2
kAKxiNGREpEh3O8+npE7zigfzADPnfNk73lPFgoSRAn4iV6NjrrpXqBQbbl0fwvK
jLibGQZREjON8ziddTJdjPinZMDmFWSznPIWvigqGw9oqdAy+owSv83rcYnAaGPm
u1PEfcD6njYjYbqlbg1gMOivozdygInNlAK6EiIbvT7p7jaMhydcufHqpszUdbhS
86sKOj0edAFTOCmfGofw9bioPxFFMS2/l6mWUV3yhz+aCsMhJvGwkFdxoNiRVYZQ
WhLTKUH/S8Qj+uy59KgnvwCM8Y48r4Wt3lTSRJEg+5AMjWjByciJYZ4bvdesq80o
cKo+foN+wM+P3qg27xGtcOL6SExPqQtmJkY3VehJZ921Gi+YPwbgDUsqZpf8ygmb
58qKR01tGVnmUOKGiq8pGiCzaFJv3UZm0k3wearkjddKPCe582XVklfRNjO4Mxic
VeiHDFKPR7RRuvPcEk5MM/Km5RhBShN5tfzN2KEafuii+dq9N/516cDIRCcrwXgx
LIB8BVDCaqWuXK2mbsxBluMDaOcZfldGXTi0JNsOrI2v3Bppz6ZKPD0NAyhjPjUu
UDcGxuVRvycuKVZMkV4FyaTydA99KQ87uFme3nzSA/o4MK7AkdCpHgZ/g5imBEXm
q79rionvAHBugay+CVtYp+AfjaRUVKO4gFZ6CjE3BZOsxKQ14NmVcg7T5F63P0c7
Az9oHaLNLgPvwjR5rN0wg6e85zrdHrbEg9b44plpktMrqeCxWnIfxjoPOIR+CVdG
4EjIpTnxxC7TK/SKYSSZAZo4dFQB391zV29w1PzJhe5j0bBS5A0C2/JhzbbmVRO1
ZXfNd40LCBrof/5H5s68zs39D5/104Jn66uONWxYGvjkiPbcdRCP95LfTVPQRuK8
geMgSY+DnQ/mTnOkKqvrm124szg580l6HRAQH+qvS4/JhekQg0XZPgGx9jCzILG6
TRhHSq1t+L7fgFbSljzAp12Vy+RhTI/L8ALRIe8VIEZ6cK3eWwkk/utdLRfUnAT7
g1k/4W2PEd6ECO+tp6DQDT0YtngmIIfdYi3iRNjBit3cJoSht4U25NkBxNvo6SYr
mQVmpA8t19+RfXJP9pMbLiOSlTpukMFKKTzdeV8FRopltANujT40cHpU1097arar
DsIio6Hz9elYeLnX8Ds3Bvun7u2MZ3zlmg/Q5FIglzs9I/pHfcUYby0kah00M/cS
Hz09ELl+cfeoc+iIGNWeq0N9eoz9GzYcJqREnrEeXCKf/NVdwRDL5xrtff9epIGD
0/vfN3tJUfQIXqKfyCI9cQSimnc18OfUwPdD2gjzeFH/VAS+/D5VEpdLb9LqX7Gg
sShsEuaM2t1f7ZM0OVbY1vAiShZPw/o3q32B/yT5TWfqzijw+zpgpMNX6mhUHNAS
MmPcJpjxOmMdkGqXxWRhIhgE5YrDkqw55TGYzXeJ1hUXLrBatnwvtDsdJLR5l7X/
EnVP55hNVUzyTtnJhQHJayfDobH7VyxEhgi0asOV61Z1S68ZeHsYrFreSgaL7E7O
xql41riqv3ATX9JXuX+KzQhC3cr2QdFWZQbASR4iSIKo8hSjwDqRs4t3ydfUl/Su
lfy39w3wogpsTA/GSbMrCMHBJnAXl/PlxYuD2dmr35TvIPrFGQd2ESU0WBy2I/BH
vbLymIDmsWRJXtfZsitZmJS8hIz2lCpsV9+t9+cirAG8/hBIpW9FwBsaPDFE+OPC
YSg2buXX0Z7/dDd0rlhs0lHKjosaZrWKCStQAA2rK5OXANi+MVChnas9fPvjEOFy
Qob22eBONnoLp11zlZfN3QRsPe84uMmjLMraI8913j7IjWGU0lbl02xxp6SVZerg
ZJ+koYthoCfgIWKKG/SF3XYAsbURbAlVon8aGdPoG95qNVIXuNbYnrg4k54Molfj
OjAAEslNvYYLZqBHrwFJCT3/GTf8r48vU8t38uU2xicZ8oMDbi+cYOg54mtuHLsE
BmWuqEhniBfmcZWuC0fYIKV8j+C6ZrARLAAIaitXBAq3Mb3czj4fejzfQqFVE8Js
JCQ3T2N7ig/7Sky1crXIwW0VFScCVgZsj6bjlq/3ZWGwkJGZhmgyWy/P90qH4NSc
LclRcqaU9QA0IB58YhzbYgrAbJVXL+7lFjnoOHkqfzMOn4xeWxBlDJlVYwBHxzJz
87Gy6YWitG76ev/T2LGjlstZ8iq13ymaye+6KMxsRURFfnug3//yN7mvypE2XUw2
SW2R7uijSy8AqmPccgYyYDpadwxBdpxcpFoKtIntKfg0uTOQ3nSg2Zfmjpeis7n9
2xGnAbGZx57dYzvFHk08gu9cpLjCZeiXBsJOs/CNOtcM9WvROEeElrROwv7DJHsa
fXRHbtE3dDwQiRCfSpyvBUUIsrKO2cbfi8P2hAjuYiPvou4ftMn3sEB7mYfhqeqf
EsDNI+zpHOxRkQVAQFgvptWnIlC/BKDR8tYSSSVFOajoq4vxYL63519PAUC2h7j0
pP2+8tQc1RNcvcAAjLBhvuugTFOxPztSVLohHJr70/0AHkgEOt/N+WPpsmPgGsVI
sKayHA8jhIBqmC1VN/VkxelZOLzsnRiARp21c8PIx+rhLpx6VI8t1FT43jAhhe2R
1GuUw2RQAM0I5ZNk2N/DxCfxklG/+f9cavVLloS27IL57GkIDQc8l4yszAzeFpMi
bgAeFVWllt7/dAjDQE523R6yMTLYJL+NJ0Q064Xz4jSOX8kB/lHRfOpUYB3b/61V
m/8CkwT/Se5NvsUiDIIPaglWBQ3Pl5uiD5Vm648wtC24APgo2qpfEeBoD7PCTWR2
QQ/mWBg9QV10tufEVS+UmXOTb6jQdRfW5obqHz6jAo3slXKC7M5rCrYb/VM0rty3
7T0PkURTP446pVyzDbnQzDDt1q62Uu0eLara5dNOO3SIwqKHbvdEqKER8aeTqNz4
ZI1hhlrqqElkTVCxobe27aAxqN+aWN9MAdcBIS08XH3WTZ7Dqy8Unfz7G67VC612
EbXGn3zLN4ZH3GHAjG2IZodaBQG0h17GrFEJu3hXA2KhJgSLYxweGiQmsXQ7Nmrb
kqk3ByhOiQJuM+rNdr7rQcjWsfV4B6wkDOSVK1wW8RwzAGSk1w/2J+EnpDzC5I1N
kRZUTYxOlkr+CGNwvKHTlBhgF7r1F4dbORWrYKkXI8r3g+iO5hYY6HfuDRoTpoAH
VwkBPimyoRDiCvMgFmtg5ts9roZPP4aHgtzrEFEygwnr+W0smLgT0AU/OL6fCy+3
HTvsoIOoS87LEuUD1WuLx/JrIgsF4i8KVVMoCEXuWd4KqxVAPAR2eiDxO+3T/xsp
ZowmEDIRTGJScalUdYVVvew9QvQJv4nqnbWJ5GsQZol+Ua6afXzluAe+eydtzKWL
GUafoDvl7ESnSUQUrmrQfiGeUpqQYp0ZgTK5QDJM3o6NKZgu2scuvi7MN32et7ly
w1rxRdncbV4KKd+9MTpEoGTTWa6XGjWt05TTq2Kcb7MwfMRS80LEkPPDQH7QCqBe
cUCCfgN15KCrHHgWV3OaVXTZJgK3Op9RdkqoEf5JzodRlhYy51ijUstCCDudV49u
rmkt7CZ8RjNlUfauYfBzLJFfSugnvpQXjvMBc+hTVW6Subdjtrw4ZhZUaVtr2N/9
NcVzT/tMUvBgclNhHA59A8pRLQWns8bTD9D/IRlN52+liYv/zPbaEYi0vr8lBldx
EdgWci91ZYLAfmE0pfb8toVrIwYdV1d9lcsTh4LaJPGrStl22qv5Cu73ybw1riEN
jxCRrfmawJu5vULq6V06aqOknTGXVfZmcNVnrJDVSez2pp4uJ+mQJklDvL01Cy8P
2BU3nMpxJWGW63xrGQ85j+RSleb1F3sQYztytgeDXfVsFGS7x6LNqLLnFeF9sY19
g4/o4haFL5VLYPOc8JcfQTPiiLtVMDrqZAA09q1Aam4/6WxjCOch+Pe/lyb9TZRU
WzhlQhUkXFEuURdIKhcVv2F6hsIhabFAnfPY9GjzzdRtuqKJpUuT3U5HZrXH71NM
/lxmQGcuRiRHqjiSbZsoD3UTHbl0CYoZUj8iEuFHXm/aZLvndhOwYfhOBFQOmsH1
yBHTHNR7AM/7UQhBfZcfhqNHu1DeTJY5iocrYKoUOScdJ2fz0lcpPPR70GlWYseo
oUbBF44+ueLioE5y3uaIoEc8+PEjLg0QE/0JtW/eu16IHgmLPqpmGubZZ0I1yzy4
TOqJEvHN8WMShoVWjC+FS5B/2toa/8K1NdJtra1PLxcYLihh3xNQP6gzO6VJUmQw
KRiQcB7PgJobelpmA2us9KqvARDzSbP5Tsfb2ifnkdVqJ2rvANGXIFXZnIVa19c4
kQ7g4kMR9k3Azg5qMpNOCCzrUDJx+Kw02xpqDMZh0Bj1QfHxV1s2wuGOs5SpQ7qt
HKMh9e0damyBmJpdSPwPqDnOakMov4wqgcGib0wrXnEBc5ggptSKCDof5YOCwi2f
/8rLTEQL55mGnqeFc/cWLf68FBzGV9eFV3uIfX4CfqHu8HbaBcfOJhuofgiyTsG5
R2Uy71wUdxUrhMzF0hI3setYhNCkQc1WSHISv1wRrx9ES4TRFuDUuHLQOtx5toA8
ApylHsVQ1UZIlU0xbu9CcGoZG2LquDTg6LDxmiW/+4urB8Tb5wz0AzKc/eopbP9P
FpAXe6xT0Cc3vi0FMQQxCDCABkXQqz10ZcwC/VfX96eilhHJ6wqk0PwUf72PKkD7
Zth15ERQYX+SC7ZJSE7M3wSTrkRPt3ZXKLJFPKNmdYW0eSB7GagjWOqEXvhI4jz4
hOLBg4l4Cc4NqPG9ALEtv8Li0kJdiqKxe37L6JYAT8PBkP0QEgnKmrRMMNdAE/8H
B5comxExVAPhmLUz2d6BEMVk4uBPWZtK9MBydHAYj+vTE2KcZ3UugaovqShYBTCl
0QrLOb+78PxBxM1GdYeRh7cWmeEBzmnzYpZiz2JLC3SmceMoJe5C/rLkxynqenkm
Jd3CzOhUcaUauUTkvsokaaL4L4zjf70GcwTgdCSoGuKfGK7FLVVBbZd+Af/0q0uK
JzN1k6On9KL92TKwJ0KUcT5tG2pYUcUv7LJkJ8gkMgD1dCUC+4JeCuM1ozO2uX7H
yBez0h1OU+vTrt0U0boGE+SluuOuqmcf4IjxNMyUbIfIwEXx3doxGmykC9iDh8Ez
IvrRXbEva3jjqaemoY17MzYLcyyq+RPSRDqkdYmIKa5PeerhwKJ0TPF4CHBIvQAq
dMxeAv+TyapzSEs6SLVuHT5ioBPTzEDsYei0Ig8JeQfI9K7cRAkv2hA2/y41rL0+
CQn5OtnktAYACUZ13nIIxZgyCbWUswIy6JBgNHAyvxQhC3yZL4VcB1cFjzJ65bXS
avEDPYeVySof7GEuQAr4IwhtGsW5E9Gjk6WldUXihTKQd9IDgUdSlYMgx2hhCN1H
dS+9qq1W1htS5DimuFw5ycec8KomgrZU92j0spkQzk0k6CUvmiFORhdI/fB++8PR
EvLtUOi8GrzVR0+FoZkMmsq68xNA24mAUjSlPJimKduHjobVTu5xFPEnc8+JwDSF
WgGugXGTBg9F4BdywKMT1mmCh/xwi3g64hAv3Pnse825DQb3Becc9jXDSpvAwQRd
wgN/HoHfA9IBoOUjHA31lo6U5mRFgwPBwVcVl/qCZjIsAne3lr+hRyqhG7tmlaG0
3HObz6wNF9OTvhdWQwn8bPqKJ6OqVcOJ93xhcFKzEbox94Do3leNejzPyNMp/agM
yG2AIGUD2KQ/luElP6QBoDMgDBsy/k8JRVknEP27tf2gWmwP6mgAJttbXGtdEbxG
N6L7aZ/rixNumgDjUgD2ZPVstloSAAZ5xNRF1Qfjx0OTMB8FBWLNDCsddCJcIZDS
1Ycw3XrB91XwnwT3yfgoa7tzcuNtSDFSmgMA5feujESFCwtp4v6I0uvB3H3cigqs
fLKRfJixf0+qcWpCXXjhBIFPjC4Yan8Xlps4KtFP4lWqbuiaH+V/1Q0d8V42/e3J
01BiA3nZVbSZiIhw3yXQ9JaQDGm7LdXq/mbWaIKl6yzGmVwz5XsNwLModFIhjsQs
f9R0afkqZv7hMKiI/6etze8drBl2nh3ZYN0ipqF6x+LhJp5glmUjP5oHI58L7zHm
EuyyZrrwM4r64NIDgE9LJCZ6e52JzcuGXYRq++GFGZr8XbhfIC8k8pbOqLASSOEf
054drxywozzXep3OA1BEuLyvfHlMXTutQOFf4UbjVCzFgcQLt6RYcgLYBW3q6M2R
ynMkeaYitRbwpHyoU6OH1jQg/WRL8YCW6i8IQP9SFGSD4kjzhFLgZyFV+LqktyYy
+HlhwJoiKU8nmHeA3sLRfyR74uGSdrCtHLjcJWUGm3tiDnZvdfYbsDLJLIvKQ2Sj
+jDdInOTvOqIeByY/lO2Io/X0JhypaBeHj/Ew36oyEbAaaUMnJwSG/V5TC+pGO/K
rt0sJWO8jZ68NyAc2S4r7sYOcewb1kVrnnmUcRyaQIRJDWWXhlBb9odL+8sPgXoz
NiHzD6v4UR2r6JtAM1H0xjq2qMIZdb0/0C62dvpSoc7ko0hod7FQcf3zhtTdNsUo
SEUzcEwBwkUQu1OdbiWA4Y4GjPTuAWw47uasbZyExf+9OZuKT0+ukE00s/jh9d29
WrQOCsSL7Dc0BFrY2r6wo4fNbE+5pSMMI0mg9A7jsvRAxI5unsdCW3G1rezbXD23
v78ixDbx4cDXpzwNLPArv7Qii3wtK9dI1I6smsUswjxZCm1klnohuFQUz9nERrCW
8v0TN5XwIU/svIXK3OPzzu1T2DFrSEeoXHLolsUAOplFsbnbrKUBQNJ1S+hka89F
4SZrwYPh5vLtKb//+Zjm9yiR6dnxezC/viskawbK17Sfb7dlJxT6DQ3z5nNXPHby
078ro4IOOg6rE59xBKktYViS9fL7cXFkN4m63Q1jea4XD3dgJQ+keb13Df+X2l+O
nWmS8z62Z8kO1huZnRdMLdGVczZrhtfuvleekniJJ+OysR9t868rSJ4e82oj0hrt
kxKXCZy7bzZJAnybpASFA1F5Pm/3b33FHpYu48yv1hUT126Y8jcIJ+zBQ5w+jA/L
1Pex/NIGHxAL4HPd5qMW80xDpULs+kJdivUnpIhp/+2tk/Rv2M/Qkp82vlSFrWWe
V+tG8zzoSM0G6v+8+OeKFHFzEVvfSWhAMvNVkQ8N7CRTufofGLvKNAhXJ2LRcm9m
3d2Efgm3LjrsrbYMa9eXb6Bqt8aBJoM5iw5iU+F4G1TEY2qkHvtse+Y4t84KeoeW
8pRvq7V4t2Rr/9ma8mEYVxjAg0Npy61YIXAnxzGQV/9jHSxIK5tCXpp4IEOi9Cw/
nY8hujj5nuKJPLsrnoZQToiL0GZ1G3Lk2McGoMjz7qmPq2x88C8q6wmc80T4H491
ZO0I1jpivItYuWZx0dEs4zL0Lgh+NXV437YOpBi+A0gyP8b7xXCz+FUdyh6BWXGk
N76LRe7++zwWjI7Osoei8cXockynUUMvrL+LgWyKa58XWmcc2vtqKc3VygBt+GV1
+kWc1ubAvQu2I86c0Ql8Jv1xum6VteQ6cJtj0J8SOTerxuyU8KjI110tEfxoftJx
1JmaRwvFKs9VA0ybmkqbPUq4rGeQI9Xvj/oxtTHHh0t7/9Sg3mt24oW4+/NOcViu
BGfyG2QtsKmKE3lF98qTQVkyAOKagoZ2peGjtMWYxZHTBzV0AchkELaC7TCdVZkV
hrq75YaEGQoj0VWLxomyDO2ZQFaZGEG3WGLYQGiYvkfpbAfaWSa2QmPMfMzPZkT7
Gkd7y7YATqfsNZesGVK+kxt3p9/uPqyWxh3HVXFvQdWbnZn3QWW63/iTCrrczGX7
7s1RLrzMSSmtSqSvAaYTQ76NM/rzVgOn5UD+m7/Ppk/PB9ZMa9JHnjW+f/0CfPlE
fbQLLt3dYeZ0Lfo/65esyytZw5wg+Thfp/wtmQ86CxgHi0mgBllLCOjR2X78AkYK
ZORFX5z2/lqyFIz/HQ9d6HwcZ4nguR1fkS5VtKhZwHqVZTdf1MA5O8ERYDux0YAZ
XTWdluBTYXMiauRlc8IptmXb/BCfjXDctWx6sGUkFETAL/ip1T1rJABeh1+xidSu
2ZTbWqwhdUJWbRlbGExuwyDrLYeSEG44TS/lGpFaJjDKi5o0v+MJszQZGZmqldn2
5Axccsdq0kWYeO27gQgKZroIKciJbN9MQm9W7DWNyx7x28MVv6oxhAtC/47euVwU
wkr4Pmp2cbUvNhfLAr8rUB9z9/VG3U+bo3PnMka9Kv3wxdzjlQiyml/fHHNyXVKz
5zcCecw0Cq3ixuKNuR8ZgK2tn7NbnCH8/vuGGpTMM6kQR2f6B/ZdcCYigDtGjNzA
FENHWEe0uhl8ao2q5Pb74g0ctNzueXUhuk+BiiB7ywyhlgOmIG7pW5dgQOgGt/wq
IHqMIveRphM5PE/PsvJ9s5o84xybWxSDDz1vXXtMX5p+/+sWPyYlo8xbIJDcQ/FS
TezLdq93dPbA0uy6m7E0qmpu7MG7mqpFXtfzk0Wk+ngWDRTeh6rru3Dj9uC8EvNM
Or2TGotSw3fDRa7Ix+q/M6hiU3B177G0PwziHWLZ0baYPtbNZNBkCbUZOJk0hcgk
U+n3/F3r9cb/dMg1k1FXGav00lWOw7q7ZLIt22KUda6Du/xIyVWKfdV3qlTaOhw0
fLtmidUQybj7wOGT8nPP+E3aqNKGeETmxepGuUKO/HDTe881Ddq52Ckl1JCF7MfZ
pkBYFRmnC1I1c3HeOP7vdQZTEo5hipjYbrl6gYj6MAAZyhrYXVcFp9brMLy1Lb7L
vErU9lwmd+v6QXtI9cAFuuq371m6BCge/vz0wc8EcyEWZ1EgelB9yn/i/ISzAWCG
1yhUagdpoZeHrG0it72ezIYONcI0F7BinrRgmVo5iFQmDWmPtUt1bV+2d00xsI72
XZ7l/mAjZ8ydqht+JIBmrMLg16sC0FPE9M+EEkMt8YZR32KviYeCJ2LuQCjVtTAS
CEx4/uYs02MIvLdVd9eCB9cpwvEYQ38Mn8nJVCWmHVFfj9r5Q08TpT8PC6SzHMRX
6Pyeip1ffXK1DVBIABLHt/hCLC39Lnzh3N+o/L/Cw/lGwgrH5eLjYqh05KaRGW9r
CmPc633KmItbcc3tW1CtM2mvZmSnrjbE1Wr5O10rZ6onPixid/vh9i6EUZ8skkNG
P5izJZoEGQRw5kkDI22N/WoLreBrg5vLCGe+2CVCPGhBP0nBRYKnskYuoOqWQ3kW
sMvGtiE9z34gnlF2dV04WW/5bodiAuzYAbd6YYG7CML59VlUrl60h2stDPQbiW2q
v0uyq857hSn5zDY+L5HwRrpN5w6pH8kJ8JCXMPZIQlgdqoIgW0jBND+IsMxNbpRh
y+/XAEfrt5Hv4RoYPHW3M4b80/qBHVi7eR8aPTHiR/S9uauLMUqjBfiyUktLz+kE
JH+awWM0aoAxDaUR4SUKhxrloQjVZc0DWDkyFBnIXl8mcDRBrGYHD2Unfk0vtNfQ
FwxS9zisuWUWzoEDbWzdS5872gp1LLLiDIqRR6Ie1gVAP8LP7qUeDPMjNGuUm2Cn
YdPiq9S1u63TCZxwNFau2J/sVQBQFO1DfKSwPmJmI11si8oAMdGW7GxVBkftLE13
zozb0PWk/i0Pi3D+oI1ZWcEobl7j5X5GhHHXoQ4Y20p/ynpsUoXrjd4+JFP41M7E
OK9H9i11CuxB84xC04Kt73A7VMXITlquiWd7XaeDJ63Wn/YOZgXbEDb/3ITxxiX4
bZZk16mV0YPITrC/mrCdWeZXzgtB6OZPVqUPUzf4R4XOUDmKmGLqS+PaF8GhzFvw
t/EWg5yh4jmBtIUiTilUhNdp5mEq3+cd4prKw4mCH1TtWnmG8LdCssJdfT7wnVXe
Dbt6khiXiflBBWrCgxBUufv6fCsw7BDemfSCSN+ZqJJK7DBhQu70j/DbDOVqPpst
3UY7QhY+/x+oas5IPS/gSMsef0+ZGOi4ixTS9tCcjRdby5QYfJ8gDxzLkYqGPR60
UhJUVkskss2G3Fg+zNr0XkFIiJIb3xUOyJyaoj0IizjGGTgM1c8dnwuubBPUbFXz
hjAfMvnogZ6E9ZqIEJxC2Tgb9g4LzJxNDeChYQz4aShdVzsQ2FRGjdUOJ4ScdAeM
XVLp67rGlvMnoOGsBOi3JLXsPAGiAKXJU27wpuDtmr+GaA/vj8LbCvFOl3UDlgp3
DAevn1Zo2AZJ7bTgVYzeTPxn86X+aGzEHgs+RNzUgZ5d1prKtuUXfJA50ms8t84u
9nldQXrqJyjPsBky82ozg4yC551MbKYoV88k2Mx7DiGS8XLV5LNonUhJ1xqco85V
OYoCZ+/FlJQo5xZnjwzbf6l9PqVMdcbjfYchLYhXne1bSn6fcsxGOY5Hl0cyBjNj
5CaTDcZJlRXRvHq3BL4bzwaO50bwx/xv/0LfBbUx2T+xLvYiwVGYhxUxy5jyszfw
vyn8l2629SoBzawueiFbz8GVFP+G5JlcbvrCM4e7K5Shsb/RVAJ6SStvWPx+lDiE
NfHMuQVSybG23giOaQ+m5pwpFrAkW5tBHA6lyKwMFmIQmEG4QJdausPvbiQQvMHn
dtUv0oT1LQyH/pSN6l5X7LWa/2gEtCWJa3AA2rKW3Q4IYpqVsCGv2xfgDwXUbpbw
uCRdSxVZsqQe894jZBQBvbmL9u61wsYjtIOiaRJIoYtKspq4m1pPZUjscUQNFgml
Znj7vbkIQbIX+4ohD4V180oDAON416zpUD2/jjJBjAr+iKxP7djm12N47+w0kIxq
Ww6O26eTP4IwMTFMMHEATCCzDLgLp0Or5Vaymm6iZX8BQJtCP9AYnkCBsUQ71psO
TKCK5KePxEu7tpbUdB5vEHzm7/fsTEG0rwA7/CCaal3QdhyWSW3bjV2+lfvIcY0H
pcFRRv6IOOQjMNdlU1RXnXKuXyfvVwaEY6uwhNlnLhabu6zby2YbYh23nFVj6Gz1
japUy9c8Ldblixj28I7wS6hfQA8qXKV7O5MZZP2RB6I/ck6NBzkbzqY5tsH/z3Nk
RI4fFTMgErQd4xEuy67S3tyI17leeaNBuV8v7IzJ2BG8wBtXkk3Y+TuEcGvFFFNj
WkDvCRyvcr19DtQMYUL4t8QuT4PURLM5nZWu81tomxwvltCOeiuJwXDY4RQvawEA
/V8i5m4P+f80Ry/1ON2laJrJXZoYld6Mg2dINOuAJDGFJJ4/oanXTHc5Navs6z77
wA5u2IzHuGMrGEGOkv0p+X2PPYW87evDr2cgAYGwr5SvvkHjy6r1SkE/D5GHdngm
qO3aZ9sKaUw+KWX+Kl6jaIzlfIWmRTxpkpIlMYuUlL6EuH8AIIk4anWXtRIcX7kQ
nNOCdp4523yKiRvSD9qDr+VuZo4WF9w393AyloUCDdXuXwbT+rH5dciP1oT1sJKs
P4w+ZdqTQazZQnuVM8VPX/7y0xbKGzi2UPoBcpJNHNqUNOMG/NMe8nmuAK0wCD22
Y3y8OuL0nzEfwU/6KYJ3ieo/gWbDIXUeWW5ez1JYdI8N7bnU6ufxl+jMCQx76MS4
qpLrHf3LYQN7Krnu7cMh2WvwmE76lUrrtWHWvzOLWatAAB7PQqmAb7oYGpKODthd
QSgJcIteRz/4/4UHN1CagGgIOXdco3nnfjPo3w4pXXnx9cgb3XLHkDIcY1n1FLm+
ZyIeltDq506mIPbwc6nDB/TxdHUqv0rdFds0wMKXlT/BPKv98XB6qznAHkJQZWXO
0cU0CjyA/x9Guc5iQ23+MZWAml2Ifs2V7NSXgr7RfiIE399t5/Z00Dx0b4TF66YZ
Yc0V4oBW07Qg8Wmybw8NZx4Dy18N4dpzf6T8AcH6C/aQgc42m8e6uAGURfwBUeAQ
bvEWwuO9RmSoB3NN/COIuVJYevx3LtU9kaR1/h2fW8jSF6Xn4k7Hhuxugh2n9yA+
SZKwG0XH1SZ4ydWaoWqLkHSGkk02zomBHO6sjgDC030vgGabx5SurOJdi5em1PJp
6aCdeQqVTD/Js/zl0Mm48OPdwdliN6OHdto/8bgEB32FArlHmkl3nJDip+xKVYKi
UwxezDJVSMKXthxDMEgswylRkAGF4Zclje9akqS61pz7MvvvnBi0qjwtsOtI+eHf
8VqNTmLsq9DPb+NvD49pT72n4fzy79Y5v4zPMA80iPoE2VHNaHtWSXg/7Svjawdr
+z3mXG0Xiq68UKuHY6o1GURZbB0HTSZHIuF2fITdRGHC57jx7VZqSZm3IdQy/byI
FPUdhPSDla5jWvd5wGfEJQMW4czjN98pk523LjCxJmidZuUhmGXaApycxsvVHqAm
tTvccoH9RfBl1y6b0IVSjvs6JeBArv9czkjYEj9P7AAVy4bnOr9tASN+L7UWSF58
mXvz71VIut0Pb3ujvGDK14hTmcCqpSDp4fOXy4XkF7+hfHZry7ijpp+mSo1URUUI
cHVSbMRemvtSjl3pMGUNad7Pp2X6KbgXLv03Lp8EsZb/OmgWh4TP3EvyrOvJr2UJ
O0BUk0N3ZIf2HG9URwyQAdD6EOe5B4lFhR0IIwofYmmhpg2VV9qJ1tY83kL8VLqK
pJmPCrnw2MZBPZzry16W98zb3lq7UghICvEHgRi3zetk0/8CjilbXCyL4NqARN4N
H9n0YjzZy0KR9yfDyC9KO06/4v8sDHbXellyAVQhLjvo70wxdOFj6QCpgzGcbua3
dfze9plLADVXrwmv5NRtyfyp7JrCNSnl0g+PNt7gC7u1okhg7Ig/SlNF70bFbeWN
JBZmOqMhwsaNn6jSeI0AH9tPuFpOFR8mjZSSbELnOO+4dLTGL16qQoYQAqK4Ln7a
XtAOALOh5wuqULrAYDlhzquV4/wt9bRCxbsw+VkZtLvNKdR4QgPKTox9Uo3rNayY
sBOTwSB0awmhNigaNedjqespTr4xlnyYSNr1yqP5kW0B5uZ+0xqWeJMbhL4q2ml8
bK68Pr+Dx/sNi9rnfOkeKjnvWSs/XiJs6JOgpvUWotev2povFeo6D1OnjQUWpCYC
9vz7beH/ylu5utx3EVPq5ia9R9xMLeupZghbH2nCj7+IDn4i7JUQNQLYhQYgbs96
quDMT2UOUn5l+nYivco7LISJ1SFGFOOxWqJrAW7tNubg2YhIY7+fhhD1FwsjU5FD
kShCn8i50CRRoxHQKyvUn/S1jb0dyBoYe7vZD8QwnCXNcYV5a3sB2vf+8M0CGVao
CSLKySQfs/I93p0GfqVAusCs2VO6ouDd1QCZI8t1vWp344O2fTQSIxh1MFjDxr4O
u95rQ7ERn1SBuiSvZOvdYep+pDYFLg17V+qsCCeOabVrD8Jkamm36gApQtaEuLeJ
ff86bViUKrLeR6nQPuh569GchqBFLaDPjVNtV5BV15FzjyNYp2oQLDRfTzPtHGO5
xSuMiz6Nht8iWIWbcONBAiCiyrVepaiM/lZWe6SPLYrlTiC+itww9+kis7P6rbhq
f+q+11htZL1LDwaZpKWoM7xw6fqHXQfc8QExfG29ck3XBmfdlMJRbW/V8wZz7hd+
gMRqjGhkTCKFIgn1OXIthFABTTuezB43Fn/2pgFwNbJENTaUuvrKceSDGsHqvyL1
5pnxG5EWoezg9Z3HHgxJTRw7GoHdsync8p5HHN94Ctfccwz5VmJSA7kbe8eJNOhu
lsRndafBpCBVK+lFlBQSLnAvG0uqpHZT00C6sVYqSNnziQQSFRrIl41lHyHA05h7
pN7p1nVJIgr0eJztB6q8MmPN+5ChxmOnOan5SMiHAaoF3G8oJMlLfrTx7sEKyh1I
pYYBKEo6+3Z2uEyd4ZPBwAWnA8SBQneLoTubaMdQvqyLocROCjfqatv97LUu/1op
0sfMz2Av+OeLkTW2Uu6RdkJRPGEp7Cwe20jKSNZsAH3+uRs0l8WLsxjZ9SE39MPQ
JFCgq5posIcggw91AhOKyvW/qj0DLyHkKp9iRvyUbq+o+vGu3tqBmxVl6qTN8Jl/
hE73Fh1y+GuAl/AK17cVcyPpXeDhg67/ANT+U31U9S19hjUsVKiq4ivGPNlEz0pL
EmPJ++cXuTX7iZA2ANvdev8RbT5nPcufhOaTgCuOillmZrLdu76psLXklpoRGG/8
FZdCTOicZMtmevUpDAErBTYhjvB45pFHL5b48BatVGQOiQyUqRtSXZFjQAvUTH8G
OVGtF5lwg7cVV8HUnAwHpdkJ28hQ8K7vcqma3N7xIUTwlRzJzz8rVYIKQgabxsie
E3BmfwsyRKNBrAlQU04AGwW13WKkEaZfK73GN3S90/k6lAHMFCzSSFX6clTL/QmV
77wS9jI8UzcrQPzcDCrxkFnP0buloTrUkn1snGy/ma6VqPUJTxUdJOhyFG+5PCC2
G6s+J8yo0XZDmP9nU8n16suGmHl4wFTJVMBEWm2tFkTm+iYJC47oRb99hDncASCw
6p+vguc/ysV4hl1gAgtITIVrZ7bdPclGL3pWO+ryBPAw+KaGrKy2964n3HBYhqTc
ijT/UEScnn1sBTpFI/ho1aMyFiYeOjF6x6bm1IIl6rqCSXTLbGhD/9cyhVPN97fc
MvYmWmdiGNS4vpv5ShdZy82Cxz0eVbEwQcYclyA1vxHytns6JF0VQ/lwO7LIi4Pl
jifrHf1lZZGmaxLGGmkUUs1rCmSIxeVa5hQ4/rwQ5pEiPUUt63Z98QCB+EAmCjVK
zbljlwa8RJ1T+EAXATH9SRMh4jQCl83KuA86QJL7b2Qs4Ob2x9oqqU8NoWeAPiIb
dXF3CLv0Tq5PLNo/yBDg2m3gNVtST8ggO25mHjEsbWvJDVvXToFQ1QuSJFKKX45W
tYiMRm8Ey7piHgT4xXZFxPIIKSko/lIge3NnCAi1xfWKs71AJD3u3jb+dh7/I8OO
ZG4xvQuC2oB83YmG5cheTGX1dkkR2LXrc4pCK9xlUaJvzN1PVpPVEnpVhfEhEO3E
q8LT2G6721QNLCAAFolDkBWKUjnddWbB7IohQYg/hE/eca/PTdYIMu0drdUAI+fu
nVwCArgTv3Fmhx1N4irTdw1cLb4NJdQKs6SWnfWwr5Nm3SQHPEN3GaILhjNhSrko
wE1pIsxi6dFqkQZJABcQYXMj0N+gZXSK9OP3tcj7AsGhui2W5Sq94otS3JSNBcYi
Nv3fjJcQetvvn8OBhTwz4n6A4PCG2Pfwgw7MZKSu9U1YeLLpysys34N8/75v3nXc
S+9xaHLQtvN4smkFbs7lV0z1b/AMkT5NhH9+UfzOm3amu03KZAnLyXFWTawu3eYA
jwaUpO6M05jg81Q2tTBW/+FT4okZ8gq+sHsdFhe4rRQK9YcTKP7hilBMkPwZdz4E
zXPsNbmeV6gi3t4HBKSVURNmiZI9AWkcPwZuJIHFbHzdW+mCKW9F0B8UJOEb/dF0
JB+i/Vhe4pPACjoVEzBNLUnuGaolfXgQ7TW7B9wrNzT7Ivejg0RVkeh/8TYkpOA2
IwLq5m+5G8+w9+il536pzJTmjDtURKvcLw4KoRDNVysEiAVyMILbkoaASl9pBNtI
sfJInStSCuh8xuY2Mwd1syvMovSlJGT4Qbu28qMp+mVPEmcV+07DX4E74st7Z1Dv
ibX1kDS1b2aktv0NLhhkSQ/KFh/Adl3UNQzn91JmL5/laBdRJ/hK3Re2DeVPoWAo
j2hnlneltVaIW2ecey1dmPYDuRCq1GfnSOQs0Nq+5iJwzg4jKinNO7z0V95k0Ny/
N5dXu3yUnJG4wpqizMhjhk5hE1UNp7WIkteXZDCCoaUy3/+MgmQI4Wa7WybkMcSb
YKRPpRzTMhn41qXvxFCSLqVPP+6kaKrJRsTxUYUqWjf7+lhlcwSqYOEXhp5mCeMC
NsdaSJbP5i+UFIpoy+9jrYM0y8Fd1IXPxMJk0XHW4+x4hTRa5qAs03/TAplzxu3f
+XJFQIt+Yu3zcetjqI7HSfJewRCKP5NE+PnGk9UALjqg9TYOir5FTq9GUQ8QXW8t
+sc1OwHAimRKHUFp9XcNqkEefne8WCidoYAhW5xBvuPHm4IvQuxpviJJh2iG7QG4
Ww6UK50sZZYMRpa9VGjK0cb8LehiIAukOhOckLGixBC5Hy5EOfdRnsDwNoTbpt75
cWM/PWh2AIK365aZJOE5BceLMe2VBBi4Xmx8/ZI4D/FgO5XNY9jtRlgI5Z/iLzr8
sBIkuknWDKyzWGc+lr3n9oLXsIhj+12te10BejXaWzMPI/mksydhC/IJH9BwnumP
HQNMBTh06eiQo74j02GrFCwzV7J3N9X/JdCbVJ6k187HfzWF8B15eqflb9LY4gc8
1L4yBYgT5LXJhs61Y20eFIKJSpggsMwjq8997R+77/4yGcsOGZTcYkvX+o8AxLbo
imVVbJ6x+NnvoGYzs1ZwD0miiwyVb7tkz2h2VI1JvGl9Nr/jCt4016ZUrZSpvHfx
/3pqG7oPBBMIO5yaQEMrP3hueonLUgAovwCIbe+NWkwjipV27XkQOpwx2aj1AUmR
hS5tAdLsPEj4coFPcp/54a+4DbVyAH8QFZ854AzpqH9iPLrX9tn7MOFaqfScY6ZA
/5bRcRH4Ciej51ozjf0/R/2ZKp/rldgyzPGglOe/P1uZnc4XHPqQ/md8XJ4XImpt
abXS+JGBDDOiPgejcJWE6tPHdhJITz7+h0S9vgZO8+iSW8rLrWIOwFWDtBxKJFtB
kxa/+yJHt/9Yk0BG4ntB+4frcrKRCe2C7QmVWvhLREp0XxF4iNxXbABqLDsx5LsW
XSskDZD2uMvnQRGmXCRG/1X1j8BB+Sz9VZQbuFFP10KnPCf8btIz0qEHQugMm8DR
fVXaALArp1JEagoFZlMwdTGTwmaR25mo8SVqNelpXMfrk5kqr19KnF2kV7Bballa
OHQ+NIodyVbNnqPNIH8Z75CV5VGIU3KbahvNXcGFeRnTR0ee8R6pVlyrGUpRvsnx
h4IwvMsMlU3ObY6St9SFR9gztH9LECiz5yaqybwaR7Kj4px++f8+EBLg2Z01Su2g
x+8et5gRkxCP5jtIMFZSZavqNY+EknXk29oEflx8KYj2OVs7f7BnLaGBfBpvwsFY
wh/A98rXDSmzmKPwWzKC/1KrfXS9mEbVxpj1Xu1KII16gN3tphIzCBL7SPb8n7tX
00jx4iT+2zJ3fuucwVu8COwn4k5eTE8+pGe5JXHk20EdMeAxUHe8kP9PAl0HhyV8
/JUOjTEZvyrZqIVqK7MgIRlfQoXvdeemg8PJHL8YMrOoEfQpNzPwBUhiE4Yi3XoH
SkSN440M8q8bazSsYPiBATOIMHeilFu3GX+Z0zDOacN0jnGkf8WfEmoauI6EfYqM
HEumbV4hQTCkhOVWYjSBg63KX8oUv61iYyqwMLGiv3g20IkPx981Mkrt6CIEQx0k
CeWMPFcLpOKpK5IEzll3tehZ/VqSa1j55bLSgh5J5psjA4K6UJLqJuDjoIxfIjpE
JolBsu1p1YAKGnMoxXggFKLRdNivnSSRpCUHmsd/FufX5kTppRv20us4rxipo67m
X0aox2Zrw/knsMGxs+F1HOLiDD0D4BI/UMEpJ/e9Qqw+vr0ujOIbBPxbeOSn2KXd
4tn/UcO0KSCnedR81VWMUY6JTU+/nWB1qOVBKEmVu0mfY4CSbD+oP+MWJ8XL7rtN
vLCEQMmBhAqfQePt/iTMggFgUnTHCSgO3xGdxlnoSa8ksMUVBIlFmHrNy/SYV05S
UWb74ol/5o7buRAEYSt4a5mUxkZSl9Wiv39I4VGrfr3lE+N5/eDmwexrVFkseR+V
g9mfGOeo9bq+x3Hnb6FPkXgGX7ySMMLShuhKeFD96KDYlojP62LZ4B170p0ZBomG
dIBRFbPvMJwvxrbayvzR8DGPNqNDqw0OkuuUYKi0MsVYX7zqW2kXwiXjxkzNSVoa
scY6H0oamHEztamht4JF+JUytQJlxx2gWOcnuC2M++S8r0jaPJhpSxTNp2bFfhpd
2iriBTaKgcH35UCRbcNMl/qaSmaXkxWkN+1miZsq02lUyEzm4NKLvUC1XW/UhTkN
BrXf89eOtp/favGi6kmhDj50VKve3Nzblki0mOg/XEfYahjfk03FfA4xNUGIIAey
UsYCWZ2Ya2371NScWAaiVcbOLMpz5FBS3CsUTx3rMOZS5MIHNbJSWTPxVE1D3uHF
hJJIaIFp0Enjj1LYU+Ahnnrzd7kVbPmN34Pc+1IZdeq3iPzdBW2RSQYsqepc+ss+
cBKznMP9+rQ3WeFWWnlJsi9VzOWqC0wvV3ADX8RRLalSiOXOMDUrQvwVnFKUUcOF
l6ppnorkhUoBkOC/rDdCbE2rkf9X2hydBAlMj6pHmIxMVK4GOSpkqKA3c8tjFOGp
9teV3l0aYyAJLW/ziidCMn4+MVolRQp6PO+UD8i5ghkkUCJQdxF+I0fE67P6BgMb
iNYtHNOMgqaktJwG5zqJmKAteEt+x40psPhDVYvwhbYTJBG/jxra2pmDSii+LUBc
COe08uRlqPpIJ7mJusnQIBSQ4s8wXh3aOKev2ct5RLu6j/UJeea0N5Ae15LWMHTT
7ZO+qI5Ri0JXtMa3zE4ShN98CCj/UgBLQ3LY5Nat9aH/j/8uBtTTGhnP70irHQcD
rtAUP40Cm7y5RL5NYy3h4pxK843YQxs+/d3PMOVRCG3zLH7gMZklrkJMaajURWlS
hXYEGRvTiaXlZlqHIKHQE7AFI69Q55Y0DQu1Iap397oK6FFbUfJSr/ufcMfNwCAm
IQHkbyEQ/b2QHoNKUjCw2P6SDO/JvnUQ+xsKjGbcXBadDzceL3BJ/9V5P9a1OxNq
2hccC4zIvcHz7nnAKNy/0mmqFrnwMfcYq0MGGDOPea3v0C88rJxdvUvVQX/K0Psa
9Ss/TcJMlbgk1gtI7ULYywTXJxhfAdTKJWW853qMpVU1NJly0E2aZ6C4DOQp99p/
/Dm5leJlmnidLwKrjk3Fzf4k5qbiCEI1dB2W/BAJLXTmmmMVTaawrW127z8G+bCZ
mgkzwYbcarKS0gXq4isJTuid8n/qSFq8Eu6CBwH0LzpWoiRNK/6//oW2B2eZXDn1
4DafAhqYgg39eDDH88f16mFIsnpFCqA3mypEL9Q9NtCnHCQaTbOd/1KV30LirdnG
SIoe8m27K5DlfSDjNdxEiK8PegMCi9YAtCp6Kq0EQUetEufsg7WM5cWveUKe8BBp
IiTWfqLTJv3FufkxcW9rgXzlLapg2uivhGCI2vRv3R7jqyyqQ/B+bJ2Ol/6f0WSh
GIsMc0XEpzVeX9GGDmVE/nL8rgtdEMcRU5QH30Qp2J+Z3PKqy4YGJEbF/DOnBvzz
YuwUGJQZ7/gK4mOU5pvfiqs1XUU2uxNBvBnx9NypCTNFKHiOkELZPf5wlM9gkEQX
YblcX3LqhKwP6aO+PvNgVinhYhBH0nolcmwNwUFOrjOl7QYQQsrWlfyuXUkAuvtB
EZ8Ey1sOyvs1T81DX+u1cuYRWtxYdsluk0YJplikuvnEAPch2UNA8Bc7sMHHMY5q
IcvKkgwYDf6CuejPRGD/R/CadEwoaMICes7UXaoqECNVpLw15pEgTwFD6jKHGrm7
Og45+Pxz+vLYWlY0/uJvDdaaOFcvRkqj9+EesFntf0nKsdX+xo0ljwvdrso9iSUu
Ir9Oj9YpKFM/38qjp23jZoj4RpOT6ZiH87zDsmmuVt0ywcPFcS8tLvFf+UUFVXiP
dGDAG+JeC7ESZLONruC/5t/N5oovfKd2ldSLKbzV7oUL2E1JF5H7hOCdYYWYwgWb
KAji3sg6rvW7I3RrVmnAUBsdAIM9Yw9m7NeHSHQFAMr2RaE9E1CnH4hsPpS4zK63
ZC8HrbkwKzG/Y0+z+NTnpW8hRRlZpLfjP3gBbieshw4t5RCSzpDSwkb+anNUVSCl
kQENOvddkNCLLyYJzG8yXL5+2emthQ/3pv4sPEq1kuDKh2QqkrJ9E52vI91JkWSS
RJOb7mtd2h5VPkDW5AyS5dzrAiwWccQbJYOTh5KNn3egJ4EeT40Q6t6YMjfLAvKD
F+A/iw20QCOIq0DYrtBtd1PW5Qg/vLazL7u1f6NX6PU6U3EV1192W/FOlEHzDb6T
5HSYglDUH3KZ7Dy+NnNUQDq35ejop6yDEMNy8W5TghHMnHEq9CnjLZNlfVrMTiOi
aJbfO5ScChb6tcTZk2RSLI+4+Nwty+gIbU4xlAvZBffR13ofBy3cD/e7HFmZmWb5
7K4Cy5E2XQHjYNuX4sAAepvI5N6ms601tomfQ3VzCxugnyboTzKVfRhfkPpSNmE4
N73KyRhA38aXKhbiPCL0cHFlb4629zTZaUQd91WDx1n5N4GmXF1G9ay56iBsEWID
E7Ve+RbcLA5fkTdz4Ufhjlm3XEeStrq15/G/XN3keG5/Llas4CtM3KLZc/p6yeBJ
rKcLODikTnnI6aP/+Qi25jaxRSMIJhfXcpOr5ux88TdeALt/zhR6cVrnyGvB1F88
ItlpfAaHs1H7sv9QeVWATvReqpOQ8fJo/8NbAMOXxjTQTH/i8NM1Gr/qt8hS+iDJ
aCcMinjNZpjbMF+x7N2gYUbAN/7r/rl+9ZEmDMloHyK3ITDQI0UF2yOBTFpkJ0Xt
bEmW/83W4+sFO81zf6PX/8zErLGS67Wrgvr9+xLRTCvyMovNY8fYnG8OjUC+xYQf
kXmCXzXw1/d4DakwhpADpOfkL6fLZdu3yyItFgh3dqukf/7l3BT19juTC/Jk77du
F+HaxIReGHz0xdJegsMXhqcJU61rx4uW+sjj31RIit8/L3PMcsbKTAa6gJxYElN5
D/qZWOX5j4n72hGs4BfAB7SH5WNjSMg5pTjYiGhQVBTE8slPlmfx+bgDGNMP0MK3
RK5JrrQCIjdR2f20DDNTcexNLbzUll8HfEICBsI1NQ/cMBJnFePefa/Yma1Oad3x
No3S4yFiiyJWkwbB5tcWiD8u3xup8MxIK/vgzyyn6BukoF4YPGYmMOBKj9DL+nUJ
Wo4bgQiIrghkkp5D/johJZ3YkOfbBZmdxObQMF4b++8tvGx4Eddg2/yRc+ilyiDf
8wsVyZfIHOFCz6sfdK2ao0RnRv6dX195B+j+l/Wq7VAhuj1Ok5SoU4X7jUoyyJff
hotJ7iwIB+28Q0NlcK4Q13aanYblN8gHyMbD/EWN4aaylS0EraevCYxZVPM7h57q
dyLJzLX2XsDfGnGUoctzDF+BVR/50XwukjnZRn/I6EdWS9jk85adBYRm9swIGeYA
QpWzOY5FHNAFNgHj2W57mTm5h26Eb016QjbefXSvbjf8Pkx4yP3CkenWX5e0JhiX
76JmuTt9/pOuC45PmM4RB3Za8LuhjMh/FKmBpKjsicxnb47VvZIFXIPFWMAVUI61
Q2+0tOdU0m877iZsLQkT6kvudiaJ9pL8Txdfog+lH/8qSCRjDt/vgtYz+qThenix
N+LaOBcd2YD9CaG8Ioadu1fQEx/9emyfklqJvpUR3vIDD+VPVsbt7+osP8/h40V/
Yy9BDrwiuMZPOkc25eBLYvBvyV0dPxVcPA0+h0hcfUTlFuxW7SZejkao+YukGoPA
hfF9XKcGHZn2TJhTgNk+7qoKqdTPC6OBbFA6BpEHaiRSMbw0iDFYnd3gXYhq3xEm
4hkaJkUDUGE1svBtMr1JxSYIe6Pcr+MLF2TCSSwHohtWuEn6thQM8NdnXinJDB11
X4a5FvY661YGrbYQRBB0igYzO0raYzVMVAHaBNQDKi/4ab12UFB+W3RVH1LS0etw
vGLmQR0Wfbm3ZB+V91dbnmlsDfso4imL6mJP8jG8taXN1DLtu3p/yn5EATg8tXmq
QJPok476/MZDBgNsA+mJ9zJUhyQiBf5BOB3O8gcZxwQJkvyKUnTe0e58MXm5DruL
iltjdFqtQdO4A8Rml4dgZMU/e7ooe7GusOpnLVR+W/NxuwN7N8eV25edxhJkF7FE
tdMa5vG/RiGwJV40LZiNUfddVacrAqkIgwMmjyPQg2IRJleVa6CNbkc25LtoNERi
wqZcYjCdz2p8AeVns7hkdx/vGxozPncAakt2mtbhznpujzIKJYbrPVjsYIEgiX2t
hzLwrir6unq/mQvq4R0yhJFZj9ylc2cah3bS9GkAgG4/d0L7+IqARp7/Sp+i+taS
y/DiK2cdD2U47+JIDgsRYIdAklte0yOQF6eZTJ/1GZ7zFJWVPcVfLejqprAUZUEz
LxjmP+NKVTEisbZLvqyx7iYqA/PVzd9qJrPVPnipheb22zyrN/P+istElEWpPwoK
UUqGtqkAGVg51VgVPxbyQTC7euwvsj3TxT+LORMFCw8cywxwIDVxx4UrkdkE3W22
WuLcAnx2TKzh2o36yLIlTiXLcgC59xhPPCHSG3OyKo152hinnhZnELV7W2P8crQC
YkBSkRmpgXytVSzw0tNl917qrpS6PL2rKuTAz7yrgWRWHRajQuqMSq0b1s4skjrG
PIHOCt5lzLIDmS1tEj/mx5lm1rpE9jrGTOUBDGCVwzD0TigSKIcBtojel1wW39Ja
hDWtqeP56zkwmRD36CkOMvkod68LLoQYaf08snrtumdjgB84pgAcfD3KMjjAUsjy
X3AggcZV3VDazb+dMKLd17B+FtviJjgd01EeOawiWAIFug24vqdJ9RwKzJwf8ov6
NASWdvZmfqvmPutnMvCNz7OEYGBCsC6P4lm0LW0jBMBQXugD9SKBi5u/P/D8SY7C
htAjzySsOtEzfV6gfGzVjETGEvgHB2rSSVSzuvk9NqgmLTjFNN1oOsJ71wtB/q1Y
8UNzz5uFehC3FjbNn1Ljur7UdS2JEfM/DM3BIsQ2T7G+bbaHN3F3MWqV2R7+XNdV
NBSt57Do4zxU7AYkHtcmWQwkvan3E0P5UzSfFnLJZnZfmDMNh29Aq1mOp8fSOBTa
PoDC9gyh8u0QjoMDGkxOd3Mkg773AOjAY2tLtk++55Sv95vLMdzN+xgrW7ECfW5N
S5OETzaKj38xInT0U4Airf8ut2NxFy/YHRfKPmdvQeej45hkIW5IGsfpzg6fI84B
ryr2pY4TJ+b6WudPqAWbNaDR5YMkmXhKHoYIeYKjLwmPE22qRJRELPT0oww2A5E6
ASjOFoCOe00CE470vHLMtSD0igzqo04qvrjdr+OeMxPdnmcfpTqHBJpMuZJzauB9
tqwo6xlBdRTG/dB7dw+YhvF+yEkft2V0NiCxPEHg+7S/5Kns1CSDMALDqJ+BG9Fo
Cq9z2quQMQP9KjncfkPQLCNAkFRQnewJ2uPU/P47r0THBkKEy0acEgjBVPJAXAQl
wsQFQ9dbH+5tC+rSUd36LN0B4SYRYn9nW+tawWYGjJ1XBX8qBv+LnmGDWUMCwep4
mhXMCvFm8TnGSXQ8MkA8yPCoBbIwTHJO7CuqZ/KzvzcuSQW154UA1dl3M7AU+WzC
UOVBO6uO6nECtJxeNlCmUPermxoU0uwGjTu6/p6q3jLLXyLLPOvSTEEJxi6/vo7U
emQRUY4tjwUufv+9h8UZx75gioh3AfFTj3X5VyekmyHwfSfuyY4v9iW3JTFPv8X/
IQv/H1OyWwpIptz9rIvyljYCeWznwGDiXwYWw7yhI4wQudZGNYYSvIrSi9b+gtUO
5J9WtEu0y96d8p6SiDOSf4QWGs+cQUaWLisQ9VLiKuTbaM2wWIq3GxNn52Gc6e31
w0jSK23tyZbn0xQkC1R+3GLhd2SrU1ck4G1TLtgI3Kxsn56xhhpYk+GrcmhWrUC/
Mf0Nv7gign8WTqSEqvTZz0ObRMoWU8hQaHYx3MphdNC9D1mZzxksfan5ghA01Tek
PuctL4SdYkbO2trVxfPng8M9/dNREt77C7f2oTgwIgR7gt1Hs+FFThen3YgQCaPb
etbSIvraO+0N3MqhWa3DK9VkXOnWtTnt5oH/YPYgKzzDclSIyHdAXbsQDRrdXlU/
wf6N8W+REHhdNAE/ns8wGxFUEmKylOgSY7N2kjfxexXKxrRzN0un3HjCUZTSS5a4
/N0oO9aIMuHMLByfdYCbaEABC9sfyEus3w2RPhl2BZiq0jnGzG/XR2LIC+GKZfFj
GYgjeUsVXXnWsnFvBGR/PMUNCKIdpmZv9hWq/Qy51KJF+J9J+ar1vXKKiFi8HzLd
GVsqfzIdtZRSVCte+4ddlpbG0Tyhfof7rOsZpx1rBnsvLJQr5QFrfkVvv/tlJ7LS
/zk+vqWquDiv2QrMFNzuWa2FRLpPRzWen9ORG3j8khcopEr0Ue9iPxdizVQsTYDc
ZWn0x2St8OSq5fJpyNQp9gDETj26tLZBuykvO0s1QOoZbOCJRkEP68Wsw+xnZY6K
tPMamz0ux34k2ii5BKYM1CLnxx+cGhLRDTHKO8AlFnnROfRJUrMly6qoOHzF8R7Z
Z9FQFV2SS/NMvuo66ivYjn9QwYXvkcAIdrtt2U1DXI2eO35BFf2V7c5ahxOme6zm
t1afXw9hA9I8TTYLfgQ0J7j45vOb2uLjsBICVO+e7a7Ow0Dx1e0PoFT7ty93DtBx
ra3LT8A+z5MWs3Zb7UBZ7WOuvoidXYsU4gVLmwFBqqIt8HUX1EH+ADDzEkWGv7uw
HIXSn3A90usUP/+lpNU7CZYeLtDsBVQgZjQ18BjUDOAgZahvAkUOL9I9Mv4hHxRm
wvsDEr5IHOvh1i72m8N0BZysvGgSVJ9I81pw/BFDmZ3kfe5RcXu+lJ7PJcw7LdGY
bI44dpkezw8Nk/m9WKO5j/u0lcp/HKuPFw7w74uRUb1A/xGOA2rJVgQZdHEDNsMn
LeWsWToYvu6rJSgOfQ1MTIVxTgkEsAx2KbPboEPRFVp7RTXut4BZWYLcUDhhRibX
+BZfK6GXZv56J0CDNhpVC0lqtioQFixfQYftQKdobzThTl7w6W/XU+qVNpww71s3
IuMIHRh8wb53uNPEnRlmBqFN+bhhLAgagMkoyxCKkupr74Yt4F3o54sy+2dG0x8K
WvjtvVVqHAzg2BFxAoXSfSWYV4CiD+oddS8MbX+DNTjeeSjFsSJr0WSfO/6p625t
EyC1yFkgLatpxDTfy4teqxKg6krlMzgRAnApGBVS0hgzg+XYKp7Fm0kQtklcaAz/
Q4s/MHKyFMQx5vxhGv+m7TV1rd+UNK+t27vxbQWZWpvQDzg7U9zjmud02ad3o4Ap
PYC/XJhCYtKaYLjkBjGk0SR45eP7IUI1KPj+6Mus1oi9ugiBJ6ccwABCv9G+pQvZ
/UljQ4Q3jXdKLLFyndvP3pJJYl75ag6XhP+SC+ywk4duK0d34StCtQvj5mfoHlEF
/bHbEwqLSpinLBPm86YUCW27KZeQn8P50FQkuEXbof3HmhSb/b3+W2QxYvE6jiGi
k45FqUAX0V0pqiaDNaHAbgYk9EZ0g1BiVn5UzhdOX9CVVi0kAerpmBAi+iDdB76b
8zIa/Oztl1IkBMbgqoiFlmmEKWb6GJVWWsFun/LJqtZPch8R5V9Gt3DMRU0dl/kc
Rstgvy5NyCv87Fq+0FNckODfqtUNuUshSoQZsTQbuIvuVbrIhTWsVB05aDuBQq3E
TG4bbT6x9s63+TbwEDHaDvrps53wPcaD7KJYWB8Rq8K1kumL4xENY9Q+5zav2nW4
vQdiwS6f9ECDMiVyljsM0En2TNbZGfvWHi01spMZP39e7YU2nLlLs/HZXULYgw8/
3nfKUIjy4zCwFLFKut5IP7/n8xJ2YZTvb4rGKd3J3i5IWAaXHvtzTFj99jNEHeXB
04Ij4faFyGFwaeWAfyhKAfdzU54zmw8bv7dwerXDFj4hbcXLZC83RFbyKGC9e7um
16OaoDRoOZ9CtLWSQqFkAq0zW49pYXuxD7IxPTen4mmTFZHthipgFOgTGsYLAmfP
36hUJkYA5VFbM3ksahpPqH3htSS1ueL0TR3VoP+wpDodypjVBxAE3WG/1BO4/06O
VACY2SjFzr/M6VtdvF8ZUqmNxBX93m3sGOLpQT6uanqgCveb264bCOAYD3R0IVf3
nonNFtqrRC96XuzYd0sddMo4bXbwS+bqKwBrXxudeyDXyOW5zNtCMGLhTh+s6Hfm
LDnknBL9AkPeUc0rkvzTcs7zw4cLcWKr/BzfrxVJ+XrAl4q4fFQLeHOjngtUn6j8
7cQ9F/M2GT2gzs1wnvZZFD0STfOdM4HpUj1dVH8OJ4jKEY6btv3VK0+DbWecB4X2
IljIML6Sv7mj0K6HzpP50voRWGA0omFcwZl6bfx4AqHbHBCWbHv0pIfhVCHbk01Y
TA8fuWhJwDk84FMPP9Lyt+5RPQGZjstaaRyiUeeVlLNFyH21slzB/k7HzFtbweqE
A8uqqUAG5aedHvIijfymb4cmS2iaTQu94ZuuzoGsEihft6A4Qu/XiRldML1Q6RPs
Netm465CsEHygzH7h1wv+kUvB/DQbuBWYeV77pokhyI5eg/VwnOkT00c+larH/34
PElAa7kaMLb9skhgo5ReoNoNIDZ7Cb0LkPCJAzvrB6mFh9H7LQoSYWcvPAAokp0J
FsSd54GfU2D4+lm7OlovWs11AB9pQEMAHX8PwYKSDcH743CpsaRDYIhQQDRpCFvN
CognnN3C4QQRZSAmLfKMjKNA0ofprmzz8pP0Hq0eCXD+xERhWYaQ3F+iGwbnegI+
Fe/H1zCBvPbi4fQCmfA8VSQT47yEAdjtrfpVDXabTR0284I96xYccIbO+6586ueN
tjEOzZjRHL2WAosWPkS9vCgQwpgkXAzg/zGHxYawPnMrnv5Rp4vOmHqedaRvwfUP
fdkheo302vH7UZMWIQscPR3XjCKIpEDhKBuXR8YJ48X/rrZWd5dmLOeby8T5CiTH
SFlm+DJW7ypWYtQVZ5/Fs/CMo7HWWUJzKEjyMtSoIoCx16N/F+x8mkSnuc3SaXpv
atRXauEav0lIe7WCA6fkwzhryOr4HpJ5/6y90WcUxEYdwuj0k6tgnrUqu2lCnoRR
3j1kaAQJZIgI7cS9nzG9xtIwaOJpwa+ZZxaRZOmdJ+aMS5/HJHRvUbElygPFLg5v
ui5E5sS0aOLXhtmr1QBLNqHz6tfjYb4xcgO1jKCEi8oGDrsmJYTdTT+KpzMP7qI+
ecsLH75lsUDUOnR4fDjQZYOuQsQ8Svb6qdFkFxEUowgi2Sqj1mUviBo22lqfk3Ms
iRzruikoP6APVYEU0pqOBFmz6I+1GKvsK5tMvR7inZ807XD4AWdvkb6s6pNC2EL4
Ca1RKnsbPbOHRGj4O0VtKor3vEuHc4ThMS5oJVk9a9w3cgOkJ00imo/2P/sew/De
L/oLyXfP2WoaJ3ChHgSYHfrpB5sB2RfK72bhUGlL1eMNLgme49NdV9ulkRdnchtw
j1lrYfIIkHMHBeaDxpKvuZsDXdcMQmm+SJRtnBK1Mxn+YZE8GVhhVJT7YIr+B4MI
B3tqRIbtr4WqDi6jcmkVFOhIjYLxKtdt6/Ildmyaq2LwVsOjrYgam/UbWU9bF9KB
Lh4gDBSTkGTD4DNLXdwY3MypvXuGeNWUiBnv0B2DKLYBsc/+TZcfWvyPzgR0V0jV
xmDVdYLvXM4PF+BPoixnjRpDyx24gByN/ubEbd2xOiogPmMeBshdD+u3PCb62lWZ
F3mTBHDWaNJKCK2aj17mkdnt17MoBkatiTJTE8FpOPGBUMT/fsgzD9EaRILfIl3K
bTrB3B6PiRe0mxA6CARsdO/kL32ctId8HMfASN/0ZGvg/9VMDzBxoZcSE2lb47VD
NSCcQHM7zO1W5QaivFfIaSMKnGHxgnCN7tpIPkdSxcvm1hIqYF5U6rNNpF/2IXYN
xdAUR4rc1jjQIGF8PtBwA9mXy8ADNYQOPBpa1ICCrC+GAVtjQt3QJsiPCJcmiT6n
IX3YcMjyTTWYsj5oHel25uKKQbdW46xFXNo31hap+dGLm5E2BtfZkq9jbzCaYZu0
cKmlksWM+2pM3OikGI1zMC2qO01JXk7Wwqr5RjZBEa+3u0ttMb/Y3U+tDy/1K8mn
/nADwQEXJivWRune4d2snLx0nMgCvEu26b8f1147p0fzqf+WWaZoFaR1YU5t/ZoI
NfvoA367OTrQLhDTWA079JnWwfNJ5mstoH9HYB8v4DCk/nee5WpORfkE4lM2lRvx
EegcvhMpmUN0wpLlQ5UUMXyLlNwyAgRq+HuzrXh9dmeXTLTfz5/uFkkeyLRim8i8
XHhjtTEhmPU9IqBaIGanm4vR4wjzOl8VZpbPcnwBF+QauD1jSWC6qhfw8UQMVApD
2yljjwPwCegA8K2+8XZVH6DPsmVwdokGAdkiS4cvpp0PB6p870jRjqRKDiyAi3g+
1xOcC6zXNSYL3b5WS6pw/JgCruNzdFmvJeYP2J1KKvxaCmS2b+z9MIZgGDDn010f
/kRiue8ngRYbtB/GZ9IaRDJ3KYP5AGVzWUQS7TH96dsJMLiVYc0MtJAaj4sNzEvr
0ONGQDxU3NP1/WXqDHfGxS4cNsgCgA+FcsTeFCSYcQzmjzecZYLk/+6rP2XgCGsL
`protect END_PROTECTED
