`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+aRJWE4l72QT0GCWU+oDccYgX5wp+Ip8OsumZfLltDqeKTsC+tvDcX7FFYe9Dn14
+7dttH+HI0A2rOJKI7crCrUIQFivFzTRRvyVL3qbh9qiKphE95i8iTJmQjLUmoTI
tyn5xmSsLRa4r2kJcDTYVLr6KghkNoXkCgjYSYaEBQkibCOJycl1AkV/qQTSClIa
wC2p4PbFZAQsq5xWfsp6MMfT0k22cEpzVDFbmgrqIk3D/aiF1Nhyz1xx+v/tw8g3
EAlAw34BjWIn9AYgpRqGx8JdUCXH7tuJ6C3DOQXeCOIfrg5sjVaNm+I+uxEbjxVC
+1DFuQOfCkR3Kwkbd4zFamTg0R2v+ApKzaFVWAwN2QgpuC3+q1eF6kG29UDVd/E6
kZCdpsg7tR3o7syyLcZ9FP7qWX/rhJ+9wuyL+4KzguVVOfHEnYjcafRcGaI9/OF3
lbC9UWaBbfcNYyzyQbTDPCNEMq0iY8cHZUPtbWLozJU+g5Zoa7tTCacfr3Q73WDo
vsDMSgWhm8pyIZXyjaqccZZ9dAK/N15E5AfGyzZJz6QYvStAmou9Ib/YZNtQXyaS
zj92kRsNprLbc7GHWLDutA==
`protect END_PROTECTED
